------------------------------------------------------------------------
----
---- This file has been generated the 2020/07/30 - 18:15:51.
---- This file can be used with intel tools.
---- This file is intended to target intel FPGAs.
---- DRM HDK VERSION 4.2.1.0.
---- DRM VERSION 4.2.1.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Intel Corporation", key_keyname="Intel-FPGA-Quartus-RSA-1", key_method="rsa"
`protect key_block
y7HVC8x3izdS7mjH30wjF51QvrOBSwoyvGRVC5oQAE5VlbbIx0J7LC5Z5ndVEDZ658fnS5GsM8I5
6WUR3z0bdXO9SynoieEnu/P1jwUxMYuGy7/q9vFEe5DcQrxe2Gqe3V1iXOVvd8ahwijiXVUC3iXr
3VYYOa/rfhfHmaLq2YYnbMworhpyr+nXmzcetUWSzO8W29oJ9TSvf8G47voSg2ry+N0IJoFg+LkB
MDkxv2Rs1Xf/uXGyfg1bvPTj130ZL/jqrLeBIsIstDlPx0oOur0u6XVEXlwLld6UfxrXWkBm9efd
KxXf/O8fKY5HJOmUXwSElcVaFhZODa/tu78xzQ==

`protect encoding=(enctype="base64", line_length=76, bytes=850624)
`protect data_method="aes128-cbc"
`protect data_block
5UbYYJ/Yac5TjZD0VeaW1o1RDhcNcGv2+0A9f2k3leR4wOfO0ZVghuRoPmAfCXBDfgbIpXiiuOBT
VfUdZaqUBzbCGl4PW5aZft/n14Tll1EWoFWc8cAqT5v53ByhQgAg8akrE3o9nlwyOzV5Ymkq/E/V
zhxbxV1d2A4tFhyvGDtT5YDmIZDRtWSgMddhQtVpfetHtfsNw1hpAEXomDuWDdY5MnOTaRiD5528
CeVbWwrxNeMk74EZDV6eOZshDuhs7YHfxYfE6yJ9teJv5nd06+bADnk6keBxbYIomLTWUN7yO2I/
wfuW1rmdu38nS9dfiYLwhqWc9waM11iXrRDBuaWSKyisiIDQv2ALdVEyi/zgTln2VNyZfe0HulQm
3dMKXqpmTtpi7ytPsju0WVs2q6y78MvQWkF7b+1ZS2/172hqJg8rrrw+xRPfXzp6kqZlWtBF92ST
5VMfBT44y0wUIwkyZfBh+GxhJREcUblXQYToNCvRYy9U0ADnDhBPl+3YTmXjlyr6FYRN4h6yH3yy
UGCgWOU3NnWOoy/FLqQsydWGOVlGiDz1ANi4mCZ8bdyXfbPpvT2EYwdKvR48Li+nk0BE3XOAmwhi
+cVUZLngnRLKNzzPahddSuq3Ic/14vukYW5/4/GI/y4y/Vlb4aNTiLYJd0AAW+RiDx6M2meUc/VH
VKqNaeyHdA97pIBW9AF39n4rJ+Bjv7G+eXedm8O5S6+A5MkvRmx2Hh2OZyudzMZOPYbclsTaOqq+
pHzIiuNGarWp0lCsu+k8Lm2CVBW4Ykj8KBwpDSx2XQbVfudZc1M2bSGi4ApanZGGWDoT7bN0s6oL
HR5QHpjuICZ0liesZ4K+6QnhJ8EBcSRv6pVeqlnXCTm4Dm2pz4jT6UA8Z18L2O09yE6lGQGa1WwK
8nFsLKoNC46Pm8SXycbzKGXzWtoEoCBq1r6pIjf2obbVfkrOSMbsXuOZIJla7RMjazwMjfQRLM9B
clueRz2CqQP+f4i2jEkb9GFyxs5fdlJ1NlFCz/ONe7A4Jga1cICWPBUbWYmtkfbcrxYnfU1Sh6Ng
QuAe+ScG1Ftlm6Jn2W26GWEMiKagGJ0+iJlsTxHaVgDkoTWH+YdGowNNNP/ItMCZUz9THBXgR/UA
znzzbYgonb1VqHnwOUug185QNuC0e0wL001+Fty+Of7ZGOkRgCletFKj7Z6cSR/IkS1boQqdH62W
S0DpyMR1FE/mx721RoOK0++rcdfYcnMW+fMUlsbe3uO6EJ/rmxTVv+Xnu+nZD8p0APH2E5EQsyXK
o1F2huC8d+A7alEcI4VTfuMCiPwwb0UDXt/Lumm4XrgVgMfKfrzd0UwNTwmmYXOgNySCfMobs1DC
UlGTtLjfNEa9HqTzizZjEJ5s6poqL2aLMcg+7VotueLKKkQHQAVBe+Zg0MKl2M9zsX/rtBcvKTFS
ksYBKBGDWrMAtI8oqnINAGCV8OpNgaOfpcBBc7H6dO1mCCJt2FwHFCAlE08tJa2Sfo2cLaAjnG7j
TfZ4Nn/EMZywFSaAQmh5uF0dsnP/27HQQlOk7IO+kqzXHtHRIvtIWMeWN2OFXMGu6IyRI2jMgNXh
I1eC58CD171p+/teDpoj3e4KdhskTF4O/wgPbF2SDAJuhu5L0gU8DhGtCk88jYLh05gxB2r4JMYd
P0H3A74DPSopywXRizjsjVDvq/wBbzlsKyXB9p3otTzbXtE9NOiQYbQRspOWm09FezV+FdqiyWOV
aqf4f8lxP9xobL8cS8H4IiVJkg3l0gDmyNQJyFqCEgst3UtF24bHD+0b+rUWGLlM/pkhUjDVZPqZ
bszdWNzh1970Ai4Zl2BG80db5gEw9/mAFUTEwAL4cLiw/f3bPty5B3grpsE5RQqyg1TzLzd6Hr4s
M4gxc/coImcxTBw4hsTED2dtFagOaq+dDLDhkK5fiGGEnjcgPvCyXE4Ts+Ee4IWTuBDpL2O0l0AG
FzgxQjORmR3lIM/6s+t7Q2b90iUVDfM6HhLn46EN6Jq8ZQox4JGYXGHnY58C3qRwiVChzqqINUU7
Y9RMlOvL1D4B+vkhw0pV631/s1jfozqKqqbZ1cq0CnN7j/KzJeljP4B7gipSuCG7is7IS+tIN0Gg
IgS+tlOQtpOxwiV6Ym/ADtA39Jxw+6IPwBMzOYFbRavYIsPu7ZYjmyKwVlA1/++8i1zvknxXGHt3
GjmDXNkQc3Br/f06JLsnICYvJmaU0LZVZpdK5AaZPXup4Xa29OVSRHEEbgnBNW32jTdDxyBvr/jw
SeesnIYDf1hSu5jmOMvdHOyLnpYZU7RN6SMpobAj82i5ClYa/kVK9NooK/fZ9khXhfzyOWTQuKsQ
Yrqt1RnvAaQ3diZ68pVLpvwb0szo+f58oLQ6Xp3WwskIcEKIQ1JDEWxtwSRebmyr1ov6KTyYS1JL
thYLSuP70raj+T+nm8bk6qJkwcQKwDqxZruOlnL5ndurzTbszbU2R/FmJ041tZ7svJaFI6P62pAi
cvWnlEieTfGAESXb8bLet9SlPyb7qU2aKb1XpDaHr9gx8mwcy4ks4gnMszeoIGKqUr059+UGCCLP
NLZvJS/3f5jU2lOJQha3aqxlF3dQxng6Eqpuwd8HKmG4jQd+JGsxK9Ij0e3nzaQ57Ngn3yE1Qamv
u3hl9LtYjvP2WH+Zpd1WPhXE8Mmbna/vKi9Z4iacz2yOm3zZcZrHNf4FojEd/DnZOC3bh9c4ErSS
Fafn+Fzg/muc9wmY0xAbqtLhs6w5016poReIFIQpn+ujDz0Bbutpj3gaX4g4rWVf7k8zmCVk0xtl
sJUannzcE2kUBmIe/qKKkyx0EXoSH9wGCixdUoWkEIGBap1IuRx6/Nnj+N602564ooSnpEp18qDo
Ior/UjrV/GRopv9ClUu0490cK5GWH6+0g0ejNPW2JB4abqT/Fqryq5vVmHA5BCGqz5p7ay39nFrz
W7wIV6Ha1xb9VH6pJ1h9Lht9VmJGSnuf3HTkWBSPcoOcvciCqXKpIDzDq6KU1CRJy7K8bk9UHgvI
sPAmPYEYfUTPbrtak1tMn06bdov25XF0RvVIdvAICtLC0+QNCs/schvothzrpP2WFIuMGO/kDRtE
imdSM5KL5OcmHiiDfr3O/9R/n+X9wsZxjqfYUcBJBwZeb7HKHUaIQ4tgb9/wHpOMDDmWsALoCYEp
6v5eGmefje/4WwdUc6fCIQDGp/PjUFngdlLUP0J6z36+UbBIy1BKzjwg/nUQ2LqIzylOW9wZqoxK
DTFmEHB6O0S/FDebPuTL6kwMf7e8kIMMdkh5LxtoIOx9GVbNGKbKhCRMCl6k8EbQ8AFKIiTLzDEA
00QippDDDG9YasYXk2FmUAteCG9IDNgHAS3bbzowr2CiCZWAJJMVrsY/v4boAJwROivRPIWn9l5X
arMLpRklh2TjzNBBGLKu/cGYL9XFoqt5kSLkS6EF97ink5x4fFx9Xu8VO+/Dqfoy0FSJVoW0y71z
89Dqcjhkpop8ri62GGiuWkkKh+vsJjQdggNaYrBq5Qnav4vs1z3cKhZAnEK97/1OaR6T5+BScJRE
ihVg8nTGcSwbJnXzwSraylO2NOsbCxttY2fdJR9fcjaWF9IAwF+ma+h557ERnfTrnQ1lOsLaNnlU
AKqJfqw/B4DnEQKHvwipz0YHFZZZ3pvR6USVz0EFGxLOPx5DkA6jjHsMYlaYLIXuMzlpvNdsoNZc
NfUS5oy/ft3Cu2iuW0PqWd8+XcjYuL29ga0ABdVDbQmKeVo6v8Hrm6wTeIRDzj/Mk3mDUUt8WJpL
CktDpZdL6LYlAWgVkVOD7ttKmUkMGZvavpenNKOuAAB3Y22a1IOlSarzh9TYA1oTarQb55A7Us69
xhrf4XgRs2U6umOwXA1m+kG37z+E9OuRxWy746duNQkistdm6ZH0wftyi+pqIC6slgOLS1HFvnrI
j9QIJ1Flyl12trZGvU+EiGKP+Ltd39pmXHQi2gCVi1VP4dU9Qp+CSDOkf+G3V3qZijfq+VGAbdDP
4bzDuvR0eUf4k9/hfDgebXUH3mse6bO8kNRlFlHo2iGI3rMN+HDQ+BMmJLbvXNAAxIq750MYp0bz
JSoWsbiWfYZsXqlb7/pEhoD/VOy0BGpqh3/W+7FWzt5aAwzIkG2bnEP72jAo/K8fYLcJD9drEAPv
7shKz9ule2gYxb20Gf8xIiCV9Qr1+N4/NEVr5ioPtvWQj4D48ULpwYqfI8lSpbctqZgOBnm5hSRW
VrjuhX+54k+6OUl4Y+2fCZqvweAb7z9xRJLdNwM1LCDfvO+5PPivyuOY0nzTSjF3DaXMlzk5p/N4
9p2Gx1ENlutnq1cy0xTiGsLwxePygYjUVPv0zhMfRWTD0jeKooNTjMMWBBJ5uX0OKERN+SFJscEK
zkcW+3kI4BsTHlwx5+zlPoVfZXxsL9m0BSXVuPq3wERBbz/URelcAJ75yJoFOwUxTutlBFZeqhYk
7H+gbsYygEuPwCBJ/gTdQ8HrS9Fjv1TxHvJqoWv+lwsMhCRFomBDupilpRpYhBi2eXz3KaMt6aoh
QyITU0FK3+YClZDh5VXpNeuwr0uprTjV2rLdY3YAiY/Ihx3ZL4CZ3cfRy1vADjOiEw2qbkbzl4BY
DhTdaiFG8QbERRQem2Sq3iRHrdk2OhWktaondAnqjMSJLa27DGUPGo3ypV0qPPpLon1Rvbz9SdWS
HILIotKXXj6RnnkWGUAdHvNFQelCi1exTMp5DenPDctZaC5S/hU45I2rkC1G2FyF/wfthcdWiRuG
j7j6rgffGLcMgb379qyt65GXhlKLZg3T9Sk1/qby81K4P8IpaJXM+Y+3x/A12HkgSjhYwxmdZ67e
6HmmeXe/G2fqbQKKWsxejuc0N1HTjjXqVYar1XuHcthXFkUKv5kVL5YUfYj/dZ2mBGgF4wJHTxda
4cQrVMkZzOD+4py0hRNLs/Dmwmi0DGR/wFb6G6YN4Of6KlHRWcJlGlF5jmrW/ahgpmdmrhvgf9m1
/I7R6eSDPsCY6LClCOhd6hedTuEElnqPngTirlqJi5vsODaQiyNyIRmegeElRPZFZJgM6MpmRb4e
nQ3WUb6kRB0uv8XQiPgVVwUyKFAki6EitQYO05u6PYBeIsxLNDqvu8fLpnU1wgD4PZAQ2symXgvz
ynQnGq8p/AqczJMGD+YhfMzdl9+I3fl++KqYdXCwUYKVbpWzatdFKWmyb0OhILAczywIAgz8RXTR
g6fHty9hVwUINTg7Zas79X2+NZX5aCTbbjaJ7o1Kb37/pkSl9gEL+OP/gUj/AM5WVFjRN7sgz8fD
B1rJerV47Vo35Kw+vQgqk2K9sjKDatSR/LJlnalUQnUmt9Kk+5/n2+srxnQMg9Erw9xorYc2rZZg
TyzQk/NiDfb35mgOFoTNYQasMBrIGuLiGbw5K32/ZEiHIQgXDEtEBxVoXDyuork+NE9QGaYuL6MP
MLsDJE2+PXIVKopys1xQnfcrUzt2A8m7Rq8ypmJnQKQ3jht60pjSoiuOSsLmysJGAXcoMkZpu7N4
he1OIjT1mpFlYhNKZ8RxdAKAh9QV/CdXI3FIlGetAEf5pilIKbO25eKNNgZ6Jsf3owRLURCk/Ckh
hXjWpPofD/eATcgi8iLwxzFmNXtMTrkHi15yIDwdGX+B4/g2k5El70LrCREn0tFU4vUR9rwUWv8K
J6BIzHdbb123XBlOUBvhEABgvRtxmumSuIqUO9oU6lqfC9WizC547xw5G1K/2sgDKr/HgnxkCKB1
C7KM4uqF0wJPau5e8Ap4mK+foqOy/HXtjFNtWsFPB92jrKzwVqJxThxIA5J0hPjw6CKykBlS3j5s
0+MPK3TTfyUpCJewvQ9wLUJkImwOrWR/aBU6dZEAC9QC4u2lQdnFhOkgxco0fCYXZjLMkulXLXzV
qR3vzMjoz3yjvkyOlJFfozgvdxrZUwFRtJLwRAEi4vYC1MgmsoZoJU/DBsxDLONqFk5bkctadHpp
W6gAdj5WWdlZyjCarIX0ibN0HaJsQQzQA0Zwle/eLipuLGcUVUf3auqccq2/4o3jfCd6JPkPOH5i
6imSwNMXcYyZmGXUtqCMCVhF8JEWT9R8wuUCCcOCvkLZUYOPCRM8xDw0UqUrvnlmb08zlFFoMBg4
wyVDNHBRWLfcyVT59qP8Bxtf9Lx9srrqduKzeAJRvDWRF6uHL73Qg5Zqguv5Gc3BnHWkMWGEdcq9
iobeyKtxW1PmELFP7DvpCIbNADjmAy8PooLaZo4fe/7wHlIP6X1HB9Nz2uI88PAo+OGjBxWiGFnZ
QDM8qqyIbKJjaa8d/QW1pOEgmO6mdCY5dE+jVTVvOhQxtBF9h59q5wKTOIEbeiIwTOGtTsk+5b6V
s+iIw3Fyuq6w0YcOgtUCSkqu7kmaV4xtYVqyhbNWcI0zH3QVt5XtHIhKCn7+XkDHzkeJg6HVgTn5
34yfwuflUFA8jK1bXNfHmurRUl1gdbuftHC40AfHQILH2gCtr6ekhaKx/nWkCViZMVIE9ro0tkv7
klnKvGMpINjEYmcxyU/u9GJdL5PD50+EloHHNngpXzvUD8OBY39RuXGmVfA5oQZQ/Or5O0srBqh+
HC8De/w87c6wtVjsPuCj8fgxMrh8DBCw9Bpa8I3PUFEYDo/9rVDqrpoPEsjHXczT6ndT9gbIw3ow
5J30t01RBcBNFDgxk7hS1fYAe8qYf1LOsQFShWW2pgnwLOzAs6rhyu1oc04dncW+PN84azGZ9CuG
Nh+/RXnx+VD9kWb02isS0Ge+p3RuEUO+nG0O/wMkS5sWFprR0IAV/4Dcfv0BxRCWz1ID0x3n1ukA
yI5iWw5JTZZvnj+wPKv9CnOZDTCfvWM2byZE2AZxKFOMe2x3ojdgXBqt8VzuJuxafi0l+JOjI0He
it4HEw0ZRC/V5O08Zp/+Kf7M7phyVJTODTUud/CXn0RseumxY89KM9j6O8RBmOe5pV4m/f/VeCtT
Vq634w2/k1EztO3cPcz6nbEcQe6fPiyXIP+4X7iZRr5HFQZfn3HfEIvi/WJzvwVKZk8vN0wL/sKx
Ahk/0/eVwDq/PAT01nXMhGvCx4YkV9UHLUZ/oR9/8yfNqTBhrbRaPYtHnTADsREhHGc5jLH4sT0F
V/Z601PcTa5Lsvki4waG49NCI2L3oAuDguGpRkQZhyavi4WqrKpcjRS4E/iy4ZvXcbzRUg/GsJWc
MTKHEVBdLY/mRbYbctAyRW9uX+UUg5z7Y5JMBRDS8uvtcH2JrDJxGo++qvXV3J78r/lTdClEcMa6
gXCgpAchCzPYWiHwQU5YHpa0jcsSR96jR/xwrov2WNQYeMZk8NCmtc3D+S0QwXT3PCzchvDDG9Cf
QUyk6+0QUFlvKrHrk80TFTcimBU7CsTiO6Gf62R1BtrrnHGBVFFYXTNKlSKiYzsTVhUIizUZgR5x
0bIYaBk+c/RDx1zX+0kGhPKFNFgvF4nunzLgGYy7hjN8F7gjWFY8KffQFAg0+gfgAe6TK4aSUdz2
xvcebfXk1GbTXLSD7wfY46J5kDzJpcigKHM9O6q2bBJ4SMj3Rl4pTOBTd9JUqrr6dY8HectpItGH
uvObmnPrderCdaCg2rDL5CQ9zZS4M3mMKY8ivMV1vwx2lvY5SFVXih/9frNvm2O/vpidycFrfhv/
nvcAmjsaraiEk1KSGRpBX47vBDVe7DM2RF8Nn+23JmIe2d9bIOXT+f7mlK6VxNNi5C0LqDFMTPtX
D0P+zNjvsmA/9fFSIY0QQn2K4MP+rfMtdJSBpIdKju/GBYf6Lb+XAM5yzCrNkY/txkbtxzxoiN2o
6ApsheeMRUqCptzwseyeGcLxclkoulwoIRlOKZPTYlSI1eIANGzL1sEPfj8t2sVcRe1Lram+a4w3
XtButmz9KZNTvsgyNfqRXS6/8qINEG6k2LcvffK++Vnm4tFwUPsKXyXlFbnpWmNsdjxybcEh6rYt
aCVJET+fSgbqKYdWW0nLTyI3pF2xdWYYjIR4sgdwO3QyHH1a8kpBd6vV1bYe3TUsIWJAhxJX48vw
cwVdgkpi4wMeAewQg21t+jE4K5iZYdqsq3XFcy5Wix/pODPAJWhBVMyuo0ycbQkUTFB0bjrv3IGQ
7gZCXFA1XX7RPBewb9+jeVKEsKIqTJ1BGgY6XmCbQg4gyWvnrso+EWP9Adqge1EbG+EjnX5vFC2M
+umbEJ+nDoTGJxQkcW6dljgjNpDXdP0HDTQm+LePjwzYx65shlPIVMM+GvHC6HYRFceeRjajG495
fxMFhtRl8VMfA4aRsWDvb9HcqnYLLCw/SG22t7BwgG5Ir2i/YuTTsqFk4RicaK3kNG8BgK/rhqBp
JR886xnV4AnxorVi6vbHRqHz9JKZBKbv87L9hY3VlgRE3mQhPe7zKzuL28t3ExjDjj/XYGC+rqve
aoiROLg6cLW8PnVEaPaQpIb6ycG+vgj315NB+HW4GIZIiij7YUngOdqeUBH74HgLG1OrpsamzrO1
I4v6EjErXc6Df8PwaztZjyxao4VNJaGn2R4vVB8yC0BW8POSzqI4ZQ0tH2mA/52sncN7Mx8IWP2s
67J1Vuuqd0GhER1bXEB1OzTEz2pwk3d8SoAaTUQ7jzo/dbyhOB6ZApCqE4wj0M56COBVtKnPl1QJ
yVoxqcp3U33Zteee0H4cKhafZcXf9KmQz8fEt/zcM1rYjk/3DgrGhlRpcKhZrYt/8unBS4PlN2ZT
csBIwCNnY8SZmFIfVzb2bkfcztDpDyw+7BP53w6YG7awwpmB13aE+tSoZVG90I/y17o3b5QYEO5Q
DTcvkYmZOduLhkTDxjlGZ/frNxinE8njt27O2KojUKAkuf/ezSnNZQmiRTvz87BjXBP2hfjisy23
lPwAkknaXZ3+BlZ7yYPiQZ2MtD6hTUyMUNuCpYWd0y2zRo9X+lMsdHjlWzVRTQRvT/tvg4l2h4E8
mUjANy7i0ToLSuQ1uANMKf6J0vEDq1pT9kJL15PS6dwC2mMFAMXQB+C8cTNBuP5WOAAD7fCzPqPg
EPTUz/fJ8fd1ANMf7fhu4DLw9J3ysaY/3dU3c94RurFjsRibzPnXw6g1RgoxJvnjtJmFBSVth77K
nwcVzFkyZDdDxBl7i7z0suInwViKIp5YM0uislhmy3X7qjgv+fAjecZK2zf8OCQqL1YmNAvyYtRz
7vVHxEZg3LroElDuN1WRwVSlojz7N3EaaWQCO2n8hxJpbmoYPMryNZtFuAqiDXsL4RhJkLiO5JAN
JUL4HFTJYzHrsTFvYLgXFmzqr2JQy6UByvzM27tn/QbrMadE9A467klWIuXAXxzdVnQ1u3gbMSa3
6ZGHG7V2z1qqBPyuk0Spp/dNMd9bIrG9v/FlRHJd7l/T2U4TuiO9ilGRf9LzYgFYtGrO5JsoOCcT
T/FIeu8FnUDoxI/39oxvD+pwlLRqZn3o5Z+gDgEQP/S8CaWOCQJ6j0r8kUmqhOUz2ecCcWRwEnnO
4KI0MUxO8NLqV39FPz4ojjjOZkM0guNvVfYqL2noVKPggWtJ2GwxyOjzL982Z7WpunOaRGG15UJV
JVg2/F/SHAkj7Ew+wIJp4pCDgDxHBS5dRhVvS2w2UXTgGgHM9E6CeXKhOozcwia10DnaIJJPE3yG
7KMKj9y8+zfTQfQIMjsbGhCg3PZnKnnWtgn6/NqR7Nast/ia2vzZdHRZrIGAeoYsRCf82rA5yxuL
IiAfNx1LvWmDn28xJpl19XQnWt3S91fD9cSH5VAMeydCh5yAqBZbYs1MmsGkdkSJX1rXn31lrjwt
wRVdKf+QRhKo1ihgigQcf3JiVEok2B754UW5cV+5w0sZoj9gtYDia3byGWiuWKQHGOWIOjb1Gby1
g0eyMOVPCgBhU0qWbWTqH3MV5lyynJ9l4vxsezQl4vRqUiDnvFI0o1TOUKc605K8qAQozpYxxB7r
uEJuhbWFe+QqKEx09F8fHlXxQ79dMXtXpbIBvDFXT0ATSBFYOPrBDzEWv3IXl+PyuoE9BShjXl+K
2m8ucT4KwSAsC7VzMGWyz9A9hpiuWwfaQiZUiptH1zuQrjMk5KaIPYRwSgviTph5lkpLfHoSGq9/
pBbrZQNokbojr4AeoWfK0Xo+Raii4ztX3CuT2bS1qOpa7jPBnab94Wq4bvwLTgFdUyw3fkDGwkG5
tG+82VRrZDRPpWNzPKNq66nkKcrPi3hjXAyCXl9ltLLXtk0/FVajG+2NPPM6OWtKf5QWCuDAaUrL
CL8x6i47Q27YtTQv8tABMh78HE9tlSELFv85Uhl2BcaK+p4dPws72muMP5CYYHTyB/l1+lpPz/gY
8c6Y0Qg6fEQ1uncqGOVHuqjSxXhwP+ereMFmBONSZrULo90uJlOEBSqgzDIaeRbtivYRHxa5Mw7+
vQzvE8SVW832T3GvFqJ43Iw4KigG1xS8kEHs/v7fAtWzSwosjzZUZzxGHS0NxmXud3NGiBa26Mzd
sqKVjqyYXIg9IGUVhtodNNTIB86QJ1j/H6Yw6c7hCLuaOvrYbbuOcN2IRtaLzOudZcNgZRVF/iaU
dN9r4I4MkXnyHA0T0B31jZ3aO/Q2xN4rSm9DW1SS7wOxr4IpQNM/4o54i8IkIvA7oM7cZG4Spy3X
SKOqhTqE2++wmQt8twUwgX8L/N4sGxg0M5td2sLztQFggW4m6vQCqEWyE283uVaL9Q+EomkLNyti
Nd/ss7DSwnkn0FhmpsoV4PDuCh86CcNMxuOw1kaYP9k4wmm4kZhCwdlSIksP13kF/WT/qpt/YmoB
g1x3Ympp8UDN54YNa4gg9ORyj8FBQ3JFzPTujsX6J3V2DyIQqHWIGKP5EkP23gVFABmI3CZvKn70
l6Z24rC2Fn1AlpvMtfVpLPbal94uRad09KxPdaWSOLnvVIL1ThREpmQ8cKb0kIHb97jgmdn0N4A0
1YiXtn0+blIjNNc0+hzQs6jtvOqvT0y5gtYz9iQSfR7mhJiRJjlSphjaMCN5hdi0fB2+OZvLgdGS
vJ1tjlGad4NTFmob7Pr8swi5blCTucjMEk5ocoyC+7h0oQZNUhPNtDlorvnA5OE2NWxobHPzGHMF
613U9qONe09DY9hrZ7Hwa/TTR1YzZ6dQpmaXq4wpDcFgTNxSzBYyPwyn6ZyfdQtqc63it9tRCCsv
dCPx3KlRRUXQr0Zlv34f3HVMn1uOxSUrJJxX7lUAb3bPg4/PStsbDSgmqW6Hrww7I+aIs6/R+EuZ
JqX33llyU8wkPRf2H8yPGQXcOlJ6oJ2bR5BfFzqMlfFXzxBME4VO/b/ellYR9ByfJ//9r+I+uYWj
ww2tQmy6S27EQyVhPHyetqcGQcisOn0v8vgQrk1Xnw8IMvYw802MwEthHMpz6vWnWmH7xQRfjW+u
ioiEjAF8dwFm4CCx+1Vu5yz1HCdg71ROUqtSPgbX6ng8cjE98YOfg2ZkOtiOrmsyDduedzCYvoP5
xOFAZ+oOveh87pS+QPRqwS7lbNr8ndtLw2aFBE4GjhZPtglQg0nHxk1ymCW2S2pw7bEGjtDHdBoq
NV2QjUJY9QEQRdNnTHiznw3YvHGf1d0VI1i5jxlr+hCEwIhSt2NQ/LN+MtJMPmSPaGB4IjzdHbS1
JjBMElKiTuXVP3FU9O+UjvLEOS/eLICgKjkSqVIommFQpBtZc6jUJa89wu+21jbzXdh/wW2reX+A
UFgnVj4Q6ZHlDo/0WEXYm+FTSunchKXaQkDdNOAhrt2RdDMbL/IhtbOLRCaACvHkwJQujQSRSgi+
Zb6Y8rnU/p6HkkWosaOld+lWnF87fF8pVREPfEOlwV0beO/oIHwjpzU6Se0bkhmyZsDVlIesYwdp
TNrBOVwc5t244B/doycJITlooBYBu9wjc4yYYxWyEJ/bsg2FUPcV506pHZHoE6zzBmXpR78VwWmq
Hh4SpER4YzgSMWhu6xjUOL7ZEUEDX2Y2cZhuRB+S67DHnA4VWom4QgvVJXoUOOllEZKD//7W0C6w
11Ei3gWxPf7+Y8xj2hp5T5ENre+fd79J/ZlznGjFLN/OY1lTy6eOl/uEXxaXQvNHsqNGJR7eiT1S
7ioZiHIHPQ+uSjW/m0vActCxUPy90cSBvGCcI+EXAwg83VlRh8Nn4/wMEcPCcJd7tUjB7f47geQR
JOLAzelUzXsu5DNRtrBfmkOVAVbg6dhTXSycU7C+x8XI4bJ1Q3FZdzdxnRXR0gUoM3N5OzG3UeO0
IcI3L52nGDpglyIqQCOmxjdzchQvMHVpiv1XGciRmZww8bEe0UQZVldtBTJGVAMNtgNBQYPdXIcB
EkaEdzxLCZFJ2fOBbcOeHg/yaO95u0HOzZYBQ25ksfQGu31JYZ9HmcapJRzZ/feqkgpLb3Ktkyyt
aRXwFEyZQTjkMX9/PgQo3pHV/dHY9dKdr0T5J4B4oXKAtleEVt3ewgmg4mrCH6SytIFXcw7kTNIC
/+7YXAfECdp1PpoFUir/3LUWaw8sk9AYe7iLw+dbMlh2dhULzBwYo4Uogs4SCg7b9HnTz1o2oyAK
0rJqWO/SMTpALo0QitQLIchSJy+ZYfteZGtmyD3SJeeNIcHzlszZr8k/zVm8kECUGbZ772AGjbK2
uMkD76P6EIzpCo7cDHHWeDA53U12xV5UrHz3WBcEAreNb0cyTpVrGRmjuCBpWnW6fHYuvMtrn13H
kdSb0m4JivZQDZrBeSbi7tbps51eNsksvXu8dkGpz4gKUVDZ4kpdetcYb6JS6w23AK+HMC195mpO
7By26z+1BQ1LBcODStI9VAGKalUWIPMnek58scBvPOkuRkyyfiDFW6682qx3ORjMsEPNwHqX9w5R
Z4gY4BEBPu6HeEB4aeOCao57a7w+4NfAwNSHDWY5D0QCD+IPE4ZaAdE//h2DT+Z7dSEXQOe/+6aQ
7ZN3oyGnAyl/XcVoyGjExnsSzl7JK4HVMbuMGuH7G2FUAO7gf7WP5L2E4k4hAa4DElMt3pc7m4c0
Rwx/+BZZMSqTVueG/IV7K86gfsE/vEuCedukYNMpAXhWzdONQ+oz2FhUzVOSHwMOKFJag2skFWa0
XRNpSk2LXet082obHgufrd4+C3v4/k3q8NIQ2E4EcDalkbsoDVRPgaIbvCUzs3wX3yMaxPA2QTmj
bXMulWhhcXHASdtsQUrkS9odTOaPdF4BLuPEO+uUsmfab7scyjcO/n29kbqFFw5eN5fwsXRRgQy5
kGt1/+qKQOb8gFVlTJ9q2MoS/cQfSk89N9Yc3/rwasotKaquAZ9+8bGASq1FyvQ8CbOEv7aIcQRu
0VN0vF4dXA8+Dr3kar8B1y/IVU6VGNEpkTPhMAKQh5wVKvWzdSlsHWcWFaTj6IZ2pBMq3FrLSOF1
ZIxWw+vNS5VpuARsSH2mFFYJ5YqXCImz1FVi/RYs7u0jbK/McHgXbNO8B+AGC/Tq9mc1WzuWINFK
SiGL9fdDeSothJfngFCTl3nUQNNVPePMNJL2R7ZZGx3JKD6dXFu6A/VAJ5z4Sjo6y7eePvwiZi+L
d6JRA3SrnVfDJnw/ysPkixBXibdqpUKh+gAMizYbjtdGxVmfSWKY8hqHOfS5fTCKCkRaemrxN2tN
XYXesPq2BzaFRfX1HHlNPzpTb9wl4y0iJeK28lptkSEIIsjHgKnZFpid2TAJQxWQ79KnUjN0NSmC
sCQ/frYR96V4NP0LpvFCSpz9Yjb8rUcqoeDN7C2Mx0keIEaLcrZEGaqg9px++/99Fdjkv/6WCzgB
anCpy3lcJ+MBrWoJqec5XO0gog1tk/rpMatQe+rH+9i2GKMFkwQqEqaYDYGb+o7mZx58hl+e28dE
hENfZObtCeck63wOJBMBWFx59Ip4rAIM8dL5eClyVtgiYP99XZWfBSW3R+jEmPODGdfJ4Phhxgnn
FzOPV1+gKyQss08kQUxTVZsvp1XDxfQfYVfhCdt+s3V/kcgfq3KOoqzIBnWWOE6DGtB7aEqv7hOK
XDiMIaaGqDH674S+vSV9/9gPKBO0Z1WO/rsqwlnIuAUtj7+PZOM1441/qPOURf3muBy3EdseV8Vx
1oOLZDrywwSxUVlf8R0XaBoIukJDZ6REoWw4W6EFyxhNkW7KHjywUNIUFA349FG65y9bTzwXOFWf
l2N5AG0uyxfIngqDhpkJ448UC5XhxZTklhscwnoYMLI1BamSFcJ9fIUfS2EAsYzc7o8dzKsiCc0z
FfjOMy+ks2oSwcL3us7DLQZ8HWkr0X88O5UHZ1WbooE5Rq5spfgldMjaCBgNCNyyIFvWVSuEgRim
fPzzEZAUwq5VyWFm5641b2jxYGiioAYATaqBu+Eoy71AUY+5Mstq75Eha6a6vecVtCSJDtZmpyoe
2juOisy7fo7C+mYUVvl4R7CNmQOzCEYpyqk1vEWn6BOA4tSzDstVxsZk4LUuZ7vKJsvERcObeL8+
zHSDl52C0RYo1Gzzexe+3rQkqd3pymmhKqOBXV1WAiQSS3E4qtsuzt3i2rycmyx774KWEBagnFl9
j7VQqeOcEZKNCVsSoyIQAc3FY2jFcVDuzQzT8/4trCx8+rhdBJo0OBkjaODkCvIoowAKCrPoT6zr
GaU0UETlMxTrT8S23xKqCyYuErRq5MTZIAiiwkdZ2tBUdwIgW5AelSWqeWTQ070Dvjoz7kCka7S9
ZNSHLRppQLMJ9M+lFUPCFBr3IdCIIBhsCDCpu7TXRMegtYa5SFoJSFHh2M3p615XdtjzjVEanfqu
J2t33qfJA86Qazc/XaKIDX8bouxHxY5x8l3Ouc5JnlONoZCtjcV5uNWRV5vnhjjjuYmfVqXP2xH1
bt7uQdxOH+J2hyzWmJTU39KwqbfsFFjiFobgQT0+U8tyb4qbF88CpzsBUFufSLAR+T6DNFByp4r+
YuAQq/6Gu7+4I+oVs51EAw7cH9Lo2w3jg2B9eyY0+IE5aT+Smjh6Tvqm8hhZctCulMiMgKh5tkZG
wrNba73DNZioI415KVe7YShO54s0zO0UOIrOHgDsD07rT+H68HeWbhggRz96EWx66hXt/Uua1+a5
aTlT7ZETYmIpiMS8w3yprjuyKzoRid1uIQ76AAQN7W1JNLq98Og40/CSFEbcuBOISqbnvexib6gX
YhySnjS4hHqwUiJHjx5CPRJ9TyySrZmEuhO/mDxw3pcAEuxK742aV5WY2XlHCMcPpFfVjOsPCWWG
6DPx05o9UxdpV6jt72rMiBbk7gjbXrLZ9ZhtnPnchM+/EwLl6FY9zHlYSyAdnc7wOyzFhoLaxiSU
K/tZdi7Yr/JIekxQ4g+vT2BOW/zFY//NRWxTNVxOmKY44mMTiW7oseXSywCcgmGn+BbusPR32b8c
r23f0K4giwhdQHLfAMnH+No7tjQJbu74sDh/19XCafEF8ekv2TX0l+38oa6kBFlyDW+AYET9GAPm
sql6eC077qeGcB019k8fjWB3KQ6YKjfltX7Q6+Kbss50bxlTW0+6XqKhFYUw91C25mwLpP3hEFrO
Cs5hFwXzomlQ/bQusoW9qmjlHcOq/YIw03FsVwmlYFPDuglgRmjf0VeqYfUe8zci0T97kXv3hBew
K9nt0wBCIRAU7pnNl8rbUtULFNdneXLphI/PuSrs/fXTVr4ALWrQyC+kdZ29SFJKFZDVQiSdnEUj
oJEEMgLzYd2m3NWXV6uh9ya3D0ZgR/WUw/uuHjLI8xiiyl0NnrKUgkZmDaWS5WNUcJVZsCSX5viD
YrpLlgtDCNKtW0FU76+WrjYAvFqL8elWp+5g7JLUfaYEz1CLwkdDpHqHqaWaz3dTE72uigNeCALv
jDWFZtmlpvyUTirAbqNtTbUCgGGWBpGDbIpjR1ouqDubJJ8SQcKix7a3Ag7zv40sjcv2w0C04tx8
GUQSecgSYkEmT+Idj5+G2rryEPgjJuSpNPBc3/SfrEEisiQCK/BVcPCb/XMk+gdL20ZUuB0lMTqb
3gb5no4oAWOUwRg5DAvi5bv7dkMAQUqRk0ArJc2LFSx8FSFVkJIKbkLEYAVGEUVGicCIIF7TPWD4
/LyZZ0vR+0OKharhlhbD7CQ9I0aaugGDVAZUWUI9cnaFNlixsa/sIpb2BXJY18/3DjZtQUQBlKZj
6nuPE9AJOL+e5z66sbdgskAxtH4aC5csKiJ+4hUAl8B0IAoq7H/IjoWvG9wpwTVHeI1BtC85AM2I
Vc525B4e1nRn03LC9EhrV7d498U8mhWIAh/LLPN0dMJGSugbGXc/eahYh1HoYVl/2wp8fktextzh
Dpz7BIPM41jGBxPr6qOB/C3bmTt7W3zSWSxHn+8m7dJ6Lx4i8WxhDx19lZEJpDoC4MDkrwbTmy9s
w0RUHjTHsdSTsLrU70CCV8ggQJ0F7I/N64E9ZAOeP3Ej96xepeOOk7uCNW8hP/SUxaYg3gm7bCFk
4MxcHiYp30Q+cgw8JBGB3ihepkqHUFJPCRnAat2ppTHVq+iLFCAp2jCaUCJ9gLZZiusX5Yq0erGu
dLNY4DHtw3RMu1SkCF+cSe0FvoMrc2XSAyLInCFWNILhRyzP5bk14VpmuHCTbueW1xQHdw+C3rOD
ZxPM9opa/SZN1z4HklS/UBQs9z3DPiD08GT8hoKR7Csa+NqMsYiTh1Z0CnLTNQcirsn0AsA4Mjb3
Gq13CKb6N7HFCOM/hxIn8G48p/Z73SJlfiHLhUSlglVT0eHXKXaYXBJXqJ1v9dTPbs81vNVDyOc7
ep6Im9b891hsGeTGNVaiYpXHHQZprVhRlUECbnx11kndBlMwJSYB1S1ptqwXAUhGVhVB4P6BgpAM
QCXWZ/vhxIVXcLuXb7fXxI6swelN8fySMYW1r2H/bEbRz0SDqNwFhQdP6iMNHp8Llnnh8o3ge5CY
0kkuOPdNcMQCiUM0FGd+3kgYA3jU1P27Ukckg98b3K0eyR++WGwSHkz0msrLh0IWxQ8/EmClTP0S
ZTmOty0kBMwfu9UhfCP/jFhDWMOWTWUJp6YNH0/xTTJVwy8d9lPygsUfS4GSJLcZVu8HM2R7o1vc
ssdtQkXHlCkvhXaGzK/izrSJkRZVEcYyZYdf5wyelGogc5BZf8EIF62sTcgmiLY+Dzz3484YVelf
XiZhgx4MY/As2RCGs8k3p2HmYWMUKXEDf+SKBQrZkfl6UZQWBPudrOW7CwGI2IOTTFmpxSVX/XI4
kbiiQRffNCgfSxcolSjXgM4dJYa1b4nTT2+epBosx4q1zX3MopMi0p+iToCXzhumcQYjJZUdQ+F4
YDCNtjcj4dQiFQMLjYjSlvjT2mw11/1ucYSA3yGQfrhnqS/inHGVhqOsM3lq0+JB/OvKBQ5cgfOq
H4cIASzag+crL7YjoY0RBzlbFWJSEcxScrgJDubJ55QMJDkrtIh+lIFWBFkYvzcSLx+d1wTS+eLe
iY711QMWll/BAenDH7Y7MK7SLOCKkWnRManCQoLlAxOztncsIcqpKXUxlSRkJUbQsAKOnMgA1JtA
rZ5LvSz7+uNSgYSE9b1ns2ktJ1Yz4n9MacUeGnuiVViO7KGvtTAp8dlP63ToSrdoszTtU8UL358V
v7WUIw6zDzn7ABYvAqA7GZsO3jL4BOPciaA0X8Ab2ACZhMK6KHfZGKDJM8LqGcwUph2uGVxeSXlo
CtBkdbO13W1FYWIYNrCH+62sNVI8kFoF4AezghzLRtdcYNnpML2jpuY93lfnGHjymJUhtkuMhW+S
I8p3mAlWq0GNXzhBHDD1uUdf8Zt8YkjOcZS2ALbKMONWKaSm8y6mUGH9fYFnN9FdQLh+Fq+R7bPd
VrZW4akyhjFN70rctkVKRqI39dO0l3R6UP9jwX/PDlSYV5dZ0dBcITw7LKp1qAC/NSFh6tdmNXjT
Ey9Tyl1KuJecWa43RCwBHsHrEOdpa+lBoMZc4vgrOIdonVlrD4rP0MYhXM9Gg/RF9B+BmiGZwPOf
dpgISpE0hKK0MMOgsftio0gLDc1nBmAt2/z3mq+bJRGdzCKjxJREKHMUMMsjpQcVGuVmdbq9+24x
rZNWgNtTsus1O0TPs6nRMyVhtWwXMGcCji557NQ3P+RSAOC6PP/6W0CDaISceiBMsI6uFqrfwxC4
3S6PWl3C2aDDLVnEJ36XMdqvV/DfsiVBPuueS5zOOAHUIQaLE6L1OfSn6cVMZ5fnE97Hwn77EeOV
ydKd7HjkYU0UhZnq8MBkQPoXlfpn44X4MHQb0lpThJ3ccAM0gUoX8XNtuH8kfrE9XGzh/GtitTXp
aWNt6a9vbx8ixN8ShTpKk2jSfYBxMg9u8DtNb4eWdcOYtJuxAFcgBRzYzqbokzyk2UPQFwkM69JT
q939SGtYTzOzbhQmckMUsvyqwwNnyySZSG5momz+v0hC/YK656I/zdxkNTNEM6XFuxxsGMpEcWkX
5qb8io3nyVugnCyb1CUImCPIgXOz1uEN3vq9s3I3mbrv0NDTAkk0C3bhxZLVg3UPhyhDMtCF/cgz
mXP2yelHXrE/vYncE27nOFKJvp18WOGDvl5cXsENe3GAfdztickhN3141Z0huHIml6oflMrajZV2
PS3jUoSkOnSq73xx96wLrEWZUUZYCTw3IGvCve0rqOCS0ZZWBGOXZ9zk555HxVDhdMnNpaP2rDZr
2KvLcXx54ewg/OqZ5xWED9OOflvR9vsprjDrz/HgXqMfe/4GVw2Dk8zYuP/kxkHuSm/XWwy8XLlO
z8vThTnNQdQmjXFP3aWdBJCu4Ep6O7zEeBgVKn/m9klm0dROiJaucEU2W5w/XCzfzleIaIXvVMLb
Rw2aCgu27tTMH9lo7ODD3VJ0N7BzBwRMSdGdsKWojKFhc5ph2HWh26DS/CexNhU2VE07DoRWpPjq
znAzFLLxNFd5lkgM+yedzN8MXu7xbPjhH/l+/B63Iqcsnu/ZRIX+XloVFVAUIAj99B+R7d1YedRG
fJft83F9wMAhAVGYXAt4ThGn3BoesJYJ0vNTnxKgc8iOAeflZrj/CnzCsvs3aPHkEik89QEy0ZfE
8/8FhgX+7bGiHC7SdKQBRpNoB8qENU4Y95y4/+2se8DRuMnQKzy9Ci3PswDz6ylGv3kVP6GGq2Cw
ynvpmWD0rcE4Wq+eBSU4xR22Zk1AAYD1Ce6jYE5qe3pwbVU8YLCud+xQ0hTA3sy9SiLcO51EGUgt
FXbjNYBCMQ+YYBcVsXh8M6erNZOc6NmDoa/U+5Ror9AohhOMDiEyWJHNB7G87BsjnEMdnxQU94c1
jHTS+K6jjFIx7JvJ0xQncbyNn9/b5e1BmKEwsIShsa0yCVh7IZGHntZSjkr+YgC1qdlxF7cyigBs
f4Mq6wPVJIjX4FffkT+KSDgbn1OXUuAQL/5LxBWpxkqF+sDlqkJNtNbxuCKHawLd+85BVpXgoWue
NS4EWYs1F68U9YmkNVEoHa0fWcfcmCL7LR6avz1cg6D1o99Uq8r/RsVrfa02R556Ji4fV0sC6+2+
lY4sL3nne1XVh+voNy8WgGnIRf5odrfNDcSA+DpU83t1/yKYbZaHFG3KUS8MXMtXNHCgnmscTI+g
WIS/dlIEcKR2h3dOzIMybszXMOFuiJN3OU5k3wDwwVp7EOSSn2WK1lLeEJzQ7gvrgRIH1B3ul4qk
kIPMXAkCsLvC3NLfTtg07iw7Fnus5ux96hCfU2KbHdhis+xiN17UP/lCUlQW/jcWOehN0c0CPe+w
nXbPGXK8hVYK87OxYrE3/O4QfiwSpJ0xkhNkq/Xm0PkYxJKRZiQbZoqPiYZgGxoiCtqySG+ft7iE
4sjBfjb0Y0XIzCDc759iGJ7vI+dLGiaoe99OzY5kiAnuSEAhifwdblDz74eRtoa/ejcr/q4kJqLj
nhSUdhMg4c08mmhoYUtq5WUvsueoghgTAgdPSZdeTdkA2MpDFfUHAWZffOnXFYL1XlZUH/fEdolU
Ob7SQQT44NyAQ0fU0Eh8gK6s3Q8L2HlVcD+yPqm3UDaNThBZ5egzbAePXg/Zky5SwIdOSvHUljH/
kpmQyC/HBN7gEuJMNJohx1XYfo7JB0+KTSpaKX7zMecTEZJpjdynktPssYRVdmuka9XY8/slFIjI
BopewTWM9LpJoFv4xTehizX/123IiiXlPoL/5k80P7H+HppqunwcJk2kDVd4R8n9lAoBVfkEoL3Y
kLiNFULDxUPKpHFH8lfL1iTC3NBxkv7zb08sL9gR5OvuL6SiQKUHsWCvS6GSx8h9Z5R568Dwz0Nh
lXDkoITybTQo4S9Jm1R1UK0nLSMlCcHCLRW8Q/iVoqgn4jSm3QpOqeohF1lN8oM65OP/36X7q5gD
WVs8yo8S/FJN3RHYjucHbSMc2wU/eISaD202+ZoOoe4rDj/8AA4HpmaZbx7abUI8nB8K3B8TpBvi
pvKRzy9saPzcTkyT8VOfOYAqasRpv7wsV9R1g4JpE1Fzy13ixWITChZnqVm/IVx1HPEtuHLPPH3W
QkfLUZZsXyMhUCqgS3lA7qq3ihebTdeSkIyOawJmgDSLhjl8bbsq705kxU1fmXyAOEJ0FOMzTqrT
A/is1HT6ZQMp5Ri7/5kEM6sNWbbPjkV9u/dbRFtMO1QISijL+gdwsqTd9aPOsmEo8Wq30uKa81/c
0riPOLd7UaOJptDPgn28DJ8hp1e+KubmVANJ3um8cgCa9+RyUWCpLibsp+KyfF3j6BOoLChpzqI9
WO1v+nv1iBek11gT9uzzQGyMNUZ0OKGc7JxCYXSp0HfRRc3jugCozIGST0f9/hN7Pyk7ciCxur7L
2T/UTzAya7rq/Gauni5NJmE7NzCFUw9+YKs+y+AzBX9kKQz0AhF4UCBW8711T15rzl2EIZTeX9FP
Pk67wzQHFJcGpEdp4DMZ80l7DIigwRAjZkjQjHJXBEmCKPt3qZ8rKvCLeQBrMIkfv5Uu/juTynHC
bf+d1LdLrmKc12U1EQw5cYalPOkfznf1j5wmhTMVc94hPSVbyM+sLPKrsP85NtatXogEuuu90OxJ
9KMvxKECAeIyQZR8PCB+pm1T1SRKP6IRosfVnt5eKroRnZ13F8CEjR1blVxEPVFaNEdAZ2rSbOde
vK1xtR+65vle43oVfBu1Oxo63S34HY10Z83iMjDr5hdW1bSQjxeJhiJj6JCDoJqO/65x/GTiXUVi
pI1ujJieUHwsX4TbCTRfbT8GE1BOO0ctIcus3DuMP8z30f8V3jinQlSRzs91bESIBJVkU5oM2rvv
L7zHS7QYmANdqnKglGGdaoojQcddaBEd1ALKcmBtby42rBwWku6zCRQoiOCilEv4Xh0qC/n7gYCt
6gP4oThgOCzH/3weI8cLzQtbiSn6UPxsJjTslyenq/nESyDWu3z5gp4C7gSQzT62eFUKOCIoU2IB
cI8uFvwhjg9QssG/4IaQQeuNE5sQr9sUomSAV5iz8aCj4OL3rCdPx+lclgYlMDtJkdX75K0maYRm
/9+Ilpw+014D4Z7trdjDyoYBJGR1Zarm+3RkS/kdM2JybwLdtfFxSAHCg/39VoJUmo2FvLm1obk2
i59h7+Vqm8wamKN1cf3OLa67Dl7l5lDJpDacEcHPHcYyWWV8kR0IVnphrTmLacdNWxmPA2TYdmf7
3WAlhHUqL7KQRoj4dCM6Akg89vg/j3QyESIEp5ygLioWT+YRSOuAIGB0/3JS+sjv2MiQ9pnvGztl
Hit/W2kpuA6vYoZjzLnfBt1zLXPIQRYga8JOVWEmOnYKh8Nsj+SCCdllC3MkabsBamRKTRCITQjI
dnht5rkqd0ygWc6JY5VhQvxDjCnzN3Zx+vIcGTzTqBhPDQYNYBNoEz+Lx8gYm+wM5x63wLQhXOWC
QjJ3cRBxVDzNpVR9un78cXYZiiKyYi01bEmctVDKFG+eFe+/YdlBQvJOXSRysG2Xo7jdYfrWUifY
PRkGfeWbjoNx7cMA8tMvLPxIh8Du/+7okRBKjKLcsMFKvIs0Z4uZIF8t5Gxkx68QLoZMoyNgm+e8
u0QJgcgn7ST/XrAeOE3hJ7VwyQIuc0Hh8Q25F8DL4BoESl+HdTPeLpNpLeB/o8Vl0BAlvh1w8Nyg
P9TzS4WVWy5ayGtnB/1NC75bmJU94ur7ORGyPnuG7C5JvtTxbbYdnMW1fx/gdYfDwz5hQC2vfNn5
fjB08bBDkR6rSNukxpcGarlQe17FXzakuLdOHrQGhcwE4gKTddKKab9DFBbsXWyXFZf96Oo48odQ
DxRTJiiZkvK5V8mjomK0EmoljzzE5PuXtjRnvl5HbBxFk6OtHNjBHLOrhyqAAkMjzWlVLNdj5aTP
ZY/dqjEROsRND5Tb6AbtqDkpPTG1glqnhfesSLmxSq+1x5F8GOCTbbP2g1J3AVHmNxIEXTGMkQQ2
Vk34F/t9jbCxC91inlp6mt0PIL7vGtVLepRtmdW6yRHhHe9mhEog02HBmEm8tDis8MoIiBqv51I5
yQZvQuafPMdasCNYD4EaSmEKECK/bsFTLJN/tehYV3PwKDTfrpO6jZZdvxONoC4S1IicEOw4vo5A
UA9wUasG2OLv9PJgziAtcKKXjeeV1vcJsAjklHJWyojutLF7TMH7yeQoSlhhzeeGqH/ozgZ6PjPE
pIAB+Uo+Fr9KXqhzwnQ9DexhJZg3RTraivP3WrTQtgrePelAHvzGWU20He4Ems4vAPJdAm/oG8+E
o4VCi7tNjAAkiksrC6P7CviwArvAzWI18mbK6EPLyaRKOO/dZGMffIxvlgPeySTs/1gXIMuALHnS
TxJHI8XWAf+aQ9+Q+lWCNTA8RIgsEPA+VzSxJQvnzJ0a7JMIKh+er6JfoQslT4aS/u+pdE6JRHco
lvDYyF78Eghinw4hrrmL9uPI6ZBu8DpGjd60POq4gawDor/QVIrA5f2swyTcsSZVubs+jyQqwGwh
iLtBythWeEc8Gq+BJ60w8tg+vdbuY53cINQNNe2ETxHVyPwvJAwLRdXRtCNIseUTPLCIEiD3tXrP
VqZTjKwmvtzs9m7l6HnBA6cWOD/H9NcOPr6kEQvbqeGNVKm3Or51g+lQkoYzTUN+sBqSTtsEvA9d
vqdF2kGY/VwkcTRIanOg42MnIra0lT8qBoyHlZ5DsHjhuYF6FvBE0wIjQbf825tRJrO76ndQrwvG
StGzXN9dtfNMzVSVJMAUxsv0NmYosNQ3OCyh35L1Ldys+WGKHj8N81EiGL4aOsMFJgFlhn+Rx5q1
GR8VeBQbDpxfxk1ySdnHrZj89kymtXci4xpJxzwhbPTFwgg53zA6dOneR9w4EhMcAAe6EhRl7scf
An/0M0oQy2RurFSI9f1Cbd5wc9xP/J00FWM2AkcpyPH0sgKiJV7yUVCRQSTunGjWMICN3sHJG9Hl
MXOslA5qshUFFiafSBwFmR+gt0ludwHzuURMjs77yt5rqo4gpMAfd51mXLhHmFg7xxLPYbF260rl
Axib+6u/X4RAVRKGA7+xTWUQA105qWS2J2aEx7RfV4WIlUOENHrGcyM+Ttr4hlCSNkJ11ItgZ5Gm
pvdaKLQ7UwmmZSU8mWxdsIAvQ4707rpoAA8HJxX6UDwCxEzrJaaN605ODs9ey5lrwPocKuGXWQgS
/XiO/3Ek6z3bmFtU51EZDzYoyET3vQ62//qOG6I6y7IXipgnknTqUqDau1b6vXBlADNc9EHhKVoT
HRdsY5GeeX3FYr4j8qytdWLPKDMfeg+ho6lppgqdFfOlqJtcGhGK/5V+tCdM/oVlxUmpd7mJp3Ln
/xEhes4zmENPSlUPNbqdAxNIgL+95H91pPkqanDCvwGzSrm5FW8YovFzhQr6uH0FrafqLPKkRLYS
AkGg0fr/DtUINAYDTtW2H8qm0UYLxA9qWrAeRpUPt+PybAEfl9qu33m8QcNxvfObsSGnwNyM1ihs
5VJXrVKLgcQAXx+ITSHH5R0A1AtVw8EAPCeycM55bEApNq3s0bFgdPacRTZ7zt4e3IebSL7yeUqx
ugUKPlwva5zLBqcpBY9hL8Co0KXyVeB5OkTgbxEd3K2Uo+g89zGjw2nPDOr9jO+APorMiCcdEj/l
j+gPmbODuoEesieVM0metTpXB7v8mE7QAeqFFceozAIedfs540PteImkPYTp9ASpmk3Op3nXLypP
fnJhl6MVyZLwH3H3WpmSc32X8Gp/Eivrtf0A7xWyAr6JJULJTcQEbF3qkUMvSYiBHlvXoW1VDWln
5K9qSONVEp2ZguBTq3XJ4uas9yvHfBBis8OoHW6RGsDFbo8dllrNA1vmXX4gkw6ugzGvw/IyvNx7
IMXk0hDighW1uE6fxNyO8YL0hR+KzOq/ZJ2MZahsBaztLHpeV0pcf1UuPPYctItnYRpLvD54maGh
OGjKQCCl09TrB9XwjOY3czRDs4nfZVaBLAxyriXIupKxXdVPbYXy5zVUhxFYcpFfjvAl8kAw45Ze
ZreXKySR0JdyTy3oBmQhfnl42Kyrblgx+FwsbSbJVHTTJM7PPWLkWCSUy/IUZFW/Av36cs62t3W2
WEqZG8sbmk+TMfwFcgVCnK7w+ybNfM+m5Pfuags2Tn0azkFTLAVbpGuNvab5j12mNUSAKzUOrjY3
/m6291CqIaHGeiODkGLIByI0r4P1M2pp/xdYz7l3cwveiK4kOhBuB5pvoeq+tKyLb8TiUDc9ZyKX
l4iO/FouQ0lqwkyp3tdNOGJCAh6QhiNLtr98eWrUKmMgPllb1WZhg51XV4Y8Ha8Y2N4Tc5xtCnWF
MesNsmLwWWTGcUXYAZm1C9fRYVdJfn43/2uVf4MMgqX5Jqlsw3c3Fw8QC/E6L4v/ZYM/MIzZHbKk
xbm1A5jZC15xkfIi9l5lb7GjIJNvKH0L65AoAJshKoMeQ5zrYn4xhCSgstOvCKMexemZ+bE8jOKf
Stg/0n7KGxjfPT92tZcBW0U2KGBUhG10xMNKfp56Ffk5PiV2YZIW7MpEHMh46uvU7dbjWjYRnr0/
yMifDTiU+1GBDWxQ2rx2xc78n0CnlYfPA6svnANIRIpBvkp+YkzFl+tA0jlq+rK62vNQh3KJ0GLn
wToWOeMvPMdh9F1YHgIsuWPPmesOexQJOksyECSXrhYMwmoNjaHD/29H/ejOoWYCoLLVhAKLw7uY
1764DfJhYnf7AaaWtbi13Q0jPndJ163qr2FATcBpjWECq4rxXtbHEq66SCeCIKM1aFcTsyvf/FOp
Z+2YXDaP1vp4F51ciFGK8/G3iYlE1u89ZYgGLrQfBk3dzjGQx2y0fH71lZ5mHXQWl3msCcmkrLYI
LRITvmbnoIsmcdC8DFkIZmGQNSw05vqdKfk9SRXJb01ZliRvelXbztURB1xs5iAt6Teh2WtkCpmY
QNutZb5luI656PlyMRhW34m6nlwcNIx0K07A4vG9e49wcv9QM40pWQvtKwWD0f5ycPK1vspi9ynp
6eaqZLlN+N598rjGEa2PHpuCAILIGf0p+HXfAALWm51Ex7CQwBouc2eCQzh0UgMfAebnOrVuLCQJ
vMNGCO4lhVz2Vl49qyqFRijtLzQ/0/Vrx1/EQN13fQ4weTKC28JtDVEDkFiQ3O4jGrGZlAj5piTM
hhkrGur6I9lOCbOfBVtZ98C7Cfe8w8aLDExl3eUrL8jWPEZmGAZY0IAXX+iwQUZOYvBoRJkJwUA0
h+KYI9bks/y1tlCxbX7JlA7ISKN90spdSL9UYtxH0tBKqB+vTM0oz/7/kVNn+AcOE4yQlJo0/RYz
y/zhsDFj+Me6Qw91zEZ1QkrJrf3Hz4xR1S9VNCMKtKwPhWe4F0ViQTkBs3aWUL8O/plvRFZGIk+1
CPKtgHs8GQw6niXzXDVTIaSnlcpM1sYwI5Wr9sKRwUte6z/8ocfdfB1YC31iaxkMh0jSKDpz+HNS
KudaT+TemHQrHMudxJXN3CB3OY2yCEQ+nWYA7+4592Mfb9qAcl3aJtI3p039f50MTykbCkxjmJVu
UTFgyFclex61kAuYCXlS1Y5AxbIUu4ZmjDEUIrLUT+N+MsAspIo/qXmKQfJnE8XioP4wdBCvSNae
E+cK/6T2qMn2/tzcEoFCi74p1AIID1eaStX2+BjgnS2hecalFNUDeDLnXFLtjpsoSMkZY4Vml8tS
FtoVyWOjSLmxiPNAg/TD0t6Ehbhp0XK6mx8kY6LNrsbRlsXxUTGSKdlSIDcrPCt3FBkYYzN3yDIq
5ZMAXi7r3BH4tNt5/W3kPlSfhig/IAWco7RnpT6si6DsheeaeQypWIpDyArRrGYVxGjvyxvewBWt
Hi/9AcEbpqaDl2C2D62evZn6OWy674h3mbxPHIX6y3l1QdIwB7AT3s8d7nSpR1h9RVGwG4+FHR1h
FY7skfb+o47KGGiQVKedC/JOU9ClgLoE66IpXAPyfJaM4X2I2UqgH7pwomVytRwsNANypgTcgeSx
1t756NTpr2kX1qRcjxh57tf//BcM657gVGjbOLCDLPAdPUon4FPyjlmtxbiqCSF5NV7jRL3hPIIz
btuUXONexyhgpPWCDatTr2TVEXlCAb4dNF9QM2GlmUijnJc+0LSvwIL1vR+cFB4Rrb6J4auTpvk2
KK+84YiZzIzJnyPMyERSPKS0QJJNWTt1+EMLd8giv+Vt4iJpVCUe/REZKpeCFiLI04StvOAuaEHV
o8kMRshtirEZtpRxoxcsqGgn1/U6zu440ps53967qOcI/ma1qZ0vfnx8ZFFkE3GFHe+nncjuiSWa
d2RzF5Q3myKaAh2dMKpgbTtFfWeW/b/6Nj6Tz6eSXl84K01wIICtyxHDuBmn04l8DlD5BMZWbJvU
MOcYds83u8/WtX3XLEk3i6/mO/JHUlXv3o/9TAN+u5+3EFSR9K5OLHLyrkII3C1ClBDyRFWIKvNz
T1nlNwnBfHyFC8Wa9vl86xKvhJlL5IivOtbZ5vZlUcZeu/4xslQ3YI/pdKvQc9mvAEaHG0CHNr8a
P/eX/8HYhGz9uETmF+npRKJo+8vnVl1hiK1F3M11h/mQoWTVDmxDZa48WsDJQkPyoaWWcRwamBKI
4H6gplLJh1AhuSNncaoS4DY4eP1JOOWxKbwE2q/HFqY2rzunN+PSlvQ9ACR13NjVl7YL1dS2mB7S
TOchoMKKlh0YHg49wy6AT/z0gXRMt/Jzjy6eRdRsI7GHH7sKeE0Zz5mFADLnDYlji2bbTTKcZHXK
jZhkjibdaMvL/43UhMyk9PYnUForUs/poOCGPrAK7WkjbDQ7ALyCVNGItBvR4OC4nNzwa1LQsER0
DXSrOl1GBJbgg2R+4MFObiAWnz4+e1NjUGoebD1i7SWuVLUBKqv4W8wqhsuaX6NP8buZYWdUB233
NlhnuuaaL2BV/sevnT2n1LRIvOAYPn0K3v8wK4gWsjc3k+YEdCWlGI0hbWSc1FSJKAJWYwbwpo8I
qSZUBa2O+A/UlrKKa3MTOpCuYHzhTTCHy5oIARmb1bLpQJzrcZLHsJsrBovYvdDqHJZs6pACWEyR
JsvnKDeJ8nyoWVOR9Wqa19Wc3i5JNZLlPIi3hxh9zWy+uqtZqSDwWZtt4SFbC7hD1rBtB1GBi3yQ
8rm1wLLlkMOCtnETQtBwI32vCC85njeisQHLxid3+b73RWP3T3UVUf4Mocj83FH1+arB9BUXQoxH
vK/Uer5OsATWjUveqYffFZWwC3AjUbaLfC7nX9+T1rIchS/DHC6CAZfBXE48q6RYmd4NYU4MRaD+
bXpcuod3mYErpzfEeHxkzZMnTcALYkAdOXROoKwOcA4EIXAXJPVUuYvtCWoiO1YdcItQChpupi1I
PdyP9l8VZFfKD42siTwzNg6UPkxVBw6LLIqf24cMVf2g9HKNfCN/ADnhFMzng9+gjhWG5uah+nrg
c77r1CZHfH/xP4GKQvdUxHAFlB3LCIrUcIM8B5x793Edce5U2Il3sfvwuPgPY1oFNuluPzSaCk32
+WEK0gECC5YsCX5UBV58izFZlb8oOl2BbU+jbq683Zc1anQx6eQRDPqhCSLnxc33q5h/x+l7ePMI
XQNY8jzJ6pFQCqFJLQqagBKa0GGq0+DuAVfjoReDuJWouDnFsqvaUC2tZEfJ0ObLRdOCbLUcX/5Y
d+N5nBZD5MtZXOZXsuuHRx/6cgcqvASr8ax4zw6UIOM5nY2vsKtKGR9POKoYFXaf6Y7gNp+8Lw9U
+dBgmRXK37w+zjBvCfTEF8bDZZDsYMToNBW34dLcFMWziyQNebvyRqTxvq3skLH+haZgrih59VtT
6Zqd5jrRsb55Lg7dKGisuMhtoMUZOOL33ABkNnguqmS/MGUNXwi8JxQSarK6vraojTX6hpYlkn4F
lMMto5+y4afk8YNyNvApFZLnfVR24LIFGbA1Xjee/tckklVka5UPFvtF5drugjqR5HynRLrzVGek
TxSCM6EWGG0N0S8ovRKy4VwV41GBit6YgHQQf+/c3nMNiLNvAGwPPf5Nj9J+MwfajeLB1s6JvwlY
eBxOnZ7pf8QS/VQfPBbFKBMBkyxj3X+A38WwCJu2mWWHoKSTMeK1ONa3uIA2GL53b8+z9gBazl/K
B9fnI/iMCeChlnWISyhSBInxagR3pEjLr+IWYdteGa79MYrSA1m4OWJ2Zo0y0kHyP+eoCjr4JhE2
ORj0e2Wte1uajioClPzURgI4hVvXPFZZyHAY761BxHVVyXxR2uL9c5ouYyZG2d0Xk6mnPzH4DG7v
ikXzx6kzxLMx+2PHlKrLppv1/O8LdKkcwK8kadi8idOIHdMxXPv6irsUsiMvlaIzILsZE2e3Ploz
dsRFgK7uVzCvmJjSMMXrYBBaXcFUSVbhY3nZLzFGGeab8fzFfViNDmVXeDK1wUYlhv7iKJOizlhB
M/SJCkB8bo0InEckX5HT+PIYrLeuky9Z0TU4V4qz/mmrUx2BQ7qieUJbQT5j/GMR1YIwKrEEnvnX
uoaNAkAhRI80wf1Ii9mKCkYqgJPQCKhwHiVVfp/Ba7oqRlIsi1qkjYxH/CujkifP4oN14YLrp00g
dcy7BHt5FMN94/Jl0FLbwrVKr8+dASE99wSnmOycCteZ2GTUsY0MHJKmF0n0i7usVt8sokl4Dbvf
0Uu6Ss5lQo9m/ytKW07wP44KFidmlacQe7UQTfgzKi/fuIW6JvroQGo+iyrNl25mKQXKaV4m0Etm
90CHAO+YZjHm8W5wbzHMfVTY0W/SsdIVOwA0faX+bd2qDnMMXS6cFVv4Uy/VIe4OvUayWL+oTsnY
PpWew0Rrq0fH33Cg4fYcCHrFhK+jwk37k0GW1/IoaOifCMtKZ9hUc/pG/W+Upd66T7NIgqnrsRQo
EsN4gX2xeo+IAIIa10XTNPCLNVy+go9soiR1mXwf3LaawmFz3ksdjbTmfHH34ALrd0YgjXMjH5pN
zdsdle3DL4H+oNMLgDMYwvUT5c0vRWJZhQrjNdZwXnJQhDInVYgqLDJ1ZVYqOwgA4xJhJYv2Q8Zs
SKMkFU0LJYHAFwrt9/eROyHoErPwObXd/N3oUIWU7WVTM+ZS5/34Urm99Nt575kvyailt9eWyyF0
h1nTdEeW83V5EMN1zsN6PIdwPOs7igPELh8/+z5doeItWhDVnFNTllTrq8/sxwUW+D/o7qnW0EaH
b1eCAIo2LOKo1qgGhJCmwu7KdziAn9MdEYxxIkDboHMdnEObnMoKRQGuQe4cP6sHGCsqiZKJNiTS
wOVox/RqG2/LRnv9s6ArkzVwaKIzupPu7R+c6WdJmu3rZlftzw+eFXt/46HSC3GvMowEu+TNufGq
GfCzIq2D2hMMOClgGXj0yRIvKzqInLGZ+uwUU57VmpD3DrRFL2TY4pkRv+c1sAgIL1TPDpRk5xEE
YeLeTLXeEvOC7mRbRkZuNF77F47RFUjxGxKjkzEC4RefHUFO+vL5kyH+dkxt4UL6te/GzFGhhdCd
+X+khH6BclgTsr/5Hlr7ikW3wazEUSlRDadG49kd5SpomaUCzGC1dWEXafeNIIRTpd7vo7A48IJT
u8pQjqIk74A9T9NnifMJ9PT0GXBiRolKMwip394LVS/1ixrieD1cKz5Q68XJWMRyl1oPNRIYI3G4
HFi3Em86IiQR+pGeYOrjjA7vgdqOghTWoTnLtgr7fa3qZNkIdIQCg1cVabfwaw4NwF8afviXLY0h
3NZLePFfLF48KNJUZoBnFN+WrfEE7UFdgGhhHuaRsesh7w1tr2am+/qdY3rDQ39NJhqwIia76izo
oA0huawtpaUOP+Zb63BL/0wBMQwxUhV4ISLDmQvBuexEvHPhQQNfQ3wqzSfR5hLu+2/RW7/HsFZW
fqa5CaX34eeQ7mlLif4LBo3NI8nmsr+tALqq6VcdS/NwB4RRPC39cpggr8Eb9EdlTV6JfzEP1v4N
maHGX97pmS+DL8rCG93uUglFXNeGKVMLVRYTIQUAW8xy0FCeutnQFnDG4LndHFwGR/MJoPVFD3eu
XdAeBICTpbLxcqQNKriWsEngqzHh/u10klO/f3vl/EaWAeUxt+7H6pa/2lv5/0jT+gM4nXli1XSg
kcQKSrHyGmrDa7u+BJYHb+BDoSZ3/nbDIYEz78xyYf4PlyMz4OjBHMHi8ZD+kzvbkPF1HawfCfU6
KSlueOvH0vNckEI+CAiv1eMOmK0MAo53LHfTqWGxK5plpEOQ5BKZI6252Pf8kCdo2X+SP+YelWSq
h05hO50R49VUgo7/7+Lo5m6yKPSRHmfv7w9g/XIwvIgOt25xZ0vqgFagp3uRchZ2dKagToEZjlhY
c1IcNGf5Gq7iwZqzRDnwaNvvYeVO5M15zr3P5IVpeUFdlk9TlOt+PHaro1l+R9dmwSqcIeIL9FjQ
YeCiuqcqWVdfBp2Y6Uin0VCKaa85Tx3jMs9wsysU7fQTwG4tYRrM90B40n2K4Y/fkT9RSaIVlHSj
ANXAat+23lNHjsNCXKvektqUT6ItBQ1lCQKDBct98ITUY6Ee7XRitUgq7trkHasoj/72o0TyXui5
EcVqh8jvpfQ7ixA34KVPwaWaKeFmQuPkWjUYfZqSEK3U9MZMDIjdUx4SZL1JL6kCKLuv41QcvRWX
BS0L81umUeTbEBEunedZP0RrcGdd1ZqDboLXstZOyPl8KOLO0jVKvXyJnm3rptpdKFQyOtw8/QnT
JYPbIpAcfP9GlLvmYzobZtOcU9jTGoTJ/pfkJMNKTsDEXHmqokJvrJ1waQttF1BesaBudOiHOIDU
VFGuRfSbtTd2kb7AnzvlunC0e+QHNsUewQWYITKwxeGudDOwyGDorgZwmdNUtdP5JnnTxzSig8jQ
yEM7qoXLbv17krmDW1yYNf2z9MCdcnVSafGxJ9sM1XLkDZlOV8swQRUJnCanWg9IRtE7MQ+Tk0TL
K1YqjXYKuh2dS2gHH4TWb66ZU8SQWcBS7yxp2lZlaoGuJoK31G42ErfJ3IEnRFWBK9/ddO7OHQVH
hTwuwqm82ykG4DKYJ4kGF1I1KpLxk1UzMLBF49i4Q9e0F0BbMLIF5lQ5Tg2wa3vn1oSsB8KlXllA
hNWRZq+7hfR8gbHwne1RaKrpVSArtjv/Fwk6dxUwTwCt4m291tf9H5GE4u9QFy7S85E8Y6tfX1G6
LYUeNxiYBVcOUPQ2ATx+F+mGwYdPLGnwJ0nHhSetF5Y1sy1pJ23R2RFlPFjMiKomIKuAHTWpTap0
eLHefNwJcT4pDCGtdnatMEOIVRx30pFZBpGz+mGPE54ImpSHuUkFPLSZr8JJ1xwh6MFhJ3IgYY41
1O+KBjqdPQsaK69f8H0KesgtFRJLIabT8yXYwxRGdPdOAFAhI3BXPDKRf7mMcyuI9/yf9x+h7sz/
qcRyGgSKoDywuZg21+bS0tbvCxioEaq+3W++NMxNeL84a/x/kiisS+GYNAGnEUW1gZaMsVko5Z/+
hZU9qNf9p+D8pJnVBfsS9JVgEIP5SNPCqKsCgkSnFCp1C6nkZhLMTOH0CPsgWK1qMUOYjD/Yfb5d
d3xvzoca+UqNeeUN4t2qE9IfSjz7JX/u9YhnLtwjlO4OmYndC2s0NpgKnT6q+7VOITtw4EG9ZaCB
X7r/wzlvpzm47/TAcNPFIGBzpGW5whijxhLRV2zWLBpAo9Yamt3mx8eyMfpxvRmulqhiwWl6Tgst
11q9K4Jbcdh1GfUcfHa8U5N28iMfZk3ijs7DpDjTPO3ncIvHh5nJETnw5gBgRUnOiCLM0fQOhki9
pW3kEY9qYBXUPvTnNQb9w8zrvj7IOomM+VBMhtSNTvx8djo3AR12QEP+WeVFoVx6XK0oxfiShWsL
YIxOFuiPIyFS5hwo95EVhbljANTzTx7ywyLgrh2w/7/QjI9Nu2s2xiIlRN0rm0BClzXemt62OGsc
TZuSriByUjFSe9GqUhgfDhDt4Yng7ik1eOS7uVgZW00nmJY9bI5YcV04edUoJRFAFMQA/xaPrx8+
/+M6e4UOk6WNwHW4c0TCwyE7EsBa/fWoJ+UJwhbQe++tzrQUueI7hEV4xPFNMUcmNLRCWzt7VHTe
Z5+Y70zSr5EjqfpPldgeMsj3FHUUNyHIrmx6XE232XGwrD5mus64jrcJEngBKbR+b2Z2TKGTZgLj
wzVP0w1ClwhhTWjWnhsdj5e/t1SNzcpV5X2MaOT4zrWMSOgVc9hIe/pKZRmHp8AfHM1YjvVfAafa
Kr7Vz4UceoTSdUy4SYc3Gx6U4TdQ7dzuUbHjWm0MhYww6rHJLEWtHJEfKNaT/fAvN20rXTJ+DbyE
O7W0oal+Tew3TPRpdCETzE2glgKbQKnSDqQGhhoQax/+rp9u/Iy6uB3L/92HCz8C4br8XIfCMg5W
azkiMDYSGiFbzkn6cBmsUakyjVhaaiQtWwqKMHSrxlqpBtUHH9HFYfcxk+gV77aw8Z+iD9GASdPJ
QBSKYNKof/dJD32fsM1VNo8ouHMnB4BEQWpTSdM+MoFSEupen2OJcTMu1vJ/3Ij7xbg4uAVrmz5a
dHUpn93jcrWbewbIXr/j9S/uhexaZ/oJq9btFD0A57x+jDYtlCLvybWwAD8/OSdqNp7rPWElXSBP
0E+LbI2M65nNNpelzD/HiV+6jfoJtHGxo4MJZ0LlMieLlvKkL/TVOsr6RU6zY6TZDsfJSiUAfi7p
OLTUbUX9bxFgRYzfaZSTxmw1Cr57uAl7NQsTYiPCU7GXa/HzPD13vwgUN8QSzx7NOOszxfwSmzJ6
zxeRJsTM4zoNiTqtRG+/KyuSxOe/Whvi3vVMq6qYXnEM/Jq8SfnjGdJ6FLsO83qungFOcHys2JEv
YFeZP5ubK2YOkYzwueWecMjCMDRcuBR8Tfu1cANUMwfzfFrQSBNoxuHYgYLr3jN0oLQS3JMWDEkz
RifzsS00hOhTgsjEkxpqDnfaaOEOXRi88R0D/0vAXtvbLfubJmwmr4UVme1OGp1uoRp74bhXOGIM
XzRS1F+RBN0Ff+0PJNIMwaeJTReTS4z/UgGSd2cApXtvsk2J724SxLMMYZ4JKwyd3pANWK2C6F+N
shWC3Ms0O9HIhlmicVYZ9ZKB7K5sL6BdxJytg7YzJMrigGR+LZbenHVq+DwJ4rUhHkJyOnm1Ytv9
vnZ6IK+c/xanMZpRBsiqfHuKXnIQIjwLYQIayaKrptK5UvPOfGIpVLQDFTwcCBzIuyC4Sqgvy2Ed
/H73fiBdcZrEWtP1vfe74fpgu2MQdWtly07RVWQb50x9x1ToGGxjgQ/CCuzYGDduJNULiyIbFchU
yjuEFNmo3VCisDyTPn5fgJMW6bsVu8mZZ59aoCMoMhjWH6GbRXamFSJZNxIsmW9VhcCX3V2HgmH8
QskBwtHBZ4el523gI8/rlESFi/B8cLGWs4aVZuw7FoDtDSWWrVVeTo+lcL8NDfKddi3fKnqDW5bx
eKskI3KxwuJMC6A5Zy8o2Oxr8NwaHEgmPlxotBg0EkOyRM8TcxB0zLGsf+jO3myIqxYFAe05XkSg
5bf+0xPM64kef7wcp7I7gSIEdX3yzXP1ecccOTlG9t17/sKBJNpWmR2KabTIGvuxIn/DfgHmfYDJ
IcMf/tbBCaY/iW7JAIceRKuFUJwAFP+SA4dyVxJXNuTaloMklcw4nSTpneymIKISAQqXJA7hfNo3
ncAzytdRCHrTgqdqoqCUZwwY8grtyUR1Uwq8YsAjBBQp/UzA3ROELkXIIAaBJUZ7CUy0EJx6to6K
QunfePGV2rW68mK/wf3cS5/G8MUslHKDG/16edOHraZhguSY+zX45DN407W9EOTHBDuo7stbq/z6
NYCGhMy8+7NruEGs4a0ysItIyrMBm5bBZsSae2wSUfUBTeJiHeC3s3S07rVzEpV0UpZo7YmX+WOG
hQldRepNaNyA+jLJirOH8CdhvrSWpSJNDCyIpxniCVCg3eGkfJRca4IT/2ByQUTQM5kylkTdnZj7
cbnwl+FKAjVTpM7UgRFI4D0O8Y91ACERHQIkMOw9KVE+uU2/LkF1TuqYL0QvJeCIAIC0t/0y6WV9
RWhn+aE9fbLmTfGi2iX17fo7AVld9N4j3vq8y5d3criLHBt0ZLu+naqabfbCAoV9JyupvFmWl1Kf
eGrbW3vN+3PJe9zS/pMJhqtx7E6egM94P3ebN0rqdvCUEvJrayX2Xo2vVq/oMSw3CGDvm0kpNWns
9B5WakPsqmlqSF4G2XQRo3V69AFqXpa/WvttHGYG+ILEu4HMl42Gbg5zk5YOSJALxsaYq9n2gNHQ
AdTFINIM1+FL3SrI658GrRLMn8jsYq/u+ofM5jEpD2tYWsOSgiVVKKnq3e1cSbPV5B0Q0lCYx9cP
LZdxq4GrPTAteWSrwuKxO8oKKh3ImKs9JcxOgzWCHWN1W1JoLz95lqfQZAgHUVAHac4/ITEnH42J
ZjbPScDXRHVoDrZ4mNiLvtGOq4JBIi45JzWVT23Hsf4e9oBiP9g/0znfQPnWbDaioQVoPVd/3BAT
lzZYoPDzymrVPBgMlHdDi7Ln9GWHgMtFxMCzDxyF6gE3H+TzZXDeOdfDM/0xG+GSyjaxV7rU+s9K
lBWx5Kj8Jba6VQMGK4JZsDnz00o8BZm2lQs9r4ff6MtsCW7z4uCgizD6rA+v8+2+bJnLN/TShXOT
fpDdolbykOMelzOVUVN0zoL61wDJDHSOZmdhRBxxneEWL7U6lVycB+gCKTrlOKoAA+HXHig2SNYd
ZwYdpwylFt5LAymU3uPb/5UrYb3B2/YPK0yXN8jgP/n8jJ2SsKhxpi6/m29R5o2POUiyb+jSuOWh
8b//Lrku1k0ZMjbgOVV8eEeUrYyKMicY2bsYIFW4gglTQVH3DFvBEo58QxqYg21eBmaXZeWSBbwT
j4pp5tnaU0iAk2stwnpxikLUCpDlUmmhrRgckCQyvLiaJT65yfW3fH163t+Bsk0ajqReGB8EmuGC
GCz1YLENPUcZRpMs2BcOIcZPFWGlumTHxHNhyXAJ7qLNzy6CpPNJio1RU2YLRpMe0RfgNhIAZpO2
sUiDAvE9NZEk7oRtCqcwZs3tkjuddc94mfnAXvMSS61shjYZhtIi/peKuGMf2KoghlpY7Cwy+43p
XjXO/xO24vvUd+znRPkUsK4fNUVUipAmP97cs7cYlqDFMRiP4qxZvTD3z6h5qnINjKO8V2Y3dkDQ
NBqsrx0Gja1agKYsPAGxMENUFzQAwBAdtqYnx2lhhW54SCwxJKoBTdJQpr6LWZIKPzfMSVKLCcF0
epOCzITBCUIeV0QrjBg7EElQkoKMIVjcWN4p8FXTo7jwWpekCKlm9jSqlrNH42EltnTEl0h38C3d
SNISWdRcA9P1K0dHu2iLsXG9adRsIithRN8yjMC0il+HETmKvBnUEP23gG2Xh9UQrCeLxJeLGEsn
/si3sVGsjNpSC0irmW+2R4Sn2cIUR0heAnbRusI03iHCHxoXNFj9yp3rZJMqM8wbVzo9+2TrTaId
UEZdk/QoeXSlZ8O4U0Iml9J4me6m7t69/+DZVvrzNA646FzM9IwepK23RjiW7OYi1WdXOXX22M70
gAPbvDslY0qJG5pcIUN5/2jcMAR8pkSQ6T7XndCNfxgEs7jZlQfewCOPaVvLCG7w9rF4v1KTPlQP
7pX9qZDJajLQTEoGsYYI4Tv1bzdZe3WDp5NtxEkMQ3ovcSFdXigP8xsed/hSDN+FGX/seETygA7q
+HvHQYHPhAh7DrRR4PpKALPodyRLSN2TOCfsX6sZlxNYiaYVcVuTK2ZhhnZQOocGytZ03WNDEs6a
AT9LAnf2abFRnpZRRkSy3ETmUPTuxlFeZp6pfeKV+i+9whHVRpRiBrvBu8uTVG8+PlCfOdE4bUlp
YyfAUa6+9tEBPRso6+i2R9av5OhXg/kkYiluOqFX24VYM+jCQC12gd8/krkvMXEAHGhxMHGXqwi3
r08/1zNJOjwPEvXRmkoEzdcqlbgIb1oIi3REvlXuVRJubnCWwGCz2EAVqgQoXLCkUqLISpSQzbNw
Zdd//evHUdbIYVi9GEdzGCXk8YQIdVJhdbSnTsP+D5uLyR/3/0ZR1o+BOrkk2GjSjsR4Dd/GsQo5
ecKdezYkj3wXrO7BC1v/bdkYgVrhqfHIPqQPdOcnILjo76fZo9uSwZF7hemKFTyRwrjbMxoPYFZK
U3jBkYjBmY0jxnA5ZCyrp4SyMSTWbEECeDV4nvL79cIbg6m4UGezEwnoJUNUAKpC0E1DoMsXU08g
HImmVp699s62yNhRCc34OAnSsVETkTM2ISsANwJJaqk+4jmx5cldvOyqSyWxacWiBLx5QaCEe8wL
521Ty9NLmtQ1jHRNmtF/E51BR6A2OzhKfLjpSuCIK2HzV2/wgGuirP4TfQaaLCb7Z3H7azBaU9sX
NZH3umMIAT+2sXip7wlyLnb5HikIzbVcI1yOXoo9UhXNBzvZW6zdjrRgeDQym3gR+s5P5XH4Q4Wq
IytkziTMKVY52kvero96fDc2m6EPymzX6FiN4KAFy/LGrw6sR9DdD/ZwydToC1HI4TbovgeS8Tm4
5JZ01gysPV9Zs3o4D5EdGDt4Ad2CJN0gf2P+nx8dKQ6xBZ82NqScEnxXTxNviIyZS1PzehhY8uyb
bjvJ+GvaEyV0J/6bOtoC+ZZ8bkD8ySBbN4CPcnyWXUF5yyKsdBC+P6h4Lu9BJWTyPjVSVMqk+fMD
pTDdaab1Kfh5NJl9VFdiTtaEcfAkBL7qlyw1N166o0+3LQopfVdN3c8sFNAJ0OUgcGkISM+M63Li
VbeMJ08jTw1i8Gp06D4I64ZcLaoi/IrUlhjg7iT1hM9mYBR80wzeAKCdCvyA2uatYjDgIGdSpho0
g68nHVaSfoMPnZWOmD2tG33H7z5lB87YyST3EtcTsbeEMq7gugjLTyjTpQNTLzjikhZVSScYP+nk
jp1P89NMPxBMnzFSDOKvJgJE0QOeQeHSmb8SuSG9KMqTcUYHM7xekiDXYHFOyjAkrB3WP901plQt
Muy1laDAjslJ/ThJxkiCA04VJ0HY7Jg0M3KDzcSgdvkITna/zLi574dytFlU129/UCyQFUOB482m
EeHos6eggIWbN6btf6RfsnsmqeUUAPxV+G149mqad/eul7z8h61HOV+CidfnpfOGsskEN6TinKfI
kAcea2U77U/bAFG3UvYRV1EwcmniNzmQUjZUA41v0BtTw3IdfprGaW8rH2teDb3ZPpr4GqBXYQCr
aUhFm9Wzdy/2sNjOQWFjrtj5S5+Ps1pTRFWVW1gmTGPM9WFVi1Lu11jjhf7CkV+TnGBFnAq1g8W9
RLg0lFjc5mNXgfayyMXdIZ44cFLuNJFfYX8XuH7Yp7wGUjfbYMxu+oZrjMKZHJZzAJB/s045Qfx9
tFw1TkvQVgGqXrdjINIdladgdOe2NXHfMUt9+gbuJMqWx/iUYvcQJxM1MkZxLurLkbrt5NOZtTNr
k2CX8T0XvNahyRCQE4fxI0R/D6wGcTnhnxr3emQdquVauXqw6s0nyLylfV1WiNnIkZRslaq3VuUZ
VUwa3+jXpG+iKiwdtyGNczDkXs2o7asfbBLO2LLsRmPOvYU51zOv0N4FG5tz4X7WXwOjKc79nU+M
MmfWK1aNnvDgEW/BoibnCGIoH4cj74zjuF/qdmgEoFayyIp+b9KKU5hjp9WhZNxGG/fJTldO4o/Z
Pv600JSe+7tCCP4Vp/YfNP5WLGmlt/gh1LxoPoSqH3WbyZJUj1vQQHP8fwa4bbSFWH8kbS24Czt/
W8VK0AnhEzKMj1se5bHFceT85jLEgDEBUeK5FcmzT7HBmluM43DyQ3EdAZP1XI/DeppaFs5LBYrn
sQArc9zrvhwER6jTDtJeiDXLtZi2pi6+w5tPIF0PfmzMlqUGKTuol63OO/4rvzlXZVDjtmxuAhFS
tghTD4QvqPrv/dkNvonIqWMbMjMe3EWsdWwuKBiOe/Z8IwR6LAIOp/QD/D+hoRv+39FmTQqnHC3W
HQGRp93Bbx1V1D2mo/Ttx+VuCnu8yW/TfirSecqcLH4rg0fSX+s8kuD5WprHx8AZW96MozRDhKPv
rPnBSvwDxGMDxxDDXxIoo4MjiqlbylwNej488b1pOarqKrgAlO/9xJqaLNQpO2TWeUTXQKl4TSuU
NHlOWp25lhPFBBJ6BKFqXEozFQK0w7ZtTGMzk7JGE2amf8XL62TYqyL9F63VKjO6ZhksO1drNb+J
T+jqhcq1Ye83f5TS/yUKfbMS+rQQVBYplXKaAAM0SoCxyHg9DYPMC5mGfqdr42W9SsRZtwclt7j1
TfJc1cOOSwNvtxjwZqRbHPBiikbrs7AvLqZ/yeu8sfTx0dxFGc7ktvpx3Wgw15O6Wy+YjipfsGPI
0DZGJXd2in6UCuGJLbnInm/SUDJwy2wAmcpUcuPtzyrXI+ryDZOW4DDmVh2TWuPISa0bVmbRU+ua
wzaEcxU0W9sYjU/prTNkNL5/ewxW07T4BxKHVbYVcmTH7SdNxeQAdDflSZOjKqOa7Dm/rrSY0PBZ
fQaGZ8shie3rH59EPN+SnXkwcLoFIsyZfm+gPeWJliRrtlTVzYmeP6uSIq5DXhS0yYH61XT7MLZ4
Imi19sJ2aKNGNMeM+FUd5s80eoRij730Ks4/4ro6ZjLilsrFuq7UncN0tdGgeypcuJYROiopouVn
8NK7kJe//krT9H2gXLNmo2OvSw/gL9/+aS0vvz+786amYE2doioKOYOSpAiB94OJ5/qnXKP7gytC
+AYY+PhLUDO64caHi+47rfRdj4UpM4CkTr40QS4I028F9WekYJzrACGbhox5DvKdE/frsNgptn22
tASGSxeqriM+B8MmZZgE6TOkQCLkFzKUb3U3ShwGZSyy9aYJXVVrwMmW739bIbEau8g5NUSxUnJp
FZBXMVWWfIpD+EIA9IS8wWU8KJuhbO3sgGBXQTSH/APQ+fLG6YOIsSD3IdZVTMNcWWRx4KXm1Jjz
rGeZlt3y6sqlzjj1hUWsYm2byQtMYhqaL1ig18jDG7D51U49xLTYL/OWPKnje0LlGdGG/KN3c9Cl
8zPJIDfaK1O4lY1CQxdUF/OF3kbIKv7Ci0vgYnoNDB1cG5DpWVCZWrc2zwMSbOQkuwIwogrr3Y9E
f/W20ziKUWZunnPgKX8uMJcmIl6JGYbBPx3oCHAOp4q4lHzSQDfRtrNfzt6kCQM5Gz6djkiZu19e
6bf4HkL6z2GvVcHWUSxg0MntfYM/EQKzs7zHPYQ6OCP0poMETbXKUAW1VS6K6dt1mIrOEKBu7aEK
dHXP1/OvUJG1GN3ZbvQXy61SmMayysPQZnd2vlRLIC86HWtFQ4PzmP/T+BQpV+76aSn/HTtzWDYN
lj2JoaYpWnA+aPn5ukyH2qsLSLoxJVAyccNDld/Dtwa5iTV8fOD1clGL2zkvUCabrUJ3ZEx6ipuA
Xh+2ENHFwPL/qAMSQjh34ak60L2iZiNNab3XwOzZmY0i2uD2/P/au91Lb3mzdg7Mkhk6/zHpO56V
vpI6ebPxCcDnuvBTMkgcZyWihzFOD9YrWsBpyatS+Gl7ajcCRwBcc9W2hM9IpKQvSa3Je42EIhde
gr8DoM7KlXMJnhQfc4VKwG/06oXVdeLY4MFKbeCZW9dILnk41yahUN6LQJ9nrBjwHTQS1s8NtRBB
ayERR3pPQmk0yF43OlNp0sa76Qo4/njDxdgwX5dLMpOkV6DCCj08nYw6Xa2htT1TVCG8cTE1mfTI
bWuCrXo8AM1/ZEslvZjGnCXtloCzPlVsvnYXdQsIf9u0ELa3FyfwOWw7odT6YcaJAu3p4VlIRayQ
lOtt5PbLDcAeIK/BaZLatX3b6h28pVMffyX+pNIH9fTHjlSebvhQznnWNlDypVC8GrKz3F3owkvj
TlOevlCutydfevTMme2azXb1EfkaYe3+xiiE/wPG2LT0lNfVkjvqB/tJSkyFjcO6jxGO1+q84T7f
4UJQlJJEpahfkjdN14kY359ZQc+bE2TvFTINuagv+noJ52YwlqChqFB5T3qxmCNsoX61EvibdArD
eaDuSi8bS3a0sFO4PGkUzibNS/cejRtkKHjwlKZpu9UQ1QLyjM0L9lJ1JYf+BUfdZbxgi6WpZtHo
r6NxSwDt5EcXyKUNNoJQaR1GYUuwbHBwT/cOLrv5Z5msmllf6dzqgpStWvo1X27gisSZx5vaILzG
jvhv2bHhiQ7en8QdBKe6vUYCWlzLemfRGF0vx/LoNpIr9CyljFmhuDWapYgHsgM0D1XWAhihj+yq
/3d6kbNodLwKqdFEQHHCeeeLor8iWJI8Tde17zQ8cPE8n1LgL0/Ztg6aqvbE8+aUQjpTFXolQNb8
G/OK1eiLdGT7eBwcdAej1cNYZdgJE1dkRM755RXpeytm8OD399I1EIkYxksoSI9dGcUlWI/G39E3
eqLOj28+9C248SawW9lgiRl1C6Tt84gaMUZJhXTeUGSWbUA6iRx/apuzbHpLBxx1d+KZV1a0FIPX
NdsdXCZfZEB/NtX7L1da3XYeFmMzSYrC3jeJ7jvYLZOqon4CoFujMDl0H5v44+GCw+l8EI3TUf6S
JcKIXGJvxUImYlqgpjOHQQC0eWcQLgKbl66UECYcjJjfd6pYHSEjJTtmumaW1N27tISF6J44Ph2K
tMrpdcvvi3BuAYxNAAjaTcIKQM7Hwt6I3/PuzgH20WkASif56C9PoJsya2uPCfCOYmBR/E8W9cXe
ICuQOfg4vx+ZaUARxSoWxFoC1HT9a6VOdbk78QFqI42q4KLNvYmx0KLkeRexf/i3hA+3S/zBVVFK
9ROuWsx9+ZuAF3+h0qN/6kyLSmuZx36ZbDfT6rb1gh9xmeUfwphpBv/5u1P6oiBfpJ1pDREZX8zN
KyhUwWHGxK8Z1T3aOwjM4Wz76onoDQHcPSLPuddwhbQNrNqNKvs7BrWZUuYb6i12OTdXjIJBGDIN
oPwBVjLGGyZxxS/WtzOqrhEjhilFzYo3yyECidGkvby2yDamPdkRb6aK7AQhc378K/7o9tgMyBDh
ukKlxsgiVLJLHGEaYV8hp673p+Kc1yUFSIDFf12Sd9JZaodn0OHckZIgPqq405PhcEBM6UACkr7p
OGKntfwamklZXDG9mWzQuMcv5rTf9gff8dAnd6Aa+R2TsJS5P+Qyttoym7vwG73HI2MRQTo+R2ti
S62V+leUn5dCVFNhoxyhDtJmrJZpzgzjEPc9eb/pR8IpmJrenFk6DJC26ID09J7ACWfVAm0qQ7vf
RiFt9EaHKhqCIIt2ZsEmLG5SVCLnsHH84nOWPfkSrTYjBzQLZTmdtSwpgU/DRTirNXSMHsgO4O1Z
z3/VRrsFqoVHKDDXYuf2IFJgLLWfofCmJE/aLnDlROBGu6iGnlBuqbznTAww8l6dTuLgpUR6REz+
eAGwT9lb5l+wXQdA+BgjQXJn/NItJ39jv2R4i1hmLDWz+iolzjQLZWgtOlw9/8wdK0orv0ldt4pB
cMC7aWsfwJGO+a6fM5denCCHm6fSEr/oG9A4uJpq8+kozOxcE4jl3sBvc7jbIrVlHkEXRvQwZjXP
DgkhJxptDckxaTidJJWl1p76RA13DSWed8IDaFam8zftxPDfJ2N4QUCN2Eh8EmdjVoCTONk2fTLl
QBrCMPXzcFGHAg/ykYPVp3sXDd0DTGklA+bkFdKzdiLrb2DU68DyL9eE/prmbPmu0oxT2NnVstEF
eYl5y8cH1d9LAQYrDCGIEiwRwxyF6CUIXmUJRNeM1zqr5bB8J1ZIO/4XYPMjzykDOxXyZ6n1913K
YJQk0jlKJSm92FODuR7MjVwwmbge286dDmBFx2RE6XD4A8pPxrs08ezMApXKaljdpOdtFZaLPQPt
Dj9/9857Xcg3ZozyefXNO2z2GFhgWmjn8tqftjLeOY73NxADm3c6LrLfATM5HlGWbi6z0tfq9Obi
DMkq+8RiC3lTEdQByah79HT2ZtewlE+DJqPrOa7NVGvQ0esvuOJFqm0Wk9xwPPwRlr3NcC2p07Ag
5Pu9n+Hs16GgahbLVyRJyvu3fh0T1S9s+6Fz3z7QGu7OAXAQrQOHFvyXL4h3fplr8QMq9bXeTdFr
IUKfMu944xaz2XZdLfXHCaT6NEugXlDy2Z59kTo6PwS2/QdJrVoJE/9mKyl2PMZw6KQSvljQII+n
vFY8XuqgcJvvPG9ydD0Q7I0oUkZ7Ax7lF/Tfgour+QKwjlZcFv/PcCE6oWpWYqSRMtPvelCUPVi6
FHVxP9f0TmhwRy2ZGGRrfVrYomnK7rfJ/InRgNFeVtOnWmNzNMfuGHUJnLvYKZtKrDvQyY/OW1sp
vEoc+F0QyfjPNNtSxYeXND7iHb4sVFT0Qk4G0u4NUASCOrgjYPXW69dXtRgbtUkSY+juK2UBIxGJ
SpbBi/ENfiJjZe5ginA1kF/Jn8WkPXj5hucUOoWZWcv4lBE5u+UGStt0VHWgepFeyuOvjtiEcz9+
RI7RUJDfrxaqDNWb/zkBlNBPW07lmImsnodmQF+DVEWOv4p6Kl7Fpyr+4LDbAqUs3tdI82uNeg10
du2yb21y1bza1D4KwCqfpOmTUeJ+FGwFfHHHpn6OeQClPpnqGziBd+NGFlNia/dHVBwnezyrXcvK
4Pml+MczMGdAqVbW86RZ0PXroCZTyNMoVWECj6YhUlve+0o4/TqYfnHHdNUlBNOgE1Pv2HsIDwGY
d1gVDFvW7drnbxF++h2tjXJBNMa22fdRSxRGCBcQJl64qYuNeeAjbGEW7NT8uH8zuiTkd7As83Po
0WjUwykCHmX5bmzWgvo0bQhdDESIMdQ+MXaF2fPn3m2wyJNbl4Ibv8RzbJLhv+RsphgUk1dDLnG5
ZeXpgwebNMnN0u+QQE/bTKVP2wnCtBJK47NG+CXHk1pRX3Qdca7M2G7iyPB/MIqKfayBKi8PonNe
7QQqmPdhauOQFdQ41fRpO5b6l8r21A2H1DDpFjVeUbbNS8ASLpRV7M/OLU7Y//POYYg5Y0+tC7o7
2+1+8bmdTgUrs9CTVw4ZU1hOb3ilpXtNnRYGXOPN94qHauXEw6olmlSG3YpHsN3rely2oVN6GkVx
1PX33pueOpLGV3YIFhMu+MOzSPcHEiISaOmWr31pM88cV9eBzRYTk8xJRVyJcc0cYHwC5sQ1WXXR
DBelGHXGcV07Dvg54479jipcYvk0uC/iOTwFtkHMMsqsYiQ8D26oGIdNXb5iwOrdZNH1jlsbMuH3
xw1xIyEF6Hv8idUwWmUA/CHEFzZlhl341CDo+kagp2/ma1Ati1yu08+RngB08O8tsZJGqbpwGTlR
p+7PRSSag9SL7e5vZu4eYzcq/LPS8i6bE1ux6tBTVqNoAE3RZ9cc6YoDE0bKTrhoYsy08WWWLpaA
F3wd51mMy0bdhX9AT9DGfLD5FWBw8VuIVnxkPaIVB/FhusTMl580ZRrnh83kEZRoLPPEn77eClrA
R9e/P2QfdrAdErrrDCV1ixToqqtSbkYvInjO3SNSw38esnV/9AGAWSVhLDu0ZCUKdhCRnO4oXSDC
WtFKmZqRmFY7zKlLLUOPLFyPDXQ9ghH/4nvgW9xTnYhXcA+2IXKqxma4L9twJh0vx+awQm9y2BJG
A+kqNanESZGCDezhRf7DBWEkAm2p7fivhBrUr5o0OWrhlFJ5nw52LNVV15r1GV4PFr5PVBrPn8eH
Eqi/ZlDQAXLrrq/hyomj/0CpNcfdKByx5aF9Li7NKI8n8cmMGpSM+DS7MgsZtIXB6JAqhnFTtu2u
8MV/usXsyt29S5TouEZ18vFgAzcSXV+QbH4yyX2OnzfsM39ixjjeb5k3oaClV07O4Wu4Elba+8i7
ycJexqC3Pfp0sZRWYMTHjOBVqCCrvdO9MRNzxx8MPnOtQ0cEBXG2AuseFogUsxoNeb6tfrmdv3Kr
LsHeLmhNnmo7Ix1VlpJykDbIyVPPi/SkbCN4qlkyDdcpFLUBsiip7zYNIiITWH2gFdh5zMhLUvuF
MHyTeD08yUi8Nm5aVwnISNfDp7n/1ImYXrmj9FX1i0VnAi/n9zs7AkU3T/2W6tyOoLcS7zCnI0vV
iRVAHnrBQqsQ4e/e/z4iL7c6aFKUeY8ARcN6d4vjHm8OWCrLr1L5ce7TWDAiCiJGBodZulu/dvv6
MoEBmylHmGhKmJdJ96yc4rDTSR/7+/3lJKg2656wmeiq3vg/UEJ29Yf/cYYS1vi4v3DCd+WElf1e
Dkhg2GULuNoPSI7rCHtFPVTsilp+zgBo6HRWtVJahSaBmW17KuMa7yWRFld17yG2VGb752Q2hffW
bDsTyGFNx3IJGT+GVMBNIP905r9kUWiMyiCsFisoENIgfHKp2x/vdnDIArlsHulnsCj56FjmfCew
RVSV0Rk9WQ2hQbArf4NvdLXfgyHjGnX9XasG6UkmGXrHtIvqNCNnK2I3iheorpugPWZoNjl3yiyO
VohB9vhUXTBlKJPHp3EVK0XOAmgbugy2/Sm8Y/OqqIuu4M5iGGjT7BslpDBTmYC9/iBgbRTYkJno
/3Cz+d3LY2ZArueD2bLLbf2357teamgW5LnSTopZPOGETi2/pi60VkRn3I0DlqB2N3TUfO6L6wV6
5eKznYYv7E2cZY9Ykj7/rCxoEJtqhuuDLjh5mVnxUS805hu4kDx3hV4dI3z6UIlkv5pP/qSGBTTN
nqB4zPqjvF1kEOS5RK/yp3S66Os9hW07zVw0bQKMk3CiK0abEMmTzLPtXiRKbM8CnjlvVXnLNid2
/kc+yoIQn58RjCEnjhbc+3gij8V1CimAKlRmTDZVoY+KoE32jxA7OF1gr5lNJlDiqT+nvj1C/SqQ
rX4wVvBApsezudJybm3MqaM3xI/LnOiXhRdhw/iAzp0qY0UnYykYAk6m3DHoUWnxzO9cpxLYflOW
l8zAFqiTNzNBnb2pCXpoyvLnkOhfKteV6iVeVmh9xZZlCKiSfnlFTa3PrQBJcQcEAzNR/q/xhWvj
fBSYTHnBF1xnT7BiOo4GsJLjPjYeTEN3V4Swxt2gkFFmn/AXTqAM3ytNidVh9FX6mxPO5MfUHnT9
XYKFerPSC0eNcOK+C6hSGj4tCd7d5tIc+uIk/EJCf/szceGVWxBikGmggYLDk7U6T5nL/ZPssVZ8
779Vqx1NyitA9YqE7WFUfofBLyxZaH99nlK1Fm46uTLoGkL9i+t+wXlkdfLWmkydQ8pSo2+X8xLV
f9QwBPgylcN2TErBdTKC1F1DksCizY0EwOxM8t3PAcALwFymbxfSOrrgCZAUYTbt19/HzcoZn7UQ
OGvnqWnFNQL1FMzn0+nG14J1ufzKCemJMHbHzXxW9bbyzKs2X8BpO2Ofop+g57o5IAiwOQVo4Uo2
efxgFHnB24ZRIBj9vLH4J5OhZ/yrmcOh7pcgj1K4VtZiv3KH9I0Egz/K0TiVLDhWB4u7QNcPxYcv
Fa5Jr/KzHW3ajjNxlymKJUz2s8M51wBBuZT33LLXO0u5tvQGyzkqEzGmfGC4edaAdJ1wmN0cxlm3
nSvGJbC0XByum+kZc1EbI/utk8hsR+MUek9Gz7YyNUKupJB4m8cDYj1RmZY+AR7kfxmdTs/r/DYH
RQqKBEoCUfzBvfLQfMT0CxAZcqWUQdCXlmEBGPB1RhXHS9DhwKbHE1QKrJsG4Oc4ewEaoO1iuLyr
UPzRWuVYuxHPdmjQp6hCA9GFqVU+8lKICKYdAVAOwHaPZzFBQYW9N+BtXDuB4cEd/ONBkI9LzX0+
bpzVbj1MsFfGrgj2aebOJvADwUIhHWK9+EtBII25kFwBzpv5BIBz0ZrdY3fbqCWkFMgCnjRHg49z
BapXT3+mZQEbWey5PcGyhSKHNSioiE9bVIifBjuase5x9tHmZJns02xDN736UrXAXpYWhA4w64tW
tqL8YSbG3HyA9/4eEhCoIMTkMgqmMHrAjJC3VNv8nc1dvI16FYX+kViRDpY5+Fde6uvBMLZGod6o
nHa/bhPwdM8yOvXDydEtasby41XzTBxGUPu822YU/+TV3+eU9pLc+ao7B1Y8AhLtsv3U3oiQYGxB
ZshUuDI0D+s6vk3bXCckBthE7Wcp1VCVbKEkrOwXl8olryzm95obdeR4FRVdLL7Ga9Z5IEaumuWE
c2JaA54OuNcUu9/VGXR0TjpOZPpvHCFQuDMd8GsPZkDthHShRRd3M3SWUx0HdtJi31w3ooX9290W
6e8Nu5GOQ+O+JqkcuQNwB1QMhn+LhuuwFn1ILFbQDw040SnQRir8j67e5pe4NWSJCEpcTPo/CFMo
kNzD52ZL5edJB68SowvJ7VZHfs2+or8M5a+GGKRhUJP7EUYjInDYHsve2fP3ClwesGqVcjn1VtUL
QmtyFIFXcUJIf0DIPLT0Ppmabj+jfAQcqJq9B5K49b6UtD9KJIA2BcbS3wLfYhKbc3TXPgpEfNDP
lE7U/hcLCSSv5HYLZcfeQtHzclpfu3fiRktiTtmFYiuxwR2GZSGgUN/FBmEr+1/Zr5E4VSUtIbfP
nocP6V8YhgLsQz6UafDNu2iGRnrjuRa6Ti+crJmh6tXKRoBgKdWIvifF/HyQ4ebfWOgfZAojI0BP
FwpdrFYctQW3rzMgYjEWQq6g5Tu8hOnxRqatvnmwJWSGlNKFTrYnb82B/4fctgJMdMuManeTSbeJ
UDhdiybDGKuMrTR8nuDi5ijEgBcbQdCfDneoUpIrsouBduQ2j5+iNSBEHgSChbqCVEffZbcFZY4r
hmjaHAbO7ELgu1c/dgB5bdDAFsyOLL7cCFt6NIuFex8iIZwwqMxxeg8BPPsG6O1sdddJBu7MMxO1
E1nbckD9kEQAgZQ1doNbLDHdE8PEFFDKIl2MG1AHhbyDjtlshwRCsxoPGVRwVOCBLIgG2zbHpj1O
Yhq3wjFu4ffgAY7X4lzP29X10NQeFW5iYkTSuJxIA+1Wi6JhnM36RKQHtlRDMoVU+cfmJ4HiEmv3
WJDjJmGnGMSCl9ktD5kvVcfOJGjYQZti7CoLY0rUsICgbiTcPS+5iVrBYsjBt4cQGvmI5e8fC8/h
aj9jUyQCl8U59jNnOacaHgeW8i/IdBV6PpMho9TiHaqbT1ys3YSzqrBEqyQkLc9xNz3Y4AbVxbcM
+6GiKd5yEDqC54RF5DpM+249xS3zOM0+vlB9L2QGPioswuo95BXNClTEWELFv13FrljfJ7Y1Dwe5
OqppVaUBHM0tgNvFRuPMMtbvcNdnpnsMICfOUAdvyYI/HViT1083nJP9D7UQbC0KeOAWvevj5eVs
w+o0FefwsrzbP+rAwBCtBGYHHJWksM8BxEpVvWALq9U07VYt2KGCcXskujxnHrP9izAqdUfLpXIs
XuA4Jsfq/u3A5nuUKfR3mpCrLGa4SdfJz/zKWKcExVjVfGufVC+UTW/qkZWPfaEN14W2QaqYCv5a
pMBjvXdAclCVcCLmOvPEcJQ9rbTIk4plktCZX5may8aqyY30AmWmcXbqj/1ABE0arnlW4OXS1D/2
fcGKb33koLMPkPPWrWNNj43Y8zaoIe1OEkCysdrW6TqrpIqxos1jjBtoOQQu8WJt37NOhbmUo4Fk
IGyhxz9PIwQRJJJNAfzOahUtLOlKRsSWEjOkPeOfAmoy/0c+oPLunUOp/AUvIo1y597/9tj3aa4Y
kczm6Wsc7OM56uv1+gw9WEdy52RGqnQp94Aipl465RIlW2Cco2i9RzJYC0VFZuCkgStfzYCZffNS
MXjCe6xb9WQUKwDcEc21HsaZwNMfH1lAs0Z/05o5SwnC9GJuYMrvMRjDXpILqJ39Grvsxl/D2pal
sOshwl/lFiuyrT/yA8oGIn/MgQcdsKhklEjjRz05PQm3Ros6auopvRfGhru5CnOfN9fwDevn/aXg
jPT33M4HjS5DxnfzzJRqYD8bjjHZ2oZQ9CnABw9TlLpRIB7AeUyBFzsRVuF2MA1rqAUW68r689kF
1s5MjF7zYpJYhHjDcADWVQ37+mTKqHHd9kpYVLidMKPxsfTOJhmgNfQkQ2mec9mxwj5gMJUcPBku
P+pbyigzZLcWzTbuO3LmbmGeure7OaFUq5AuhmCcLluzt4kuSWl4kQqf323hw1/Kg+zl0d8iA2HJ
a9vVkw5ibsUW0j7xDjxtchOF/a0T/w2tDvGOb7Rk2AAdXTcyr/6bTc4Y3gbhzuDVPDegwNss0qEG
1kaEuDOR5We6fhwTpyMqopeXBrudIqfsYsG4IQBniSVbkgkTaXpYwjPQkp7IiTdExqKWIfk6d1gW
0tZZBp9BCcWlmFxoplK71jC0S94FM+ZA96r8RsQg71ECf83SZtbdc9t+BNummFsSdEKRFo0fOPab
FvlHkufxtUvm3hUxFQ2E7pF7Au7XuVzublUZl6MKK0CPF1ngp7xy1+Ru8CtyMSoYceiMQEDbMy/j
2Fv92v82hxU1sKGCiYlAIM4hBjo6z0bnNd0CDUrEMFTk1td7tk4BmRDLIsza7KP5vXi/3Zu8mA02
7uJULon6LlCO+v3nzeO1fkZ0DAJxjVU6VfLRGScNSIgLMNTrRBdPQtpwDYPYDm/H8AKE69eNP7aM
aKtE494hH8qOd1K523i4C8Ej85lABVFgyZUHnLJmSh26sCL0yCCKpWNg5PmvIA/d7HTuR7+5otUX
SCDESlDnLEX0BWT98aXxJlMo/qOYjGLZCZVoRkTPQoerji5Q7Y7kUnL6rZiONxEqnbQYZOrSMA2m
vXVpbDSZeXoVHwJcld8XziPyTog0ScGzhEXviluPTHY1z/fmAKDosJ4MdmsvRczw6sULMsA8xuS2
nnzpxv79c5hE8B8tebLgfB7MpT7lYe1toLRn43SxVoQRUYtjItZhZpGFD2cFzPpm+2tv5WEDcZqb
W0KoULWFqhIxzpsLeffJPsSi/yYoNrYHF1P7Z7IDFW4llMvHJNXLL7cwE7FC4MVre39I0i3IZGVK
RRamsvC/75Xbbggoc3UJjojdQM100cgL1CdIi9SzypQEKJ+EEgm+J4QX8Nr6Yts6TV7Lh9WzgVze
GS/wS8TY8KUmAGYlqcd23aBZYyd02a5Os/Jcti3Xw7XrdnTvsF4jFCtPTjTeukfZoL4bWeGFjukc
tbxlfADCxYUh0SRRR8+zCIhmjzKRr+01q7H94rXlZJaDWvTO6SdkFUKy/IT76mYytzRP9kgVyfqm
tIKItnq1y+KShBr7IK3Jgjg1l7RiDaNqBS7e9SFgV4n6ejwok7GFawHartfy0j0USVytgDaqcn9V
6LhP/UDD1HKe6mwai3tICGaTJiERBuOafJ/BMXqR3FHDBnQncmdIAmHIUCrRwE3PDAIhLDL4oZH8
YAjmPHBs3lL3Ar6QbuiSFpaOOtJtXWfiwSXLpbAx9aw7StdY2sHJlSok6/s5vNzYQrvORolw5DX3
vtY/YRLWEmIfFTfjP5wElOQTUnBK9RcFlRA3tIfVxaBnJ1x4khGJBQiZY6KGpkp5Q5VKxh4JVrOF
qMq6cfDSfXBnkf2YwLuXnUsymRDS47iVY8yaR2FctpqzIjaVHnmf0cXKydTF+oqRGSHf6p0N4JOW
01Xa2Tc8E6Me/aIoBik0hLO2PoJoj1svIlbJkSRaE+VBWAaj1QDYah8rKM6+G7IjEHXBjvoio8+D
KlnjlOJPUj+XK188dd2dCnBg8ZAiDPXpYIVX0aLiCtmFNz+oFAfcyviMqwefL6h4GYBclFhrD2Xv
xrwGC7Ugi23OiSWG4dIelH8zDBXsUlC4+I6wI25rjVOcIckeHeQ2NDDA9i8SFfq5chH8+XWqwH4V
Bc+jl2khxlK3AgtiwF9IlkVbFuef32FCUgieey/qDbRoYLx35aD2Kzny0Td/cjImvKim8NV6/wAF
e1l2nmY/r+TrTv1Kh5SzGXKO1MjueBlLCXonMtzAVBUnHhmHl0zZMpnKAukyJvL6+PEeGTdoYP9p
TxyCL92nXhHgJ93UYl7GFkDIRa87vCVaQppJo0mLLrAmTNDJFjhfoQsRVeuMGz7QNaca/4y/y/1p
sEzr2ngDl8bUEUJ1wCThPD8S6+90waTu5K3VTr9w380bwY+SnZJ8o8ctC1fep9U+bIZJsIUKyrhU
kDSeOZsuNzoarSXiAkwLI6vao89cyuSOGArpE4iYkTXHhVWp2dbISSSclRB7QS6nZdtT5x65WwRy
LRUdI7mhfKUH0hT82XwX+dSOy4LT8oF2dx8myzroxToekoyxy+uNiDHxJioS56CAnr0/CEe/uJTl
0yiUfERes71veW72CKR5jNFJ45N/bTsXO9pWWREk+L5W6cs5P/JRsK7DDrIbaxj7NYYgxYajcHxu
kdwuvp3bsFy2idRyj32+ZGtTqdGKqr7eUv5jNn7X/OY45GCvQw/gFiBlggezVN0/dxAnxjFL63so
7pCohx6w4ETQ0NlcuO2K4kqVxcxTj785IwBDByMY6QDFbtnDBYJX4Y0qbSutSXCYJpTV/FIv2Cam
fkdg+BBlpYmBlbtQytXb4pxRur8jS4StKDUa+8IFyQ+LFAERGy/nq6M6ELKqAWHJB89XYyg3jKEc
gwpDe2qpD/IGEfU6rW6iecjP+dfuxaDvSUVUGKyICE/6TuaIMyh748lZMadBv0BxdvBmifXmebzy
OJfCoiCi0P7Byz6fxznopoDYVOkQLYpdyXsCyW5Dbg11qQcQzd0uP47bBEiNYmMdh+hQbMXZXnp4
Th2YNgAXj7gLTnBfOjoIqROLCuwZop8BNTXRbBQkydzhS0Aj/JOOyhE2Vo17Ay0IE8FkaA9coN9x
Wn7x/oKcXhWsWg6sK5DF9PqLpVx2ApQus8hsr01vxQ9K3zd84A2a+oCjdqatWx3MeoKvxBXGC/GD
f44H6taOW9X9H6xWONYw7cCWqciSSf6gZcACixEjmaHQw0JRmRjeDY6EUFlIOy1HRw8pRR9cpvu3
OH3+8B0/TyoNnvawhZ5Z4tqzIJesSPVu04PlHFTciTfFn85r3e+sStl0Uk2tMIjZ2JdWVXo9LMoV
ZnROoOg0OcvtIgcGWv/eD3xMCLe1MxixPzNZRKC1dkooW2/a9nbLE2w2LVT0hahL9aDv094AB1fG
k11whxMgvfWtDxup4qTScbyjW3qkYYeskdQqu07fg6mahjRFO9HPNTUHgenRPokTbkjjE7S0DHD5
4wK9Au9Isr+0V58LBnCR7mb/i09yujuZnxoIVEhDNL0XA1DgUvTjBGpfHzYOkaHapgeXyvlpLdtu
wW0u7Tc+erLjDbD6WaO//BsyescjmDSHjRC58oAbJ5ekSs04gZ5n8DqlCIXjzdHsx595hm8zJznq
1k8lhYybuHHnyLiWqcekY05Yz/PO8wKsZOPC7aDMlzwgF8FAMARRsJhmRbaWZnB6utfADLAiOWzQ
PiUC73wX9O2iFWnVqdlZBTsC3cBDYSKk4GFkNbwEegqqjPz1e7J6CsTV5snDGZ++WmDdjFSyd1Th
aM4ZaSwhWAMHrhvtpGXQc15IdWqxXCWIRwCkNjLeBRZdMe9F3ak4BWNkkOOlcSiEjxC1EvqAtItC
BOWt5wpqV3p3P4Lc9lM/OCH5QJX4gUT1SINjZ6Xm8IpoBjfhJHBYOjTRvrFhVJtT6NBEnlrqNpgK
p5u2QklcmE1VWipp0LB6Pz8zAd0Ek+CprKRpxIbmLAYaKZb9wGkcy/9sR8BVyXMHZPe74HRVv8UB
VB8FQX0emNwFpWasbk+z3gp0jtrhW59mV3Mdeeq2OQ0XPzLMffCby+3fFmd/4KU1j9ZKVsvW2qlv
RauKfozI6XfPgeHx4KwZuJl+XHIeufY05SAOBZWngz4GDZTgFf1yhZucVemRWpgX89d8HkJfAXYz
282sws7mmeiqncr/WSlvfd2vw7XrP14w1Vj1vhaga0K1SOL8sEQsuxThSDVsXfkbZderm2YJeeT4
/oBbSmQ2Jm/B9Jvggl9oyJe1M39fCHPoSs65E2OqHX5Sxi6DAerBi0Gj2Evih7jS9XyK7Z425IYF
4kg2P+PjK7PRTyNAVmAhBxY50iknKxAMgwoxP1znjZbL553UCdlkz/uEDxFWc2f+j9rrz2Pf2O6p
GMAc0tM9fjZD2qv+PAJfqG3j7n85x/2Rf6xRV64bOBdsjFL1fo9Pz39tY4U04OYT6c8mmakwR4S/
WeLGTRCmBT6A+bvEjBGuWoiigBWxUAMOHIJaeW7HJeDN4hlY4DMbkuWAuRM/Tju+ltJXitR2Yfe5
1ucjkFvKjXXYhNR0oY5zev3C8Cc08QVsovF2lW7qFqhP3x3FM5x/9TTzZhfTEU4W6MYxUP5R5iPw
uVWXDbuKLfjM0BCkLPx+4W2liOv2e/O80Aag9Ncz3PIJ20m6rmiwwtLqs0QTC6jHrSP6j7EbBwLF
EYHI3bykVD/IFWgIuN5d/wDqSwJSJrCYLrUQ6lqqEYNGPgsQqj83wmobYooPeRELB7hd9nz2I6M1
KCw1OAuavkuMvaY/w/ZbzCXzWHSyNgdbrMdaFM/HbJVFrtv1Z9odZOaDrwYL4o2fw928hsm3UpG/
jumyQUtLERzuzyGxtvjbNXxbWN18tV710Lyi8vMSjSrQ9HwD5L1XUdpBoP1mCQncnh5ulfWXk30M
B9l6VnlM7ZAsZYm7OEzU0KzLHxSJebOBD+A5Phvw4nGSEVXQ1UK6iJ9RROjcaVXi5dkHaVGnzW09
racYaN9JITZd+v7JW8V/CLkuoBpWQ3Spmy6OBqUWdOpx09IRoE6cl5fS/euB0+49qU8tT6BLUx9D
yNpKARhhe+avsis0s4k2wvdLkAPNjQG0iTnF/4JijxdCqlG2wil2yq6/fPMEb5v5Yd4iM9mgFK8B
AhLWQ3Ur49P+x/BMOVCqavTrb3JxiyG9XXNyFO4ffxhuV3r37a9IMZheOmEWwwQS8RZA3pZCMCZA
HWcrQnV4KqR9D0DUAzY9ZK9L14+km1OS11nZAA9CT84qGN5ewrVyNw//GHbNlF0rflH7H6ojDqRP
qxS/HB7JWjRjIavO1qk5HDX3uxtoDNLZyk1/Gc5gMT/6FL/Tr4nOZoLSE6uhxtCdX+3s5hKhmE9D
2iLn2GVVrNrKl8mYtYnmfy5wZ9zrAlG/U6dQoegdqwA37mPIKYYJ7dPwfm44XfX4hDTu6Yv7Rtqm
Hmu3wvTYRvg+7jlmuTQGBOpogMDlwL56XjhiAGGFw4Hz/73zO15KBUR1xJxkbM+s6MR5ifPPONOw
kM22fmxrqeCxiducH/3FjAxLSkfIaCv1uSoHxP6eEJykjlhBZg2sWlhdMj0pXBmtWuvZQxpHQF+8
7mpmEtXWQPI9fIX7JeCqeOhXiycLB/oX4irw0uo8p/U0IP8uzZAyAyshQILLIQHAczy88B+P2O0g
l1j/5pG29vUR0iXEcdvfX9j1Yv1Hyd4/IwGk/Io7PYgGs2t1cVr33qUNUJFZ0WCHVGCI6pUz96P2
bcH5klHpoJ8nu1t50GqcTD5IIFovGOZ1pjHznqQDdu7n3/jjhlLPtUqqjrUK13pfD30KoKHMgtyq
GDrSkNsQd8vVgwC4slJV35j3VqYC2fd8u0E4k4MCIJ/pCBf5uwzAzvck9yIdk9ZLjiLQIdw/xTO+
JBONDw6C/a3ZpLmJ19hrX+/vC5xzmkqhj2o7wtx35D5lc9GffX5S0vc+tGP33xnlvS2H7Dq+sgw8
MXPtkc9kBLeLg5tkX/Vdaj6BbAg9/OQ75tREFuqCoS5qylW4eV+UY4Rg9gnz22XYVhzfSxmrjisb
XHmyUaTWLadxlotVRIFGe0//DwdjEJjghdLEqbrouExgppuYo8XFmVrbYHP61txUFo47wAJQeIHR
ESBTza98sV/29LS8hh6psH1EE8Dc+JEu2NOWgmZirrv7tMiVjuMzqF3b7ru1t+H6rG/GN884TGvy
OdxDw7YZ1VjyaAWi/qhDtAESpSuqPvle/qz91y7Z8Hpc+AbN8w6J/QBZ+hLrnjB1qhInDlkQi9vp
q2/UUJEDqmJk/wRYQzEESjwhoVhw4gO3DbmF/z/EILzGg9i4PFoTJUch4i9bbBYZvLXJBzOXV4aG
GlKTttr8utayXL58GFYrqGGptiHCMbxe9tbiFPY2ZVzewE2iVkID3HSqciCFG361Tqix/78Xvscm
JJ9kyOhxf8SGehHw+olTCrdikp11HsEUv3chDMZ4LUDcNQsZp85Oas8Q+TDd+kmpTCTRjuow8nTO
jIsuW3+cSKnUQ8M0i9/Jsod3Vl2uOmZ1RnZaFG1LQDFBLFy+9aN/LLju5x9ndDBGEv0kbW0jhRGc
L7iASRxZziqFAGdEtCoYMLPgy5lcpDJxEa40Y1c9J8ixCNE8w/C/E6OKLVp0UimiJu8Btv06F6TM
oVE3b8yEUpv1EGfpKUOMysmc1owXhH/44UMaCnpVb/wybzmpHoNCeS05gZ8aahROySTjc6ESl39K
Vl9zFHj0g2zVAeZ7RjOHhM78CxQDR2Yc/xHj/Bcqf2vL8NFJk2YSNNVv732K9CshO6NKp5is0jiK
tb9liS38bgxbsRn3FkOZ1R6nhruEEijIBl+/p5PCUj0jeBjFr4S81T16xQxycvxQZPNxEx01zp84
ZpBo+At6gErx+P+ZByBy16gSjk2t9gcDldu2Ww/wChFY0EZP4APHTtfxPoUkbSLZsRZracIh0i5V
ZhykIV6NmjqrJz2NHi9BgZN5eVkT4r3HmIeTYhhp3o16BgpubVrS2rTjrYfgRx5sSyaART1gFLry
P/uUb0YGX8ZkG8uA3+elzvtpG9SiznyhuLocd2lZw1H7qpC3OHe7WXutf54YiM1fnFpkhhVsR9H1
gcGedEBaRU5n1oTjBna/qsUGcgNI6N2xp+dU++gmiWhNdcjYOw4qeeD7B7sE163MSnEN03NrXpI9
5afExIMRRtpquOGp/+uXraE8QOZjyZVTRjXnr7t9Mt2s2Dt/i3IfQ8U6qjeyNjb08vTs/RD1qUyV
jxNvyQB1ACyucUtQa/q5JN4s28WpKlharm+/iV0mKO28gsRIb7sLhmID69u/3DejRI7HLj1yYEHi
Pa/OXBNFbgocNX2VjJFsp91xrAtks5HjOebHOqnFlE1PuEPuOXctp9v7/IGz0DSFxtezINgypWcg
bm6ANZts3TP1UrW/ifaLsWAMycN7WgG6HB/cChoNI/FWnqGWJN3vfyokdfjokzazVwZC31CXmb38
4S8pKemX6W/VqIrLAoIT4TmLaFoPrjTRHVfOAP9gRM0lPeY5GvmVlRxzvSKQiIBAvd6PZShJOdx2
ek5M4l3aG5R5lBJijhlBYuszdYs9jIztYS9xf0GbZHGINEv0iIAIZbQmGXqyvqxBbVMltLHrvned
E8KYlvju0gPPTX6F1EmY52lKTzkoR4y7lQusXslIkKo6njnjnFwdujUI1TLwkF4/4hUKhNnsgK7u
yFsttI4iSKR6OPaUjZEDcVscXlAocEede8LEVNpjx+nyzJ07BxDy0+UeNNigbBgQ56um8uMYcG0H
E2RGK/Wn/TrtaWQClI5Wkc/c9L3lF/SnF9DGaeG8p7qotA5mPtSz8FmomWvqSR7ZPqJyBbCi6l+0
RqKECc4EgWxiYJBqb5aLQpEptqacdpdwthmWeTuWzNH8M/hdKrK+mw2ZOVO/+TEGYT7WAOTcutJL
w6lR20evnOk5OeEdjeOkEt9JWjNrYbtRFjmVv9Plktf3Wi0XzcRAivm3WLE3751uCBAy3iy2QVtc
jtHO6S1BMDFqAfbcj1l4CLX1+1SLTRSqbtQNfuw8zLXR9fuEuczD7J4K9kDwj485MrKlCLn0cEwc
ltHvTYZjLvbC2o1wT3eLVGS5lkYOvuS/kLvjuKOVlEDaBVa85bBfdP50ndglh5T1nOiua87kwGXw
AlZHGOwNWXFbhjqcjlDHhL0WjBtN+VDi/7dQ6Rpr2IwLpIf6rQen3VWFnF5Ulc0mrzMJX3dsQpA5
2nI4IGPEmPAufTBAzHRxnbTB49h0G+B3CHTyvkddVlyLTSOl9JxwoqCxrz2uqqk9ByGwpTCagqHN
w5TdUtL/dIFGnjHbs++BFbkNSAAFIsAiQgOwe2GT4ElwuTq2dqgQyusZW8X1I1pbNkcWuL/XgiIK
WHy1CGRTn63bRa1S9QNqnRP1kFVlzAlUeWuYeZ6FdDQF8I/aS5p3H6FkNxGDRRDD8SIdEJlyIO9l
hpsmhzT+Tw6JqpehFYBeFhTJaCIT+kRlMzq/hzqMNkb6VX3i2+IB+MJ3AbxPKrCcLM5uHCvPld0X
Ts3M1MPl55p8iqZBeBimaZQic3VxrwL6OKRq+/f4nyG+tSAjOYT7DGaQLaQ4cDROYKcEKCR4t4a9
r/01JJmNDdT0eahxAMZrwibYVcw5ijldAD6+It0qAoIx+ew84MvmMW5xuovbRz7mj7ZZNLWa5OEW
B0KKFlJotZRw145BvRyQrFoyaE4jS9ogT0ahWIWLz6Ysul41aXsLp9BYU9WDxvsbAcZMozA6S2Ko
9ZHo8XwiFe8+HTJA+HuE50PGtQKFrJnvMpr8GsuAlUUzxvjnPrk918Q04fHo721yZHcyDCU9FcRu
vghUs6/EG5323n59w7eUnGoRSTpRRHMi9wIZbDHN0mq+Oc0JWZ4j8PuHy2dbm7qTKtqULYjHyzGJ
wXW5kFdfK/KbA2stFGA/dlpQ9VUIjavAX+XFCUXZNfNTw8t7tVo+9v9tzgtWiEmClb8M6wgkN2zq
F55+kxyrrWVDt3v9G3Zzc0lZsM8b2Dx5c5XEWYY/JnSVQ4meLgOKklOUg8fM60DC6qcExXICLv1A
DE6oGqGUOSqVltsTDcDhfFHc5/UGD/BhdNJPIBnPGedFBUsFrc9GvgNqYw51gLmpkuJ0IM7JKAGK
spRS5R6z/Glc4rQw1iI0trUT+xNm2QG+mHRtKlIqxgJcMUQN6+glXaya9WCVeMlNm9xsk/iglp2U
dFpqnsNWBPGXcCVGy5LshwLeOs/HhJDbkC/qMIQteL+nz65bbykfpcJ6pXLG00FgrgK4GUIr9XzH
MhXC2uE6inlfVQwi0vKcPam060PzivLJ6jEAdBeu63RqEeeNgnELkPehrM9OiGMfOATSpFuq5SCD
3hhyP/6FSEyfy1J49nYrcc/dchKPheAxkSB8vzpo4kkEirjO1zH+oBcONC4jA7OwzTNIwhA8LSyz
n5yCxBn1leU1Nhi4c+v4iidpGU20HlUJ9EKhFVLC9/yYFmHC7579ct1D/MWL/SvNHiRdrBsTyYH5
/AgRtq4Uy03uvyULbtYtjQ6NwNB/7tcs/1e2Pt8FOgUmM5O9Ku/QF2juPhDdprjC/PehDxTh0uDK
AGOwKwFWXrxSoVKkghhuCmrpxbdRNmR8T0DRkS5rSpFT4I84yYXz8fRt5uOXSjQghtVlOJwSnaZj
V6h+J+ObUlkfmT4Z4fMhoMQ9hpSIRvAANdWuy89w98hWifn3/aj3VYb0nZ+J4B80C2w6rhDpg8LN
IWSIu9esVZgQa6MYuK59kXUvSDKGEFbbeFvBQ1zWrcj3d79d5pSuxxoY6dX4Jz6rvVpcJwAh+P/L
v3aW/WIo+3z54iYDVzRKIQK/58V8IbW+obvRDljrPnEv67Cx+McCm/LYBiwsFGgbWKQ35PPP+kCN
96eZbd6OW6uoWQ1caLjL6SFc/LmKHMecC2fGmdTCS0WoToAfrnsrslm2t1uBES7XJVx5Q5R7NOGr
AUH6QkDhlUPtLTr6moMKiSjMWQ9GbPGfvUIIlMqta9PN1LwBvqEGIPZ9tl0MpRkE2amWzZtQQ8cD
oW34BY/jxxAjdGWFILCDqpM/5GOLzfvvZqlKHXPcqyGvV5CLf47/dOLqDCibiQTl5/5P41UIO8oo
zc042jZ/o2t/6lXb8JYgLvu8oNeIRSpZx6ZBYDPrrw0Uuz7u4+sz1Revu9ko798NU0l23duT34hx
ViOyjvCIrJ/3mNjcZ1YZGMQz0yYcnQZxrmlswC+tdSXy7u6rHTi0roglB8Be3zwIzyMvCynB+LCW
b32LnZIIVLWVdHfZmd1ZfIsXCpB21gFLbRnOj9M2gZo69ivJqpDoz4joRRy1fh5Mr+TAbr9ly21O
j3vPv3VJdpSHlAg3vB2rv4dnNX7nM7eXftF0Nov/p5VGxcoz62W7b1kb11K6rrMQq7tHFSVGwLa9
3ONceKfMn+6GOy1Dzln3uXGh1AO9jgJWb59QSR9xEJ3EK0ou82MIcVrUtGmnczuf/kk1gQcugRxH
OLjRtvOtukT8Df7SldAWuxxdT448pc+wJb5jteP3QmDdoEU3e2IQpKAtWuMpjst9j57ctP+ifCHh
7We91BlL3+xIDkbn3TL7au7LX3kIe8KN41geiyB1pg3cahdN/AH+Z+jAz3wqHaVdusI/l1k1DWsY
LBu1QEAKVLHBQscGfka1kD3z+e8looSGKGtat4/JntwShTYigDqUXNLwYrtJNfvunXwaIYUUm0An
mPxR7N+bR+OgH2MaibDXtzuXT3bYo1HwFSvc9k77ykeHIClhdmW1aS0Kj5OLVNXLRScOI417/+v7
iz2Vv2dHfLaW+bl6VNJZGJLdPzyec1ahwpcqXou+KqvrN9LsNGX2WJfo2MMzMJ6FVsk1je+H1ZEL
WF+bd7W52K0NLAuiJ9KMzyu431aJkEYMRUrqKg36D/lG4pwi54KdRWCI4ErC0x67YL2rwlxi5P3C
+iXYfPo7HqW2M0NQ+NuDL345ZfIEjMxbAi/5fGru2cLncE08YfpA8+lKtuw/2MZ9kbMWTp3knjT1
k+sCl4g5Zb4NVqKJofDaHQrNHLrr/lOuw9JLrYpMY9kT1Cz1yNgLQ0zjW+F4GOvv1fx5CzuODQeV
6zGkwFwcNzZQWkJiVUoJJNMAip/hXSyTIO77M8RdDK2kJUWej9gN7jr7Mym1BQcoYgU8kVroxRx2
wziiIIFRFFJOnHoMHw2MPWTMtYAPPNRgoV4D5I1e+fK5VLOp3UfsBP2+qycK5mwY49PkBg6Of74z
p06H/4BrlKzoiKiyxMNFPsfvC5bYat7squhrc0GO2BoqvEUK5oc/NLiCdVh0mOXptH4G8Fkbf98+
YMbeGk9aUC98vz4uzX0vRpmfpBa3LL5DS5Ysr8zQOf0LYKd2TXZEQbbkNcoAVKBfKTyCTA9avXrS
7PWf6e0W6G9BOsYepc3KkmCFXphUMfCtCxH23shLwgzMGYvrfSKN5ww+9kd0uRrNYRCqdWEJvdEA
Ck7EWav66aK8siPrjZB/QPgBipAPRGgfCsmJvjMOoUc3vLho7M6sXXrxjehgVPuAXvJGs8cACfbB
n9NpaPHp6JcUQvWwlXHCcyGIDnJTpPB089aSNGU5jFsyy3Yo2HPMM4RjORoTuyETZJQtsjdUkTw+
3Smk3pCEkBmxEzajWsYxCFmtLD5KYDrux7ph818WFsZ76ptejc1Q2/3ArzG+l4+5tPywerLq3M/t
++QSQ/jQvy6hfyYgVOxOwCUIZxu8+/1Rl9d+tJPx//8YNa+VEAerlDMUHmQbTzvkbKxoN4Xv58h5
kcAXbHqHQO2aI4eAdRqS09OTAokzJkJU0BkS0eYpF91TR+j1jJOST+ciSz6ibEjXOMVfcT4pxhUq
iaPW2G03BpMTkkcy/Fj8H3xEMorssx/FQ95Bt8QG3675SkoGZlIK9ehiadJXq3F+nJYcZjqZGMZM
9muPArF7pVq/CxfCEv6NUd1lhXPxVlQF6PW8BliW2SO0Z92ZpT9/3RdqoR2iLNkHXqrpkyDu2YVO
58dQvz3XQgmpDOWK+MEOBIbKj99cLnWMZnqKLnK8YM4g3RSFK3SPsGDY/Phl0nNah1ELPpDMg04n
P0rcEOFI90i0uChqibXIo+7hlXdJUXvTJf8sq1UMlTWbP/s7m6u2XzUmHJa8yn1QqeUcXadJOPGN
BCcqDhSDM69HrRjw3izIjzVuCPmEZr8bOpgoY2Fj7aJAC2VmPseRg6EmwLkv45H9I8Yoc2kzuISS
ICO146oIqre9/05ebEOHNjYzL+hdUWPGZBRBKwBYMViFxInRq5zRYlx8Lrc4nvkipPeGSoPINIGS
hmq56IhPXICuCPoGZTdf/GGN/DIBqgvaE4/JiogJh19GMI6EO9LWo2pbPuTS1rdy1SPjKJWr2YSi
6thHeAvKFrdYbneDjBQYh7bUdE8KyysgtZEu6gWH08WM0INhgwUUPGHfM+sp6t/i9tDgCNo60yjH
3/2P6Nwy8qY/74x7dZtGlebTNPeTGK9Caf4VGT/EKCCUhML9c7FW8edyzABUdnJTQBX8T0jP7FzC
G517fpMpvI8jDjCN0Sr3zUP0hEIo5kKiOVX9OMZN8yKDk9rxecoDJDGfbVZ15Xkuuo+k7JPHk32L
Yr+bUIy6/AxPREmHlrNIRGmp+1RCI8VdfPuuVEIY6LE7xORjdBdfp4h9kq1LpLNnj9rlg734QlSr
2J47/ZbhV3pM1FWABnwaJha9KqxGm6k3RF4o8D07bQEEM/FoFVzgp7qkyDh+PIj7Kxiywj8+Kq1l
hXFqlB4zxhZoDoisGaMcvHwwwzJUnYoHqw2+DVVx9m4qRH4gDLTTDXgzBLo6HLNKZyC4Q1hJE/Q3
fvNtJ5U9pIUoHH5iIPGzx5i+x8RUaB3vIgZIBGlVXAflrBony29ceYlDGUFnI3/n/IUOJpJPipJH
HUuy66GPkYO4kFSYMaW8dO7kC1oRd7OpjwyIkFiEQ3YErrQptd5e7Q77C8bOzL2181QVNQzMyMvb
CUIscFPpZ3NW78g+3G1CgJ+wHi76Cy62zSsdSuTcYf7R/bfovMgPhzziV0/tRX5CoIL+gYuvDCyj
gaRIG6Ker7DfblHaoerbPTY+ZhydCISWDRattzuxJ8/wirhjYCVUmDNlaU0/eHRdQhIVwjwFJsV8
2DeqgYgdtGIMCuDd2L3Q32ta9xSQxAz2iHG7lJrcD59NggORiu5+Qf5kIc7aAWd2dryKUO0B/Wv6
3rcmwkQisoeDkutA4sSu+UbBHFwg2xlVv5tVOGVqvh+NcMsrIDPFBtaGabkF08XIXVC5ujdiNjuZ
eme9JF6gPrab6GEMLQD3Pb5ubOWJf9/6V9Ol4a66ZCF9t8pW06LzGjiRp19cSa+L+m4UIex8EpEd
Wj6Q0VcWhEfXCVRfkRmatH9WmYDBA7U8YZu9wx/Q1ghueS5SsO3C+AV5BzfMwgQZ8f61uqmxeoxw
B8aKUuJjWCMYZpfY6ANvJKpxCLMZH2CVArxAubDbn8ZUVwSvM54AjcuQPj2AkAxWkyUsZgPban/k
nZt/YPpx0GR80qaFyrfmJB7xv+TOqvL4x0vtuo4tAoAEL+NmfFq0dEUo8LqFNAhY4FGGqxWPFlS4
T4Bb4g69Kr79y2yMI6Ry3ER+Pjr8v3bini8X5OUtcL/ccWINQOfsOY4EhXQau8+ie91h5IDdA7UE
Y3Un8dhTkJGQIkEU9uWIR56XPuvqE2/iAtu0z37yt7RZlJ7xCtg/VgGIJIFkJBtZSwNilFlqx+t/
T+3O8oZpmaOwUho/AI1vtPAZyBmkIidKCNLYmCl69RPpaGJq8BDUOMn72ov9AKGSLXXxOxHbz85w
8cAdLX2VeCDxAzfTD1wK9FXgecsHrwPt9U/fD7/z/WysmXKpcDi6X+Zm41YCiUxrllcmhwKL9zhU
7YRze5dpH5/mVw2sUym7KvKJosXpq2PQXNrVekVHsZOl3QINhcCLN/dgUfZCR0TSze9mbDMi6v4b
KwEudj8/QIoF2HQRjtPsputHO7e/uvcKgE6YIi4/TH6W8mOGCJA0cPE2DKgAR5N3xH3hXcBcM86M
x5nnYA81wu5Mf1pByljW1+LKPisDoaS3r7q7k6BA3HagQEGO72wUcmPvBoaIGT9NrPpcvZTnIfZJ
KGEh/iRAfVg+BvDtAVDu0jdzwxJmyOECLGBrX1lb3SwPuQu/sIuboaMY65/hSzY+K6uEAe6/yZvk
KwH+xuW1GLn6WL0AMOb93YVXqxelzWgeC+buVsbv8JFylVCzqlkteSfYuS/KSV7k9Wn9ChDksMqB
+BRlug3FNNQ536E89/i10w1eVr1uXeV/mDF92gBl/i6g4LozTpV2A9mcIKlJoZCIl+g4Nyq3L5ui
OnPf6r+cJIJr1m/fHnDlMOC3uKLVsU/eBAlEripkO0J/k/DN5T6tMB6BHXfmETYmFtKlkYclRCSZ
M3tGixWYNe4IYAaang6gbgD1HB/JXSs6SH80FiILOgZ5XzAre4LXZTfPzFVdBzaaN0+7YzQEReA8
VB0mWflyE1jGa25s1UON5NQwg/aIYOXhjodbIgy7x5YECPZdaNXodkSEG8I8U2A8cKA3NWVyhhE9
uAGS2CCJddk/G7yD1idx5zzS2YkRDjUZqveLKc65hzpmfCo7KJOGAu5B5CqbNAhbIFud7ZmFX8HM
dj2ikcddvtzMv+BpL3V4m+VSDCukHOOSpj/szlDSck1/wKg6ZAIDbdHaWP27ftwzIDhdwcuSgM58
hPuKh+G3jpXCJH3tjFkbomxdII8NyCYpk9TGwl9J/g/yc1A6VoX4J1JHHguk1eRA6Q2PB4vNWW70
mpZ+ruVuQ9jPU21mMg5yNB4ZpWQsGrDZ6WmGMD5ViWuRSlBa2TQAZkxUJaxLM5e8DEpgSIa2b7Yn
7DsJ83TzVMgz2qrlDqJ8IkLPLSbWrsRBrB2Jp8mNf8gJkQS2YL2GfzdSbUBp5aCaXcKef7DWE23V
l0cgCeNLNVkwnqc5x+hLHwVT/1LSRay/+YKwUdQohG3SPbln6MRptLXR/YTxLku+peKfAHIZoN9l
rQFWEPjHHpqmZ9xQVo9biVY6Vzsx8vQ5yFSkHN1eofjN8OdvRsuROd29XNKCL00TZF0Yiwk/XvVu
KoPj9WQkkuUg11zZVIKOWRiWqAfCGTii9agWlqgrpPlE32tPZaFB/VWono4VnA1FDXhAvExQMNOy
QQtaXYPhPv8TGSxB2yqOkEu6xto4QXw96nCd1vxic3/hYXYUKa04+0z/HepsKTNfxQQPq5z2rIdm
l/s87DNOeO6qlAUMCs4Kus22+r4ZnbKDjvPyYMzTd9p5eFNTZ7PUKTEPvAY66a8vMvgZt3qvUlfl
c0goWLzQ4L3UKuNSOwgWSe2CxbruA4B6IU5brvth39YqrgHa3zP9E0iWmMlNtjsOeOMjGuTYQlG/
GG2aKUZLZ2SEMsh++F5iNtHZwKIzT4DiU/EL3dQsyZtgHcBnPjRK+i1ThDIa6MLk2wYMZgsOdhN8
8xJmcGGIuntdipY/gKuzsDwFfNDbbs1MYZenTp1DXrLlT51+xY/0bGSUXnVpCUWZCnSrPWdTrViS
mo0QgUh8uV+RpD0Hb7PYVcBfHlVmeH2+LKa+nnAgQaIkL9Ct7DRKc1XENfBIFqADgbfpPChrieVp
ck2EpnWtrxwjfpVEmmCmM3lpHUqEmkdzke6s3Rhnqdz7XfZ5zXeQYG/wGCZmnmD0v7tZF/iOn0eb
1wr8/saRCnjg4DAOKLZKIh6+AT5PNYjMkeW13qOIgD3BSAdIRTKQg68pOWnzhdeoMv++EXPCfhnC
A81b6SuMzJfmKpnaa7zM9B1Cs2r4pTap85/b5X/evdPfUShtLvnHq7fjMm258sT88GiNCG1901Vw
hdt+ZUNKYGUpOvk3Yrup33+g7kMQLoBzAmpYp0cO4mMctIYywfq4+vewJFJXxAxeCqyQnoTTNAf9
6wQgJX2DqD4S0v/bqGZx+liTrJBRalrOzgHlhW1l5GiISjcxyhnarbgfh1iFF2geeIudo5MQi5oW
9XS8gbkSDGTbnHtTSMLc8wxvXgCcWbzZIlHHwwZ6wbnbFGg7QKmFTmLQbSy3K8yO/agSJx1WkPVe
R36e2+s4xFkD5QM0bWfilbXH3Yrlhzu3NpwlMwSQOBljdtWj2+BgVuPj5LBcBJB4kQMPqHGPyDkQ
5gA5jcyLEDaTBeHcfvST2/VPcUh83PuhcKy65C2bKTBl/Gd3fdlxDIXjohSvOEjAH3AJvu5WAahP
rMObIJZHugvE0UZfvaCB3COjrgPC7hpC17XPEA+cYa9yuNlVsaBAoMsNjnh37XRsxjBCdZvY30Qk
ZksAOqwvq+5HWuLIIdpRc/QWY2RbYyvl8PRdsnZM9gpsceZrmEI8TfQfwQh5DqfRFYjQd5KBWWGp
FeRcDw0705S5Mo1fBqqJ3jF7YO3bHOuprPEMHBzvEY3NpjRkbNGXUje5CK05uR8jMFoRGAi9cCAI
TnFbQxvQDQmxcqM+Wxh2dCmO7EA+qJaPvTSNhdrwyPFsIYvLjfc58OUZdEQCqdnSO3L3t86Rj6/4
f8oMDSZ/vk3tq2U599NLsrhCagavHKYglFttUDMPR80DbzwDZrB0ZrCipfTAxk9KV+TxPeXDYJt/
o4oiZ1z2Sjnffb33ntXU0QUkxPVxVGI5AXrxBigjQQOd+ehoGX8xKLeNsIat5G1bQbFkT019K1Mq
VpypiMENcpFpKdn7z431c+YgOWlfc8F+Z58LCBY0AVxIJHNrhoiczFxkX4+fl86WrIXrDGeriiCI
OcBUPKjvkruVr3/4ODkQVNOiJZBjOn3g2Xry8rD7lcOLsP9g8wePjH1Jm1o9fe6a1X5t7iVDpEZC
fpdzECaE+WC/fyNrRwpHPoZFqZgj11GoMq9e6ZUelmUW7H7jOzgniFbNryuN/2ftH+JLybK2o/uj
zBeYMNxqh9a+yTbLiWR4E2hzOKTAw5CuM0ycykyF6rZFmQLmuR8nLsq+0Z40tglAU5DQ7yMnyis5
QRN4EY3hzOvwLWOwmbf8fAbMzvCkRS/hziIByCh91ltIkHznLfoI9/pPlk8IPtuWKXPaWk4okCrM
xuRETEv6WdsbW1u4zTluqIDLC4fEkRFBOiuH1O7Wi+TPu602ucY30fSVGeQXtrfZ/8K3CscTKqwY
uwb1aaWEuzPvWjInDwpvg6L7DuCmO6KGxYKzJr1VzDpzjHl6gZDgG2Els8vHmJjITwSTDNghVE6U
znBmUzNyRemOWacspMrzHihtDhfYARYhMlgG3KOCxyO2QVnz2MomB/rLfWisQdXxnZmO9svH9lmF
tfRju3YtGeM1tQysTdvFP/gdSdNQtzw+C8lVXcFcDeSIyYvJUS3GnZ6Viusc19zyS2pePDGXPmB9
ePgaNRKDJChtQ4/fNc40mSyu9nMj/daA96+49TcVgh5kQaF8jrIhi+8mkHJV9SL83wKZvTp267by
52+AkeXu1rYRGtv52yBXFCAnA3ulESQ24gwSKnQgXv4AmqreKHWq1mRTRVxIfxXH8ASv0J6FOEGx
Ne8i+ZKRv2RAokQjNmdsUUMWEDzYG/KTVfVsZcdJYzkbePtfFqoF1pucGhXs2xqFog84NoNiyuAw
PFLqE5psld3eLxi57WrQWHlU+Wy8GcNvb6IXqhaM6A7tK70FmtNvgoN2U8XJPy2vKdzKcUq5+crD
sU2p2s/eP09ArTrhV+fGAkZZvbB+p1/Ku1DeDWU/gYjKqWRjJ83nIpDoaIolOU/3FYJvYptX7k7j
Y1sVv+EKOqjyxXlgxO+4wSEA/7tFUWStshnSp5x4uu9oTyYxGfeKFy3lnuh4eKQ6ur61vTB60/gF
6emE8sbD24m1cOGvM8PTzdlLVS0tcxDOo517YhS9FsvAer7mTrUHE7CWGEHX/dEtICHizxEZnM/P
SRpYl18mSCQxcTqJsS5iTC0LbmWsOci/h2WwUN93tlRXBfyIu6FtYzlzZ4uWFwmzqekiQVyULy6q
XQn1XKWXmcB6VzHW2G+efjYLuPNZcl0kCSJ97WdlBondwp0yusEkVAjd/e4Vykuiq+nW6LrTe6ot
1uqxNh6biF9cjkaUzPoaHvISn4iNy0M6UQzNAQWKw4EpDGkLxkmh0x6+4/T4HJQSfJCcAR2+R7/g
klYnkmfwhd61mMODWncpAwkd2z7jsnVnMd6NGf12wzTWBmJjI0zPExX4rAf9Y20cHyUNoGpY4+0/
W5/kTZsJowx3KzETPnY2cA0woos3c86jDHQjjdhX/XtgqTIKw0eAUB5Jb54b0ieWPrtyHpSBxAwY
pywS29pgEhEa/V+mQgdQvsoHdmZSSgxuevrCmBI+ke6tE3jWOqerrASdTHknnuTJMEryuMnF6FOJ
1NUC5CXYiJ4WCcRvECSbrM9iYRmzU3/O3YyyNnJRWJp5Q1kKLL56x7+EdzziNGWSYIliJqJBFXM/
P/ZKghdRpK0f2/yVLtCcU6lW7jeLQIpsX0RuCghPU4sMLpLyQRTs8KiB7/mnCi/4Zx5jnriPgK1x
txgbngcwXYcZJQsD2zhlS4D9Vfm1QTk4D1+b4boJ+D93bj5FoRbRNYuCOxyFIdm/ygRagKO1LzIT
opO+varj/PUEvZI8u6jIbZpllCVRlcduBuulZyoia3o246wRRsUfuxwpkpGR3XRCcL1Xu7IbAH3I
/y+YhWCjo+s5cCKgMKY01rHyVpgVQO32bf5VKZ7nouMl5+72rCIidISIzOxDrfySlTNYmTSGcjXH
zIz38bj0fx7b4HUcSstHExH/FXpQ5vGpLw4LR5LWTMI0aWf9Y8R1KUK9tfaUE3WLF44sW7jvTp4e
lb6lPSP7kcM4qxgreMmG7bOVrzx3NiomJeVOrdu5NnrdekgMcwmHM5yLrpA2jycAMojujSShC4Zs
rSpAMmJhqWY8yeh0G2o9dRUvg/BWZQbzrIACb/Fzz+XXRa9nEX6M8IwfMeTXMKPHFZkY/A6UM81O
oldmAnPo+YeP02C7OM6HrZU1pepOuB70jJpcQuN9avLHGTdNpxppoCMRpwo0h4tJFiSD4tM9dp9B
Rz5SxS3juhXFVrzoUiHpOl9UA/BHr3S8TP8GT4XZNBUB8NFRJiQbv0wIYfqMddX5SX+Q2HeYXXh0
KvOeocas6mxafEmRbhz5fNfAQyvBP9f7xEqZj5LUWv1lJNFUenGHXDj5yKtBOKfupMBWb1RirIK+
VEcrocnBYN/B1hT32IhT0tOtXzfBRPEGb5Mq2BnZy1mOBi8dENUNoaW+P10PY8pW92LsMzYYNVLY
2Z5I5vWzoyVw7k4rzCPzjcgrad2Bjf5S+iyEEWvAQQhUqMr2OxCoOAG/vPO605n9HLXtUSZLoAZS
u2FFhTgSESwSDclFXLQkem9ltdsDRqJKubx1fUYigblrFQDlpIsRCYpVjeRZAj46vdwmLUIUdNft
Wj3QrZeuBO7eUPm3NqTELUtrxj/oDIJW070T0RIVD61Cxs8DRvaym8z/ObndpwDg2i/lq5qI3EFk
DLAcnKLINlxVAGZ0ApnWb4igUUZwGpqu91CiSqC+7DEKMu7uTT9PVPAs8/Neu2BRiK9HEYVFE3Fv
H12ewo16wp4+fOuLU8J3Uud2Qd7I9uPagg+uJ5e4VNI//LlP6Ianekw5JZPN0Jy4gk8K+jtzBokV
l6jPLT4bIDiY8cVJalp7tufe8rwNST+4Xivi+Xx/L7cBkETH3ssKY7qzlRf98sRUH/aMAoP44INp
bh4ejmEljfBbn723+Am1+O9/nT3sbckhP3s5WWfvzkT68i+35/JbpXLIkLqS1/ZLxEtoHhdanGzy
EJgzI4shFB2hjrmClkgV2ZIQbphzjgyYxT2yh3u6ttLB5miTP7Xs9c54RQR/M177Lb5gTMoqTnnR
K1cxHcnqMWpPvq3XStY6Zj3DBFxqLdz0RpwwxV3F16nM/s774cmoOuGs/yxSSCQAKRGjELmHOc1B
YYLPvH6CvBytTlWSFu8eatnTrXZR48TkvYH4Lcz5TPrSpnDu3/knVTu5TzaWodEyy+Zx8U8kLmBY
ZlgIfbW7Glxt/2RsjbdWQyPtfGDspa08G32dazgWGQ5alR50Xzz7duW2hMeHnZ2kOk9pvue9Xj6W
ZleK6g2pEVgDYrF4B3YgsJGkFZc69GX0RxVd0/NAfa2w1OYUYF4ARLY04SQAHVVz/olub5U/705t
tPiAHr6yJlEH0OCQo+0CJvM1CgvgBk4BUabRlE7omYNBcKjxvMbBlRix1NYILWfM/BlKeNRuiGF3
r86fK8MKfEbuI+EJeHHM0rG5jyxuRcBFWXQJ4xvLgjfr4f9+gE5iGvyJCKMiung2CDRffaFrSx5S
BOWZOqjlo77YOB1gC5V7AOJFv9PybBD4NsI9bC1GFT0+0/8BabU5VLTt9CyOQFVmiZvI6F9r8Mc+
ogvJJkglIQF+OsF3is56ToP1AwH2EaUnsY4FohQo+xHysyMsTIH2tQnepd96TQQz2ppKzZY9VTU3
bdWoCDHGTVcIOja2NS7oevGU3XsJwZdzeZPCcc1AnRN82UCqj9FbUV5DEnK3d5b/ZAb13qErc49X
KgDv0GpLjH+r5wJfLUUmfJHkyyGGKdgkLYR2Z8u5GMBeUNWwPI7EWCcaR3hKuywjGjc0f6DOVY7p
h6YKLx7mWQTkko1dLWnUlAZsy5HGnWSjMTvuUv4iGTS7Q46h/3a2EZBOhAEgifwP0gIEe6fWQ2V/
y/Yk3AoeFdThKJBt0aWdrItpgmOZOqU3UJ1yrWK2rY9lHuBzEPcED7mhG/h4e45tLcIcxsbN+YOv
AxnEdaAZWa9LAOxeqz4OUJpWt0HoTzZdTOjxoCfykmUPrk1t/VI3sWJJBfjuGl6PPUhEBuhDZIrr
7Gyy/nXE9Ln3Pvhv2lzqICTKo967Qy5x5LklvvrQHUCKNGCtuFUHq6PvTOPAVFnlOJhX0oi/xNod
uLkJ86vYF9i2kxHQf3VsS1Y5DPdscYPqApb0Ka8f+30GWaZysBVWSaUz71fOHjqjdsaRUt5Btem4
WEB5vqC6NiSiBpkngtUWCVC0K/YJ188/OZDeRWTUBprsKIni3XfHO3tRVNEWjcFaCUhNLaDU97jR
80eDcv2irxsCXwZWSz5kb4JmriB2kw7yM7mUJnpk4TtlE+gtlLY1wq9qCouKHZZESJIt1SbTcGyd
wGuDaHw2GjsY50QcTcLbUgBqNe7MGyoQmyv8yuUnhLfyj5pysTfw8RPaKpKtAXSb6NwQE/l2s1ps
s8TNDdnsQDcyfEOeyacafQWUukhcrDLKLfL0DzsQ378WisLIcu9ZH/PKm8/CzUp0+Mscb5z62tJe
KiPK/SxUO3BvAuUjblc+kIpmTUupfLM/WjypIU/YY0Pe1xSQbwI0bzNTJP9vB+fz3akQk3UubFkF
VzyIZY6BxUN+jwDpHxaf6Rw+4Zo/SlWSRInO1rGGnkUYqxI3zyIQNvaacod/yexN1CatOMG3ceMU
vL3z+LjE7WRZNBKYHJ70VgCVZkSu+U+aE7w3UAdb5xLCjhb2bVsuNiKpDjVyHM5odcatj7ptO+gk
InnWWXls+v2fxYZhhst/Fx4BN4ZXwgpFq8rlyujjmGmrnK5UUHlkrdwv2cESCaBc6dlhM8GhhAGB
ffk8n9tikWWRQmpr0u45HfMDXULPVG3ylFC6seSbeuInSH9YZ8zLOZn4DB0T2sGrtIFL/Q9kFCbs
n3rXl68iQWzEcV5Qyg6RdNoy3ZDIY2qi3wdAQ5etZtL5j+j3jK+0Wr2fxWjG4J6dFk6+UgU8nwxC
euR7zxnc1UAmqglWCvyL42lkN/Gv7eDevqi9novx1bNQu3mCLX5Zs4o/fgGnR9binyMMWhuQiwNs
8ie7sBYOsUeNN+EbA4d7XFZ3eMZhpY01qpLwQLd0M3mAAEYVhuT/3Gy7i2rV1LJnfkr85zcgG17b
zb0ivO42xPsgLE+C0Xxpb0CJn1Yb7yL9xONviL8vwHv0Vx3Mfs2q1+27Mus8NwYKMTbDcrVP66Hw
G4GKVHZuPjXP7QUWrpWa522itvydzWA7G1vyFUgOmpCCqxz5X/BtzwBRfs4tEYNF75Nxwmx/3Jz6
JxVSvbuYjwO+vmQjfn5ajZ7U75kg+1ZTVSj8wKeQ2ji+DgQK2b4aFIrLMaDrR7IRcJSoUsLceUm9
ylfMiPZbBIXSwJo1AkOeCmD5bi+MjgR2l3FvufyXXPJb/33ujUwjYziLdMd96mXlRNkyi8Xq9hqi
O4NHnyy57R29USBRtOC5hQ9Q6YW11tkhnjbRZNvBlp/Fk23nToV/G2jctRLaHEU7d67SMV3C7MFe
5r5rVPymXypvFPQQU6RZfC6tD8I+GfU93fUHi/CoFHmyMCem51IVpCGxFa5NVZcW/XEUVUn2jgoj
xcdNbqqQFkOrkW43637oCVnl2Qx8Aj+Mapme0bjv2mAAj6IZFv6lWlxFceduQ/XzPLNEWbti4u9E
PGf4WEAv8BXhr75u9+RmKH5RAZxVZgNH9J2KVrxyPS3EsBctRVvsK3U1wIk82gwQQ6YHZthTLVCR
diwmF/rgzRc+s64nanABb2EHP3YiWAxwK1OZx33pTJNoCPMT/wgwtvjQtm8YTP+BFG7UaJX++6bm
tf1i/pQSPdX+875CaiVlCGVXKg4PMLUSwRlFk3QhwFS4BjO9r5h/C+NE31eWZGrEs/yDp4yzU1eh
I0qAVc/vzzw/HuEdbet6X5s1cXvM5Hh7gtZ8MNZgCuoeDvjYWdt17wzAA4LIJV3WTZCm9ruW9xIA
xaWf8yr5ShMC0z74qRyA1aMlAuHcAxsbC7KJzke4DbebSFWBUXqKzZSKwQ17whN+lfPfkEx3UoOU
uBlPg7j4v6tfC5TqNOodFsmH3Bf0tLK2Xa3mW0sEDR8G3Ftjp+tVDqBgMdULKp6XylfURCf0rLm1
jMGatTOZbLSLL395MJxAt+rxrcd8XeOmODkIUpQpgf1YpAh6SNlkd+jFRHaZ52X2RD7j3bX7SbXu
XtpEgXwmJo68mV326WQMhseZVQMiSm+8LTiSxm1G7I3h6HFF8Fw/wPEi53HL0uVydPIUEfsKHjgq
UUaMubgNBt71jwonijt4ETbZUbz/ZT45aX4HeikN30OkIFYf3GHqF9w1hxqXUw03pmLKIja77G02
x0zLYjiAKDh8mQI2KNJQhxme2L75GH1j3cPvrxJoZUB6smQccIVTimrFCKtbsn+cb6c098KbrL0T
gtNUuH9Qvc4lKI1MU/OYzWZyAMhxcm/0rY3mJSz1xUTiKEZ2dbH4Gvd8j57gg+6M7J8jm9s0zS/i
E9jB0GA0rsbFwigcet2CLcIBGEhqtH0gHEY3xuyDgYWhumwbFLJODgp1gOsNYqjbRyc+dc6n8dm7
36Q7TEPmb05TpyTXcgJuSUVy62106x8qT2M4teMPvFAjhbgB77Owh3AjmuJbKxnQGJAFoPqFtXc0
JHLhSGzLtPzH7khybu31JWLCAtHLcpfdFJ+At7h1mLvRrIqe2fcP94o8YCBgQbj21Xgqwqipb56c
Tde0rkA7kJ8EwYigq7aiNZlYZGiFA92cVFuliRIklQyQZFv6NVEsuV0OR/u46qW10IBe1qGWa422
wcRp3PDeNnyIgMqd7glZ6fw2XE2h22xb9aBhM9W8de6U8ytSA9TyGRV6hePORFCCV0W/VQrR44G7
2ivQ4R4vZ4g+RmEF8CEbfe79KVQK+q41k1Ik44diRg4sqkAVgt3yI4A/YfbC3qitNOKaPc+wErQw
l4AmfLoJrQ0/OMH4Yf1CQetB81yWZaMqGnkMeSjdo5tYBn1YtcrlYnvEenAb2JxG6LOQqbTdvpo9
9yugmSc8KkJ7CbhCcrA6Svg/5PIQURmFFMZzWBxZydWsXjXcOra9iDEmSrpvdjV7UAsuPIiKqaCk
HCQucAV7o0efgZ3x342OhgkEgRrJ32qZYSNakd9jsMWmxUSM+8Vfa1GSB9DOVXCbY5VUrdkVGeEA
3pvPlsclWiqhGeQ8JvBuY6gtJyxzSe6+GvnsgOB9yBWowS5qynQmrr1o2scbPw1pnwtylzJU3+A5
hYBhe1LXpeikBDCda3ozlFpRM9HAW903r8SWNWcZsV5cIuszZkntExdPzb77iE4WZLsGIV0DJIsD
3wbDz8tnJzvaXFokNxVGczFru2ovhcVeq1Da2q0CxjmGlD35vgV8KM5rNDe23WCv39TJQ0bUPPTd
uJ8O1rSe+hXn0Vy/6HBugKWcicmZAdOECQ+kWOeEUtBKsCPDSi0RqlU4ryHqSnqxCqE5cxUbS/bc
o/QijXsrgjWoMw9PfihOBNBL5tUmMogftN/2d8eR3KlrY7cwBT/LROwVYp9/Ond81c197Biqa1yK
SyMFXxwHq9IH3HukGHsXv1/WGhdMj6r3nov4+BRMT59Qwto1xgTGAHMcx+NAeAOFzqYc9Oi0mjMc
TbEIbzaZVY2gIBNCzT7ZIvNnXQQ6v/XusvB4Mcr5AbSIq7LsEJhsakpeFmUveXYNYLbHUtKJwcNc
OwvKxZl9pNZlLx7upLGGVHl7KmuLwzMchQXmAA6qqkl7+STO8qtc5Ifu9JBM+ISSjUE1/SyQZtE+
JxBXNdJmdV+u+7Z3MKJz9ArXBds/r7bMOQlmSItMnX6e/pV/eAg+jps7XG4AKZYxusyQrRxooo/P
SPZyLOC0wADizQBLouS0NK4hhqr+7TES+6EuCt9wRJAemE3/JrRkUq+oZ/h6dl6qIOukXdGq1tF/
eqIaGAjAkZwu/exhHpS/RrOss1XpzUmMGMsqvSL+U2JsNjIzDb1JwF3EAjvW7T1Xjd4pzcCIk1MP
+qZZOTbOacWXaCq2ld0N6Q3WQeZv72vfydYxBoUYSTMwjtZK/Q59QqSh28ATPqVWiRUOzEDbCkK5
PzccfFAV1GM9Jduaqvfn7sAkhAJJ1pG1gle0ArDdgqlablu/d+a4Ng3irlaXfJkap8pHU5J+QDvY
g0YtNOC5g49H+NGDL7pW1Wh9CjZid2XYJNI6jSl+Eru978xIh0/6SvnMAsqEc0k/++ZYsl8qOhlU
dLNUd4+bT1fZz46IRvo89anGtj/1iskdNO4FMcO5VTXXaA1GcPOWH0NH1DqfrXkDB2iTnQpiWKWC
lCXTzBe+cSMkLa1PRVyi/lZPw83tScxs0emGX4nU3e502P/S1nJjIDtlc639VwHxFq6gs3Fl0aiP
+ya+sVXtvYGVtogG8+w14oPaFRF+t6PJZQAc+WGnYoYf8CBufIpLGGNl8tb8tOYo5mDGace30qGY
JSmDTP7ni0ZydZB3yvVSC96Yfe3x1LJAsUfcxmvD+j6SHhdipzlAoGSS3QJbqmHbLgnx2mBORccO
ExrR2DV8b+fhA92M/GLoln56GPn74WWQazLWGQg8n4rEM7L44CMcFIiJm+WQkEowJht1xin/0Y4E
5AoBspUqs+dR7iNGyXku7pz+rRYFcAdD5n6eYbdOlEDKm/tyCgLAYvBb8F5UtqSm0jbeLIE947In
3qrw0L3NhUie+vSAOgQtPTCj6DCjvKqw6IYI2umJGpMT0e7bwzsZv1BGaz7vcsuWPhqA02wd787r
/56hQQCWloXMvGz73+3BpKmQrfWAJHc4RhtxB4vWQB3vGMxw8RB4s9WCrJ3HwPDWwzA8pfPpOJOW
wbjeUtrUWmZnxltsstuQ89YdqR9Bx0qIo/+nXciqEK0+UL+uBCEMyCx9Q9yLjy6NfxCcCLzrm55i
sbUXOa6zOpg7BXpzSY5aTsse4dsxbxQHNTvjgtM95S1I2Tcs7tdVwXBWplkiVUTgcYRbacqnvgsw
850caBhSJXlN+xueNKQvx9pkWm3FpM2ESCDW15onrbBZr9d/6IkGbkmKFD7f2zB1lXFvgt/pVt0+
4JYaGKXfN/rWqZxyMjfUpKq+ob48YlzuZpkPDe1C4VroR23e/SiOZmXXMHo8faPhb/Y7zTwHdwtf
zmjyr35tjLVqo9lbOBmo1K1ZW5HknLbWIajqI+vMRQqerDdEPL/bgAzwousli/KuG2y0OLPwlfqL
Kg0OBW9f9ty76tjk4pH0dr5Y5N/JPwkfkLoqtkNQ+P2o+e1Jlu5U5gn4TMWcd6K1jVjw5uRNe6+4
CbfjdYYiXUMGKWdNg3Tm7CsJG7I8YF/0Ac3bnlZeXaoJuClM4yTXsJCpGfXdHchUMIS6RyTRqmvO
jWuzh5RplmDEOp8N2X0/+aSS7QksfxDn0bbgfZtlDa6IzMAm2B4krKUGlLWqjcy9y2aYerzoVjXo
kbXq78k8/RBLkP2b3EbIaq9F5MMJhXX5xcATE7qObfneQxIHxvmOwgOONS2QdXbyog4DzH90sf80
+ajWRMeiLTCNM6qOkJ7tKSlEWXA3rNlr1w5/2OWyZeAOGpm7NzorAntQ/HFL4badLnSjF4R1Lm+7
OYyWsoNeN501SriWezy+bVMEZHtO9M8+JuJTDrGQCoajc+tvTQlM7JRsJt2C+v58qbuZNohBmkMh
xqu7MvN9ZgyRsnG8sUCxhg3u6n9P+XMncndmHeIostfrjoo4VzGWAxBe7UT5cMzG1uJis6p6/QWK
EpMISO73W+dMt4qRmnv1hr1Sp9ZS9liz+UGKTdoc8kTsAssVXY4uRchtOieMiVAstYDwDtgBMwv7
EQIthZr+UzdrLNKRslCy9B9HMDpGqkKErrG8+koyYa6/5PrBoYK6/tdrVMVV7RQScUlcuUanlU3F
slvIJ/h2ABGpvwwBlI/dEUjZ8nv5HXTIiM/EsRBzQZddYxH3aEAjgcSn4qttwuFQHVeLDIqcNhDt
TYHD1nBAAkzcTzNyPosZW5ag3wdFSuKE/SREMChAyXFp5gq3uZ332n2FC9/alB9KE9CHevxvoydV
XlKGL28cDnHLC2/MjK47OPj0q7sqSTnc5We7qmcYRlVEUOTWiQCDEHVQOoZ2iIY5BGfp/yu2VCO/
FKaU8c89V+/jiaKh+oSs89BrYDMhIHZyJ+ye6jZAlg8RQDA7pw46alaF2E33JVjeqmpGkibcRdPE
skxfG1r61R+bYRs478JdEmk7GkrGX+YpFnPDphi6+7qSpVI9vac7JJR+aqrAClElMnjvygb1uOHa
5H5hcp9B0h4hYgXlLTawM1mh1/VAc51WQSc0Yt9xzeqy+VQzTDm+f/XOW6C2NTPKKoR87k8vV7Lz
EaPq12rsESo4/SPgg5WoCVC6lnO0VdGpj0o5bfta+R4rEvpx6sIQ3IehpNXc0cW9GR9UcegIO0Gk
MTLSjyVpkGQFQ1pqlvIGZWhLSeghEnilm9bik+7aH9JD0YYrwPmLHIB3tBfCW940Sz0avimHJAVw
slbqU4ldV+W7/i+F75IgC3UsetYnWmL1amXqB1bi78J1QU50mrAMgIdC+59rc76pMcOc8d3CZzTV
Mtip/ueVCwbua4T6CYWwolgF7PavhJhOQMNSxpTdCZkkFQ/dv3XtYU6NtjqgEmZEDJkirDSMc3ta
SS/wEaFO3dEBImwbxSgd6ppYKCV90WvTQR5/iBJlhHvQLsEanRzOyATaRePVX7uD2oY8Mm+Zeryb
Lq/JrBS4tH4mJkAOGl4ymkEEX7jT+I5r2XH+qcmRxgKCqQbBkpN2k2yWkG0fDIv2iASO093BOv80
D9D2DqnQ3Wxu2Q24EKcZLJUE/U267GCUTlkIb0sWSwQZcrNS36hMtn0euMO8H9sIYXfARaGXXzS/
3Ws/zKhsMgcclmU0zjjO3QAYecbVvP8wmPGmvNrnw8epnjyNHkeeaudxBVC4xXYrD6fMDruLi/Ez
qmJ4IrBAepRz+MJ9Gkwk/Fw4KoMT617dSwGW03lT8RevSCQmxfQq/4+1a08nGLpIJZdR3fFGp6jI
2RW/a6dGTrx+7mM9OPEAoJC+ZEXYu/JLA/+I9gsrNsShcaNWCZCOCFewaYkJ5Yw3GsdT4/8yjyLP
IB1YwzuRNeuReJ7FgeElFS00vQwtdIuIVuR9lmbpYXmZr2ypyAqU/FOkvd3+pcr5YbN+iDCYxlWK
n8/9WGIq3lpeZHsGtoPDYV837JU3umLaAypUXBPQ+g7P6RNfaeWLFOyBWi3K5A9XnOGOfMPf4Oee
N5gMOV1hMZAgxLTZv2r4lwLgJSAmOXFiR5CSXBcXIBPgH6azJllzL/zzZgPSSlCdkBIdmBlCl/5w
XnDl49y2cdRndaLVL4VSkfpBp2YRocA3kseLaXFU0gu9cU4ARqruJMIuTRbpBIuTgMH+qa8TImV1
mKfDR6G0mjA36i6hxcsJoHGirMdbedRhll+HD+U3d0HYjruVP5x90Adq0gHIic0FgA1NJp/cz+RZ
6wjI74RDbYPJooyiJV2az6hV2G46bym/j1sDUGI1MNgCcXVZYyW9h/W0/IhahjcZ7GVGoB4v2KeK
t+OhS1ZjdBgvFfaSIslY85IUo1CCoLyZwv5n+ivTakUgLNe1nTtEQZuzaTv7Q3Wgb9GVB2UyxOGz
wNjHI5BAKTkG7V6n4uCNdf3G4KVYlOPibx42sX2oSqqR3pS9JlqnF/WSsDplZByQKQVzPSfnsNRt
J322EwRv468AhHmuME2oAvjZMILgiKXjZghmNiCz74E8cUQUlm0nmUKVeVfFXMDIvVPAM5uqvm1W
EOr0w9HPYBX3LTFwLjUEADolmcklJFvC8noaKdl2aFdFmqZxQYC7ZLKBC5GwhklyLhwjtvjcKsIx
HCPtbCs0BkZFMYbiFhEKnN7HQoKVHF9JPs8l4PBFbnfM4gXcCeObyEGREH7lPoQ0yiP59tbDi6Y3
mHYpZkw3J8DX7oZNaOjwQ5w2a2uj4TCq1Zr9fpP49svRpok7NIBxVgxiKUYpgk39h/07JUdB9IjJ
A74BGuQ5YI/A+5BN69XldRssDJsYgB0rSlXDq+6aZm5Ek2RL1Rb6tmzIpqLOn020mIsV6Jiy0CqN
QTFCFwPDkETxDCu0TefL/QRUXVWfuWkvPb7afhcs3kxH9LmXYLm96MWrw/ujCQz5MB9ZRYV5EQWZ
3wbP5qrT0nOD2QEiR8ofl23kLeLeKNGuoX/xUsGrqzs9k2K4PSc9YbBSwpoicQozDJlIfiD21n8h
ih5qnus0ofUEG3ld/5WmW84sjsUqwJzwNS0wghentXHsecD1/Db6oR5CEg9R9svM2dgXhll8MLLL
eNFiAwp6B/PuM5/V/iwHmkDkcWVIvefQMB8bTX9Dd1tgS6iac7qgoMq3fT62JPeSaNSyXTxiPA9U
XtPfOOY4BXgM0Adf5xJh/twx5BbyKMRmq6pf0AV4vTXHFiPG/xTaJvrkkXvJ0a3IRCp/0LQe3LAK
xmgsfxIY1+CIbNBjCSqHr4PWY/tAMJA5nHcqvJwnH2JAq00C18ZB6zgHJFcGI5LoVE0MP4qYvChr
7/+puJJLimqR7mBR+6+ZWw5y6NZrvOTbYYZgZBVhcunWa5cuZ6aoWN9DyM/YQSy4d7WXrHE2pYi/
Tcf2KyQ/hBaFuFfO0PH56IvXfeQkVP0mTxdIz/j2RWVQOSjRHkAyMxjDLVbiW3UGtimwB/pxn69f
sj3SxorV3wNBSGfQ8PWCwn2Yx34mcFjuCLvgXgdrEItsIvPyH1vNoV47Yil253sKdVUpMARCz6+I
Om8wEeM6LqSy5Gb6DqjepB7Dirn0Zr5SuchrvSZfQu/dU+K0S5kfFEHoLahIVhjSK11GzwSDc84V
P/usPE2L8OcGdOg3XmRmzDVQB4ca0iTGujvCbJt9PM/y3mln7CFGAmKK4u32tsawDDITwBE0CySx
UsCrfYA1Ak0/wxWlHbOS3mEbzh4CDKpRhtPwRl+iVeANiKyQxYQsxcEEoHR7t1JIQsQfWdnb0LL+
I8uOl7jXZEkuCocKfqfMDCplFQsQ/uZ2PHIv62EgsXfjpOTxrS3NUzcwrcEt8EXlXl1yPOMgf4gC
r4yjwX/3h0AFgkQAb5ArKw1GQ5ozy0h0vvpjTsAJDHrNGSE12qxaE4L/DN+Eirg/XM7LR0c3log4
9BgKbxK2ag4NSWLHxzjK56IfRknBm1vulweCgLDlIOURZgrLeW+k/8BpOWgJYxJlvmqqkrCK2kzS
huu0sRJgsOyyz/BQp+/zWxa5pKSW48LyRKfNu5mYer3eUByuCK9UzYBHOADKAaqUcaaujTO1zut7
CYA6PpMEIpVjZ+xNi4kXb9KDbIU/Fycdof3qza6gVbH6RIp8ktzTxXtmx2igSfN3pQnobPkXclqX
WNm6baNJiEfwMivlTgqbIjR1IZ77ifVFFHFxY5xKUPdlrFLwp8OOGPCZkhzlZXnxSfJ3g1O+aQl+
ITfWwmzX7mC2HEZYsNMnkLsM28gw1wPFi/SPRBR4SHpr25w5SwYXQQvRgf+LyKt7DErSaeggCBnr
w0UfTSXp1cT9Q95HaBfQHdSyil0x1PeuNLiRspunDnz/IE3BH282XTnjsHTplLxOGKm4V+CI/b4R
iMtvmkqF6Gq/XdbqnPiurKCa2FG3MQwmMrDrPtIS7oQ35PZqBkoC6w8InyU9FR8LN+9Tt+PbGseZ
JUOI+dKRVSdMpRTTKiL7UoCG5u1DI3NALD7M57n/n5MxmIge8FRj/xrG4Un8qwlAnLx5uLGhIBFH
s1B1PTdi+5B2Ls1JUHqhkJBimjRhTP4tjVIRGqJpaxcjQzjwDR0zQ27OWAvDuBbSeJwwrX39J05S
P5Lnxp5O7FjUZomgBcA+PQznlM5vA+4WXDl8Lbb60OYyn/073FbggVTOAQOBw2YFPfuW5+844/Kf
e3dUlKkktn/nSLg3sgylRPpo/6q2CwVQRoddU8ESeDd+zL0goHtsPyzPHgrKdHHDDlhT1leQJ+58
2MMQtxp1Gwk+Uj4qd2EnS/ouTS2wNpWTNP20+ti7xJ5IzKHAaI1BVtqMU8hzXzgjF9YA+Z7lNLv/
+4PJ2Vrzmc3WcSAe4nnJZ91h5E8NyDug2sA1LFTKoWhc3zCZReAbdxgnBgNlvzYK2xDjzLqisp4O
KrBcURAK0/fwKocnquAy4ahds8e8sF2ddE+Y2pYXm5ACV3HoL3f3ile9xyyY4IztdDHtmMbSTLtw
/HtGna1uC2nkY2mjVW/pwhPc6D2rx4YZseHqI8fTHv4ECYmZ+dyLiciRRnbwmgBFiCCv94KXxuaJ
t3e5eWOMmUORV1LUMBqbLk9qor2qDnQogaVttdDAvSVAf/GZjj37Nm/bTyON9hWUslVRUejlOrE1
JNFS8Zu+M84ZhrSzWy8buOr3kKOG4vmyFUevc6NJJuSaJ8V4OtJDrLiw5z2tVikgWdCSkT3MKeaT
wKUxef9Wogs/L4+lzXSP2iIIds9tfBzEkpzMCaKBrWWTRos+25IOfER5Au/+ZqpKrB0AbVmXCsw4
/murVFHEvmviTyPhhzQHKt3+oC3hmPatTh7IyxGOLITmcLDRwWM11YxBveD6e1g9fIfw68Otl7Wz
NCvDLaCKZImuJ8BzMVRgwgQLzAENizgpyJAF805yEr9InsJpYAb8R4sI/wpw7W3qyk0ovTCT/tet
n24CkGlj7hHuLDt8ngUWimX7Vw0lqrglKq18waz1g3bqlARkQkJnlmEwZmXDIdsUH8sgP+rx85ip
uaKbz8omYMZbaAV4ieUEi+uNyLwRd0UtK2R6e+B0wf2dC5NgOt968I1e2I79xETPJhBPNsBbsfWQ
bqXTmV7Oi/4YthauxrO8dUFN2uTYZGmZ1uxo7jnHsVrdgX/eszIUoSk/8ktXZb7zxhtkYMrebrFy
PbV2IAzqBNUV3Ep9VmcOitc3vlk0AhJtevu17SMB1FtmkzHHlydzUIwHcs6E19/1xtsQxjtoRVOw
4xB5FMlJqQnw6FQhhL/RMHrDCTiMNLzfzxvvAvY5VVMOyOb6farVyWIQ8TBo3V3UnXzN8vmrNVZn
u8cbMIsZtF5psIRh5qjb4bLEduUWBw//xT1MLYXQ5CwoO+eEuu2QEevysF94/pHojiYlKQ1elNyt
iAYAzMEOT6r9cH6EEo0ncgtwMJGAE9bPD40k2sTwHlw+fX4gHaB+tLmOMRmuJ/hXOiX0M1psVyeV
+joUz/qEY9osZAN/Me+o5u0G6ys5bMPK3nYXetd2bd81v7rTUqkwuvYgnhVFwXSfKXTpqTDTTNF+
ZTT42s5hGkYd5arA/87EbPD9usGXVZnyGsxZZaTdsg9eUnOsijW87XUyIJ3GjcNmJIKJKixgKtjc
gOZDTx+LlCrIk0frdHBJkiaa519BokWzxHDGW9dLION4WSTzu0918Yn4Rg6JlYh0QhGOswmhS6xk
10LS8wGeYaEfN1JDq60fHvJ6HcXKM3mLgMO0HsYuxiTuxNzFdUiVnocMEQqgSnggXrxYjvYwr5YU
GLcRCAWxnac3xzPmmo3h2ItqkXiuKHPv9is2pmTdGMvSCVSZpoAKu88iBRTZax7iL951KDGoBQJV
i2zRT+BbANJvHg8U57fRWSEjzkIaaQYU9YMk13P7WnLLuQxR9TGt26v3JcNCO5evY1cXkXrCFqUY
kTELb0uNdIFlvVzB/bz1VNypFDtbanL8g707qNodcpsJcc0gHn4d+haN82QRrp05NjKht1rzuFO3
oNGjERT5rAJzoVP+bY/PSBZtpj+BPRtCEezesUWgDVWgG837WFIJgFAQgkU0t+eIMMO9TzXo3HlY
UCGZfqWMju/B3vCBsMfCFqmqZbO+u4Hz/rthZYoxgngQVyon5Dn185/dcYTiHvJuJ/QjlNVEvZXa
7TAZ75uN2/Gs5xB0XIybMoLASFtQd4WmYUQZ6lBFLZPOIZYoN3uLIt8t8cOtagGC2eU0ndlguqb2
gWR4DHgw4dCkQIXRgWlX92jbOgMTkRMqyvMwpg645LE8CQTOyfEQilf4XahZ0YdmjsYYi59uHHZe
3aPTAgUZA61GqPLgk2h0Fmexec8ICcC17eTxImLUwe9SuOfHjuA7sGCoLQJkCT7vaYgoFi+AYVhi
TSkOT1ZDA7e3nj6NHrL/f8GggQ+uUxAAeTYBMZRTHgdbC72o7kLN1Pu9pP24GmzLKGCx3xOLM3/Q
BddRIqSG2LNPDTh35DV6LLyjkAydcOH5BnM89gmclq+4SG46dMdFuzFen4lZyN9+D6Hjvl1OQAUX
OPO9B9fhHjLiaWqO/QtHu6j4OGz9P+wlpEN0zJ10yPzkOZufj0yjumE6fUozKd91aMqkF8gVRGK8
teCFg7AZm/Z7OEFzpVZA3QOAEaYfvP/x2v5mh5xna2yoL6yqTMLhIYfzNBmg/YAq75HsM6HcvfYX
H/XJrJMT0s2J/qNP/0iOmP+ysGDIA2GVgnEdJvCnjQ7yvassfVrEgXfLqobZmS7XPtw1tK5BUXdu
RzFCauA+6KXD/0Lex/Q8ZVLT4c+pmEQHemVVizhbuADj9n2CQz5FbWmC/Ckihr8yDXteG6KNvSHR
4QCrPrCCLsr022dXyZjYUVaq8ChfxNgI3ROxO5x5ZxEwnXqywJe/oyWcULWjbvvC6SqLFz3HqEST
nDeO8IPTlzHFb1x3SN5QOo4W2jREPfhQMijInJlwceUgSHJoejP2YJt4kBB3c2Rs6l+eGSHzaAFs
xJ+gHN2qrcULviPcXed1MMZ6x1yFTQGqn/iiYtxAm9WC9zzb5c3apWdQUxFWzJ8Jd4zfQ2ds/hxf
acWzm7Dp8nVbsQZrd5GJ/Auwl03dKZVhydP5aTh5y8uJFkzrJhkvG0j573ZHEnVy0A51MHgAR1Ep
5GcaXPi9OcLh8biqhhhATmu7cieWvRPSvso7w3k9c0Je5ThztkNZS5qpQN031vGU81b307vqMcje
j+AH6wYpbAJwxs6sJhq9X5rRqAm6QwU1MySY8gBFn/Lq5rPMkazM9hh7/Hcw11i+bzEhUTpdvI2y
+w1zZhNLQ1zKI7VQEoHaTIYNxDmmqK/u7YcuE5teFtbcoPB5MY1EOMuCJtkd/VlRWaBsGx7G9u69
d3xS7CYNV6UGSZFGmPE2gHGfrmkWmBghxNtL6L+XYsxUA4LJR7wsvzQOdB2fjAw5nQFVQO5LFoUw
9WmZqAPpMGZ8FuzeleZxoLV+tyih4nW8GKCsIb1IZBv480LG/8tJ9U7yY8zoN96lmaB0lxnfr4BD
MqmDuyAHq3QWzc9ZD75VAvDrA/22zF0YXMpKKmFLY7Vz/nwunlQOHxqjrHA4iLZIQE2dlA3wPmXV
1HGLHjsCW2jk71ybRZKca+Is5B3sVkYSNa1G382nwbq3s7Wy5Xsju0QGD2vWh+A/7yFLkl2nEOB9
AwxGIDwXTKBfFq7BSIn6p6NRdPgAF4s5qfD452ZTmIPIrbN829jfARIoNEoFiNn5YNzezGZ1G9ZK
NOLDMIxNf3p+13GiAvhlahiwGQeDfC45pgVaQZifOeb4wwlpYoluPPnn4tmtgFCmeaVfYSxGGMxJ
aSHJVad2rFHOWDPrqO/HdkM/nWodF8zx1rJ8vc4Ub32t/4c69zgck5XQhkbV2lmRFGMr4IiPEyG8
79SZGbjo4tkzu7psJdWW9gY0mLR8OQeudIihRINsVg0MZhRZh1k4Rp+XTBMaXJW8xRjzTK5j5Zfm
kuwgrdVpptJpUTakMhGx8Dv1T0hG5E1IOdd4dO60yFuvX7zW05fe90Oj9+PXxB8bKlsf1d05vYT+
sUdilVGBiQctiovHUMdT7fpMDnQSg8PnCnsR/GL+bvzrJURt/DA2KrSTaIkhf/Go0q562CUARpQl
Otlya42BZt8H8V/+MqM7yw44vlT4vKFcoF5nneXkfZhjKkTnNTW70SPpzVlUCJaH3//lhPsTqVfx
F/ztcvkJzEh/2Ty9rwPXj9bNRaFFXkpu9pUXeWRTBM8/yRH64dg5xErYZeT64xKyiBURJIVczffc
jEw3lCStWC2X1epc7mjOWtmSDQFPGPIUfjGsGjovYU0MRys8ZRA6KcU4Yk8jhy77ZqQx3HxkHhWu
PGU1TN9+r0DAPTn/4zlAalGjJyiG6tHlCCaAJW4UjqPRJYBUNZbvpXj+5q6PXExTn8WdfJ7kqWbT
jf/t7npYjxtVkHyKalXhrVcJV3UzVEDklPbMXaCGzeotHVI0HMrBMY9/1bOUNjBYeJKfFT4LN7d9
JupU5Fg+ZwFMrjZtcmmBvPnOxSeoNJx+LJxaW/tF14Z7vWhT9SucM338swOJVQqkToU1Wj6KmqPk
jhwJh0i3KxxFRMIgknSODePXvpvphwfaZ7eODJbstIo3ef0YPc8RKAo/CbAR+y1OAbh+dqW+6Vsp
4ppJqFw6Pjgcy+xTpJ9dTnyPm7DHkWOhY6vfBSAjzysETqpYmxK62MQYQJDHPnvaLkEqMauE/5g8
lzmrZHPMXFU7qlrZ0O9uS2Qss3oct6o5Tw1XDO4uozdHee6i7Q5fPhEwSNvd4RjFzUS7lP3dWxvR
Rk/Carbv9/6drDx43dMEXu2tCdC5VIcZ7ZMhCM/6P9wbJVpq9WkRRohrvj/QkFgM9CvHTjrbV6s3
4qFJ+i97fpeAqT5fZuiwAH2sTfikOEtO+HQ4Ukz7Hs4U9LkWAiIjWmjldmSJLo7DBzTBcO83n8Jt
VrNrWlnmztwpCPTy9LcL7w3GjSmHbxrfTWsuRKOzhJK7oiV8as9+4c9YuUMYAw+QdYrCinWvhGJp
q6ZY8fubQcjFZAvktBeu1N3xrcypTZmrGh/8nigZp8ev4ZpConIAFFdQhnDxwnpS4LYr6pR7puiG
jdJK4XFGMYYpSj/uoruM2Xi14AtwFvbUNqvbOUxcZGnQQkQ+4ABA+ReU6CmDyFuKjbV4bF5hiuCZ
xQxB4rBrQQHDhe3EOKrD34oeVBMrGaOTat0UnjoBkK/GYt/YC/o/JRQcqgNqnQanBrZYsWGzLMCM
JSUPPdQfO7FYYrDMfg5EcKBYU4XX5qw4RQ0TvRIhThzxUuEC2/kKJvxekJoZ26RA9gbpwEM6zb86
3PbbavinpQ4zzHo5jo5r1r6YVzEOg6Rr1LWctC4Q00XkNke2Syns5q1soxKMgez9EJyKcKYLksB/
r89y0jOIS5Jy0I/ANoyygevxf+t1STjKeIHnwnBRB8iylo0g+Pg3GtLSqHNABX6CSr+PZ9YbGnr9
kYjPT8wFRASSWwaZKR2iFPjgABkxlK9p2YKrB9WOmOeMwBXeVVivbY4tRn2vKIMIjHj77uX/NQry
MNl8mdA3x402UG1oSzZmOv1hxdsBW1VMHnG3663S9I98HfpfPejvl8ARtdhCoEVPJ9O0Rgjaxe4g
9GbpDe5cv8UCEra2eLQXgHqHoYiPElLV7V3523MZllGJx0f2bMeGWbqc5hbIj3cd2m0GqdZ7zAq8
aouJlyaVpJJUA5ZUxOCqG6UItqqHnVDijFJbNeiFUdncFaCg6xZT5MUsaNZ6ngfIHTK1QI9d8ycS
2e8ELLu2K2z5tqZmTp1bDqYiPDocdEhvvCOonHsTopWznXPs3M/l7nkd6SXXi2x2/9cwvvM3Wuju
Ml6crHhZM1dX85ouvCL5x66ZJrJJlBn7DXRIspAVCk599WXE0rPUJHng5CCJMy6Bz2xg8BIW8JYL
eHrQdLwX/A6QGXKamUNUv6aP1TqSNYHb2RqYyaw7Wi43oZ2vefox2wsbZSmCmy6Y8WhZZvKunaUf
SeP5WlKujkh4/f2UXvII/hzSFW3l1hyLHPP6f34EfzBk/frBrhLcICs93ZoQhMc1CCABlVNrm4qf
NtpWueHbCOp73esXUKstkyaWbEHTo+YAnRs/fwEE1zvWAqNpDtk5zvoz323YGZWGOgrJfGAxPPHD
FkUV6zKYFM5BalYCeGlGG/DjKp+bcIx9xa/R8Y+8A74Qx3kgUg0CN4bjl0xrwd8doMcpl42e5WiJ
3kpCGwmMG5Kg9mMNPq2s7BfQ3s4/QJyQwkvf1VGK8FP3z07/s5ye9bLZFsNCOsxp0bV5zV7+8+20
/iLEJcyRhHQWkcQVMimJVP73Uwb9ObACttuvAsyjcS8+9o0BNsDwVOIILgzDA55yo1t0NQzktZ/F
NeOKlVdYR6QrAjAY2nDHA0eCiVp/IDb5p4vcTVCglCBdzsMAqzpMvZngoZRXshZ1f63AuNel7+Bu
FZangavsHrpeJp5bWYHrYbdwap6o+s9fX4ECIM2wGoGoOQr2Uqmr/XJLdSMrlQIEiGRYpFdSP0VG
kjedvXhLCNXdGO/tcCLlj2XHD86XppVxlsGgpI4577aCNaldvufgWk000Q5wlPsS3crkAGdRw5j/
a6/Od0RWg0QrXamMw+b5nwh+TqMCiAi7pMihZ0UCdOeoLnTJq5oGxx99Tnoxh6G5XlTe00mtvyjB
7to23BvRi7zXrkvNAREXC2GQa50Bxw/y5dqRInZhSyT17dNonQmFAEEFSRoguheCDSfshlsf6q93
hl8Rx/KELWdGw01gpDHvliS8oNAGC2T1NODhWw5UOjOWsTe30gL3HmO+ZVKv4wji2Qs673kZzz8X
0rcARZElWfZa6vsUtAUBpYtTsbWdhKUqkzCKf00uLBalx4YbJksk1i3fA2wyQMYt24sfNZ1gb42W
ej/+tErObySu+FDrCoLuzPKuk9AeXCy7HBqw7uzOOrWw3q9v3PygHjElC5iqOTY2qotRyrGw7Qxh
ZbPKGFW4tToJJzlByjWilikQ+UZdoQk9C02a/NP6JEFvkBvkCESY1LU9jROhnL9mKAYx/r+QJTDg
hMThHDd85Ft52iuJ/L/56rfSpHcg6FPqHC2Pq9eqdk1ZrfyCW6S+f/Gs7B0q4YxGumkpR0TN4B3I
O0nio7AUapG6ZeQV26IUJrW+ztbxrksDU2z6Vp4/Jl3p6sa9Mhs4h2khHuNAMaHf4HPAlxaT9Hvp
b1MXZraQoeMh3dM2zS9+m+BA/xJpmGJ4dJs8LWTIrCHkng1bPp6l1q0HdXfLCSnOZXmLkYl1/X0Y
cOvndBthWzauPT3LG5QE2fbhlPEyH/KeSaRoUf9rtZhjyWD6An0UDRUFx8lXte6hE5KJZOe/dz+l
7gCcuIIQ6sauHfjz4DJUpECoWDidpONrZSXFiLLHOyeclLC92p2DXREqYfPnB5mtPsu8YD/Ibw6/
OEdmrGcWneUYwu7B0AD5ohbGxa587Q4TRY7CMSMA1iIJaYq8JZzwvp6bNYx9l1eRVwl+NXjgWVMs
p9ajesROAvRRyQ8jX8ewLGE9kfhn7hMSLyHZ1KOGzrv1TEQ/N0kAgOyO1sCvZTDlCE5gBQXuy6r8
WZDwCCPKMuUG8aLbYK2Ns8NcjJkDxlcViKwKjiA2Bm0gHFYZocHZotspBKWbf0H638eFc5zllapx
ydluE4t9BgcI/SjAFv/mJZldhQWt17LbjyINrotyb5MXl1WSvukrbXQtKvUXiOmTQsO4Ph7gUEK6
xjUDrh6BUft2dewGETVDZ/9VCGehHGShUU2j5CVhl24wRZM4vDrd9r7GkogqzBfHBtk2WuLD06gw
XnzQZSw17BP/bRnY7jXSqXAHSChjuH2j3iSMCX4OJiwDdINcgbioySgMmwMAtRappN228F+oHCrE
YOxJq6UC4JgfGW2P5LWFBvvqCzUglmoAqfcDIxr6vUm/phwaoBOQwu85TbmmPV1ihhCujOPug0YK
Raa8YnADodSqGic6ivW15CRJxBnBL6Y2iTLf1OBUl0Qg2cMSKD24uZ/e3/Q/qCJbimcWtinQqqI6
Biv6O9sSnN0R6BKkT9zw2+HrA68lcGqEMgNB4Sze776/TkMyuxW13ChL3pVjz6Ad/ozqEvtH1lMy
jehnDMkzm6B28F6/1FngCfojwW0ce9pyidPySJBjS3SvJw7d39rMcb9IJTnHo6u9zozuEKS36IOS
oLFcjnDN3FmC3MQIevvuaOyTtiAWsj1dvTD47EvZGlM0rBUBuQWVH+KxWQStjmbc1OGDAaBXhkKY
JICR8hJP7S1tGuNXOKpWKssTQ7be66GPoqWipKITZoak43tC6OkO4pE3E2pzaAynpn2o0+PqJ/mc
qKMn3xYLucf+AC/qSjBi5mGOSF8P8HWN10q2Cwo4XnTBNCFlDFISJ5GDpFlqDZpCPEZkJijS/Sqi
kfYfN/m+3j16U0eXC8IVxpIqq2rZYm4SmufMaJVa3PX0j66FfnBrSc6/+fMCzZimYJI0KpyVuQ9D
uMO5H3WSkfaAnye/++rTRyRu18u/eLRNXdR+BND6pHo8ys2znScoJjnpvCNsCb04HgWs3lTmwCXu
CTQxcLlPi6ChjNFEGEgGZTRBOksMeTEgmJjpWkPzmLczB5G/9uPGReAM7iB4FY38o4OQgjHV8WLy
WIT21RihNNcSvrd9rgKhzg42lnh/TCcfAOhtrwUXaI3R5e4AFxBVzljTbph1m1oxXwg9YrhCZrUb
0C66uE3IaJraSt3R7qJ5Lj0Qo6X3nSrkA7T9HKMhK1SjQtVkOrOHivwOFF9eQcrt6q3DHodVbTDE
rP4q+sqdwU3KnrzqQm9Q7scU49p50gUvoDW/NJLeR4iyf0S9VlLFjQTCX6x9uiz4AedzudY1gFDi
vS4xyDOhYv+wQeA8LgJ0b5w+Wv9RV3rrpnVGr3UjJ6DOdam1VI9hCjsUReM0SvEhXZvrs/uBivnz
8YIvSfEIdQvnYUJOpwvGRO82drqNYJm9OeBnJ6mP3vgKXp8ZT+cKJ2BCZpK0QUNMKFdG1GiwKxZO
7Ly9ioHRDaC0PsVlm22HGdMldZyVRZ5KyBRy+yP9Lcogd2VQwRzZ5q29n0QgwDhThznMcRi01Ew9
XIAnngFiv1vCcvnEx/PWK+jhQ6ytzNMPZ4B7imwfTNWyPelufFbpah+TECMJYIrYTOY0Fkxql0ps
CJPIU1pX4s/UhHKedQ5+Wq8ChLsvOgPXHkPZlmcog9wNr4A4WGSO5qGcNcPX/b5EcL1pBbsr4A7k
2C0MxBt7dbmtu9tsH9mmKeBPyk65YhkrY/YQ3Fh6SVWeB5iHyEYl4tTXEVGugXP8N6OFZoCcXSas
xl7wuqFW6AmS/2EYUvT72xQRcYwFYnUIkyie3gVs26ijw0up7owW4OSTZlpcVOSGneDbH4fQadQq
42/A7vzFqqolcCwsulASNhZTjIJY8nJA38wgrrLMk6horq5msFGKDPE4cq0TEu+VshOoZKryy1FA
aIHUZBjUxGJHw6PZhgXZqQQxBJSE7xXTD1T+y74ddctxUslwb93ZW61YmWYoDlhMlTCBtce80wyA
+8ogqEEcj/57UdB3EBVzuza2zHbRimyHEBAX2BmsLbBmoTmlr0onp3yuEyDhPZdzpO0CPnEHkocG
REfn4JszBeH4f6W1eq/m24J7hSdr+z8Sl7ifluiVrh7u+e5qyxW/4nQJj0lI87vZxh0IU+4PUf18
+3W1kesMPLXlcmXp1ZhzPV39NS0mAHGtEEwsF0bnWB4IiPMnu8e0Uc5K3GzFf17EnGSJgyH9JNRY
K0R5QW28Fm0hOHdjVTYAltV18UK1VIhunI7xzv/m+Jn+HDCdZ1m08vXnjoPRfoi/z7Irnii3zD+J
3Guwjkcb8K0h1Ipm62i+o9Z5xtHy2UpT9/wcvIEh4VWu9SKqhEdmsrkBxOzbKDvttxZp0RuCHffU
693mB6BNje+m4uOxTCrvHzv8Bme6t3UR/OrLz2iA5wzJZmRzv0+VFLWVbR7asFDOPdOyGKCa+sJY
AFoNj2S70gHRpYMlOufy9tPnY33cq4Aroqlm+yl7OL2p8Jhcs+AHbrlmiQIknRnOLc7vCbfIlW1g
uyWkGzyFEbdf0MUYFx+mg9yHJeqRmSnQNOZ15s8veWuQWwmIKcrNNLXGdE6lgRKpfAjdGsK7rttx
1rJO0Z/kuVlqePLt/rKhTrn+uDjGCga0Jvd+1uP61h7I/SsFBzvTy/cZxz5akiLScwa/+tRmy83y
wkiEnNuGlBbf8XOB+WlXLllsPASDdEoHuNILVtOPgfg1OCp4NuAnRX8/ii+yEeyiz9fiKWsQs9Qm
ZqcU73LnJvkTx9/oiYW4CaGH9TJs7qCUCxztjyf2Cjf2lhr01v0gkWWEfblfXSkoUizjRD7Sx9XN
ZETNNNR+c0o1UvBmzntqjqWuRLHPmGKCPwINhtFQmt7g5hdWg2DsE07gBXtzrECyD6qzMO9zsGAz
lO7UtcMIMaNo9w96O3j8ytgql47Qy1MzNbMptJfJCNi6Gj3ornsCS6mEr6/MtwGAiaTTCzjI1YOZ
Gq52qV+cXxPGS6cRzo8oLjZ+2zFzA5lGR/J0C8E1z7OkHmuTCByPQqeXvmWAOJQo21SNQNmPFT2J
KmvNuiPRnorihP7mRq/dtTzKyRKahQg8ZYtC7I6r2f4yI7rvvaTYm+A5AcEMYz5pC+SViP4nBO6/
d0MH0+x0fhxjh1U+V2hqJejdsKyhBwThSkUJ/FCpXMCM1ZGgRglnbw9h6kehzuBL+Njownfb7+3i
9QxCAurXAX11fKPDnE+DcMhU7FbO838Gd8AttnWI94+j+C4Os1zxFMtNvhTC5EIP5gHbC8AOsK6t
tFSSPBRr01endupOAY51kiVuTusBdZQyFMGs//sxm8kf6Go0fz/dqPoZZv4g57HR/mCCfJo4Tk6z
qPZFSlaaNxPUwfXT+/EjHGPjMnPGMEQM4lqsASXqfJsWeh/w4Uyd1O0gExaynPNlprAaov9338QG
GS6jppMAMjnsA4LOcuq/V04xwjXvSCAAzXBQ3fpLaAhaWWbQh3JYJsg7SUojvIoVZk3tO/2nHhk6
3D/C8hgmr1BNkLMhsQ4utabL06BetZBWz/WSdvPnhtiwrA2VJzj+JDF0IVvKJcllfEaQbO2VwyIl
/nOq4ma6f6GCr5r6qALaMs08x2uQDC3pF/HYoT/9JuzIf1bswFCoImzzY9ompepTLYYqFeXOjHKi
kERLRtRTquVqDyN6y2IeFBEwSqL9stOpggXvuxBJWHRn14beWuyNkoPwFktgxgpMUd/VA7yMUBlO
VCo0DMa2BO1LoUdzmF4xYNi0jEdJDYKrZQIWEC/9zgWyN5jD1IfSWSseLCvKjk+bOINZjY0lC6gK
a6G+/iwhY2yt3njrrRfTyGj8gdn0AbhuC09gLtVIChT3G0HXNiHls6s2ZRxJ7zCjUX/AedZbe6+b
8qCJaUOLsNUABeLtoKrjL4PGQA8eXobDzAQ6qEGtURjQvXSQ962ERVv0sdxWwVBgiKpbTBIN/j0e
nZwT1G727l+36a7n3VsAlKvwOEOQ4WBJ2LA9zqR9CY1/TyJQ4e9bvD5m/ovM2Og2xnkdxeTgRiFD
hcYwb7bEWcXv1ivZVOhaQNiGFH9UOB4sUGDZrb97FkdXdbZcMyAH0WpQG49sQkIxhnZeS6MAm1oy
1T7+5k8HUHi3mvS8Fxwc5agV00JJng59hy9BHM3FB7BlzVJRZgbma3awDBZQqHI7/YE2izuAn5X7
CO1zUdj6RQwyxJTsXdBMu6ydBUW0gJmLB8jz3ewzohBWczMjO62pgubkYMlb65vZqcDxdYE64kHS
DWa2Yd9q1abjWa3J0TCs+AOreidVtyLRTqCqr9G4rRcjL2Fw17hr53Gx1SSolprZPP4qiaNt5jfm
NdwElvV/GandtWUDpm1PUDvVZDAStDMxpsHCCQDjRKk6McH1k9RGZvem6ypJcgrlJ/bpwvaUmAzL
PhYoIZ+pieJb+XROID+cLyB0sgL0kM5ETTgtw4Cjg4uGy+hTi+809EgSgpRdb98HP8lnRjeYbD4f
EodpDt1TAYSAWGvLV3meiredhSXNIdajGAo/xH9tkcG0ZnEZErTRC0aoEEkyAzLHZzmpW1w8hhyg
znjSrHa1KuVd+ZM+WgoUtlI0RJkoApDi+3RFfrBGWojR+jhmUPxj3wvwYVFO4DozTtouotlotrGO
x0U+2mAy37AAhJEqL4P4VUIsInXv9jsFcu/VTmml8JrSp6wgA4/d+vS4yPvICSI6KBwCTcZe8/Bg
GJhr09Js2mSfXqQl8xqfWu98LlEgkTqrVk9Z4PhnmRYMaZp+6/5g3QFzAYtPLcBHRW77xkwwPh6F
SfHLOtWtplIYfu9943wfKidYBvvwF9YWYSuUzq4o7FRTuYjlO2/sB46rCYa50P8fuNEdBjYGi6hM
MpybkKGEqYwmbIujv9J0TWo2ZLVSlrxYxbWMR4yLSFY91TWesc1cbEiF4MhKjqJZsdYIKn/MyOfA
cLNlAdr9Hx4UQ/1e2gN0Uq7uONyoSTy4K+4nlvG7zxQaCYsLJk8lF/rl2bcPYHJnsyd1/RLIgPsW
u2+s5Xt+Yb6gE3dbbNLUaH7xvidKMJPjx3GoBOyuq62STgGJK+V819Eb6atCuT9dc46SC2PXBQzP
mUsEzgV5pEr/RxmVP6yLdlIT0Q4ec0BLh67eouw1FVz1AOERYS6iHUQUJ+r/pWDSBGQF/PKUK1bV
a2iKgvCOeA087N1JFWpbwA8XW1IUOeCw3aTBIiX6yb19NPI7GXaEqqHj3YYEJtVUhfPic1rhmZxQ
nMMfs/5WChMWehiyZ4wNnbECv+V8qTw3fhdCIPjDfb/LXc23JRrLiemETMcjhmfi8OBEBLj3doy8
9zktgbLn4GyJRksUko4NXcWSQ4fWHNybOKnkVMCstibPTdGsA7HOfX2pMKl2DBRdGp4R0hl4OZ+G
feoUOVErgh2pVBJhSKkGwCBHYTq+I3y+baebytTEFfgGWkeeYDao1qc8bXEI8VZ6izc5T3O+1ac/
eMXGNHhLCJGsuhIxOmqBWKUHMTnSCtYLhvZ6dQmu0oHT5SYjPOvN4hob7aGFfHjNu6aX3UxB9qsz
FnM9hNT13EOZc0l1c/Za0d3gti6RiOyNwIEjTRiTPp3F3OzqfbAi8uA/zcdQYJ8FScAPpyAhqd8z
Hj9JP2W/ePsHVBgS2eeeotq76wOf7wgirBcqA50aQrXmeMvzQZ6lcqNbsbs2i3/3rMsGB3esWcDn
6Gi4sssdiRZrysVGLiPHjJGzsCLQISDiFq5T+Kb5UIFwgHknCtr7SSeWy4s7053DYhib9ot5S2Ni
pdn8VyatGVBqKmkJPVY5bTszs5TA0wJNqqQrFHpxJ9qo9VvVPrlFLVS5/EGBVfxWvCdvSppsUchU
Nnmx0FPETpv00dIcIZP1q8SR2F36nzPi6R7/Q2PzqP0RTMU1SNNeSHe5YU2N0eHNeZ5bmAt7F86G
6N/ZyGQXB2rGKRo17/OK7Aajuk7JgKE/q5s3cMY8d+r0SvAMb2TH8xn/qV+XcOgKfiXlqa4DbAS2
sL7FN19vOSsQ/BD2nnRhMG3BdNx9E04SPnq4nQKBpyioayNYbM34Od3tSIjGnCtz4kOjq/NVqKXi
EuuXRo8OritKZIYX674np+f1+hJor5OMMO/hXtPqtADkmE7Y294Iorhn0sKRS17VPoIFmLIuN+UQ
U+hUJ/UQxz4hYmuXhdW5VLvEPxpfcJMCNXl32pZ5bjsaLruAjf4ArMu1VVStV/CdZHB9skqw+b3g
b0O/Nrci3UEYBeRixYNDGSzuxLNFm02+zd1uhgA0uenWNraXFylUbo/L3iPS63f0zh5eNlUjlDn+
uUPBZCwNvG04WB+wSdg9Oz6zoPxPBARTzzXujfyoFuyXW211WUKAqr3ZPwAW979V938dN9+fMlMV
8WUXufJQniElobT4wgqaA5Baue22r9jwHVlkFw/IfryRYgW3zhZTNsM+x7iqAg/hlxrNk95DKgto
6ucjZZECaCV/yxRB4zbkfBYtvEwxBYaFcd/emOw+R6acmH1WaKxb+01ekSF0OrJabeh7Dwe5XgJn
92llgBwIOISDJGb/QNPd98djetL+LNDAl7XVVSPJ847sUfLYsZkKvmHcFgz3QLVDy4WYx2Ghe2br
mqO3NIs3NNG3d2Xun/oE05JMklciIOW6v7KQEx9ijxioi2gbEnYEtu1D4OtNQ6MmmGuJvbmPyDj2
+5nz+TwDVqbreU8rfhrkY2bKksvkxJeDZT+PZgBj/OH1rkASRJbmkx71vFFtNbsSnNE8Q1Ctd9fR
d1TiDESCY2YI+f/0PUF35NI0H+ilVjASMbzNWqk14HfIG+dh/HT3HkxSA+xHYHStKe/1pb48C3Km
99P1PQW+G3iLf1mEPVwfSk24ovkD2C2CtAKdvmlyCweupqsofeWPUK9GW7oBTervVi2m317my9it
A1LaUpw8UrVgO3O8Lzvo4nLMJ5ep44z69/+XNwLZ9/zwqU1IKZgoaRBAAEJ6PWwGKR5GvzXBLbLY
mU1je5pVSvvmemAA1fdvuCWoO0YEqvmpAihIKwRIYPpKUlA9kzyXozbUOBEjGgUasmfWY6w2U9Rt
dRS0IMPVB7XmXwzr9HZh8hhWLmcS2lFHj+w8iZaHaYzxypQmGaXYmq8ZBmpVE8z3irYj6mSPoeaP
/RV8kJHCSciG/IG5N4r5hCKMs5uThxm8eWkyoNvIEZ0p8aA3h8N1r+HTMS2DgJSNJ00fTicf01Fj
4pjFBdvV2ZTUCUqXHtT1bKsQIoGcetyvzs/HFbcfeVCoyByMWtCUZcDaoekZ3QdMA3zHsrWt55Y+
7wUoD2Ir+CzFqWvOLxaAnXqz2ohP9FsFsmZTkRGhvdy2LIHgY/F+dgurjJX+n5Selklm1TsXy0GP
gXfo978LY21HRGU9S6+2RrUZqME6ST1YHeiyja3djJR4nRuYu6peVl6yU5Dydf1KRvEdBn5qKXC3
ta/r62vw67xH6stiaiZgKuXBar5YHUtsMp6wFAtOaXblXmVgmvpc2O5+qConM6OB81FhJOm83V+V
qLgyUBuxIbIyhY2MpURUaDIomDtXlG4lM93kuRY4uo+kqj8VqOGYME3yHxhGS7BpQvfUeVualm1H
oI1/7t0uIDxv7h7WM0RHPJ6o8EURPm5jkcstzr9E9j8QKbE6BEsERPNU9sHNO1gXTlvN2rbx/LBS
JrGKA0ZlJFrEWUmdQxrST2nDEXy5C9hMVEOR/5X07BI+/CLAC/r+9DNZkb+dIlTpO6ft+c5uwQEW
9DlxCuB7DM9mTnZQmiB69PUa7FlK9fjt8fYL/6gQA1wjz2kckO2GcNnNh9iqjz6rPbNaB2HAjQpy
17m7REhPCLqc9j/h48Mch0XS0YMTP/wgotwkN8Gx3JgLyn5ncqnni+CgI01AboxdNfqW0Z/TGavh
g+tXCyUoJdx60L8PvvoFOl/zxa3e/1VnwtCwW8NQ3Y7CqZWB74gj0lA7X2B9LHmeA8QcGf28ArWU
vI/fx5wC70o/Z0qqZ8bUXw+OLK36tiHvjxqlkI90pmjYMd6f7sg6QjRBkcX4+ngr51nx1hPh1Xy2
1eFSRaDZfwkob3SaQz32DPIlgi2ZrLrFpK3lqb974byqkNf20jU/aUaQHh1ry62FjiBP9wHkyfvP
hz2yfR08yhD1AelWOIXtJD6ymAFBWpbz+O/K+BLn9S0aqhuo1aQpObm/cIruysBAGnorfImaEdoI
nRVIK9EU22YQP04pw5C6l1dUFdFmiKrNTMmDdrp4zpnW+uBhyUc8uS1AKDLpJzwqjIou25i/XIOh
r89Vzlbi1/umz3mW7QndBLED6bNkaiGcmINfRHBa5Ijf9SszW/u9pgBiSIktgSFAeEBz89plJ8s2
8PVdW6UKuM7kEElTvUPaKnzpd6jSMgtcZMNEK0OeG3eQkHLm66XZFumJ+jG+p4am5Kjc5efUS3bW
jfB6Sh4b88tz7Kd58sX+yi8Hks6xegAf8MrTeP5h2bvpwRjshsHyzUlNkaj7XNa+ccvvrxR6jLgw
sjMmMj2UhBsEPgb542PumyU9WiFh4Mrh86+9A76LKCzCn1/bfxbRFEN7cZm2OsO9HaJ6f9tO1Eyg
XP7OiqE0mNt9GcPlWkDhGp8OwzcfOE73PA3y+YpDrI4cZvBxxpZ3JMEtsk1cb8magbRMBIo8KvVf
4qcQx0ctuEd2ObOKBVF99YnBXy+lCyDWb4aLpKRx861odklOJBz82czcwk/nU7mgJJd0mCSdiRmA
PYCVT0G7AbAYIeI+3Hwe3n1f7K1MgafP0OVno9NCZyMztftu4g8cmzlRQsBfzHIybp1iLEQR9dB6
Uvg/XwxrqBnx7A85MNQ675HiMxWWmlnbTBa2IYnWoUkIqLArOfWerbgvuwMRmTOJ5kS5kb9Q0AFb
vKpJGnsomqeWEH9PGsknbQIm4HNzIZ6ib0u2UXS9ONZOvFHrlvsPeyAWMscHL9ragYGiZvhZGelr
pWndtT/7g/XBN4O8g/6ArT/7vFPtq5a+hlZpRSL1JibO+QdxxHuPuLi3zUg4U1s4RaODeDsrlNyL
ArU7kSmmUWbXe1xlneN1Km4Pkk2JvOL2+54n5XGJtjyMQQX6HXbfJEDFJ7O3HN2XVd4sp8qF+gkF
G8poXttAVK34tXCzvI8H1cTUDzG/uuQvZbGBW7WxOzA43+3D/+bNqw3Dhjl3fZ37f8j9QbHhPJc5
cc0Cp7LbRcG5ZrIcjL1t3+jlTUfrY94SVSOq9jY0IUMAVYfnZLnsEtinDOfa+ineabUSp3jXUPQH
jfj0viBZXWNqoxjAK+KbybkiXL0UJWhJ41CmaKnYoUE4bXxBIGwxqNDxJvE4qPb7jAtrp7xSAkA8
hNUu4d5d190KcT/mAps5jVfLTTa60MVccjxZnEsNhsrEdK1L5TzQM4Jx2zivJv2vOW0MWd33hlJo
KEemZDttz75hc09biFWq6Bk5rBSCJHBsJxq5vCcgb0WTGOVoreJC1uJbO3coFLCSTTHo9qkpirBf
TdeE+l/OW6lgWHB90LXT0Fs1z7CUjZwxozgFk0F98tXVjPKOrZYw/nQ9PbMsD1QdvhoNF0o+7S1K
aA/hT1bHL0uMSo+5AcIQ1t04fGk6YTbaPBZ03aoIjN+9pTBeZVRxh3eifh/zo8SFpdmDIrSY0zbl
jVJY8+afc8W/QAbxl+fMBFmymSS+oAEWB/uykwSPr3pZZ4S0XCDdBueFK1Adwx9Xnoim57Vb6U36
tuGOW+HTLFFYXNuOFrUtRdRNTj22gE7foyHKotr2WnRGDGBMfaWMNn3oiiX40x+4CRo7cgQkvCJD
9GMXNldcPUrDQENdV5qBC7YK5ZW/LgC3AO3tD8t3exwR+VeN8w61k8UCKd5tMoQfaPZ7ozYZa1mg
MXhzlojtWFFPMoGPSCo+/8xaIoVyeM/4bMW6f1M8Ho5gpn4Q8CNLmceUvfS5QMgF57qJKuc2nwSq
wDQsXoL0H5HjqOkHRWybsUfYZml3etrlEnYAmxsn+nm5MDefaVKI2Aw2GBosNkUlHoYgAlJ7K+ww
1+YDK4jBMJbwm+NWIquYqMgfGh27wnb1vWYbM6WDTkA9w6A4QrMuUqRp7VSR/+0b3/Od204RDrVJ
lxg9mHmjRQ14TY9HmwXR3Vr4t0dCyaUR3JSMobXOblJQNnoVTqk0lsGf4zu2kv8k7iWNgBoAo2O5
56k8EcMYS8GJKd/jFGjWj0zd4sXkBBI/wpnEE3x9m5RElggn4JvHalPIrgkMctyAeDWzRFGco4wq
DR4Gf8dVWDogvB7Q23xOaRu1rDb/eegZ8XumUO7YCu+QpmYzaEd9UgjsI0iWV1DsBnJ9nhCjM7hz
PMQri46VNrBBeej2Kh6b/lKRD0H8e+6Xn2+w8E1//jyvoOOYzeehwWd6Kxbx0pEA2LOsjLkMY+vS
Ihr9VjcFTv1BS0vmtSgoCEEyiWCtBx9PHvKncsMkpwR5CpT6jj0H47x5YiNVoD9FOtDjQN1ut4BH
cCWOwDrQsm9GL4KYbtUSYesiX2KWbF9MFPd2Gnw7nZOqjT/+Sfbq6kGoczI9G18xH03FtlJAH625
i3GDTwNUDesi5ArPBTCqo0FFD1a2bvUxgLBZiYIzLFR09AZgJRTLX0R2pp8pqhbspx//l/rGI4c2
PeiXWJWr5RKirYF5uNrg9UquLNrjSOUMXpvJ6sewAub0xckId5wP1m5QYRw5E6aVgeih8O+zp/Cb
+2Vxnt2DaJU8mIdcKAfKWb/ufvKbom3/uY+IWF/oobCF3M7VVZzuJ0ofDjx7A5HdneF7tjSqk1x8
O1bfDjB15NedHPC5aDbjTvqNcrYJIw4uHb0pP/mtewnYoZbzs2dmS50/fbY7Yt1H61SJCdWX1Dgj
pY8NlvwcrN1kE/PDn976wJVTd7roIAmFM8M/sIfbSo0m8bLmHz+dBHURMVz2PkgU1XDIR12QVarZ
7NyNUwkXzKrexI3wLaFfHVAH4yp1TObMjKiFge6ifjSAvSGmyGrTsgaWMTiCDo3PP4g4PQ1hEhcR
FSX9/YCQxY9YmFqqoXrWjSnnG0ddfUsl91JwO1zveJXFW4w4nSMU0yLIrJubkVHS55U3F/BXz1m2
HbbN1fL/um6GTib+75i6AuYMzgjpOTm3mtAXtSMC2c+7dKQLlRzNHQFkCRtfgvEF/mSy1I+hj5Yc
/6SUiervKEFf//STeZr5yHxJK1UUy2AnqQBL3Xdo+QcwI6v5GTY7nnOf99xFsRaXMcct+1I+/6yO
L9k9hv1Ts/yfwMJm3o0ikmdvC7/VwIifdDJE3z+497AtZAYut6D1zhfRpc1mJ5NwCKVGDOAq0/0A
IXj2qMe3uY2GHk09h9o/nJRMiZbqh8T9YV2iinta0c0QO2hlulg1zyRU9RKLivALlsjbI9nvT6ri
/l+jOEZKJK3s88LEyeQtXP6YogQqws+POZp4ktbV1FpQ39en+TLNfvDRzUEeoEoLLSnGUJpHwEOY
zLcunt8QCtTn3kbj5YUyOIrx1Wul03brz7omEQVmsaa9cVxPr/K2rT2orVn4aYnkvum1rEUGDggO
YC0TVPtVCzfjZGf+JyKKAiFX4MrGMlrvrSpkAoWOkGTY8fuifnxpSmP67ppcmn6nngYaTp5zNaN/
DvB+5KY3bt84eunoNnrKzshHGd21NjK1dAKC7ElYUSaLrTerYJtu82zUy/FnODQ8NMQ1H1k78QnB
2zbYo5AOxCegAflWfp0SbiAryQSVbIXUoJE3HXnxYdDVIc5Wu19BX27L26GqDLiYSUe4HYo/sysc
3ZH1yuVzCcFwQTt0yp0UmYM1sEaKkA+QHSWEuJdQNYDbyi+DjmYviAfWLqnP1HI7lY0stXNXAr3Q
8L6V1Jxu1GxJteXBOpvN9GUCGP5u/q4jhDVjZyC/ygI4Ucfyl17v5ZHir0bdxNnkm6eXgiai0zoc
Xn9m4A5QrjqovbrraQ86PmfhSxgZikwtW0l7rX1CN8hMUyuKbKC9bPfy0bkuJztsf0i6h8FYC0vn
I0VIlruuUw8dcCpuMZ27eyP9wkpqTLi9QAHykn16vWdObMUfs+BOWBRsO23SSzI8sGdFtntMY6AW
vrInbNwEpV72vvsEX+b2/oKdRyuDprUA3TqsVuv2f0/vrvXcfFdi/FCwQ/1Y+vBRcJZskp+pL4IU
wa0CZJi0FDItbv6TZd6ClFWzEf7MYQ+vIDDIlatkcQ5l9DeTh96kLOZnnHSPLjhJ2OLm4V9F4agh
gZG082A84/RJU8uqYy5t9uigFCblPgE5N0oAIGLC3ccPkJwWaarzxMkqRtTkk5iycGVrAFwNDiPS
7cexwMHgnj6DeFLcMuuj2IyDr4mybc+JHG3OyOoszfqGNu9MvX805OT06JrSK340G3l76Ta5FTfl
MK9is5beSoIg7ZrcZzgJjs33hHZXjxxOba1ve7hItgFskhLOyfY5Q/S1yiIPgTXYxGgEGLp6uqWZ
8/JL/U4x2s9Rd59JTeBdlq5hbKq/+HUsL42prdlfuS3qqpgk7gBEWiaF1p+KvtQcqfw4yZHBYsbS
aFE7iT3AgOwRlYhqa+wIa2qZvuafnPwBPknhlUvdtEcyRhD2tM4btU6rlXWv99Xa/czIJaHELfJ2
97jysq6zTVWrfaVBSr4gPLqjMUzqsEIskRVntghQn0zZTPorRAn3KfzWUM6FzoL5cLl3Tk9Gr9ew
4W8XOCY7VxridHvD+j++31ithyKXIltA6UszegTXhVV92CMTVOcxUjf2BAULQ3XUPwea1t3H/cZg
lMFAjXjoNz9hUPjavwsqJVx45mLEF7ScjmkeA4Ac6UKYZ2DWmBQdmZnFWleWZMkDCjrnQAsjGFoO
iHW5FSKhcvLG9kA44ULcxwP0+eac2KhhkNVM/ekmzIWZHaK5IqXOSv/B9bZWAx6C+wvNGulE/7CH
GkQ24KfueW0Gl/AQeI3fJWlXdfF+hwKa2AbafPVpqMoLa97YRqzCREnYA5Ac7wBErdgZ1/ZRyQ2i
EHKbyqwWG3NoUMLL1SdcYcZPUS6VlnHqkEmfX2LT1QfelozpkQ5/HHjCPdx244/8pXAEho1RPOjU
d+Ly4VN2swXHK9IswfmCM7QtuvoWpKs3ysSKWKdUjc2ERptiZj3BH7/4iSqAgIPUEJWKNf5MjbWa
EcPjlpzIHtUqeJ3wjrufRa1K+r5WT0ICtLqHq1PKEKiL4g4JlPNNXNPWt8H+taviVo1Mlg+qRy16
otcgSdLPPUB/ijWBbwRRdXpB8XkMiMdk2zUwIzAwTBJ6lZ9VQ/gPobJdO0AJC9QFd1Th8l7uV2li
lzNf2ay5ZywCbp2TP4uzbUX5xVyJJKxRjL3HnvMty5FV9PFsvJMT0gQIdVDiF0aMsF0nGrkrZE2P
GXC1UuG09g8XAMAHciKYoS34H9TbDG12d27qf+pG2yTjh/psTY8GfDL00ovi04sAoZaNoI+em9+s
IfXx+aWOimFDTRrWFaVm2acul7721IQSVrwwj8aUW+q1vjVkiZjFBRGBKO2G6r/ecqPnLfCgKkgG
gnwClqX6U4rta3aDktk1EHV4Lcaoh34NbK2A0BMda2x6pmxYuXKpZLWbPgjIPiQZ1yI8c8EZz2cP
Mrix2RW+Y4tkqaryfMpVGURkAGESxH6P7g2IWvIcZrT5IZBtUTOp5oLmBO3L1/Bx9xtv5y6REgGp
uxuhsgyS4YfyR/zPoKfPvK2jajhJBhumNVeK2kWf9JHiGDLIPmwEft0zOTo+kn5/DYWjqCCr36h2
M49vI0ihuPdden6psNoQzkZy/RM7r4SMw3CzumoHDdOLY64zXtxAqYtFtQjUTeF+fTVaYZtaDFku
j0IxqWcT4h29S+Imepk6PH2bUGAExuOMAq4MZ9+1IT098KHutjcotEi6yuFQWCsd2m/RGU5IMq0h
hu5z9sbhYmw4MFzPJ8/yNJ1iWJS2OGFZfF5OjCJs4O/pk7H7qU2NqD1xj/7/U56r2bx/zEfd7wNm
DXOXvuN/JEdlPc/MPnwI7JacpRSEMckZPiCEAgASHCxQZHPgDIkm0soUh/7F8bOq51lJRZWOl+QM
4muFkkeEtV7RFs4Us9fD1r6Rnmw0MKkHa241e7YVjGcegKAOF5HeWAsRCqsLkBX9GjBuA8m45OWV
1R/A7RLJLQDeXke5nNq62xnt00K94Mrm1lhflc/I0c7Aph/q6MxnGxaVNu7MPLoX4aDQHcBbRfxJ
FX5xmPBt3hVXmkSSkNg6G3boEt0Hfjsd9nbKWPqXhwgShDF8mEJ4tj/iTtwmel1fElmlaV/MH7TX
rnxH59vX+dLDabFcn1EDLiwd15SExbdWKUDz5KdDCLkSxaFQZZz/uwLiGOL+cFW3uSgqQB0yE6U/
JSEq6W0PL/JmxD4x7CrSDw1wri+PPIN886z2giHmjxtKVfJsplRa5ZMiQwTiNuxwbz6uZ4bfIjph
lRo6pdZZCi0PUPHwaor0n23HpGVc9nMZDe0ptBVyBV/ZBuOxz/jKMa2iW4doyqgpfqXbP7ppYTsU
K/7hsNOhNcNhRl1psWJCS63jd/4YLf333YKhrIxXUcevhVXvTcE8BlO2U8Ay1OMVuJn1Dgfp50/m
r9q7yU/PIHos9+xHSBX/aKmJFXdqRPRoGjvd4MoZpQsUtzem1NMGfOuCkGsxSR/Kh9jZZWrxp56e
h3Eulq+5BKFwp7d9U0jmFOJQTuNs5nEfL+9/+KjfnkqmF6xvTr3zlZS/BfX68T/Cfqhl159hsSsF
/SY3YzM4sgKAZ6wExIYK1NHpMzSFl39bbocVblt498W0nvDM14/ecrQDAXN9p1fttCy4XDOGuboi
BgGPLwRiUH7rML9DsdO0t4dW5sof/6zyI9iZUcvaAX7fQVMkSjmecEcm0TD9Ff9eWwoNrA5t9GDx
5vypPUk140zMbZCtT+EeogExoa/YIlaPDodEpbnBtiDPR002fID98iUonjVguJk6OkP6BdgVEXRL
UgOMYxWhJFbRiJDYmU1Lxjo2knPm8Q78dSh+R1eFHk9HB4D8A/GJnSlYBh2/VfryrJcupBU46Q93
EOvTvqXm2tb/jBAtcsr9u7bhf0sA36Al8MCcoGsYG/VWnOYJWTL4P4svR1xwgVppy6hSs8ZibKEh
SxD6GlCZz180xkzgMpmJRl36JxwtymKXEjqcRpVEMOIIA3qbeY5oIA660E/zxIh3WnQFZVXGw/me
ObU3gyD8x4XfAxR+dXLCtZ+LgScFkA/ow+XpoA7LFbTCoslLlhBp6R+6cJZ4ylOtYfg2hbBFNcwb
1s21VFaMtzbcp2TBBpATdDU5VPKO9Kp3S6NhQ+QQTeaPB8oFZi6HS5G/wni0cfo/LgbKnTm2KSKR
eszBpcokKvU6zbE5B9uO1TMuJRHVt/b3lmEeRZaDLVZgvSBg/aaKKoV4fr61Pvri40twdltSMECb
xk3slmfn/aEIu3TOssTnV67uhXOu9yK57flhHd3vux1hvJw9runTif9lnhIbmbLvC3WAP/rArKrW
9Xa2LkYfsQLwi0foh3I5k50ijbIktYK7sWzGukqNexiRKKoGqItKMMqwRWEshSWs8CbNJUluaJiO
polRTqj07zWoTqnmEwQSwdvjPBABUsD0/SpKvoA7aOFHhBsMqYdBxworkbbwpGEmJd6XDwUs19gY
wM1CnNU58s7DIEsUf8e9zkSN9Ju7ng0mtdbWRfRS3g1nY4XLU8uU6TvTFgZzJ5NccRG43t4eYWDQ
ks5Nu+QrCEMGT40i+7BZ3+PR4ByEzQAq1PoW81Mwpfps8Z+5vgFrwIJ965lVujQJLHHai0Gc8YlK
NInndrny9X39aCb5cSMvm4lVqXml77sNF8JKvf2cFy5WxdVvvm0xJ4zK9I8VtzXkaSCcK9o+4t4h
SiN0CQlEaggbt8S8Dk2i6toCfgy8+iMbAKL8G3TPPIBXap7wn3gzajyAkX4CQT63xdyPHkKxOpGA
Xtm1/tcf9u7sbr52AM5Xk/4MOs7GSsFgg+MusYCU7CI4Bo/ZthYL5EdEKQKFJElC/ZZpfR4aBZuy
IVe6WGQcTWX6QUO8sHbSW0hnMjptJ/6WQpiknkLEOkxD1eR1WguahiiIxOHyBeNepOFFzVUeynfC
9AYyCfWJzovgu5tSsavHkqEyMLsQrUgrfSNoFM//c0uKSibAm3ys2rAx8o6yk4U6eeefPHzGSC4j
PZSD10VGsgJyNF91Sbw8PLgmVjNPB3JzF9tjK7cWUz+IPTf94eixATwHb2+/bKLWIl0fnDtmkKfc
TwRh1AypfC27Nn/+FFtH/NalGNeyxT570nEUPjx5hv1ZmvJAgykWcp3wwtqdTCAXwCEh+ku+50N5
th4OTsoue/EjGrXLzw8Auroo7i+r3+YZ/A8NKaip3govq8eXsCCIRKypqj4FQVoApHkv4C1JOivw
WZHeBpOCR26Tzj3aOHWKbSFP+VJ3vMG5QoGMaI9oVd6dCT6lFzmmCuW1Zj8BvqJo/mtuPwSmzS85
wYK2Nv4QrQKJh5QoaNs+mnTxsJ07+V/QMst4JoVcS5FdaLJQgx6PNqeMFyDCkKepKSQp9FGp49fd
BjcT1L9WP0IUDi/5SiqT5OdhGTUU7D1wMlRX0ZDe5jzDSVdNUJvy0C4vtHydK9nEpfFdyS0BGKln
h2LwKFG/E4/1AKDXq9P8ILcdaZZaWftYd+vm8ECdUs2mCfYTnNUwfqWfn6NisPEvFLXckCmY9riR
TkNoacBQYWjizKkiBro304DQmcgq/MhNiD/ArravjSpJXLocHSPqIdRWp/3BZKiEEIUK2K1d6rtr
23w2GYutxR2xGa6+gsYq56SK4NyfMnwTNOQw8ObnZDGO78H0XyumLrPY+QUsGfzNk0seEDMgiYg/
ZYXlZOcZLvf4pYq07b4HjKVmOBKbXznRIWyjKd4Gi+LQVRyTENGtB5fdFcmJbYSQFL22FG+64cF/
bdoSgJ9CuiADXV7+J+oMsok35DXVaCSHeUiRQ8fRILs2w/rFMX1YjDy/H/IBib6Wb7HV0iQGApaz
enIN1Skh+2k6T/s59vb8OdKpTPxhW6Gox6ccMrIqn//smb0oBy6runBDhHF1OFZPGX1qEMTR1Fnf
TOuT/7/zKvSAMFaMiYmDb+Z7ZGqzwEobu6U+46/Em63WgZ8bwGusn4CO0j0Zp7RUfEphTTJT5LVf
NlnO29hoFpL1k/MYvQlgRxQUhp/OtHCY+IZ1kLaZ4JRkAwhEw8e70ksTyaNaNDD5KmbIeXSBqvjK
eSQ9PlbUVbl0ORdlw3rd/Rg1gAyfUZU2GRXLe6Hn30+f5VfayOlUD0TX2rjlbRY/xhHHTmmaSQTW
tntVgBXGtsj0tcGxJ09Ih0qacb1izU5Yjl/lbIm5lMZlUJVg8dtJ3YFvO66ju9ezFglo2/TQpUrd
eLMVKptzLusjzLs44StrRpUjw1tDozomvGgrqrSimo+rQajGmatMJqYKfl4AZ8Ude4QJ2FUhyURg
d7X2rcMzLfoUWMioYjpBU0kWbe7cTzeuU4PwUMcfzD12YcG3RHizPnZZcpl2hLNYjngdsNTyqa7E
Mxbqi+mlnKJwuKDKyM42294UFEWHkdNuiPEqATNHwe4fYDMNrGZ8WsE2EZV67eruNOC2ZAoM6+Zn
yctD0BfO5x/y5tqYXBnSs7+dy9P+Et0dTpsSNP8KEsHJQTbgGLyG9/3CbrbWXDHfpqSyxVkybkOi
p1ipnrrisw98R4P6CGsCKWccswzBdj7Z0PCnNOHcfwm9EnlMttBA80F+RVPykYDw0mZDT3v0MRNp
8K3t0SLTGO+gCukpVVAqPcZaF9UOeTsmj6YLARUkLeq+q4TetpSQ8McByHmz+mOr/cszo3irqnj4
sxw8cZ5ji0aaSaoH1gku/iDuSgZVNu2ugJeFpEuhuod05KuQjrlpD7AS5CJT7IWCMz3wnIUX3Z/O
JeMB7Ojy+vGDTSPeKhdCJjf1x304Tf1yPvKXX24DkEAlQPOP8zy5vle6wT8QU6yzE8+kZ3BT3iKz
N85jLWOS9ud9tQsbKqu8F/SgAqOSCvlo5VagRQMEBExZ3kOLgBuUi9SrZU5fNbJGIIlLVzONeXlt
UUCQd+bonJyO2D9DCQizKQauHUjuDO7tv0FHt2XEA23aoSpal1/fzVBobLoQTQCzoXTA9FZnGcxM
H1IXeHOiX6Qa5TfdAp//HPCUJeDcyswMYMwz4y6xYgEexSLMNwhWgng0ZnbvaqitfIu4EePV1QLD
QiKGaEiAAREhCwT0nemSDDNTAZU0yAAH3JjJ7k9vbPisWo13uTEGG3095/lC/HisKgO/9K8dyzhM
4WaspdT1fXU9YFuoMUA2m6P7tTLwzJFJpiugL2E5CJnGTc1l7LDTp4MC2cw7IpvLaR/7zLk5tZMQ
5Iy94jZ0UoC2a7sT2kV0fULSlgl7nXM1TaOLdvRt5ZMIzGGQ0kMm9lVEWhWtiY0lRNhnsKXhbic6
L5E/SeLoay+HihbrzkmPzVk90awMYYdqT+m5voDlZ/umDWTBdo7ePBQ6iztDig86yepYwo5Ekbvk
Me9dyTNxi3JgfpCr6z+t4T050R4CUxJ/YiydaA4BvyqEsrrmtx1WKhysCcXDyB3dewmfdJ3Ng9O9
C6uTdhtSRCI7SvO2WSpOfkcmva+ZtOImZgvkwNSp2S33bLIaFX3VLgRVrB9u1NfwKN/12W6/tqkT
Fc/2FY66uNP9pKGjjfFc2nnRX9y+NYuxX/ZhQiobTWzyeh5Jz1X04hMpD8nqCsPBClJpvdLrxZv2
fP+2nmgRBISnwUKQ23ngxxqq7hHvblXCLouCPRCfy/Whd/+MDaLeoUx+TBUia84YIsktw+/y2BTK
h3OxT2Aa5xpQ9fmmZuRPRTOg4N93ujmn7Por6t73szRcRF1GD+NRtIoHCYoLHbxzuqF4/byqNbCi
9/IOwiHalfyIte5fs6Ism3Wcx4I58GuK1X22zhH9h01g4nr7NmsLRRPAFiuwkOZPE1quebMiMpi9
KwoBJVz/6Qu8ZMHAGgl3nRLfIWKXeEgnzi1W/mLPTut6i0IzfS4y8zGt6NAty2KWKwa9OMxEEhls
BbCPiNFeRaVQOMEGmu3irYyx3swHWVPlQC7lXNf+dxFIvnfJlJj6SySzNmrDWoikVHpHs9+7cfxL
+FsUKd16NFF1xvpJbBMGnSd3X+0fFVLuvxWWygGh+AyudorctDPdyMlclFtA3gd/SZ2KO+xW0BZx
3DMUGfYrD8Och+yXYeGKoWK7aaSgWayudJ49e7D7u2vjr3JRR0CVjuet9Tz0gtTS/FhIZdq85yxQ
abgSQDE0pqutLVSPNLmCzPjbpPkIfO5FMpfSuEBeBk9cypH+NHhCChzClKvVa2/mEo5TWm/Knekq
zu/fcmKbdM/AqX5L4M4MEOjZlwMZXBwqvh43MTI00sC6vSttCL5Id+GZE57XnxXCNO/McuGdV4UE
POJUIbNCJ9rl0MVhrerBHnJKAjo53BgruA/k6VwFNuXCdxV4VWhg8XX4Na5qz+mHJFiUq68vnmq7
cDhgS+BcOtDzWJIjH61m+CZIOVnyGi8zJ4hL8dtbJ5GO7NcMzXLZF0mdwHVm3qNOLLWx/19EHpvg
RhluTewrl+7h3HRrPXiYOVSZ/4H5fjnkfinu2nf8ZX2Uai8p1drS7esumUbwIJUDA1+uSqSQq44/
SQ/xT1tpXuzGiaRcVRWlVYoHY8FVH/mznItDoW64hDzCbyfDKOeBDLzjEWBnWrUM/DBLWQaMm+Gm
cqm262fCcTq8fj9Hlz6yiIIGw69lGpicEiWhAunftLdEX2CtHo1zjA/JGf3gCcB6pE/AL2tBIpZ1
xQkG8vVHt8mEa8+k9pval4T7EcZ1FSYGIR84C8HNt3Pav/pSTi4i4vrXSkMY9UCQZizyRg3t9fXB
8H2iu1bSj+Juw7/OxvWQf5+ywHHTpO2xlWi9R005SN1JyWFMpObBz32rztO0QhPfAYm4C9fxM1CB
UFsi+7Shbvjlbi1RViSa5vM6FIGxN/DwflhpWoXdW5FFOibPA28VnShtGap4zzpg2YaO+XTkVoyV
1mYdKDeLNNZKYqd2fJ5IlPiEyPdSnfSFR8ABZuRkI+7tqZT2PHtV6RbubeKtdChOdFLRmbhiTeNI
b/B0QRJ0x2A1NBri/Q7w0YIXE+OnxhIoFRT9KYJYUedkoze05hqUrO+XIdk6l/GZmfT7qMQaLVl7
I4A8YWe6RfmiEJejDqVFcyDU8175pYGdV+AcLD/8uOPuNtTwr/R4Y/QR8MGtqPZ/B1ipUyFEe9Fm
j9FCIziV/nAUlqxwozElFDhTY01L6/SZMOzFluRPa+ttVkc6KI5Gm8poqhvKoSfD/GmFDQfgIYTN
ALqlPLKZ0WM3pGbB6vIQxCfXWtnqJbCfQqnxs+87IC2+cEYpakIY+T2sV9lr0Xu54AqXqPkWHtTF
OqaZeAUWw6NzvcMRsb3c/IYVccrLExg97zINOVgxl6x/8UBx+/0KoMY7PetQ4usDcWWQePo+vkuf
Jbtgtyv4S7+6iQzmOaQJTOR9GGR1Sd101Fm1uvVG9sCmKsTiS9ZsQhHYvgz4jG7JTlvqgdSpDZv0
/F/2jR5BoGOdmgVb8bPL/hYPHSUEMfZJkotzkOtzIqLmQ3D4ugWReWa5Xfo/D6ld9AzbVn5XTG8t
HYbArY/bJuJ+EaGXBsY/t9MaV7IP0DoqQW2wkfcYYSdkzq8+bVXoJB9ab8oZWSH4xNCZoSizEieX
RR+4p0gn55kc58niYFAdCyGlyxoJjz61+v1B42emh7nfsw5T6169/Uv/E0gnXYnX1ujFILHqRytU
+zxzvZ8uYxWd6D3Wr7fJ+twYbDPWSQlG12mZhbwm8wKfAVxtC41R8EGrJOe1QS+vzdNNBXkuNGD5
BjuSZMyhWg2BSOioSR79mwC1QGcchHIB7k5XT/PkDWEErdZAzLuQlhf5XLoBJkKxL7cXIFCfE5Az
f2v1fC1C6qaXN6eDSXVamjWFxt5jftGejpzsYFCfwJcfNWiIV5np65o9z2pzeOKOA/yDd3zxzEsu
fAstXpFdCGVQaJYhGjLwh6uKNSLU0vwwYfro2Y5ZNsskejTvd/H+Hs3S8n0n+D3OmJXGUdH/puVk
XY0DYBZDzXBQl9TW7hMeXk75qT5rXuXbkn5Xan1Z4QEgXfmwhDXjExpxZJ0Tsj1KuaV49/GmdhfM
wrdsy83HUhZ5MG/ghgM1CPF0fDFDjcssq801j37xsFlSlZb81WqAaP0/zxNvx4+OQimRRkT9/en/
HUzC3h5rPSgW3IPztjyMTEdaSTks6aoDvXwOosxTVVnl2gjTPxuVXj2QCv/DDKgr+krbi0wO4XTa
5wx04vEteBW3jRYEM1hDdjTnUta2P9aIk68TYP1aYopYLUKq3JIEUbJnSK0DdLMcyFyoHnMnUHLD
7HWSqBGOcKestz4upkjzjRxqPU3rMqVZL6QNZzdZWCMIGFR7eHwukHixsiL2rDxWvjvtP6Lz0g7C
0lPVw4RNlpsUlDCnaT9WkUTdazUV9vKse19h7/+KVVKy299HwXf528iLNepcpeFY6p9OBjpJLsih
1+TNpHeCGi1g5KJCcxwSvYFSTdSFafYjLVEYcKuIuedBQin6+kj2L2U844KXjF+7mOmdwRGxKqmk
Izx0fK/oagOjh7uU1W2UtWs11oLVeCMK714LzhAAypN88oq9abVaXGfxqYVKa/xNL5HHio+UVFTN
i87FzFjQfTnZzVbjykaiBN2/WUKmW0+tkuX66CAHuvDLHedK0T+yo+2nkQnyrjPmOjE++qiskVjv
2qgL9rkPZnxYGzp6csnK1ojhBMop/+3BxGjxQ3PLAZ1AltxRnJE2tIu5eg6zzwGmRSKURO6DGsaW
3voE0Hd1kZnfolAiNwp3q46ZE+SkZsjTeYNS8ji5J4fc7cBSTauNcp0J8L0r0/8OhuWGU71TLqDU
jd9NLzk0rptETuhrLFVUpiKHDmBIO4Q0SZtbj6NKpbBak/uhLyw6y2QVA4tF1Z5w+3K4gBD/UgPM
E/EOyjC8v8k6QUEIP37Lnc4Oe6EDlXhuQKH4XYGreRm9ZLiHlYCHttSsF5mQ6OwGKTbpLKDFp0Er
RvfsIMCTmKjfzuIV00tQwbkmOMVAPngKZYOGI7x29habSXUGpeN+YUSvgueBazIeYBeIy1yofXKL
wFpRy4Mp6oowqX94XuL5a117Y10UpKf4dSUYpyp/a21jb6clNl+di5/VDJ4F7CArmQP+d0K66KOb
uV3lIYUoEPc09xBy6QCpA82jpQn4B6wVea2A/o+e862s9xQ7nNFaWZY9bWE5tEFhJc+LNREPmWIf
thwck/5lulf9Ro4w8z42rNsCxeegrOdwySaCStxkffayDphAh2w6Diz8NnkZje9UNDQvLz99J3hK
kVrs1vmbNG6BmmLC87bdFifaRpsR7srnVwYWYmavKSFwrSeafO7eLI28K4ol42DI5cTPT3IbBFi2
gf7gkkAvDLxsxAf+Gh91egdYNwnGxryFNkycu3ZzFtLmvxF2SVP/S8imwFo2MVrVFHUt15Hoqe5e
MQOdjUd3hPY0w+b3hkWaZIOzy5eUKzuqZ+ShYILZ0zcO/2BnEUBW0PNuDFd7KCKTCU00GTfT8/z5
P1XvPz8zLdKWv3e+1E+LS4qmyn4+1KTl/eUUD9NZHa5q1/AD3UFMvZEhRC+/rwFsLHmfV7kfgBtE
sxGGlaTnfcnNNHh1UYd9rqAnRFGhaFHLCRAqFR+vTfWdqS58jb4lG6gpNYbJx90riKjeSGO8j2sz
Ig6Z+R/6BY5u5UbC3ZEH+EHCebQBbVRkrUuRpj0G+/96ZoSKyKPZnsmT9wlz5C70eHqBos0f0wQh
Hkt+Wb+82q4bNEW/+KbQ7/jhSPpXODI3NL8qc5bAbNT9r4wXzeem2oeZkBBXg/XI1vkuGqKX8bfj
m24qJB1fldDskFANYpmEYzijboY35/bSMd1s2RKVKS83vqQGmpXw2tm4JVy3jSXf2uoydVoic50d
1Jqc+kNd23lq+uuB4WwirquKxeykLX/QFEKe8FZ8t2C/TPkv405OfOIlJoXhbQz/vNQGSYUW/dA4
Tdx3UsTGQF4Ace3BeO0HcciWLMUZfoaQAuGVvtPzoiVqwHqV+UcyzAiQzynupxRTCp6enH9OxjOm
TYKMDhiQUxgA8yLJXXrGfrcMvMN+uMBZ9lxntH3f3OrwrQ9tvWwTqhcyEKfiorTCbF561R4k/q54
fUDdabLX58a/IQ1LE6STqniLf5a7C7iy8UigBhnvNfcagzLQS9xD7wzeIs/hNFaj86tueP4DvHuN
wBqhNsUu9cGBsRI9Y2QOFoLxIAT57tfoUQ8V1cgX7fZJmI5vQ/EO5mUKXuAbhNmB1TaiD1ktX6i4
kd0RnPXMllRN2VsHtGBEmcKPe9NHqgxNevW/rDfpJI0Y1HlxDLtXzMwrnATEiU+WrSDkXQB8fctB
V3eM/OdmdqtLWmB4g6RNtQHc4lwC8ZRzDOEiJ0yVmlcdYj5Zx0gWuqeTeJ6jeYOhYjciYOmabkbE
7dirCTk5lVIOAgBTT5cKL7UuKZQk4UFcTwbDFKA3KcFBe7kX9c5nmIZ+RHwKwouovBZoSutwaH5K
K+n1JkKZO96/Cjld6+AGDdcCWlCMYnJr4OuFeaE7409HujYHQcyctKY6JF8BFOTDEjpO7BYNlujo
+TuipwkCbTgeB3Yb/B5ecOkhwmuPnRalxXApGgd1bwqlftZHtdv9ugK+rhwwyx7AuY2Dj7soCsb9
43WQScHp50QqBUbT9AqFXZ+kOPlEuhoJ20F7WXDewDgqZdjLJVx8faY0YOTnL2LrqdbBU9MbDu/L
IFsh9MU77rpIt+1YqAZYmctVFNDDMod/9O/ieUwVvuanVssgV6GnIiOeicRew83q3At1F6irF4bo
FUfDr+HfMB/Jg+bwvzXsWKdBGraMwsMKOxXsH/Id3lLDv9TrEBdsyK51o2I/yZy7Pz7RdUkK3OK/
l6QgtuhSnxjnqJ5WwNs55lRmQyLshYOXjvy4KDgtz/9vdDZyabzZhPfYhV0Iy2GIojZ62I0Z32v/
Lb/xI9LYXJd3yokdx05mvf90jdon60HU/4serG6HmveI0IXvSDEMIZy0p6oz3cYHZ6xRVLpwioKD
ivpiF8vqh0l2GKP//o2u9wJ7Dgl79DVoFlY/ALxdg4wtHoR0E/z5epoHxAfx3srZBlZxwjEeVXzU
W2+lI/grDaW+frUVTWLRZGVVio1ZFwAjo02uP9Xns3VQRG4FbZD99SgeYR/n27hE5CJAnUXYVKEZ
m7Aqkvm0/GCliEqpGd0hl/8ps92v1nQWLxF4o6LUFA69WUA0aUI8umtOa1Krn6qp8u42wRzsLGms
+RtNy98biM4ScQlNz4uqZ9tkk+H+m4TC72nnPmyncanDMG23N+MPipFlcel3ZgXSkOAwoW/1Qkjr
tY+owLk9S9h1lMevZPC1JxFqHT5KZ2Cj03lDA/m280vJc+MPvtK7CSzgPRDyGeo+LHVGDtf4zl7n
U4kuvbSDng+BN5vo7Ef+qHS4S1ANOUZOYnSgHvW4MoKIMjc2M41khnnBjI1u/TjKPhrTb2Gngd3q
JsgbuHmDRmM1uWHDs+G9RSy4nAZEgBtmHrcPncbb+BfLUPnRelqfNANo7vQZiqEd30ZYJ26AZL3V
aF3QwqefB7JSiIOs1jkakDahnucvx1M0NP+kR/z7bRalhtfow7qWE6+b3k5wB52XO2khT2Y9aySd
re9/YhKaMVNJfVfjtZjMX8nCedvwVvuknNWy2xQQQ9M1TDsax720trtpfpPM9JLPLaqjn3v5ZXp5
8gyfdbVJWoS9Eee5oz++//afM4dppeYPkWzJtrzqSCRWxlOpcu7+NsfzgENKYI8wjTr5xgflUV58
3+axYJWC2HFSgATHF0tGhKCNY5OkU7wUVwdA6USHRF00FdHmzosXJj9iKphM95RLWgKdRLWEjYso
IGICuWYkq3F5mf2rQyd/ZxRyBz2y0oFILwa1MSAIzQRgYABpLbAskWPf9/bLOYQdgsLDcs0GyG6X
XnfHLEkIWtsg5Kgcrgm6tgB8GAxpffNbr+pNsd9a4Up6eM7AJwGdWqLw7J1ioXal0dHnTO3FdFds
uh9Mq9x6eO9pL4Db2mw9Bz8/cFap1tYISasQ/I2U9Wvb6iZAlety03oDsHw4qSslzXUdjUhQqEcj
xZ0GFBu+MpyW0as1mJP690Iu5tlVoBT1gNzAAv90ncebhNZqFuM9teBB3h0kNBdnWJnQOj5jVVCz
dm5MclyWT8FixJMpuAQuvwnxV9RV6UkVaxEsLZnOCeRHj1dJxB5/sWQvVHFFFZ4qLtZJF/7aV1KY
3t0ljDpkn0dwM5c0APMbQx+t8mvGgvsfjCCt229xyW1DvuqA7JKjoCGEA4Vlq8ZtwoHagEvQsx9I
u6vvkKVG33mZEZcIt4qjgWQ353+8OqN65MG/Q4jA7ziHn3Uh2irktQ8kgTV7jHA9+XpJOo1ivNom
uf8il0HBkI7tdEz0E1rh3yVZiMiUw1treqOKtJQSE2PFCX4m/hpYJJ6N0yAU89zBxeZu3FXePkB3
Nwvl+/6l5zb6xoMpWYsX23PZBqf03tgF0Lmho+c4bUE9mjcrbBB5WekKvD0j0ID5J2wrIOkH57sB
bY7BOmx3j266Cg06GOVoKO+OT2O2RUKDwb6MqLWXeYM9dn95LaV9pF8dQwPDCjAAtRMzr4cSg+eL
QhBeBeF1LirGv7IxQFrUk3Zvl/KaBEKGWvcLF1KiLJYko/icYd+oAHZ7iayYbPguvOYIdNVh0+ao
I2IE57lgvv/LKsWthFALaIf8v5VOsAFupQXzDlymii94TbySEASQGHgZy5rC9YN2xar9S7Kq45kR
DWIUtICVbuUQsDEbyblIw69jF9nvYEb4notU3EkYdfdPXH391W97M/MATSrGAzWZBuNd7RoTuHad
CKwT9VBSmsBG2ubE+EiLQUzfVq3NPo//8UN+U8/lJHLedutv6VEFCf/5+iaoFWtTvUOzWwaBfvdy
w9UprmJdI7f8pV17glXuwX6qXrkDZ+Kqw0M9s3OYaR9U20OH46+WUJI7QQRAC82XSsM3d1EtumKd
IXDYCLgZqT0VuKjlKPMqHMnj06Wze46aPR5Zw64bErQw4DfroTevBX+8FhG4Po//P1htsxlnJpwi
603A0NqQt3z25u4XFyDS1Fr+TfjIjnoQo1WWI3E5xrJY5IYFAl9C/RI6SYy0yQsszPDhczC9u5CD
8t/Xr+C/aHO3AiBseH8Hagjde9V7ZIDu5zEJX3twVVY7ccLJ+b0zvPKPIHpvbccgwuAotlOv11FC
0L/O9rNZVG+1+cq7CJkC1aKjFmys6DOibyUxhL9TeIhSoOZ3QcOjPO8bJUYJ4wGucfPAKKFdz7tG
2LkTGZW8Jk4IxtZ8fa6hbbfzJ9N8eCx04XE4E+7TBhu3pRrNBIUybLjHIsDZtOLUf0HJoANuUOOX
nL6B+HQ/VnxF/AHLa83EVvqgqgmXtChhrl6zwJRR2Yeqcz68zcI3i9lQqzhhyhIapgraViMAlL8G
elv4maeqtW58MBExqST+ZE6l8xSDTwdwRimEMdN4RSLzxVohr9G27H1BHoTZRdAk9d7cpB+Yf+4G
Ghyg6RL4FngKf+wLDxffI0KNkDWytT3fn23xpjyksLdM/keqtnixXf5wZciWt9mPPddkKhvRhC+P
G2LQ2W/ACy6s5p4HhRLjMN/UcT8Q7aKgVWJVWTGcya42SUQSBNr+iFvtDhIrlXIR5bEEbJS9K+CO
nVbfSlkcGdZ2C38FWEThEgCW/errkb1+lJKtn04KpG2gAR22xRqhHCiAr0egYPcgF9q3KdXLZZxi
IJ8wau9qou+AnGxkGD6/Qp3s/2W2Kw4slbunfJ3QTLlG5454drnW+ajkoTFt82uTFemOWcxsXOCq
Mrp83SSb6DKf1BaI9TB45O8T9bRGQUoERheCpXrtMn7EiMp+MjUYAufDuYjWsuORxbxTiqWj1My6
i7egPMcE+SMgO17VVhw6wstQUiO7+iLYUcxB/Qr6NGG5m+cWd9v3NNuOXJ6PfcBk/S+AD0fpZ9ZS
AsdEee5BTFCHuXYteFhV1Q0ayDDPYpZdVnVeKY18eIF0UNuYnNU69XzDdDw8GFLKodRl7npgcpFx
zVM5WQrDn6zeh1T90YUZsfmVI+vOCZhEh1MPuy21cZBnsUML1lVTmvzVSMRdyLKTfe8akPX+OOJH
AFe6XlLiqHhKhAS5F28Zt3MQs3PTvdksN+kSHYkHhK1rWqWvmpDA1P5rrAnPnpyiybKkfzu4wqcI
CQAepfOAWMKTfonMdUt0oXeNDjPVVUJJtlK0kdix6k7FbjmgscHAEAavWZcDAHs/5hDBTEfunSTx
Adsy9GHJS8UEUJTWa7nIg0VazAWU3HreARP4TvPnFIEfrCOquys3UlTUwbz50KrTe8voqrzasc4b
KhnrfQs1CHB9rCYMCuNadf9iPhIZWXQQZx+mCvYuLf1TSDcNXkP36NctoGsI1QXNWmHQ45T/BD0M
TIhAtCG0n34gjDAK9Q66Vrh4tainBAjELkdfXT1lMQr3s90l9ucHpKWy5fmslfcKwOeiJpaoOaV3
Iat7MrMO3YjTyiYw+U7uuacahJjAigZxt6AthNN++RURTf1IXeA3Dchqw8TVk/Y8ao0h9uQ5Y0It
dVn7WmDiYLVCxcb6mYWTNig2ujGNTrBJpyDaNnTuaW7Z5msJ/wK2rrDDsc6WPvlWgka/f00XNcTs
BwD5JZ0zfIpq2Wsb7XNwqnURYb4S6dhl361rxB/1goUtsJFzeuN98TgUmUSB7RZJJ/uQvvcwVXyt
47vlXHfRBuzLPLE0Zcgz8YRd64b0rn1WOuT6RT7JrmVRjRIWG4kG4gs9UuHrpMUyIdV4P5P38c+M
IdnsRpm7GJLP+B9CawHOHZNbhz6r+DvaDatGhQIip/Ue0Ou3oiJLZ1Dsgm49e2Jh1TDUasCUvoPQ
6fq14rqsyl//eeb3Sb7B0xwrf2X3ukWcHR78N+nJ7NFmLux0S7QXuiCEoC5IY6K7JjJZ8hG4Pz6/
RmxWxhw6elYQY0yWOxd4t1y3W+lotzeh6uWIqxfH+x8tuFy/3XM4ly1gJm4l5XEVpXiLMslow+3G
NBc1wHJHg9RlsHS42HLzrTuAgmFMzbNU1VV+phe15KxQeoig3Uu6LJKgfnZKfP2sXyvI2qb+Hf7h
94G9b1d8YuUQJhTda5L1g2McCdFZXJiC20itqDhQHnNEjSzHleIlcmOgC1RUmg7tY1/Zl+kXsqBm
3KXG5RfXKYdjfM3+ECMVcx3trfOVwQGFsp6WcHQYI7j28NupPg/nASiS5Xur6MQuNb2VJDOq26Op
4IhgVJCyTie+j5nl6EevRn3UXiG5XgX7RudNKr5yFR6d1H/cXpu+KepjnY46s8mGrh5CKMSqTgWe
j0Wb8OUzz1l2ahMXiCowMW7WzRUjobSbL5Xe+Zai2Lc4kjIU9M4pe2XU3jQkIlyLutap0UdQo0MV
eJC5uNn8drJxlq9dEPtgSlS+gXygkhRBCYq4BVFuDINDVwFKsBDgqcfw8N++XcOtQuAVTHJJiCI6
TbQ8UchTDjaPRWBxqhV0tiMv7lL2wkt0SbtN9SOVjLEPgtd3huHEq84yUTE1U2RHaZ0mtxnR0h6D
OJke7A/CBQk9jT9lG4ufHt0ETBNvMKW1Ed3ZXx/RqV86TYyRBMM5GngPZ/6f/gIAL7PAje7ce00M
hzgXTUQ9+5FHRnhXkd1hhZ/yx62bZLZs6KgzkzSOwWxrYiLl2LuNgOZ5fdxeGyTCDvlxaYl209Gy
dbmou9j6JrL2UDShaJJUOTIf+wAz1VU59xop50ZsXJDWjEoubiVymHSRNXGsil8WLXhXcA6R1rw/
kojcSCGnYCVvc4xH7GQyvED9Q5fy1QhR4dwkwyii7Jn0+bqHo6/JebN+DzuVax3E4JFYmUlu4wta
o7lmIx9hwWTuTSX8kb6+qndS7j/mNxadOhlIrDpDjqy9EbpazoY0XjPGtFLDRxqR2sIXSuwKpFmR
yAK/CtfnUaYCXHfg6ZEpIBzZBgo7fKkHDm8j4W4P8wwM5dC5tcSk7EJkCnhyj69aBxuO8B914yXP
s9gFJzu+N1nblvYGgIkRmixo/cFOGhkXmhcP3rtAc5+H2psq40E9PLsq7UrUwb4YIgnSfPqWlhus
LNavqKs3aiuTetFdlXfBE4Tfbw2DoKPsMiaNysvv94G9wVpMXLsjcfX863HJ52hMlbTR1OyPKrwu
KF3k9FsX81RQtSO3fLI2C9k8vTwttGTF00qFNThSVMlAgK1oz67lcOOOS/6tgzQyDLB+/sNS4zGo
/nAEC9ztUeNXqob2heEHM9QQ0838/L184am+Foy1UzEtlYrbLCaPMN3Q4fUDTrH2xuBzSaffoktt
SdDVjUFCdpCNfRPYEqYBqHR4Z/wxwF/l3gMnrZzcFbDmL718gtaOCWnYQcyPGa11ZTbsbw4/bKP6
j9yt90iZMNOqsMd5TSXfcZiCLAsebQfKXDkPLoHunuFcDakTH36yY9hq/vQ0abQIR0gB658eLYkm
/0ZOsX1d0uZt8VYWXThwU5A4c/3IiTVF/8q5A5J3cecnCFUkvgPXRtFICc+oBzgasy0PccwFiQPA
2iXPj1Gm/KdHN0Gm+JZt1/VuvncjwWhkXphoOgR6vKNXZQms60UAitxbLw2wolQ+HHPv/ygVvhPl
7wqVmcjMMJushvVNWHvuJgvxzDPtp6gNrfo22oiH4av+4drwA/RQaw8vnsF1hOZdkdQBlSVznQ7b
IS5oWP4rjSO75202oLkfYp36kYL2xJV2wCAtKHOCzGp+YLM4x1+jdna/ptFrB/eacGR1ZLRuf2BO
Gru2uOiQo4uCrZ3vEH7TxqI/cUADEjfY11i0k2XVMzB+R8qHJsivYZqmW2FqOW3EdBjMa5td34L0
0EFhmCtEVAC46uIP6amUZBIkyf76zoNMc3S1nh/Ju7b0GqYkuzn8XfMetBEFwDWlW/zMNJniAfWv
HThGTs8iTetDsEkpq8mo0fpbT2qrJnctn8sBG+dt7axDAkY9pkpkBHba9+eKaUPmX8+2jVogvPpj
uoXTte3VEDtbYlvDp07fLQ8F9jyuwlOTWAxnlhoGkvxtXSzEhCOFAgcEDVTy6cw7TPgrdcF9xolN
icBni8T4xNQ0eUQOT4CejIa+Nejch8Q298K6QTdCrAAfV1L3IcYRPIThuyUO6N/Krt6ekc9MRrT9
m45sOfPHBGg2WIim/UwlvB9TUFtpHnnX7jZOoDr6+fE3kOgIDJo1yiV1G0FA3b6LBw/bM6qFhYVO
g9QUbsrpLwD1oYDKsGj3ilrTCXONeV9Lq+gIitKDU8JUygHe8OTaty5V1JvIqDJdPUBp6QgTXX3N
QbwQNMRXCFTAg2ZX+cfUf5m2hj22PzDYnCF3eCsj1E3sQq5D/ofQgNYSZ0A/AP8Z1D9k6JvI+I6f
k1KsCawlaLs7fOASO3EBcwkFxVoz1d+6snEPFaFRiwCa5QSATFYi7S88Hag9bCn2U+Ujir8SbkTg
g1nqsAjZqLlm5iBIyon5GkuXE/lvJTCgJX+ntyOZl57mQomMfYSUU+sgYbyOIHHmL5C+aaRtfhmx
tsSSrGSkukMsE1pfvatj9AdYDv4ReT08Ec4NGlY+OFSwb/eypK27PsmBfk1zOxTL66KE9KUCp532
sX0KqSaKI+d8Vr0Tt1NY/NaKNYNdMPmzcbKoMN4yjGzj6ymzvTt8TceUOQTKtMHVEUOra0j0bBXL
FnX7G8OoWwTXOMGbXjDDzXaR0tNDcYA5qpK5nXfoM8xfdmWos6Dk47DGUj4HfcHIB+19wgwnKJaf
QD8zkjzvgN5NUo953ubVTEg8Sf3KthCHsRWk+lDVRm5pgaIMWPwicJYdogN58eHdiWfiT/EGEyR9
g/bRtzqtkA/ZjlsY/Zlq+CaVjhRy7Pavgku1ul+CJ0TIKsF7BX8k0lLWRhRPTW9F2Y2VuemdfV0M
EYFKKwqLiW2Bt2CPr4d78MxR9TG+ePLnJ+Wf30VrQszKcUqNQ8npC2J1WzlRprCcLWUQb3z9ZzXi
bDVItzvKEGN3x4gY3odP3RBYBKyvjyBcxbe43oJ4sDPP85WsbkM7zI2idwkj+r/3rs0MVdCkMg/n
9uyVYbHk728xI8mr+1WHRIZAyA+LsMzsiQ000IAd2OYaUyXpga8sfvZBVzIJe5kfrifDKTKejWCi
plmNq6m6sWrtCKJiKyyYenyvzXdN7iuE3KjO7fcujY5MVaFMaX20pCb/Frp1G1QNyB0FPwCZJQ2r
P6POYc2sztAvZRc35s5b8KK5wCOZ8Ygjdeq2wQEX5ytYWfbMQZLW0V+O3Tmiy7PToJxPZyjWGKCJ
PDhUGMuf0g45b7rUWWPXiz3+Nr8hfkIBoBHRXznOgcx2B15aGIsbTmrskaw/X3L27omHKNnJQ9Z2
7ujyonfF8zY4HTb5Nn4m8RKe2/8FsAGIl7A5Pvzcappsx+ObnJIBjnsk+YI0Uuo3ObDiwmXVxIqt
53+jmJNB1Krz6JUXxoDz+gWPka5IvujFKI3gs+Dfa1aHc6hluM87MOnnc38cexf4JFOdwnsHUgAe
eXwybUKL+6aGdkyg6x5RZ24S3jdOf+RzYf07CLSF0k+xnYJpvSwjXttxnAipsjseHsu7iblgjuO0
pJMuppXt6jffuX1Wzng9MDuO9gwFbm/53bcW15QrH9BgAJEBceAT+raoCYMv0UtpFJxzJ1AulmZR
xiaq5Punl6AzDoGVOPPlJF8XLgu/clUJR9JG7qg6em96Mcrb+tlaStz4xppRAqkHBEuT9jkOKgSZ
cnqutHWiOUY8WeyyA0SCcZdWU8R3XkYCJqWPEYYsHRtcY4MPKEe2xFiWNU8XSC5Ko0hFy9ayrvI8
XK6kazjTnYUxLkcpOt4b7EsaaiVpsMRuWRx8fJE/PmiQ0/V0Pw/cgBv//Ia7xfWohxkd4UhTHw6c
sA1zLnnVD8Vjq2iR3j4dWaxySPj3sVaEUWi6KDHup2RZPKgQbZYA4CVPyf/2bF90cohBAFQRVnYP
I2TQYQRMUGq0g/oHj7gy4uVkDfx5AB7562Gl1tQmMjHmLkjuKPumzZAPPvxfNxsM2ULpjlS1ZIGG
oUkXlX1DCdmkHunO+hnukijKTtPEHyXvuaF6RzuyNA7XTxkIfhlj0+ykBs5Mhdqlqo3LCCMtDoCm
cpKonA6KsE+KBbmyZtxYkP7Aj34hyuViFBFKYOoNwUEKq+OX6zLoIO7Ssc2USHK4Rhkgs3xWAUzG
Lo0oqaT497MPA97/3/APek4aojX8cjDulRWsrwbyyUMBmR3hVpcKNS4x7jlSUF6Od17vsWa2ftBb
YkYrfcOycqkNxnwCCwWV0xMRLZsa+oV3E2BhmDx7iWC4bcwb2o0gn7P4hNRHBgGCLYBEXwDMIl0J
BzAvagEYzw5CMOI7aBcLS7Ry+uWVkPbFOOh/YvLcHpkwCRo+LEuXIChJPTiUqnKTc4gDw+30KCHC
+lW20ROb1XAHarT0a+Y2ZlCgYc/1xMN+8z1Ok20mJUgnhk1FCaAWSeBACkfKHXJRV/gvPyBYUk+5
nQSl//kjy4V65l9oPA1oc5MgXNu+rayilJfgP0WtferDx6ocv3tS1doBj39rK/du4MH0Wc5PUEE9
DnDHvGAjApCk0O0wJvj0RU56RqdgVhQ7tbJgnNmCKWrkYaSg8aysfNsPTCRwC6dJaxqmhBuOGP9x
q8X0J7XddIvcbzr6kFXz3CbX6lsAR27XvoR8o64FpA0JhsbHjkbTXUu7iIk9IFgjWxe+2WiT5IkB
VbtCV9SOszeYTJa4lGd15xmDhov0x6T75t+46oroQ5q/9bLq6SQwlmv1+JeAe15cj7jW5bj61ZaK
1sX9iEqoAxALhC/4NHt5JkaFRc06U2JCul+sJmZ2OzkVu0PQMDw+CXzZUulPTjBJ3Q4tvCnDu1Yx
W7NnzcNO3a4lCIo5OGfz2Od7bb4UBrwPTZLD8hAKIl/KrgEwtfWRSrI5YaPzP4OgqrRiPz4wGdxp
9EURO3Zu9l2F/sFiSMqgsNrAeb6aRQ6rmRkAAAht1ggpx64qYdhSXg5dmkcUHBtez7diWpFG3veA
/4dW0xhOs1wR4vFaP6PXMSG/Gs6VaVoT9bJd8HK0oiD1DO1v182UBXuTtaLXX4mAjGIMQlnbi8rZ
Jw8nwx7b/qP9v6hVciD9B2PvbpRxSKtiWaGQXlGyrq6mAExZL9vFYR5jlQag+RL/OJzU6LNap/oe
z4s+T7tGucz2yLNRkvTNydDHaxSeQ9gaFFByC0fLfL3uLayOfDEJmZ52kkJYxpct+j6OtkBGlLJU
+6+iduR0uPX59A9hcgoTQ1dtq78oYTMGWnjl7h4pjyav8S+aEOwd3aagaorsdJDh/bukfdIJ5+Ih
ESdK9IwVW0hvgnKzmS9tOf8jjQRC+ZFgnMt+hm6mKY9Q+Hflg+fjBI0KbwJjW4zOC2yl9ts0Olur
PEG4oL8V0W/kKMPtfupeLD/F3HqlYenCazffRurfE+mtbRuZKB4rLuap2iq2Ci1oGKoFr9QChIlV
S9pYe+foni+G+0N9Yl0tZFwccZ1muFaT5YaIZ/DJe2RYy7Fbyj8X7Y/bGvMSziRTVFsTky+CwwsR
KaYf3TuGAy5RTqb1W9i+KARlqY0Fso1WpLP09krMM56s8Jjx9G7KPOWG9HeJ3Eq+nUOc2Uk8mZbb
9qxAQGwvUTFkCFikOW9IRlE0UfCw1V3+cOFv2tzDl+EG8RA6e8RPDbtzsnVPahGXcPhLTdXajGAv
asjXSljt0GczA9lMz9EIXiRvELtiKCeqLgXQ/IUyUkYWlCVPmKMB0WNB4pntV+0ZvOB2De/SATFZ
87iLfTt0Kjsn8V76JYluQMHQMfZrLJRReYkNeh0TZF8vO1iiC1i0+WBuhZRhM7O65DWifVH8oSl5
oowcDWQTCKBOsYtHI7tWCEL96YAQ4K61ktWNz3TalLJXIeOEAiMlyCHjNA0bNTbT81qfNiPxlOiW
U7ypv9eXhlN0XMUQCP75kXdMsunvuQTGqMnSWS5bwo+YWW5TcqANfEX6KlV/BvMGJEO8Xo+SL7Jf
vvznT3Avf3rtAu0j2jYqT1c1SvkDkCs8hjyRsTiCe8I7pGm4PzuNxw6nnvbXfODE/CmWIFSxkuIz
5+Bymst9rUTKS7RTieu5OUf2hU6jk/OLNSbQwv8ibmHlDClc8+vlWHqhNIYh58L3E+4ujlFLr3Fw
7//c/0/yrSb/tsegudxAVvbLy5lkOruzZ0UtXcNprjpap0SfOiU886ufvk6y/qSVcdfDPBAwTwwm
L7aRuRessSE0XO14JCys19dScSbjXlT3LTkZqra2Gt1B1yhJV1PuYEHSa5x3w2NyL/C09KySkYQv
MxwCUfr+OImsiV4vU0mn9VRzs+FX0Xlh3HjrueHa0qfwKbvuhWjKLL74RsZwbLDsmUUHKtnlnJoU
xuXgZIqaDRsRyB1tiS0BsRpOYcxA7Wiog4QfN+4JmU2kUcB5TQY16n7i2X1zUglguJYtqTPAIkTM
lDu5dUHzb9ykgYmiItaTOAqpnlUKYoVp5Bu28L7Lz0hH4v3sKkfUzg1CMMEZSdnpjF7+aaAOfUW3
0McTHgsPuXmRksbkta1ll3TUJ+mYoGXvGGH9JxHYWKwBqYyZnNz4Qn0maymo8MJoderkEarDt2tx
VrOVrHCHY+VofBNDgzkTKugAEqeTnPjhxjBq+0wH1n5EKebSKcZDUerhuBo/i+7SZu5HSNO2HJmd
ErmRUQUyEgf8gRO1uzstvr/R2hmYcGve6l73S+7UA2qMmHFJEEtZWAUwJM0vUEpkmgX+dzMOK+8Y
5GoeJkejU6jDAWgq9Wya6JmoZSQtGoMSyQIaIT25gNAJ2XILzkMXzPiEVtIUHKWcqc38Gf3KArH/
x7NKplAztOdJ7/acZRNVDDlxYMV2MeYBij0vwGlcmGoXt6qsFG4IF1NB3WY2nnaJJHcV39i3n1G6
90thi5RpnBzLhuzlz5BKYVXlcw4LncCIwAJX6FyVZcFC0b3rVAC0rHlhsA13IorRnhbmQRqWtKO6
jAWwSwnZzz/Xn5+Y6Wq445ZedQ5S/3ghZmGZeuNmR/xc03AU8I0FhARAJ5Iexb5ToIIbU4Wei2D6
UzwWiVxdfer0UL4DfuVn1sT5Jr7bo26ycRyqaygU73ijuH3S5s1S1xdsprYi+k/eJJAuDeCcRvtb
v5zc/4POCDsJA/v/lKKt6ZItGn7mV4To7oHgB7JWB0L2NyL7J8Qxb43UqqOk1Ab5CX44cH+ZrsHd
YTq7YFX4ydbmuXKM1sp3oUZMZVTGw+5tbW4NsMGLWgewRDOoEqDNQXyKcUfFm4uMJWZaqcKWxmd1
nMImmujJ0qbQo/MJXUHBNE4rsCL3zbDvJFyXqG/FE9SU0eyArNBoD3WIRYlMWEmj4AFi5/Flyh/o
vL4rFR7lWhJlSikR32NZ6KaIT70+TITD1gGEuwObsZajCco8WKIOExR+TA/EGN/1CUdK7fSdahsP
ry+PLReI6yW6L9qSvN0Ue7ODXIG5Hy+eliw6e5mIHiGXRRa5qFB+Hbo4XAaiVqATTxqNDr40pfCh
qFxSAKbzyJ9OWUor1IG7AzqjY3T/rbKbbT+rJkqLfm9P7WaWjQ63zJn2Uo1R5+7UzEhWw1zSfRdC
iCYsSAI2SdeD/XCoT62YlsZDNYKYIMFxQTOPqWCjAgSzWIOmpRUlkT7y50lDxpPPs7zhTbhwqQHz
yCSZLygfVXK8N0b7Htwc40rVrWSF8uI5rmr1YpOhs0fid+kBEDbXuw8JcrvFyrMlUdGfCfFesbyV
evJ60HAyMKNIS1WKEXof8R0iXbZsjUEqa3q5vwDkiFxlTXf78tuFhfTCbewIZQxh57K7QPHqFaIp
/oZEt8pQr/FIxBVjIdJzJ5Ly16JW3BvHiTHNDYpnJnOaurwopL3RlqGQIR6n2kUGAdnmq0Nbpph8
vzf8vvhzb4dnRKWo74JA4JpXCo39RkW4f1OMguzvNdQAEKmTkg5rA8rcOCOKCuAQ9zAx4kppITsC
dLAAzus6aCtrZqhNE5ll13/KUmomqL+mYigA6WJ2xsN9TS1KpG2ftOc3LKAYjSdYWoKg6vTMHJJc
LswdHzDiBivb944K5J4HGGpAvsfaDe7f43NKnl1tndUvjUwg5Dc6ywv4tvKA4SodTJf7LuN4lJFx
inG3shZuzB0ezF+JS6j3TZvUIt0eCTyzZer+aForVckNAjxxdnGTbAbbpK8ibvNGngLJcNEbpEQ+
HCDeFyPIDyjc88bKParFhUwsAnSiUiS+j9Nsih20GCWRQOR7IobyT9kOg3xYJzoxF0w6HR9zjmOm
HA69lPOQugN/ftUQlBKRwhfx6zGyXnIU19Z6wF6hmVnXqo3ze7sJ7fB2Ge6aZMUbtT6lrOPpHa01
V9kQdXEXgCy4r+syol1E47PQzN4putUpWgCnfb1fJueunnQTlW5xMdBPaEaJgNHHkkf00nZxKviG
4WGdb/C6o7fWpG5t8cEjeltJ/1HYV+/o08dL1NUa4/kbc8uYdCiGORwoO0wxQYbwC2uTF0pHsBIU
lJUduTNi728RdmCRjSLadZQ+lHz3b346qey/Xxchsj2J+y6EWvCUAkir8Bfo1aenc2zY+DxDquKU
fh+jJki5OORl58JZHszjEhLxIqLhxQmPgnmr2iJhIqCtKlYTh/PPMEM3EZ3XMUS4YGkiYFejaZPS
v0KdP8iqQJe/O7qNn+M/CKcDq4Ham2gk9zOIFHnqvWOFI+KsZi4sJGkcd/0xiNPbQ/ZETG+jPCbc
bCXTrNTF4wne++WGLaiYRG3ZAGORgfe7WeYH1AFjrYMT5LfyfPz7ji6pQcrP6mX2EYlXlma/KILx
w/KtTZJnv6xN4hi81SRtmaUoeIJKGTFfLIwR8N8dPyR9VSp9WXSIxSfRZtqqs4Oi/+fkMtiqyCjx
gUL0NRw2cPLVNauV0+jbhJX4qaamxieok0avdumHC6lasi3evaLlljGGyyjf8wAjNP54LtOnLL+C
LFbQ7l8nj8VO3PKrEIhObJbZZhhswaokwe8vtz172N2Yz8dxEokAljM8fuMs+u1FHZTaXAo81hmB
PI5Fec8DSx4phoHAnTFXsKHD7BAXjefWVcNYzHuK9Lm04vuzCnIVZNqLnjhsQ/j0/BGpwekDqeF/
fKmDxqfNp6wJQzF2Uf7+GXKMWPrQu8UYRV538pjuMEdYOxx+7YZ/qZGHZSxvNwCDfpajbjxdyF/d
OJg4QAcTPCvIXrqN7msnQSF/SlTP8tw2QeYcjfssk4Wm0502LSsOpETqzmp5lDhGahVnD6q0f9oS
nVeYgAbimEfLS57HOEi1yH6M1rYHOc/G654dw8LrMlJXKzjarlLRKAuOl/1XtQk/A8DsvFb5oV88
8JWxQCjHeVBPyx/sr7dxYhlBkoblsDeyP0al2IzHSnLDRNOsrBAHnH0V+Q5y5HsBuL6eN08uKgbP
x6OaGFYXWE7ZfMPVEdyVpIwwzCLSI3d7uAMWrHojvEMRfQ04hV1j7wHl3m0d854IDmkFfwp921v9
jSqSzG2bj0xc/2wRplc8YTLgCFRjHUkZ/hqCdtkLvK2W6NhrhOow8hiXQpCF3NBeWaoMz4X7kxd1
2d/U53m6q7GHI0ZOKcpvK5ahLEY0UgMeXqoWKEPnJj24zzwHqoaukzd3qtHiE7cTnXhCQrK8ONtQ
H+y2DnOe+i0RXLNM6w3yJ7cGrBqtiLwrEvLg2V2DoCi0E+TvRQcjPNGD1a1NYstIZmrH9C7Frh+Z
Pk3jP0ETkK9oxoL8v5aw5ih3FzyO6sEjOwPN7G5C19O8wm8ulOILhw35KAiWLzq4Jn6j9tkb9Hka
61g2YKk1AJ219QJfP1dcHQDWolaa4AHHes0Rbl1Fk4kY35vKX5DqJ1/jr3VfiR7Ck9S+OpO3mgxv
cxeIKii1ZSGdY9GXkyIMebr/reEYGT7+QV8dz+LdAeHXU1fnKP0PiYwNX56ycwPUedHOWSgrFM7k
Cf1hfo0Slmwwd4FdOU7qiu3TQYad1Kv8Vr994vZrXWTniwn95mhlHW0fq7AJq6Mg0mJRufzBj9ep
nk1GDhSmF8pwEl1W9LfOnt5Yz7hmK87+SrAkuy/4k48Z6/i44h7ctlSy7Kpz3CZ8FsvwfTvKCadz
LsCHYShwEcB/VXPLRJ84NtjodVRLkQVQeqY92UNiOMygx8tfIwPZescw6xyZFAMkBaRKMyTMzksr
z9r75RXC3aydOp4u45JeTiZoELtNUCAM1U3niHvvpvjf/zglzFOvyLyi1u7IaSmip/ZPbl7m/g5b
bU2nbXBsZJD6InHxlMMLdd/eOSr70xHmUrHmDIoEfA4dDWWGyuqzBIYNA5KvnH1vu4t/PEOhAI82
xEkQqJGTaYZmRwTPC3mEfUCHWHqq8NWoxw83K3eCmRcatVnlTF+Kct4UJ5ysN/XZscEFVWG4br8n
C/y1vFiXJMLQwkWqcOXKyANwZvBk2g6TRxN2KGaWJvqi5lAKy+hwcs0UR4NynwfjA8X/rf39ljdv
w4FNR6rNzcqqn3ZWgbbn2P9tFHD+mfy27Lzpvs+jGdrflaL77903/LDz7hBFAYg65jALHcXC6dN4
WPwotwvqBffjK9eKDRRf7u3AzmRl6gHties3asGCQKUxFVa9r8GuP95A6hS7WM2Jy7mYoxbRLahL
r/x1VBlCvgTWHi4y6YAQjDBLNqRvpDIRwvIFlSpKXnFV64nU2kHKoNy+3Z4Eh+Pler7pwU/g4hxh
XeLW9yYn/Uxhbj0m+4Gy0zBm4RtST7NNarEEoR6UGUVxrKurPxTjDJggekcCOyf+bV/uirYD9vUF
arAJbmH1vYEELmHoUQ7eS+qvMh4IAJhSXzAZdbk3s4Z4U7LPaitl1h5fEiX3Oxg0Egso1YTnZaTA
42va0VXRNd8iN+tqsFzN2ZXVDnSDMOXyUrd+hdHeZZ1ns7Rp7QToMhpX244xx6BM5RPJqcHBNQ6I
1Yg+rFd71oEa5BHd0EdEGvKroWKDGCLDRgAN9WiR5yLvQKyFHHHJq8JSHPPBk+m2pEXXcpCCVoDN
cXqMdR9sEZWkE0FfUXENCYYLIW9kC8g72k4gaerTXLdTqxZG8aysaRb8TbEZEywWdXduNG+G+UYW
SOSIhT7MTmzApmYqPFLJcbQL+lYT223MK/CKVJkCXMQZAMotXaATZ24YUwDQPpCG9Ubo4PhcYrJH
g+oaa4uSU3AnChQOtGfYkFym9poV+7Z1JZAaG99uIqqvOrSQpMhzMr5ktkPBv+VVDtSa+rmpCS65
Y16ANYZjRva7d0jXQ1Ojr0WDv4qD2mLq9eqsLk3CxkKHk3t8JefiDvQWk8Zxq08SMxXj+6wcFkUi
K2fK1yHLXUMVSA37n7P3FMfsoLw6oH7A/7tnCPKluDoLIp1a3WX7OLyFyWjiBmNt4eU2QqanGT2W
UjAP5Ge9ECcOVPQAbDCEYMzYjR3HbPEXS1YiNtC323nmKa48et0egZErrvSE6MSgAqMSItm7DHLM
4z+DcjD6DNeX6x76seR4lkuOjh1DLMDTc6Ll4epoe5wv1ylqK3YyrwhjZlsyz22VNbxb5Z01QBU2
tbbiC3reKuUwUqRvkFAQn08xL5tbhop5Jo5HuHCwNdLv8KNEBfhoyafGX/XEZJBYyIYCgEcMpLSh
qmzKiU5zsi3tuYSO2Wb7R618pX/VyqY3FVOF8ix3ULr+r4NR2qjO7tL2VyidkSOocZAtZbhPwzX7
dE8CW+xicgOhZpLzv6YjQiC2FMOKx55bkyCAk29zbMFhak189cikb3ZK/KHyHYYaEo03EjHL3m+4
CNIKCCPWueiB4pRHilzDSmJjBu92o7BNGo1Th20GUefpu9EzF2FejqGw/mn1LeKRj5UfsLjVm2js
fZ8e/xRLYHq6M/5xQtkuOXxZ69lSRitYWdpT13MYnie5w2t4BT6PClQmKTm51K02Tq3hIxCcbkvL
t3GJdAp3UKwo9mtbG92ycD8XXaV9Fn/NzQlc1kIZJeQXJZc3ChpNpgbesGfoQ92khnkp6zsrp+5h
1qps75Tj/AAR9I3bYjT6tdua2UCYk7TYf2zkLgC/C1u/9jkPRUl6F7Ohsy1kVsHHYiXcOV9Msi8r
G9gtoJwYoB463zEaUmvQ4bRviZkUc/ZbN3eiGo1jB9/Uq1i3Bk0fj5co5DwwybKbgHwa9yYe/cGn
HMZeMMmC+sWlJXg4Pbl5WxVmUdY5L+C0f3m3On6T+m62/nnzCbLhxBER6QvnghV6gpsEJAPfO+rX
zAVSEEow1C3dNHbqTEk/UkGd4RvJBA7AG6qnJNjBLEPWZMwQoDwT1nZWxb3ZOSKEYWcXNOr5J1Ho
zU45hoA/VrXHSvqqQO1X2nkfWBhtKmtq33dkWUfJ5mFzo9sUHYG/DjY5+bODFBK9mi/NX0ZndNbG
KCOKqWtIoQyzIXtx9qmcOw9BvmNZ3FmhpDhsWxZasCTUULVxP6jR1Ioa/Z4h/2B9XFrsJ4o+f66e
MHEnuziulvmOn5jsd/SvCdA5Qk8LbDzRAdJv+QPqyGgtzhaAqiT85YtxqiX5JvHUYqQHHtAqMWn1
vZgSHj8UYK/+PC7rpZAWjBczlIsy1zQ6BZra45/JmlNsXJqzc3CXa/KslrnWDgQ89x4LKWknLunE
NA7uXNniGOYyHUzNvvi3DYH31b8WIEjXiEicTNbi+F8LUYL0MajVjocUgksWWPOFpDAtQOZqZUZj
F6m7E2oJ/fguf/sZubTTV9CqSTtV/R8PKIGEckZcguBwySek0Qu/64eM6GxZ+FFxq4QuW9bZFZUH
eRnPTiSjswdexvue15E5VrJSzMv40R8is/jm2JhSjaX6EbzyOHTg4cPGPQwmGnCCJm/LQFs2mL/e
aLnjtzXbHjZgHQ5drNcPb/rV9PNcXrc4wZ11lb0O/S8USnzRrwOnhCsK4Pj3bn1JwM6Z+xjtfyiY
FGf8w1qNadz+0DbuLJXhFcJy7O8YLjS0TacU6xIdTP42ZOCxi5mDzZPdvM180Vgau0otBVFqFWMt
XFMJS1BPeIJJ9clC2fV/8g7uLtsHZV0D9bGXrAYf2a+dBlS9P3sR5BevFog/s7SS71ei7g2s3aCb
w35FyHASr/hhBI9czYBDJ1pqhKcf+8wEaile5XgC4s9Lr9pAFrA7txmtRxxGdxPzMzj9ZWREDZGy
xGBEHxXHeFUTKtRdFvXF+pow3hEIDGkZX7qH8PqqdWSam5v8WR0c5cAjDJIO13lnx/FMeXd9Ss31
Mmmp8hIYlyz8XXaPiOFU0AzipDN2TXUjcjPRpCrtxAUpd4vLIk8GWvWbTeb9jHhpOQIqLnQPs+8x
EQ1sIHObhXt0bL993ubjVjiIJdfuuFTZBHyB3R0crSyKMffPvj2vyjSWvMhlXjloQ+B3HXzr5ztl
z0ZlmtkjO6GKXAfBHp1SUBPMou3TGmo+3+27Y8JIuArn03KTwmP9NGpXRdJNPp7So4zkQxV0Oamg
Sz6rDyHsK1+5lV4RzLqdXQ9w/Zf9IvABwINmkTCzwP5L9ut1Z69cQFJ3AsxPGnzC05JB3OPeQBl1
eicu3MQdHbf+v2Jdeioe+DH86ne44UTxS5zfeuHV0JVUcu7qETiTI+HlnF6XLzd+VFT2zhjzkmOM
ic014V+1g7afGmcces/tArn16BE2QIPQ13QP/Og1fpt1SUr0cMTuZaSb5ZmSGkpsXxxmXKUCztFP
QaYVXtQm0FkPiMirveqHpS6hE25OuwWULpRPlfc44t7zGSevIa2w2WV1vEF0nXHITYoUm5Fogen1
waCR2jzSrsbj4iOA2ByxdlNODFIIe5lXfCwNTqcy6n9AQKIplany5osGgOFAf9oaIRGDbX1c7Ec9
nn3osgjpxF+X+jz+z+aO2upJy8yrGmSrqVeKLIjOVG/rGXJtLnOifHYYwwrGYiTxpw45RfImQuiI
e/f5iu5u9KLV1BP1ZfNRXasBj5tVOKK2T4vlj74wQxIA0mPonvbZvg3mXD8aane3S2xAXI4TmH5U
pXYnLpgKSRkI+cW702vOCvW0jdizZh8pz25z6FxCGcgm737dKGlNWzLPdGaOrqctFztfvsoJ6FYO
sVpYs2OhGoCHeoj199KlNZZf4y6ZGe8F+L2un6I0ci6PQZrWY0wmGW7MPq0EUtPLpvFtzZZP13CW
p3tvcAX7iE1SZEse5//SpRBxANv3gs/H6duawHypRoxfPhAf5D0f3aRY27RywRcPYpBT9eZ0XHym
+aEldbfmcqOOPhmDXu4Ur4KXcLK8t7DGqgpoSksW8eTY+I0zb0+SeR9da6tLAnMPZjSScFTicUNG
xHHKjDNfPQR9dNx1Q1msYpGTILG5YllYLHjqh4iht84mEiC0B8ozqAECrWTe7tN8VuzSvL1Xjpzy
sNu7+fmPuucuOc7pK2sRN090MwqBjrhAK2tbbSSq27KAw/QnuhtQUDP3UL88idfUt+ybX3O8g1e0
zUY35AEuhigZBcDwFjMfWUa1E3fdNC1pj0TZvHxmYEQG8VyR/nFMTallSFv0DAZLI2d4oRYWUuhk
9sOjRIBhSx+HXlchu2eXvCsbcfxfgi8S67govPv4ZZkhxodePfQTUjVdUc4ZUXH7dJZ6nQkurZi9
Fz27j49OCT2aCvsSQhsg0vT3mzYfrzcojlORrp6FKQqwYgut+g7ONuls8hskVbJdJCkOJaU4/hXt
S9oZdf1V4bOTP/ZfvH24oysO0qwioTg1Wk2CX8aVSUegRLUF1k4z+7XJB2tdBKFE2Nc0yEtdnCcv
+Vg/3QFzH96/OzTc1NbDF0w+BxeIn1MnsndzhXiSK0SJXJ7kXG3lM7xnRlhj/+Cy6rHnbFV5fuFE
u6xEn09Wn8iSG18p9XjUo3Kag0+XquE+KW0tdyEfe/RbcNab0liduKwip/qfIVHdugBHoQKwlKhB
BW+4QZNF6QMklZJT5bQQpxfZ1KBf8qincGNpxOak18rw24YA1TyJMZHDc/8nMXgnOMWm/rlDBysj
TVkm9KkPXrYCeMM0dj85t7nHzDWxe1Bc7dEXIhZNbRpH4XhEVM8mPAPvUAXJYmF/ltqvBiGhAlue
rsXDOL5CtPGfbWbHDHHkK6dNFQma1DPMElo3kZ8o2V1nONLA9Hdwx//9rTbP9P8eyQ6sWoIvWOdX
20Q4dCSxjVF4psRTuGjzzFwb5C9i3BjOsZGB3nf3mNs/slT//IQDugjmNceaR8BlaA0Stk0q18kC
VXFMN0lxmdsvrRzzAPa+65DrCf1vttWUKBTuTjLFIys6fiAp/NfLZ+8iyVkgWJBcKAUw6sjFImyl
TDapzrLzEuJQLLevApR1KP/kKJY0du8YGBo8QhceV6R6zUf5gIn867Fjm0JavTWqJleOsplsCkms
0Jb9fIP4oDdwJSKr/TV7t9W68//LLLQzVEV0X6cZ5OTihTcfocGBgnbOALBFBE2ijJ+Bf4O3XuNS
W3vrmjW/uEDzA0ZTlO7j8EPndjz/oKU6MDK67CXwQjg68tLZEEbd6jt6O9NaybJ9vM7qfX0TjxEK
DuSW3h0ljOMnF5XbNUk9XJ0Ap6BgM9lT53l+//TgOVNp3DKjG/SSYJW03t5Q+i/YORaB24CrkJUw
lwhOI+Pil8XzTpAwNkCAPkhQKefoWHHfqpRQGynjBYtiqxhSp73TebHdFIV2oKL+eF4PTGIanENv
ehSEzgq99DaL5gt9MIWacTCzeHHX+VI+upj2IywD8Z3hHyHOaRZYO4APljDDkm6v/7UCdE53mlD5
b4ZHNPk+QXVipyi42Q9CIWJe6EefXrkVbL79RxzIUAaNMRm/twsDiym7SGLSK18m6hXzMfh3j5H6
IyQLFbL5N6blb2OIcwrj/J/F8UCF2mnZO5du5/t4HizIntSBp+4x82kjDpHtjgLClGcex/mqoUX2
DRAafBZAKtaMXLkmumVMpha3zhtBiQDvkcEwtbyLSJWfPeL4P3EKzXMkWv7W7hACyodDgUEgMwVr
o/gNBN5lpJB9yZQcKDUu+SXHcuDOxdRQLuJsy+lTFJds6e+dHhV6aF1kr+FWarA/tqKiA1KUp4B3
CV/ZTtbFPlIljjSDTaqeQaVr7M1JYBJKDdgFdReJwdyedSlqwUTeH6bUFAgaMC+64gC0Sl16qYAc
PFrCRSFpCQcsdNN/F4LH6p08Q7F1lbtAgAu6c3iR61SpOeXThTbJBfVWl+rSPM7dJzETuf/WgcY5
NYvpW+rkcpO9ik0nzDXr73+LuhVZUOO6whXpgBISdKgGDvzwsbYt7d8b+12090s6hu2h29HqSkG+
29MiLNNpWdJ6cMiFifoNy93sYtb1IVxsXFALgXhXvCYJwRdrCFx2p8PCftkyq2R2SP3+O2R50SCH
ikwFEnT9tOHeKwtg2AR5uDObKlexwmBoT5ZazGer5r/LEfNJsnalINdnpdNvn6im+744KMfghL4s
LDn/LCgdfc+uyu84hJCps/Y2zCJcirUPIbmZRVTwMXHWuDkLzPt1QBlFs18tj0Q9Cx6waUqQu1VA
dSvYhUCqlfLUQVGqNXw+d/A9HdvfURSmC7KVaSf4WYNg2oo5fhugvCXy8t/P4yvvhmj6DryqgjJS
GJUKM1l1IuCc401AI0GCQYHx7NuEff4eZy8fTackrflJwCHWS8DvszhEmRbDEaejfpCcOdAhPDKm
aa6e2sHsjnXWINEsVltqJkixXIrscdIam31qWOboJ3AIGkvB1yuf160N7Bh75gF/Unft6TGP8wZj
VHIA7sl9y/ae6qTfFVNRZ2U8DqYSdEvRb8TljqHmtHzB3cD5aePpJYpUpIdenyiMepfrbvCFbo7/
ZMExlfu4eJiBvMTP/Kz/ZYxR68DUGgGnuKtsj3S6UyIR9mSc4NcpreiURQghakh6srj86KNVa0mK
AKoqtaW7ZYe06j2TiR1tBzZc9/q4CnbxS924vzj3cVQc6OwblbwJ7NdOFNkVpsqxcMhcf0btZ2Qp
ui6UxfCNJdb5MnTmKALcZEXR8D6lnCjhGDryfJCn0CuElBaVF3XgIBx1ElY+19WeLihntWB2WD/y
tDG4Tu0Ny37E6WXk2MZ+3rrdWd+kPhdvLv8xVPSjLi3kN2K2NB1lRlk3SCe0EsMgRQ0hsphxPOQI
M35J/kj/Rm64vZyO8xLj3+ti0Eh8n75UhUXjSNlOCly9fOdjs2zOFPfz/wliWJINEgGLoghFcGx7
cF4BdpiN17UqoQm5KQnWDfSzwJpApnnQozFA9OHPkmxByHXWsZLO1VLu7pUMPhrY9soxaojpc9/9
59U+mCi5hsGUffaOCqhySMMEiE9HiWRe9PqNyfMvKdl4V7R2sD3QuI26t7wGmD7hbxvorU0+JnV+
RFITsIZe6KzRywXIgK8nwyWnac0CtRAVrXXsWW2htZXZi2Bz1FSYS7esJiblyQR22W5aM8cWO2jw
Z50YJT5IBfjiVvVBfx99ZoJzTE1nx3tLlg1NF5EHbUZ+DgcnsdIgTQugOVmrCxmgZNrvOF7xTwbS
pCOzw4cVJ/jvdGtYZElu3ksnVCoqdkG61RRQt+Rl+tWYBTs4Jgg8tsNTjRf+x1acUZaPiHsNVzyG
dV6hWHPiHJtvgLfN5+JYKGXnGQ36qhKTvMPIQlkSBzdvZmKG2p72T+Ck/SPe/XuY5PsiT4mqzvCA
6Fktc+1ne6oL25Bp3sDaJ+xfs3YKIbyA0UtHjJi6DbxOIWRNcEFoialflAfiPQhrQhfW4BABl7hV
/K8MU6M6RjhFuW6kEF6ifp0pBDK18P2g64DVycKYlKyOzjTtEYCS9radororRjHX718bDwDilG+C
/1/dbjBtICJBhbsyGMJegbAkilTDQCw4GPn89pZvAYoKEezUCz80TovLH8DG3M1/wnEGtFzCsWx1
zcXSNcNtmGF4Z1AHLx8Yq9ZtNMtp/1FIszhD6XS3IUKjN4WLGXOSe/aTSz9hZFw5qg8wE7NGpcFB
P2EKuykHoi/eUAuZwNXhg7uk2Ca/pahWG184VbmzBWvBIJSse/7WNfsf537pnVUkYPeXaYe8U42p
+fdmkhVwxz7tBVam6t+wrx9JpnTmbIeMmfTNheD/q+pYx9LCjJ+poCWXvh5NRPPHyrn1buRwGZIP
JS9wJD420CqtZVndDPi00eWCzydoHywEeHRLjg4G6IhArN+hMmUobT5v09YVHzMTTM5u1Z0+0UUu
/b43K2OZTuUfLdFDUX9HwLaK5ug9LiGBhnxXRDknFrR68eAB2RM8Pj/pKs4bVCSKNoAuIgh4AU6y
hy7+AgugRok0IUDZFnLzqZ0MPV+NuPWqoOqjruoC1ZkNATeC5l7kxszKzD+d8mjEGa5cpEDR/0tl
1FlWqgn+RlImC7USBKxJImZ0MuzFQB84jgTwXRdHqkU6HWo8m+k4VidIkZQcAGbOkOGwvQQ+OyQu
QoEZry3yUh512B3pmLhQhuM7BFxcs1G0AJladoJhADNLCbjrE6syaQKp8dcsCBAWhJaIDfta+iiC
1q6x73u/uMOLpFsB/Qtr0y4Bw65PnvK5WzLF+Ff70A7NEUS6iDTjeS5vM8hEkcA44MJQ7QzD7lXi
g6466fvFTofg2chSh/XAVIyxLbj1Hpl2UdpyrhS8uhXHT8wjrmL6mptByZpp00XbSIU1RhWH+AEK
iNYqcarb+QuoOE7hLLKiv4xU+SyLBH+fQNvEbq5o8VCcMTL+mLF8HTzhgzumyEFfEYM2uphE6fd8
v+jo9CWmwLHrNFQEi8XfTAxWDGYmwhBayKbOUifcjmB5iCSDcrTQaFPLd7quqWhzGhO2VqN/OtHF
aYOoVN73tSs/3RV5krTXdSwBkDzHk0GFa711iOaVN5LG8bqbg+/KvYxUI8fOpbxLTYErz39Dyj1q
TD5CllMkMTmmOfbqJkxz38I1aIxHr/IzXD+UfLQhvES+OXTAg20rGL2Bt+P/1t3lxfsF3FejgzlY
LJZ/ERXkuTb6ToBy+XLQJcPteuRFHnwjYFEvBImN4rZ5MLZO2XTWtGrDQzORmD/vjeDzuklOY0vl
dOR0NI7SuCyiDd3WZASZmm+YOPTBgqmhPfc+seUi+xceHFZOqYU380N/sZuR1/rTIIHM0IRa81gp
AkqP1ThkqF3xhqFXdrKi9b2FS4F5WhuubaQmupeLcgR1p5YpaYfIsWkmeOpcZoqFA4qqcRHP3s23
RMEv1VR987NvO/MWDaAo3b6ojly9/Yc2XHxXmjJ9MQ081dUtYHzZu4BesjFg8eHEbLZk3u91V1iC
suT+kmAGapg8St7pUAhh04DyB2B+3vt0pnmKpdGs8Cx1dd+P35YTEWOFQxWGRbEWmBvbm7tb/lIU
W7QDTLkV7EofaWsy4exgr7uRp4C0hSPtVKsZWw+9+EsjD0jU/jHWdyj0RMYqeHqMuhuhaXcPgZT7
LLsSDGzKaLfb3B4LUEZZyPIBtYhFXTXvg6DNuQsnDCFhhmJ0gItaJ4dkntjQbo9xU/aDiS2ToHRj
u/rXRyT8QUHyjKA7x7G4CtQ8DfDZ1xilIaS23QLp+QdEbKmTwEebL72Pxd81gVEYyedy3L9nVJn8
x1EO+mdb/wzX/1ZzEoTOqtQYPT4Z2k8nm2wk9BjSZNiYaJRz9XosqSeZbhADmeituok5clSeJqDu
aqo9WxiDpYNDF0Yul3vM0mNtiqdy78ggYx1WyXrF3Oa5cnksodHhTpUmRqq/vJXulZYFTezghTeI
Go39htONyz5FqfdwzgIccGqHv7l0nndE3ptwuge3V3v0mrf2zj6SZkTRJKr5//sRk/10evON/3fl
MdvqQaJPAZdyGyYY73T7LrvuxoBwKSIWur2JJjt7nq7xeOPR9oGEm2vLXTXxKZkQ6bpINZE1v/Xv
gnKqIuR/o7hRA0tfhnG1Bzf2BbByfyAsPtER/Fsjqku807X+wM7DDiGarMi8QJPVOC+++h8TAJ0+
sSSgQMAiKi+DZMPvYeS3cEd0RLHvlGqTe/MLhNmv2IjMMtO8Dfzy50Fsv3XYR+Gzq+3KX8bWCsrv
LKYQIbDOO7/hKDUWwQy4xe6guY1AK4eCHmCU9NbVNEX2iBglqkKOrtVPdfV2H5jA3/bBr2neKTM7
V79C/l6G7KcrgIj/P4B2bShn6Ua4ASF2tqOtgKymQJhYxz5TCjnp273YKzKS5gxJQEs3RQxe+IqH
pWUdsRD5TJ2NYzroliRn2Ea5Exf/YEt4UkDTSueW4xcgR0kfyqt3ehXve5vfXnGRnGJkSqyyP/6P
sDFmDk6WNeF+OgcDkqY7r9LtTmYA3OM9jkZGOcwarv/6+QYKdVt4BkQcWOshfsfOcKP1D7qZ8Bmm
bbp7z5DzLhV8vE1JD8Bvi3DVj8+Cs5/kI+qJ6zEv1yT6GaqxRt6a2EXMTzrboMFeAfoEDuUtup0d
NAv5EvQACsDJsVF2HOI7HwN9wWcmWvfdi5hSfOZCZNNLBv7FP+FWvWzmQMMhJxe4CGSrcFnXIZKc
wOa1+9TmyRPjaAVPPq0x98hpGbRmR0IOAFJF3l2CeY/5rfy5rutdbXKOYPyaD9cQAVQ8CsnwoDhd
zSIdEgP00LwnAvK85osL+bagCwFWo+JOZiK3BuqPkRd3tYD40t0RI0Q0r7kM1y+vboIvaGUdnAk8
U7baUFoZZcYHB82tePmBs53lXOytZhiYIdtZLc1wPJkn2seoilv+r3dlfy1wTI9rRPslFSCZUYrI
lcrpwOzm4T3urz7vAFrjYHqp/KxA5VnZdvdblySoXBHUV+6ePdVgUnSQTvAnThLO9qotzERVPOuc
eNcwpUQyRd9UFSggH3EaWQOjrPlUAqFSt13eYxFsgZtUt51gDQsMQ95/8LUZ5LzONgCbeDkAbCKA
53qN4V1/1fWUUf6Ay1XtxIzdKQ1YhQgU+1LNfWHWe42/coBE/avcoXosnMInH5ZtqBBvKHG+M0z0
7gtDQUvnfzuFhah+s9+rAHSRxkWadRpsCoFfacplxgkyDCuVmZ7ROZoiVFYAA1lcHWhxHMKM3Ckd
zMpiN7EP7zXI4b+4RF7OXwYNSUdSkf+dz79X/+0M7r0YRDkBRKqrbRE6Ub/qw/utXb7QmRjipYIu
4+ekCLp+0R8BvsLq/6ATpCWsfFUzW7pN7/XIMtmFg13DePY8yP/tLX4jhsJ/TXSC3g/ZgvrG//83
Fzw0d1us0QSUNgbpGKbGwIix6CdNTtjtouF0HL8gyS3/x1vy/BCLwX5/th0oEcY8fhm4hpxRnPkH
366xG//FYwrDtCy03FEzsgc6a7TiDf7khfzsUlz1wDlsaWVxyX42u87fz5Ag8LDQoPQ4Ck6JSjZ4
0Dl3u7HA//scewLnsMMIgC0HnQdCA0FBMFn9mr392bZT/Ga3kqY8uOZaqrn8xdTK4+fuLwqMDMK4
Aogob8fkyW5HAq/uQI6jCbUT52PD86ughumvcRqJ7qkS8DdRBYhe8v02D7vVb7xhGoYJxkeH/kba
8En84eo0oEe5BBaJF5qxcutKZtflkf6cLdG8MZ4lx4P1KjSu7PKdZEcQNZ8ayXuNp+HArNsvhEBf
9yZHB/eDP6RhqGwkqtwtERAnIdpNxmjPqhDgwgDqblX3WopGuD/hW9EeoONbiqDQfVajSZ9OzrtK
l/T5szZPnqvQQNN5nvYdOvHC8xD+MtNML85F2vMpuXJpMR1tdVw9SXM5ocWTXtB4TqLQ7p1/8nZV
cYUdisFpMrlDkLxfm2iHeWlu/F7rxKrFnx4ZHaBWs4uobn4S1iZqaVm1agHAzWjtDseKUxikj8WQ
V5B669rJHKXtcL0DcBbMttVs4FFOzlWzSCT59WO0hzsAXPVVHD4xijKd6pQ0nqqsM4fv1CpyDjy/
dF4qn+fQqJCllAYhGtmbpLaPxKpyrp+QY4IpOJHTEylLZ19WRMisf/lpjInR87V7Kev66tuiIa9O
OGKwA6vKhdMV++2BfOhLn4X+hhwUgkyHhY+dMazhIJmx+r6YJy7t5AivqBJwyOo2ZGpjmijgDV1P
Ehqr5hqT54w8+ixBk9qZ5A0R9hZQ9+6c5cinJeZOILzEpqmXRo6PujA6FjWU/mZHm035kIhyGpKt
NceHqmhsfWJvIJtAhs+o8pRSHHAhLGqBqh5jr9POZ8T4O8Ai1EivJhav59MHgqJrBIubrmJA3FEz
uanulIQRMdt39H5QjTl8eWwqX8Cq6UYmHLcw4lJamvRwc7PC47hgNnZAgt3P1yFbuhQjtJ8OAmA4
1F9jS8eb0E9FIEmvgI38xTE2F8Wkjv0acWK0l0jK36mMXRpQIpfdWFXn703juoJK3hEt2YooFI+4
jJwYBlHDFneFK4GWDqgCpghUlv/eeTjccgc7ACkWZ9dlvcftt2iaokLLwRdqvpjhGctkY134Buxx
dNwsvf2y5zCGVX5gTeiczmq5FhD8RufIRdciWUJL9AhqQhBWykghfQH3/dBm4pdWwdHrobym1vqp
sZYgzkjoZaA4tuMHD3B3bP30Fd0NFp8G5MDiVYTwMngp2arDUGrhX0wknie2sROf47Vj6P08u3Ki
CxFekm+TsF3aT9TkNkIbWLSn690mX7v2jR3Rx+wGQtFtysLd7kayLgG54lRKhuDCzH+0GCa34e21
7l3tacxbfyQdoIXZw3ilHXIDvTIHxxSH45r2u0M1TcJcpVDsDDZdwO9wh0LdtWZgmwHLKMlXW595
cEblxx8VfvCU31PLwQZZoKrErWCY7rIMwHWggvmeGVRTGiwygXG2yLI80A5p6kI5TehAfkX+zOnl
xmNtc8xUfznNKxK+ERA+XTgfRDzyaixQBiPn9cKooqpflXMCorDWilH2VEGHy5scmkjhnm2Qqy1r
gQgeQnixypuxILUwVIXMMJGHhTPU0W/BvBKYxuA150dEOxujer8cq8Bf7WNVGGpwBbTjQTomS9nQ
L3C0EUpaEurON2koSbw+yEfm8zOlvHdhmGoAssbJ2TnyC+E1dOXODHDchaiZYramcsuwhQKIqR5c
CUj3Mj1l7gd03IABEjwfRKihpYB+ic5bF64ig89FtX0yNE0z1Uqy5zLNkugiEXf/+6Hpak/IY/K4
CSN0T4SCXuY482sG2nS8UglAP4dpZjQdZVYm9s6HmIyKbOyQIPcFkZQInj1wlpMQ6+HWPx5yQGMA
dACNGCmpnDQ7026Le8zIsci+xJudlSRFkNoCTzognbOmG2gxfZUdDDlFn/bFw/Rz5v/UkdxRn/Yt
fIA+cL+Vq/x2CfFcSEyhSKoRSJMvU3km3yiDQkcPTZtyHTm/OQDP8K4hY7H/31bIRiCngCR0EAJk
D1lQZsmQmWaGxJ7VFPe+1tbxAX2KntPN2oCcJ2nO2pWu1JWw2T8TQ4kxqX2u/8UJ4vtp24KmAETl
w7RsjphfOhcpkjRcYpyUgs9KRi06rCM6yDeecUrhfUPFupst51GF9eawNSvjaFZIP0c7yELMhmtU
huVzuMZcSuxUZ9/GUp1yzjWV68Px6gS2gCxS2kg+86WK7yHVmF/1o6JvHJbbFWbtmX53Sub6XJ50
ih4LRCdJZxOUQPA9wpnMNWqMceDjyRW9kIHhhfdcZqT5Az7O4B8SQBK6bRfeNBS+gUiXSnfLGbQ+
Y6bzzyVgTjo/fM1iFuZn1Lr4C7Uy8yzrc4Eh5yT438z1ACzWZ+kRtyuWjnB8zfet4NPeldkc900U
hJSGMlOBsGgdwiw+kxBzf1oHAgKbhIMn/cWkDD3YklNrIeevFbRHvSY6+iooztQl+Q+lmv6ETcOD
1/jsTStR9cGmMXBLzWZwHc8C6qP/QVsU7Fcrc+JU72rSqXcIfrTnUmGg1evDKAv3t8cCybJXajyD
U9gZydshQQc3yd4RWY88jGF2Z8skdkgh0wcZTUuU2l2QC2/W57kXKNuuGkujE/dVEdu6ppC+FFu9
NSpPfKgM1pFq0dcrq3iB7+Pq7TFkn52XcIR+K70QK6aEhs+M3thxdPZjFdNacIsSJgY2JGGtX41J
oDPmlMqNmIogUbW28GjrIfMI7h4ZlhujadOw+9k7Vd2mbYMSnqkzthO0wImTGKnnsrcncUe7CdQ1
hEeHYqulzjQRF2MlefW4saLSUL3ITvnxAvozRmwtOL7IELROb9fvdSQKvPOthdLDc7soy1/rhwKr
U9khLjyEjK0z9RDOQivmubTNtBrJQOxrskQ6Ft7/1nktnBNdizovozJ2SM6rMVcfPeHggIvgZJ3x
1rfw/hj39TfOZS2deXB68bg6pVaeltyArhrk+D5HPvHVehvv+VGQwGeyBM/0OCYRYYmdLAZ3YQHb
yDDRmO+Y/9Y+QNMPxP+mXr6dKH9JEDRPOZcS6LBieL2B0YfpgX42drdl3PX5Z/XG/1KYtISoCFQk
T9goX8pDC7A2Wweo9Q1Ex0XxB7CXAEjwHVr89hdwZqx7xKccTL9pmVQ0HhToMKa3Y59bRr7O3OB2
7y4eAa6cDL4H6Km777aK6MvVk42WC9fXLqYFZcX35Iy8IY9eNFJLJzIb5Q/ivtn6E5/F7rFQHiO3
6SGNZZwnrtbu6vtgIzOgWliQCRGqbYdacBdmgp/6P857rKPoTJrU/a5nXlo93QkqjPf4MYJUMgk3
S0u2bWgcpk4YIipCqxVxUN2J1ioaNM/2yoMwzpUgzU+kR3xT6kMXxF2GtZke+dM0ahodNrQqW5Wx
gM6C3m9SEUcwyckh7bi63p4hnFmloPwF63BJdb9N+p6b9eCNZ7SpHHsb9NxNHD/W3mB1DI2Kh/yH
mKUQO2S3kHJmaKvLJJmJEbqk1r5mv0ISHaJQxwagB0Idfm8TKc8jyrvBw51NXADVbh2K8i/Jf2XA
R/rnDe+9gw5J/mN6UjXrg4diCo604qL1+JQHKGNsG7dBV7df2J4EsVnKfFwSRGunkYlRJJHM9xrt
Nan+GG5F9P6N+5qDD2xD9Df4IQ+PBewKoSvfiBVfcXRNuMIaWSJT7vKnWt2ggBVkkNZIcw2A+2XJ
QEmXsgHg93jPHrPRkBdhyXaHX47ivKnPSkumeVHUiWWEc6vm6uTstEmD3Sg8iqaqmxNrDobzzsC9
NUMu+E/i40mfnoda/y7+hWEuX5hKTeg4YLB2R2OctcRwZBMHoDrkbIcRZ73kxkBRdp3xnBEWBy2E
AQJ/T06tArUtYlH6EZERfbj7bgje1icu4OmLWuovc5+/mB3GjVMQ9k6URbIN2cu3jT0AJp8Ax2ac
oOu3hFfsYg8Jd0uDwwusO5v2wiYONJyFSp0y65+jouvpDJUDzdKo5QKdA7gGbiZ4UbJPhPjvtPqR
6Evl2WYuvGIS8U5enmmpOAR5+lJd8xmKIHy/hyB0f6WXDslmyF1iyPXRi8xHpP8SMrfXfnrPCtMv
J3SVklhMhC1MdTsDGb+eA9sQIOW/asm+dB08Y4Et8RChxuXXTdLRRMPCG3PT+KgfjxtSgRPxl4Gz
UlQr4nHhcGZhyXSIjb3TNYNOONffnCUTjpwQGBg+qzD03QejwpkGiPZhIMJXnWo0EkP6vyZR2xUd
+XoKOMxbETrdiIiVRv7wQfAItmKbSU0L4cUuG/DvG2TKBJcdgveOP7BKnDDvKlffvTmdvkzRLoGF
veqvP0YQIoEPvk4pT/8jCvmeiUFLG9sVFcxjSAhVpyCdrxqnQ86iDqL3P3HrVVO6jjqKSTl6ge99
KGQYZlCVkrqaLroA1IMkkds048tfkJmFika5awErW4eECJFJlikaroMNVXLtwCua3BmqVR6SBRRU
mhRT/r92/oZNVqkOjnBhyOG+H6fu597RVO9QLRy/Id+G+RT+lJ5JmulG71frq9Qmm1+ACEeeuBGi
48NyUKmE//HJIuXTwBI1eRZcdUtchbwdGlg5VWXJrJsTEv0mgBzfokf0xXRaJ27CZHnecpMnz8jQ
XhzfLGu3ZGyLILLs2oB2GOpaTfC0zW28uiLz04h0xWfLVLoat+RWpYc5DohqKIblSNlbrcmSfjqT
3lg42iBfTkfZzoHDttq9eqANiPokqeTwxE+xX11kIzAWVD7kpGcFvcZWqL00j1B7c6hXzmQjMa/u
qNn+ZaKEpulq4Hcz98q4qkh6JrSUxRE+qPwoE+G3Mug8Hg3dZ/B407+VwC0iNeWlu+IirzxQJCo3
WM+IBSuJncBxCVSzJAp8ZKpG7VDXkD4QFsaIocdwdD5nRPFO+4OtUomB6qp5XwueX6IozVR2byWM
ugc/Vndtw694aYT+tL6UMNjdpoTtA8h6rnSzGfe6sJz7VNJQYJKw0WnVp6b0timHN1KsEQ950fCO
wokVgA6Spx82RArSN7BQPZskrknfclw8Eu0D/HWbm/9nsp4IfZ8iZrAYgVHJ2i5hMFalJY7AjAE8
HOuBTo2MkyTKlotQT67V6gNrqa99Ol3nOX8tvHf6cgMGSjuVExBEeoTT3CZJ78IP52/b1otk0lY2
DXG83yJh2/OCRLhMY9gkGXmJto4gOYHWqi09jppodUNO+luWygXsTcQrOeY8G8zBeKHACchI3St8
KZmN+71Jt9zZbegnFLKqc4x382HbobKIOM2RJgZpPxkqoeyzztVd0lKCHd2weyafcoc3qayyLNJe
T8dLwCjCl5an/ttoMO6UN+fxLNcVnzaMAP2wBO+uWLJ58PHt3ZOBPdJ7ItfiNfy27Bi8QrtcI2GZ
3FS5l3gA3eOw11NNUsOnj41dVGz/IKlQSFTMWTI5G1skQmrGI4gwq4XbA6ucsrnxSCPvaKaRjwIg
boMrpK2yqb+P0WsDg4NvcDDvZC3L66iZ5OBq1lWvIjaChzaIToenod0hz2At0dNRp2hoDaI2MtK9
IXS/Bsgux8Y+L5PTCF3PtSC/7H2S8EIvi0VE2i39Q83xteK/p5mD4H1bpKxAeUZ1YrWP04LxODIB
XsW+NtQXij786XZpGSsoKSyPlXlz2LDJKSbf6RJA7SNu6SB1Hz01Z184ldhRaalR3MnWNyboPaFM
M2/NTcTk8bYk1lfNFgELZcCN2Adk+559EhHqMBX5N0Zk+HwWmq1iSB/dEysx5G0+ETygvO4Grdvm
qUalGgCe+gmYk29j6n2i6kZNYNGcWnvOHtE0BOnlE62ReZtLIHhpxTVS1SJJvosw3KxUw3bZBBoQ
HsVNxOm8gaz+fYJYF+5t0MkASxN3Wkodi7v0V2bxpep/7IQ53oZLUGGy80BL+puXIveo6Ky0dGy/
l2dONeWsZvkEoHJ0tIDQGHn4s3R7y1I5MIiXocVYwW1DBH/1ag7wKNwsPMS61C1MzxsbPOhiXuo+
9Bh7yFYpWFwf0x4NrZw5MopvMecS1Y097xSSKD20N+K+00wqU/8Tbxd9z23nSIEY22PN91U3XEW2
XtDi2UfrMS/RQcqhiaVL/ljpRqlRzdp7jVzGgDXMg6a1kfL5G2FEzvzdr5hHB/92g+KU3f8sJwzv
mOq9XoM1Mewn2QBCrkHTBFSXUhoiFmtfxspCKD3Wqo3+CgRSqXva9FymBeYy59kfdJ4Rm7nPSGp8
JaFh7aOwnxYezd6fU9bAuw4d+Dl1xdb5iOHkDAHDiCvfmn5LyYFN8Ycuu6MZdz7eQ3vv4niEkmZo
jc/fOM2bJuk8My9MFuzffnixi25hV8BmjlwoX7ndnxXMRmTIBp4uNELP8488PjdoRG8lBdmxdGVv
eU8G0RKU4y/h2UGEMeieY9BBHdunbSrmFpwokfaZblR+WzDebLywAUaP+nyJiol0JNtn/DCjOwZW
b2z3b+VA/+I3x9HOOGywh79owtRg9ZD0QxWIIpnSa5tFLadsjASw/PLv/AyZixKHU36mTWY3PZXT
Dw19UPSe4hjx4sDhoVWvU3aHqHxKu82gp7niYiYbZ73tYJMkfy0mWHZQ9MebT9w9fWlCmsWJn0eN
y5n0NwQBy2E3RWEGDA5qr9rqCLo3wvfpjFLipGC+esotUiEG92srLvFeJIbhuBcJxcRVn8qj/x4E
eIbQcvR2aTGc+jNwG9x1onMQu81BIn6KKyDzc4tVDkqnpS8ygMb5yDsmpZznOJe/eNqgbU9p8y6U
kPtsgiclvWamDTtLkaMJfNa66IGoQNZbWsYxYLraqbi4+zK3uP8vQeCfJqrCUozyvz9ajn/Nx0Ta
XgMSVWgu6wZ/sPwOwV5Du/HVU/P2pH//jhBKMbl2gmadVrduC31+RPBLiv1BcCW6U9qlhKUV4uVU
uxLOPvFMp80RRXATuGVWPSAGflykulQh9+442BGl6jx86GYMhrBZbRHINy13gxsg42IGJrcpsbxr
YC5jLPgzNklFezmYlD1UZMz3BHMyZJCrEO+qtM4tymFhKQqMFc6uq1JlIs+dntWLGhZAEesWZ/Fr
UAOYyVLyuC17R6YhVhdAXvmGbpMDAcBhVMJRJnoVfU3mA8cAij1sRtCzLa3ZLf+8lXPyjlgpqLrK
Byqe9RQ0zFqOM2jPbDrfvxuBMIJ1pZPiMRPzEcUV8j3nWXj3GipKvVKQKTO3hE2WAQUBoPprwdlX
5ggpOwGeWE8Ea9yvpcNs6D4Agaiz+blsjHgm4trFdyZom28oiZu2eEI4ch2kOmvjx0yXqaxPS3hB
hd65sNYX70IUutXIicNe1RWoG2AiMFWZZ5aMr0EolqMv/IDOjm+pYczPn54jXQEgfAa+bH2kfwAA
7hzyOpnM/l7NXQ13T0hkbVW+M85wFz3YwC+yKBGNxWwe5EM8Nc3zaKNcCQpVJGxvw9SsG3094VWb
DZGK1lA3I0NyA4b/8y1tWxVk2hcVyT4e5r7v2iimOg+EJ/lYIryeIN9xYyMiAxFQw6hp0cQbMtvZ
evmKYOf+xuOXCYA91PGmiThUgjlrjYTIpQMtLT1FAijzl1Uski5zycZPOCn+fN2SmwFClvb+S0RO
vsTPWiJYOpuT+pON5LJT37aB3xGRfbuYK/ZvgBPV3N8BhTpqM+imp4lcGYWf4dJUC2ho/dwhIjyB
bBaJZQEl4r3bGCufZRvrypfE4Z8pvMUAJyl4UDsqw3cPN5QV7SWNCLNI15Uz/gNinSK431b6kw51
CfoiaKWp65Ei0MrUXtQOxgOhSOY2SbG+8J52z7nFBV+tSdbTPYIuevJOA8LfRUFODfWv1ieg1+FT
NB5ZL4Faz4ncgZP1DotVPazRX/9e2QCvua+APg8Ov7EhOavOvLDq58JRH5dXxEzB+5cV3e5M4efc
S3QAKrw7bUQ6vD1vX7JhlDCGueFY36a4A0dYzyO9kjEmccodAOcOhdjdWiZTjBTB6G/lofSUl3HY
7JkZf2cpro82Dr5qMXtvwf2y0bLAheIaZ2K/ytC/oN8tSizQ+la2rw/HpywDM/OCe0rTrVZg8Eib
Ew8QuwJZKHHfwqZyeN9kr1piNp1JvULquR/w7meyJdOedKr0d8ogkvL4uN8DYv9nFifDO3OYQo11
1q6E17gdcTwSNTXji8yYm0rs/nXJSqrJJ8RCi/gvI0dkO/SvhXfJtGIWHxLjbuIJFE67KHuXhMYf
w+VnN73tsCK1IRZz7iXzD/PDhc30w5ZAeeqNttiWDlICf8aqCWHKh64MdEHsjgEq+dio/Y5oNG1W
KgKIfwa2xeNmJv3E1O7fb6Qj9RkDGojkhQOOXwl7KoEq+fU4C4zQ5Z+zLEyDoFRZgdViHxp56LlN
JS3SChnJQkaPi7kPXV66ES9osd78WtozH/v5bQH9upx6qYqZsyU44QI9Js6W2cQqPYSoiymGQ0Lk
pIB9XhnWqre1XSxXLULgN02NSqg8eGIw1bwagfHlGtUXd08M3T+vIT9Ftzex81zvzQBk12J63H1x
wOgDlOsWc2ueuIJu/L+8BdrB6MGtNY9PucDBXpw9l6TZ97LxG7aWbpGXvZlxMW2VVroOEEwBTrqP
7Mks+k9aBupMtoEK6CPPbanJx2N3emGQ4DtEkZQDwUBjjzZL+16nx57UvFkin1K7UeaUOW/3EPUd
C7uWkzyRd29or59XrZN31U2omJuRSJX6zOhaCRy0qt0uqLEBa03UO1OUYEaw2FpI0D91TCdIJFV9
e4bJwTEQl8GZc7lbFlGxD75P/YGzpd1j5ITPtl+Q92Ybft0ZyfY/DT0l7AxdpECcEQJ56Jq3i/dQ
mXInvdcDj3tWuEdE55ymQ/jbimVgrmV5QHgg7f2Nx5dar5y6Pr5/QuIsn3MS9McruDauJ8WWaIt5
yv0A57TOvltB15CRqbdDEnodb57qzTrkb95uRrrWLpD6MWIGRK1xeK/OkR6Xw96cHEyrxYeWS16b
Qmv2opH0REgWVzjzszzgD++t4UFE0dc6mkOXMjd6j3XXq5R/DEppBvmDD5zsb4lUPf+zwshvaKnQ
UelrScg6MokNbktDTeDjIMh7xEjrbL7tnd1vEYPasXw03Pp0Hmn+F63829mn02PsHhWZaLbqjTH7
Y33op+MGCYlypkjdGGspxYi5IteZfff8aTXUmwSlNnn0wp5P26AlNFV57t59L8pUs4mpj/iWaHXq
h3BrLMQ8dWOD2ksPcNUpphkPvBXJ3A/l6t/XgNo3PS1LzhFxwV/O4TX365fLmDkqVMzhUSW4afrl
w0WBWHyGw45mEPaL+lQt0KNpyr3JB778eLGAMKGaHiWSdQJuaCO9qd+mCxUQh2beDHH+cgsaTStX
vzqJjD0QRIse7/ctFb9kNyMyQAdkleA//fCKKFgImntJgZy+UFmv8QtX6n7vnhkAIGvEw1YWLF0N
L91rMUP//jIDsgtLJR50OYgRXuaZnDKRaOdkRQq2PIMhW8FGn7/AGQyKbldXNZ8+XmSq750uO4fO
jrTDz3rY7t6l3hwgV/bMSoJ0upIebf7NIxXt1TUD122uZ9GVCFQCPDYnWHiQA6/feFaHZvI30bE7
uO6EK9ZVpib01Kzhg5JRF0B8Hd0bRcY+ZABoU+eN0KwldQoYUlrNzgzizxLF2gIcAWFIYnamC6hN
PRgbeXIQsLnKVW27yz7N2s0/3q5bAz3wO4byFK17zr011QVw2bAhiOmxNi20/p8O0kU+7aJxZ6Yh
4RSF2f0raDXia2oAaHZ6Xb9CMnvYeMLKwRzZ4pSCDov8tyRIrMwVqXY2XkbrnsVEhrbT9StfBYF7
D1tp2TmaWuGVcjg/hPzxia7q7lUOOec9S8oG5tR6/121g/zVrNb0xfGwZC02d0OBWKhePd73AMw/
lzqZ3cvra8hs+w3qJnI3kwu2zPgL56w7iPZWj0diHse6DoE0PVa7vyYyifYtgBxEZVOZ5iggvBBa
bM2rrjP9VWEvIB6wFyHHDz7jEL/3NgdzZ2UrrNkPHMEl3fBivBGOclGPeNVrTKABo2hMrymjCK67
ceGqnVIgguFHMDE+cT7+s7TpNcEJksrfWM4ireCn+FJfA++cboxXieAPNw/RRX3zAMqIlfZo6Scw
MF/x6VLcfKreFYxmDPx1KlEofEsmI9d6GHQMNZNxKHy1052BO5rxQSFbUHWYp8eDup6jk/BGW45R
WZPL9HxkQ6GSh4wu6Z+gjIrE0RRqR/hQgZE+cU0buqrfARfJcdrKO9QfVOFQsHVQ1LhL7oivDYoA
lxO+WOM6F4lKBmrZs59oGIooGI7ihm4xyAs8c4MCQXci65CLlBj8nT24vuvcHpOalgEgXCsRr3pk
YUSwkgWYMs/bi5GLqOfONTZBQNWHcvnJ1mq4s2Zd5ddMqLOVdCojxVTf+BtmPhU0emzd7yHT5+c7
t+qE43NYD2BkYI5KqIe/IJN1fWvWKRQphfYBTZ/47io1qA90vw0SkEQEvP5CSaQaUV4xCI8yNkB8
K769v7Xs/BseTf5GgLzPLy+bnZ8tJ16igV0/cIVYO5tnOvDicKyVwcculVdd3IJp+s3HJLw8uiIb
bZw9C2v/JnPG3BsLl4P9oaUVdJCATY72O3E8/oDM1CyEUMQeLi43E1dPQGiPrDO49qmkaG7nMXLh
6/lmMrceF8f41tRdMNgSglUusPpWZMB/z4rzR8gxTGk5gJgjZ2aQDYEZC60bLix6rJRQ9rUqzXim
RCb0Q+Q54KLlBd+TsShp0ruOjZvonpj0Stf5fBACxjHjpWYmcXFNQrctfL7Wyza/qkdnpvQ6yF1Z
uJWTRfL4tllwtCt1pIzUoJ4LCFHRa+4rYXUUj7UHKxrcd8cUt4pYDg212dwyeoN9z5ldHklAtifR
heJxP7Mzre8KNoaBZ4yOJh+QaqDjZt7lHMsEwTuzhkPJn2DPsp7PKxB08vrH8Rh01c10jCsqQt8w
CF+CITcVYPc2IX3cVsuUjoJdvxLJHOtAR5WFYZEB+QvDAXOa9iC+TGEa3OVxhxYeo/wSBPASzbB6
RorpFGKA1UIOgFmuKBlkhk/bAqYFPNSuzLAkIMcwxKJIrDeAt4I7s6qv+ru5YxFzpXXCIhdJ+XFk
lxvZ05PN6HadKaRKdkq5eDNCV8mXUJPz0/Ti7Ei7NsJqlnt2Pvk9TBevkm8D23wATcemVYZQZLZN
grXnULei0NN7yJd+Yc39PZpjFXd7GhT7jp5EiYlOn2bjYfZ9eUbDMGiPp33XYXhqV+O7UL3ms7b2
Qop03RXgXeT7Fl51Cxwyai/0aYcVV+NDXYkAFtZzlII+KPl3N0ft6/QszIZY9KaDU3eEe2N/INXY
ptGun5Ei7se+/b9BijEQXvJNU1/7kxVELOE6lpWBqMERzWuKYYZuvF2yk1jycbB04cFApDv71OBA
NvUi4Wa9hfaAKrWpB0vQG20wicbXDGrgxZuurlkRrz9/cCYFIPty54hIL9htVTtGAVZU15ynF6Gr
6YNGAfNkTkNiUq4vCYorgOikHsYo0PyhuL8I/nZEL57PkjeyWP94BVfKiwpyMof03C2zlEMXSnQe
t7/IyM5WGX7+oTQspwmrnXFEeRf9OvelZ9xPXAYIrOvgH7BLhfUQnzYh2Q3/cnHgDqfSPgzy+dJj
7EM+fYg3kXqA8oYYKxHavt/Qdlq6S3k63DzTCZuPsr6mmkexaHJ2hjvhuszH9TWFzIQM9mcDHGdU
2GS1p7fhLuRlzQ+tUZdtHWCeldANCDR+IrEqtV38ZZLwL+I4A6p7HBOwX91o94MQKhaeZh349GPu
16D8/LXDM8+nUT0u/kr6N4XEpyJ4vASntPlxlb2tBdSr5E66/P5fSwnb8xjwL1XcHBXqynzmnZwe
5IbGqpe8tIZvQwzqluvapdTTnZeVT4R5kVJjeqw5kfij48KJTlb5tdmz6V4XPTOQ+NUINKaeYfho
cGKnl+2Y9Lzj+BEgzTyJzni9xpKJpxuSzuFl/95dvznFF5eYDvQSySHcQt8dM0vqFm1YtyLFO3yl
P+6hNJP3hG0u7nwc7Ddts32XV01bNhotrVQUY6c7OruC6Yl4AJTrwXmAZN/fe9Qe5tnFyG5p3p1Z
o/RG3J1G6fqF2O6r8sfGgLhYZA1MkHi7NXgil0tHxtlgBmvy3uoe1pRIPMNuJ3Irg10irbI5KNWh
KkSPty9+x0H4bIX9loxtRmYzdWSREEhd17JzgZeMxyNh7gDdTpIk2+VqpzdlccHFpgdC+udtldqK
hcU8lTm+a0kPyRZ0hwR5xdDjTgKVy9G3DH0buHwDe3bg9cShI7u1SpOLOcwVI7YU+y3hDPrtu/I4
ppW3d61CJtAV59njQFqv0F0R5J/r5ldhgmlyHmHUCMeR64GJN9YTPzqqNaglQKzYwWlIy9pnDjCp
vx/3mFLuYPXc65BtmJFSlV/K6bvQsKhxiISSxEbxFFrwgOe1+MD0yREidgi+xdp41Ty4R3K2JnbC
3HGQmYzrxsuSitV5Q7Ic+/fOpb3U23YKcF+wOQixCk4nLZtAN1Iibf+EIM46VJgKGJFYzmCb4LG+
CwiSSeKlHjygcviD4Ip/+KdUvlm1eKYg9gc/XSFL2UaAb0Pr8m4pysJUWYcTZrYoMqxgb2AAmRmt
zHZ+5xIGpXxcBZRiQUH5RdlH6cgdbh1WZmnpAmlXX9X+zvUk4JiNytfPqVY7Q8Ndt8fChhjniCCr
eE6WRmQrRm4eZkUQ3hSDXmujbADqmGDrSKtVJSBb5qw8Rc9LR0gzT6e94qx7qw+EUoNCpf+rVwzE
r+iEzuy8/JTJQvX+hNh+jyI99Q7sYqVTFfgDe/eurl5obheSWDbQ/hy3YKAYMfk84Mo4Z3gbirLz
m+DKeD98eyfMvLO8iOl3THbn5gXCUPbi3fn5ogFHsqSL6IVqI34e7IitnLmbuoo03pADP56kjA9l
1eUiq1mXOBB4qMqVl880YG4l0JBqF9cSu+B22T6Y5cxRWmNRgrV6BXSIELuxB//vdMYF/URq4IgS
glaBkXcTl3wjd7kL758Kju9tv7lrPhPc28WJfELMDtXcmBJ5jcZ2MX58SZKYnxLwuwFr1LX/akQ+
03K6TlH+/4ynw3yBGGIsFQX2Vmfx1DMatj+BV5q28prMeDrcvqJgWoxVdryPD7AnET4N8ijVUSU7
zUgZ/zpq15iT3/7O28TCUu8DnGseHnxoSf1IQJL0qQ2tOuULx51JzMJ82B0NuNNwgNS81qgfZxh1
XEApaKnlK45ykWC+oxl0PGzJzd19iEQW8p5gtBvSjtweLQiFmlfICMDCbYEM5T89d1yRI1brzXvP
C3ZxH2c+SVpAuMRvjDo7SBRozv2gvTZG/1WnMZVgDCeoDy4NxPdIK8k0ykIbtkJ65B814hI2QkkJ
gZNxeqt1XaMtQUeBQyPHoYPRzqvlys8LpSoAXSPtoGShV64ZsYIkEmOvZZyo/391vfBnLRQ4XazI
q8zBZaCiU+WtHpOjUUM1BDTIvakrI8m5kDH0GwUY3GETgAxcbYGWnDJyy/pImomD5uQ3h6HN8cpk
Pv+hI8vGiB5XCSF/nNo4a86J2/R4a9fsVakrT3znQWEA/cydiRZW4CemcfwVi9wAVMglfAZiU5Co
cBhMIkrfmAC2lSTlizXs3jweYzHUKSpLZbImHAaB+WUDJLj1EepMjAyAb3KoqpydjkFZp527Ivac
xppTBeK00iYcP96ZUEBIJe0aECI2h1dE/y6N5eYc/vB739OXwfrDXGyipPdH/0fO79AE8yhWE/Hu
M8xHzXhqW0K9dVjhJtnpjt+zaQeOcq+znIDAUv3nFHQJ0UOzGHXjPL2/SqaDdeyUml1nQqro2cGW
VkL/P3K7CuHI1x0PRPsCalBeCFMBZrG0wmvC5eVHOKt0xfB6FLRrmiLMkJ1smf4dtpYBueoqmCpl
/dRCy6Jvrffc7LpV+i0G3tb5Um4K0XDG4QysRVnN+C0IrJ9FcdfFJWxATm98s9hzlxOXmab7j0dq
EAFyaKMYKe7IeOXI55XQ+xaJVauWzVLSKFBjPwZTiCn2Pj0TQIPufxCRl27760WEMId7pTFe+xBD
aTuxALaLmHluskOKC8DxwKs64RfpiKfApSHFycGmQ9JZA+AZPpummXbU56n57cp5G61xJ8tRhTuj
MFE/B4ge2jKQ49MlfHkcSzY3X3o92Rq+97MNgUXkROoLvmV9duFA1paAF/vpeG6ynRVaKLtHSfP1
wpLy4J0xhyejbyCIIFjLf9KvfaSs/McC+XQ88mGqooriFghbRq7JpjGBEJ962U+Y0srgaYEX8Mnr
+w/nglMK54XpaRJHuzgpYw3uIPEwL9X5fD6UtEtgXlR/FettuiZI8MyM0P9yeVIV/DYffm64dpYa
uc8cMqegJttIJ7DNxazVNpRIG+x0F+mee4pLm8SKvPMpGsk1KQJHWmAgED8Lmi1vVFJ6t7ZZR04U
GWFpyJ83kFPwySsgLV5Hy7RAhjOPGMWMM0YXr4IXwcw5Nut9LaAPHcS+TF80ce3azA7jzecSgcq+
Pd0fz5yFXKP4eJa6EaZiI5ceURiNyeGyrDAehdT+uEogpvmv143nPQffJCzGmmLvXTih4rTWEwWO
5xuVbcdYPFvH4hQGij1i6u9sNaNjuX33STmwlNPRpQImiJ3W9dzA2BXtqiBDTcWhB5t3DCV+De5R
qIkODPQ8sT+YmVnPsaUIThxLF4un7ZWLrj5RJ3UD0rcJMEsDCvqzqJqqXYGj5deRxPVOKyioiQnY
AfTs1ONbWN82UmuZ28CbtzWJLaDYmCqJxWFe4Ei+Und3kISCaA3TE3dpsO6cOR+de+eFSOr43BFn
5y/nQ4URePkPYSnTIWpAGOf52yHNxC4nHoF+7/c2q3aK4x36V/WdGKRI65VIKI2ce9Jaf0KATxJL
0EMUETPLVUS/a7ieJZxYhTP7oSwJmwPtlRaXkRZikiWEKm5WWtWOu+Z8+Q+2EyNX1uOK0IA/71qT
Mt9JTnEWlCKpAW3ibiba9Sc6oRpCbKIchqe1MNJwpW/3xpo/h/EpgKjyYzt8dUUYn/l5y1PU+jB4
FhqJ503vKL+Ydd+msSfhfNThaV0plilCVxKSJVzZ3ns3Y0IzmGbL/QPB4Olk8efcvK3/JovA87Ya
e5NmseJLN/HocQQIPNQVAKLy9wNEr4rZ99YWkhb7eHB9EVjih6HTeJUe786hFlHZ37qa/KLy5Dhz
/GkWU8yIaJJvQ5Nri9DO+OZO0J+KjQoP6NCDc+q/fNhU9u7OcJLyuMB/j5ZqeFWPTiyR+fySYP5q
2GxF1j3+gCvzCm62+bnaUew0BhKZI+a8Pf7+Qrqu3X5CfMO9yHejweMsGD7MrkKAX/6URg+XVdVC
BYk7puI7eqk2x/vUZQr380hGQJsTHbL9Cgf+bfNhzivO7GjiKEpFv8Hjvu17eIu8uz3FCLCrA60I
lvO/w1CLrOb3iUEkgPWtgmt5Lxg1QCNTjZrW4s2Wd5uj4xJt0mQUp7ErKYAz95VXIpcWwR9ajdBw
9gXmjvaogU9+KrOfVQCJVKTGhTlWSJJaAJksVDb47DOIJmz9ikmJH6L+oq88fFuwHy9nTFIHMdVm
bQqo3PLvH6A3ADizGTvOot4bnERkxtBUPtYBegJa4S3ai4mZHxpMYoPYUsV8j9HnNVcgtVsTF9wz
V/0YxY7nafAS3pl2GXgAk5d8ZLLUk5NLm+dYmg9HzAhpR+9tf03WzsH4G5wbfxmBEvIQHt4KWrW3
9PN+xAriYew67JpeACQQXwkjXmv4Kht/XqwHjNwFS5lVny0+fZIdHlqjMNWNtBmYUFNFL9s3mSMp
pRWe5xSTUgjzHMNEdul4DvODHJzYLpnM8lIr+c8j7uJC0BfIORzDfoMDAjWE1ROkezXcWYdAbM4y
Imnau1Tm6tPDbR4vjeXGdJoL0BF8yGiC7VZQPjZ7WK0enBfKsiN2jfWWQ2UCyKA9Bynvxc58ZF8h
5ADDj8v+YJBzFR5lRi1+G6j5Z+lxLk6ZuUJ+FIPeIvbKlN1P44Io9dvD7wgAmG5djcbovZYFqC1w
PVOT8IHdCfGHzaAvVVY2dYLyCSgWpNhGVpehLdfvMZnodVdRY3lD4Be9/QpyBafBbj9NGyT7xiqB
V28PU6PWT5kTedEAjd9PmjKn8hRx5i/Pzdh3BtRmCuzXd9y8o79LE/qJl9zcbH1z9Ko+fI7l5g0W
FbB4x0uMZXSlR1E1gdw4xKTibBUCWHKmDe6ZS8vYdsHTSXDzNIGGz4X/ItlddJ39BtqL2GhIEMIU
vVJEsfykn1w8gFiU2x9Xk/4VZiTEEEotLnAbTPmcT9tZrrhQlTvhrQWRs/Spm+kpsape8sUl8qij
QFsURIde2ZCkzBQxULLzmJjuAAuQzFEgOAamzbqsqK4xS/6Pkkl9p9dUTpMXrpMMcOELgYYO8EKd
JgxSyWuoeDXnFiDSZr4lO4MtsyZ0Ldbg0fuy3egqIcmaPuppiigQfSO3IAqdkxSoBMxNUQQ0q/Ov
dhw9azqSc3wSrsXDuflP/7BULErK7+A/W/T6E066y2IJ37h+4uXrYlQqPRsfcuyiQSZ8n1KIF1Mu
KFocIhS3KckjiVNu0OR9SJF4SjsaBEYG/5SSNa0NaiyyK6tZwBhIYmbmVKRnC7D8kNMTpLqLQhCC
+lLvjAKD3XeMSpRmcjwfODBNEIp4S1wql0RYgKO0S05MFhJhorFmVsi7vMgmoX5S+42tGNdKT2oV
8qJ2+43R1PZKc16R38chulkg0QoC37acb8L7u5wwQ/AEYgq+gPIwbGro0Ssd4vCiwd35Hv2hIzMG
ThLu4MDkM8qS3s54v3leOtNGBLRdihG0wEktq43ITwaUWoIDVQiwjDVVgQC+TOkG1JaW4OUfF0XI
Xe7jPdHkI9tkDjhttkxsmCrhAv/qMcEANNXJXfKSNt8IVZYRvX2lXmUHdFJ59fGiNzL15jt3DJ7S
24RuJptux1D/9rXBjfWj1pjQtyQyR73xDsJQA0d+skQlErqHMqDiHRBIws/gWtq3Z713oNUMdkWw
NKXFCr7qOKxYTjdMr/WYf2LYI4//kQRqUoe2QbZjJUMQTGDjwYryTtSyvEW2BnVJSgoWoIUni/6I
TSVyhTEUQeytktlp2G+r0pJdB8ttJTuFcNGXz+ZCPbW7MOTKZ0AXHLqJ/yjXr/mSCxD2KUJYUtn2
3hJj1u2oeYiyApEZZeatVJkSTabiW3m8c9XC79a5N25bvmKLKU9XszXRw82Sf2gxphPQcwGReeTA
tPOru7l9+CXX+QM8v67Hb3BYDRLZKG9CL3aka1fTrhKQSf/mHAIyOLyj7YlnjPyLaoaSrd/fO5RM
y735u7CbWra62/emoiW0CntJcjC/VUsSlL/o9q96L3O8Qp99kn1UydAgsYgYIAspzhxiZwD3Y6dq
y1/jVmirepfZjbkXhsJ9TDJkFEgnxQVLtSZ+ilPKc2ZWkMsI8MMYQY5B1bKYJpvaixQohWgCxzwp
II/iKvM0B8Nsc41JAoEbzsvGU1fgUFm8IXvJkKGdPQYTLwhYRf4ygffSe6LeWkM+kGybeDIgt0iw
fA0oYYh1K34mz5KJZFm/RTRxxyWvlOzdWVeEoATpNACJVxU+QnqDdc+3uOWmWx5SHCUWzKYTs2E0
PLZOSWl2Q39jSwcrHa2cyF0g9ajgHROnNBTO5l+EOcYVma8XHAzxjfHduSPdSqKbvNsHpJ7raZok
SzjJ/wtJ7b320j7cONcvtXw5NKjOAxuWfpKyXv8ocpRcg2w3xfstvk9gL1jd4xhRK57BRWBQAUQc
ZtOIiLoNO4LWZihfsmlIgYesMzX7F8/Ktnri953r/SKCNSHmEkUxFuGpwMG3K161zXCvS3MbHKMN
CIb3xpcu1dtcZsjDLqIWGNHYkEYMS9dasU/FnI4rL74nzWeiVNO+2x9T5AXeJ3gBLxzjth/idGt4
6XWLxcNSkmBFJPhKMq4WA/wgSD7O2x68QgDH7eMze1QzLmbAAmQn3HnufKWvlNYg2M8zFbG0YhDi
QVSOC5V9PXF4oNR74wILW21bWeCd4z5yyOX1rhm5UX4Z1kIcJ7wcsO7jPxvTY7m1vkqnDzOrguKr
8R5Oh9Kh9aoC1ekVe2Ck8mCuYKFUmCcxhiCB7FxXrxiL3ol+/zlnUXKmN1xbp5khc+Ok6KCi7BPC
wHAylqebSWoY+AF5Mk9ZXBkI1gp1xcRbbha+061P3sJT9ctj38eCabmyrfAuhlcAuqHnwX2EpF2q
+ymqjO5KFK4rTI3I1T3D5DA6pRLiysCRxYmn5I2Kaf626TbdRbA1ij9J/IRZxhTYfY+5zTtAUQKp
GJuoY1qJu5Giuf0bC/n/c/5Pg14ZxJi9zWdSNG/e9FFqr+9f1sACbqTkbVjaI7Lm9sTkkWym3zMX
aOhiBvARWxqDypF90CnyCZozU0+vDh0onQr0JGzxtzU049maR/+1aap2LZdihKtJ7306HBbuW8eZ
JzD/tiMh1ejueTjPfd9LpM/I1//8cEqDtMnysO/2btm9o6LoDMAmECObZkP3fugYDiyUEDa9amvm
PoNjlSoyHxyRaPVvieAIBrz5hLaAx2AHGOs/q/41hzsXwkBmT/Xo917XI/qcokNMFNtyBtJ5EwXW
JSFXUoVPgi8pWM2iFHxJMO4jb79JOFBF41vrRjtFRBTl3itfUbV9UTgd87/H+mbtSgm8XimbENy+
DeB+PA4zJowxXMvv0fHIU8Zgvy2DLuiHNaM+hNMo0cUg/ePo7WArHeJ9CToTqHS0rxdq3DBcpsa2
WXo4TfqeludTPgFcT/no+XRMtJNv9bvfB0gklS/gay+we7/mlnNB+QnqvlLf88m1dpK9hpCjdxww
EijgNFIrEYYU5/HOfDTW4O1EmCZbudmK2hQHI/Myjs8UxDhwwblMpGe+3aJWh02YIL3agsqZrI14
ptnsScdUmJCW4YVYFJvmJPHHQVt2NIWgFzG0oDY4VTFchp6cK9MBiR0LCNjHZ1ftwgxo1GOUntSG
ZR5GGVbQqzHWRAyKVOauktxMT9C3q66O47VNGmFvgaKM3HnMj5TsWLEXCWwLPjpWjICDKG0MSOnv
eTvAsMjWycl4cUilzo6FJtSb/KPirRaR5hpDR7MNBFsP125Jt+y48YePvDrA0O77t0clCRGHqVI8
RwaZQ8RcW0juZ0iXCeD0hyMHGHaoRHMpp6U/lLxCUH1EZ8xmvRqLrfvDoACE500p/xj6p5NDcMZz
4UffZYFrewGR9pHypVKyptcdHLWlCx6KJM1IxxygJp5pLvx2adh4vciBzZ4SSm2Q13fKD+iN6/Q/
HEfsxDffNZWzTWyJWpQVnYFUplBTiujcQ/cMYgWw8lR9o1SI4mYdRt2O3CxEJqGbjIMuGa0v/QWU
haWGcsjXNdF4pqkaQsJI5cV78PUFSIsIysMk3oMNkdjzRWa538xqTR4DefKsiR73qlwp4olWK4n0
JITOyYO/O6kBwWpJrKv1gGGIUimV+JPZt3NAiJrjJZw9prTvfupxwXlDN1DUhdqvx4vmMdXkS+Ec
yYarJ6r9WxB7bQzKyizAdHJDBBP0x+nx2hYdZF4KGAO9lEjEcpUfv5owk6l6R4yPRPB3AV7sR5CY
djgodAkb4TDidn/UTUlqs9JrDlTbqSgM5dpzyWHey7KaOO08K9eUV/LDjqQqrC3T/sLobHYSOMeu
RhGryUImw2XNAy90NQMirYuqSkN5voWKtBpqfrZdtWbVQl0olXZurHl50kAvgl7clM6G0Gi7T9Nr
6e+P4o7AzI1NU10fD3CW49td8trRRfnFrgFI0+ac7Cm7F8GZFwROet7XQVmt0LMfBMIhUkRUTUlj
oOg3O3pFqU6nYfvJ+7MZjIkd0Bp4n0h6Gfr0rOmorEMoqsME26CStUQtNKik3gXYgZv6Q9MgkaMR
6yso80LNCxC97h2RmE8K7iVWqf6ZvLPQOIZAihu7zsQ2+Gb0jpSYfHTiHBENEpGr8fqq4QsbM1Dh
F4aWnrSazxq3V5LwLp8mXY4M5qFKjOA6PjyNCzLYzoILM0xZyOozKJwJYsW29syGoRYl8Ya1Cmor
JLTRzOcsoP55Em3+2AvFJVoEW2Fk+xIPxSOUSmkVZTvE9nk6Hti81U24zQuiMV8osQCkvbVt82AW
dVM/9YN7z74/b/gkK8v1v/Gx63RR+pwcEh1NJvey7/X1UPPF0zIL9KQXlitlgrMlWlVu3/aI3Eir
YTtJftiix6CwLsazmjr+FgMwmzeaS/rdbjAzzd8UV0zv5Ln6z/YyxNqZDCRxPZxtHR3BzGNfqGeM
w5IZAjUiF/YGXxxVweavovCjK2JImqysOuZLdM8s7yepgaGZXrb7TCF/7Kp8yr3AopRTQRYLguXP
T2l64bHf+CH/E2x2C3tYDaQyzdaYagsarxXtxZkyRRBDdAxvO4j1hlxG2I37s1iqzC0EQJrtCfGE
wccqc5BNqg+WEdvylI58U4FBA6T0w9yZCIZkYotUroV19YJkJuuCPv/vupEyoZ9Aydyq8+UuoH9H
OK1UzseziHU3Ko6jnRmgJook2S26PGIujrzQA6TxT5SrSYtCxgbhPxs8pppyYkRDujJh1fA+gGCD
SQ/BAkdnPNt/3pR7PwxlLkPHgj39M61BJ+GAVllGZP0YSVhlR99rcJyTUx/nLHb42wPRZ/PB3t3z
ElG8vMc9NBBTqMplqhNv+bB/2tI+ZPvRT3YaJV+xJmU/adGuWyUwuCOLBFP8lzbPbZeQ5gBsIPAZ
hb/CSZcKYetCUJcfc6qg6FqtqotheLjfwOWSatK1r+hc3foGHHH96YIM0xWU0w+x/xBgNIwnMW56
5IUOrOUkOtPBcNR+jrnL0MJ1mLK4oQ9O49Y7+RQB0ieDzJPvkibfPoKWTDVk8hpc5abd1ZBNRM+J
N0bhGYvjI8FmaSCjZmLBYuai5cY5pcB+x+/jMnRjHfgajEA3/GOZ2r/qgBUcdcjEeDwO1JVD9FKZ
8JMlySveioqc3OxPFg7jUqr2m67xkliU29JpUyKuTBIlPE8q/iMQ/vBy1w3YkIrqIjcF+y0o5g+4
A3/1h/d7/lHuECYDUqtxYwupDJy7u1gwOnascUx96TagHR2GpBaXCa/cC+SDIvBFxu9Vo+xf7w5j
mUz4LwUQXLgf0KmtwdRwowAYMre3KqElVh+EDymfueZUFun8fAmQ8Zfmh89Q/erFMAaZ//iN/L0D
ImD1Grsu3439yohFXQl+VItbk13LluTKiVurfj9w0skjEesHSPtmt8t8i/obStLLWZwvPSMDJ516
2pCbGvdObOZ3kOjBx6H5cc2A88iL8767sOolwBjaQrif7zqq3a1SvS8X1gF7H/1moZLnb3gBmfHl
FyTrmQHa5FmEXqK6TSUyK03MCz0fvH/szKkMJb35ZTrRleO6cEyRl2e8wT/96lCYT2emqkmpwYz9
W/uBVqdwoYpa9ev5eTLDqMWNA/VvlWKbPPOJ2DC59jiuALCy9yI600I0N6VXJuW4xhPczeOgzTmp
56VoEojGty746S3cDlbXjvmvzbsTo+LU6/uKEDGEfh5vH/p7jFt10mvNOPAdz2GJMyO59EwzxFPf
QsWJVBJ3gjQvv2Knf2JewtAOvEznsWgJJ6sNHjQwFNkTQwyOcqQHer/wCKCvhHz5Z7fAN1pqSuF8
XPK67D572AoTSwnGLwOZif+MrYLeGGftr7HehDJ6FWSRaWPWUwSNHggDYLRgc7q7lhQ2PGZFf/ii
5SjwaxQ+zWymjrMOzfkcA8P5JUnl8MmJQO2oprmOBMEZaEizap+A2PNVbcP5wzruRzmrW7fdVgF7
WX/jIYvuSIsH55PCPMLJyblaHVNEL2xNgb29CNFPOeD6SQLcinwosdQDdq1A1/U5016rI/m+ESyR
pkRQ0SEVrcoJlri9XEFMA0QYWYKD0/jmVzj5J9YrGXnWVkp6voMtPs9dx+wHKgjv86j1Z0A5Dut/
WVWcc+SmnEnDQw+qa5HIdU+nDf9iFoDQidWlUChLKM0V1VpePME5kVLp2vDcXGgdjpls6sdop/81
fwwCIviN/z2rj4lN54BIyrr+dyzlQZVSKFIX2ma9zyKdFH6zl5eya8ky/15fKZ3wjWG+l9xveQD4
ax706ZRR6XG6gAisp0Bu0h4gv30QXden4DDpnOn1b79A//c/S5TEpPDhevKtrm20JOL9niHB82Db
XsB9ErybFD6IyT58LVcYnDl3TdO2eOeYTWnHFRtkouuL26h2Ym7qDR8BLgugpQ5KTdt6vFDKB2iu
wUaefdoYaCVjgiuObg0Sn8cBfyTdUvAK6FswqrZYxs9iFB7gAG/rYZbjHXurhYTR2AI47ebPHXlN
TWF9rrBt5erHZy0u7loeLvVGCazsccJ14Z6uuws+411yu7n6kM2mlIxNB3u0+Z3KW+SwUsatNnjT
GSllHZJMv8E5i9PUKsa3bYGntaPkn6oGGv67MTbCH4S1xH1aflFvOmpWGmuTytpN5tBo6bEU9jp2
rW0uIAWORNhQoNO3F4Z8jd8FbyW7yXJyLf6atkCxkxuoDUrYhW+BTdLIRMvBIbQVo/7X1yw9LWJM
HzssfmtKBGGw7y5sChMpMhHg1UkqCG3b2Zmd2KQVAHAuyYvyntVozgNSqGLQz1PGJ60caWuJ37DH
xUy5tYHJ6V2fx7Xi9jV6aSLx6DrcAKIoRDuGXTGejI4qlu//s6T43fhvr+qfbb28wMFxkL9PHyPT
bpmWIXlbTrGqi33x8eLWVTgODH3A3wzGamTyozQRJeGNcWfyCmMZAx55O0XylO/Nn6fpNuB8fYkX
DlZ37rImBaZG0cUvrpELOI1V6v8ISPFlfg7k63zLNhj2WGPv5vAwCLKbZ4XeFzsfYk8k3jc1o+rQ
tYtesWDYsO12EGsaC4nVJECHxldmmHkSlKPrhpfP3PIDw4vIVWgHAVbXACbSFLyR2yBBycW9PPq6
xrHtGmPuleILRzyY/tDj2YVHZtUasooSphGYYaS23nFvZOdh0ICEzC/r9o6ma7BexnQ979g5ZUHR
l4IngdNtToyaUU+XS2spNa/SOIL8pSNGIGLUpOP2WOaAhcJMDKWAzUmFOz5/bwT2+9Kx8I6Rn/u7
PVAdF7605IRltnE6MpFCzOXyN6IMjP2tOoTvljWe8Z8fvOkGNeMfZO7LgI+CdjmrMHGaYhmLpSHY
EdXpWeHj/ib5/q6i6tAFLaCP9ezazt1GHeI+cGEFiu9XatDNmiUTnc1WhczLtfh4YEydKjGbjNsG
BlAEYiDkM5RDkzx0hOVU2HEjofs6MgSNoXRrHsLA91vtsG+7tuAN9k6KvrwuJHSjiInRWu8ky+/w
5bO2tCiDaxbQguTEZlKUVYwSHakgVBGS8yccbq+q4hGJEyldr/lwXHLBFqEC++5Gju0CdJ4rAgol
o5QdSF9LU5y+hj3oB9G7PD/AKVA6dW/6HjnWRp6M6lk/4rO90d68F42G4t9uUTRGZDSeYfKnp798
Nlz3ERFhJ4gcs5RdNdQuXsOEdY9TszVPR7AOXGG4asvvxjE2X0g3GzCYR9S2oNI1hYtSDnuvULCN
kPLJ9ZcPeYns5pcNVwX43KSQ3NlD5o3sQm3LHhk1falSuDP5LScNakEnwPUHBxX05jNZ4TdGLXaS
0qe+X5M2e/rqcgkNrIxaYwXatv3VNqxA1HdZgJgyOuiJSMQTaJdU6N3qwFXlZ8xISLOMY8tiXuLP
walKPGV9nfxu4BqHPVQ35fMmf4LHpAwxHcrXIbmn1l9RbZ1//+QI8GDs5aYhiVPkDq/kXyxnvb+g
cKtGp/VElHQLX0nWjb6sswyJN6bqa4SvlQCUsU/+WuPJ0kD2VU0lMwTUYbM7HyaA7E8ryxoy8JSL
Rnb4t1B1RBxOM8K6Ar0rnbEo5Q+K+m6u2RtIMYmPm2Vgly3NvEuW2JhFjy7KPeDVn5kwAI21+bBX
Ner+R3aX31GnVbVXOFghU1La/rJVe3scpA+v5xwANvFb7ebNIn3cWf5dZ6Bc6XFvuDQkUTl37m0D
Ynuq+K4webwo0Rx3YQa17btd2gVmlcaWKwohPF5KcOA78uAjfkSxu9FBVdNlIAFrhzUGWHR/l8Vo
e87gy8oYlYG/SeCgKN4Wg7b3w/tjsZkg7J2hYhIxhmRqqWO86m1UVmtzUiXR4G7TflFl1nYvIULZ
QIArwQDssrU7lFKPJb3qKJEISasnJ85eWFZl0Go0eQb6977go07Iwu5DpWOs3zXPxLsZkd9kf4CD
e9kh6+/yFHQlATe2kOqVKxKR3AweDZwqTYy5mo0WJR2KMPZUfax5d3evP608IE9R0yQRuGTFkVLJ
6KQJ+lRJW+O6DNFYIxOcLAC/9g/eMMXWhylIXMnttcOaK7imOlWYqTbttRte1P1TTUsKnFZeXosj
xf2MF8fSgZUsrow+6U3zG1fGNYDX/Xyau8Oqgq3w5BzdSGXYbx2LUyrPCEC0/OGn+IGQfK9/LtMK
UbBGo10Kl0zdhxMRm7GyS7jmc4F9Dbn9fnitCWXI0rMrMcQav8o4t6TmSOnMZTmpfe3mIB07r4eC
e/aR9Dhvx6dg3GB+wD5UCJ3htz32EpT/L9QhWH8wt7HOmMmBJHh3NO6qAJGke/aHVwUWMTYGtS+x
AA4/WBGj21f3m4BWDe0TprZHVTS1Y/8khMuwOppD+gRpt0+E3RuUSya9v4tJsIYyVZtbnwveSDXI
h2OCLtxCM2jibD0Pvjwcx4BjXKeOHmkKHjx34OtsmE/8kuZ93kAV2QuMCheNmpPbj5dAeNg6NLbl
rWBvYSV35DxDLBxlnRvd/StEWfTnBG9QqtIUNfcwZl8Ndn2kehRFQvkKv3ZqHDh3A3jKL3k0Uagd
ZHFRfbsTgiuWajgRTnj3boWbyYYiz53xk1iSYYH4f2r32JUx2NfIla2gk5IkGvpM27A9o7uw/dMw
s8DFvQ4n8PAXnofjzhd2gWN9uddWsGW7cqj3x0I+CJbzfZ4ae/9sUjhvUO2FGhnrfv8HdKrcoFql
MnBNIBjvahdEQpL33wXHpcV7ufUohQSm2U9SzvQIm2n4YBD/BDBXMxv8958OYPXB3XsfZZq2x5+3
FzzyBnFiKFCch1v7R4XviwtSHWQAWOJybIh20Grxh1PwgfYbnfUJKMsdQoroM+4IOnyTVhQVuCwk
8CseWLPY5aNj73l80Npi0AgJRG8EtNeDz4XT5xVXzOYdzguGKmss70G3Y+O4LyI2S+c+e2YWRc43
aE9mAgGFx2JSSp51j86vUHDKOEeZi8filJ+xzIToKV/2kdoROfpe01ZpbBHGPZ1vwDii0FlBxEgs
losB+P0Ji9hVxyS4SVLn9YqKzYENdeJGovGY0tdxKBm0Y+i307dKx/aQTpL2/zZlQQNKj2F/MsGW
dRYByU61SSgGXGrCRnJgmHCMxeshiGt1pEMCLGV7Wtut/RJZKwaXSrFRfRK8XWGYuOzUkN2Ylryv
36khZRKDGu/X5XAM+HynI2KLvRQ8A1g0j9h00bQSSvDagpDT9V/HGGZn3XGJvDbpEe/MdUGyTA9q
La4nPwt8NAyCYEp+fPN2ZQeynVss11ZD543jSPNfNO6xzJ5+1D2JgoV0qm0P+tx+jPQJuQPUsLIr
qzNQyJwYUmwNW7prBSMWHfbkFeGYOKZXeO94slEeK3kQGofHQGv6vcfKvPb6AfVnyR3BYkDpm3Fp
csSU2ygoo9JipQuYmUGVa7jkWC69QljhLS9oy6uTXf18zlta5t0M0k3XJmkEQCPED0TCKaKJJjvS
QC9ApXA8AV/+hfCcG9PZx102SGnRGK4s4rBzfDu7AtyQwXGPBxTRQchhutq/D96xDV2juDFeglfj
Imof9m0oBL6r8DMn1OQYrCiW4ue0UZAHqBAt9lQu+v+z0cyVY6URSWFNjRC0fQUHypqu4pbFmsCN
xokb6Ba/cxVEJzTgjh7Fqv6dHsGlP0I7Dk/BeOR5cqFWMdnJ4ErNwtsZEwnS85y2z/qsuASL1REB
VoWomMBezcx+MBtaUgBnRLyDuaTRfRdmsBJZVMaW5j/StBQCacCHyrZhgfhx+vibxODRs+afSa1i
nMfVMHqz7I3uIG/x0hCgsm7CPjM8y9V+k+QpG2a3MbVH3JB1b4mVo5jboWmTZXLfTTElc1Bxaoe5
2+EzUN2NpX3m0pnf/pBTywwdy0nS17Xp2XLvVEHJ1Hat2cLLjAqX1EJIC/dReObufdSiLalOM5SG
6Hlr6kLrffoW57rNuHaeFJSHOIb9r+5j27KnAFsoFNjSeckYRG5C6AAyGmdBuOpb5Gls9jbDGE18
/0Z0sJFLVQ6LLYHokqKYp5kvtgtZVDJmOtRAqTqSHX57uE8OJE4LhntOXY7S261TJgFKTJdi5hh0
4EhlwtwspB7D7cAsJTqeutmgvStXLZ58xbewTFb7W/lZBO6+N3BqsusEEdq+jK3qO2Vn8fiI8iy3
fUj8sQJx1QQN+pxsZQe7vwY0U5/5/0t6aSJsVRypmBBHXIOOdnsNlR/a10g/PhH4jxEiOb/jkRms
Np4yBu80qPcrI+458T9a6ShFJX5O1XMujnt5+itX1wdTMbnE2O2rv1F2wnmYTKyB+0te1UNAOR30
38pb34keqR2sQcA8Mfldj8mcKqEQnySf7SE2Zr52RaYNqc7uzdb1dCGmZErnY1ZI7EjNnldbRizs
oJjnDIutXNAj8LrM2a1tpPCZE2qInJG1JE2SKFcAtRKflCqV0aHABhoPBWIfhuJmAiyghZv5DHRJ
Y/r1jMhb84WzEsBbMyHDEp+QHDM94LarxwcDlgxZUfa6qrxinakZWGaAkDTl/eOhUxTYO3ZJa1Fh
7p/8GasqWUBeAdK7c0B6//8pFdhZ4T0d5S3d//z9C1ZywZS0Z/rd3yh56UHwxV1xyI1RB7E17Hbu
cXOWW9ct9tsTwr/LMNcnCvRq+OlbuCkPFAw9tdSllFPAeV0q72JxwmhAwVg7joTWQbJXTJPQCse9
DeBUvDoOUrzVIhnREC6YhVJXHaAt0OcjLeONp63zJ///gNzn8M869Dr+gyZwyyze3Yl5axZK4UuD
8sqYELm+ip+R4KSBOobl2T/L3q29yeDlrX43VhL2+LuuWP6uByruusyIw2v+RjnRtaMisbKKhutG
EbYGTk1GXuYCyhKAeXjShxBH0mHvv0EXLSKqBogvdPXCXIJEw5+3IX3t2s9P9d4OdcTccWXMO+Kp
YDZokasltJExkxE3hcdV6bW8TOQp6qiPjN9cdx8X/ZGD+s0Xdfz8jCmQSuLirX2mnL+NHIpQ91ev
aZ4CaLuN2QN+UtWEusAcFg+oBVnIfNMyXfprcGJtznG6aAGLiVaRppVWKEEqjnSgPGTOK3dlAOal
Mz+z1UNLvxv7xQG7O1yejzICeO4PfgwOblVIilPooRtHS6X4gx0kCdcZ0HozxTScScFKedUeigHs
3neELpl46K8BJIW6O8J80gfkRXJrc83lh4dZv6FTyzegiNEqOXMKn0DkpjKWv2fA12r8A03wySiy
mshOtjsstFfs1s1N/WaRERjh8dua//A4q9BmyAb6mLUZaJimtPNAdozwnKYDYtIuwGwYxBrEHWFQ
yj6jxRmZuk2ACg5dmZoKDNkyFztgq3BPwha5cd7hg69Ao99YJr6uU0tzb9eb2HpLbSlRHTQ1/zeV
VFC606qcc+dbSdzBHy2MXHbcEcI6b2J1zKVxGDox6GkylKBZ+d9X0u1ZztX5qd2141xquNFJlfGg
9AuTith8rfMhimhv/z4uPppn30JkZpU9WXX4c/0mJOxpH9zF+fudLQH2+EecnLP+xgUyZ4wZv/Ko
IF8w75cw5iT1ZC6XVws8ncnTMW+tauYznN1KO2rc6CQDsfOGQvkv0Jy0TxbdivdoztCsEaOaAGrV
9l+XOU60xDaJmiaVyPdbwpcofTB2WuO+V0wZwvSTq6uQFQtJaGXmZ+hKp66usefstaglnbnzKJLw
r32tPubHaS2g5c6gPGjfrwIKi8EjPXLZDs+rbhNlbMdbXZTLZGlHHNxNP9TQraJ9ZnGFQYyGb30V
4tvHvpieHb7648FZ93GXdzro3D2kkzBUlwSG/4hl8nNhmf4CluounjCBciW9cSY9wdSJ8EdP97kF
hS7CTIUtukKGif6OjNtAmQp7u4ZwF7fP/MHvrjus2jt7citNCfYwPvoHiqZT9DGRld7fvl+z1Rl1
QfYlJl7ftIZPbPMTQnYbyTD6pjwFkPngVedU7+zDDnnt8+1nvEG8rz72or2IKUHS+zvabgSpJRL0
4DCwcuBv7Cz0vobOZqLeMgw6JsRHKK8JbYJ4TPJUaTxeeK5HAwrHIV7I5RlBBa0Ufl/D+d1L4eFM
8y13JDYR5uzEVIkaG9BgO62x3iKuKBVhYQw3kMvtYAAW6FOrThOPSAQyR/zac/vc/xT1G9TVsa40
efBjwuLs/1X3GgVT/2eBaIPseSmUg9pGkCYhJmfkO0DCG+fpFT6c3YkGRqC7Cccb+RyLNNt6nRc6
8SUJg5Vp5BuTE3/KtIDq8PKMjFgIBcrvbY3h4sjeWIaH6uGclCDCg41mgkV4EDAggSQRhVsGaZhP
N/0cG4uBxebbO03d/KXUtsQP0MOf5zAi3Rps4bDwvY/hZoJlhrpVrYfy+qjPWW0oxQJLsEcstHBz
YRW8EH2ZVU5ERZuVL/A1qrVNPRwqHRTDSJpjHGm5gkXDEqOlIGCfZAyQHi74jK6KpdZK05MezqH0
Kf5Qh3xTElANi6UbH+ZV+HLeOpHn8oWaZxyv8Onh7CRQz2ERwUHd6Scn/lvmwpm7grexjLRYer23
PYPE3RwGa9J2Y+UKLMuBfOLB2uL4ZV9m4GJfq8uPmt4L2Oiv7L11DZPsxbDtlw5thg65PSWOm7xb
biQLv/oIgIQBKcPP/4/WPdObJbhnJIoIYIbPJjIfSDdAIRMwD4qRewZYa1QvZ4tT8TKW6qPyQk2z
7bWsMunYWkVbExTrmz91yanz+E430ywq+QwIEEopLgPBXHTdNp5sPwmJTlvifPAznO9OrJLrCaUT
E0xqrGbLZRENgMvLndFgMC+/a8lrNhvJdPTnclPBF651LjFL9/7BkeojH86GunKGd2L0kjcXXLul
rxgseTfyYqmgHht0UqMS1utnqOmU8+LsS0fB0VOSDLKo+LMqielv69VsUoXLEAH/rBxeQaszXgzs
aYXthBsMXRq3v81OHhN8YHtpBK5ipX7P7/ddd3tyuL4OHZvXa5FyDVizHj27jW7yaSPDjt8A+70V
T2g16hQqUSJQcUX2yXgNKxY4cyutN5wM/avrIUVq4ajUaQJcKroDfuaeJLgfAHY1X3JjNlyqFQHn
JG9EWBApb0s6khSDthwe6NGQGMGf8wZwWoaU7zfE2TxQ0ocermL6cqPzUxhz+jOOjXH7s2VtGdHd
+WWbL9mpfrpT7wuEOwaUhGf+mH8auAuk1KnlR897XbjSfEzeF2NDKY/1ZzjODQ2impTnvjYbHCyN
LV/lc3vAV65qmXQmCHGkCl3tUd7fQ9AjmssMMBgRHSx35k4fvL4vZP6LI2jx/W3XQbf+AdkNpyXp
EySYG8m87gOYCDYS5dlFCnZq71PzQb1AMJhfNqOhSCvExDSEQlTCgOSLZdqRQ7vdMycnUpHdd1O4
HctX1a7rugccFdzc2bQsxWddfF7P3FbQebNTDm40q06MuUPBJC2t77IfQN9J8kMqJz87STSn8XX3
Nb3rU5hgJiZLz/MGA3RHhMJYIXTwXvZy6KQOQ1KGffbphSsmM/gDRL77OQhzuuk/ntUTZ9zNcp/f
plLUzjs/AbvZdluKe7PTLcbPMPrLfDiaCH0FJWmcG0t5td1IphiwpcZNXq4vBwYIZEZzoa3AfQ+b
h7tGri83aQ5x+wlS+/Y6IWGWwI8Qe52p40fT0Mi21LRwIdyo77KgW/jDJeVGu6+WaZyFRg5aQvpM
OsxL79kKnjXhEJDMSwoHSE1wVPynSgVRO/E2PhHc3Oni/0aAU5DlAahK46ggg+L31JUcb2Hd2KK0
mKz1XbWpaynVw/OqM/HpML0HJdEDhwIWgSbROhtVOwOpcZFmmIdcXD2+RFzSJHAvLIgDt9TW3Dfz
HuhGU0bbHmNK8utHfUPOD6vRjiUj6pozzq5QxdojKzdhbuUnhukNi1A9NGZ8Q3EdjAoBfXdr1loL
uf5yKZ91Ihr2RPSS4KxPXLgMIqAB+jzUfMm+N9CTpeR7l+Vaf9HPfxgJoltVliKmcP2Sl48xUMRt
/1SHjkLA7kkjrCihuzwnbaxWU6yIEndWs5i062LQ3F4ulhgcBX88NePtqY5wlXbDuKNRvUSHqFSE
b/Z/Z6nUJ1MxC+kof5/TZ80dXhAuQoB7UgzqbwG9tOmUrVlX1fIV7EQf2KNEJg3i/8lXTIkrDluz
zqEI2PVzG58g8/b1kSEjjV30avbdDxiPR8ItnvU9omUsUuIxCtz9JzMJ0dCuBiU3jxwuc9Uy0XaU
pBA6plpHQ3fZWdPSN60jABvad2CDMo2cIvFm07g9TH0u9sS+IuCn/SoSMhCVDYERsIICCZZRCvB1
gXvDLRGZ9FqMFZEadYPEaT0/v/Jo1hPNr29M+vjwKnCXBQERcq9/qgfQGYqOBxuvLIdls6w9s+oD
19IuNjaAc+mOQyeemrSpBUsAl/VzlBtBZlnlkGgXLMXu2pb0DtwBoiwJtt9e4sdzc5Z3PgrlltDJ
aKXQQSvrWg9RZ0oyvkeJB9hfsoNDgtK3jtH7SjH99glDox0p9clCH7iN8rOkjotJzqFiNuf6ATu1
uaSoaJwbXzReNc7O0tg4M8jo3Esl0pBRXyS6TRxM9drkkEoajNsmlEphCWMkvcqa96bKY/QY7+QQ
K13mwzdDAGq/MmK683ds5Q+ywpVRVAT0U+ykeDzsAIBHVGZyHL+x5j6FzmK3t/v/PQBb5bEgPup6
IUyi3jjz2T5dGNt6IGrVRvEM3z+jKCjwj2For1wnSRCBgb7XAYwz1cZ9a+LoSKyp05TzCucRvvoZ
RYpC626S+pHWXuz193X4/QL4jhaRCF1yNUY89O0v8mx8zpAC68m+5k7+5X2+vY8yKIAr9N9B3TO3
5ln7Uc4S5st51+N2EjCu0+84EfI3x0aMMWp/sRUOV5EINI6BPg0btx/J+9ADiLCUuLDNhL58Ph2p
u/vqVN0WhonVOQcRNkrnvmJ0PG2C+jOGHZ+FgtWAQkbfwejxeAXDKybMCiPpwMNjeh+hanrgLRpS
vsgm5AmJfebQgl3eoeGXee4jZJh5egGVuy5btH6Oo6AtUKd1Xr7liaqabW7EyjglnUNBZGzY3yP8
6E0hlc8/423Pj/YAPkkFUYx5QZD3QDWeLKmO4LVWIJueShoXQ+D2jVV7vLZZH6/kkFneCG5DaYKU
dhS1K4SPLPXmTy70x+098J5cmYK2QWxxozHy3tiL6hfhxBE7QHqBKVdTww11ao5SP+v3zDAkGati
oqt9QwlBsrHZsV/7eaR9xCmxMeI6pM6lSbts0zvs5mnl7L0sxJPZmCIiGnwZ3ua+7AL9BL1Pic4m
oZm8V/k6LquGFFa4e7TQ+1O5LULNtSbgwwT41zOdtYszxn5wJeA4zTO2Z4uKJ3dfOPsZusaXIh1n
r70fv73Z+xpHdAUFUU/oaiWFuHSwLo3Q7vPHn9Hixgn2Vi2CBek3TkqQhVBHMdKnaY71AuelW6br
OArbqzL4585BLj7oRK7a8l1vYsCYCCgtsm32LVys7Id3uMEtHkLzXhOq/eBZcFolKB7EUNhrKEmz
BrkezcQx4qKpbV+l4J+IwKHfrLqWDiI1f2iKKmiO3KV8IFP+NgdZDSYxYEleorjL1T6l9dTxrhJY
3gJQht8XFT2UFJlbqeHZxIgXJM1B/gUgRMsMtvCHcOP8asuWRQvMg1CS3Wfi1a5zZt9aFeBVrBnh
cHuap2dxj613aT/5on2/amlalahUlgWnsET6+I6wB8EqUJr+xAiDHHgQEJgULpN4iYr1spbYZgZX
YQ1suVkKW9VRZbrpj7R2+zardVQF+Wb0Kcs16d8r+ALj0Tzba5WjQjMdMhFqhZuBwx8bShiCK0zu
ROrXLFZMShTmEdhtpCAmqYL4cNfcHxekvzXcfmiw96UiB21XlBbjEGPnV9m3JgOhg/eP8yn4j/mO
787LQxwr3NIkdyYCE8gDWPsHXuK/haWurLehpRJjdfO24MyJQBuuyjKF/RgfJDKNu87KTiGWVipA
2UjKgYOoaq3XPt2t4frq+OOriB81mSYa8v/HcEItOMmnXH3nLuUQX1Dq/w28+pJOwYkwN9jh0JF6
zpKrbOXkNa1OWAbixpVHv0A+woZKN2NIOqba3SjvQ/Mz3Rv9Tv3IdGmEFwkUJfhxPWBnuohZgJXG
wAUiIhQf68/eqdNkTgXDcAkz+039Rylh93XZdl5ZfVh05BQbXTey2a4M5KKimNzjPl7hT4IE+ez4
pyT163TYPhKYOtrRgWoOPFrgVdkg6xXF8SIrQeWfPIiMgA+IgpCGRnWVFjtr4CuVvG7QOGBTu+D1
nGhLtlyayjqK8zuhcderA9pVOb/FBdx6+SvSPDsCKr2Xf2iHz1TcYwthj6P219b8BsgMNV0KO+l/
R8tEGZ2YOtlid+ammLxLpv9IPcsEuIqYX3uMclcpzRgQ+VrWqcVRfOM0MglxT84VPsHPhgjwKAQl
8ig1U+pK+MY6dxtbPLJedsbYTq6AV1uEHUCrFPrKNEPNkqLWxHcg8ID7hUcMtObIXZqqEAOzcDyE
b6Y4yIdkjQtHBv1micrFKwAjs0/e3pqINFagyr/B7+H1U6ojs8l94gfadDbZAUaHOfQ/GW9PUtQF
CwAZ5LyJ/eoTaZubtDWs0ToNKPKGMC/VgYq48bXdca5nxssGCFA0z3AzwiHLL9fciGh1DSH3PB8i
3aRgS3bmXCQtoVefta9sCzylGmV64WUNW0bwmsO8ffyll8GNGKWthvu9ay/S2dRWea4QU5u8EPAk
NCHxDOGiQcJdIkAeVgy5Es/aQaw8Pp/6546ZAcIEPZX1G8HXv2/Cis1De/WFqtex3FEAg2tlcqf5
pHWa+h6pblgB4XMUPyiZ5JqFflZCHrddD/MdSdBzArm1Bx+4RWzqG24Hz29b/KVp/dtl+mVSWRT0
wjfOKnlH/F1HezEUlj+K/M7xFKILd7JxVSpZGH/kQJcR3Qx7kMj2cDpvKbJ3XQe+XGk4mfj9IGco
kCj87L5SFHrVCS8Q0vauaPXhdqxW9Iww7ispiaMHeD149t0Hu7HAMIqeg3kFnEDkomseK5OGo/jS
2dgarpPNjZrP3zhszkHlEZAm/PWktuo2mWVJknJmPA/RR6BBmyrsiaPpD0Hc3pPDbjQURdxkHx9a
H4TYpamaId6jj5kfp1PEw4rkIElUuwfK1LQwvDalZ6WLigGGblouA1eUjH8ZRJGc82S4czJBlmPE
b+6zqiGo3gH+EQ21NY0Fk7OyOc+nCHqfTgN9n++Q8LlIhkCT6WKGIrTvi4pH0SbI0+wg3cIMAPFA
FZ6c45/buXOD6OodnhU1jkApvvqehbEjSyKdn/kIaKTEOFZtrdcGaMWhfuxo/aVU8KpjTnJhEWkL
eD+1mec3VhpcGItsfD050vYOt/of8CMf7REisCY3g/hSh/B/EeZmnHkBkFcow6aBgl1uVzHXrASI
BApAH9xA+mMAjHOoVa5hgD+e8ZRAZOuYRf8+ZOw0fljsrCJ8ELmo5ZWh0HS86E98Y5Uvgc4sJ8+v
4jjxdF2w7RVI0LnnFgMiyccdd9GGBKJMRXTMgLiKaVIl0+gc2XtCu3TpJK7CRU5ZQaPTXkHKNwtO
Q/8nihYMigDsNOLxTLKIuITZHQMT9DiGTEbg3RhYviXML9zk00xLTxtwEVXht11fkcpXHhErmVgy
V+LQUNFtXS3zR4iGlDsjj8lqWDStgyFhXb4miBju6kfVrWZSMj84NxqE+sWqfycA6PYHg43tuNT/
sLYN85yics62tzC75/yYRDq6A/QfcI7y11IzEWq6YkiBnpZXc23sFwxEG/g4za3UIIA9KDrGcIhA
plvX/2fzyxbylPlg9CrQd1TLJ9b/1GGADepewlXMo9BGFGnplum2lBcRHO1ISnXBr3xE3jNMUYvP
7aKiwd2EZfiN+6ZibA7Z+q5Pdf05qRTNImbyXWU6335o6tGN1SXXjunXKQrwoNrb5fWLN49tVSkr
KmkvVjxVag8CPPYSB31xMTx3pmV+vqEpe4gLaxSOUktmwFlecnvE5xVVezBRFicQkYbvdZddhF71
2VdMJhhIUVEtAl2rBdxNVfXXFkJyU/QBr4sTygqOblfk649jMgwguoisCFVtWjusDjbesF9nrWp+
37zdzjThw9TdHRmJ/i4uz+4SJhCsNYS6+jkF849bhDV4QkhcfM8q/Gk/vR1bmHL+67MWEGVVksSV
4Gw0w8EiyZOe34VrOUopMoNXxSGmhZ87pSrkN8i6/69UTAK/wVbLsq5YnYLMPASgqHUG6XKtxC0T
rtWqq64lBS9cKvPGUcF0xeeac+fKEyfEqJ3HespR21IaWrUugjue2P+wm2yQDHDRzew9Rk4yApxA
SFsK6R2RxTSc0jybJ+fdHh75/2xozvsgrUL1jbIG2xjfeMywMmjxSHKKYBdNaXQ4pGYh7idDMBpP
/oZRtMLR2Dx2V5MNfcnvuzdoBgi5UQL6QOOGfYN/qhclws1N3HVANaaytD6+r3CpdYHU+WQokue3
sqxUJ20IXVqBZOZVcBpOrLQbN8XxCcoBKYr61fGFdMvf3lDRia1t6td6/xCOPzXqdHa2bDv24fc8
B2tF3g36W3adcbvoaXbQFRZk5YKqMDSrBahqhdxn39FJGZYP4COOE/yzmVL7H+HELmd4ejtXO864
poByi44rZry00KcamDbwNeNrIl2Qv3b5YkXQ3cP66o0X+5cgitiHMJFeiPdEbkJ+y1K5fPeDpCDI
j2dibYv3ADwQIRE3vVA46yDgV70az2JiBt7dFgqxJmVuk0Pdl+xWTo4g3aVsJzRrtmSXhIF9Hi3s
qv9YqSIQw5GlKDdBrz/b/9VgIxiqyfLpTEBOjkank8zvjXxKOasde39sD4muCQT8wVjUyN0vQpUl
xLrPcNmx0Dxw4YXvkyUpul/GxRpVA55euxRtLPUDTRwBuqrHqqgahdY8UZm8t0ZaoSdP24fuekSv
0GESkUWuS5RpJiXJPABVG7uEm+BbNMCgnxXDhtACz7TjT32M1+IEbvl8G2RkzH5+SLlhEbgHCPTm
y5CJfSFALJdjqD1rt5SIZ/avf2XI4LjzcNv0dIx9QG06YXnqdvkJbMwhDRCba5eFPcTmoNEIN+R3
oqJHjeTvShD1QOJaggsZ3zCGHExO2why3RHr7DXLpqf7/uP2+sXuWdP/7M4dmG/y5oBomJNxYdga
OO9kUsKmmpK96K/rg04gDQUCuIdbdStboVWxZYRettMGvMecwSqQvoSf4mkPly6XCfCMZqC0Jr/G
ckUovNEpxzgYi8mcijkGjsKwy5DmQ0omVRhy2hpEyikTykhOGphoxkeJ8HAi4ipRWTn4Moj+C8VQ
2YMKKXMRahJLlT+St6F0o/4khZI3VNkDjVUAZrKAQ/0QJa0XXmmjlo1WCzyMOfoALcJm64HOkmrN
3vr5iX0SYbdPwLTg+oNEygOVWEiMDA+ZIZjKTFRpNBxuK8LCBGfNiizWVOozRz+tQG0GzkierAPs
idocK7UbCpUDfo7IqG8w+XHw1RI9dY2VP8BRnAYW4bynJ26ZVXz7w7e5CEohydgzxMXTSeDFxEfj
bL+d9gHJF3asfGpCCdmc5DokXDBbWF4HFaSyYCDh2Lo+fPFnwSHIzlExqvA2OKUq6ibRSledc9Wh
Hse8Z7IjXEoF6445pLDQk69TloSEaMjEpN87IfBfEokJM0oc7s9+eu90K8nvYbujgbABqGfodPaE
Hy8HVGHqzg+wNmsytTeqISiMLzDqQ8SnqdMCWoJL+M60TQRbB1KGgeLjrc2HM+QxgmJR/kJSvhUC
CihGWs90ysyJeIFk06uAi+a6ZfBWnTfcGj0jqx4W05JNjQhGolx3ofbYm80qkMLLpbCbiYmDh5/n
E1XI2lQSGLzjPfvUvF0vx3Fk0txGa6qNYlyvFaYf2OW+f4gojoRkQCM7k4KW6II7l4njD1lWIaAF
hGSwwqsYIiYEwrwyOu2VQXpelYzoOEl9uim1hp1YdOrUG6N5J6CIrGFeJAa00odhG1cIGn2IHwHc
2MtI0iwFNKrgwpQ0k7HGCFjmcxMY9i1GDb93fDWYWLpON6AdQvZLR3EbSKKKnr+a6T9GfpsEGoF2
ntWfovZKFC7CAlDPtocv+Oc3uoc0ICGDQEAMTuckFTwvP/O5u9him8kTBgUNOK+1gteTrZPwPhfH
e7zcF1nKmKIPSs2z6U0d/HwTvxGYInzZ5nY5vgfeDFV2QRmFwuu1LIXz+7vPhDfMalleTtip14qp
hE+wRCx6qYcm+gW3UZENDY8bzDICOhQgN8Glj7lAGLbY5MHuYs9GFFxuL/5N8kzTSGdfk994ai7u
XUwpSIMOILmS/VPYvk7yJXF0U5kMTJWZCXJgk8QNyrveuGhEfSMBY+JmMKpESXY/zPRACcpWimn6
vHb0kHRVFs2GOOIHHG0r2VOMkFHFAnn/MG2iNgLklvwPRrLCh8/Gpl2hwsSJscSYzrky55B6Q+dA
M5nPOwFbpJMemTStyqMTgyvJiEV2QnORMcjpNafuZlaZkwrx6r+PC8OAlN015I1oJfo+boXBpBzK
zLes1SzRB7UHYlLmpj+0KhTZheYVhj50t92Rz/3bSUzWdJUKt5KSORFk7R82s5/whrtpyYcCy9FL
DLuG4onU8SBE3qVjJarizf0/E+fPdx4quBERn7bTRruoTOLA06ja/tIHuna5XEHo1PvZ/QolN9eX
BE+uBRNLA3mUvBdH0EbPajNRU3T5E131iQSoxG1Q9kzaa+eOXjs6vHCSZn6+jRj4dZuHI5xRYW5v
OcUUm5q/kkkslGZanTAzwP3DQ80TML/BdMBQCPsoPBKF8fj4MRWcd5YPFaUd8kEwMIVwGWmw709Q
Q/lYAWpH92b7s/W5ZFYb+OEKLhYzHphYeipv7z0dz3t7b4bJhneqi19CbLXri/zYHk1nIXjknK2g
Y/u5gDadKWPjBfa+qN8z9givh7QCYQ0Myb6VzUGTnTAy8h2nmgj4khBUm6no44tcbc/icM+nwHf8
YHA2GEfNN6W5Y5/mCtQmZXsVrQG25tZ90u5MMLrNC6v/bCmVLOQvYl3vz8vEYp5jmLN2VrijA+ZD
XodsBAazKNoIVY6nm+RRT650J8Pwlv+GK3xmevlKudkSk5zFY+10coxygQm+xtx3aJaEKMggY52+
+9D0zo9AhQjaJQCBveEnixX3PVvcqPG9eEDgvGOWQRvL+OdFMB6wwPLLY0p2kfXEx6tMw4EjsVAR
VoDlsWCo2NaoP8lbsN+a/XQV+XqhxKF/0JhKdy75288fK78KyyoBpHUinmEYVU8n2VmEXvArwoDa
dbRXMRfP/i3GPfY7F/a+u2ccAeASqGZGxxu4y2XxlfLuDoBXjtUr0q6S1XyLXBCIoaGCeOfgF4z8
/6r8LLPMCfx0ngfQ9KL2A5dUrB98X1bIWEeXyVNSVcAImbZxaCmw1vlOAEJjyV/sScc1UMjHkFVP
QKanGknMZ6O7VpKlWV09A/iMuHfz1c25u9eytTkGrnlguTGyTlw6al7vzSs/JeYmHlAIv7pvy+Jo
rEl0/W9eoPaijyX10pxIAi2EaOW8vdy6CQc5nU4CsnjM0zrTFZBHYOreVAChB+20M9dpSwYtato5
le2aJsUh1G824X09PTTJ0EVyimf4xRek3Zi3buDz0UFjejtpo0XfKJv3040ZXQMDeV4NVcPVnat/
ljhxh+tOXWg1QGqi5mDLcgRZjWDm5JXTggzpiHDXT6VAa7E4U+yx6248Jaw0YuK9UKADD1wPRGWS
mspX4vqypUksmH3ZiHZk+oAEYnVdndeYLrhNcprTaRaRX5et91ywVsJzIBtEpIB5Kt5lrJenUX47
hUjWUMhCzTSNeZ2qmg6fRVmyR8ygZjkmauR/Z7xLMF3ZwSK9jzoLyKmVe6bEKkoe3Ka5+jJtAdDe
0MzrYmceLS1LkTW7j9/p5lBrhghhJBLJFC9uFI8m6vMJbRDSe5EZYmmyNbIaV+gSdnW8ES5WAfce
JEMz1TF0HQuLWS9NVhKVCLZpCByQ/tKemdhsx3yPw8VR9FBc/Uk6txE1Ht76ZYJ4lO4GnHXPfuX/
qZfKRqUdgZFsOQQJnmMaNLT/COPjz3hxUhjSgXw00p+GCmeABixRErJ43NdWrHY7oanthirk7+U/
MLdYAvjiWnyjj2mxmAtGGHzjR+2fpAOoJzHWwDerZSHn3n7LikztcBgWQFFpRvRdPfTbMpJywmYw
3W9cCGoUhdIifWDhK5xeILQAEhOEwSL4FUkO78BNXw1lSG5bZXhPxzVtNvd8QfTehLK9/DzYX90E
wV36pyQT5k9XF5n5IgIb1a5WlZ1Xx2c15bUmjjQJC0hgozyFlPBq+dXITax3oHVSOh7E8uANYteC
2V16tEXsh22XqMZKYn5CGnAPyPyUkdTWNG1lw8bfNvanANqvUH3+mvPWObV8vGK62zkxpIry+l6k
VuijQteQIHC4LvR9uR9ReN6yFZBYWH2mxr23MfbojTC3fuUMewaMcYdcBn/s44x6/fIQKf1U8+QG
d/l00+4/ZqJRJyB5A3BoI6NAXz2uC07TKEefvs+v9GPHRcQxzndBumGoD+PCBZE3ype+CjMkryKb
CGtPkaMqFJlSiVFGa9GdJND1AVlzBRgZ7mYufYCcJJm8p9XTRbk8cgme96zIajnCAxqiZX/ItQxg
n/7C1IBmcfFpqxOOmCJjVZD3kCq2CHSszJpgNAPbaTKYDqHeeCZR6LMi4/VX+zm/NQvfEr+lToV9
x90fDMR1Xem1ab2e0b1p89oTM92A53hsosSSdpA4PyRakyYFHzcADTKU/EVdtavXjJCLnDMa3l7X
D2ZHozLNIQaa15XhfFPEVQKA7pI91IcNAVZmlTAhwlkOkKc3hwLkGIFM9B0dKe0dAXLBLqqTTUnk
bj+n2C08E70J/AoUHF1JPNpETmqQ7WdwiJkePSyUTcWKmYnoRDopqF3IaSvUrWBT1rAaeYGNZX65
flkzW6TaOzdJZRantNRAHJ3IycJeEo1G0PxjQlBYjB+EbBkfjucP//dPmNQX08XAvZtJJaDTCk6H
eT90DOEPkIHYw2GjKuFOq+Trle1R3Ih5sM9zI6DvEZaswAcXhgOSg7Fc3KNW5AZ5tb6vIwnkwB9Q
ThRd5KNxMhA0fGAU3dXZealRI+gK8J141waMN2NRMR2upYE/TEPnGPR5eLz0AFkv7ExCThicpehz
/VJuM7ijebgyFGbDZEO22PGk6Ekfb/MLr2oYMeM3jD5pRMoUeAInUYwp3qiwhuQoX2CN+0qiypLq
qosfx6QdnAxX5psk+7+jDANzeJrdp1mnZ3KCWhKN3c3DyPHx8bnHS4nD5NZirgnqOGLzrStW5mP8
CUsM3Bj9pe9/qhPG1yYxaI+1GNGFKQp8fbWO7SqvvVdEjCrnWMNzYc/1eXsnnw1Xo3h3ej4UMRae
KX29twwtBeyYVPgELuxarStvyqnQmaz5/mglAYyBsVQ2ksxiQwSSV4TAnqjpQ0XSLknG2NDhNH/K
7PLMXz9buVcFIrNqDxJOzZgvp+A+43n8j3mC5HcvzvtBhFHESRdiKnLcbR9P7MBkHunUnqtkA4vu
0lmdtz4VIzGv+jW/bklMThl0zBuzLIWE8y9ZGZlwGouGexAFo8ynrYElH3KFKDKBRVyzWwJaT8tv
HlNgI8j7sGcwjwW6gD4FgYokjCoMj/6fXMn7wDlcNYO3KlYuE9GJTLySOf/S2dfgg50t34lO7Imd
j/nS6mjcwtFf6CtALQK5IuOnigWdJow4N846ClW+DSDbHj+8KkrV49OGEoiAu9t0Ik1zdD7eB57/
6rjYDk64eZYRMAMwXFuXKfTxKIiSO3DF2iZy8ZQt/CgHc5L/V4P9m4I69rZ804TeWMio6wAfGFTa
8EkrBxTVGMSdMT4q6ucCeT1yVtDsGqiL1JNRy9q4YGGESZzEbhpoLyQVEYPemCYg/Q61UBU+5lGW
vNtqO/KbYfRJsJg7hPgRcLKxaG70tmTpJaGZoKayDfrlSehdVd1viKKO9SUdbitCpQe8jqTv6AAE
LD7lQLMeO7404wDiDiNFAuXT/urer69M5t2FGgvV9upFF2J6IsZW4R30Am4HiFNt0+7KqKIDqg2V
u1/DY3bPTm+z8ZP7h60gA2kFvG/ZlkbAwUtJdkbwyktSalREqMWw9nCDAGYo9GRjpVYXvtUD6+pb
ygYWIkCTggO+PTz1bMjrZt9ichFN6rQ1bvvLhWK4eT0AP5wBggjjNxV8fxnr0+18cPrkSkYz8naK
XeKK2Yh3wVhGo37DVgba8tTrXALn8ZdEFu3A+fZwaERVCfviNzz+OEMMQoeFR0Ky/wIsIelN3qpS
O71yWYHJSTY47jP3IyjMqXmoM1FxcWp0Zkip9pY+meu3dmIaqYeRmgiKStIe4wzc/lkb+w5G0Chf
KsCVjueCKBYiU088uD0OesiNZ+K4NyLsgsJtVNEslBDO7kxzHDuQ1Hfr8wQ+b+mCKnxIBxwbD58D
N334JOKIKBrx9+WdTu+TG3lNhTBvduSUquExtxv0nfEi/v5mEUHqcU7KMhD8SnVOzk/1i3HTzDrO
Uhc7ybMR+eNNm0UESfLqLIq5MWvVLKSbmz0jyHfrAbALlmZuwTpmpJhsSLa5SUJ37Yv60UP+X7rQ
aSSA239My4RA5WF0SKS/NWHMyuleFAck2g+Q/JhKuN38RYfeSnanFHrJ1viTkr0o52ZWcVqS3Xap
yMdABQb4LS0+hL6X2awhTIKGmbPzoEfIlxKJ0jxAcZe4Nk4i9MQtH2PhQMVX2fqk2D/UwpesmPQE
gJvYUt6Tra2PCKGvpRwnZ/nJ1l7Kyprrju6S/PAtbrUwXH1AHwHzDUij3/ysMhKGfRXmcSqohqHS
QlbVnNerDmIzFmkS13eXQfwahW0YD6DKkKzhq7/zCqA+r3GciRc1Ty5IQu0LZelrJhGxQdoGIzkP
GTQeUHZPUVRAFgonkSQwlTCCN1QtiBjyRbxl1vo40uqxOZzKoiGAuWFpnD5wiToSj05hJ8Ri+Lh0
VVtllyS3J1UAbqNkAvKlaG4oRAPzNv0fuBZpFBPdIvJpCZ+h2zAzrmmooRKljAr0z+59Ga0FiZb8
UNjknnLMtRkwBVRBUjcbf8R0sJLlgRLWB7UAdsSFFLEj9jNDv69x81kqDdSkfOF5QFEIk+ua0HV3
PQm6TQVMjYerCZhq0q1uei5thYgoiCIvBI1cWU0tr/xoFKpet9EOmuWz76ZgzVbvoNYxnl/KDTpH
Hv2FqYFSCKDbNSNxe6owU67wqbyNFSv9x/BC6vEnyc4ui/Dk6vAfhBofx0cMkPYDUbT2NpN3++Ej
GmLQ15F667n+8kv47iICcANTGXgl1m3HFnYKvTFNyerdGIn0rN8lynDQ+S2uE0+jgRjhsVEcSRa5
7lv3dMAWfpx/i/63SVRr9CRcommiuWibxwoEywUCYH3MY590TQvRUrNiEVTiRW/ditOPXTM9jp6O
VJlOL3SLkoE5/gfAHJIQ4HqJsQFlOVT1XtzyfjGunqAh0gDG2T4BjcAm/oM8KIEMotD9uQyCf/jP
Ibk6+tSFxJXna9GoqWqcdWvvlE2KIurBlnIyrhuwV6WktjWNRhmuweJwsWnkVh/ops9aTZVNv+qm
vmwXfxdtwQmVo2IpRVoc9sbbj04iJQH7f88/LBaeKPJzj29lBBMUPC+u0aKEoq4xDpmuY1e0ub2o
fO9sLk8QWlumeLuEY0T5+t6frU32he8kspjGHPqekjvW0XeZEIhUuRy2K1A8DGBDRPj0+jWPze97
g49JNxF4HBIwpg+8TUq03YCjGMMkJmXyi9RN3omlcChhyO+Z4JXrfi9q2H/HjOjvkHtEliofiH1w
7hQaIM8V4TiBtzvD2WchxTVpf7u+OdsFXrivtwQzIAw5KYOK4iu/MaEXx7uncUwFpsK1zKkU1QmV
+rFoH1JmoE/ofOhYaaV1EKwPdxubQqnvY4x69rfWaX5qDzyK0nixoSdyReBCV/uKi286FpiV+dwR
MPDewkVLK1Gp4WjwguIcBKIvE51QfapLnSrQuSOFin8RTjL4/IyHBMAKI41pngfXy+hEfjP3ImCO
9KDVse7OkqSXNOdMRUjK7cGNZcJo/G/pGIxHMOTx819qhv6jJstiCkqNTxd5iQqwRRf7Wypsl8Lq
FnZ3fqDzUJJVIHKZKEEJe3GyzgrwY9rBKgAcRuSC2dx1dNlW4uA3SC0En96euKl0/CQy6loTZB+x
KvSl60/W9q8YE1FW7gnjRVkF7Wqmh/wmryXOYignBN0Aq7c6MdRbdoCNjjdil+rUuEVO3YQQiCal
5tdqpka17CK2qVw8Qp0tGCSOlM4GJh0qPJyhuVAATaIeNFI3+RECuZS/wTrtM3OsunPSvH8OFkCv
HC8ajTNKaFYLVZEb9l2OHmgfJKhM6Nn+lM0CtlDphth616DNWGd5VkB1AbVcFgZb3u7CPxaoB52V
N0k9SB2jw9qXGmEv1w9pmgostyAFH79tP2o/r2LIRLGWqMmMH3CvI0rnUIUZpX4fBfwLb6r5zYXe
oP/3TRQygDHWSdmQQD6w/MZGadrKzTskK109t6sTKS5S44Nb+BCKBb1d7Q9RHvmasDioJZmzuFKj
7yzylOexz3oz0EJ+SOd3UzDheDQu05X7OanawF+/EBKJTF4zr+LWb79rsjnd7m8Vs+vDn/gC213t
GlrpP/dfHfdkp4TCvfp4dHU8RlPeBNhDsxVMh0VkF0DsOFs5awTYKlnUP7wIr8PSkJq8Z+V4c9SQ
IPx/5K4Ov5cJCvrmm1dDtT0T0LwnPqrLp8N20mz/xaP+/KoJhXKln+wiVQEStpUrVgXQYsLgRxwp
M7v/eFhAPKyMtrKWOMw5BLQ02Qg/QDHUIPxVE4ytJZlQJgSl3Oo2XheV9SVMqKD7PMqCcbc6LteX
cl78vwdK47H6MQKpwoHNI0NUbY4AR3mcCBgDaS5+Tzrw+AqgaXnuFkH/vosLwyrqzQWDmoL60wLa
TEbRtAeGIK/WrnihVEikLal46mXDyuzXwZXMytYBl6xIUtMFKBirn2j8jQKqFiEBP3072n1HMa6k
Fd1Amsw51J4fnDJ305fIfjJV4Vc7s6iFKINBq/4QuWRTpRuPYncxjZQrRf8pp/ZhBvoZjr5iDMWZ
jdD8ddt/W+d+3kpbnOhs6oOF0FhuKTUbET8XMcKYVEy0lAnDgKcWdn/003/CKg44fryeo3ujsfaY
BojYlUjh09bK5FRZyEHQq2ZcN417rWXPhW/YHxjsNvm8HBHkPRsFOJHEhmFZ/eglHNoySvIqJgiR
5PgdkKqcgDdbcUdZnNycx7NdjbJnWogK6xr9D0jRPQqz6zrqxA6xURMT0yBVRUzz/5u9XWKJ9J/2
b/4vPkBuZu1cg4iVVgx7BLCoQ8nxiwNB6FPAcdFmmx6Y+OQohsS8d64qqFMvMM4TKRHNKlIcH4Nn
ZwPRzmH0Sem8Z4m2Pgaf0lKVfhERFU4cPXs9RZr4qO7xBFSrbiaNj+xy8D082NQx42uzi8LPECPd
O6OdJ1zxqj4VzkiZnKNloQ5IbmCTL3AD4Y3do8uZCTxEQcRcfFyaqZaMZUhq9fDjHY7nQFOywSIl
8OmbRJS+lXitOnpxleeNwvscceBQq4CsJ6rz7wsW795AAq2LaEmKCgrDW420MyBgUu2Cu2tq8X/M
x+U7ZaFuwG5eKvdy2VT7dje5cYr1EUTz9kqYmu55pzYdPnGm9zjrwtbjwNvBpJsckff8rSQf02PJ
yDWwBhoICHMaLfgvkggpwPeS+dsgGkXgYOupGOP9nSNGk+eSlz+66LXEh+JS2WPGM/5ymU6QXXHD
T1ceTaV7SZ7YvMLe2+AIGGxtZhY8qnI2XHEe8S5qQxSZ1/++NhxWto8uGpTCnqTw73fS2ags8cDF
AcOPZ0SJlUTLtdWKxkNUkAhC68dlsmx6r1sD0EzEu4f4EtH6sedswSXhifY712RfSoLejRZ9ulvj
ln9S3DafRfqH2BCXJzanSOz8YbDGPppXpc8+ZACLJVnK6K285bbxaGxY0fkPCdxHKsAMXxdCA/uC
+pcu00fUDyd8H6kxqqdnKZugayY1XeOvQFBAxGVNN+exjhN8/G9RBfTSfANYLIIod8FRTce7uB6q
vCZTtF+9oqM4AkLgXyc9v/1gwuaIhPr63zRyniRU5dZRcnAXZ9nqIPwy4OSWZLlKakZlFuprB/cE
u7XxvmYwQEjLPAipW+Z6s/anPRTTqajg/ntIOpXvsRz5bd51DOeA3EPRE82b0mRerhNP5qIs5xX+
DRGNdPo8MrE4X5obuMS2ZbbqWmUEnRHHOi8V4ifbQDNImhRbVfa/X49jo9PslxQekxR+m8g6mTZo
F5qZQDTeADS4hpAhjNCsiKDfF9tr9jEJwXCWCUT4+boPJa0amgxK8nvGUebaqwLesg9Wx02MSTdW
Y9gtRC/I7wKTgLPm3ukWxd9GGAFiANsxG9ho3b/xNHzKJBTaiIgPV/4ic2oxiHKMTk+BmK9dFpEy
wE4vN/Ad2/mqavdic5TA5UtqpWa0oFvihbnvJkhFBvwwN3gphqVUrSyjRLSBT6YuGhH3377Urhyc
k8eSi4PpzNk97ubREVIaDpyR6huf0i9acrM78PBZATa7BHTxUdMkqo8Hooo78wxbCOQaglPEKDr9
GJNktUV14TsnO0xFPsJIK07jWzJWMsDc8P9pbgfICM4+aK8XfclHOtrG5pTYawO65teJbf77ZLQy
E8WqG7rq4qO0uW16I+KU1PR0nsdQpZlwkIpXVIcjg+BGvFnXmh7QKowy7ZXYLEdLTl40xo/0Exal
Aj0dEiNSqVcoFvo69PCjBa5ig7aFQLJtwsaKVstwv5sjOCIufOkv8PTJdgQT7U18wTfaaNima3Y6
dZttCGlNa2I3HIlkCEiDvjjw4ODM3fWr98yXoJs1ZKJ3Wx9DkcnXknhBP2o2ON4R6nHwv6tPvroy
b/g/hK48Mg01kmEYrmxzLSIHsCxISIAjzlDn3+h1yrPGN0JaYxuR1VJNrcsB0gE0DNAX2KKiBh/j
M9w9NV9pC7yd6g8AOvYvZuUZHmCWQq7vDT/LwuSYfiRS3SH12WcEUMG4lLNJUu7ExH1O3HOl1z/8
K1+hzhpWKLRUO9JziGLlLSwf3hiy4edfTVgX26d9VXcoCvyJCqPtRotVKIf4Yp1nQpp2s7iZrFX1
ootIqLi466iuoBXBgVXQDlF231T1z1XhaLwlhJhp9a/dlmTwkR+/lORkmFH1a/94pGjxsHNEZ/Oa
zsYxLZN3C67T2g9tT4iLAtqRmkFMN9TNtfmgi8IHeSOhgqJ4yu0tUnO2yqF6sS6rbwoFSkWgNnnG
EADK05Vj8LqdSP82rTkz8f7xZPO2j5bm76N09EgOtIIQRZwAO4LzvDyBpMi6EYMj3m3IbPNRa/He
b+408rKKoZdCS9Pwf2dhFYFN4883r4tjNvj/AvqiuQOy39tHNIm0RV4XMIncBhnmSc3JELWfUoML
d9JBRG1dF6tSOArianRlMYpFf0kFt8RpbZKeXLPSPtGu2nrpXpddeD3aCxJztjpTA2rJr9dRUBrF
4RBGWnq5kr4plcllL5Vv4oI3uvKusv4eZKGzxCYuGBukhZZtp+EzSzcrL7t1C82uNiuqcaBQVcID
4C0DNN1pAbZwh9OhNRhS3uicdto/RkShL9C91D23wCeGG75kvjw6y9xE5mMvVvEfaQevuPx8jZCz
UEaTe0FCeXJj9jBPSQXbYG37szvm/NbtawhDlIPHFW3QaCzGwO+TXn1T+cMJjdhu2Gp4nuHrmiXW
ets7vvsGpKkx0Gf20LIjblVO/Hur7yMglncAn0lih+BR+4gZUdLvE0nc6jYy5/dJXd18nmRXqhSm
Q/eYWAY2BjTB10dxuyb9fM5KDQOgxVAuOHv/2Sve9CQ/NtD1EL+PrvSZOPDsDi98KiTIrO8SBwo3
z8xqYmiuNFXvSHKbZIA4VMBhoO9FG2IL8r4Xz0UnZAuWeWl/vjgbsSn26tAtjBSSy8a52PzAb8ac
jr9BWlUuoRWZrp9YpGrSI1BUg4ZlwgaRn3Bsv+NzaIBIVhodnHMBJYjxNHWpCfW4BTkhpwlFC0U6
XYonThQuSeMoATmO4th7kByvQ0wvEOywYmhgUGN/Z+m+7P0I4AQaqBspdFm/f8BoSkxkhz2WaUDS
zQT7pIc2C2KLDCiwvNGIvdlU+5BS3j06dU9v56H9HQE0hORL1/qkMFldyCVvxwYJpc+RgMc+KkGe
Z4bKl37NAnzXxRY53BVq+odWD68U2CLDCgjauAs3EW0Q5FnnD+zl+bXB/eXvyhMOQBZPGYAqvT7W
4TQv+k7b0HxTnO4Y1bY1plq85RG6AVa+SW2nc6cOP6Qf7z7RGfPxxM59KYS7CTctq3ZnNP+k5zt0
nNGuopYq7Oo4XR1TGZhH+wPwELbCgOZsxkOSkdT9YAY9tS7wnwqmukOY0KdWkrikG46ws/bVupx7
6BKMMrJg/YYb0Xl7SvUtbbF4ji9ykl+ASaX0KJgsal9gq2WkenbyAlNHbs0syCExtvTz7UTrS6BP
jlbFvhlXSH47gUlv/+wGpeRBzjLmbZhV2+sYueNpochvNHASbll5Q8S0Duc8yYpd/zHkqv6CdVCD
S6lTkEzZaAFyaxSAKih/xhoUPfqmzCQUiiouVUSfDqpc3kfzZjT1l03sDajnBt4v0JU1fPRc5tjP
cW4ytuqCWcjoBcJYal2+codt9xseVQ/eO110lKjQ4ZFqB94yVHX+un1ASi0m4lMznmYAh/C6QDPo
JPJr+TITlaY1E7lEaR3uck2y/ee4hIQpXUNZ4avnYiboa3RzZFI3t/rCbxVEpDzOA/XMTMKTROLZ
Uh053hKoFKQu1ARwkGHHjf/EybFdy4imAppRwfCM0zUsyB52XI2QBIeg0e1t5jX+x8BNRh8+qov2
nP7JL/Fa5iNO1RppG9WQVRWuRruUmYSHCvBI0syyaeLVHdsDQK6TXv0OnDVQe6xN7HTiwt8zM9uI
/Ci8l2S0txjqjnAsMkh+RnbYh6sSbTtRsd+AdQPwZR/j5MiUTc8CTWHrQsnm/SqX2mXvnU1aR3xR
DqkWKT3yRn5WCBFbKGzg8Lx096g3Ve/tM7XrCPGBTUVjwH0oPf7APJrda0BBVXtBy2CDntxkBzPk
O3QVwzKzx4+VHzCj84H8Xdmwqfp5AyHBGhlBhy0a9Gbp/6mlJ5yGNNM0AdqHau3/ijMMB0x0EPMB
MImAIM824GEfmFZDUdHR/zZy8N8Q6mZnd0081dNK3P71ad5YKBmOB+qsEVo9+k1xa+AO/uusdR3O
kmnVDcil/sTfiiKWRkukSQzo7zJE45SDhxBMCbYndXYIM6xVdKW1fmdzXUqg6FJNH5fwt8YNEaZS
zqQJPOFjccsmiQhmwVqmJV78OsaugSzIUYpmexMVlLqBGqQnPsojvBqOFXjdE/J0S/9x6rIQhFsd
H/HeCBepodksOkX6t+055AlCDgNUHSKQjFCLWj6ygBGRWNBjROJBGbNA5+b9x79HGM+3YROLmN3i
wHGajgv4/AQTIztU1emLSqrfQVCKWfHVhapyst5EwtGuVjd3Zkm8gbB2sG9yMBHcvXFXzSspg0dZ
Ay9emB1lrEJhJ0IKRIHVupi11t5RKtHRFEkvuAVYsiYs2fdMJ5yiD+OD2AABBeFjCJgSGzWGRH3O
ufbu/LaK/0GO0R8bM41ZAUOSdvX+910pKmmtaKnzLPLlr8NWgfEqUJ1wrxrPlHchidVc+GFIFRJU
9UCotyk12t4nEDCwgrPMdvM5XlXKep67TD6xXUzvd3FaXLFjJ9ND4/V+ym+wegp6PHRvkmLNqDdt
uRxXszQFe7DcwDpnUurzUKujZQtX7k4vMI4uuneJWuqZC0HHfqWN5q1bpOmWV6CBrvFPorxpTXJZ
dBF9Y9JUsbf9wi273q/C8i8lhriUsz32nrmD6r7sAdqCQTC0ly9J10IlQSVlOoY3ur1PfOX+v/WD
p6ocCarwIOVtZz4xVqGbSxgfd5COK3lF5M/Efcgj75TX1LJPgFSSwkOob/bjdNoXEZwHoiEzru0J
2oq+/qwMbPJQhp3ee3IelkdKPV5ac1RCUwaicnCXMsqMRMUj0NETb1N3pcmfUFKJoyMC3T6f4i2Y
Ugq4ByXaBnc35Kn+0sd8BkK3Zz93tEQ7l/SepbYYPpAiWNrXwxa7pr2OECuyMkgU2xkjlq8Do4zQ
tNbRM5SkMYt3RXDaMfb+OL61FVcCSgigxUceKARFOazLC+YP+phyWe5L0YlEo6L+K0pKdtO4PPeU
bz60FXWHgPawC091ieYFgJYi2j/FShMtNLYespUXFLj3pVFdsegBdmNMpTaqgvQ8WFEOpmAnBzQc
Lha2RSPfBFOC8uC7Okjz+nF+wg2VGFABX+1diuEox3YQPPwXPlDkV65jNDviqAl/2ayi6vNuZkY1
HS5WafsD9gZXZRJGrk7OnAqbBvPL3bDYJqm+nDblKsjB+BBHScmCuqkRZqDo3TwR/be1D2LCEbWD
FfY22lWj74z6PWsWOPrFA/JsRtL0wLVN3t22iJTZt1nhYVH6e3SrA2cxtU/b3AJKRggro+ZNMMtH
Pv5N7b/bb6ESmmhkWEQibP7L8J3/H6orGlu6JlQmp8PR/Y+1p/NJHpK7Y3pVpaNEbMXgQjLEvfqj
2fQr7sCvweJuKvVn7g5+zi4lQ1cDsEwa06M8zZbrwOV4RGLI8Lpxg2uchYTkwhyjarGRk+J2c3Cb
WwMw+AwrEewJHjnArjMPYCoGQClEdRrT00NaTquhat7K6t7xzp5+uQcHFrN1fuWUqwRvWONR2McK
qfnBKJczfB/tGQkOBIpu+AYVV9RclEjva/CLLn2IneZd0TvKxRWIS63ivVvZGZRpdSyPGUEv2VRn
EnREPSsCK5ZzVx1IlhBfJiKC06G+rPsxu7Vc7ew4WqjrBQRAy7IZttt55+XE0ijCQrX4WYEODFe/
EUwhkFsDhJxwqi5PMPZlFDLgiiJSkkElNnwbS5HdV44n+/ZG+Hvn1+v3s6JEifVqQqCwKHpkJy6I
ZVCUD1n6mHh0DaW0jqzfn19Kkc+Yj0+pBHNt1/b7mJjtiJ9P9DrkVN4sCzSoXFTWTyVZS2Rir1a7
L+t2UvrR1qj2O18hmqRWl02g2wBKDsQ+uEChnBn9NwJQnmkFEgbltnQV2bhXgLRJ3HB+TbUPvLAG
URiMsiA02NEzCYmRuBnFynPULKPa6fgG+Jh6dgoKglvukKUzoksTN5WJZ0yG4JH+4TrWobMd3gOD
c2hsJez6+1ZBS0yGdquYKyF7+MjNIfigg4U2X/5C6EtqjGwyqJrytPw1cQ7WOJ438S5EupztgA40
dgOt7GP4xVuNM06VSAFdUIHnfil5WjpsFQ2stATm1YpOyr6h1E4cqe1Un9LpCgtQOkqG6lCJs+b/
/jmVCiitVjxDvYtUXVciJMgdqsDwyldsCLsmSTUjXjnTmY4u2ZebQOldSfqjEkXYXwKvTK+c5nIu
EmAEM9hHwTR59pXoTN6oqh8ta7yCLLRwZF/DOw6UoxhLxT6AFvXmKaLIaW+Q8YLp0u2SCXswy4pu
2LR4jaiQG95g4PyGvWZMpPvNd43uy5iQJS3DxmIAn3dXqj65nL0SMDg5jmbE3hzX60fKKMNmh3mm
RmUjG61tK14MI5szSz3c/w1vL28B4Bfs2cKGJqs3UsKdLvlB39Bpdz/kMYoEA0QIv2sZ6xSq0Eci
Vakzz33yajgUrn5UPaceEleW8ds2JopDS+igwlBpquitLLDC1ZCh9CzvM1fz8B48OwELZmv7807c
uXymUzEEYt5azIb1CuB0Cn6kxOuIBr36chmQDD03vgHGrftfvDVo/Ryazk7DrJaZbZ51fJ62SX/a
RS2m1N+b5SyffEu2H3JP6ZCRcjgKY53TaBNuthuyoJtLme44K9Usz3t+zdD83qiF57o5H3SqhZma
3lV3icso1XGVm206p+R7xK8xza49kQ4/ME3g+mipvqZi5CfLB5w51lbiEfqLbCpF7BVc1ztmYtdH
KwpDLGp6PptAr924qUeESeywVTEkzpcsMah7GbN4kbENFqpwYddWXPgB59pbMKFI9xHgh/gL4OgQ
VaScJ4j6KnjAXxDOxRIer342gcpHyux0N6suOu6k0SOIBni9okswrylumOj0Ed7Dd4eYA+WElsYx
VZh8bJSin023cgVlck8CXLKJGOIUR0tRh6ook8GQDMF/pbRChJShV0/xg7wW/67Y+eyQ3sr08VqX
rnq1y5fsVtKdcembYdleC+jWDRs132xYu6wPqpZVI23axFKWocSDhybefHLmcddUCDseo2zl+Vp7
qUBO6nZJ5es22Dt/38o3Xi3U4RPj0K7AinLjyCqkYt+Ngzk61l0JOTwx6vJv4blxZf87jA4yncNH
lJxo/ENNvni1pIj4+qj3xpFxdmV7K7T8BR9/5c6Y+IeKRVrbIQOWlvSG9GbggNoLwseeHA0hp6AX
vOYLdLX7v0NProhdvyd0SHrosAxb+AfZvLsxTXZ1eF2NHuP7o8U6ZZsMKLX0+Bh7lrD4vOQFb6Lj
fQs3GfF6m0yaXE88XZL9wHq977SXHc5RdHpI7CcLeb6orqwK2/XOjNQidhBbAQcICFE44JQJ+oxS
zNCDJlNbELUYElS9vxBIOUaytPwzX2u1CIyyce3GL28fdPNh8iGjNzxEn9tYdP5OexlY9eWYyD06
Hm//ZgyNVPDu/omZ7CEy13HD5WtkwQ2BOOzbh0HFgWAJAcvhqnVfL5T+y6bJyPuxBJjetI0J1or+
YT2AQDJwOclhMr+rHw3KDhVIQ2jLo2iyGGz/R2+Kpr+WmOudx36VBzBAJFTyX3t4biN4UGVNIOa9
kDyN5oeBO6UWVs1yHnzBMvuEV1WVZXyCUNRzQqD6xp8YWOG8mSjlc1EcwJmndp+NNUg+FIj6JXN7
+I1I7UKYJ4RJbSevyJb//XuYgETkiDD6w43Jib0j89Ekzk7yq5sazpyD5qoDxTMCcqJklsvwSj8g
fCLHN262bv9v8ZABBUdDQyJ38jIkXBfJt2gXZKNBFFtTjrJ9XMKz7jrJOwjkA2S0SgYh9czOzp/r
empelt+BPbAkJ0el2zWFpUwZWOd43gzLKhClpJxgpbdvpyqgcSvpalqOg+o+0u7znhLrh98nHUl3
aFzlguHwL0pyiVM3q79AqItUD3OvxMoZlSNltyge/4x7zFeNJozaTzSeUOYgBzChcTbVZ7x/kGiM
P3WJpbeDnb/zcgJMKVE/W1ROk8As255/eAiqWNoj5dFJ52sG4dKjVfGVT3hdX89o0eVYFPokyRzy
y166EJOzjp53h3oo2cZVS68dQWwnwwlXzBE2S32QNGrKaMIUzfbAeBAx03GTcr3spKMNGvMMlzN9
4OxFMR3OQ22n5V19Ui1XSelPKr8m0Usn+WNvhg6PgttSBRYz35/yTL718hJXMRe0S+81GnyGAk0S
RRbbyMXuBMQGabaqUGkdOmgnzh3UdoPJ8dhdt3I2I9mk2sSf9Hg+xzLV5JiBIQVqM4CzLxCNDwgE
31jewfdlSdllJkMEWuJI5EEqWVcbbfZZ/OCrA+wL2Kx7/nfyQkpCi8qQx8qmQPE8xiUkoKN66vVu
Jtnuf5Z2NE6177ycMnDLo2NHHwHeCREH2N0RuBkiXpYAhlatMZNwRkgrRwlur6u1w/N4cQAtA7JN
AhH8gsSy5iip9RNS591h4iSn6ad1Yjw3KS3wWLuS13pHW951VbOmB36zthQQN6rbpV0PHpkFfLd3
Xbwe4B+XbV7jTRY0+n42LQkQ/RhwbZ+70GrFEbRnduOKfVZQWNIIw9Efz0SGqjeXoqmX5ACnxqqa
fJHgdXD9DP3D6GgHw2U2Py2FmqCpeUhIUFzcsAAQ/YeLkSGP0rqyBa+onuaDen5md3p7gBRv6ZiG
k2BeHHMfDiNG0ZkYqLQRpr2w/KyMRyoBIAQ4kjs5DH5Vtr5t8CMLHUhEBJ3mwM6Sc5N0yPoHiwdT
j1lPGMJ+8PVOuun/1Zab6Lst4D6J5QvcVcsH8G+ae+rmaBYdXUOQv7LBACQ6rgy90GS1vV/ulTnc
Wplh5OEkNS4t5CNlOvKx2hi4nqNapL4JG2qEsNaXeqCHY6qn8xRSBR4T/T3dMnedqkfQZUM8jWnw
JW664wV4oNdMdEDdhk4rbZcVfVcjWArwVo2GkAlUQTwvSyyilY5AoH4x2Ot5fXsU1MrOj2JnZh7D
+FkDUhoeDcoIW2nAqdCkt6+avGvgD39Nb1VgNq4RO+aRozvH4i0zXibwUwVmfVXjfOtIVRTZ70/x
WXzFblxJSfAbqAk5wgOrDK7yhMuVpSTDlF4wlUBkkSoNVvsqXGJBnrDLTne2tG33Kim2013XmYXc
gCHBL0WRm6Hk8M6XR5/uZ/kjNa8kyimzl8+wauClQZCLjD5imGr/kSHpsLEN74daUpSdISkMaGfs
1+M7z/9IgNg4784UJ3xbuh/nuGAig4OA9JYKNM+cxtJLCF2kG62aHdJdcQ3mlnvPibzXHAVn9jKp
MRi822LcKE2STH1oOWqBdaanXd/uh4mvm8SL1zh2LlUWkmtYJxBtEiom9HqD5ut7kptU2Cn1mcWZ
pZg+VhM2cIvcsfD+ydTGoW7ELq6njyoDSoWOIiGBUONXu+/QFxQDmyKAJs9xN4gQwkMllePGR3jx
O6ecLd40HlLkUeoketlS4YUHn7qbZsHWldk3dq38rUKr7obCwk3QCO0rbp30KMaYN7f/vrdRx3Le
A5Vjz5hWi9MM3AFnxyW+5ut8MGBK4u21VSWoJ4Y0XaZQXPGr7JOdLkG/RNiaPLX3fRsPlT5yAMax
ywpBYOekRLC74phVYJBjMxpvM+zbuzM4BN9m1WJcBsCKx+xYIlcec6a5GTOZGF32Nd1+PNEQVQzx
+OnTafpP2jW8fyFmewHD0WlFCCCJM2PxY9KbDaA2QxXWgXjRoWfLvxWawyeQpUl0URyz4uNSrjJ/
N8oqQzaHpFkkxJT+fKwUGtXORfH+Tc5atTfWvv7N198acLQkObxmTHDDjt+b6Do8IJcrfLx9oUj1
FkG/8P6lvfAJtJpbMdG1mW7CYWUCOtlTyriif8RKVoKbOMfnWhco8hhQTYUJppm1Uw6hHaiOPZhV
iYlwoZe+cGRlp6o4SaJBhyUcAfgCZxPoqT1xFB+B99F4/hWPG2r33ll46GXv8fjevfOmeNA+/W94
0aD2uLnLv9khtOTD7T2+6Yd43EI4h7FIJUYcO0AXA65HLOfUrhwa/Qs95DukjWj1S/iq3INZxMuB
xNJRN/Ez7gw5dZ05bZu0DK+cKkSQ3ePFp3CDRg0Lp699Y7ABQIZ+73BE9b37YyOzzjhA8O2d2+gF
mL9CxOmuq3mBHOAmIEpibHWTDWGCDOM/+6zfpecHvC9/1j1Hfb/dy8zb57tjxACGck/MEKENvYH1
gSRo+YDkYQXRKOQPryQ92tXhNxqR+J4wtSbaXRJE0AV5PEb7dYk7fsHP2U+M7PITgZjt9CFw5kow
F2b+58gKxwnOTo60qAPhUmlf5sZ6HukmxGb0YBKfzuFLoXelh/9nFwyY2VrTfdUn1l17iu1F7W4V
HXe/qO1BeEUSkBrZRuVukWYMJSKiOJ3nulk4q2M1Ld2RfKo2357aYrY6gQg1vgpCfzTybSS+oYR2
HWz9snGSysYOUlHZTSHnzsNvgvOUtp3/cCnG5+tne+3FdiPLYVbMBmFknA0zR3A2YEDc4LmXVoXI
TraIKVwrsgKjePiFe8a90sLqpJE+Q34GnvjIgPpyzOTrQy51bbmW3zFFFc7R3JJCzpJFASfKZeQT
8I66sr7FlhNExso2CTRVKnO4tpRoAqGJQZ3FCsq8fjsMEZPfFaE67BHF3w35hgl9cHDjEWoS6cmA
k5P1arFzMi5pyo82qBJ6/eldt1oq3yTRO3KXeJm4gTH3+KiC3aZX1ggzFCz2cKdkwbKoXtR6RX96
yv/9x9yz8DkwmqZLJZkPFhHaZATfKpUvnoG6y4LR5VBL4egeJTDt+crt85rC980/9dUjui4EXdLF
1dpFXLRcK2Yxtpy6wjp9KSs0OXZPUCewlx2Wli/f65gs6kU2wGJSm3VH1gkrJFsqFDG70iy3ifqK
hfavW3ZylVvnu2iD8HB3yij7+watySPYAvABCG6KFOIDENiKejd2AH1oT3zvh3to2wb1Gym4lopD
OASPyQjrZJD7Uinn5BcJ9Mlyn0pRknSWsl1dZBdgLUOfi9uTmuo277id2Yrz4WHypIe/6oO4z4Fh
tx+GTctvke/2fDbBSGEsxJOQWDcXoOe8wEjAzQASHRQ6oci0nTzLSoEzxrbQwHAOF2UGvNBocwDS
CZSj9/x/IU4xMnSV85GVvp5VxquhppIKTCAv0t9QX7l7lh9yKJpoSQVwCkpxl/QTFm53Gqv5clKh
WcBFHySPL1vpwUTgK4f6y6AEP0oJQ0nM3u6gxWwNT1KDLRtrH5Hmc5DpxLOUovMzbCRdG6FVPogW
fc6GY/6SClvklrthp9FN58fvOpDfsBWR/0fEWc57gwImjbh2waimBq4fExBI/9inxNftuQHYYxcC
ROKh0ba3OxjAhGdwiZVr4GN0Ix+4n+G5zLK4HUGQQdHHHOH7gsmk/F8KOY+xIuhZqKO5x92p3HNV
ksPgpNvhApavVkkvxFnmkDcdAQN89YF+iEmCJFap9n735kEP+ipATE8j2Xja8qt8E6WgpF/Kw0kH
NaWrjzYdNi1vIaaHEzm9yXIUY1GZO0WvtGFJEhqAttlbBjRe3+yShhe5I0Ae0yx/50df8V9/YMFZ
ACdzUtsT3YjlMO0IyFVRvBXiYn9co5dken3ZSKL1w6Dcy+4uq5bt8YtU5LDQzquMlFvYJ5oSihbM
X0LCBZ/TP/ZHl5Jrot389h9IsLiigtNFQtFC8/iHViwqRY99EUijzEwun1FrVqbgX8NsLjmsAOqN
6Y91sfKEWfDDDLBI2pZk2ciMUlL2JLzG6PkwmK2Z1jdbu9oZB1lj7ic3Un4X5Z/3lZ5IPvD919G4
XgFkfQQ6e3zmOmIwflNTFijy2KZQpA8hE6QbUgn0/YWf7jGcUamWwmvQQrQvYXF/PpKNn8xqHmDF
RSBOCYV4JRplsv7Mf9Q90iEuvkvdtKx9uXYQccSiY4ti1h9aOVMmEtiUNzF0saxCkiE7ScPwla0/
diwo5EbaOuukKNVF8WE/nnOBu3dlqjvhLfJvU9Dr99MC1Nrn+CuaOcPUjTguo6TeBtNzche1LLeb
WJdt4+A2tNmVtyE2MaYUporSgIkJSTQGQUi+F05zRltrMEYgEUNa/ZKawreHt8u6ezoEYITuxhH2
CqqhygzUwsOg1fKA/FyfP3SRxVzY9xXiOseYtuzjF3pE7WHJr5JpMz1QEppy0LlIEGB1YVa/2rsu
d2r3HwAQC/PZftwAQaJMVRYo9FYvPlFN5z6RaNTSCp8T8+O1Nn4fRn90m4t3TNPSExeonNt3C1wL
MAB0URsOXRQu/kyKpBnfezvMNe7L+whXYPU0jhlGvUpMzedXLVVD3j25cqBYBSWg6QfTRn/3MJdP
DQA16uY2A6vqHW1UdO3DfT6gtepKEED2sYjJ6xW+huzEuDxu5oD8oloikTUfV6kh7OWm9qzakdzA
5bufF1evTBcHqJ+e0x/nlgMPlPk8GmX0DkRSXtyl8fc7bPi+KxNmVUvBExbhoDnJga6dAeZsUNza
A8vUqP3dGDYjOUmcob+i4VHySW16ehfeamobDmwe0DL4wq8lx+JicKi0XhvpWRy83p1iv+Fdxln4
ALHjSVTf6pUeVWPgmweSC9vh4zLGmiIONdq/B2ne4kTe3kzIOlKJE6EcjKTfLw20Fx0n9UbKPiEM
v9s+PaOlnrQAjU8z08uWIy6Nf/aI/we0JR8EHDXOHXxeAOASZFllgetN2g+8eaL8ZJib5sorIcng
WmRrdZX0cBc77bOrvbJhxNeBJnGsHKdeln0fhVz7AViO3O9dGyYtnkKMgcFl1J3/rOqflWUOgyUc
EfKFWVCbWSQQipJEKjZd+a6VtCAe8QMD88o5nFOgA9+3wEWsAoZJxU2u39CdFJnxFYeLUqIAVVur
kaDFOvsITRUd1RUCuRbQoDtiiw7xJ01JB7Ju7eAFdoYt2bB5PwNSi8FsiBbHGcIWv/wu4eLBi3xN
t/ncwzgUw1ZgJqvAKhiY/pM4J6OT7tO75VjYb+4oL/J1nGUjYeKpuszkicyEVujH62JWxd2s2igm
AhYNG92GOwy/3d4o6e71HRdaPxs8sGWkxPwQuUhNCB7JiO2yp2PA67bF1Mkk59K3nNJKt2RedLED
6Gtkj7w8nmCYKiLMznu/IRddvFFIP4nadh34si5Dfjv1N3TphVUxmFPi/YTF6hRWDrgNDhnJl66T
wnUsdYocU0MBOn5nnePQK4sozBkePxSX5tPut3GnxA5e2COUbB//hoLzcw1N/8TRjovTZgCr9Phy
0aRDStwPlcZEPNnvyjPKlIC2aHbaBGaXGTJTpca7jepD1lgzCdEnBRdqFVq+jH+EuHtvF2yGPOuq
0k2IPmC1RKFL4IsjKweEVL4O02ee1ULqFcYnipI4nvaEK9IXjQ6RUdhEPZywO9Xgpcabae+cnmfY
09hL6zRmEW6EtEJQlh8cSdhXliNGcLpnIJdioE6BsTkVXxK+/sieDrGWZSPAK86UnXRxb/eB7tFJ
/SpbnrgB8/r7mkFOQVGnWMOk0v04YolZyN7Uf6TcACUGjzyBiAKAEI9ifYcT5RnwqHhpp4IKLss1
PC3VhTWmSd2dHJr7kkXn8w+5cnmNhpewjj9VW3JIKvTO8Hc/CvzhNSkLVv5VuRSwbyKCc8Q6Iexd
vRYE9D0rEJDbysL+tC83gdyJl9V1jVvRtCQzNzlJ2HbXe7Gi3JEXyAWysVT2MXuUyIjfl9J8gg65
rHsjMpZy2DAQu2LpwaEq72hkgtlojutLIlicBkYcEYMs/Z2Lxl/siHTGPEsJaTD9TfaaU3MLRqBs
O7k4yL7xksFV9SWaIHR0qIJDBrUvw5iosHf/iiZLGNs5QFPtIgBGeWj4q8B2w1WKT3jJxzNDZTBP
c+/uQ9rROP/F0AbRWdGF5Rxte6iTtaZIp4pKELyB4FvEZcnJ42gnfegc+naVl7EwUCoHsoaxCFvV
y7cTU17P+3YRshSsJQYkMn9OOn3rD683IH5P4UNKFAKTj6/8/Su1qwCCcsIBmWonJP3MdXDSWZ/p
+YQGLQilIr1TzBKvMC30byka62WeZ99PZdgojRh5/hEPtfXhPvi8+5JJGsI1Kob72KcRbATqitd8
+jaQzLUIJuftERaMXRScDtldNnni22bmO+aJYgSoWN8v1gctkUPnQ1hyqGAwVZS5RTL6DxkbuDPg
cIsR5S+0n6sScUu7jL3AU9LUaMxHNrb2pj4X/bilxRx0n68W9n7r99nC6i/w+gOw73mvlVjMzfpE
giuEbp4Nkj0O0TXBA9VIH/4NVBH2l86PFawuW4mhmwQJCyzhZYfdhYQEFheIIP3jUKEljztKtB9Y
JUZQUmFh2F/1TBC8BR3EQyzbBOzQckhDmaL0hvfzHWjGe3FZQo5oE+pPHvrNxg438D/4kR+hMAS+
5uNBe6h4rhgQ522RN3TVdezbEoKs8LsuhF3mCybhjY2EThTQEyrwG2Ggy9a6E/r2FQ5ocNLi7FzM
21T5/gYx4FgHqDQudWuPSxUwrp+w07W2d5jJpQ5ESGv3+mJZ/wrU+DqzTX4ufQigMpPG/Qh257ot
cBlp6N+n/Mm7MbKK8Ezn/7CKk/hxCZXLWvetVQt3E+vZ6SKYecLA/z2Jsg6roxinJsI7ahU7aVHZ
nwvLnHnaNTGV3sLhXrG4I2m+Ewdjc/4m/XsbB87YDdyYyM8behKFDgfFUPl1CK4Ah3hlTmIm0QwU
PgGjy9smM02CqA6u/s2NxrEYQfZ41vz76eVp8fcXc1S/5NQZz2sgp7ubexyV5dGkke+5LKQjx1D3
bxtuXYiuvuxqBsula89omFY/ZTdJNRak298Op3qk/kdTqPVGuVhwycguAxZ3JVjxZe50jhjScn8T
XNz+sdnT8aAPQZ+WxzbyBLogoFiCJvK2/aIY3cV7fApzL4ktar9fLqc21+bptPAjeg7LPgpTerYl
00jShDges3c20diijc3Fc+P6MRxjhMwbzTApAv/6dmTVKaiKLhtXxf1GEnUCzxLAwkA08ClV5ag8
PNF/opC5T7UznrNP1nQJizobtNp8pxfBPt+XojGylq8eeoDydjK+zATY5wn5gmW5BNiYeTF9I2eW
Q8L94ul1lkuoonbaYCwvzL5rA0MbsjXVMsZ/X5Sq8GuhW+VnO1SZNvWrjQRIftRQYf3Og17PsuPz
9JipRc2IbgpLwWF7ursMm5xYQn0mgEHzG7aGHzZ8TL/7tP8jjSKek5qGRebnHZIqKy9mQMkJ8hVp
QjHCvax8aPGEU8Uhmi6ZTHpR3hZpLYbcRUqXiO++DHYcPeTD9kVL/w8ZDM5sS8VEWKdLgt+gEXrS
6TR8d0503hkbTGAYyTOhXnsE7+OaNkeuvFhoW2rec4Rkzabpj9saGmY2hWRBP187ex0qT/0u+V56
3xvJvYLF8qS0+1WwANyj+GzvicyNuN3elvplbBzR7ne9r8gvpF5IEEEDW+9oals/21yq8wrZS6Ve
yKP2P0HBr2ErzdA7JMaXqTMvdbaWG8a2zWkvTos86lZkDEeGdD93DiuliqQNP4p69P9r2JfTDgo+
6S/mn/pKdIyBj2BrujyMaVIVU231dEq/syI2JigXx8JwXNVT4Q3DulGOhVap4gv3vejNvA3ybDZR
LK1zwmLh5aKA3Gz4V/lzZs4veG8hKszDK4++ssWoyk2gUqC5dgJ+oaffys/vws6Cc8DTd1+DAg1w
WdwHMHcmhxHXZekZKhF0i8R4WOmKBU387/PYaeXtp8Rw5jjgbNtmLfBpUmmykb0ah1xvxGtbRcw1
D7ex54xlv8ET7OnZ15AgsO8kCA/PoH9EeZ9j2LVz6LrEyYpzGuSxmmApMgskKkOjcAdMh1X0gHYn
4QK0IWFCh2lNasGPHp5hFjE3D/U4aYpITbp7Lo58ATjl0rNxpFDNf16PDBPFfexkfnh5rQKMnxus
rB7bVXIk0Kvilhjg2WlVOLDlhSXkx/M8JcuFK5It2yo3mBUfDvzG9wjm9jpumWOLIE4RTI/TRuNS
OVmfbEcxvmbFdQHACd29/SJGRI0D9cO8ECJ3YmmUy5+9DCHAtrEsQ+rRMU1LGqLnwZEX95UXoX9N
G2hkRiqijhQJdJivKLvgAe4jFU6zF5TWX0eW2STCUvgwn/anJaM/vCfWNqwTxN1OS4IOTTMEH+IG
K+8ukA6MtHZThE/CEa5U+wMqFbc+LqIF49gOmdEyFI87Eiwr7oWCERxTO/3Stzz8DgrQE64WSkkL
lzNhttIre84/OezHSFXaRrcPV7mVEpgSWDreL7zzbvHGLS1+tjsb5CfGUJoNfO9doW+dBwoXCqzX
tYws3Ze/LmZs8+jCNAUNKLoxGU5cBGc67NUHspW65Lo2D9EqbyvIdVcIsOYwmePpo4CfbDaHqrBj
N6ISDckEltQirSRMDEik/gtfkaSTshqbBIbLpoumcPi8GopWOCuQ6hqBLPefk86Iggu/HcDzF3Br
+aCqB5vsqIqSIj/sDMGkY3CtXSRkPUFezd0N4jVoEiAlApqw6bgCeZfy2ulNgD2rm6Qjg79gc4ia
yiIEHLj+X+nRudHLGBGotir2VzzrjMz9CqotWjhgPy+kYL+jsl3CIWvWThWbwXB2VeU59yhWyoEP
quFKh+jshwqGoCV2l+pISJc8/oaicZmfIeml9q95tJFD9grKanI6QxXAWIzcNSpZMgua7K0BNrjo
YnZp+mTmLL+JQtj+dDgn3Qrl53Vv/6R2Ricz7soNgu7L51Fztdu2NoPziCbuEwMz9FZFIJhfavcC
G83bZx/OAGMkLfK2hCh9TV4Z8fvXxp1GEcX4+5WlRn3VJhdH5o/nSZnfxFSQ13P/eFzBzEpDz0h5
FXjeO1olkkV9UpwfFxJ4uaVBehJ4P57nzfWh/Fw8D5wgnOjdim7OUuoe+H92joswDHCTv8Hi4jd+
Fp/hmF57jMHR+HhvU1KoMbm3WXI/AkbzCfAM/5wXjdlcD2Xv17DIl1BMpPbtE6LAcuKPeRyTKS2z
Voo1gtjoeINDU9guaVvCqxhhflikuhVHUw5FTKe+whOnrlsIFUop7L2FaSJ8c5bmnoavXTboZwPf
kIDkV7c3znwv5RXntro016bW7n98JCoJ1daqaAZTbQu0pufFdqUkKd55u78KNvher91/K9KywNQ4
zzf1IdrVsHQfPT0zzB/97t//A6Gu3CYhFY/PtuR4jjDQagytiKrur/ESZUwJTk+si2uoGHbaEtte
kgjRD7oK103eeBHlWtqg9PP9emBOsk2sN4ruYbS1d/L7PDHq5Au3c1xXkUjOywnJYpHyJqgajulm
cjlCt4cEebIjnlk1BV5OEnwHzL6z4byVRK1gH9eL4wQ4JEheMao2QlA9QWXY4JgAR2HNkDLe15d1
Ppebaa0pYvPmcWC+fgkASpKERb6l3LhGm39Ky7DDYoHvMJb1ufXYNWSuZYrLATuJ0Rqh0bO/Whv+
mxeRoDV/39w/KBY41+O8bytcs/qtFwgC5o4Gm69Z1RnG6Jk9zjb+BeMtP/Q4VB+n7b3ujoVPKzRW
2lVjspvVVKDwFbBVGU5zScNh04MDP6pk7wbhhopoahPkVwwBsjM5Fsarm8JOFJOewfVyuzXjCfid
qyDoX0DjTobPnQPAPZarp2Kp97xkx+8Z5H9emE+rmbvNZThW2cXZJkH2K5sUoeUWnPSCC4hUPg5e
PPMz+bf2RG6rUyoqHSpQRmYOaQ38u5+/7AkUZ0fjjRQMXqT4Y66K04CdaswvcnqTauUDh8hpySlZ
b7B1Fn6jlfO3GGJI/9qyVH7eMB6+gz8mSIUzU6FiLLBMR1x9ETnGdEkiuDxaugYcJvvnDylYsNvr
HYeVy2vBn3HOnU5IYhGTbtRg9+8XAjzHEqayuB8T7e2OSb9T1DCI7/TyBYPPSswTZtgxGplGxjLS
SpZ6C054bH6cfh9gPpx5J0oCZWzeCuUFYQeDxt4Iag2FCTQvGGW/DY6Q+uSgSmc/OOCUcmnVQR8V
O7Ch4knol76IzhOgpmNtkuMyePZSWS67n0bV1eI1vz4WVrhveMOGj9i8F5FkXY9NevNMX7F4RRp8
mxTut4KT+eAh3rTaMQLFT0+iO9wgvBOy/JL77rc52lqB+0ATnK1kC1pm5+8xeCjZX+PNymAxW4F+
94CeX8D5ooIPBzGLwQ96ZtBTkYhQRlAuGc/wqvD5V0WPwz7y+eUxeHi4pWIDRj0F0frAzsc9QkIW
TJCX5sPvPqS+nlQNbaEtU5R6/bVFQLkVgTyxiWHSCTLGfsmiYlel1calmmk90suJ1GP76GN+JCb5
Xag/c0tRPKe+u6Hc/Dr8zsDbkW6RU2avDUjXmLZJHfS6oqGGb+W9xesabTMUMLzFZEJiA+hi+QoR
+1fJzEOHo97OoUhV4VLO1iBPzo6mBfkhWrIAf4VdAaMn2vKGCpKP659UK8AM+RgaJDorzvxgfv8Q
qsEgHrIMAxAd0zMK+efUst7+oDNMgwYVLBoDQmk8eNpm0KWHjdD6etud1d5CAlBys4p+TLpo6iFj
4ezrbMYf6Y5sXddvgCJZns+zGopQ3nERn0vhGn2Dd2Eaa7nwFiV6o9XVN1LmD6z0Ftoj3oSAiA6f
1G6Fu6uIGAvH7FFs0qaZmRljmteMvzGxdK16xEInZAvH5ST0EBtm8lcHfOY5YaAPU2RcES1Z2uez
KpqR65x5s4aZgr6STA8nybhsEGSkFXND66SD9gayi7IqIV+H5Wym0T+ZonjhJmsbgF68xmCm+T1I
AOaBGi+vT2+MqiuLV7UwGEK9NhfOrWEbyLPCtxwfr2nyMqQGYOtswLzcI4NC2/KBCfUkgbojG7Km
vtLVxdCFnA3XQXiKSav47CQ4JbLkJ7poZloh9JqkgwOVjU4A/6qElMyjKuw9assO8deGlY94Md7h
0gb8XPKUhRd2BkEqkkZB2IE/vWy//Dy3czcEkrtcX9EjxVpYXdGO1q4DvVYJySOsdYcj1mZukP3D
sLoVwbO0XIY0euVBiP1cvbjS4YQ+cICiwTn7Hr/Zb1VHXPsLZLtO934qVSNaLG9oJG3psqLOTjQb
GxuMKMrtS7sOY4OoDE5By/zOYW735G1Wd4oGeilzJWArW+1qiLnM5FQbFyNsUnt1BXfnKmeKwVQK
sKhP42M8LYKjRfbc0PxozHM2bfZqky/z+cW7tzSZECJ0mPbaf/cZCMGJi0EJ7k/Oi8J9Gj0cvGAJ
jvcoDUvIjwW86K7shYwa1oOaTVMJc9WL1DNshuOo7c8ATOniYAZno8Prw94LIajS4NvLT8lscQ+Q
GkzMTdX2JTCHZFhkvYfev/lwcSPTry4t55NTAtj9DKHhCPAc6tG4MwcozIZnqSMTVB/6KpY2jm5f
930Yj83dfScymYJ8z2BEeyPvaBttxwn5QOITU5vTSwUq+d2p50g8Qq0+AGatU4oFIDG5qlTdCzV3
o/iC4Dg4PcvQlM0YYEq4raq1y7k8yUJ35lCaSngSuMZBn0Bxq7BWJmf/miQAtE9vs2HBkjI1UGuY
sK3ZEemXYTGF9VC75DACQa53wdcKT0TD2YFFkNA2lY80TjBN7j/EwIc4NhrbL9Uw1L3OARumEeYi
jHDPFHf+XDnA6/JXek1e6lSNcgCxh/zzbKWVhb7ywhKHCBoRfvDlyfDNgYAZu9N4XNdwyM0qLfii
22eVMEi0QK9Cl18NBgNof+0zE+O0ytz1MHWjM+TMbN8co5imApw17JzEbkg2jdHxJPE3nQUXIV2L
p6C8mLucQuPFqOqMqFmVP6bU33cmVev+c3yDfughyh3PUgFZuKfcfx5eLqly7mGORlNoULKmM8k0
s0s8tw7k91bwAS94EiG9H8sC3QOJcT0pXBXdEpVqVBMtBVVlkN7YyjENp6Anu8HWsqM4x6z7DiON
MFVqBxLKBhc2XG2BDPdXaaCCF767S+JuTNNULrVYzUX67cxSIBpXUVum2ze1lq+Ww+SUNXnBvRMP
WR+GmrSALP3A7euD0cjm/BWaTNw6RA+xPq/wFJpqEJvF3OV/4DvtiTey0nLSal32Fmr8WeU2r3Pd
+fIAhALxTyP5Ns3iuJLB4LexG9UmV9796I+XYNrkabu++TvGuPmbrupnTeKpanKYSlG6d89oLtXp
U0i/WiLx6Bv1quQQWmg9vsEYrw60BfhfwheO/DGLRsWlgQMUlhQMYjLB1FMJGBxSj2cjAmUdVyHg
fvNwfWuq526FiGFsV/gwMGmrcAS3EsM9zQ9YAuNObN4oOfUf+4qdkdWULW2OjZNHCwXj9wwU0fZm
eRBMtj4XotgMVS/I5rBObkER7F60H0Z3PzY6UU7HvoZ7ip0871E7nuhdw2fT8URYd686eCIMBXVj
DkwkhTl80vbPhFtDAYi/7axAP0vqxjY3ONH5crAu6z6JWjwVUbLQYjcSfC0t/w6s5xjZvKtsnelS
pjPiWvDkxTlH/NysnvrwCl0SOAp7/gQkiAZ7zHPksBvJ/IwRYEp24FU38PEiP0Z7gW7Bj86T82fu
nKnEhku7rb83hD9kMxSfjxkjtAgzU6MV69c2mE4UsNBdiGHuYANLOGBlkgE6ryMLonrcjwoxb0sQ
fzPaEGluKEKcJCJc9HVIY39xyxWdGkmqYq5AGXJpNgtfxiOf0TUT9rK1XO6FtPsZ4fN/V4BMICW/
dv18lE+jp/IUH/2330uxzNKVyOvVSuBf/L2X6WYusxE7ungiETybXreut2QGr27JpXD6bKjVyA3H
PqXTy8uomJaXIE0p69RX7L3jkfgwhKh1/qH9HAeBDN5I+1jSvh39u0DKk5wwHSfHuCkUZXGb1hR8
KV2PpKox1G1iDeRgtqA+/17PxEWA9iVWcOqo41pSgklpxb6rEpC7Bw9RxkEmEdp2l/iyfb/vL7IC
SbRqKipe2hpiQBxDvpGDWSojsZUPtuTdmWyTh0TUKjx6gah/ZSfChzHoBJ7nIUgZ1ivKu4vdlvV5
jntisZLeEEPElBOML8K9D9qmamZjw7Cc/eY7/OBMCUu4uklIulAVMTKfnkwZDc47i2vcRFSJ6CU5
62aqQyZV3A2HPFZNakcucOdxERDT2VLLch4JArAKcscVJMBo6BKLLVkv+dSEf19Dr0Gz2/lVJQrH
dJmD4z/tZmK0lJccqK5HMvcqrEphoo6u9c4B8G+0QBMQzmKJss43wwpsperCbO8o5TDQKu3JjFSM
br3EVuYtAYDQO7mDazUxI2Mh3MYJlVj81ejH4TqIHzpjLVmcjlC/ZYdcOvQdFBAHt5CDpiUmtW3Z
3JZub38Ypnsz5LatXA2mAF7tCiFehp/IR2wxLgtPtV2LuYibA0b+vRS4stgjQaZuMz0CFOT9vMBA
6X4dNkZkVq8RmaA7m4qh+ew7ejLie03qPNcGg98dFtoipOOi4fF7nnJVWBQXo7Yc62kqi+qXzxFW
8xCfmTjV+TrFwohw286B/crUHCaq4RMBLynj7OaAo2bm53jgCt6b9kny0EwHI3Qu8/w3NG3kLAZ6
VoMCJbIRbDb/tT30Tcy8xjM/5p0fFgyjE02WpYwMvLsvLGs4viSIcqGp2UhMy+vZCSKs6xA9Ri3x
PMvKEwUyosTA9w+PJYOIlUtQRA+CHn9MnJ/2N8OhtzXDqaRXSe7EjkAgVpeSvtXspDI0Fw5RBYtS
hzqFqu9waFpHxrIt/gTP0blf3Rll5sSKWS02PnkpfVuR2uW6O2Yu63Q/NLc8PLQjMIP1QPVhJiF9
jDeKCtkL8YCd4pRQRdqir0/BYpkXMJPwtTip4h1vUz25eZiJuqjEGHZcEpsy2EdDGopQgMOlvUC9
0m8Xm2am/0MiF1P74M0rGvmu8WSyZZWTVXwpylvf5+B76erQgrj2EQtoIJVFVN68lZoVkLtsNzcP
d2OGQ7d557aq24B22soLrnsokH4lvdUgHZDhPDSwmQa2f/e4bK8OKkwVQqZrQSHnbFhM23CtNDRH
jKXcbNNwwfLBSgg+YCE9annWY3XjPAYwu8YDZLDykYRF3NoGIp6tJUjU3PQiLD9o61ng+XsQQK7n
X77BjDxx/kxe+OhuZqAwP3+Zx3PG/KAEth7eyGaJpQb7ET6bFkBgDFzjLozCD3UaO5LsiLwP6eGE
bVlm5MI3RZYMcyvtf5XXuoudSoONZPif/eI4JBfdsc8CdcOIxrNy1+Qzw2pr7gjJOuMLsI9Giu0V
iW3GTUzLrfQYgd3kiiovBlVlUlpM5MoVFDA4fBPLOI14vVGjEfmMmdVFC9+aIVwofyGRlZOzs10O
Dz7foFFkjlvWIkKrqTWZ85RzljzalCdZI3GYe6D+Pi36Lq66tVFutyt23F6dy5f6MMgAw9WuV3uY
/k6cD4jY7ySyDcTel9O5obQbJq6eQ2nGZMIZUtun32AbYdllqja4hVDPD50frWyj0AG0M6Eu4wph
MrbfJ42xIQpbIVChXkjy3q3k/mXHpKFbytuycIn4Y3bEOESYvuEnIvqnxKale+1hodL2DXAvx3RP
oNXMgy0j79ay9/TLgCKw12Xp1GMcLEKLjs5T8svhbqOzTwheIXl8a/jRMKmL/Ft63nm6zLkeoP3T
v4Q73WRzuQChYlsMTr8iTMH7DxIx1SMUN4n0NXAAa/1XCPJsP71lbxeJLwHDRUIIXAA8M9ThjoX4
Jh1CRR8cIoiFqPTLJz1uu0c8e1CNKciGx0yYoM9oRlTbLWCieuvKwlJik2hAw/3efTBM/uwTDl3e
AritvqXb4QWZ1/faVylht68WdGllFeIafb0zWzhTvuSuF5/1jCv/Y+CrPuVYOik5QmDeHmWBAVPp
ASXPOc3Pf3eb1ArLS/SkbYge9WuTJGDhgxY05KQxwIe2RYvK1ZNFu6UGMrZg/oosN/xa0APEkyZT
uzWXGAysaA/0DyCBhoRlBo1HK8X6n+ZWRlG0WoGrqzIkOpPBDpwa6bynEPliTeYrOUy1tbK+j/Eo
Y0tRWzK5Uw33zE6ENDzTJcyy0wS6B7tliteLq7iQbEROfzypOIuUINgFeUnr01MI7ZVluQduscVY
6KWD4GGVTAjjL9uAvU2nX0DzjVUsrPs9/J2knz1Gcw5wvBZgziTV+2rjH4TcsqCuiR1wgW2SfVt3
bpQr56j9Qm0rvJkQ1kkv7U+jXJr602lHQ4ZVzPFCaNRRf8+jVHiS6q59zxekWv9Uxs66QfvHaxI5
eY+G5WeTS3y0LMNKF70DzVAsMQAl6ngR2OjcxDAEvgjLk3mL5Die0MxiFBSYCGmBwgZD5qBONlL9
NeUu2A+4Q9Ho1IkVxJORny4voyEOJLB1Bd+adv2Spp5pPebK0Bd/O6S8lZKQ3PZi+roqePxzd4ot
ZgcuFWNeXNJZ8j+IObtVS+fpVfUpKVFi72MkFgn9Dma2v9NpF21wFXyMNSL7oRZofqy7vwdRr/O/
lCWe/pL2NLJHhfXNSZ9sV/T8Kc72jdywMRKu5up4/1xgYFIu4GyVEoJJOxxsl+CSB3nLr+5RzPZA
7coy6k5wke1b6OYkbLXJdzPbqYS3iHGXkgkAVagttA8c1Q+htzFek1A2hwSfNiunXRYnF7Kw/cpu
AoLuoPhpTcn8uHMJ/b4ZXGFvVHBd6EUNA928r96HAdKgHH+r8XE5V0qRwpRIro993oszmcHkIete
z4O1X4Jwdiz50ZV3IKWV/ubxMaogKU5HNpwInsVsBIDc/Q5uAUNMp+N51QRPVwZP16WLoIGctqlG
AW2scxICZFXMYaCEmPKzRwa+tQcHIczk4bvCVZMKSUwvnf7lvonc+zMqdU3ycw+iiqaWgJBSQ1wJ
wWC9XaNxVfWZuIg2dgSncy0K68rltptCd8rgLTEpHmhLRTRUaX15KYJHAX+fv9bhzHaX6thz4wM1
vjIbQ0LnGm0AfE0qoPp+WMYlDNgK+kvvjVrtLD0hxs2EUw7yLIVeUI9uWRsA1gIKJVgfZnv637ck
77AMXqp1a71WZ4nT/hc5+PIOeXvJKhlQvrxGGB75VEaaEccglajA/oslFE4jb9uS3JVRNGWdbS4H
WCbj0Q45l3W/ybVFtBR7n7wtD1o0T3X/I/t/A50c/c8B9covIvXvlroNr15pe6DH1UadM/gjk13U
wvqkTYE5i0gz8u40O87fWui2Pp0mXdKtOFBaE1kH7Jx0UZEMNibDPfLOvE7RWL+Cn/29gnPJiSJw
CvQbaexrmQWbjyZlC8sb5Bp9UvAo9PpxIjh1465TRDCMGiIs95RqHDqxiy7tDZNs/VdmqolvZxgV
TyviARSQ7SNt+Bhsb+zA19d+EyezmDEl6sQM3w57rpVJOkPLRnDxpX3q8MTZS4w7JBQGkYxdAOt/
hBw2cEMfgOEizYc2YbkHfaDUocj8IDfMm1DQN5HrpFS3pfrFTfwR3nOM/UuE1vuzvljy6Yrd5/Ho
sV0mT4wVfy2awCMlbrbESr+EOWLSdXcFyEIJ7VcLt0CZKEsC2lJnC9d3BANe+FtzINvRz9PZX+u+
cEMrQ/sZuU0CoRHXip4kehO1T+QdjEuxTLOFzWOLz4SmVRaiffcVHp0R5EXOTPVlQIZAzL7hTWBu
sZoqkiPPVZ/5VUB+zzAxR8tQPFyJMSpN/OBGnMILMAZJC7lRMFt+9lLB2civO/6z/WW4uALQrubc
7bohSATDw+rJKvb3yUX/S4LL5tuYzrTAWp1g/DsPpsHTj542AsYwPIQXKOE4dRnCG6Jtbx3H6O9d
k3QV92PwcI0ed9ReVcslvp3u9xBuP2reeMZ6LaII6rHaRpfN85qHtBJzgozLyhsh8bGiHAGsAXO5
WpiuQuPfNIqs3YllEDDtFSUQwNbPVMaS6nXdqPtcX6l2aJVnXy5QTBpLKPACwedU1bRAtv6H0Uez
urP+DiY/KTHntLX1EP86Y06lrlULwSU11MbDerLdq8qah9h0TVfP0NPJcUzctjtupWMFSfgEnu3o
bJEzEur1NZPiBlOW6C03U0prGpOcXFT83eQDpeZXws6aBhTFaa6dX5RRL6fbaUaOgBDNqSf0jC9v
zZZ7g1NE4wAVRk6O+AEdziJjuX93zjgjMQevpwqL7+BusHtF4XMt3uWd4cOPCWNs8Y9Fc2eUw8h4
xs4xqaCYJEnOZKFh2uPCvpi6jm/magThEo3+g6ptRCWdjMkCA4a30fgCktIqLfuHH0HlcJE0k757
qmx9u7tC77zSBXDqZ2HtU8eXVSBM131e0NJQ2LaW7GJt4Baf/iTrVp4+uOIL0CmSOSDtscBOruN/
zBXjpYQCI0PdPt5XJ3zHvaSHjpRUjb7IArchD1uFHUmlwnaq/OcbIbag00AUxJd2hwvFlwrNj6Rs
2TxSnvHEMMN6wuY/OncxcTNk0u++Xic5WtDbtmpum94XZbBZs7mx1cVQ21/p6ZfhBh7nThCCvbqX
May8jmNvm/ROkwfeo+qUoOyyXfjCBi9HHYjCnHu4Tu7pZ7nMfQKhuoe4gA4s/3NK91TIeBfwROdD
kNXWEM61zoASAJ+SifgVG+mJ5KvudTlyvrv6oJXXeseDRqscOiMKry96ohnJQJzSlTuMfgRZ2xqQ
JQnQphx6wa3ShYWoU+ZiIiPWyKOIEI6X3C8Goa+gHj0V+0SrMd+tNMwMmTBquO9E8jvx66LVPuq3
rhIYUGbw83nsvqrZBZvRSghLLDrClPz7DVDMuTmzgCp7G2VOLHOqEw6R3ZkdAr7wEsYzSDaM6jzE
DmB9lI0oLLuX9oMa8oI2HhUzUfqMJuzhWDONePC/83/6pQKXwymgU7pM5bq5YcT72LnlZjo0Jsue
LjdXtxXik3oacyg/6u7SaGZDtowYzT0La0GkkdHgPs65+xsOT98W+7JCkeVZ4x2aCp+sfTKqUt+C
dZtUNRLk1Sq4yD/K365Ua0+2CEhCLZkoGejCpMOvjtMRmWcTgTk/wgrlFLtgbYJ6+cGTK10crk/X
lX4CyAYdY1tcBAiyfq/OR4ltYkymiCObgp41o8HZoKwFc5U/rysW99AfGGKk5ZAvKW5fXxeqIMMq
07i8e/ViH/SAdiXmx34YqcTzgh9Tv3iNDvNs2RVUTRziY2pTTk75w2Q9AKP68va5jHODoVpnJNrb
2ngc/Lq2ojbN3uYQDYbITJ2qUz4SlMCVHJMe0iawm4RxCHJ1IxhQ/QZuh3yqSndoptofkrSxabtS
GO5zeSu/0I3ydx39SKNLXURdV5ax/lRV3TQ2AZ3XpWOoLwtpn6aEJWHSU5SiAk+SvLVfqoYBJ++B
ZIuVh4LkFtXCTt4eKQBlyn0KjNnE6AZAK5+AbPQmP2HOVpj0vWwdoLrMhELVsm+Bo0rRoU9LhOEW
w+/DFRMgMSiTClbCACQKpejwb8bQ0mkjWjwKgPeh3+0JAB2VKODomLKxRvUxo8TIM4rUoheER7UZ
C25WwG+4Goq7hgN52mNNdrcXa7qj66vu3USIGjqLmdeRlNh98HAlTegFZqc51/hv5r6cm9f6yhCl
o5i3qZSaVP4TK+B9PUiqdZ/FnEWP7DxgaAvpPI9Jc47LalRqFsBrY8u6KeBGtpt0XtYsxW6U4dk3
BhxVQNCpg2qvQWlVpM15s2EmBcaOmc3IOfnOqCtoEUZiPIsxveKo1jwQTgo5DLgFnnahbtnTeK4h
Eb6rQvH8ML34Q2M5hkayeD645VeoxXZLXB0b2ofccohpEAuJ1wrpVbc7DvgvNjpHn2vpVNurGQVH
B/sJ7vsy/FtXIw/JwHw5fXKy+db48i2p56Ip6VvPfi1tNKK3WsHOABvjvfS9ILDCPlJqDgh24S2G
PZDOX85cuO/gyl+OGeL6ZJrOb0YO0bADgBugS8Mf5g4OgH8YksvYyOTMKxUabmZlgxZRXF5Dy9Q9
/M6g4/U5PtC4NsnxC9tVDY61+BWpV18vt1eAgN4F3IAwinjteeZ11aixOU7nF9vGOb1lOUFcWS7A
WVhLiIWO6schNgAmL0i3H3vTfapYnU41MBH+dc12Hnn0kRZ/kVlPs3mBcPQEF1Hu6Uug+pwwAxY3
1XDZiG9t3xAHJNxuicobtAyikWvk5yBDCZ3g1NAnYthvBhvGimu/l+pa8y7lUfz3gndo7zuNEEU2
VSa7rrL5RN34NLyNSLIk0GRD6i57Y99j2GICUV40c814D+fdtIZlc5Jf0rUX27h/ZYAZagPxUZt4
KXTLXp8r0f4+NbbqS3KsMgdzRmj7dbGXqsfBgcgyslmHcjcAaXZVg54LTwvsRp+vLRKvpR2bfymo
Zg88pPYeasMn8h66XFu3m6eCApV5BmeRleYlelB1MpDzmEicEE2HxwF0EBIyq1/ZFEhmwaxHAhcN
2DOUIaLvLX4zu1ekyqP3Cq33XcLdG/FYGp7b/sXxQQOLlLzHhFSefifcs5TslJhpYL2i1s6R+P5E
Bk2btIoyUY8fvOchlnSk7BPRsWiAW0ydmuyNBCKc/zCLKrTBt3WIuygh7rVooa5SYLZUBJa2GmGy
80xQqY4S7siZPoKo2dz7qNUtfE/cpNBLi4fbtB6CeBvb6wk4OZB071Urhoo7WvdXtrg3kPy8sv40
uo9ZQmtIgKdyJ52MQBKFC/o7zz8snd/CCsKPEymh37X/cjFMa35wvuhBNaKJrwljBjQDYVrjL7Yd
Ts48DuaWyllsgqlbz9ooXxCHJcyc74p3BFc36BslG9qBtaOP6qHkLPW78vWMe5xkJkkSSHwPg/i5
eWKQOXvEbVioJwtafu2ULoLVePavAMynfgwGHbIpEHTH+bu4csj343FzUNy9ohXNXyfcV1ftQLGe
NBAWO/Ewcab1HP4n67ZDaxo61RoofuIc3ewLBMnblapPzTrt6ddMPJyUMM+nhd4BmGAoWjCdggKp
KLx6rf62MD+3eSD1Rsc7Dr/10NuEypjesybGYxFSnUjLnLIxI0QhkT0Dca/5CWY6xl9YLU/KImtn
GM5WA+cFQOp8fSRm6BU6xAk0Z+NEc2HFpU6tngU47MGv/yff7GjFOw9xKs63B/us2L+2GJENa30k
XUXvb2ubRBLe4qW7kDGqBj+VDdk/fWLeXpxoILjm9HMv/R3oem3VMwrh8/AmXmuMicvwD0Z5fZJU
Li4wQZooU+2gCAl4v1cvrSbBCzIeaxu8MWIZWFCfK3jcVgI876WUBeSZJxKyKByA0Z4AbW4vM/ZY
HI7TQNrvBoNkh63Zgh/UMRjiDaSwN4wTQDJFIlHTvJrP2EOqs49wKtjChBzOjkeE/QwvsEdTvrK6
puQ7msqs+unM+9GjRiOy8hawv6aGc/dAqqBoAS4KqINXNQgbOnKqBzcO8U364P76gsXhMnIZd9Ug
7Jak0ZMuhHbyX3q2s/MTm4aCgf/nUTJZoZosl390sHi0xqdXWgeFyew5g/p3bJIF9tParsY0QjzG
sOO6O8zZaTfOA40OvzzNwnCFn8jwEj+Vp7Q9M81ToeEI5zOauisUK1ehkxQCbNeib5LeVEPie7oB
78YjjI4xKFNHTY3+SgSdJou7bU19BL8mXh9uS3M8g2tIkENeUizMMmLmWBrUcnmW8Ok7mA9EGuqm
MsYHXXm6V6iqxicfMFpGclbZxYgZPcfkNjPZ5VmaqXKjMFEUMqHKlK7tsx3x6mAP/I9rDkszFLZQ
fOfv42BgDVBOUGtHi2tKNYXksgb+IDhhI8tJTmUlKjV3nzuhQsb0G/1z2vhC5+TGxu2+QqMbHQkJ
4cl6bEg0C/EjB4GWOlzo4j17P8mZWDPbG84dZqg//LLtNbGXQtS8sLC9gUBfWRAtCGgNuzrsPnRc
BLdB43DCYSP6kNQQJ/Y2pklbIRj3kaEhfG4Bm7Q3Xxw5NMBh84ulu7B23K9BN31EAhEqVhxSECpF
v7GvXznOznOjiAIOc0VDYwhDvnDaN33FSr+J1TRRTumvf455GXcbdxJ8AgdHiK6OyoJLITBxmHxK
QVBgsqLZj6kcWbVEzXWbG3fIK77f2SuCmCISuwM3PAgSVrl0bcmUQ6svqNUwT/NGB1QzNguolBQ+
qP9FDSlrs+J4ECq5sBzrfi0nDjvfP6c5qIL+R1ya0NzecV6edUyY0QFFwGzyByuRcw610c9392Mv
nrlwsCgd81vQepHM4ZvU+rSCJuwvb9A5aGEP4TPwgT3PBZ1mKU5xTLJs6P9m0RvmRMOUzPeX/kfF
6Y962zmpBUvX2/MsfT/qNIK9YX/xczdWTmQTSyXG1rlKPqwMQAECUF2LHlAfPPURGe31mDoZbYqK
9/E5yvn1OQbfHqWc0CVLogQMVSUmoMVqz9CpLhy0L2qVkxWvGFuEtIfILDjmTIBiTdSLrkYNGdij
L31PDqzXKto5P47vM48uuT+PnDwjlLlusHKlIXusFkhDjk6AhwWJuNNjrnnJb4HHKzqlNkiFxWsw
Pm5llgoymkMJxzVADLDXP5aG621NQi1jCzrJmD9NnrhfQdss70W8YSuWL/1bcWKgxzYhW+d8oIql
cNipJnLVbrv28pjg4ebTEXvYim7dpQ5PMTCNLuQB33Pu+r4R8X9L2N7cDJrmXEsGXBYPfF8pVdFk
ninso9V5W0tH/Jh+og0foLRn9k0pdce0LplVVwSqTnBTDoRfw0kD53UzOV85j9UkiyQIytF8Bi2W
/It8RUKlIAbo0QHQGJc2uAgY1VLG4AVpjoyriEJo/ann679/eRg4kMPPQn5sRD1FBy33FxlAUSNa
g949vWwPxoPmbpYPyVHmVl7vJSZVE9REWMzP9dF7+NAv6BFOu2vAJshqEvdZgUiIV2+An7jWTgCc
i7Q0mIyptH6hAErqmb5qW3TKcPFVMFrFPTjiHW7AHlKeB5cfvFzAUFlk1kN8sgwAhvk1JGjKbxXy
qsIB3hlT8tvJgieOrRsb2iUWhm5/+uwYdoTYNo4LOcetP9JpuniJsSyhhw2DtohKqHDVgO/udW8B
UuvIJl+yjnKzvh38XaIGyAruLn/+mfOCUvhopUeA5r7KJDGMLpY2moMGa3hUBUc4V9qrLJ6u/m8l
rRE5uYmwOa+THZe9H53z+1T7SYC7V/muU6KKi6RGlZWibCVaHh+iF806o/Hhil3PUXLw3iq1T7PA
SEh6+mr8oz3b9+IyC6pmDO7OrVBAJVwCrvk/+69dnJE1rDOSyY9QQVinACmlMcI++uRVCWILhryG
oEUnXJ7Gp4XMdOdaaEM9EeRXc/pSH4PnAJWWt1ff2BYU2tHeJuRrrm7sehqxuK0befCH+RcRV6pa
4h4ZSw2IEyzjSeyu40yOyIPcA4z/7v+bg+yrdYlM9JVkJJhdSzNicFeUo/2Uf0P9BFPbzRB39wtY
Rle6OEfOzbsS/Xkjl1Nh6oF6d5TN7vjsjybQ9w5BLXLVBVDoNxmIDhxBB4zpWnFEnsYnfiZaKRCQ
uVcB8xWVyXnCbetcC0iI9IoKUrMicY2u1guPfEjquM0WJJiMUJdpl1D2E0Wz8I36hOrSepjAWopm
XlNwO5nkpHnxlbwwrEeo7KocS0lFUhWkvuytthf6IHR4isCY7sRd+h3LvJlWrJ8w2mVxQDjllIsD
ssC8aQQ+f9GrIYLmyZ799vfFJNwygLBuH12lfOXUjKuez+IsDEXx2wM2zMu3ui4ewVfxLnC1O+Sc
9T1Dl+gGCTTuzAcHU9iGUf/50p1CSCmd97nWx/dfzWCuyz82Toe7mG5BmDnsB/Q2q/KhAzffqp4S
obQOqDnbn7ryp4SbcDfmgik4OHORUYcgAMe/PMCKmzRaMuycomty0gWhwp34GZdfqFYn4H/qYkpi
4E+A/whXmgDus2VGtD2dd9GGi7RFZz/zJS/MKra5YFSRwXo89tNMJ5Rnyf4y8IIHapl+ZC+iP3BH
9LdMLfhNMWIAHICkdl1laOWf9tLeg1KoG9dYpqGKTUPWx64xpTPfVs1SO2PKHrEY5oVX4p+AG5a6
hoDYSEm1vLU5S0lWAWtgb40B8DkDsVtuTFvSHv2SJCbgVS14UoSbomOyCcB6oq03j/7jd+XXqK0a
pSElRz4I+FGa0rqIRUv/XesnlKqT1Qw+6NP6uxZNLNG+eL8esXYvZ+DduPyJ8bFN13nJdN+s/jZP
aRT/bNEZkNAx8L1K0UEMuR0t89aBDZsoEYc2+irGveFABtrSU5hIa/u95ZSWfp7yOy6KaU+10QYQ
CPZphM2ghlwtofQnkhv3YuvmRcQfsisEOCDUipe4siv3RwaEhFfO2OOJvwbgp7rXH2QEmnMAYJpY
Uupf0Q5mEQZIVVpaH29ze6bYTwAeLhD77mV35RI85zJqtQSihbDm+/QjRWB7/QjuT8S/BvKkcXxK
DomO5aQiKL6EwbPUx9RuH+A8TnbUq3zxBl+Xg/ADkpSs6gOXp9Ao3q8ypAGtYLOtQzlVHYAw2CXq
RETrMg61SJwRUOnA6N+H8IUe+lpiEhwyKmamlKD2gLqxpMB3I3rSXJJJMM1JOfrVD6xYQdv6PwoE
jKgDxbOl4/Avv9Sc5kczuTOq/0jJrNzbRpejG7oeA1CFmFOL+OMCsk/wm6Z7tEj0BkqkjDS02rCt
HDP519hkvoHCb9pZt0nTDKhra8HRL9oFdOIKfp6U+S9ng/gDwgW+Ug0D5I1l7KvhsnCLQ3vh0L++
TipMnjK/gtovr2EJFcjjSygdArqJ1UuBpITmg+e4QMLFiDhrLQGNWyzlRulV51/t8+ocISGLZAGU
ZXAT0ppUzPhmmHNnFFdsLsjB2/1+lkIKylFS0ZcARHR40WNDkNzBVu+R6htg+enUFu9Cj2WgH0Ld
IHYc7ahbQq7yyLLv9LnAB//c1l21DTNA8M3ihG/LYYSmsuA/lRDPVPgDI67D13nXf7Vnz0GfU8yT
EImIbd0W4alM/e8c7/OSjn3Gh7XBNiQJcRP91HJxtx09wWqm7VWQcuP0VCjOMNE7lhoy6QA5glDb
WinCnGaBjcR4YfXYKyHRK9g3lb+gZ8NZKnWuBfeD6/bUSNendcPpwMZGGlccnY3qjO5nEKuw8Aeh
4jX9J8xjIa5zJW8tR/fU845dg3s74+zLflEyd3kyRhTgI8L8Fp78xKxHk8N/dmq+iLR6m2cd1syl
qaiIT26Lgj4byu0ZlpN+8RY5LSF6AfRgnMdwehVtvlT/GCUCvI8YR/aUcCKy9inPFlJ5w2OLuzPR
578ZXCFj2VgAnJb/o5pqtMjVF+JNgPDp4uHtpq0xMJtVKijlq5cwaBpL4DroSrWza6lBqJi9fQVl
3GAQeTtxd7hT9oM5gCz9hpBdTOlwAZ6nr0w8wJs/xCYBo0kuV0Pgv8Bxs0t1a5LJzrVHr4vncDUb
+BRScUolnzt4tm1IIbrHa4eLofn+4imCHjQ8epa/ZZb/ogz9/FKv8ecIftYqzLuCSfaIsuVgBf18
5CaRsdXhPvjZ8eSwczLthNaDkBX+YbfZc7EU7b43VNzDybH9kKUBva5xn4AvE19hun7AHCruRdKg
f8QlhvQBQ2RBE4YuhX2hSao7oacnfhfCUb9iLajx6FSuAymvgrsKVyc5JkrTeP5TvrthkwqyQIR/
uwITxOQau/cXEZr5+E45D2YycRnjz45JIVJSFvJPThujzqvC15Exkrg/VkBlGGsyUyt9iWsGGOSb
8w3txo7fDuVox4KT0fpYc9b7QoxGqj/pZZfVd1jvFV2UDa8HUNjx+B2bzc1bTjCqrfebZOsFlsn7
2ti9qmKA4mu1a10CuSc5aV72aruStxLF2sDAT2DrHEOdmO5OCwYEouSRtwb+IXgCPyt55n75Ke17
L1WmJ7gro//gPkgjlC741+gA7kq1D7VB/Ddefy4Cs/kZ9nOHFJ8SEW59eEMtQy4xrYEK/n04lkT5
UsCjupz3udC4/Hh0KYRXHwu149I1qGg8BzuNdSBbm6BL+9XD4wU6G7UsvcoXJvpY6U5OoHvY4UTt
SwLdi4P7lBtyb3UQvXN4hxU8wvUZPbsXX+w8fE+hHfGcB0ULsS8Kgr5B6pZmT98VCq5yDTY0Z2AR
QG18dNFojPNkOG1ZrDOxTiC3XhjaLGfovHJ+/ucXLTKmKzwu6rJx+1gHgbc6QXs5rBtL+11xMZGz
7O2hedQ2Th9ieCuuthqthuTiG6fSQIjCRrpgSlKV4cPc7kZC5/Ml9V6fm8Vq5gk/yt3rUHWOcrNT
7ZLCaBh8HqaPmXTqAhbQtNQfTr2VRd6RaUqOyDS0UoswsgRwl8HEqECeQsJiz1xsDvuQ78/GTM5L
RU07EogJVRQjogoK40DPsfwVwq6lpt5uiZfqABG33YFd32fKWa+REab1QWfl6bktrjrvvkmzm3/W
Lc1faWDZ8A7itFQcOYvRJgcbnDbQPs9oyFr//xkaamYPs4wAi6OAm0O1U9hTwciydnIZGm9hGMT4
6zg+mg4a0D457HhJpTRQYZgMwzvs5fpP7zJMIIlWNP5/nZrp2Kiy+l8ydq+qJlfj+Z23PVrr5Y4y
QlKkxAYY4sq/r0pM3kcWqCAQL0s1Bi7KHF0YVt6juQlX6Eh09n/Shs5DbS5LxbLrjbScsDRE61bQ
PIPKpkwFHpWOiNZlHEUVm+HuYVLFaBnBjleOFrxBXE43CPZgw4swOnbcxPQjjHsYJQyEbelxNr/w
n6eFrNYqmm3mvvWsPkyKakB3AazH9xe8kh3Uzg5+efy+uLijIDYVxNyEpYu23X0guJL8lS1lel8L
oK5ukmpxJSqgoE3y5g3ljJ8ZlrwwCvAoWDZxNEO/UkiZyZdt7EasJ+gDz2skAdl4XnqsGsnH62X/
p3VEBwco5owWuwYwYagF1yHFmF9Hvqc07XIDwImaAwY3dXKQfNdERzVQg4e5jxXDgctikvkNZPYM
5nuxKxoiERjjs5ObC+/shWREpyz5E5mt9AHm9GGKg81OmqtdboMPtPb59XPMVdOSloBS6RemnvA3
jXxgWb2F7+w4IfntaEx1NR4wMyfeCnm3aHC5QH00X6U8ithI3XEAC5NjgEI8UhSi356XbnA77Cjw
LBcZIzABASQOSXjsDDh9yigbKhEb9KFBq7g2sf8up/AmLtKuVlwP9mJrq5JkNc4PhoFZ7qwuaet4
xo5B6czWeLGWkuuHHIQF9+kjmxdk7OSOAdDmAi/AXCuh+4aiStW9kCTOfn8sBnXlMTjPpfcnPz2o
i9r/PShc6tcd9naDZ9eStcleHaq6Tgh8nlY+UgqYdoetY8ezY+rKIaCjjwLKTya2j8kgLTgGzS0o
pcEskjC2NZ9cCAf02rmLwSd/Pvo10LYNAsp2gYC9XjnQsfamgjxh75O1TNG6u0ULdq2/99cGVJGg
aqLdYMLzzzK+11VwZ/tGWRQO9eG3Xny6zwnnuBUhKI6NO54wXEYQvVuiL/GzmbKU7yqU0pcn/KXS
CgDNJNE5RQhtlbyf/b1IIj47k6xHnahmM7toJUQKoKo6j9zQ8gqclCDf1bWkh4YVDc/91MVKZN5c
hVHCRE1ySvLDa+jaNayO9r1TW/+jt86eutBgDh4wMLsDFqycYgoERQJ5y3sZ24oLtMwYzN/3XA8W
bS1GRNoex5cMlLmieeqPbgF4po9kOAB75qSrGp42x2ERKJDzqLUGYWeWbiXQCuhynqwT0cfIuqsL
sYMfisFRQ55BnT0DCEIBm7y0XDGeUrEAnZY++JZ3KMFZ+JIat4cqJO0zjODQOmpp9M3w+MNagdyW
0QwMWzPOqLslTWvYtfy7DGDWZ1EYjkwlGGGI4swACPU3Faq0tn4mYFiKLhRhDyfKtCDApIFIrC+X
Qm5+7AR5vbNbgkAxbnKCcdQUJ5n74BX6n1apLtjoZELeGzzCwxHiXR5fQFfbyPg1nUYJ/1VfgoJK
AcwLdvJLzSZFFpIMuzWDGf2qMM8whf2ApDplO+BgvWYOqmwUaJYT5v35/iD3kZ1AAll2HFjy4dfr
BolVni3UogLyyiPgfDLkbFRy1NN6QRuiC055HP12WCcuxaFUKDV2MdIB/NLTjYWV3beyd2Y/1Xv9
dKHmDWB9D7ZUlIRiNNdiSTv2kCNFUFHmAREZLKVh7+eo2bk294uvwPi/olAB3bTNNMDrRt5l7zr8
le/XZ1rB5TQVDBG9PCJgRHruPyHii24XE6NHhjWtXj27EopQIe5udO3E4R5pFYcjadD52mL/cbYR
5hlxDwveSrQfgg4BLRKlZuSOhpu6J0e+EsO0OVmMvKI6i/qQ3xE9btyzdfPyT5nzaFJRdp8+CkPV
+ik8RjwURWXzqWguFVaOghDTnvbdxD9DUY4JUhzjNeb0JQgF8i+dhHXRiqh56kTerGSjeplk35+a
cVW3rp4qoHzlKRsGT4qd5U5pM+50sJdR730L0aVHDxRurxHLtmSlIMRLCRg5ST1dFExYyQoxx63K
CCfSS4uhCgeROeRrBfEUO6T+HH3rCgjUVNdAZu1HpbdeJ8q+nU6xZQ8wL+LfJ7m1mg+NP7p0Q8zd
euXWFFbw4mQCd+H4626wVxImCdxfU+c0c4XzQeZ07JZNIPzVEktNzT2LHO2h4582p6w0dBbJeNoI
BKOepV0SbYqWcMw7A6nQIn/+8Pthe2LGPEWUlXis/XZ3cirY0VEjHq16GGVIHr6wTvJgLGvac7i9
R2pmQWGPEAniiApIYSIn/4DAv7wq7GkTPhs3k9QPEpClX7Cm8ADB2hvMhDLsJBr5g7fMpjCKBH3g
nyqOXC2+pWfP/k1Ru7T1O2eNA3xNE2ob9yg3f4OF2BQZEbVqD1ePG10HWMK2n9ZjAkcBmcSbkoMe
MIhvR8iHaxUHFq7Szs4Xj2sMKFg6KTz2z+DLzypuBE0xYDHMaCqpixqaP2lsc3LRze7NuNJ7AN7g
al/uZBnofM2gYIotlEtYezBFqVcL/NrDmISblsuerBAUZsvAQ9mIqUKE25naR2Jmx7rKUbbW04FT
JEo4CL297zepWkNwiuLkzJr+qVCjyBVjl18BLjcNl7j8WHrbFLRDV9yaezASl7DDh3Nm+7uKtVjL
/7VhLJqbIwxtzAmEjC42cchUKk0By9YmxVlido8JEZJX/PasLH61xFzYjC4+lJvEIPGty7Seg8Mw
/A1uT376Q5KsRjkMslCs2m8hSWEyX8Jm2h3m4DyejTunYWlmrbtxhsnFc/QY8T33XiZrBCnidQLZ
XGGFlPh7upRnpiQqf98K+l3icycrRIOIlKRFEv6OhzEB7Bd6LykM3AW3k/EbaUOj/QAQMfEXdC5o
o+tvrJdD6GnUBIjnRgazph+cRYrPGK6ffT91oCyGW/8u409X76k7WXhRRyk4qe15BW93N+gliXak
NJkZGL4lIBOpQWBlWRSAAcGfTvkNqxRL0rTN2Lm7dGYbKguw4PaUYpkXlbOQx2PW62RtN+qoq0Ak
+poiXBYu5RNzkWcIDnYZaBuVCdyVGnK1W5grRFYw/+DpejFekD3SbXSl5t9aVqrWOVZa3ExYZu3q
LJIBlMJom/pnt6uNHeuZx1ig9SpTGMwqnJzeVdCAlVpOXlTcYgS2Bxw91uxbJHZCW7L97gbc24IF
7wWIXVs7q3pPyidlnhdXTnPcrQDkSTF65/hfvaSQKMs0WZ9AwbdkHlu4d9fwFi6x+UcqH7DHrjpC
SqyG4Yhc6lsq2PLYNvevk3M5jvMlkAAsb/6BkNZfsdjAYyIgZIy2yGHxEvEupuh0jgiEH1GJixw8
23Pxj0VF13xD0rDLPyvksZzukmZ9HbXlVjBpeZ5iAZGxPFu7lsDCgk5tLoNuVE2lLUsRQcjt9osJ
sDR0dmvPAxEEEQ4AgZfTedY0vvZ905IyDBXrhJVzSounHwGqumRbKrXiMpfHmQPTDwko8ZZ24CZ2
wujzQcufBxYZTC3WEdY1QHXx/TRWxe4uNYWgDC9D5AWUeZxOSkrr2E32DzXlyauQc/qE6SFq5kmM
3I6WMgNfI7veAfNx93Hqdxtq7pVYaga7xgw6dont6x5OiM7mdsvJdTOu5vtAhbaw6LCfq5DyL1bp
zua7wTccpZlH0jI7t6lY0FIci+6MA1PhFmvViS3R5fpqxWp0GApvvQIkTbNdOCuFJ1Jd/bbMRYB7
eVHA3EQc2zVeTYnFwvmFou7S5XdZeRFfgiTyqbzN5CRqWhcnQeQjVo+d7810bIj/oLe4nVu9OLom
MnXbKvzfQUwMvO03fyg3Ri32gBhTAeV28fy1mpoAEhTUyIgl5WqTn4wgYWUU/4AjAocWgF9Vl5wy
RbAfBYRWkZ+lUOjj2GbyX4SsB8KOObXoZITphVjVeeCunLpM+btLWa5DeMhe6TWbqaEa51BdchaQ
MzBCy/ELPQWemuJrBDfUAmNVIB5KL0kYIvo6+VB+SjN5SjvlcPJOpouhWJaZQqesamyCqkMeorlx
yOCOdkW7NlkwCCNpR9kLr6SlcdSDAJ5dR0x6s1Oej9EbVzAaRXfRLCuS6CoCcPgLYv9AQaKe7fir
3Vp7MRmnikWYbHpsi9DnDjJ/ACJD3VCoww5uJkFpTcsMORNkJcwFbENZY4t4s20HwQAYACsSHEyo
0QAuh3Ev6FcEQxds1TQf6wdaikV6aaZt8f5CnXwsaOJrpvaFFxt3BH+Jjy1dMpn50PTQgfLQxYEf
C/0MbfFtIfHhLp4tHYA8PSU27slTkD7TYAObr0yQuBSsxdRPtejovMwpG1jbCkOP3y0OwY5g3jVG
yLzOIIWRQH3k2i4KJPOurHHmcxtAFx6WmXKL8B23UkMgZSXtaod6qBufAIYZxSG6AOhjfT3a9eXg
IJaRCf6xyBUM0EPqTu7VTtKZl8Yswcsf5y0Mg3DJuto7CX8g0DLpO2gzIeuYXwV6yjNus35+W2nz
Kt7IRtIdKOQ+bfenBsZUHiL9XIM43xFiOpDGzAvkXL6xtPHORLP5KEFA2FSiUpKp8U8y0Fb2A+xL
Rq2HubP/sXaS0tqoq4N2UjLE6FnRRlwyVwbF+j/EKC2vUN8WS/fXiQ0oD0JnwnYpCVtGbffh7nIN
+KItLl7oSflR1XNVqHC5hREIxLNpJ/y+itYrNhfcYYqTr40scrqAPlPhAb3b+ic0/bSmw2lUq1Mx
aEVupMmC5QF8dvC9jb7M25WCDVDNu4TRTm5mLYxiz79vuxAKDn80vsHCz334hbm2UVFvoggQOs+L
aeLkM0wXgQorNIvVmKt98EsitC1N/i/The21px2/nch4DudBvBA9jCVzuyn/b3xrE33p03oQHhhN
jrqBgjMeK5cxErXyZPuyrPokp+qQMFOdDe8rEmrMRPSOV59XBX7rgLIzeUEwc5HVMOfMfXUey5Jx
84TZ1RQ1f86tqfmVJHKkgOuDqOyKSeJNEkUmUxpkyiWuXUPmIQZ1HFHfk8z8hkRjXP8Bi6XOExeY
JoG1SD/7Y8kCf6sOwmaYSrd7v81InxpqwmNZNEMr37K86EowluKTjMtd9Ltu3HbmHQPU99aOx2IL
q7l7kZqRNk0tE1w/r7tm2DcOUZx4TsOuyz8AFofLJ0JKaOqQQUmnS4Jv5XeCoUjwyS/v4hsDfZTu
4WZMSJGhQTlvFpvZ0YDRAYhWUgeJtMC0/6g9z5FNAgiiyBUHQqf3x0TL4K/RwWxdXp2QwxEsa8VH
SjOcS1wE1yh2rwcGM+y8PZ3L3A4ztIFj+IHAZ9SEMNuYHWizhXVSfHzPsVxHL1JZ17MNapUkOxRi
Q5lEj3puek+bygu3Ggz2/y6u4D0JTMhiMV5ZHgvHu7FnE4z4851T0zNGpJfs2X5w+UEBaMxU2FiY
a8gYJ14RFsCeHtIOHDbU+IaqtIUThNqZOTIvw2LZwHPedi46r/RfwtbiugjUyzRqJl0r6VPPGpMn
fuahnTZkiH4wBu183p6Uf2hYoAdz4r+e9RjbWETVvcJ+/r9qAPZu9pLOQisOujWl3P7B1Ra3opyd
LOrYC6OQrQhjPcxiSw5wleVQuNKprd8PP+thOMnN+NV9hIYeq6LqsyM1+yrO8opGfclnDH75FIgz
3x56gLdCJjPR5Jhej5hYRRmr/Q/RJ5PIkKq5+qAMRUk6vcKnfincWe0ZNhlEuryAySaSwpc99Scw
Tb9ljgKctkNlw1CIR434FE9sB6V0eMif5cJedY4qFw6X38kzFQh8HbHkk8xH8oMWjED2h6ZU20zk
xRozusIpoD5B+fxqx6s+0tydLHTUGMrBMv0WNckSb0rtEP2OvIy3vmsOsP9h8i3McgbMdMbM79WA
PMopGqJ1w0CbZ58yUCwt1Ajeks2u2DyAWfif+s6mRzrlwiZHJg6PDAcc1qxIJpoFnCkCvuu6N+5S
lKiv8FCTjVvUvv8xta7C4+bPOiLqCL7cRm+nL4ELmBNGvn24W9CCgoX7I3InVk+KrtW8hYxu5IS3
SkAMToj1iBzRdc0WHbz5vtEnrFZB7iSUv85AHmGGryLt3RDaruHtRFDPwoouibik/4q70ChuDHfH
hqJVUQ9mhNspneCdkhy8cXNpm2g0lUQUrvZDmg+4x+uzIT5KdZ5qNgy2D8MS1HESizBDc8ibb1IE
cFSq8ydpWVngcADGHVf9HDbhdcV8wMMt0U5DI56v9YJ07TCIZumiQ05cViiuPJGyILnGBvwNF1Jv
Db5pqn/H8Tyt5+dHkwtkMUFjKVTtGkBfjHfum1/0Lg0h8G8zfdF0n1skqCHka9hJjsbrA71wSTI2
/6tYX2NMRllDb5plKKCWeUtSfvhrGE5cNjhRlrlHeKzSM75+YdfJUk1/s146pe/3DzHbWDXm7eFn
+64b/vFfPenrGh9nwLAVPgKpoSH93df0Pet70v6/3GXwz5pS3UcTFgyCJ+dStfjcYoYjRY4vjw6y
4fEiwVeIGyC3CrhP6r9Ezlx2ZRMdWtwusaPCJ5VPol84066ldsMmntKiSu3zuzCWhV71HOeRVqag
w1EI34Za0X4SpkYQvZuTMuHSUvh8pLht6E00aU3gKH3vQImi471gc7ZbeqkF26dvV3QT9hjnyYoS
Gqr4ZI3PDt6W/eRNC7ZOh9UlQEzpm2HiMJ8j8xBxZAiKVfUZtPDKO2AsAvnPSL0LMgH6/wCgJENe
tyZ81hOm5xsftVeVWnjvt0CuyZ04V2VRsomczmyLq/AU3SZMQTiVkGrdye8NhuyuQgN68RIqFXwm
LEPlQUY61nkbAGEMm92TsMHuoHZSyAkpofhrTgiwT8jBRIrnQ5yf3rd68Bljn2uj+3uiLtt96dD5
r7dZjxtiSe5CDYTGocWo+u0uib16/mMhrat/Nff44bF0sqqCK6H71n9Wl+iL5bO4aOZLRUHJuVA1
oWPfE6Y5lI3IbVUTItTRP5B6dHkS31eRdio+tam9FM+h8RXXc/QcNv4BFXtVcznJgTDLOaHecIG9
HDYhoZZqZsjCkKzUqJG1tTtybszRu7+tjhiwghbyNIE80fyG4sOE9aiHj96hn4NVowg6K9edAWwq
DDdrHSYbbYA6VhW9Gp2u516BE3v0zem1cTs3WoMBfjyAvnnIAzMLu7c0yRqZPO3EPfCAhDGIwq0S
iDT2zUV7yYMsZVMvnDTT6OqbHXM9eOnlzFpv/VGUoGOK5i2189e8OsvObil2DqAeRWDFG6I5hJ3i
vfQvttLPclastkcFC+37ijLEatyoiJUvulrs9V19gOqGlurlPz/2vc3M02Cgppz/vzrQWYZrn4V5
Adpp4eq+RonWbar7+zQ7eLXu7EJhfcZXbc+ro9zDnCxSbMICT05k9ETS8Nd+hky3QhKEcyrWG8JR
3E7ecjGlfH9SrL6Q4pdlMTzsb8e6UBy2snpEEgg+6pzrOtxlHGid6/3NBABicM+gGtW4TmdW7Q/q
P2+8oOs4DlGB27FVhMXNMOD1cNEItL0kifSDEr1Zwejj+UgVW5HO8Grdt3AidboB1tMhAYxgBcr2
iKD5aOhBBMAUW7ye9DvApzVIomitYhaMUAFFYBb7ppusqj9XrB80jcARm/KpeZwxd3Mc0x8ytf/2
6aIpLPnRBEqllSwr1vdJyi8lmhA7vClV891ffdkfrCDcjLbEiP+4PUmdB3s+v8KlRxmgm4UDsdes
/EYWqXPXx5yZkEXIMTxtwlBsBHzXWufIKAbDJzEAfsOcy8pNZrfqw0iwOI0TKBXyMjVqzCwIePHW
IhK9d6ZGpO0BzixafV+zP0oshqvEChsfy2B+XkO4/ZjU7BJSVr0ETn5VPx5QPGEMNkKV8WyJabyU
rpvQMl630W2LrLrLD9VVn4RYkFJBz/CuJjunQZFOh8exZupszquThugWuXlSIzNpEPyUYz7BMG4l
kMQaeey79LU2N4NlxJopZzob6CC+MINUf2hS7Nz8U/C75q6PhnGfK2ceTXYWO5CCskWfCoodDBw3
OfYHex56+jULfPjkW0sNvHF6T+NOQjxeKbwEAQt406bP4QAknKQovBtBpjxrixr3dEcZqktNc8mY
aThbrJ06GqZnywzJOR8X+E9YfuM3L2+lD79l9sU2JV1jL0g2dR7IjpMjHina8bDM5GGcqMPu3U58
qwHsQLriTA/PITrc2HxjTwXujfXv5zxmiN0D/8J0pltR+w96lE+Ngt+q/+c9l9Cp/fP1/5aA2vj7
0rRvlIRVTGhf64uxKIvlrNmj7HaPCVsnOuSZMExdqyW32gldevHa1wuj4Mrj34h6kfwK5SembAEz
wgGUPAawqHB7nTU9WwatcKNhUqZCYniamdJRhLHOuiwDvP70e0f1qEls261gdynCC4Xm+UVrbpfd
+ZtxzHJgwMX4UERXHqOj13XXGQY83YHV4bpRhl2aWIQJf8AA6qhqgn0r1PQQ5+jPvIcJTWObLgmJ
QVVAV6+bfE72EkcA+AP8b9xCJNzJmmZDDB55byPWeWM1psqzaoD+HdSRI4X28yoz9lLCa8PcZ1qx
UY+HzLfvFT0JWmE77VwXGCn4Z5X++vUSDUaUyU8sCJxlXEslY/b5aIqHPHdmejeSAdEGRzvHbTUs
R+k/wH08uqCbTg0YghAj3LmOEekqaQmzYqnajqjSJ94O0cT0z5FqPSS28fApjDgLm10CpynHxu2O
YD/QHQCyYVgftsOgF7cJNumZtY95BM22P8i6fRsGFfnwOUcr253BAV/O+0olR3a6ZzG8SE823Dge
HDl5H/Cs/Mtb1Zg25aHMLnO7EnEQFLT38Pe7OLvh2XJpx+MBcdxJ2DR5gNkip5yE9OuVyVQPLxjy
6vqgVuB+i3ORt5J/rQV6oFOAyLi3qi9s2A0rIse2ql3Ka+1/WuUOam8l7FY13KZrPO5eNvAfhoYI
xCHd9h+yaiomrorOO/3Zgv3pxWG/BEaK8GwgN3kyjVzrGLnswAvItRs6/m/WchQZBobtdMbAa9kc
tLxF1pZ0eK155MkkdjtRkYO8fbfamqJZu7om5p8dBL0RgGeU+U9V7utJXw8V4E9XP4pK0Vax4qzn
HN77wEEeY5MvwO9UbOTW4mFVNHuY1pNc8EgUtAMMrIKgccCu57niHgQvSugoYaIQevV2g2G//7al
2ETX+iWCkALd6ZozA7nJCpJlsgNJ9k++7OOypudNh6n9p+TFkxOcGKKQ3jZRpoY6i31zONq0pMMb
nlCWINicOHyv6f42mek/lUmwVTNDfIk0khi1ILR7Hq+4f/WrpaTX8VfAB4wZzNtVsEOUiFOjHNq5
c21UVYZD2IzAuhfWx6u7wJkrF3HMZ1hof8EIaY1jp1VE6Z9dWcKv2o/EcpCXdrwFGUE8WdI4ga4G
cQT6RTsoa79QAUSvlCaHLf6ULDU8aH7ec4Y74hnFIlyc50gvmIg7TZFEYqIT55R1cT3ELgXRntcd
LOiefD9ma69MN3qyWjwmzq1MqAzCFBp2ZHRQOJhp72c+gJ5Ar/cWYeHAfvfseK4uXqhZ1JoslVqy
cAea6rpcSvolWaErXuP/bsI9lDRXt3bVXJ1752aJDSCqP0sy0So1jSIV/H9XQsC0yw6/pNu0C9QH
yAohg4IZxv5Qxjc2SLLdEPee4g2F+5sfU8CMvSy7PwHlpw2ngttpU8ixJJOaAyA3fX/lQ8SAaghs
EZhz3bfAQOuqJUn2DW1CMl4lH8Hmwkgi4Fv9b3j2N6iERpTh5qXV5fitFbjLaJ5h7T+8cYvez59j
nLgYQK+uQZ8vdCCoXELmhsVSSm1wQfR4V9DcgZEudjqv+ChN8CVP7nr6UhI1Wu31K4QWdxpLeIUl
+GK074314OM63lcyIzY7kPIbU+rSmkKDSYc6I2oGA5bOc0/vRCRJR2i4yqCoS/53XbT8Uzlxp1UR
/KtL98e8hjJWpIBw8Nt8Varyc7VpYOa10WcB8HtIaGYg5i0UUtLZSajIgopQhSkZFNMIsHBzZxz+
4qUhfOCLLsoTneo14dpb41kJdRL8PYFJjXLaiTSe8noUsYbl5sFrB0FKof+evs0j5pi4CN1DIatb
tqjme9IaxevN5HDt2kfkIDsQVp83V48JVfFZVkRDIDHMHU3pFH3i/JFw14jEQMDZDE8l0bSQxIQY
jf8F/h246nn1kkN9OibbEFL+qdQd/UQkiJEy8XKM4E45p9VdMLdeODJtWjwO0FqU2zYFsnG6day8
WYeHPA+PPQleryJLHYxctS7HxUBRSpgKB/T9ukkxKTFB4JLQIhPTL/HWKUZzJas7OL5phB0J34aU
eJJ7GYGdVmt7Ej90MCeDjqGDve5Eu7jzI2aUV1NF9UUGaD4E64jgXdk3py8IJ35SuJwMp+pRKY90
V46gDIGZcWzW6AqYXZMFCdUo+HD7GbL6CiphhFIRBQItfPcIflRTtRVNtxkIwZy5wjpI3ZMRkw+d
quevT2vP4G1g6enqKLoXkKl9KUWVJoEB984Q42rb7RnzPSI/ENN/HIMgrfP8kcO4Ziq4B5m5e90r
ELwRR/4lPGahqUpEpETz+kEJ4WgmKZ4eCE/USjP5Faj/KtUL8JukQiywTI1r8Ta6+d1Zdfnfm7Xo
XbRP+2CPu9pKaqYKJHvx0F0xik4OdueK+rK6vMhsdBUhmjitCar0XT/Alxlvgp/2G2ZxwD6Muafs
M2VBt4ToEHrN84lg4OrpLGsNkLgR046yNZL4zoqL4cvCI1qVvKgXbM6MTAAg4Zt1ISud4+J3oeyh
1ofuaeYrowETZywAWGAcCsOHRPLxH87nxFurbuua2sK94qWjnsXynsoJL0rc5WQqvdVWDcdIjfkd
xYY3RMGAPi4bxc6lyUWiixMNf/+m4pu6eiqnv0eQGDS2ktvNVIK1HK3KeyCCJGsOfrKVnX+y4mSG
sK7uhQr07YbzuJx4p5f8OGMD4ehqaxmCXX4Jzuxd9OdLC7ttsp/iRhJDK4o6wDvXgkFaXaS+yJB7
X5yilH8NWmljVxGF2OBx7Hpdm8SIwrd2cDLGlG5D453R17glbX7JGDxl85CtugEFBvzufgtrKTBe
+sO+SaaT/UfLewj4WbNtdbyfZVJfJ/A3zuYusrWxEbw8Tde0+64lfLIR67GFA6ffVth6v9VsJ9LU
0SnyM9VwFc++O0EAO0miwoZSTYBeo6tqD+GoB6sy8M2GM6E1Rc5cAgPeDvOTF+VGIx+HJ1ap/u+W
7viGBzw0SHJOexQC3Njj8J/ZlYLTxyzYJIGAomYof3VeVbptRwAne+cwXZzvvvhl212xMeMNplZY
Z+VcnjajitiBoMXN+iLQ1vvEIM34HJNFogg3l0HyRHLXtUDEpKp+ZhH3K2AKH5g5ZIE1Fo2CjDh6
qhfxinHY36FqqBe32393kR1VHnK6d1ubw0TSX1uPxtSQo31CPfK1NDmyBWnj9DgCbJhK7PCbvU/d
9MRZXaA+EQJmPe2pTicKIrk2iFWo0HTLI3ue4xREPBgG55vMYKKCmtEfOLO+SvpQOJw1rPid6yID
lHiT0bi5vAc99fXcWA0dChKBqvz4yS0y2tG/sgPoV1VbRT62zgZrsISvR3QqX+YjJWYHgcuLu3x4
jyPNOGOu81ZQ8ihf3DRAlkNrDgq1dN6lTfKSATBLJ4H1Q8/+mc3kclsHHb6qdWfdVxjE0xc/yK34
7pwuZGtMEQpTsg6vovuvS6Wq0t8fb75Rb4pyZXgBOzzMgJtuZfUFyGr4EJiA7j35wUG6M4/7MDJ0
FIBp7e0Wv5jTV7fzfVznQstr0nO5BmIWv91M0YaJNczzXPOdn+zEF8otzk8sM7z2dUMjl7e5igaZ
ux2ZmXuPBSykebXBCoKBkKexS3TQw0+h/yW2YEPVC2r1CqPBVXrWa+ofi3kMAI0Nu4dUDVSZNxf9
5KM9FSD4F986J+mjCbCKwoKOwc4JsNpUPWnATIKqlZ62Qz2u3XVUNLq0vexIpgdtdzCPfcQTpnhj
tI9ZDLFpmec5MbDnLdGpSCtdOjgTLgBFtVyd0J5Abd7V3lOg0mGALUEeuwzLehmGOd//zKhFXs51
YwRGEjDLx0+OFQcpa9LNgrSn6KP68F5B8fDUL/NqyVtC3mbd5evtP919Psbdx5s7UsPJsbxPgN3o
HY4r4HStdAXDMoMYCloSDxbrhe+CgPXWBjBtOb5EJyeZjh/NI/o/jOLWj8M/gH/4PfWIsIa/Wc2/
4IyeIwRVljC9cqZBTJ0S42Aap+3WqMJWxA2CrrQio0U/ZNuNNouQN3lZW3wNDqPil772YeYoT0jy
UAzP28pDolmTkwHgGdkf9cEqDsSpzjqftOq2ubmKyj+G9Zbla6uUall+uuaK4je28PyPJfYkPY/q
9FwWjtQOq+XpRZtaIh9uKyAscTExOXL1Cho6d6XxPyH1+v48VD0mRSGXICbqzOMtfGgqSGVc/vaW
r4KdbcelvaWzxVFE+LnH74lCWpW++Km1GE5QKyFUTwLzGjsP8USeuxj/6EdXOY51YQj/9BQUYIRy
e15LujojrUCU/uU16v39TtFvzg1lKKV8O5XaVq3Ji3me9tzHcIVVbtvffuhlplTdkJzzJ6EdbAiX
WwR2KDJYNxW+F1Pi+TWOOYv0elOWDSUGkgke8fvuottrTzndE/DTiiiwNqXJtuhp0pvMcswwKG+b
A87E20mBbmZkhWfBGrq522m53mpeIXo2vongQb1kaItPi6zEkC1yiwYLJ0CvhD97vT01dOGvCGwR
MERCzYFosSSiMtx2nrPQWNFQebT0EFL1njQfGRrk0bC5EgkJ+PGYHG1gooxaoSwOtV6WAqjBqTi2
/DMoeS/CkKEEtrqk3kg/KjBVhvc8waZlKZ8BxFcfk1nSITAPNCbxpNvzBX+xvkgdQigF3nIbqC0P
kpDMqwmr9mF041UN8mcdsvY62njaZGKOepAb8/0GoJIQ1OjKXPNg3NAMMf/KdZirNG2iRC/yT80z
itrW7gswiMgwAFuu8fFLIPWn/fC00u+5S9vlDpzPtOsZD2JfdPixeDVJnzQUMQJIGdRA1ft1F30Z
1xIyUp6YiiM2+Qe+hqQ5v3BT7NbXAF8QfrhOiVB1FbZ3Oa4H7DYALtW0FZNw2fXXwBpO93qC25iK
pCuK7N+rnYorcoLn5scIvOr/EkNJsD3kLkdquQo2oyEEF9hbB2FF6FBPkp9Ei+hdAQmkQtK8c7oz
gV9Erwd2cp3PCrIe9xQVtVQF1FWEv4GtnIprV8kZ+f1k7TbDF5I8nqzYr5BQRG4TNogX+9Eswdhy
4e3dKF+OK0cDStGGqoIIcxRI+hi1Rw9WJ+xiXFmdIrFtX18hxR3gOhLB6EmwzvRYOjWGsvmoKZ7e
T+iu9VwsMAPEFh5aZ1Dv/LK57wALvQiMN/alOim33oTlhQh2c7h3Qx1iBA6WXaTVA31qHb08Gsuh
HpOK6aLp3pN1biXcm6YRAqQKAsByw3pPBkpX2Sd+LaciXjD7DkhJqP66U42wM9knt+ZcgM5zhVUX
XfURJDucBbFVIxKhFJHnVmJnCDsEkm5XJk9mZpA8Luf4dKHnEd31Ns86uLfSSgvs/QatK8L5DFCY
K7mBusH4WFZkYd0lgsmk0FnI2k98tjG3sCw30H5HTpmdQGjuC4+AOrJTvdoYca/ElCtpDZ6kH6pg
Za7kVVoG4R/sNCG0DRDGbD2eo3e44aea/wF3s6oDGDdY1lIjdtAmqtAqA1IdHmUkt9nTnE2zIEmk
j2TZYy1g+RRpeltKxcnmZXDRHI4wbGvymOcKNviYuXp9e7SpLi/zhy6O3W+8o494lql5/CidYsJr
u2hvEkx9N7wmnSih3O/8J/0y5PoDjsuJM90b1yv96G6kVSSv6WdjfamIuZOgmnLFEMTzimMu+C8L
wr1kGLQyVZoTWDadd9zoNuWp/cRFjcDPKhx9+mEFRKrBeHHMlpMzJOzy/Te32YMnjYblsqJirgnL
1pQfgWAU8YYrJw9HmwH8morCwfvY/V45+7ggYMvrcBza4Gt5NWsr6qnDoyRSoHANKWHa1/75vT4t
xowBww7b+Ii1ZC7sIF6cZ69C1PKWgAQHjg8Uuzyse34yJ5Qmm+EjU8E6aFv9hqdsVyGBvsA6U8Ov
DlBiVpC8Ao+groGxOOfypWEPT2cE35nCpRxReTNq+X2WPXDQvMZO9DLHqo+AvUY9xivipCxH0py8
kTTTSbJMEK7aqOZngJJutzd9CAzBquj4hMmPo+U0Jan/LXFISvvuBvG+HLxatu8eHcVzfuMU/7p2
FeusiuRF7JbCu56azbN1coOoY4PhZPlGUPbJdWKspv16NqKzNpYd1wdGcCoxlUGt3ZZc2l0hrmo7
s97mY8uq8MqUTbQyZQq0AomVhmb3Q9p6m5VSELCq16vQR/WDwUMgYQd/XNY9SlCGHZXQMA8tfJDh
x8K6FBDv6q+/LW/AKowwvscVAsmys9hI0Ietg7fYVmLJ7yP7snBlKd+/LUR2VEdx0jBS89RjgP0D
d9enl4S+czdlUjnDNPihhUeV0gp4gmroklh0HpCCIMrTi+rEoR3lQeodzPcZt7jeIycsPWwOKhps
+3q0dCpxSXOHrrqofKO/ohtm42n8x1RZqbTtc0nFLNBNhePYDcvaV8uO0+JEOQMKNznUwuNt7+1U
LC9Y5WS8+Pye4O4B+farQSrdCjODfCy9kb+jonVGDT4r5MkrPmJpQGoJ+0z0x9wZ0jt7PcxiUvFG
Wm8mJlT5XE2PGCT9+SXU1NCS8CNeb7dUTou8FMLggzhSKtFKvwTaeaCjvGzYRqSDHAk6+st6bDKZ
mu4AmEEheRToV/WLE0qx3QSbv0fmM6uq5ZsQWvQGod4M3alH+UlEJCicfBq+v9SOtMh3zqupwLlM
ipUyribW+400PpiMC+H5uiRtqZy1fzF6tjF/uJ3u1pUeD3vIiljtBdMbYO4ezVRL2C+jgLE6z+0u
BmfMz7LUwv1/0Iw/lWeRPdl8vPdrgr2CsLdkRc7dKXZu0YWNMKtGAZe4zL1hLYLlPRZ6X8BmR0qS
Y0w81UukzIQYiZdHJmPSZ4XtILKOmXBAqf36kUTwTaLY+CJceL1XJXKfZTFl01gJegc9qlvD8gY0
QGWKeSz6vuUBYktTXF7cjBPeeAJ2gOHDPZ+eQjMF9XcTluPuXB+DKhazsWpUmBZvhp5eTcCq1dW+
RQLW6yLPlAcgLSiyB+AQRHW2R4WC2OqXkOn89UBVB8Eq5tkP7JBZY0g4typfsp9B5SqkDDd0qw50
xIYZXzoGhfyr4nc3Nj5G0+FPoxWx+VD52FSkkf9TvGoBs4W3NnxIDDSpsTCOSYNw19mH4ATYvgMP
WZnTIL0rOsPpozDdZp4f+HR5k5zkFZue423evvxq2Ukau6SkcdVkE/7BEwAP3CrMaQU/33hBOMXw
SGwsOOMVjOCip4bX3jc0+ZGWQYgWLssCzLwk8862mAp+SpsqkQkLpSDWOs407tqidNjzXyoT6lAu
QSZ0Qr4gS7qq1mNGY8WDexjquWAfwPrXlqkHWHZwSvFxZ/afT4Yq3GcBjMmL8Ew76uin6eoy2G/x
GyYtUy++ff7PzIHFhmFs8jvmQ/rMZdhpKbTjA0xoatkcpFW1HaQqQANbCozdlfP12W5LmLXHsBON
VvxBXDANBXNEG8UNYUxQ4CokBF0aHmtFet4uHTVEvNhOspSznekSK+GBCcYXtwwIDHPq6iYOv3/u
QywawIR/VpICflwTM8MG6JismLMbqL1Sw7RhUpKsRdA22sAKTQ5BctRMcOoCV1ulevwMlYH9V87Q
kLY3vGu9pdMyS9P/nRrp9ueDPUKe7Puj+LEVafdYhCo6L4OEoYePNGG7qGvVQg8c0tI4g3RoNayW
+sxiJO1DnkSDSf54XHhBqB6eLipzwfKQlRVyIMnB2xIiFOOtmY2VtR4PWxkE3/YjAN7HHfYg8fZz
lo1vKfwk9nPjeyXQa8Pm5G7+RM7Mk6SkgrciVE5NTmgqU/d8Xl/JwCnOPLms4bvIzY5MjLg+38tk
8pPy+AmjzJlh83VCoVEcy5ONe+6Y7+zaz2rVv290nH2QhIb9Kby/JRtyFepHbNWuXcUq+tgroRdY
hcdMcBAu/MTqmmgXI8ufz/vx5NP9oVtwMj1aCnh1OWiu9bYNVTjkZA9sNjfBgbqKhDyyme3c2TA1
lIGaB04/aTnc7G8MJjlO4NjnqER5iyaIGhceijwCYpT73B+PQj3gulD5FIATR3AHvpwH+eVdGxK0
pZSvsmjRrWQDuaYiGrit6UgqRahEml+lzclW+vj5YEc4nH0EKBTIB3PXu50UJChiPSKn0YWTfASe
XJEIag6pXm6r2Ej5wXIXZdhBgx2HVIeuKlzvg6DnAboooyhQ1y9C1VPxCuCkk9m/0klC2wDAQA6I
5XhV5UscSKuFoGmyCo8ouOZ1132w5c1BVIsUhx0EZ7O3krne60tKOavhSZk7lM+GauZjnULJAhgn
ZuqyhGWlm8yBIAz7DMeAi5y4KlVsbJyYTKNghlGW0D3T1yrWlg98mPGzpkoXZqUt5xnYKpMR7VTk
ostyE4jzr5EtHkqpNza+TAzKTpjIsSEXQiItKqdeJZO/eFlCCjnntZTwzYgzMRuiyym8s8jfv8op
f7enlUbh2ViJNbl0VHAu40T6YPHI/pIDSM/Vy5Drj7TlWG1JT1Wa582zXMccuhVBOczrUr+fJCIK
loHsh328NhhzcRUgZ458TQlvJouYiq/lJhhuqF1sXkDXOdpVwZ1YwJG1oBukv+KQQzaMRpDovsSI
KAXgF8eK6VZw1vZNwIPeNpMck8Xx0MpbX/8TjhRELyeQuo2EpyT7MsAZpLhAUUK8GDqgK03FYbc8
KX7qGB4WGbkTzOicauq0sgp2BgS4ThqmahTfyr8ClAkvnQ5pJcxh+xvm3YCN5aS/VyemMz9bTdoa
357vz7XiGU72dDxfpVgJU1ObLxtgOK1pptlmgsmNZ1TYrT8ceZ6JGpmqjfGjlNA1Da3k9sDGCRHk
6Lxz+ZNCxibnnaAkssajpKlnXII4AmVgqDMLFm5bYB85bkN3k5PXtPRffw9XQz39PABPFgBxG/cd
U40HSYoIFfPqZwae6/mfLNPCN+07vea3oRnj+Anmsj1Pu6rP1/dFo+7RI15nG+OqmBqkNqD0sn8/
IOlK7vrgTyfxRaoS0iu/FL916xRUtwQi5EUlyuY6V+nBTXsA9qaq5AdS9urQ28w6YIbCzuh9PDSX
vprmBnzBNVKxEbTDuUi8qIoqFuzcEYWms2xORh+YRrJXhV2qYyNY5RBgeT4DFS4mjtFbRCy/yaAp
t9zBUuZtcSEqmVOxX28hZXm5RIbDcPO3emzKEiCH6kdArvkAh1hp8p2vLskKqBKmafX/KzNnIgTx
DQ61u6Y4jpkU1vLRcdUflStu6HUHWijrPf6GByI5gdvAieMtdaE0gF1WBE4GuSm0lJzVc653z169
oOvseFM5mcdQ9cGvKy/feqwo4Zh2zVjkHfTs9B69yOmPf2Aq0F9GIhqEK6kOHYowiqnvpMYcA1LH
4X+m48tDOLKlqJau9d1TUvwWZP9FVIe+4iEBeFutNh5QXGVweTq2pCxrOZ6PQX6acuE6VM+EgmbO
TF1Xe2R2ckiS7xKlerMu+HC2yNkCVLOTiO9lSPuMKYJz1pwRBxg375whJmstnTziYYy9zzFyh4Wl
jFek8A1Yv/IFrGuKWFozwfTxMqKy8c+WtLEgf6A/W74EILaC6CgfILMoo8bO8UWfUVFT6y/IiIz/
MON5FVKa/C72h986BJaLbSCj1XHlrNfM5yDqoHq4wtxoug0X92u5qS7ZC1lztUFLDRrni5Vc3MIQ
tI8k2cBZaD3p822Z0fM9EwHK7OUPiYfFhEBQnLOZRbY0wkqmeibqb/9o5hTgm9py2lcmFahCNegx
zXdE7a6WWy0CRQ1r9Usum0HDUuY/2FdW0y/mILedJdr/RTOO1l8rWtADIaoN/WPUzUbyYpfur7tY
GI7aIcXxuB5bShLUtdKIsqtP5IzKPCxIbzgNyKx39X9DD/YBD2JYn10uhsCAJ/yj/7umUuDWKNRJ
kA3MCAZmJCcMfckxUU27hEOmiF2l6vol2C8FpNoG1+cumloZ3Sc5HEgSKu/03IhhVgDnpqjL35kN
znFL0cyOmCkKWvO0wkUWfEdJ+mCV1Eeaj0Zn/Tzqsg69jBmQFGSO8y73/1bjrr6JvcZ7YC2/Bkpp
Rw/PgA5/vVo3q4EEt5T5zGYRna7KMGTSJNOeS+7r1cj/6r6uL+77V8+hYSSciDV1zvKfWYycQN1o
oBGlHRnQvCOpr5/uXO7tBKbdX7RHHMGyKil2MEQXOrmEVRJhAMhUMW3c1Ug0ShHzGkNp6u+OCR+D
EdjJ1DKtSW0v20jPrt2IktxC98fJxxFJaDhJrHkBhXu0/TaP1bcGmVdyf+hFb8T8vjjkuRDBBG7D
reRbdDaL2JPM6C3X8LFYZc0fnPt32AyTjJ2wz9U5hQsSy44aQXH82Eie5hxpYciWJ+05391TF9md
zkfK8cpEXh1aJePhJbLgtBW5EhJzScP4LVjU3gyh5QZdr1DgE06fpy0hm/IqiQma2Q7axKx+crIE
2f4S2Gw8wZ3k96AS7aCxVw5uha/wwy70ZusNIq4Sr9HkOc9VxbQoFVrYozRbhpjqBIpj6vUim6tm
RNvZ9EWcnvKtb13ZaZcemLUPiPyou99P4CKlfyfLcGZsgJ17kBgSk7cWKlXKoLXvDOJrUD5Z89c0
aKJK060yms/lNpuTM4rgd7o5GRNQCnUz1U4uNrVWXawixpg37aAEuigOvYwZHwa0yMoZli8cKkUv
diWS/zpyoGp/mkBgaNIZRXqRHVf7w5CzrcdeTny/2lKUnzF0Y986+hHel945dQ98LhBLt6ljR0oU
1nm+lWcT7oP0njWxLAzp4qofaSErDIYz6Y2emx6GJXBNeaeH1W5FszRFzeWrEfJb9lQOrKxNf+lT
STK5srHNH/JAZsT7nZilAiftrN/yoouP04OhZ7WwysxlcbQqO/IrSYq1nkzuA1GaKpJQ5ZiJ6fqv
1iqZCvXNcTw84fGAiB0Isqns56+PhDXOsACqBgpI1MO110qzkpaTqd6MbxeXqW9XshsAJaw4yYkt
lq0moAdGak15X/XUwuOUW2QD499TzQxF+iK4JVXaTw3+q7vHbalk50408na5hlRM9AKpsy8N4Fym
UKz1Kle4E0AMIEnOJ3eX0FBz0bUdPkCD+lPQJzuf093Y/TfxuZz66E25knguw5gfZKtsi7cNhWGv
AmFtWYsNz2qbNlovejG6xGbN18GcDsF5S6BErdlGBmuMAGrbtQOJbkH7+7HRmbtz5O59+OkgRcwQ
uCuybzamqBoMBVqincRNRahb/DQR+7ABwct3mz/0fdG2HnXrrDGPfzLXUdHSPlI5Al56PaSk5dxg
CbVAm1adGi+156iFh9Dn02Z2ukPbFd7naQYraq6Ri6vjTMLrXjwA7zduYG3Pa92jSd1tAdvjEQHH
FUy5W7ZakoSeABoOFGZe8O+lR3rrmmXqNve0Ym+//E/GVBKS4W0nidcY7atCkrJlMRULY+4fQZGL
Y81WqXyhJyoFU1NMSyd83WIe1dj0H7qofJVvPtUdEwz7DSdDiLTWjlz1CpoW9/HakdP5eBqk9OEt
Vt7SAQDEiGUPr+MjOmWsHspgzaDPvRrasMC7KEQzmqfeXGCIDvUyh3/faL/QkdPn+9F/odmMERzl
DfnMlhLgKRK0iMFXGuIQvInsB2LZeNwT//kQIMvNnIrEXr3C5Ka56FYJrLB8Cls1Yv9F1+5AkpX4
QShrHbGdY7QrfWaHVgwPBqewQWpRlfzOH3fRZ4wMFZ+lIfyjqE/RRfBRWXRZfu+8/pPXPiGc4hKk
u/eUl29nKJ00MGheP8Q+uayEPl0RL52sxfzfTCtARMhWJHOGXULSTg0R7ciuWw91JxMTwOExpXil
oSLYAu32JeuYFSuDSxadJxv17uG58xpu53WtynSHZtNadI1EjBpBQkut8MBb0aAr+uTBnsg8rpHB
G/VlkoVd2Yd4KMrGu8tlhmVqFFbASA53L7G/+gQpaHDIe3HEllaLSxJaI3q3Pbx/5ooBS7Lz36Py
3F5gTL6WPRy023xHQTf2R6/91NpOBQGu2YBP+lEP0LYbGrgZ8LexLkgfSQDLHyQVcokS/55Dv02V
XsMOyIqssPuO3ABg+oUvDMk1AMjSg9XMcYKGtxeCbC6wi6M3qvRl2dxe8o0Yga8vwJjzsf45z3EW
l90Upsugowa7x0mfnkjR0xuU7o9Ws9zjA3dmF3doLD95R4DmfkPUvZPUOgjcm1Y0yPK4Qv82YJ/H
fSnDT9EucI6fXjzsYd72AbWRAaxYEdYUx2J5JZ78Oxs4vWLIHvxxi+TjfPjw1vGuIwe7RK1okYUb
CuuMxRnMcZnaW2bG80SFKQElYhqaDjK80yr2vJE9gE0pvdICxkQkVoe4AR2gLmnBlBpNDL7CgZ/P
ADr3yiTRVkswW4V6H8WpU2i3eUIi+tPqgunoA4k+7AmGr9/ZCrb4iHjJE5rjA+b/LH57yJjDtFok
x4G0qsNxX0uNl2pSTnPZFLxrZviJYATWSK6Tqig6Oe1QTDjU5qFsCAiRd+468JXLVqWOYG+IsVFx
hBhWuD9YDwLa1oRCnUPdk2lmVxZC39hvJRNIa29jOKLkPeCwBBenKvFn9T+bjxPxHbV3T9rdsR3U
mVJUBWoi+K2Z4Icv4huv0dr1OuKlVA0x1zuhXEPZEyTk695rz7dJ8RqsEc67vNuVRZzxz1Lj0/y9
lhoop778ktB6Wq3EZ6GhjoZwqRTHoyTtAGVHMkUj7qDw0bDAEYAAFzY55kVJ2r1M99td+13o42xH
FSfKN5bZAB6ePPznK8nNvQ3D71Z/bBBWZIYF05prkc/hCOsQBRDl/Gx6baap2hrd8z40QawCCZq6
mhuAC5a/aJpzKThPUoiHZmOMXlLR+rfXV5vhivAdnaBmxoiSI/LrGviqZR/mCYsaheAjAbe2ktJ4
VhScj8b81GzwcHFs5RwckEcgfUqwmsV+hp4Se1CDB+Mq5ywzjIpmIFyn1Iqrf5E07lv0cMvXBQ8M
CJEQqR7oUNacR5v+ew3OrxonaDNWTaoFC15MUkNf8yofu1r0p+7Vdg0AmzHk58y/OsXBVv7pGM4Q
KjMzJqo1PC6zltFpYn0GgM+IJK8XZoP1m11XM2ZABWm64xBrsBxWnGN4L7VJ+bbuT1TsoY+sPY0Q
i/oUFEVaNlomRtBFSC1AS8c344gJSnKC76vxjpLF6o4YmOGjkt0ZsCxawojCqPWPB2f1JZZIrxfv
9DrG85byZzzyOVOOfl+OI5H3wvJ/amTCgRSw6/5VzKtJCYKMrzmGqXE5D3IatHVWKlxq6428J1tE
D+qVA7bPjwjPABEXHMnHf0laGlArKW3Vkcq8/5wgc+Doa1CQMVIiMwnqnH4hM33YS6P/OHFBVL5h
ylkBculFpHuu70iRRGBOfDmppuhm0o03tPPWm6kuV9JxjkEt80+1bfbhL58Xtuzr4hsPSG/Tarvo
9IJJAM33nWIMjUZaSXeYDsAHtrv3UPvbfuwRwoi1GgnFV0ubl6qTt30uhKLB3AqW9OSAWEhq4og7
C4D+47HLL1h6pT8A8sZJZlnZD4RmTg6Bpp3p1211qucZSi8YaP3zLrEF/JzICYHVfZ9Z4mN9KHCF
P1vKkBhvWFF1WL2ZXDwkPbHxaLjexfycWqIz1TDE3WE3H0BS9Z5PhTnO/JUiHtUmw+wqDWYLZTH0
ARaQbtqThRh5ajO6rX6Z4/VWpvHAN329TTPiAH+J/wsImsZeAutdPZfYQvh0kFQPNaqBSYZbRyh8
Rnk9MaLBpoy1jze+wDZweCDKoRH+FHEilL5lx05U6hkrza1yQ0OIeb4gqH65r8pNHP3RwS2V0Xyd
ADEwaY2AD7oTI8OeimtRCsNs4lpCbTHJdyvGTMe1E4kZYWLnqE1/AOgdDydsLUPDRJ41XM+TGWLq
HXpbgStZI8qPR3HgZTpYCXxCDthG1nIcI2B1o79tWIaw/O/SP6F8WFA4HLEGjrN6p5l4xUy6KIg9
V/mwTozOnQdxYJsLlgCw1YiAy5VM2IjZqXZk5InEFiBVSBKQ3iszKJXAHx4okgOJgrR4CeAU+Lxh
Qog106u11f1z5YsD/byuwH/HU5pjVZDkzuoPpuFzKPOCiZieSfkS6T+kFaw5i3zxJtqU0vSeHrSp
BfBMH2xf4iCje4wcsxVBXPbDGkHw4iBKSXdVDa3WZOWnNYAY+SxKxjNif1C4xoYoTqiSvOPbBwZf
d6uwhiCD9YML8e8+kl2Plm0mNUFdJvEUg5q4sSghCVX6Xk051iD25ZEPfK+oo9VPj0FmXtGEfXxU
qgLShbr+9dDMWKFzFMnEA7eLSGV6ZJJxYxQ8SKThrlklklNmW4p9EcUKphfR4I3z5MYQ/GsAEcdU
R+25foClzFats1Cm5mX2e17zaLhlv1VpFsNv+BMau7+uJ8BGqlGeYSV6jFu4Rc3yOHGs5R7GFLUV
q1hiQbAbnoq/otxr8ynxU8zUmVbscaSr+SelAuiRgwudOIm79IVhAvPHR8qDShi99DdGKc0bh9KQ
XJQaeMsWfy05sxzMCIxQiTKgF5o8M5nMVnBzFUNfxxnydRWm40Ri58nZKm9bE4P0bZtmHrRLn0eZ
tLckf97GfnNeCUf0IgOq1/JsQX9WDSgkrqAhSfCQhxtc/9BxPHv98XAPVmH/30/wh7505NpnMLIv
mf5wt2+gQbQ13gFjssdLbCq8PWSHOdHOFcobKNdyrcVMcoZagL2emAej+NjVD7Pq0DBRbv8SzVeP
ZK9R/o/dnuOQi7CUrhFC33P+RR4YMF4Vhf0vTKS8ktOojPRa7o827ROUpyhvFvfPOEcEde9TJDWf
ejvaGb6RUlnMiFju/ZVo++fYkLLnHLePwqKy/rDU1MhY+zhMwVijnnx7zR+jZ+ZjVa2wBnhU4P9Q
KVITOThBQ/5v3JF5j27w3HvfBOguIE7AkcDnFA4Iiwz6qU66RiHwzMCTVAOvLSL7EPCwolNFUOFN
uSdf4aalrlAY/7k8oTTcPRZnAncyAhZdTDwZvdFtExjYduORDX8hUJWdZGzRosOSjuDN6ShiK3vO
ANSR8FkXYqcNly695xZyInI0+xSFLfdP2qt8wyQyDsPsIP6sUVN9YmurHLo74u/QlxqfERPXnGxj
VewggGt5XXZr8zFEAeK4gxfwsFJQNf6MqgKj4QbYdTDe+HEnTnuz9WzdB2HAtwq2htahEOOwkdMx
NeURQMvC0s9K9FkrZsCv9i25uLRA8mrLsQh0gj6AxpLj0LxKsnXpRaNhawHAFRq3R7puQxSjljN8
cejRINg7okvUh4ULlbttRQPAtWpFe3zHNuEimp6LqT+r3Qf3PegAFJ6uEXfNl7abo2Q5LfLW3EJR
A5qeW/q1sB+Q69kS9e96jg3VHCLufGnIXj9k0egJeKjTv/utLJ3oBrULFZxQAr1wE42pDDdS45hP
X/JwfMKdGTBWRBYw09MAs/Cz6zkFeGQxY5ejTZFkU6nS5dQydLbPBslCMPZ0tMDFNwVYRB+AJcai
sucDsfhxs1qVRe9X3gwwhCuI20xciiGuaxIQR6ZJoWAXFyKEds4MM6j/rqPGLLAXjS5r/W47LgB9
+pC6qcOZQlfH9fCCDwN1t1uAu3ohVCfyWcApj9sNhNcdR16O1J2TfqdrcYNNNv6MhmEZ/qKXK5dr
fiRMTFo5OFIH8VkUhCM6ZvHgEL4dV1NHiBOlho91fw0+xiqyjbDfr8FmiOUGAC2Mx/d7L6VvCAcG
wvl+jjBpYf94WZdajWlmA525yh5z96vsB3T1WMeB3NBQDJ7mie0GKCxev4im97/3Fg9UWEZyAU6H
m7cJauO5h3G2zRFlMFzJLq4jVvsGLXgQ4dA7TJKS4lib84H0TuimK/ZicLO6sEyCjeB4mK220+CR
6rBs0a8ji7dXlAY3nQcTLELHn0AH1lt9X88TqGz7diVO+Ifn0iQ023x5BWl/sKZP+CSsrIw3qhDh
f7FEciTSV9NLsyf5D81Vk+I/h5rKvJUAuh+x+RlUnxV5V2JufDuW6pyAjVkATAqQBX6Iv8VpXYVZ
tyJp7rIyePNRpeQdB2MkUm61ZtZvUAt+aTOEL+zWe5ZxqLWukYOfLxFBwPiP8/bLlvoaYsinWaPu
aLKwK4wniOLbBJMzmxzPO0Zfidf3Oer9VFZWORs+XGMzmFUDPxc16PFrvfAgUnF+6gBTgB24Co9x
OoVCm8ITsZdzpW1VVpU/+sRsVi3/84Nib45gwZVgog6kxuMcAPkGtAPspJ/pkmeNZEINh4YhktRt
42c6dX2uMEyvfK2jO8jvarH+E4yqHQ/rYR6bF0vzhu8ZWlE/nMar3GVWuYHcPlgxKS6jwnhH2pM4
Qf6b31dyCFY+EPX49iPT3Y96MXBYD/Ovx6gF4+FKmmH8Kh0Z+6FW2JuybyEXI/OXSt2t2oZdY5/b
k589Vt60Dc4/sfBjSPNO7UQhmLNIvXKJzmQvXckFeHQ24//EMKZI/p9supYfvmr45UoNbOlOWiOu
PpD5Tpv4530wpfOPNirhFzv7F3mMsbkY5tGE3DJn2W8uKOmFDbPRbLd7Nj/VRxNH+mGf5mYmjcIT
FoaL/OX9k1KNt4+MPkfrBUF1GWmpRzZNH6A9Jwj9/Kc3123mnytcSNNsZNBZ9qqfV3DTODqcNgnY
IxOW7zwsvxjNlHJA+hf83zHj/pzdpFEDK/LDwmVqpd8+Icu73qcsOmHEAK5K68z7VuggsqrUqGB0
Rfkak3OtKyOzoWQc3UR9kZ6CZRDXPH9R0iVPKsnMzv6S8112HUTC8je31pr48g8SkQjkK+65vx+I
8EHHOrY4ZDmmgf/cNgab0p52R2V81jMk9skA0T9NKrPhUFkQz9ciX6dA9GkrUIrGqCskGSGpwcGj
Sz+JdwdfEbSMbTBuE3nHNF1LSmjllw3/D2W97pqAzybFodZyy/W7ybCyTipCFc4dBPe3ACyXs8nR
G376v2SlnfZ2XNH4mF23+CCCd16uGO6YqcCAuhClJQewYDxx3Y9FHVheL9eyYu24Ws8QnHoEnDzu
UqvtpKV+KxxM6gVRr+izIj/A+He0htOavs1/VOFm492X1hWUKpKsuk6Vq/h2yF6Xlyzp7xMRA66j
lTKIaTrklmjCo+Ln8TqF2Dw76cqIC2EjbzFkQHiPB89HmMaqVgiskoGkGUYcMw5SQtDl9EVqV37V
f4vR8iMdlUooJ3zqdDE94SRXVD66mkH+bbqB7+8jWnXdM1YU9XSV376YXwn9w78VcBlYjOLiz6wk
sMirXzJJJssv8y36l+qF4oz0v0HO3/yCkrtd8uJRwPa0VZSoVemKUjy4bDj9zobq2UjMKfk8X4vP
XHQzq4mKzSD3PI5S9q651NMQI9rvjlPOD+RcW+6ztZg+vR8QSCHo0GRNg1rvljpUWNnkv58Exnfg
14iiJiSa8mcNXqfBrbRDTVr6/2OWZDAMcwEXrPM8SJiyv/kWrp3jQy72dS+CyAbEnXlQnS+v46TD
nZm9hnh+yue9pAr2+umeekdQe5CGC+QuN43V3EleScxrJzZ5pwfAP4hhRHhFKv9PsZUl41JlNdhf
DyRSpS6glSAPKIzaZAUixpAWvbrP6hPUZW9hIKdOMcgQ+/oS3QLRkVOmLd8NGgY7UHycPFdBAke5
VQDco35SdNZA0HMuLZMbXZ08dwER+sOdCCUMLUyCF7nGkutuqTYLcxn50pLEOIcgmbwa/MiPIXs2
eMj2ef8UlaRoz8ZjdSJep4/Xhpcrcaf6xsQ9Yvo7wi35H0wdbjx6mODzY8Ii3MLwdxu2fJgsjojt
fhGTmnQtcm1QTDWhsgNrVs6XdobOb+LGCdbPQtZBdq+pZragwpxJkHH+X7TNtgAweTMZ+DoN0cTj
HzoN1VGsBEN/K5+Pv9INTuluQm4f/BCt5+BZiZfmWiVuxyjvMaUdQ9XrMltfeM70TycLeOYENogi
q1RxX/H0IOnlpo0I0YcHYAKe7cI0c1ycEgQPkwobZY4Oww8P2xu5B6gAGzCx0NgzXHs/c6CcQdRt
CR45kERvC+brcgKq6B7IALJYjVMD1JM5oZKq8xvUz+rlegGs31Wd2UoSGz1vIegbJZXZIeB8QXB+
SKfGjwhmYPL3ewGEMhf1DZgUCU6D4n7A7eJbeYy59/ND/k++y54px9LgsuqZL5is5fR7Sn33YNNV
gjHVmcniHxJuBYp4RSmoPRPU9TEefVTphLRmqQ03qCIqCz0Zkziu3xrxCUgck7cGbcEo9SZVqd48
OhWNsmhEwV8SUOOQjMu6zbkAEJguvxaTbAhRGqDbLcMOAd8asXv0MebBuLGvJyJYz304V1jXzCOR
Uba6MWbAX+wmspO7yOcxOL+gk1CiTkEfqC1TScHc/1m2iso4hRLuGrMJvSbr0Fwcxr6M2DOa/fj5
tPVZAzFzLp9U7Zg0kKRZlt4anE6IR9G07F4veNDDwZCaHI5lbQKWinOxH/6FOFuPe5KKVohLE0HW
E0X8YKtGm44hwVbs9DogRbdJ/vEY4ddoQUqxkus1WRqLQKI0KtSZWQmFeP0kWVJ73SPJ0gljli+m
5RaOMJXxe+q/YZ+XHkEcMxQe3fHBPi1iuM9cZtKPOVsJg89BcKxYerawuKA4J6z6xgdSLaO/8CXR
9eJa29C59U5Ny87TRhYiEkCcE1AybkI/64kKI7Fc21Sa/rElLC1oWWUKKs9RmaRCyjkBAtYS6QaP
qckzmUlr8lp6GXjYR6VTTYZHmB1xaJoVjW6bX2N7lwlr76fwrUDzetji4y7dphit6qq7VRyQAZ9q
H5o7cI/OhKgxUBxCf80PxxoDoFjTSxObxDxEAz+X86CLcmsq9fB5kyMS/wgcQxFJfnu6sN/i3RpL
fxt3d6uO3JMbZewt/uhsGgcj/PMC/KOFjgkVWQ7tO25Fg5SOOoNI38uDoww45ZTHGFWUC57oxbiG
RaVPP2x47H+GI01DB4s/K99BAKSUwzibB2K8VXOfgzf8Gupt5GeAg5giHI0slR7TGJelgu2nMcdm
T87snI3WM+7+BTtTlHR1CgN5gW4oEHT7wulNLecha0vWbbOX6zzV5qDQoLY0GlKfaWFh9AGSGVd0
ZpX5DoXxIUC+LOgN8wlLcb6NguWKPdUhhwRPwcHTnKivaPc/m9PYe/hDaRh0iC1CdPWGuKsWJh6C
iX2wgOWDdlWZ+fZ70xkCjAy2QE4n0NuJXDqkvJiVA5w1JQ81xpVkW3ImiN8mKPY5NbNoyUACY4AW
BNx53TVCGP1MDh31RiX2AYcwZrXdaqLz3bgnNUsDZhGbaq8tFKmm8xceOAt5bafdlKKrAnLa+B+x
CTQSxCJ5HXAIYT5g8OOZCxUkz06Y1CinnlAsx+GZKlMpv0XXkacNU6XP5BwI9EJCIRjZYQPCAaL7
1oJDNhnG7wKvy/9qOb7bCw2KiLq1impBH4r9BMphzNqth1o1R8hmP1xVoJOambBAvMddoEKYQf+Q
y/DIOwM8fMjsqwZ62UNDLun2u+gJAmrUB2ZRcKD/XPnnQyJMfvA+5/CgJ4ijMrsDXsqk1bTVbt7D
CX98WEZJ0wahshzbj3dfKnSTRCA8lMucOrxOcocL5JjvP8z/RzALThRZ2zkOrzQtsMf5mnq/nUMz
JQ5tuOxOyKgZ7tV3CVdEvwKjPU1xLy24DEqsp61I9k16//J3Lgy2oBK9tKHRw2SsQt+O+Su/I8FF
Rlv48JHF7n+DK9MUCgoHsuSyHmAvkk9g4nbEIfvqJMdIgeujhbgbxq5d+IEZ4amGbxUFyJyibaVs
nEyd4qRIrtqY/1br7jHpdommoMDqJGQyeqQv4h09Y8NQpTR3F79qRjbX71+C5MzE5E4wvLKxurwZ
sN9YFB2ttOZ1jzD+iJMRfQh1RLYXOhEzvTUDQsnAHL8e2fXqEEFdOTOXN96AzWAllNyLQ62d6xBi
S3IxL1PaiNzfKADkA99+RpMznWwEmLoojJxElCumakEEChgr4iSjTZeajsL8fxkEdmnYp4bKHu9+
v4VN3bzUFTLhv0hjY6XyvwKBUG0pgjjx9wmjgRZjdHaW4VNpH7C0pmmJvDCnACbJnt7KrxdW6srh
B90ZGI62rnB7XMldAgAX8dzBpaGZnkAcOd8eOiTXM2S/ETJA24Zz55dsLiI3oWPKjNC5Guuyf6uj
7aeVmlQI9eEW9mWqfzDm2JQdIWVn3BvqlI7a2Y9HpV1/df+A8mmNRAjVaMsjVSyjuIDH0WTGwKoX
CacIjk3d+8Mp1wThBDPXm9HIpqBpvkrIGJecRWnUeReO1LfY435GSKB/2AfpFt2Bd04MyihjsXBJ
lZQOqcqKACVt22/Yquyk30IZIahnfLLhIxXdeWGX4AOoighyngX3hb56gqb+vld9BxRn6kbwMIUN
3aglifGHYgczacGrBoACCwjcWg0TCEFX/1atrScO4Q+nZR6OpH3pOaAx8AN/V42zQ+bAaGYnv2HE
uQx2TPNXiLlKEZmou4Z7ZTuLiK9Hqa3NdMXO85sddKuL/+Y8+ZNQLyzxQnHHgRugN0rHajCrqTNy
Rs8gfI0Hk26oOCWI+fF7yjLDxtiYbL1tx3iESTkQBnui26lpuWOpnc1gERo41WM0HemfiYzSbW6s
mJjugU3NPwYDXpITERHidCLm7xE8QxUieR6YNTk1gHeOpdgbFPKi4y0NxOk9HgrHo8fZO+kne+A4
GCcqupsf2y7PE1Puk4gOoR4cGL36BBpyly3c20c6xTtZP2KrkbB+fDiQcwjHk0USLDvG+2CiJPZs
NyelyUeKYEisG5bZt0FJoQKh3Dcbzh8WDhw7uKuiqvZBWwaSLEdm2htp9RPTw+nsNK+UeNO9XWRF
yxD3TDjjUUNVLOMWZsbVN0GxmkMOywDzZd384t8ib+HalmlkUTF0jdSoSPnkEO/Hb/MVrx1B94nG
cE86e4U49Fj84CM+8d7uhBXKcTK7gWQncijdQ/0Aas10nYThD8nLuwu67tmKGhJZ71MJKYMN8IL1
KO1JkEi42jXLYmx6n2xH5umtM/nrQW/lc/R2t+T+c5fQYCitwbl/reWVzX4PSIe6KJo90QLM8PSo
D79uc19ZUmYG6gY9VRqkTeEQSojxyxbICZZwX1gazcOBCRc2mm5JZQKlP8RP2v8v1jGLTTtySeHV
N706gRWv7eqT6yxqjWrnMj7B6JLyoAL9TtOkdzB0D0EhAresDzUDozlo62aDzbWKTc2u6KcLRLUZ
6VbFshR7KEmJ60Iabqi6vlKP2RjENjtSUZpmguMd8mnyC95KF9RcEY7GJ7m7Wk7keq1RjMzXi91j
TBDc9+eVB0w09EGaW7n5ViRzlF9QSh0eO798ytZLxiEGBUhtFOAcjOkxWvFFNKdlq6METcodGlUn
F9SpfYzoPTsAcR4RhwYp06zEX92HKozaQVP8zwel4Hs3NKJASliecYGZj27IFRTijetA50xJffej
dy51ZlhAYiD7YXUb9UBj+4xiIpVNHlqIdJsCUu7h2De+rf4ZQKc4bxDSF7Eq1YLnBEXsVElKqR65
5aFoRLJ9AZ23rKmVBaJ3uaSb3nUTJnGa58ioA3+avQzCKqKbHGIUgQuAR6Z1NeWbXdZr5Yb4c6Uq
EcVSUUaTXCpLd2phLVXtOh4IB6HK34MfKBMZGrmvlFFpADbMRiQsd5vcFS42VIbqcfn/0Rd57jFH
SmU596X46KLuFVOO1y/hhWcQD51FCBDW0OLDwOQrWGr1o/sCMzGaCpS4FXllRQiGbLgb66Hs41F8
QP8mLU4ShMnoe+nlZHrarmYUtzDrAkNzVAVtjLqlj1B0bH/0qiVsWrFZJErptccRRUJFajn9RZ0w
2xjs1wUmO5rLaJX0qcW2EeUIIrCSpXB2+AquQy/yOMR+OaiyYbvHUP4Iqya1GYtsYQtJUYY91HbI
fKI1rKREwucJU5MvF7e89O9pQJXEkDpXYjSXUunN4QnkgrzjcI9Aw+zt9u8mn38F/dxB8M3/JLz6
PFF2euHfqXIc3lgaj56m1ZaNQDVLIdhSq4rlR3KlH1OZsxz1TvL38/lReLxsZrr6Ax7vDi2NhLW9
rtKJpz7RXJ6LWVmxRmSO8gjDLHZ5WqvZqvodtpUWgaW2pEHlp26B3DXYcvoncjVeRmDKRQuDfqiW
ZYUNyIbc0dNdenMWu+Cyq/CRaoJQNdFLQejXUhfwUYCkyjIqeMnbb16lCL+zhf8ovVr9uH/J91oe
2DzHeDsRDiPJW1BBh0vg7t2HmBHL+epCwZyrQ91EsAmxVjFvh25fAXH0Z+k2XXveidIspSfAz4mn
0qdO1oO1xC6VRcyK0HdEnE5dW12brqYpkroC4e4AzFykvd6SRHqUKHY46L06D8/lQsADypx3ARWO
HTbXa/1bduFQhRtK+4HJqf80vKo9nKrE4weqFrnuvTSfwfzc/6SA4ADcGuw8hyc5e45U6+NNtodN
zECr1qD0jSKVbx3tHJU37FNEKBprGWNqOMscql0ccE5dObyB5cMOxNQfKaXlpAanmqwHfPE4G+qF
m8gRl1nFPLy7GpDE7e7WEQV7RDq4ZW6MCwqj5ebnV7g+XrwpOCYmn/IzswHyINb2yIFVOVM3bUHj
DJ3+fM6IlWh25s0aqmQc5VCcTN93Xu4yYMAFkNTWGS6U5TTbBo2Rd5AInZLhcst8c16Zg6MdSoh2
p1kfjQUsPSIsnUyI7Z0/JtBNSQILaE8NMwy2lYtfBIes/NN6HR7D7KCRIoIbzchcMaoJT12BSDD2
hLffyPwWjhH0ITBku/D2su1KDsUh2ussk3TBTJpGYac7kFx4wjQk3V8Ckz/biSgJiJmDdW16h2xJ
n7SsW8kPa6AiEGP/TGJkTfBrc0EpAbFv8PALg+m6p43Bm5TxvHDTtDIV1lym9HcY0UFY4xVOQaeZ
BPdAzd/KKAz7gpJpFRmFhGSp90fwYnWSkGmjRu5pNZs5sr8DthBNcxMePMvqVJo1reD8VApTDodz
LjELORTz2fM/WhhfC12fwA9jjGglw8nPpix4+J5q/TMqX5tamC4UJxdYOEFf9d/1wwM6JtHq5A9z
kbqfZBXekP7sQVQ6YgemIiKFfw6d+cPoX/Z0E7B2lWZPbfhCzoXxozEor8CiadCIk6IJEC0xfi3f
rvptgTUSMGyLvabmKAZpBjC+OmdQPYsc76G7UwFHUjEvA+GloicY6ZAQRRnJFY0bz+5f+XmesYiO
Rmwve8tb77y2kmzHrB2PXBbk0Epm9MfEsdB6z8poEVOe1Bli83nouLLE5PQR9TgN4sCkknmQWYcz
PXBrn3oT01wIatMuCVBjnIoYQOdVPms/jEdCdHpNPIjCDemQxLTUUVVA/oaB0akJNqF5999dF/QE
Y5DKNRUYp+C5vK7Q8mZUaa3TXB1uGt8RM5bbLh4xS0zqBV/yPjVwuaPe6BIXFsafk52LdYDMp3t8
KRve69p99Okbq6SV1w23lHf7KV/mUYnzPVkd6a1pgU5O4okEno9Ukd/3DUWWO6+2BggOpt+PFRl8
R2AF7P94NPVMR2ddbpO6XoTLxVpr1ALquMUOw4J5X5Ptj/D8Fzh8KUpZCzDCzGgPorWe4mwgEbsp
Od4ESrDVRXyjEZKj+NG5RPlB8O8XPHN/g8oTw4CHSg5mf6HcdymUah2t5cu4PfjZCRxfLEv2S1cB
Eajd3zPpYT5x8Y7b67Uf3aM4IOK+54VsiyJMG0ptewUXXlCtN/QpUYVh5iXVZcdUPTGu1eVbmVGr
lzERJrWE2os+64r159x95lHbXgri4Pii4bG5t8zKxDc+zbsE43mkPiY2vb5a6lLB8IDMP4QG9bvc
tUbwFfq7JJbFWmQs1FIstX1mD3UHiQ4gAKFkoeusv3dQaXQj/dfnc3SeqzdT6Ddd4JUVFamDti/L
Foydymz1w72hJx/7SUtmb8TUS/SOP0D+oSHh7ks9K4l4+HLzEKzlwZ05eOr09NnRUkyAYcnCzZsS
CzE1r9LmIcUtgFdaPgPdQcV1tumIEClJ0aC63fec7OYSF6nNxD7DOYiIQY3bgbnZQGlj+0F6lRId
U54fCYeiCSvkH3m6J0cnGFd9W/ZGocxrA6CWm6PyuFd3NSyLHYxUA3ECkBXsnkVvMiJjt6/PRdsB
2DecfVAypEiEi6dx8CZ3Hrg2cu3PtHZz1aSRpfeYFpfk1jkVLmigB23bgJq5nhajcoARSv/lnq2L
PF8fs9lHTumLZ6W7vveE8a+fuxYbr3ExciJCpWPqX3Udunx+6SQ6ldUOcBrFNbVmOFJ1/GAqEkcC
diTMsH5Xg1Djl7tHvgNNa9TZi0j0v5TliYv2O6PS3/mr7LVxxINjGaQCsDhh+wbIGJsLLLWt550S
sYIAWJrrPeN3kd+fTQmuDLpDdjLxsEisUiEszMosUEZkXOiljYM8bfYkDXCH5wSR+H2Nd5EnB/C+
sBi3eQryIlImSlx+ToPju8KjbcPSS6Gvy42hxzlKB1hNnbaryuTsir3EQm6AFeVXVfAiv0Arddl5
sO9F2SF8IxynudEP0M7rre8TPBPJBJVbK3adTxe5roDTtyo4kMUoa17SIncvzDXXMVh/zGlUJYbK
NSPRUigGuz/taGKQVTt3i31g1SaKeOiGFbgnorTy8WJInHL3xCOQJrYBIwBSh46shM4ABQ2EVE73
8iAvY3wAv4hKTGDho8kri9RM2FVNK1KhQwb4N7XTeVcR73Kp4+4BIB1dM5Cc32RdUXbCacy6Ncbw
i//1y2cv2/WpQGY3HXBHyZEzgULM+hmoXpScuD5ztwT/SeQn2+EqGMVRJqRb1m3i9qjCtswPfN18
XKRsuSdFnt9cLPLYAuNosvk33fx3/d9llbJgEU+iyMELJ0bXQvZFDTU3EPnr0Z+BMNUVS7CdIiI+
rYwQg52UJD1fd2uRl0x1pBMR/l1roDOk2WL+VvE8h4xM1pMcoOGcHZ1NHRRFo2dbZwuuxQw/spVO
JivM9JKR69vMyTqAHrZvanS9Z2TIHgoaZSzVb14tgdY9L8fn1aRfo+x6KSVL7nP2db7CTWVmhqfN
dUysVqpeuzcxisCNOvXDtWe3UpMrQQiDcmeSC5W/0fkuKoxTBHuELWEEznb69DF4OAACp8n8OFF0
Scao8KyWlupXTG0MFnNhz0b3TVhVNKZMe4U04WUd2zV63onjuapzrNlsm+dxoS6zHOY/XL+k9OWR
jnD2p2wDL71vJouGIPlnzU2TUepxAtP53dqPg3/rFJcm/DTlzvYlJZ3lIrrs5FVTTEDBzwp+dz+b
aiWb+AKLhSw2S7Wqdd5Xw2OL78OBrZnYIRMQF1616NZiLFigXyk+0L5oyVWkI3LO7dRsed555dM8
oqHi9sU6vobSYFYMg54WD0mn03+4Olm+g2YkiEgMDoe3fPMHWqbcbZ8ax4p3nEhgqLizFV5lfNYN
o3nawy1Yp5WJEo+D0LQyq2ErSW71wcIZCp+Anpp1/AOVY1XoYYYK3q2TYf6jQv+HHTpnjzgBg5Xa
9uJpuzg8PpDe7ZDC4N6A1P2t86oQiqsXQW0KLleGmxa5DaZN3kdRvQ1CFgnVduQXL48MJN3GqMmJ
lDo/UvnCkrztVCwjZ0l5K6vIfWPzwS6mm2+ZvdzgjH+hbxiaSquojhi+V4ZgjjrkoOesWZ5e8jNq
F694MaXvuILr4bzF2gcawGE0lp1bYchyd4CwEr+iqpQTE+WEJBlrv8wOhr/mjVpD9qJAN1TlALTi
Nmmk3/S2FiUQBCdgSvgB5TEnikmXQjdMzOn0KMuWEFl6cadqEBL52xpR26vP92QJ8tlfPuVCqiQR
fAaOPOJXd6OAZSuNq6spNkMQcI3swX8fm1jtR4DlY+MEv2zHlwrEvCbG+dXTCY+3N4zbHrK5r7lu
QhAbI1XDxwP1jdcfVujCXVbSe8l2urB0OZCCauu3hxKaGoRdmVqkH2VfTMHY/twPTJX7f+FRDY54
Dhe4aduRV6C7ZFXhPgcCZ+sh6mlamBMF8KldAyF0o+B4CXY5RcLhgaIA/Rq5SM5PmMxB2fzWMsqz
EJwXMR1rvpctKPvsA5cdhUO5xLEe0RKM7lhWHIuDeyeXjcBSrAozwEqbr6R7xjcjIKGMGToIEVTw
7HMXjAzaChQk4ZCLcaUclhRIIMcV6M6VaD9SuZf2u+POIeYhpwzP1cZdaFJ4sH2/2+q+bV72Nh5j
MTb/+JMT+ow8t84uPPxJeLiHANUzFhmf7qZWRSbqLJTAiFf5jC6i01zotVAZAc4LCqPvgEo8Qb6O
XD/egIypWT/dCNQilIpB05tE8Wx88YWLIGKJy11KVQayBcEi16Lv4mFkZYRba6WAfuMmNLx9Tstw
B4UfWxYXEPfxuknvJBUTC311rV8fzrOe0t2t9R275onHCsjF0kUkUhQISEm2YH4h4Aau9eXB1agK
2HbPkV5go52udjEBc43byab3PrElxkBLR2Z2qD0caoQwKeTmoBNUqrk42bL7Y3wmsQVfMiPHht/B
P/KUdzhVYQKl8ULjfIFz58sbLvnWQc+LQmYRuxutIAU8gOiJR8zBCtI0qf7tmC86dUJpw95lbZpf
WLgRrppr1Vm6NiQPHEDhM+sx8aA7H7R77RUxigmUFfV88GqmgNTql9JaXlgGBECezLRkXeNeTPxg
QA+kODCT0jgKjflljuISVFd8JvOvaGXj/OqOt8vUm0/rJL/r4DcHTyrzpEoYHHBJgsi5OCvG8fI1
XAJjYCFCag/31NFNSZaptfKk+6feVW5ETzVoYxUdLg93KLpzW3ju1YIk/EQpJ447a/VTQ7a2cGcB
ueq8ZSGnK6nF+188G3EFc3fq8fF2+Hvh4lIWf3WCPClUzSrW2u5eg45wbnwohOG/7+ijSnMV1tTN
wuHBsL1RWJ3h6gVrzikhdgodsl+/Ey+SQIZOI5JSzgDM7ak+M6PEHPAAs9KMFblpRNJVX7CkvOyN
rtlSQ3FJoHv7+7zsVzWH6v0b0uiG+XuksFnnPA7sX1xs+ig8NtCb1ONLYCB8655r5k46yy4P2XAO
MQTOGfv2Yk0S8L7W7+oKX3w2qcIqSCZrYLNjfO1IV72nf8Rf9oNCFAPrQiYHIa5PLKE1lhWc166l
I3Kk4ico38DR4+lW0vHL8E4i3LyueTao2U273MIolMFklrRnBgjcfiEoP/ENKd5Ei1LQTuUna7n7
03pbFbaJdO42VxahT8or0/k7bhunrhquv1GK/9MqEQsIyIm2NFlBRWiT9274n1A7nfIeyQg5iXXY
zlaQvtdV2arA+u/00jatIz724YcJc5636d/iuwd4xlyix9pdOLYNzlMSjRrvheHQcP+q3EFv2Qza
nqs3NWGrBu0JKAZ57t6uQ4tbSojd1lNRO+My+qk+CCI06uPg64r9Orx2DerlJ+XYVFug0NwzUmG0
r0KWnA+ngw/nQra91t/qeC25sMpf/qF00eIr9bUc4BRiV93wTRhLS1jgHIGB2Wo0ZuT3bZg/7WIZ
yxzjRITzW5xq/sKDOCjhtNIEClS5hIUkHRCujFPgpRutdudfDrCpJ4SyBQBTmT5LFEToNzAAwT3Z
wdGKnlc1Dz49quZBThF9gq64dR3/yXsLpcgMtsS1X8GLIAY/XuID0yRlU4dFGIk5P1d151wIWdpd
6MofvxeAAjpgQ+qdTsgQ5PYmKgiq3EKbduJKCsCLeAkhV/n3jRRScqQ8t0OmIpJMcFcQXfSap3bu
iMn1zgy5Gfh/LPZlYL0+UFZI25roMBUSTftG66rafU1AUXbekfa9mDe8xVVmWl8YB3Z9iKOnmtSZ
6LLmZ7Wi9dTHXXUiQH68LPrA6tvcYPe8mSGm6CR9j5YW5LTDWXQBnJ2S9PO318sHrkABIc36qXa5
O28Y3mAreJHYSj8hasxj99xdqKI4LPOfcIRbHtIm5hc7A2iTKBdt/ROIJNMnU1eMalwX5NI/iGJa
2ztWfGY9+dE0s3xEfsleT9WSLZTA74LFrWm2NHNaKhqvOA7gfEPM8S4Dq/x5YZJnMG3dzD30KZ4V
2Qt6Af8K8tPe/MoDZqW/qswBKiDGRzlN0of6wmUzQ9dH6yXL3Cum6KCjVIzUlqafkr4ZWyqixdWK
D9be53ytCSZxC7vboJY90fuCGYRZn2cfk+eko+f45wjoCJxuLVtqJqypTzb9LMPJHdkp6EXbhV0v
X8m8ay111AW1YwE3Thg7mTJ6EFNjtVteEKdDHUjzc/BJw7ir2c078SGOOrNlegXHdi5pDelKF34N
1JHbyXsLRQiNFZgoAypq4hniK7okpBkiHgmGmcdjE3i9d98kHAyhLC5xyrOEBN7z2Cu2tKWJThVG
yrV7FRkNZqb+qoegQKbgDsqzOgHIH3FYqczmuqvwMF8gWtWDaSTqtV115/3i7Bq4WgauGzntxHqv
mkdCcuWGi1vHo/uRh9ObKm0GTUsPMTlOLjAphyP7ckeKV3NN+GdOzFeHjx0N6lfgCdcRMNeeZtFF
x875uVUVtoKWc8rvhDeTsrc84QMqGBDjxK1khvl1y+agiNh3C+SDQFG3S2bLNPSLWG0A44e4j6Ty
IWh4IMAOOTWj4DvkXTw5RmLh7CEaNe9zQCRqEYDXqLdLnkz5mgwspNnqruBlofyLJBkDPwoM/xPz
MZm74vptmTDUMt3+ey7XJFcUIc+wuVrsEyIvHDFgSxHywfmcKhh5P3MukkhHZaKw+N6elYivA4re
anO1TOuWyFlw8a+z7xbTApBsUphykknYZDEKk/ZSHHWvL5FBv/rbp7eW0MdriuhTU2MVpZLbJsaq
2DAEbB6W4TJEVmLiwjTo40P3E46KVGEqL4g9N8liyEGe+cFXhpHn19sgZwnxyH/do0HB8FEXsFei
dVggtFgcni+G07mwtM/UXbliKKOBYHmIShIQgTBDTqV3PEY1CXXsSSn3rIvZNaJeai5Mn3YUDTsI
oF3IySx/apSJS6xZaPXqHfNfxoIfHd2amEzJfiwPX4wWvSiUVZJjU18eb+qfYKybin/zgCrPevT5
85XAk4+SHFiDjiMBXMqp3eQrMFuG4cimBPXZuG9AHwMWsPfCqx/fcHGxEniHrjw8R5BBmLkJ5Qj+
Geayos341zxhI/7ibx6NedVmNjs6DE68KTvPd1EOJXZFaNjPI+BMtBh8VzeJFCpVb8OWY3qoMpIU
A7bZHao1EZEIXi6PdlzVJCRebwS2TQKPrxAbRTzccTMsHPitzzlvCiymwO5/gLOZLpNpnM3u0TEF
bMFgQtISBYBgwLxecPRMPnEfXziq1PINjSRcsIoq6LKsddR2KuXzDqKHEc6syb7a7pwkwURy2Kjx
G+8VZRFdlAgk4Dsp0GrSHfKvBj4YqJvo/kg/Ot5paC0bwqj6yM26VAr5NauK2i/j0PYApN5d/2b6
Eccz1bgNqYAUz464XRl0REc5S7CQsF7E8uWauxrPr3JYT1aHqZzQntrXkn/jo4YFEUYvB6PhSXjI
YDCS7AxyXO+S6jZms5OlmfjUjuv93hvryrG+RZwGIPjnCrAYBTeMoaEaCKAQK5JecDilLpNW1+ii
h0/oxmyusG0Ppk20xm1JkNBhe3jYANjXJTRpOEfjhesPKucfC7HdOfgOVsVhmyeRBaUeu5j/wYfc
9F3bKedjyAvVIGsaVzqYKt1eIWQU9TzWRA3CGdJN5f4Ln+wdZbMXRkG+PBMWOjxqSQmuzELdVKXC
3UHSx2kLyrF9DYuq37hxUsM3609b2ARYqd0jfjzSNaipbJGzL8GtxheoiM6j0pyoJSpUdCYUoFUI
vobled9GINsFgNoPzniwiYKUMIAZRMwC2AmtpkCFF6SfoSauFeJ6y/WPLw37NLtMJ1NK0YtCZWBc
BYpsHakunJKyNkUFEDc63JMw2aArIGtgagkkg2OVYwSx0FTZSedCP485Ll/p2Hv1Pw5ry5uTXWII
yQI1o/jhVDLmXRVHzKfyMB5LQKgWGBXAXf4vEaJ746j5MwnPVRoovSb7bw1Aadj/iNLklMhgQQzL
1f1IS9uY45VSJWyo0Aow/pYc1/4Z+l1GbyuZeFnc5iAjV9g9bTxY9YMpiAgTASir7UoFM/R5Tl7X
PbCk7fM4gpMQR++ReVeD0n9T3sOdbV83Ab8cPtuTL7jrJGQqk5zFTTWwNGLTAduump73im7KX9zF
6B16H8lTwEUAC/imlDJ1aupVQ+LdpwLvJoRbWgou5lmj6k3u4XQ4P9ieI/BmI+SgSwh4axlxtpqf
fn68BhzNe1+TG9B4wlVtIykPkO58qs1tp/XQHkahp31WH+ms0B1ODJrg5uhGiRYAnnhp5Dm7ftF6
4qfXsq/o8dW4gaNXdh13djDH/JFJR4+JMdAIP55IjLcA9WYnHF6N/r9UIiDlqekYLuiysc2+8xea
VFrfuLof8wMJq7u29SuzAgamdUHVbXiug79Da5qxhiOU916RBpmZF5CNdMAzEk5p1ZYTBNx0Ndbb
FNjtSHms4o/d3ytaGy1CEzvOd1x0eSdDK2YUZXXE2VqNmhdqhptVLeafB6KzzkjVtpvl6Fe+N3f+
AuLiO8nDTd8CYjzBWKVwhbfgM+7GeO7BoLobNuEcybSEfHypsjA5L+9EBa/nzxr3sMiYkrramUQf
s5zJD/rV45KSgqVsE4hn1DPCnJNHL1jd4d6u3KyrOcd5yFWGfp0Qx3fTSPGdyuP6U6jHm9nrdyY3
diox20q3f8Ow/jd487uPF+B5rTqwym8vyyZPvnen8V/HFuZyIfoucKs4yFRunLVacgY/Q3Bm51+L
5xm62jJYr8poqG48U70bCWb3JgCuJAIGMarYBYdPkYUgYRYSZwDvj73GCHfM66qilDiNTFMTELgo
3Ha0WBBaAdzrN4Q5JO61ejwCNrb/HQjVEdKIFgWz8NP6JNLF2a6yVLjCpFF1s/kERrWTLd4z4PAq
VPHZy8Eafh/t5h2H2qvLnzvKSCZgfurItrDifAtd7797NUUJAFqQfcNiySCHavo2wlCDrYrHC3Yt
JnCdVRyo3iOA1NuG+V5fbt/QtWaa6EVL6hvLaKIC/zuHmum+sv2+EB+jQSF2G5+N2QhZ0eQ/w8hX
ACUygYCzMEpNbnwl4aTO7dAstlsuNtP62nrku/joGy9BUaJJMCGvDAfGI5dN7uzoZetSOj+u5sZv
3bHHNyAlyKylXJFOGZKNI4m7gThEg3UD1+49dxmdR4AqW7vMRFqWcbHDLdisGdsumkkVNdgILU/d
+Ki4MwP/eDweOLMx9urM3+CAVHThfsLf0v4mLAXS4orjHKbwGnchgjwYxF/xexE7vXI3aG0gpjdJ
ePHHCoB2LWlSzJiR/5+rHhlltp9ogb615ItlFnYp540GYrlqh5/2ATlTpneSE8lwmoBnQ+PFqbPk
a5688ijWktaet4RMmwkCwgl+naFG2xFWMDy1pjKq6Dy9mTws/brU4TH0egzJlx8FMDvfxZpCBWad
IXCZp7hzVvHu7/RRGUCAdZREQQTr1hjsbhDCPAeoI23FGOFmEQCWY+REWd4G9tbiTRahU8ElmdyF
C/6qNTmRaYaGIxaOGAFFb4J9LbWcBCbJgpVdZK8cirCnuBMbmxZCWHToqIADPXie/c25tQ0h89RA
zEYakY6cZcGPsXkts1rSazPEtWDYWhIgVLbru5OVyHUyzX9GvDEsp+O+eIZipTqbd36ev7WYDOBB
IJkCwciJYQlO1LaypB4zXZSlIN423MY34FXf/OKswlS5j/4RFwx2MpsIqeHUVUrJqtOiRQ2Hy6Wu
gBulDUXeoxCp1Dlxq5vFrr3ZUnqrKM40uznNKLS+ia656i61G6pHPn5gDnZeaoj9SE5wDVl/mQjH
GSm5WGXsoRYNPiYp5fn/GtoFXOdr6DtHLZJSriv23VETtITvaTHSKn7XQtqVaFaUSQKp6AXDsMl0
WMCFHiq4DCJdOrXaEpfvVgONR6FelbVWSDBkcz2W7CcsGoeaMIA0sFoRQLaQat/9HOou3sYeem6Z
sCQ2XMDCBlOnQ5yX1SUxiy3F/3Tfz5UrNlBB5Fy44vNzWc+Znf41C7B+rHKif1t6dEsp7vn/webo
TiZRZnmjNGzvgr62VWnHPuqttG3KjOtlSnYcedHFmeFZgHuAGr2XYLkLfwaqBvKjW2yx0OPvLywh
VTwN1PVgNKRNROT9u+vGD9mUlP+miiu+KpU5V7YR18RQV6bZWOyJEzttiKcMlVeopJwmT33SEKaD
7nXNu/Hk+347+sacbyDAve97L0pMnkR+yaA37yFVDI2ST5Xh/bCR32P5WqZVCUe3DWbRo8n/R/wz
F4Uy64pNkfntpdA9TcYVQPqBQc/3k5SPwdQY8BQilj7WWNq04heDXFfKr84iEbE5ZGT9/HYY8qPn
lkMzovlGarNimDMTSiSbR5RQo1Wa4Eh6SecGkilxq6mlLNIHgtZ632+FBqNYNbjxlxHtM8M3dYAt
VffL/ffJ6U0b+yfb7kcWugheuFjg55W/iqBFL+ngaD36BUhd6swPq93vUaB6AAqZ0S1x21HN20YX
2yaboEwH52mYOPivIJwpsW3l107OSXUjZkUmD1F9Cm9vO9iqx+mNBjVLpAQSLG6cmbB2uCLYN6cj
KZgufuXxRSjGlrcsJ5ZezmnSjEi3JxG9QcIMRCzRy0linK+uE+nHExH80EvczAAwqCWGgXgtxO/O
ct7vFXiohIQbzg9rkEB0+d4E8km8apdwbOKTnYo6rmG4PfifepvSQofVpNyIsgM7xJZt/m3CU4Fs
Y8uGyrIL7Pjxr4OwMf8EuTchj2ZVc+DTtTnbYcAOvx+Fg2uKqZC1MG/5zbahCz+9oM5gwm81PwiB
p3qQO3/9wUeuzozuk/zHYaPNhIQNwxgN0VOiFwnOR+Bg2ZElSe4TgNMiVxCzWn2r6QyuMBVx+Sdp
xtOPzAZr6LM/fz2Q27d8QVaaBwKPU0pLH7HxYynH89Iq3sU5A1XxQSXT+6zEG9N5r19o/koSTNzp
lvSCqe/sd10fe1a+SXiL5igfpb99vGdyWu39c3Cp1Xl2naIHeYiOZL6yam1sfiL1YOKEJ4tymZu0
yqTxpps/2NYSC4NpXy/XhNGM3HXJeQDy+dl+bP0oaDKtt2IVajkHcOaVkcbs0VTXoOFaNj85ZZOk
MjVuVsG4ij+YfN8dYh2wirVX0eFRea1ixDuHGvHL3jiV8SLKanngFM87p94I9KzoJ86NxYUiyzA6
uVL3e0TjsuhXjt5uCJJB9YGdIk7JkAAqkpNIt1Xz+Yjda/6oGI+Cg8IH+zwFoqk5/FPtH0PwpO26
ZlBAlOykneKf4CQszIONQk+WVIwOJDR5BJRUmWoxF91cswZGBBfRNbgRwd5k08vrUFG6vfGfSgZT
J9hV0ZN3fzoFp3Ar/TDGVg3pfeU+kffDDWk9gRPlKENuGJeD4PSsEsQhnPv/WO/wnrkAIztVOjZi
PpPBPN7bkAQnh9CZ3etZC3l6/X8VShysibDUNi6FL+G+ObTa2KVV/c44CBQ0HrCYTTCV9gdOA5aB
FNugEUakWtXm0FIEjZPnWx1VjhTNJoTKrNziXK4YyCMuLd8fGmsJaFtpOWC2wBzDu/tHtdev9DHe
0jL8xO4ITkw2S4fl+hnmq97ACynXNCY+JQtoWw8x05KD3+3Km30ooqYpTcSg0Vy4TyPOVZHV6ZhR
DfWQEBfyZ/5uaQtR8cwer6U86LnERVBda56bb6lEeNh6Qg/PXL1huVMCwWKDMym2y9vpC+Aba7Nw
TSLQZxe0uycilrjX2vA2p3HcxQYDbcRh2aDQoySoaHqS4W4WFCPZcpZCQNkUCeRwsQWBveMKLnC/
MwJg/93/mtk45N/iUOuMi9xPBIJpRFLgfmg4tv5lgnJ3Mjv/PiRuDHc85YbrjtTRFgsSXfwXT2Wz
OVDhmED34QW1r3yLNkR/xekWkD8ADQz4LzwvYPOyt+cdptNE7a/N8LKd4d9R18UGJlX2PUOxiFKY
fi8Ih68sL+WEAhfNVkc9tOJJZzgnNcGUhI/QHEOmXPT4uPPX/ukS576bPpWScVohurJ/UhA73OoN
40tTelFdejZ1ztCwgeO9uoTfnej+D3vttCwB+0v9bm43W16ixlSnc6bPUtudGVuWGJJuC7e+kr+j
57rZm1FbSyfcHWzPaeGU2gY/TIVczN89GGIPB13NcoRlaX7cNB6djZaAYWFqJgpKXTurvU1+nOrh
z8Zii/R1aDT9Ogv5cuWDqRdV18n5otQRLT3ArrPnEI95X17g5AbE1cTaV3pKxfiu5JxvvtYwvLcn
LgIyku76Hw8+7K4zLgkzrhtqSYKWXa+5jvYBgg7bB5aluSJZLSrIn40ag/24l3VPzP6Y880Q7FVE
ZbVcZWt3LEezzRLaX+Kp80oEtmPVpzSmGYNBjPAOpI266/QumAf0B0vEqaTJtmWV7xo0kNXQMcYq
GNMoC7J8/cRFHP/T3csdXqAIHeNUP0vJ0eBZRrorrGFXkxtPBAxweSehTGTVywVXKh1srMs0XZZ2
U2QRL7HEziul07B1tjIRyfHuynLz1e09MK9Htux59De4MW/SeSfdlwSBTrzs4WKXQ91MpLS613ut
73Z3cNUkOmESYY9o1NSeMwDvRCD1jZwRX3hweQ279DL/Pl4dy7Rct5OI9XHOvF52mjOWRf9kVa+n
Gjm1BHRT5QYka9siQVL2BNn1D+eaGqSTfJ2kYDMqWY5MCBZqiRTcxTO/zWHpQjCGjUCbD+REeexY
6vHI2WlN4Oc1f6IZBVmm4yZAX4U8DOtYtP71ac/AHgqv3TvmVXRQTHf8bYXzfftiK2oiTz3na2P0
jbLE0BCcDnoSVYdXKKAtyQRoD5WnXQb2r+kcGAXIDh2ESGiOSAYoLuT04X3MUIJnJleyVO/MsQVS
ewOX2y4B4ZMS9E3rNfzUDqJayv20zIqEgGAY65XppgXkUOTfAzAfTw47kZC6Av3tG5JBnLMZpCEp
fcW4xexpwJWwDaQr4Nls9TsJ+7dsloR707yBVRsV/a0d7DFmjgF1OARvE8FlBWl+XkiCgcPwwz3C
NA3y7qmJF79B6Lrrw1KxkAwSb9NNOzuITnu4KpEaWqF2b5KTQibxAYQkWV89llYe3Yk97lQCfigv
9/WItER4yYRqM39VkhnywHEmfhktC7+pimThOwQXoE+nQuw8z12fN3vUYmFFjUwEXQs2yihjzM9T
EzSabdAopOqzaIVCUE61MEWlCMZ9M3MWNFFNv3dwQU57WBpQXZBGgKIjX3tNaEzqbWD4YacSkZEy
mYJz64ApFB3ZrREh2JPQvzKP/4h3LGqREowWx/c2vmBIURYe5vAD53egn5XMaQSUl/3+LzMByrdW
qvKvzboOfWM/DjeIQCIZb/H/HduKi929O3gTzcUI5S7wnUHSzqmgJReMWCcIfPibWfcFkB1mt7iP
N1X2Hh8MpIvEmQNPZJHAuNYJ3VtskYFo5TkpK2qsUPlC1nVe4W4Lvr9MZce+aK4nSFAFbLLnBbKk
T3T+qTrDG2aeYXc88rySMMvNwK1CnKmBYexhVWFSSOp+ES1x7+FoZNT195ps6j9Ehw4yExkBIIkO
62SkEInZODXmZDCMfkhDSesG5D2/tv5cN/7zfWgLOK5NU4/lxK5lZ/0MO06JCzAe+HBNuELL5cWN
Y1kxzENu83N+qDe5hcAB02xKjITSGSrXhP0wdypzs/47EmpwnjoApza+/BdcoF++bn1aw+ynWoe2
uR7CymRCyRxyT+hkpwwkkTRccfsGgAsrRVLO0exvReOetVMZfZMbV1p+Qa9oSkca+eBUKGQRC3cM
ODwEQcgnahegEwQGJ+bbwDnEYcinU13etknfrIQ/6GM0v4sbDxbmD0txHv0bRF6BdB15YXgZbH82
MDSfPvZaqnne3y87iL5LWXeuY2jWiUdCDeDk3nOO0p1zCabzGWRVEtsv6XtlXMOQX3brEQNQdc9x
VcP7f/QeWBtLOCqQTpH8WSnRymYOwex611N5q/lvvmFn+ha1wYYvUqr2kqeembEXofhpxmnW2MlZ
dAoJ6rf/2ZHCdb27bHFOR7qBqr9526VJsoH6M0B+KjMt35RhIcIUtkY4AtTx736rwC7LvLrOyBFY
waqokiFDyFN3jRKzKPSKKGBJo4RwIyQKaqN8p8y82cgvoawOzOb8LxL/CfhYgq8KfNFrY714YbNt
Sn08sEhrWNTJhW3B7WJoyU9nDgVNq3TKEu96m7zA+aNlMR3zj9YvpMJXpxgrq3Tdq9zlzbeAJQ9Z
3auHztFTMCuhM/hpsHIE4OjAC8NZ5fOPELryWEppbOQQbuqNhC4QL6tplUFqdRtN8zLkYJI73BaI
pU6ORbeorSDss11uAQdPSNsdS6KY86sFC5kiHjh27O0wFYbleWilLUH5o2mOcmOiGP7vFbK4Vygk
xQy5jb5hregpo7VjV979nBdau7JQoMgt8iUVncc4licD6eM84dDhkUQvvQ6r1TWHV5uA0zhj6w5M
5n9Zvp4mQvCJjOHyMc4ygztrxu4lzGcrPFR6c13k+5oqKi9hLT7/14oTQyCRqLVOM1vgOfraThH+
8I8+jWvhKyQozJyv+VGr4pMVOt3ff7il7xry8QTygPC6XGsT4Yo4cXwTlViKvlx5W1SskUrh67jS
Trd27duleeeL7jOP4v5GJBKqgD4h8u/0F38/n0xzSZKqTvRC60duQY3ETu9aNHhrbKlWwyY+Qpn4
iH37397QACjN3XjacmtIay/Um7PHH7p0W0lDhx+cSzxBLP9Yd/cYNcI6jCZz7qUIbCORqQodz4fA
RZjafHayLkkIUVK9/o+DLy/OZzhLtGlxeesh8AOdOEyiisWf8uEuBD/sUGTrrN32njp75J88sI0X
VJCwLmuiYYevPG8inRWrpCpyYJmwBeEh0+tEFsl7XiEUVpiTuWw+WwEPgwjWWzRMVNZ56Ivl3Y8Y
dQHw3SJPk+vMwI8Z1ws55u6dsmoXEqKgsKUUWDg58rlhnX/VJI6QtrJMKAhXCLZei04pnPMBBbX6
ofobYHOI6wDf3wmi5eIdX782906B8k6FKFfvmI6k946U3p2EuzY5kX7EheiNl6tY2REsdEpMuXjp
9UPYX1xrlrFh7lNht9gKjYtM3ld7bR5RPk1RqGPf//XUHhXGCGL5vRNoIIlopMDBr+r/iL0E+8E3
mN+nWIZiIwVg3vaRMCzgzhoIysgcw0dqb3D4KLpbHCEIMkSRM0wPOrlAFwGPrzkI3XO9sR10iYJ5
FODxkbvcj/BgGH9ftrubVAnX4+E/xlVobkD+DcxPHFRQwNDLObRXKscbp5HQ7fEXOWylTEUkMqwd
5Unx/YhtPrXSwKzp+Yd0vu9OkNT5j/TVVA2wWMrQwRu9dTSnLWww/YGboVr/hXK7E4hOtNPpuY0R
6+qBVyo/NMkY12F8cMMjzFh4iswn/Ob8jWHkpZig2yZMFoSHjGlnreX5tXe2YR/efst7Qkqt+xQ3
zw/D9a69nTF9uKgRwavrzcJRBNBRJygJjycqjC/vgQvntWCn+vIydEqmPoKXaXzD5OZhJMhsZwBA
EbdgOljVURJgV88+efVWNF4WAXAO5SfBiTfarFKARzOcE21/Mk7DAry1f3Feng3Uj/opAyPr3N0N
Y2gs7vzHekS2ostYZdV45aK1wjw3TAZFqovaewAaYVnkQQXwk892uReil96qwmhQ81SJCBgPJiPh
2i4sDSG9O53sAlETdaiJm2nmHkDNmL5F+WVKRshAsDI6B3FXvXlBndyplihonHqaQVTR+uyqWnbH
gg/6ZV8AamheXBz0TWgM9tawyJpKo6RCuBAtxH0rtUtmy/7K8hbbqSWgqHUKwNhJedwxINJVXcGt
pj3DjRXa0NJOnQJ8R/NrbIbePoaNA+VsphtQ9je9+QS40/bO/ISwfAz+hgYK266+mPO1v7WYc449
+TD9ti/Zoias3SUwnm6FZoSwgMfsgebMXHyeM81niYDJzo8VFD6KSEvqlNW0bSpmjG6R+ogGPN6O
zWU+2a1b+FfnwVznH5UpQZtrFmqvT4Ltw6RZGCwH5ePmNAgSt1yNrRV4lrA4TuY/blIwgD9KEn5M
835F4d0ScY2MUXx5iGxTH6LkIDv7ISyrf+8fuZSnuYsomHKhLcKdFcR66W66FDxCkbQx8my9pqh9
DnXPlgP7v+osfg2izzz98QECI1jnACm/0Od5IAxP/gKNk+83BXkN2oxd3LoUfhGmDfwrgWbz+8jH
J51+id1ImJd1qoYb0/eHW2yZBnSesEfV/AZ5TlxKksHjLccxZVm5gFHTCADti+fUWzmBUv0NqRxL
IsaS3JIDTXs4rwhXRQ8BXYHPjfvt0rsc/DyRYQuXTDtgd/7OvNSttxGgkmkWA+1ja+nlZKZB2ytt
YbtwhJMxZcq/8pZWa2mdf/moKnw0gfjcNK3MiifB3R64dDrBnd22JKTVMvh/l6pB4sbxxYeZVqLh
Qi4f5yrzyIn4P4YqDNkWkGWRQSQWO3fRW/CpDCDB02xa+tcaTUoT7PicVMBekzYWefMe9LGY7q2Y
fUlYjrFwFygViTXATolX5lHYL3kW5XdXyZyGXN+c0MrgI2j4dMhXav3iIvK7t3mHv99SKUd6Bs69
vspljsiUG2aee/EOCGp19tW96CcwqUmrdr4VstA+26v+Kn/9axPIsraLCiZpksS1DkHdD/Y5TK5n
QgQ17dgyLy8G72GDAXnrfGBp07gHhZxxGNR4iCsyyQ8t3CuocHDpE8ZsQ/5HREKUyMSbfiLCURsp
fribnAInHl6nj602qPthW1IN+fogWdIBxsz9pEV6e7tsHaX5fQuu9fKT5JXhv+HQbEHitl4cXyK4
HELXxVnisSP4F+O4RHL8/XHuOBayQPyYPfHl5qMYysj5Fo201NyyTG7HQMl+dtmFj8aHEZX5xBqM
Xf4NrgdhkgCvMyXHsNn6lOmKqY8iOah2slnIXS6Uaztr13R2MBtISd5glpOeQfQnYmCt22jUsHqH
AYiVNB2TYWHmphSSpfHffEB6YjPmsosmcAilzI5LdBAJedNq3mlz1JBaqxzPqKiLDV0NZf5e+a4t
6KLu/lAjhJzQVhazlCjX3Pmobm5Go4FU4R853dzxO6fvjsbMF/XPkHQYM/SkmAOcGPGI+ObbJ4Rg
jnzFMZYaHjttFtVi4smeAAoYnq2T7G9edskA8foSF+ApvJOKbThoU7GAfxnIV29erEmdpMbhAYcY
MF7eRjR6P+TMtyCG/DLhh3DQtdg2hu9CG8bcrL/iN5BkUJjdT/7eUvBkEByDpDDSP1P7jg5l9poE
vPppcDWDFh/IfefXXRudBdYxDrOXj8vk3kTZn9DgRHNQn3iW2a7uYtl47PYKCGvLiZy++r2mYssf
JawRUiaU1qoQAtXMuWK3SktOiCureqa/jGs38qYC76HVMnqOFYryhOYV6MP4u0rcbhuZZDxKKNzZ
S8fxzwuT4se9JIvn1y48EffZzSmMSfYAR0iHwhaMTV88bT8qyYW9dnFggtyR1wF/McOFyq3KQAgZ
JxR0ZASbo/fFFLV5DVzSF0g06mF+dCaZbDClGMIuk6Pq/fG8jpdJEj84Jd7PyZiWU4jG4sKEP4oo
F6/2HG9ggszztMNGagkrZytBQn1X2IBqcRmphu6birE795zuBj3r30C5SHuP/bRsO7EQ8+HR6Sgd
avJBp+XW/IY55BoUocJK+RzYl97p7s03PS5A9dwYToNUylYO/z4F/wuzNOpmliSAnt2Xr4aU6iGl
twarqBgDaot+Y85EeccEWynW+vOIxwOBHxIEMQfY45Ko+dxC7DtXa2ygFz2iXIKX0HQnE29FadbD
wVOYPCPhdmhtjz6fyskejL8QxZA8Gl/Cv6RJ0c5ZlzhwlA9WLGje5qrSVhouuD+Se1mTcKkD/HRK
2U+fh5b1g8V08QpuSNQVzWBw5jxB0JPcHLN7C8/ZBF+WTRgwQtsxlXviW7SBAehYNQ03D90dLrVq
8YcxtDxPPboeW4kiym43LyCtTsGto2L7kEe5xrerAweheFb5qt5bJ5BI7mx0Vh90TuJsbnwPSjF9
koTmfXyLGNQV8n/E9x//vseocGFKae4My+572/ck9M/UbboPkwlb/AijUhv9Eev0oVwziEjARClU
9IFEVcQd5Pa9jZgf7KI+HjJ5YYoK+5q5wtP22kHEuzV6seaakDZuvQOwnQ68+lwEO/yWaWHV2N8F
arwNFqCxYZdIDF6SQtlhoNwO4xMyLXDgiUv9a9SciF/iYUSpyY5C3fHHWSiGj614VRYM9uwKx4Mw
KBx5Qdpwokx03oOhtFYPiJAmnL7aHrcr82PIdMOd1kjc3XnWdlQ6I+7TR+l2xa7sPzZTVZC2Mo6H
zshiLRiJKv7Fa/IhiUKkgV9nYcPWxd/SXAjJPSa5rFJTY4Q9++HE1CjGY8Kvpfkv6xxtSfTKLgi9
BMLuoEdn9mrelH9akT4cfF6zXB+iR5n/cbIIJ/5ADyMO3xbnlMRXAqnM8PrAp8A+gXv1k9/sGaX5
/LTShbjXZGCrhQeFEQSf3lx+UteJgWd92kFF+f+VmB7M0259/LQxD1VxgD5KyagyLrw1TLloYbme
4x/3s/9IMCRtdLBEzBqQuGwJEkAtyotb+NVeIcitYnc3kxqCQL3q0Ml7BgoHen2w8yHH6gvm8vq/
k2UaLKZkZ9E+hVHKsDK5jv8xwK7IT17DAhnlbrVn5W6cmy5YRhY5es/dCzBYps5RYzQ3TL4q4VNi
1PoiJFgpCLia1ABhq5wNZksvlAaJYk0Bhc7RSRhIIlNosVG6OPXg+PcAB3J2GOtW9qLUiJUvChfg
Bxkc4dopTGCNVuZx/YxQLEX71hN/XfN463wp7q+v7rhWfWzMXhw1EsmZscJGMHShWBOCR55rhpmH
cT58NmptbXasqWvB5PsCgHxwO1zSGJICSruxCKZWIhvCgKnZgtCqdwkeYvv9G7YmYMJV86NebYbu
8YoQ/1GtTrbWaXLR80FHN3fpjSRK1M6pzwVOftL9i3fhaSl5wxodTQ38Exw8HqZga/JpumXRG9N3
IclyEXMtOebVB6ob3mcLrhsaTtZpxgsp4vnnG9QWoREgWp0Xv5ljZQnYY1+7C4QBrrQ9XhyH8toV
xYg6FeXZK27ou2Tfu6JqHcN27QK0jB0mUO9Nsmaut7GQ3kd5XlB0DnuxUDMt5YVVCbPaVkN5oR0o
yiiuFcfd268o8YQbYCFbme3ljq1VekJBsFJdXBrQu0ODblX73/Or49hdnkVh/ZPtNJCkmrd5s/JH
EKQkzaKB7dVzslw/nw3Yr/FCeqfCVpuC7K9gqnsGLypO9G86sEFG6K0j435qRniSAe11stjSJAnE
oZ/EUoWcHlN653G91VVC2/jLWHdy8OCURgJq4FoX3bZn/C6gDjzPZ9ZZwOho2MoPRBqyb79F90K9
MujjncOyYS5IWhh1867hkxwcxBAC6zUnzU71eQJNdxYMh9VjsJxnB1rr4x9osbYynEp9ecYDeAa7
oY5CbBjaxza1B+GWLXS2B0kjqtEKcA4EOgpOBTijH5Xo8grwDGKOW5570v3JfUNpcKhSIA2jJEB2
Kw/EoprFkexWNVMMIrtlVWOjn0hsyvSqOnAIqnnMQa1A/XzTI0Tug0aNzZYDsZZR4DpVZ6BBGYSi
vKevc94Bc2OgqUKmqRWgYuMUh+Me+VHtTzbDhHfHjt19hThFaW9sxZvqICcV78T9u4v8h+0Mm7uG
heLK4bgh4/7mpaIqa0Bzsep1LzIcFFqa2umtLDl3oE6J++XX7U+sOwouevP6BwsecLZLMvC6jidV
ZFkcg7RkSSWW1nDVXJhEJpiICFEEONi2G3XWffPApoE4V2NA3ou1ziSKaQT/um2l1Tu7GIRny45V
AjZS8snzxdgcY99M59wnLPs7SLWLMuZQt3JoaQp/27gr9Wke8WGbHybwR3KQRS2wYQNUR9lOBpGv
9MwWiXBtaWEPPTXMrXND0qMBWujDaIdabe4yQk4YrVLvPI2iHEF5IhrO+J1Ws9gFIHv2aGf6vP1k
1E87Spkhm0D+nSox0hRzUELl37piXhzc9ZgOwTR9TE/mYIuXaEWL3Zz4I+7pqA1VwUgp3MINyiJL
8ZROQp0fvnUUGKe0QAWtAm20hTaUhaHDX3YLczrlJQjCkNUF4n9a1q8TfsbF0jquABtE0v+WWYqK
QmpfrMUsNDBUvszNPD/4buyi5pj3hCo/CIl/dyLflO5KPbSdp9riwjLc67vVZWJKcQYstiKvxTfA
kYPMbNUHRLBEwTUuzxKkkf21SH5x9NYZxkJmGU9aB2LpJEZXlS3AIimASJpwUgDuZOlPGjG0fCCj
y+mWZhXywseCqudF1JrF4HE01cTK1P8wTp+DCQbz1V3UWwop5tMqfskfaOI9l4wklUAPX11hzr4E
XhXUTNKnYSnLFiIAPmW8zSpiN8CLIe/TWXLCCG+EIQc52CpdJq4DUWTP5AClGrCuKeTYiGcN1Zvv
lA3etFqEETNkEAOOPm8S/dLNPgzd9yz5NBuiUpSjJtgoQoW242iWgIMOm9TNckNHZztk6pkjTSkA
hniHnIbin9YRUY+o3UV47Tjlusfg4M6X0At3e07UEHzNXDhhN1gbpJamugMXB7nBEqtMv/UvFbbo
S6+qilKHg7GveZm1fqLpXzDUjMo/LjgROQ6BDI7CQqPJJ4fDMZWyKAxki9hX0BXWPLLaWgwYpLr6
Ohs+9q0AsEv3XL7pVQjKTQxNI7pxigmMhHOvv6Kh5gYuJxRqObIGyUtgEzjzSm5G4no28wWUn0Sj
cZ08u73wrjtCdAbu0AUYbx3OjdubowYz8qh0A+3J4Q4up8R2k85449lG/wPMdf5NoI2ePceaialE
ZtGS4pblws46tEXeHfq6ZuLxl1lDqhCnYds1/xcWsnTtUkYspQFzglJdVdh8+CPBir56CSjl0UM4
hB9c4/fhvxzzh0i1QU0R4jWnW00ruK809fKnhaEej/SW4sXtCNW+A7Z/oAtQEbgxu0+da732TdL4
TktPMDUOtWeXNGhVUU7pjRef2UyFvZZdA8wRwKRvPMUtAQiutdhHW1mqAWeMVA4FP5fDjn9zrEEh
9yotY0iBP8dh4QpzgXcRZ0h9JfXAksURUFNyUqINyP99MssislV5XZnzP2FqcUw7e3bufhlhsW8k
2+Ba+HGWCSwFvjp3gf8tzoaT/AgcGr7yggrDvm4P+QNeGq9pVDe9mkNw5w4vksf/Tejr6w30y6Po
fHKR3dJQPj+duxHxJx9UdhZzobMl8Mm6Ct/m7C49an6YSVXdoD/kQ+mSNBg26epGhNO4KmUSDCow
Oz7BO4SqVTh72XolMcflJFq65FkCXDlwfPZDpDeX+TD73lApt+uTLe5Vt2T4DD13kTHwyD6/9g0s
AxTtIT6tC4gyBjcHPFOl0hnZbX7XYiPQaTndMDQr75Rx+UXUiePs1kgIy1vZ+WdMDQ0m4R3+sfxG
EdQysKUMS0K2X+lPyQAJYTyJs9h2gvZE+9/GrO4GarTyUKgXkJjZAVcfLNcv0LhhEPflvM203qGE
52T8LXXL+gW37wJnYZJjWYYhS/cBjGaX+4W0MMxyLL5vx1f5q2N5P3rZ75kMkT16zkMatJ1orVt3
xsu0W9LWI18WD5RDenHbIo5a+btNxz+PclT7H0vnVpu5X89AqQ6obOWJWT2L6LjWmmBZ5WM2Cb5b
g0ULMIG6QKk3DrTIuyFVfsGqPSORQQOkOpfd9wdRI7sypnHjWUqnYYFgSify7SUDx9wJFA1q+jUf
UsBlZbOfGIJd+LASY6kjh8SIyEsxamtZqZ0CRdTWtP8Frt5o4OnuWp/jasFq0s6hJhGOoSeStTz+
VVxCuXARv8zykTjhu1Q6mS3sse3zAC9X8JIX5O2b/h0CIf13fd9kdaMgf7NFFMV/m4pKNesKJ6Lz
l3bgvyYh3/e/Jcg5gL5RNAp2Nc0mo5fsg54BK1iKP01mL0yd9yuQQhqKThXxLk8so1cOyfmaRWEB
mg/ckXE07YEVkN/AcY33/xjkxPhWapbcNrBJqdz1MVvdkGQMLoOL8lAcVO4blc/Jyv0I8IbdwhoI
Vw5yI8bXAS5AJNEh1hDpu2qsne170nJ+OmpnuX14HX0/Gb+FeAdCYSPgiJsJEtzLmwtmDVK0wQMM
zW73YHCFbBB7FzvSnCqrudS3ygBxmqjhQXnHd7WBMVxNdFxzdYMgoY78J672g3Hyt7l21kxwZd8S
Z4K9mPHrxlh8jw6G1Be7t3qbWYx/Iyrr0uW7VbtJDjpHEcLmdvSmXDMDaJwK1ZLBXgQP9IAlNy8r
jc3Jyw+uGgZZMybEzEHXkPhOwNAHUhzStSfmMPTAArWZZ1pYVWonqA4delacu5UI5LHfqrjow/DS
cwwX7zRUqP7RqxR8o8v3b7tIVQV21FuQD3GF3anTdPbmRpKNx3dMO7PzxfsQga7O7Ko+LA3wZzWs
WEEgT0R2j7VMejal1WKbL0qRSD7eBiLnRHjPDQN7a0VuC3DsvlkEsH/3sKWxYiO0Te434TXxasg/
rRP9VFGPb6lT8fhi0NkMOpFUaAx3JQxdrWN9SeOs3t4jhGpj0AXzqs3WRB/2EKx7BCYGECwyzVcA
zB0zgrdVJYa10rXRdQo9nKXFO4QiHbTgJ3O7DqOTK7/L4GpURaXs3Um+KH9FMk7uqRrZFoFvici5
F7q81YCtFBv2ftkdCuQ0BqtP910dibz+AxQYWpI8kSSb+GIHRpyJYOrG6GzMdrr7ErNYHUhnaw+h
h7CPjDftyKQCTu3j09HhcYavY0cJwnJJ2aFNjuWiU+GL6BWCce1/eekEPJ0ckURPLVTygaVqjxK4
y5rvPsWC+hC5xjsq4Ms+sQaKvBRwnKTorNhT9COKI92+Zy/oDSSg54/yEuz+QZrMX1+Ry1lQ6dqc
Py8MVN1lqFAPbu6QFZTfPfIWdl+vTAX0D1W0wcTEU2zLhBuBfGtWb2c9bCfMDqROjyC2Fbva4vxH
Q/JryOZVZTMOhwrbJEncKez0k+XAJnlMbqY5ywQNEjFR6RnY5SdXifrdGgDUntnh5vozd6Jpgvyp
jWqCqwsZcNJLiVIsDeUQ4/bkSrzN5KtVBcmeFLj3czIXtkR0f/MVTXjkPBNn3jaMLub2HtlFwV3e
VSsyk+TKYJrzYPO2qYHl1HT6GDtCGSASQZwd6SsCDQlv6huUyrPQlCBmS0+RIwbVojxVuThs19My
izqKiY/I6Vq7d0W/W1xUgMRvzdXotZ5fJU1x2mADKh7E1vscO31QyaaSZzQGAqvmgRVe7ryWPHbI
57oSZHZ3jYA3jHXF84JD6aji+SeijK7hsyWzXyG/x6szubKD78/lMZfmVKakffGVj7lRYsb2TxoO
bK4v8mMBBhBjzdicms2mOv8BaFuClY5o3nBXWYT3ZxaGM9kZQOOX3wXnSY33vkEvm0m865QYpcxB
SD/6iC7mUIroB7JVBbmpEpoBgLPC29pZWG+K8pj4kglXityh3MqwhrfT+UwTP7DxFgR4pCrtdu3G
epub7ROlSnDys50+/6dIvHY96kae9r7qrzKRO2aKSEjvAU4aTnzaDD11dguKIRbEzHLyO+nFAP1F
06uG2oq2FptJqSvp8s9RgNkoJnrZsn70KdY7QDjBEycg5XEKblxBWlr6d0OJlJ4S3yRnfR20GelW
TMld/wYiyDQPF3nlJZsT3/Lk7XPgYaN5xD6OTnkpwKDaImi68zNCYuo8uh1YXB6jfOnjZqiHhjG3
ucVJ3vTwr1EUivji/ItU0rNn/N8+htll07eMySWY6Cc/TO898GGvEZkQCLnNo2WLCLmZndB6ZkN2
Rve5ZSC19mvEE6I1bEU+GxZJ40qKaZASBPNQgCJfsyB2b+QvSj/PqAnJXQtTtR55evk01ffmupZq
TS1gEdNyyNCsfDDSydXbGKeSotmGG41o+pkH3d1HQ6Am/AOfwiHJYirQpv2kF1yQl6a4HZCUOSOu
tyhRVMVYsXOY5NjnU2BDZBqPZKUawWAp4xQNHddk3pGMZ95KT8RBXPN/T58wDWo7pK85zGyo+Qjz
A8EtbJLB/m2KdL2wn1O1wBujV1JNpPZvtDTE5WBnsHjsaO2R796WxvTgvbqVuf2L9Zf1UGs+L9gd
JG7yZHlONRHzbei1aglQTjQGiltJHV2bhhKnPBOc1VJF3Dj4ugrvJAIVwgMSsZNgxhdzCcSr2h5r
oeWzRrmwBsaWH/qBdr/Gh/wuMYjVw1on1dTk3GNsYK4EGkVcdTue676sQP3TD3/B0tvTh5A73zct
Qqj5a5F7rFg/MUyTLZS/KEOXEajhuFcupxBaVPkKJkdWNHNbez+EbyhpEAf5PIcNu+iEBM3QZqaW
b86WiRCWd1hS3sZfInBDeHoaCSuHoyOMMeXPmOBCLHv6fAwnwE4RuLw5NMa1Qwe4EgB2VYuU6vL0
HZ1sMNr87uPXNkh/wzvruNeahPilO5dMvnC7bvun0ZKsMRfsYeDquXuDKie34OhhY3/C2L6XH3Sb
CUvm6udA6f7VJSj3BrP/bdY691vqorfPZkLZDHeQuXB+aBblEkiO8Ns0TxXuMbPSKmoebBlj0qHO
isUfzCNhlNdIip+kGw5uozvaLnToo56zddp3nsP0fveeY1V2d73owf3pNISpup9ozesDpDaFyUxS
nJjgqvaQYAjSed835z+zx+7OBxX81gdEd6Llk1KjBhzVxBLNPZGQ9DApmpy0+lJDFj2hUapQqro2
xeZbogJHh3UVpvPLl1i1FT2YvyA9upE8CcsQ/ikSistry4gkR6StmUbSQ9Jsk85Z2gx+3BB6aqH4
aalu1Sz4Gl7vHTqwgtRRdD3zG5qOby8akt/jIpzukYONYku96Pqz5bg3LaM+ZgKnrwJPDL1Qz2dP
DG29+aS+jIkHNZFvsex9l7b+ci5/YjWiJWl+4h4NKE6U3SVwq659z275JlShCviNDZZo9+wK5eal
TYoZ7Z5drE3KkOQe5uiSRWJrkGf9CB7f+X3mnfpv+2+PBS1Uy086W6JQ/WGKwWyybt+xflbmrPWY
ulGaemkvdcK+d+BL1fTcAWI+nNZ3vCMAI1cpJ0O93n7GE+cDsMpkjsZRz3qoGbTxENbnjkRsGhSZ
c2bb0n///CHXmpdtn03bL4VXIFstWXnxi5Y/2ym5rHMtQbC/rNfb6WIGd/Qz2T1RjeGE/aQ3Y9n9
Oyiz0Coi79/Z3ANbqnKn2D5jOSRhyL73fSxwQLJFkkwQXLju1UajFWB1qrtzBzvi8a/Rhcyn9IGs
8iK3Nnn0o9WrfBBHACiIVmO1hPIELq02oxcWlpOSZ1pLQyWFvXXgFBTMiivzU7SyJT0Rmm2g8VWR
4bM7T+qF6hw9yXwRnw6hHatJDN1Hue+IfJAOcx9TUxzxzd7ePlRSfCDn3M3g0weskBPEHxSQC37p
q8hfY2tKMTiOCI/VNIeTwRHOCfZ7PY2V5iVw51+Y0zlmYEFVouIzF6afb2wz/N1jL8B9U75vRj8T
S0GFVyxou/DawZ7ESpPDWC/e3IcbhSha20CuIgNikJMOFLUeP3XZtcQNfwO/09TmjJvxzB81BJuD
lwk8V2IYhdDvmirXmrOqjyoRzKmQUaaDuX9Ba4SA9xb/Xl7w/6rxaTjdxgjhZ/rFzHXtVv60o4ZF
Q2jiBvi3rjXFfdz+C1C2y+4NDda565LIIT7YBI+GKdpj8J/yzRY5P6D7KBAqvfP69UOEPLpTFZyV
4oamPMBCXulSuHgXlMZKSdAdIfVKGbard0YFM9gACijX2bErUIs3QQQgCw9x7jjqi7TBsvCP2J7X
19gV1harwdZGRYEGYKVYdCueFzH41Vy26//IAO6/AJn4vkebHfWkP/5sJhAWBpdzUBWEtDAsXJcg
+oSVzNYvhM7VsgSt9/Yf6zmG/2eTJIbwCSDj5KNCQ/kjgLf5R37PxArILGr+UyRYkWjt2OpYxwEM
htvMo4SWtKz1AF9xPZG/1sa+1KO2FsWXem5sQYXL4nLHHrwpS0eYHz7YrC7U7ns/hJsOqw9b6wgM
kayxsfLsywK7L0tMG52KSI98m1E6ZXr/aiN3hKoXNSGIt3u76ALVNJh/4GHsYFuVRYVflQePFzkb
AJ1p69drru976cwy5PxyQ90Z7qZfv1TwccbfIyqMC4F3g/ePBWkd/z15g0Qb0ite38pn2cqyojbM
3V+m0CzUwVx8qKLCRu1jJgoBSUmXwtQhZFInp+XdPDJMS65AkOY+/mjqnDFKyw9qtW85HeKypVXp
fiZaEbbVwe5fY51WVGP2jRU6gkuaWRVXzB9egUQi7Es5iWtEM8ijcLcitH/5wP+epLFlZJDEfQnS
cuocpcn0CVn0jMJCdr/XLqTyJzGTLHTDRuIg+jKfL9TV/CpjWtlw1OWT0lHHx4br36v/mcfDUW/l
9YgVSXYssj0zIAyw3OuUBnlkriiiqZJ+4iLmCT9D1MPzrnQV4FpR4IO+Dxnmh2CSvv+HNh1Ms6EI
vR1UXqB8zELS8LBoCRlMKmO7Gql0qpK2phv5Ew+byiUmPkGrWnUUOfhGg9uhf4BbsSwuAVLEpOF4
p9oA+MkDc7V481kC/JYX3e2gTRkBjVwQSaVeqn+S8FooSJJBeG9i22xIIh/PlegrOwnwvFW1WADm
afPBCAkthCtCseFY5S4Y6d8cpz7x/VfwMbJyo2Jel977C6W9CJVbNlCAd7pce9iYrJtzUiKaTB1F
5zPbYZBfO9EYgaDcpDmZr4Hm1exqgdQYMHYGg9vvPsF/GA8w8htFoLhsePwuXPI0GhIKilbaq06P
4F8BMtN83KGuOngk2x+TWO23J8GBCwoShoZX+8T4NuHxYnBjTLKojq492asSygzyky4GsLCF2Gc0
zMdR0fip92iKwYFiy7wbp66EIhV2rCgXblbnYa1rejjdIWA2PPi/MhPPH9jgtmsnPE0dSkB/cLBV
rAY7HNhN9LsqMcSAujOC/MoNemg5KFuxCsVLY7SlhtB700X3nVhtIbQXYkfD0+PrOc7ORO6Ine/e
iAmZ2zUeiGodHNbNNccxldiELfPEfL5UuVTrXZKN8tuzq57RqdkSeQGey28XjIfST9/8l6hp007z
GAa1Aqe0fkTYLOlNQpTewmOJaEPqatvnZcPkRpTVQ2O+fI4E1dGvD4Bl/Gw1jc/I6GSe/JZBFj1F
OaYEKAStEQGAhSmsBhsppevL2+9+4yupHtf6k1nroKq3F4O4NiuME6NoQlfu7Fhlrqq4H5X3XkUU
WttMKLXhDYiAZpGvjMiAJHECHNLD3ykVvxlHHz8ib0LQcCyEMRCXHg+OAJW2kzZrPE9LDMUG66yx
ThqNumR4pxeI2Q95M+ioIT4rMnu57cq7HZ9DbYp0T298Qnwx2f/9zyJvDaLw03JYpec4d0/FVZwk
If0/59wYplvixdxdBwh87agmgISx+NBztq2jJqblkZBlsfkQe3DOSOMv1VePQ+7oPcu0Oq7AKAUo
FwDNPAuhcw2NVVISylvKTiBjF8TE8nx+X1qMR3MIHoBFMehYte+v75MOWG2xVp1osYwWxCSGljzq
rqDlT31Pi+4W9yO0EUn4Lh5Yw3x95/wd1K0+fUXa0REgMAaNrP1CjaVn2d7QFcuRc4E/vfbkVOh8
uaG2+zyV+ZSwJ+PdzJiX+q+WJF6hr1Tctl1x7q8kfmgWEmBLZecqcDIlR0sY1uzoHiiDfUgDWxYg
V545K0Uy4iLRdcn+x5DO9Qrazm9uGVPRCMK8J0KLolhEuqleSaH24Z1rMJL/ujwrcZZopmd2teoL
vDLTKtsMbBW8JML//3m4zzVPudbW+GRPYOlOLn+C7UTNu7Bqo1pUbV7FipSW0jvPIqF4Q83AidkP
6FbGika32wFCTiY5Tfcq7f11dPNsB9yRjB1k9PFzz/D3r+zMiOUthkjPGrdmhrHjN5doN5pid/k3
bFWrX4hasRHXtrUtym3TIGQXSxjonlcUwlvA8emkRqyYPmvgUx2o6lAz7g3ry/5UWQSvgAEazTLj
8psz/ZVHKlv7PRrllbUooTyTs+zGy6qDOQGNSLgK8SnssWAItbjKDHdbSc4wdUqtzADsOHiGZwZN
poGbyr0eqk507R9QN3YsjSfxPfp/5yJ1BxCkv2Xu51uGanJh7gXd39VT+CXE6SrxDnoVOY5NCCtl
4TOknPaAa7Z8FgQLBxUXBqq+o2XwDV6d6duJgtQa9j0CZRUhutzqbn+keXZ6eNJgLp+KBEIH5COm
wCttgOs4P27jXawd+y0VCLELYwBktr3bR8wuqXFOWoX1SGytF0LVtLQRX16LXK6N1JJWmG4aklSm
VQEYX/UuSn8SXgZWe0hQ/xJolqCvd7dxSfntz9jCDA7KoTzcBgdJQBjnBdNV3L28tXGp/TIJlyWX
c7ULVeLJC2FjqxAddOhPSI3zEO9W2E1G+hPC8vkXwYb06A4U4pQ9mUe46R3JEPWcRD7y3hrLUCUM
QWD0NwG6LgiRRHxWBgFQv6cZV3TCoYOiSGi9+dLxk6o8emG5RttAjRjoXsA1mEt9DLX6UdMyQPsj
7oLhZu95MtgOHpE78QpOuC5hIDLi4IYCs76PbkGLNTV8bCAp3l/TfvU1uXnUa2e2kgCTx9phLr3R
juiCQv86dPTTDzX7V2Mag7zNY3oJ90TL4eHTgFXGFlfWFnIfo0oz1Ap2EUAU3FGGpJdsdA7b8V1z
7X2xt13wNitwkIX4aoMg8sNaB7ddF0bBxMl5n/sbOH9/Gn71q3+ay9kP65z8Z8dJ3qWeGvNiW8xp
o8m3SoZeSP/ndn/tOXQZSvDB2v53mIXkH+jy/yQAToDif3HcJISdQGZn+BT6m4Waw+VTRlUShhAR
q5ECBrLzQ3S8B7oIm7fUiCKzkyTQUrSU3hCSPolPssTIw52CZH+mmO5kx4YtgtDEgC3orTZdmh+H
+2fkXfGqUoKP9KsKzrfQJuyOGdx74D8ZM9oTVpr0buewIvlEsfVsjwnKxqkqHw6zRq0PiZtO8gXN
Wz18jjrWOAUzbfCeP/UIPMBIaOGGp8RIQmhpVfWEZBNztXSGb785Zdags+kSnbj4KnsdQS3jYJRm
QELL368CxFfg30JUiCf7Av/w4YTZm3EuZcy/MhNXhEwKju4bUVgZJ86pzuuul2dBbNYLozb0hR4j
/IaOqBXeVnEh2Jkygo+RKHv2JaM929YzdWPfoqaueQWgr/0guOjlqwujkPaahkOMNC7ooNIdk2wG
xMyX1QcPhZmZ3dPYvd9z4btHLv3xpG1E4mvp1CEJ2o5M8Z0dneNH1ujgy7OEyNp/allSgbisz7Js
O/ORo5Y/3ICuE2oll5nvbrA80B4/pXt5n4KIrRMidA1smXVJQJshxeOuCQvcxrpSL3WKk+QzxW22
9VP12nrGYNnt1un+hsXmhhI5grAgjJYiH3S9Y2VcRlA4fxMgZ6NngmmtQqBYo3HEtfXNMqeVvjTu
QtvWhSiKXZOlEBniHid79kUBhLDRulD0QAthK8aBHFW3PifiS3Sn0Jb3SVWh2t1E4poFEOPskr3I
CtdH9+haHeqsj43Yq+gEW8WoTZ/Mp+4KJjYM17xsBSA0aNF6fWAIbwNVabnmM+igZrMQj8F7gD9/
yFeTYKFmDtSgEDwXrSvjzcZWS7jin7yRk9q8yykn8DN4oVZ23dHA6dec2XVYrKHpcVPrizJe4loH
c/vgTdP/DEYMnfA4KwYC4Vld68YiecotZjXZrVct05XxvKdMoLrKDrM5AQ0YMsHjH7UWS+cKhJcx
PlPj0soowXtOIZvajQ730NHgmlLl2GarC/tbb/lIT9PLPDXUwugi7Xe6Eb0CW69UdvrDZAmFOQGI
j1e9VIpxZCyXgmYq6tNyRcVnkGrpJpvL+EwLpc+7rWU8QAlRU6jdRzZKdkaSLQqtePytPKuxYUOX
3I313DtY70OlooKf1mWStsORMTMxs7atCCcZhdsBVt40Tn6vSjcw89GqWAllPskOfhF9VB34sF65
hs3E92C3aIjzPCre5uqpJ84Ix488Cd8QLBKO+k1QyDBn4tCJZYC3NAFWxwzEt2mMMIHE9u5eJ8E6
sMsU+cEl7aPEx617Np8SO1aHfsUclwkgbfkSdT9AjYCkTaMGDaWLHlwRdFiWUfsH6yEaKBLSvrq3
hCeDDbtsHcgLL3YjBY+kX3821wK97tnBnRcwn3YfcxfkYrb+mPbVC9W0PqnBoOrzRWwErh3BUUGI
r8AyeGyaAJsrq1u8W9WlL8jH19awJBe7o9vDTZP1DCvepkaWJoqwse9OnXtLOlfAv/8mz6SHhdQn
l6023PoHUyitIzOV3f+qEFWKVCtd5hou1MxPIlsopdgZOova6/4FqSpiCiLw5bPJfrl1GsM+arA5
mKNW10YKkURD1OmetV8suV2NLHGQ4sKQn5YJ/jKLPPxxoo3Ag8lf9iaDtZWhH4r1vgE4g8x1k0xc
QrUn4zwrjzupbjBzQAQh7tfChMYcWXnm/j4BXHAMr+JFGRmA0kUkhLwRHgCcVIaqFDgyCLFP+Kjp
AsTfj7mzYpr4mY3k5woY1s9z8DpG1JCR9GW9UlO6orkUbiAp4lA2N3wJkkoSN/wiTWZBIw79htWi
YAfrYfZwyRrLcGwIvozf+rD3tpwC/4VmkaEB/RtKr3QmakbFIujTr5blf0S5PmqDMjMB8ZMuF+2S
3ImICOnVTH3I04j6LH8uXAMf7iFKkhnP7fU1fkTLp4R/B2ph/3n1ZjU/6AtoO8FB0XlUj/0Fvg7U
Q68ZwuZfrkZpYfzLsPNw+YfzeuASM45VvSRiZ3kjEmNwJkppCBSvTHVVmTNce+ewu9XGrODQP5ZB
NJiPFrCXAE/wVpuqUXxn8V1WMcTsSch3kH5k6hyk75srYNaY7YSNQZ4pFu5N2HRwvoqz0epPuUDo
BLNnkd+gWLhODGKw9+iyOGifWy4GZ32TSThHInIN3gWwZM5kBssfhbvwjO71LHzEKDfm2Sca7Qu2
DCJhlm67NZl1XSnIP3eHeOlctePoGFua2g8ksNYJ8HQJ4V4yxSzGgZ57pSmGFvrUUf3eiY6BpHjw
YS6U+eucfu3fiE6CaB7dRLmSUfwLnEIW11+gcdOv/iUYfuNOKMyN6AruqoGA9+GJEB/EbMtrU2aT
Izw4jw0+00Pw8sMInBxJL1Xs2ypg99N+twikxKUzAhI3tvhhtfFNVq4k+iQV2k3J4mLnR+dukTlg
OMXy8k1X0BheXKB2sKjLPmLQQ+7Ww2KFJFVt3q8nyx4XbAZLV2qqYClr08Lx0Z3hgrrI5K7hGntZ
+5Vc/WQMFbT9lW/IYXZIDsgQSOd0aMAIeuWnwJDDUuRSGoyC68e7ljS28w8O46goOpWT4y+cW3LA
+wWG4dllEttXL6eOrUH2191Xm+1mwno/as/bn1Kg9SdGRS4G/oi7+cSupG1UCCLUfO2XVqGwPK6V
rC+d833xEECr0KqPkQrTPfq+DUeBu5T4B9bzIxP1NL82l/PamUdOXzYq2FqUgbVPtR0hCxXuglFt
8XGb0ZwXrcAOey2zoirL45LwIQoe05Ifx1CfgTgdXh7bg41HFpsDH1/0gEQB789tAoftpswwLaLQ
eq94k9C+usXlrm/Wpf1lsnbHP7nFZGex+CvcZBfK+jgp8vFdfRf+EKatsV3tK5PCMSIm5llv0O7l
RSVUfeAHPJVMm5/WnCcF5DN0qyDAPJoqW7Ivsjgr0QMiutJJrk6Guuvf7shv4pyLDyN2to32Y6Kl
iXt0kb049A8SzN21YP9p+y4pcCTy60NtBWDjvfDnPRIQ4YP/M1tB3m06iLy7RRVIDe+ZTBGjeoqe
J18X4qpBhTQNOkQBAYrwZzavJNP5zapLaN+NRohrEScwZuDMnzE47cZNrPc6Q4lBQsSpGbxyg7zM
iG2FlPsiITJLfpK6mOWksmwEWKcdrNVg5og3Fw2gQV+nKR3fTFRsyXDCGAE17tHNcUuG3AzMzJCF
CDRtLPNsgVNEkV9wcmdgRVRMYzgNMcc1hlg/4cAFccTr8qriq4uzVuD+BieNYV0tV3wQIYwWADiN
zzWDT8N53SoEeYWfRfsUHvO9Rdb9EtgdszRZKV6lb9ijnkY6PHv3OPkhmvxJeNrc3cERSK1lA1rE
gmSKMB/0mnloRT1rsqjHkPaLUW04cieV4f2W7I09RyQ7ATL9xpGodjOvhyWUHx3Ir+SRYe+twUOw
S8+sRUAUNWMiPsRbmADso+s6c54eyOVsY1e0DGlNvPU84gwBT3XH6PvqTi8g3Qkf8BJ3rYZfxzVA
b15sCS2beJ1yxobAdvVJNE2K4zVKbj/rWe87xPj+2bMoiwsMLajJ+MA6wR0Fyf+micTV+sqKW6V/
fdAMhcY85k4WYFL233hxe2D88/wOAjd+/IkeYmIiIdaeT+l+a/Slas2x/tVX11eovWWE6dWVnV3F
LYY85UFVOIDdTc/tpev8FyuLOsa4JkHB1IdNeIzctlMh76fbhLVy4FmtzeJY8nnJ2ORNTyKSo/EG
Ov3vZwDBrVhtRmNLDdIVHfDQYZt79SeaA8KqbbGXI9sNMjacMx4oZchPYZ1ts04Twu9ZnOMiImrC
2QYpNFOWertUOxvyLf06oNUQ2Lthtto4sol70JpcRp2MspYyzT5aiWPlCFQwqkL0Z4XfMsjuD5iA
KqDAysLPXIJvqXSEHA7C1ybZgLsHoE1WyQOst+oLv4jCbsHWjMU1KoSjTLLGasMvo9L8mIGz0NGB
0wpRZojJwUsdCC/C9eb52njgqdiXQ560fB/4Q9YcBsm2ZRXCh0FJRPR0W4JiC+HA7gExv91B+Kls
lgqEZMhBQsEXSze563BQYMmMB9/KA8Z0PmUbTpu91nZ6LKfzihZUtn6BhZ6ap7hF4o4w2AoeQAVV
mGWkB5Xm78+WjyPCAF2QLCcsxdaxhw1a74NHpNGryff3Cvl5KRaxmcQSGqdOU/9bMkHCbX5++tID
N+QGNIWseQdfJEMgb/XiyB/kRLxtBFP4W88whwXtnJ6fY3DqRUGAX3dZBwQSG3NWbj2cyShakWyj
PkraYwUQgqtG18GOzoS8Ko+NkomW8RwjaflLX3nwbGokLpiqe3ZXby5GDP2E3Pzy7VpPG+De+jMD
uY82AmUjaPfsmiH51kcJ5K6VT0eQIQEZiSAIAM3AV2tBPCTRfZj/id3cjme7OVx6Oh0aVMUONS7r
LhOCj+QRduPOGvFgEK1I7J6BE5WrqT3wm2DYaHGZRtDGDs3Kx7NBaaFHkcUqkNo3W/OyuJE6M9ck
SH2GC+0PR2PDBRFnaUusj5cUpGKiPM/VuUp4z4gjdcF5VJrMfmQ7uoNb63mfs1DnNNZii4Ip42V+
on7nL/KaL20+xW4ZbbEHZemaKFfMR/eXgz5w/XwVcfTrZv+btcGCyY03dvZwqPCxXliZV40zCSBc
W1nU8vN5QVWF+eL8HNGCkwMnb2pVocvM62ZswAQdwSzBjKKM7pwe1lSKOpOmKhGibiprinEyDvUH
HUWnasIzF5L25O6czXz/+mdx5DXYwq+gpOcbstbTBHhY6z+SgmrBdPLHt5xkvlqs3v1UDmIEE2nd
PSATqYglnkDcDLAtfFxH+FNC8Vn3ApnYaW3eMzeaFBl0tMftDqUtQ9IcHe6QyNJqOlAT9fHO21uY
TlrskBtTS7QYNsC7OHniKZWlLKY1o1RxlX2qysMl5gwD+3QJXHpW2KeOrhzTiHvOdXjfAxi5+3el
Yh/gakk6dp6P3r2emBi+buZvmEV7rXt7nNXs1UGyQYFOUBC8yOoNS2kD0iCJp1YC2tu5ed86wdcL
iDubW5k4t9HN1084Q/lXoiBglGcEQSnRT22e41YgFYMrs+jhadQXK4q784Nfmooj90ehTwOwVVcz
urLLLrHHhpxqsKVtNxDzqZIYs1j4m7CIP3hetN596Ht3vE0EITl0NX2BnMqfq7mtcyeY6V7c9sUX
KqYyvpx6a+J9DvBdTz4nPJMSOl7AGSKLzH8eouts/6MzolfjiUQv4BHqD2x9z3jOp47BiaAL4MPD
kpfbB2ic8xUcd1ILe6CBfWgFJjnZxMA2flZc1H705l2bUu3KOldiMqGrTb/tTJbQEsIFlxjEw/1o
exjcXFW1CnUf5ZmTcLrqE9mzGr9XaGr47U9H07DzXnvJt+QEzsiF5fIYHl6jJqcb13VanbRtXNI/
/klewdLvOhSkrR2XFf+iNt319Gc4PmPJdoBD5I2TbwA9BtiWmoT1lccw3SzkRc4trdWrkuh+6Vb0
XI9xMUAPZRbAL1fqGqvYe0b5j75iTYTV3Z+bQJXuc2Wj1FbIJeZ8TjQUELpU8rhn0tsb3VKALcX/
0IK8l5RfUrTJ3456/y+OLRQ9zSRUQe47VNL3ssrHqA6GiIGst+3e1ztr3RS+YLivaEJFaUsBiGg6
FPLVS3Qm+Erk2DdVtbgSqIAkz+ZCrzhKD9qi2+X0ewP0/UIekavfVKBGJ4eiR/6DDjvlMn7+TQny
JRuPKKaBBdAOh2b7sQa70wsgK5Rpvbuyyv+2itVMxuFD/e8yEi3dlbpuTydCrGYyU9ycYytTXjw0
ukKMrw6lLlRvLR9WoYbrFK+wCbHe1sGTHvGEQ1bUY5/sEgMvVebCrqzsPnymNwpIy886WO7rWZLL
mTh5fuTJVPCXp+T85kh3zioQZ9ZuALN/pGDec7incE+afok9ELwy9EIQ/GmUAeeJnQ4hV/2KmowU
PbGn/VbATUbYLBlDbPhKs+Y86RALjMlwvSERaeeigCWvyGlQX43wexNySARYYYG4/p+wAreoWqtZ
whOO41+Bid7C8jMgX1ANvEDkanw11FfAx1m9rAAYJzFqDaSz07kRa0KdPo0Ss0KHPrVFQiuH/J2d
i7VubV2JxQO5MWhEsBJzzUeJNe6q3rUgQk49yhSPhrmxgQcLE12psLrWWHMn9RNvlFWABwiDNtn2
Y98OC4uoQ7PqMHCoIlKIpG/xPOcIqrBmSCA7Hk9vaEaqalp9OghRFnQpMg0xNTvwo0cNTaj+5RL4
SPC7/jTWv5CjiuFnzv7SP2y9rH8SsBdGhORGvUsM6/o8asVQEu6ZyIb4uS+DxpgsN5AEdRuwIdOW
ybM49FJjUKSlwd0CVMKb1OA1LC2S4qaiVrZPpiVQkJswzfr8kLhic9IPvrVgDe4/YxUDmuL7Hgq8
i46oXdimbfNUW3CWvh41sbKpx6TOwVmGUQXKM3plfTsaCeMIL5GEb8DWqYD19worbm3YPkEqNsHt
S2finoCn5RowaalhgfLJ1xflL8FiObAGA4X/+eZ4Wp/E2c9izPLTgBVab9mdTqFNpJO4bLgvtmKT
9A1o6HRJmQ7CS2mnBv6/ctwncYxuteKZwXDXuobNIbkS9k3sNDcf1E5Epw2NIV3lZUbOmbw7pLhL
XuyUnnqoV18Bu39EvR043PbZ6WC03TV5dto/ptjIfMTz/XIrFuZ3IY/fmuYMat+C/DwIsqjIMT+V
taMenzbSyRku63oK66BqjmpE2RSaCaIuMzObzRVOqAhjXLiWrRDsulZHLZpeuzbns7VmOfQR2AkT
GGKiveGf/6u4PHwLZ1R4NvmVPPHrHMGagnQKRS7qwHOcgBRh/uODebHXVNA16sMY+o73vvVY1WzM
tGFcMfKj75F7kGW/KkbXx/y5tBufxDfI3pSGJTlnpjMREXs5pzbSjlzHm02JwB63daR2uQUXjTmy
yDflc8SVTBGfAQLnt7GmtwTQMdwBf+DrlLZv0/8PWWVHGEU9Mu2wcNYWXWBKjOcJaRkqmQoNbbsn
csF9OJDsN6vfWKcKzCRxqWFSDtDeEYlqeC4y4DleP73jQcloCFB7dxQd3ZcPwaBZQw06hJydkspq
y0qOfGKrpynEG/ScPachuOLu7jjXSYqi5vptlIDgZ4TqVs5SRViPJdmtO5YHCDk5SH+4RirlkLD0
89Kk+N3kNHHkSTqO+jay5bK7fSN7ToKheFbfAjs6z5qFTWiU8ObUBgnb81lAIy1IXDPav2skNCTr
tWxZugVpSP9HhDf5CHkB4SNV6b9cYeLka6GM0GaxTsbY8b2ptsZvfAepjZVte1xdIx12iwlDzkvu
HUFq6O0YcNrzQae9CGYs5/n+FQ5I+AtB/B5LOQcK1M0hv+ZmqwKWHjObnTbspwY9IWmdP8XSo05b
bHs8psPT4Axg8Qmww+KQAE3STA8yWSIlFm2Jetj5oXrTPZjQcAKIgsPx+4pB6QlIlxfcBJih2o0Y
lheNEAzN7Mba/0t3Ka1giaQrcv/Bc3lIK+XZpaxNXXHabQmstn/P9ZFqc7iYSDqrynwnqXKHghPw
siVu1pxRL1k3x0aS+ok3Cp4BR7io4K/WGX3h/LQU8OKI/J6eBX04sam+HhqifMkZS3vPQT5xCB86
0+GlGmhk0FCIy6YOdOG4VVeG+h3itxn3k82EcOOKGpM5+TP8ItaduAqXLJ4Bt8h0HlXkIaJ1Y7al
f3mzee8hw4mzIXrSO2wWc7RHR97RVhIWvXUHFRTbCcS49vdvdL50VysBvV6Q9Uc+ELb9hMIlJLp8
5217ElrJywKH8G1l0FY2omqvKL/OLksuQhuzYrfjIEWX3xkivYo/G5KXlOMLeXC9ALLaETcKHXCx
a21oP07jN+MxDHlY0fNXGFznOchJLR7SrZmPyT4PcaClizBWrUN2R6Ee+GBhjm6W4LLsJIGxKfPs
BWcbFEgYR4Oq2A+9fbi7WbsZB5lJ9eFWKuh3pHSxn5K0KZokMhy0NOFMgyiACf3+Aldj3N/UboG3
9gAv/SUWmmfPJMsXbkk2NNNHYYS/2S5fOtk3WLxrq6uWIX1ySR9xPlHYFZXmN6eAIFI2eB9on/OM
BFR6tuUB7i5/RtKjGUJDUWIz/eH2s0Se1ED6u/Bz/WbSAVGSdqjRxN7nnkEifccIPA1NTD0dF9+3
q0NVO+CEYYI+E/VL7TlX+XzFrylC+0XKSnjVjVqfCduGn+IA3iRyI8F1HU+o/Wn3kE8lzc6NGw/N
gwM1g4QwtxXJDoUaK3SShVKVUFH2aIWUY1nkfyj/EFmCIq9l/r/QxteW7ytQnH6g/OnY2UHHuw3P
7FzWyOpGD0HYvBejPY8FeCk/U9xgHoHLUe0H8KnsW6OR93U6O60GME2pn+TWzbmFyD5JP8HLb0TU
sL7x/DJfFrh6NpMbvishTnKb9CYApbXCXwcYPAMjRIBT10EwnH1yb2s/QocFwWFSYkHiL5d1pcl3
lOlX8LbdkNHH/p2CrhUPNXsAv5g0V3Max5wSs/mQyjkuxiufyDVboPfhii0bN43ZtipkjcWAJSJn
HSv1Y34eH/xiL0rV29/A1d2tm9mZFYaCi+rQfUnYzDn7q50K6+wup7mtCaxDzlhOxeZBitVN/9Cn
hofvfA7vPS/5n9TFBizPpZF3Np1Gvce82IZDpWeN175i8GtQ40Cs767iV2C0EFr9zgD5LPizPNmZ
DCESO89oPabkoMiuJ9UOEUJs5CrFU/Rx+Bq75YVVJXqroXLCVhX3q2JMxYg4T45QEKP6WEx4mYYM
F6CnjnHqCvJzQgAQD2Bb8L1J5Pw9Aj8DNZxX6IOO6SDAphYKE0t2sZRIBdEhXFfYxMnRNmyxDeD1
JIjcGODWNERSNAzBlrVh16Y+l7lJX8KKsbvZnEjrEJWloVuQVaLPnit8cUM9OKMrU9X4qFzWBM8w
LRA2n3tbvpjOmKVQZpt+qTWRZ6Zbq5tOra0lt9mfgOyKakmgIqv4YQnT9PvpTW1oofzOZTnnApr2
+EJs5hfOabRZfTBfK+RMTorW3D02lM5rf1PWV7cEpNqblKiCTZJyBaZgpfdt/abxf3yFG2CCHHyj
FKCogPt/Re+uUYUY0D5y5B+x2VqP3SzyratA3WPZ8/4gk3KFk+CaVrDfiNYKVerW54ClgMVn1GKO
w7bgSDOaBMzIQnhI/fraSRii/MHROivS2r29xJfTGzFPGmjemDUymto8IWy/6HLz01B0lC0AOu9E
/O/Dvp9ygFvEMYhZw37i4AXddFH0s0A/3KreZWw+6b22R782V7PYHUvFgGQwW+HNiqi/fD8VoOW4
72eXD0iWw10bGzwmzRc/GzZ07GSiiGHhk17pyBcY73h8wtQ4ma38EcvAVAasYMl3ZC/lUHO/ypqN
R2+w+i+iNNs9PWzEZvNkf62wejZ5R/QFF0ZI3i5eeJpLCyIpMgV7UVIq7yPH9kJgFfJRkaU112Jq
qIqY5IjNFsE7i4rDjJIrpi0U+SsvvXtaiz5n6mxPHD6oGJllD1Dvc4wudIodwu97FGmwI8kGRFel
sagoK3dTz/vuYWUfkaEJcKcElgxrDRpWdFqE8Orfsk9xv8qUA1l/NmfmCLdN2ne7r7hk7u2nSl7I
PR9wErjvg4i/+n/u5yS0zhfRf6z4K+MJdM4EiMdRtxI4xoRGYj1OAwbWaTtD8s/z/OqjqjFK5fG0
4buGcKSQcCdX1ogetXuansojijb5srJ8CDEXVqYlJkjN8IV41zi6RwWfnQmNm/RXiIRdcqjb8w6a
nHKYhrJMJwOuY4UcbQ4WQbLwxbbp+oSq5RNUJmvUSBxsQkH9s9q6lJX95Kx2kRw0vuzuMZFEwt+h
wiI76p5UnD5wzghxi4dVIf2orpKwnTvNG07SyeMYq+PbzZPiAAyR8DkS/APPS9MLOzOhLtqtpEjI
47TjqD991FoewgUZachC5s6OeX0x8u3OXXAn4NbfeyHLJU4GY3igpYyu79+zO6igNPkTfjm8+Raf
xkqEVU2JPSU9pwPWPpcLSm4ZayK3QvtmVlh1bQ4wvDn0XfI+4qG3/d1ZResE8n95zMa+xxlpgE35
3ffXh6OAv1k6xSPuOM3riiOupkCrxnIQkiBhlviGFjOTTZMULsnFUS3ElZRWjAuC7PYZ1G/w2YIy
38CNn5UEvOMV25sWm9FMHi0a0llc4MVcP9n1Uz5ExB68v8KM0kKqM1w3KOfHYm86By2IUeZVALBV
dZ//SdkfMD+09GYCDM+DNeKlkBpJizGSkFB0pc7HrneE0ZGkEGetjQlf4F9/CqU0D+JrHMOK31dc
CCBfC4EUXf36WcDQc9fdWL+PQm17rI6Tx2aCrvnvZJMSCFi4+ylFVgcssji7d824k3XgUOEN+luJ
JOnsVEugDirx7khxEpPss5PrUaoRYQob5eoGcAleNvnq5IDIc6oC/xsCQZr1eQjMB78WuATghmB9
Pr29SLJl5iLk74vPc6N1JHco77TOergUk2mQzdfr69wZu222LYjYM6wKYW4WsNOnE6s7Ri9JtLO7
NOwdcJXEankcT++50vbjV+BfCqRj8uLuPIdle15APdWVPUXneYCJ58SaeCFs9AkiusKDifphUy3u
CRzh9PTzK3RVxoNnAgl9wFFPRNr+ZWuySMIobhXNxWNA0Sf+K7058wYHVR5JquN6fYrKRKFF8zE0
9tSzKrQdg7G0ZC1onA1b6/JibI8JsJWo6ISlm70eka5sT5X135laQGni/Uz3d5CTfqB11oNVykpM
M/s7GKqDmWRicmrjbixBO1io0pV655UTdq1e506nc5Xcsnku2K76WawOBg1wXx940hFz89/JwAzB
fRRzaUGxc1IPN+hBm9eX/k941Vn+/1FRce0ngVkcvPboQkgWPw2XUMGkIT/inurEZfdlE4Q+4Yic
fwVjqgtdNsoiIyezCyhDIDJL+oHgJxRGHN7pd2wIatRQHE0yfkjC/j3j4CtEX+QgNYHs/y2UK3fq
Z5i6VdI2Eb163U19bt//08iid6hSdyRB8Nt9jmSHttlxCsd9ZWYG2EC6Hp4cLtTTN8FDEocrZ3FS
tiuznSFAoGC7uMt7+aiQ6gs4GFq8lltSHfr1p286vx5IcHY+o1aniHVkVCMaqiJFu6NbgXU2Sf1H
dBKkT7VihFqPqsNDXQ8F1Yes277/2/2XlTnoBkCakiy+iIAZJZvBPRm7TCgTnMZ87p4FHbGYQLFT
PA7mlmNHP6Iy4XJL4+adDPx2diXF5EIIWM3B6WIb48YdvaAg2gzNWg38hcfSMJ6bSa80CW/8gAgb
2HBn3vQyOKBYsK4N4Hv3Qrod/nUOd80foag9wg1RYdWlJjT/KF3cFLvLoRh/EJ/l9jvqLCqQKIaa
wQLoudWlSxCQcrQAwHvqvMAuxn5jjRIQxfLExGl8iWbDErkQ4ykKg3bB1ij8FeaQRIZLvdUk6NMw
XqJ9sacgQrv44ZPU+A26YS+JYLRE1tSInYK6sqS+cYmF/BeGv9FafyFI6qTaACZwJrbyOCVgG6gP
4uMc4jdLGYBmYf4jQi1YP892c5JqNZCfo/EPEQ1KTT0BnlenXT4SuFiR1PkGyzzCrUvFlGq5JaZI
Iki71Rm8x3ybXW2VWun20GSpVgcRR54J9Xz6uOCVEs0BN8VnvSX3MPReRIozGxGLwkIILF5KFsPg
Qw4l2WDJwnNygc2D6DFSGSU51LYeQDClrIQPM6v+KwuOzPXfKhpUND+rccM3i/zoN3Yx2Op7Txuv
eeTiAuuJ+wuNp1GW+UCUiNdIjiUMYIcklua7GBOY1hYNDaFGSqBTbiTK85zgjAfdVe0mHh3dq3q5
zJxmgLo84k/4qN47cyIrPKBXWR/lgM5jLzvA72cq1mvier5m4CzFSIr1rpZXyszQ9x8/PdeUvsgX
jCgWsfh6CWt3onpmCnShdtvtxXlkr0XKszW+122UISQBSNVlg7hTMs1bIVqoihcsKCULKgth9z6V
C/vM91hzR6sBvLDU/XPS3EhsMSiARTRMJvxClvlwF4VAIXIwiX0XJ6sImsWUqqzMll1g51xRgLx3
R2p/7wX2GRR1MVLEWK/SdsaiaB++u4qXR1UxA0Y6x8SmHk2sygaRTj/5OYZl45GDu0munyfL9I7z
QktmbWR8oMbWFpJzA3XMAddBDNmeBRo2d6+DaiFbsFBWuRzwaVb9dH8uzvqlpAXwn3d924KqyVbI
5LsO5Tjey9oBHVd8XrA4nJ8aHhYXkWSut6qJbECMv+nWK51pejFJ3XZYbYFcaQLzXnSlHWw2rtHM
M5q+gZSswlcC8zt/PcyhJAnpQa2gdbKdyHlVL41tF5l0WGV3BkVcO+XgDek4d5Ck6Rd2mEt9J81U
EbD7I1FHgmPeUWvhhDxyLQlQBHQQzyeOeZgAaJisLdiKWA2p4PkiaPAPHcyvpEIyTcaR09+lQkJq
ndlTDsg7TWHPYUiaP4OXWfYrQBUiiV03HJpG+nbhibSyK/yNVu4h/Mv7ckf2czhJFHNX3pfvSv7X
YPph+LIxmQmBMkvVAhMVqTS1sDkWg4KNdzZwR+zy4DfON4o4Eh3MxPfwM8VfLzzN7z4Rr9kgnfkb
C4Izy4+fNuGu3Qa5oSGPqqi2subGmSvZKDS5rUfvcbX086P7XC+6OZ6CtEJOinWVUgYuCuXOjINv
Nex8LTi0DTN2Ob6uUzjGMmmW2A+ewLR7fK18z9dYP6wwrOvDYAKYpUc1bxPpFmOR3+wUJmb7UPDY
xw8+I9c+6+oL0IvpIcb7/EWkqPEUv8PtsK5l7srcD8nkNYKLdYDABtH7KGVZiQNTwHqEz/24EXnJ
NxkjiT2OtPJWVeYRW/DVxQ6Y0aeytDsIMJcvzQlEfp22m8sbl+dL9wOlPCkcLpMcqwPbjtvvR+Cu
4OqiguQ2k+/FlzRCet6Bqy/MlEJGxhOq9lViMTm+5V3F6vX+dcf7zi6bTHG9YVEAJLHmIedILFzA
wfmnJk3jcdr3QKB1LbIb//dMO0hnrJWwcpZ7Seny/uRad2Ctw7rcZuMukccMxjHWotOTKFbydO1H
W4f3k74ds3UtI/90CF/IbCVXGkOrlPIeydVmVf73E0oLoVUMg2k6MVuFUpMySwjcwDFiRDqSN//d
6zO43DgiHNWxkYJmihxdKD/BW4qdxFOL7SDn+o2iT6jhCc0R8N4hNEHjfQepZAUpCq1McxOMYZBE
cX5IfO3AcmjIkBCF4C20H4uye35HFf/zqL6mN2noJwTNU9ri6h8J6B2RoVGOi+3Qjl6a9oTooLXd
mHRrD/TyJ+ouz7hLqKzHF4rBU4XmrSWvltaq4W7DDDFRrVvsq02NT32d8NX//+F1oKy6qWHUyyjt
XN5/OPxTh9tcBHpz4MoBnEzbqPJMpuyHz6BRRkkMhHAycQVhbct3+bckdF0MGgsGQW8tQ0tKLjYP
v6n/HIrxFd74m6vxd0QaSMYQAPxs9RjGHfEo24ZdE/1kkDFIqFp6UcEuz2hPdl2xH1fA0RLw0iV3
KkhyoqQuQfQXZioHEqYzk8tmpISBJjwpROB4psYpWat0og/vCcLvj0I03MhksXCfQMGrVziOOBe6
VhnpEY3Qp+9R59aLFiuPiSE6zF/bApkeZXcCi594nc7I4uzk/bpYWkzTD95wxCuHX2T6Y3Ygd+Xu
YVu32y4LI1kvze5f3Ke8IdMKYhbtUGxCQqNOnW+YoWRsDzhQgC5k1wmwnHmN2wviR33ITy5dAyUv
PfPzQCIlXXNjbNaUdtS7bOdRbB/qGxkjZ5cBM34fMkaOcajGiQBtm6IAod+JCkamNpybyKJRjeNo
zcU8/NfUZBb/ZMQHTy8PY+SFIKAi5VooZAzkzuzQBx2xMcz1m3w8ILaE6R8B3d1zkFCoGW3z5ud3
BurLQES2YYz1pFfhj98uy6G/FOd/dJhs9Un5JFuQN7diH6glK28YycVNkOlsId+Kop8n7DMop5mY
BrCnJvP42PIVyfwy2IatAZUKxx7jgfCr2VP+I7iiiSH5MTVV8JvDpv1hj+QpaUsTeNZa3zgLlsZi
OReNVu97scG6/s7IqfQb+u9Dsijgna0867shAY+gRreNmtSJGlMfCW1UWq95ypcSv5k7hTR8Vr8s
R/Tp0VWkzT2dGOUpNnnOq1Zj92BAq/cZ2yd5t8bsJZuhi6E1prcx/ikmSMRJ245skf7iJCs99BsM
m9Hkde8EE3jbQud8jr1SVSfBTYb16/YuirSYp0i+O6fFCro2EKdhKWWm/HPM6x5JEF5kCEk3Tzx9
qdPBiribsd/pUyHoLNsvBtgGIidMB9sf8aIB3aBTepPpg3gHgXhIWRBYnjZ3KljI3vqRp0R6XVIJ
9+oMR5IXpXUj5L8rl0nwvZ4GhXXnmvKn7gqoJkZHlige6oSmFjvQdBAJ7e2PaE/sw3xrGWOT+myW
9u8yO4XcY82JGbMkmkKzFAMs6MvwVavcB3va86QgQ/g1n5A4rvp8ze6mZiU6P8jdG0faBCg1Lcth
nLYZTDuI6W+01mxB/e8FLfQwFd2Su45z274ylE71qvFXkxOc7YAMrS+e1Ce1VmRZGGXnb2ISKcw/
F9oXH7IIAH5kc13iIwgPTWB3KiyqkvnbzCLCDQCqdqmXoTA2+lGIKKPiVSjLBYves1yhYVxufNLB
VCGpNy/jACC16gyKyXpL6jfc20nSRVE4ltQVNq8jlB0U9kxralOFFU/xp5vQgPbjA0vEH97ZRA3R
FNUTEpo+FgiuHFyWlm7ivK5pbP4R1XBQTe33IXkGlhgfBvyAEn51YL3Fz6C64CVX1X+dnNAOC3rv
pIJK1N4yaKqWqQ2bKv7G91SXAOoUWq/j3M5/UWo7Zf7G9I3Mu9AfplFzQzgaHe92eeI0FOmQ6vTQ
KdLYM6ff0KcY2PhHtrBu8bKFOtL0E9tgU410sL6WhyWvYd239++nOhn0OtvDSNMaq17QLIdPKtkR
k5beHGfKiZVTerfSRKHbGwSfn7cLDbs26P5PLwLGaq/3rfuMePe6WAR9JjAHzvvN+dqP9Mw1O5hg
8Zjh/jnVljjNvL4K5R4ZWKA8ifeMPNvhS92VY66clyRapY1mZCjUl5fb0Z7i2cEKltszv1M24S/Q
xhbuA+wJvIORvpw+s0ebaJm3tHXghDEn6vaPjHC0vFIswPokViJlFYm76KTsSBb9ylMgipr8rv5v
6jehRUWZdSJf5H5FuCdisWBwjh1pMvzsL2fN8k173OeTlQUoa+wdXch3NRFsqp/8e9YeU3mXi18k
+tWb6vX7vZJMAu5b/aG/2yQ8XCunOifzm+i+TAwdUc0ufarbLJmEKiqOEwYX/jJpWbUyzk5KAL0f
1AUucJuE7hwqWQ7lD9KHOx90WGtGM6LORQXM7txrcMOpxwB8PpsqiyHjWA6cYDlHgyU36sGZsCqS
5YO7WbpdVvZ8AV3U6Dmvj+WbmVpIQlRn/PUyscxYQX4/boTEX7ao47EKRCbCJFIb6L9i+fHJKNMg
lwe6jzIl1GAtLoJ0xD4BTwNvrQ7uJzkTa6E+gbmFPsOt8BXSAcS9TVrtDaNkPnUIC1A5cUCkGFBP
JvKzRrQhOF8OkASg5PDgfe1T4bW4gzqrrHr5tVVpDCnYmw+Dl6VKONXgokXD/pgMu4M0Bj6vcftA
Qx89vlyjInmLj56aMJfwnlcQVxUrH2zYVAYtWtJch0XYPGfnIsqLcN2/4yne/LhVPWB5JiZxgJIU
gnos4e6T5CT2w7RyiYZC5iYRRmJqX6P1a3/dqCzza/Lssd9xxmxYCJIgwQmuhn1P5blwzBSaBhpv
NkqhO8ypRaIHB6D8gWo4xlszn0OOBHy3TnKEhDqF1jOW7mpSGbHYjFJ1Zl6sembgPZhc75W+bnqY
pNNap5wuvyRwdhFg0kHv1IJxlHZTyfsnSrbKd++OnJp9Z13LShBsVElvs//ALqwNJ3oLZLJ9xMTP
CXJjA7vDyN5feppY1ZXfIppI4KhqUTLqIQoj7Z/RhFdIPXdbFRtSLUOdUE0sEf2oRfg3WUMzu8h1
hluIFkARIDbYbJmH0+14y6n+IPvPveyIgZo2buV13n+4Ezm1SNf13Qa2WFAyNWdb2ERrcdBY4N/U
VFgp6kxlO1YEs+2hyACOtHwhaMp9nt8JjwRdJ7mHSl5Yld3SpywHq67ary/Rucn5+LQD+arpGjZ4
s62QSylKPnP51A0C8Jd/XIWCB69jy0kXiurVFkpU+EkOiSBvp78yhpKGPwoW3LRCr3erqAHrb4GE
OSugyTgPaQMyu/1pwRtg51s1AIpgWNXMK+UUS3tXoYfdUMRLAdqGzzy0Dc0diEZ+53VNF6zik/k5
xcnLU+qIbJ9C/8N6Vtgh8HdQDaczucWsCLA23PMbAYLhreDR/3YFWsmS2dYIfb7F1XvRPtbHM08D
G0GtoJ/d1mggeuzCNZtA8qimfDmxd/skFZaKkmP6+cGJUPVMJJbfdFj1R1YUcrlJRCSxQWyLyGNv
2YW/N/dI3SCXGDrOHFfSEAPn9BjRAyY8Y+zKC+hsfC2EA3Qof7KKcQwQJCJROzYdDbugxdH0vS1Z
HcVLdapRtioT19sExHQD63QqzzRDwg9CzB/9aEHvCybKEP7MedH0LZYE/4pj9dSONcdaEwuniU5j
Hgk4DG34S4v7mn/jNfXZHeGoL+xfVZBPvwQp3CoHW+lHZYGeG9WNw5aUz+k9OLHcOGOx7ltHa3dO
jexIzwmTJp88U2BlNNmjcKC5XDvzuLkuPHxb6jkPcE6PxJqtShYaGdIvgSA3MMdU94Lj+vH5B7Fe
NI34t3ZIv+IPLptDDPLlMcbcSZPYKwqMuem+estcRzkUytrq1uya3kqlZlZN5SBS1HRk6dPohs6Z
U9vjIRhBTKLM9lTP/PfgoYrgwmsE0GCOuZsLUlGFC3UNP3TOQPdrgdvjvducT+xHy0NzbnwJsUCr
WVQPFI0KlEygpA8HfpBKbVWmJ5SRXW12pbSalKaCEoM5DsEoJjdcOrdADfIDz0zKvLjW7AA3ptCC
Z/nyzGgzgepO7ZaNRcX7T2cZZFQFW4dXXphrquHL91uNFrJPXTm0KYNX/a2z5cx84wDAYgwtmVA1
ktfgJwIIBfLK+c0UOkxRhuf+PxGT6TwmHJSvKEXMdv3CN6wueSpmoJfCTEMXuIdhLB+NM8YNqs3k
AWkzByn5vtb8V5kT1wr4An/s52S/Pb4emtBwv6UuQ8BVGPdbUHqeXXY1cA8D2ouINvUjz/VUx5wT
8EBSEIREoz2dxnB2rliGBDC716Hz9qb0iVwA3NOxAgCNIggTZ0DhjlCNlzyLS5ay5pVYHzJ347d5
9B/0IbLngE1OWlYjAUOHIuDNTGrzOJkDlTE20+zcBwBQGW5o04C3GHuS2O2F14v3yBK1aSRvFXFy
zWqd9ckjt1l1V9r1BaAX7LSJDs2Aoqx9O/NrS82Kn8cSB8eyloEIEhBmnS4DRqR+GnkK7g0vCPe/
phfYgA3mqqrvBfXzSrsY3Jywl+ZYlgVfwL4btXE2VKq2IVS6fj1s+8vAFzVEFzS6kb7N7J//4FM7
+3Tso4ClERqcckGDRTnqMdotPrrbR1teNkMTy+AugZxd5JR6cXBB2qpJIlIzGr27T5znBVufWiHO
zp3CKNQgcCcfH6kQ8Tf7Un6zt6nu2eEfe96XXXUumf2OhwUXaCpA5+EnGaSEZhFggIJfDRIYUnBC
Wz+deOlUMm420fx7BJOBIvYxf9X0pEfuF31IdyPoG0bSC3SWLybFktZC/gU6vtM7Aw7/TlOfcEzF
cnUMDAoECnllroHBNBMVBxSLVUHzL9ehh0Z5FbriYhPXQ3Fwg/+raPo9BCegZqnfnbVE9KLDFVMx
vxFG7KX0BY8Ywlq2PHbyDwfdXDg7mABzGVm5MbQsD8Uebs6XGx6+A8H8QgQeK/3cgS6oIw5Rp5wh
YQaJxQicQ5J8XttRH1foYS8SkbHAvPpXe4P4FT4DaUf0xKKuka9uLFoisRM+2RaRYWKebLAii3UI
us2dpKLXQWfGktaG4+YxmK7JTwYeFBZy8zKOKhK1tpOAI7VR7OKyiMUijHhz51oxZIXljFa7C4Hy
67NMKUM32/sIatW7nK3Wl4SBCDbdrTdiDJQG8z6HgXr2w+EjqOf2v4f0+l6HIxy/IAugtR5PRU6T
s4OJPQ8Kgn7SM4Tiy/F/bkOojjH83tZOFfqo5xQoUFxF6wnA0x36ntlCHGAIgL2w0MqaWXlfVMqm
c2ucKxRVqiXd04Su/do8DGVMXlQexpDFRfoVNCxa4SA8vjEy8dZvwXFvUbbmDEcQJcxRIwSlavb9
peeSw08nQ0lboVk8bLWJ6sDfyndZHE0ryBsPk5WxXgDHoaHgKR7DsdNmsGLHgcQsfvOh4BNRnQYC
JZQIheJCAxqZZFQlu6ahhVkRewKc6e8rTuv5mfmNHd7Qk7h9Y1Vn0tasoNSHs87rUri9iZ1ZMQdK
e9e7C4jPu6lCNNkko/si3e59jg9lYDJ9BbCl4UBU80n1d/f1qHTH9ACDwc6va6MmEOx4SXQVmoip
pemE+iFrhCQapq0DAxkVwc08sUFgVj/HQj5Qeg5voOSLYjo6KhxIHTM5fiV5XJV9ek0lnvNvWlTF
tVYDWat3PiibbN668wBFarXBXjB7r89Rw1VK3frUpPZO7Tg0bkmuHAnS2TKSfxMauMMbA1ALkVfG
f7bU1OdiRo8jSLat2os1gt1fDyyKHAuhA3S9aSNz3YvJZYGyQRNoJiXVrCr87DwdBTeH5TaBqdNs
cXi0cVWFMdt6pRdjuQJctKn8DYMSwRTHKfSdR/11v9k8rWYRwbsQQMyXWmiDeZoDOm3qSkLba4x+
8JQQNGkVzTbZpqtIZ2vDc8t1fGtJS+CLeoVJP9Xuv/vELEaqVO4k54iHYbYTudxh046g+E70cBmH
yGobiMHIaVKtHgA/Ecs4TFj7KsAoSqWzal6D7PuRs+d75FxaJB0JEUjGiY5/PVhPe3Bf6I9nkif8
vg5AZWv0TCFx673nK9oV6M9Eg2p0viWZMvSy5hP5e/ErNtrAT4ZGx1Lc8KsN7KRZU9yBs3pTXTyy
vforr8lM7ELwiPY6iAayjY7mi+W8a1m+4RnTPs3c30mhoMqlDvyaFewpmSK2Zn2vo1xJDQ1vE8TD
y5+F3Jc7UFalTqpQFjS/O28B8OgzzSui0MG8pbQuMK++LduTELNpTOsULqEcl71pMPFA/Xsm083t
aUs7tjiIMBK3Tr4oALKUEcT6tVeo9nabIN/4QYJ9qdy7u//x6a5pX9FCO6sez0xPr9YFeT9fFcwd
ZzWtbC8xgcp/XTFVUd1WHRfq9wOpQj514HQwuDKrxKvWWj84yubuVkyMiucUAsCo0aNzSr4uGFTB
WN7bnNLmP/DZ3KVyuZ93TJkFtuUbzrXMRdYR3xC9zqBl5hUJ8DauoGeq3zk4BEehufH1OUMlDUYe
lTetSq3h42h0vUR8okCCr2wwqVOXb1sTLZEU6KdX0nMKgSGkFa7EAXIhlSizfK9yeH/SfpLk3+R1
yojzrVqUPTo/7XhuxN6nOf1kRq8OE97ELol1cv4ABm0JbmsGwoP1lmP14sbHyh16/NdCt3UVMhjW
cpvq5YAWO4R08PzFV9NNn78C6eLiD5EBGJm/m7LXgWluCznOBCHSUvhOANIGsBz6mC4QDN/3qtxY
Rllg1WcETFHjxSsbnS9on1dld694vnTNe93NmP3WImQAWSp5ez9QK4Gku/JCLOjLOEKzCmjFFjl9
cKZj0C1WdayEgpQuGUdD+2glkIUYIAeBNdpsmBU5GRFpr060uKaNJyh/6VuoqRuCEjdD5MaieiEs
P5l8Kd8GVzb17AC9x2D91y5F6dHflb6x2ILAQXoVMT3hLf2nS/E6/BhemBPbswcF87cqjIKsOnkN
bxK47lgfh/wPJ4gEymEdBO3fpCKhCduVdPx5KHLZFOUiniHpuG6rWkewJSwycm4dluG3i8WPOPbF
BrZkuhSQZEpyxfEkCIIy9Ma+89T3bDrS1v1qDFx450QBKw/eR32ZdPmpGK1uJAzQnOOIwiYf2vDS
wL+ofU9QpPM7r2aj9Wd0NcZhY/Evrnum4doAEPLEV7CKfQindQPNxHFrkt0VAAnRO0qpoU8JuV+/
T2DVc8HoBBZmnjeYVjf/j66IBUQCj2ZKUkbPpJhBKU2Lz+utzx+fsYShNCYLwMOZV4zxOPlhOByZ
UQaG2hsmsOmzqF9HCuQVJW/XKOi3BEI0L16S0VbGA0viZ267jTRa7qLMhusSPLrZfW+6x4Olz0nS
d7Baw+Ki9zlqUgDcBOcyeOz48PQmr+uNLMZBDfuyArgia/Y6nrK0jKL/Aujz5sRg6JyqExWJGHIm
6rF8+/9INMsRHdNniaT5d4AYmQT+l5wfS2FSLLGsZwMkAPewRqhV83uh0mIC+/lOaXGqrAAkTqjN
1MvEjmVkWzRQ6ABBtZiF3X2kT+b5eK/Aa2IN4rd8Tpis5MtUgtcd6U0VKVwSQhdzU+8DgQNlor88
7mkpmR9kSfdgR5dzX3h6DdEA6rhWVqHiEVNd2UtJck1dDU982TtDKL3dPZBiZDPzknss+FsoG25W
5O0/DFijCE5WK1h31pzGX6yloxsoOAVDANjDkPL5SEhwc4XsSj197uVWIjjSUS0s3xhGQLcmTf3F
kxy4Hzdfv5sb1vDRPd/kH8m+x/fQmJVQxb7DUskCEmir72FvbLLwG0Jn+2jsZSAI5kH8Z+jIiXPf
Mg6Cy75HCRA/VNnA/3ub09wTh2no7kH7l7BXifhDL5dJrDrp85pbZIwcU6wyO8xIl7MCA70bW+PK
Ow75OP96dnWWRlJ/UAwFkz+cJJ6jDxsNt1Pz2faf78jn1sRy+64A1E3wasKOZOUAKyhEntt2Sr7e
diEasjDwGwkdwG4ZFt1yQ6iGBjY6W6CkeL9hBGPkuKYkCDwlFxMDz+eWQczJX/W1ulb0OOOtKUuL
KYTYaQfFmHf72L568r3tskBWcYLUpJM7dP10JewKZHY0PyPpMxVmVZBVghe1ZXwMBQ9tbBaRj66f
pBaaYgsCNfrDCjBkvzBy1dKLeV5LwPvM0ooHAGlXq0IhG11fOW0WSpFVenwymN9uKNpG9UZpGgQX
Ip/khnZ2pLAtR6I9fPiuSoiw/r0KilRPAyc7CHzvpinzcHqP3ge5fccClxN80OtpJUif8evpKDQM
GUZ08ngHQXkPjEzkzxqBtNdQoZ+acP7hr/6cJ6i8vc7r/pKHE26cNzgkxft1oc47pAKzdiou+AyU
nmGvmpFTvT0S07ip26IQqEAr56KDV63IXv1djrwxDnNMQZUF9Q23iGmpEgaQx/piMJoLdWu/a9XT
DMlVoeS0XjLrmnxC4IL3w0mdC0KMdNe8G4ViLobP6oOMzLyFUFee4kNN77jVpCJINQSRJiVlaO1L
qNLV9ylZ+g6l6fdpfe1gHx3suXHjoZ6AVl/GneOhnxRGJ39tDefQZ4M8tCLtl/d7Il89q/5x9RKl
bO4q9y5vCNqQoXHVjmMj60wrzZoDXl8qItRQeEZDmuqR0owQDxm3sZ8cVOWTHuPRemf30RWuXDDE
zt6RcvhLegDr/gczyiNZBM70xOd3fB0Zsv1+N0eDRTuWOGwdkpGmEPD4Fq5vcq7R7NBL5NtGgIbT
FIdzJsR2Jtx72NmU4LO6rKe1srX5hl3Z3h6QL+ZfAERVMIgaXkuKy6ACGid4lPqqL0hWE6bnm3Ec
ugJBqtdJSU7uHZIv4BXsic9pF3blFpk6OHEefGoevr6XMYRRC9q2HMyFFyT9EFd7Av2k1Wtn9MDH
vhI0l1c5VeLhdbq8YZvq5o4jHXpWL5NOw+EUG0KBIg2gZW3D6X5tYZMs2YUw/ohPFtz65q4ldHXj
/eYK+lsBmwPjNK9P8Oiyus5CE95IV7SgjFU46rfc72wnLHZHLRTqw8Np0JF9lN1n3wJjMpoGj3+I
mVE/Xn16NkeE+Vlra3+kSTxKfDxxcbNLrnKRduKY0qkU61vIuHCOXp2gdzJ1/c3CNGU/hq/yq8aM
WuJntlWLqHE+FcdShGA4N0FT6s157knujMofiV3Cw3wSqMr/bqwA00Kd+9hRWZiR3fCfj5iM/QJT
DuXX0oUrHwBDyWFuqeAnvs989TlggDyjZWKedFuD+7soBgVivGw+hpCUfL8fkWETg1P1XmYxc8ta
FHhrlq6yUYzQJaYqfB4rZNpbf/pBFdnFMMdtjR4i04U9g5/J9IxlDfwM/tlF5hY1hK+x8YAso6y1
xBhqshzRedN1nYBNbG8SzqsE0aA2bSCS2X0BqvFs7bwq4O9vW/ln28Tqfl145XPqq1wCXKmKP9h6
0swsu94odX4hKkNCJJisJY8/k50fTsypnghajrRXTnxBZnr733P5McGKGDJmrtsOVFeS7552ivV/
V/cd6643Lhvmny/DWlBayKFBo/vPpanpGXTFh06ENAY5/j5+vfggNxUgtTuv8WuxVGR18W9LaS+/
KJb3kXKtups1DTv9acrabVeY8hAxjYMJma+UQ0sDnAMij/+C2mwXVx2GDogObBjrnTZWPqxk1RKm
Rq+ubg8WCCvdVNHLOD0XF0MWjvjffVp5XcikvGIE5w6UgJZA2YdkeZuFdkQrpCO3+4G9xtfofvjp
jJhbg8WehehNVCpTcy3Ux1+7KKyS6T42nORj6v0kBw40RAXPtlTVh+9b0Pfvp4yJ3OC4v4hEM5Js
L0eOcsSoIX9io9z099QYg3BgYGDeXi1OiIuNJGO+olaAmVR9f4RP9Kngy1E5Ymv8/ss/p/pz8Ogs
+UKnefGnz2/LO9+ha/T+gISqNWipcU+qIsx0Kcq6rjCHp7ufEdribbArC4wkuwrFA+2/M+g6f41u
MgF7VusdQ2Je7rz57gLw/f5RsILPxIKpxOesCnDywDpZBKYf5HR7MrLS3pYHcwBpX8dntlCozcHL
yL/yBjJLm8llWAj6+dQAg5hJh5Ga6AscioJ7j5mv0vEsx5E7Zek70oIhzZgHufTl4U8yn/R/WKRB
1A45jmt12GJKdpYtiRCDaqc9L2dbaIQ+DrK6yvDIgiBf7Di5EOb/QwqIVnHNToHKnQiR2NwoPb7r
YQzShy4AR0q8Hw+Pgfl1SSutDsdtssICivlsAnLTb7YecYzeq8bi2J9nVTGw6eK791MSvlpiAD3q
DcDm4+jgoJ+3nVBGzefcLq0M1XQV7zq84Zh15gfqv3Jd9FO0pICmlELvlg+MVdm4BMR0JY/dkltp
5S3VEdqpKu0Xr/HDRJJYjLE87wyofhSspeeBEyKAk5J13hlwu+3WJKpPE9Dl4qLVnvSKvydS3u5C
YYRwmlQ+EnoelCVA80He9C28vYhaWTrBf+ZU9dZHM+jm5+WBnkvLtNCuuTnwhUgB3p/Z/Arxir1G
1fdcsyk7k2T8V7HT9tmCs80PxoOn9ctZx1rsqnOG/H0g2Xdy0ho7Nm7iZ4Fh3xy/7V8AJW64+URu
rHQ4aaC9IsJBEfatTf4dcLh/bCv7TG7HJusYhVFUIpiY3wY1geY0UZuuGt03XEXJ/zgmzdTIDyRq
D6lyrwtppdIRFR6DyLcOYkpDBZkMp3tFfyagDFqz+1GKvs6/4ksxZIi4SEiX6LMccqy3BVyNIe7K
/r7Ia0HJBzfx0gFH4R0w9GD3cSUww1aKi8l3060urGnjN1GCJZCO/nJdQ2nY2b11Woz449wy68GV
YUmn0UesX7L9EYq9DnIkLbmdtEFra49acmXS9shLEScOEjGxkozv4QrUW1uDj9Kb+t/5kMRzqdN2
qppfF+7KxVmocSsYYj1Dg28R3rOUJ+MHe9L2CivukSkgsLk3sQMjHHS8sPZY7Ekdjlr/nxz2gu8c
0QBkuOVH+K7FiB22e1BlB6vAWCNGVJ/ESjI38qv9XCwNlpXlJSnAgTOzW4VOC54Egy8RvZQFrumx
UUFLc7MxNLqMAVncOMO6hGXWAd86eiJgx5wHSb5UXXdGjBlAVvuX5lTqa1JcxJkmn/t4pMT39QW3
RGlXthN2CqMWcniYKV3JQ6+/UsSmXsycab5XtjuXlEZ3ksUcUqgpG7hYv0Fjp3tj7B/2BXvi4R0k
pZQzLNn4WYR3pZ9kjlOTKVBEZHTyxAH78FpDU9yjOLK83Tb5gMVAJkSf+xCUr4brkRCkyebFCygR
SBqW2n1rlt4/NhP++W8OWYs2IrDWg733b2w/HnngxsFNzAXpuEjOE8tiWI/VQ8Kc6Tzn/E4evLnh
VBKUxD58+gAF5tKWWJzWRo+jtuNm9ToWwV+q00otlFZ2yVopSBiTrLbgOzsYkkcpvdypFm79myX4
g8ObKAhbO22SmVHrK1WC3cRP/7dyxLiYbmpxz/+VdLRfIosFl2mZbkf1Apsgk+iCJJCPS3HIfeVr
Unrdy4PUsC9Uh/3Lpnozm8N7Bs/0CeG+GYiRE2epTQZ613nJ6OfL9aGzls7ATpoiqmckOCPAL1QW
q4ANfkseg4B/+YN1RIFPLFBrmE4tBhbXVmW9xPqyLXRIyZFs8KIigZUSvcRRZxsjS66IgJypR3vq
0WbGnC2Zzus0XiS6Pb7qidh4n5ZFaiNqxiRy8OOooIcXdspOzRDAQgfVevJMB50LRQ3avhdl4BfU
nPPUdsgYy6Ae8hyWO+m11rS6lfvoRjyk9h1HFb0bRRl3gHCu7ZJnHkjlHqp6vkw7EPr8eXnE27ND
hvgfzmrXTdsm/cxKsCwRe1QlKkqpXEFXiHh2f3twvTxU0o5Ol3DwGMcXl0WBXCuLfCkuIRM2TpHk
VLct3/q3/MivimwLtdHFwJzufPmNzPYUs7iYuiJpb04rKBwzd4PwGWD+Zc35JTKZE25jHi0KqRJl
TIA1m/YKs3YX0aUKEK8PDmm87B6qSUpdDXRdB8EkB2Srva5/5apVJRYFxm6ZqP4Qej9t1HydSP4O
FmLSqkZLNQc9QgzCCFS92IJ4kaY++Se7DtXTE5CQhdTC2h3iBmUmN+vjFOTBWPGk/Q9ztE+dii+r
JCWsU2KHYG3+e+rdy9wCsksw1CFsBPq394heM2fdBlWvWopb497cXt/nsPQRM55hpjJETrivNMI4
tBop9O1arC0DdXD1sF4+0QzyoK0GZUxXITcGBSDwcbsfSIJp6EqJtE5BGH4SOoCdI2ZCJNwA3fMi
VkokNg/YiMjtPcEb6fk55FgEs6KTfLi7zxZKX/8JQkXP7Kae8wpfY0LEG/mF1gbABtHubgu9bQrK
lnuYggOnCXdvJq3LAEV3WZFdB4LMxRXeoN6p34xtvWDzyb/R2y5+pG8wL3cXbNb+hXp2hJ6ohvDv
XLoFQQRPNdqHPqM26GMT6Krblgh1/KlOU1lMm5AILrqtwhwXcjqh19maVtR3itseXK9UGgC8AGa1
1g7H4r1SzF4gnD+QN7NAwYNKZZm7fdwkHSehI6NxjbeJTp6rJP/ERToBTzjJcg2UDTm1Dh134wcI
79qbnxhYFYKnEUuCUrEPcgBhJAe7dNTgAXX9rwhFRw8oWJv5AzwVX4ODnN3Gqd9Sh7XWNHNH1VOS
QBCksAOkG0n4HVqgoCMpnpl/xDp3gakuUEghYNZD4/O5qQCzWyq3e+hegiRZiv0r5MGbVr7hiVT1
NL0cTL9D1RVFWl4KMKRof2ylOJIK5mFL2U4rBwhbf2ASuARSHwv6OuwxNg2J50T3lon46GzqyOtl
ZXfvRGkyLA8ENoW2Ql5gvt2yxKJYo5tBTInQ7ZGabNFiu/N9MzasnQA4GwyRCSrPqJzTKAqivVVH
8i0D/Ly1hInj/evS9InvHI/PxPmPMAd1tJ24cIuDkZ1RIeQvklFnvP65lXTB8zyAZPpAd5GvMe6R
jkJDrrIZILHIQL95r4m1QFb4mCAHQwcyJKUdcxG/JFqM/FRLyXYl1WYz0JVS2kcJ+meebLRTFeTe
s7f9PV5KAGzzlfszXZg624zsVrTG4Yeb3muk4d0uu86Q+56BhMJ9Y8CFanNQk7zes0fFbaiXhMAL
h8BhjuWLB7nq01HJmEHxdci535/lRqgQ6SZ2E0LMtlr5rSv3IYW5+fAvG/7xg0IuwJmclAMFGTGq
QgN0+VGc6opwBH61T1YIcMUerVgpbE0gpFIN/lpWp0bgrt40EkmqvP5hDrmueIojhK9psh4j9STQ
FGwJnMYZPaFYbOt/cp+OEwQlCF3TVPETlC6NKgoj+xwFhQqfSgMzOl2PkYiOkeBeIGwzeR1mIxnr
DWCeMgRdPsbIIYQZPuA1GvF/gzguDyVROfERXhfEEoYqn7HIZKGONzShph7bFWXAoU+xwdUuJggV
R9I8lT0K4S2W/b83mggtLiz6NVBxLzYZ51URWqoHF36UGjbrZUYcx5gFVtyqtD/w/49658W+CsK2
7YNLYQJ2w1CHBoYVHtvmqtJb01JrLSwsyPgdRxBna3+t/K926KumMmKyhPPZbxsdoroScyhuoU98
Z3wI4tKod4slICSSVMGJm3anMMfVoElXIYJ3K5X7xWz1Tf21lMrhVf4acrrq0SZgiKrPdSjd3fwC
r0js6prSa6JvaQT6mVdGALociZ5otsJfZ9pLmvcZbEXKdSiaCcMq8hkrt+0Dg6Qdo0G0FkHfMdU/
Vb9m4ZuJzdCYZKl+DccnyIkbe8gPBo4i364BhGs4z4b7R3yswjf2UPejoxSB8Zz5tKVGo8ZFMChJ
KargkSzCLMXlIXWUQNjoRTAUj7SndAIeDvzK8JMLhT/fbCEUSsbq5p4mM6dFgmFA4k2lk5otFGQX
0DVYqmpRKGi4qiziNILHdX4rdgSR32PnmeWOOkYPP8IWny7RBGRM0gn1Rq+8aulIOptJyObtQU//
B8Np1x4DTLb68yFxQQMvi3SnxH4dZQujv99+YKVHSdVwonTKF9XAG29NRsu5s0nllWf3ZyzatV3+
hQHTfDDSaX4KFm2QG68v/eIl93vmCMf9pyx3Xvyi2Dj2aZxy88nLsjzYcLb9ulaZChfZhQjY6w5e
fcAbqs5PYVfwIfJJee2ITboVZ6RppNi3+dxW5r8LPs0Lxmuv4agF4fNa2Vf5sKtlxWro6n8iVX5M
RlZ9m5Un8kRSRITOya1p8mKi3fOU50PAhJ74leXnihm8rfC8BZJhgKkJ9BdcU2xiwHBgWfHRC1b4
fFinuIPK7pjzx9T+m56WOAFfgBkH0qJmukQs/FBqzrIxBWzLCoBM5Z16DNq//cGF43GqcKv/CWGw
9Jl3eUxQod2sUzPIG6dlSEbv0VW7ARArM6auVl/uhhLQ1+PkheBAOzINwRQJ22sarFnFdCsLObR/
XAnAegFPv4FcZv7ZRK0BV0vBHm7BMaNnnb6wv5cov9xXvxr0cmjpFFxdSD4vhdl2AIoEdDSLqA5u
htXtFDs1whgiWqvXDMEwax75qzuOaGAND5xr7n+c8rdofCQZY8AV/U0wWjo8lIuTSSouSdaPbCjI
7hTU/UnaR4dzK5GwYmR0s18yWyHcy7pJ4rmeAGaAzjSY2yej6sE2Rx7OZ7GVMEGeniTS571We2Mg
OtaQ0kHykUSER560XEGOFCW7KHGPedgQYuPKh/8u3j6T7jIYiDCiI0OG8inWCfRbv7ecK2sVb7+R
Kl6vjphjJMG5u9nukl9tbfyoqEngM67FsXi3oZe/QWk+bw6jDp6nSp8PZESTXstTES1il7ckvIsD
1NjzmHNrDF1lHF8E1a8Vr3YmmeJkyO6ENDdzgaalZzTSeuh6F/PtR5ipXZ/23Y19/vfFkWzm87zR
Pdqhu39REXvJ4hSPWUuIKZHkhqc7w4IiM4NGa/fgKwCIH+ImYJuYMUAQ454S0A+56wTeoTHI/QJH
S1R0GcRkCO6hNIwr9DhJFu20RaaU2eN1bEt2tl1xOk0dOXMm3HoMxZCq0q11J4S+EIUNiys579a0
vN6Eu48G3zPHUJrfvrWzxA3jb0tB8sjRUk6X/8UUYmHwCuucnWkbsBU1FShfNI95Yie8s0iwHNVd
QeWAOiB9mbrrUi5k8QCg155Uww3WcgC6ht0bTbYIw8Btls/HpzENeow9nAqz7rc45LIGBdHUh/Ub
pG7InCTd6xqB1dECgSEYrbBpElVXtiWWKDWVg2RwG6KVnfHJf8NFfBD6ZYcEudt0G9SeVIMwIZka
TmtaO8DCDCuIcKD1slgVFqOSY3nT3NJ2vn6A2USaMW+SLBx1IHM8Z2rv6b4Aq4FxGApjyvka46UG
+DetcMBHVmNDN23qXToWCYA1ndpkkYPnFPVM8IAPqfedGx5v8vGg0rmUuyIrqnIRzXrjy6/7tGJX
4U/TQQy4SqWStgZ6vkmJiBOLwZvzZ0cprPMTMGilTThjZO3D6YGFMA/DlWmeMX9T4uAlftNqAsMs
kn95AAss0yw8CZVNFR0KV9FVWQtPwH5rv4XEJMprdqd2E9dv3aDwTQ0lhgfmJUaa5f8Sj8CQK/DE
L8eFhQGxKHxaKgl6jf7DvUrjMHc+BYrplSyb88q6ljLReIB91p+wZYCx787THf3Lg+sugM0mUNry
n0iKTJWdWKKngWeqirNeCqcmSXNsLDoZXNxVHLIPEnTX/41k/vzekalQwo4mkjtpjq97jn4/6aKE
D1hKWsyNXaA6KTYSxXrFZiqAFfj4n7t7y3qZ1plXc/jL16avsmTUvYI3KQZjv4t6ganJHFx25EaY
ifyfyWZP5SC6QyWuRm3jxJ2PNpULVr5aQwT4b1hN9scoX9jkyXLtA/uqFtfj0l8JZgEz93NMniOW
dL89iVFvzDAZrVqY7T8/ss3A32T0I+VdpNHSDqTP8T2UFjUxGyUJZ4zfhIoeqT8qK8ZqERKKUILp
cVdDY7IbwEXUwGfsq5NC4MIPnVHdablGGVkf7v2vYUSf+vS5j5Vl8prnEzV+ePt5XT6RZ5Z8gexw
GDGs/lhTrqXoEFr9w1o5NW1II0xKbMO3a+INrDRk1q9ya0E+gGYNgPwxkwhGVRdgpm7GaNangSIG
DECIwiW/Qm4Zl5InuvJaBsrE0l8chH8bhkRQiCuuUXXqj7el7WuSr+sW4zJeOsmj21W2uKDEc0Vf
pBZQsTsaAC8EozMQBxS+/QFkaAt51dOIHu5IrzcvCnL4WCazf+CTePEaadOWc7MBCWpyxDvpdDte
EQ88KRsq+NMCs3pigkC/zK7Z/jBP2lhhOCCQA05wMzSU//DlPl3bE5ew+QRPkYj51SNazv5o/ykK
PsxJsfDyHoe1X1Tpb1hH1xwk9Dh3sVGlUB4NzSm181aGrObCmz22B3EZSu0hI6YRADBUgTUmDsga
v+lA/3viIxM1heerBn5sRFM7b6n56c8kLbzaJIHlNW4WYuPg/IubdRLZCNQ8sJYXoqglTZfltWNQ
JRBt8E9SRRRGaZOJIlYgAuAtFrk7tgrrXz0phi+QfrUGyz67rFiCC0RReHCVDqscaMuGgUrdeUnl
Wjbp+CSTwc+CLpgcxFj/kFPUTLlhf8fFgOZkxiVxa7zSrUU1q+x5Iaja4FNuQW0KnPoNP7F/fb/k
wVPqaMEXWofoH1mnswtZYzljUqHUjv/nFXkwZyuW49JVe0yaozDLytg0nCw0o3L/P8QsaMDRlcEz
r3R0A2VJTrSbuUllKQbvXX+CX7i4IE2HDapZUb9aGakW1oipIX7d5rm6tOAJR1ztnPs0ZrG3WNx5
ZhXWjmyKMMci1WzVuF1yJTgUPVEVhXfxGpCiQPRkVTgMCR5Ev8Wvd+czNxf/6UkwWg69t/TirX6a
PWGgysWiv4tP3F3s/yZAq7I0qw1M+vzULHJoV9xe3AOhJlrlQy/N9Dgi1lMmc0k/KdudQUAwCtAe
odz1q6w/JVf7LtqrvtGk6F5KmwtenQDGS2UKJqVN/l9NJ0xXrSN8llj57SxGI03DLxVljevqiESq
lOnw/yfE1/zJyZggxQYgGI/HXT0FgtZvUbl+uu3HoiC/sgxtLvZXLYx50TGWrztTEQ4GjBWdlthf
v1DzUdxtuxOjky8qQ97WF/Ed5W+fmyphb1sBvxvLOBIn3XIqnGZpqazMSReY3MAs+9GOrVAWExfp
8s/mnOdb6MdDohEz15a7oOd/5L0uzdZS6cDA9cnbXPFnjXWUwvkKyJcpkU/vT1qipc7iw/EgT43M
l4k2eFMMUlqsGVVtVNF2QgvbrSgTDltcXepd7HEvzucLsnI0cfHBuHUxpPpU6VY7D/4UMBLjySKA
3JOc1Jw8b5sy07z+wySphwRJPMTRmOSz/TYiwWi+IyvNyePh0nQ6wicR4GMNN1YJtxVrwD6CMyWX
SJAtR5U4qSzZfZjZoGBPlB3IONSyNHCYT+6hJ0jAUXigznBdGGssL23UDH2hnw2c70vTR5nx+h41
Hm02Ww8ri/6JIuWANiPoRrtBZ0smuaIrMlJucuXOgqdVFfYyfA+45coq6edvy/VVCH+k8pwojRCV
E3J+izyszlSYLxosCfchiaBzgIAMQFQygUHs1SlHpxElZjDEfMOpKTM8UAwdx/T7M1uYnNGfE60S
KlH7adyrUZbsv2O6UxhNcDWQu2nwtSYsW+V71ThJ+3v2RrSVntsNiY8opsjs9huUV46QUuFi+oll
K9Z/UP1L2qnwQRrkaMQ4AIQHUa6qAtJbPryDXjsedA/QsURYq97NXkEFGhKfkc8CnZDV5K07T8VL
O3yn11Ub8GY2oFHHkeJgd2KEyQKwEcDPBwJLH6yvxQPvAdI0RvmOB936u+a+tg64AeS6Z9am5z1w
G7vjKp13+QQ5JQjAQ5KRhM187GjaYACKx6kIhsvxLxQXOUbjF28bEZ3B3YUQ77bR9hWJ4zdwORQl
XjhZOJDAW3WqM5/NSLG/mWwEVIJPJqXKDaICJQNnwLtCPPbBF7W2HcBinVOSgJJlMo1cZ648YC8d
SElTyUmk15jEIEOTgcaM6/lXKjEmmdDunfWaJktbw8kw/LMcW5mdgcL9kpWWtI9oOMy2sbwKD5TI
B67Mj4vxODThUYTd+AOT94J1czJgW3PRTiwi1kRPdPBxlOZcGz0ixR7sJjFDjQPUKuUc5T7huNK5
iFlL5eWujtXPsD/WxahH5bP61FMFt9NErp9Xwp7gtbP37EKqRvu/rs+ebnt5hWYZWo1fWML6vnLD
dNX6ABH87E/CTTHLndfjqbJKgNFZL7Y42oJWIVo+uDRNX6qlVGb8oQq8cF08GGIJcTjFwDHj7/qW
BEddJjW2eIA5a4Gygo7KRZzLEfNB7OyefGYIn/RXpladeZDDsydR03Nw+wXyYKeeoP56Gsmbee3Q
nhtgp99okbYOHZUltEiINfqY7Pc6XF+pAS0pCv8nxojFa2ozm7vLdjDYWMlqixfUz3kzi+OatSqm
x4MlgX+3nLB0PvE42p7TNWhr0c6GZEFAyVBLPGBEx6ofbureL25s1oCP4T65iLpimBZw47lnmek8
I3kqWnonbdkmFfJpq3TOG8WsIXmj/eHjAiTP0xXYv2OTjfSynJ/jO0COHoWOP6N4pSnSuHi+e2zw
lnHtAELDigf7e6RnzxnbY6PKyzwugYQJcruTjFt35uVNJ20Eaax/bqWbK80UvPECTVMrpxKckbzo
qbGrMrjGAvm6tWmABmiUTLOgpLJS+Y7+etw4oO/WbTSNFSocYuL6cTw3QaWfqicixORxwj5p6+I8
MZCslR8uTSjMxf63BV1EqU9C3VQOi67WDEnSHQZYXLQ8Uv1cxbaAYkPc1GUZF0iVkK8+olqv9VNo
Hri0UHrwYctLQ66J9YgAgVgSm/mXwEyUWDEVCUlAwm/V9G2wlKi5qvLMqw0tSE8LzTL+iqXgyCpg
81RG61In4Mb5Wr3Z4jX6RQAOudpfuqN823UbiwFehgBmeUEXbZAUgceWcbWYW/Z1JFGpMYul57lf
IF44uPLvVdDsBy4oON4ul/YcCzP9RDUBAvRINt9n59vS0AZt3zx/jV0qlvhmR/PdNf6dYGj51Aw/
Ma1hg0j+5imIy/3gbC99cBLB54Sl4vSvKIeg5bzvyL+4KhZrafHUzvhBRqIbvM2vKkf4u3tRmYsZ
/PB6RdamifCYxzTa4YVUksbcY5QfuKkDyMQ/7uLP7Iz5dIrJbIPK3UjDlycDYVn6a9BHHpaUJWCS
ylaJZqXJluTN3HmINPx/b/J928uWVJFxO+yE2QbdWSxnNonk/tRSfgadrT+ADDUGnopvM6Ibk73H
Bh12haBfECHUxgZk+//aSe6cAUx2QnlXXtnguTn6WXY65aZ0DrCgnn8DbdAexRkgQstgwrcQtV8W
DcNGNjh1Igol/nzJjuUdfctHhTLnkPlfiaEIB9qObFnXo2+aXtYqTLKIWRc0nyUuUmvD/rjs29yi
Z8aX0sP1ZVgPceDHm2BecpE75qlPw3PlGdhakNHEC9JeCaEWxERimuxgrCZ9nhIS3ydUJDBwzAC8
z1Ln2m7LTZltrH0WQqBif6kawMNhn79b6hvAWcFTrwmj2YFJ9nzIj1nwZ9ORJVvK3/Sxcy4JDuVu
FAT37zfHBgFkYPH4UNmCrisSnOMrBLQnxCKAuGs/ZB1otZwea6ISFNEwJ/8g8Rhv75aC9blG3nir
DyGOqsMpYr7ITtND5Gaj0T3U6tK0YWIlRNn+9xuWyEjzP4bTp/Wq1oHhXFMPrMKbfwcH6zyh08/v
wle+XG8xMGHqviGc9pAGbpQ7XSlFYrtylblY91zRSWnLpOirTa2QWNIbSeSocVfuXzPQbxV2b925
nRwgLHDimC6W10lYA1s4XvdV74ESEGMdLQhtks3fERHtfg7+URGXYSRtN1ylpwYx2OsuChEOfxso
IW1BMvFt25hrNTVRzMWnq7S79AV0geTt0WISwiJbAos3EH3Ah95o0XUoebue1G4Jw+6M5sgPW3Ik
gtchHj/puo3CFBzdMxzeQp3hoZ3SoAqDaB9xXf6/L2++Oj87UwdTDl1HiA2AxtvFWYv7IfeZRZei
NDMJnp08cnha8OcMm/TP8HD3OC6IAMeWHWD/j23BsQcUyrm7oG9FYV8H6Si0ZHm2umtNU49p3Sd2
YPrQvwIKdiXlBueUu3pO/o+2C3kw6whgEP3FAkMA74J0pavQzGrZ8U+K+p/z/4znTHYC0RD5SMYT
nAuJGbVMkKB3RyChjM5OdxCOMdwDR/QODj8JKbogOwcLIznf/aKu0NwlmkNmTBb6WgV7SUg+HBMl
1lsysxrsgkeRzR2F0fLO6u+laii/JTpC7XyqAo/jyypTFF9y3lUbFMM1GJAtd1QpoVfk2jb9m5dV
1N6iM2zC/l31qz6ml02kfuPXa6+5OUOW3prGtiHc4g3b8IGM0hw+p5Uur6KihxgnfZfvAE7qw+L+
sZBxSYnhSPgYbSvA8R4GT1Fp7cMAl3uQgb17oSo7Wb+/7H+J/zzRaZJPsGZSN4M9XagSphB8CnIg
hD1PFWfZgRxHhPZGSwpEx7v9h8KN8U4EzX78O7kS0sjCKCozSKowYTc0EvwiCN7I4A8fT5BC94xz
sBASIeSoXNHH2ivfSG3sN0uqlHN9QECIvgNrs++s7wWoyuQTmfIbJm1E4uWIzTJtH+zOSLkXBJy5
PwTlr7nIQjJlUv6P+yvnMUvtaoHYTfTK+iPrWe4e2UHbm8pTOu5FCMBYujqYlVjVHSST5UlocL66
pJnpIltRFYmdsrxZhV8SiCnMt62KOx0pOsUCdLlSKa8fpTq5/HipeiLaPlviJZjb8QeeX22C/RM5
G1gYHJw3pOhdqhrulM2MT1pRo9lS2JJ1cXKX6xamNpPCmdlFWj4q1bwyU5Kq2h5Le3uYO7yU3kB+
vqQib8RzLMo2eUIQMxLIAE9DbcG+7K2BXCeAjAe6pE54oJjmJzV0IupGdQUv0+eT5nyYWAZSntLH
a+/9TJfJsmFnyk9aQGI/W9IoxMH8l9JSkUKQtLN42gso5j06/yKa8XqAZrT9OVvJMjsfR1F/drKZ
X4XwOW2HecYH9CUh8fYspzaIfHPua57xrFdsbLZKrwA8hT2FQJgZb/yO2xWRaXZrYwz8zfRY2yDn
fT0UPSt0NI9wSYNf83IUmm0vEPDsWdc48FBgjuAFRlMtSqcAbzvR6EVE8irPJYAYNPOMGRygJ5Ny
iHn75eGLxpBD3eCUGkqqaLzduee3k0jlXyPjoijGt8UJVH3QcLeqTvHQVude2aSIZestMkK7laaH
2rTR8pQ68eF8dn6rAQgWd6ORm3oMY6Y+Wv23A7ZZGNYqW64nZp9LHdrDQ40/TspMViu6rllR3BUb
YgKLsynU5lGsgGeke0pOKTukvSE3vvyXVrkHdfFtzb/akKegzqckGqxboFQrARHYX5mf4iUkMNqS
+1iiGEV/fPtPgf21y4+csH7zPLyFUKYvonC++XoA8LJG3tHAhgt2k01JHR7z+O7Xkb85VfaibSGI
TgvYZoO3kNlMTdOtbf9SLgHZtIGoxjKn8Z9sHcl/m3hb+EiiY76YUduX9JAmqMY4JZwrF4301RF3
LKGkVZO9cJanZ9J/kMSKM/ynJJjmugZNN84ZHuvJIPDk3OQIyJ5NJstBIrQvAmMq2ZFSDe+p1pZ9
2h3NAWr6STY0JuTJVGHArALE56s36akZg7C1g204JYNUl+pCYg9qvdkXg2FUd9Myg8oAhJDLeA9f
15voUu/pLT90Uwotu2D66fejDQS54HH5SXCZabCcmKUkFazArJC2dZeIn9QlqZtghqBa5ibT0DW+
zTKliDf1+0DBTAxqR9XySyj9Ekb1jexnQeX9um05pBHmMOwOuTv3leH/RYO4KER/ZfCOxsj+vhou
KBMgS4wipMzHbdp1l+xrkvohQzG5KlekXzQv18y8Xb+1/f61imGzfitxX67A+tXiaedIHieS70KF
lCzQcJ7DvTu92LBU8MGG+tj7ULEjIuTVaMDUgrXzI6GNqD8eD8UA+oPdoIoJJer/W+cq5Eoqt/Kc
xl3uf/8GqUaQc9NimaWfyMQcWFDK2kPf4qeje5DaNk1yZaxk1nGJfXM3rR9hTk/oFCsVrhlQkuie
ZPoBujvgrOLeduh4dd+eqGBawcSPMJmBwpMLr6GzxcaMuHiYdtyQ2dSlY34GFfj3yX8x8l5M/JNO
LRPB1RqSZ1Qkty4etcjDTX+Uzc4LFIR2jGhsYZ3A4VymIGiBluaj9ImI8HpKvqrmAzCedlz0p/Xz
8YsfzYiQxvdngebWXpHzy9NMc7k/uapeSP2rTlGc2kk3amhI+oglZuQCs4BzGCcvEzDFDmGNusr9
HENhmbH95m7+Q13kWhamZww8X1JN7/t9R9oqXTz2RBOS7DbCk6PG6MeLUbCnXug/lJZhjWnnHyaK
8dWYcuEzS11HD0BHN52Z0je2kQKExu56rPT0fd5s+ZnhlJRKweqwcCXPf2hhqnbZogHKUNXX3Dir
5QUvdUhNQBnsb4XgXtTOFkQJwe4AovbYknlwrfq7pE7SCrZTLKg6rI9ItwX8SnqoXsimtx4NuGe4
yHQh4fVM+HQyLvEi5HWk7a5UrRyUW5hgUTK6zlQmdiQwtcUN4FgXEoHp1JgJ7RMcnSBb9Kj6RmI1
YNUJvuqDBPK5Dwu37SAlCl60ZFlRWzW/2sflyKW3o06lwiBIfRZpg/ou7siP85qKSu2bO5n/vvTY
KJRm1JGua00xmX8afJ1a7BfFxH9MEOpBpgJQuVKWuivawg1NiSSwVZ4fvwa+n3HcBblCJnJfW5MO
wCmc0qalvr5+l53iCqIaKBhNfpdyc01YKNahdwlVe4DGlk7Nw8ViNu10x2E/zaB5krAUjvRe7bbb
qzc3wZKhWszImF+iDb1bPhKYZzD2c/Ufjx1hG8kNp9FGnG5MmElwCMH2mygFC9wrI//zTwVFfiXG
2wbjQ4A9b+0KDMY1Zi2K4FTcR4lavHNXFeoDRq5XGr8nYk66HKak3X/um5P5FniCEl5mPN8j78hx
oGztfg1R0jGxfM0qFXUC2eOLk8AvNqz8PBLvoefRkMk5G8Gz8y8Iqoky9VRedSCGvAP5Q7OE3KOL
VULAe7zvPX2ZgdZ+HBSdFmrOkXccuruX4lnK84jqIfrYu+rTp9Dj6wGr+2PB+ysIbfqQWVZ1rrBn
EUdhvGG7OuGKD0uDWUM65vW5PHLjeE2PQXnG1LY5WE0407Hek41mPsq38NzGziVBnT+iefoby0mM
j+gMPIiRcISonyJmuidj2XjkxewtwfHLrrzaIc3H6h5r+XELUo9uaByVfudegQM9VDjnNkowBvEC
u4LYTXhjDLNHpwNvxYHu4eVptFodYefmBfEBhCMBXTS3DZyjkit+HKQ158ik5FawdqiuKEhQOEsT
zc55DtfOTLZSCUPgVN5hWAcFJqYAk9UpZT86hRFUIEjVaVrbpjKn+CTSAhv+tdkhL7bHu7o3Uo56
/dj6kWQEzk88JcqF93gTA5snVXiDhMQ9E/vspi0pvbgttO2xhMBw4pE7Uab9jeIVBsYtlNq0AsF8
awCJ9M9esLLd+A0CXZ+7laiOa7zPMuOgr6r2yZ9qHcZ421x9c5LFlM+4e3MJHuhnJDtNTCb655/T
MkcdjTa5SXdgUiaS5CUxeKEgWm7G9knyk2WfzptdGqaMvlV4gG0SGVnYVthfG+2T4+YPcYKCuARM
BbutHO8bCcvRJF15oqIBULxS7Jmh+qh9PFnJj8BNRyTczCMVavlU1ENWPgnCbgyZ+YN4FHNZvK9n
mvQa6lElBoh9xRHfcZtLTt6VzgpMxkM6UD5wm8/q8gDcEnzkgBdHjnyPTO65/c2AE90gdo7RZHw2
8AYJXZBDrv5yimf9kHgILU7lEOoiaYazNV3WBAxlf9UUKrmLZgx241WNQhFYPZwOkirDiv4WuxZp
iPau9VP5m5TaWEjuyhI7W+adBZhuh/GzSbI6CIqL5XmHC1FdH0b1l3CRw0XVqakgGpowujNXjlAB
MVh5Iac6YXDmi4IE+e9Z+QGbA6n2pSQRmozOhSk0QvLW/1mCNPnj7qc/qvohvOG1OYT/kKefr2XL
KD7oMFJpstXxCP+k24ybhhzHHdHZ8x3BWAIUqnMI2r4VE7s0I07QrTtoAJmF7S3jVzwTvQeLB/O1
qLM7dCu+OqbJxcvtfP2NZWik50BmJQM0DdT6zrzCr7LRxSAjdE9tiAWz0oLh5h2eOFcTPkY01Nl9
XlUQ3QfS9t4pqK5PsrMrEmEohsW3vqhizkSase75j/Sac1IgPDl8cDi9Uk33bzHMMcn194S2jqss
u2/DSeTbalIrVI7YFwm6OIoE1+8+HmB0Q+5YN8BB++d15VufOlqAA2B8tVC7HXlXNJZKsCXJFDTV
TtstlbLUPiKuXorJVKe/tgdk1HRKOU+xL2VUoBkZt35nk7wqml0UPEQ5r3JWcwS+/zeG3A69AZRg
xJAEtbjLqDPGaoeudArdvU0/XpficRQAjMXzvFuGVu1SvTk2xJEm1wqbkLgmj7TWk3Q+vlaYDFuN
2/jxQSQNKUgz0rIRH/5l87Vt1qT9edQ5+RUfgEUs9wwIKHzXtoBCkBOu0/H4eHgJWQUuazMK2jOQ
fdntC4zrIVr2OGmY05fheM2HhdA+3ig0ZcPGma6wUY+XcU64XOpBP+FGbTbWqF0m+PFmNrw9I33J
8vmpBmVloRX5wMHEIaSpKcWeFlhvoJPL7KEJTssMJJIDy1ZRTsQl1/PEf8gdPgCYaaonj4YiME9V
mdJwFtz12nskh416pYefhHpf8tjHCGDiZN/4JYCSE0jC5K2gCMZtce+q9H9cs5bk+7CHBcXIoI8n
S8fvcajAivRRNWCvl8xddozcsjw/OKLn0nUY5jfV8xGdc7DgeyBsRtaSdOYDEMHOHu6csaN86X0F
pvmYeFwnZrxNGUj3Hdz2yOBeTzKD/wLK8S+nfgqWAzLW4tBTOJgYgBJbOjY1v6pAqaw4PmyP8l5b
SJUbmvtXrIHs1/J1D3zjV02P0O83Yr0C6SEbDjFMWKpfGVgGu22XqBvzOngJzcrbtc5WXdaJw8g5
VAV1ugWFHl4w13pAgnUNnLYH199GN3H1alsjCeQbxcQqX2EAdEUj+Vvwj8YpenceeISbrqzhS28w
IfnUlZm3s23GgvsqJGnlTVsRjajy/d4fArgI3I9lYmTXVSVwvFoRrkBNmyxRspP64fvXBm0TeoRH
70dJaEoU3bfLlonB8t9YfsNj2NmXE6D6LcdyWL1droYCVbhiLcOqV1zO0hIxZffDFH0x8+xsduFr
nMfCI8sRlQ8cGINsESETxsbzajFCne9Gjv/SZ0DdYw4cDwcBSteXbX9rkPgcP7dLz6IZiuK++2mn
3hhs6UC48FFLvw9/sXEk8KMA+JxrU2jmuNWmKZyBIf5tmZpd+sKhIBxx7n6DHV0wsoW06MBn1ri7
M01U2hIKjXYQ7VpU+KICUCq9TlFc+sHE5LsFiYUp4n7bBcMRH3NXPe7kQ1UPh8BWJbg3gpAfs4jV
3WsCUQqiK/46hXzgAX08em2wKRMtWxgdb/LH5tEArzNaNgtnf13/T9P8aTqiL9pJ3Ej++r26Pu6x
BdQBThblY/i0cAyR3S/EzHDiTYWhebig7us6l0qc1uGfzhwNeOV9DH1rd6L9puUmHtmNlK1zBW8h
kgVjZH6l9YZM5b9WwOk5mFEtMZoJkrz1bs2NyxEFnmZUZNjDNPz+vIGkhiFnWHydzZ1pB1SqUW4a
7LrMPo6MuhC7GxAaVtDdDqiFR9IqePMde/GY4XeOz2Y5vqiw+4mACqaIOmYUZ3FXfWyWb82BHc7m
3RvHq5wFyhL0mwid+pZ47rUscr8aPeuVGZpZaE9aq9B/DNtCZdPQyY9FOm/0UPI07R2KlfRUp2iv
U2ZuVXi6udvyWbg+GfydcYK75sSYRWhcNx58Q3+hwTQrMpX54LRDhpj8aYYu4JiJIA5vyeJ9JOw1
vfz1w2R7MUV7TGxdib7dAspekByQgykVwrpSWYt7wc45n6OTKSfcyn5EAyGGF+nSpQ+6hX2DLLfR
oYZZ4Zboj/rcwjAHim6MY1QuMfgrqGaAf8SPFnXQp3EcSBLtlIYPU+UQqx0oAAyroXkk0WYQ22TI
jSpYxL7qa/0kMohleIhngXnD7ponhjnV7RxapU26Y4yCkOz+nARrf75FW0FmwMM1OnlOOiaW/wli
8PrcL8swG7HKZAAkUbcsNg4nvd7dXVIG7kaODFhyG1ekTnSCozfhYsWQhoWL53RHWhF4k7SS7HLl
MYxxcyyeMOvwS3qHY0Tpf6TaWa3bWrYiHmnCjgHULqyqnL28qi9g1tPVns6ZNwO1Rw54alpM7dXE
IKbsR4JSRzePauDNpfl0HIenee4yAHA2Pxdms9Bpns+X8hZxfca+bFC9WYYSsy9AC+Kqx9A+okX+
GogQ/M0gdvNlrJZSz+Tc+/dfrfOBReSDTgHpvMJGb8x/OuEzlU4xy6d0yhi6rAJQSiTiZBFCHmL3
8NLDGx9NJI59WJTttK4HRUi7uOUmuZ6YhuCNJ1LFzw/n764H4pl9QFXhzSAJnsTdho6dY3JxM5xX
dbWdFRfMH1IJuoyJGqnHOBVchAFKsB79vl5mZ18zDJVuu8bmaJMbG/b/WqG8RWH8SfjhWbybPa/o
LRcAmwiiamwzv2RBwosW1ojEn7G+ax8GOkYC7l6rEYhNi1oaDPsddGe9CBSLUmle3LNTAZ1jUSCw
8SIL77ep6/3LMuhBFb/GOuv8uON2S/AtH5LUIU/NmwNbbLrESyd03HPPol8bk8D7Gge7OR5PITIi
LlUybsw2lg/JFmBp5eW5wpJHZlhjnlGmLKrprWJpacHO3AF34qVWXo6okYTvMMhnEQwb/Z/En3m0
m5bbpvJwITFtse05Ze+jVLnRVnKWQCM+zYJ51bTm+sEFCFncxLWAHcA4fZTxR+6FYjBEdNa63VRW
eKet3QEyqICIQcUvs2HvfQvyKLkLhzJuAn81Rn9QMevxzSHRAJbnop0m0mUXGM1NUkkP6E6xzrXd
W4lWMzIFi/fBOGTo0ejZF6tBv7c4klqwQeFr3+C3Jk2JE5EQlk8uSnTL3C7TN+ATUJuKdy7If0uy
HLM/EFcSFWe7ilZ0UHEg0Z3E5g6474mtFgvRlcmVEuVekYdkpm7XZps2p3eCBypdEX5hcEPHu78y
XPZJfYReHMHlhwa2JEmmz0llBIwYfeT1OC35iHkE7mCh0NjJuazgsvJVXGR0qXowEcBnE7kKHsuZ
fznAf1f5rUVIUgNeulpPuH+lnGYRmrmS4dnCqTrIeYWDdVuYof34gytYjgup96KBNWENiIIr2J4p
OphhaQNbozxF5CJpkWAobIistuwWas/yBcGXYET3MyIvvq5KO1Hc+TUV2cjbkcwuwDlON69ITb8F
dTodb5HfO5+3ZJNAy48esjdIQU+u9dM7T3nkiUnc8khXOx4nuKASkHXSxaOZdDML5Kdtc2vFFyKe
d0IdaGnzWyQgNPD8P3rKPUWhdWHwbZP/B8U6GF4uhHAUCJ1iFxiiROz0WSK1MRrFJ8tucZaoAf4P
dlxh5FBCPLi3UaRuszTDdf25cw5AgsXzKf0+XYGhqpPvi4Ks5TUuR27ykqybV+MpC1kPOzHo9nB2
6rRoQNJgoXBpBmocSbMegaqEloI4AR9w7Tn3ShSj81OMor3EZktFk6aND7AyLywSlfg58TL/KFIE
MEFTFkOk1zOXrV10ZUOXyDDfxtxWUAGrxmX3eB67g1kaG14l4eTLtlaUzfLgjaOv73FqfHn/PrM1
w0V86Vt72DhC+oBJ7ikDKFp2csssH7ezoqEmf4/almBEERdUFHTbkDmLwL1atPbAwC0pc5eLn91j
LR8fTERpxRfuAJW5+g21Bm/ipeDWPHrqoNOwBYq8eaXo2s0hjfQVb/r4l5x/ZQsR8a655F1IiEHu
GgVHBdD9VWbWj9WdOGFL9YPLkjuA4YJjYKXbISdhYiyO7a2yljenxJLUz3u1N0lHppKlZ8O6m+Af
Bp9ZegTisoqygtN2gUy8j970G7KCQLPJvLkI0XBcblF4WauRJxFVBbK965gzsuPGNUdYShotccJ1
QiORKhQTmo4YxMTSWiBkeY2uy0Rpk5qGG73I7KmuQvEAFcYIaf4a2V/oQBWqkVzS/F7OKF6Z+Kb0
p92jVTPGYm9rwH8FxMP7ZoKpUZXmTqLjjllf20CKiExTOg/mry8jJMSiPq6MzPuD4GTEEyO9kboX
MkNXpNGiPGW3dT9FbHnqNSKb6g9VK2QBhVlNUo6+6B/W7YhN3NpOXk/aivSRnq4Cl2R9/lNSYGJP
eoGNppRGrYOVTdm6xS2v8V3iyCcrLaowsZV1FsEyEe4JT5SXqCL0LtSW7zaK5J8HQKn8Njg8w58A
FBAJ72ITHnURecfBRb0YgH9oo1NNIjfCb8/lfngGJDzoLvQRXQKTZXrOGH+qx/SU8+NzrLJYmh7D
/jWmG3WbLL0GDFn3WSoTfddud3ZSXOmckaecGhVtxfsdyALAAH84IdGxxBQ6dBgJSI/hSloB6bMn
kyZV268FnQNxf7GC8QArup5Dor+RIIw6JGz7NzLyqivrGhouXTgVEjZCh9AdusdmpA0cyRGznjvH
Q2ZdKHLQL2/lZcANhc5JYohBQyV3H4fweU25EAYbwEKupTXBWrsOI7i/Bgs1YG8n8opGrrum6P1o
dQ8Fbo9XfVRMxT/AM4lSqs2MFic8hVv/m8lOTfmyTGHnjWhEK7uxkcSmHYtL/MPcEfbUOVvo2zir
/2o1uMus/5oo4srtUusMIE9OZ7ozXj1lfLSDD7ZlNECKr2M13+AyY0zQHUn7eKzHL/UuOtD7DYou
SDGORSmmZL88kzJz8AyVK4v83K6EEXm7h7xOJWtZKaJsFX5LrJEB3wNsMYdIgsioXpxOpufhBmFi
JGC/Re36cdlH46Hd74Sx3A+lFNpGjT4s5bvanFDVK6+dhAJPgT3hwgxhZ6jNIdNS+jfdAmh4brrb
h+FHdJvoZavCVEnsGL6DM/boTkAVQpYtxQeAtuvT9sy/WLvPS6bezOTaWI76dmiH1UPIElToHRXr
BfaaH2VrK12pZI9RWKM0opRUhMb/Xt8RRYxqzjdpMJ4t7MvR+pLFqRbbOPORNW61sKm29RVJfoxp
cKeENZqEHUkbFqUfEdegGvX7mvQ2ZBsvja/NsaezNXZ94NiCCDOvDhksDNjRkT5fSr5C0ED/BL9T
lCjuQ6ZaQ8MV/SyaNpNnIeltaycRQnT1I3Cu879F8UVFedn8LD7QHf7cdXFbwsASwrArGh9ikY4C
zMKXT0FQBgR/NDhDv2dFgaeHyX7rk1dsK08Mwv4/cZI4z1tToHgquKIXiWIuWGSaz3TjlwvAEhbU
eyY53HStgVtzP5VR6ZlwqqVQPDqfdx87onRJVApbNbRbHprf0FLtuQu1gjvXsmkYXUyNpln+gNLK
2vanQf87WmQmELjfiKT5xJC08ZPCNwx2UauFpx9m5s1N0n9sg5Q73Vgs4wMYBZQx/xxJyJyg5hEq
lEUb3/R/3C5vFlX9Y6/X0Sl01gc0onwI0Qxa/2pXmXNcQG4va8pkpAi+hIx8rEBOq/uG0t7cb1Lw
WrRxZp4ck2OdLJWU7lXGtl3K//XMt7odJIfC5vz28YnErI+lX/cyTe2Cwj+2koDlTrUSvYvtK3yZ
zV5wsttd+rBA5v/Qck4bNd2qPM0GNRik/QW/W6D4S1K52JLEOMAvtDVrLsn+VJG84OmhYgOto2X4
UakM/2cURGAn+zhkS8ynALkGM7hQbSYnAT9Vdet89FGOLT8ILKXIPkrxCA50Xxdw/eNB8Vy4X8fu
pS7WK16skYjA8L2qmVddui513o0w/z2dk4ffFsnnX7lpp8AtNP+I4ZwvAAmZ85DEM8Ei89GX2pz3
aNE6CL9d1MULqO9+HlqK9nXfsupIZ9EaMdvRkQ42carcPDyehklEqFCvmNuiDp3XCkOpTarjyOG2
wYb5Y+aC0YBwN2icoK+7lXQ/C8IszunO1jEDMrTUOEUmZX0d1oPdbEgUUFeFwcqLapWZSbIlVQyg
tnofhhrPQqYXDP7wWLotUNxr5U06tOBFsxCy5QZ5dCW1nqkV2FK/0JMSKfbar0G7o0sEe0lb3np6
mWA6OPSjU6dJX3NHV7PB9Q5a7d5+JbagEVZ2ikdD4368Sc5nqNcEdWxpU/L3/sUy6Hzyti0XyPrk
kt3Z6sNbGAekc0n7u9KJsKTZhmuvw5RL6km1PyI6bRSZkQjy9rzZpQa2c1UbNYGhk8Eawyd6pdd/
iYHR32fyZDcucDJesOXoTl+g7U7hoWeXHW+kbhjToylsjQePqlrJHZl4xiDGqXHwRhczxnXHAMts
MSn0V0sZXcsUupZ5x6eifeUfgBfhXqkaGrDvTcx1/9/07g95D+Cp3tASIzXGUJa2s07lxG2hZhz/
kW1nTMGKo6JgduaQg3EPUEmcuxjwpJJ637bkQF5U0PXoHK4XTWnJ8ODOvRErm/8jyYao4b7HrKzV
rTI4pO8dRUJi+qCygx/5y42uFa2JcRTlAPmVXdsLnZEPee2cNZ5iqUS6/ofU6kY7imXSpDM94KlL
4j4WkeMKzy7E5dFlFJABx2/wyUjbX3Czu7Wlq1Wwxz3jBlGDh2NNQMxODqZEDWMK9FFsx5yzRBEe
DT7jU+l1jhInFlGLyNTf+50dl9Rhxu4+uaX0u+1i6MfLDomiPGljK9QLsVabT+/P00OHkkEVvpIw
B8j9NhBoGwDwJpV2eMnyLMLap/KEUpQHUaa5Yuzl3zbA4S8JKTRy7o1prs3vQxUlD/dhV4EaCGmG
3bOhx3gwijJQ17TN249TAQ1cEjP3N7sppGRiDZGe88w4g3YYzu9AdkpPuxqtGqZk8YB8e9kaZJJi
k+ygY4W2dLv+YcQefgG8k/o0BaXmjWXiijSITWoiPrI00NmgfrLL03N3iXwajOte5F/gfaxyffIM
CMv0vB1rG/Uadxdt4VKOKhQEyLigzvqdE40xLBxn6oMGMwYZYyr/ELbyX7fU6kbUX+CKbGwjGJMB
ANwMklRLJq8Yy6kLv80UZJiCQn3GOOEe4foJNhPuZvn+LTfeSLSUZ9Wcqr/LPTlMCHeH3ZqXFKMJ
hotRxLn+Kbr0zu0OkZfoQHQAUlTgl1qP8Q8oxORUUjb/TW7OmK3xWqQ5wsZkroN/3SMNZfB3XFmZ
QXk3IB9Lje2WnWD0XBBqDRwfr3Mq4RgfTMFqOGVQO5uvWLglqL1UCl2M8casNi3kxGdyHzJMLqUN
HJKLhNgbbfxVa2P/xWZSrejbyoQpniM6Rytp0DrsYSTYf24dB9L9bk1AyI5+TH13HNhjCw+nK2mt
v4oSPMlJc9x08eRc9gUlU4Q6ZnaMlOJC7Low3ZO2Iqvsh3VwmKxuhPL56z84obTK3OIsz2UzK3Xn
zjW3t+4ExP/aDonTQ0ZklQf9m2hy8GxUP8OY26PkmMrlcp6d3F+LRKMgqfJ/7dixAMvhPe33e6O0
+qsjYdjsEiVDWxrVBYnmWi9UqdB94HNWQYGQQjmqDBMkbwTBRL8pWN1O6m/TnIDjFY9KWDfY9y3h
sQTG3S2AUH3lrKsvbAObCxN6Ubt3ZEQxm25jysUQXK2M3QIjUrkSeOTXSB6mZirmMTWYbFUWjId5
nLP3BO7oT3n1Q3tvpj4ZJ242ulL537pcZ7JrnZdDHb6ugDFdZD2FdbL40YDh7ujAbwXL+tWNWCDm
nMYydAsQKP95o+HnykLZ3JUZxFMPBjDWQewiPH6eXpdbIpT0HLrzecUNJs7TpUrJ7sxciFvfuUF8
7TmXDeFghe7iTEOtm0UkR32gwt1qjKOCdGMc+EHIJS73feOoRz49CQAcaENPYXK9RBnAvNjVqhMF
aoosiJEyMLkU8KlLP9AV4iFcn8oXI1m/gDx7DPeHuRPRBu+shjWKI9y6obaFR0Wu6xggSM0BbQJm
mR3TY+LadOFLd/h5IZTT4IMlz/dsO5nPG8tBc9l8u8I3zPLePLFCrREW2Ij/b8qfERvqxV3/DKjS
o7EzHICr9NatHn04QVOFOAcIMNhqeg7lr+JQyNbu99VFlZWrYNyuRpCmrXdJlkIXH8o2q//X/kJi
RR5MZjrqqsTEs5YSfkzldcM3xu4qJR3y+7fIPe+8FZ4KcqXZY94zlCxBAfUlFtTDFZhnO39tvGx7
xFHhJ4C/NB4GbCgYPb1s713UetnPwoMoLmmHgSTrhLNrfI6EzDzFtcHV0cmiLLDPUT5rO+QcRaIw
iDyLjgXZlf4MCJk0b5VIKlzolPvyPYr7bAgvI7TJ6QZSIeWIPZrjDZXcV4ADnMYbFPnMpqecHFnW
X2yxrPDFWVdQWlMaIBOY0j6QlPOyPr5lMmanOBGQvjkEUyIMm+xlTHsMdC9Iz5g4u/i8jZ3Cs0zc
PFEMX9LFswVQuderQ1oO9SJ3uYo/Y6f4jzemDuVNfq73xXbV6fdX6kU05e0T/7wKFMRrPSIPBj3w
FnUvq2aVXMuGTuKTaF3zCPe5YVDhhtuxravJu435aEwgT5QrjZgvNMQUUfSSqmvIKOiPmdcZpvMl
ji6MbLc8RqmD6xOIhxyalrUKCUoxaLYatSt4NQz+SNltGFSFwumaCtBvYHmTMJ2zzBHNdr4I2q6T
rl1gEuHZbxrQu0Q/hRIxsg7+iqAvK+dsp6hDhVMClC88YMC1lYBUD7kJpDgTEM34gPt1dF3C8ZCS
/FSWYYOb8hKK4leRcK/01/jUw12wr8OKE43ZMI88uQmotcvkgiw0laqO6YMlyLg3qJz3pZBBsEId
qu2QNNsD1VQ0ohaokDCn5WehFydLTJRZC8jvP7xP0pKOfwY4mdB83Go5qjR02zAqprT/F8zUnfki
d1ehpQTBRqVQ9QRIneV1Ed0Ljh3JJa/Tf9trGkyn+bvIsP8pcnFgGLaJnCeokRCAaAL1JFyoRN7T
TJVzcbf/4isvSFkJgZtaiJiMEBhXOnzBuNAIPQ5vFY9FJl9QyA7qR/ydb9hpgnxYsEXMtGFcX8BJ
fNOuwEfwFpXOnfeKTcO2R5Dgu5jMILCxU63ivb6FMkoT8QLK8w/zk9qLybOwyblEhZvBZbRxtczq
4NLwki2p8ApIWknzeCjC569sRwtTCHvW5HHVRHYvJMb0WAkcY4ByNJBExr4hPWpD657sIHYVyOVW
2h78hnfkCeMheJWa1RJGkVsp5N27/NGIPB5eC3bfRbsseA32+RlmigLZEt0Bn5/BNd7Vn3l1ZvLu
ryAtTyNtGB9sINaBgmGZ8/iPnnnhzjPQVVUb6tG64GrxvBWtYxB4oVvLjU8JrxXJ/H69hJxlN4T/
2RltUhJj0CIqIexIZsVBLd54VJB1MndgYxBSdoBgjQHg0hzcQ1OFxyspDShaZO4Iq/qvk7C0aouV
garx9ZKE0ZRSmHO2NAl7+0AVS+yIoowj9DclhZtnyvGf+h902rk9TFz4i3hirg54l7dABin24/Dw
mNYCrJjsd66sCRq3OCpQVZ8JTcVqKL9BsPnhjKnQOXHkXrFfZU0tvdbrG7QAqVh7yDyf/sWuMgW7
EdO2G4zVeMe++SK7uuWbpFwnUIwHUoYhyVRAXmvqK5JI3w2e6CVgO2tDaig+DhAvlI0LlZ/Cy7YM
sPm8lGQ332bI84SRV0MzkQAeYQHPoDhpDaXqzJaDOR9ijGwuw5hJZgq9vym5bJqHFuyHL9X0IYx7
Ja3QDRLgLyqDzTdNfmu2MYGbSH/7mtYCSw3u1SbOEfrGJB14uVOZaANx2QW1MbbroUWhv6hFC+jo
/yFzhQbtmlsLG6OAwvOUUkJFcyJNuiYjIku+XmpR3Dg4Sj2wk6eXeYSDdeOe8HEGC2YjHmPZExNc
PoWmQtKoiR/Ug8foZNSesShYLAG9BOdenMoXwkPCUWeU/ATyh6MIE3/zaPipQKyXSwODXMkIBT6K
Q1icJBbH2MjwVOSsSFEkQK3i0b1YmQoTaVeSIzWuBVWMWzm+H+bTOwBUhAHneNOemCtdack/+yP4
AelqM3fUPHR3mRpkUe41IqSWQ6l40i0ccHlSPwIRbCpJgpggUHzLgGOQidm8oxoTqRJIYyYBIl9B
Ug2KaQgrmyipFooS+lJntTkQd9a2icx8WhzTseVllbEqCOAdvGEJhKb8gVKlH5XpBtQR5QJKOs7n
YOxELaBHr3KvKlH4b2aZ0kuHBq0aPX4eadN2/uCgyTwosxJ0LMbtA0LewaEx+fNiX4x+Z6h6wv0p
MqJI4d5KNXvK67AivFBFESScXefzzuHqskcseRRLtjvDh9a4x/UeminlKt2rQqFhQoqHi2wRMyIK
Rnhxqmt6Q85hEmxtRHhRMfxyguBwhcn5s95O3avl3iv76lLq3ekFCj1NtWEPLw4Ny1rcBFRu7iTV
Thq8lEzeKOIUGsd00CEpPhSc9qXx+a4l7RJDLyA/NDOsaKrg33bU56h+RxUfDydP61tfVLUoj5sQ
es7fERvuGtAw0kvglo0VKzb2pR7Osv2WogfAfe996cXvvCYsMgjwRWKrc9+KZM+/m7vdm7OAyAV0
7MaRsUUu4UO9XPvxB+f9/I2+Vuwoba1U4stqLC9GIsxS/QUwOxB4FahvlW5gpUP2RxZU5/dv/P2B
9ivVuQKrVSob1NpSSX3iq+BRFbyqNx7k5pt53A/xI7B5t/d8nAqAwvemzSY1UCXfA51rPS8I3RNm
zQoUXYqg5LTWaKaMdCx+U/hdhjJKUeDE0Cf4vOWGy9SCWMipLcgp7qAgUHrqlYIEOGzgGZ4BpSOv
N3U8PejAxPafjq/0AdwwiWbDHa4swx39Xrg/kdxjlldRcM1fgonD6Oaxtvna1ymsvQHilI04VOLr
r0nZ2fmlS3VxUOIo7dbt6zKnu2bD02sUsMw9JoENFHzpLMEmwWFiejpysytnz3HdhoTzxa/w7CVO
3GQkIvYvvNO1zyVEX0EDs3bbjXT8cBjzBFTJy3KWEqt7OT06A7PVYWsjOyXiGNNxj6LhKREHZvxl
8lxlKJ/EZIbqSvgEFo2uV9FR9XdrEEEheheN4JA5GBcuxqfJ9d0mlhoNOvhfXbelKhDIFppmJUdC
D1EAm7qsMhP3KEr8p/aq4J0btYZnnkGGkS7+PfECmQAM846xlR9oe8LkaG/xA+HwmbKngqpn5vah
t+lbw2fpnXceaKZ6eQ7EPw+4iw+htpdS4mcAu5AAI28uYF/R8F6hszyIhjkhtvIm0zm5dJhG6Jjh
pWylL53CFtzjFiQEA9cCdkxvxLYP579QMVfBWdt6Z1rq/ENVPckCTaucjdC+3feXCbUXfq2UHXCr
sBXin1LzcgeIwKqyDubjTbI7dfdgPLhe1BvN50s01RQ+AFCDVQf7kk7KqEc386lfHjlnD7tj8vB+
p1qWPSMhYws66lwRpr9BP8KqwoXSzECuX045p1ESHRZfk9MWeGz0DzG3oNpW1oRJdXdtWDwH+ipo
68MiCrat6/rUh5Xj+r2NgiEW+XvVr8U00njBkvhk5Y9hVCL0mZ1XKUsuKNWKkIpsyaKEAWzGCx0G
3Y6P1hMt9GIPAj5CZxpNZPrhtynppamSGdLLpITx4nSHSc0OScmafvD0VT479Nn6j8SImVerk/zv
9subg6w7SoYeI6C6gjmtmZQvt9MaqNUZ7YYFYtTOvpOxBDHgPWOH8b2nAGKt8KR/SRBfmRNIr2et
O2zEE3IcHUtL937nQfXKFutUwPuVFj8BY8oVjEeW25kegBjCb6Y82htiKMBsLT5Hsy0f0z2f5sEo
eCiNhWCqalEsh+MJK3ivpBKhNA5WsFTo8UwtiLScwINj3iiw10uIT16fjZGdeYaGUlzfWSQIBlzi
yI8RmCZNN8m2NTOs1r6G2yVPhYKAK3+e5eqYhcvCizcjkllXWZaKAIEUtMFwXm1NZbXpycefSwKS
5osElcATyF4BCBcldNwkZkhOvRwqEumbhiWgZgi774cbkcm3eQBgrAmJd09HJ6jTqvf96Axn1BR9
tAuS2LNAqiMSGsM5lCMbuqHflAM5gpKhcn+fyat+eqeXOrybGiWsuD3NNlcNoWLY4JqqsPTFRIYg
hIIHj5NRLztp8hmApFD5yFa/lUD41Y3AXg0V7/nd4EDrbhh2Bm+LXFQGoFzm3RAhY7gUNaxi9AVr
6FzgzSeSXRdqbq2kBX5qCZK2nBiE23Ixhe7PBhYhGJlonFZhSEhBpgRjc84Y2D3MDkuZZHFBiFrB
8Phxhlcpmm8rmWhJWMfYyVOmus4bS5NxBl0VXTIbfvpB5AbjAuA99NaAb1w+hYr8SVBNPgS8ZJB9
uELcEeW4HUFYDbMOpZhFBQEoJketRbECO4gHxdJhtrWvKx6crje3m1ZxWJS/fjqbD9cp5+pAwiQ0
6MGYPGWgL/kam+0Sk154nwNUMYjH+FcUqCLtNAYOeYE4WvdwsQiKULPQNRrdR2jcJj8+ueT4bT6l
XJXqLlnDw3pXf7Czh9a0/ZBb9DvBveUvzGc4ZPZ8tz2bsEzSXqamtJGmJxEEy3evJYH/r4h8HrM3
aFePA/dJhjBMSwN8PdDCwzndBqR1uZRD/Jww5svwZuy8jxmZjnMdShG8DNbxuThh6n34DZoNIyvA
xlxoxpWPbQimKcCpy2qhiqpqkII9Dbu/knhaNPczat4V5dw/QWpmrOeR8PrRGHhyYgtrgTErjUre
Brcs4Wk6ERfwVLq7kHZBjLFazQmyEB/hxLYuiJ71Hg8eFa4kRnORZAQxqehBSSAOgUq7aQHg/Wxh
wB+oloP9tD+lYhC7kN03XIJ2t61wpuziVc7WxT/jAdkvf+2EvusfJv8c6scmwUcHZnvenOOl21qk
Q3hXCl++Rghf0T65oU9JpT6v5OrcZUGQUvU71hCGIUUPNtqPRGz9BT1vB8FE7/AQnSAhN+AnOQnM
RhKC6meFqYkyHxgTA0bqTJNevlYHIgYesyG6NqmKAu7EAsKiFZiXQC/GJKzM8jcQlAsB/EwZLklK
IZoMeub9YAxIiVePXOHZeKi9z9tB6oO0LfBd6Lnh/l5/0WU8cYZEVHoe6XhEyYwHVkRXb1/KSdq5
w8I8LA+AKyMpnrZDL/NCWskfl0u+3JFlqzkta8b8ZV/XL65+Wh/uzT6yLBYCuripyhkQsy5oFIwp
Bj6gIs0ATNywEibUZ1BFhf8N5CWgwUR+6h1mck1cxSlr6cuL1mGDRnfDNa/99GONpjjEjKcG2Aer
Frda06LcoVhiEm7ER/mUSW8xtTZNstQvpTonkQm1buXSuF3+Iek0eXT4mRaPXkL8FdmqnU7sI+z6
dF1GldQXM0PLPZk2GNeYbsXII5OD/x3cRyTHD4K53JT86mlMIKTphJTYmgFr/XAQN/t2CVt5JHGD
El6n59uwPDCdSsq8d+aaVWhsQCgp7YKpxNbipsL/aC/Q+GQ3VzH8n97mAhLGqiUP6QWc6Ln9Xs0X
xToXMWs5jvPD8IGHllW5rxOCrYmoy9Tx0hiuZNvxhC9YBAtVRBmhDZAnAmQvQpd1MWNqLLMBvsFt
BGj/X3g3zg0arykOkJpeUFPUl1qYMujc03NyPF5tQ3WHeaEUvc5+6X+sF5Ny9VOL3eCkCsGxHRpT
tnvvDG9iMDTyWyd6xD95aZZQdyIVrp5KYZcbsnAv49dnBjfaWps+mbekqIWF9jZABGO29stStAyp
X9nhs8p8Q98Y2hBY7tYN1lisiDYXfs2yDYomMuyK6yuo+lYMtF9DOOP2ddP3DR2RU31AkIcCDBOU
5tPUutPDspasmupW7ORxp6Br1y8w7wCSDhBvU978L2QDsdv+GgC6QroTy7VGyJRA58M6tTSEUHxg
rIcL1XvRdy/hDYOf+sgyhzq9hjRnynQ3mADsOekX+srK0DcteJ7W8/6wWarfANfcMKuwXP/uKmMf
3kKK11nZ7i1srV4kDwZXWz1LcueTnFRbNPmsb8I24t2+nmNG3WTQFgJM97HPAOsbeCpm8Y73zEDp
mMXKcmXfvSdrE+KOcrl1Jz9hrlVYgpB6Y9v1ttSKKtCT3F66EMz1lFv9G+f4kvR/g/b2IKmVi5us
XgN0Z6cA+Fx3ehp1WzCdX4mODZU2MX4Bz3rmQVI5/Q7t2kaAwoRtt693BTRU3kU+8IoWuuy6P3/R
1bzJ1cOl+wfWggtsNLhgjvNQXb+FHlDRh0pnzI0BWIgvQ+n+FGoaQQ666QD3YeW3Hb4NYjwFqYPu
u2uI169zSYyEYh1jBWQ0gH+st1FkpHHe53kZrUapVXE4D7bWQuOWrq0y4cQRKmXkd1H4XyfBKyOk
Prh/JShaYHM4Qwl7HYEYrzy1w3ZU5FWgBk7oHbV1h97VKexLD6S8H6X2VTU9i1z/UFrOkr+fD/XR
VoIRmzjYcc1VsYrWZI34S/F0QIbaI4EmC+uVtTs6u0NCd18mneV5wdoxjxYJz0jhFzM/QWsL41Vo
u8fdlS0lHsklj+1X1PII0viTfTku+YrUR/++2XEcWcnaiKBPxdnbZ/Ktp4vVMm30DRhlgPUFFeoP
MHt97q0+tRl4xhMdS5HQNe87fYKeZ6jFiFI59zIHe3UOcZ83cK1BhJWHTkczALMibpnFUy1xwq0l
BXiGZLfiVZMQTxYvpBPnrXC+UDMagKSn0L7n7svmx5uII3fXoumNFN/A85HJ5jQgVYq4e5/DiiIo
nDCPzE5D6BALfQS/ojR54ME7n9FT4bgEFkAy8I9sgl+cVELCaQy+COtC5MFyltXkQsQO2VNYdmkU
glS8Hvmrqo1NZtKzXGBPcviZnYTFVam1/ga3+b5PX2cinQL4UPhPNigt6Dje3jzb772jKxXjZjCS
vzEFlbkgR+VjW/SfGPH9E1nvSU1qNKY/3KoLXbYq/lnccknByzaAyu40roTDiZKZE7OTG3Q68KWo
nOolKPCvEh6GpoXBHVEJPdTleDtA8h79F176ocYe9aSz83OHwinntS2F7xwOafA0ASc+TBDSuZRk
b4OK/IGBHsAS6UZuh8YcyRA4nttnsyJ06pgSY0SGLZ5uDSyMWAC0+vi4FBUmF4AKkXkpvTpgXdWj
aKORjIzfezgxqyaC4VymdHW2XvNO+cRp1PtpAZSM2PADhS7tW5FGuj6vojX+IyTFl5PluLuHwR4N
a6N82aF0kpb6EQG5+LbQMnKPzILZKtwHVEB5NCcvoMG36qK5ijIW3Pb9AkWpfUeBsYJ9TnVQgW/N
FMtu48gijUT1JW8kqj8VzkJR6eWgm7Fa2iTUaECPveZRqfKat6rqBW9a8+LbSOzZ/Wk+CylT2PRL
eAm8Nu3M5CJu07nFMiUWXQ1CGKpymdMQPTM5VWBxCIJTHZCk9ftL8GXzimd+Ji/r3HTSyPieyzu9
Dp9ezoSj0VXc0kFC5U8baftFSC3gtA/QQyqspgqsQID00HEa07imOKOumcbFWNb/7SVRe0gxihat
uNfacUOP39uWIJIelnoRAp+VEqPOQ3/QxOclkquWG2Rjmde+krQm43ym5I7kotUW0R4ZYzT+O9fz
GlBwH9AOuHv6W4o3Kv/Q+N0dRwND/gWUF95orCzsW4fPOz6gbsXhIfZ0jmhVjBSkt8n08vCjZ9IR
ra8KpaORM7ietl3lLo8YWw2V4ZZHfbZBmuYrjjFa2GcTbxCkohvGn9bs9KyqaAnwX2C08m3QvDU0
cpqBA2n6PVFhhZVZp6vpQlbXAvUFfG9PUzFrbZJW8v7zcdYBXi0m0Aphg7+PkLoj9qkxUsQBFoou
X6oEnthZ++eKqQUuDQkdBUbsbP0k3f9Xy50pMRPnNnDVH0Bg/zhV4tCND8H6WRoDfZYMs1u6Y4uP
U7vDx/TpmOYiHiVXPLvP6LJJ7/SA41Q+w6SWFMaxp2QMaDjz/ixZVxPJ1RW33SWN9AmCtH8UhmML
dHiofOw6rXJMqbrFN6jSruAdJYXf2qBZQER15F80q743NxDa3FP67VIoyGL7+G2aqxdPoBeeQhzu
cNmRRzZWfGwkcm9GsrY8cNvw+/KMYJ+3Ejon5z4lyBXUz76T3g/FN9Pym6Q7plVlnxX6wD9R4xnL
p61PW6p1Ce+luO2D+HleDehVgBdbB9W8N/MyQCZAlGgSXoW+dytq6RJRh5zLyVcgcJjTTiwFt2eV
rhXz+sjU67SrY3JmdfXIZXWWNL2i51YaGSPUyF2xuI+g1+1FTzr8b7lQuXq+YmiHN44UUfbFagFt
drYQ1FpOdxE+qwDgMOTtGS+9r1FfXskrIfFAdWg4u/eq/YD49XOcTazNAUU94Lj7ASFI2T0d61+T
bOnRYfNbPMkGu+CzLTR+WanJ0SarKWjIW8iYPUQ0xFzGGVgpeZrX1DctVsSRa2NlzvCl0MBa4Rrj
7z6YzeJv6gNgS6Fv2b8lAEp1SuWI+LaV0GDDD0JwWeTKiMhT2uT8E1mztlFKE93uTZCGZA5BKeLY
wgC71noynNlb+N8mq1lnWbZbcZnqDKR9rYShrvzWj9ohN9wXDY4Dsms9ttbBFW++jH0WvK+NSmba
OtaiVNLn8ojUi5JBMy+0PPinSJFV6r22gZEfkA6FUAZ/IsANzsduwqVVsWTXn0bQ/hqiSN8Unkqa
LVk2OfeZFZ/6UvmRqaGVBjjjSdStBPbJmcRja31PJLowkr4Xew1eZTj3BS1B86OUY2YZnJishRgl
JHPqQ6Jx9dgZ1/o2sL0QvyL9s9tKWitZpa1CjqVg+jF6ZgAzFVlky7egrN0MfneF94apUDcDqmVg
5P+/tmskm0vw+uPD+i548vjJFypGwDFB3gfBmEpLiqiWCl+qTBDnHZNx8AU6MHh4e4pKhaxTVfm9
KPy0X1cqm+oTSDnF+57gLpMsI11NuBsxmAoKRbyeW6VbKYjNGfblWkZxI5fRn4r6oE8i02YuNd/a
MUR8QaqDiWrgDWaOZTuXtBR1rRsl5UPEuT/wgsnxnibpWbBDa57Q5CIOsMMJAXmoqkiFPtp14yxl
ARn1s8OvnuryWanBE/ikA+3N2BB15UMcoNTmsV9YJJwiVzWsb0Cv93jcP+PAS+UZJ5SbDc8sEZif
woefWhWj8w1AhcIjo1kI+E9b/QFkjBuETaiNWM29QBxddSlGOQHHN46OzyjrzQj5XJEEF303S01b
ClN0S2IbBP6KFBLu6d7riVMcI2oMmEVRwlXUmr+qVYnFmy3Wg7nOWE9xDXeD5MiVSbbPspBErE99
nT7mt5YQ31oAwOP2LTXosg7lAQQHwCLrv2z+f/yBB+KwkV9XlW2IHVtE3aRjSoH8sxI3VkFzTe3B
7dWmDsCjhZozFg8GWBbIEsufngX3fwGUzhAQD7mrZv4MErmaLpq1NrkoO+WBCazRfsehYz28nRVN
GpjWpKHWNP/NwrBR4mjPfCpQUEok2zcTRd8s2h0v062Zhf22LH9mdnn3ESq3llKnnXHroLj90tYF
HOT4vDMlZA2lD88Km3uZ9tvpz5SMB+XTFwceVvxVq5TjNrxkhNYyKxgZtWOFutQWcO7rfPnF01+D
WsdYpareHCwJdSl+hSEyJ0z0YkWsVjCnwvK0Dc0Upn579+PeJOlqIMnNASfOD1mXRCkEwvMJ1QT4
HTd1ia3P1YGWAJaSFjqddI22kH156H5XQ9vywmaAieZpzfF5pwZlIhmaElsz0pZ0/S6nR/M/lsq/
tzoXjQ0qnTVgtiwnepzQZLFnFAdIrKJRkE41YgUP5clXPhslVMIw20KoX8GCGJsTVw+/HJRSvFzO
7ZU5SMK8ObboL2c8GxJLZRHdvZXDOKxRinFWEScNQbAIrV3ooCeS/hlOpnZPn+5aFr+AT16GjD/x
/TqHoSRifFdD2w5mL8yB3Gi3hANKgxkgZSQlwAxrQqKFoFSVFQUKGEXu4llx5LNUNTj6pLU257eT
dLk0CjBMDeYtw0fOCGvoJDYFQIwm45Ev/PdN0tNTp06jQtbfrMwbdgXwzqNgaQYIxID9vgBzFQas
o+GPE1ersXKZD/EtMBlzpb/uuCL6SbuAamAt1GuVAPPzO++KBgLSjgDfVP/jkpZkP1jHF8kE44L6
jIXipaGHImlDWXkytR1yHozaBOJ5eF4HGK+eKszX2h0w2aqhXuhAJjsTJepEckzqrJFcW1zoRYjm
iWWj5TvzpQSlYP6O+LZxWRLicNuj67IzRmMiM8bBt5+hHzQl3Zp8h7NMGBniVcRdnLkyzNg5XQEq
nU17rSNyIEC5YdNgO5vaBv8spe90ldljCY2w7h7T+SzQQeOZJmaYI5NJwD8K4BpX2zNAtn8h28a6
od/lYJd668QNSZQ56Mt52vSL5uMyqG0w8b+HcSgEaUDped1KKrDLAISEF27yClPfv9sqGv27ytEU
uYSlTI8ejNCFyzRROfQq6FgnWN8LPRKuaZHJWfpZVDWr3VEt5HtRhP950i+7PNBuH+uXycGXRzR8
19xdWyJxqVKV+aOt7OXlSvK8129adfsuc5o0hm2lz4jTFzQE0ikAh+gDrcIYweSNwO4Rbl8Uk992
57vkLz2TbPoWLp9h9H99NeGdWlzJZvozbSXCzIB2P2DrLdFP83v4yKwb/M6AQo3AAWFdXEtW21Zc
wa+xGA63RHS++n/GHPHi05/HeqlNgX83GUHRZ88yB8TXI/DDmKeiGwkkT5R22vJtP80vEhYSSwl8
haSLvhsRed0VnYdE9WNMU5M268aFbsZ2Kvc/LGtMGh8M4WgvzAyVT9Lo2krNXSieXoa/bRVeWRMU
KRMwqUuvomPufDv/rC0QYE8w7xKbADcJ8yRfRqXZE9kUDkrKxIJcRZ1rP8UUtnb669dICvxhExWY
Qfo8hnKLMJXfHtHy9PdWQk44mr8MflcU9+buV+72NzdNFtbQ/I4K/Uas0GxSX3bD+o6Q6z6WglNj
wZUrKHREN/H6k8zuGj0EJqYfhy8gL2PJcdf93zhkN+LMMS6fG9BMBP/lakIXQIdbUnYUlPGaW2A/
frYD7xwk5HuVUlFVDLcpVbvIqNIcq6PCjl5LeNPVdDq0GrafKoylLuucfifuYwpGuxLe9ol+YE8X
mI2CDUfGYlHHWThgDCcHFianawzjaire6ze+v7tIuiB1DZX44rAdb4P9Pp6pDIjfwfdx3rBsFOWl
1xvpIPqZwcGf7uJ7ErrbnTZqnICAIgdZed7glMEWJ2Zn4glq0pSO7LHUr22G5CIp5OAZkiFC7Z9f
0UZAAz1rKXU5Fj1LOuGIVDGCnBNtQlVxk9kbV2EIR5tLdr6IPePKD2OpZzX67kXezba0bjNoR3/7
OjNTECagIdb/9lqILmzndPMZouD9ylUPCF0ujjaTl8goazvEUyoNqRKBeDIwQHO1B4uUhaJgqsKa
175/cqBHWFCHmLMiv6jx5fisJJ5GvX8b6EcQyK9ILrb2vknNgmkEpTVfd/zXC2qnN9wKbksI5BXM
p8XUk48zulXjQfi6NxfcH0nrwwPjevkMmoQYQdCYA4TRZ5F5/LOYuIXGQrK9RRHEu5SqG+A4lbD1
BlsXwclTflpqDC/PqJq1OvmrAPdwcbAMrXfEuAnOEtC2Rrq5qlhD86LczIwVRPQVXJ05qYWP1quq
CO/I8BAYt27QjzEGrgdEELbeKZ2kyFEaf3NM84YqPcuEcjEQEQ1Nz0OdDVGrZiwcnhhbmq+3tDqO
l4M8OVzvXq6Mvw0w1bh6pgV8mTXhEzSoXktiafU7ew/qQ+xCWKod6/WY0e7N0NkXMvkOYNdJXF45
EZDLflRgD/NIeLPyTpzDwc2MImPP+tJ6HEGQFRHoEB7Me2dkjYpkYRLCfgGT0nrcw+7ePsGrSUuB
60ZXy41bVX7oWvV8SESieVU/IDu/7KF5j8Dc6gUZDJKO4kI0V9bdQIleA3RNhXEEVZZLaVNympt0
idQwJxLdgAtgnyVEgssMsVWFsW8F5MWcRj35egRiLndSZYTWZEWNH4OFmrXr1GIZzScY85nzQkaG
Vfp57CEd/0UU+eaEdl0hd4AMrlYQ/oBRbW4U1q/2QbjnDnYzkzC0TJUZgHgRw0YWnQlZJC2g3z3U
ttqfZ8GGtDEGNhR4djvLO1hR6KbA/ThXd8WNuNGQEvtbqZ0jYttoRZ9JHeuwovbb7nLrTwDPkqtx
90MkuLdLetAKEndHyqdvRDSrBjJ2DTg6stPRz3RNqTvyk3W3sszdbEIxg8XInJ8pMAUc39i2Lplj
TmgZyuSFDPfdzi22J7CpRTbr94QuNHACZ/KQCAb3ZaamKhYWiPpL87TQ118GhpDrrTn+Xb7R9iet
XIjZtmtnrCk5OnZOh+tSJTdQdVV2o/XhH325t8WHKbEpPjtVq5eybEc2T74celccRHkI5fmA2DvH
V40ukVTtH3VqbIGoLUghkvS70HUHOslcss3kkPxYz43VV1mfzzRuy0KI1xe31PPd8/ax5Q045mjZ
8TvsmB4OGcBg5UfRYoe1Zh+nxBd+UAEex0jZP8Sc0nMxIqqA4ONv9W2Rr8b1/+uFRdNTHVDOSz5m
3To4cu1pHdZP3FuechDhe4IkeVgobX0/H5G+bLWr6QGDKgOylqyjkGNCQxuXuQXYqSrAYZxnSrqZ
2tjWRM2UEfr706dP+r4/JDn6f7bQdHP1aKvXIvUztvbnUfLSNrdIbxtra/Fq89oUAn553BJhJvij
GFxNyRxiWKN/S1EyoLO/9WFpByVGnZgwgvLFNC5Q6rKQCqpmNIaN3VBYWh9aF72vWS3PMl5yqXZe
E4A9o92sjixCrhDdnc3aJZYd6QkiAmgiYtECz2wNAMKhvfLV3PSeNXNHzi5WGJ5XKIQE9rDK4xi1
B+/X2M8kswM4hJzyTJC5VpEpKoEUPC6WRdoHnJ6QTma2A1XllEXupLTjOL1PMBclkBnVNGLv321b
xuxt4M8dmnFS9+6eFgiA3jUIMJWvcCRUia6JeIhL03QdGaIEAEeOt6iitF+OFyeixSPCf2TdBAgY
cdi0c+vzJvnGKciruGccMs3lgOz9xAMbseM/tBcFk0ZwCNByswRVxgwRkrnoUAFp9+E7//029uyh
O/x/uwwBWE3ZtetbRErRouh9fBe3wYP4k9nxyUEqfndjkBpUqyGcmaiwYzYX5SX6fp8dXCUelT0r
vwoHUCsW99FKRU/TsMGTYRc/2RA9/1e+AlfJWEjkUGfXdhHq0VI+2MkpKM/knEcJgIgzNdf/pPXP
K/eygNGnTMhO1ZvoAu/cNEEhNqf/9QHXTbCtJYPBGF4/AE2YLkTb+D/PFfZW4WpGe9Wzfpwt2Fq0
6vetpCClcPlrhPZdFujjzt6eAbD2/dvnPAj88bAlzfhrcnaRrvTTPyIiqGQWFHjdaZGpYC6YL36C
/Xl4LjdMw8N+bP6Ju6xkztntrTWgzj6GqSOtB/XXfQdZABSFS1nnDDeKLRh/MCm0t+WB9pNjJ00s
hakk1g8pjN4KH8Bk+2HLC7CbFpdl6WBwsI+0FYl+bjIHmZBhB4k38duDn78MZf2B5DO4mSgvQvTJ
1tTXFtBvOV5TltXcLCw4iF3+NrefP4xIF32Xn0ftK1bUbzzkrOFC79MTl4j3Ksn33h4R0aGVacMm
02S12d83gJMeTU+THLJs/9Ay8GIc4ZNY23qsVwQ+nOPS7FajXRJ5RbQrQypRMGt/nFoLa52Z+60E
1YTDBU9dCZ98HrmCQ7z0FkKPPK+oxrwFoZ9y07PX/954qAbT8iWn71iqQXYTWgoLNvsqBs8H/dck
t+Wt1K4HcapZ4TunG0OZsIy8E4xSsm2umyiy9AVJVphyA6e+AmDeOdgOXNUMk1empfw7aYdbIc4a
eM1FJ7r2rYVssh7F9nX3+i3U7zrllOeq17q5x6P8d50XeNaljj1c2KzrdUbaEhcAMdEgQkZOUd/c
RjttM1i+Wq9dpWgSRDSxYu6vwxTZWrj2z/lw+kP3qnhsPMoQLqbgbMntBaXyo3vd5tIyMFQE5vgY
lhMlIz3Or8CSyRAfWZ20+hkSPuKgg5769fGmKSLUxNfGhIHb2ynbiMZPBf2owcq1l16F7Ah0+QCX
ZaOiYAEjcxqxYbpEhsu8uWF00sIFkIG52TToVJM7OWKnPKVbUQIijiRMe2NaQxl255VmmjQihVZ1
m2SFx1FnG6nlGyHT2Y96NY35UWdGTMdR/oxPnfHUDzqCYGIEH/nP7rMEizcKwd9FC41X0fRGBM+p
UTFVyC0GktZ1n8j2vkDjbS86AX7z/aFIyO0rjPDsoie0gQqXej+PEyi8hkzTWt/EE2fBGpFNsl96
AxQwdvucNPeKSqxFUgUutib+O+eIV8ArA5kEgcQIgvqwT8AJ3MgWGlKCv+qhKzvW864Ib4ajiDlJ
F29lkTGVF0s7YSabHV89txqMEMStzQOPTdlCqaP22XkXL2fEx6XQgRi29OPgaZLN0H7QBgBSL3S2
GAQ9WHmUaqJnGgOTsuD6FLcf4YKg+6PIs3xfKyRgGPyUaPljYz7V4EkZCR45W6JPuoQuYkxACM/e
6k7GS6KJdyJzTlQjXgtcD/Bs4AEGrZ74q/sfbSc5S8gX/jCE3p5wdzsPTBtcme0g5gVNWlxuEzn7
s8ARX45WA+JudxhnJ3j1MukS8fKmD7Q1LlSOq3wNShuKYcwi/RBYp4+0qE93ZglIRMpPFhbatgS0
30L68p5LVq3rccibCstn8SSEtkdSoBVjRwqt+Kyav0yKLsid+SxvT/Zj6wjh4f/BjFLAPN8xCy2R
nxxSqYUx8NeweHAgyIbhUVJEGlhyHJFhm3TFRgBJz9yEqQw6FrtN4xRl0iqmIPru6FPSfu4aC00c
tcja4U80LBgBlJFZVAI3OV5Di3ymdIuH2/0SwpbHYdV2NeEs+MVwpD3N12SAuSZckPClxArf3L4O
oAwZ2INvA/4HlFxxDYVj4JGM16FGa2/ASfb3Fpl4NqSuQ1XtQD5movu+TlFois8Wg5P3ud+DVJE9
bgmXdIwnV/3Q31kaz8ikZZOLbXcgyYIeRFb1z04+7UiSkpriBSh9y+QOp917vFy4303NDdcVIYd6
l5pB9RSujkBzHJ69xThBlqm2tjkKMkxDDZL3YPrWgII/r8xdQcJglyvh2KG5rpo3xiu5ZQ1uyUnW
6ntYdp+t0r1HXfRy6IzZYtWpQy/Ze8+K3zeDQYRrXbNmwr87mQM/t6lWqQ1jt9V22kqXX3Km/cKJ
96lnl8rdrO1Fi6bj0SDpyVJdoPbNIGh93/nndpmC6WcfGOGCWO1DQ/8SHWvtxhWu5RFr1805rbN9
GPucH/wMc7jREjNIJHbpm/K89xszO8kSfCG4UiqVK2GWnjE88qJQEs4wtjDZVzk/BwEqeVya1+ut
wT4XY6Jn5VGqdIWuH6kxsMD2uHA+iHHzVUaryumS+uHgDZzfG3PJwHoTAgps+lF1oRFiDEaG7d/e
n6QRSaoTU7ogKK2ZngnyXlEDZPUxkfDaU7UJvoEISFEd3To9PpBEA8ou18rSK/2/+K/J2gPI/oHL
SC9gO2uxO01ndvPuChTa/JtO6EVDJNke+WtVGGoY5d9FI/69hLjsgnXzmKZKd/qH+D5klNWNjzkd
ErD20mqpE8ox1drYbqeP6ezmKmPvUV6QxNR2IX+59pxR/K7G22aqCFPid0OZ5pSsrckmZaqszL45
bM/rkmp2mjOIIgysMVFOfCTmf2bPb5UYsifY4VXkDEsQKMptCj9ctuwhMK6EA6hcfWHaqpinKrfx
0KJl0wGIGKL9vOJoW+RgYVcbA+zoiJh1llCXDv/o0ViuJODgQcqys2zuxYgL7yDbXK/IOIxSxW3I
pjxLWxZSiY07z1fOY3qUPhCo3exHNYb1kNbQ4XfgKqkmcMv028Ndt3OAJ3sxBLC/0Y9o4Nm2FcaP
+VBjHBwDqWYPVcqaG+NtyW0mYPc6NFZO0m1S3mOGNtNAE6Aj5siNqYLXBp4vKzcuZUwY6ttqqrUx
dx8gZwpKzq/14ci/Lh+a37sAMZ4SdIaiFfrRZRAQKPcsqxlTR9skQK1srRPFkB+0kEMspX6o9PC5
Ek/a8dylPtXHQFkhSqg1y2YcmmEN9w7qdIVjV2ZU9nRKSkrJODVBVeT3YqL9k4Ab8so9Vt2R+TBh
liH1dOuoXLam8WtYEseUqWe4AEfWLTG27h7KgsCf5yoUuNiEq5HtpsmInflGv0WXzscj3VoqmxEW
eY5bKUqGOBvqInkRdm/dDuUWYQTi+4FxVMKn8KnjtLeSio9fRJ8VhoUHd5kiQzMdq10ZseVbVJWE
99ykZhjYWFjOeu9M1D5Z/jJ+M+MsnG47oNLV7UdMOrULL5mvoZ5vgNsrMTHRJS0MLbeyaeMG4pmP
Sqq363BdsK2p5Wxt64CLy4J7keBlava3Gqna2xQM1LUZjfHb2eH8NIcgdjOXu5Y7pczIjvkjy0K8
AkNVe9vFsiBOh4raluvxRHNCokCzFH8ueqh8IhasJAOVFOMWzIxbuYxDk/0MXst7DzFx46Sxkyr3
fWGWV5i3uOQl7VJXi8G4lGDAZnN92xOM3JFmN3RXTjL8izrZlWU8/3oxjhzTvBE6zfRt+VV/jjpt
JLjxxmZ4DuTcFvueO6e/ha5R7ct05yxCaYPeot1NqMR+0lUaA/wKqZpS6A6PqL1a4H/fij4mxTQb
RXanv+E/azA41acNib5PX3h0QPBhjjggyja5oflPRjN5GDCoy9cDPGzgYX3EntRr2ljoXM6gfgfR
eFaoyRkGdHPTY/qHEoGEIDGMSGgQRujMyEqAJ0rma9ht0JlgHKuB47vDQtCHE/NiD2wwN7UJFyI4
fz8TZuJbdjc0ycSWJk+uLMLuWVedjrdNCOoQhu5yjDZ1qQAuemYAotIJD5C9RnQdn8KdP7RTDNdj
tTiyoxUXAqRMzMbvw9rbA8jLCvqi4yXBF+HV7RJycpEUczcU4+DP1/WeXm8NI2O4y/1+BxUnw4K6
AuUsj5ZFkKzO297Bv7kbhtEZurj/9xdZ5jfvFlDSMuSY93GN8LeZ5+r0WNRxs5BJhnxFeQ68p3Xr
qRkS5vQ+cQ0822fBXnXh45FV5OTygvefZsTqeLXhZkU62NoNIivQmKPw7deUQhF6UlQOnZOZ/VfB
vHwbUxgw26JviS2g0SEEyCNjI48ClM6w/2qvkrRYoRLHhqkHTn8s6qkFsa+Ou37pSfWKPqoQxhLs
Z9/hu6ZRRqb6Wcys2mRjCjE38qWabU2n5hIVXILvT0ABrNJtKffVKYQHrcv0WcZJUwxe0HNh92cM
ANCTg4u4fhREMgzE6jm6LoQgAWS+ritl1B5/bImgVz4UbHtaC1be8n6LSHXTkarvY66VOC4MHsI+
FUqa+f+23CqM9i5+hrJnbBqNwpWGJXyaMYfzFXmitZlomuxKvkEWR2o/453tZmFvOWiCT2eMo2LH
hQJZiBpWgH0QgSFowdEay++l9+sfIaO6L9CkfTh/HLPa6dKNGjKIHN7j7lwFH6Y8POZ3DriuLn5a
L3mfEnkO3+lY8lrDvdWdwzoRkSCg6frO79sGi8uVRQ5Lr9Jdv9JxDkkMUpdBRxTZfteFdngmYJle
YSlaF0yRGvQ9nkS3k0NhY+LhAh/SDp4ovNsdpeFNEQ62ZhrptbUzC07MLsY9pmO/T2ieobYJ8iW9
K/kCM22DLLLIMwhCp+8ii5K4z3Co0u8veXhxGjYdGWvFOy0ajsrMZFE9KLeTLBiPr0DOysqBHReL
ygCy1hrMg077ZGCgiXwMwNKsL6CyVloUhyb/okiZoM3q/OHeshVs14n09HTckyQUk4B0aiH+Bd3G
FgCDrbZABAaqhqr3PwvAn7iqlR1mJgkSGw6eZzq4bhuwQY+iaTF3uzedgFsIJHsNezNZ4JS9OTnN
JnpuE2udgHTXGmAsEVv5hlo1ayNkrnnQTTJIs8LjVi4x7VLq/jMN7shPwdYIqcNUOEXUbxprHVHS
5bN0VMgauWUeJiyowyhhpB14ZLEi2qQq+VriDOQx/WUIH5BIjsb6D3D1gXQib1GqiWZG3wOCpXl0
rWfzEKXQVxeR1X3/XJCqvVC89k80qsEX5Q2SIDjOlA3hl2WlEDLZ1Jq6VINIM92dWvCHhY8jc2bW
PECYOIZJ9YviqpDz0iY89J+xcws6bJ9UzT3Z15lJS1tYzRVFzvHVseDHp+Jy2LeEKAK9cd67F5dK
+fOdpW+z4GimYTtnn/dGOrFIqKaryquaw6YojtRfs7rCN8uZJQs1F7F4fjImEQXtMJ1raMh+Ew5Z
ZRjAqa4WCCTzG6vMrP/e96vX6RXNmh/dEP1eAc1E95ZNSV+3wxVuCoq+crEqBptxa0IqReHp/FCu
lh5jkhBBqg0IYST6HqNbZmaUjKmGY4UM1w0vO3GFGPmeaNindaaKx2P9xvKK8rLYYEjA9KHE1Hfm
dOMPbQawau9HzIBrbPWqeZ+1zB2mdyffpDnJ34vcT2LeWz56JW4yHl2YXq2uC5SJGORNbuRKnd4F
1VztvFExHCG0t/c/1IJSXIXJiI8vtIm12a3R03DVYU8Tl7ma4FL1SOPW8/XxXGoP6M0AAlIaGQA1
ybF8iVV12ZZ9CPnz/dlHGm8VQkaILNMfVHGEQBU/AiED06VzGaTdtx9jItIZqfvfx/M4xcH1ktcy
YO63nzlS8Mfse7ISrW78wlWyyEIS27y15rR6BNQmdxVl6pRKDTBIQp4n05dnTA7bwMRt6vPbeOdX
YErJJe1RpMK2pQl0YS4ohuRp19btBa1TcLltNMr1gBDZKxHb80H0CEK2h2u/J0nhfysA9A0Nhw3u
MXlEbyUsI+MdrNiqwsnWxSXd+8vV0bzNwEi0fDzkVtTs9ixN05qNyWCQJn+hZ//ZjCDhJ4cM8IrJ
Aa+j6kDzJ1ncDrRzWB/jkePbkSgNE4MnRoxanymhLqXuad/Vg15YbTXzJZVGdOxsBl70NHAebtLO
Sre6ghGCXqVwR9QZ624jeLFJr/i9O/7aKpteh0q8+9DzA2nGak4iyHRhkQhnEjT74W3+bMbpj8eI
7ElzJFa9tp1NqNwr7wZC7qm5BtGFQp+saJAy/v9BoMrPBTyj3Fg4tj2AyYjsFHHZkqZ2hqfxUMCV
wMYvH+CmefVK1kJXtG6ciwgx7oVGR8dlPwqQWykIGOOo0kNqEZbV3KkptGwCbwW3869iMZD1Ie6G
Ez+kzL+hSpqs+rEMQ6WlhJQxly7PNaqL5/mU2elADK3/2xPow+kXnBoZtpRjE02Qb2OnL6vkPIXn
RmHRH7RWF1SBM6dWgbZjJFkCoa47XPUtyNDBvIwTxFe4dB0N9SVmX0zMT5LmF4HcY0oKz1mJgXpu
lX17c/x99JIB+CWMip6pQoY43g8VpdN4MrQ3jHNCE8JG/kl41klnGZcpKOeCUvd349kI/lEptGf7
AK8D6Lzur3M3dEMMqJ4YJF5Fg8kNtFwmPTQsflqpHXTk7YZJtrLbUNbqJoDHXAmqsPVemBdxNCva
KDJe/EvqLOTbsOUDMxCoBqMhl4wfuLOSwE7wqjjwhykDAi0fs4E7pJz0s2ohe0s/PFzGUKiB7c8o
NdCDIS01k9FvN3VGkiJZCUEfalbRQ5r9+YSKaqwLcHRB/c8vtd3LjlNF7MRhsl7wyq1IG1RbJUZ6
CesKgdESbYw+VkhX39za3+DSpt780EZTY8SOEaPPVXu6gLK444hLstXW8lNfKWWzrWs5THySivTF
Q/AgQhQTJyWMz/VcVyWLg/upVnJ4NUNtuZnF8gjDwiBJzZ3okTuDdkuiZNBfv4Tx5LTqxnWEAQw+
TYDJIR531NXnPtFADOfx2/6Yn79tu5bOl/sQH5XDS1lqFuCyM4RK9Kuo2P6MEZrXVIFDMxcb93lq
5wv5LX3U4lkqKu5f5Ef8FFHQnhBgPPmaHqBcndHBfDCGRr9QxRi3xZpOWxRFf4wTf6JjNXBhShbL
w3n9hEy87pdK6bd7y7l6E4pm9HY6+gBiKU9MZC5kGY1nkjnqYKivuEQA3sXvbpBQFsGOBHjo+8Gm
I9Mikw/xFt5lFXmF1iO9EniIBWHvsiBjl5Bu3VAy8ACR3S8cDK50YiLvyWCLFQUdpqRqHhRoNOOc
964TusdT/IR62BUN2UxCZWgpu3L0++1AvZ5TUIUoXB8VDgNuD4lo+IQuYuPg1h5gqUiBqJ0MLhfk
zb1n2OdABKQh76+bGYuQz427cBO5lQM+fYzMveFal6I6Ss1O6igBeiBwtCQiD1MAvxzVimh2lq2n
TDccwiN8/OK0TPkjVinXIR0/4lKTPNNcwC6yuQ7FVmiccKMX2FEBpJRte0gQB3UqH0tAf2gqvrhy
jG7Cc8cdbzkSEfXBE3YCwbHYF3UtMXlE+JqVsgOmb+lyskFo/m05Mj+/kZjJ3quMm28ORPfalGGG
xqQRz9eo3nU10sOnKN0N8mjuUnawWNBt6YikI71xGKvggQn5wqRQcHPdK1c0/4YzqHM5YzNpIvW5
RL0Ym/WV6y+xvB7acPc7jWIlt/ZvMofcGWhxqRgTMGSMDtsT0GADMci11+Y04g1C2oan4iqBs1gN
Uyuzd7Eq4ETUbYe2AHLqUiWpdvxxNKlQPlV9HKd76WRPa+QCNuPMllfEJ66gQVCPWTxmZZabu19W
oWtzJghBiZaWmg94Z/jLW5/bRmR7caLbNtycy2Y3wPqvOr2gS4zJOr21JNDWgcZxJQ9e4NbM0Kww
C7Sx5tMxKQ+icaBJB+KskCViMUfqLmsKUFS9CFWn7fOrL68+/7wEceafzFCrDeZsIJlYIilbtqOK
DCLqDK1DUpVUDN6Fyv3RZXWPUO1hhC/LSdgNo1SibMMxCwJY8Bz6lSNr0gUNtj64Qh5KKF5P7KtH
u2wld8cc7hqQvUH81eui6i/ONZdqpoy71okIh27qfb+wRhfTpa0G1LcrFNxWdQdua+NYf5jrfKVM
tOl7JC2G7Kysl8vcc000eNbFfUEZAOr4VmddsQ/6G8+Xkuo9B6HpJgHlWta42+z3dZtzqotvoxZK
N3e9I2VjJVEdKERpRqPt2m/A1BvuyDdppRrDiE545FgKLZ18H1fniuFoXVPjstmtM5XDhzrAzhTx
BHxX3bV3qUlED56oRIpPRI6PScWUyJu9ZZ7FTJalfuN1fg19Z2XFwYAA+8TDXwkgE4Jf7IEO0p6g
UdsKns0C7WgaNUh5mvIp98T+rve7H0Nvfi2WnVA3h4cO2L6KtLJmaCO5veYJeaUuWBlOniFpsLmK
/0zQ9E5bvaGR2X7yL4PUbFAwm5v2m03q1NH7fGVWC4hsGbD9h4JukXAN+VFMobSN0F33VJWq/zJm
r8NKKTDIAFxuvJrE2xkCt0ZfBdKuiuCgPZ6vbeNneFqizp4Qu3q7uLFB/eX4hDbTeMn1fLm107FL
4hHHlPefnMtVlRX84B+WVj6xsYW+irkGt55HMvy9VP3q+buwEh6dwbdCuhlHIe/8BqYeJF0xl1Rb
On9453DDcJiVtnOr6ElvJOjbStzXOZh5Ru0SvxMg/DlyiSwu1NFQpRkhaRpmjrfYbFKwG9YZ7PIP
IDqZ2Kk7qe4+GIQwjyMPUsKqCmFF4Ss10xDOhUoB01OKxj75qXlAuc8L0kfi6ledk1R7K82XmHUP
rtnTz59UYWB3Q9D9XrQ0muxFpjip1aLZ5EF3wgR3uwQMC+asQzKZsDiiMKcGm1E0Y/aI9IPQg3oU
JCP+cFh3gCq3usL769uAOz5b1x9AAqcYtI5JeJCJ7vIoBMFL8X3/aB7JyXx8XccotQUJNlDt4DFt
RbPolCRxzblQDiCrVQBw4SyKdiqKafrSslURtL1d+UjuTTcz6bbhwPH8wHFTGsD7r0q/L1wLZK6p
Cc5oopXcPWmiDAt160wWcgtH9mZ/wtIgcG/ZtnHrVc2xNbML0Br8e1hWsyO3tjkhShIWnabMHoAn
m/WXKyL9S2uu5sm7q4y7X4Eb8d/aULIwBlqL0G1Lg8gqm+B2H6v5BOg56nQmjO0u+z688oXRGTBq
imrdMDc4dupnUTu0OkVlpnXX3qyMh1IzsQd7y8lZhSeyEoH6z7jfpED4x+ijneOc+s2he9ykRB0U
vrcRhJgWatXxsfEuXA46p3LJxYwBe4j5tBB2+CuIEtRkkoWEVE5Uw0oY/jXwUKxRJpNHpUp+ePRa
Hqk9C9ZQDRrzyEX0vgcIg0Lg2Mx5Gq2uXDpPBSIvNahh1oxZwTLEWQpCbAnDulQgnOMlNFDjt7CL
Ls1cVS7mDdVysMIHMdBGHZK6d0reZmmFeXafhWRYLtTYJHZMot/3ys9QYniXCQcBJfnWTiOLUGWR
q85kqaYB/e95Zr+vnBuMVU2+30p1G+d3AmwP99zIjsWiS3tY+99vVhie5PQr7vInCYL+9UbCYl8E
iWom3iYi8ynUM4WuB5mtT6MdiLduvPYuUQzU717DhdV/7OmewKblIr8imG4hif/bFXL51bjeVtgi
O0kUEbYltD2a5VSK4Lz74HGu0v5hmLPDz7iQfgMtutohAejzhNPWDEHVVzT69fjlmiXJ2Mr7fXfr
nBaQqzec2EUD+xAhlBB1wqA1F/mobNbP0oCSQdTdCB8nf0h/ZHoJjtQ631AfiQ86/BasAL3MDA9V
+Wo4AbRxqjp9SWpLF8FNF0rgl1xkSifm1Xzb8BD3kAxHVF1z9MQZ2bBIx2kmXir0HuvQNpgW5Sys
HyK6Gw8d9cgx8Prs8PkYUGhZLdpVgGXL0LOFq/V0uG0iCWVRa/hCjNiysTZdupBJKNU1kgkFJ5jN
/lS7f6nLViSHc2JsIjggvBNIEXTx/TjuyrqQt6fsGRkDDDaURyoORkXdReISB7C+nnZs1qyemcN9
6rPgP1U1F6+ziNuCX3sE7EPmCb7m1GEVH4CAY6QQhOgg4Q0bCeM3kIRmfrbjUpdJYhKT/79VtG0+
I3OD8b6KBWPag0wV9DuFjyuM+6Amp+ABvSsOnAul8nKa9QVCXlyxB+ZIsr6FRXKJUNk3tEuINqyP
8c8czK8emLgSqBZQRiAPYjbyDO829/GgtFvmW2MUBW29eZtlR0bKayFhEtKba1gzYQBrs6eoA6uL
rHKLLRep1yeNmDw5qvPGh9fCSvXH0STYMeh/3BOrGU2LOJBexq+eH7pOY6Sg0OjAer+xetgEhunZ
T4aeMMJvpP8PX/0E/rzFsnQjaFKjrsZDoD1SJh2kJLb62d3WFvkhJIp3QgtATyrzQNOK+8T1NvHd
alPRIG7LJv+dpXNKDogGapUVXJo85V+xetO7Gd/xwTfoGCN7R0VNCAt91jONdnYg4HKDEn/GlO03
Y5JlEvsFtYDJ4CVrySK1Xi8IWwcqhPLj5xB0OK2Bfcy0h52cha+cSbH07C3ncTNWbLLJMqhxl5f+
TyS7YAW6m2yh5G0J7dnUZK5C2yeWMFeqv33qqNbK57VSSohqdX2+65Pq18Gr2cq7d7xPVe92QSik
RLl/PFZwu8RabN8WlKa+HIXl5LSEh9XhGxQSsBZF4BgYoAY1acj5vbn+6QNhumi/jDU3i/4SPbPM
ps1q5hKHvOx76reZwBn6R52T2PcxyAICYdKjxKAAPBzmrKYZu5ZWQQ8mr9svgX4c8WtBJkdIt5uy
E0oApUSMBwzLQ6lgDc1moxwUaBH5t3Wa7amu1A5nydo1F+XGehYHP2yMi2GKX8jSGMHYjJeexPH4
n4ZVY7TfF8SHsFs86Wf7HTjm79EYcGj+HVMuAs1KKt9ikIozbKKXOoVPSmWKb7gxV1ii6b4ACDMJ
ZHOWy6w+0zUTQNxYYq+k4y4lOugaXs/VMQdbZFlQml8etZqFexClR8Jd4HnqmF4vgjp0t5ItFK/z
eloLShNI/VbK9mg/DATsCx3iezHx+Bm0PYPnQQFQA76eQkuG3+MR9UxPDBT3kPk5VP1b4X8De5+t
atLwc+wcWS2sS3BhE7JcS2+IwiVJI8qbjtsYP2dHeFcw5M0JfKSlenhu2WHCAWB5UgBdbM1hOeOO
vtOsYnmTl3rjT6T54FBRBbTMhnfWQXZmKkTAf+sG+qAJM6k8pPrDgmA7tEUc0gEgNvE4VYyKdAns
q8jLHoRwBD3wFTJyBO5kUgBo04M9kYwPysOsxb+cvDJNDJFKxSbPwqQaLkvuhHG5NsKePWzjPn5z
ejeJ0U3H4waS87+FrG+WKlcubfhzdMrS69pPQCIqy6uX+DXPL8XvAkW1C5BlPbR6FBw/pQFwWWdc
36EhJrX87gAiVqr5NZI4LntJlASebio9k+e+ly0PnPENV5l0TTaXaiZYTgS5+vcpqnfDri3AW/d8
trqsE8gKVHdO5GkoQ6yUjuzvBCkAuBhY8G+f1CfSS+gwRwMCRXna1Q68aIICjoFKylNiHfvZCTiH
bg3QW/K+Sq8uEa34Tte9MEQP3VikJKmFgypwHHTpdujvCxR8vmvCS+BoFeV4OoAWwglypNirxz9L
07m3kS1XKbyUvu9i55xicFDUKybvT2IL/Y2RDCK6f/+e4qwLezLWJmBiruzRqIS/SVlDGaI1gSDw
HOfJfQGpGhTpz8Q72GK8Qoj9Tti5x/3hB4PxkYIS2abQ5pl7ACbAfyLCe1P2s5y90puZRa7T/OYE
PVBQQubstRCzAvsFFTDcBSVlDJcivZO1b+2eAIaiu8J0K98A6OlaNsRUWlBeTA0r4qRrQY6Yq/tJ
zIzf9TTOt65yA+aDaVclDmglqjJ7EpbacsGDaiMeM+Uy0ZJ2O4XvN8CeqQGzIbOxU0n3d/MA0MVR
u9O33ZgFvi2MrZl8lRzCwsxBxVIME6Kznjc3lNHbewTzOi3nKbI1UlyZJre6EYa6XN/hAWWzoHof
GPQA6heuR2DlnxFLsgIJe2ITJcK5tvW96eCuLIIOQfLFtMr1aFfsGYQoq0C6swbi3lAevZDp7MEU
WnY3jEIiHTUosrFUWLWXHXdNWFjtLHxyxg5pHDmslMJv9mUwaqcknGc6z902NlLRSncdBEyvscjq
ouTjWRWH2MDyfbWTHKupvGys6PPcIFB1bhPXPT6pnx/SuUPt2ii8sYD/EshIbozC2ZziEbSWOsWA
NxUakBzeXYNK4/+1Jv3fQooBod3Gr9RNqQcHRz6ueBh2boaHelMI9xdkQVfb4i415SbyGh94VrPb
9XeQEOVAGTy2FB9PN9wXLfx/gul8U1KGWVw9rPaab2hWbennce5092L0u4t2YXOQhj8Y3hjZ9UYF
QuI269qtMa4dup9mPkYaob7moICENmMuCe6F1janFgFP9Xxy6KsQDHzgU+ahMCgxXCtcZTh6nWYr
lH11FtbxnkY4BMsf1yzIjyOoFLCBbMgSqYQ2iWWg1pcGFOVfrD+a2uqZXcrjcD5Dmwy6vacfavRI
aC6hy39K48U3N2btjbiHzBvW8L+Q0jIy6uprvfSmZwLfnds0LyfsjJWn8KBg5mHnYJJnkm/v8dns
6lNuPBqyPylbxIJXpMCzUzAqj19K99KlWoMS9cPIyGBRSqxehAHOi7q5dH0Pzv3wdpOMH6QNqad8
hxI9dY5sx7IeI3Q8nuWM6SlzoN+QP0Da3ATParvnDAL3a1A/rkBjs7LaJHRJbLRRiQ0UCAzevReE
HMDsjrZnDJher/adssMXntgHZhRZ61RCkrqQ7IY8FwMZyIKrTtZsbuFeZLS5CV2x+1Fz1QLygZ91
x3ud39CTfZ25P72ZGZI+MRCps3Y54LInFceFkXlGglHAwucbmqkrncwOs2XGzSSwYyBSPseYYVJW
Z+2PSziBwzh7YeCcaFSzzNRgP6a2CYeNoXlMuUrjqTcEV8EXeFPQjKyBQM/LL7DJiKkxS4yG60mA
maCqyK6BPZhaiFypAHQJv8n+k910AZJGL35OwysjzA/w7XsM1Qd+oShSjDCTMZjTbQ6v2iGLQp/P
h9cUpz0V/2BprLQc/RpIdpQqdxkMnvUYjYcS2AnDFN4Pt+2GBRloheAajJNTsk41CZBAzdRz8iq3
9XrW3xiW03B2ylg4zBXiKzdhCiahpGnHtDoT3WaFhhj9cURsT1GGs01tIPlJdWPBtqYC+VVs2FPn
wWPk07gMMM6m+RrnQn9ieWv84iGAkmCloO9By/N7o04ZxGoKKb5Pcw/yMYPoypeu05k50QwyDOaf
I34CUfu+MUnIAs1sPU27BJvyFS+CKOCDzdJAmVBYEXr94Uy5Jv58+dC0+Scd+7TcvCBrobr1qT19
oolVANceYh4xc4F3FNv6nxBrLg3QTKqRk9G9V14M/4ozQ8Nqf6p0Mf/N3aJsrGKotY5W01mOUt2G
oSqOrxpP6EHt+QuWXzr9EUkX5xmyIX7Ar5kqVqTERJMstVFGGK2G4I64i4N3tsGucm1QsfCZCOKu
w9CbIqpGvxtr6H/+aUQdilexVWwjndQYUjNCCd/UKxiILxk0cYtvKDrZ8I+9NMOTYzuf/7TxaXRt
ER3DS3RM2wIru0mb9CbZGJeEoax6nKE7mlRxrNP/9xB23w71eOPISczzipTNXxlsx/nVx5KEvg34
42g4yodfgM4RWJTFO0/NDe4jEz1eE0l6gWWBAPcZaF8W1oFGA4QEgI+1F77c3RnPYnWxSLZnzyKJ
D1rOxdgmBZluNT2EUocOzaNHqWRqsA8Q2zYlKQ/fRoFG/3G77jFhIGcAdh4xuraIWxBmXbSFRTOn
FUPl0Zc14SkhgFnR0drHQFTlIyVX/P5fCeKYK86TG++hxzGulYOBp+AsjJjQlGcy/6FF64xDtSkd
nJHXomsxZ+EJUJ1iWakBifPgdOSYWwG4hpbe0cw6AU/4GYagcdDy5GxiyUZS1mFbdfkth6tuYglt
zD1Yaw/lpwBn9c1GzJYVnMTJ233yPOrxa20jBLJDpyT4KW+g7Wxi352YDLJ+1M7dJ98z88TBvKB9
LoenIeMsfnA0lQl8SYo7aaPzZYafsjT7E7Y1Jj8ENPiB1B7YoLDIzDRPy145NHh5CCEdYTc2tKfU
9m9d5d5r0CYtw9ZBW50zkmUPW6QGzXpGbTBhFcvlQKCKv21UQQ0JLld+K7S0kkg1SXp55xQnaiVO
q8iC4E4apk4Gwc2kDnqaPyFmdTl9sG+dAyeDmH1jLROxe8KKhDW8+VkNmU03hNzpxAa+99v0NZmS
5Fv6V9LTSv5x3BznJcJsCEX76IVtJy7Saj0ASIQ5O+6DB1gfQceaG2jnpKpspwymqlKe4kkPlBZu
1DZRv7r8TCeP0alCpCvfcoCn7d7cBKRZimFIVxYxK0lfkMHMBdUFFYIh+un1bJpP5WQ3S96A1Fh1
wrBbMkmhS8CgDtB35ObJ91lXrVN8ZXyO6ay+TcPe6UtRZqtoOFIt6RD/TCYhNXpTyls4HndAAXBv
q7eCi+VnwZ6oHyTujNU+cYYjpVwdvLEeioQgoAlCOtVkDVDyA/LieHkJUw+Omx3ERsco5q7bfPqz
xfxIp5Gpx61oTCdlABrGqfgGwSQ5fCJ8dl3oM8FQBd+jnUvX1vBRrICrDef1ytV6ufdjj74bkc7O
qSBSQvQu7+JV0AC1WklzuMEMVGqg11irlVS0vn3p4OFmhBX7mcYup5nsdLcQtyZhDELB5PupIoC0
jH5rPCMOJSBnDTj6pKidcnvQSND2qW7UvygAsAeOoHUUzyhtJjnmi9xZIQo8JwtTgj5Dm/+MSJPm
9yqlUwqzcGM9Gj8m+O70liFXEiSnoc4kdYm1s4Utr0+UkzXkYmirdfo8Am8x7AzPNTuU61B+CO0i
4dOZm6jASiZGX2c9sQC0HNWz+yb3T/U0xXp+1vIPKk8/YzEwLQS4kiiHPLmQ6eVU0uSmlisE056S
HUPmwPi8lcpNEAIBhcRkcpP4Ki6dwcRKSsIipWw15T5vQhjfNRIDKibwV0q7wNN/v+ZUgXUt6a73
bGElFewkK+T1hRUaRGG+x/W3zodMX21IgcZfoRDkSnLFYAUEMl9Vrgm2D3+aBOIJJQm9GECW89v6
nXu7XN3QI8sKukSro9OIOFeFvYDWQShQhiWJQYZyahMTZzLHFpU2AkqTgjIj5OUQxs3Sk7/ZeYup
2YqTK2+d7UixLWJKdbO5YZGGMopd2vBUqxCnfr4kIWCNBE5YVKvEFaybA8M8CbyaGEcWYhkRs/re
F6InANjYTIxJ4xHWccFrDiQvUZLFiBtkY5ccqCq0j6ltVHPf/r/EaB5O9DYsgK35J1HFGS6OUOo8
CnRKhoZEqkpCVCDgv+yuda3Ozf4fkIKDhNTSezCUwPZgC6RaOEhruopX0RT9FRfksO8+jxBYEwki
IsBp9Fm4Lopv/WcrNhSqz3GcMPYF94XxwYjG9Mv2BuFTp3JgGDFDPE0el36vB1bKdnewv6Cou1bj
xrUfcFMCvNlRRzROFunR25z9ysIz8keZCBrLlnCaKsTlQ7wpz+afpDq7OuYh2lHHr6KSL//GxNk0
tVVA+xnKN4UBggy6kJbD1mttAfLWUt1uloHc74+B64XYcW1ByOBz+PVxshap+Ir0T/uKVtaPrQe7
qc9uuwJIHN82Qgq1Dl3T1E9BbHpVTk4mIcf3p1X/+pK6uNhz7s29Brv0BNSA5jdrix0Bz07BUU8O
at3n4susUpOvYCUdOD/RkRFs3QGk1qNcvanalBahI6n1kWO3AvlG2kveGtkHMyH9j7IkzVpp2r17
Gv1/clcTyeAyxAFfqHMa7ANIY6DCXWrkkv/VbdfU8XoehpdRxe8zXFJixQzmUttI6S0YRVqwx/Vt
tjROdsVqT7Sme1fL0aZzImtfBL0DALjHF7RKL7rXN/JXCPANBjSfalbr0MwJnrThw2ktUzVnxD1g
uoWrwr+MPgM/VFSRrFCBahJk3BCwbUH2MICcKGsgvTmdIaRmx116IpTMz+iKuGhYfjR+0Iwq62nG
IHlOJONMk1PPZUlAI31A07CYtEYL+qtcaUBVyOyQnpo62xYYW6iNvd/TyTOsU3GLcvzOZILvsBf2
/U5Ix8aIPrsIYc2NvcDId/PlIGAFVA04FFSNMHspG8U8e4wX4tje80BpnT81ZxFlsBFcq+yAwcPS
lMZMG28oIkt5qta4QxZCpy+9F1nJl22ZmgWxEDIeS9v683OgaPFxbx1oUSAC8HWTpIZjtNBa13Zc
E/JT3it5F0Vr9DYPLnKkp1IBQ6Rmrx8RTt8CLE2rj5CShNkxE1YG4F/acNR1ZWLDatA2aUSu3aNx
lAhnu1WeOvKEMj2+5fQJya2ssYVqmdD6p8EVsBPN1L+8PY7LmlkEW2Mwdts3aTr3FNv7ZGS+fQgx
uR7wEjKEM/Ll2pbpLVDIKmgfa1nwFHEKuon0ZwoO5FXDPTAy4/V+16JQHKUZz1YM6BNdvWb+kZ+1
VUXi9krnPW6G/cL0YJRjyKXg+cn6qKX+pu3ZiM6oGw2F5fWKk+ExTY/fUuq/mTHVGIU9gIJGx9wi
klZELiKo1t7nwG99H/yYHyX923B0P0NSvBkVvR1dcC+0LL64wh98ZcUJ+QauOs7BBL5NQ7mfK+cL
sKqgI/Ag6E4MP9z/F/YpYXR53Zs/SCG2ngbQoFmXPISH3B9uxW9nl+bxxjM/NqD1oIOTb6w2CAym
0OeCkrorQs4F3pyvi33jEhCg1sU4AyNVanQoM2A0rqgf8VkoI6elGJ2zXRymglay7uV/fUsM3zaR
o7/1oHOAA1ul0vWfUYkyLRQpVoMNWUoXBa8iFRDgog2dWcW4R34Pw6aGMyaBvXmi1lQjdNgG/mg/
QDAIjTDFA7bh6+Fpx5b5UBHQ/YrgA4em3NLdxvuZZLCPjYyzMbHmGfn5iCyvySyiAJMCIU4IWyNo
tUi+WjO/4yE5IMsetnhvIUb9YK+Wlk7MqzJ387xoHfnhBqCigFR/k1hMPchD1VI8dBEk/ckFKOVY
IxSbno4DIvoSx4P2jS7J2Q3gOu1g0LadUkFhD1YnkITfMZeKwuYh8T4OTSTAHa/Co+NB2gCfex+L
Hd5T12jaL4lXzIhMjFbHe1syYnKTWE9kNetvGtt3QbN15ekOobVzMDMM/6Nr5pM0nG6dp2I78jKY
BuThap3KNJ3V0g5n1FOwoBBhoIKVh9CaVtHQNsIhwp4E8+Y99Huu4LoXKkCjUZoVmLxBlmuqLeF+
XgYcsMMPycNau76NOwCP4/y9DYTyJvJxO58f/bsIZnnE22WxXa463aW+FGpTOIiMi4T83M5FC0hV
djcexvZsfEfnbnv8YPr10WKfaG0XMe8pHGBjjN4MDcQAh9Yc5njCYllBsCCB8FeXR1nxBym4bvVT
VQ2Yne4YmvK/z0PBuaGI5tBovaJl+7GBkwJsnS0YCNJBGznvbwmUfL8yTP0OFrDwlN5xztwlECfu
0EANZOXhJk4F4joTGfpkbHuHqjVtXflCoXSJRrkdjWAX88Kf4/LY/An4+DB8vFa0EjA3k9nNgunJ
AFUQ08jmzOiYG+FJespvJabKgbdn88HsUiR3oNxiXHimcWEjGgKcAHy5XHg2JmqfBN0fkrgbdgnP
C2jq3W1EEHhpiEfzGarRNGSWy2ZboCXsCGRszvsKJb2WIgXXiqeW9LftCUT4bYfTwGEvDAIiaYuF
Lwm79bsgdfGignbpQEuJ8cZS7IQAPewqc6WBYauLRI4Q3hFWQAGHT5iWd4StoeO7WjK0ckfNjGYb
49mypOK5lHOk5032FhoDgeTyxcLoFZEtyklaLwIsiO72fX7vjgcOvU08KY44nM6yuYfnGLO4Mn0h
jvHgiOUTBSUYOXad7QGINfbtE3XKxP6mZ9ZQMo5VYDq2XvFx1B0EBEQr1jzLmuSgSwSEM9ZoNycb
JJTWiVx4U4aMHerXM1CAaDguggft73Z2k/scOAip8uhZ4ZTt4osoUe5hRUaJsFMcjdfh4wjKS6p7
nNwUs5iEhorSRQrhZpGopEKR/q0nfHU3G5PT9LU8Q3fPg/cWrXu3izWlx7SjFvvbBRMbgLF+b81y
NZgm7WrVfOA9TpqaqxyBAgkfLP5eo/+sDjnKaAo9wgUWqPl0w0z0AgWQgnhWrcJDPwump/MHpok6
NcNsrt3UxbyoU9nGWOQM5YwX7bAeaLwwKJbofTtTB80Llw6dDUSp83rMjBIMHPdyEzlxoTfBili4
ZJYi7ApLN8BZ0fvHv4pKsTaxGyeTQv/Y3AJ9i6NcWvVfRArrvQbLPG7Ils9ux2dBBQpnHZTeqcgC
O+Mv/bxRI/E+amR0cPZKF+mQ8G7BtLtQXHFfdqvZm+Sgz5CUv7/hykEkgRzjHyT3mKco9yaHtBYj
2Cw9cTllJyYWdvA18LOtX3GhkxxJhGc6GzyPkUfX77vonTphwP1vgB/J70Zk37O/dBjfcU0wkEVJ
wXyB1u2TVhJXRpHmroT8wI082DNFb220aTG1Rc5dAfsb//a81pOzji84A4g775aAV2lmfG6hQSHv
3p0bCjYcd9IGdcZ93RZH2muFGxsP/zeTyD8sOr3w6YjG3TkiYVqO4JTPqG+PBSfEUNwen6cUOAh1
BluhA2Y+S9PN1yNdFbR5sRz/mtPglIeB4ITiRUV1YsexEujhDIbbTv9RZPtEKbIjb07C42WAS34f
2C2rexMiVcgic+29Z3RT3e1qOY6aJVbjZ351nv8kTZ7My2EFbaJEXm8T0gYyrwp0IJcgRS1CVygk
gKkIBNJtV3KbhVc0sdsFCwshx40roaz1wNh69o/OGcUcaEyhb9ZSvYuxs+qmBp+UC1SzgafEHUul
m/qCziSQg8zpUCC2ykql1sBB0NZO4dh1sthWUT6SONgZ8pRBvBNdES4OIUGIK+5R4P9w21CyHGEd
zmdwjXrAS+jCfziUwZiNvah7ZL+wX822JrVufn2BwYYucopmJ6IIzJhE/EeOyOg+apIU+3FQ2G6c
8kJYxD+DXTevqnfMD+7g9SdmriH/hbOEOWbyf6/CJwzIf178iUq0l2BYOIJpFRaxzynE+R23FdNV
J6+itTaLseclhpL8E4ubYom3evfqhDOobK0HmDxCWwKFp8PkIUpBkHwrTk3MulEdMIL2bAmNP0g6
3dh5XNEPoDsAe0jVcAeCJiWW7ytyT9DWws5T8zFdQSS6Eh+QoRGyQbzWxjMB8KiIQ9ar65YoZqt2
B9jjv4KljTJ9hIEX7Erem6NZ7AGf2+P9gjQehZ8gcLabtw2YBWQvH6nddIHqbI5lqHJd0V2lErK4
lWoNSjFUmaPKI9OxjVqvcIIiIT8ntIU4jbfzywAzJFlITCQJk9+RVCSLVokreZsJg+ruiKWJMFm6
UVEyykeHCN/fPGqAFdT4rUU5Er1t6CFlTd8UIZP7D+wpTN30//Tzr55TqSaJLTGje7rTc1NI7cta
xGdnnYj9eAKkq9pbmHz6yyFQdCw0h5RVQKdXBQwCKvp6g/UOsl16nLrQhsORmW7CtfYEp5jH9pvy
rQuUmzo/LMeKW69ARbT6J72B7HEHGoMbg/rYJ9Z4DMGIPp+xryv0PBBKNRN/yZYSD+oOjSklUxZ/
7EV/KhG77c7IuQ7prANNKLHR7181bC8k+vsGENMi83YG3RSpK/NFn/0LDFBmHqSLLVmDl2BLkKU3
8RGgRvCVDfmLe0LrcbDcEhEs00zJInOJ+qaP0rd+ai916cdi5/H3aciTtaDOm5b1v7wAnc9Syh/G
1VF4CoxMxAaMjXPGgERRsApSENJK8NEa0Oq5NsC7MZai/dTitzYGUXh0YkYuB4LgNTW8PFO1y0sJ
g5CUfFJyYr1LH1m9StP3Y9EtrnVuZjqt7LvQvb3XaLihUJBQfDqFJXGP+hen0b+Q2PDVB4Idz4Mw
TDPez3+cqSp6mIVb8Ut3Bd1Amd5WUaWrlx8fRl1zvTW7uOOHbtbMkbsySvhJGtxPlQUB0lySor6j
x8wPJLXH/NGVAUFcenPxQESbbZgeO9qhd4oK3AgAmFerxyUqTvfojGTUJMUV2SIbqm2/bx+Urxl9
PRiQ4t2ydxwstPRyOEh4VARIVg/TgN93hTJS8fGnHtzPT6AYzM6iI0+ttEEMCdiSBb1BiKSxzGvA
XY2wFbU2vvjWNiJ5FwHsJAgWYm5tZjCQorivwsnlbvnWPyIrBxsIQ7AbhHz8Dg0YnDV5uS2OWijq
h2UHFAuORY+henHLntYIUGInDxVQKJWDNpSbCh3Jclc4/jTe7jwxCT2bm4JhsKG+4nNBDqFcMJpn
jCYPs0NAgye9i1TF31+/tG1g7dNZ3kcMevvgfLUOcU4kP/shWgbVnF85LZKWR3k2jpFl0sUEC6P3
pvzJDjMI5BRY+O7xrwpnNOuPirl8kxJXhxa75SgzNRAx/e8ZLgQcNMYCkDBG/JhO0D9b56tTfcgU
XGHYR0zLkwrhRELtU2VDZQu0KS2BPU7tpira76TWb8LrDZwJ9C6jJKkMKpaARJIcYtvmKxd9wr4w
YFSMU9DvUivq/feGL9YWYSXKuW6FIB7LkSg8q0RYhxfXB1TxO8c2teEm/zdhpfF4xc7BDTvYJgBo
+55Q+t8I+0lgU9BS+4hpcIGzg5X2EmGG9yKxov2j0wW2bpoiV3STVEj4QICyzPqHkjherNl+PDyS
72B3l3OLhwBjmhsgkei119yZWGkgZTYzUrNleHRSjqm/tzAU3+k/ys9IQh6otKXi76S/nxqX611Z
d6QmtI8E96eU2D6vYcTIQNW0QAYFqeRojusjHA1fA9Nz3fuGWo51jTiMGKs/62TpcAIrnFnvQf2W
vVTWQWbGSFw1jMGogw1rYA3LPZXmQLeeLl8KYTrcuQpsyHF2kV09774CFXNTQsTvLn/7KoKLYLAi
htXxayzsws65XNKCyrZUSZonilseR/JXi4M8P/76SN8kmBf0YOzsHGgIOYoCpWj/Vdob039HhN9S
idYXzzplkBmVbzgiUt6Xs0ZpJnXUf2xNGNYi1K8Lo/DViH14Wj/rwwEG6Lowa8dCN9y8sC3t8EuJ
xHzDr35fSOtS07ja//l2S4/Nf1SAJt8moGhfOxejq64Q6r/vtf4IPzQkpBqAU95sVW7S0OXSZics
LUxEzseD4aWq9OlKdoRdHMNp49t+eByRAIZ57fPubLuJCEBqV1n0w+XNlah1zQDGcmO/2TiHbnI1
UoQZilzqn8GeJ+5esa5/VANjaX/cUO66YBmn7IbAwiSYqwtD7uiAdcOaEME6ww/ZQmt4rH+5uO+6
VL0Hv8bsEJR+5dgIkZ+Q6+9MBH4MyupI1KJmRIaBytlUn/pTz3+MeTJ2hWHOkTQrx4tULeqCcC33
XcGnJijnYBDXlkWn5yQSyHBjPGhMG81/GaPTnKtv2r7iygMYfKgh98Pkp3LD2zMhXx2mppkHZouA
rEcInMMj+Yg1IpOj+OhacoyaWBCvduQhvq4B2kKmp2EoGChDYyOq6jCB+6geb01Q0EKQ/qVSGEaf
1SqoTCC1c0y60xMf5TY8Ri/w66Y/1qr9Bpo3qCM9yC01yxTtCPNdt4sz1pFTWtKC78Lx4v0FT8i3
9GiY1o5Mfq4eYynGfe3VKUB4XkNnUlG9vG3kdHYWgC8bDkdwaWCsxjKXgVox/FeV0vj0zDAZk+4P
CK59axIL+5ISbJ65W631z2jT67hmmsi9CSsdBhXbUEaScMP9W1F0PsUz0Iy/KKtNsBxIUjv7potl
pq7qfMSQCo10le23mNjp+skIppMjj/2ubQIpOtfC89xQB2+BALVxlAsWy0Yb/y2mTHLdH3+Y4GO5
ZNIQrLRbTrFFwtfc6uhI8RooFEjlS3xOk7by9z5K6qg/qo799NUCVxsxJM4VexTJOjZehnRsJHmz
d+UL2iG+Q/qXkluTqGO/DX0Et/VKdPMdFjqA51+xQRG88GSp5SZIi7Ab/JKMeFn5B+QHMg27I771
xLvr9DKWumRbetcM93GR554oShsbhNBmvLYDn6okkFw3OBpHh/2Ungu8lXey4XygZ4gIyarjs3h/
Ww8MzPtDnRn3WnrYS12mebgDnLvlf41MkEMpFBGlEoaaWvpdRKkiYNEd5yWLnt3fnnTSCEE70tQA
xLXYA239RnJEcXvhIJ/ul/shMpOfHAxOIu4AWBup2D6v4UJT1uXhqNf8nBYsE/0vaBb0vxK7GG9O
u7+bVtLkJVl6a1WIxBP5WLMEHDC7Tb4rPTMSUcHGJp3UE4Lh+ta8YGnoEUJFtgOIoUez5HVARvyM
cbvgpBwYF4YEv2kWxBuwdtK7T/o28CmQWtk6/bS4j8UmdtAMC6CuWcNyPEQlGPtfWxe0DzRErJR0
r5Xiyc1Ez1oHgNvH62bb7deTNarb5gdV3G+LeZaHOOH5SNpC1DSrcj4Jyue680S2YDL7R6DeuqjP
JaBO0PuQso4vmyyBwZEoTJQ3D6oRYG8Gx+Cb9G8l4q7V/sePDwXmtni51orGtUGVmRmf20FmFACl
Oe+0jX9aXJF/X3/lwLvGYfrIUX3sRfSw1nqYIFHb7HX8z+8hG4Lnz78yqsnOE46ZcQ4uqcxDqgg4
liOFfyXYT777ARdST2Y65GdObFUtUMDDJvPDwepssMigZvfFLV9zEgvWRYsnLCazFmn0RiPS+jfq
x3EHnv3TcYG21FbwB/ljSE4taDdvwL3KtjBtbGbsCVEpK64MClMZj618xF6W5wxcS5DgOJILTxZL
qXV7jFLUjTwthWxMK6hmwSeMPkIWSMh4wD/GuZ9Jwb+Dm7LPhoq4fdHbghJ0vimIzgoIehWFJbMz
Y/hlaa494pOHtoKCFHulIsLg0j90C0OuCtaqMpBQ4RCOW9QXvcytc8nw2YQ8Kz6N+bzqbI6gltml
cFEEkOuUQ0jHkdZ0TBoDX0QqLCHp9J+YdEzNdDneod2ey1DxpwAtCp9xFhKFsyFBJU5/iIEkjxYq
0cPB0r9/RS44WHxaRg02j0ZlGMN7FNWXu8ONAzO8/KGA0TxZqwUUv/zABefqqX+ayIwJfaVe9kst
T2xr28eKEJW4gJlxI+rz77N+F+JJ6uDfH9pILwnPwuTDpV85TnA02DIn9ccr5VTbL+T8irimwRwU
sCGxXsVvA8f7lkNjDznxH+vH+eCATuYZyjz9YvxfsUsNIpJ4UcdCyC5l2ihFpiVuTR4TGYI5dAXY
E4CBvALDET0xr74pSVVcr0hLIgU7Xy1WxEDPb5vV8tnzYtAaaeRfroCZILBH65OSmK8Khg+k8oMo
7v8FtX1sPfK9g0aQUGd64bkLcAsW0akQBn686DxSne0I8hUDx5HWSId0YLkS15jLdY+NhFvSK142
NFAZD4rgw3+AOJjx3d6zd93PcCRv+QlhbLcR5pwmtOPDWBM/D57Yk2J5aMmgv9PQTBapSbQD3H4n
yRdje3YBWnzIEzbF7ZxSaaPc4DkOkoxxOntP52IEI4pfNX2A0mVl7koL8WQZ6CacobQQ2zYEDKb3
Z4jmLSDYKL7NQ1KcUtKWyQuCwS3iyS4bmVNtuk/7bZbI8q9a5SL85KWJKxthmamw5roDFSsOeaJh
GpVWUr6GqmjqR24hdI4z1utwCQExr/4jAFAcSayrGGM6ru3Vb3A9MnDWRj91oUiFsq4mYIkyIInz
UGb18aOCJRpYUMyOkUE9e8Fazl2PLYbUns1rn3kyHMpeqSqhVRUq87AdSh2695Oel0CrOcbDcRcL
78aEOiJ85fJ8sOYfN6dbKKHiOMDrGAt4N/R8kPIo728nBb7RpUzm1l50ZuF0GaqAgFKdiPpGRMAd
+tdFeNqCcYUDz6RM6DXmtyqHvIxgQNfdVWXppftVeWLVQ1TZstF48my7Z39T8V7ggSGwahyYYvFG
etAzqHC7jtLEOdOAUO3pvMljtJnyzW1+AIlKJo3DqGp48McsXX9IRGI3Cbok6GSxQ0ZN8KeMP/7I
A0+rnflt2xFuM/9WyqpEw59MTgX/1E7imzTwKeV6CsrzZUTYy9yRjeTXYLCobGJeh4qU5ZxUFHvg
qyqb2zep3amhOkjoFIa+EXAlaz+1UJ4nskktvpbtqTCDaCaH4SSHORMY3X9ZY3XKmZ+s4z9ZKr09
fiZiL+uk7dKo4H+MlEhsptdg8TFW3sE0RnYHNzascr0/I8mOxdUZBFN3eZ7jXS94PXlUfzgnqsNK
OrnexKx4shC70fz8M5S/BQyX4oB0xLMeIOMVkKXTpm8ZZK/rws2iweazTNCXnoQ7IfvzjWRJaE8o
uLIDhrJRwFbbMX6T8TVc6GidRDVEJam+fagyGQVowc0ZGP1YMlo7Zx9DjdSV3Tw1eF+LizT7mg5x
AwdNKeIcqPhyAlWhwGFamsL9p6WU632WzPspGy/2ESJ6jEuDxn9cKfC0v6/4MnkEwdzoLhn4jhrG
xldgSIIEmU9bVO9JL2DLzEzbwWfvAtEvEsmLEuBNs/77k49k1OZ/wjJc9xPojCDLL0toycDxtNXx
6i5kU0wOQJLaI+735iLGjkp8vbARAkbEzSjcnOYVRp4+24vprRbAlnR3VbBwPtcpz6y2kuldpNl2
kA9UZF1DXsUK0qmcZlmE7Fxd28EIFGtQrTeLNH+MvKSP9fX/kTuSJH70pGZgiPcssuMzeb+Dwapn
WHmqm8kFZ3+FEUdkfAtM9WyaIrarswbeGMez6KSuDuTQzwhocTiaj7Hk5TziLjS+tqVTXjZGRvLv
vJQ/0If/3Rv7EZPArmuexoEiXnGmL89UD/mMTZForrG2Sx95URezgigOjNGKkpjkOrsKBfQqkM8J
bDmOyFUWNt85bMPu6FbqMusIFrkDKC6ynZgLRc0VxOjTugF6xXeyFlJC8afZLkyTlT9rSedgVpuI
8p+Uwy+Te09cK3qCZzk38xHXdcIh17xWo3bTfz6JFNkj4H1CD28+ls7iH8BbOgChsoxAqw0GLZgN
z7jScKr6yOMgr3SrTsLepNsLIMSn/mGERflrrkGJa6YLQYYy22OjXg+NjonH/3xLCCRDrRefiJ2E
0vqvnjJQW3DwAq7bvVoq3C12Df5ZWIF1JmEJwWhe45oJgPfS0wlnqzVfLfmB7z1IdL+TU0Wg4FIq
DZN+t1G6iseEjcurqj2lyAqzTsm/kKqq53r2cSQwheppm3Y+zFXGcn4WqwZ1bjDEaT5mwy4eBftK
UbFdo72r5U71IDc7eEOjzKTk2pSjZmsWZhhnJEoDdSx/2J7EeM4KI8Oq0u87cBLRKNvgn/jYnnAa
einjxvTo0IHEwmykLxHLTQSo6dPPdHgA2Nl7uWLIz1CI849oZyApSGwMmeZ4AWJRI4puH5trKlEY
L1m9WBMLvNdRtFCnevfyPMapk9pQRH0IssMi4lE4XoxTPS0NlTMlCGhO6I07HR8XwSVVVe139vDG
ZASsx1HKh5gZSp69s4AUZ4pVIPXLUwkmfoF4gt/ekwzYh6oZ42xDPtsMrINydOZLHfzN2Wbt+xYe
QTlIweuNOiBPh751fLaxCkXkxxeh26St1qQYX3AlObYea40iyxV2WWhkz6pvdOp/7BBHHIyOsa8W
6qsVUU/7iyDf6zrei47CvC85FNrIPqsKHZIwHaM6MXVUjJMRj/AmjmRDx5fLJk6T1K2TSzPWNX1e
3qzJ0QJtlYin1BMayoGE0JhQc11PYjGfegJUnNAXf8MSpUmzA7TY2/+Wkj1tsG13dweAaY1deRDX
fvpvYaILc17Pjdppnld8bUdhWCdKQItlSFVMu5Affjl219cjhc2ZeQSbkfEm3U7WnFjjLMOL4p3Y
OeBKym0BMQgXxFaU2EoBTqOjVab1P8+OhboeNXZomMJDmVMheQeIelZNZqP6+aT7ouxbFYmvm38P
btB5qGferY0hJ9cQGH+PxwHLvft+LS/yCwoDEszKjTsYQeHJIgC+dqG0lM+f4+lDSOyKBGch48Ty
ZVU7/vtJl7PhDbYkRCSJGYtOhqbxDgWyAc6O0BzxL3oeoXJVTgP3aVOtpdYZNTG8c6CH0bnLqGRf
SUk5BjOZdbquDwgUsgA+NsKEgeKY3BOMJkMjwrkCIdVRVm5rI7ZLNEgfDGFgDk8xcxKtyYRwYoq4
b37NMgZntq02VH7W3XqGsMoccZXiYEIY1ucsNTkXuxD40TSesooBfSm8Epa0Xg4ZhhriL/5LVuHy
LOjtg6syATjABgpe5WtIS8P9FNZNN8Qxkl6zjbVtNzYvtP4Zy4riKAokLfpyoTXAO+kQhQdI5yv6
OC/TcU+qtMN8EdnjEBQJYwVYL25CxSqHapgpkR+v3cwzC+lolrzx9tSyW+S9VnN8W+7EyPOGAqEA
rt/aZrFmkNoFK92WchHFaqBYWi6dz7rQ1PHMpf+2DlGnuasleHuIXQj9GZ9VO+Xd3HD5ru5bV4Ig
kleqV+rEiXXXaLjXy3pH3Mqkt/GY4TQ9/iBg4g4VyX0Mmo+sqeRUqHXopI6IryllGXNSeXK7KQvB
4ZmLYJOnhxubPVE8xJIOSZgRjiqqL6IFx2gxKj6Fd5NAN2P85wHY2pZjHXysRBlj2S4cYg4QTcLP
Ql6z7KBwqthpKfnz/h4KHdczfgphOKPzr7GpJ+A61N+ecTWLS5Pny1YIUqizqSUhbA/N9J6Ff1NS
ags3UoYNqFXQ4U7ovSs3QJ7IWpVR/tCKVqHUWJ717Odz1hzfzwy3iYviRFNiJ+TujLaTrnF/uHyc
c9L2Ad25RKHMbcHgRIkljJ6QaoQWWUNdxAOawlSho6HGcv11YibkF2cOZAmDvAPN23/FKjxsW9xC
pFbIBy0L1ddTnTcWvIheGH1XsG/GzOvj584qF/p/VUgEJbULO2X46J11IiAhMBbfXxL/1NJcr3v3
ZlP4KP8saGMrKGrw4XYhGrM8nx5o3JNicK1qnc1U05HdM+Hqh8Vcxa5C+mCEhYdfKqVzh+xON8n9
P0ZwXaD05vA/5T4fH7mbm0DTXZDKWJn9oeU4ypD8ivKJHhKInNEWAMk1jnOQ0qzVTDYm0uApTu5w
KLzaqXd6DatljEEt1YoIq8uYo9nvtFQmhOFA1hRvGYd8eo67poFSLKZjpBaslYj5ZiyBA33Of6Xz
1N9WqYVRF43QkfOZiuZ/yy+n/1Eg3bCJLjsHR3tKF3LD+e7le/XVilfhy+alKvFEWZfvlvkdErAJ
qhYpw0qaU2JPcWwjZ4hUvnq3wbSZ+U8n9Umw6kmQkFNsPr5cVr63lP7zcnefgiXfdssFDElKwNdG
2royXQ3NzMpvZvlDSd68ypRymkP2w3tNf5rahBshwy9XcRDlqQihsf/zddH3zBcy+cJHttgeQWvJ
BU+3RgFEnuqVC3ygnqX8EvwI4FCMkJ9JjsubLmfe/g92y6cdiuRv4Qh78kD1HDTSAwyZ+h8FF/V3
76ZYtRcAMDUVgiIBSB4qQtFjfVcH4vFBPNW0Z/ZNFiAWiQWfd0U1QrTt2wSZUFA8xP11JwmIVP5t
1V9F6dBcEUYqq9Sry+bqSbmPdDxztRsFKTpyIPo3xuW7+z8itCvfKgfa/6j6K2C11WrHiO0T737H
zf4BJcLFDOUgem7i0a1zZE4EvhfZtv7WmC7UK+i1+8BvW3VtdcDmakeNxIvg/0IfdcHn0zDmWJCO
5hj/DjUYm3NyQUmVITkIGvQsQ9AsAbRxZr/fyi0r3XN6WGzIZC/X5iJeVrI0YHlIXqTMN35msnuH
r/dPSvIckhO1Fw8BPz9MM81rW6z1mruGQwUOuNU71LILBD8P2tTUzB1INQJl82GKVb18fX/EzY3d
RQ4dWjKrc1PxuhTDniiFutQ9B0fjft0L5/iWOz6QE4cQpGcZ8D/d8fATT0FcIXb+QU6O/xD2nvkf
JYVHrBEsr9GHcdKQg0mSd5sqFyYpHy+kDarYDEtsALnYa991O6OvMrOe9XQyQTCDGXf2Vw31kY3O
zig+8cDJKX16IMSt5WdBnr2qg6+4olnaLI097EfCxddOdZX/VKcsn6aOZtnaDM6d+FkWPbiDtFQf
oQwDo7icKdy2MKekMv17bEDOHY23Ln0YUMJRpR1RVOfX8QaXiPf+LZpy4DaVEsh1pUOWGtUBXm2G
JobpfzfJSaU4lqdn7aYLWav16svtiKBwslSF/H6X17aDdgRrhOviNjzHK4irqx+AHp/FF+CWAk52
3jPciAdcl9LiR95YR3CLAPsaWrT5aAGMIjx7KrmQyxztJ+x9nUcKKRyj5WODZWRREFVQopHyJ4nf
anSe+Chq4uHzLU/I63vBX8IjXHANYS5CTTOdylssZ+ArmsOBagbVLb15He6+4EtMpVw8vUkN1IHb
ZNpq4LUZnoDr/a4p6L4KUqajzTVFTqggeFsHPmP7CChB6oZ2XMVmG+PjGh92hFElCgCbXRXfsJDY
JHObMiVa9QRte6UO+/iSqqv7guwmlrsJ/WTXhzvsMDdCDwusaoP9wA326idxboQfewRgo9ZRacnB
IglIaQH6n86djBuW44tBjtNS06psryQUocpTNtqMiYvY4kvjzbeKMTrgg2+J3sMDgXVsQnBl/Nty
S4Ksv8zQkbxCV7VDIKpulrKCe0cwFFXTLXGzAlfYSKnQJf7rpZIMBo30qveqnbYUKGSKHkxJpElD
KPKGtOcaIJdbKXYQ3G8DXsFgXAgcVhi4wFq6qmh/+2zdKVBljiRqNBI8iHkR6xav2HJub4NhPpxv
XwnmdQe9HBGaX7dl4Gj0P6h8HqcgiCbL70jFcJWHfxZQ+r0k88MH0EYpH0JywTDzlLNCQDULwNB8
x5QyPV0j+udNzZVN3V7fYfZxXC4AuwGnW0+WmZHlJGeUCtTTgGCaDh16ch9xLJtMN9hL7h+2G7Zc
APOoTCgC+DwkNHzRWa25AXzvHviPThPM9wMW+07tGfSgYmpQIMJBLXo7VjqOjwLjtOV3hRrJskYE
0GAMQvtwHeW5wk4u71orLP3O9zEsuzYUgRFB3+J5N5garLRVV0AwoqEmjl93ifmUJvbe+cf/4U7n
igPLCzzTuuCyNYA+KRzkVqL+IhSKN1DYBi1oIvGue1V+DEAWiq4/y4LdtLpyA67Oka5N4kN7WJ3J
sQd4sj7AG5GqpdymvHIFtBeY3wgcnyihX6jUaVvkxwhEiKYBU9nd8XkAwVTAWvpp709NM285NNSW
bITuPd13rrsRJVbQ2DDEUkZd/nN/LujMhkn/dreOJKFK9FDmeDSA52vGi9Wp4FmGs/e7bZLAcqqp
bcivNUnVRrpC48H4o0NP+uqBuN/P83cw++TclVEknnZT4CJgFw4JuxJ6iGHXm2DOCU5qSWbexusb
IqY4zl5qS/leN3ct8Vhpfn12wYatMr571XWXqijy5ziTFHCKTzP4aSz29opn74ujnee3qBwbCvBQ
04sbYBc3ThleSmw9Z62yUnw+QoJ77YjT56RWsfSNyhV9wmpoJD2B6fo3H085NoRjW9thkNESMZDD
w0CpG3MRlgJ9UnNl9UmrV5rejni70oJjlfpKx5M5bJHBhybiliAj1dPxc6o4pW9YjsRl7EISxMbE
0RrrzTWVMXSdsExkw99W83M2oPEsKPwYJ4KlY1ex80oUFF6LqhzeXqKa2jSfpSs93brxU2tU5FHo
FeKxVpoAAfs67xRXr5l3L/SDrVVSiatMDtKQCNwIfflISqqO4vbW9uRgdEY5k2Hxxd0t+FgsEAO6
tZe+idYjJN6oq+JyCZT1J61L8Ly/Mp6ow9LucluvtuHiqO4LrIy8Uj6z5and41Q9bBU/5JKE2DYi
jXMIUbjfTgatt/cY/jyp1Vrq4zhWTAlRofYSwjLl7vYm12VvcPmv3jdaXMCgsJ4QBcJwp7LI6D7J
9ZJ3aDMwguYRYaWXPT3vhczQ7acRqrISorkV/hOEcsnMhcObOrOgGn6APgfNq2kmxI+rrCwZmwYY
5Vj49MDAHeTpWQP7GOD69+r2RY/JkW8ofNIvJqqjen3D597ybi6AlCppRegRYT+9qIfoDSQycixn
g24C/8CiX/UyUGOD363bI+OELPGvHbtrh0OIu2nicfQBlR07shsq3v6JTLYmBpH3lEbEviMVIXIq
dVmq/dN4qtDwOph2IIkV0GLu8jdRW6f+cnqrV9RdsbRFwefzrV+lUlY5N5k101ClC85m9UOrmbL0
KpBA+nK3XWNm9u5gifRDBgOzhQGqmoxgxJq6UUkitYDIxkfXIMZoyoZq43LYXhIuOiWDpfCOnJvL
cmlB0HwCIUOYRQn5zThD6LGtUBnKM9OdmaUKMLrO1BZTm4wuIA5z+xmlMuZFylehT4cJ+eOLiEEx
FrQ4n6Gv6uXhY3a7xP9blzmGL8oFVTvxoloU4r1YTZr2InDhIq5cNsPzDmM47BxKqjinA4xcL6WH
RNJYscA9r0HyZLdgI80ECl4g5+ok4H3/M+UhN/4DdBBaut7E7CYfD7CV8o1dUc/ra7AmE3MwDPHi
nU062my3a8RttH5mIDu3x3l958bPqWA2+V9Waukeuzkshung1G9kxkkEM+jDbHIWiXmONOgrG1Y3
qiuzeOXDkEkoh7uWd1YfXo86Xf/OiKCDshOFB6hYfhJXQB+cywqIQftw8bwI6FM0Fr85DVEX6F2T
FvJnjkjdA0kZ2BDXM+uzqRLfzsld9eRkqWnyYa9JhbsiaFoKG2zP9L+VrwjF0InzLace+MeGWW9v
b7baRrygoFZ/PgGnGr9ASk7j/bTtnzq7dce0tT8+b8KNlY21H/pRfR/BAZK+/4tIACJqN7nFVS8C
hKD2xRTe5WsupwP2tU0xH+PdEOvaZuOhLLkzhTuYyKbnX4uF0cikoSkCkW6uBGU/F6Tq2JVmTMcD
GXRmkfIB2N+y9Cp5afV7T7J/Xv74R3TB7yD5ORkK8+zKMAnqyBeWxKYEHY2BGvdCfnNtDqdou0Wx
xP54Iqa2k+8mvSgp2plTKrn83nP2PKVFufojEfnq/M3gCi2njoeZnM1Kr+XP7pq7/VonW+yYA0FN
l5RT45PFqJJ1zG90I3l/9RR9HJWxtz3nlaeEn0pblXXJo/rRQmlnoKAodF9N/jVZzJzXRXOAV8YU
q7MhwxGcw0o5MpUatLWoL7slnE1jw4/MMGKaTnfn2K560DMFSHVitxREwWyP98KKvuUdevy2ylyt
ykRUei1ZWNawNHG5tqN1AzqZbCRlY9x77i7mjm3aTkIPKusnF03jX2Mt/0UlEweDSwINkX3T6JN/
DArewhJJQJNZLFDJXaUyvCGFjN20C6ireDgr4cRGS4LwPG9CZNNkFtsTDPAqbFzdZld005LyAdJ0
aoeSzEQrkUFyg5372b6+gOWxgoXRyEnL2unpLohwaX71R2oS+70g2bF4kOJKu6px8S0xQdVcbS47
mj0T6vELiNxkrdlrc9kZhNrXNM9Ut6cw3reK6RXG/eWKqIZRsnUTtYJABbppZJVwQDq/90srqSzY
TP85abB7TZtaIPmYu8dF9X7vnfy5WBf6soM5xh+zfi8oYU7j9GBIr2akjaYsSlPUspvqORhVBpv7
1WN+xXpHBtxAe6uN5wvP3gSntkidZsiGOtg+0CFSeNnUY36Ps9XH9QT56Fr1DOs8tE5q3Qe+GN3d
tPwJDrldiq5bRNsgKTZ+8/imDSRZ5rWYfpujBm3oYuDgfUc/8+RKWHeg+KLYwkuxrbPvjY+/3QOx
a/QPd5n4bnj9XUxcfga/eTw4Vnp7Z4dEbNS5zPl5eMed2wjY+PxsrIcZvH1ajlhLniWgJQ7vgM1e
rhDqPKWsHQistol7QPI1RngGnj5A+/erWu8ZE717WvP4jw5g4uQICCMgFSgk8p1dFYw9BbPjVa3/
GiSplcvKoWHa0IJOiXbzJLVChgMzPhp85TU8f5wWj4YurjpO9xyJZLWXCraP7k9C/0fCbplo1oML
Uf9m99Kovm/3V5XJ/ZBhJLAlc/MONJVuxqgh+cUMVjn5QFCR101aUGEn7bGT6JTCY7lvwuaKPoTJ
bsl+DETfbMC83us0Z30gZx6SJr4WPYtN4Pvji878WwqW0vsBHDYEjyyJ+9Eu3UZjU8z/EVOZfaYL
gjDnxED0so9/prQ1VJtjB2i0AM+4SStH3iz9CfQsz7K5gNAlvG5Edvj5qpYzGfHyV3FWLtwiEHKs
tNAdKeBZUdYkZWuz+rgwoAf89tYv25csQl8u7ymPx1a49I5FYEYbSmrtGUcln4FYI9HVY6lFH2YA
iJntSTf5TUrb6UqljEE/opE6Cvu8au10IntTzWfV0gp2JDmSEAvKKmXgPZvL6eQVcSTfNPDoom0z
5Ujhz+LRfz1uubW3KJq2qlt4bUaWeQsgi2OzNB+1LLY5mYhsXwd7dK3Jn1OVp+KeEeyHqrWIuryI
rabqvHFHjmPHMPB5CHf76yimSZBrZQtwyubhQmIS9cQZpI2d/kb6bkzXk8H1xD54Cn64PdjYR6zj
Ssb3HUGpsB67Hn6Aldt241rpLbjNBaM8oaoeopeoY9ri8RLP/UN4Ws4DJoBe90r4XZocIg1JTxvX
oTE108uAZLR0GRHb8Skxqx3N/+734fChURLWKf7sojoDSA59z1Mw/81Q3MtonJ1kLJQSaw7PV7OD
I/5P1e8GVTQ2OlyLngyfY2+p/hp4VLB+bZz/TIZROIZqchGSJxi5CLFKnXigEeuQauqchsnBfSAE
fKjbel6qgfOLlR7zPU8WpLmAW/iaWTox4uNfuUbnAGgL/+IRXVe7P+eDyQ0wcXRI51JtUlQ2QlgJ
J2oILtnipS44BmGGiFLadt7avFjqT/EXN5bLKCONPB97qEgUFApf5PZSSxeCzmpeQk8tqndv4MWT
Lol5Eb9+mVY/IURX6UpFChzJm6OCN+EjqJbYbHHtgyhwq98eQenzBF12INQUZdCeEK0VYa16vNv2
6J3JDI50j5ZgCh+3QSAeDgpObBge/mW8BLF0x42kv5JF46EUFbkQCgeiDGMK/oj15pdQXNzzTIV0
0js4xVAU/h4tJivP1/KKt/wfZxduF0BZ1Vy/ZxYpV58usUejUZfCRpMYDWrGMvUw51XrytWzzW28
DpLCoh2yBCIxAUU5cX6pIEUj3jfaJQj/UQq4w6PDBhEcnOEjBbDvK5ZR3iR3dY5hqR18Xvfzaseq
WZvQnaLtEYw47XLcohxso3Cp/VyqgJl6U6zdsIJNbmzljnhTXhUyzv6YFig26Ew+9TKQZCwEWZcF
SasAmvq++FUQcQNE1EO+nNmQXrqPU+a/gfKBqc6kkh0kfQbDK35FqMPScHAY7UIuWt615Abaam/m
m4xwmrNEtAGRNrCMjsFNdd7mY9muTWKQ2awFgLIh7V39pNGumai6c5Nci+XhRz/7R3kuvn92zfGl
CDaCxIA1r6AvClHd2ybeMB5nKgdRKCuPmJpJc45mryB8kM89bW6Oy+ye/EE/Z43VrYrFtG6a1+Ny
8hxtxiple0S7+w9n55hZkA5P7eR+hl9B+6VFCm5OCnGcIErOj65c+KMuxLo638FWCRlvgiW6gYIj
4n5I/x1p825qgKZ2lk+GU12Nssr66ayqt4+YjQDhufWzZZ/MR2+PFd5AckfJqwASiKpCea/bdsjz
IlrkVB5u3cgZrTf61rE+ebOHDFczfikbuaeX0c2czeF+VMsEwkLoVbPgMCG/oEkYr0MtuvR8tRmk
nQlUNfmUPjERbPxwxSyujJA0e3/YC+S7zQAlfjtg62iU0KlrZSDvUL59gXrfgCjU8fQurqCWwcoI
8PLzioKo8eYYxT0NTYV1kR/VeNT2akBnhLgGUgtj7dCAD9n85yc7XgVtndV3Z3iD8sBYmjECiQBD
iDYDXdspmmNzb6ATAT9Nn2aM8wsJHLvpWZUDaGfWGIqb85ah8OHkOEcaEBRGId4hL4d2sfBbSwoI
hbFCpFCy3R+y55t4q64ZwlOsq/f26DD20sbCreCpinh7UMRdYYPNcPfhUTr5DR6gxUckYwmEpuqW
0cgA7JFajshMSQOSJnfn5F3tSZ3kYXYZfMQw/5E295KeQrXIefjgIrMoAU9bDnkK9awONhAAV+4L
B8qehbYN5N3svf8YBtp0B9cXVm7kZu2gMm2JG7CxMb7ScWNTAjI2mr73exlq8hFRVXJHxhTMdSRG
Sprp8nypKxpDzvDWPSZQ4hDRFQL+wZLzgCQ+6jWxLLGPPvqPoRBE71z30r5ZiGfECZKiqRs7mLOO
yGU4u6V0hoa6de8QwZmIb8cQEvl82g4tl5X/e0yfepL5SpvaUwMV8PSJMEM7L8CPh+1HPfD5780V
AyLl6b0MtALjk2b35LKRcJlNWM7IFRbrSaYORbmrsU2/tlDDCfR57m+FKITbGjkNylGwtEYsTjHt
Srai04t+Us2PjPo/BxhLG1rLUoKzMrOlHJ7fFzGsoujMFBJNVYncjIyyBaQ/8DDWqSaUlcM4dKDj
4q0O6wyl0SFMcz0OHoF/LflgFQGgyGjqpHjxo3n8gQm0IfeN/Y9Rz527x2ZfGldvt/Yvkfp08Qib
fVELe0w51lTgWUNhyFhs5VVWmgVWPWfy7KNOE2T/5dc9pzLk6CRsm76wzkEt4w1cx5HjyLF2lkd6
XhRpu/xaJm/IGN/daDn3gPCe+T8S5Hjvh4t1rm2a1F3k/JdPkId8JruDGy0YDfj7seTi6TR3K8hJ
aZ0ynv8vqjHFXzB85ReL3GFXMS7QBHNVfs4sKcp/jOHnNmEHXAfyWkRynuKDpIGP9eiwV6YwjMQ6
wdDvlEhsoawArlx3//5qjwHXDLVHPfq1byMC3VjhTxL18vc+vm9tiOAVP4Wl1KOKfzXwE1CWiiVS
U7t/UDoH4c7aW87iFRuZKlZ3ONfBaZzrlCnBCrAGc0h57XUT6Ow0P9/A8Nzj+EEOQg9wSsKUf4C5
Y3Jg0bNpwXeWhKpknkW62GwOYgHhJKur+berAWDnDqxZiJ86ukhvG80JgenjfYwSNnDg16yXtfwL
ZjVYuCTjF9azS0mioKWq0unzxnaBv+uFICquk2Ase++VMs2nVltPVPfajxjT7Zl49X5G9rWyAmqK
ZekmjCWOQHJFKyvAgtw+Se5hDL3A2NaS2KoVV2DCEWaqCj1HP0KZoqfEn6RMr+vCFZ7SgOJcdEbu
ivLaT8DFQPkSlPow1FzG9sgmBdGrvTgQMqigUzqhcUdCq46cu/fSSNkO+3q5gUUhhBdNZjuPoxpk
WyKIlCULF3jwghDZBPAOqUUMxOSXT4juyfWRznR2j54/bKkaxmw9mjiJ4IWKp5O4XBmY6Svcynsn
pgckkYxJMO4Z0GWQEm/0AQlUCa4zriM0I8JI9FXyDu4vLFrOt5QW+MQe9pGxJO/9irL3wlIgPWG6
Q4I8OCbVf5QllcGgHq9ba453W/Sx+AyQokSDlh3UBa0kQk+XSm+A9RqqClgZoAz+EQa538dWkw6/
aB9ll2I9VlO5XPbC1Wd5zV5aIATKhTJoZpLn06kX4ARn5IjDCmvk+3tRiAituwQ6EX2R9cWoIG4m
flOiwDG1u+bdNfLO63rPaK62BIvmcQsYoyO/2NdRxsRarwxd2fOjF0hRn5IgRbyZV0aIrua8PytJ
0XZuQbC+BQwbN1dvXL1/VLc+gMkGIehAlb+V7ehV40oD50ka7dOzTHQop493h4MKjw2tPoYSBo2s
xkyTibdTwADwnYYiwAELMwqBes32CwJnjROmuvPs4Gvg/PlJuVXXmWfEOS17DWtivvcump/V0DgC
6EFxmF1Ct4vxTd0Auklg4Q5mGRR8QvPewN/NWU9BarrXg389dWNB1ISMnAxhmw5TiJao2qWxudrU
qASUWiNoh8FurXJgVteE9cX3DZd3/b8YVel8XQkZS/h8AzFpilDIPiKc2QpFGlVpYmRU5jtqZMol
XyObOiz9JnHj+ojw8iH+1SRIRu19K3ImT1k8IZS3yiJDKeoNs9UoAvCmlo5Pd0dEerIEg5INDPMP
yETFDpsME9FRPs9sKfZqgaG0SqFpsIcTS1AtCsaQwfH5jiL0Q8NcKxqxYu1S6HDs+DjkqT8qa+me
mGm8+SdAJriRWUaqtPiwSfcbigpfV4UhJCwuxBQx7sVDkfjb7kVgI3EYFy/6Kqyg31t1HzAMoxvY
hzofTzab10OP0FOJaNQwy/VU2W2PE3Lnet3v80D795wPoJVNKhtGUOW3eP2PJYtJ8pBpOFUSY+gN
Trw3N3iXmjDYeMa7N26Sw7qL6+1ZLaZHalFeSAzlcVaKiYruWh4lCM0wV5pHPD3YjLQqW0JSXS2P
a0Go14EwqLPDYTNKxMgv4xFgwzeO5ZEHifsHMWladmvclyd/4yZwIy/Q/KLzJgq0ueXzr3uXCFMo
xvmYI2pO7JGAYl1XRISxl+SQwtvFBT2W/EwGSBdfdt9yfdmoFjjIMan125QzxBM64S5qISc0J3Ka
ZsUg8d4b4VUX3QSzaTUHce8+XqYbl/s2rixd/0Qo2lqL1j9iYxUeHY6+gA4AcmuAqPAS1T6VUNEq
VarjA4dI4siCze6CJeWy+U0+5M9i9PoOU4HTReTSUAZXQQOelg7KOLpLm0Ka2qoScv3/8FF0qsHg
UmJ7RObTGbxoEQBqOAnbhbi64BVsw49EYaYh6MCiAZR6kb0ajEDeoTxhohEi+xrs0qoIvKVmFCyS
70mM38hHIDknyujORure7lZEjhu0Ho7wtXhw1Hx9LUxDLKktvRwuBD0UxGErSqdoQKhuG1DzEW1W
FlgX17zD1A2nLoAPVH2WSQJ7SHHTpO+lvlScnAzrlzSwiB4o1BuKlgVDMZPLIo0G6PNoXZD4NVG6
ZenaxAyVzPbUao/MVHo2XL/HTk8fKNxxyg5WcnRJ3lakztXYKn32aiFn4neNyVoJ3DZxiJ0eoMpe
/XvKpfAWsA8Tc0OnFyS1jG3C725pdCyWoX6QehShZ+AhZkIXXs5phhkitmmJg2e0lec5pNbH8MO6
eD0vT/eNEXlOv7ewxnkDtpdkUBKs5VTBJTGIsHLYLFvqoF1qlvzz2kPVIn2RNyRgztR30tv85vvT
EQp+nqSw6ImcXQpiCFzHiiOfhDt8XsL7ZK1lvo4Bb+ps7G/K0/ceTZqgagnk4qENFLeyCHfOkkWF
qt+y7Qi5IM3repltwQfxIEkpcjqUFM94/rf4rQIo3r6Bu5BV+ZXffM5aCMm3wfAzegdJCk/AeSCz
+sJuty8ISx6KAwpDN3q0fJyUt/hdVmwPU2/mhO/NM0xGg06LKFihFQ+oB5ysOSAmv+N3Y+3aLZEI
892+kGww+i7hMx1xiOTVU2M3oVW38/Qic/sL+B2kPcbUG4ZLg5B+sQOmliSmj2yknfaJ0Uvm/Bvg
NxDNd+OO7nRNJ1kaKSznTS+g8ID20TKSsXujUC1AtHLn9rFZODyOfgPk7Iu01L1PKuQi87Oc347P
VVIq700ThH/8uwDZy1QGWLGLpXTZrOv8ncoqTN8YBYLADz/iagNomrecVO3+3ld9/MHWIwMoCG8g
/tAcoU/0D/S6zh7P6ZtgShVciS0tD6xA8R920gbqQj+oBYdPN54cxm3axc2r8aCeG5KuzUGIj0bx
j/9aZ/zDI6vfbKREnjLyHn5y3JdwDsrvY6VjAwJ6qAJCbw7QDN0IQloMAx2N7cToXiIeUrMm+mqA
cSSP/8PlhEiQYy/RAODjilqqr+9thJ8GaIFv6FBcHyWRc5Gb2FUwW41Qib/SSU6Of5cAPQSlW36d
MT2v0UjAym2dPPjpKAP8vlyP6iW4xuLI18fwkIO35mUs4cmIx4gzaY2JJoPfVMW4fNc3+k7aEDH5
6xO0OaataH/6+ryaj1Fc33FO6K4srzIUn35OX1GQ0bOIZ6PUHMuhOJiST1jIUuDgc4ELeImjhOqh
aWQWOPugHJPC0de3LJ1XpLqWMxvYW0jVOoTaB8DA34ZOV/O+GHsAhUAAQtvvzaRdvRmZmXNtFEo9
+3CNVkKtY1H4I3s1O3JMCthyy7KrIl0b27qMBcAr6D+derIbllrecP5TLXARZbaqpEzSmdKoOriC
KjBMsoIetG0Nj0pFnq1aiJBo8NcCFq5/kWxKelxcEjUojVArrmouqxzdj+7YHcidPM9HfsM2utJz
EYLuFZIjUSKGG5yHG/VKupANb+haR8wNMAWS8jhpkjplv3LKyeu6PIo0OhxKh3F6f1njF7YAvtKf
Zpy8ZWu1Gn55ek0zJ624hUgWJMLOEeMzUIN6h/L0hwipBj5eehsURit7D4TkVJuJbesfp1rPT6A5
W/URRCUHLzJe6Y2pzCk3gk4CO6rLh0VEnxyIFBxfGdGZmwIfSMHR+Pm4nm3yqGyaBP6WtirFXfn1
QyZoENv+LAuZRwBxn+9gAuHGNcTFkmDhsRrNxwelzhmFYS7Fgnbcx4qCAG9z0AwKGRdr6p4ZTfz0
Pbw9zvtnhrAx0VJjD+HArNbHokw7IKup5J1dED9KNgK90Vewu468q4mLneNutpHV9YIFJz6uWSMO
DGFM60pKGxRiWotXBS00WogEBykJURem+aUPswF1X8mVe/XFlnOJM+0K2XDtb6kpHt8p5shNYc9/
vnqMhGX+IbWmqsrO4ycRBJwVqigg3BXejiaXTx18dyVlXENNl+/AdS3a6WyzgZ8GVOCd6Zt2fxTo
lJCGSD+m6dQPTsBKZJbBak+FUKIBKhPxXDGWgkp99gYQ8BrTqZCMuRKyW995k1Wy0dIkCO79aq6O
5M7COzS7Tm9jnf2oEwLLpvlPFglx+6PcA7xDRBNn9sKUkv8tLq6/14JwIXfS+t5sls4SMU3z32vc
g+y+HhhoMrNycddMVGpcjvqRmWxoiFa39NCklrOHipCBeNMq28nUiqGQMr6NjRZMrRxZ5ayFMpLW
xNnzazjVQXU9pqlYBdnLjOZ4jVQlyC9TqXD+9fxoFOVhLHtqZBKk2vIxXPoDOfZRTo8HdTiakijn
+kFsy1kS/G/30To+b3b/2JmaWKImQywoRlwzFQSVSXnJkq64xhl13Ox2aN83K7yw5WXx+LH2J1By
6R+mtL8pJVD5vdg9jI1yngpaKtuRn1M9RsBpyxbdKEYyn8i9iC2/26J/KqYi/MOwl1VPKzYVpEby
gQtshNQUsPTd+mXxSvNURIeNxwfxK7vErNM8AdbHmcg760YyDCFRR2hn+lG903KHFlqm4+DnUdYZ
KssstPtl3IK8g6Ota9KRt0fSxoFcRGMtBZaUBT8c3Wr7I4rQhN+eMNagzTWLEAtlA9ABCNw9S79L
VI/PtlSOI9a9N3jOwolWAGFsNoEh0gkfy5L4Uy3eCbBJxNPjKG6SAAjHxRmjoEMdMj31MT5GpSch
k7kE1mqybGkGeLZ+YMADSpd04TBmoTSBjm71VdR+yNS8BmRKL4eP4mypXWM3ccG0TuBQWjgLzFSE
UnhJnG1rzMnXAGiYyMOD0E3yXpO1BIHgPeIMnjOK0LIW6nu6sn60sd0bzt3wECLSu52zioJc4Zva
0QB5zYE9OaamfSx/L9YN697Sj+Es1eBagOLAZFCqDlcQtg60jZAUnx4puhW+TjQZ/QOhXFKGUuhQ
kB4vIlUJf/sPCaDhhV9CXhSwhGhdUgxP4dDT0qLdzlvvHr1SvWK/USijfc6TtW/Czv7vVCnpTu/o
IV5pHTs5OwEp+AtB7TVUiYHWVGYn8UrVuI5qX4BrtDrzmpmAY/9a/Rnsh4dofXCkvGvadgF3TRhB
TvHyI9I/mqAKuBpZjf8TFSCYShfGe+q1DArpE4GnDUCVABCuW9MjsCqmO93rogjwtYDmed4Js4iz
8P6NQHzcVNq7Ptp4pkkIWjX/QLOBBgtJXz3W9+CegDCuTli5o3EATjc8bgyX4gv0SQH46VhLlyo6
H+noGhZatm/ckHTCKIl7adIO/VMocbKVQWuqN6EAtVCzs+DT2i9GrmtNxD1xSoDBSCIJWZB1PyP1
SfOSRPbWeWt/zyD2nwZk/QQb+YR6fHPwYL2RUySy7E0txAnB3dbDXAqXVevCtEGBWoPncCc15rTY
A+Ngit/7IXQeoI9rzk0YHYVdhdfuJegleBTAYypbnofXjIQ2qi+B/T72L/jU3XH0qKs7CVfy6Loi
J/j6MI5ZhczcF02uYq3kHYui2uSqafYOhL3knUhLheukqoOBiYYGewXARUdi/EKbYMTRXoZsjqLV
1dUASnvMEHFoZhzt7E9pNfpsn7kFuyH54txUMi4lsDtSnTM6pPsVDs/GuI2hY/vGTkjg1mZy76sD
1TamLVWXb2DqF0daU/WOKkM6qsobTcAtjmICjLZeWpVoULp2fmCA8IsehVAuDkI11EyEvAZHqaHc
sb/kTcKdHoINvNJ1l5YMl6aw2Q6Ni5+3mrodedkxgXxs2fSHHWIitSmg9wsBGMkh08SuMlayV/y3
6hndb0mNu5h9OcvMUt0saunqAEkMN8uxOjfYGwqvevD9u4RJXps7YvORux9m+pq3qaxI6pE+gaby
XueN+xL+wGjnpblJoaty5X+HgUi+tsB9RiOwfVR/JTaOTL5GbqXFuxK7eFMVXX1zR7Vtb8cQEy2k
JHXoJV882ZAvT6eJpaU55QQz5f2KCcwAX8r2035/I6decw6EWYpvcjugbCzdUWFvx6+3YVl9CGQO
1cFWvLqaZDzdJhHShSNAtB5PzH8bA+miH7STM4Rb9td3y2MLasBXE+t1bs0u0PDBukNplWP7CrZy
UxNuJRl+8KumaLO0a98l4yh7tyticqiJDEnrtgw4QOz5a1UXXyM5b+VaeTFRCAfGCMt2L6TZbiP+
ybBnfng9faHB73mSe/Gmgt6UpyUCE7IN1Ehs4nBFcBVqLOyqnk9rye4HDTD4Fr89dggfYIkf9w/4
WzyedkCgh8viI3Fhtt5bNpKWeTOjiXozHpkbyd2wsa4OpbQbF0D/F+KGZwdnxzw656eKoSTsztF+
C+RugehTr2e96ACXSIrWA6wDHGCGZMrY1U8D2JutxHK/Q74AaqUkA49ZGQ8eD8b7cW5A+IOxAWCS
hhZspT2XHjhAH1LJdv69Z29ehnKO99JtobD1DbCm0Xpg0C1kRSvPFm6GAQdoP4YIFIFE73uFk8u+
twGKj8OoRYiPE3ZMXI0lp3lhJzS4jw5H9Ov59xOtEXIcvolaHZ0i6PbKZJrIcZvt9RP1zzV8C6vG
eQtrOG5flWTwE8w2nU2ZjOo76IYSinylRIUGTdSN7RW5GvzayIx9fwRmICdeVNiYgf2N2msSmEET
0DDfbQfD1xhmA3Itl2re8htoYG0vX8CtRKe8EY2bW/GzKf7U2PQjzplA5fs6dRBO6Fb6kbO9+7pu
e03ikqUfbHnq+/I/iloEg6NwFKCXqLVIPeIBPEIB4PIDZEQMK+tmBL4Et2lc4fps8jWncfGmECCa
5IwFpeXgO1UvMDhXj7ueNYn+WNoDwNSw9HeImL0zdeupw5gqH8gRGBVo9KAFaNqxA8oajg3ZABZj
ZhLJSKPgk/9BDeFm+dwVinSi54lpHL0VW5kKwpaYHQRLxEUVHBZuovN1a4blI2jl2m9jLsNS2dIf
8EhEZB426fxv8UYXaMOopxKW/0PGB7az3WmDebeYHo7Z5kBXrPD2ceN9674cG6VKJlWUJLAVPqbd
jUAZ0qvDGmGjrdLj9CHBBDtUP2Z32KpMDO/3srIZylElw9xngQCoE0VQeYe+dNY0chKWE136+X6s
NQI8SVhMAmXuTDLu1E2R63onlY63iCKF1haPK3vLKaXTNfB5aLfntRusWuy41Ly7eWJguL7DC97M
VyfXrxZ//cGRpsaKbYlZyycU1EXKd8OfkJfZ8AqpW3mn3cnNcKyfPuuqmPug93tgj9eFDGBG/PeE
pAiyPT1yjpJeiziYFnoWEO4++p7Mv8r4FWQex7C62sNYMZqKX/ICOH8yAUPyAq8PqyPcXvkCNl3W
5rsls8bnjAtoVohiVUYk2VaYlboqO/hAtLMOv+NiVxzNhR4vZaU7t/hwcvTihEvVmzlWTxd84rBE
7nST39TyEciTusFEsEyi9+StemtvMymJHNFBXJtDzOx/aYfWnBG/1P3JJ0HdbkNhRjjL5oBDKxWb
9paArlti9N48BKv2ld0IiJwP5vnqAMlMN7l9v1z1V3HWPM0Xw7d+Aw0lU7Qh8z+Ri2Z2uDL6nZTQ
UTePAlf/oqiqAHCVzmRRCDF8PpjNesyWqwSLHBJKTtDgOl+3wQ1UBEgGspfZbsHie7xQU+FjRLg9
+49QaLhH8AbH37fX4iP7WGzdNVpUpJc8fyJQhiHZC00BenC9WZcbd2pCiEp4ozto0gUcoVD+qZg9
4cDBsl+k5/sxFNSvGuTFtCodqljDnVeRb7y6UYEzCOD4WZjUv0Omd2kDUeseb+4xirOeNlpkovqm
oIBU8zTvcQZ//SpPZ9UGPkRxqKWRuhHWJgb5WsZEFTFMQsUgkh85vL+1hW1SLq2A26CATGwlVqrO
lI/OyPExPw/v1LZqNWAbfYQZIs2ALGMj3hXxe4jHpZx3I0Un3fjtK+Ci3j1nsD5x80FLnga5EZH/
fImBsBenZ/88r6fJE0r2o8LucjyoR2F4ikkL80lt9h0fU0xB4DfYKSN7lghDfhcNToTF9uXfH/jk
va7TkZHnRW5YsSIWjHdvRC43Xr52Wjry7hwMULCwgldkRnaCiNt0grthIxLSbHcH0oDIqQA1BPKF
NjDs5LjkfxF/V4/ki7bpvwZDEV/7cgWU/VTc2S/bozcQSQyqYY1/tWOob7QnF7dwLdhD6/aDMLjs
dyNebGf/zM3kSopIW3c7gp+lvuXsMGrjFT9Qe3wUVaRPFcIuzz+98r1jyuy9s/QnxW7sZjedH4+m
fbG92CUsfJ/HqDDEkMhDk/eMO1tV6e1UQBRcF5YJ0CYxOI9zUobzDV0eSSiyv4NNPgffptaj6RWd
x55oDHy5QAAYlSlJcUngWRwrL8rcMhHWiW93LIv4u1/IBUtRTWyKalAb7VlY0A5ojWBEcu+25OS8
haYEnxHL5FNF9FiCLo+GR7DKsgBk+mKFtYT1HvVFlHXwiKZgKMVEzf/eVzQu2s0nG/oGTg8G2Q/n
gSx42nalrC3L3lZjQ9hN0sWkUh07yZwFXiY8kySHZaC7mbtxM03T4Fero/KOl3gUEx5KpTCK3fFq
cETuG7wLr7jPLwH8T5qq3rt7QWyvPd3kM0SDeuByev1H58Fnxl05BUhetSkFJQej+c4BTw91RRJM
SKz7t1dcJ7z+dMttN6c2J3sq+X5BRxYoMsFqxu9SNRrEH647p2URRSs4FdzdGP1uupkeqRx7fnv8
9VqGMJ0SF3cPInCBfIggfWFbxkQaduJHomVP6DKXB8SbIQs2Dfy1LrDSsqA/jXB+8k79SPMkm6RX
n9jKem4GYKO6E723rchm+d2kR/wlrenskFUMzSD1xwXDrPwnuvbSw3wglx6NKGdli2LRv576M1LB
ZSLLQiKPZfwriJlF/LvPrCtGqaMEaA4hBPQ0TRoIzg26PJGmY/nlgDjNCoP4u62SL1YW8ID6/TQE
CdO3oSGaBuBT7U6Ji/Fx6JlXbABrITn/hmm5+KSyr03MWt8jw6+7rmif5May0JKTiX/PlwW5Y1pB
ikns/Wk0d1EfhUwDe4EaimA+dg7nsh35xJORMOX4QlpYGq9tERrtLuz5ZEnMRXT7ZU5vdrzTfpo4
ewNzyGvSJ/qPRNwHi4LUOYB1ShubALsnh6vtwTZhGW0Wt+u+kaEzO5KuKDPH9cagQ+9riy/Uc7J6
V3i87luJbf4O8R/DcyhhcrPLz+DCnnWuGw51LC3ZBOUpNftx34QwGcFv1/tTcmBcJiDbpkxjuVA6
JtGsuWdSyOzrqmvxd0Zi0aW0J2vjzbcHWv4ceH0sQaWafGGk3wTxwCGLi2VTTOqZLApLuXtoqdOx
1gI8Wz9SqCB0Rx2v7ZspfC/BpXkn24R+zbiBH6ZXZlpLh5lrUaJ5IuqktdHQYUfG5W5nrWl+a6rW
oVBbTx1WP6bGC26GW2crXCXrHpBhJYmeE3SAfWgZT0QPesJDgo6aIbgt+4qjrojxq1MHwZ26BQXW
jcfWxTXyZ7fKJXuDXSh+fhDHfTnZ9HPRokzjjRK9h3oadmzMafD2cn3iRPHFGPRYI2QFfGkaVLpd
mUfB+6Y6psZGwzdxeFovMzxvyI0zD8sawS8rYbmkdgEbjtUB3U3HB4XRFQTVdby4qwsHjVRlkjHt
/GfCYRauxgCKJhSQ02zBvytGxC6vai5O4L5vQCfUCXAFbaepXCMdqfuPImuM/liZreWZjxm3kBtv
yUMF7j4ILQMDDlWJgG94JmqazxAUBJwPdvnQgqtKEgJ78dO8SidCkbBly27F0agDzOZDCri9dxoE
lC508G1NKYVR93Ra9H+JdSzL6h1yKd07ENzQ44O4BLYFGL+OKTj8pUsbT74/cc/SjnuxqvD1fbfK
ultaBp60GsSlDlMG1GiUF8MGKhRjYOriTA1Q+bcz95D/HTBxxtl5XQv4ijOceUnT4AA3eWUr1bhU
/GmTPTmd3yfbD/VNdjI0WuGc6dKIngTxWQsY3FWjdeRFDcx5CiPa6nlb8g/BF495OSL7Qp9HsdjL
eAbGpUu0zKXauLAnS71y6iCuqNeWiK7cGuY4s+foFv70Dj5Gsaxn7LqsitOCysrp5wsNQ/dodLve
aLvhM1Uekif0VG7DzKZoDYz44zCu6kDAXt2iaxHLA4qyhGMAnz+n8Oq/0oYS/ybiWF90tXe5Kzx7
ehEbM2UWi1SNi72n0BMnXZeakRozQ++EOd1m0isMdcqy0tf+Vl3etUh+k4+abi9CynQTQYHzICcw
SN5Qdmb8CVw9WO7p0LT/P+4FOyTYZDRhy1kWvMj5s7W55sRRsMQ2kYH6a9c4xlKYeiOoppPa/4Ig
0KmuVY6232gSYKuRZyZq5wA6ep2w2GKlmeWXxGlJ2bxOnoKCuzzJ6OghRilwu9/TwH9GVIlwE5xi
8MoK/6ZURI4MWhiCbSJX6aFi4i4ZJzeMZqcJtm7WrVTucQDYnaSB56Pm8I3+8jo6Toq/0JAD90Rq
L2UbXaaNBjIYNH30WgQx7cycbRZVJqkfwBG1c2mA/CcF2ePJYc5Xy1FUOYT5jh/X9jNUiriPiKr7
4a/fYE7qWu1l/lWeL+wZ+01mDfUDvGdMm5VEqdtDhNMcuXOryysrnX8rZq8vLuwP+HVZvOYasfyP
ThSZVK+IQgaEn0dgM8EXmwbrn44JkyDT0TtgvkOMSXz5GC39Hl0gAWFQDDD1rpgc6s+NCZgDzGZy
b/HFZTFFDQ1gzKKxKvwrJY0wKwQPXR/dc2i7uTbTkgHirILmk8idxObbA+IMmrlSovq493gpQjot
M5KUNFmteppZ3A2GFCELT976td3zmOvYiikngPAdMEE0yNYtxECct8XNV4szBf+Vb1fRms4Rr4ev
s126fPjnntVEMmD232eVH+yuk5I4Ojr5VCjxtwWJ69voVJllAcyMYQUOKHPu72p2yFOwUyNJhJ8B
Ta4aCpxOvP1xPss7/hFJNjEuY1gLCow6MD6vAz69ZlSWQLa46K5itefaj1P5k7hR2drqPKdKXHpU
tzyzTnTMPUFTxPQEdbhaYiRK1cBECeccvxAoLHtSx8zLf7PLNLRJLkLG0A2J2VmhhKi73V8V9qVC
U6agfgRRP/Ne4c/6Pg4rXZfHz+vCWXwDyMQMWhu2vz74bDFs9Aug3alq94U1zIL0dgHsYLkM2ms/
Ku5LQ8JzrskcRfemtMp9W/zT1awZEuBv+5eOripqsSpmmJQUneU4zv72kA8DhqCdl14OjRDO/SLn
cDnQG4W4N1eghZMFVq059gcKjOaGUBMv3oQ23erTjHd6lYiZhl29x9P1sUgEbejm7ogvgxAnUrO5
39A6+RbjVISHCI/hh4pgAV4P6kJY1LryjKxLIUP09JFk6JIaBARIuDedJ3FKRBOsCgBGVqDbxkLU
AJElWE/psda+jGKwvbBb/Mz1u7pzA1icmMmIwFIDgruiKb8DhGu49e5umvv4gzJvg0hxvwsN05ti
YUtiRYCirMkehCiWEzuG6xoJFI8NZ/pMOpYXsO3DT9EDIJT+IaFGdIf31iQfJv19lAAE86ytf0Zp
ILZSyFMv4raP8xLl73LmZTCoF1kgBwLzVUHNoczN26z1zuENcPI7Jsz1xJxoE3GxBF/vonps9tjf
nNH1GjjyQK6fJWLOhC2t9j65fXQXAZAuz3EY3PJZyMzrVA4ftN+cYSZ4NKOHGK+KvVKGYqhlykGI
AARkVtDiPfhP4JdiVu8Cdt7U+QuAemqWGHoJAY0K2x1R8Fe+pvPMfbMsqT7dotN7v0fwWCp5L5rV
cFXl1IVxFUnNbGayJb5/oLP6plbDy0P41JHo7yTKwbFATqyhLJ9eyCK4ey2/4erFf/iLIciHNaZv
HIsbqHzGtlpaaUrIhHAaEIE75rWlqSFYI3GFj6J1bX80oPCH9qPs3mFOKngU1ib9+molJdjucAFM
bqedBiIg8wBuIpHpmGGy5Jm0cgVlx7n/aqYJUjgQd9N+TEVhMrbTP8/VIB7WhOrDhtvE9x6XlpTF
maONEvzKltzxO0ipIPm8tBL3VK1TTgAAI1oYtL4+H5Z7KjavhnIuCBMqfLq6yf8wSUJ12oncFzSE
AOiqpRSgFKmbXSWyo8bN7YgWOXzvI3AAe2Kg+for7fvggLHQGvKtv7oh7Kl7Rkkylh5roqdiLCds
ghK/vvaLjv2wxAkBM4cT7dlcPwxrVfHaEObUxLHcbU9yJNjV+2Xjs2DMfRAfvXurwqL7/ocuk6lH
vPK06DJZhKhKlO4yGGFqRcWTCP4zZC8TQCbWRIF3PHm2A0dwNlAg9Rxg+RgfTms9GeppBSZIO+6N
mVTd6PC9ZlfobYn2RQhzudeR2LTpyFOShuUiC+VgBa7W+Nobf2lMAR4FS7JkJo8ps/JVPfwAL1hl
1ZXWd1kw4dESt1AbgAAsfG0MUJsHnjCm8cBDVJbqFHWet//RFcVLODIjTvHQpIdqgoKV5100Vg8v
M2icRLD/lzycw5k2xancfRSSRVkygt4f8uw+Q7tB9Vpr4kktgw9sp3C6lfRyA1Zxmw0MSPHB3LPL
w8rWfAAqdlO1q+xsc+zSNkLobyuvvcFa4tNQSQ4FVCPCgVpthO44ccB/fquINJwn/S6V1dDN1FVy
Mm4pXGOg9FxsJEWrJLjWwpUMbBxPeeogB9gHI2+pIqdwaw9r3UHa6qF7cNudaiLTBWP9ysUR9k68
tGciU+KszTLBBINKg2Jxb/LL0fTYfrr00K5Qhu+1RpDqOetzNQcKIBJIEQTEfR5vWvHl2Z8tiSgG
OWskgN5m7VQEpoTZxRIVrbvlfmqXWW+XiY/zH5IftzO0vTf/kdipjRYO7G6/gbFFgRR78b2wOylb
xJBGnuIncWkbGSaTJ5lGfX1Pl5la2qfPvs5qB4QfJwnJYXnz4U9ncjJYW5WbKp6vt06iLaFloc1d
nHeofaWLgLD23PVWH3EHy0mHBCjk3k9yeImvFHoNh8STCMUbXjYuXm5zciBkggjaLrY5iwRqQRX1
5r5CaeCk3sZX3cU3iXjJb4gY0nQVSqgUYV+DZBSugRmbSCK1lLYKANn5nsOPAi2g5ZEdm5M1JWSN
Crr9kTpim9cYkZhlBhBiyEAHizOtptwLevLn8kdIFsILdvakBcYrQA9+qyGYvMMJchU97vAOYyQR
f1EJ62Mwl+jr633HwqxPBf9QzvKs9CH7AwpG5Y7svQUPNA1v2TE3Z6taxcun+9MCT/mzUTuVVGfA
SDJmaRlrI43AqPbzFN2kfy3E25x12eyv/XGVM+z2vL7L1wMyo4swLhqJYmf6zElu4SvwfzvYRzoO
MtaUHvJa7lRoZf/Mykm3tBuxOA0BYUv0P9ZejhXIaW+19WwGWzq0/mJU3Xh7NvuFB7wm4ZGxDab0
khjqso4jjgd4AW8eow6pXHTFHKaBlJfBuF9NcH19YwS22XYPFlKBxZ7Xp9fJHahXizG1yzo4Gm47
Yyz+sOe7rFLJ8iEocY1AHFncK3TgUDwuNBLxFx6aTi/1xvcTkQf+ksMGwp4OO7+UcyBWUAGMmDjc
nrLBAPTbv92EaO3ZIrZqXag0DN0C1ZAOxeBihZswdiGuSAvqjfPYD84TsQfFio+SBJRyHeIeP7/C
XN0px1XJZN+xTN5jj5CN4G4LDaqsrNDx7eegtMnX1LRB5lsJ1w/MJIlY5Dbu8suAwTXNDNun29vB
2H4ZV41QIb9OPoRqSKEGCeRj2desglFjZuQsnvo56QeKKObf8/pgm3jM3Wdy/Zsi/NPaeIgdXaNX
pR1bz5u104tKHMoZlpyQ6kH1u/d+NakC7zrjF0XiA3d/QAPAHGXIpwmlhDiIgQrBIvTM9OIEXqBa
/TY7v6rM6gE3A3rQEOueTtWhMaSXvhVo0bsJG7QygX8EureD34h1ijwwMYY91jz0GQAcD/VYltBd
lvHTFXomaSx63RJZBt6RSq3gRcBtVesbNyMRr+U1s3Rn6agd6jpacPs4WWcpmYYDM3VOz0D7nwLe
4h0FXEhov2GeDMS7JJSw3D2yN1K52Ej6RW8IPzDUcF7Aqray4uCs1XbPkbo+vypfl4IP8aAL/oxN
WDNjjvChSXrLRjZb2ZSe/FfYcFbFwu/zwebt/RiPP6cIyxqqnO5C8SarH72/tuSYYCFJEGsSgUP4
lOw0IC5cBZayWWRhws3G7W5g4haQXKvJkQkmotpY91O8KKKU4wJ/qn8SAbrHEQ8KLipvJsHuxI/y
MD89+Xr6i5fTchYKQy5N6LaZGVfPXth2urAWOX1MTlephEaV+MEijk6w7sztuwAFima1QufE1lJE
tVJMegD6xdU48/z+MJSZXWvRZl7ciON0Pdl1stRjOvXsi4cZ72YovleMaUPg+xo8+e1CuSFoVLEA
AVMzLmLvjsW9gswe8zARC82F1oAb30LlAsYL/ITp8iP11fhhp7sPzpGgkQIhBphctCn2iKZ6lGQ9
+Sfr83FJcgyEOXOJJg55+8y8JwMS8K4HlYLSBXTgRWbvUvF5zYcIOQPpCRM1w3x4reQww/xj77G9
+yiVNkLS1LPPDys6rRw3/OLJc5eOaJNsFRSzHRgMiRIVXlimJPN/8+FRDB1QK9bDNCty37z3VZgZ
doWynSkrQ7E7fCJUP7+uA0jtJJMkChS4IYNxu1KWmUpzpsAsb4matds+wnZ+dlZqQCcdn0kRxJ1k
49onKnSJJJS0DFj55zvuEuB8XN5dDkd7EkMSQpLZAPaNzAv61jfakpYufWUNNwWCHd29wmKlosa4
hSV70co0t9PsM7x0wHLnWEGp7nuT8MmO7thbXBgG9uGxtq5rSOWMGPHWGMGtA5bYcN/LHkncKtwu
/JjlPzniUMHpVwjq2p8PDWrFNdvMFiaoAebMeE+x2BZ8LLtYBLVw0y2oiKBT2buJwU302/Lu9Lbe
ksCadAn0GDbldrTFGgdx5IvahsnHbCH57LCFE62zvkwnBPPpCEmreL4tpMB0ckx3sapnzvxluWVn
NVbB75h2NN8c3JjmOtFO5y1LgIadootLDRKYVSTEmVIq9iGrx3dycLgFyezlxQXi3Ja6aZ8RgCw7
Ec76MfSeNb1JXFekMEfh+vWl4gT6pD9zlN4io7Z6hC53Erct5sv0V0WH8F0THT6zby2ex/AfFufs
R70qHQNcGGcYeYxi7/QkeQA9thoCjf1bAdyqoL+RtEsaLP688O0x7TvIP8OxE4GIuymhe3zOm//M
u9A7bQ2QV4C045cRlkj6M4crvNO8P6d89t+waPoDwtWl5C1QcyC3mAZvDTRilykZTe5cACPc4f54
s91lXoZhRECEQPf//RVvxkL/e6UISmE5rdcPeIxIQovGoremapm2JPK0uoeXd8epBKmwqxWP0CAK
iDiCFnOTjQWzQHpBZH0L2Hpxa3pViMcUK9SnN7dhpzO6vzWzCw+xmPNGPZnZxI+Qz1NwQ0qTI7lN
qpH7Xjvp+fmAXDRaJndrcplLxVB/cdOZBNXDouQdqhtW2kqAwm7L6EeQ9O5q+U2VhNEaeoMWN4pz
h+ACo0ct9g8mUc+Ac2xea9LBzu6Fg3HAQgooNBf9lFQ5qXQal2dj2RObiahVvtnMXbnbukKTDPAr
Ee95jPcF3WgSBUOrfyg90wD/uIeGiJM1Qt98ZVeiTYvjXV7yt6eQN+OCrAQvwGmrlWKGVsEvx6Cz
gwKwdww3OcVVvM5yIN6g8qExHiVfWU1PahLShHt6/CrMiT6A51Kk8JygJ8Z2FJPXXNC1yS6Orw4v
5iE1EcrKpBXFz4MFz6Lf17aUPRN1wHVoF8DKyHw2STWGiZyAV7DAgBAiTNnfHZ3VVOliiR8z8XGo
au7lNNjCJ4s6r5g73kIaHOXVRthpks+Pyx5Hf5J3yxy2LhGZFGR0BeHE7qx2E31N8yLc4/kJUxh+
M8WKq0SMjL3Nd8NDSLScvuT9CYj7m65mjdewUKPJ8bcKq/VS4qZry57KZnj1/llgh6h+o+iKzqD7
Kb9yofIMYHSiEUHB8fl3a4arf/zJuQoxXG+eojq0xsWbvixLkgfUSZOdvh0L45ljQxjMWJyGflRn
Bhvz//gOa/u6nbl3DSESCLm20hhUA/HK2yEbCWgZyy9+VWnQYY4R2Sdv2lvADv+tY6Jx0qlTv7Zz
tHnhUTNhL2uCHnm9sWvvkZFsEvk4udA0zSzMn0LeulsoH3E81U3Hspf9tH/1rWEhQVp/xLGjARLi
0flVCGdmZ1aUypznsrQ1t4T52qtQgCwquSmsg+X0f6+3DJdut9ziX9768IJidXh6R4gWBdndIJnV
wWy8lpeTGt5kz6ZKRT3lqqcdGWakXonMVVVWZIjgGK2vgCCZGMoapt6VF2A3bohfNMyBCNWStCq4
q01nZqBgT9t0xhkCIX5nUfqeW2VyESKtolq+eeXbqyMaJW/VvdUsYqg9EY37AynYOFNrz/W+KQNI
Xl3HkEdFACJUCjoHHj+3QCK/yvTYAyAKjIjKEjGceWdsItYdUDXeAwTjRy8G+lOV+2nweqPdKzst
lvzmQwdtn3BkrdfHzRAH6f61WwrMqLxvmjEs9waCPIMQ93kdM6Nbd9QzjRKOp6j7C0tjxj9nt22H
BcW+M31uHK4vB+GOspI6H5YtNCdKj/2vhc2zw29aJ360Z+hSZeYq6E1WP/GgU8a0w2GjltvtO2GG
4oPQxVilIJepBqGjYZIVJvtBDndykh5ry0hLOnBhVy6kEvAAxhSdavQHMKFrCiXkfKDPgSVYA8E5
FivScLl9Fj0wt9ZCFICexavkAd2Uekto6i+9W6ujZTUKTvpngDejJ6/0w7SWxXVnOyTNWmjmO31X
vCo1iDKpr48EzpoQbltnWQcDDSze+EDk083+4tMA7zoClX4d9bTj8UyQM3rm5esQg/8bNOgaxDU9
rMYK8crhjqeLbi0Avpvmr1wh4jdV+mXggQJtHOJBalANHJb1Pwu4GPaY6lANuMmXoDc1n0dWqcbS
c88dKx8hrhFvZIURSjH/b9xJ31pXdb3o8H6Cwi+ns8u//XihAraWdoAKwEimBTSj4RHKvkkZ6iPH
x3OkZxEqEj4DdWfuWJh2OOQqnlAQEOKN7SgnJU/xHo/O585ucc1dr3lPRTpKYl8UBeIMe/SEEqTj
eJpTSCd489jMtcl8awPnJEi3Lh5xslaKTzFdHyXiqwlCq6WoAr+OhkprnzuncJpNDckKvWG6rjYU
beOsjifH0DQ/pewLLzg0oqCjVjnourt4bPd80LFwmnToMv+LEZk+8hIvGeAaFX4eC3i9QujG2w9w
0TtdshNBXE7QV7neehRdKejh5OeSXzHKGe3XEbGminbeBVgsJGp3ZbbhqmA0FWoQjaXgZuJn4c+X
6oVtA2qWvGpi1jf8Wf6jEnJ77+ooCUvXPji7a7QWxg8ODLhittz3gPt+kqG9vRN5L3Xt7PvMrci+
sLNWupjoomhI103bs6yUZE/FenYzwat6IElbn/H2yiD2j+xpCzWVxAF5sqHgeKzho08tKLgiIlCa
ETFc377U8KWJ3XwMnT985o1TBOCDWDy5P95lr4mK9HTMuxfhbnfekYxTJl100sxxdZEsADN8fAxg
84Ky5NVMjTX2dREH+FvW8ex54JhzdoclsUvkJ2uBXVZXNrc4fKbRB5XKGmSM268NoP7MBlVc5QFA
ndT+L+t2022pNTa+Xv210FIegkgfqHtMCCI7HTcb6kf0HFp8K/iCKKGeY2fNqL5/dgNWbbG4OG8E
JNBrOmE9BKJjYZIwowIzLRkji7s62IQEjhPvRjhuxKkZ2oPMELplYtLB84epCUG6rfbDWQebIXjl
W4e4HUqfavm5YDKvrAY06hl5c8+OsXTkjaftsM2paBzwccEfZh4nQpGsZ8zJZBMBNYq79igAw/3n
knNJGUIg9oFXopuLTe+V7Pmc71n6z0EFPZ8Qf4tyfSyKjH9VMTBr83RphNBP8TnVuKX2weBLi1Bp
Pgmj1tM3XvOXWNvZnBiCp1X0FBwS39o/vH4ncEGGXFA3CemmNdVlG8D4JxslahLpYfVytXlSYau1
DyA1gtYcmobn8nrKFxJnJecYW77TdcbPQJL86rnx0oefsN7hXkODceOW+f7ykzbQhIzu1ZxeNN7O
OheJFYC1D+GQeKBfnxNDvvOMBZ20YCm1+RgOkE81es8Xjm1OZxDEI+qs3cSQqDaevJiHywK8qeEm
8FvX/pASy3Vzu94nomajGiiwMnfuaGVoTn/CbqF5yNaJBbbB3jB1kq4cYDdLPflLEMMS1pCfnPLy
dINRRZ7N4ZlrIC5yAdEnZTDSIg5BemAjXEWPgoNgNRW/8LfZCc2N1/0zjh7EXByrcvCDVRNroiWQ
D3dxDzVYtbxV65QmJFBd7SHHIQb/swhBiOzpTGZ+vLsugueulZYYgGMEIGkRBaprc6V4UVAhvCYW
kxkrJNQYVLe5CW6eunmO+C/5ZcAJVZiYCYgQZo1GI9dk3edqAANM2zRlHQ2bi9qj3J/abYXfD2UF
J+QPPq4EycNKlxFlY2zn2/TSqm6EvXjq7CF8tifHviBfYKK0WIO2LyyN9uWCcQnLzKFVjgLwrCzn
6e/Woq0cwfmjoP3JGLOHufZiTXRgEe5ya7mijlw5NcB3ZRkEgHTnDH5Gqa+1TfBhYsMxesFDtB5/
RqTAEQFQUO0/8+1iavgrXBvDePBjoxDQZ1VSGrGTVblYMtbKDbd4JOlLZvTV1bS//mT1s+VCjswZ
VHjWWT2Lzv2nlBwGkZ+9fboja9e6/S+uXuIHDPS14gh1ZyPQIRxzXzODSlzpnQokqQoiDoOB5P5e
GQOrWol4ciSeTp9a6ayk35q/ap3+RmoNqdTP6T6Ru8rkh9fUIGdx1fqKQBrOq395uoppd8WkCacx
UusEMP6oyFF+LOwKIJgMKuuvn+XcFGGWRpW+Dvny7HZrT4velcp1JKo2gKmIJsQR6rzJsB7wGnaL
A9eLrx0iBsgLiiYfnVT7sI0nm0cuDePdg+hBIqg9lUsmOQCqTeiK9O8i7W71S3NEi7VQQHp3Ufe+
W4cWmx38AR049oMt7CzauXk60BV9ZST0uFtLjqcPatnVeqQgGYPDSVd6cg02N8USAXe/Do0+Mg7V
CI9qsIb0o8eEuicX/ZUcgcwAtlgdj5iOrB+0H8mdz+5Ugm2eyOAcLCJhfgdyKOAzeyF2cDt2QJmG
TqUI4xa8utG0qjD/AuUSr2u+ernE0YzzqskWy8Z9mwF93jNLTq4/iMVx2b34wBNHFwgDexszFBBO
TQoXsQyVC4PS4ngoGkPPMbYE3FoqI65ia0fC4nHxv0XlV+Kp0FpezGvxaD/T2C51XewsvPfMMV2w
VaOSgmliF2KwIWau+XC7Uq/us1goBcjtAJTMZjyxkcYDQ07NC4HcVxXdJF5KEmXPoqWbZM8vZMpm
cG/q/UdpA0gLw/1FdVCq3wsEKj9/tttM8PCfGW+S3r2Qhe3hkY2yKPg8gm+/GMMpN5YTcyl5WvwP
f2+LfcIpSQJpCz4Gmz0Wv14bF4wjMadm77KvbOFszd68eMu5Q3KPLD8eBf95Ca9SLLwRqlC+dZRq
nf/9D9Z2x00Dq8qG6WgT06ie40L0onWBpmxCglMO/izSIphSMbixWCZE5nVBXbBRH/32zGW9JbQ5
mGVI9CehU944S7Yc0ishsdGU58OZh5vKHE7CSx+gTNAxWNKNvKSEawvEczj3+Wr7PXMONIGn3tM0
pxULi531ho5HyohYeb8rjdYCL0Is00voThK6L+a4fKven5LVqcPNbsj2zyAHTANIe++hRf9ounCG
QJBmvBIW01FKE6VFfcgy3Ug+BSxnepCffVGEQIE7jU3XeWhf9vgkL0kw5j25qUayF4zoAniX+6Bx
nipYeFalkfpVUjwJYslBmV3py/o7gVOYuIZGh1tIbhLDji/sUkmIeSBJBVCH5vgnkGoPtjJHpooP
SQ7CdDj3NwF+MlrYP1bIUOyQuXxrTHXV7x63X1qKqaE7LP92l+YLn/VgTaTKpV2aMCxPxDfgxOAX
Iqc61YyAk681j3EGllvFPgr6UUMUOyX69EQBIzDwEeI6Xwdb0mWr+C6j1934NS7brr53eZ0qcm88
I3YrstVKpisOM5Jk/DOKvY2aqD3svAUIMLeHbtiJZNYb9ljW4PoXblnP7H3wDJYdphX5nDWETMNY
gu9eCQbanYrUqkqBEEJXOEOFpuddR0fqX6aJFh9bpgytBFPzMwXdKrnOyuiiw2ZtJFC1cbEVtn4d
1aSAY/P/f31LF1lDzaGzdO8YQ1WCC3Tf1DYe87+zyoXJ+u30t3BmACVlkXU0+UqJjoaH28LGwuuB
3hfSsdLATvBjSNlXXvVOAlgoT/jbj7WCJCRN4qP3nZpdujGZOGLXyum/RNarBQAjEOWDdJEgfvnb
7+pN2ogGUfzok0oQaAhHp7Y57gBGcCcbS3DazQRi/E7s5ZkQVXutzr4dDXr/foPFtuizdNbZ5zHS
T7WHbGhvkyYCSEEshmJyW6aLeQhC469Wnx6B3IG6xTC5aWuv6SkWaw8q1wCoNH0k9zMxZwbSyEWS
bDFwe139FzsBZA7JO7lW/6Nb5Z4u8ocpKhPKVO/F+vgFxkLP5wHbyg7z21YH4ADmhg+fRmCiMsuN
1Kwj64TxHQuokYjSej2DkXSL7k3hy4RRuRr6dKCvFCUq1PqDD8LRHSSA4JwC9HeuFVlvZb9qGKSa
oJY0EBPur7vD3XwgfSgPFFzPiSU+ERjcnJMkGU4B9clu42+H3GwsT2AnEZ+dSz4XBUhArybNiqed
KsljRGcdrQ24n+1k4scXdd9zV32ujiUn/C7uxaWZa2sYppX6YMgq0aD61XkOr8IWeCQQzumkxeNX
rGcmrJWlMjsiat5cPVoBtJZRkagMTs7oiuRlaVC2apcYj3/P1Ycd3eAvuE8h6hUmT1o5d2HrPU9X
0+XcGZ3iZTbdCnFncx8hSrgRMZnxGaiNNeWGq72xiiWYoJI/AwJEyUrZk4nuoSAc/XKul2nq1iEv
vM4lsANJvmVF/pPHVEqQIk+B9tpU0plEPp5OWVFYcaBYrVtLXdiOO/Oknk+aKJpZ2621pgwkqp1H
MRbOGKwBgjRHaf5+ZqbILoBJpL/AQUhmmdMJXsSpfcJb7T8TYkSp5+YhZGw35Skyg5/ZjCQ4jPOX
RpjZSFsqYOGnDrK3aL/GwqVEm/fSP/W+SCST1V7KUUUHp5Sfyy0tOoM90LsDBhaJUWMlMxi8NbJs
EWiLL+2oAfuUnhvkz6WUj9x8QPKm4WxNGCWzaCH3EREEiJ4JJBaMUpAImCTN5+hEZDFGWU3a/kFw
RMed7QMHszcHs6seP5PpPbqtfoa2VAVUeWUEjWuizPfexlwgSTcCpgC5zVCQslEkW49gBIhDB6i0
QUT1cI3WFHVAwYzzIkgTjLFJADG1hgnwwMvicZ6lTSqRFjfevUEdyGBW8hYvTyZrNaLFGBA1mWnd
tZvPXGhPcpbgkuZuQtOZatSRiEamOmAobyJr3p8ngI4WSdU6qZYWOAv4GIDrc1ff+bo+gCFfERy1
D+b8PTpSzwreknFAzvkWmo0yAIQmmgDBLjyTji8lbM+TLNHx6tpOTXZNXwCMIkuTrCOj/oD86DD3
q7YwAro6RIrzxC3hfgXiJoyn1Ch4DB/s3b/HydWB0PfgyeH/QFjjKmDp9A95na+caSxvSjTME4zi
nFVovmGrORc6N0obPEYLYMuSOmAEPOEfa5Bm4eEuFP0qvWlIhmz3bI8IA/dbSg9VfgPuh22Z+RdR
Lv3ii/1CfCm0rGUl2nwprMdcNkVLE/dOJ7TohMafB8p9hZO1ahsrFk/pPes7fOSemclWFHhHJb5H
VBmIHPrp5fTlj2G/ZHjdP/COdEklIoiqR1I/yud1HoCoUTqGAfL8i8NXyDHikp4UvQA9+TjeThpP
5s35rpTtgOoJm90PavjEE9dB4mzXYJUAkXz9S/S4RU2PoGhtyuBFBxFWYAXsZTyARIrWpF3wwUyN
sRJb8IvAZY954XOQ/DvB0nHZkAJpS0/UqcDsXfIFXlR9FEkwQvQeAB0mpkxBVwGsEUt2s8szCnf+
LLF+FHeGvRpHDBfsmZUzBRw3g6ELsvJuCbX2XuRwG6fkgIMn616u1gGnYwYr6AYXPazT1aD/cSgI
d3U/z3hThVokDif89+iiawYdIH+3iqd74NiQVbOBYtmLhyV8l7HG49s9zLSzPxyHl6gQkFbn8801
AUfpK6xfZ+khtrKRGW0qpnmW3Zpfbnl+FRqgva3SIDFOHjKNWH2vh2zMMgqaIQ0JBCIPXZrlybxP
3egSSNlCJ3YQwWJAZxT2OwBHnYUTORUuiFxr08hCTtV4G/VohsHRWpfTfSS5cPdL3XHp+1x8mxjZ
6lplBVNnw6JV4GY9uCsnJ1i0EzYes2Y8iiugiLbDyWMLIn42yfTQdtXQI+bZJn1h4SqxFyihTvg2
gZkQ2ZzUY61vekVbyYMl3WY3befh7rxdn+02rm/6qPbqhmJ9QGoVrpOWFNf153PrKNTE/mc7Zi7D
9xk820mIzDtO+e2kbCNvBwdGRwLi7SAjmEaM6VK5NcMzdh8ymhovs33DnVFouO2bgC5Yl5uY+bkL
MR9cKnpsbQ2+DixbOhAppH8lYdWJL6i37YHaQX4CJydGcQniUtbVzGudnkD/5lTQAHS+6Vm8oUoR
CGdEUDIhBUdKW2jBsGLTVgTBsQKiK0X4Ni4RvaK6qJVvabpKUwvwExWkJ4O4rtcZJXgv94kTeNJ3
DYoxO9ZTBP2DoUG/nQNn6mA1ZVatJQXH+0/rx/OFlg256Oz901hP6DO3R2TJpvPtFXnAEVNJqdgf
zb1IKK3oLpZCc65C45tJyv7Pptxvx+g+9Az/CCYXaIntUsWitJ129OXn0O6BvtrQ65VSQXVoex+m
s3+/7UhFjQ5tCisPW9rOuu01AIT1Ca6nkJaOYNJ1fpVLsji76+knoi7BcB9/Au0FxhKF4nn2Bkjn
1wTUtonlYc8VhioRdaXOlw7ApvdfHyGyzN30wPfNcHd46r9JQbKzEu+n3f9S9+tITUynwf3AITN3
4wwoV4E5DSofrpRTTn+Mcs7Bz8zUVEoe39SsSY/ZPWpk/YKEoHMh0NOgbol19sofJm18Qa3xBmTt
loigUaJrYjVnZknjqH0yhNzx1cppZFpdv557cPzPCPrPlfv9YLErGOlApWHAqWSh/l5N9kpBKHXX
GmWmPtrjhQhSyWBaOwXGFuOnqgQhgVynGQlbTPtABh3km55qaU6/XGxk1FBSZ0VHZge7q9PvIdsl
tG8KaDDKbJ+UTZM2eeJQpuZoQ6g7Fg99GLMZ+vFx2sg1T5s72mxzILs7F+LlG9bNR+nXjqG2Au62
KvnWfHndbokNN40sLw8PYCdn7MMhW0sbXLjuZeg446d1rklvCu9bCmXn+5KKQfmOBNEXScakBF7q
IBOXOyXRng/pxRGIBObjMzMsSFADw/4KdpwCKm+y5kUg49TUjy09VOgHpHkqqGJ3YFhpMgVQn/kN
nZ6tNmWZt4vFZnlLcssIgCO1NZQkBXDAMKK8QQLImDXLtxS1+7z5hQZeOZalmW/bw9Li1GDKbr0g
iS+v2cRtM5LplGe66V9RdDyUtgaUbuO/0ObheWqc6u/wsepc1Tzw2XAjcn1NKX4euoNfVpOSbzJJ
beQBbo6VWD3LDnE1uMLJFf8tYMpPkjiPdddQlC9T4lLxLhKjTjIcoyrlsXztgVVYOFvOkQNAZN7J
4R4g2jESmtH3s0LlumjxVZtG2Ch2SCPr2+VxeYhL/lPyTRPWItVq2J/ZnlNAG3Fpjagr8BbUpVLp
w3cGFpfJmjfvga1FMhJmw5m4QhX0NeqJ11XF3q8ha3UaPYXl/LSPavKBEYjDsdw20qgpxCLaWzUu
PE/0V5c/UulNpyeWYn23oBEboXnvzlxRUyl2+0Gv14lcnvi0aTBS1sdXGLtwf077cae/UqsqaAM0
TlQaSLGoRkLwE4xCc12cfNBbzIlTaLbYBaSEZOKFctgHrznCIZGRHCt86WQiFUOROxdPkq1eFjTw
1+ui3HxhT2vGla1DmOibwZvDvDPKEFK5Pob+LY42VcYAKLJdpu+p65DMAas3guMyqvCcrxwF1B04
VCRFbAgZa7LwGK07LusvUFeimP6RYE//3lr9dthip40zeLm/jmbloEmiC90smtZHLTqwH+LYCCql
88Z8rY8Y7jmf1EkBw2UXX8DE3I0mm9O4mmQ+8/pIrPR02s19dWLSszjUca/PgJCqtA2KTrzuMf44
xRc1POze+DAoZUMx870DMEykGG0uiRNIlsb554/NcAJm/cZPW3nb3elMhBI5Hds8giX7a/BqfC9C
JYGeKVtWUXVRC6mtncIbBxO/vOLUxuLEb8mwjz1S19zPUeKssN6OgdQqx5Y0kel4lOeirOUKp+Ut
Luc/CMCADKwkiNuj6x45OzAtmy9+Lz+5Z89kCG9Qxfq64nTF97bytlCMcZDOMSGnOGLZGNR7tG/P
hTSX+qFlXB8/CkkVVpxA4QL2x8l0DMBXicL+33YjXmgZ/GQVxcZnWePaMT1bRFQX7BRTNKsABMIc
Obr5Q989VsnxwEX1V8YgirfR4sGZW/0qJt2HBTCPPkYidUFcPLgpnYSAwDu/iQr+rF66OyGTlotQ
lmcsx9ZdbFjTvyi0D7vZ2BDn97ObRU6hLx/P9Ob4aIp0BSQhlfJkPEARfee5YIIx5hoBO/Dp3HA8
+VaAiXyftNcBtW5NN/kFdmBa9F93c7TBXMLl4lO9VqsS7zHLNNVp1evQ/pm9jk3F3UhXSWEWW136
zupgEatkxiuI2jYaXDEPRJ107GBNEuIIM6Tcmq/p2TxGBi4bziWR8n6Syn7zuQROK8dOQwJ8w627
yQRrczWycBZej+e4zeWTqYdlIdFPHic9qrRMkvhsmVTggAjAX6eJBgyWmIMSyNop2WEY5clRXx54
Xn8sW9i9vJ8DSJUq6yxA3hI4FyGscofG34Nc0eJ3//XmxrMssbzVJ8zixHLXeN+W+7Ojenbxf5CY
DUAcyTUKow2jHuCHtq9jXdZnOiBMMu5kcslEZ9LplAEQEW88XEmujicZZC7XDEimuyUXoJM1gLqr
dZPexP+h6qFgfEjhH7O6pnp/AwF51/xKR4bQN0E4WuoBYmW3F1IHtSgZneHO8tlKbTfyn7goUT7Z
oajavBw3ZsxQyCUZZpDcIV/DduKS1DYzJA92rbd7l6BWJuQs8rsJ6d/VlRr++yNwUQwnmfMFn11I
PoGo2J23p6liaLpLaf7LWMd7Gm5wTUGPFEUnAFxmcg6Rm52SNjhEwD9EVlReUkooFT4374GMlktk
a2+N0K+JMHBy8+xkj31WKmXeaINJ5y1M2LQhlwOpvEZ3gxVTPRN+DSlLQNm/lY37ZeIrWXsijC1s
ctMnTH0yCFEazw0oSCexyVS4gOuaP6x59t1Qmn8lfJFe5X8+8IINGxroFY3/kbp6PPQnQoFOFuax
4ZqjXcXKjWv64lZ69mTndV0ntPGEYeYeuVovFkwXKuc+iPxhuwNFN0Lx39K9vvjdfhTlY2YfQSYy
gWWINgexCLdv3vYw9bTd5Az/bobXc//un+upTxR9ZFlYdU4Da3D0LEVAnAciQvUHR3s3EOZlKTMq
X9+UW9MdbMh6+rXUy6wDgrufkXmT34araKaOF1bLBC+D8qF0rJ7GGJJc2oMhQ0EdTlKoP53d59E8
a3cS1GdkdYZ1XTVroc27+Zw3zXaPLbW6ozGkw3AGkrGm0rSU4vAXO1wjcnxc1W4I6bfFOSZhyseN
piJH7CK3cCGPc8wEiIiC5/X/6sUExeLdQzne5OWl8Rta+oMCEjYo6Vc4Q5qDvd4K94b1/uLrjxv7
U4biV5wqjvA2ZeqYHPP3h4NTDh6uYaiwO5FT5Xwrt00oIhjLMEYWXaCI0oHhH0sZ46LzGLqQq4Bg
vyX/bYzRP03fRtovzPPrEgTSDqgQz1d+F7jpgd6Q7GMwucWQnRFcVFGRlHW1mdZsEVbedn3ZeUmi
bx25CnV4mQF7+Zyz6ffjO/FaJ+19itpI3PIp+hzscq+iVRxwqDjc70DTb9zDMO9EUw9B9sfP50Qy
r/eCZh6f6vrggR0YkJqh5XaBz8PaiaEj79iEKOp8vRBzcEP7afLZCL9/ZBt/zz6wlfoz9TyLJTp+
WLpstRG0OKWgRU+oHvz2CQ9wUZ1bRsOpkA4oSWo7l/Za+Dq80NwusPAY2fJZz5OtKrMblhEGDN+K
xvpyGtxCBHCXIg6tHlHQH7E5dVHZGFMEEpRXT8TFzGve0wgf0/sg7irrh/11CL3llSOzfo+gb7rg
f2UiGWt5nbrMD09t8MoverDBRXcd7Mg/6txlq7iD6LtP3sqLdlvvbv+ftXa+lCXGIWxLMG8D+Rtj
VGujy80IKxkTs7BSZz4/Sjc9NGna/g6iQJOt4fJvUtA2HecaZDEVeV5V5Q8WQo8FW0dqpoaLQ0ne
1bTcmERDpkZQClWR0cEYRniX0HDfLWBFQv0K0eL4SBRipymHyyrxZEWrZa6KbGXkYvqsMtQBDAoi
qZyk0NCU8lBjM1D9dzCylrFcfiFKgU6SxG8oEAR1ozt4dCP4+9y6ZBxT4WNhtHJkTv8oviTkcETk
akMCptudcp1IcqnUuJw+8tEeaqefSjpGeocCbHZ7x+WTr0Gwm26K7lfWF9QolgY7IZWayYraUnUO
+O40A6sx8WG92bCg50442CMucyzTyOuMEj/zNwTB95VQ3u+XmzvzKNYF1NCnIwKpUTIS6vQlqMAR
T1fky/SG31VHkg+rDd0fgOeHaJeyxBYQtOZtTf1Tx5tUe9PDPfsBFojqxVmSqPwW4YxF0lFV5lUo
MEd0Wzmz97CobOkjctANEp7bsiFSX08lWWCZpzFsI9wRr+EBJlFGn4GvR0oD41LJgrYelPU0jzi2
RY1h4tWyeSp641UisAKYID1maVjDqk5kUpUnIEhnmZeMo+3pe0VNfZjAMJCSFdnUFoweWQTM8L6M
R+8vcdiw/JLE8BHzPZsu5vAEK9mfSTPGMLVJx4ESx8668FIpkKbGnZIU3+8nQ7ZTYfztUKB33LAz
434fkrzEKygtvE0Hu1Shf99biHUWHopAwjoF6Emy5ZtC4W047u+Svz4DiKFsFT20UY/Y703F9LuR
PSRI4O85BzQm9mxQSzMv2WeLpDHvsuxBKrRqRUW4J/AkFE7SZsBzxquGDaWZfi9Q7q8qUTLlGr54
RSiU/7l8abmIW+LAEO1RTxi94AOtjIpfXAWGVFPEUJxeTQo0U+ejJlMxIVS37FkkSnXHM6Zns8I6
IMqz6WJKFL8p6khdB5N49WZKTjU6FTSS9SDiWm/WVJo32Xbv+E5ukFYXJG8SVGiyAYvBsPOVtVUc
/mdfSh+3EJQ/VXkGZCG9MAh0dM+ZO/NbC+hYWfmfPWl57fcH+fn0kTmaj8P4+yZCmA4fMNC4/T/y
mdHnI8rh6cbZEYVMJhY4qmcK4B1xrhV5vIADkzrMhL//YE3ekaI0AkxiWdg9U8mY0znnjJmFWMY/
jE6GiCQdxRmpd2G786AzSwx79+zsESgkGYeZXb1Xw0h0QwJ5DntoTMdnISPlOJbadvpXY1DeGWDK
41lmS8Qyu2nLZAoCSOvDJCgArLDm80r/NVwJDWrw3HQEpWxAcQGpXDqTv6AMQ41h/mOdRj9UK+Dn
VCQgRTQDiLEnQmJhnpez8CgdhU7P79GhtvF1aKnkb3yJHB7XVH8gJmGQJh0DddqQVyG4bLRtKDUh
nS7qqxCVYgJMJS0ZGxJ5JiLHvIE9JjUIE9SzjNr6OPxhuZbNVdjwkavy3OHnsrpRNyW8BQSxY5Cp
/b5IJgPQWVA9jonsNDWvOvIs9FNEgk2H9bL/msTtY+6VaLz6eG/Q+wMgRZOtw5PHZ5io2RbrUEEF
MlIzFU8sS9OxF2fa78yMBFdbHms5yuy/FsamJel+/w5q2AK4QUy7ItyQEaFiOXmlsa7hrexW821p
uGA9hmi7Xkl5duvXI3YYcgTDP575zQ8WjFwZ4H/PfW/S5LlgN1fPG3NvttOLK7utQPcTZDgbIG+L
0h8qJ/wxbTe5cQmziGHdsJ8AkSiDqgzj731SoasL8oNllzfg7gGoAlJBOi0gTe+b4uYxgwTgrE1X
tmQkvmA84mNZoS229/OCDakbCIKTHJ3eWtZe58AdgsrDgNiyyIw8APL99hNGTd0kwBsl1W08Dt/V
Plex27xT7+R1RGQalqZVVJ43D+vvZ/1koYRSkd3xJ9eb3i1dCo2LxvvGcCXJOxPfvkTr+/Jt59Yf
Pd8FxKWjoqufEvouE/sLUT5n10AtkaFplP2WWSbrAiPcsxgka1wEV+0yCFBjWanFCgIsvSJIGkw7
il2jX321Y5UdZ44KpaeCDoChA0Dpf50Yn+AQTLVQ9fGNfcKcIK7/MU4dDuf7Ac9BepjZ7hDhqu2R
kqFWsMNbKAc08h58Va/dwRnm4zIoB2hbcgd4SLY0pvhGQ9axMLh1hfZm3VDB5WT3Ro+ub7IoKJ2Z
/96mffRo6hWQxcqyPJZCoU9T6WhHwEiSB8k3z5CJbpPRNXyoCS8Zh76Sh2GlTYeSnv3PGOMTg6+I
qqgaRRsbGvC7WHXVHNxJ3Q/TZeMNGYn8f3s1nYIHtUctjfWlNaeoWkn8f3gs3LmeN21FQa1+XmOj
ToQqEycj6c+ZAAuWrmZAQLi2N/Ww1KF6clUKCkErOuEWVf18oAo4iwX8keqz7akh6ngCtbfZjDkt
8E7o7lL1quKRugGFG+uXY8KAjq3xeK2xbvLBosvXZwiTIMaOgh9n6D0BrQxxjNKsEloJyv9v4/ng
yzloMH1vlpTXxdT99ilBX3vvDxH1QHl7vUzpQY8Tnl4uk98ThCiuWUM3dpFu6RTFpm33WhMVkb2l
nSxignSK9Nt0m1mzZjbkNaMnJUinmFzmP1lg5HnWRF0dcosjfgWd/OW4kKbvtWvPcJIhaeTyWv6f
oXNzfVQ0NO4ypY0x5RZTzEUz1OdBMaa4/q8ID3WdoNaPnSBIqpcU951gBz9HamRShFIoRKEiwiGN
JbPIV6crjF0oYOiO/5IcD4jvG2yPwQo2obrhE6O8oowMd/p4iCHCPyu1IpHW92CtsTaxTGdjWWTQ
1K9XK5VxmYn9BUdvUqS0Afz1OWW7zGhlicbCHbyrokwbBtlpKS5D/zzfDUmqnb2gqGJTgj0AU6wo
W0dicyruhrXs/0dJyRIJljH8Qpm9Ow8xzPpyr0/BMnrWhKdVM8Jsn6mpagGdx5VvVSMLLE6bmXON
shYaY5OTP5jVCEM/iUTMF5HcR5V5fg8av+VsrZ6ZqtKaS3WUdGxxw4PGd4DYPAaP+1y8KcM523ls
v0Kvt4y30TXt4bfZMfoqZJylEewYTP5thP59f7OwFI/LTvxXO5a+5wqGAQScQPSYxvXdajKVKxdw
9ek0em8Oh61JVWGGcjVp9zuezagZlj8LHBlSZXsrrhKilwToYq2okMpJsb1Ct/c6I3L5BmWSCbGp
QArGSe6k3VViiYWboiNnS7uO59ledze3zlSS/A7s3nQGpBGFBSIFMs1+NBvshNl8WdOmPDhDKPKk
mYLKkQFWCqBe/YfdZ5Bo/wM5qUZ5MlPnKqRJQ+RHL2cMcwFyb7OWKHztIaLGfIxT5InhGTRiDWto
mWpqcYtk5GAKiXRugW93KoLCj/amKT7iqu0Q7zI7oxD3e2aoOtMvjTQfmpVUWeVN7MD7tHKDxjtv
QKgQPPExvLEKSKD10DpJeU4b8rlepW/CiU599gxYsU19grdz6qhd442S4tEuGQbsfRch45rc9uCG
5Ndc3Jr4Hvh5+4HqYk1wxJAbXH7R6N43tJEAHldLo2nVsEonmaYvUFYsmN621oJpTMo7InwnnZ8p
bIVIDkRmXIScROEeHCut75stBWNHDd6M7SIytqGgQ+T99XvCBAWES/nIFVthPFT2T9Wa7j80XEXp
AeHLJ45ZSfYkygHD6kjBCUo4SLJYfxy3Wt5n1NJhy9G+Qz8BiFx1Y5kt9uARBye/LSwq45JWM2JF
87KQ0FC/7mQUy52wGBrmDK7omaPj3YE9KzW+LyVibQoPJsivlyFCAttfdqKFND457lIKv5FtOIOc
0wwNh18srqKXNJYJqi1KjO9klZmW6NTUu8TIck9p9fRABUvwQh4wANwUz0144Lyqux+fhWv5Vwdb
c1MrUZuMyz2Yj0fpAetCLlHkAlIouZATEujZfT+ZpQIM6HmBF3ORLOkd1HZNUINSI3UsHjEVOC7L
DZOc4/oVHZupJy/pFufQeMilt3whlHWZFisy0L3iKYfsQ3KZOgVNpI/RHsOTTXoVVTudKeowNwSL
x8C9cZU3WbiqdetCjTnkRjprSH3NeAbuni9DZNshA/vBpaozm97tpvj+MBmOyV6QQKVOH652r+DC
cduZKrqiDUhfZr6poxlBGMxD1nr6sIqO5/ylx450mFWYhpyYP+0i2PD9wdb3LGWIlgCRV6c4jSUk
9o5lXq5DGY/ak6/P9oUzKl39MW0jbZWO7NZ9cuShJCBOZrSOfdV37r+6tNyneD8bfgeVV83TQDsi
EGdTOrV/kCol8cxgFP0DwOzwIqNNAZVduAv1FnEn1giurFrxXRpgniSO6XtZdsybI+cdDyEnLWTx
WRIWXstRPUrb8MU7TzTC5ps3MavBS8gUOfaDwoMBp7KH5KnPtfInT9/HgtpKE+oFS4a95j4gpCFF
4CbXdL3mP0rIG6DFF4hrsO+7SaJvgw95cn4JmKCa666YGqZhotlVsYiCEyUIpgPpY3xty/iQ427W
KDn5FLffRFGqbNQUmKL4zciv59UWpFpF3FJZpaI+FjilFOmgzR+XC0FaP/Vkl8GacS69qI868r+1
vJOXFEIjP30bveaywfeBkbHqQkBwo99C7092FuFrfUztMldMi/eit43hEdQPJsxjpRFlyS4cJrcO
O7nv8+nwEmdj2DMG5OrukQS4XpVrxuqBWkgp/c2hGcd6bqcClXhNClhFLwy6UlAVkF4+mZp6eYjV
dsJpjY5NjXogYRBJ/FFABpf6sesvedvDeFkeu5tT/5d8SLldcVHI4kgfv0k4LIcVQZ+CF1Kv5ZGG
ge/ZR+DsSWNlBkj6wYOHXZvLDYYiD1qhCshp4svT3AMiedSFisXtgvqSDzI0UJzZAdVlry3tsZvY
J/XkhpL1+44Mr+H8oUalTBr6lMco534YLvY+UaFlkcaEEVXxCMUy1srLjW3G2cJ81lyrhTKTY9nV
jskOIs1/0CYi1tTxmk8BCyjW3n6nfBO9pxpIuU+lIaR2m8N0wnOuZ+gcryVmHieaZLxhRJ2zsauJ
+5XyoE1+/23XDfp7Qz1X296lJwj7PeHJU0KppgfpIiRaSKzewlKhH8WHnB+EPsNGjPtb+bQ92Buf
hb03ue8C/G8osxXQWXmUE8/wkGF6ugb02NaVe8dNVqviHUElvWa0Bqp+ur4mi4u3b9kSTTV+3Cuh
w59otAu5tYqwRQBPZMpDZUq3Vx07Xs1SgruNIoimuFlWrxHxjxJxLCl7JdYv/iwFWceFR8DJVUfI
Y3Djxcbgp/FNu+JMnae819XRoS7VtNgwOxdhw70AZ2qhrnupE7pNOuBAHjAJzsKg0xm90WX+iHRI
zcfya7ab0xl6diau9jwJkLaIKYC7kKbvdsNBw5jM03/fJvzBgdEhF3mT70QWcj8WMqf/YcaZEKxk
bN+nCnZ0yITLm1T00unaiQ5ix8AVIjr7j1J1cPbG8gFoU+nHDng+yPJNhLI2VNhHH6W7POt3tO9c
CKhBIxcx8B1zdP4h1B0OF7key4j6AdOIf3WKVYXKnaSqJ7STcHLKOb3gtrUjdefYtc29WlmvXPBN
ZVkqX3DpkX/2N4v+XQo7YNH7w+QZoHf2c0gmDJVFnscD9kpuWTyl5AWcGLxqXVjSBmjerRjfSUMt
nO0M06jFIRPRxtQfdjzsBHbmentctBXKXsMvkLVYxFXjVz126hG3F/Bzt4KDPf6bIDPPSeC0ZfZM
ciZ++8kZdo6TNo6iKc4qNamB/0XFOQha6DpUSMNOue+cGaU5sl71/UyUGv2u2U8iUugH66Czfbui
QB42aweNBUNi5j4R7avZUnqMnWaDOoJVA/LnaYWcYOiVT8iSn95/eBXLuNIG7RHMHRM0FHJFC+cq
9GVwLFXVcWfaSgyVLwHC91k6oAJc+5sK0QxXpdRhUZmLBdO6mf0MVAsJiOrTfr2P4+OQIqGMxiDu
IPCXBtxIK304F7xmD2xJkZ+JflsHjdY6HRExNi5rdCy4HuCl6tCZcOF5ffJdXqZUjXL+ForXAvZ8
pD2m9n7h0gMlx2wilnLiuxqPtPZt3UDkvnF2FsXNNGLM5JXFUqpK6QOkevvXwygdbQBMKBuTthy5
0xjp3119f9b+PBwYQCm1DcB1zie2stl4bNEBAoKox6P+BgqzEXTkdBHIVONZMImBdt7Secq9Owlo
ohH41bPJyCQBNt+G3/7TJj1sMq+dBxmq0B68Xppd/SkDIXcR+/ylBUPQ1w1OQSKsMMmfhts/SXbn
6N5PpDEBbkMKO0amf3b0TMOaC5J2Iwxz3Lvk+XZlVjaSaIFnAQvDXwacARvLNQqDVC7mNMNZ7abf
P7+jkeVnOhtWtIevYo+PgojHcfz9xnts0pG6ouBUNmmdkY9Lh4215wN0oZcdGwdB7TO7/jRd0JCp
+aWZKWZW+xG8xDqScvxlkz6fy2odgTI7XyXcaFQYfdB8kMyEsf1VxD/Oullw1bVBX4JOzdjLezu1
KQMOsG3hUD5e/ob2+sQWOxC3rYYlA/1H/FYkxJtgPWQKdOfDt6uWc/igJ+KyTRmNNp45/NttOl14
I6BI0LP3FxBDVRHE5seGD+ZEdcdLmynJmbNn1zPQu/BcH5H5oOgxjJTU13a57FoJ3JkAYYsie2XY
sFSQmOyghsTzxkfoYzZ+OYcl4afaDBRPQTkMqJA1Lk1eZACoHy0YZ2VAMjzmRIykh5ydordnRJzC
j4UGXSVNUjlRIZmHwO6SgJbgJVBTf4azUFa4tsSeaK82xCLtDRApKt8BRrTIXFfBfoMxywGGDUz6
U2chUxoWbJ5bDY4qgLySijgQEh1rLIu98KjpxTbgGpVecSXtQ6SFgF9fXZdUbV8JMwz1jKMbzdlh
gps74v/GnJ/bkCcMeIA/AIn2/EmoWCW2NKGij2A1741xrudg1we60OsEK2ItJpo1UbyPxsYHmg6Z
z5NR/Of51ZfHBvZQqf/BMqNsm4nXF63CVfVTK9EvdSFM2R+3OY+PgyCjZd0+ly4n4uRJVdSjkj0o
lA3G5oyDCvly/6EecwyMTw+TnMrusoXNy4Hv65u18u8pOpvH9M3yoWrDoPWDADO6QdOsfj6LDgdW
UFpiz+tGn4B+vK8kMnZjX+g1yXZPu9IS/PUn9rrPZm6H47FepaZ1ls589u7hRht/7fWD9fJrVn27
oqw3xVltxBS5PvIh5cFGNoC1Usv+/7wp/a8YqJWfNEAJbpz9FA6cHCStio3UoApAWxQUsZ8geVP2
/CUJsmUJvP2/kdNaJIeTlf5moqnhIXQ+c2hzB06720Fi19cn4bm5gBAe5nwOFsyFXUKtI3y3B5I4
4VKu7A5cAmLIqmpmoQqA4waSNDyv2B9t3rhuPhnJyWJ6wcc8XRQlR/z9FMnMBbsd9K9UWLl4h9oI
DBFwM0X0T6zcz1bJ0We97QJgI1xDCy31qL+TT+272oZpnSSoZ98HztRk00dG2BksJkPT9i5MBklX
X4OhNQtnX2yWuIx/UHhCAGoU5UCfaGrjmhhYS75aqM3W8wI0gTtg39SXjdn5vGq0bSstQgpioFbO
Ry+OajIP3HdO5KOYXJ4GMkBlliZau3XHWpumpclPvGF43qBjCCLDHAqJ22P0roRTuBYOl0xUCX7F
zmO/DtcmucJXsGdD2LehW1IcJL65Zi/Be+RQwZDhv+5snZgY77JF1MTZ2OslfBee5LJNH3tdRigx
FPstqLcgYOCkt79dTnaX4S11oK3S4Q69C9O6H+0ICzkeeAG5LUk2BYVySGxhNwRo4DrNLiZk2vz9
tJG9o4g5kd41ANTFrl+CBsOuen1OeeiTFaeILQCdgg0YXaqn8G23FLM3n1xVV9BBEjvz1oioUPfE
JUVf1N09gd340Kg99JHnLTwx/n56NULGpPL/jtDs5zbW78HORm0Yk971wh4Sh92smoOt9bZafavi
TlVOQyj/lZIlaJerXXKQblscyWKsHpr1Ma0Rf2e3PB1XvppmnDzgObX/t7X5AtXFuMNFRYeo/bl8
qFMFXWKfY7sagH5keeIcZsx2NRAlqteL7/FdfjlFefeDzPB8EokawM8pYXt8nAaxfvnjqKile7WL
t46pbSIZjhdKYEG9jbHJtaS/qQj45Kjl7oR2wmACqfSHAKijeGjQiH/T5pZj6n+kbZZpjp/biYPL
vmuUhwHDzxY6514WLq457oiWW0dOALwDmzdLntir7i0mQwfUsPv/UOYsYH/OUVXee/GyxSQd4Ndh
3FPM3Ie89dNQC1lZ6/S9w0YTihy9b6Uf9ZQ1dZwgysNzbte4wlzyQ9bmGJlbl89STVgK5M59UHa8
OX4/m1BZ7AvxGph+4NWRML0Aqcs/eeYkLhLyDAXn7311StOTHJq4dnsT82uF6n9GGkbo7esYNPmv
W95FD4TWgyy42Im0e7qWEpLWjpbzoJ4bGGL7HpR3jZXTg+0OgHcVARM/zOUt0yZy66tMl7PEtekT
5S6vJhiwH743XuInNcSEiODYs8toj1sFGR9VeM/908p9HUXDkhxon7ROUcNIdGpNmPtxEn9zWoBz
2rvygPw51MsRtm2Lc8UByDZaE6tYOMVE5bucVVDYyiNkLmQZqdliNHz0r8KudmCHWtQUVm4CcQDd
Ke86tHFzee6sJWaW+Wdxc59Qk0LNCbQiD7MVViZNOuEPT3wyDwtHgqd5kyXyfZG+LVLdNVmluXnF
3fosW/7DPd4y0XDNXv1+Iu4ZtqvhC+6FemQUfiDIySF1pgLKthy7xP700Xofu5O2fM4TG2L6gZmG
NB4J/iV4SLgLvdsKMOPL33hi4ivzURlOX0H8yS65HC2ABe9JrhG+nEiznuD8Nbs/QilacTeWwus5
JlftYUaAqu51IVEIvEvgiLwUFX4zz1D09Y1evmkNg0bHxHPEIZ7BaJQ7CfPfhOm3DHwwxcr3vnPO
uhEBaI8TtzMeR6JWm5cN3OuKphu9ko+h4mCZ/k6x/YJkXUtFfBFCXlYubGGeSKXAjNMRB5GjHdHO
XcFOcYO6ERMYlIbNEo+Qg8MsBLbLZRehhxhygAx00gSDHAu+PmpPSy87pt8BQcDnlfI0X4JpVrxp
t3qz4pVdGz93V6lRzncRgxhyJajmrl6G/Bhtvo/Up3fb4LTjuoHm7RR3ff4SZJPR/fBB2T/CdMsC
iDUJ5DrpWOhJNr5J+OQecdDAHuNkThGwsdznFifpP6Q9pfgR73xz2PC6qr5O2toATIqOJ818KC+7
+YJt9VUzGk236vGR/0dotgorzM/QqocxxUugJAGUKXGvQHQ0e9VWHOCyUXo22/OmrZrclIaKLjLt
DiWiz12ZkD7D/IX1bsqfTDpbG6OP9snMi+1Ftq8fWRJhoaUWzztMMnQkoVpehmw3ywkX4GqzD6nJ
c4XOPqfCkJyJgmryIB1jLnjdtZTGTNUSfKkB0KZb+J0NA7IRWHCXoBFswnOvmbK3hRG2hhcdTyP5
PIJZSJrd6bveg/i4tqTykiJMcZkcPHD8gMs2ivXppGi259EpT9BF4D7RRWdT/lLwV3QQedecNjmG
zRwONaKEiWrP82IyYJo3+H6iCTk5q+oPd9OPX+k8fROIOWH/Fn4z979uBTF0qifEfPoEQoD/pA8F
Cw8A0GmfpNzo0cvL2w0YlNxpW5chJur175MhDyzWb13ILRIFrDgTlizVLjXaofbSM17XWzYT3jZk
w+0c6+hMxdHHM+5f2Krj7ADLglxrTuwLZcJ3MqD8OPJO+/bhbRH7/7wYN2cVfC6F9iEOaSJcDlp5
x9m5vhJR9XcF1THM5KXjVAzZ50rAvdj+j1Uk548VBU6/i/HurQYnR2GrB8H2Iz89WDjZURb0skNy
g6+FzPaE7t+2FLy+VS/sbNwtMgjPDc6xRnN+eBEshedZAu/XpEwTvTGjy+TDN6w5jVk97SectLSr
d4CBClWOnlceatKms9FQq52Sbw9j3LvdKz1QvlkazJnnfuIwIm2JM6gR7ljbcy06zvkle4b60heG
ZmvfwAWFnGlTfmYGQDCAALaDp3Gsy1TZlfxleVy+2gBdPTCJ8CMxpNbJSrPAx/i0A8cmuN0SJZEC
MH5HdEvaC128SrP7NCbiprdT1qbMR32xV+BeSrhvvD/HSnWZ8OSc0S+dRn1JsOEO3lmDqqB7pp4H
s1LQuXAUUmllNce9I8T59xsmBuljmGeI3u9vnMCVRZkTWRB4OQfhYQ2JYpqTLMemixS1xKhFWeSB
frI9NSzl8UZqHWoY3BopANK7ghHwhiAwFHvNV99Zm1dAqLYzUkjRqOrFK5IDeTL4dXXzyroxEtwA
9qzfbKfyz9fo0Wai1O24yixUPsG5cWzenlimfM1PIyWRqADZ4Aj3qvIgyuCBdm26DIMxuzFWun6R
4GiBu89D1akfZ1tr3UI12EdaUwWazpSKle7oKMegJNOBMoiep+ytjKNiUJBJBEohOXSNQnPvBjKt
EAzCFcNIaRqvpjem3FWC71axWRpUrYp32GefMon5yBD+S/xbzNJ9y6q+l9+29Pvt3r0+Z+Bhr1qO
UUvNUNENuyyCwV9lHqAf2yllz+hbRjph7RMt2fJgUpgbpGdyzaVDwzKSL1ab2M/FrvHzhKq50E/d
L+lhBDQNBfY39c1P9enM3oYOjlDYz8Jr9iBWUoPKh++ynCaehj4pt4t+yaKheufGY50FAbWWP3z6
p65n1qYHOqHkzfzx+SyJ1X/hLHyzQYfz7K9v5Zv/+cxErcCcC1egHfGR1Lkzv1rMITZDSYvb8nZi
HvOXDZ7fNshWMYXL4AJJetp52MvsBZx04Uq/Fc2PQmDoXAvEvDbFNnfBxJylQl3qAyNCF1DF28Dl
JtBUIwmmsSSdEOmxmbKRnDujKuzUYqei40pDgsXLAB7YN+mKd6TJJZ9qNx9WlqKh8hMBtCmVD6YK
IdBQV5X3Yo6mwU2/6EeyursAnUVkrvywiG0D2jWOSc5aHoMJdd74IZpWE7lPNLN2kL4IIUF3t0GF
pcKW6UhMWFFAQWYwXxdItPjsBfbTk0s0vwdD7S7Mt1DtEmYfPjMpS3sWDK1L1wrwmEKmwW4s2cCs
dWA9kUrh5NFF7MStcgl5bpvfgCo2t+Fw8bwaHQQWiDc5vP/4jdhGnu8eNJwO+8X6MH/zODUrtHQV
XEl9iajmyBecRFUFz6oYX0vj/DBP68UH2F8pH0zlBeRzV5/iywCnfw64mmvdDnG4r56WgoitmIH8
htYwHEkF/HIyw8X7j20OrYgYAk9ej8B27tpmlhIyBimvD7Sxsb4c6DyJi/n1sG0Mtyx/itxJY1m2
+pyUYRHFzrs2e3sDPVBsK6yOmQ0Jza7y/GEaBlflg2OV2KALcg2s5T1t53DqqPswyQ/TZx8iG9Zg
prJZxEcVSgoQ/fWkzV1Z0GyS/PXPN1oRtqtaHlWZHs2xJZPAJaCSKHn1N96uj/zIbk8jI8kFGU+d
vp71jQxC5JElCiJxs2ZhcdJ4I2/C0pXh3Lf9Ca1d6PTcJgqXIwyLk97qXOkr2FQRAIqTDuRwch+S
dg0zhy85afTEFonAOF0v2DOj7XcVCwe4rOiGHsgZinfIsYmyFTP2zkGyrX1iTWHOKVXmHm88mvNi
tXCPmjCYiB6Vc3/mz7jycsENJ4HfLvFRw8Ydr4S/lGg8vFO8NUeNU+QbbI/skTYiZyf24DdQ8OWg
nVsxuCbCw8z7LmI6i+1IcssUPL1w9zUng2jp6yy7uEiFCwlPCWr3NnMGqu5MbY+KcYA1xWnpcxme
oOLQ3unFOWkOAKhOe9iF+HZG1gUkLCGntABqu9Uh3Kk17Uciiz3Zi5Kn5/NnDq6wkPqzcMwoSLOb
LBdrYRINju3IzhwU/Spq7D9sdonA/mZqIyL3Mbf82AF4OcMUACZY8+PNjXgNQvOm2EG/t/VMQfM0
DBwtmPTzCPaI/kYrSKkb2pKdvOa7YjBWd2+ehGtjyEsYNlVgqZ2120G+gmQpNtxlQwlfDj53NaOs
NghbeAdWBKW90gQ/XkNSwR3STPg6iqOxHYR1ikhJv25qKdL4Yb2Qf1a3fgpgwDvxkTCE68YLU/Ws
PtjRQkz8de6uqcqt5dlIIaZS1bEdP6c6HLjSLgfOmtWkFpR9itQQzZh+tGn8nY+PgZyZKJ8iv7gK
I7eXk7eIW4TrfSMnuc/ZbC7DRYeVBGaN1YrbnDGtUTjSQ/2ysg1NH8wMscd/pUgBAXAAbDZzh+mW
1j+WvnHVbTJzDfyL9RnmxCqTUFqKAtq4wx5TvufG8Jxrm/pgc/JwnQL/e52uuUcsD5hv68t02n5p
CiS9bY/2K1iGFXSTcSPYoIcSpmJnVERABTkNlNp8OaTsMKAk+pVU0iZmo9SHh+PHnl31s4JFMli3
/oFSJgqowL47yMrrW8ncRtG0bV+S1cE+zX+cnKi6YSvkMxn6FXy5pWWk6X1FS8P0cKzUIZ9zvZB9
O/DCFSPScqCCBopRXthMw64hZkmhWqsKBVwnHD1T9WTQ3uGnqVfbugkuFyAYZ0Iy+87iBjvCi/JK
uCL5WZzEybRm/ohzD0nCCvSHPCBo6Y0vDc+p2TJ/gUTvPfZ5zfP/WwLA78Cswx413RuYaoMfaWHK
ZCEH8M0q9fQVtpN4UO25ZOmvbCzcjT2R/ItW+dEJdAZD1ZSt4W/fx9HfwUhHgPQbaeCs2awvV9pj
5ySNjN14i1whnFv9vAFZ1ZZ4XN0GvuuS+PgT/4Qs1L0hG4V+2yF/zo6c2bYd8BTMWEZH8vN2SJI8
SKTyxOC8/nfPF8yp/6NqcK2NO9X4wUWkqH0ADUBxNOWe0tVlscgVd0Dpvd1WvLtM84m5GYpbpxX6
dpeqaszoF78YzAPWh+m7ja7+vEUd+cybppNkul/YUP1HvEs2nJ+d+k5ZDkOS30Y2KO/Kf0YvTI+X
hbdOfD1oBZa9u8lqivs+xK4EQxkmtttRT9HCN956ukJ65qdoWIHsNIbwlYGj1qwKtACydWalMoDt
tJK3zEKAoUFrh0m1zzas6jSW4HLISpmSvx7DajiZSpb5Aycyx5wHUdxGU4PnPCMK59sYQ/WGpwgK
jsCUM6BuZ8DKelLuw/Qh93mDxUWYipzPs7K6UGTGa9u6xu9gz0Mkxj1dPttOO/irIbu2jbH+ynDc
/RF7OTOOewneUWw4FvfbWXrpK8GSm3es8ANlCH7AkN/2HPSzxcGeZRsC88Y37nlo/5cBloc5zeKY
9hsBPthjMkxvl05kOHHNXTP3A25882m1etTO0W4W/R1BKyJD7ppmyftfLDg44AXJUsQmy2ytSHGA
sqDMwlhfoKfrdAvwVtOE827b+7W4E7dmw8QSoLifPUqXYXUnPUeictNDn74jjtzfzB+nG7/rYFWF
wvsqw8CZ8DyPKXSPcu6D66jSApYENcOC0R5GZO/9FRDdibChApebSFwIk1lc2NOdrNc49HJw95A0
QSZR6w+KRiCdXrmVGb+bt9WHytRNXD6f7Yfo2mB09NlC+DBbzhZUXXEQNGxBDEI8i7GdSQAYE76g
p/6g8UBQypkCJO9+Y8nHecBOnVBnv7WPxy+GeGvfyNyjsWudSF138GE/xAwCfkkOoh6vnpgA7eqb
rwUiNrDI8p8NtCWugc2gXFuMfK7HTrIfa8sopq269YGCkNbpQ1zG7Z+AmrItTnI8oUF/v447FjDl
unBpAE7RBD1Y9k/Yy2KNQR30ypogWO/Qs9aLhAKqWRr0p0hpGIEFLMa3MwSzZBeGfLlgoXp3d38t
3kQD1CVrV8o2U6xr9EBGThAPUiIhnhFtzuJIOy7UnbPZKbRVIGESXMwG02TINLrJz7QNtOKzsp/z
sdBrGjTsd25nY5gDo9pmiofKIIQnsgqIQ4n321aqHrj2N8iKyBbxTL0gcfoOoLyBqNwqvW8cLJhp
1k3L0jqulate1MoD2/Q432mz5iupMce8bww2oZkrXlp9cRy3Vg6pyRB/Cb/U2cU8vo3EdvP5leA1
suesh2+oQQxrMs1aaSEq3OxEXrriewbjUOOVEkUMhGFjLVps3k/nF9iaOygRfWHLpelbZvGmCMpu
bxK0dNjTC/tCe6AEZQnLnJZ+9G11JNfwZMaw0fOba7gt4rGFqJUC4nwA44uRZj+i5lQr3aAUNMRw
n5qMUq+37TWp/yK71IRk/C8cArHEUJ/4qAXhHSaMME8GTvcv6nLRssOhUypBJLNIHjnNAqD+ihCS
WX4BY9qv9zZwnMRCEE3INB60BDuGQ5BJlWhyscmZD0KP6em/Li0ZSaBZfewOpNB+XAClUmDTJnWM
h6iKN9GwI7ZPPzMt4dOhSXhdCVJlzgLcxM5LmyIRi2hQDzIhNGNXOWIB3fF4eyfxuB/pwBJMyOHr
zwm5leseW3nws4zjygj/CjHZ1pVgIn3Hkm4FCpO7ubesY1qktDK0TEsw/tYNVMp+h3J9fvdkffGn
iKV5d9FdF8rQm9FzPk0hyQVdLSP66de0f+zF6DWhb6GPXqdbH4b+f/UhFHkNrR3grDu+AqiTsMqn
3jZCS9RQlsUqs4v3cmp6WQw6uM33oBb7qezKX2pXPGIYL22DNUSsOXz4OxJ+OFFnNGAZcAJZsqsh
IQxIdDuV4pxRrbFKxkfq0sftwnoDZHx9pxfArPLSiaSM4RI5e+URLbbOlcFqVC7rWoJTkDVI4rK7
HgzDx2R7DJW0gCzb9QKQ0wvY9jv4GtMKsyfxVFlVOYDHU6znjbO0ferDVS+XxjFNOkKdcvh9i8oy
E1FRizo7OmFK/miqyu9Le0zaUJJ4xjlCR9HlN8LLKol7aKyb4AYHdvRuEmZhAdEBQc+wFkS0Bhk3
oXqrRrKmMHv6E3IonTmTfysfyZdJXr/xHN9iyOuLB4nwEliOMglL4YyHgNppdAHieEXuscoeGb03
dbNEKDmszspRI1rySJLUxIKVqBCbGWagHAvHPcN+xwmyFdc7sGw18Nj6cl7J/fzf3oO6HQoO3Lpx
idLiC2ayB1x1RtQd5lkejl/hv4q8fmi7WqaJlllnKufHHXZ2aaoN9qncL92P3XH8eWOJ29TU0N2a
KGrm3DgKzRVIpoqttviBIPzrRY7mGPfae7JE7ugArk+rKSi7NC4YMYKsBCoB1UNe/OzNZUr/YeTp
im05HOKW6C56hGbe/ZVkSFwglkqclrBBqZOWUDll/vY7uZowX4UeREHvfcyrk8zPzCKur0Ass0+P
iMqKccDZ8NLbUlrT65W8miTLuNKfW0td2PQ0Pb/HZOINnaLP/rMhmwADCNMiq+BAV3U9ESQNYMeS
vvRhQJjPm6MmWwEsqUPk92kORBCEibFitE3ANF2swED6sFlZObz8v+7KukT8Gn6lS+C/V3wpj0bK
N3ww8kG2/UdnJLaufjN4e4sP9BxxjAYXaiabzvSsMxImKoTW4VG+4e6FSDiqXNfavTMisWob9+Ku
KvBKNxQvbxG8lFs1XnZTZWh3b6hFg7xJpR3TxotqwzznxjL3a/nE+W2EOtQQr4dQFTLq1kxwNccl
xNBofn7iiI0qRAZ4c93cp1kN9iYlsYmmsHnPjLUiiabtUTobRLbOALXYHOt/tKZzA0wx7oH+gmIy
joZroAY/odKHvBN/aQctmIHU3AvDSbAfMJ1J/R661BOW2Q5e2d3SLW2Q4VTzX03GafqjQx9LpvBZ
hoAs/H5aDQO3icKeACl//pWYbqYxqApUv5aYiCOSr5ileAxYC5Eh1QsB+iqM2BxRLJRGGgJuUTbd
Xs2TvJTU8CuF88zAQireNMd1LtUyVqbmfHjRTHdJPyiF94Prj9F3mlsZx038lgadzqJtFqxgNvgz
kJM7q5oEuQXCF9SH/9o0yRc4xee4s74jG0e+1oZ9ECzITzJOwEZ1THQBvl23p0FXxgEObnbB7Nhx
CYJvg6AVxlQGxRcR5Lxo9nNxH2U1xWv4QnR4mMuP3Hj6+bhsz8IrdcR4XZ6VvTg3uX0tjnHpeGur
4cqgNykNThMZDBAmcuC8PCPaYWclhXMK6EJQ4H10d8PsSpiNFpeKt81/xMoaZH+PryIZ5GcX/jER
wj+Vx+JoBDhiDT38oThNSIKglCiyrNVnsRV24ceg9Z/cTy4p/vzeVQ0n6UzuBI8faJbubNTXuznR
3K0zo47lO8zZATYhyP/AtuY5i/fLUwYl2gKS6fEQcFpBfX0X7PhfIfJ2RADwpcSDz8hRDNfO8w/D
36r4DHVE7B5t0EgDBsYsvZz6Yz3D6hnV6uSalyS+bnTrk7Mhf9DXbBv+mNkQsw2rKtSORdBmkvsN
5BtxjasSfgQ6R6vMuuk9e7wGo5bhqrmAqXdoItJyTa1L60N9leoRO51B8KkW6SAxeyktzh4eghCM
+LkueM904V/x9TnbOX6d+jPfDGnDSCupI+istGh3fl1DoxJU3HbewTZChfSeFXtHWkrxuZCB1E3O
2nI6BXaCTyDvYch9IwE/OxiW1h8coxiAYMMN6tKpncL5qK5RdrPhhWJKRKhWLjZB806u/2sJkdwS
KdXniE0/CZAO9VE4Eu/2XVT8kdhTlG3gR9xIvw5qiDrcU7SZWAuwpwLIsDwocVfwMBxvDK0yDL/A
irSgbJYnTM1OdCkSlQ1dn4jRHJpEc9w009xfqQTvqFQO/6eMmWjYmR6o0UELa9NOrbv80ZPWG4q7
XmUCNqTWHcfVLFqG5NUZ9fg/d1sYZT9Ya0DyF9exvsMj8g4wxXZLECwk1TeDlm8MVBHho3x73gTT
R0/91Mnt5Hnmx2iJ30+O8OeAxKbB7gYHWJj0u03bZz7Py3AID6KmBYccUGdz+FwSSXq0yQ8pJ2iW
7lCIziq4MT2RIlzgKfnXal9hU7WpoCnJqY6MbHAnSu8lGLL2gTrqAZ4lpjTwd5tUiz+7V2iJQROG
snAzjKHRQElbfYKvZewkwCgRzR5V2ATfe3NI2AIwZAcQ3La9AU1UK0hfRnu13Fm3nA5pLsPVs/pk
NwrFrnk8xetAYRm3GmOyToHqfOSy2uNDdjNu7Qlxdp82Ni57H7djlpqRo5897sxUqUMWPjx/29WJ
eeulGZB8fPUa0Sapr4iHyObWshm5gwSjxAv4sqcII+Z2w1MVc9qL8DB9PRtqNKPi/+ojL7F6/Znr
a13PsBJIXN4ICckPqwT2+McsUThmicYts815f2WCFHuXw21ARmTacW9pxLBatImDarhYTmu3HaBW
96cbHkLAIahyINIWe3PIG0K33KNI+/sv038fnEQCAXDMEEVXLlF0qlJTew4xJrXR7W4XuVLVYCFa
pi6InNRIc/hkLmfHbW08IsM1FAFJ8SKSmrSrT659eDpQsps61gcSNdyZH4/vjP43vC1uOaZpEGp6
UKq6vK5DmVcAeLTbvVVy2SaFgzmPnwEnhd7jPprIgMiCmmoKVsWNuRTXAQeIXbpCJJwiRi7+WPmJ
cmOJPn9QHAzzAyKvDmEV3JSEOpO4R4peDjffuoqjiy5OqFpFh2f0TXhq3d39Yp9xr1c4EjfP0CVy
bl78Ze/a+h1Ww0xN+WPKRwmV326bx8Nqn5pigzfGR9llwD5lUxr7oFUVIwDmt4aPwuDMit18SfyE
Lfv720Qs1pOmY7+eiIpHY0x+kg4+h4JifGl7DFPO5vaSErz/pFc/guN9ZrsvpEaN8uIdl7sYgKcj
q4EkEsPmmicJfpTHh0nk/sDM6wVklWy2LKCSmQQ216KM5T1+L5dbuzgRmfMUe6tEBNA/OzU7C0A+
q3VnJOaID8lLTcaayvJJe3kDWt/lBVmtZ5bxrSlK9X6GjM3fWF7CK5/cb42cQlQ/5kKDSpxqFbQ5
eDzCBnvt5PgIyq7naiKkRlceBAfmk2OKz8dkdf4QbABrdjaWKfJHHZy/y7cjuT06GaYMjXLgfYk1
nJBtBgP6atTS6+dnWTpOLn/Lxpej9bIo7t013kwIlornKTE6Cs9rOWMZoiJUW+9SUoBYl20G1Awy
TQ2MA2TDXANhf09bcn8u+YfM+s8pcKhIGs8NBVP1W5S6ppNuaEdsoZ7zfRakvDkHAj1WOnic+kwp
xQYgIOnyCoAQwZ7/Exw3DPoAk5ZEBl4kL/rucc8YM7+Fi/30jf9x+rmm8A5WOKj00n+66xdjN1oH
pbnmFe1v5C5RhoiK2G4inXhcx4yQfwBPYYPbZYhC1MHVKR7Tgw89ikjlEelUla3SCjiNN7LByY1g
ls0PobaCyqzoP/8an0jXnNfvLI89eVVMjQwDnhNrgusGam6Cc3ajrDa/9a0HUIQqneMmibOLtl71
NsTufmrKye9QMbENWtgJcar8pbT+QI8L2a7KylpS+0z6Gb+/ZO4bslYKlLRiw6Udn7Awtq6oJWTl
R37bsuB9jBC7xGiJK4pWDCAgBEOAdiJgSgXmlhM6WUFcRM/nEdNHRcmcH2265U+u87vtorE6s70/
fomLsBDg8R65UDWgFJ6HzROq7q8hhCWnvIwuynrxZeB12mTUnqlk14dfZ2rRmCQ89JJdykgfmimi
Hk2RJgIgv6LK1sS8XOn/fyaXyPlqcoqFosXccxk/it6gsjGLYJBgEvM8svwO6XBKQ7smmIzjhL7W
np3f3TQrxhstUWmpfoqtsnYwYFHpj0GKhCBlFWBnuTY5scjlv6NoBMbj0PeGoUOfigLjKbkmMy5c
VD6VLMrq2xge1gnQ1ZjPhFEGS1ZU7aKq1lqYEyVP3uKAUdwUQCV+m/RVHQPeG8vHejJhzh4a0EyN
9VbEeynR4X4vucLRQNxQ72sxVdnYOAmUppUbwgTBdLbd5vAbCpyEdzKZBDMRK17Uhi/nPUlqZzqi
sCFWbb5jwOeK3nOAfly0uQdFKioaG6+8T9kTTTizT09NHiKlRWR9sz7AmK8vxAvSN7P1PlFS4NfL
kLfhKCaXPdJKEHJa3fvN2MwjAiDLPMkDlVW2ETcu3b3558gzvYq5lL8FGu8XKgODL1r/NbAy3/qD
YEAjbu+BTGFYeEwmkqWvB3JNkh2rZ4l4wDe0SDnli8uRXrkWUv4K+eaH8y8mQmKM1QXytMDQB804
5MC7LgaJtS15jjFY7ZDNQMNg1ePJR2C1kMUkX2Tbb9SYe17CHvQhuM7UNjvNN2gxj6KZ5qS1s8oT
/j2Z9RY8f6mrfvtoyvtI+S8luBe8zCvS5+a/zvQCkAd1k1FpuIZAxxdmeVo3pJkzNkLpOU3FtJQR
xRQFTN6I3WtI30pzVU3OlYb39nrgddNkEvdqoJdxlClmCFHFsgH56r8QMsAHC9EykBgQsKrUi3Ad
XQ/cj7SBpElCk/LDJmjvloJVtNhwT4+wqlAE2Rwbr+OJ66XKi1TpMIJI07fWErFZDAL3GPp6z/wp
OSUmy7TdyF6bZiEc+djStEAcvjBWwbkjJtvd7ZeXSQjsTQm5EYp84b9DytSyBPVN0N1SOvX2FdmT
FXg3yrm26ROOoQAVMS7W2G9wNh7dtWy2pXGosMKABDjqGY7Fh57Lxr4wV+WcCLHM4c20eyarKIVu
D/52EISFq/Ah+Pxw8ZoF6j+0wEotUA87g3SJneCSq514dkjtRIjoTq91b3t+d/zEAAUtOMFONEvM
VWmp1ENEWo2arzadaP+IshB9MeJPkeLxbjNwXyh3KEVcT4x4Fb6ZIob60ATuhvEBrB+iFj0mjjv5
0EpXYsVD0ywdm0EH0tjJ1MVUDWdrcF8DTFYzNwdwKYW3XLZk9zuPKTRmUUfUWQtGFJd9mEwjZcR2
0lP1RFX2RLHWadibIUSXTfhLRxEB8QG7XvcqqBdtYN2ITU1bj0fb4rKvBK50jafNwWB/5Lkd4qdR
PHbyU/6jmaYyAfLr212Tw2d3J1kb27BzAjm4w/Tg3Mvt4omMKU5YtWQMCq/oy1520CMPsaYg1qMQ
q5ZNuXKZMIopQP8khLazv0zDvYEcsqSpBYDbp0VXbrFYJF7f0uq7wDcvSEewX0fu3kmTPFLS5ZmA
Ty80553cU+Bc8Xv1C17EyjcaTfPY8pxvzdprFNDaG0DLqwVYmKRJqpWcgHfNESigvcpGuRaYZ2p3
gjku1DIu2NWZ0oaxpW1czgbdNoDUHFo1gHhI8AxX3WVPTls0qwBuvopx5xX5Ck4B4vTHMAN/O5RP
7lf7ZkrSi9gPvYZOtgrtmhcjUwqMPZL1TPHSkX8TTRjrAIfQUA3Y2SjWNr9rX6Gq9gVLZOnOcD6z
JIK/AijYGc9wKYOh1+LNFxpYBzQNP0yapAIyvUniNmz+Wn9xCGCRMAr1y4u6tIoDzfFCt/ihSwf5
sY3rkYX+T+dyIhcF1xVdzuMhQXkn4gv4ak1W07HVGQN3RgYW+fROLuyHIF1p7WZc1AdBXcSHJIIp
DpU7LUB/8ZEQ+Yu70Gh+w9ksw/H3zATAePqGbj8aOIeOX6STZPifQpyNPYtFeACUMoSIX77VQWzR
0x4EfgnpLGon4+qFn3NY1yFq3EtPUyej/Ao9aTzjmpPlCU3IzTcW/ps9lbjepjvgvYZzinSrp4QR
clNqK1/OKCnk7rjHBftnsPYrUlHZ4tcnJwbCl1yFNmjCuIxcG35skmWS5xqPcMWDHhA23H/SzVzA
Cl3lnnOrfoLPfS3UCCmzc79hwGszkrYjLg1ImrFUNIaKnklCmCNzzghIe0usjDMLYwUDowFHxmFG
ovyf6cS3x9e7Shlz6DDIfi5sY7XGm8Ty9k2zna1clkX2ZKKOZ3RL/VeJ3/P8+bclzQNlpugHaeho
rW5aUJrhFjqYlXawPDi6WaDTRzXoynNRniIzKmpjpozwXXba4/NYZkO1KfnGObG93Y27SA7zu3rt
jdTPn8xdf0rCKaUZGi7fKKaCnRGHM4wjDRnt8G4RDxNeDBAu9thEBBUElzEw3tgy3eus3jnu9+2Y
qdI2paQbhwhoBJ2uQAXHA9w93hPYyPJOd0+WWUT05N+iMmldQrldFIw1C41alH3rxCezsEGjg+0d
EfURiCs2mQt4ScGJkahcXc7/n7SzAc4mBu7AgBbqlctg537o2a1yHLhSKTN1KZkXkJ/gfjYLNbCx
bNCAWfP61mAVFbVOTfRgTy2aVCdsmpZRkisNByW3qySyErQSBBO8L3pM+o+L5Jn8XhQDPULb5KSI
Lb9m1okzoe5FHPHG0uNNOA1w5mJSHwbDqJ2I6M/MWmTM4UAAq/4Y4HA6Uf/OoPXAkbLILV6P5VSa
8duuWgaU7mpoWZwXrV+Mf0Zkq5+7kTWm0qdOP05oHJ6rwHq8c4WAzrw7jSii6nxSos1fViH2c4s3
aSJ63Xuim2tOzA/Pto1+vVjoOnfeHAx4HynsBvlcfagPQNUeou5aP/tiziTA0FXkSB/ts6irrm/a
nR7cWppO0Nd5qEmgMoq1Yj4CjGzi4wZa8lEGc3+UgaAuJwuQ3xQZn6c6T+HDvFTy+ee2NZ1snyUv
SJSKFaAdBWmQ5KSf7wfTwCWncXEqJg32+e30ZKtxpb9uVqgYQs18dzNyNEa+PrvHBR7gx+9CCV62
R58RXD3Sw77hwXqBuNkf8u+zMSctQnalC2oWYYMDR43+oCLszRVYzvtyNb6Bxqp0d8hmiBVJjZer
Cl70gxKvpChozSytkPxNuSsi4cJ/tCiupJQrFiIYTgdXP3xSFtGeakACpvmTKNbfP4UVa/1s8Kug
i/T9ZoQG5N+cj5agRbM74wSjSVEYhoTcoIPKwXxRGw/w6/IwmOvERotLNQHWqtusJRxOd9OD4cGh
x6GBMmLQw5Tq0RXTD7dR2Sikay00StwMWxXbo0KQdkBFWlugqUzcetrHEXX02fzLptZ/Oye2uCe+
we82e38apoXLgSmvGOjdo3ZElCcL5+WxKFT4mb/6CRRZvlJzm7Zc8EtleJ+iibBu345N6xIVzQfu
YjVApXvOMqfucAQkLCrobwMnXHTp1kTGcVpTLgE6N54O7i6vwGIDy0V3I3j0duyeOPjqMzY42w3A
0VGZwTzpcdVsJxr2c2PcqY3FkM23QR7NWaWP7fgTVwYTctEbRHg84pQGAgtnkOkdmbsRXKQUgMp7
r26lc0u4l5njX0iu9BCHuCln6Iw1/xhgibUoUCtb10C9Q/CV0oZVrDQI4wLwU/3rheA9wJdFndKG
yyZR1fmZP3kYT9G0oJkwn71V560dZ3ZD3nZpdLdhULL1LOlcA207UaNp8BRjpsPcteJJbMavHPCs
OaJXImhyddlkPwVWjeQGQEm+onO52aAhaKTtL+vaNG+ckn9JTSV3SEuzuoigHeteosNBGWqAu8t5
CiCcdqZ3xW2RMj3hmNcQaA1bVCjnNjOFkRwW1rDGooDw5aubptOiW+sbnvyYtD2EZHzJIJJNChkE
d/ewzvCwdxvs0En13h9c4+IVQolpYZjgR7R+4m2pT1DCuZ7d2u/KAy3OBBtEP/0gZ7MjX6p/UR+o
dJ+/6adw6dC0P+dLI6UZd9Br5mLXU4spF/3A5gPaUeLTb43zC4whgyLoFFhbxWqN7skyAlNNKDEu
NDu796vpi68H3nD/JtiWMlPgD+D+jTAQEVJa3l1ushc/wgi+3CE/d9nPdVSkr3YUUTEUGgmxvP1l
RvL1U4Z8enX4DArO7bKHd7QmXgrVLrXuE8nY+/ubmoDPb9ap1CKIo0zhyGa6yvZhdunvdGR5BPNk
qSTIDo2u3lF25nC+2FIaej6IFevuPl3nmYWXwTzoNXda0R64bmqVU66ExHfv9wnXXEamRYY8ET9+
gwXg0uGqv1FU5jXMXkYbqyZWTUazOZEOdgTuC+UjIkPCmyqsuz+Qrtia2oE0+cE4Ov0iwjOQQ79Q
2ToTKWP3ltv3kfiAnYfenOLTi/t+8zAqZupQy11ENGe3BW3VbrsNcLusOEVxzvQOCLl3ptx6y7G/
MiiOf3UyJI3FZ1zkpe3luVapEkmcrGFuR34e+Lpd9DpfLnnYDUF2RUWaOzjnkyQGvSXh4aj7zpqL
YCi+g9ZUWRgmODhecy0iY/cP2ewyeVWqDx5lqZgo63Nd4dlnjSGhdoYBEm1UcS13V90JtW7KFN6I
b9XVxgZ1s/J+9srV71vkCYLAoOvvDVYlR5F7t8c/v+3M3VcZb7/ABQGy8g0QPimTZfIw453Z3gbi
Gk3RPf9xwSXifxeQKpt4NR+7xPtUhYy+eKtBBT1b4Ps8W69nv/cpt7hHPa3r/xIvk1x1ocakOoJa
o/yrR5vrXfm4lsE7s7cktaQgKuNEPAU+O/5gnhxUCPz4am9QFDX0jwEBb0wVnpsgjhRH2N8P99v+
K2yxHoc1/zc4AsvlsKWI/bLJErUuqHLl2mUgMGreOzw9k2NmZxMjYY6nBzoCyf0GEj0MCdX2o6z8
PSMmTFzg7VnkUz6gHmmJowCC8EyvNSUCvUij3mn5P76c0U7rImxwRdhhew8FRMbut+DFSq9HlNm0
eWPCsDk+PUYgrlXKkzm2rZqWfbrXlavzCXUhXKGlRG8KneIjZ2idzmn29aay/mYvoDx818rJquAN
yEUP5jMbxG+Q5f6248IHyDNRDTRjlGGhkip38H5NabImNY49utIeILosE0sfTG2JGhwBhhGWXe24
McAptOQK91t+17BhEDw8VdiwbVOpJ6ua4E/dXrTqZ4Ro98PU+3qgacX7TV9fIGxAxWqSLfVgqLac
WLGDM3mG9JrfgnA9zmBNbcwwaSsMWTpraXz4hyNwAcahvUAutgVHhmLx7UYt7U4eA0C/m1+ljHxz
MATnd9qaI+uUHNzOXgPPuirRELZAwGmF5AoyoTFxGZFIT4wKTNu8nII8LRn7S/EJDn0GKtMz13hk
BCEWvwASnuJSWMzd/8nyAGGAxHBUbGvw6rHmD6TpKkS/YOpCbWJp6Uj0ccQSFNLQbD7bnVeQnpyA
LG2qq5SkBCgOSNaHgz0kj30BdKKUGAr/uU5MTCUO8wRqZkRAl6ID3yjLKEfyRN0trT6TIHKIDt/t
eKYfv8vXoRnlrxt51iQl+Dt6QrI8fHGPy8LZQBeuMBC7muB3zLgjApJiDPcbQwFFT04NFVOAwPIa
XdYemOE/W+NtAggkQDSiNEFF1q8w8hTy4j3Iilof2d0eaSrBA0/qCm4C/mZfdCAdyGEkyvVF5HOn
6tJq9VjaJZ3n2RjZccnH4fPgnLykJjOOsFKB/hL7eZYVbFgQwkoDTbjafCOIgInE5GJ50LzDSaCk
2EZ8lCr/4x9/c21AH8nvVQ1mZXeDKI/vHEGnMjnwzd0PQeUP+PUQJTHTz8XxNfgsNvuO1b6tDLAq
eI9+W+PGmeHKMIU22M7qoHN3BpPaMR/0dzRt2mDjnUfRIIaIeihIunLpMx3QTEucSggXCqEkZXBF
Ikeu9Jiphg/kNPGm8b0xUWYXX03Pv/UJYj8q4buV0bLtrRPlGzQjuAbTyk97IDnhCS61FScw5J35
F2yds6eJKyeYuim52rc2WT+lkpKgzrUKpUCLd7Xb4H6XWy+1ot93obwHOfrp7h26YwTtlFm8Xjqi
p9RjbkXWugHWWsBqHsdbvUejrFpwOlGgEmyjqUtBpA0tOO3x7UvRA0DpHxlmSPfOsNENswonAyXh
M32n9lnmC1g8V9rlB5LYmG1uiU3v+EKm7gTUFMoToqUYpTQVI2PTEZ5u4gGuhXxyJ/Sp1tQ7wWio
dGMNfJbGx21kQhuar22zUX2vCQClJw/WQewTYwHI5hlIfgyfE348E/ik/6KX8PQ+X3T+xA6alSxR
RoO45M4i03W7X679LQaDhS/RJj7O7bRJLsNm0dIV7VoAEfvTHvdPHHaYafB7LdEOFbUweflRYj5V
SCAjjdiq7/FOhnh9UaY95hg5NnRdnO58AS63w1++mixWuRZ4o9+sfM28H/hWFOrYCkZQZq95Sclu
mqbvSDU1SJjo4X0SA/QnXvh2pj9nYVAoiybQzeajqxPp5mFovFWxxY+2EhkdYSL/uPg23Ed1vOCZ
estSISBkYpto28cTzjBS/TmN6EjqoELxKCDaPmBh8QDeFjWjLq3h2JCbGcH2g7lor7dlSFX21aC/
RLA/zIy8oY1ov1TETi8cKuPVaz6ikx5kR8Wbq7TnxHBaLtvlitdkJKGl+udqcwG8wQwgHKVoCzOW
W9nnCEzsKP2mS5fMgqySA+eDyrhlZ7o2dc4lRYs5ayzz8BVad7bozAIdJtFmMYDhgPZq/RRvIF5G
0ffQmNw6xXU8vVKvTr7d6/4+wVv+Ii7XmgZNt8yTJh6/c+nBvng+pP4+YS3XWC84lJPldmAPE+xd
ovS/78EoGl46qJiztr17xLDouN5hFnJtHBv+4DDbOyhbXIe10Ai0GXE0L1hFsYm37+MlDBRipIQZ
NnB//kB+k0iFvH4S2IbuZAkx0mLAlFjDh2U2kGYg7P3ZVkKkwH0anKc2KM190Hmnh+m6uXhMUmfH
1uFrVaTe8HF7nGHRMtGvuwclOlg4TgpbFEk7fzH2wy2BYZwTzARiWWmVFOdVdlk46mcKKbvM9Idm
hL4NbBEWV8vVAsirxCT/gVUv+gKbWCbtFHOsa0ihRKpAYbMFxaWMDwoESIvoq0qae2/6+vu2fKl4
CIYXAzhh6NNxozYiHqzVbjK7B5w3IS9ay2u2CWZSq9dbE9R2+zRClhbwwlSAwBjomvRivfNAv/cu
WVlv6QIe1t4FXSkk/p3RhNGGzdW0+lkJPAvhoahmvNo9SN3Tb3Oux0pRHDw0kIj6bPkO/WjCl4/T
odPi+VysDFkiwWpHRyqkBCQgOqOtpaPRm4RkJv/V9mpOLoJxhOq3XPZ06XNiGDrv4ip8ODjQErKF
8A8l98t1yKhQM928a6F+vVT/Ghg/4CdUYLL0a+Vi8g4LGQCfGzZHYjoqnhAM1//53dDr6SN6HOJs
n9n5nQwGKveUZFcfBJfyqa7HrYFdbMOrL7Y3iuiCv00zR94R6cr4tKKuaOKKiIROZ1IeAtR7BXBh
WfKsdNf8nNiEaFGNZw+6f5mnrkD4YOCPoK/XppAaXAQsLixS1l8OXMnG8izNJUwLb4HOaFoj0pu4
H0OUt/+YsIfVbk88aH3+6DlB/UOiTfUJteDGIc2Ir9J+3P71HODvyA3AJHHzFKhkVPAaJ23v2S+X
r/blLE54XzFGydetfg4QcxkGYEtv2xAdpVsjakwpnk1YI/oJzsG/XC5SoAONYY2MldjmBkGA8PjS
yYfd6FfVLMFadXVSHamuvhK2NEbgEZaSt1IktgRLtV0IPH0BVVyc3N4eEZxhtgPv8ENjBigkdAx7
FB5zRuT31dv0pOlqaV1fJVpQWz90RPYaq3SCI+vV6c/6Xhyag3l1IXImGlpiEODgkRElH5AqlVHI
gWsx3XaHxuXVzSWp28TN76yqBUXPoK9JBdOhMF6htkStiWSl2oYIesG8ptXIFh4XLuE1K//SrDCX
fMZxGlXd79U315oDSyMH3lqUQa4Mjd9QI7xQ34XvgDnfxAmG9V6MMJRn4oODb3tBVFwu/GlP+kfa
2F3ZagCf6BjO9l4Q7cNteS4/rRfcQUmjCdpWV6TvHs8WKURTKN68umosVGrfEF5dyCISMzX2QmU1
U1XrsrDZgXuVbFrbhXUETIA0fR2mPv3icSWUx2RhUTgnc2PbeRYegkOgPGtc7RTQ7yT+44up9yle
I477f3lgSHTCr6ncjjLI/h+cSsfGEIRvEYiY7uOYWjXgyJVcRmLSRrD2AqbJGlyOLqAsZGZ8e6Ty
LC5GxS0cb9H3rSkZP9gWl0APQe+fLkocU2ABRghbndnQ8oJtaVoCZmelbsHAAk/qS2/EmCIxA7lr
zPvXv+3ZYmfQGHMgG+roVlrkANfBUVupK8s5JBKWX3aKAtEbVnH2EhjgbJE4tleTQKdlhRufiFTh
JKxzM3UB4I74IZp1/QL64oaW/GZSgunfaHnDU4HNn1fprFtjSmSnt9jK9KYvQm832uI/dUXFVjCE
En1IAD/bNnDtlcltkhTauwmfGntChzlrMzf16Nm1/Gqy5DtLl1t80XNPg2p6vcxBZxzjKHjDad7b
er8HiwIM7VS6nhPtJq+p+SbiE6aB8D0Gmz0g5ZBlv0j9HoE8EJBiPpP5RFKrWVMpS4nHE0ERXnG0
amuu4t4vNJPwe3kTQ5Z0Of57nfM9DvEpcYDev/hiUpvkLjzlKxHjJbV/pvufv4Rt0in56OApYpOO
rIIbCISTvY1YPGifomA6VYSJFwVEeQctZ5qOeWAZsFjvNPj7WbHkb+agp6o5BpjO9eT78w8IrdTv
8tiJ9+1FdfMJounuQtZ8+ZYPj/yNpoHY7+CKI4aeSQ9e1Ctb/Viz4XFbnFiPfideZYoAyyCKBLAn
iVXJxQjXC84choPHY/BVo0n8ce3wHUIBMx6oEkE1PMYm8MjRgLeONLOeT3tMatvIDwNPrU4D4xuf
fUot4dGP7ZVaJlO4KJvi2nmRvLdkCSW25ImobNzrIVa1Dw3v8FWq1Shz0SW5XfiFKXVP81eYx8VZ
7eb3QJsBkBbGWgYhUsWdHP+JdMZhtCI+22NWE0+q0LOCLw6tDA23DZ6WLTjR55DkFWUg5JW6wmr6
3iFT0w1mtw1tPKE20I1szUiXNRgVkNMK4Eo14/5d2/bQYaEXi6b07vdQJ/qgKuo7knoAnDLk4tvr
fO/ZWii4g3yQ1i4MVYzIrweLC9oQ2692YxKXLI43t58flT2UEa+ZIUQWKHBvTJ5JS+p5mTT4okAP
tDvJSVKzd7P4nQ5U+gCiH0Se4JOegINDTdUPUipraWnMznMOMai3euZX2e93ZCJ2+iPpaCChIDLr
30IVgsxO7ELmh08Z9eutwvkpAFOeR77ZTWBIahoiU8YuQgKknb+7/9IYtjVfm3/urHfk0yCrqRl2
2VEGuGIch2lzxb6fRpgCFYsm5rOtov9L/16/fT+a2upOVUDNSFMFAJSCVD/5fsb8NKDEolotO9Cj
+b3qCsnPPQtA98oYUVVuX0sIgYq5JejgVYq7E5UCflXLTMgXsj5LtPTLwQEyHofJ/JnQuJyrGOyM
5P9FSmADuG0IzRTm8598a9yZaEHHJL2ci2tT3avxltAD4WCQ914rDhF+E0OoKPRksvilFyFE4dUL
2LRL4wYPbt+c6KVOdJJlo/z68nHr4YGWTrkc1MZgzKU53BX1lmSdLBaFrLlfE4LdQafPB49PUZTg
FT+hiHWEa33WgYcR/2FolD1VCmnmXlrORKkLNlsf437F8XwAGXZlK3o7JWc5qQ65k9h+n2xmsTtQ
+BnJFeVQgwyGi34s4Pvr/ABBdc8pgDD0qIARdbLt1l1o4w0KPp2K//C3+U4waAVkaEw7+ccg06TK
Xr4nZfVsrXeHmg+Ez5xuIvlquM6jibODm4qFdCKgv0bakWWwZPDtsG3SYXtYHTI6ta4p0aoLNx3r
p6yry/HtA5prZQH016+m5GSGyGRz1AGe9zD69aYiDOVMbDE89/jJbdHefIpvsDEVQqXEgWPqZp0D
mknVGw8839pf0LaWI1SIhcHQL9eHtapjN9ApDAl+MoSF5awpyVqhPqIn6f809X4vTlg+DyNLfcOW
zS4uSwovCnxVo65g6EyRh8et/VFLCNyjMrscVzplAmHZl5iTK2jGwweb7BdBWikXWdb1R3y4Z4j3
7E/4/YUaHcy4CGK+2sYvkNDOoyx8LFws8NyvyPudFI84VXurn7Pbj0jeccm1TYIdjWwku4NxTRWP
Ev2uQpqrT1cGt4XDV6d+i6q9RAJ49mPBl9sbyTA1PjtLigY6L9bw+v/63bH0cYMKJMZXRiTt6cr0
rJTDNIGeQT+JIj4ov6xAqrWuOAo2xUhWJoKxS83EWrVwqRBbWSpTAw/zbIGeIuzsbjLMPQGk3fHr
Lqm3Nhfasg7ABGxrVMMfim35GZBGh+RBhfnEW2N5CzmUX6K1AIBpF7sXDGN6Mp6Pa0+LgoxvNNhV
n5N6GYChXsGZuuA3SoJUL4TBZZ5M9uQu4oLguXTBG0Spy4LIQ8ctoqN917B4/gjGXVRO9UCB0ru/
JZspkX8I/vR28wTKIQafszcqenMvR1OJmKxn+E5Io3oegSCfUvO+L5EHqUaOGLUty2w2UsyGJpMO
sIyQtCpQGUTdE7pXCsP8DyZ7Xgvavw3y68VqV23zLH9fLrJK4xXec2eG6TDPLWq/rciZT0vPO4zD
P7gX/+4eWTfLekx3+cAQEh315geJp/AT/M4P+vPmoiLVJ6eJqXvqX37ujLewoWYqjdEcZzaIKgoJ
7mGXsf6aEziAL6bx6YKzQilPP0RFnzvKf8T9IYCNu48rbf80ujoMretOWX7Y22hJ6vvcp2BEATTp
47Luwle1+BzkTk7Gx+9i5ykpVybaqKudRw1Rd31BwY+uxs0d1q0vtz0a6qs4yMSNlUEPaXO2ykHh
448wpgCbBcSRwjiLbpfZ4VwGQVBQ7cUBKIa1rhzXSBdVNKY7SD4BOSH2kYiMidFoLt/AUk/U/m9y
Otc4J+rVbey9nj1ANm2PPVDZ+7prJxGsLn9q29m2j1a9cTwS9hYLcN2foraqeCJnfY3z6OyyeFt0
JbRy2+g7/UPD3FGOBs9yuUg6lxJsRQGVRnkrmgNlkkArU+ZRm2dkiMkXbelrPfILXfBiJnmNhdV0
wbxhb82du4+hAqPw4RMLfcdjwDonMMVSHhUHG8YLY89YHQYbDcCXG5WIxOqGbIxbKo3RMq8V6MWf
sJM+vEjURmTzkmLJlS80opuRgRgb0nVFCQyJSeWc/nhYRZIa1rsNrScuOraZBMP0ye2TcUjx+VS7
u4sngMhloDlkVA+CodN0T9gjZtnvbnuPTrbSgZPpe5jfMVjH9d6few9TIpDAA7xy1qLKatq33ZvB
bj78KgvsSJdaLUcOse2j0W0Ft3rJbpirjhNbaTGNSOpO+wKfygPg2lZ+FA15v1BhQDn4/cLMsH3u
1CcCXcDjKLjN7SGQRQX2GPkLHU04fLejbuvAJ49fYcBfdADRUW8Zz+oC5RDnAexnaesPLlqAb2+P
T0heCjHlx1ZTUWdaA2i9CxgUgSk+FrRzmK7kKo0R5P92IlFXILhJ5Fn1V7usOSq+fF99eAoOvCHd
mGbP0mlXkw6XiVIVOzAxTrk0uJxhJdxESkVeHclRimfFzysYvNw+zyHoqIhXJGUB8xG3OK7YQoUf
C+ynxw4cpeprNN46sCMpY/KjIACTasWeefGQgRD3t5UUtq9DclaCU2bLYYvO1cNx0Pd5wyL3z5T5
yFQTGrlhE1/5ouTdlVvhINgujfnw3mHiabIVEMvO4EHzS8pgqEkILxPIJjSCktt9O+yZaum7egtn
an6ZdsrY21i68ARBiGWvKz2RK7q/Asmf39IvuzonWen58bnWbi6uRL9fAoPw7Bt9fMW0i+lvkCBB
+UcJXnHen8vhHkzZ7kqB7qk1CCD6p0araf8B2RZb8vMH0vXcuqo2zHf+5rapucZBrMRlBembR074
AO4zBtdrZA41IsbqE5e4fWfgcgsFfqVAncaQTXQUpjPYqvR+GVK1if2PPH2VphcWQJXpyK5KChen
JrSKOsmQ04fAcdsN6CIUTCE1eaDGXUFHHpvLqW7W6fXwYkhhYsHLU4xkkM5BDQFmRTT9MN7ocMmc
jss3aF6dSEtxIyNmuv2inz7box17MroRFLOFxiC12HavStwI5yfEtzPlg+R2Lf+lyYuic+mldVb9
ifJqd5N/yb4BQcirgM96gU+fhqdHeGhlqjlsXIlvSSo0JlJUXGgjR5hlMQmVlN2sdJmGSOjRU4T4
sRR6CbLXrCrXvMfkiNxIzI+y+8sxmFZEXcWp9v6KSQyjj6kDQP/1vwlaDHHgfaeScD6RlG64NfMY
+XXp2FxjvJ5TPta6FyF2OKNl91ecNNLztQ+bC/z7R/UDjhln2Panyf4N0NQzUnKlQL6NClaPugjW
0XAPKGlxC/LXJa+tk28tSA4VZzcGbj9QITnOIaQ8m3///ThmsZs7t69TM/0CTImOnIL3Ss7pgMtO
QAWX5WeGWXsvCzkXIDNtf4x+SZxRO/4owiCrHN/3h1DvKTT35FVt8u8btpgike6rixHGscee5d/j
avNHNnbe/xRhJoA8TGRygMFOQFprCV7Q3x3C3Ku7pLkU9Ej4377Q0EM8L7uS5MIrXPOUoZl/T054
u+IfD844r/zC81spfQaeJ8S7zNgPMdRD1aKggiirz4axgoUXxzpqAdA129k9InFeBI+McmRzfkRy
WPPQOtAXuDejrDO3vxx01RpFZqkMln9Pug8XSzLQd1ReUb05F4awKMhcLNBe03QhdCjk2V2CO+Rc
h2sHvWy6RNIxelUXEduAB6lvPXHmJJfzHMbb2KB7LtB97Y5/gbU7iGC4J+axUHKSHVpISX5PvCOr
nNiRGOMXBXZh2+/I5BV27fVZWUbAlPo4rF7xgSv0bgZf9QMozJyso3OIvjzIIb4eNWmZkyBaT+Ar
sw4pXWIDSvrnAny1nT341d75K7sH6pQLxZDcRJq8o3fYCc7j6AEJrTgNutNH2F9K/0oXx13ipkpc
7jM5GLX8isjVvtYmFd8ZkyGnMaFxguMFtZpDD3RnjAQNOgsYWnTxt9UTL8OqI3S51E3y2SsV/emm
54HVBQ4jZ049LhdKXIXWWd6Se6Aw7Xtu/UONPxkDYGif/PwgOtmeQamPD889xW7pjZ1bfiHumEHa
miEdt5abnqh0kkal45ukzys8DVn0E5QVZi2Z72fdqtntPv7KNQsIO2nUC/MkfeVPwTcqY7JlcHAl
9tpaU8bc3iR7dB4Nf62r4jrL2YlZJIrXtfElIRrN46J9yUS7VeNUZbLoNiGbqyvc1mkHC0bhe0uC
GQCZ6UJm+2zY3mzcK+Z2Bt783r7Zf4oquWEtibGQIzU3XHM7USjsMhsAEbdJoCWpmLg1ZMddHAA8
Ka2FlGuD7OdPFaf87cxVgnfZIt6I16BM79afHOrNMbeUbS2Y+t7VJ9XZA98mZRz3pyTbO69GIkzl
mi0zzMg1TlEJsJAhvj1CVc0dXuc8RfkmCe0VEj7AJ1xIuqUG2v33MxuEUqAkcWSLM9RCXzOCMl5g
YVfJwqAnPEfJKbBt4nhT0rsWj8aQJVMOORPwstOnGWhLid1Pd0DevwtLpMURHuv2TzQN/9P8qfHR
TcdAWOE6AskQ4eIdXbTUMOQaX67sB3hTraRApsMI3sWWKGZk1Bz/OqgFYOBQjEZiSQBDLwV4epOG
qtuhiTAkBWWNeoNF13zKfaXK3yWiJEjCCOPs9EkNQMUaY9Th26mFthi3zzdwAylcRqvTZZKqn1C/
kdx4TGMA3kYhGVVXjszC/WxvizuMFW0qD8Klq6m0GNND6frUrJw8yNqM3pujnI9J2YTRGuJbj1C0
bhHLP7DilXynbez/X5D7oJyUXd1qxN7uCDFqn6Lnc7ioiPYAvnn5MprLdKQGjVwQxrejI6Kp2GV2
MNoOrxXMaiZlQvofvXt61TWo+qUrVbk7rILWMLXZW0s/BaQyYln7gSkib+h8eEF2lnLNV3jMdry5
kDIH2xrPEdP3uWMQctECXuZ8uHJoKQ4S+i5VWWnND+567GeQnAUMp+5Mw0awuLSGG8J+Hm2ly+WM
J19UQz5ubougAHYYqiz3y+S6K7kQKivkKLq+dNvtZx/tdaM3WyyE+qnOpxOuxNZfusa4BOKdcExx
UPxK7AD2kuHPKS37d+elXryVyNTX4kNIzw1v9Fw6QxPt3vgKdFIs9jhzFmfnM/vwXMFj+CBr8GWc
UxGHNp2gW5a3IAwOZB2kKkQ5GTnLotrBb6lb5IDz2r6bgrCVeEXhvF+fEPdpukqMFqk1/oH4lxgU
oK626fwAmPD3SBIIh2U77tKglmXFxDb9cnqoTwRQM0rMlpiN/gIPxe6W9HehAXYTahle77De78jR
1BfdkNdDRt1YdS5c9q1tdYL4HQxDvacBlxkTKereukbM4STxCh0+393p/NfjkgmD5xSRE55nmjnz
c1DVoa2wVOJLXGftkL4AAByQIS744pS3aoOqbPuLdLKwommEo/m0wCdHpydkLXsc/0JEJYA9u/XG
kq9fxA6B+N/gCHXDPTE7Wogyzs9e+w6cmsTCKjzIZOumizILKqDl2oUta17fLu+5av2eCJSs21EV
gyvI4+AHktnG8aW/ozQwf5pqZYaXsq6tc8jXky00FHcpuSg1BbCpA0KIEs5dSZgo2nmJwdh85QGg
ljmCT3mMymfGy30ydT2Wj4GLp4ucG6+Tp+w9vmcXDFgHCQWpAVVGDV1fwyPyMyRMS4AKNEvNNc/9
d4Nd/zcXrjCb1C8D/PsjCQbj1ypwPrws0Y7xDVp1ONlPlcEb6xZHKTjIODLvEVnRmJyG86jSvEpM
HyRErG3oaZXJlgX7zzwe4IkR8YSM2x8fUrzcPiFLIhUSYoMYcIjoI0vsad7nGLJr9+Sx2V2y61ai
Ufy3ZZn4/K5YdQLUl/noNgkHjCOEx8qp/RSbOZsqv46An6Af5EbbfhEdUy5QPVg8M2m4uIFI5uMa
/1NeNdbnB8Ih3srzjivlX8PkWPBV+niHXL0CD97+OynbfPRErA8+xD3usPmg2PBkYbY0U/zBujr4
YtGo11jG59P5zOV6dRw086anV5v0OlrN30yGUr/1kRbLtoxdo6ghVJsJMQUhhMuaMczRuClwseVP
Fh2DD3UgLTHsC35eV7WEm3vdPi0/6qICahHc3hQ/0OfxfAi9Pf8GUi7DQ6Kq9NRcKACqi06KbYMC
kd2QZbD72ttwuXnFcTVy4tFo+XTMQjaDjF7e54AOh1P76x4vJSXjs7Kqcv/fQPGv2D66W0j13xBL
NCLgSID7Gu1sLkR68DC7cu/Y6PSe2YTe08N1P6bTURSDmYuOW8uBlu61erX1FLjErk9LkO3NzLC7
E/eTD4VgF6P8lCkvl2xhdcTXFLbtrTzkTSvIaaBF4MhFKCK6lJ8LCAR2oc3MELf8ihwbhtcXmf58
s4DftemzlditPPtpXRJhrO2v1S6B0aZ/RFePgvAVWZaKIPc3mkZkYwsqUxs5Fn6rdHzHuZqeTMix
VQC8U0DpMToRotDEZhsVTNfvtLo0V2YrqP/ZYI+x/IkYGU0uIU4jZz90lDi8qgdeAqwEIyzS8arP
5mO2ejAs0s8ZNbZCJUrq1siwEVL+CfF80fdvPUivCU5iepRMPuNDXqGVi/r+Li7irYsQFb83SXCC
rGDNP+PdgVrVa4eLSY9XqY2zGk8aHb60TWVxq4nbBAvsth0Dx+m8YsP/ZSvkZFYvNVyatcGdg6by
DTEq0+tmJMtQO7k5bHMnnc6LrhJ1ogOeFuta3Aw5JBOHZofBnRfmexLQ9ShvaMLT02RiqTAuuHNQ
LlFvtPSzcmH58wViv3a+p0SwHqIIq2a5i8OmvRrYD1MX4dOHqfBccujEnZzzC/raJFxT4+KMpPBX
qxURHvB/8e0ErJhabQrDKFirRvhD5w3JIdmvLuO10BiP7R5dU4AhWmqF5NMOdZFe48esDJEmi0rg
vNQdxZSmyYIh7wKrLDc6RQN6zLwoqWQRgKnymVj7fCTwr8neE94GKFMFmSDbGIOetX0/2bfbte39
rHa58J6SmfNTRbJmiUPErewzI0NKLyPLzMCNuwXNrfuwo3n9ZKI/Vhdb9H4QLHyXME53Ihb1YAjj
160kJuOyYTQG3a0mYW/EYj0vgFvigVCOWoabPBfMMyjkhO2s8+S1M1V4ZhjFQ32wsNk3FeX1WGf/
iU8oCgIHelC0cAEFANlCX+baDoYCfFa8UylUvF1UPfbyRwsgoHAFA0lgPKGK5iJ9ny7HonNX6tUR
cybGAR4sUFLOX33LDbFAq+6PDiKbzxmrjwjop9mJ+7LZOjUuoTRQOm3rElwyxmh1gCtMHifG71Q5
miKuD9+VbMuP8XOahaQO7LNnpBIfGre3976Td8I8Qn8VpBOO8dVL835XgEy4JGEwc5sPMy0ult3S
+X3AFIHDBrrgEmZ5pDSAYrysjWBKs3aMY6xc4htvJRc0QrUnxnSRu3bXWrnaWjonocD8cYNM5ik+
m68/APz6z5dyX1fezjKEpLGvnPGs6lU2Er3L0gQpJlg9WZ2bgsOcCFIEECzubiQ0QrPiSSpOfatz
55RHyJmY+gXb+GQx3xB/MeC7+ON7qdDtpI5fzJ8N8D+cdN//c+sBp8OXAVJZSHHK8wAEhiFTrrYA
vZMiHubTOSwPACQizvgCXYYp0hwQxnYg0ePLcFPcl/OjercEceZHPDZgpYgot7B21IgSmu6kPwdU
/BNY5FNEzdCAV4tDy7AWT1mYIOkc4yrp2uSx3UAp7FZuN9B9utaBbq8SX/OCxDHVPG017qdUHHsM
vtsVS/AJREgISbhIECazKY7r0W5fX5WpIiwFurFnw79ebj39LEJ1hfEXWjfU55kZZaXBNxmGClyi
R0V3OgDAiFVVbcJ0VjlFpHz3OsmOaQSZLyHQmRyjM69J8jKD89CCshWcMtohSh21bvvHBh770cud
tAPIOTevhiLqE895g7QsVABCEBYuy6UtupHGfDbV67px1pOusk2zjuVOvlj5YvSDB4Ns0jsMe5Ci
TKWlZCpvU4BbEPo8plMEDJ1J0TRqZk4uErOlqiqdN9C5jFyElRsQVSDQuDYgmqC90kThjkXRuhFg
Xl9J5pftI/soc+v+7ovEgp7eZs0I17limJUJnd1SDd5ee7pUAneebjI1RfpyGXkNCEF8RGevjci6
tUqBpr0zpcot8twtN/W5HO7Kfhxdbn0ootXH4LjBGkwJhRybdaINLjcc0XDV77E7PtU7Qdo3PlQV
FHjV5RSC/HUZ74ktj3Mf0yxUmppZ1DLeQeN3vfc796rWQr7auCcE5wkHBUXYPRx1GEazwvn9Lmpu
8Gg/dxfaBQJIchL6tHD1NIp3l1l+rQkCGipPV2goUyHZ9zI9G8c9Sq+E6lVfRtqlueMSQnyM++y+
4U8x1L8rFaqnoxlM/Cjbh7VzAeZBvMwocNaPIYh+zt3kbuWCA/W/F1DvOB+K4OvWNXKEFubUCfvl
Q34mbTbs1t2rUoBOYJ10yGhOZ6VQjI28CM6L0CowbNdg9oWMbLHVTxAE7SOjtJ4HNP3AYDWrESjg
bYjwZzyvlTXOMBmPAGq1Qt+rAGmSwyTDGoLXPPpO3bdJypdJQGITrX7/JAUvjhZaCYriNT74t315
IqyIkadtIqu5AIA32FfNwAkFx9s5uQdghpTM8SGG2OeL+VEhuMKITzv7PmfkMOA4CzA1Tktkd5yB
xQyqipzEg74TtbaiiaAnXro8di2EgCY4eHVueo3P+m32Q2RsQnRSO54AG1ALlxPpe7H/LQhd22r+
v3B28TkKiIkxvufGksMX52J2DRgngayAVVAfVhztV/XFYGLon3/m48uGeuI3+vkLC0iB58AhYoa5
E7Z4FANG/k/jSBHp2DwIAWJLpppTlKPXXh6G75FBAcgiyVpL2Sd92YWNt/O8kF7nE+DOmqXoikr8
uQZGKKognhkF9FOuyyVGpdXrtRtm96gQcfwKSrL/mzj2GD+BGSBfI1uc6tcBR0bdwhPRXnosC/zl
oOWuo5aYFgJw1iM+XpV7joOk0xLJpRW1Ve2bMsEgCcF+fK2CFT1kE5rI8aG2q6f4NPf6gj7N2xlF
MA2B/oJ4Fam08EFaesIPPOlY1CL95QqcMQpIs7CGaDsWCeVYu/+HWKdh/3fncFdUHzlVAjlDMEh4
HS/5F4rBBXO7lMFbsXwVFp8mY5PXFb2u1aNeQLeBHNQp8YTQXEQ5FlUH0Mb0DlK2iBKAAItuZjja
94+p0uJWYdiTCSl6rfp4kjl759/Xb1INnfueg7HzDpzI5IRbedYiEgy1ESYngGzZHiegfIux5lHL
NO1yrPfYlyLAiiBGXhSKfSrbmM13w52ag5JpdF4HnPlQuabpXqFDCBrTevhkJg9WlEFsFtqGGst/
olAO3OUtXUKmm+T3Ll8dW//0KdWAx0BGKU4A43y+JwzJpALE3BAMbtUENyiJUbbvu7C6wnG8HV8+
CwXW/RXo83fnpZhRU0n5QBqahedo0VoM1LbXB0fkj27e+TU0WaIBHNOW+V+LtaouJroSj95PxJym
Kdcv2uEAN8pfDlsJnA1FuXkpLs5WZh7XOk9GluVSVfKgDI5xxTfTpNLPkKU6UR/DKfHmpDSxb0Cr
+kqK/qNW+Q9SdgkhvHcG1EGd3MJl9qmfdFkSD9eWGJUM4tsj6Z0kK/ClyI3R6xNv2FKrcBXgGQzU
Kr0C4SwPuY1h2MfCNtcmlAfAxPbNA4Q7dWtqzQiz79kK4XbEhdfiIFE7dT7kgFAUwXUTDaieoasf
Law37PIMRYPkwoZTMmrh2w0soVqomhIZ5ZaklP3eSp7dB9yDDOYjRh1h+NmT7Lay76dLmVMIuTTF
kCA+SLXeLQcawYcuF8TfVCXfbh/1S+t5PIlVI9/kN2xsetNLs871A5d7TcoaN0UqTfWfEa3Opt7Y
hnKDIHqKb3335EoVZCedFHqUi6DmCAJ3OtwnqB0/0vDXV6HJm/JmhAgbyJZq87Od38bTGdKiWbWF
RnqoSPx1aajLOoyIDe+vDHaaEahx/i/tMxdfK4XA7VtEYeohZh2Cy9zmRowpw5Qy8W5Sz/rkw8Xk
6bp1eTyy7B77zPpt1dbW9VvaWKCRsmWY4Q2gq0Xqr1bfbjVcWdhIwDc1XHF44KnPqxmH14j+9BTS
tmTPLjcwb3v42jogjbZhKLvyvxAEc65hkXOfUK1DpHCKmhw/x9eW2W+ayTiY2HUFZAn/b+mumliP
H4SoUo6fMQlOhXLjTXtpyCL1t4AiSfd3HIavtjWp/JvAaD6zISWwReRTY7J8+A+ADHmUlyQypqUo
6A1QqlTQrZC635rVhexZxGSrJyhETMn1DRVTPMp7oxerj2JfhiFQM0NiE0L3hdYfEe5XtI0MuHFb
Fe+iOreHfmIRfMZVc+8rpKQxh7ol5VAaIcnp0EdnzO+VXWSx0v/EZMrVDdxjEyUGvU+Ikf6h9lYT
8j6Sg7J7NvK5bW6lXZkMV0LhUgPE3vcQWcSCuBNBx5V1EoaSgXZoWF5pz1P+ANX78cOstjLzhsdo
wgE0gmQVaRk+ndKUr1ic8usPf9IScUir3jbph24xpz+L40+k3NjAzEPe18da38lvJKM66RHVKbPi
BMO9CLBoDbqTA3Q3o4l1sGG4pnuksJKqGeCo4D3tRejdGg752CIi3UtUufwoIMsf3Dd14MjMLiZ0
sS6jRfCGcSyJj02IE7L63LZ5xpLmPVpklAc5vqLHR9YpNNmj0fnZse1ZvQr2pGShjQIKF+km1eIx
e1aotQGzjkk8Hfldh4v5CKBnMG0rKMIbdeetjGEMJntg1ggDZE8rlOF57BvIod25cLuzGSNWJG89
mK3KY3EVd/LmKd8tGc193GyC2ZanPNINs94CqclZL3UKQYg1xcuk1ddjYyA5vlfoABkERRgoV2Eb
ZYwunnULDCc7exOmHvVGtvN/USVaR/rhYuEilj15Esuzn1n7D7ZHcReHcPKWN/kJw7CgoleOKaPg
41dyz9Aj+u7IRzHU64/qDLObBd0sHVhGjxNgeCJGVF5cnRNxW4MGPHz65yJwf4fzdLkiPhQ05KS7
+F8nvJccNVpZfo4NgIMVwZDPBBX8EHUVSJNMl6pABVlwoEZPMVLSGE0WdjfRQXm6YtPgp6A+Q0q8
+lpXJyUAUQ67PsTw5nstsOa34lOY4+YpvtwWpLBlyFS1KWNXf2CDIo7lBB2MGkrsxivRRip5Pfrs
h1aSNnsU1BsNlPZSQQJNLrxofCVJ9mKvJp1Ukne6U2WykQRLL5AkvHc0FD7BLg4NsaqIcjV8EiqS
cyUVjmWQXSJvaZg1EE/0M6N/rpMIc7yoiKzXAzXnNMlyn/pui8HppQDYGHcSwROjHL/72TNdUAEf
4ptACnAQ3DxKFP2rmU+dCJ0e24KyE9bA5XqWPlLp9xQsxAYQTHhPIEG3TjfwOFNwi0Kt8tKoagsb
O44J//J+YrODnpwhfbEPTHviusO7QnHric+DXDAvzizaIn1dKgWZzYrHUAY/XcbL/858kaAiiAKp
txU9oZUBDokICLzflB5BuOGgMX9H0nViUS386+tND3+FOSpURmNl5UeO+KDBaj75/1sBTSIs/pVW
OY3bddjkQFzwqNdfiMypeQCuppVwpJvduZmZq9HaKCkS2YTIbWDaq9F2WBJQBH4sgJKzYxg4UvW3
XDhM7HT+rUUn2taLI9O2Rfg5aAOT2kxMeEQD5gSv6UPq0TPtkGdwEIAErfpqJ4ZnwhiyJxSyI6ZA
BYFmyauIG7wn18q4Nu15dwcLNArnB3lrKJfE92SSiC6fI4u6FLiDlS4g/N5w0Na1CU4/2hGFBgjw
KoIDH5zKkKK3E4GDnByGSE9q1wHAPmgD6m1X/qSon/LKG4m84vBw/asgI4tDQVSIsFmcDZu4JRik
mVlSsoFD6dUD2DirhaqktXdmYD3Z4gkBhVP4aUyZZu4Ch9PbsTqI7F35cCRxvbqOGmgvKfuO/X9j
zjWNDeuOt7/EOPi1gaocWerdpN+sT/4yV010oYkeJSa5xOv6/H/IO4K0ao8fxMJ2lrUkCjaVho2n
Xs1kF8ZVX45QfKe1cCs9WSS6u3UL2ZtdVgjX1cmuVLfhEm76RNq8lD6ope+Fj+7U8tK0y23RC0Vb
RCWX7WTaE3UBNdE5SorH68R2so53Ob/zolSPbIWm8L0ck2/2Rt0iTVQItU/c02e7TOQq0crX0+sn
1iLokCswBpc7yZnUWAy0ga2AUj6YzCOKNXZqhWoeQaVWtaNxicPKPU64ZN8MuWhjDLrgneut2MdN
sm5ZAtjR3wTb0Sil0I7lGJ1OrfjUeyPOVJTL3vU4/jBOhA5AUnD3wqqbcGh3xG5srzZ7rV+rsCP5
3HSUo5uDM3Fy+jZfPo4i+e2EJyV+u1lTQ6sKAcqFwn05+MknJ6ERu2WBaBNR8d9GwJU3+MVGLaqM
cwuvoW7jDSwYVJbOE78eT3Sf+oZtcrbyYINJACtnoOXZjcfkZy4r/KOZlYigtqPtk9V9I/D8tHVy
maKFV1w0sXTtaQ92ne290tc1Emhr3c9cgDqcEUXF4CluYKSLdjhuCRHfpcUvWqJUTlbJLCtNqEaR
OJcZMwAVEofkLoPMP0NGcXWC+dN6u3WkJ5V4Bqhup59Ra6mN8sf7E6d2JNvHkiVew6r0xguk+f2i
PhnCI/rfc3W2Jsx9vCfaJlArRXP1dx/b53ESljU2PbtIPFxqwyWdHOEBmNbMiWRBiJGZwQOTVKAp
IgWgd02qCFvAU0ZuAYt0jXCC52HRM7vW6NeSCVggURmLUNbWa02xioNzbbxDtv9kaPeQPud22kFs
MrvD/b8XNwipQB5lky/bQqkX7UnRR7JxyeUsTNCxNqBT+rYawAX36gADadVG7ObGpChDn4dwnGZG
3lTxQ/vykkOKgI6gUWHS6ZgpnwP0iv6I4As5L/sNSX4HRyY5bDm1/6/CASCNnSQVYyFlS4dnhg73
fJgriydSF7ExMfmt8/zU7lD3b5yQDbIjCie/Qb9S3zyF/lziU+k0mvI8W6h4RL90Xm+yKS0/MxvK
yUiZ8jEh/bKbzXpU+9SYL8Gw9o2/CVVWtbG9YeCsmRqnbDuOptoHOF2F+dctJiA+i7XJN1NxIFj+
bTPCpImPyNiLshMZP3BxBROuXhEFrJOgWYB1GX+0X9JDkUhbMvwQFivfPirLeblmoZZT8rcsDcvg
P6hiPZY3RjGWE/tDUMg9BM5gAz4RX2eA4G33SuMXKqOkiVekLLjdwqK5mpy6Zau0jKYqS/4pq6Nq
i8o150hv3s6S2wtCUWgJmpoCZnBKsMBxQOZUOv2ij98W8BuYJT+yCyJv+boc4/npxwdZSf1O9La0
wj7tWDbKvjfksvMFuM+tv1xUgcWPq3rSFtzxIjwrfHH2bWRQ6Cf7+YwU7aheE9++bcAtb2ZqZ5BN
MEPauFQGA2nmndr9RG2qFLjQ9zm7kegrJ7+k2suzAL95UEm31z5sZmaLAoOVd+LpLLf8BPTQbw2O
NPB0ezRxtT6tvKtEupv3KCeyI/mTWjqtt57QAOUdEakxvmHxiwngHmuMiENmAT3ALzW4YprEw57z
83u0dWOI4nbck4L3rzcLDMFZTRLCfIQOUm7ICmhqO4iBCUPhxbfT5ERT/Q88sVdtQgVbFweJG4L7
vbsIhXAVXRXIa2srP1MgXJrXNYs9lvS426HZjJzuBCH1Ja39KNR+X5L/gA0WJfzJ/snumCvVukd+
+/KuSFxOGm0AysKyaKi1XJ75JixPYs9Is4n83mQiMHEmJ3D44m0kwW1rHWRfH7ka89awQJHWBSUO
XmMWzqr/D3udEvMw7rB44e2EY3AJwIwLK/kjaHwA8wLZ1ooQ25AwEPsLQyeMagdxmVtGPmddMdO2
+BJgO7egvCyTdf7HiT0RUTUzYlEkWhzTyoCFfq+5AyLToKxvpz6MXRlRQeYuwyiSMVep3DZ6wU2V
iCOpQnSLFMFRG5c4c3ukctKfVlvVPizl2PG+yiGI801ULp3P/9fJNLhF5EKg/u5yevExWwpbpSDm
iZ//LRPKjCmwXvkf/5NrbAqssHa2e8v+41OnerANKIVLKrLp7U1XwavEzn6b/4ZVSZ2HRy2d1X9y
KK1qZfavcjB2bnTNJ3K8rL7tNwe18dHJXZMRCKcXZOPuksaV9KBHb4/y2WGDwdg3vbQjXd2VleN0
k43eOG+qRtLXmAHCcVr3BEPOLYz5T5/9rNTqoE3CH2MJ8io+cgXwVXsWXYyBTItkYKpTwh67AmDI
N0Ck8K/6AbC44dVNjlHHijOKniKmmD3Mo1cTzXgzstiHX+jGXqAe+zB24HXzI6ZY9Is8MMdL2PLN
AHB6f+TijKeyMOheYlXMS+J7Jej5i/kMpQbpD7HFYdGNxdiV4/ibY+0aaBOOqiS3YyXkhZPE5Gn7
uYag76L06XDIN1KBPPjJCm0Ctl9NsjBR+EEVhs93FbLVXk2d8Yw43/+8lK59B0k/BnaszRfA2pKn
GqC1ufNg7BZ4zZH2ZUtzOe9q1xc4zSyTxH3E76cL4rCL8Bfx0buTChAmLl2+c8vA+zJyNlNEbC82
JNwiYlhjqZvBijKXCtrYliM9/n0zm7jUz9K2uHpujq2gFOY3jmcButaTzol3gvFpE6qZ6RVfHMg0
XhDZzTSChPWMQhM909MQoZvhNYlM1SuYmRnKxn3Rzv+ruh/6YOOCdrgITdQDp6dTuq5oOSBa7qFB
ilXCjmRrBMDlgGZksr47BjJVunwkCSILJXJIEBvGby8vJXlVmbRovBdxNFmHvRs+zuGlYdkd4KgL
crj9PgHGvvZdaxrZL+V2NlbQ7vR11lxz9M6g5i5pdZXO4LZ6cWcigQ/Oihy4WwhTM3U1IB+xtun8
6UDvlSKxggukPdwEFpHehXtpxq9peqSIcKXQN9WUak/sgrx+a+vTfyy4SAYywI1aUW4Si5N6OfH2
fXof2XmHkTN/l0Xpauk4SKaT2qrS48fQFdZtHT/uL5frzBXSj4XCF4Jf2kVxc2LlrEiTj7lTSt0K
0danbC9oUJkVQv01MAuN/GiYTSLxmjqinQhP/+CLGttWn2KJHeXH/gCH+nvXxeYGtOtoXC4iuFrE
Ip5LL2DOeylacy8XMbsGhVtqxCLMrxpzOP5ihFRT2axhzABFxnRHr62xWP7FjIjOKaiORRvvDJdP
ugFY1XwaW7BOyEKxOEiE1rWtQdrlQQZisWFaJJmsjFgPftYMJlbF6/cMSYV4jbEpARsJZOJrmO72
ECZ9wtH/d1LRx9ImcVEmoRuuU/NDeARJ2rQEZwltqYisNxKOxXFhLDy/c2defjie6X0Y/pR8V4X6
N+jAeuBytv34X0FpA4ksFD0uNiRmfaa6mOzN6MWlM6D/emtu+xldOTt9dXVWVs4V8QTBHbKTTD8i
mDGF7Rspncu3GETUKXiuKQSdDrxXPlflkATRvtxyFnETSOQ5PqVArYxJ8A1EosEjyKVpw25DhXan
VylbrYbdIyL6MvAh4m56LvcOY27PadyM1FL4xyzWPnRZqY6L91cH3DaoEr/0xH0vDw1P9EKcGdfa
neWkdLRvCkwDiBoYpnLwkCGoCf1ZJv8Jr0PL4bI2efJoCw2aopT95pFuckTw9NmMIdB5ZDyMZTgG
yaYB5Vi+vDW+2VFq4AxlQtB/Ia+PUCiCwqJevTPjrUjVYrPJ71CYkfxbIhDJdBfnNwLK/VH03imw
WPIx6MRNTifnrT4Rrhxacq/3DzmrcRgS3th3ihPAdvR3YfHYknfcSCZlrJ7C+pJgdIt8QQ6Y0Gg1
CQddeJl9FT54MNQ88y8o0e8gvqDC03CavHvDLmrUWfGbouqvfP65+CTsH0zno7WXJqdOb8i1dr0b
ufRSIrIahQDEksg+URZ+WF0PYcxMRWcOTUrNgExHR2PNdYeiVL/yW8bMpyaBe0YsURc7hlg/KK0p
aXqKm2wQbgmM5TpEg60fnMImL5H+UzYRF/ck+OYl2lddiRIOsOR7RQjp6wv9R00DZnq4f3GEltul
0nU9PyBIwaypDYDxUBz9k/eHb4G4Id/tAFzGEFHEGN5bn90bKz/GiJ+n4NZvpVeBJUcYAzcNtr+m
z2vKGHLF7foWXdxio0DzQHbdI+u8Z4sgfz+PgghZDxoHtdwIlw0KQAfaenu4uFTL0LYHpWUTf0uZ
e8yR2FqFBtaZ3po4lOr7eiGUwap80RdBuG/ibjt5kuQxqj0NQMHp1ixp37nyCUlYr2TA4u28zNcm
mRw3BoLIaUfXXyDjDVzT6HunuBaBVwGmQNk9fDGtMW2iPj6j2SKj6mOoEza0gaULjgEhrfSutAOv
y3HCSVZXzU3WhAIza++iM381G194VafDhLegHHgpNAXxMBwdWulbiEIEtk3hegxvxq2iw7gm2pyB
JanhyqutkY9uMA9ff5sQNwMCe9+IpaqgXMclpL0z8U3S2mVw/T9OPGT02eGouwFQ5RoO7dM6B2PE
qY147ozRrCDV0BYTZD5qqGNjQQBzwpdYLJyBu6+uZRIKYjQFEkfd29jp8L+aHya/8ybXMeU1AoQQ
wno7irxjPbgxVDpDjDRY6dPM2rOjQ4I5Bo07cMWlVfaaPOdPTk74jrMequvZUv6e0ukYQi1Rg3+v
xSdS0yE3wo1KK+U5O8WnpCEu7iRwfu2v6do/z5p2uLxQRztKn4/2QLO5shcrD9dslNgmBy0j4MDG
sS9FkjeVuKH3xyGQUW8WH1WMP48bmNYm5IkjS2SmbHKsd/nYFoDTKuFa+DYXUk9HkN+VDBps256B
h9c5KNtQ/edtfihe+x9RKONp9j2mo4e9XhG35SjkS5yx9d7vjp9koRnldRUqoM3IsgS1vtq7rPXY
EZvzvVD0tUPvzQ3qDSsKXOo5TT3VjQreXrLumrYwVaBU5HWd9pFbE1DWOZXfed3utsvSMALgdMWU
rkpdoCMj+Savc+QqRH0t5RiWvCn94z5etoz+WHKrb+s435xcq/ewUTqMZq71LY8LELsXimdtdUdL
e5Qt4V8igs3ZYnGSGwJ5AWz8yT1Yn6bEkspY6gdoQDW0Y6PaVGK68R9cLcoBCiHB5vPlVJ1tlZWv
oUjEEaZED7/H5TPaRTavDlUI35jece/LtCB/WvxyNkJ/JYv/orrt+pd/oVRMmnWTRz1ePWfbn//9
ZJ6FbION/eMDzXlNbdfQK1UraLuaG3/WMJbartoucvMXq8vdI743KFuKdAN1KR+ixLtosb00sDSY
Qy6XRbdZYLSHPzePILOqmiKQ7C3x2sd1AjrG4Aj+sLSTAnu9sdBjOVUxWnYO8D60dzieSgouGCqf
Yvjnt4pMmxc5vBSu8r7RCNrCK0u2W7vBrc3cejZldO1b27jT+fY91Jk9SI+yCezZpfpX5wMWB5zE
Kw+V8K/MWLIlRAQB2IsRAfGNQdpNMrI1WY2ECsI0FLs3djohRv7s9oJ/r/BjTVnoqUT4xwuVuEO2
RZvsDs/+CDCkvF31kdjQyTLaDBP8nfWiHXsgmOTKD103y5+B+XdZb9RxQE81JgjBQ2S48O6yQNQ0
KmVPb38L4f68+SnOoRnYMqUxZeUnlAO77GRoXFv2TpvszhPKoo3c20EVWWEMa3rwPPwbYRtPCgD5
TE3a9cXarnvku3qB7ZuaC0D8EZJ9uODDVsqD1619yseThu1fG23mW87g6G2ce2nDxut0DZDUbneO
rGdqLQlEygYG/1O1xAmsAKBc8CbrUxgCL2yYc++rl7VIHGmMRsbuOpC2ifklvaGS2Nf+Qz+5nJ6p
5NF6+hI3tp5OB6pShlnGE5aO9DCql7Q/iDjA2Lob7IkXxy66zBeGZuo/At+50vcuUmkwUrZrKznU
bkZNaObjHOG5ms5e5UcBrLX4c9hZk/z5QzmmIvaS35st3VOkhsf+gXfelNqZEQZ88gcn4G8D3s0V
NQwBYYgBUznHMM2FeWbkoH6tQ3Rl/HT2B6EDVihKWk2aAD9NKBWP/7Rv93kTFSCOLcYLXZ9oeeMu
XPDKQw/VkSGG4dIpG0JsN7n6Vzwi65eKdDIrRNklipAC3yW6Dy+rO/PHantvQxhsroX1+4H/MiGV
VsHLTOVL1oxNAfwfOCWqysV3rU2c9VhyhC9dE0Avbj5+U8l+dxnQaaB7Xi9PaInHbbbTtat9g5vX
BZmfBAxdLaqfIsgwq0ep8cY/dtrffPlP0VKPHXrrE7EtGftt4BSGEZno3o3jak7QMK1muGavalby
qqaJGM9adQAd6KuIKhsp2Bbf2XaUwmVg7npzenZ+0m1gXDy8kW9cS+D9hsJS0RGc81Y9myaZQRjs
1YuNgtLMZSMFQzcJZhioPy0CIIOBzTL/TNw82Uzvh4Kt05Qf8uIAHd/dpErj+VyDEpVC35g8T/KS
E477vYxJvX4Xx5MfW44cEHTZT2ho9FtsSVMDLQyflOtDE8wddi6xHG52CRWuAwAmosiGslYlpqqD
hJMUu+zDfyxK+x+zXV4iRT5f91AOSM7GxR3AN2LXGr5mr4LB4VH2NGAmLYxTsZJSuKRlORkFRSnV
V09ScX/UEw/c2tSh1GZUn/YSi6hq1c6DRLjKvjNpyL6qmBSnuyC7Cp79IZ/j+1JPXUXvcjL/Cz6l
GFBNnpRxVWoRkN5XfPKoMU/hEqfgG4tpIfEKfAaM+LfUrK7kscHHDEY1azi+LCaRazai8FM7mxZN
W1VxKykZpVf5l4gjsMb17aFf5p1AHjGJ0Ktn02vMZXfnPHKxqoMcgLf3MUUPNWPulOPtDLGda7fP
aGwUrAStiBYP+SjRWGXpbCGdFb7JEkXdGXtbxeb1qImG59F1syBiQIFVTtJXAYwoXtedCBeAPsvI
LvxmeVOchmv0Pnjl21cAvr7loZco1nFVx7EAfc9UTikSb1SMnGVFOd6as1wtjnIHnTSjYXoOVT+g
+ndJQ7BSgaXktc9KiB9/KZtDgBBOwYLIdEpn/CJbR1ngi5jDN9VT6BDMQ8wAA0jn2AaOM6EyQJ/D
y5YWmpvBTCNri9X+VwROcZSu5ZDCdRLkGZN9/H1KxvfnKOgpcMmEewDEqCCzRoRnUeEBbV/F1mRh
hnVv8pReSxvnkc4LFrpELboAMBSoEHw8Yx4w0WayPzngEitdR44qnXtRdaw9l4hxgAHmfCXQtz6A
+ujXA5eOxz/wl+iF3aJxXkQ+rofxPlqL4mBQg/+cnirkx1liyS/1mD3lca8o3AWnkghJeMKosN7X
f0p+nNn6Lj1YIA8zB6bCfOaBDYXQzEby2TBUwsHoexUv2xMKKx3PiWxl6Ra3fLuz4X+1qsMtqLu7
KIJ1p/gFsLXeW/ncKh2kqiEgmRCUR9J/xmf6B5MX9MMmQ3f01gl9Zy+TB5UdYZAWeYUUKEtI3rsY
CmcWcAaTh3gx3K5e65PRN2t4a8Ew0j4/Wk+edeVXZbEVn4/KWGhhHmZyYL9ltXyoksuidZAHZ+XL
z0pFbRAvlvS7PNdA588Ab93xjYsIIQDalJ28mmXmSfkc01K89HNu0Rv6LC6AZhiAsEL3Y10rCG5F
B+QZnD9pn9Ec4qwFB7WMcE08s5jhvsxzkFlR9CWEPhlBBC3PaCWClv8wjTn1HIr82l/YSStShu+0
hMOftZLvAmc3S+POP+mQiYV/RwPJBXLMSqhJayIWiE46Dtvbc2Fxeq4CukqN2O2JGXAvWdH3gc10
qDh0tXfWJguCuZ4uNC7S/jXxcyl4/8g68e5uC8oCZ9K44i6L3fO1edAfK1kncLnRX76w7KtMG7nM
Fp8RYGsOEhwpxmZypoJzTZRfmp17tQ+iqZCymX5QXiWWNJt8jAlfx8NjUxXeRy/yY3G7svYVWJvW
H7ML6Od5rVbo8u8uUOAyAk3Whcl4jYRVdomJRp1p5hrWc+48XBmVc32ZXcb+pNhuuKG0JqZOTPT9
ZoiSMajd24lvbA15tNlRd+5ZKnXaE9L9gsST1bXtQsiX5ggjMpwv+kZBl3Bq9K88fes8gM7d6Zo5
pDUp9IbAXjBROb0W/Lof7iJK8yzVPR8D2IGSjDOIBa75PbPMTZK4o6ceEif+zuKjqNNoEYkyX3HM
Kjtu+dzYR28JMVhJMG4agv6W3oJFuDz9hduT1hTHYCkLSE44x4u3l41hVVA71DvDpGAqAMe819lS
tdY1NjLA12uz5vu/onIXwjww6paDXK8CoTTJolQQZGgQkXusujRaSJhzZnGN6ZF+kVeT6DkHa4km
5jN7pNv2mcSNVw/QflAWhrmarGPYtWv/BHIzZ1L+tq0IBpi4uUEVfInwJfMl5gw/cGWrpfRlF6QT
g0Bh5qUtnDew5riydqJ8ipUX83bGqThvrbwQpoDQEQN4amRw5JG5mjxUk7sk/31408LRTSg2zvJa
Q/+HYJq/+Gy94b123QBze5KrnpfCxm//OzL0auVlm6cfjeQSXoHN3WxVcvc5CtfxH8dWIMHC70V4
yIkTe+/GxefnVKsNA0PM2imcsusHRXHiVCdla6e2boTXyBEBnm0SmzUxnn26KRN9MmxREhTjG5/i
a5IkRqv7R3VxfcLJ5Lx99ycWEwsYQYHF3qbKgpvWDcR6VUQp/WjvFFMCHLsyJloXPE2fEkUy8E/C
/pHz0UOAcBDNDQOyeNLZSZFkuhkpLynk+jPzd4sWJxKCoTbPMoSpvtx4CuYQ2bb4xY1sZJiiXhWa
FZmPHzHRhswUnawifsezpKt6R40a2FkOn4yBlLhPAxJ9GJ0lZrIelNE2hWl3z2h2ICtAEjXHeulT
3fnnAhDsZpKS9Zmm9dR2IPh7FlV1ZwCgTFD2uSZ2dJQtMr2vocMfpCdaUc+HMJBUz41xpCEM3GuK
56KHjHX7AX4CJyYzBkrzC5Mx2ykNXFYituoU83sMFAwX2mCDqUf7U1/dnHAF4E7l7OTIssO+9RUB
VLPAMvzOvMAAPXHaPzJCLUXyv9sGLYLaVXel2ZMrn3MY5z4lYVCr2ZaCF5CyCUZ0vFNwgcMElDIY
TN/UccN6dtVuin7b9gU76fICTboMBcB6OOM0Bx8cJKS19ChDgwe91dQHcKyZlCgFid7bmbHFMSVJ
UUJI9Teowi9lTtfusVqb2WoS2d75H+yUCExg8XX+qfvg/cWwCE11fMu9IQT0oZuzhkZvyaa/nnjj
o03qo0+JfeSk/oKZ7wAQfEXD5T02DqezMqjTvKW74yFyngO+KcNJUIfPutjZVfQiNUjdQKekBK6S
rI4U6o4uvfGr0/5bZJQzeeyw7w7L6sP7rfpI8x3BWlecOYSWqNOZslp6CQtcUju8nq0U0L72FXRu
3211au9+cEAYrKet0Q2tvnS60aBwmgYC6YXGTHf++a5ObmbRd9vh2eDjMc4QNODkhHE2/GDM2zvh
EOa+5rTwlLJP6JXt8pdznBlK1ssjqan+hoG4H9AxWnn2Hgi7kaQgV2oEQyIQ9b7eQeyUUucLhErx
5pprQkv/Gu3L5Ig4cus50wy4NpwABghLice6TIG3YvUqybxr7BehUytZhlO39tcPA0NXOFY335fv
Wkn1d18BWIkSQO/knyQjzPvJRkSEYK79kcD0xaMuO4oIzTUs7Kf5MAyAvYSbEmnRADD+1gvwie0P
IJr8oeOyPH6buhROPO8cGvSfWKXtKM8Vk5xyagommxIVJB/aa4ak9FqKpUxfqzaQMNvwgAP9h51u
XQTqvA170/4fDY9JlzBeSAdeXuiWhmd3aBW3viv5bO0JAScygpSO2RKLkPCeUMIqQ3tIBa+Ik/Iq
Uxf4S5c7NTH50MwjsvGyK6jlTEiVP8go65g34E4p2zV6753Pv6nVSc16sGdJpIN/AKYfNZykPheS
71SCwIp2xPKTbodjVRbCCuT0FnDgFbhqRCPZqaJyD6Ebwt03r6B63Jq/oYkypaVL526xgS5Yd8Sn
Or/Zua5BHjBdAEm+cKcwYlNQXCIS5rVk8JUalMkpOudhhYmceCFEIynvtXnAGtoH4rD9/XeP/e3o
ymF7lEAYL4RWbP1J6gPo/YtkLCbJDOMLd0lMXaiXSIZfHfm4Ws42a/4TIJd3SgOYeDaZYkfHsrKn
znneAXGov8Y5ARWuiBtEaR9NutjXvvZl1/HkHdXZCi2CQRpNmg6nQx21Ky2g2NFIHv9DihBCyOcW
tJVQ1u1EAYk1Fp1jJpikS1H6vUyPuoOPpj7Ge2UQcEc0Pbp4936k76NRoqbuXxICZS3zlv0jyQ0p
t3wAfDJm+WIOyybwXo8v2SW+OaAcAsoYY/HYpqiq3Xbhw0fPdnev35g4OpmW41rhRn9dU5nARR1l
IiV8irjylok0m5X5Uih3OWjyHmXU0OvgeIaU5gMtnYcqmxVp91ECrBRSXC9l0Ve6EidXfj6w/Vb+
8/44sTdeUzsf19ZQSVyV0IC+WktIuhVeFGjU0EDK5YaW9LOmwjQCdCvZDM23p5RC0lE4uXCBk/E0
UK9O4QTMrM0XNRpMMGmkMsN/xSEN2BQ7lhenYxxn8Nium/34kYsZDJrG1cj0HCCHWZrWCTxMRm89
dUfsLBwfMDhvaW/+fpsXrsXx65FWfGJKq+79hELygyqYSaiSq9J8Tli5nSGzmZ3NCVahJ0s1GJMB
kYE75a9Vhx18Ulr2EerR7zxZddGXFr2We5mKx8vtpkazXiYxkld8QWBnTA1/jy0uEj0STHu/UKRD
kkxrzIvwBLjlokDi/Bal43CxxkFtIJ/mpVPixuoi02MysdW527MpDktOD4aKVcnQWE+Bg589yfFM
WgpNFDqhyQa7W7cZIIF67uBgMWz4n+QkWimiBRS5SQKo9107ZbVso9Yv4aj+dGp1b0qK8+Z9hHiI
SxZnG9pqJUFVeTRpioiV36IHrwPkKFuRN5/BXqyOFSN4P7OyZZXz6FaGo8e6n8o3Rmbqs1HrF60N
jXmWwjnsMCGVeT/Oc4wvkW1GhYfqnB+XgyYuqwtkq9aATph18Han6h9rqWD+9xNpMvNIfgrr32GL
i8BTwg7eruGxB+3Tr6UEiCwcfBVPHqJJPbSOVkj1dAMtclsbOuCi1pN+peOyHwowsvWbMLBF4L+J
Fw3vtjnDgD3Aph3nYDWeYR/4nHtq+aUio9HlZ5n0rlY9komVb9zWqSg+iH3ffuH6pCAiW44Yej2Y
EdOpsCzvzpCSwEKVr7o0B/OFZnu5gN4NwnLjewc+ymXcSFz9E1gTxQwXGBjWLkxicILUsrZ3BRFP
gUSbpcR1J63slPzZfRvQZEUmh/cmFkUKtUBUNMw9FKnkaxzAXoiAk6LZqVvklUZYo+VNA7DrO7Iq
Tt9fbfshiGR8iPTyaK66Hn+FCOp2Wx3PFt91CgGtUCeX1eSUMWIQK+x7MofKaEqDOmaehgikED/i
ZzY6J2TXNihQBXu/yAAVtDmtqG1WEopGcJD63a8WNdxvRwx/i1tdKSRSWaeBu7v+F5uwfJDlVmXz
ubVta9jZML6NVrl6Yg7nV210PX39T24Je9bLSXtpeHW9zn00N1bOSc0RZfRszYkpUxW54IRbkqp6
nz/5w2IpLUgK2GPFRSkN3O9BcYvRVE+i4XZMYLokEgwTJiaCCESMqXg2Pkn5n87W8GAL+OcDhBHv
iXqiCDChipr8/ko17YQyXiloo0m58ifYYjhX/Genh9g1U4k7n+/MMwqyBHUARp9pR/y0siKq1Kkl
oWZspBXRNsPo/cFjqLs/lGFk26VpR+V66x6/iWfFnit2O/c+v+zxwFDitQhiMcpAd8YiMU9Wwh0s
sjs6B8wrbKoViAKiW/fTlM1OPdw6yx6pPQu3iy8tByV+wq9d3KhzZJrBKars84gJcttbH+CUJPUT
s8J3tZsVp0UUdaFLlNW1hJSiocnP71dPe+1J0OJdPUq4324I/SNvjYnz6Vels4HyxwX7f2mm36p0
iyajzAVkALEH1/icLVWQZJEYuvwwvfJTiPzu2nFks1A4IwvC2mXT46Y89dPJ3ca1eOWtF7K2KJwM
D9QDV0BdxNGQ4AN+sty6sgGCh80U0LSC0Nudv5oa4X5+fHMd++wKcMm2HuyMmYd6Ph1hGpKYL1P5
eu4ngc0WdCaDU1Vi1cDFCu1p3et17DSBbfv1nf0viiG4F+wNyCUHDFlzylTfSlAXce7Ck++cmLaF
OyGWP1sSugKu30Y9hMI61C5Ap8MgvKjvLei5UWUJ7qdKIsf/VJlJK5rJ5rNkA7yByCpc3nO3c1kW
U3UVDuC7CKfhxjMgglPWbqQAPJHUG06ZEHYefiB6pxh2J87QLm2yhbOkZ1MclrcSV/vsJQJ9GeaA
hhxB0UW2fuXt2IYROorby+sWdZHHHSp2u01i244KGaq66qvZC0/p7ogdE1Y0ptnxIVeS/vyfOWj6
8JMrd6f7CQeNoydW5iUmJRTMWgapbgXJrjNGxcEBXYGA0XQgvsH2jKV1xQg/ANRtK7RX+dVR+gfX
u6ehktC9N4CXsAP4kq0lnVkn+bduM9nF1NF//UyIvc/fhfbyy32CZ5qgfFzn5rn0ODpGi1H7qfzV
QXRh0nb9LmSzNglQ2zqT/VjxgchVdyhx+ZI5RjnHD6ukbxFxiVTVqvb+Jdrjnt4F30EpeF1h079p
51mQijnepsYM1Diy3YQF3fS2qkgq/xpd1toC5uQPuV/XoStiCS6Rg3uniHfxqCAE0GT90mQOvR+I
wqEEisTFBdNKW8oYmrjXEKzXjFlLeERhZxxtrQfm5/383HJ+xmwE6KgcUM6GqAU/E2baQZqL++Dn
eJgiClrMkyP6TJ0pFYFZj6cANiEDwFimbMiG/xzeCZ7CAgw0KCVTTe/9OXgC1u04maTkSb8nqrNv
ksoq9uDADKCVIEfL2GB2ga3Uktmz2TRIGq7PDGGk3PCDgyerFTfKszNX4IwLtGmmwS/gI6swp7va
KFdRSpGLtEw9QqUVfrKp2+ShpuMXFUkSzwc7CpZM0xy8/GZ21Ds8DjWWvg3LTWswFs8bn5R8eq8Q
VzsYhdL9/ivC5za6Of6ZTS0g+aUqIt978zivw7Si4OTo23wQ2My+ze6gNWOD3FWiXgW8sIBjaP0w
hY5QtBcQCF+FUP0H2m9z21aDcwT8AUSso0k8Ti7PBFLFDdsb39C3tDt7chfuAbzhqZ6wsIqCHcfg
CVRhG6VUWI5f0Qvl5FVWHv9zrDXjVs3mIZLZ3uc6FX/D9JSiTi5HBvg5XAcO8JrrBOdCrYtGVg0u
lcDXuYuolzUBOnVgEJqomHVgjWb9aDa/Fp8TYEFSJyEHw6k6Nmu7rddwObL0UgFoKoD5UeSXDQwO
MosB2KtJR6nWgsZHofw/wMCb1vyBRZyaYBtmIcJhMQD6DIT8kb78503RMatnB+iy4UkqRSWtLEI4
FcqA68KgxBqDZsV903YkLLNgK4N7fourDsSgF0pJFF1mxfqIyHhdVqk/hX/nJrNAjP2/zSsDlNPN
cDYUNavltg2eeTRP8o9cQRBsegXZrPePVcqaDZjJG1K2IO0uMkoXuItgR1awqTqwgm7hHaVlZ/Dq
tqSvJwcRj6twvT97x6HrNT2c/4MtTuvyiwZes1bt6kviG/7/2ILF/KVgKFT79xD+LwTSzlZEcUwX
DqkYJot0eQhqraaXtX2QNiENLFzDFTy900RNAeLpRvAluujMAnNTXtX2N95qgaQQHOFbBoVhRQT8
/O8pvMBa53jVfL+sqNwNtipsnpyPQhu1I+aoNuCXJiYhj0gUZm4z10s+oARtN8hNvBOe77oOq9Sb
2xGYkVhBtGEgjRvIhTrfM2f9Jkn9ijcfm/5bKGLj4u8WOw3IGvsGFeus7MeaRnh+z+q0j/xuDLwr
/paL1xzq+K5o2sv7aHBs8fohYTy/ikRJ/VZ6QaUC2Y1vG0mERCzq3PDf11RBhmXrbLg6pTQWvQn0
E9U4/AMTraSsmTIzCULVvLOtT1WRejcCJL8GBheTr+kiGKEGiWdZQEnapcDCbUifXyf3pbMkXFwg
jWP0xOHfrqkYkJzFDY91e20CaR7In3Bq05w5A5JEZCOCwWcojg7+kka5o9iUg/MI0C0M0qXwgI25
WTN8W3Y93WZsrtw2cMslGkxKJfxn7QHj7mldaDW222ATsAFo4+hW4bw8YkVnPuowPd3zIbG1zrhv
rw0AKrCaPUDs5jwAI0E+tjl9wVadth6rFyLmkmPDuRgA3iG3rECeqrhX1jKtAH7mL5E3n9lOO6N8
pwSQJXLKwKcXycyKfb2QiAhX5AB87TbGcFnDOBabp0+VJO8QLcjx+17A91SHTpRfd/mXzuWreM/5
jHQEnDD/YvqcharPfwS2BRCKEz9/0HQtIUlg/2UQy2/SouS4CX3ZlWpI1aE1zoPW56PKI6dc1k7R
ozx2iG3sO3xZ7QHU6jIkp/+rhsQ1LtSEk9pgErt74u37LF+VdovOunKMzf61sY2oc9bZ0ZcTPfW5
JWfCXpDBlq6Bmar6pzjvdl8BI7k4a0VMWS4Y37qJnf8EGYErkZ3MzoyusQu0fnXkjNqk9bE5MHbW
JvjNAc9Ly7FDiU57853M+9VVGSKvY+XKRJ4Cgim++COdT7P5ENQnTHuWCgNbN1vT6MWRtOK6jqo3
N2esex+j2/BhAago8ot8X+WfnzNQ088/Qf5KzljBfuw27Uo/mJeF7Qs0AoYT70sD/I2AtxwfVrKx
LGDPKKiRZalZD2vQW3glvDqAHuMzR+D1tYWJOuIrlCoX65KarzivUntf0NGJKVbay1av6iIMEq3d
8SAVgj3BOyF/YjI0e5o0HfSHRSL5ZJtQtphg3lZrZiwcctYxQIGPAWz3qArg5nSHh62LXTV1bX2m
0+VfrQ18ve6S6AykVAbtU89IYBFbtqJ1szcUoybeYysTwXu3JWpcm7tmpAz90h7WtkjxgGZ9bsOx
d5KRuL7AhOhiewIwyaph/Kkvlyrl+cR/AIxP9dbp1A84XZpqZuf9KV7fMLA5msgVfpEdD9B4HEhh
2oIpw01BeBmDbE7Xa/YqoNgT5oyU/z3bHQsz8ZiZejcaPMbMMeNBdfzXzM/V2WgrIIqmMYcyQHgk
7HWaVsFUpfrz6cwxNf7++Y/skRokePDVOOJlz2xAmogGK5moscU8KXhFNi9F+HEKghlqDZMVULRw
lz8C7c2v9LvEmeLstLOuUrBFElxWE8gAPRmkI3qQfVvYH4fQhn4Z1aK27DqbmIIEhDBXlFAE20JM
l55pmATt5WA/xvqoQ+V8HcfBPQoqGgaio6JfMMNtJdDXsN7sQhG2mrvu8uvIqmEhUshK8lFr4cuz
+KNVtGbVHGBuAmc2SESiKAkfxl54LyA3lCQpdFHOA9S8hm4jkNZ9D+ljDenrIZh0ZEbNDu0KZ9cq
sRPZArnUS7sWaU8tTHXjaPON5zIMmr8rzGBDc7UiqMoglDxZgen19xC94+z1X1t2Aw5ydGq0VrlI
a+LyAh5bM16H2USULRo7QA3tnmuDDV0bKOpwnUaeS9JkFwc7mpX9Dclcp8bNoK9NKVxiEVNg6IV5
m/C6B5ykImN3iPhwJ8AZZz7jX2PNqT7c5Yf+Rwe0ulIqtfxThzoWRPjuYFxeKdYdT33MNhpV23Mx
lnOzcjA620tZpJ2gOyVe19GUcBEVR1BJGPL9ISCzWs9TDr881DeZzx7EZSaDXSMlFOZlEkMGxbLX
gB75eTS1hnQrS4BR61MzbGLKAygocMF9vOR/Ar9ESTAmRbsuJIv+TpuM1DwM5Vqy/O3bV69fjm81
DG+VC+ru2gjL4rpKIibzdwOIi7SjvxJR0R1g7b9NuABlKcXvTaOIzuEU7OCcqmpHw0AgoQbtaxWy
AEN+NGGos1KERRSMnIK1TIPXmlvgi5QL+e7anUyd2c0xKmZtnu8qQ5ks+1ibqdgnqi/1ffIgJpF9
JLcJiewoucZtvW9SYUrw9N5Rv/7RWsguclID/HLSCPufoZKQ1VANYhVWKQP0yNw2HKDHet/BzgaW
JLdevXAsk9/K+5Qo2KN7NKf9ICAEQXnWiZ2mmUlts5WjSj5gttRSshaaog+rR38OWqsRxow12nLt
7cEaTXHOr8tUNky8lVXGyelS/JJJCCuAm0AnlLKRfrF0t5EmI5yLN9CWtcgUUQNP0d3M+pcXskKx
aMkJWr/hu0sKvdQAeoDNABbTPZURpf2FMDRaMRtXmTJMzeWJ/VPRqPIgQNeGKlkkSDG4qHUVrDuW
B/z9d5sEvcL8/YP56kTG3NUhpBOzH/zsqgkHz1H3HyjgwMwviYdqdMTyKCJNYM1L3YAOrXI4MEPH
7B32xOziXhHe1EKO5qF/NcDRFIFqtzeEPL8St5RfbiPTmM569t1yzEZdHP2Y54YQfewUsBUfuoAe
xER4A2Fo2kcOHPJjwVIUJY60OCPCwWP5pj2BLzCP2vtSZtSTSXqIeGixhAcUc+nxNN1JPeqIsxjk
/BZ3bySKw74+yGwFu35MAMhLpRm2e8hq1aO/4dDupZ7IWqAC1P196f4VH5BB783bv/U3lYaLa2MY
+PxSSGSfo8AsxJMY3HsOfRzGXZoMWHqLmI7OFzepo3D5zbY2IQGrcX+VhGUbTojNKZuauILLE0JA
y2fIOY4huX3bBY5J8KmIsV008ZxdfwPvL/CLdQj1LMzlUHhUXYHR0z1kTAvzG41hEYpMi1H00PGL
qUHRNQW58FXXLnq1OFJcz80rqDUcEnQZMZbBMcgC9eovI2fOZB0Oo3XN66zF9tURFekTyi4QKNVg
u2U/1H6CsHgoAkGDQ9CTOQ5LBwj+l9L5PTn5tpkNTgwRC7kIZQ4a0Fh0Cae8yTtY9ycyT/0zJfZw
CX8t312V9vAUoj06XXjQdgiPprw1sh7xIKqg21GcvQyLzq8JqBjNwfO+gVItJcAWcuCaUgecJd+g
sfgHNOpNSF4Kmz3df6gz2+nNP8JMLrRpTBB6n708HRmGsTRuqsoj3DxiWGAkFxHuSH3sqxKHzwsY
rVc6k8a7YkkstJ4kH49l5g5Sw04RmDDPVQRO8LezuMI6Lymp39h0JPvqriCl6NHA1c1ZYUL0pI4a
fHEPI8qlrFKFNYwWeMN3oc3L7hFjrvjY06XHbOOnfjZoJhvffEF390Z4/oOy2AignqHChqn/aAxn
bf6M4zeDDtAGpb2JRs80SmrjvPwsyONodNZkWtzSRYrKas3H60/Xd1yHw4UWB1zdKDQHG81CZHfd
P9+P2naKxXeuBuDVAAlBXG8PuW8kxhDTpZWTF0HR3F87USAtzqacvq/6OqajMSxDTBdTTrDgQNls
LaZGrCk5gc/ltbBN2d/lndCHdH4mxqShaWf+u7QPEnAyZL307cVHSc3Ul/BQ2BwJj9ReC/ZMMnnZ
t8/Q288nzJx+kWUVF12Z1QDqfphsItfJ+DVcTrrj9IX+oSHP5kClSJKUA3MEq/z1s9TYLSHoErUV
xwf/h/fFpTxDWmolb2DT0iqD1nj0IEQCMmoD9F5Y/HV/DPaJGZF6nzXdgoEWfKrWblThYg2CNtq8
v2aOzlmGqSndZiIELNg7a0vkyrcFxk+gjdQWo42fQww0kbzLK91VIHDh46wNljUTp6NQB1+XDjEP
U5ISV9/coo2gvv5WFWxGr32eWEwuddNZeU7ZZt2bzWxtTWRpTAGxLjiyf7GLEvrjPSSTfaUIqg+2
jJytoKgZvMQEscaTV9YIx4xV6uJ0XLE2gzZhgcVYOASC6fPXgDkUMjS8XXYYS6E19mim4eNN3A1X
IzApNlKn/pgldx3MRx5nlg0VtNcg0+ITNAP0aVmAFmcDfAetA16Q4sQpKE8GakWrixf1sFbfb7qp
16rLK+ly1Og6/j4/f8/wsYDAVTPH5BaxOrkFXMos4Olmrcjm7slSaiPrtwcNeAg32xkjJsKpxQ0C
vy0+cZQt9JKDiYyUy2WgixSH6Pn5EYc6RhKGrIO2V+6poK6vuSrllAbDepiI+RvHZ+AzH4JXZoQL
tUElr9OljZDoo2bajRPbZKfXv+hwuzH4QCF+5ZYMJzumkDNumhnZ+2TtX/8x1nxkbfbi9JSC4Tal
wRj96ziEwhZH65TgQs3V/khL/11+xDEhgLIZWhFw8oQyoM2WRx9dW4PzwNpvahcSn4Gkwb6UxtqS
4UM2AXnfBsjomOfy3UZ/UJreYFYzsHrEXV9taa+McE1KyN7xgKvI/Wv2mF8VDnK3HEmY0fbaoM+M
RUhn2rmzT/yxmhrHVmT6phnRJ9g1KHP+bCJ9VfA2BnSqpyEZQtucI1AeWA/XEkpAY+qkpw+bxCu9
70ftDUIUB2SEUS9MN4gZmBnSLuLDGsk+XAXnYkO4cHEDb28O2cX0V73Hq1CPlfAHENVlcnAeEORg
ktyM+UjrCTD1MsxvNXDVjq580ztwgZfBC9gKEU6pTnR0z/5WO0JOJWqhnsmWWHzkEUz3PuCrFg4I
XkehjXpo3787xyVcNIp2ITJY+VWLTYLsf6B4RN01ct0OYtpWBdpyOa9//Ze/VJkUY/9XWold1DrH
OyxA56+FJ5W6GgcC719zmsZnWq/s22uoZqbnmwCcDNWZCVaqdZzD2oTL3EKIOpE1tmXOtp1c+syR
NY1mzLd5YAJ/GkhZQZr9i0QmRNyZN5GGMbSowQVa9kqx+rbz/A0lItluGn0MRW6VqgeletBGw4/W
sCGRRVqUsAnJ3ilEzA6rsdVW1ZbEx2FDQgwOFEuR5uSYXeckQM2BMc3zfre3a4FN5Yu4g3leusEa
WLtkGIFwQ5rQI4vrBsAFUaLH8M3KSp9d0STC/sAUBh1US9EplCktct2sm7BKrfiJpknXmZbiAl+p
9Ne0rUOfew3ZgJrX1fYWgDvoT1ZbId1VqPueIy7JpJKL1wE0LrkvX10sCEOsWwr4UuunZRvwqSt8
T3S101Nnb9bxjgdFIonn5l6uVUeqLD7nGHxY9is9oz3klLuOloTg3atFDrNtNpv5EWEt9O1fJoyh
Isin9FrFCjitligg9H4YtwkoA38urVoLGJX5822A8yyhlIxtsknrl9KPs/UTMKq2yAoGs3ucdS7F
6263uqy2+kd0mvDbHjRRKeX+QHsv5KNO8vYL5Eu4g3BCZhg7n48TsJsQVVv8mG3EM+4GavkEWwMq
5n9Iuh6Uj+1n4aE3QgUJzedItMSbUsauVwXgXJAGs+cM0WNGcPRK2W0Zp/7TIUWC6e4vKxJwIl4L
ylG5aTX2R2bZcQg+B1hT1L5oGIR3f6+BlMM/R7Y1uM8XUcW8094nowgyNyqvlJvmG9oZdsprbNbR
3IkEwGetJlO0DXJnRwlJPn8OkxgINdwuuBvO6xs4I8KQ/pIMR/H0Jy/JtcCS7W248jhvUFBaiD8n
LPfbMeoXruMjjRsgtklvKxgGgRp+pzSuv8WJqlSL0VXp7S5Guz883qFVaG1T/5BSPvjSV8VO7qDP
OynwnrThjoEduwe59W5e0jGBj6j5YTjBhNeOFCqmwFwxnHl7F6f7aEnzQTo2oFzIn+4A5ZzAr2C0
q4V5mbsoauvfpcjXg70zgjZWIM+HsL9xcj0/WLQAbZjjeWomJAkp7gqJ1OoUGfdhTMQnMZcz7/zU
8uL3UPrwJXPJPva+8Yd/ZKbCnBBV4EsVt3qmvpBHiZM01IJnjb3V7IbhRqfdfpS3nD70DcY04Obq
WL4X9H905+aT4o1Gu6h2SyZRu0UFlTjqDCMUfXgisq7VkUUUgK5LWWZ2K2hiuahmkiHA8zvnBp/S
eXoy2yZh9sVyyQm2fYCk0+3ZoQ37gmqTF9bq6hTvwjupkrnI0xXrqOQrQlCcXBLX2vpSya8sSasg
R1N+rogyZHDCtU8PKx+qo0yfudoCIG4gZ35pmNmVSBO6/HQySSuhM0cuBfRLPChMsSr7LwjjOCCF
zjI1mqIIxN3uBudysJ5lvvm11A9HkJNu2ZpBMxqYZCLYmnHUcWr8nH/45l/r58Jm5roBzztoeHTF
+RQV8QAf5W/d3BX43kq8F2K4jxxzM7GQ6OReVE5V/LcKg2JTUvVARcCZvxQPiLweG4/ulrpzA67s
I2icLSxO8gY/EksdbQZ5SqeARvhGb9Z6HeEABM53Gbk4XELMgLjaWpRaJwA74/gcFZbhr7B66Unj
qUrBTQPk9Jb+p5bwDHAIzKT8+1ncE/+hjSJXDipzVHG2ubles78ROWHqImUFIJR8eDdmk8KBs17N
7FuCzxWVYRn72mE5KcANsUV34DCvOzwSFYfqRdoCtGFbUqwJwvMu3lDW88LZDFyIleV6wP7B8oBg
AU3VdnOoh+nlcd6Sx457agKQWwr+yJqPY7HRT1EQnhAOutuL2pBeao7xKfDBzEkMLTZnQKdqLhRk
38Inc0EPF+kqYcsEMlqJMN7YdRICsffkg9ZjZUNmFt9t30H4hrycw9b8yFToSH3xlWCRGo3//CjP
sNBws61AoewSqooM+B3pgGNEJIaa5OSP6a0JI3R//T+8HM3SWwGy5Rt5eCrN6ShZViJEwTli07c4
VIG7GR5Mpc8FzEixnpV/fOgGAYuKf9ikIK0pdu7lIYGqJR250qNsq2ln//5QWy2ak5tT1rA/4vb6
706JDBjoPTzVeOvzKDGi5oE86jc2f+NvDW532Dbg4ufYx68xnShHpSG9IyXWZW5uiXHn0wy2qZYS
1zFg7DjQ+ppF2haoWKkiXfHjKA6kgcGjRWzfDuDPbTuglQarec7jJSo7NxA2whA+jMk9oLQmIRUs
T09+o2j9vjKT2dFf/cuFndHWi6mcXS5LXL3plM2vqOdP2WYWwbbMNWL6z16Ppb8c96A0ZDm+9Xrv
CGys0nKMJu1c3ONpFp9ZX28jXuUI/QIN90Q9Ti03QuGd4mnXSpg0X6lTz5dBIVpijPOLRUDW7WYu
OBuhGVKjxhvaNKV9L8i26pFRPRHQhyGB+YpgxKmdVi6ZAOrfib5BOCTVYJmHYa15269BqlOcoLfd
Iw6xA41P03Thd/QPhbNFw6t9gXM1NyI11w2AXgSe+Lbj+aDaCV8H0MbLrxzkSJ5CkI6/M2QxLwAL
3/oTZm6knLAcAaIYeMG/4qngR8fLVQBCN+xt709uyT1+6NOF7YjcRHn2JoPZV1eFlQfDVQS6/W8w
8ExCpAEgYXI2EG1n3zhYFQo2qW3mbYoByR2SMv6FtYlgo53qdximJQG0u9cGIdQdslRBRWFMOjMS
dCKctymbb0y4YSp2w/LBsyXElYTW6tRydIkHw0PE34u+OSdWjvy6ayi2XbrO0RvDcozBgjmKSPKg
VvTSBepvKy/Ci1JLAgGKjtODiNNQAUU6OOrBkd0oQofH3Ne2vRJIIk1rSQ+qoBNZ7AKlo03Tj3LM
Fd0CYyw3sSr7rwe7v0NkIFDYlztjFbfer8ZCa5vn0AAE6zTLeN8Du91v4IJXZB9R0WP+HpClxMdw
cqQBVz8LTiCM6v74iRjuE0UPCT2AOv/E3hGtkZzr2JiLZXbJeJ14yT412dOHqZ9vytmyCbJdLoHr
NYlVucZLVlk2brjmHeh2c7gDCJElyd+RcIhvQASfXL+XXxeYbCvzWN184inCzevZDvBP5ii7BcSY
ZtcLJWG6Xqau978L7SGXyZsDo/D7BAzFJsMu3tD4coCKa3IJ6qV9AsscCGdWnBZH8SAcqdlqRb0/
91pHkmNZ9ysEc7mAMDfYXEy44HRPG4d5CEJkhu17iSO45bPFmEki+jPb3VPB7yQYGORj8ckOpCEQ
lqYk/kRhjlPSmGuwpeb62rkA2ZVw2+0oC261Pf7uY0I1cYr5xAITlpfXTIMvdtgoVlbtNQFhYws+
tdn/772BceXi9ZW9POvm95pxLE367fvJmtXVEf3NnsOJYa5RjgzfW9F6+mOJNU+UgJRWD9GJUECX
N7O4bIfhUyOpGCJIFnD8ppLcV1IPvv0E8Ve2MDltFdatUXANVXPkDxKDdjmCK6N9hVzN2s6P+SdU
iTXClaLnevmR+RDBD0MhadupyxS9+hhgCJiL5z8JHxmBQkZMgE8Ic8UimkSEQPVTSoFzbphTeO4M
TZ5Elt+UA6hURXjS6Siy1eSfpALdoctrizlQoun4cgRhBkLCGqY3JjxpgvBl8H5CAWImQZiRx1U7
21yvF9DH97qyAKgwydLZFu2uKAmy6pARFQbUfmCq1Aw9j67gmnJxq1DBDp5ACMnTPjfVb65SzHHE
tFlHV3vtRKPelE/1193RsySSx5csU1Jc62nj5QL2w8erwdOcvWjNkYhGKtRyrmTYb+QIpw1fWVqv
Fl2TzslOR5DMpELhn8Pz+bmphVnSf1X5nkl2mwHXBSauhvpGX4k4Hz5uuMxrzxp7C/oZELwiELEv
9Zn0eVMXYlm7IJM1DDkPPyAY6IejASHuBA4d3qEfIgWCvRXeTI0ltgrmUXqASVbbk/6RTgzfKf9o
wXr5eaO/7otnkR7J5AV/cPXlQ7XX71rmU7nTYv1vnMAFPTcN+5RjPqacp/5hQsmsPV5+s1VI69Bb
XkSQMe5+Fe8JtGZGcjJ3ra3nGEeiNyplxpUxFu3nuA7oET5ECu2xfTjAI4tqX1qVtP6RSZtomEVw
/moa5neMIgd3HZ2P7AnxSk3k5/BlZoetd8fElZBWcHF26dwCbG+7gbUU79NH0oqyjU+c9jQfLQGQ
Z6W9n04mhoa3rxNseaz35MLPYq4rAUtsCYYfCBlPpfWLQd50bIUrKgV67Vi2J9pjq5M3/YHRateI
Wj7hJSBi3rWS7Zve6xqZVdJLTU8tVJYdS1ErxV2oKVGJQt/a7s1v73K29bF4LhQb6u62OjyTYo1A
8eXBbPXFO8IKPlZtXv1y5yc+K//DpqyBUMmPr10qJK69JqZxn4MWo63yFeViMJ2wBRqNKZLbifi0
PRXSLeyn4hng96IQOYwtywLHh6jnWhC2T3pt7CZMyXwNzgDoSTKvi3kKhUKr4Hg/N8+gD1qxGL5D
YjzyUiYgMbYwvIQFFjIyJgFT+veY7CSJ3yDGAZhpoQiH0fKCJ3O2iHmTe1YWP6edDHYQvPKphCKj
JvgOtEpKDdA3jnZ9d7pVEVLHjSH+V0xYaS2c9ZCAo0Jc7O/tjheCHc2T7gO629X2sjO5z/wRB9Vy
RzmHRVUFcSExKlKpybTk1lzDFIxiLO+mnXJhAln4R9vW+8Pe0FNAJfWlRayQTqte5HnpOaWMLP6S
/ORIEfTjwJMUyNjDsELDuQrIH/zZ8+9fK9dF8QKGpi8WLu+ddkUfh0hU+aizrNzcBYlRW0Nu3uuG
M4k6JLVq5rnl9wnMW5TPZ+dnjQdU87KcB8eB2a5HXND0sJq54XX/iNzkmIpwCYvwf+QnWkPSBaaM
Eo+Y7qmoP7b80Qk9LCspVKFMVctiM1EFIlUxc0Lq/Mgr2sODIRzDPnpLpikQwx3tRkca45s7RjCr
5Yq7tLQnukT4DAr24OAbUxEA7nbdsiqL2TNozzstNAviS1j0LAJL1udZasBB7nxIh6TSEEjXkn62
EQbi31crdM9a0X8YSCtCLDY2j28K7HZDldtxp2lRy1B3JDqH8IFUAGOd8+esPWAbkK2FpNwqN8d4
WUk1eRVDBt3JEuzw01XQR+mMw6wpErWGfV9O2jFWAEhn0eznEU14WZPFJxt8QN9OCgr/wT/iX7vs
QEO0jVKMm7JG2vtDAtJc2DOhMpAHh4s14V2Y/wzIaK0TkRC/vT1HfGSuf0NlJCYX2Kt9tXVkU3lw
ZlQ5QwNqlRyB4SUSAuuEoutvXbYZgx3yviq4vy8N0GkcwBIoioKdcFmtpkEBkAyGpJvoy9gHU5rR
slxpe+2QsvN0fGeZVjV9ly//mDdwS5oJvvnj19bHZalfuSxrRBQAej5ifBE4dZyHYU+AoVkMdqhj
opnTejTi2Zn5IGKWdtZUOF9TI3gPTXpb5jcZTeYxWXctbCVXJGEwMyHDnm7xRuMPdvmYwtPF9esL
QtuuxTupmX7eL4mRczyYJvXXlMo8dfz25Q2xdpgp+uuyFBpcPHNct7j1P2CezF3te2k6WEv8RfNX
geI8Slp90hsyko+SWXSimInT0h6bdPSTyzQ0sdwevvPX5iyGQjX9UufopJyQIoiY7dyOviQnvCZj
WjuSuwj1AvVFOcTF/Nv5lptnCxbHHCviSCKgINEbywZHCgkViSxG0r9YMQjw7cVdKfGrhVAc6ZKw
OKSRMNISkXuA/1Uq/DY93AlK2x+TyVXek3hxG1sn159h9UXkKIwB31e4QieJJQrupwZRk24J+EXh
L+KdTli3z/tX366doOOYD+6pvAxNsX1Ukt6TC2RqX+5ujWIA4vDfekQpE+4hBTAHWSlBxQjxQURE
XP+FNDPaH/tNGwyq6PzrMt9YskV/pG7qhxoBmEab5WrZPj6bSrnRfJZTzcxGCw5z5fIx07lJTSzQ
tyFYRDE8SlWw6XTLfCNlGnRQBPzH6ICvWDHTcb/YXbn6jROhueuwSrrvWeB8PHCInA68ntKvY2Zr
uC/ERpg54fnjYkNNPE9NjMIZ5KLHgn53suIggQ8vSLL3M9J8IINnOpbAPDvvNm9oSa91BEpnRir9
IMEjSOhUmtfGNFq2BggnSGEJqh66AbN3xGePkwdxkYpU3wWBzqcEivAyBjvcMEhAynQNCWUMXEjz
6fqC2TTBANTngY3sXRZ5vfOLFExG1hJxXv6FaBmfWaiLQXf5OITATo++DcaVyl32BCPJa+veg8es
kSj2XgWmc5RZu+y8S/SZ5fEamarqNOmUINy4K8swrmn65KYPe0PdmsbX753ON6UcnrRCrNjs84WJ
YgRMJgk5R2V/8Kb6+d9JcJaklFuQF7Eh5bB2CcnqV6WMivU+wF1K0XL7d08hPFir5Gq0qKd2ZSMA
7saUR4PScmPCyk5UZRsasqbmrtRcGueZT5Fsl85yZIEqj00CSmHrYAckgpeC9FuLyCSrPvQr8uKY
ylT6ri5WEDGMgvQEPEHENvM2LA+CPyAcqIWkuZx2ELGqiAfXZQPFLhe/iXrDmIhEFXDHs71I28Uk
BoaPA7+f+nD32vaf8eb6MirNzSbLVjyon1DkJof/Wk7yQUepEZe5JGrhzq29/OQRmnh1I5WkwGVB
JE7ANEt13b0AOKqMjfWiwyVhcvTNq6ftYkKUpQ+jF0dV8rEQOudjFddHC6DldecnyyFmy+vM/B7l
qRspnaFIJIBAgzJZ01vcGAEMIBvswcgSvo66rFi5jnJnQdmF3+vsVjN/XP7BMuJwdKab/slNHAa3
bj2oHhtcryelrZMTLIBL9GCeLToGfoZCCIlzUxQCyFL0s92gdLuPiSSLAi7++JQ0uBTqqb8VWStO
Jc5LCvqI561qPYjDg9F9PVxWKQ4+T3RVl/+nF23BAJhZuWVNVp5zvNFXXPP28Y9vhl70l7S2viAs
kD44RqFMAI7t3HeXaKPtm2rli5BYD52uzK7mkl27pN4yJHxdm4CAFDlNqpIfAPXHPQGgjh78APFF
3THk+navagj+6hWXT4fhRV+UevZCaxaRS7JSIR6wC93bnvOxNIPmRtkuYwSks3yeRSGR1rUqPvLB
skA4whQZxz8L24gL+6eaIMZh63tchcxNMZ7AJVe4TRLSc9L68lztulScirBsuNubewxyXKR8osvZ
KvY82elL8BcENYlI4STOZRg24urn81gmxB6kqye6FKvK8TDzxq87psV2IktNmLb6TC6pAjfYBf27
Pk8MWMe9BRMnuqUe2WHWRbsikuiZU5rTi+3npce8hO4oOLxSryP/+dHGeeou3QUYRHtuvfnutZBg
PnsCr39Sesb/+SaT/tc3grdQcUwnbvQcbwktDHPIHUrx6xmPRmtu1Sl4PR2AsuoOmet4urS1UzSO
7LPS4B5KKK9lrE4nrABi2GoRVU6XXi5RIzGEa6UReMWEtumtvJjsf3PehvwKfVcvuZsxRDbOtCAq
6rGiwqfYKqU2gJNqVId3Rk6nSdGdIx16RAzEn74Ue32ihvPlFk884aLLccWAEbzxoKiBShDLqF1c
A03dpGnzk0qKRGdgAv42VIwRwZk/IuG8CXMN0wT7RYpTm/xwvSyD15t66co435HuA5tAMBmAHYxa
xcpBjeKDwTUMsuBJ/UXkzRsM/vp4XfQyaJHk42+cB0SHWkYcYudgfkWWW/OkGv/qAk0n7RxlRiEh
6N27Fu3Gb88JXvKbop1eCL5j4iVprXFurJk+aeu3ygyER5G1GZEgzjKPfQ1CjgJbBiPQEuAcsPJW
cMJOKa5Nb90xn3tKM0SvJJ+O6y3BV2IB9aqw0hPCDOnhPlIXu5YnYrubsASBxUGGPYnKwopz1CeX
hOpbQVIl1RaMP+XsnxKx8eZ18I8JxCpBCW/0+avOdIpvbTJqEvJjP07cHn+yXo/OAS1LYbqh9Ngv
CwC02f5Jl3VkwgkraIdpiiIjHB9K5a6T4sCCzMoakxaC3RTIzInnyzSLel0HxboAuCRtmdRbUepp
kE5t95l4t+8Tf0S6P8SL9cCVQ28FVhPbg10xIyfUEr3d87nXr9/CJFBxEMyygHVLzmV2MdRTncPB
4cbCCRj5CdFSA7m0zJ/3AJv6uFvTmJGnv4CaAd/CoaonQIVW3UqChTpeaRgJlRcPz4gegnq/DNAm
eQiXqCE4XO6oWlxGRP5oHXPUj0AfbSNQhXaTAmVypeeWM1ulBMcCGAmFIhpIbxnDC43agUyUuO7G
O0SMqzmB0dtPGqhmXbK4qEQub/fU5OGVVGBef6xJfzRXl13vXwsSuiyKHL+xW19Cfd1ljuR5fmq9
a7EvW17XDOxD53hEqaeFqS61o/+2f0W8Mli8Ae1bb/TtCRDsmeFJhAncVCUV2jsuRLJBZSEmNurd
UlprEKC81A5nboOYIbe7F1hnS6NGUw+GD006OpNR9EQGwta9znj9g2yTEWgayuvmQ+ZW051NPHsC
GK0BAxGunFtZZxQG1R3KfWivxbHr1dYi3MnTSzQgaTxbEkTgHWn5Ot86ynF193WZZ1+AF1w8qLXM
/Kxq3sCeQSqcOH7LN0tly+ikgGHuAgV8TB/6U25RRlNbGC+sQLQcvEf6s3zsKYiOPGAb6dnec1mr
3YeA78LA4TS95rcItFYQ+ToCODALY2aIts9vTJwN56FQxAzqYhiYY1uWPXCvPAsb//PE03sGlfto
YBJq2vo1cVYl+MHx6BzzSxKsAKNFVM1yijlhYXcNPtaGxXh0q3JWu3IdIdx1H5iGMn/GHYTvGDSv
ppixz0IC5b+fg6tE9dzRisUkW8/BgVTarm20UUcj2O+X11JS3Dh5KC8863cB1cVD0OTFZPIVuYuT
GYfvNODI6bk1q1RG+9LIyPTeJFf8xPmpF9Yg3EfRw9gTx3IoFDtX8u2YFJzRXYhU994ijA1867uQ
+L1LAf/rEW3hiX1S5G5xos1HZG7qW/AWda34DEoK9R/Xa9Q70WkFjWSSvCc/VDSArJuxjWXanEjt
D0w3wfV9qSKakzbfpu3LMbnqB+jzK6qOuPKsoPGUZsLIlOBbd+PK7+1TFezpunOk+NXaMMTJKktb
Mls0SThxpPK1cRGFUrpMnkY8Mmg/cs+98mA7RolqFlAXqQxcIoVNDfRzY3Te338oZpVQcGHHTTf9
FgckaRmjNjqMrq4IA8+ukjGfwsJ7eFHF0s7xULO50hof6t36fsirCY+PddKILqOlxEufwrKG6Lrv
8IoBN6DUvaiXRrRjaoXKIDae4wiZEuU6uyXB3MMiBLIUQc32C7oAjjURjOXc+QXL8Pp40ZvSxZcr
baqVJGicGwjFEfCBCwZqXQVCy4wY09Dy0e24GGOYHcmuFbQGm9H8PemkxXmDHhErv9Kt1r9q5/Hs
tqdBdA+V6yrlsmHoGHsZJ0JYZN+8/IghO2KNEauBvJq4MjHn9zHGRwiY7evWeXHFQbH2oisIStq+
rAeyGKQfdUh+2Kx+CPYYNNsRUQIhyIKIHe0ACBsybtuoxN/cA/aDPE8U2Rp2RGyaTcZcQ1fidnfI
z/7MwLq3hR5VV9awUc78TmB3Ij0/MCUPkmEORMGk3yW5CPA7E2WI8CCOocF1otBlcW99/HzaaRSP
41c34rUSkAu4YEewDfHWyrUsRD/N/JazvIdu58F/wrXSf1aqGSqhk7sO+rVXml3D2WaY4j4jbBhB
/yMt1cEuB2l+vxCAzbhgRcA9LnGGjdNu9NuOR/x13Rn4YVqCKG2TVhUox/KdXdsp0hz4A/y8fBLV
If2NCktqtfdVeYOiU9587t77iKOX/bjDsI94gMoQHjyPavRbV74ia/cGLXTZX9/Nka+Oh77nOsUC
O87RXgcGavZhNuT5TJfrsfDgfjjHSFXE2h5zN1SMdXu4bFp6g6UBt+pe5op/Rzzkkjr3tgl3WV8X
gw6BokALJN783+H/lLBV8TNyKuSBmJt8jhByKUN1cvH6YZ5ol9Nzk/R5/6QewHa4SaaN2ul4V9+Z
aHrrwMgLXt5y0sRFzZhuUGueJu157u4WgkI1poThl27Ql2NpQujY6k3NHjYgOS13O/JesYEgC7pT
d8xb9YtVy+Hal8HP53VqntWOlZEDNydlPIZZrK3UF+BdXGp2BwyE4dYVwhpYb2kXbKiXoQlUIyKU
9PyAcyA9c8cUl+cS2xx6Z8S+Xf53/QKsENaFrx3azab02BVO4ds2Z4xAHUTiUvIiVzo5TxtIwPm3
+ReNIQ1X07d52iyP8wJ01MklaIr947bMu8zy36nGud1EKWJRpN9UKo7SVduGDSUFUN2alSCMpYCf
kfgFtAu7+fduRzo4ErdWNXXTkHH21gCjMahiMGXZCNTfuu329luuhhNmIyL645tdJuMOhVBb0Q1J
K4XasAclrX2dAGSKxQJnOFUS38D2a5hdF+1fi6IFZF/0Hm/nvjA75oHdftISQFQ2x3LbejTNIt/D
Lp9O9ftYd7kfsp8FtrUDGXAjdAzZ/xWHWFBioOCObrwHg4VCO6Oz/Z60NfDYw/ChwpuWZ28/l18i
8OYWb3RHX69W7shLfoD840jo4JoitU4LqttmTIsSqchfSgGfXrpKHAj4if5x5EhF+ilehLll93Cl
saLG9+7Z13VH3Cw+WZiKO3kEhavR3hJPjMpDYHWVIblHYUQGEezYKyZHmeyNgaZALC2CWhlaBZyd
fZCN/Hfmyx2Bqb5XXOdiTA9vNvekaKKZoXR+ICIosc8E4SHTjbkWy//lDpVye5VNMMLciXTp2htH
S2P3M0pa8hth295tJ8fwpIHEEQv3fw1AAF1cIR0x9n4AusSXFEnF/0wGTe3CtpsNSaB8GhrssNJP
4Vm9JabjMgXUPdcEayHVKINCoi7CIhb2K9RD4ruyPbV6QAnhqfEdcFU0xwBmJ2d6pxYDOxc6L8ed
59whbVPHDcv9np/0Tu4Tkd23DAnrTsQIgrVyW/m2pBvzTaH0+/LeLIzWcPZ8DEf7sw6YEVKNfIW2
oClzJYEz1DmPcI9NFRLcIU/bKd+J/Ue/fViW7HH71UBVBwWYrhAiY/4L3WUDiXOlRZe4Gv6LcyLH
+3BODc/dPbQK6a47nWkANGHlOFDlk55spO+MyPsjE/Uyt3w6J6nxCHTEjFsyYXVOfJfJjiX7HRND
ElECZNWQkyqCzbXVqmpaW2dFCxL6qhCnEvuU0anq5f578TNSwKmmBtj6m6U+6HF7/vxTmKzuw4BC
D+xf+qqmdJ6a8Tgz07FSsxFsGIswzhYElUjAvOYhl0Wy4ODovY333dy2NJxJk/TC8AYETiwB4XbT
Fz6MvEOQRoMntied7V9RxcLxJeLtVqoRbo3Guae1jipNBi428Ven/ZoScT/mzeimDI5k5Ta4ZLiN
0wdYUKGTJcuUQ5A4Wh3KD4Z/bBILwxDpMT5okitLXzc+ZaNrcg4kuJDbatoMovu9jShYLQZu1A6+
tGm/ebYtHTaTw3kbeuMph6TdndwifRqym8cK/3lumorT1Pw1XIpKPh/4xFqNulPpteQ2h+cl/OM6
DCvueTwdba5HjZe4yFKO8Pk02HDkW8Q6ceudx5GhxJj6VasoSUYUFwjbnsGzkm4iFAmDkscnywSx
CQGnyHeUGoJEkMmzLltemZQFeG+oowtVyvABczT2QrFgz59NDjnx2Pcs8op9szMNfQUDLocmECJZ
jjkQegCT5ciwANw0Wn0UApk5GHM4q408E2YuYvOyKxlFj8PYbS9EJIbTQbLELxeBIQTMI/vhYoEU
Ta1W3m+BmgtxaQ5smIpqF0bG0tFq0Lmc8jTGyAiRUawtfRybaWOgFVjwzMxu4O3lSOUyekulXfXe
Q2pRjTvlTu7fPu3BKLApsSUFltvDXVuRo/je9BOQ7hnrn3tEMsc8wBWO/KvTxAdxNzsY/bds1uBd
TW339q/RB36DmJWZI7iz8Czf8Yl2j05iBnwzQThR9pSI7BDHcdJg5eLH6Vb/VbKxL0DB8d4DBctj
/KdeTe0Y/0rpPqU40tAqhFpaKBYZ9BKtmae/wPP6uCABzJvqJkzjA/HQ7hsvsV/HEs9hFbxMfH7Y
Zq7jYK+Iwcdupj5qBP9pZR2ApE+NaENsdmTNkRwvTySbMU5/DI5ZaV4UAzwK09SqQs057CsAqLTg
e88V+NPfSxt0LQO22pZaN4fetY8sh7MvC1hV8BehrkNIs4YmvCNz4dWeXZCUxCQ4qk8HfVRyvmZf
1Q19JCEnnd1Yxf0HtOvwxq0xS6GOAvTFwd6hX1SuA94d+dl/C7kOfDfPIqjPyO7kOH5daLyb2YE3
u6BjJJz2/U2jC0LQNx9tPvb3Es1l2YISFZjImXqKxa7n5xjx05evdI81LIWUptECJBKn92Liwjkj
2uIYFBaqQX6edBU7clR9lwVtj0WlsMRifqhdfnZ4+RX/ksxeRpK735C5s5oPLV2QfvOv/hgVGeuF
u4YZdz5+FmMZ+rt1gKc7w/H9qLx5mMtB5clbMTkhJ+sSRo7peNeLTSfw+t0VQBFeDAHV/DWYcyIl
Xv84lAN0Ng10+B3bwkGlyuXtQI+SSSrilUI4vQY8qolsNNiZyVG+RGK79Ja5QDUrbthXE5sYWeIr
3ddPcIlBEaGrWjolRmMzy+DxPEpLlm8Ixx1l1X/e1j0TyoPpJWK3cAXaY65CCpGKbY+Sasv6zTYz
XbC31ebIRYlBNPwijIg6EItvYZwwbDDu+jydjVt3JiCE5zKnyh95wz/4H0/Ye0S2vUi1/RkPecVw
BP8G+SOwwoo6eNi7Wl7owVgYzWyFYDfwfUSq9by0YIOYXRjW+tbB1MEknZhETQyJ0DYyxLIv0tYH
P1MSPPb+GCks7m/THdpV0JXaTfojHiD563+t+CCwSvofZAdSCHOv4VbrME6RUsznaFlfWDsI1woi
tAwtPETL6v3GbQ7zkuU/+IViUWjIFAaGsP4y9R392Gf9IrxTsj9+fHwi8fF8e+QHeXEkpgaLcVaB
ikPnlQJduEgd6kX4vjqFRL4nUsg7mQ4TcWdcrHMnz5/emNafxk8TqMu16+5touIJzgJ4rjbTy+ic
S25tIizWmWvLAYnOJ3lbW79CUZsa/2xYq5AbtDQPTKbdRJN9/jNo5AkdF/Bb5Gm3Qc663qQqiDOH
dhHVMMFmsfrwGWIRT1iKnXs+PwofapY3lpZDHXQafMuo35/zOmfu+cSiwVY3JzRNVeXmS8fF16Sf
I0PGZkXLLGXD9gQcaxBo2lG0ZsbtiX8sLmZ0/QJs/55VeyU/M5i91FVFqSqMNO21AM1uqN6RMvFl
UOQq4/usblYOAf84oZ8lNSHpmYRmvqDVq/KgKc3iWpoYOqzT3xk7HqGbqlcIZGcEtjADMGHMfTAZ
B5VnDFxI3P9Vxly5s+mW4Q4fHYUioDZNFn0Or7JU18AJ97CxFUz+tcx8iaEpM1+JmT0O0qfEqrB9
wCe7OLG1NM3h8W/omBwcevMxecl4qkVe3UUYdV52obj26y0Z8FjssfXpOr0kRVVDfw7/012iWIy6
OPCycz31wCelI2eknLOvNjRlua9Xp6VLzaEL1pG8viVn1y89DAOzvUM8y2ZAb3doW/zz6Vc8gWXn
7vFm4KM+5+oL+/Ca5HlsP0r4ya+0Z6Bt8e1E0zCjTPoNGHQc1OXCMndL6JJR5GGdgI7j0v1B7w/3
591h8Tk/MXRl6VRlglEUU3pNmtcV6yEqJ7SevgY/A81z6LP8sQPrGUxzCLnOMsE+J95Q5m+cmw2x
5Now6aAPDajh+Yx5IObcZcenvG5gq7SHEf7tS5UZH8mW+BZ1kK578qB69YGmIIzo2GQ0QfFZlEyO
2MlYoTJZyDxtVqEtRLSON3PHyftC15mNqSn3OcQ69Z8I4rE9Xl4PNvMRMdf8RaicdoTE0H77VI9X
oIysei0o6XpJf49cIwgop/BLM4Tct5ViIfOwKYMKOHsVKe/zMKiak6GLeGxV0NTjHlzwsBcyfFGu
tFCh6uvTHaO08+WG0TpwcvDE0Ab1vuHV44354/cLN+x1ZRhvAOvYT9Vv6ekOjEVh0w93L2W/R+Nq
AqrU1j08HHyo9zQ6Vxyr15HNBeabDAdRzBahcs/RRGXtkBEn42B5ixVTjrYbv1B0bC/9TdyT5e2L
8I0hTrh7zrsjIYDosMCYWgW2QZD2GPgw3Kg7lf0Smc0wbRRnXrNi/5mYaPtejwh/VgolhEFcRZvC
doGK8VLc8QxlRsXa79JzBAAVRPa7Z6vt1/1wHSUSa45mHJankfk34oaB+1G0k8iCTlvL2z+6zxxu
pT6BQHR+/mIxQI6aEafpRA3KsKytont5gdhcQ+CqEt2ak2Gf/Pr01Qwq4KTxAKsD+XlPhm3bzt3/
ShTqF0Q4Tm5k2Eutf8eqs6+Sv0nV0OuA+8MUxPjueQQ7psWeO3ILGOD128LuNHCrjKjR2xvig+8F
Ora10gb8Emqs0enub7QnQtHqtVEI1v55Wwq78n9MsjM6/Yll4q2ZGKtaEjJMKRTpMbLHLn2KNQST
qGJhYTboAZVxE2KNniCRo85OnFNrGx0dSS9iPr81DseuIVqFrDNZHCc0ONWruXfYS+z7/Ul1bzdO
RODIiNNd6xnlAkB+sc/Ph71Iy9C2dNeCf5kJNPsjW8MZb4EC7l42xxMNA/J9tcMaMBb4GaTR+Spp
Q8asmLts8NO0Qn4DxiMQV7wVSaucg7qurNdLVAdLJt1Cytbhh3m5HECvEHNI71sQ9w/dJJ631Pm7
JZmB+PpiDFeWXmVNz3h7DqPk1eAndte6eCP6rR80q4pxR+Fs1rcuy0E4sdP6AEn+ErxOY/GmufO7
2OZj8mVf0OLkr3wohB2sZmfyuCLUPuKBiYwIZvtIHIY9HrNvu5WFfLK3IpAoI6zJb+X3t8uo0NJc
+djlB9Crr1u47XyH7IIi26pZfRAT9XPcSFXAMzWKNF4WxlU+8u96XqrOGfZtTCiHvfszZHeFO9YQ
URKungO7uClOFnj9NmDhLeULpkoCZYqUul3UaM9g0CYIzSc5kLU2e7gHeSTMQ4lmpeBjuKcIvaLr
xPLoL5NoSvcKBSQftjAv41RCsFywHNGhSE12lojem6o3XMvppJ3uj8zp+D+44hCgCTi2cOh+AfWM
c/VYKWCaZ9K5AN6be/V5NfU+LQe5Mpm8zQYR2hja0t6X/lD0/jsQ17fHrcScVpRjljQOsAHY84Vi
fe5q1iDPnOCl4CRTHh3TQQ2w5zdyCtn7ymtKVO/05ehJkkuBujkAI7cM1uvY50c4+SOb4dbvDx1U
DIEqjyNlWAcKRckdmJJrMtEaedYDX+XnpJRO1RAQoF6Ip78oAphQ+z3eDwcoo9RqDoNPuiCeiTl2
YDziq1/gA9Ju89hakYGeMEA4dVbjhd561f70MN2yd4M5bB6AICy3zdtd6FxxcBQns8RMDQ+878AN
Z2Qmt9MsOsEJ6RUcxitxmxsY/9mKEHC58Z37M3yHaTpUC/AqjbXkerw0JfbVSnwBPxExyCt50BDk
di46lVVtLbNUl+YOyJigstPxmGHcpD29GespqNtkaCKZNFWQr+2BB6eJJE0WDBVu+iCjQ0ntFFRg
bRqC3GvcYjFOmKNT5RjTgK7B2vwa9b+OBdU3kgCKjVrNVTSDMDOdBiuv3Ngm8a2DrwnKsJN1N6zL
aJtDTnaWmPxdmkDPbZaudhTxslct5svO6i0SaLi50HtfFDxtuij7AHTNNdvgMiYHel+ljZYxSHBU
bPBdbFoOPfDj68dGE4cZT7sI6DQxPnvrOOgRBnnr+2rtwHDWchTa0a2jABgD/tf4FUQHi3I4w5tP
JVFTEhRXMVPLwdYMynjoEPJ5GSmH0QCniQdPYyBo1IRCBd7tNOyl/lyz3F8ibMpCpZRWDaiPL40y
S3Q1fu8axbdiXH8aGG7GBKx47nrw5jgdKNjU42I3JeajLtmmrVuwCw0We+qwa7N2KXXUO6wkehru
vZDJ9IBQauvQfkxbDySbVFnnkVb7h+Xp8HU3yAsZbmqzhvobqhbL13x/WrrKU3WwY77Qu9wEkojz
DNI6pkzZUYr8se4GexST+kGOv8Sqw7wCm18MPfiLx9kOaO6tvhkaiGRlQVsSD5qCRW+XEFGoBwMB
BZOgaXzXu8m9drMEa4zRFdpFtU/KR6P5SG0/cKQbaRiOJpeuknpnO8//vTkJbSY5DRU2jaB8FCix
nQGTqLp7jPujrdlgL1eAdCI2lihRsiLYnXeiL5Epis4NDt6uS8x0azPgexWmMLRQNSYlqDMZyFfn
IZSMTblKSl4ZnqBoDGEAZPRQRMfpM/IZoyvpkAX/Q/e86Sl4y49OmZgHtm3of2ouby4Y0ABNxU4W
oxQeTX22dT98VynUBIfD+/kzxYeWXxcPnuFQ+yzxf261Dy5dFEQy16yDmqYNA7DS/YYl8Tab5EjG
HoPrqXku0Ukth9E09H4qVLxc88MPXlC17pjXgJ0XdZ3zIHUag+1jIXo0v55FLpNY39aRwGabNCFl
xLafxypKgWtujmt5QrFjawBjYL75xvXdxs7MlfRQFm1qAt1oLuANVYWX6Eq1X/efvvBdshEuAS70
4R38gao2qS06n4JL5MO8FN6HxQXCM5mkZlVREyDlh2DuPb/odOC2lI1JMgYQZZGzsTY7AVYNawV9
ip/cy7u9fOHPLyYlo5yNaBz7WGUU66cUoNS0LW+OzWQKQjmyHWt/jDGUw9NWFfti/IzwwXZD1RVT
APsUd0cWgoBCE/g4norXs9b7yNJnso/PG4QQxR5r9tCYhrfC7SRg5WmHKjbA8w9hhV7z1oFxnKCv
7f7FXiCOmw3Z4R1bdgZheeasHy4jLsrYGdiiRMzOhq2xErOc1ZRno2EUyPqqhaQCBKcqcSw5TQYc
WLg3BdbuxfBj4l3DbpuZ4WUCtoECtrMiq1QGcMaHINma9pdt2wNLAHBF3xGHcoejgSSYgcF4YE39
hATcU0c+qynkF7nwkwMD+7swQoUhQW3rFt2Tm/fhL7RK88K4+71dtwmqRAUKeise2F7wzH+KjDKb
ViJeQFy51fbGpi/0sIK0ologge4AhQ0QgL8zTZvtdtHlIMIJ3fpYFsacLqNZC1BssWgKpmny57U2
VoE51mansJ2+NW3XdjzbuoUlhaljJIk8a+GWTr9PlEPKlhOZqfKyeb/moXFmwJWPJHGLTTKzkt6k
SdWmArp18AqKYjNLmIOWI0PNKarIfbaNCq1r22q8C3AGVvasZignz5bltsDD1bIO7ZxjYtamEi/n
2xKLvMBOjhksjOR1P/uXbYGxYjIEUdKPPuwj7XD4TglloqQHB/SmENQRmm3Al05SW+Xh0j43/hwF
ytfvO0/F1yClrWrA48Vy0uoqF6FtCXQXXlbAL5M/SnnBcd0RpCnDVoe9ET8eiv1SP6UCctEe4uhC
34Y0tq27fwiVVDmTo/T+80UPT0mmqis45p74nfn9n6DsgG/Rb8EzPFAlLj9mdTAnXNoXBcBxQhVH
SQvwV3kkSzR1hDAn/A1g/5zn/JpENC6tODPvYSW+tl0sjbiXq6bZSr/Uq3GyIlfgsUwJhiAxNz2g
/3gdOe2BexQIt2hsyNnhMRscJHk8y1/1rOQYUPwMovRfxPtiHpwdxzAg/TJgBu+Q3YTLw0xEH/l8
ocEf+g9eSeTXOW/Wk4bxmqbX96BoAJ46y7AvtNaLKmWqrq0tD5JPDeUU2BzXq5MGDKoU+uArdXL4
RBeXS65p3bcHGTjPLGW8blq43R0Rrn6olXb5j0mJ42QaeUVNNYJimWpC1TuX4wlweFKs3bVLVKkN
R2S9IV9zll6ii4jHEIS7hJToVGzPoKTYdFbwfBSaFhMat1ZbT/9cPtl8KAJqHsvPvdodp3u3VcFB
Bly/jwHZvo+KZztGXISd32ujQpY/JXgO1FMWAK3s4R+Urwi9jeXEb2OEsAsGwsAAmlmlfUvMDAFQ
xePamYyoFrrWLWbXLdRWuefex/MTHgL2e0VpvCEeAazSaWX3X52EJoTwrvWSPwa4qF2pF9k+ZF3H
oEuC5DGIA+gZxjLRJYJjFbxpgg2XcwVAVNEFGj/A6T/YjxNtjDocIZRhuk6nRYWbsz3VTeDqv3yl
b+i0AhCckTAv5tQqyBMkDtLrGYmw9Z1ARuGEv8BtL4y7R2JPwnA8pUrYoQyOQPIiGXx27At5yfXY
I8DRM9zqv4FEkIeoZV127MvblJUcRlsmysT5Si7Mvyzh4Dw8ZAO3UhNAvQcOHK7T2/tGF/MCMnRl
ueTbufGs+z4wI9zwps5//VFChv5tCYO6HpnFdUVbjT3n4KJ6ZkhS27sCoSAk9Z0yYIA6RaOSsS9x
4dmaeG34eJBb9HthpIfKTyj+sfdqF2Qqt1KrRcBHpLLnQZ63F52LoE1zm+LFJ1PUgZI+a3BFumYM
7PF95YjbBQXOtIoKV4loykyk4zcs2dKKWsvSHcl1lRoUDIJLioVVqXkt8G68Zzjfm99AcsN66UKK
ka46fUCWO32ZCvfLIcR7E6Eha7tfUU1gKPl5vNCukqbWCUflqaRVpsF3qEWD+DxoW+xUNM3BQBo3
6RgyfKp3yXHSdUnyQCWMcBtu8ckZARMDU6J9IMm3JEBtlt+HU+JSOYbJxU9/R5IaH3WtXMNeJ9IA
wk0c9e9bmRGP3EIAt//qs9Du0dOtIR0uRLW3lT0T0KefVJq2Y9K8KlZkraQFKgfpU6mUU+sa7o0f
DX6eXpBOJYbwu8/eaysNBISVfbrcVHCT2WeX5vbtWKJl0cPhnFW7cXY7dBVCgZkRydvWWKGjzn4z
+R8XuIaSRDo14nxsn9Tk1ZSFxHsYs+n0R92Sum5QZA1QT5b49BZRNo59GWOGehFJ+yP5wC9I6hLJ
5ayYjR8lBsN7o33f23HAaA2kLiZzI0fiPXV1cNGF5HEpbb51btvha20w9KpxDezVzYJcK18PI9aq
5WVcSExL1QPIQyPLJnrpYEKNUFq1OEZYcLPZ3L53pRcD222hgP88Mti1fXAvqTvViGvcvMnhKEU2
C+2k6HR4BxElCZT7I7D7J9vVx1zP9CxbmkTTh37Cs/eBV1EZMcHWgXEFBWd6ZExUkhBHC+C8Z9Kj
wOBZomzc25GX8vD4T+E16SE+CEiw73yUwXby60KTezCAt24jbK64rM0axwUbZlpeIAiJ8aERHQ4x
a5KISgnPlx3+Y7cxEdgAZ/UrATuNzljb/9bZUxPgJ/g/9Xzu9qpjqf5j+dEyLgP+poV6x0NpksfZ
PvZzA07nTV6ukqcB6UCiYLPulng3MPSrfhnf7JCQFxZBiz9JhF2nl2xF9A3gGSydu6eS727wUNiU
6BTk7F2jYXyFzvIJa/rMhCiWIU6ujZVF+QjMM1WXstkeF/qN7Rv22wZXj4GSUIARv1YOH3TFsh/0
zX+k26MDiXZZkwlFYZMDFf8I5FG/6Lgx8RayU7mUe7w8rx7byPGEYm/s8ZVwfGN36gJXScbtNEcI
IonZ2YE38oABwcC21KDp29E2PLx6bJ17VrlZXM3st4UW2b0dmZG/Lul9z6Ap4Wq3qBPXDHdJ3RuU
qr93dJjTtaNhhySZjGL4tkTj+qdQFk/CZKhTU/qxEY5uBLU3YjdoSRca1snGxhVE6VoxohLpIxJR
UuHhI+OtmpWeUQqpXeJCntFwz+aY9yqklQigEmhLnIijdtM6HrDJz8r3Ll+WyL+OehIqmCV9TvbT
vJYLEQKffm8gRCcuLPPuacPHn8keS3NRLObQg3O8aCU8idgJiYXq8Dr5YqIF5+BDdOMsYmBXa/zk
e2GCWgcZMZE7RWF7MHNTbUf1Xzd16IhB5GpJ4fslREFe1mLGW6P0tychP8KFYQtejtuhlibJ0RNl
l1xMMC5VHOJzJMx5eNIesHupZxnwjDZ9SmluVBFygKYDBbgGEHu2w4UOlpy1hf0I9COw16yrHhfK
I9wv+ytsZVcEsgN4HJIj/SngEVNJ8kLhO+ojYeq3M8X8q0j9nj+yuRiKmR52KnjQUpms8Rwz9Y27
3J4zZYHSAK/vLlDGYtm2DsdLBuH7TSvEX5Fv66awIbEXEkXs596UASS13xgwsIvpZAIP486MJhUw
nKRYxycBy1BLzNXIUCIi4gdtlt19lH7vKLGakIYHgiCWcbQMR4Wv9OsjjEvGI+keji1OyHrt05xi
3aWNmRDgDBL5tLwZQbgLlH3rp3v3Hsokpz5mW49ZCFfhlNEdVNMssh65WyComQ/Uo8LofxYr1KZA
wPxKJZsdiW0a9MBjbjHCNswM0vnkUUhBcFupUkcTa0Ej+KGfZY8TcpJcdr58zsi0BvIb6SEgiJSH
IUm17fx+aK7hj9qLTdVYKdZ87H4IuvYhd0VD0qjGrJSFZQPEtffQV4nqfcAWepXnhRnp5YItX30T
sehiEOQDBaODvzuh7RxXXfPUO/2wjltarxaLHKMVGIHdc8poizx4mtHhboLmn/GVe0InmXCru1Nz
Wi+Gz1Bj2R/MNrUMexa+r51nRokqF+y1YU6hOzCJQQFuoy6VscWw/jiZiwDUQCDQZzO2vIiDTovX
jAvj6NWF63T4Ewcr6M3xqrVpTgwPj32VxBVILy7JuDjQ0TAl4Q0S35WzGf1sjXcisyNNYtiTmUTM
hG98pHqf3Mhdp+HUAZtqYojMyfyjiK8ttxOxUkPhkJm7VKUDIs+JLs9qmsz8SG92WKVDDBAX36/A
/K2q/ZLYeEIyWP/A8qbOoGKTv6z/oP436QDHiQnbWy2CGAU/Y+srsaazgxjb0l/CdPXr2GCGjuPW
6NUpBOz2x7fx4mGzx2quz8avx8Qt50UvQeIYISSVHeWRvN+GUP2bmgq1IDbpi9QmsJOHW5juvxew
nrz/kzZslO5zrYxfPXWBLbKTf5KrpnqVOpbTziyOEPJ4IWyQSDPm6rTxrrmDTs+XFjYjkD58+tEr
lqY0dRMEWupt8iPqu7MjsBlkYfh+Z91/GKYYVThRaUnslCOiRscGLbiuHFFLHqYWjwnVUGQ4o1sR
lf/ShzHh/mzupd2t8V3p+7mx0y4ATQpVB1v+YzOTGwjLNsH3I/vjtyIS3AiEqI6wL07Rs7lCQjAx
gaYq0b6ald0GkR+vSQh+A0qbeYBseVg0pEIdJsw0rrKqOg9k2Ew7JVFWXl3NpxYGKDiC1jAGUBCh
X9+nUSP1FO/IwKtoVgd/NJ4HNe6Uc9O2eGJkr18T1LAq4GaWzAQbWOTG7YT7eaJae/dbREK4yz3l
3OIqrojDiOlyCc5HrMKdwFFmzsrNAW3YMY+e0jVUBBpMPaSKjKGz7v7V93LbgBIuNlCAXRPNe7GK
5X98rslRkvoH9lp/Nl+1Ls14LcoMYF2lkjG7LPMnvyjMEPf4o0T5emfix3O/Szjz1OXtRr5o6CSq
+ukVEWeSyDAUbcAq0L5Lf+1ImxtLxWd9vWGOgmVB/+o7xWWbQrZ/Qmp/YIBjGOyjUFikQUj6yMr+
kxcuXT77iFYuP1zQb8Jg9fnLVnmG0rBpr65bVErtiMRx3HXGjDM9699zGyKISzRQO7/Sf92nUGXm
PKJQwTmmILuV1ApG90msUnU6QTYtusDt5NWZiiYhAycTmb1fnzbZjAEvAOh+O8cKwsiPn6ho7NYh
UdyQaw5276G46xmLymw9PtodRxBIKnCnLXMAw9rLQQM8Mb/ALN9k6mr8xujnwodhQYB9gt0MXQTJ
OcykEHiGgSKCOkTHbxAREOYYhpyBC5GN9CaanNQwrtjbDwIhrS4lEC47r9zb/3pPDJay55H1tOVa
ypWvi1i5REs6sUXqiTuZt5QC5pBFC36vA0BQLyecGZbCVrOYxIULQeXEkwviJZTVaXlzwDrkEKv9
9IViWTnWNKy/ktBc4xathNWF4ZZv/on/R0dpmILRk58V+yE4rnuVooAW5QT9ks0q3+wqbFrGYXEe
8QCm4gqW/3yROEr1QY5zjEYm+FUblo2NHW3DwF138m9FWUrbgBMbas0yvc7g+L83Kk6mfm/De4dG
gDPikOFjSHONpKRi0wpPvfirQN+TvhAq1Mku+jQ/ii0hodoyVAH5xjDqtaesjTjm25Z3Kj7oYqh0
ro5xlry2sq19u2fRC+YmLUEON/WzAD9Yo0x+sKNXQ9motix4NrGa3IUlOwMOHKAIG/gXJCLmh5r6
K6ZTsAnLCjB8CUH+697P0D+xjlQWZe+/XQ/QrmTbnPAQ+IZ1IpqFuRxUVW6XlKH0E6DgudCKoET+
tC1NkxlSkOmP9LiVYH5dp3HxsmVsyxlRn5BB9+S7sgt3Sc9veCxJe1/6S4bWaY04V4HJFUu7fxXm
tBPf2suMfQau8w5hX5kGhZXPD59kMU5TOh0SV2yZgitz9KZX6il8WIY1TeHJFrCdz76hOQXxwpPi
3G8/Clzta94+xeOIsXuGP9wwi4y1UMw9rBmoSLfNQ9HVFJsN2FOCbcaMao2dHFSMz8se07+7rFbC
eVJ/3Vi1PRRO+y3PBo9JTG3n2AVGf1H9CKHVVDEaNV33KEBGsWu+Rt44JE3W057JyUsnSzqi4W6g
KpVNEcUSpusQZrCZ8BLsq8ChA4pns6I7mpCNDFWnob68kGxoJpM6pTo/HrWZsD0FcKWrnXcvo6Oz
TIVOjVm37aB/1HrSmGzBOPzgut4Wx1+tFtupy/AdMyI2DA9WO8cDVzzAeCyG3UehcwbbxH2NcJCr
lENEnkSU6//nYMEdmjg6/BovUzexWnjmzx5NXUkuUZyTFW9ABbKsWyakMcL1uMmx62+3bb6iUKvH
MGLsXeDS2ai6ZWByHL79b1nR5xizupNTU6pvicDq3PBcimaOg2CdTLzT+1RgOes95hkS2VxYEpPf
DE49lSNa+csveIx1xCaVHneYaNrFBAMv090RXFRxg+JvQ0GfBMjqIvKwJyariO7G1eCfdOHLNL3Y
kOE1Rpr/alCjTHXD6TAR2q+KB+4DLghVLLEZ9BFDUIez6fofi5XboqIKMZFy6JaiEy5S5ddAM6ob
zDE+c6yscbF3fVgrEe65SKrL0/NjQNCiU/sD99GKeatpsBucL75odzshse0HMUseSM6oSnIZtzHv
aHB/HhKDXOJUdePaqDXM3ciFEGk8QNFe6qMOOkRKQmcMscExWd9yEp+xQT++1khInPvREgdBY5kQ
7W2OTu1vU0wbAywMcdputgjACtNLTqJVR2fWjhKpTV5m/x32UfCoRNmRq3IznliM9TqjBIo1stjB
V5S+9dWFwaf6FbCUxYtsYyjUOD+kC56oOgdXBXQc/Y1s+2+uYtk3Ik4KNgLCB7+DcjQ3lA4f3I/O
n0g4IkVp/QPFyD21MMWEbkmUsnbs4VwIO8Cpt45OqN3r1OYNi35VBLSyeH5coPGggf0+vrR1cBfZ
UB94VFspg+bZ1hORrx1dgC3s9NKBc6jBCGQvjrV7UGo90keIWj8dXTYcrQpFnAa78xIS5UAd2GQe
uxT2WWrgVCWFpN37QKFwTLFX3vM/q4W1LC0olRAVAWlkyTLN/+NgFkvGXiRYMolH2YQsynLn38v4
B7UtTOG6ZD6wOmgrbVf/xpS/j3f0LBvoL7/7ofBCgp0NQTn3ZZ3mIvan24HkPrhaga3jn+N0a54z
qhmWuB8piqOMWxe7ZQcCEWC2QGKthiThIqP+MryRVWj4eiHiMPARikIXSQ5XAp9fLDUJAusww0WB
Xc5K94ECu7NQLlYfRguf7M7TyUjGFMPL186ZsA1ysFlYooH9EUFSNxGtkr0JDFe1YZm5N42fu3lz
rGVyGn5syoLom1lMqxPHWwo/MqX2iODns303TLxuQGaSaNgzJnM4Y7ISuiYdl1r5nLBxNMmcLCTl
U2G5ZTKpHXWZD4FHX42H2AdZDovGOWUDwPfWp6DsHeBa/UQW7zm0P5W6vz1LnV+o/sQhv9PYme9V
34Tj3hjv6XF6Du9p1pEx8iIcX810lPPSBWjOQQC1CCKD8PZbhJBQ2TayG4jby0Q/+CUjs634r78r
9lI+UGqAXE5Bt97q3adAlrlKzqzEFfPRB7S549GEQEFMd1yLagT4UQKLpq+hvbDVr+0pEOkiB4vM
rvmm/LKz05lOW4SJlFZr1om2bdXRDBi8YpDGzOHmsxWnqZld/yx1DwpLnT+6iZZtrBfnlBukAKP9
VFNFEGEWNI2F/JVCl5p1zLcRfzit+awBjrpZ1P03Pe3Atvi9M7/31JfuoGUzOVGUTgZJxD6HR6We
hc0MgzMujTWhRcg46FSkkHdeIbxFeLem35GqgZZSoUOZlSQmx672NVMxxLrjU1Bzz5gXJHK+ZtRP
E9UlVfi36kCnqgkIz57jFja5qEjcKf+//23ny8Pj2FPs3aBoQvi4QA4P/yw3fTnKCh+v08xrj35T
ZNmhxFoIbT6PkB+ZYLz52EfbTWePx+mpTx2mjSQt+7hxZGFpFJLXbqCzXfylwsLR3W8Ehpq/NfgT
zycvtdHTBHIK8H/OCNfaedWhJRxyIhAUgPkd4mvv7kZUW0QEKW+LzE+WLB8HuiBHzgCAy8d2PfWn
uUfBb/uBjzcmgUAwyQHEXoHrz+k0B04Dn1K48GimVArVwt0XD8WFPnhxv/ZNL/YBqjL6zBgSBwsQ
rZ+n83VO+C0MMDYYWu2L+MadLVIVbyzUZgqJbNYuWkRDAiMv/gQ4zIB6kqZYTGelJd8sxGgH/3Tk
3/hMpFbwPBjz9Befamgv9Q/czW0GvmU5Peix4j9BLKXd+v6H4aZfdkI3Okd+R33bTLWB/f6UFXKq
/Ew4EyFDG6+qhPDRiaOVOsJdcG28brUTOlz5WOPPjC4j9BVDtbUOxQOeIsksQBY59ry0EoKQ4bbD
l1aM3T2ajgXLeBONt0wCBmavrF/O7o9S9Jp73IgdAUcbZ5Lky1YctN30tpumeZuYt/hXChg72WAv
Aq8vcMpkkiLInZnLmZ0Y4F5EWpfZL7sWJz32CPUwxuNq0i1KRDJ9xNguso8tfSdvB1tBwXTXYYCW
hPyx8JjJT+XAAO0gu+1lS3r4J9Es39F2sMdN+mGVcI8OIfUTQmXxjua1RAXipDZaXhnVQ9GcUpUc
7YzvUEa4mJcryRAogM82wWMTtr1SDeKqwByMX9/Lo50hI/YPl8q8QRi1j/ZNfRxe5Eayw+Q7Km42
wZEj9uuiV+SRlO1Wi2ejee0pMGHK4LGDHJZBms/6Wuqb1DWiaAYDcMJf7Lc6Iw306DMNcfe5IXil
ovtPPdlHHRjJyGPofFapEhMk6W+VwWysRIaZ50+e+io6I/H0EzrT3zWHZFhqDN9nwthN3Uu1hWUq
a4sHDrs7ld0hbRSd5/mUexhVUaV2LaRD/m8N8sQG56WTPTjBUjrR8yfgDjPfUbTZ3k6RoNenjBLW
qwxc8rpJMvGs1KO0f9QmevLgEfm2WCM+xuXz1RQa34v9z+6UQQGKu06UK1MvIKCEyaQO/G2zpKkS
wUZQLcw0wVCSzs2BO5HQ743T8Z7Rd0Cs0SJMTTooV6VAL/RZ7sptjesezjvaznGFCILys5ILqplE
44DdQItChenZ5m7hWM52JmdkSVnGnSCATeUPixIH64edQmemjFys09ZyluGbfbycOBpSzJuvYiJe
NZm05V7iYEj8qxxk/FabHFO+wdzd34Gw6Sggn2DwxS1rY3GVC6V7a80rqUD4OAB58jOtnygaaS5k
b7l9ZhU4pGmSrcrRvMx8JQRWl5sxO4aIPwgM5BT5Udi1nYRm9yJcVskJybaWqEDvY4wyKRGhbJvq
msuEHqdxEqsdCwB2IEahOMZhCAh6Md3MOgkw9USsPwSnMD3EwLfqFZsf/aTL+DiC6e3aItgd0F1M
SEKIIMB51KZKxonIEmrcXNs/S2Z2NWAuNVejbJvTQl10M8FYU1MoPLG6GE78TfmcMGRK/1WC5KkQ
USkFoWUUjMe1Yb1q+dxfL3SytO7uQ+gs/0cu8zP7+B6Nz4WbX32g0G3dYYUj3SjuOOb/C2/huwzK
lerECDKA0q77DxPq9YZd4C/AHbEXVmoUTE51KEUKhGy4inV56yd9IY1e47UKU2ImMutm3A2iqpmR
RL4y8BfffDOY+jYPM0OUFECx2TmEkkGqSnRNKZQUJysRJBknp9QrCrEWjCKG5j+9Mgwu/5CC6Xdy
FpNmS+8RVYcG2eg9Ukms2ED6YE1YOJNg/uKocqSLMP7D16vJN78wHtpacl+quRUkyR14S8Qt3+d/
w2x4rmmrbMrzCGP3GXMr/1yEI7JBba13LB9bkQ5juOTIQVGeFPzozeQcZPEINQ2y6+PDvKOQn3m7
IVYuu0T45e01Fm4j6mhZPomHYQJ/et6HhJPrBXESeJVkOnVx7RD5R98jycqFhuclQ6OBVpisv+nf
0Gd5/YaEbe9jFauavOpoXuooJIoda3+ZZiZhDb9pcLoNEjYjKChrCs1/al7E4QgkgAcIShIHDZ1D
mH3JhMgB2VmQk3ezkGKau5kGcKUoXtlZ3PBm4khkYTWGdlq2JxmubFIGKeai4K2zfXNEiFqJETt7
vbN8C2n8uKzpNSQ28aunisgAnCJAxg1U5mKN5i1ZvOwYodVGv5sKa7mVeqaRGU3r6myS7UKudoer
yJKWBUnr9Y7B9USwswCRAEQzOPl2AsmitthoMjjk5Upjp9zaYyMUF7XZy+frGsCPMca7Yl9HWp8s
H16s8svNbwgbhK9hntJ+maIKdoWG79krf85v5eEnmpT70NPM80i7zM1yVIxwHdxEXIMjMkUKJ1aH
5DjVAcE+6WZ7MvFet3c97IZa9RDWLS0yfznU8VcR3Kupm6/lGrfUpXI8UZvGUwmVInE8k0f/AVy5
mR6VC8Rv5xBpyme7CgmNTLN5fbM7MJjfoCzz7G2VZ6BuVwbuUGtDSemZc87c1hO+pt1/xbf121WD
tccf0YQqkXhVUdzJurhcAIHUrLujw4CaeCEHslXi2gfr/3Mwf4V38nh23KBByYZhFVKsiVzbUcF4
5HeUUW4QVihHKfHhZ6TQFclri8PjSSHN68++ceDm9rnfYJtP/RCrVglslDS9usLjBIZQaKhjncQy
vsFjKEVMAekTiIMJd8vzGujMvo9LPlGh6IBpyBXx7AfeaSocAbyGX9zT1b7oIMIftr07zX5Z1RgG
c93FlKZlJTG3s7lUoDSWvz8rPO+05pFjMRYo7hCc+/JknqM4oH/LBUtVQR70/Ep9o43jiMITzib9
Ta+JbhY4//iHzRyTC3m/V5GRRw3jXoXuGLdIKBm2QyAUCjUGL6oeCEu7X9ynxNI9XU7cG7YtECxe
6sTzeiJqN+xrU6aQcin8Qfdf+DXiYX60BwQJDE8X45m0W0s+2NUpOsqItizXbff/0EBX1evMymx6
D8ZbhXKJP7IPmBbqoTAlRXRD6D1BulX+Yj3sxkmVA2bJdCEOe6Nsie3cvU/kiISG3LxsdJKfiVZY
qFZMoQgl/h3xetjISEY8ukhQjGK04P9xrkDot2C5CMdHFWP+v3T7AXGu0itlOpVd2axlXPCM1Rp7
67AkAWrCvO1QQkYmbrP5HGvjpwy16g6Kd2CP/AvbGsw+OHM1ow5a6PkIk7T9bnUzyT6CIY48ReBN
mL4dY4qtNPfj5G2J6LrYuo2iFrxKlTVh0yVIijyjPaTNMoR34LX8wJ7EfcvPV289S5sLVfkSs7pe
yQuorVSDHTylF9llDanacVHCYo08sef+U/FXG/ZEOfLm07KNdqeuG0mFAwn3Pxncfa/k5xorLN5q
+Tl7UzIl1YIkirlf6U2O7i+/NV8HFDI1z1bLudFVHgRu2aWx3N+irH6Fz/6o+jHT8oOQMrKtREtV
a4QIfcuc8kQztjB3G6UhFBYCLUdZO+ASeQZyKJ0BhERq+qOUXimjp6mk4dITp8GJ8rVqJuPtY/uK
PHA2t02eD3RoOltmqkW8qWHOt+u/oarjvhfPw2yyOMXsugezZc4fcIf7LOzCUY/zBv/QKkWMVK/0
dn/1Br78akFX10dHOerQFEJS9stdY1VpoGrpInqnVJMsYi4SCzZIUIZPlNvi63x6qlcUoZI6wlkb
sFmGnBPpxP8B8tCoTf/Ck2AezE9LjOyFRBs3Zwnw0MBtZO8GVQVw7Z+3djUYDBTFtHl19mqHqUsg
wU8VWKN/18gO9tbkWlFTeA6DmV7aIRmOyPXruO/zjqumPT7gzzYQdpZ3wOQM8RutEoT6TbfoYilJ
kwFQBIy6fuE0mLdwlSivPH9pSMa0TGMFo/k83uXYnvTLJ8Ok7DOdIPY0B4YMP/dfLoccHL6cjSip
p9mH0mVse3wlCPSsbo3UMT8S9FsthsWFcbLo12yOIUuGv1G9VX3gWai1suwNOuNtTYCScJNk+Wmp
HaXFXq2sbCmBlIEUT9oNFmHhQL/rzE4YAIN1fJRRHFSrAWZXNqdw0zD6cRaz+NWN3/PEpSwZ8jls
ZOmDoZrRWyqdwAR4oBw7rl8BPhOik2Pj+kA1DcQHuWfk4vIWT8j+F0agKu/umtsGgvzTGWi9XNca
EeH5CC8Iel18I/xouVN7a2NK3S4VFcxAn1qNC51El/MzleU+JtU1GAH3QVAp5qOkv3/iII/4VM4+
gBOVWElP2yURfsHYRIQZzZPSUa4hOxy51z3hvEal7uatcZX/26lPdgJW6uK00mOskgjJSC7jJYFD
dfElJhXkpU9tmCAILw30kHlCHJt9OaBYDOJ0oTEFnCCrfkXVnxrUsYf0StPaR5wSIYlr+Fm2YzIR
pcShNPPoBChnqeBiNKjwv7ZhZ/Ogy0zZzMUPzkN06AtSaajWe8i0R1uGWFrd+mkZJ//dY9zmBu8h
o+As1ZWmrgsUtyhp0V+25sIUUp8jrdRYZ4scQiLYFRKvECo9J5qk7CNVCSGnDIbR6QO5zJiwc1N3
FZ09dmtQRV1GqwvV+v8RKmGySx8C2PV+HX0ZPFmmYQ61Yk5xBJMHG58orw7MUHSqreorINgnXMaD
ekttRM59hCzB50n2NR86OyJ+lreqRSQuVCYbWeElRoJxOYiwDn2SRuhS4m8G9SeUT/zcS8GeqDCC
fAI+e0pb4Klu3/kaIfms6DVqleLi4jaaEuUOAZXqEN/aJLpooLC/dFnoQwlSL8tJcp2PU2OZGas7
Kz1nsSEv9OeepP5zMuu2mA33s4IKWDKYRQuJpFOGhtS8wIFtxCDZmaE3HZ1IkUfGqOU7Dm04upij
EBotZslsPl8cl+rTbED2or0G6oYNvcaitb8Ly520RVMZuuRM9BatUDUxuaSuaRHvMts/ybAzLo8Q
rmbzJ7IJMIG0HSWH5BAtX4Xv+qvM0ZyYiMJXqELonfaS53fQg/MjFtddNCs5Is5dnn6+Ir0nu+Fr
rYXArr/RtdsgC7gpKy+sv3XYmCE3z4TTDKSbiF5QyD/Rigg+hBB7q9Jn1dUEg/AZBaEdW1U3fNxF
YFWjeiaRvTDlFoGRzfoHgBoES7gzVkfgrzQtn3SiH9Vl2nUHakplybcYZWSzvnY5nX5TSLpw52pW
FKxKvHgovwpyNOOiH14Kn2DI1pOPp++tsO/trtSyQV3sA6PAN+LFThXMdJRmdPp/IUNTrrwa8iq7
Zgec7WUZDAH9ZshSFdBiVjcqFHQeit4jZJKedWU6ecP6eaHoTbyCp/rZRJP5G27caP//DkXD6Emv
1vQzTgFL2elz5g/fPP+oRdjElpDRnTamKH85Qm2FfnjP4JxqUk6Z6OZSbkft1vfA4bUfmAhalrTb
HlzJ78L8uvst0fuCcw7vQ8amPp/XcZYGaO+VE/eIVSimIgjyua6T2xyN1vCOvLYo2e5CBc7W8ejq
6995UcA/H+xUi7Xrn/vw1IaE8r/UA3WabRdZGVP+ZKd2kREPRUYe7yI1Lc49U3z5cRutJmbvr1lY
oD7bdNGIIl2bVqxlKFlHq8hVxwIOzH/EsbaQ3mj/uUPbQX3eTkBpwTNDJXzbdacXnePQpPTv4uZW
U8UeNO+EkQzR9ox2012VdUlrD+AR+r6B+ZD7pdfxbOCu8tqkkr38Vq+nHoJfgP4VsDtZ4riGnTwD
gyM8oIDwTkVAvpH2EsjG3H32C2sbBdVipVqUySBPREAKgBEraPSfeZG2UmlUhzo97/LU67xQb5sC
ZwLZNDLq+A1ckgDq6vOpCKnqIlT2L5f6auy1XagP8vh2z3eX+OnxisZ+s2Aj+Xao7w76QrGNnU8R
WS1NrPCarQQuyCW6Cg6xVh24cITt7rLOavF1P1+HrhoXHIOhaVP2Qrc1+oreArSO4RPpJMBc6X4P
EnO1vpbTfhqy5OfEkrSwlORnMYGbu80Qlpv804sqs+XplZ3KWkWbWGPhEVGvwMuY9dOu6SbkWKcq
OoIjuTza+WGJcmzp7KZ/5VnSCwNc4QStbC0zJn5oJB94JaJ6O8zeMcewBz0b9H+UMn9yvUMO5wYQ
obJewUHDQfXktEhHjkFbOA4MCGMqL3doqafPn5Kf2XhOvnLdqtrHtTwwnhGWNfnHNSBvkND2wGEr
WFA8/GOLpLd5neOxKqYLHPR5Q7EfH6jCmMnGgyodz5TEGzoFFZKKLxHb+8uj0Akw6sEUtLp+tMqN
TUR7d1vw701XdrQAZDc0cydFZvtzzyQ8MUVHQVkXkC4bFIwg/cWkBHeB1n9LqtjBL5zMRZwt0daO
O+JB0Nf7WTkfcEyV6YnSlQU1mYwUlVxBWUMMbyi73ZmseoFXWQpjTOlitpmvP6l9SldG/+odpCos
S++DaC0f8xUBMW8kNuYxIkMdkNx+vfz28A6pcPD5x041VCybJekXlGpta/ByoFcdqN6EVO5jXzIS
8VTFpzd70PxnJo1UAFJNWoqVVa3nZngCK8wq1pv07/wfQ0crWj7BhkCpsaleOg//CxkIXT4rHKIE
/VDWBhyX66uvsi07gE93169lmEA2yITd9OvB5D1PCF3iJKZoq4QTl64mzyn/AvpqQfsmbvn/nWO4
BXbZZIsu/cFyoQI9wW6kdB9N2LkfIES6d38hGIpseCWNt7cbcsjp4zFNUMoNBGFjLEvAZrbGXEkY
cF69gYilKEhmaQkHd4vCsOoeHfdD49f5lIgFU60mc7drGVSC5CL/5IzgVVSEFR2QZQR8YjYdoXNe
u0AnwEZ/0orwma6LtQ3zLCaDmvI9R6bGDkElg8a3lPyCPzS76+AfTvnimfXNMBKrhEjr6M4Rz9mU
ZI5akCOptgKg447j/+7pbDTcKUiNCaywtViGMwQ8S6uCKh6MD2M46AevLBzsnR8ZjI9YP8GNnuGI
KFCkkOgvd8nJ11Wkv7u4ZaJX4w3FYpcITzzpEZvPzpiYQuRv8CuefXoXoT0Pr3/Buk068Zq+avTI
Qt4vX6hqAiklcWRt0VCPG9zCSn53Msbw7W7mO3X6ILAzyyeofcITXbTkaatEMzw5sjCXqCvVUrsh
pTsR+jpEIzLKIGxakw5Z34PyUE0oYPRxXjypdp69Ql+FSIUJgN1vC2EjNgfzJo0rIICHccqbpNv7
KKfuPlbCk0oNig1dnAwJAOInJtY3fYzs9NQHNV/Wp7FY0glc9XFYjCzQM4symW5uz+oLkkIqHn7L
xMvrVtgCnSDwQMNVHGuHwlbH5Je5irS/rspQYCNr8adLIUV20gsBbv+kKU3xvojl33uJMeZgRfQy
4eeqmKkrJo6rG0j/tn16pQeGc0CSmUOQSa+3n/tRfQpy+xjKSlsOKUeykcuDa3PoGvnVz65KBs4G
7gw5bkH5wXTxI2Zmc3gTGK7/FzlsklVUct+kCVMb/JEiY7qiskz43rr0bVIO8yPModj9lEr5FRcm
9PZ3tZZUD6mcOi0tNJZR7gQX44H/mZwoGUQtD+4NbKZ3ggBKiwPToi+t9nSld3CblqIlMbmsje6m
nOEnqKjrjl6UP3N8DgoiuM5xPfuv0roANbZfl0RtDBgwR4/TyGjpAT7aShP3bCg0/KUKX0GU61uE
YwQuVEWO24T2qd/o5+xEYDreh51g3Djxr253+96Mjq157RoR1pAk93XugpemMgJxulm7d3afKovK
W3tCpdjLiHQScQmOOwyOeYdiTTm7qTnd/q+3CmrzfhSMEzQ7iKB1CZOD5EoRjX7DzLrCrQONXz/i
IH0yPFz6rV1Xj5NrsrwjC/M8qsoAbzBiAgWHndCCCD7TJzjFrvB2CMdVGmGekqsMDUabWtjzTb6v
P6KU4gSjS7WzO9Gk0yi2znWiOS9u0Me9f7naABFob62+buI3NJzKaT40JGn1T99yVrtfdJF35WSq
psnTXuguAkDJ5Rs3cmyeNF7JiuSzHLKn9TGYRZlheD6r63Z9KMnQ4FtJAmPiSpjC70va/Yjv2eTp
ETVtS42VU6mQMIrEWGzfAl99IOgoz6RpFonnZPZlXtpx9uqQp68UyqspDXY0C5MTvwK8Sx5USZX3
VS0HP5bNcMR8dzuphYk9E2Qkmz0QeympmynZaE1JOJtPrh31qdkN7ncX7VzOk4+0F9/nkqVYFS7S
bfDg2CFlwcVTSPc/zs3IedU4BxDwJbTcNcuajVpDRerOQXiHfHshHtokSRRpVUoX+Bn4V2SGMnIS
dNVxB2E57glrmaVhPUwV8DMtNyrPjzSGOu+8NPu78LoL2lcFzf/E6B+j1kt3qVMKF1hmrZyzGw0W
E/CoATq/sRxxOTfhXtYl5uS9ahLnLks+4CcplZ1ltrL/T4d8vSlry5xw98RglCRbADTglm4JB6mZ
5lUPCedaGIOYyCwzGe8uq80hoO6CoSYTD6ArByimXLnZdxSWAX0pqNodCADA+yJJH7v3Da9Yucps
GBQa84Upf0MSuisIF3C7jFXEfjKHkcm2rZvGXft9+BP1SjXsA4degkyK280OyPUUXRkX0egLzT6j
H9SH30IWYvwW0FeZ8XJc5RZQgpw7xNBmv12xZ6GB90+ALAyPj32Wu8dHU8hdjwoYzBGjxkUTMY8D
eKxTzOO+8/l4zmZYqXVdBvZfwAV1qo5Hnyn9HpbFPajdSq5LELCMvf9k1SgbvAg8Q3zIiOjO+JJq
17xdYlRbOGwTQ+aGNgD7Iunkpi6EOiDtlHKm2+X3KAJtHUTryhhAjOFIukxGHGAGDgJzLpQHZkHp
DpAgVhlCxLSEmZyaZWGsiRIlyPitOTGiTtcQwRS8cF7RxlMJF49jLmZUBz+CRyE1jy9Uv64ttO6z
w9HtUQx0kFQLhicIHCy8c7tXKOSKRnr7WPwfmebINDKfLGKK7VVake77TnRd8okHb/RPSgPzL4OS
p2UT5z4Ex+jet4wtvDlwYpI0faKwTu6TT3Qej8GGs3egWOSQLOi5duRD1jn5UAW0C6H4awFroyXY
0LVp/hXH9GdX6GTh4lTPDtRbs+3W88GUGBjPNCLzQz20mR59Eu19yz/zB0sIwWNVZaiFVt/s7jhm
nQ6m4uafDK0T92z3WNo3bu2Q6R0MTTSwZq2lgnXpIeBUGiSYYig8PSKAwkiCwDnvkAUhUH1z7Bdw
3b+/oMrYxnQN7gpvN7KUXkILn6m5yhZqQpwx/Hq0lq0wsj88RifFe1Cvo88PozdXFlTaPVXr6/Tn
uSCOYr/YiGYAGGkdCm2ccel5J9E1Zv5lo8ZUFOK1mJf/3PXQ2mv0f45b4gm7K+vVC/fowBKes6B9
UuEL9h3tqoTwT7LNrWDvVSUgH1xQKUgZhNfzWIBukF+UfkyFtAAh9DJJ7Y4SEQk1kMtgEeV6jaR+
sjenXG1Iao+4mKGGZm3jmEZKT6JdcuQ/ByiQhJ8lcJQEjjZRDmtZSG97VwBf8OaiD3gBjHnjR5cb
qFporfW9aELbbR2rCZe5mMR7XlJkfOeaeB3FLaUkqzU8HiElt2zpsnUAUZVoxs0zssVxrpxVX26M
/kbkntto/Jz1GTOxdPkcX6+gBJkbHEnSjkHBnUPsjgapdAQjK98+NTyelhvemhejbCHNZjoglE6R
I0mINDY36rzom8mZ5lF70mXlHz6wpEL9cPgxJwbnx7qcGnwy0R4XU2o7SST6etyIOG8/GNt/BRRR
NrAtV60qOmG5QmVH/an72aPWml77tYXAWsvrF2Ms0io5iuDBmF4G+1+I3XJhk5gM7hXqZI8T8T0j
AD2hGH3R9H6Yhb6golci9CGOksVWFHG/EVOUMChbpp74pUcIEZ960n72V8jcfcrBN115g407y3qB
e3R8PmRuI3gtfpz2CKM/D1uJIGaVEoYxQf0jo1c+ncw1SwZEfV1wvYqo7uhiT3IkA1sVAgjIortk
QBj9q3TVGBsHgL0oQO0Ph077V4FdPeeuBX27p9VWBU0oADHlZnqp5jd58mVqbrlYq2LtwW3pz564
FUSRYZBox5KtI2T0Ps8r+ieN0NfCod9mEHiRxIeBm9vxHNAFfU6rzHTw4bF5FtnEy2lUEWeXgkxg
AVetSynxbAKSBE5N6AF6BhCbzwWOwqKAf1bH7vkkepnmHCFVNeL2qKi2aWHYHi1u5LiVRscO7peb
9BSjuqo/PKOBJf0NfUhPbog42wj2+Bay/XQngURbGMERK3VTniJ+ixPDQ2RNzC9olPhjc9T/wJvT
pZoFOHn7XQhpIi2luMZHC30zXrzhFUIFG/gMMSs5otWurf4tbqDHKlWTVEosbBTXug3Pmuk2zYtY
qR6zcfCY8xZ3E1gJgH95rhdVO1lr0bKn6Wr4OALrBNX2A6N7xlLlanqDxhlyRNQXPVFl3GubQm7C
Cz7G52HGtqXFo9XsxRbRJJf7OMLPUPfb6Ts4eIw1C8uj1Dzi4l43Iu7C+37Oz8QK/sUhRSneKwpl
eGF1sc5igXZvMZxvkcxsbOMMpdLi4GROdZ69Y+vGoxsCa9TxnAkMMx4JuHPOfXlT+XvRmJQDFTG+
ie4hkQW31ICb6iQvQovuJ7VberY4MfTdjjEMYIEOF7xwG9Lj1HxvO3BZSVDpeogrfDlVTuGM5Ag1
a6dQGFF+n33KJX0meXnbuP0/+xoSWS4t2NB+p1dxzSc4M/KSdTHfAqzR6feVrBliSLytkq88Ll68
fZJNzzYBJ6ypWjd8IEKXTg0Q/MYN5oNHM0sGyLISZciziqRUEOCulx+nMajOuZAonXe8gsE0kjLn
M2+cbHhguSxiltQT2uu2b6aEVWdTgKTaRwTTdT4VEEDQPPxWfHXRFC2HfWDLzYq3nggE4RdaH9km
R8bOHMqjALSt8wxL7QnbcnM28Wih4Bnn9PJjV9dxMeYHeYPNWLoaEX1yoSxAtZwYpbe/uyhwSiC8
ofEQJFOX6OJuZVzC3wQpWQ6yph3t7e4YBBj9X/ASAnX9g9NmFKNyHsoMh2ckoNQ/QZjr1/vlQbC1
03s9Wbbzdv66Q13IgPwC44iVihcosQPmtM16Y2rEfxfa+Yw7rIx61YWoZqnYFIBATY3xpinGoqoT
8hVA8CoYKFsZEF5sF2sE6ToOv6v7K3oyK6RIYxLwGsyonBUKWC7VvoXv25q5bu6bLMUeIkD0ZSlq
x2bPZCupEm1BGRFvh1pqpAwlSNgnfZJ8+Vdr7RXhrXSZnVtZrONhmDlFluOl7uTx9OOBAgqtLIsO
EsqCXAdILQ2m+4v8GLxGmWR/4jFzlq1ts7qbByzpqDEoTHIlojhHJuzjBOopDvcHJeOYOzG0M4mO
mSSTftNTvVWUjEjYJxqlgNXkT+EfQ6PuRbceR/mhCqybpocUOxPmODpkZ5XiWoQMJ9qWOtOz/ax0
xh9y8jY3TDUYEMmt79XihIg5Lpg+dlfnmP0LuVDe6ALC1fg/jpe+vU6Ix1usUcnVSm6wKnmjVrKt
D6UDXS5eLzoU03fUK1WDNZMqc0nG2G8CGmUVPb/rA/NpU6/FINCYvpyI4ppV/mPEWP+swzAW+KfG
fL9IjbhtUjO4qqanKF9md/5LDvRvU4RRZIugvK7WwE2Hmfq0pLs/8cuIL3SKqMPcUyOrPGo33I+c
agcdiOCpM23vDr8qsW/nrQN7yDc6oob7qQ4jAp4hQ28vCtBi9QJgWbvIALX6DfDEmokF94+crnGW
hC/u5r973OpKoIAAn8bcHOsHTuXvebY8DJbAdD9t3LeV3nGI946JfjEbu7G1WFEeDolGginmc3mp
0al/PTOOmoWjUdbnflsWZ/aHUlQaW0gi1CUjMCjp/JZsIXo5BFUcsUNQBwWsYaSvd62qA3XNwgOd
RzRYOKh5Fzr3Aim3pKcPxgbmZFOedCpcG2eKHPX1LZIU5rHx0hNDafh5CbTnH5IYEbDGf7k0t9aR
jWSwGPqfse6tcXU5TbUOze6CaWUQwnmU+JYTrSqWebXMRLliI7yW19Lb+5I86O87WIYtcPSrqVQm
SVEwYx6Oz0bP2LreIk0r0Qvy/dZydb/EB99B1OF9wUQd19Z/2Ar0N2qYRkILFOpC7U7cGeRchXQ/
1iAowiZ/VvyYcEKtuHXov/XuXURS/U4QWhYYhMMs5igUbt0MUMct3DMJskhsfAXpuU6IvCbeowot
ZNEjYiqSvOrWEla/gJuOmuKljEhh4y0px0GlZ1f6jwY4Yfdiqg6Mc7E2M59C8QxRtZLokQSZHpet
MgUgenVUYXEZ/Nt3LyYlcEm9DbhFpZP6E7LNMSnjTUlLksMQTr9f6ENfka0fshKsCFiv4bVejTXk
mV1xaAy9Qq0+xW4RzV0/hcb6NFL1Woib1ksDd8pOut2qsXRi5PqKhdnpm5MMD/ZLfMEZ7r/8eg00
7YhiJfEjDJtb5mspfqjk+skbFUkCljKaWqiE+jPpD1oph8Rx3yXtNBSbpaE6f2wt85LRZhn+wrrB
dNirg5pauXyRiIWw1XR+eEZ2NwJ1DOiNCoW0CbF/Oeq7DCTt3arSERosRs3OjCohUKnPzACP7buQ
GA0+NA/l77eI99Bqo1BNiGaXQUI8K1xo9RVKCnmK8ISFR/YY+loE71dHc4nbm6hWC8SHcYcZ1OG4
cwIhx7nrklIU+oKxpeX/Up7AlE3rx0UR85KoeSg6ScZVRvpNkYB3tGKXkxoY4Yy6TQSDpaKP3VgX
Knxuy4QT48+lqo9a7EvcvE8Gz9OoaP4pULfOrFifmSAFpS2EFDOAiStXlYcIIX8UNWPoC9b01ZsN
1Q5/SablOYLQKsxbFODgSSZCTm2JOQ3t2KER8/T7HDRG8c8wy1rTP09TRVi6rhx76vm4HjMC9dai
s61zQyMFT/8bP/skpDTSAGm7E1zynJw0/cQ7uVS1g5nbMJn7aD+pWWiNfXNZcrS7xpoy+ueFTyWU
aBAM7l55msECM1JnU5jHw/qJYttCFYttMNbssm0hQTjH/EQJxyUlU/tslBe0kvJR+NTaJuk69nRP
zvW6YQtHS2LbX/GpSjvedNHxY3hro3iD3rYjqW7m/J3KuSYIH3MHsk6xlmVrLqF6nXrH80Brn23z
x30oogAJnqjf2EIZrlcAJMj8eMvv/35JEIAU0BUhgPkhINMgSEi9/DqRQkdUjkwvUlLTj2pHYJ4y
G5qs9zdmRIJQVH92kFYup4SVZyLrj2oEz4DU1tTHCUGjTGiAV4SGAAPAWj96p3aeFu8FdYZ7hbmb
6LU5KY5UE6jAOgEJ2ebthEpyKV1NWDxmG25qnO3BxPM7OZ6zy7+6zClN/RrSt0RUnsL3eZ5yA/bv
shO1R/WnH79ikwH+dXRckRJll9SnIpaan4eciyviK7dAmq6E/2flw5RnJPkE/HjB+Qwx/+Tru5CM
W8Bl72NV++6kSIuykcLhC7jH39dvQl5AXKAyoWmqARNvRxXbTkXir9STHvSDuz02U6cQcAydd+CX
Ecq8zHlXp1vxPBoLcha+YWIWvc1OD6OY+Mw2ZUdXL8kOuWOJclOWscAmMJZLmIa2IA/bEUtSceXN
0chkqtJMbzX4e9uZEjawlJSnCNdu68JlNZYUDnGpkKEuHyqRLogLaZAMhadWVEuObNIQ5bRpEqoa
qviSnd6lWpJ4fhM2N68Qk0yzaw/B+tABJzAVb5UVVunp6zY90GX9gj+qX4YTW2jrTBRlAZanaE3n
dGc1pGSDVPMKYgrLc4EvchoM+KtAa+qITLADLR3jVhl/JSsmCyIQeaKjeil8Av++N+vlqUFtJORk
Dp58G9hPIqpuQEyzVYS9wpn3nqz0ym7r4CX3nJSwQtIJcx6fWJOIsQnKA5lKJeY/Ancc4o6TLCpL
u1F9f9RWuunLByq8b1Dhpk4FGfjbqVsmdGf139ttgTqpxW3bbPQMJP0cl0DBZGXwmLEDvj/KBdz1
gTaAf/LAYKlOEJo/vmindVkGE2A2zMOzLg1wCEL9UYPW13Bx5rN1ubmwxomINt5LLeaGBizcWrCp
CpcS6weDpeVzz9dGTYUuFcaqI+8FjvzMeYJZUo1nV384b9HwocZLu7CLFd1o5oAj4CBeJASzDa0L
+GFIH9e0LJ/ryqNCz5HFUVP+kfA/2ulMdkD6QbleoJW+N0dfGidet4PG9O6o/VRxr504HfpiigoN
Cquc4gr2/mrOdbbvu1YBiS0t1sCSli/m3Ni3i/v0jALow0WHWiPeBak8wd8Ou2LGSyRpz5d5ctpT
0u7fltwiuGRFtm7RUpYMxuhO4pechWjvOTRpXet6YNNvdkER30WBTZuh0B8LH+eJX9aHfoxnx12N
YyLe7fRbUWb1iUuXhuFkgIUp8gay7BpvCOB4e7tclxWudyiToS5WV19jD8N29QVeMJU9zJy8w0Sm
Sbu/s4Us9H3gxPxHXQf70t575rtvbiAf0ixOzILyUT3g2VMyNI5N18UPIxGLZToyK5Tr8l5PVUy6
aPanZK8k1iS2FpnJqL3nRXWV6sf8+8QqWvo2H4Jlsmu8dip/sjwWJha+KlAXLzU1vdYspxErnb6P
EZbUVQk1Jn2qRFvxOhFRQY2y9nDyhramWYiT9/3EvrCp9bpWA+mMohb1p5FKMIw1iFeABPr4nmdx
Yg6sZaDK6X4N3RxB4SQZ96Ux0GdIF+yDbo1IBnZwp/DvLigVRvY9N3NLu1HtaNb2OUU7UnKdTIns
MTQh2cP3tvryrQb+XtByxH7todZ8ITZRyk4XiUqzsyddf8Kq4dWVv42TKfkHX50E6pmIdvW5JAAl
VLN3yyMjRgnksN3SEtqFqyKAScEaCJKcgaKB8WAPoY2yChMa/+/a2XfE57TH8D24U4j6kowL4J27
epGlkNIwumIz87dChdK/ykgpR1VlE/paTvgP8Hmb2SNcxgDpEdZppuFRql4QNeJwMlP7PLCLFPjV
m+09eEqs7WhhYsYh8WF4aPBHVLqyhK/tEv4+ZyjWI5076FVHedmRgyqN7wr6z/uA+yLLtnXt1u48
DoeRr4SqrIKb1KFSLpxFz8Bvy0I5AjiPuG4KkHrfFn+JDWfQPPMKntJVK9xw36kIvaDnBndBkhd9
DgV3lB33ehIhYXwBHTCLR3V4zMAyeQiOFdeTgeJVy+eSllOFr2E8DEZ8gqz21ZwuIqdUYPOCx8op
zhjrFueUa77fB3lM/h0ETYBfWy7XgpJKZ4SJC8Xe3NC8ThQB6MgL2id9PUMOddKXwI7JN7388ZeY
NtdKxldUuuzz7AszL6O+8+YjBstL6NWc3I4B24aYgbfqBZkh+bJkvM3J9GjoeWiERS/M0hhfreI2
9HlMaqS4RcEgBZxdPUjLRSZcIVhKejCu5GjI03suLZkKi1lM6PSuVpVA5sqN4VL4oG4+JHA7ilIO
FbZaKuwin//+J8kShAcctCN304aA8cMWCJXXO8KQ+7INg3vVRBOjq+pSlZ0Sqv64mL/nJ8BfJpqR
F7R0BHcJDxLPHQdRz16DsPOB8famb7p6g/i/ikRrttLgiZMGd089tuQXQigiTcesYeUyEBUs7PIE
PEg1QYIjcQOfJTU7WyF0Ry3sJKZJilRR/6Ptbd18r2ZtWph/5hdeQSvBZi14okDqST9c6RU28wbh
msGSMBtw9wu+enO9WC57bSpjaef959owmy29dmtGs4t8z4Mv+KKIs/qCw0LJc4ndsRJfgaGWJxuG
cYN9fkPm0kgndqmjek4UJx58iBoVCZNBlUJ9NOw9a3xoGlytrt/xusxvVD2zOjLhvc69MEz2Xhtk
+sIDaUqFzREp/cjQzUs9nK5ZdWbvlcRNO74xMp4mpcdU4jpIk7PcwWI/Sdid0SGnJBDj+pXR3GdM
FarVK808uRNSo8ZgPScs00jlJsXmoWEUZ7TmNDxdBEHxTxR2LHFgurwThWIhP+j5Q8kXp9u+QXXd
4pzNApqs7YDLuiBmiEHY7vFXMCszsCwCV36342WB7hTDoj22x48Efb10fUV1MgATiALM0vz+SyRW
+rabTrsWRS0A9jiGZB59XryizibmcPf2phIXOX19acIqxmcJbqXgpYnKGqUNHzEQmQvud1QZTYgE
eC7BEERs1wPsmMKfHQFZ9hR51mWLj7uWsY90+6tXCFLIrgYBWeVdepiGyT7/lxI/km0EoVCqRIwP
OvWB/O7pPj0CDXTWCoYE8+4v5nTR7Bsn40Ifotz/Ts5SlHESY8s/gzrIqq6Paxb2SMNA47Cq9XgS
InfDcR2gCCnGhxvasy10n+vbyDa4gQPZEg03JI3fcYzCwhexJ8Zkr79ne0/3PP09luO7THGOmxWS
ufKX+AmxEeuq5m8qZB1dQa3PbG8AZcuJ7QUYtGmSGB+Je02d1/Tf5khE2YpAxKwON1dVigXo/wJl
CmSIJbHLAj4h/DrWW0NrG0aWLwHHylA2qwEqnqBAIhTAR593KYwCiwWoCCYtqOYceOXRIKStyL4a
p8e/P/N2/akm51i/T9qWzYQ44eVyw2OmBzX3boH0ZYD6YHStQCgDJ1e0IheNCKbyp09JAUlfmQu7
/TvQpzpmEtztQAnkq2Wchp0rvwT+vgPGGtWOfgPjf4O0TR8+F/Gcy3VgArH3OjYqSMPa/IxG37RN
cM0yMkvFDz0viPNBfqiVKscJHP0q+WWUc0BpCRUQy5apOaRgo9OKznRkrWJ0z2GIHdUnHNuGSLdO
PnEwKQjncc51sVIVIRTRmdvJEeinFE54wPz4Hsl3LiYKromjWnXWPz3B1HtwheOgqgGDMhRsjTxh
C8EOTMVNJrod59s/Q2AwatCJVmpshs1f7WJPhHOLXFqRQ9xLBoYaiaYpckaZLhS7HdGyq+1W4qKj
HDueshHLTtYDY+s/CIRLderCwRF375IQctfUKYTMpp8ow+4a0bWfFWBRyvxajjdzSQuJSXVK85eT
AknlXrt1gqp2eKGD3+RAdF1AXMIcP51O66beYAV+HnIGRPCaKYNXPRNxO/7miHhCR1EhY57LhL7V
jJhiJJU2ojbpILSINaueR2Za0Ad4fkYisYX1lG3rGih2ecjSGbSsROLO3BTewGNIi3SNe31kjA/f
HYKq/AQKjOgHoEO+lx4GEbE5G4I+L2iNy63z2WvGbn13YWBmKPfCoLtvVQrGNA1rU8DA92UPjeU2
ByN4A/wpvuUkANwOZR3QBFJR9jvSEaWt69AGl0QLFVO9TiRvcTAPVnjGdsyT1rcxOig6+SRPVjcy
u+WlgKH98cIHYcjUOvzcdBHu58Y/VGEfhwLTzdqqhKqtcSvLLZ7P2KxTJicQLgnTkFgXjtl6VzyF
XuHPIRJoqdNrfWrmZYplFsK3JYTngzNJ4UhR/N44+wleppn8NcrJH9NhyYBE4C2Wb6n4rsWx+x4E
RC/YO21Wbfcybjb0c+zebLqYua4XMHMLxmT4bJJTWpnmrIft+5nCu7KwEJnI5FyTwQkuAjnDxNWe
6KP4pDABDP3Jm92GrYdWTrj/xdPKA1AB6kirkPvcIIp67JokX6EssbAKIa/T+7hfN0MB222kLbr2
kDDMxergXTTja/pTbxb5In3c2mlcQ1oPHkiQvhFi1h89OKXa28DlB1MH2bX2yRxd6fGvUM/JuHcS
EFKzltOBK22JLMj1+P/lKIyIaF0gdIbyVISIdmeXzB4cFaBAUygsH9u/SxoIhpt2o0RpZsEzbQY0
KQILav82QzqX5tWHanRe7RLxrt4ID53F5+P1mrSKenukIvaTzxKvIyPT77AeRWuOY7irjXzAQxrt
ss+TTsJmaMYZLiKiFu1NApJVUzcJp1/drmSoYOLdkIJRJc9UVR0t86SmtfLJfqSnp0EPutzaWyG+
FZsB1H+SdFzUMeHv+5lUvuhNYJwi96d7bavM3XaCNBOp0BLJxLzxHjzBGyO14fIkswAPbDnow3+9
Bdab46faM6sME789souoPRmW3EgZhJE4A3wYMbd1EBoWbMCTxgeO/tKsMIPetDh9xKfkPcihREeG
/Ca198wbQzrIaTTT0rTCYRypsCwGlDeHkiVQ4qB0YRny1CTEtD0mrZqdelxPrpZlahHmwbVj2jCm
gSQM/3pRqj3MWu7jG4RBCqgQRn51+wDG11N7UJJvPTi4GC9wx3TfY2v9B75VSEtM0+xe43jUSPFb
FCi6eQSews+sNRC3CuCS8hZTHE0GEZXUyaDKQEkMLHXkpRvv1aZeIittR/BOhqws6NcUF0iJzyu+
tdckoFN2OZ2baILGj9rbSUMKQckg7zKhjT3zPVZ9E/5vKZjl9CaE6VmADWFMjVjYbhv6t6lJvUI5
G5UJetYAqMGPjDViEgIHW2flFUlgFZjRTFFmueNEESoqJym3+pG1kYlJdmtk5ut1UFY0gGy5rc9W
hOKC6jjdo/IpU0IRoVk4Co434KQ2NNIN/wzlWA9AVe4niIe+Kk7nffMvEJWhIf4bQfEPkuH75cZQ
ziWr8296TKfYAGVub3MzIK7YHohPyIt69POWKvpD8SijCUra57TzH4FuLAsJtazGVN/btfUcONfm
W7QnZemWrpD79Iolb1dJzEFoUwe2t4lpZUwLZsdCgx41YqJvtRAJd3Lvs3zia5eOQI2GQj7gRNgS
Ij89C6DBsoAiiImIUjoApAQUew2l8069Pom/m7qaOe3fZfS7kafQbXW9YFfs6un9kvGfFK1AeLL6
04WN8YUXyxgCmMONEbeZ0LbF7LbRLAjUt+CBH2vn61TDcJ32mT08MyaNQP6ELrtJgpVjL8hp5d8g
YNT5ZE/Kd5Lfte1hRumRhNjr0jLKdcpg/IBwNsLb2O2KQFiOT/IAMlzG+VRKM3IDtAnRk4LvgFDp
m5VkOCaoOsjvFsYP8Trb6NnZ5jUB+TfUrvngKDeiU/QAML4JgKKNxKZx5AveIl56Dil11D6Jlyyi
7ADQykWmUVIq16zzXZ92CCbC/BTx0E4UAMOuuUUHscNv4DKfUIPRXptLvAjxQzETFP/XpLWYMI1A
EGI0xcQ67zamNwVg5oYuzYlW0I9hcfwOBbBMCMVz4Z+ePk04JFfgas5XgmcpVKb7+G+nT05LVGVr
eQm2+GoSeJAuB6odSQ4Nd99vmSsZh+7R9Q6JIFVvwpYnQbOOr0Lk5ZgIHGmKPRq3JVWTRI8DRP80
ihKGWeFN+tEhNasYezVjmWUuo6AEp4EK7OwhG9YeFLWjKKLRUQ4WKEvlc9zTGmxHodKtAW3N0AC9
yqkCr04qx6QepGh//tC1VgFjnu3pC1gWAzuoAEVFxGwa1fPgy7m+6Dwz5ekwx9fPoO+gnDZUBZhk
8lgtSM/hbgL2X5L2UHXQ7ed47CUdy9odJTo4XZhb5PD4GhIZOLDrmUkW9bCh2A6Zojwt2htyWhRv
TPutwRw7V9D3F7buvjYvD2LnUvKZIMslQezqRcy8J626g7kuftcv12tzEfCk0NLQngcz9URrdRZm
y0za3cNAbazIDzgcNqw/VPSBA0l/3WI52Kqync1XC0zge64J42Oo/7KUTIM2b/aPpNIE+qpoFKA7
DtHM1wFmQkwZvEaJ/SaXAtFbOtANz4UME2rQE8Pe+cBnCkjwDkRWyFxjGgSaLp9Gdo/qlR+Z0lpg
ih13bb+9ZhGch6ztRagfVCjy5/1PNyGdNqOR85UM3QAE7xflgUCgAaOrI7mcYnXs7rPnGBa6+yNY
/JqviUjyDhpP9g6OisKrJIKxRf0MeBS6yZFETN1gVjtnak6jcBKlQcsHEbrHMGOnprtIQzmtCTsc
eRoCL2DXUwqLm5K/3lQrJeC71UMpGp0PHodvpgjKOyrvPd+jjkLvpCERXpCNNcsFu64zdqI5nyd9
I+xrJ1sgpCblmce6bQs1nqR9fkpAyrhNODy49cOF7AUqi252gCREtGPHL2Dh5i7Dp06Zru9F2CAs
FzmaSwsX68tcCMFra9p3BjXiUFyxRGn+r89464cMaMZT1gOiCePMyzv31ko8vGDE7Q0xcYYBpFg2
1/f5NXjXkX4f7Uj8FdbXIebB2w2hE1J2fUdTtqrTFeWdM3C3No0jUWr0YOCAGVTvx2xraT6XzYf4
uKQi64sP7b9+lj2BBYGCfRoVBqxS/tq/CtzZPTXJxrsoEf3xFrLyGudN+lgI/SbVDI/KcU7yEafK
j+BGj0GRSy0F6kHAJ5sSfP4aF42HB2+k/R4W2gnQMOfMZimtcFwDfVVwTqw07WuZwzrpzGp3ZLkT
hgrC1o2iypHLWCnH50uMT7caH5lH+JU+d1MV+mqjVEXXHlb6dap3SATMg6qh7D/9cDV4ELD6Dai6
1qct+4dIcevUt1t4FSQd//Vf1y3J4F+Fb+7riAQ/L1l/BqjpG3kSUQQenBvF3EhfnVULMSpIc3W8
A5n5fv0TdHj6M91rhFae7cg7L1YbSQ+LhVwMOmru2AYgada9+AN6+sNST5GOrLlHC41V7AyDHfdL
5ayF1puLqRFNb9oRVP+VEGdkGkyKB75esuZFcU6agKCgOE4KADiB2QJJDWj8sT/wmUIaQMs3wT45
GauhJhkaiX1hC1Z+bhRfHn7J6/AlzXHH4Wpw/ERfpOHsYrUQMkG/nc7U93P+2nhWSioTMNSqeNca
1KitXg/BzqbK0CCiowMKV5aVMoZfgRGrzGeTzEiRaQYyBBbJawY1bBpsJ3IJmFDynod2BjjHo6TC
Wur5QpIiHqEQW86x75WkkRy5mD4gzXkrMJbYG1cHGjTdIe78MLFK1/a2fxA7braWLqorUIAKz4st
JtskhquXX64SyG9HGmKPxiiBL64LrAkuTegKlMW4KAizuZY8kMmzPzOmaGI74nBs3gMhPLf+Dp9n
41m01IoGSbpAZlW1vLt9R87BAFad8D3Q51zfLLzFCFZ7HqZ+V9RtUDv5c28/qaGWg43XCYnBIb+J
eYNIG5qWIQC2SVdvYV3yCmX4rhcrzdT78G7bnBRtNiVkD6IRQwM1A0ABPR9V+Q9cw0b/KFmHxRtW
5sO6vXb/4XO9+Psh1p5i3FfQOdp4gDt7bXvf1yO9CZF1D8ul9tv9UWGgmvJerGiBNyj9M4Hk+RU1
psaMqjHgEIW75njbnpjNCVc3TlPP2cQuvWMEhFjqpF4opnCgSYv1bzekSfbAXYxwtxGFKBC4U7lO
/xoXzziwydWLUZXYm9pOEpAbhfxSnJYqKG9SPHKqA8/JCPTXwdfPum5l4gqS785Ds/WTru79ykyj
l/gjmvSlHu5XGd7aeZ4Ih9jEgfvcd0aozdGGhypzPOsBrqMMovx4/iAuWTIglyJif8pQ1jlAgM3R
/XxFAZIS9w9iYQAGfYWQdOhkGoP8xHzmzp8BGlcQ89iwtDbNi8ThUWdciZF/V6D2BM/ljMaoQUNo
tQieuGOqs1zOpqSs9Vf9SaC9s542w+7DEtr+EHKBUn5g04E0WV4qSS/8C180aOOdU62kWSL+W0Js
tr1rIGL/iP0aERyJeIn0vUYhnayKoDKkHg+sGyeduNYhEbvbcV5c2tYdVXJQLH60D0H4vMe3d5eo
/QZpU/5oV3bJ30MytHHEvMMSwqlwS6YjCOnZK1X3ST4rvWosU6b3rA6w8VEsJj12eVWJ+09xJrZf
EyQ5XUlXVYp7/xpKkKxT+u1DQl/qNAK9qvoTLr4r2Atq7/li8M7s529Jn5/JvVPwuVVJgxehy7Ex
jq5Fu702hQsjSn+vqsExo47ZR52fGIVTOgNrX6RjDv624t5Oz7Mh1o+SrNGVgBa4//FVuqd+BgYx
RZmqweohAk4rIUGTjygjFAtM9idz7rLY3n9bEQSc8briLLeCvNAwtRWKz1vC+DzH6t+eWTVN3arO
tIzfxEz2odIrEiKQocwNdxhKhCVnzPvBofcQla1ClO2N3vTedr1DfiR2OoXmvVPmd8kcTocN1gpV
hlrddyEOmDZk4QsvAwzdSVjDU1YpNLCGCKf6rSfspDOXRK27tR+2qKn02GOn1NvRwb4hqnIFkPCj
wCep901UKyr2/0x+nJ/AAw8brPkg8twDj91Xi29ANtmiRqZdpBa5joJMXwsRTuMs5hmV2CWRhn+i
1Ox6zWTpNO03tiE/ePjc+60AqZmRMANe9mPJF3WfgQepeE8mEH2Djpf7vO2VBUGfFPYMe2eRv5Bm
SiuI8d4PHx2w+OdSfIxn06xZpPB5I1/3/MZ6NAhL1lNcezUqucxl/SgV/ZFUVuRwo7GEA7T9SxCo
eqvJ9+kzHfih7KC8SPNpEuxKWhy1M/0BL+Rsb72nGmkeVKLvCYfhBELzVvWXWs3IRnSJey6WWNTj
DZi1+MxGyajb8jqeFwuAGCyO7E9KQMz278r0JITUjClDZO2Bk35e7I06r0pUM/8MV1YtWylgPxNt
oufvCgx7y52sh/tot6XRkJKhM//e5j6fPxKETPRyQoISkcxPTiTRoxl3XWOglAbcDeTTEN+H8JPN
Vnri1Q+CzeNvKLzLF6sBg/zgUFXOwTnlTncAZVKfISJJmNp3DxTxmyBmKLknYhZZW/WD5yXbiC14
w0ODpWoGxamDCoHJ4RYC71toQSAlnkmUHBlS19Q/vIONdRzjll8C8HAMPZti3PVs8bO8Umt+ihJ6
CZXDJ9tP0MFQhHWYclXlfMXdJCiacF7zKagCEJDVCfW6be9bHR32+x/VMOlhwmpdkRPrwEqAq1MN
vo/539v1kCpoWYWfhwShstt4jSuAtdo85PvgsDEPhEN+8PMxLhD+1QFy295IaCeVOY8dRAuHZNPZ
xA/zHsCMX0Rv7TvDjLKTYP54Up+tXunw/KTs9MjA55qRU/zW3v3UgblBURIJAO1WR51ZNb42/cPV
iJOULyIh9vaKdnk9Em3UrQ+a+g9xbahbvumLzGOK/ocoCz1HG6ULF+9Fj74OTxlh8KNICyle0LiA
6/5K/RkeV241i5WzzSSFlXU2+y84MGdUYrRxkbQswrfyd2/r/LfjGriirUSer78BsbDPfbFZQ6pw
YKbsgZc84zH6lqlcbRlqweJRgTD8Hnd6hE3W3/3paoWn9Zt7st0HSiszv022m9mVchzDmFh7uX8J
Vrz2YKO4uqzOasWo11c03OYsw2g/Q9UjiZGys63IpOrcyxGgqqhskDBZtA4XKzqebDCSiPwF/MU/
teiKy2ndJnf5L6VAeTLT5fkOyui2JyFqPL9m8ra+5DqX9O89L2JZf44JJlYL5iYCwjR33boShm37
QiE/yVR2wPVlsKvXisuF0ERSyj4r8Lytw5fPPzVUwSa6bNzx57sKH5/I8hC0PjUTdx1caVB4SLG5
0taJo13uopZxb4g39YpkjGvBkm15oN7y/SjUdSXR6jH9icE0AZ8RiTNIymzy7SFypbPHPiPHvorb
2nkxUBgffs5bCPNDACz8UnvfXJ8WVi7nEF9M1bM3W5XfyNmSzhmgN5OTKXrLXphUMajdtoVKlYVQ
tQuaHfDKLvYSx0cBkpDMaHQk59ADsYF0ubtdFESGX3SiHypAx4Q8I1rihpvJGAcw5EcG11e3fP+P
9fJvHtDyL05KMUmAE64HyaB/157CZqWabInpl/hVwnh5m2qWN+Z+CuqTkQL+3G1x0P97TPT/0ouf
7fmlcDlBjQqtIxk9DYM+PHzJi6cYd5naVUuzFJC3w0xMrOsigTVnhlJjpmVugJnvLagxpd57sVvU
GVMVt6wpCBMtVyOcaU55JH1I8LzVJLxXbO1BuMQDAQVSTzKejD1bDzkL8S1trpQdrzw8VJ0p5aLp
Qq3S8yQAELECGvJyNu9a61jTtF8oz3FFuwc2+b4UR2zpHIUwc5cnfNdjPTFD589rcl1yrcqLrweP
O7OQnH4WLU/cCYS6cBJDM2R2MXE0PiLxYZMOxt2KRwFfh5J1eOHACoP1MwcRrOMDBh8ubiPuJ0aI
xaXK+CSOjq9MYiddDEiCkbiNt4qVoeQJnLYhRk46W9EZU5hKZykOSFF1IJvoUTZkF6Ir3o67vHf7
JpD8YzPi/28Q02bevhNRqvFsU5Ul+2lFq0n15BsTquiQm+7WbCmnRkyCdtU+KmlYRJiEI4izIPix
W/R4raMsDgDYtNy/QarMjyOUCM+uUgQhxS94fTTQuA4BjZwyFM2V4xX1QrpSPCvF2qAeq9N+jUye
B55tCqXlxUjexViTvUdSv7MkY4vzgS4WWH5w8nIXOOkc7vA29/mdOMxYIoxdYRWqBdUW54fZehZD
61JGwf6LkRbW6x/AkHVL9TuMlYm1cWDogL/qzr+WCOlTGkSPg46O3KEEFzis2vtUSMUYBrA4951a
0C+q+RV89Ju8yhrvDfhc0d8BkAtMccUvBAxsJ88PyV3c7154e2s1cedO0MKFNeaXRkALgywcfBpO
KY/85GxvtHJ78afhFsBRBsNOavc18p9ZHwNALWCNj7Wdjjd8CIsni69kYLlUBg9vxb0pQ0jeSIKt
u8FxYKPQDtnOyijDD29/ST9Vo2hUVATCy82UJVisfz3ukaz000E9BnudW1CpTXVWVTETcUTUDqRS
OLiC6L9XZ88U6ZRjplOAXcCJb1B3BTuxNEYN9DUiCm1Aja8A0j2g4P3/2IMQmbpcG5K8ASQJIEJ+
eYH3KuAwzrWoptycVtGxf7d9QUdz+ri3AvW4/hesBGv3vrYPBWGKZkeICPXBAu4XfB4/Z0eD+Br0
DVk2uP4evwoCpf+PPe1dYHVBTG8PrD+KgqQMhGHuJ78H7NCACAxZJnINB2NQEUfFc2BBqLy3/uV4
sxAnTspsRYAMb2UoJ9FYJ0dL9cCfZ+RbwtbGJEfnW8sZBM5jTSDQfSRbbtSonFrKdKz4JxP5VRmK
dpw9izpR9jY3MeWvlCcaFwIa2gVKCC36IyQ6W+PRPAr/TLMtbCwplvXFDYGcT/OdYfZXZsQoYTVa
JtfjDyCV6kijncEF8+JyxzxhZWK1GkeU1WIw80COpotC0I8rjbWEK4xGpkxQ8YPWYgQhzKjk01fg
1mK/1nK8dIn//HGYKId6CGdqp61kvQdYyh/3Ecb0LMP9bF6UIW4LcYa994FZEF5Ma6l//7EK4Yog
dD4o8MCEB325JWNHmvEGwL0Z2iybY+OWvxavYtIo7Fk/yhasbjlNHxN0COQ9Gxlw7q0FpyfGozgL
aTPUWbp+L3MmqQIhnpC3M0qHNIFEp+f4yHcjGVgp3jcVSq+xUh0vDnp52lMWggMuIzp/js2aWjXF
fiXO1532ojs+WorYOtRI5B8Us+/setT/6SPzsTEo3YdQk7vYONFhZIU74/d2WWw6kdAnB0Ed+IiN
cGqnD/ikfDsKNecvipMeeKVAVC7WuIeI28CRMOTRkyJ5jJvBthD/dgLR1rAouIZe9cgb2dHs+q34
QBx8ZhH2LVEL+IR2fT97vR/EYhR2hG8lpUpbrbpd/hCcMC9Wo0OAI0DpxSWyS2pVtwPhN3wqIALf
eIFIYROXDLh5mCr07UIetOgVy3zBhPxokNvgLd8X2TVEbK8TDhUSnNBg0q84eum9MtDkI4iLUwlu
oh0WSszU84TZBdCj4k4qLlLNgF1y3wZzmNyyiWTxxoXICmUh6Sk2SQj3JM5V1Ip1z5t4u3+EHLOH
PHedn7QvVEKCG7J5MyIVlrNCO7Igfa1nBYsxesTUNXlubUPV+e8uJ8k6F/+KxIy6GkvidnJpQ6PB
sP0eS5vdyruA+dBO86jEh59fwdYnub+CcESkpWqcgTj6W0H9byVmxruh2YXduzSB2PQVpAgM8ogs
uspMiW08npkEauxDKRT/YjPrMBiWUOZdI7KkcdQ+S1axFN7F9nA+JPCt9k66xD6mI+eapilb1wEL
Sgxwq4rH1VkXxpBlD3hW+/HtuDbKxz3r8C+u4jwVT2OXU0sEZqwILQ0KDhipCLW4p9hN7bixTWOs
PCG3hBCDWkTqg5UjV132n5xE5C45Z9ZVpF+DGks4WMZKjKdB8AMb6r6M392YZP5wluKr6ZRmoSGo
qmnrlyZV7zsE8n0rdvTdD2YtPpXXgcLxJJRrssGMY/G0gKLvI6XoTIYRHNn+b9/m5X0IQTh3ZIMX
McqRJRmiGJu5+21W9gfcfDSd6s9CMbEJ238Vk3CZ10zvVWzjHlNMEhIDKQ9rRTvoLpkbDYTGWvoO
40YO5GNMfag18RkVQz54sx095VsfhP3zaEdWcD9TsouKbDhk3Sf1NKwsrx3nKgAsFCwob0Dyeyka
ICv/DEYUa9vpzrt+94/9odlQFMgVwaYFHdaZ6h0oFjUuXhRn9Nme/VCJC40Yd8H1zl6bX/zh80WF
dvVGTsDkWCibQeMWoSBqP0imsuUFFl5M54OpZvouP8W9DJKli6BQEO8PIk0H1pUn2Se/rd3oCfKg
UwbgzPuxYaB+kcsZQrWSArjXeUWkexj0JAqhJ1fKhJZcfjCrkkDe/5m/bquELGqW+Y/bwHWN5kLq
EXNHAkpC4i6l8GnpC0SC2CFPBoSRh1KGgq6GFmdKS4K5Ov5L5WfG2rsV40qgV++FPi6mSg1CTFWp
5z+Ysxirb4N7kKFF8fgwHM0MoYTXXN9wAnhos1/Z+dmk3UH96KalARZqvd5OUiSMFu1t0bSK4lm7
zA8qIcrCZWoJdmMeLUi2nYa5w+rNdfRGa8YxASsw3EQZZsvnyVkDJPaS8SHY50bf+16As1cJstTm
TRYZnj7IotAL9FLTabTR4APwi04AxqdjGks6igXG9MFf5efjtO7gDKHiFWg+iZ4prwwvcHG5bwU8
EmlfWKnWcRabzNgnGMi2HQ1LngJCP1DDSXd5FXoyvNOa6c6842dyAxd6l5fpvaMKyigMibkMrYKG
aK8M+DrWrB/I+DFunp9txBaSwVRIK/NDwzidi+OWWhqMC2rUC0c6UDN28fHS8ZDd5G6S2OtJV++7
EYFw5/jeshgJSE3rfY31K7miiVxij/gDDbFhuMn2NVDwFNR/u03kbI1MbgUsEWR6YrAxjtFooYWt
eW9jeE0gcDgKXG5rF6WaJQiuPFUYg0JmFQTYPrKEKyEeV+U/pHQpu3W8K13UxvtpEFCYMqg6RY5E
B8NY7WU9TCfk880OF2ZZlTqbTP4lCPje0XLTBSgHV1EZeA1QF/ldRBhU69aAiNHSteYCKok8v4E0
pRziM5oPVGkaAU6j09cN0if3VI+kPMhQ0n8qRjSkvgbcmdIZ1p8hCZWrZZ1K8FpKft60F8wei2aF
uzuTfSn2f2R4hpT6HGLUxWxv0DxxrRljKpxDHyBGKllXILFA657HzHbUikUzlTonilb+MTrEhPe8
FWrRR7olBldeViP0JjJsUFMy+dzq9CgWKfyIhpO5uFol78K8ZLxbbMD7IM7SovoZToncVZOtUegB
JhHfio2mKrDwLrxAuzXAukN+hPIK+QR9gIYfnhBiHhPyZlW9T8F8n6Mxirm1fCcPGjvlxQZc72sR
pODxKnUmFtOUHTlpNZowm8b+0Z1tdmrdv6T5/wOMx+7wZ+Vkil+emNPuSM8jqgT5uM699fcHhCru
V1iPlSfFX8JeVE97DztKJUWjixyzTyhZ6oxG2SNk3vmehtkBUrniDkib9QHa6owB4recadffwvjc
U6Ihegki8S7SplEuZ2FaJb5PJIJL3YiZkKti10eVtLOyS/opFndkA9h2lvT9avL+8IAFJBWjJjru
AsLUG+v42S8iEk9ZN2hqooQ2b1uVQz5ekLCTNAjM9F+xOVliIHW8Qp7o5JdRxiKDMuHYHHViKnXb
RHzekU378rgerFcWmgBbwLNTuweDZnizyqEDS3BEaDEfbNzGUCgbHy/t41wpNBW70Nb9rXB5XUA9
kAX3ITYzjChtNNwldUn46s/ZNug6vGJrceEHjSfgvXRmjIRKYI7NYb7rpop6dHdAzS+hc2ErD/hi
bhtmh5SfOxuJfyRw3YvvHO7jeslqJcZDEPIiCXae43OR5bv+XrT+vfYBHaB7+Ow32z14EuxwFqth
iEzcezVl57Z7I2XdhZW4M+0XXpX0YMRpxF7FSYLB3txHEShUr1qN7TiIbz8Gwbje/ivSj9wwT4Lh
8Y+AoxSocc28VMYBjywIsEQJEwJVCb0HXl2aB/KYxIX57bPaoKyo2ZuaiLZsgY71Jy1DiNWIzKV8
oGCnN52jSDx33fBPG0lnbrLzHYbFoXTZywCR+5jAiw3r6tdDPEc5mNT6y52MnR/fcgxPgLzCAclb
F4lhzmr8oUUgap4sMTZFVyeVf0kPiu/Ku/2Tr3vAx2XO8f2yqlMYZbaLCAy5JTOpcMx25oagOKtd
w/8FGcSm51nYc/AP1lNoNFfhgAP8v5lsN4LeKb+XwwIb35gwEf1ED+90jtqTX0o8+1dqhX37eNX7
rWopTKLvhZGkDlVJSWKE/i/ypPmqBXPoPaVweLFFoXmsT8h8Z6Y2s3rgmWjxsfk8VPJCCeGbqyaB
DtqUwoWbiHaY8rjJ7CbSjcTn5b6vbObWiEDvS6pEbkOJd/yNlROQ1u+210xYZUWPZEGl6Hmhf3ua
J0Zex0zSCFizJ+5c5EDCdv572hxD5/WEwwLtyMRe6HMth5cCsVpVq965arcv+HH93keS7N4d1fEW
/e/dY406ZZeLpAyRpde9p5B9ppRGS97jTwskdDV1iI+YHH0EcFKhcelTUDSB8EVqe5V0sd6ntkkn
YNSwnanObi3//jgNyQk+Ac04OgN26HFJWzWHbGe6IYjUsGAdpbP8GMEIDL+lJqymieQOvt9doWyp
iaBmASWk17YK6js3yfvFalS4QRqbCJ2LTc2M8/4m5I+mgjM+oflEOr8PCkzKE2Tph5SbEsaBEhBb
l9ZKI20bw5spe5HfmaXNafJ6zVbbGpV0Nz0QscRt+LjTUVCgUA5BMbwkZ0xjwyYeIFcAd2wD6SwF
fMrNYHsuvXMlYVGLgENEKzUr+sJdB7mJiteE/lOVwBXQ3ZcyEPTNBv4SlVQz2NvmL6u01lXk+jsX
JXlULyuhP1KvLI4WaSCwQW3f5bybSRfCWXbhZpvFe9f8NqW56FsPOoSrPN/mh/1rpcOVjlvbYAte
IqcqhjgApO4ZXORx3D4qGmaIg+nPBjODfUzDgeywAC/I3D1YXE5UrpIC1EjkadEUph7Wgd8CzWJA
Vv+mhaAjI7dAOk13ltKHrIkyvNzceD72pjeFBAS1iS5re4YmZji+xMOs9wZpZX3reI9Foyf1eDaL
vKYrPVc7jOVNufIfy5pAq6kwoocun9I+opY+L3Z+B6ikICIzzk2APoF0jBVpSCCwUbTMhMEghxku
9ZcIV63cfUrsVEsAKTvJYDhIjDa46apn91JohCQ1HMMlVejX0trc9ToTDChMA/oTByNMNVV3GaaT
HNMmHCqu/w/Q8EOc8QoTAQ6IEdyr2LwyKBUoXbOHK6wrwzk8tbGYynXoRxC+RpdWn/iAmMSrJulU
JtWcRERSpyGqHPLdm4C5WUPsU2JPftd9jtizFLN70JHV8UT7I82UKt/SRxUjGXwfFUGWaDMMwGLR
MVnnYuPCOf6DUiVgNgxv9UkhclganJWpA0IzmI6Rhzak1fwBR8cqvzGnir8JnCmvwoRc7vAYz6jd
kUbveAgRoPHZU7k7hMvbw6X2wOUdXYpbMLxMQgzTNulgUUl079I0fF1oQqHN8xDNScMFBHpzOjTp
LD6bro1FmXZosWbG7oMUdbp0VVEVGRiU0Ygd7k8wklMDTrX3wqHrXBul2KYKRSFhNezrf8tnGoq9
NISUa6+Wb1zd4i1NV8kKBUHnuFkwyYpEtieffn94HaLBsuzLzNEkc99NVl/eSUmRIZ6f0Z4rW81+
NYAJT3tXYFNgaDyWqcDdOEv4xzs2eJcnBouZZOSpKJQ5K5bIWFa5YrgJHKsKrutZX9zEwMI4FVaC
6PC4qPvx+zqUkK6cIXQfadONeuNjZLgptkzZmmO6S+9eOQ5pX35lv2izwiPRXGpBOUl41jo8rZ3k
lCNVBItVDFcuIyzetEVR2qjMftg0rW2AeFph4PC2FZBht1Dwsv0XmmEF5o5slN3oktDPKqXLpH8A
TN//wJWU5IWvx0XhwhLucZYKrJh491+CfTfCaDa3giHRO66PHYMGYa47YclWA5hOIXlma3U4xD9k
j3ofRomgIHbzSaiFXNuoFskkW7GWRdlJn5vG+BTgPWCjcAaCVmhC4LhelWrQMcfI0Dlh7t+3s01r
MZvBosRCs0aCb0AFebXkRyeyhjKq7GP60LAsU3IsAGdHkiwJE/v/bZ/OWbXe/ojLAmbsUYliA4N3
jrpXCcV3NPGQl02NuzDLgoaCZaeWn1H2OwJTXPERRpLU8/tmBoe2Eqr93BaZxGNEC2qeb96qGvuO
9SaLilb0oSXaP2KFjCY0ND7oq0RGKp77pnq4vOsuJb3VLjoM1hStsdlTmoqIDJg2lrfgnY2JnUK+
a42L32KHeX1XHyIxuzeltQpv8lqJc101MbxsIuhdzF+tARiruGyzAVcZFPNZdm4SdyFW8gGAAN2C
L262D2RE2mSuIoFzSIzDgyyRqk2utdOCtKzavtM7lwW3Gpmpck/Py4i2WvDqcyypnkdxGo4bLt99
u8gsSqpbP83uREdCVD5mlOktAm5MdpfbZ0QIcHjr9qybQeu4BZIuK+g7REfiRoFLl60qb3GvbRhR
TwSeIX/TD29EELJJYitkNKCreNl4vjWG1XrV9Ag4itBNmMI20VzNzMC8aRKGtGNSix5j2/1l+0Jc
eeN3O0TINpXW1lnjhTrZyByKM0fEOhsH5FzGrml4U4wgFaP1FZcClFPWrBVS4qpuYTJ7xxinfIxR
1W+ojkuafWzSZafG25LFxQnEuMKMPgVq1s/PNmdCbKO1frj6wbzH7zqSYp0HJ6pTBV1FsTmqZ4eJ
piIqJLESGOEWMhtnDSLQhHL1Qvd6XEBBuwDbl4KNLVAR8k4WlAidWZ1qGOqB/p6DwCA74izpF+U+
TairrByJYm836D6CvJTIoXjippDQniwgtVVXMAdKyXvZ7OLEZLd4eXiIuGf0+MoqmTI37sVKdSq4
cvchjVXg9QPE9h+YgZ7bo7f4NQsVtoLa45pV2l0Ed8MqIBnDewgweBLtVme4BTgan8CewwKKni0h
qv7JkxlCTkpdgt6G83cX0mwNfAo/sUgZj8SofsoK72o0NEk0dGzAitXryRjbncZZXu6eg330ZgV7
M6ACee1JFHC3kRCVBLnDfxBRUaqbSaB7gtV9iGo1vuqvSTRd2aRzciYKywywOSSfv6NXRX0yaN63
78W/BEWrpFkfWxuCJnx1Qy/eGN9d90QsbTAkcxdZrAkG7NPkXmk+hSeMD/ulE7yWM5PUmLLv2BFs
mc0FTCd6eBdZM9SNvckVvLjVEfi2c0+ws9Xe/vlaI7qZRTEFwH2sdGvn+2EcawyZZS6RVMHzM7t0
E3HtExrLUXszMt2I/8jFliRdM1nB+KIOYV654ixrVzg2lAIjSNtbsbAu3z7gOEOpGqwqrUA0S7HF
BVDMHpAynnMQaCUjkPREk8YIm3Z1mtAqhpNQKy3eKyLk+oFbfpQKEtcwGeT4EG7mDiA567EYlmWw
IyCqSJZI+/BMEfmXmXdcYvOdAL3z6iZZSWGJQudmQ1n4g2wnByhym8Rw1QR4j3b+wU/DNitLZ4e5
Lm3c1MsoGxZ2hnupeUXxVhwxvblzfpYaHAkhfDXHwM0BqBiJPNq0zp5xseAJJOXyRl+uP4/cGQWP
vbkMIG3a4r//oRFccVA0lRsOZXwTIy9FOAMPMbnD5a/Lg/vnuR6tycm4msPDDGHkWEOriGFI8YbD
eElYny8QXoGl6XqnQ71TGaRTDm64fNR+3G14jWHw4+mA3vvYgm+rpq5tWN+YZTSUMWX18o1mYJey
zuYDLCnW9vaecoXi5LhQYN9+FAnvu1F6vM5mx2sy3LhTKVEQhkxZ/es9Oxa6QCCSnhoAvMlVHO8I
410P02Q7NNWRmqZwNEyRbU57KVyukw6PUFf4chmEWVIz/hSB9EuxjZX1PITHGNRpU/gM+qM4B4Tu
gVmKJ8K2+vNyAYEuKtMvY9Gt4hkLcPGSp02JkSa7eOZvBFzC2V81K7gsXV5fBqA1dnD2S4ckqKo3
yKh7HyF7/veW5Q5ZNbJGxfp4xjT9Sh+bqkQWVubWrfniyjtRYs/cKSsUKqlUTrzDt/+OJNBMZSy0
1wg1v99X7AsQqeyNuj4iSmtgpeJzd/B2u0La6geXuvlij4uQrp2ZH9NaG1MZZ3xdwDOg/tr83tNT
S/v7D6nwIhkoHICbcUuIfPatlNvO0jcgnONq9pInNJcy+ici0PFB7/Ix/Vht0ko4OMTk6ADeBYSA
fOfY5tSNAKn4bqw2+2CMEWohZLEiAdi+MVWCtCDFkxIdCti+yz9AeLKiKUPxu5htzM5OTsKa8vJt
nDny1h/fcas01z4BdlWkRGHMEufqMFZbUu9DRoqucDt5mNh7gkrsu512tI4cz5xZmB9kZguz2pUu
hpKXNb8It1RfBVEcE2WZf6USHK9Dcqe3MmM+BjBNi0BHwfcKRaBzmAvXDUJ5S1OGTW8Ldqw78lHc
tjoPjuC5kivrBnd8m8+utrAmfj5uN2G++z43xC33r2NdtxOF1F7GX7gfHzM26Y3hI1/n2DCaVmwt
+rqH+7GHSfXrbQoyI/YDHSkOfjsfi3KMGop6tIVGzGkEgKN80ufeRAmwTZOk91RBSAIW5CIZkMXe
cPsS50ITWorMeWI8Nh9Q1WvVDtQULx6AdyZR+GT8pWbVi0rY3k6st6rM4oDULiEMgZ/hTOVtTxrj
+lEOz7w0R1kH886e2aubDEObPcsHrsgIqNijgAN0GHdHpXpggpFqIH6nceO+5HjAlQHMkVIzMkGZ
biG7VcLAyAnfVrs13cOMgLrB5NCjXxzKpV8KOF7TQqDI9bi4LE2f2lUih5Ri8I6CyZcfXikPO8sf
88eMquMRWRDVRL1XSTF18c9UgvVxkD39zjfSstnd/vrtOzzhvg2345oLZLLsBDcp56sNyC7Bupnl
EhjNlxsTbZnwK+q39ORJckrmCW3VQKUn/8ndhf9N39v7LuVpGnUtAaGzEwCnvr7LXJHBgANdP1ek
psY7PexqEVbJh0md41oaj/5lsKrqXQl/omMqDpWCFO5CigNL80tUMeFZI8Pto5iDdoclhkVWHkrJ
qt9ONjYJquNJkO+U1IuJCqKsEMtZFEUSpEd0w4x+y2WUCKpTgX3wipzBnjftYXZjhgoQacWtPuXx
A3WV0HnLUgaU0ytHkxZqYTKdRUuQ/lcu5XtmEvtJNVD3DSzMTeb5HlVViRf1w/O0gDKkZEDBjA7h
XqLlEGgGJRan8IVL5sHO8/TSNpePICwOJNZRNmN9k0p1JQNtuXsL52pF0Fk9bIODsZS0TaZVVEem
KurorLEN8fVHyqLrsNB/2WaqabExfLRG7aHPgY8iiMJGLc5WPjQshqqIv3kuJ20gWKiQsO73c9UH
yvqHQN+6BS+Kvitb1FWimH8prWf1uVftY6CyQEbE4Nko+Q8NOoFzVDw0/Jux6uZHAkRJ4xthoc5X
pwhsD8xi4F9mQn9DC1sZWSjtLdVFvBMsph770vJHvaeSEx4kD1NpZ/oKllZ+2XSIXfJNCSYpMJTb
nMKxzELSHC7bOsLSF2nD8MQRO2LFrris504Mg2f6zXhP+Xzqth81RVddcczrNP95ivKMflg34xDj
xCCubSnAwdKHAwwmfA5c/OpI2rd+Hp2JIRmByJxo00ifoyJMmLHXiq/pkRyjl5Q5vf6/RJ/72UNd
hQxGKHSB8gov2PYan13h7cEkABlImZvq4YmiUimrM5u4ui/sFDc36hsNHidMLojTkU7UCizatRjE
gwRQYK6QuX/m9yQbZlINi7OlhKmz958Tee0etKaLzKVn9WBG4KuL/fK45lH/aJF4CGvgVw6vOrCz
YZL5dhCgUVTrcsmImTLbmQfux6Wi7EjvPR6+QbqXbJFP5pQukqNJRj7fW+7NbK4OyhOaqGDy/P3k
tipfw9HjpPpROFMhAL6UL9JYmQM8gk0BIXzbzFUzrrsZ6uGPx2dlrSmLgK0BrzmEctm02269/82T
pOpJTpkg/aVqkkqdXRjpQlON/1uiHApWsAPPErXQzEBi8XNqRvZeVam6cHcQHpUbrSskbNV1Ll3W
0dT2ICq4ZUToQL2zUZA7614Tdty4BExVPpKFa9Fuk929fZNgDsjJBVFOuuqA5EMRFa6oBdTwayVN
BxBVQDaRjhIa6QTlgqmtu78VVRX3Y/eBAb/l04dBHm1qpd/ETxAr9NFCEVB57Q28Zc2Wl6oHcyDF
AqRJp7D8uzONq5QO7zZMF8TL5K45e8EKUL+vckULYyySPf8L4jCvWNNytXbnfWEL0VFlodY6x1E5
qvdDobwMrnkbMl0H2Hzh99FjFhdeQYOG8qBYizMXXi/2EmMgJTbGhKVHcaSj2ys/sveAiwm1V17F
KK2EdsOjuLtRCkn25wKCmeI6akl1pUkPSeJj1MIDwt/PHCbgswrh2EhO5mULyJajEnwQwpO562LW
Xk0x5874q/FGSEywYUlUc3IIgrYPu4MGQiMx8MlVRsNmHxGO34FTRtdCaU3PWq5k1liAzbJcvA/a
gn3HfvFCixiZ6uAWwEOlF2CJC9ZYEt8qUQxeGO6rAVjN5y7+79o6TTrhb/A2zUm2Cj22Tt1Jw+i5
F8VMNFBUBj/gTkEuk/tZcoByiWKFQ9Gi5Pva0gn3b3XOITWowCFUeRdDFJp9NQVuZziDFlj8gtUz
RWM9fyiEOM9sokzwultKmJyd4OVKhLzMaZuBQPHq3wBfcmCyTVwNO7Tv6ZjbDPk4zMfTwAYc8miy
uUqUdaZ94rv+Zgc+njwVrzdQWBNHVhbAgNqqX5dOzqt/HS5SGtPw+fX7ubFV3JVTtnsWVSev7I11
EPAUcV9B1+pTS5tGhhlp1/lSsTNU7dyGiD9zGGMvXRB6o1O4Pyj9a4v5IeLfqqiS3djJCz3Q91o+
v1IispS1aWYrR3WWsf7F0GwtiLY2dvDDHvfiqsWwtktIgQGFLL6stfJxybhTykfOzVLnifH6aGme
YgrQBcBxX2TTsxE6lPdcZli39BCEHXUIcz2XfR8NDzU6ZMzs4jrqgTIh0TIVtDjJ/VXylJ+/z8df
bAS9tms6NzFqHtQA+Yuca2qBRIz6/1icEGHKGTb+YmKh1Wwdi5wBQ94SDVJ5UxWprSoT3ajuUXrb
Fgldvf0RxbKpsrPwZmOPf7NVqpZLVFR0ak0k4IPOr/BcihTzekfJsK7VXjjMhFGzIQ2KV+c794iC
afkkX02NLKhANCaLaPFIBE7+rnNRJIF1SkpaKT9BeIMw5ezJdnPNkSQyJf0WcuT0TpaRmLiIinT2
PZIuVtH2J0GClEYY0/LHKA5d12fBo+mbIT97ApeYFGOzOtqu4qtZpPpTh+zxFrQ/vHEPNJv6oqDQ
2yIhht9IRS3bhcjM7o1IRdVAmrlKFFoH0WeRyEH0O2Sf5aWBnx3SJ0QLIZ+fwTadnDD2MT0NGy1m
P8tkCKol+bBLFgBVGAB0CDqz48/afabGMH4J4sk5EGwZSo9H/zjbmthOVtJi6YYcLhbMonwh8Zcg
9UJ5jvIYfWHHaitIRI6mB6KGe4Xw1tYkz9gxQScx1/SCKjbVsscnMUDz47A1mUWvgsQ+MAvcNYjp
cwbT/s4MjhiIHu+UBxdAMa8CMlfgVYT6J+fLrXZUhsJV7AHpMEn8wlRgy7CCYpe74aw281ZGBJSU
LrhwEeNe+RQKuhB5DfSIVBfzbnlz/DZqMgQvFzAzVFfIML7Bx49qEJ17RMKVPXKJzcHzVSX8MVGK
8kjhQ1ZsQwb2mh64jcrX4sEdYHdc1vevW26JcbI6DNKc1nK34a9uFBSuhUfux4ulLBgnkigkTThE
SXHL/mhbcN+ln4zGlPr675SEHhCHUuZxtsB5zOUgtR1tQ6zUJequ0J7ATu/G1VfW0xApsP8P0VwE
Ilt4wT93xgWyxvvLziafZesY1Suh99MV55KdpKTa8WVMG/lWFbYhWFktPEhMmFs6TzxO1XwIXRu1
DWz3pgnk8aDsOvgsP3/SRQgdjV7iz/O+TELRjaVo480jH5+wzUkJhmMtkvRZBtrGI7DugeDWm3Rl
H1B4JyEsOq86V2FBhs5EqP3mrSO2RIn2Vtdf52veEP8PvEpwR5GxqzpLCu9+ZOjTWOwpLLH+HczY
x2WX3+qZTMayIZNLV2Zu2snFA5T9bNa4/duv9eXCmGg08vMQivNrvymnlbAPWPWeSXTLFHnqokhI
W7fKZsc2bWMwywfJHGSDFdjQzmEzivCHrLvKmzPuFgAiA6Ll2UapUwL0DDTyeUXwxPkJTnJFK3cD
twb6XC3Tw4zK3amQtGu3//N7xxxBH80VR5k43pgTwUIYU+uFoHGe7mUC3aZcXcjAvwj0qBjQbVZp
h1tyTxqjJy/GZGssiBZ4lzW5iOh057j9+yBoiTngLq1UMpNCPVejZYfBESZJJ2h2CDXzyhf8DQPU
7JLO0MMLCnhiT8v5VQiP/OCcmiltoPVBR1/W9PDhtVpG3y7J231JT7piRP4z5FKLktz23hwHn58V
KFxBG0u/yt3Cs/Ma74x9AlR8ZC2h2Q+OsK6m3JJW3XadlF4emYiO7C5x+PdnNCpbU2JP44qHwrxP
zLPZEAPvwoQQag+WMFLoAL289ysOmu2hjAC4+989Kkq+6kxPLwEVqJfoBQCGxQa8ddxDAOD9/UQB
d+ZN5wZ/Hr0mRFZMDRbdzsaD3LHcE9/T6FBS/ZXdeQjGPT54kQBmmI4rgpJCYx3lJP3A7C9yuzt0
izcgtA0diAWy3kBdhfs2tKKByjOmDDZDYe4rOf00EJyD6vfVKq9+uYKAy5XlUCudVKDJobwbXkXd
r19NV3UjMXfhl6PWIGqw3sikJ/zQB0ar/Fw0ajinarrnFgDRvhpjuTrQ1500+x36f1IgD7xn9fwy
nbfcUCrrFHbEYs8N004gwuH+fmTFqqyKvOvQGQhNIC3+zyByzU6E6rril5BfCuecfncz1BIUpcZ7
sHAH5kgI3gHi8E3ezLai1hSVtLjWOxnCHdc9hXFo67jRshyhh2j2kEPKD39pqxT98sKePoyfCdhv
9GVURnBhbfgMEU6Zmet/9WmqKXCMyzK31lTB5otY3WUjkFykx62Z3d1cc9gZgkr/q1XLydrM8C8k
askyGn9S4bEvy8ZWTO0lQZjftEuw1YcBHQxq8QcTS6lNhPdfH2aUmeCKO59wbNfHIQ3UbTbeqOIu
ArAi6empbCjc6f9YDsuHTrNfAdDSLSt4piKF7n9zme0VhZtvjiLQYkRZKg3Ec08OleIwbw/WjTKq
xcwKhTeJwR7RRHTDPxiZfQzlZ2R/kPGMiY07QhmH1Sh7wmXxD4l+HwNcSgaOjsHILodXHcnFug7C
wBGWq3afdK2RZRCt2luNd6ByevbTOTPLepD+Vmi4mKyUQSvg4xWljH/Gl5LveRzfP7l4slinhhoc
XcBkVe4NpysAO9l7Up6EHpawF82LJQMxrAw7wXoHRmF4DGVafn8fMunzZPPbZKlOyqjh3fvkVm2b
OBmu+gdusBRXQkX0HiCV9sbH8LYpSKTYlpyvkXWH78jlSItiHELncfmLs7WQNkWSWr7QNJ1GOzuJ
TiOd33538DuweK5kLtOvP08sVPDYEWEVdXgfrnSrHKel8NKXFKPNLBll7AeWjK7XtJcDXh02rJYI
twuq91741+XWoLsA9DikiCihzq2kZxvtEciKj5LQAoa6cVtkbiI0h3/4Ta2jLqMCB/ZVjHr/HzE1
1vLdarTOwS6DoO2sdkf+/sGlPWm/Y2fwZNjpaPTjdWh3c8NDgfctrHj65YSUfkhPVIiMjUTDtYDb
dBMcbKZGH9sMktas5Kw754IlEsYHjtuLmGyZ2Zlj1tZcTV7t82zzHzkXc7YbhVTX7lNrArw7zm0b
EyLNU/fkL6r2+Nm0yQ9yBX4bO8gUmYt5CSqqJoh8c0BGK0PZog+3WRNPE7BPz+pRD+ExQ9wYZMa0
n7c9QqqjuTZHrpO4ZYD5DLR1sKihHxcUc+ikMQeyWtPCUH+fdu4It7nKuhwFbZtuE/UIMqPQUeMw
YoPa4CmTdqzz9X40Ubhan6P9Ns1kQEFXnI3wzJ9s8RyTpy2MkKX+XojYX2h8Ji8NS9UGekWCnF5Z
yDI/sEbezu78FrzOLn9L3rW50Fz5M8QvOEq+fuAYtDiVoFWzh9aN5TxwLFNga0BWZ1nxSkDAGoZv
JgsS4zFLEpRrJox7HKDi2S8RsVnWCcPTyqxTxNx8h/FgDo2462nmgojNp9zMRSTZiZWLv3C0bHyP
2OzKHvUICWHq3Qc4azOrgmGhCwKV9xEX0eIdv2BR60qSXQjMCVbvpeD59XGmqocjT1TQsohdFYTB
H/A8XYXyH0CaSMtiokn7r+eemRSmT5ZaHOvldrni3D6ww/H0NCjWsfAbWTk8/YZ4UDhTP08mNSc2
6tWre68te3UWIKlCW+DSna6i0WwH9lJUvyEg3jF24DKWn3r6mvMHhCGB1Q36HdZbcmIBT+4OBb++
1vwbaqosWsCYvYygbDb4ReVHYzpNqQ1WO2e3k4UJaLa8+/RlpLJyJS0TPfxcWMMSwDqHKWAbxAYw
z6mBF5Pqvs4BZrGTo5lUGhbN2Y+SyFTW6AgttgLrUHDYTH3kNxb18fvJsYqFqmCW01x2QadKVymp
atvV4wpPw/I4ABewsoNqIjQkghO7ERn8MEwEJJLrKkiErbR6J2OI+X+TYSNVUyzplP++DPkX25Jw
V0+8DWHWUkZJTOQAlQz/xz1Q9lF3q/hFR76umoQiEWeECyBq1k+WCujWtGGC6XrRzAzVqNRT6YI/
WIwJHagPmXD9mS0oNlOQ3fU0mrYaGDCtVnnSHHACz88uSBxNuvkmEce2Twf9DuVfQNG97W42ZsxA
iG5pJnGYp1LI5Bb1zhABxEU53zyJ7UA60y/R/5VKrekCFVOrVQ2OwIvoqasGhOE/NY6uaeNt/2QJ
M7yyhsJe3Odz+ZaoiOw8O5XEC9EuVKskykUYO08Du9EukkhYikCl64nqgOVnDAFVoupMO2GEWOWm
eGQE24oyuAAOJUQkf/15KUwS4z0l6Z6r+njDjguNB8GWp6wWXslz9UH5nTVn2PCOmoZaCbsNnSrA
lyb0eLwTe469OCvY1amsGvDn5t0li8+viI4McZBqTWpHUP7okyKDGw2ssGKbMwL6Kv6bBlDKxSVD
Y/9ZEX2U2qxfpXbjJOsrPLNny9s+Uj3yWOfD+qpVmR4ZVZDVKOHQxei4KtBNJ0V9roSy/Y8HkLpR
iIwuax1oXGntKe94gXXk/HH0BYUWM7Ppn4acwCwzoU5Z6tjN1xTxm69wDLw3kwDTwPudvmwSep1+
75EFhb78klGJTMwYjOU2Tb1/WuTQzJVPXF59yq0kO+RBH627B3E3G5+IqdYlft/uZ734AP3QKhlk
51WFn1qDrx0/SLdc+KXJRZtJzDeTOwN/WY4Ru0CCjS8mEjENJFm6dMwrLuFwwexi5EL1vS3AFZCg
66GNRs5t/B73uLVRihwhrVnfSxph8BfcckdMlShPPwr8wmWm8ScTzRQI8N+fAz9FqTsstFqyTfeC
lFb2cJ1zPdppR+Enkg8lIO5W6W83gAOYmsXc7Bc4Vr8nEunovLeb4tncnQlu5Yg2ul67+lsZtxWp
8SH85U+1pvoV2EANMfV5EugPelQMcpwsIB4xad/KqfNURiQlWrCmcDPlChhDjL8chR3f2uye3s2+
u1SpQNRz96ppUBFvdfRc/IFjmuo8T7aOpcG6hlq/J+1ura7XREPfrFFovCI4I+ZDGCMIEWJN1eDm
2VQrE9DZ0O9UCeZnjcWpJzHy5XSliXwIPpahV3an+q1NVosCcXi4fMzGXfwQAlwFretLSYzZIkA9
fBItCyisyYRaHWXhvhWyIKqtn/MMq4mvz+QXqFrC8z7WNCTlVwschOqeYgWWzWBNlmYg8d5Xe0u1
guYNSsGwxfx1kEjazF10Atj/wwoc2O2AGZlVGI2tDRj/fllbSWjiZfTe1sP+avYQVgQoyS60WsNE
3d30alfR10jG1fUohIkDAWNArlisS6jAz7xPIq6lGNlYobUC55wu+judIL6lMNMUJh08x0fBMTxh
rC8xg2IPpqZZYvSo3omjWvjzvvz4YPYDGNo8hXU33Mr6MiJwJeKPkXnF55ynxoBMLbwiLZdoC0Rn
l2pxdozPaklogzP71h0e7pGCHKkJPD2Sue8zei+ZrzOEQ6Zz/1bcHsL8Wg7SoW5nzK7rPu0S6R4r
KY7kOZ7rCBoCRbbBhC1+bs7UaXAODALwIgezk4yot62ASaZnHQ8DzVIeCgQIPUgPXBKrHzdWOYOa
vGSbUenEMxREppH9xRChdEsOGbOMwAFZ0xY2R6q284YtasMuxvYBad7q60EuIajMzyuQ3kb8MZwQ
/wBh3vbeqnzHZe7NME5f4E9Ym+UA7Sda1S8zXe5oyw8FoTkBoQlLXDjuQeVhaXa6JAYu7MO1dkY1
XMXXr56ETSuC3XCRIYFxTDzcya2AaVuNL6X8/65Y8O4Qj9iipTvS1PPWuehfzn5Tgz4ncw9X3xi1
K36mvP4KY5lOPmMc4ekT2I+pMEckGSyHS1doIWxceZhg51lE/dp+eGW3xMQ+FlwxgeML8b+mjZsX
RoSn2TliqRa8J0GD4krXxt4uFq7TFlNXPYmsAbPexeqSH+rXRFVpJcfG20dA3N8gJ2ckGsnUsvRO
7eCDWGiwSMprmvPILybl28AxL77lbRp8MgnaJQfSXdua5vh6oHaOsjXMnDW4SQRBUe/1Ija/P7Ry
i4ukx0bMutw9ytVZQRBOZ88xEihYoRS2MCAd9q8bKNz/+WBBsVzQjiwwH5Qq5mNr7q6PO5qCDIhj
aJZkf4AZMrqUxsT9oK3yzlEiZMLFqKLaSzBE3aFxXqPtpDmwRrji8P4QECr3zdAu41YkRCxof7d8
Y59rusdfQDO7dry8o1EBU/5mdR8AVkCvbA6tX0aDzd9fpVrh74Pgc6nr86oP310wK9qEHDVJL9ZV
CrNoBi8OX1uOJPrj++BMNAnx/QHBYr06Lzh5ooz9E4T3qJPKjnrh8dfG92Lt4jLE7HDSQIWjuUkT
e3/IQxs9lopQWMMnNtRXkEri2hIy3Tjoyl2r37L97Edpbaz42vOZJIyBkHoz77y3AxctM3vNHoHr
RldPTIcT/uvRl2KXp+138oldtAqJA3RKL323tj45uk+0teh0ky3UywleZ3s40wwYSY3+2cHlTbqQ
b8d2yZbyRZB9W6eYa+0bQtV5byVLep2UgZ2mkCzw9DOFA+aenTHb2pOCEoSpaKBB6DRe26n0LQ+S
n0pXGMc4JFuxRm6JhuBJD0w6b8Ca3e2vlDZmQGIsvgxRENW1cJDOtcteWw7aEmQOWNAYRtNb6bCY
N0d8kH0iIawZfHYWSpACokki6En7PclbbsdMwHfBIHmgEJ+MXaW80KoHJMdRPrRsdXYCSu/wPIFN
Ow0fbaZLFyfP6K25qWHstJLc/NSGRc1wuxNRlEYPoC/aAx6fk4Gyug7aKxNRkjIIE0WVpM67ipNa
3E/A8tMO2CF3rQwndOHhwQ1LRtPB4DfW03QzAS3YmHEvQuBp6v50eQK8OM2zP7mIZLvHviR6hkJy
Y+qlCQdITWAglH3OeHXrJ05dBhF3xHjyVyi23bTDhNEAfOs0OIh0Pi3QbK4mAW6WoIIjIvPfGSMs
4wj35+W0RYyDqZXRIh0LEuDhSIWvl6Kmvx2XTIBjCUawF6pyJjwADkV3xcKR6ZP0t9gAmxQVAqNH
WxcVLZFRAXpidma5gk4IKIZszEXiwl2NXsOHCYQkz7dtPng2jWYhHw47XA4vamLWjZQaOe9sbLs7
iWtubh04BR13qC/3X1AwV3AaKOCuUYkNFE57KpeId8izXL91jwJeJSbCww+Ka6PRBFbzr2S/MMiJ
IYhW+3lAIea5cdeic21R1btO2xyeQLNWa62tZrobBgP1cSz3k76u9DZW4dOsNnrD2/L542cl+mCF
EeY/he7221CBaEuFaGlxleCtdLIHR1p4s41+bf9kA6bMj6Kax8/N3tfdkOdqIBLJsfCYU5UrkfPA
7bGW+/SBcAh1t8g6Ehj4wWaMH5QCL17QdqVWRxXIZ87NZp29pdHVUkNZORGYzxQSivhyV7r2U4JS
FuWV3iWrwNWnK6zwcB8AFezvYAUS0QF+ETGzrxWBpUiRuWMzmsfo2S9fj02cCNc8zuORW8AHWNJj
ivrMZ0oQaIX75Tn6ii0/+oAZ5NkMYAZWpMnfna/i83XFSeSiSrHpYAm+s0KiabFOIccWjyJqBq5C
eqIfEmP8ch0qbVBxHZ8NPFnTONcZCPX5t7YYnbrdBNX/7fk681ZO47bNV5hPSSXOGWM1HPxaXUFY
FVTo2gy87G7ytOXpnf375OhtgvH9psZAXQlwjX+l5qFLEL0kFls1nv38fo9KFFRHxPcSOv6gCtJ6
uEuzLqtaTsUUtymbVAVIKLF8AZuaIPOtpycvCWylvfZGjkweA3wBQyZY8rXUBKDyTddbYURmP1zp
G+9Lh8MSf8VFnQxnB7LU+MqqkUwWcKTrkZs7wnWfeZK8PxAloV4XGSxO9K9/ZLrwcZMG7A/32HDF
2qp8YSHn9/8COx4TBiLIzF9oNnu1itJa7PiY0IjxK1IGOvUEdAfOm/TaMPd6zvb8NhL6Mlk1ys/M
WuvNsraDiD/BLkezTi4oYfQDFIVHkRRC9SGVSe+Ekv1+kfn1fx1hKjHXvVLOeZz8VzX4KBrLq5iG
0y5lTXePMNr29rn4rzoyxMObNbhTWcbY6vybW0M+QXBoN0CnNhJvXKRu4XGccU2PEh1WlbLcXgkX
djduUYnv3TjkvyrCXoRZhstjr1V3pzIf5WLIqgsADwXFMTGpdXtM27zpdZmen1aoBt7bSlwUDxS8
1bPs308KiGsO5efdmsIF9HrLamcV3AfDrYWr7Im9vYOOPw0hCrhl4+SvwmdqMxfsmtFv5SeK5MFu
IUbmo1URG+TSoDTtnMb0RfiP8xKxK5/2Bc6RikZUy3uFNg/anaKhGV5gi2vbVj+T9vB61HWKDY9Q
KLKZgly6FVO9MzhB7KK31WUT4sPzrGYqhtwXS4mFIQ+OvpumQjeQJqGg8z77qXd7yeJDMa8VYmuf
hd0vnFUdQsl9dTyQxNGINRXtljmla6qwSz6b6P0J4GkK3h4VUWk+/CPO7R/krYsrNFN2AwvRu9hz
+PpBnSFCqtODxy9cr1tlcUyfdy8ht8+x0zD6PX5Y6n1QMqfx8/4SrMy3zzd4i9voB+uY6qamcoe9
ocLcnY6A+6ODgCKIbFfb0M4WVY5N//O2PpJyeAFb2mZ2tZt8XzVNLPCE4M0FZurSERAH/Et572JX
723IHJD2xEHeKHDsa8wqIGmBkHbEqg7VKDY7ggH4no7jgw31AbVFFgkpAyt0EnTZ/wb4xevOjDdv
CoMLyFK5mXeJ+Qh6CGUzIVWhB+RrooVD/lRHHNWtUcl6Dj1ei4dWeszlUxmA08RbhVTR3PLwUp8M
fJyExcEC3ODCjRqkwGsfAfBSYUblebhrzoCDhwpZ+yjEeH7GikxBykKHakskbs+civ1/Z0MSlBLZ
RVSAQjDQN5VQ6FFIxsFpPA5WyTcZiMFK9KSK/0jB3a9nTMP7mfoNkMUQaiBDDNS00LqfzGd9/Iom
rMGHu+ok1gB6vr21JQsOTBy89pyJOu+7NH/XX8wTh+reDzgd6BUWNpx3XoHVPBfRWdtgTb7W6cxM
jS/9/5Og4aJPiM+Z3ie/fU785ZvG2No9lv/WGlgZqSEmi760VGeNdd+WrUng4JvVietrNCnR7kEF
lrLOjT2BL4sgh4jSosuiUfMzlcfF58RKnFTsdqRxpFopw36w6uotTLSLWJwzB4EF21VsF2oWyTHF
3PChM9zeLnNv5Jhi43nCK3caPh4IdOouE66nZDE3s14r7wH4KViRsu+8aJh3Om35UsomFzuA6pFX
DxZN/bSxRI8Wz5lC+TpKnt9YTFGAVMV+n+jSDJ8miwWCe/L7c/M6QyEIgCz3DPO2isdvblDz5Mn4
6bBnmn9c4ijsc1d00DCrz/UJOgzMkkwT/p4nzSi6/vL+ICOCGWFRB1cvSijVPQmACjtPpbVAi2yh
wbU2ZpYFCuVeGupu1DEQ2FNbdWgD1zQSdzuCUcqoO9hppKfFnfgCC3Qgt9h8gHTsQ/kG+x5kXcVf
yfeNU7fl7tFurk7YrDB/ohHxSEMiXMRWrc34mjHx/XqcjDwO0DhtW1ZOfcXic5C3u9H+WLDr4LQ1
6ZsCF16b8VqFJTFL35weC5Ld02F8miM94iVsvPNKUtOy3WI09ndCB5OVRvZYLNP0hjxMqoJdls9k
oYnbPLeQwOR7aV5T38eJuG92f94ARtm8MUiEFmKAqLdUSphF58fwzKq/ZLBF4L2yQur3IRJojUnC
+T+o3NncTsA/fsHwBkFkd3u59AVaR1t8KH+XGn2XpQj2vfCLgE+HivY0zxZWGbOgq2kx2gKxeZc7
RwuHcn048fGUIS6FT+jDfjglM5z7SIYJ5XwX290iv8vmOjMPhvjyOzuGzVOrQT1GT4kX2GJBZoVm
QtsIYZLme6QOTLM/9pL7n19a9USX/2YZ7XKWafX3Omujd9FNQe47I0dfiQHmG7rL/iSCrmOQ8fd3
aETf0JNjxOe76DtPGYGi2qlFEPgfvbZJbUa6f0BW4oXSP2lZ3JMbzwN+daJlZh8vBOHX0cD6qJU7
1Jj68xxTz6sx2rKg21RtUKG+EFA/EMa9pog5PwM1teJZ6RPAvKINfCZpZogd/3NZemlO2sF0c7Nt
L+1W1ESn9sUw1w4YPB3rvfN7vWpk+nMPU/Y77wWPhEJDulfOWK8pdkV6rAEcgla3TpP5ET/qb0wk
+l2iK0HkpVzb5J8OkxrUsiXE9T++MBRvQqtJf606W9ONFjeUQVuab+NDzMcz96BAfyThJ5KYeJyd
jaPoTCFqHh1OzHWjpYNI7jw7ajypxjHFfScbCYLNj/srbKI4SOkZXHNPFROaLLK+sZ4scdQXfxJs
mY3rJPjwGI21bm71DxHP+h7Pi8W6nupvn6Q/QFIRyyD5JSdXLnTtGRBl/DuYzlQtxjpU796ZChTE
imXkbfHSUbLLx7Ka1tQKCWdiur0KFs6DTI/Jxsx0wkYuykU2lEuFDygEq2+ytIFuUEGdVoXUoKfc
eWYwGvF9uGl4UaIMna0ZAH48baud4Tg1jWNRPHFMguuJ6nG7f6Gp9xxyQVdIJ01dwMjcAq4KP8Tl
mXsTeIxinNczRN2xMPC1nZlY3U5+FV4GcwucKkp3CgG0KReOTSbeyasgq++BiLXkUhAZm1D1kdU6
/Qz+0qUt2zR5F6oIzZ9PaLllL5bu+YuyAQ5m3dkHuHmbHqrMH61N6RI32IELFbrqQfXLmD/lCy3O
nrP9EkJCZxG2qVwJm3+XjUwnTCZlcCSNEU1vgmc58S17Hl7yWvmvfNRzX0yNAOaS+9c7CWITjMO1
2LiGiNQatQC7XTZ8ATqSfTHJiHKdbTm4WuD4XWS/KFoBdGD6i2Hw/YxEp1MLjvraaW2kzPGsQ0Y8
rnGpPMJkZtUV0E07b2AT9SRJQc15k2XzxdllCftBZakwFZSUlwpU0i8S9p36ymzJUbH86zxW7KT9
HMYLmjNQ//5dtc0zYdPYttDC1XOsGNzWSFCa8Y/dh+5+rSDdvgWqb6sDXwenA3YZiWm3onXQM2EO
OFP2P7+VRTHvmYzFM2B7nLo20PV1p0q7FSi29t8AfCId9wh3A5ocTIWv2rhdPluXoYJ5DMVZOOir
m7t9r/5SVenPElrJyAXqW/wBaQGjAme0xgMqNKm0vf7kMnHPAlNlee/PPiTTGClE6EihA7G2rlff
vUL7JuFUbFtiJ5qz7soX6tQ6AjP5zjE7qUmthgIpuavsx2jqu4L98tsyimWByrQFioXOxgXj4vkV
Vf1ZmycoCnzHWamp4sNSv4fJm0RKoxw3Rydajgp/bm9lYkkltXkIqMmb6+B80hUhbQlOZotMDfVq
C0syVSHWg/DCCnFkZ1U/ox77kNSe4h6T81ori/0612KvAVQGSFiRhx6T/G7uWdUVSYlHsoIc8XMR
q0DYLrIAUjMP+CVuMkA/DOsmCnMVW7TQRhjxEG/GwahfEo4GZZbureQKxuOdER2wZwChFbetbFgP
qV09oMUHlJG6iOaLyVbEREuf3SKCA4b1fTKCPwis2XT/lUDxjWnqs8pWryITjtpJJPaBXm4CiCup
+uHF+Y2mdn/yI5kC6ZRSlbOes6yieuNQJoH6oZmrbeF6zBfDAjf0Ka/L4tgVTxwJ3Huq4oS6erqa
UI41Ho1c3rkB9KhJxtVWVRvte2T4ZQi7Wt5XKdtjAvHeoTDYuJvomRiC3MR3zBsEKEseI2/fZQIy
vWndmfSolRZm/U5iqE22JExuRDzXcjVKX9cWQl478nvme8Dwug0NOj+fNfku7KhSl6gw5nTKg3kh
qlFVmz2S1SXpT80Yiy7Z7pCXpDCzvg5bXFfueL2Kll4hJ9XAEYx5qYxNW+MW64uaaOQQFpxJWTvF
spTuIa460U0iycwHGx40NNgYlu+Wz+7tPapRxo2ebtQZ5n4lQLHshPxiDO2LDfqy96V0JlyNXUgs
ca/MwzzqTI7cSEwMghU0iimYyiT88PYJgxSH31whzViyV2C+VXVFRG2JetbKFhKFh6svOBIEvxF5
dYt+3PYIBazdEh8ojmB6naRjDaNJuDu1HKpcJ2VKTzo/fiVlhL5oupApTlOAeVjNGfx/rOV2P5Lg
cE7pX4x16we82eE1gxc61ZZxKXsyEog0ruKscdjwDOZYmkNozy2u23n78NAKBDaMKRx8jeY3aTBV
fD8Cu2NwzAAwBTxxUrTCZchstaTZZ9/wNF1q/wsJcabP2uPyrVVmQGIk5OCrtFO/KvbyLDsKVax2
mrewagdAQrs/ybTWZ16F2sqerUgK98NEMvZ6pPcwBfygSmQ1TVRku6QL2ivlW9ZXxrkLPixqE+ty
0Et8d9aicmEBBQp8JedQsRb2f9bjSYO+ou4P483VQ19y4GurGpW9t+whmHPWrilbKDvpdJxZeVl5
w9Q4vR0jILYhoaJ50KQoqAKC+T+WkW9mJUe845reHirRtAipOO8Syfmye13EP8TeJbZ6IQcksIB9
u8gKwQR1S+8173cSaK0O6yI8Egeuxok5WJ9inFRkEf2jottxJKpUeF7hZ0yxGmrafbux41qQuxJD
/ASIcbwpIOqNYSbjMo1irE79kAJIvGhQtPhAQPF0BiNOpO8OlpTyfReLrtdrvSLOI/OR78iDONX0
5VAqLlVc7yEPo64dlmPdxh0DDKReBJdj8hENKjj+uRs9QzI3SmvirLfgM+DdrFKx9Swnb9WIXMpT
jsqHyqCGy6w/fR5QZ8sGk5nnj6GzECJRjmRMUWZ9bkbAoWSNI4d2B9pDPhKPEVwU0r0u5JMidsrU
YAFaxDc0cwHdPhgnIsu1JR7IPTaMn5qUnT0TujRQQQTiTIAe9pPWr48V9fQBXmAy5wh7jgv1Ykdk
aGZ5pY5dqj0aqgK2ke90XnwPjQT5CoxM/fn6iF4c8nZKoh6Xh3WaiY6GpPa+xaf5bXSQKqB/sD1d
kDRGRy2z/k+krn3IQUl2RH35SUU1yw2/fAjSKufyc0wtbEugFHAhdTD3HB0PWIWB+0FgzeYuKuHl
d5D0d/B3rp8SPqj1hwqSo7q1MSBHuZJZbQS+Pl5ii4+ITgRTGjYoCUsPZA4I6PFi6+osJTMCrtta
dFXdvqGr0oi+ETbJLpk7thZ75Qf8A/La7nQVb7p9sZjini+JtxGyDkwa+ZbHgFlhzQ+EmtKa9Lkp
wWa5EJTDC53oVhnh+dlVL2DinNNxbpd8JV+3Iii15HwSo6iKpnOrmyuR+S9XDAWNaOPBTUMzy/e2
6juTviAVE1SUt2yQoH6bRpQmcQK3CKgukPrBJDOX2isF9Ba8xj/sowuZGsQD0dr6wROpQSkSPrlZ
B+2kBRMZyC/rKnV1Bndvx+SnITXTRFbNPqRj1b0UKVLNuQDpjF3MDWPY3wAtiKrkJT2/7DDaH/7c
JCmoU00MCEgBzFO39o05tyMHYQMiyuRzvKZetuJcexLHAuu6on154PCN8aiAaHHhrAk0ERItqDO0
TTHq2EKslebIciKSMjJHq5VXlYZ20VS92Tjlk9qzqmKOpvsb+NYsi6Fr+esBUCkRKt2TEgEdyEGf
Spa9/Umv6ebeX06Ozkk/NrfalXhr6lRQnyuSoVCHzajhjgR+YBsh2ZuYpH5WAJFJFDP8yUG2DTyZ
w5odUpSTJlD6jsg/e/FztJceX2az2I5S2fiNeO0WUTlnMJnAz3RWE+K0PDCco+CT+wQFBonymJNM
jI6w7KtD+f13NP4SV2Sr5vDrc0Xth4WKNw90O5USxQ8srdV8Ilwkmx1HcTL2MqarytCjdez7AYPq
734ykG4DtMoUCFrjYjcol5AlaoVkiOeLHdkVJfaB2btzALWrIEThELwC1g06QEjB8mVuyIXqXFSu
EIWpCS5Gi0hlm3MxgLxmreELmEMX1sw7RB6tKKCa4a/3yKU3fP61CGvBqJon5qoVkP6g5deLGXBI
twI6WX6cvBc6kNvg+rOpYs8o/2O4ET9nxir0yJpxIuME8crSXEoo8UQ6xedd0g9qTSxFfrZeq0xC
rfUr/co78xJKLPwrl6azq5TaQhYl91ApJtwSo4G/vwrCF2NdAcWwwCOC1Vl2FUDPZtGDIKdlVdvN
zYcDyC1hE61GWX76Bj8W3o8uR3lYH/wjRzm8ozgNzrcIT93D0IWwu5qKFugxYHxA7SOuvLTtuKZ5
1fBoCvCUSr4L8XoiHVzx/3D0cKcmKkAG26Gj/tmxPwcjk1x66WhvMpLougVfPS/VbfcPDWLFYWaP
BPt9vnF87UV39uFdbiaLuMJnDtZHCBeuuOu0n1amcbZ6X/gdgXWjuTzKgVMsajQoGr4vRihMam+a
GyVfZUTAv9XH1WUGEobaQ9t4Y5BpbVX39khgVQsBuoQFa2zlGD968YHOK/sKeLbqybES1aiiZB67
hrNQMNwZenKauBCa5LMXJEd9icLNOHWGNk563keITQaL4nYWnBBHF1RLcCEFXNpH1RvgoQi7Y8MA
gL5pjALIl9LchLHJvJwrVN9l2izLAKg4VY5SH8Fks9I00ihTkEbTzpHePRJeyZN9AGRYsj1ZytzS
gbF8JVH/xm/0iRdIaVdjqRrWEdM5Mj4H5xvkyAymxU37K25k4FQuGD7JwWgwcpgZ+1MLfClLLZx6
nxK02ecJvNgnRYnZSA9ZIRPXh+bb95usQBmhaNt7Fu5qsjYDEX6qXbMFpQLX+z9EjP81XNfnC956
qwYkthBT/Xop1ntxgBb4JMU08DduAoEEk2OjllQMElF5Kkkq45dNXwvDVB0wIwiX35q/WUyLHxdJ
0NxCGF9BhllyLTOtA/4BVkVnp83biBmFLm1EruDuCVwua/D17cyxcP7ug7O68HMF5ills1K7Gf4D
4Y7XQCPbDJT9i+pzghV1nfajyrNXRQ7/hns89THNrlXBId3Ccf6RajA7GBgP4VvuiiF2ZLrftEBL
a/vrcE78a0uTRU8VVH+TxjBMVvJCxxgu9U5VsZ4B3Gdgb0ciONRh3XTYX4H8UOlSD9m6gK02zR6u
VCIW2kgiHUwvIuEY069GgbBnQNfydKTwZ5snisDEERRlujMEW27UtMGirvRP1y3yqG9XE4fa9z/u
s1HIXRhwPzL1LX3eKUNFXNs0IHL9TeWZCGvkJfDUMt3IjkZuCgbdEcZ8GY6ngWHXEww1S6JvF66f
LxzRTJ553nyVV6pYQZSRcA8v03c+jZZ5QBL1uYpp796WlT9OijH0w8G/FTsJ4RveFM+fRgFJCLZk
IRvsqHhjIfTgb32czbMVGRa+RyFk16B1QIQ444C5jNhLurXP2gbXJu6toFprbXAYy4FIzCZketS6
bu1Xqg7C8Hh2kVxtZjrNyglKMeIshe8F/RPETAT0YWJmvJEy75BfjiMVPu/Hh8q2Y4w/snFKMRzu
JWD508FF2BZ/CIo0XRRR0EslW4voNUDr/D0w4xLFdYuGMpnWoRthDONEE1mYYyWcwTE5rlnuGlcQ
5TdZF72xkN+7qOKtTda3RmWjjCJcocgXEa8I0IEKrPHVgvpu+ED3z6G1R1nXz4C1jzXtRtebt/+j
9q7z89RS9fS2T8ojMmAExuEK2P22kiiMTpHIAplR5XWSpzWfR8jefAUIuiDiNf6n7DblLwJ2D7Wp
S+nVoaOZmrr+xC0skkljxlSvF51EMXLN9eErjMONwWSc33dQaVboZlQBfUpV3l1/s/0FgJqmZ7xR
VPgsq68+hqY0s2NRaIVi0WOEncFTQBK3oF/VX6qSY7NE+/R78lwRAoXaxPEB3Aw1THuuqRymubRx
PLEMR8qLRyp8294vh0VtKo5l9KzdmhMShzycdmo27EeiG9cgHWO9AkqNnkCddJtZmyW4OKSm2xZ4
bNMuJfwPnPzTA+Zmh5ysVvgEbbopCGtaeAxLgxw05I8+rU6SqBKO2eNgXBgDXSMhH4RheahAM8AU
cZv95fL+CL4s+2ALiwDb3mUwv6fPIyxSfTPudDg9RuFTrkPxTDnsGHrz4gFb3mBzFZzVboPlk1sB
krn7CrfKfYiQ9pwIKVFRWfald6ahkiXRENW5Ay/Xrc6YX1j6DvOLa/wgd/uTgV7c0ygcauvyKkUN
L2a9O9kvMbprxqYZydB6Ipg6CkhRWSs5uECSJ2Oq+iX3LjWu8iPIb0zTesx7JGcs7w2QIjenSlCR
yjPb+Wg7jaT3BeOZTbItmPuCo7tGL0HGIO4ZmXKwBpsf3Vr5bLpgGN9pl5E1naIKR/OfusweRz4E
UiqHy5vZl02wcadMyb6fopbIVgmxOhrb7UDDVqMVfjMg6NAxFfAS2bTBOhxfd4FCf0LWJmYMUD3O
2j4uOGrdbe8O+7MLMzrFrm2qM2m4cqYd1Rx5Y4TvW+0NWDABBXI7pdVyxxkGdjEpPV0jdEK6X7H6
mEvSU1pmMk9+Z0Ckyk2/oT5jODg7S0rc00oK2oJdUiF48JwZ1rmAGUL+5D10Dpc4t2ltxaRX3ejp
Q34ifLrUIaAZjgIy0ID77MG0Nisek2FcNhTcPrzAexpAGyKr2sl5t9+wWTu5KWK8Rat78E1YqlPL
cmqBTeJu0v5mB0gHZ5zpnr+zashJK8FgokYLczU40UqxPdY6+SgkMn8OBtWz8bUrMvmAFzqtpKWd
4NqkUj1mkx5q9yTFCdvmJdihF9Z3LOKN8h6OhoXJY8+CgIbuExdMxvs405UTjIKTVenoqj99KLad
svJHsF4H30N6lJ7hxwoneXy/IqIihZyfU/iPFQFdZTY1EdWi1YyCxrGoHRiU5a/a0/dtIbFWy66E
G3j/eqYqp+5Awx6rEW67dsMGJ4/txMH5J1xu1fD+g+ElAVrXMcZfxjPQ4spuxp797xEfJ+bXvNNK
7fLVJdwL0wl1btdbmObnUgmQAgEwA4CKY9BnwipBLKeg0eOfqFu+k55QpnUJzZbL95R5SoLLr1vQ
3HEPhx+CFtgS7Gt4ethm5lHoZWg/UF8bmVHKA6zCzbnrddNgsnw+Y1kJCbofLcc0WrDnZqyam2q5
1jfbqxcViZ8EFAl5sidRwkqw++2/Ydta7Lrn3TuWzGVcJbK7K4LsovQcLmDyi/bjqpScTE9m4VuF
vvXUYxxNYTNxphaVQiLShG28HRV3yMuODhfHKJpRbsiNriIK6dwHHbyjSvjThgJ6/LXuOt4XnPP/
cT4W8zTWuPavP4Fc/Js3vMwpB9jYACCHIvnP+rbhRcrv6C2SW48/L2kI/1NioilnRkKFlBqGt/No
hEHkpTpnGIoHAVJCDVmWMKqRe/zvKfPBFS0GUYQPA7q/6P9YPRufhaEwLV/D31zhlfwbpVqxsN8U
OUP8gcxHhzWmitLK6Tz30hZcBIovMYTDgKXXhSvs6yj8JSr4yxQ5xrAM4MDPpfKf+e3f+Sn8SNf8
+I4v5CRNWtvIjt3y/Bg5s0UHZLphwzkMJQCxx8vDPLzCpazYbbHj4sKZrUk1mD7xmvbT+7mU/4M5
0sCR4Wq8lP8XuDKBp9sLJmZLKu2WN25mXvjarajjA8auMwdF2vEhRub2HXCVbNix0a3n9H5AihZO
Y425RFM8Zzh70Iti7LnszMKx5fBBQJ4zC6TvHPO0y+zKsW3IRpZPL953XpDSyq7a/XIqigSsmnDf
UuZDr8cQtSEzKrRxl1SRtUzbQms5uhl7ZTZ+JC4C69qt9EAuDkGA4nMy6Pg6degMfWZ8pe+/SGxK
66WJmXJbeurQP4sagUh0xQqKzCHNzH/5S3m/g3AFJlbFRdpRm1s6AgPmrWYTay5U0W035IaGaEaY
NUmsoJFYAIkD9h70dZr1W/x2UeewFNPAlC6drnnkGiLdM9+TDFrqzks8SxLHJd1l5vMfmqhgE+dU
6Xxym6kLld0/haMy7atVKZ9aQ48CUr4Ai/OpJ0mUs6JodOuO6a7WuAiNrlrgTJAS96+N8paIe3uR
UsKZtSTbRSUrjlZgfAxVF0HataJFg1r7n2Hw86lQXeNVRQAu826qfBGhyYqKaJUlE4hybYDwVQCP
nsKlY5ZfVbWWj1bqkAfrTFvqP7vEaGb8K9Iw5US4ljJrzEm4eN3oJPAlQ4vgJd4ugdW60MiuTx40
L+HY0ghuyOKEw2D6NPTduuPM+IDUXs7JxOXiiAmRdgmHqJwO/DmlQf4vnhkS0HRJbUdo0a0ItII+
PO3SoPqz8XFA4fjd9VMtvd+wZLC6NOr4RKiHoERLsu9W7n8kLdRhCC5EjAEMtj+nJIRAycO9dEP+
ceid4pCfqxAVMhG/oH6xU9636uAJsPRxWosennjWiH2ePDb0kN315/SGXYtzSyTpTyb1A13ZaNN4
vM4r8d2ReYV4v9B1lMtADmv4e97Gova0GWSTnOKzf4WD3+W+qoQfzO75c4dtPXmZ6uy3Jow2bGKy
rW9H9fPi+QQw85PuGtpgMVEAeF1uCSOuZFrFXY8m3Fnt0hX9Tj8YEuDypPKcMIV6z7dZO2PSEAUW
iugXYPp30qj9duvLHZVm2pFtWKjesMDLDe3utjbCFPXGNIFheV8lo0MhjFA+rXfeAXpugaFYDFZQ
Sj9rV1hQVeZg3/N7y/R+g2mMW1fTAgPQwI8oocCGzPKqxw/87moEOL7JOlsl3e4PcBzEiZUFII9u
+2YKMTUWGqPK0AeBP9TcdTl6fizdgZ2rbZjyKte9TNbPkAuiG6DHxfEmMol77p26RlfTtIQ/Q0gF
e2N6Sn0DiYmESc46rG6TWj/JOYbbLsXIoBMeS/KestUwszkjQR+e/2P2/F4WueJIWi41ipVtWUuX
V2+6INwJfkbUnVJYQsBixyGJxSmdEPCV+Xa2BlF7qgXm/jIBAkgneLuc0q5DIs4TCsbVMqBEpRMT
4rI1kFQaXTTEnW4KKvuJYAcC0tDTwHwRf6IS6S4YiZ4abvKsFzbEQ8RdbTumsIHT6d97cw+Jl0V/
9Zv3CHasZBKo6DvHPGyUBEuQoS+eM4bO9D9ULolV9Hi6qEbyktZnivTv78i6OQ47hgf7cx6okAX7
c/nZ9qSK5fIvJv4dT1hMdv/iA7Jra0C62tHQ87riFasx17ak7iuRiaDcuTww4HyD3mHB/WTDNhCK
Lf44QOd2P4gil7f8eUg9ikscoyXnS8vy7EieRPuBwtRCyUs0Kzp8g5uoT9gPPeGjuegpwMhCRwQg
um9b4EHsOhhEeXDq8WG9q1AcpaGS1hmZ5jGP/L7kEW6S3NtvgndCPO4SW6eshEFAnbVGlehMzVZy
iPRS/JZnGe0mKLA32oyul32eb6nCod4SFYb797f2Z2EFudreGil7sa9w/G4L9dSuFkuE813I9hCD
3A+TbWczBAQefzuR+4nwTaqFBIR1NTbhS9EKTGsuHWDui5jv1i0rZP9Z3Ld4kxKH43cJ/1USmI7C
0rg5GVyQc/FnOmRW1BYL3j29Qy7W4XnF74La3qM3QU0VoHw+D5luCBVdnm1AKYzUxpQ5SK955S5W
keNRa63X2NCoTPUx58wg8Ux8sJ25dvZ02pA+oANvyAFxeyn7bi9AoywRgobFzF/9W9t6KOeTiFK/
M80+ftaPdScgC4Xz0NxbEZaIvE7qNXd1A0RukfP1BtdV0zg4Auu9baL6cjcS1x4MciJJu6mb3uue
tvaVRRVyHuh8V12G0YLaoUEJYAcgbx7OMKqzrGYO3l0N9pP1Ab7VC9MEVbtgQWCnHSvdndU+mq+a
WTCnoikftj9fTnA8A6eoS5sXTWC3fNClasoIh3QLf5EE4V01aVNUMmZgxjheqZsdLAHULjgczKi+
nG01CLouUZV7oKoATTrA/IHgBGMvLfqe7e+mZfrpEKSqncujLn2QW8urvD6iIsMezcp90l0+ziRf
OoR61OHZs27nA5PWEtSPaqB3QFZ0RfqwbDM3VqORZbbrhSAz5blR6BzQ7PQmuiF+JMsdTJsXvWhz
4MnTaK7SLuyYfXmRHOFugwbkpRTGoEPbrLycSEBFoKtak+NLwVFTfmMPTU6NSVsZBIDwk6AF3o6v
u0PxIG1gBxIvGR1l4S/r/GbThQquueF3Q1P2JEhXpXW7wq1AoEx3bxFLs1AHb+mYFLA3XTK+5jAm
rGYTOI7IbOLj6fqhZyhbBWD/Q31hr5nVhLHffyYtKPurQ4AaGa8I7rFv5wry6L6Cr+MVBnZ3BCPL
ITab2M3ZG9iezmdLHSJKFlARzuQ+MyFRKmbp7lBH5qF47TJzSN3j0Uz//A7EBQOHIE8ehoFWm9Q0
8Lsf/MGdJ5ccEOczWC6LfOR25QYrZ3cvLQqAfLhuO69/tnu9oTuuToSd0KKsTNSuS5hJqXdphYTl
9Kx7rBZFUhl9ZIY6bhn9Ejn7JTuy/aaN+GnBV9s5KMAmLc0cqz0Yrc7PG97qebbdCHNMVKmO7ohm
ss5XqkKsmsIPfNjyh76NlTzwuDW5Xw9oZ5vnIFAolgteW3NB5wGUn9Kl7UY6SRsgwvHIFQ24xtyl
5LF2iHuhQb7KLdpTGm0iUL2gNxLIlSeCu5gAzb2QKkg/0ckwmkSIMmcEody9W5q9PZuvTJFVZO5/
x0qlnaJRzz628r5LvU1IlyQEeYyi5LitbbnbQH4ndd4zdBy/Qr/EMRtO7NGeVLHluTVZaGHkmfsX
Yu4rsoD22iCXGhvsQPhEeTVEgnjwqWFx1hTzzUmXRTGXNH7nSBRGyKnDA1y8yvO5s8+8ckFnQy69
glq9fNuQWxfP00zkVTn8h28CzGH5rQo7eKDshQ6rG/o7AZjyF5cR6dwLu2cyj9g3+wP+e6Ptpulj
FcV3YRIkpr7csFaJ4bp/X5FioNL4mFPXTGbYyr5tb/5P7Tcf1OfZZ9pJq1HmJKHDHPXR/m8T+ajJ
vAspAbBCsJyoqrSlxbD3oXyMsqQ4EqTqcGsRFy4XdkWWvSFzH0ejbXSe31PyIiNrI6GyCW+9Fp4t
jiMJZx/nkJmlox8jq7ShpCe5VC96SuBgR+py6LQHzUVu/fRkx4KD2wGfXEQVEr1YqPjTWmAM9zSY
8x28/oHdU8vuTkdKZEui2CJIFWQoL99W8k+XetsSx+BmGSm+2iyse+8ziHb6XksB3dwikhoCLrg7
D4XUf9+Wrwe0AajhnfzLFk+f59f3szsF+3LV1NhvL6RJy1ZrXG708Ojoz+6VTVo9Eg/1RajCuPsP
UYjEHOoffcGKCNzXdsSXCwdRufUcPukGIQ0cZeHA2FzPgwdAaJWuoMWQeatkD3mlos+4cxlTei7V
UFynt77tnZpyp5eJsfS0RENAcpHwlcPx+7YIwjOnCt//aicTc2Ds7tw9gN1vTmdFKQuSd11mwbxs
oILQsxuhKq2WsbwPSzX9qsBLTqRddyCKdte2fXlaw1YdpXEmcv87cNerzNO2EVXYarcaeoHqNik6
xKUTWeiySpQn2K4ygDetMcDo1srXvuWvmw847nkJMIfFCbTafFLSmWMcZxvK4RnYvi4iRoZcfVN7
FOThHMVSqIhN7tXXsKXpB0oP2GWtzCbAeNnve28xH1kepJ48722FU1dqBcVPqWKcRQfWkd8CPSvf
+Cqa1xV8L17Wn4Xq4TEF+aKYzoOyVm5gADbLw+ou868K8D5yBg+RrlIzblXRTGHKuzWLmrOOR9FJ
MKpe6dAxcOYmfHK/lpT+oc+7xl6NMBAGy0QTph3jV/ywGgLDjHY+MQVQFTZApUOqqiknMBKkAEVx
2QK51GbrpRKo+yKYgrEGnZeQ6bgOfL78Ysf4+GwZnJO10DJTxNztQFZvsILp3YDLf5KzZWqdSTHr
QFv+WyF4YCVukxjXyqkv6N6LEE332uIhoi0YSqLlqtol0ZX1h+3nvTyDweJWDdsRQKIsncZD5EaT
1nV57YSz3Krm7XtOU3+QG75mham/bAt0bsLd45vMkU2iBkJ17dvs2e0Q0TXLgFxz9FkdLDSZ1OTw
nLGHwOpW8iWjUP7yF3ftUUzVG9p+nE3i9Shy5phYaXsWJ9sjP/BFZ2sTBb+mPL0MIPs0bQNqqO9O
pnIBNXfeVlVKxtkONinN5DTIDgILnZTiz0MnTpndry+URxSwv+Bjex39FPbIDI+t1nXKhe2LPf3G
j17nvGu9iFMgh9PkDcavJvm5S7OTuYMEXSnhSb6SlyvFPVl4qeo1qj13lUY02fgH2/uIlAIaliQS
47amPVaBHkpxF8kRT6V0cv/pPwk+vLpm3/0FRoIWd+SG6HZKiq/Eqe5BjocvSP9d/TjYxMLXBHnr
ZVAW9h10s7qiIeIjfslBSBHPpN6HmMjLVSJw31ij1IRHEPTxfUNxhk/TVlZc9X1uIB+awWAIC6ad
0gu7BZk8s0oin7QxNeD/yFJZhMz4SVjTX82tmDA0BDZ/3Q5VVndPvOZ+AoYSBkX1Js4ZCqscyJOk
NWmmC4nED8UYGdRT2MPUzvJjxR1HHM9tXkNIYJtaqcuN5qJpzRL0SwhSkKEZNdp9T9t8+4ko5FFY
5i7Niy2HUQZDuA8No3z+sBxWZq4aZwih1anM7jRj1yQZDj43pKSsmjMKjyXY2TW5Ud1j4HEW08uG
paxKi2IG9zF4qJiSi/20erPjfevbRl3lYy0d9Z4ENFcOuipd+DU3pd/60n7hdfSx9LnwGqXo35wk
XbHQ8H8f+3VNzJ4rQD8tRQgS6FM+TBfXAkVPXI/2E+uY5B1SyTSaXTeYCPqHI4+GbQehytKsj/36
ClfKscsT8pmtJvVvv3+y2z1n9mzVNxh/O6RqxMJU74KC9Hc1lvqOEB1fBcC0WyVDStvnwK4tdbTw
9f/gtuZdOEu1AlfYyMWSES6EtUr9JcoQ4YjX2n6eGp5fOIkfS/VkH12q6SATUzKti+JjyCFoT2T+
fQDCVqquuKfVwDurgbdrOytkanFdGlugIWjfbhrKyureenMBqp4Sarh9wDlQHHczAfmTbF3rveKh
IYwunpRXGilYKzLu+pPSsg/2UC1khA6wHXhUvtAit3YBi23le/4Ws2m2mK4m9d1Fk/1ox4uQl/eI
SrEu2a+PeXXtYZZ9sJvL8Ef1BQdLuGnA9V5vV4ilEXBAKnEKRyeQhoNtqhlQTPC1/nqAURTVI4LQ
gZJkrM03xNiVaerqo/ybggLeH898H8T0yb7BZ+lCSPqWjS3d+rSyTpa2NBOW0OadKp6wg/YdSYQI
KOIwNcV66M/gIGY8/xi4L/5Az7UJjIgQgfuubo8SapCkCppV/wzml0h7asVZT+QJ5UcHoJHIA9UL
gYUhjt97mJfCpjBw+vFz4r79eYn1gwbHsZ8Tr6l2q0z6bNU+hC/ZJz8UJKjKi2yK/IPs/tlpk5FR
mHd88xMKCd+SLuKNlCwmR169HNpCFeXylj/u60Omgm8qCjKWv8NqzPOMFQWvWmgkKEkCdUiUegVq
siQB9+wSj+D2kWYOFgBnKZvKeltSfUS8aPvTDxSCgWBUiCUiJyh/MNgGTKGX18292pU02x9gHzhT
LzLh2HSN8Uixo8yzKp7UY1cR6g7Ld132PLGLUObg8cdloNLwaJDFYWPRcL900KJsizxm8QlpRD8X
4YoRc3iK/v1Jjkc883if9JVoPjnMJzjEsn7P53gJ570sD681DEuLRZwq80XCRdLHhH6J5vmwhxG4
cEvPUfLVpa/Cqy4JdLo6LVyT67GEtBPqh8WVXs+VZXl8O+vd5A6o2LmrRX7ianhBWNgABGGqbiLv
TKmotmxuD0ro8yXdPp67tAUMKkuGdMVQBFDl30bJtU6clPUhyS125kYu8VrX/hEKq6sfFnaswEL5
PcfzWl6Z8wQexYzlWKyxUPss8qojdUZxf3d8nCLeiPhTQfYG6DZG1G2vJW3uEYmuuxLbNr435xYW
VgjbUYLf6Q4wAtuRLCnsU6FtKo0Be+5uTp09l3FouO9Vwl+xgNXfOhnd41kL3S7XZFAOZBX49fyz
NWy5KYnZJVgGkIGWBNAH+BNBqR/+NAMsBbvzTu7eiiw8/7C+HHISRI5S/HBhZKrvM7SavXgXfVcK
1CYTTEc+htu4Zhrzw8KdJYN1ZhGqpmoxSnBU3/LcVyk76MIaR3qaV7ieBlsUHiA523aeF65r95VT
h3M5WYLxesCZFmNToQsGSg9Y7Hk3yn/tqFGmj6jhBEOELzuoMs70BU7Yay2Odq6o3c3LksOt8Jd8
T5FZjDM6azSDwdhrZdX8tq40THirNXWwJ85HUEc5OJp1DzBA6HXKm9N41ixt9L1Fmf/Z+eGsa/E9
UmXonn+pHK6nuF8hh0rNtsPcaf6ryRDH4B/P6l7LniGG8uUKrZN8HiMy50RYHO2gLL4g5Eu4JE5U
WI9E1FDJlp8LgC36QpC/3Br5danTrAgXz/E8CKKmc5Rw2LipFos2HD529DatL9xf159R5jdrFMAM
zb0LNtzV4KSIqcPizh8hBy/UXWgOpYFk2Jdtsug5FoQjbB8ud2YTIMVJmgel2jnkUCXwvwE70e2X
13hBG1rLyuCv7PVpe69/8K3IAMjyVqLs1mvVL3n/nbVDtOitdGYAr8bKk5vHZ40ONPJfiNeuLm7X
auDxc5JKlxPdyG3fZ8VGl7BbmlRAD3AZIcAtmS3yJ95imFNhr+lUGVxpzLL50dyfXKsn9uzpUcpQ
bdFYrTqvFRhc0J/BfQcuyuIxiT8fKv/8JvHQidlNuqIOIVMd7n9fznTtsgxVg9poRRFn3Yxlhom9
1s/MJfNSV45mxpDyhENsc0kIXtIUXsYGrLBlVZZ839wGPMC8Dd9DZzoz4AG0F544LnY3VFG6mqFg
crrbRK81jSZKTwMiXSYQUkHR0ec6oNuaPERq1KI82VOq20oLLAqwdzMf09H+f/jTXyq0gr11FetO
dGKGgCO2JD1F+IBn284dUsguMzZmD5LNnh0i7+f0DxWELHRzyaZggZ2zcXyt/YuxUTPmw6DD3/ry
cqL1IlNNLy1l08y6SYzcBdcnJ5uEgfT3+FhNdbzzl5cqmqDn3V9wWc84nrN9AfYNloVxF0peNwk8
MkMGQwHgTNfisvtdQLWVr8yV7tK5apg0gLXMxqrZ+e2VvLe3hfYPKYn/tMMPbneXPkoHmp9o/7pN
zjO0YpTTv8uXZkl/nq0oQ/rH7D2lYFEnIaetRMPlWoaGSwZsaBPa3kj+DEIu2ISnLQQs4bWS351B
A3s222SxAAA3kz7kziMzy6f9dBLY1vsPDKQBfoy3Lj1W9eD2EsfFy7idwihyseSMw+HtWzura8mm
JOlAy/CGiAgpdwlWjjQeS77mGs+X33BmeNlKI0FR1cpY4Gm6khjqdE+8evnWNvYzDZafg9YWt/v0
RfQYi3Pu0JrCbS4r9TTnKk6rdUpw/ksmmpajMKDcNyb5jkJPeOZqQzseTks6xks6U3mk6MPSszQD
zW3T/HkSSUHJcDALyqc1DQpaLSRvfOzfpVtHqmj9sdYXYNgPure2czn832liMDTnik6IHErB1rBh
eK96zcjgVjNHkIL4Pmkma5nAL3T7vcfv4mf/cFVEJk7+8wx3OFP+kTQiKgn8AHF6oVKK/XGhD00a
3wjjFPe4BC1Nynb+5li5+OZyipR/4SkzcEH+hW2fF7bJFmc44tVGL40ES6Oa5I38fcMrrPCNEPsg
mNf/PSBw7svBUeUp7K8WUsbQjdHs/Ca3s1/f/5/UsoN/uP8BGLKyoRhbjel4FFqfLJKoW8Ted95a
SAOR6RybAWPFnhDedwp0asbBhWrtFz0px8ghCWzIodrnTvQYBeyRCZ9fXATXPYFSkH7EdItsc9Ak
y6Z/Tqrnfn09cu8W4tIbQZQkKRmMB8UbNbPUt6S2JmmkhBCDVrwWHHWcEPkRXF9/Qe0/9PzytVaV
wtRsUGxgB3JQ0CsaWDYl20dxpFqByX7oyWZDMEJ69Gs4iSpjTxARhSYIJ3pbm+Y1CEXMGd+mqfmg
xuhypMaToi6nXHclZb9hWuIAv7vVcXf5GrbrmKvK2lJTYdpmnFaWDMLhnW1hNMtJwMvjESqdN0ux
TcNpRIUso9c4NxbBZqVr2oiQ5rP2ZcSsmCIqu2/hbkeyiH2t+6dZ6WXLdejUy/hbOYe6AXGueaB+
q1t+of9ROQ7jC+Hujihd05dJJ36OxQ9vjO6YZ4logwCx83PzaaL0qmMTYQ6/Z54lSmQ//lVH2rUF
RKmbSn0oUroxJudJMpld8up0J81i8sqMAWSzZDR7QW+iBVlklIVQLtlm5zxh0dDPCpvcgZkQw5lT
lsHkaANKZjIOKV4gKkiGNonRWiNdlp7M/w7HkMmTVvTBNlqVnIbKRbO7PRTxnHNksSaDgz9enaTm
FOgVgfciprZvRoAgx66F2ACssLTpCb9zE3ugNWTxifc6ZICCYbofFfIVyWry77MFw7BC3LA0XsdD
8/RdRxkkFlr5w48Z5grD5uHsxlBFgJ8pwCJhAI6WWD7dew2i27XSR4+/1WZCSbWKQBBI88WVr4cJ
+Hiw0HBgVJazrBMp2Z8A8GAy+evvp79K1Zbzq+TjC/6wu7D2fg2Fpoe+x2GEmN0RZO7jNyu2oO7g
DcEzxoBywtK04i4h+WYg4Y9xODXWhHXGoRp/gD8fjw62l9DS+DGbv8MaAMxw0A2SC/ptJ9xoedAL
miNBc/rgJ5SVQvbiuR3tMctNbvUJp/0ugnmriJgVJtRUl+hEpBEBJtYs5/7egENYRm7j+zXeXtRs
FBGZr7lFyaIOXfJvwCMyniEsAv1Up+0zZQ7mPxibOyXW4nqwMY6L7SgVX8BLJ+Frox+I9JG9a8l9
wTHsy1SIFFX1esutyza428YZAe7kwQ5oFC21wlthVLGn1nt6k+qUEN63/3CkiVE3+zvvA4yp05wP
OX5zUTqHIglLJ+Vr8VG6VB1B33KCQaL3C6GM508Ae9azrJ/uST/vLH0kuo/QGhCwjBb58Ya4gDhQ
47riA7xjKfbNk6qALUHMLKaRKIOWXPtqfrUdGGkYKCulTcEIEVpxoGKb2UDoEq6D5gqZn7qBsVNn
Qx4nLiK+JVnN8TzygmQEf0Cz7jGwXq102OM8/IujXM6k6fPdEDhm42oeJ+rWwrHIUklfShtf3f72
8VO6OaDxmHNitKr1LEvqiGvWRj+USFdB3ywE2PsKDeHcQSx+E5INE+p0kgDKRsneQ9RXtJZkESmi
wheuzU8BEanCYoX7Cmen3irdst1403oqJ/SwbiAL1dxZ2wS9XBsAG5kHC0v0eZnJZ+f9Bl6YmRaU
uwOXhBVoSSFRCkOnsK5ajNRA7+v0edS2HhiL4XK0VvbK0Jq9tax/p5H3rNUyELvNMSVZ6hUMPpOF
6ORLQTsCRskVUSgZ5uK1Hm08iHDJNbyOSnHqsSro9PUV/fmKdpo9jk1W8H48EFiLTqm/atZ5uT3O
k4exyMzZPsQHxqHrfovUMzX9BiS4SSvba6WJVOxNRMh7Rb8og4D3KXH4FzBAxi7bL/R9hriS29RK
BSX5b/ludJYP3PsUvISg96GRUzneVpAkp81EMekgmh4Go3uSUmeNwUsIrGUwjk9Mmi1eiZfWiWHV
qpGJAqJndcWsxQqfGrNpjHhgLRTkt9DZfoipw6YFyNvV/jSwDEZ6r4pkbi45jWdXN5lW2bHWePj+
ZzVLVrCSuFVCRN9etd0RWhFmnt5p3cG6CRr/hJGLR/KG8UjTLWyd5LqnEh6k88AA+WXzhMVYomcU
B++8ZXwJXT2KdE43eNjRDqpkoGjB2M5zuaOqNo3+yM3F0bCd1d2O6y27/BVOsMT4L5BBC9QgCdmC
/2TbgWDZu6hbAvFL4WxKjFxHnevn9kQiurCcS+4qcEtWBTahVqUH1f1pqK4pHf1poV7mJdqrNjIb
+AgNx2tU14LfpSVrf+JpvSgr6Am/5TUVh3bbn60M3mtxunLfgfaN5JqoyUdQn5pC32/3AOwm7sxY
5dEpXEFR/9r0R2pH6cFyocOL4X7XZR35HnRmRzyWUhZFCTye70n+jSRI/qO1hEU9EAuumnQpjX3P
PlFwxaCK/iX8s2Qehbw9J629sYiCRnvQNAzTojXXrxQYVpJ6E6Q67uwA+XxOMya67cW0u7ulPhvg
bsG4ep8jRB7o7ajAQKFsXBRgM2Pj2lM/Rd5tX00jJvxS6to4Bo8UxerKH6INt8f/mUZwak6bzX4O
OySPdaHVKX71uEIpP4/MehPQ/9ZKaks3QX+UpxVIxI7rt5YFgW4UDSDgdE8fMTVkHQc6jcRs3cbe
6HiMNOldk1TtGlDQsDmfZLhLJMEPIzNUmPmG6/1pvuv0iCsFUHzf0pso04mNgPC+3933/gEVezxO
gQ1I1xQGSga0WynKS0MSGGvt7tSsKfIAHCn7NyuYISxVgYY143ZqkzWHGKOH8LRWiPdlpM0Sq+Fk
00nGA3JJDsBVweEZazy/KV5QfY2S59UQUGXkK8Z2WrtTB9j6q+NzWd9srTJSr63eD9isE4KruOTI
xiv857kvyCsiYCU1znNFFf286pmVX9wM2qv018zLvjAqOZN5BXVR1KocslHSSEjQaajnZBBz8A43
R5yvR/l1FCq9neGDB4fIXmby8iI3xHYqFbzGRviRlo0lvvnaCVOoGKFYMsSVqrwdXFICc64E7yGz
9bhVa8QZ37Rj3w30pNNRzY8ev+a6lvXRv5D+yLs+3Gtbww+Cnnziq4OSzYnPKX+wmu6FHZ/i6wKv
5t6NZX5EtHgD+5KX8lThOKqcTOB0bstWZ0+RUrKEn0IR1e/Z5QZ7v1E0Mhj5B+j7eaUmdKRH9BSr
3g2IZw2HaqTXcuBuKkvtcsL7ZfbVZGGXSXFN8XpieepRPEAC8Camho6fcWBjA19oDgBhnXUNl3k+
ZWWg8k5chfMb02soZiS9kad7CChhTV4GQDEDI48S7g/x2qv9oStFHjs7Z2tlvKLgUfvhqyNCk7kD
GSH2DIg7Uufn5fye15OffSkUr6IVFY8imzO43mqDuxsAT8tJRNlj5q2ZfgYG66C0K/fvHENePg9X
5WiCap7xsxEjac8onhSMbugAYPgvAVgLAycTL8jGEGmXn7x3I3gTaGAA3Dgc3I3Z7WeMiU4BpZSn
WrdksOiAmiP6ei4gN1lhSyFAb9btjsWEmsn4b7xYWJAx37IvtFVycq3uSsPvErIQR/wSGXtaai2q
q/qwujZiKn28dL6wKRYv4KAtt99ydD+7XGEXpaWOLBmkVg1lBuhVusSN6+hEw8Sbzr9/XIv/Lnz7
lEEu4otW308Fumu/PsRExC/ymdCALxbGNVfmibiasz6nYsGGHrXv50SzO7Q8Q7+/zO9gDhigZ5wC
kdlfB8FZbzzIUCh1Pd7TRf4avDm/cr4ojsAutKr0IcuPS1pywoS5sWjOBlmXzq5wPlTtzlhomSnF
49RrnXzWAWVcaKP9J5+7cgG3QJd28lMAVRYyPIDfXesNHOr2MOkx3Zl09SmPlzY/spUkLksF7zAK
0LZSFk3akf7mceDIu8usO+jCmBxhGrsSwrxwupld/won+50ztGHViqGav6mY+cqdfsyc8hAl1MQ/
ROBPAIrPQ7ts9ZmdqHKEhVg8+o7BiojQqYfEpDTG1wKnQE59awgu8EAZ/X8CmFIw6ExQWXIpAXLa
Dp40g7B4Fmb1xgljMbbko4zeN+RYSFYRqhHCUm4Jwv7SJMaelamtQbDWiFTj2MhDQVLTii8lG0Dg
ZxILnRi4eSAB+KdZRQPgjo8TCyV7Ur6mrKevEAqXcFevgjC4dNyahvSSBhBcrIeu98qI6Sekmdk4
cfXwt63kAPNQ7EY2wsnvhU+WncdelWqteXeZiV60AwSunj/pgTVp+Z2pV9hgmeBny7e9kIOIMEol
HRqjD7sScR1wbhOUB+Gla2llZyETJg3FXTpepC3nzsBfORytpOtg2xO5WzmId3cGR3azNKdJ8VYK
gvPRPvZRoTKv/qS/rE9VtlP7Mf3XukHhal7wOBc2NAfZafOETbifHntLLnM+jyrnrWZY9o0y5GW/
xACqOuXCRoot5YqD1R5bJvkPe+87rBVT/8CTCZmZsr06iejD4XnscoFOvpxJO3Bu7qAvonS6z0gL
vVdEGae87ltHKtzeb3YnZTZ+kdU/b/3/cXZXd1R4N58BUqXm5S3NFYlpQKBMINkuas7sgBxm2MQk
baR1TRAuXgDV08ydhRMScGj0N3sAk5L1YKNWDUwJF83adZrJ6uqACf4ZQeIfGCiqMfJBfy42r6f2
X7CQpSm5SRZZPuPuVQdRgmbr3OvvqMJ5VgmkxiPVUhN62GLmAG8H32AEXJUO07XUKaTLqWljbIOb
MaZoBI6inIvaB+VCxA6EvdM/wKSzq7wZbgeuMDPUp2SdAC9ojEAxWoVz/X9AXkmLl5Pd6ZbvHqwP
e5wU5/s+PuShAynv+BvNUH5/XvpdDJkgkOspjA18ejej8LuwaCSQDYA+/T6gZ2JZIskw5MlLB1gZ
shcQP+/ZL51slrxExZ8LV35fQenLxtUwKGiEVR6TnlBUOdnAWeEROD8NKHA+LNjEzkdGOJQBlEz/
peSJ8f3950QhPXSoTpsm/Fvfd7QZkX/YLNm3BTUCci3pDZtE2Er/PDCSNdtSRmxYtC11bmUSHbA5
actzyWYrD42iqz0JRO2Uu6x2Rj8NcRH6JCg8Ujo9PID0AkXAkDq2pehEAWWFPo57NPzKMjow9cLI
slougt/5JSa7GrU+6lnFVapJ4t71kmqIsGSaRpS+syJH17gh1HAq810IvVHdyHpmTsrcaKUJblXm
o8Nw96CnymRlgZWCzcSKgHaLojPyzCvJz0PKjngAfF1jNULMEg3MkPiFs/hxSBVI28/a6G9NSzRg
d+b43JpSKzY5uL0MRMoIvWZh/1rPm2LgyNjnK61+GJ4SUn3iVOjXJj0DFaHpBSz9wA15TJDhNh8x
4Eb+LceVA2ZG1AiLQ9yXsAEM0TqC+ECTsOnphBcyZJshGAdItUrsSOpDTzWoMl90ZgmVj76QK5JQ
5CH5T3FJ7cWygSnrzpb/1CbWVcXY+tEwTbkjtrZHlfEJW1WAaVbJ8fYav5+VCxuP933yiK9uA37x
BMkL09jgfGi4eZarBz74c0f+fP+rZ9rYavTKukUPQ66sIr3fJ1Rn6zMEE/SA4ffkAS+jddJkkemH
hk2wvGDzI2tKDuuA6Hzb3PCkxiGTWE74sIEaeFl2O3Zxt2ecNFa6CU8+kD1DyYp1zuBiPtzKy2FQ
DLLvtW2A328gkbrXFZ1Y/rVEBzkEf7X/UPrRclvFSDaXZLfnone3OrJIu8DiQaXG30+KDIR2Tnq9
VhbMedxDuUFd135XSf/SU/6DFKq6E2vptmRjW3hzFTO5081BmBQ9TFRpZKS5KynDjPTJ40JIK5z/
Iwp5TFimGoPjlgjDoXvaLIIouiq66A07dzmdQ2/kjIvvFM904nYf5Ydf380D733KUHETNrEWrZHs
SFlWCqcQEB5zs3v9WW5pBjXhUAKjqcNecFdj7fS4uWka4sD0TLpp8PXnGeKTCU2WZTh2Z05CBpTL
xDSpeOINouwV37WjIpLyL62BJiIpEBzbZm/2JYbSfqa85V32zoFCwfjP99Qw4FG37fm7Lrkw39T/
GPTAfYRPac0IJwlaSRBdL9u5jZAJz42qhwZcliJOy80pYOTo+bSMBJ39TEtNNAhRJvHRxnBnEBUV
ritX4lrdoHKNk49EQcpj9zoMgIkEObJkWIVCTjCZoX3tsCwJbwcvgk+SJAObUWq+US1Fpg2d5nhI
N1URXUEJlbax8fAeI539be7yH0rJjCB3+xVRn+xm8GmthgNx9TD/sq6sR2OcLPv9LqP7Q1r3gRyK
bh+41sXp4WcgtSGP9A36Y3ww1Agxz+X5/IpMTOmnYY5bWNY29xZtlPndVXkWvw1wSExOr+jCJkcE
o0dGf68At45u/DJOIxI1qEBOR53Id8Jv9SFT+P6iBrt9hPtbGGCOYaDjs0pn+VyPWvMSZ+Og2NXl
VW3v7rJb3HcWhadWSh8hXkvtyNF35+o64qmFBuLB2+NlSSHTgjXLKziZ8pDm6F20GuMQaDfIeoho
yjwdNgqoRe89Kk1u4MPcECne+TjamDKxgOgpnod3C8xBICP4uPZVARvu9JeRgZ3l38p0gH5dOnNd
WKuzooubtocaay0WflhClhQMwstenmvLYt59g6h0UPim6Kdjd0JOZ5vcjxaP/FLaXKgkVgaPYS5f
SMORHnaezlEtShg1uBBwePpFLtu9G7yJDqh0VK0SmECHK1YgCHJyiOUdjOYVqM0hIbKsvTsnNcCz
1SlnHpXWWeY1AttSmwEBLkdRYTKbCknY4K7ys5q/PqVuO6suSs3CUCFVG8uawq5VQ/DoMeGV37KP
Ed0n109rFUvcELoNpns5dVgT1gYL6nnofEPYkplNJamgX4mM3m4qZvxLrnI7j2kkNIliVJzWBj/M
h48sTWYhAY11u3geGQsuB//2c9ud/hgC/xcRz/itGyy2DURjyG+/6RBuPKOXQhG7cP83x54WxL2i
tmmB27NatefQSTyrbEyKQZdPAj1G6Z9jMe1DHeKWcGVOgYk/MawcHmNL+TkWd4D9H8HCng2nqlD5
pOLtk7W+0nydkrEbG2C7tFQs/YadztMYo/fPOQCdHEGNNSUH4CR63ciYu1IubqCh9/OvjfImAKU3
4uy1LV9dovuRfhC0GFi2ZpGCxxxLM9FhUL0jn+unpC6GO1mQQzlqGTUnD41NqBV84C/Psgj71psE
lwqqTXJdptptXwo0eM618pb/8Uj7hRRyOTPXm7Ob1GliyITKccuI5q4/jSofI5r6XMmPlOAk/z+1
aXWvo9O9dz0ZIyP+B5thbX/2rbSBOeL9Q0d9f4MDPvP/eWGiRp5F76dpPNRLkuuGv1fKApNwkHSI
zWuY8hZe0DKROEzaaGRg9hTKJx0yR+G8Lh/HGyu+z4tDn2kQEet8AuNwCi1ckBjP25bkMfKBqboB
WRra3G6qihfq6Qg4x1qb3d8GNj4gR6gnpxrBy3rivyg9dxB5eDuPBKBijxjlGSsZc1yxwy27u35N
f1LzUKc5u/2wn6HixfmnH/F1UCUC7C+RHjA1xJ36D7cJKELJ5Pq9vLpleyhaYLnJxxBl4SAt0IUZ
B0qOcVCbYOX2/75J/hEsxn+HvRT1Loxvaw1QhWZzrLXmgrOQJwbMCMZvnHlGAKIgFkd12g3IlxAY
KvsrTCwURLOmRx1ryey0v7x67Y/3lb9XY7THAhvYyG3j6QMhpOkKkFd9iOWz36mEeV8Ua9rp1/pe
MGmS1ekKVtKm07QuA0M2RQ/rwSASJ2/7AA9Y3VDO+l+8D4JGS4jO5U9xTqieDR+zyRz3lairzBS0
InrXwqYB/LEdDR/ktSr3oqImrzJo10Vo3kwUW+BR/a57dtykqcsynvMJlxtdHihVgeEUWJqk3Ckp
R8VnOJjflt7vPcW05XTrF0W7FEQb7UZmbjEEBrtlUFPtTsC055F4gEhjevXOkIHPt6OFivRpNxaf
/E2Xz0dDvr+l0Xl0sFaHSZjPrxg88Iu4iexuPZUICiCjoI8XESSVr0GLO7MO6lLGSArH2l3Txme8
yn/3it6vCxp9WXluAdS3mQWeyuJBQ1adbb8NSYICoHjZQIdtg4QXFNo13TqGsdQ66a3G7DndiQ8Q
9slKWBqjt0m216mVPh3J3+spV7B4ycA2PkEjRW0LpjXMz/th+k3ACQhjKULWINJanaqnk5gESSox
hQYkXnjhnor8LdhqzSgC1cfeZUqLAZOZrLdwsfUwh1z8ox5vcsbdImCQlnoZyyNTIxHAiJwHRuUG
iCR+g/somIavujZbahWem3qBLRgm1EcrxzYgx0CFvP53/puwFMd24yynUCMRZPVB3EdGhyN9lCRz
/RXayEpWC08IfaXI7iUvnXaJNJOb+XNnso42lLGOGUCSLRO9rJ7a/6d9vTFBP8TA7+4BUt37Vspm
9hZxa39IW808uy0WO+q/6aWS0JJuHPUZxFOALjTqjmbtyAQ/ZcmvrrbLZ9bG8V8MyW4bLd8TH+FA
XUSuLe00+KeCLTM+Dvineh+Fv9VBn6iPeY//raPdxTuNzEX9N/VN6ovTWIZ2qkLvAkEpaicYEOuk
NPxmtoDiPNIZoZ1kC3wcddbZ3I0+r1L37lC8Y6rXPKIj1Vi+IlSPMnOXbH+RBIeVHyC3M7V3LqHc
BYRT2GskUeGeoXc4cSQbJC/vrMPuya51ZzIFR3iTPTdaDVJLccQLJQHWL6akQT6O6OTmO4/F3uMk
pDgxak7OV692sZbR74DE+noMBRKTSHViOwgSIENp3gMULK48efj/F7IjpJ4Dz+xQWud+s1RmXm+Z
xfv+hk/2QsE7xyrI0oOxWYc+7Zw0C4Bw7/2TdfKKlWZLeoMsNEKbXpmM2MY3TrgSi63SICaP5Knp
CeRxG7mn12gJnghMSbtd6KEcbPx4jispR+RyUwsZj6GZYhFozO3C9UajakxVaK4mqEO7stTdjBGG
+4GiEALxA3f27y5EKReiJmTsgsO0iCCukibKbmC7jrXZRTnIHmJMFOpnar8Waajf96a54YAUWtRG
L8uSvSdrJUNsjx9MXWEX4xt7TLVOUwYphaKtAskjWlz+S9axZNMIHPnL5B7LEZLR8zL7G1KlBdFa
ilGuTYnhdZMTISH81P/CtuHHYPjeHBq+oHZOeVH2qAzQnINsqf9Am++h9OooJ4RmUjmiRiSz5GVe
6iNTlh/csygHLX/YQVsYGq7fieV9pj1qLzQ8XDPLeCTy4AB8RP4ScKo4iTT1o/FRqxoaqZ5QKV5k
BF92PNZ+CURBnvbwqs4j4KxKCCmeu3acMoGEChEmrkQRCMqnIHIoFFQeSvSKAvcWvpFMKECoF1GP
PhSmh0jks0myjkvVY9g9cESLQ0nOYDwDk2TR1NO4HqEAUlqTgphoYkc45nVh8OYtDerB/3KaHw8k
kAEM8LdUo6cUNoqkD7CVVZfgFBODlo9k9SbKhp/Xaw3R3XbMVNA6Nm9ZD22wDmcTYNvo1Vc+N14P
yZAcjynMOzwNq9bqd9Wk0fmVeBz1S887T8iqqoS/yLW4f6/jUfxk332I5+y+PvpZQ8BYya2QAbeE
Ds6miAkDHXWT9MU39KkZ2Ww0IUY08csGz7T51yn4QLjtxmeM1LAM0OoAs953QV/irnTCWuI2U4Tw
tePnwyX/5gtzKNYlXgaeUrPvsXGXXpMxjGUpU6XRXEPIZf0ZlY2/awaG9t/SEJr3s5JiI7bQ4apu
9E3ukygrJuKpEasqCF3KdrUppfTXC/p1r5WV0hD766eCpoqATvL6EX1vi5NB+IpqAIue3AtFKyJK
3U3WcMlxlKKt4Cgh5jdSjGtrAPh+Nw2vBQMA1OKNz48zJU0FvLG6mkXnEI398WfkFjCTfkvf8rbc
oSzCUJzl+l5WSiIHvhASnhgHd+N2vOegxGDCpumObGHWLzgTEnM10XkDFUfZ4ifSn2TskBNLQ8yw
TTkDsTCgJv/CzG3XrKgUnwwyOzRnHd1n112zR7LwbQl8qdOrCc01ptJFtvCeqS6nMSddXeUE1w/A
vV4304pAulVTouPGVOvRElPuWlh8jXcf0OeG9jobjrMQ7bLlDN4wOzFohxPK5W6cvurYY1gtQVrB
KwVTctcVjLSI+L9l7SAjN7elHHCoFaH6cCugyGMQZIyae2pj7APUBNhjW2X88m76vsIHQZx0wilC
yauSOJDQUg9j0iMw5m0snto1BiO7u8el0kgJGkpPBH1F1Cgo4rsfjrk1y7DuT2h2Uh3duX93jt/9
g5vr7cLkpcORIKXUMU98NdDfLYHffBp9dRLcMFNsv6g7NKX1vkVuCPzmEU+FAVEmc7eEgknoFFlq
dF3UB0g2lYC4qQC60nY/NJlwenuguhyeJRw/GhZd+FCF9nDV7eCkVzNkZfSlUjvKE2lDe/kkf1nF
gnu7V3+HYn5t7JjRMRzSQXYb8ph87JUjn/UThp96yl2y/LI+phguPGygo9KzA0Bn4o4OLt4KTzxW
soanyrjxJB+0kUD533AmQfsxZFOHYWUVBRVYVFiadqkJnHLB38KNYM32RH9U+RDRFSUO2EM3OOJs
b7ZpeCZrAHuXcdqAvoYU6lCm+ZQYCCQmd2HEtpSZ9w+E8dO7Ud+OiX29wK8OVXplb+Z51gr7gqcL
0oyj9xI82TQf5BS9ogscMHk6uRciY6DVjUZGuphoCML1QC8vShJkSU49TJufg10Grp0AG2W8DwGS
nkL2U4VaG+rRq0JhTPAfkXHZst5v8oRCVYCVlhkVDlumcrGGcubay5pabHYny1D/dXRnJxImvFxE
3U8w+1C7f5b6i0LIbVpWrRjBB98KhCVNgi4RdH/EEJGKDL9uLRz9DOutb1uQqxlBJQFpg3XvcxUg
lkiy5yVM6cUd0oVNZ8p0jioFq2o5p+WtkPrfK23S4sH73E92NqJgEHgMIR6pm47G5txHi536ND6E
F//nYPCk8Xg4rNxGc3kjDj4vwrLfCBhXB3vKRdPYbwOiofbpfrOLEkFp9MdFgvmI3ur6mZuPgwdD
mI0Wggc30xH5ZR40qkUg2bgqkb/6D4qDDSC/cI81DOLpIc6EATL2wle7bAYHl2GczsTp5bluQWxC
Qn+j4y0uMGZR8PZrLux8ylJwKSYuA2gX9okBrO4NrvBjVQ9xEKS0UfT3RHfVB0ighi0bQtOemfDB
ApjRXjtnmRUIFRrQABf0vKSd6hLJse5LGmlvt1gmhLZ6njy6kxOD7FQfXc4kGas58nZyufgwkK5O
8sA6DCW/wRdCBf3NrkwnUyCPjTJPIYQwQ67Cew1OG0x3aqxDEELpp9zT0j6IlQj89gJs9IgDC8Bm
fQjJg+2K7QzC+KmFX3PE/YLK5zo57CxlZUW5qVb/I9yrsQI0hbm6a8NVadSsyaX7sp2nzjclLtZK
0inPFOa49/LWoL0URAcsPVf6Z6v8ybvrnWAAntNbdO3UTSs+tiMr/yb+4CXvHZfAWPT82nUF8DTp
W4dlxer/QdozvcAZPhXTzuGIGJlewGMAJNkBKFqfGwZsezcri+eEY1EjDL8/S9Vk58JLL6sGXgs4
vCoFKyQD0FdIlTWIvmYFjkZ53Yc1H2T8BLeWiQPxvOS7G6LMLHN3mn6jEqjIi0vpIg88jkyvC0yP
00VbexNehKcwqLp4fhEJjvYN9/q4FsumOskn+PKPhtSB/nfaIY1Ub+7/tF+4nEyu1nj/9hjxmQdu
j8jL2CyPCIF1ahAaqX7xYvSRqYY+JPPFyYMU4rPQ/irvbByt9bfYspozMVgRzQS7NoDH8GL6DIXu
pQavfJlCF5no4nXIhmZdYyTkwxBz8NyAPRtLNNZCpfLLNBcxQV2troowhAgQydZOqvaMQbz4Ednm
PZuHkmrxFiXs5DKEmoz1Mei20oF1UJqPS0uxJKsCQAydvrXyU3bEpWVXZbuWH9lOMSBr207az9UL
URHbKoO1Mn9EBWix7jENKdN9IJOF9q2w3zSfx88dngAPDTAFINZh6dfIz2myh36yeg73jGsVhjS6
k44UlkYGxXe13D/7msWm/AqvY0ba0BgJZR9Ph33lHZIw29WfCz6aEE7J0n2BvHPWBZ51mVaPafgr
PHXXXzBKH2+6yuFy6jhoFy6mLoJEdactI3SZzXmSH9b7WJhNXcoaBNm6WStRAsWrqPB/YBrtTiai
MN4tF1pPtPF3GWYd4J18AzXQy4MmwZxre1naqi9WBghkflElJ0jzjw6S9gBGX68/eVddTV6AoZLo
59wAuNaeyGTHC9BJyMdAFvipSbdTFGlEX1yLEg8CgMVVMn0ys+khhzRpANgdbmLEYI7FRnJ4px5m
Bp3bvKut60QaXU+fc+XkbHRsSiZQW2IomI263fKreuo8TfYSuo1Z9oNTBoK/ZyLgsC/abQkOgJqh
vJnKPm3/MpAGMFoFNglKtH99unct60Bn4m2NWa8ZoCv344QElP8KYsZqgUwhLoz2UXzYYxfsaaaD
Y4SORlquotrQQQIahXxOcvE04IfFFCBWLLlq4J0lo1kiiQEYZpVIGQj2MOE4PDSPGPIC9UoyZIkq
QVUFn0crTKuQ6hwkxKxoDBoeXRaSMKRMMbjv2Bf9ZJRDBKEJjFNSHfXAsBGds/Y5ovwy5Eq77Xah
aInhscMyi/27Q6wBiEcR35YfnUglCdh+LvfeFhobAteJ4ywR/KpxcRdCXEkGsR8uGap/9PhcNU0M
Pg7Hg2R/YjsIkB+Z7rjfvnIPZGofTaJawv2t3v3pR8JaS6SdHKYkG45oTaEtyrLlCnNRQXKRWM9e
CcSo++qtl9wlDqEEziBJMliYY/f7dZbRBTgo6HetFIPbVqLHKov+5dcNmPK4KuPJ+a37RvmFHGlM
UxbJ0/QXkNIjmQLo05pplhp/bJ9OeJGKU+aIIEQ8tILuQQbBCL3rZ9+7vG76zApp363LmJPMx1ck
cVQqeb3w0xmADMlbEt9IPI9StjC3HcVpdjf73lLG5IXYwNSMAue20R9SqDSDmM+SdZvT/Vx37Zs/
pxpNQs6y+tXl/KUujJGIHAidWZH3fXqol27eGc7dgxFHF8KJj5GqGCaPFUf5ENApCFC8YUOLmj/E
7p/5CDtU2Ac/fOiBIXZJzr+1new+x742N0lAPw5CjeLJVvgScFxkFMa5P4BdDO229NqNOw+GyWuh
nYk7JhLhz1g2oUW1T9L+F0Pp1L4ziKYHGGqURKGM0PMHrXvTffrqNytjJXBR+SxXfsM3B+cZmdxS
CNM4/CgeSUeT6pJSTj8fy+XLrYXgH3R3BFiRBoK7JY1btIuphMwhrEEBBKzjm7W6HpRT6Go9LawZ
3nfNkLMNcLFAJi1pjZLysy/fISY9WWzvOLZG3HIyQIw0dUawDgxdhCXvpdy2aljTqP+lIzV2GiEN
G/8bYwYtNxWEJdUaaUYvFhzmduxoNVh0GqF69ThrvXZU2JnlXw9Mnavvur3pXzOv4RicWSJr6XF5
NnDUxgK5iVbGcqnrNY1djl7kjmywNAVq5w2oJwcHCVaGTX/4xZLoLZ7217gXsKuzmpXmqqkZz7Nw
qk2k5GzaJjc7kYQB8GgvICTmm46cwae3HW8bVAlaNCtdoD+q5/hb6/0s3W2nzJran38sc4hdjmsn
wdKlkDvpSDj85vvPb3qrDoWBSm0EWscKVTP91nyiJB2I3Zy5V9BueIrVH8tW+v7hIjSrgcS/XjXp
w7dqeMDkrizwNExz85fIaxmmtYkFPTPkJboSqZ5jkT/OEM5Ap5F/gAuSq7aF4xbBbIrssDzv2Wm6
1FIxlN9YjqZ2yAbZOOH/+/9y7zboZDprjWFDgrrJUlxImjEP+r7Vn0FEjNwEim2SIgJ/4T5snyXk
VM6IQgWQyoW5y2FZpsfNClSX8jGGk673CaMsorqE6/hImHr+f6LguMBaQZw1ZOKE2ZsKCq+7SoX/
APtOO0x4L42SjwAhVPFl1ex1OvCILmXvkSO+tfIYfdAxCnJMPdSs9wl96QdhoJQwFHlgZfWu+DrA
pYqfhvF4u4nXX61yG0ZPZnajhenJv8drip0/sxb7RPNPKfTBICjHi6OuZabYaX/kxvwEwUJoQR2J
teIZpXu39MQCWBbHvZZQgO9AV/z+KzzCcLh/gw/AIxnZZsXtyVGdX3V9SEWXKo3DnBYhWhwBgjhC
oWKiUcnbyej8LGiFsqjTIDXpBWqdpqiDdPDTfPBMjHoeeXzYxHfKOuaEreheZJXoAvsdonR3gf4z
lZNjrTMy8ypQNC0NbtZpCiXXDQCGhRMXhkVdB8k2/oB5PR3LSV6hgdwC1RHAmANcIWl64kaHZ9mB
ke4PzdtMx53gTWqt53VAZciXczu1KY/zF7GQXhoXL8RV+UvgB45409zDL71fUT/vFZTlZRYoWNa+
t7PTfFborUTN9mhyE/74NZrIZwR8Se4DfmY8qNux8e7SNEhkYjmVOx9eHQWcKkV72QrnchqbkxZ3
b9AIQUk+V4ET7q+/jtKVlA83A/xbU8R/FLEOvniqoUxKBT17QU2QCE9/mmMUSqiAfIXMaBHUzi3C
EFnKeaKyA3XWzVIMuS5FmvBilL9ueSNUQMoLaAP3EJELjJp95V856pyeycN8m3PqqTQAieS+/h4k
zuGSX/FSTEasVen88ES0CbrrwFVNqSGgVMjUefZ9NTfzUWAJuEomV/d+rx9ZUBoLkOmNjE4DMWa9
pLMcfZfH9vOOwusG9K7vJJPXgP7/8mqwZWNYtyraVIb7uxCg6cS1XmyPcXcZOPAZ/tQ6ATqE4Qpy
JoX7l+OCvGzQwWkhexDHVsW0mpVO1sGOAWpgZeWePvn+ejzNhLnbDDZDk/ipWoNX7If2AhRe+QdM
iHZZlbrxTIzdQEfDkEl7TPDFR3oS4dCEEyWwQFZvlmuv5poufJD1F07XlkeiHpgO6Uk0y1GX2eH4
9OVodRnrVp7/RY9m4FVN7lbuWwhpgiQBoaUkkLMGlzaqj3SnmRm1isBbTWM57uNb1XZ7w74WGEBD
B/C5SiXAnkp6V16bVPnnzl1lkfDAuljGCCUpIZb9RTHRlD3pKK262Rq+1PRtbJb1rR/TN08A2RRB
KAriih09PJNbJP6nMYZMO4yLLfC3ePXYX/4NDjMxNu+up5hps2IVseAxAvkpsk3ixEuHhprVicYX
RwnAI+MTLUSqWD3kkaZGJfcxL0ohj3Fu0tpxZW6V+2PdIKDNRvL5UHB+H85C5Qwf0xEYwiskPBUT
rNi/V/HHRvbXn1BGWWuDZgD7B73mtxBfQkFvmCp4xIKYBNajN2TruShX/nwVzRETTKZ6NNyTCeKn
WIV79tQzUkDtSpSsGlu2UxdsYOZ9aBzdgc3aHOR8+DO3cxJLc27cVypxqHZvqxsWwy1RUeQ7c1kC
Zf5IgGq2u1jmYXIHAkNdmtFI6MxVJVPlCe4lfyEbi4Ky6Tccj0pIjElC2EK8xcTx5UeGpQvaESfv
ZVkALZiR12S3w8LCUEAfuT2awNyflaKU2dE2ErXY29c8at1IJEeE2K2sDuICxOwfiNdlLKlPGMGD
MEZlF/fA4gbLjLh3ckfCle7OUu7KEcUuAjYgFQH9vMo4NvmWkiLpGlQwNA+gKGVVUaXAYpq1jZhj
IJ+TmgRn2m/tixMP52hHOPo15m/yV1ky5Dgsmpmj+YWpCHdcOhRdD15Q9wqkEW+1wEQ2Ni6y4Y2K
fZkln1v7nBSmAWf5+mB+pyoeRF5FkP8CdRzmMwVa5ZFFfoipg3/x+iyIDxtWzUZ5Qc/mm6nmGTel
Krb+SC61Ckq1Zl1ZfBryyiCy7t5Yphx8BHBSXv0LUgRTxwUDj6KSwWl9MPOQ8mHRi7vjQaaXx8YH
2Zq7cXeAzdTON3DVPRxmVAiDCPy/K+Dya8WJZPNJmjDntFzYCjpUrcFHubzNv3UNYD4V3ZcYheSs
gSLSgYKqumw1nRLEFldQ7A6ygrussStwUW2ahfL2rzWNtML17tcpJwpuOdEJMatbGHBXz/AExDNO
xGLiQGoQU2VCFUSXmLaYpE0j9b7APOgM1sJoRTRz67a2vJiBc19qvRm6glm6aYVDoxqa9kvpWyFF
GYfNpxmluIRCLy0UVgFpb52khgKyYyxAiCzxTUpRINT8vmTHs0b7igpEIngxJrNUcACehly4GsTT
cmoeRFS1JApuN4Bku5tCB5JSGsvtxwp5pmB5Rme4QGVuOCq81Ayc2NluLJUpCJTaRSawSCFQ090F
6VfTj9ZTA4QF4WE2CuwSAP+Pfrbwilbj04btSVyb1wrOMpb0o9bC/8HQhhga8cq4e45EcJxkr5tf
Tw95pVWpNeif7sIQsuunJ8xx/PIC0Ni1l++j01MdLpStQ8SwCnHpsrkgrLGdbJ8lZoso36/6E6dI
W9WpuTf29o5sGpzVbnbd00DZXUmRnXNmRvC1t6Zt7A4HKBqwjo8umoJlxI+ZcULB40Wd+7CT4nXk
b/0k/GxU93BhrQl2sUGms8bIxkaa0fj3NxZKX3UCgADYEa7cS/aspfsnh+EX7FWur2R53r7cRktw
lmAgKaqNqenRz68jy8uxY6T5+PXNhdY8QYgABG+dQTRF0di9rQ0sPqYGuHLD0/sUwYzcURrTmoGu
dZH5KmNwFUepGzcF/UzQsb3mI6UCrM2eBcxa30HVzU70WXUwsQg60t3TGrpQd3W3McUwEz8qQDwK
+Yw4JG18kfcDOGQjgDOl4lsDG7MZa5iDJBMWyr8QUEW+2vXUxkBhFfJAZgRiVyipmVt/kKsJ2AdT
g3+WxycWPIMBa0pCHtOUUtP9Q3BqsIwCkGNgc8Gz7d5+j3yFaOlRuwhwOfwsvnkpFCo6BuwiVBhI
ONICR/lIoKlJARZJMzP1Qj9uyFgP3bzPwPD8Gxce+Yy0gxjVXMlOc6MLGrKeyPXemPgkCLYGHADh
PLFmSh+Etx8CVBKB3Va/6Mipb5hLK7SLP7mDX6RhzdlNBBCz0Gnu7kGyLOOAbbJDR4BqNsXyiSle
TgrOLm6PXnV3Hm9+Juhg0JSsWKLBfsJgq1sTrIMYTOMMlPeY4+IWWkyQ9gBEUlPOUaxPGVz4VUnE
7XXi0en8tVKBWWOAV6LRGcF1c5mGGsyE9JIJn6kZLuJx4bnUhBZVEGXp++54/jpjqa3Cp98/uzug
CSCpSRtWg5ZQCfrkHNFj+6PG3ZL1aYNdBqLyxAMWDwDFbbJIRXTaAde+xVSokBoJ630S7FY52IPo
QNZmCWwYHdOVAedCsFFm9cPFPulabZQVTjoKI87yYMLZ5gKBNl1NRO/CTz54LAVjSOoZ0I/bBdJC
mP/mGW+Bkl4cDuBUS5SXfjsGPIHtNfkSuvAsJIZUGFTdUyEkri0igX/pgzmUxLZlMlzNAGz8JVcC
sopSpAzHpO5mYPojKXdqjY8CCBdWMeuh/AxD3/0QoILmJczcVJ896cqXD+7JWezMySz8ZNqotFdw
krKsaA1zQlbv3PKILhnmDKNbm7RBzN+8J8QkxNVtfh8R56J5qPeQgqJntBMd/FQCUax9Ybe/xv2u
Coh/Qxz+H6zn5nWhFX/W2ykiSsyonolx3fiOPrk/9yRZAyVtkVxkw2IEThh+Un58GwLtHFHtvR5P
SW3qnYxB82BqJQXlSIb4XSkgmwj4dzazWNHtD47mNc41Zyr0ymQVAyRY3w9I4CEzuVFH2BmTuk10
O6U/DZPKhECjt4LFACZ40xzv2QOhnM+yWAJNNxfFMOEvNrITsrUPZ+dBx4KZcEoPtf4KNFURrRZ+
5Yd8xaTwmpVPBQrzRHcxTvgA6N7RIFNfbMS1pPW99c/F/cDP4ElSqkK4VsJHZy7cDQmk3zLypkn+
8epeBjDzm7kCSpk/bCDsB7Hhq0ozc4r8Re2l46qsNgBr1z05iBqqzc7+ygVsr2AtEbQf5gAEgDJP
mF68D5qo3m00WvOFZx8EL66DMVUpR9wqeHLHyFG2A4nAEaJlLrmvIym1XOiP59ReLSSepf33ekug
JnljnIyRyUndP554cW6R/w2Sck8v2AiedU1Gv5rncEEvT6PS2cH6C/w5DgvAYwqogtzqk6WJTc8V
J5v9aKrR94/zSKgnxdRjQumU/R9TubRFuztVShc2NgrnPlkkcKoRZhIJB1v/MVehjA2dlWthM3cV
1N4Vgzj4cE6vjCdERbzRLD4KfGGyn1/O5wadWM/s/9+ebTy65vZ/6iC3WNHu4GGXtxLb8/8/lAEd
fb3Qj7dMcESnTViT3E1y4S7kkCauERKY5YkXG6ZdDjQ+tnxWLOXxOZoHNW0CVlWTagezn4mHTdXq
fmV8Rp+d5HFLivaZoo8WUyFDitQ80kfSKjXnSIO8E7+b1KGp4fXqI04bjaK+DDAuUSNf6+PYjoHz
gU6rIUKNTdpkvbQcenYz0HqEK4IDhCr3qNfKdroW5MEmYm2hvBUPp9gyMxw5XTTk52Ps4hH05kdX
iAiqYnFqn6btEJwByS5NFaHVQYk8k/HwQ5j/F6Esuqb9HDOolAz8dNMgPcDZNOhaPIn0VBJeIIm0
dNU9QddM2nGRWIh8XtuQKXIUOOzX7gBJwakFrRxMeomPgtJf67f4oTuzs7muNhc7LjcwBri0c7cu
4UUS/9OatUl8mFKog93NLSTgiiz1RqpVHCjHfvGLvFoRYMe8shmnx1Rdow5xrp0lmJBw+ftxL0jM
odZdHXjtmFsy2nnL5U+lIZbvY+n6wz8AdFFywiVkx4NcfUDO+x122JOGDfY0em9iMFT2tTZT2kMa
Nshr50rNnmqxnZr5/hDebr6/aqK5/YpfYMgFxsHnrCwgf903w4VkTXTI+XhkUWcTI6+IMVTzjb3z
tGhymJjTWO0nvbsCxXP0ztqN5CXct7LEoaVa8+KHslsWYxAAe/izAWmhf16NUXcYIssUYSq6rmfe
vMizPnc82OLQfauo6UwMGCs+WDg+dC391AW2FaU6WvPuBVxCjWScIflwyyooLlCu/WYemI/PQ8rv
XwP5W3AGK4WbInElFLTjXuD3aIGIfK0jALt6upWBKk6mSyTS9E6CFNBnw+5QnOrPEyUSZZmK5NJi
JYpnI+qLuTmK6qJkr2lbaOGCyGBhCYfyg4+81cPhI3v/n/TdnjF+ocaO5hv2g3njgT8RJb4ebJY5
0gJMIIlmaGUhyUKmY1Gd8KZJk3hMePnguTyymjnxfBxeppnOkCoypYMdAalcB7VSR2Ph8IdvqmkE
V2A5Wx3dbdYIfl4j3v55HBYYJ7hlVjDy+M7n75iGW8RatECNXk6fRsWllyOyIFOZtUlqbG1wILRK
a7rdnPyABsXvFmkZuEtqTSzzMev8HftxjGQMcb7eLH5/Ld4q04V5DAoCoDO7NAlpwumgO4xxf7dZ
D8o2oeyOLvHAqQfZnnuJrvikimTZw73ZtJix/XDdZlU5EJ8rgvhI9W6n9nx1HHJJ9aMtaASmYQrz
54rlZZh8ByuTeksVFt/xxYALyVeGr09wewmRxTVws+GUT28Q2J7u+uYeyUKjStEiYXCxJrEWmXCf
26E6EwfkxXdseEGbMpkpN5j59WupK19x8EbUHaQWACg0bhI0HtCbCO0GiWyhoGWLFqtEj2e7DlZJ
JOpahXt5n/KKhB432PvFDe082QjRHALXZHAsYCFcD3NHc4ZrOv3bqTUmGV93gsfi8Kpu+pIR4Wxq
UtLi8u1f5vbcHs4xtrjZbirpoES1+ow8JN5YSwV5Yms7QwWFons2TnNCwHWYBOvh6+P9eBbG9Wu4
85KslYGId9GdUT0I/qYrmnir/yAWzMBC1K1BZBflqCU3S5AJYK+8ESq9IQpWcoAfKMxQXc5N8XhU
Mk/zs64Kw6PEcZhIkFRIgT2BEa6NY9i/6CWqATAT5xsZF513LhzhaRm9fA+iMPrA0gmHmjqZw76E
K/tNWHwf8PddkaIJpSlriDN8c7+fxdU/0BF7xRsi8Qr5UaW/ncSPqaMjLP4DF+DDcL/Rz6pFXuRF
5nDl+hpK48WNRp1KUHt8duLpHFXheIHOHRP5lgjYqqlLRY5NTTni3QxQL1TsNMWhsqf6aSXH82qU
RokZlwMthckH+6jt5JXTGRztXACnTq26SYgr3j1ZqrNl1d/kuOLoBNDqulYzuqS6EpV0NlYLgJ4Q
nSuo5PxnXl6HwbVfWSdlelcMg7DZBgXsrBZjqG0/nBohLX0gJjj+K8M8xqhRHvb2lCXlxKFMJRBX
FDzmromtKFgygDPdWuws77Pkprm2d2DLuiSs48WjUI6dzXpTspW+S4n7WBLErGKoZnJ3wPB/XM3E
YudduSyZv6OdOrjyX6ayAicove51+QnxV+PS7ynmQhd6kacBtRUerY3h1HQi+WunqUqImuCm/ZJz
GDrBHbO1QALdC4p9dcJxFbuVVIiINAEGKkUqwWUpBdycroKZOXOreNvUSMJUaYbhMxoCcdAWad8k
vIwM1GlY7a6+MiY/EduAcsCvwxUaUXFyKtAh0KcNIkxb2jWNhu+QQig2cIX763/lyEZutFpvr0C1
2dZb0kIqBJGDi7mt/VhGZQz4M4wgxkezZ6kN6fq4X8/zzEt/MSqRYuYpxHw23vBXR6W8eTjc9hI9
X7jwv2rTvOQ8GNFVhQJUT6LkzUUbLPeq8lmSGdA0L75f/AD5oggHqOluOl23v6Dluyxlc95aWfaS
OIaiUuyHwbafMbZreUHv2KsfUjwCGOUqVlhPTvaQuTpAIuZTtRmLc9pGOuqk0TZL1zL74/yYVjlI
HtFvZEvpzzhIfEUlGr+hu+zzSP7xTDYaNVpcq/aNnOqT8vveQLuHoVFqZyux18txiishzt2x07U6
AXnpFxAMID0xf3kHdSPmUJaKOOZKO67vFv+C06f8XMLy7VsZmFy2Rxq0keLGKKqSgD8oNx+1NFQa
HOhNCIPfAhq1gzCzJ4ojLE9C7gdSRnyw2vUKUMSUwutza9Cu8P179rS9uPC9RaGLDlYdG3ViBB9e
uGcJtC26rMmxAZ2+J0+MhnjlQXbO6AlR8oXy+qvaqcLkdIPI4ULbxJC4sJTju/udOYi8RbD96NZk
A9mBNYpFozUkyfDaMSXLum7NIpGxk47OV8tJ9nDLaZZG/kO1XSZs1jsI0W2CW5LrLugOz/qvNf6N
FhUCK0E70K9TWp8pp1fGxRlSxZhDae8lKkxIkfCRCZpvsGVdahe5xWPKHCQZq0oBfDBoXG7qvgBM
mcM1I+KMrV7KBN7+QVssYyPBD1dtRC/WQpPFsxTsG3akOU24K9TSiTl7W2x1upHCqHbMKZ9bIwGw
bpNRG9I7PlUmors5X/e2kX3lxcYDItv0t1VqxsTV/YNbyXTuPdGyrVw8cojFG2TwHzSIqXcjuipt
K7w5gKrkc82SS9GaNlMzytbTPJCWLqEzNtGHV9QUt0SIPqRTObX61TiIf2FF9yX0TmDPPcBvJ3cy
zWFQrK4Wa0nXq1SXaz/bqIOVAD1w4CglWeczCXmzr2Egn1NRRFOkNyPLI53ULEsDw+umF6K5Aox5
Ksh+Pb8j01j5WnG7QnG2N53OBKm42cJPVBIKA4pJhDQpaSkWKUQpti8MYWITrN0Ww8Au2ElMtAl8
DYdsuTc1S3GrGX7oxAAJ4iTUGPKZ8Beq1yeeZ7nfCnTG4l31PFSKeCZERsa8xaoAlst3Qi0nz6Yc
Ldh1Xc/vkKHccFVUxJxZ6JEUw8AHHArh4iy7irR5T3Nj/E10ZZPTs08h04ZSN0e0B9vQGJ6eeiOT
MrO8Hy8PYzP9WAsNniG6jpK/mPWHDEtEXcGjhhca+JGA49S4EPwBeGIUVeHjHuJ0yMouMB2wL54L
VjgNA7k9gPTesVUWVBum44Kv2SV1F9aFXT648gRB9v1jClK5K0dAvA5p648gsS5Ntqj/JMRPDwnH
xE2AHR9FJq4/JLYe3nm7H+Y//AkHSoszkm/UfE6h9fDXGsKpkCUgjSnjJU6SSi/fo9OidmBtuc41
kzV3LpU7mjcyyOEx4NSGVyrnjeO9xNkd8mBu7vtX0E8qjpsaXmjAqQPkN1cZH8dYH5OHxXjZl9i6
ysqEYuFnFQrebIF6j/n6N7lnq50V9rM2CnZneWAL8Od/1PXBjdV4204EV7hKb3dmpVbkzOFL/9JY
NvRo8S8LeACcD2DYND37QyyFR3/HuYTYqvNrNyUR6MqnEIHJ9RqIZPOLkke/jy0d+XPi3Ffja8rf
LGCWnIc0Vqu6Z3wsApPl0nh+QmR3+U6QGJIZaVpRNe0+7Ky8R/OjXBxpuhLro5nmrmvNUv+D/8Uu
sicrgxGcgulyx3NXWy1Z03xTS1+C9t1h154gf9BLgk5ABkYJ32+kaQSXOS7jWkB+VUECXyNx44TE
8hdmdnK2Hw9wH7RyoU7n+B/efL4L+67Xt7RVJrJh/a6E0I6GMKnh8r+MknqHhyMYe2pNOyh9/7x2
H9PzY4pssS7Sy7StTEF09ZANyKVGQp2T6q8AOgihTAVGQ4+XBJX40rjDYi/w99tNE9UJzTX1VqGA
P9Eqc824JQTcSi38SxOPC6nE1Jkn1WF3/Mp2hC17M2hZd+AeMJ0fxsYKnHwiq1uoWmsKhj9oGldH
xq4FpGoXRxJ9NrPzluz2BieOt0x3CWkjSz6oDfSDSqSKOkMJlOdxDUyULgCBMhoaed+mhhnGyxAZ
2lZvbP2mbAfogpB4knnkPbbDF2wNleNI6P3D2C7E5glE4+gyV9I1IznQ9YWznI6NPFWrehHYpFp7
PY5KZi5DRCIW5oCw34G0qSbDwqTJXTPAbXFba2D0n5EDusYvmlZROkMUV9wmp49ICEy+w5x7B56p
DZcjQMS6Oi5CoMDqspfWJ8otBxEVXwyL7Dno30EFrhWXoObjaT7cIIZRom/fEPJ2jsYStxCQa/gq
cBeqrnzQ8MnyTMwK31SPENBPCbVhMBotiZfd2NOoKyRlEL96p+GNEkIzqPZ9FBj4urVG55nYY9FQ
0Tzc9INkTEk6iFgx1gNTYjJOV64oxEqLGGw9Mf8dptmP9VEl4v1fr0QX2G9SuDtDXBVTMYZjkuiK
BzkGRnNVwpl7gsUkGBqJNbP+c4d0cc3dkCC21xJfnxtvg4Cd7gRyZ1m7SUYxlg30wtZ23rMq41Dg
RUY34DDA9G8ek/pgob5pARGAzN7iXawfftUZS5DGe2qxlkoJAfsZp8DsPKAXqWMuJmXsDvMHV9kd
NbOYaQ/1CwS+VUftQ3Or1ELzDNeX3DFyYuBe6iTI8W41ECbLgV+Rv2MaGLGWSAU4xRQ8znSSrf0u
Q+i19FNgAuHr7xYDw5WzqSLlo9IN03gpBLgvsEgukgK7d1GgtVpdd9jKSfugptS7SWDeMfChqzBb
7aW7RpJVAGPNPTQ+9WPss3d2UbS8h9q73uM4gBA+bl45J2GsAKfLCM5Tpa9s7/xEsbMVSadWVqGO
zvISSSaOy2yPmeHeqRagupUqMkpVkJWgZtGWVwXNuznNY9WR0Z/+Gpa3/WPSOELzYq9ZQ2X6PFf5
tb+uj2ad/qgczB7ui3KPMqu6GEC31nkBvmyyd/ce5PHAd6s+RY0Z1u3NoIbL5QLs89OwaKMtyo+3
jiidZinuG55bZPftHTQw70dHhjHAxlEHYwGmP0n77e/z773USaOR2V5SVEscmJ15NfMIOfrBhnGO
C7/Je9Eak3RGcrl0QCNBPXHUHRGdgLjPhbUk5VMXqAVcXG7yijRNnjgHKLKgWZwLBux42f9y34Ha
DJd3lpphT5BJ2juppRirEZBooZzB0ttfKrEfNrXM24bc0R92f/io+eBSnzEf6OqbKE1TceGpbIpP
ub0Nf7dlENXoN4VBS9k2O22hVrfn0kamiyD1zkYv36Ode3wIXbX4lTnsfuT2bpt8J/qNrcB2FG7u
+myWjyQQRdHAKmaDFTlYFUh/6AJA5jjenOfKlcopSUw/lcwyLx9p2mCVqlLlYfKr/7ld0JxfSKSR
9qob5HyeTYwRIiJz9x8B4TkH3n1o3Z/N1/L4e3SzN1ZIN6wjOI4o3JFH/CBhgxcoJjwKzDMpa5ed
N3x/oGvEkF5chSsDKR3U+I7N2dHTt9jQMGMRyCnR5HzdDHfG5ettLRw809yhqcl4gu4lvLFrdf7r
jC4SAp5XnudaqfHsqJWuFN/im+x0Nd2rQ6tMGBN7XxdktXVAb9HiSvfLYNUDLJVmmbKUChYe7foF
EjTv3HxsSx76cCDekwzF38b+ZGGAgSXmpVa2mynUj0IF43C1C4NSTzOucBwpq2QXNQF6pWFdSx0H
u7wZcw7JGM21RY78ZdQKaMooLyhcQycTAF+DlkzO8QeGqeK/fwnorho1RlzoJQ+g/9HDYWTl2e1e
jai8Mr3OfkVCHrR4CLd3ArUOzMEBaIOKQx0Vl7OHwpEyfsMbG04udHVwCCNUaEpbpylSJs07t+yE
OAJRgd/fkCCb3amzKZdj9UQUJbzL1dDavqip6ijFO7EbTKLNTUwj8uZCqqc7JZcUcEHP0ZpTNm7t
Qqjk/gW2IBlFFgv2RVpXSksQa27Wg88ekA0Z2bXjH8neU2EDr0HR93png74Q0OFdAqm0/MWUcVLo
1+b7fcqWx1qZlRDGDq9bvVjERiDi6w3lj6ql0fXwQskF0EUKSqI9GZMrG+vGR2YCmWtStR78vRL+
udh7zRJ6y1/wrF8SuKlTLq+14rmi/xPmMMxxcaRvjDEqGGhjKVgqrAAYpthT4gdEPcuE9sU6gXuG
V3R7wwakJOO2b7AMMN7Tt0AUkooGrHoAbQWfTibOplHZKUgPakwuQTDkgUE1xAT7tXtuLxv5ehg1
GnTjMXJxT8hAsgnqxFBvpAy7F+on11UE5gjWbbgXse4B23m/lQZvWDelHawvzIiPekQUwA8PDXR2
dXSCQ+0oXjANSBhtA94ESvvAytpYtDbIcJSlA0QsM8dNKTkrQpdZk2BwzeBC/XimedNV+wsdDE6E
bA7sTnig3268LVlLdgeI8wTMVVQWLzM2E+HPK3htDSOCPSaTFWWLJXYsXQpxkrQgaJTZWVm2cblb
eqvTRgRYo3FRML5MF0vEHuqbztiYg5sU8+zqsgBhlSEgInEtwqzuHJmQLqkOcOR1FYlobEPS2qzf
Ym6ZSsuW1w3CPlnvRYujw4bAOBPPQP8QdVImmR2KAz6xljl73Bz3NYrX1zwCpW/ZABZlVytdm8lS
QeskKXbHkSlkXHxQ8+MXi+5EQWQ8zBN7J2M3K6GKyKDRaTs1cnYDnHJVjDp34Pl+Myfs6gEymFYY
eB5ahu9zbDBDqLan6JDQTTuo6yhEYcxhS1joAoqzQAng7qmUHSs0yFro+USVSmp/RrcscvKXEebz
G6OU64tXtd60XPbAndfh0pv7yUPFFOu3ZIpbOFyE0CVdjHz2aPUALXa9RnSVCmuv8Cbo2HjFj7V8
IXrQbNaT55/SiUj50H6Vi5WbkNg2aEs9LWrTHrLL8y52oR/MYSPvrJ+jqvkLEnSTcrioxs/ZDqrh
ay6RR98NvNefN1QQ9t34Ru38cSQL3NTYdPcheI3vLjy+WxnZBQFBDFk7/xvZLnkhJSJYuKv1s50H
u7UYvOjnTs7Q/KKRA7nrb455KHrHjDFlpRVm5zyaA/HdZ5ptz6oUbMoKu6PaeppgnmjsN4MDunj0
Th24SW56sAS7Ji28twMxM93tG4PbWqSBiOvNzogATM/hneRHjqx3AaWWM1eosKF2NT+CY/q+03pL
a4PDNQ0jIM3W04UMc0jZzBDtUuVIEeSQBuZC+b9gXBGbI4xv+G5htQzCafD6YQtCjtCIIgyacQA+
6RoKBPH48zz4aW6xhN6woP1KBcl1S2Kwuu3Jso97z1H+n+4QznAFbFHXXSyuZlZq7W44EDRwIDNK
bZEGJCmDL4CMaPbXzjrKXjgyDRd6IqXviFcoRqfCVrZv0E0lfyqi1vHZedptdziZLq5bFibtT1Y3
5yuW1lX0Sgx4ETvTFpLwunyZJnSL4FA4PxJ95jw6aG1KC71bXocpDz5yEIE1RcpJXZJwms6oEZJ0
q5hFnlup52SC7VNgPSN5SiPY6MgmyWfn1rriSZnDufdkQfXXooMaVOxBd5cZBamZwzlyPpeJ121d
N9LqQLiVePi80xHGHkASFUf/h1QAgrsm9615+YnLagn+im5BrnKv2BlmqT3p5kASHkQYawA4okK5
w7zVG5YPZCmi0RVBcUhguvzrWFLzoXnD3563JmWeqjcGO03jagiGBe1BkP4pMakBILjnK98ItQPf
w93/u7A7DNRkKdEzLViRi+AL+uP6yaFRKhYZY4YImcomsj/EAn/y7TfHzyPyMiuymq/yHaPIIArj
b5ny39OCqe/NFxJEjro77GRIDjL1zjqAX3SCj0omi8omwFsMPv/AEG3gWV0F+Pq07seS5IYZ7NHM
RAS6KbH3D0vvcQg1N29JGnl0exXb97jh0DgfR2H+UAFUkyCN4ITiK3XV4KXLAE0njuzG0TsYSGck
sKi99dkRm85ZyZ/Ih7e2G+nyL5vZTFcYw9k/jjwAEWHlIKlQHVFncaMW/0vAKRKenLtI3Vf/zsCk
Anxm/l29ULal++7vi00EJn/HurvcHQiOHCDSgPHx2eC1M/KZzucvNF7YzbqPX0B99OdL0rV9hhtG
Y/LmjCJYSv4B+mrcE9uYKSGilPowj4YUHjsprgj5jOG+pxufWrstvwDVfMLVZYkSBhkgzO+Cd/Zx
0JHbFkCHI0OOqXDBUe0biwYD0KDqU1vl21zzPKCwDZk6ZoPLpW8qaxby2UVmvLmZb12XzW6cDkYO
xjUmzDa8Iej7eSnWprPPg4H1/hnJ5f2wSQvNI1URk/Os3zcupZoQuXG5g5ojEkWA+S5M657TAzAi
VtaTMRIFW6LiuSmdEfvwwzvbD/n/GbU7veTfwHx4hpqhSsxUUNAVS6RjPvm3zvgawB1hTgxdtXJ0
vlXSqNe5ILt++8v4wWlKHWCSsRO01fOwBDr6KiX2qT9AzNYZC054fNzXhGwzKdb+zJyFsBqq/Dyk
M+x+ntDk0HpqRm/MbkPIKn5juuu6qjs72BmLkz7zG8i0rPsU+1Pu7V265VrLh5V6Md5pk4yBvL8k
CLeRLQbOyBJfgFsUFffwS55Sp/OmdqEvQwKFff8PhJ6mCzy76aNR31hzbgFJjqXOY8GuFnTF+mpw
ElaUqJ8weJI9p9DK8C1k1X+E7fi4OpFa/Wcx3qeLzohbNbGG1tOGDkQL8qHKfmlBhs+J/5QcxltM
pQqoBEgeW7iAvZ7m5NEoBNdFF0PPYz9gwoXJDergYdp8G265P7fS+u+D3mKiPm4DxwRtBZLzXrXe
6vnazmnxpB4w/ZFFcTzQYfOHXwnviae1XKBRNwXAoPLzRLTDQhrcV6Ytkmd5Wu9FLpCkiJahinkY
FaJ0aRNIVCC2Cg7p51qkhWzr7I1aE+IkTOS4h3qvk8dtwJTEDOvjmRFMZHhAJ58600VSW8FvQ7Ud
RKDLr5dzuo7ATR/EOdukK4MSfRluf5BIzt5bDGAMJCWubKsSK/aQwImIpgLGkvp/mO/5HXW91cT5
b0UM3duxWihPQqjte4x+Sa6MzXFBPOxjGoZP4oJSKTrjKgk6U8kgMtV0lqhFRQSMZooqhe0iERXl
VmA1d2fKVC5uYlWlVDbBjaWSNmd3CXkyJJw1NJNQUBz6EDEr4iNRJ0l2Sw6CjegYAZCh/vyHk4bD
h8gpi/FP48cKn9op6AIey84kY+hEg3LrAFmnmqwSqsv4IP2mw+8VbSShjq2HP7RliSuUuObzETg1
XxwVJ69TxOqglcQfi923/XlEMNr0fvBhDk7wvJ5TYCGfRnKtrGS0uc7hcDgBVbR8fZbwxIChNgc4
P0UPGeRxajvpds+dQPtxlHcsUC3NarOCyUIglWTLX53nL5Znpsso5BgZgCbEASYs8QUvXmggDwZZ
160BMis2LHKlNvtuSkxTpybN2tivlDFY3Tc+zihTjxq5Q5a9fS9vzhPp6pz9o6FLTwmfayfe844+
/H+EnrWBfswx4c+nSVNqBLteJKnNnJzFF7d5Srh9t3fcVpKT4xlcNq3bcg57dCHNY6fmEEVFaAbG
LjGHVKjjq5AV5nAykKIqArQ+GtURpuVo7gqkKTsartrFEX/KWOeLKhzoa+Va2FOobyBmjCq+3ap4
j/8Fa18NkJY8Z8ihj4VCEOjvZiaoMIz5rhE5kVNrrB9BYcYA1+KsrEOUQZVoddZ8CUFJNdooNYZj
q445vAE7/go2WbQj3XZ3rI57mZkUQKCHhgJ0fKrPOqhjTzYlu25ISTgPCuW+o1CEchMmPoWkRKHP
nJvQz++5WxlHah2tl3v+gW81uvdDVQY0okJsN3X6qMdVi/iOxe3fq4BFaMOyHRwIW/AS2y8faszw
pxzh7evso+HCYczdW1w5TttJFVzZKJHf0srDq80yW3umgmBKorcZzWuwWaTbHJXNDjebBl+VPASa
/4tgvrBwEiat2LZaT9i6VbeFA3JEtchotsynzd/WFU76RFO5DkGBOW9kPSRwNH7DGamA8BLMbf7i
d0e3vrjlJT3ss8T9rUORSkYrUaYra0bRvI/JElYme3AfB5q27tgHXXcAnTEnKCLEWW/Wbou6qzqW
VQQbtaG3mIoCVJR+mp3mcKZ7zsVtFEzLKz85yUOcaZYuP4jc2w55MUadVQeFJbtiNxnTlcUYTD7F
6uFleeQ2hf+i3EfXlYWXJ9vomRWWbmhgZ6x4fdE8TWGuxhWng/8sieHUsdBueYQ5ZH1soRsx0P3f
9qkP4FS1mm50TIxsoPnJ7lBZUjF0xkiqcMh46JdmcmarkSn6S4mLPZBq5WtLAT7HWd6EjwGECuDI
I+dpFOAEU4RjluFwu59zsdKzpZTis3szkGhk5DHAXRivirJbg5mIfip6TI0KTptxAr2GxRIAZfvn
LEFdPifoICLou9sOXwvGiILW57+hgtmOGDoFF9vTHf+Zt2bgJJc85Pe1qoxAd1+dtK5phfrwXsnL
+5ZoUWgSSzA5rhv17d1mAh/Oy2rcHjjuxbejS63MJrr608/cCNt0IvEfTskrdyPeCf5EZPseNbow
+M10Z5sAoHx+bAjS5pYg9FEOYaNdO3eByzhZhDJOVGoD/B+6L9c9/CNSItTY1cr/tfOhZcI8t/ZX
NYpoIRM9+iUi1cJ9ovxfeo+HWw+6Pqany8B6NdxKajufzauvMpG3VaG3S/P1NzK060G+xtkwV8+/
frQJrOHnYEw8uLY08swK3rA0NAEhARANaF/88q73d611wcgWAKy/+Ndl+l/ANdfxb8qc6VcJs40j
R1y+Id88BjoaDhVmGWLKxjA8aXA1cdYwfv6wYSnh22iPx+E14ewY0nS6+JZJpox5phe+ZX0me34j
0HrLgNYQIZmj47fwjWSPMOJguivNDwGs1TiLbPCZITDbkfHnmH4row0Kw8j5IHNTfpp9gCoB34Fa
NhR9y8viwJsQ824ryTqQ0apTxrxYbcQKsstQe96IR0f+hM0R5guLZU7QtFXhxDSySbjvnNEd8HjD
wybouySDl3XKJEMV8OnE3yy4IounnCm2NTP+0uTsdu9jAtGDnwTmhrmpMCuhhTsFKgpKTkbIktBf
mYEHYUg7sO9v7pSmZ9RwnXS1U0dTpgyzYcpC5VUT0qShQyb6x/d3Osh5l9UwB7IGq0kaqrwmYvhy
aenBNkwPxwFW4Vp+IiAFIiFMzve854dShxeyIr3Z2omNgNo6ZO9wYsbYvtEhrZhKYpDwV7V/qHbj
cZjMDAmxgKDdXiUqb4fQnmXXOVs3ZhVC9QgLQvaViD8ZxyjjdnGXGcA/7DpPeC72UvoP/h8SX/sd
d5VSAqnRKY/DyUxv9Kdwol+pxHf2MCaghohaPxLH4IMcc83T/Ect3zQ2VlrCPG0HhGifWuvuD8gN
9NPmMKPUKpCejGffhLYAQjzwKyjkba9Th5Nbcm1RmQOLDQBw32ZMOhGPoSQXqSN1cHKftBpcjoKj
VdXb0pn9etKce17eZVA/pLWGjNn+/LZwOxoHj0FiDChSJQErTo6OLo8ebOo8V04+fNEqxdyb+8TV
agfxOd7eOULeMytpukkxYF5Kac19DmrmO6+5hu1m7Efv7MpKEMX1A5APyVyOFVxttqBLBed9XE2h
4CSFFmtoM20+5uI4ek6EICt1E4NID8cWuBeWKkEj6dM1X+7gSNaC7FjG0MXmQ/gBuNAhGgQoUz39
ua8/fE+q7MyrXRhoUqFPvdheFr7OawuSKwVA7OjeXUf/ZgaXGMaxpFVhufC9m8W3Ih4IaSjE/Z6Q
2d9AUIkNxVaUPJ7TBDBkbnMEmAm5c95DEqbg56MsJY4oqQ/uAuZFGM5AySMtNDNNHQia4CcAMoCi
7waiGU6SywEBc6TIVjM7AGlfZ5qV8LSHr/pEM63XbKYgCTyEGtengebfAS2y+Sm93RuQ9JL3fE3Y
71WXV19ViBs8OOoOO0GYr9ORBp3GMg+1rLjxhaIxC9JgN8+GJ4A4NMWrI8MVBMMZSDsUWo31Vis5
Siked0CNWFQslHMVk8kYvJtsIvnPhBA0Brx+/0ZsWtvmX7N9/r3ZppJRSJ7wXb/+X6H3ri8B9Tqe
GZe3q/kBLvFE4r4V1T4/7XGfUqxtLTIqqa2TyXWLZ7JethqNVrSpxdfu6LfSuu96WDusa+4IesZo
gK196Py6Dviheqf4dhO5St/JgZx43drTUwuVJIEn6HH8CN7YsRoQITasiokf4m9npMP5uTA6+laj
+jUx625kziMJ2BEiSu+P7jJbj86k589HcuLDsDh6sB6ZT15Yq5BbbzuLUTXl6CWnbgPn50CK72Ga
lAWX3stL5bd7Cmra2HB6bTMcavZYQDvT0Ktb0uPEqbLbTdgOMJr9DnK5GdgU2cX8++7xDpQO/Fqh
LmTnrw78ykjkd498up4CzY1NhoYwLczljRETCLzNzH1EZ62WnsVVv0JHOb2Hpa8zmCDkqfvDxIRg
vBp5JJr0OyrAnFzeop+ZEOG4paHybITmd04+aOBztmBtB+Nhm8AY2bp+zmqsi4Mj1g3+Up9lvwBZ
mnTSyNNIHgsVInA5LKF26vD4UEkms2/LiXCGMdgMLq0xP2Y86Czr6NcG5q3ewwNm9C5IcJDE5vkk
vfQA7tCm93yYq0FbHRynM3C97EajnM6OBKsin0dscmh0GDInQ5U5w4TwhxmXrevfZ5k+2rxvZ6Zp
dfPWYvVeRuJFHCyeYe0ckm6MHuBY/1scaMn1RO0nc4cbdHNBKPATRBPSs86Lkk9dN1WEXJjLX2h/
vhbkY1qAzHxw69D+VGp5yAUA59bUWchrQrWVqEEulJYbNBK2iZJlQYiq+Az5vDy8IirbpRfGBPj5
uRhMUgqLmlYKEgatojbSgwryDcpsdd8qDu3yoKB5+84YDzUqaVRF/dgBC9cR+5R+dB4rchaokxPO
/nC2BmMhApj6Hn4TRnsmRyGuJpyYT+ZVD8XFc22etk1Em6WiCU1FA+ISlLfuOqrv4MIPtS0SZ5/5
fI1CC+/SVzZuJO5iRB61gTjtXpIRAwc3H/9VLU02RtEZNe8X5A+i8rWjZQsPgZZb0S5TDcYNngrz
4FPwog8jGMYUudgLJu82xrnRLTCqXuApSVnVAg2Tcdsyeq24YM2PZ48Xtm1GqViYJoHGbdRkQleg
5LfE6grPiimwXXxIBLGm1xvUQWv2JQIHxxCtqedX+arQGK3ixx0PdaJfFXzqiuvQ2hNRRAijsciw
HMDjIxvUEq9KNyw9NIqh2a6zCYNdbOuq1dmfDyV+1DR2d/mMfLO5voyky8EVkT+PNVUFFKmCn8Ez
SQHHkNnyBVM6UY2wejmkIExENWBORvA6ZLsB8UsNBi2La114qt/lvC5ZZdjw9pIpkpvN1OFxqWNi
tSM4Jfz78O4/NX6Sbo46qtgCwko3qsVGrFib4Md1KUhUyqR2VCYPuWoKw4VWW4fSIWeUAQvwJLuJ
8YLqxbDSDt0+zwE9TYcMAXenO8X6IISuuSAyPX1cOZH1lbXsAiA3tvuBlZh+FDdtIpGj3XPobpav
dCzkPCkoLxwkCQ6ZDpmDpy/NbFAir3Bt4r8kGWXP7l8ut5gWIxv5VOXjLVyPMMicr63xV4PilLuv
hS7ROWCoEKNIYKi1333PF78G7U+bmyKyvhSwHj6yMUYBQD4y0ODUL4bCGDhD2vzUju6aU8+KCbWC
7+v58G4g4mq4+GfhgNP1BrL+Orc29OtccBAkPxmV7groZPPqrWtW76A1Mp97/mD/BAtzDoz1kh+8
IHE/X1HRHXSrw0RICDmNfhuxHaI9Q9kURjDUVR8hasp4DcXkfF+bX4Rj0SlEfSz7mEAK493ARBt6
HsJqA/4gYS2A6gJre6Z5ZvHtd9MqF7eVEN68SNE5WJgoeo1gZNTDkRdtPh80MuTTgFKKfFglYpjw
DO1arSkrA/EK/65xQrYa8N8AINq6LvMuEhDZYG2besXBGCx1tsjRUVJqkSg7rZWAzpH82Od6rciD
Z6uwFT5nuuVaAbzHCvdMurQ9oCZRliR6dETW8XIjSQSxBP7BRopBDOXNfdpsVU4NDlAEyiFXtHT2
fYRZ84BltPkF/1vKPDylhSaQO4sABiadLW3aAvrIyz/dgXADLAyeGA14MWxDEECXx70sjOIRgQkA
lPCKJ+mBhQbvjBkw2qHPjqGtQCii4arFBbyqmIgwYSdW3sZ3bu/9r+fAPkYWvF33x4ZVs7bI+X30
TlUYwyNeZh5zPu1MECvDYc/lWWfCpYgv5SwwZOKC/Y2C4dMOeS6SIZno1vKqOb0CaxtfFTrQYgjW
U+iOS9S+LoJV9xZ3mFC1BpDb4RYXyR7pbgRypLCBfSg63H75dDvwt0pED9r983xuFgudwXMt5VZs
jFQxFYRinFnqV85h3uP3PzjK74CKlNxiiKLdZ0RZ8847k4Uy+mkUPN3O6Pvi2yNVh8aE+EV8xkeS
o5S9nMp0fnMQ8X1cr0jEAmVORHbcCvByzdfTtrv4Z4VyxdBn0fb8rYCNaepj9Rec1seW1M3NxMm5
jAOBnc/2BdqFgg/+UtwIjC+6U/JBCwyxMoTdGk09ykyWJLe0tjaS7NHlebIDoTF8PIQId0ZTorPG
BH0FeVyGnWQozX5wweB4Ehu00GhjJZ3hbqVA+Xq7beyq3IYGspnOSXezSF6I9TtvvYFrV5Tat94+
6EJ/69YVn5457nDS4Ly9LD2t5v+misBZFUr3tzDBtbWryt3GBZ33MFQXxPkQC1jxfjvTXy+0GU79
8DvOIhs4aJeaDPcs33CG1oU8WfJMpe8Z8a4Bhq9ibV3at4sjbyke86BULAKA1tQK04GZ9gA6viiy
Di/wH0QRsRcQiTt7Tj9e278WuIeE6g3SPeeGvDAZ8Gpxe4jxjmchVKOBWJ8w+vyeh/wFYQNubOeE
0iUmdi+TSAtOj7Xyp0XxL5rlT3t2FYja2+bfi3asrkzC8Vm64kU/1CpiGBdm6Re5M/Gr0PJu3N2l
CeClYn92mBhu0/2n8SxtotTtlzR5KMvqkIk73ZnBHWYX5nsuslqT35HSoFu8FE9e/jpbLRYOfK9y
+eeAuA6E8E8aKxbrFb7IOOavs72Oxy7M/IF23oPm5mayTf2UVxcjz63B/zEjpa44ileoGqmL3zVb
mT0RUVmwzKvP2FxL8pbLXttYYvBKAKvqC19/uFXAvik5GJ5tlGUCfv9r+XuoPKfvyYiYT6+xuGpU
A2TvMSvgrkkzhfL/wJYZkBjBicFiK8WtTVcUjbav61BDDoKN6CzmQhmskWzthGRvlNmikXPe3tax
nsuyPZMX2lrXNzyiuwX9eYgKMUQcnzKUHMtCRcTxR0TcvlkIIMblApbu1jpVkMA4FOX1BF2W7Pij
WN2tVdTpu+G03FqAMM/I8PZ7829UYNadCjsmOyqcV3ZfLUkoGNrOE/tcScb2XyINrFFrpFdeNLPa
8lkrzej2hyf4B1gb0o1JTk9Jh5f4n5BTkwasdxIKQEyAoITdipEdwRyDpNuAg41CW22kIRV52hLk
+oxjVFMuruoFeFJZzc9oDCJCo8pk4rjZGfucCbago7FQVo1zQMxthuyB45t5ZMImwgBw37SsK04H
FSOTo7swgAn0rj6YwE2i4IevBSJs22UOGavR2Y4kK9ppcDErdfnBUBpFAoGrvkSBTD4n1YKDb4Kr
BJzwly+O2sffjaJLHWl+orw3nzw2PxXwVhrgB1FBap/zuO/cJ1++8VNLOGdZVK2ZUaA1ZVEx1m+C
nsHB5xs+tboYcwl4ea42zo+hYyBk6vy24H++RESMfd3jm+wFcTvheETfpYyPl0DOMINdVUkMoAW2
abiPQ+FU/qr5D7Q2nR7T76Vrw8LbTvqYGqSdZm2Mw6tVDLxDazJBtKz4isWV+luDKGoyYB+nIm42
UkTeYX/ObGm9d9/Yt9AraCLMh+a166vFTlzeF7JUKgw8jFheD3eBB648Xc7VNlHXumxmi6sWO2fK
EGff6A9eyaKg7gKKkE1PZKJD/V9RM50YBPTx8p2vww8BUV1Hho1ssaB7iYOlP2oyhI/4P2UQ/KJR
cw5rqBdx434KMkk8rlM3echr9HPvDjfybHPzs6n0k1ALzn9/M7N8urKK17W/Gs/EZWUSRANsF2Xi
O3r/hD9Zv+ZyLWdDhgiwCvfckdbZDo07k0RY5qZN6UQHimV3BV6AXNG7WbfDYmnQQs292KbiX40V
vRMuoDRKI5S+c3YEmTVJCrtKHdoLtwZZ29UhCp30Cd1lIku3LLgDqlpdryo9hBfGTJ+43MWkbFTR
RF9AUadDzf0xEhR0JRylXk2yozobscwuAJ3K83/dlXYilkOqx5rOyRkB5msW1oK5s0+vRINaSJ2w
Zijb4ozyiTMHvwKSgodbc79Gv2bIXAqgwfRaMf/H5ucKzQNfk4cX44GZ/FdG/BQXY8UiFPhjFaa7
MzyFN9+iM9Uyr9p28cwkdXLrtR6pgE39r2tu1TdidKwDyWU7aEUKqeES0pPQI72/kIbYZ36/ao4x
TbAeBVASIxEoHBCFBHOg8oAuRIQc/9wJeRWQZAlibovwZVrpZV17lg+bsGqcBT0aMxd7mi6xn4/Q
zs9vxlqP0ybfE8ZflvyT6kJX5L0W5lBpD0L3Acw63or0cYJImwn9aE0jnLlz4cqyUh7X2Uqfdbe+
LmDlpGKJXwlBwpf5Ps09RufG9pJbjIidkhv2CQpUU3JkNnDs2UpEcbrqXipRgoy9eQfj0YN92BeP
irR3Ngk2HnEvByYvZ5GJSnovqqEf27oPEnqGjFx6O81rbrO9TgUEhufS/EXbn/bjF9q1OJaTaN0g
Wb9jA9wo6+4i3beMlT5mTPgmgNyRYEG2zeX7dYNZbN4qE/PJJemLHZ7phmxIlVQzeHfW17pwH8ni
z9uzjasxyMTvr4FUmhqsOoQiBV1vj5u1Vvs7AbASymX+gq+VQ19LkfUz30+xmz++A4Vc8x439G3A
GqkP0gZc0pztdx7dBrTYXss8/py4DTf8zMk6QKye5lO3IhxgRlguGPZGHqMGQsX/JRwvdCXn6cDF
tccUa5nMpM8GAOuOb4JEkDk2e+PfB3gsW9XNM30ONgQEtDRnalMHSoELWNiAKqntr+cfTU3k1/s/
/xxLkZelAao1le3iVBFz04qth1p/3TN+6TFiMzR30J7ryuKYfr/AScXOIhsmQ7gjvin2YTwUlRej
8ksrEXDDdH81PaUOII/v5Nv4lCf4TXxcs8o/LqkaarCnIwDOCEEK2iY/JNLMhO8tITtE1+P3iz+B
WCJfdvXalvZtUEtgNCDKloYjwx93IfwQkmeRrkxLsPCU1PiiVIrQS1mDuVVp4S81GKOQjVlDPyAx
JckfxAufise4p/qdHj5EUaT15z3buFW0JtzwNeyEPJbyqxEXL2cDdCC9p66tR/F+jIOCQtrYADy+
8f6wJwL/u8p5fcKgWAeAMZZ5THxOU/HbzHcgCXp8oVjXwpYs97bK9LHCaEjZlb4snU72YwLjAf/y
KFi++2Fz6J5Ltdxzpoq114CEe+fG4s/gDRzFVqT6TFQWnuDJtiIGTPaXL5wQt0ggs0+5Ke82koee
TgLi0t5vlGGLBV7cuZV9uJyiJZauhUl6oxeLuPTeJT9PMs7cTCvH4SBAK+QGhZPoEL8gUmDT4XoN
WBKp7Uhhj797S4JoujYWaOXYjXCrihHPG9TE+pavtkf2+giLldsQVkAjID/V/QyOMz4RVUDYGHDB
uz+GEWAH7gFlL3hjQSUwrxmK/DxsYRyBteB1EfVaOkrgpckT+FmpljV54m6o+U67Q+BwcyAxg2KZ
C8Or2Sp8LPPUi4Wbq80EQIT7cYpx3V3vWkxtH3JXRTrLrKxpdE3DCPNuBUrX7pe3O4jIcXAkZVlT
ZI4QGXTV+/pHVKW3Fmte/oTVYA+ramimhtk3ggmu/NMs5wO2a70BYMBnkNc6p6gx5l+Rf0pqIemM
IQ6CDfUEN3oviK1jhUUapbCGGvscX+F2X5Uocy1BzkKMrY/wwPPb4IlV/3ajHo3keEwBm6yI5Xoy
QR1gA3CG6BJuM8c/HH/oyliaeHgwmeBNDigyeqJ8SeQE88x9+TVaaZDy8gyZ3yYJLQtnFM5lkosP
Zho8T1tYYM81EId5EAnvKXVWbE2pq3Zvjhs9f033C1EEOZ9yzkTtkOpwMJE0ex1lhTt3yGACGHnC
agrXRRwd6T4VtFi7oxoVCztO6HevSlRvgVE75Q+zbtOhLOW0zKQ0Z3qUNFMamMUR+9ovFs12r20j
AvWAHfHZX3PK6emQ+oEr24fo29PFcy0MMk43OgNMVbtmGvH3EHYjv563jkZtvAWWvysfpHbYXB9A
QU7NXPXJVGrAX5IPU0vpExzumSkCehJGdX8F2BM8wXMSD4GfS7bAO9+fxa28aikquw6gLcE3OFTu
6pXq3CO5ZZOIZa9vv8+B3Tnet9AiZ8gXLviVLtRIy20qIetmYfhzxb/Hq9cRh1ICF9nCA6MlEhBi
YJKUMx7HhMP3nF6Z7iz+WXMbGDXdRedJMmszfJ487ShYzLwoZyrU18yTGVOnlZsBu84o+if0eP/J
ZlCCNSXLnaYhls8/+hAwDRxOt/sjoFVOqJi7slzV35HJIyvUgSAURyP7hpp1884nwY7Elx/Qisub
Dl0qdbp4ucT2lOR6Rxx07D917CH2cxYNpniLdg9kp9e07qnQY2sY8smZGvYeBu8fM1X6jpHbM0U8
l7IdTrNe013rBmf+5MkzV8ItBcri/QzJa0PWC3VqZmC77x6s+tcVjmu+3xzdha47zjLSITCPCmTC
L0VxxtAD3GZ932sCs/Tz2Lf+3uNTZKIRphBPJUE+I2e2It6cUkXbfGflRHTZzedmJRvtbS6nSkJ7
2LDwk5zWiISoK5cmpt6kti8kGfTwEYLM9B1CdWgu2yNzABa5WOWo1rTHc2PzZiW5Z36Lo9XajsGR
8lsDoQXBG9rHzcFlbkuDhfgiZ3PeUPVE7zaDqmMTgERHYDAcPM9u0y2ElpDcNUeZ3N9Kkqpw01du
IpAV6T8e3jmLzGmtPD4qdv8DTYqlkV7jbIzbsfZr9U/gBZQTgGmZhHETBExw/0K+aSd3mkvBqaNT
bOnP6WHtexiQzA8YhCRNinZgaUQUfGcqa27qeFGY9hD8988oI4u5Tu/+MLrEC73iHYV7Iyzxu4a7
Q2NRP2Gl/pMs85k6OH0V5HJw1c9mjb1ubgEeL6FsnBWd4TWxlOoXgkfX6jDnfT6tPnDL7abxQmHQ
wiOB5spKvetgOlhq7wL60RbEsogZuEYZycSYjqTsp+ZoGsmiMprkL51l6UeC1+2/U5qfpev9zdKs
0ZVherwikUFTvqRdQd6BIM104Wim7ed7JoQ3olXz3nsciPJ4cL3Smh6zY2upuapXjLR3g8nYRGQU
8GvyfX5uwJsjg9KIafEgZzm0aUUa7jKOs2oZqpGFC+C/bH9df+9ITTIvoF0N3B+EBaftVQA85Mg9
JsHCYLtiHubTJCLyzpRIU5lzBy3Aaor3pkEkoF37mra8McEPPyXOspAxo3L/mB5hCsVV6gEPDbkx
UHMIfjSI3WiRsFZiPJ6TSjYFpSHGxZiBnpMFkLmiylL8AED5vHZ16n8vVAJdzp3104kB/A8TBSBU
l1JKEKjDDM3Ni6NeASQYCJEhXxtAGxcpq+zgQWjw/1/J4gfyrO04md6tVpMsZhDTzrUgFedZlliB
ACCXZ7d5edzto5PstGzqdFmVbhdi5JNNIcjQvDeyZOSeea7UHoW+E1XYqOztV4Y+4XQuF6WoV+ja
tR5S7hHwl18X9z8VlvxQykXuO3j9xESOPn8dzrR7beX/dBu/zALHvueMPcH9CHiliQHwNA3KWeSs
wsmXcUJB+jQ0mEihHeCceUrtCJ0ZvJThrBJAaF1wytNPkdR5txdwtuSKhvTrhM3OWXum/6BDk9TV
08ZDT+oCsQWBSnz3aKpvjp/KUt7QcBZF/lFD+lBB7hht0Uc92yy6DfoEeUpTUHvd+AzNABeVdcOo
zyrEBu6sJtQFgGw77DDGHTozzrJZUakO6DOUC9z65W1hOIg1NWgBnVrIC8aPg3kcIwmRE6VsCDA/
zXwwfhu1WPcR+QvYi5NO8IIC/s32STinMeb1F1k4QIYA19dYbyie1miWsgQY3MBzxfBUF8w7f0ls
WHOqlUpT0MqJNe8D72iP3oLea1sRSGJkB8U1hVUONJfqtqEZ5g08trUcAq4aEcMqifGyZ8L3yxAq
3lldoIW0WvzQ3mcDjm6FlZtSsQVJLRHheybL0/LPHwp0RNhhLnoalXj9ZKRSYxLEH/pUS2zrfqxZ
L3btieKA70fWPL72Ve6uw7nT0XviVKsUWA9MV+WjZ7Z9cmevb9NPn4c9IgDZnKuNOQLkiQB0resn
IxuADH6wtQE4YDKHlfdeQdtwPjEWOYvtZ5dYRlwoCoMxPzr9zjkm9XHuy28uwWH85dxvo5I2lSlK
1KgMIorojbBbhCk/cw/JSu84wd3+c2On4mh5WmRkA0NsrWSp6dFbOs4qxACmfjXPD5CWmgFaBPMs
9/byFQalXQDphUGeETIwUGVMm6AQOIPLkP9rPR4LFEi5o+CuEWnvDr2P/fHRMMAJQn3eIAFV4NJ0
fYG2cU2rpJr0as+o9438OhbkbhQtGhudmhNbsWLeRc3yox+3qaBkrdVUigf6TQYT1fffltjpyS46
yukJI+rp/+8rcOnN8hud2Q49nvlRsISasSzIqAueseP0h5u58jMvwCJoJy/X27xP+W/LJ7SKWurz
yeEZ/fbjQF++KtYXAa/+UcWxJIBCrov34SAGexVEBYJIp5pqdHLAKaKyXqJauT8n9IbyOx8XUClt
yyPRVUMWpJGfSF1Rues4AP1NqFPEv3MCVQN7WglnEMvkb0/AnV9IGH83Sy+9b4fHXDN2p+eZE9IU
ZWEbWyt2uNV9kqoTUuq8PL3ciJbAgmlWfEY/o4vd6T0RmoOUh7mE+NB0jJwNABhv1soh2YFtrms1
6Sal8TOyqJdtqNmmGucBy/W3qLRe4TGYCKlZIyrCo5qCwkC9Y+sf3mp9qI8gTkT098cy8dQxCzAR
iIF48Z+ZCmWuNcOYV/0m0zDnK4ECMLdGn/jC+f9vYs04Urtmgg0zQiqf2XTqX5R7QyrLSiAsPbzV
achyIxH2S8hBezitCjXZ3YC6Qux6HfcqSkavMZHVkpx4HqWmdmk6KLSD4pP3yenVaXrEGxM+g5Dc
BAA5cbxtL5/7S7eUxmg7puItodlOo29Z2XmYJDSKoBWpqf2UyrprY5HZ8oIfq3hiKhEk6hRRKbpT
ssHfeWWrkR0rJ3I9wAAFdoZc+SoDjn/q8Dk28uKv0b+1HtM9XDrCZ+GI4KNXn86m1pbvnRsAl5j+
JmJDFf/mgm3QQI7hpVrCz+vkCtjlj0SzPXF15gLHcjCl+EcdKyYEx/o2bAZ+l7Z87FDU4/ZJnrCq
UgHJ/ulYIbAplzicTeaz2wIWGmrIZtk5xTH57GllrzMBj+Y3HCTT67e8DfWDMR5Oxb/0dWUJa5kH
ixOWfrgIgLjDgugDU/Vav8Tsh/CV42XL/x8sXRkbilY9kZVOnWGJ3huO6AK7uHZyh6nhBm1rE7JD
6aMrWFVBWzqCQki5rGIffDST0yRhByx4T6a12IAHxnFQBPqj0aBqC/sbIWpLK1ieTRTCV+TChNvC
9OKNBGFVw7OHNk/BYtjmlB2nf2wZfwcHUQ10k0vT8StizQX23TDqdA3qTewxuvshcNLFAIj76GEJ
T99SB9PYUn9KUEg2+rQR3AELJ1D04DHWt/79loH9D5LRQkUnb5SxjjmwerZxz2h9gwPjy77Gk/IB
tF6WFrr4Eaf2Cw8vXIfNvEt1U/GCDSbHzUeuhB6shsbF/9xEPBTZOJvwP+1klRR6Y7JmntfPKZa0
NNrsjpnSVbJRW2V3UyeblxJxrxEPBCuAPS2j7V5CRRTo6DT6HBFDXn+YKf1j9QJnv2TyH/MQ5RLV
uUzTIvagmJkQVg3SyjVjHgqiq8q5XbLei1+3bp6y5zbAYhCEKhchCGNS1L+6+5dIK92OUekp+nIP
P5sfhq/i/v0z4fV/p/LNqmBXs0r36PuzZEqC+X/BCKaFA4gLNc9mn12PoO9Z0piB6EA1Mxz9CPlA
NkEgjryEfgMfJkip/X4ugwN7XMRxd4jwyqyVQQFOZIi9zyocjoW0DFAqA1zQUu66dEeWxGFDTner
SC8DuFGqtDGqvIcMmPvHfJcszqzkD82KD/bjonkrTmpMf/4UaVTfOSWJ9HzomQGmXz1H7TlruUIX
5BllIDa106jU9Yg5zeoGCduYEkAPz1RG/Q8msPP496kvqLxPW37OykxqYMd0asQ+Ols1+fB4yBeo
6Q5P0gNuKQFMkXllDpSGl51i37vSmhpn9RC624hxKmgYk4GdkF0AJ2Fmf7tqjzNNR6eLwOTPLv6z
97tYRBhXl+PFXa9koIqYgHM86JfPq2fw/NXWU4rr9XH2eIR/Qp4A3cqPLQd9APRj6YLcq6U8hg7h
t9BoCXeRE7vxMcn2WydgbHcV2N0/3dbjEtrRJWfQfn9rsJ3zLzTODNW4dFNAKSFkQApehPL57m8n
XRzHvzv9eM+UL7sAAjdXYGoJmXzR6v8vyLQ99qFcd4EeZfgVptk9pKG9PX0XY19W0tZFyCIc0Fsu
buSA3JbBF1yoTj30AGRL5pKHbKEyEIfh0vV707QcKYnt44CR6CQWn/uGuLu5TvWBDfffHOMGT7l7
ngDo/k9kmuzAJvW2xiFXwsrY6R/gSH+8Aj1bWKTz3tVCHXH1cly/FfyBaA+Hp5I0YQ1Zo32MKc/R
6j4kQ/K3Pxu7xLx+Md0FNb/sgZ1ZKe5l6E2m5hvDIaEVNJ0/aFnrM+Ub4mJQafsBDNU0CSwMpsnm
RkjR5La8xiwThn8dzcUpEQVY54z0eDOC6HGJz/sentQ1juHc84p6iktT8lr3VfCwpw0eZVFf3+pP
tH4xtIN2DzcTM0Fx9dkvsJGbI8Nou3AK1kMVNWgRMzJ4//teb7Q/B8S46vtn1whAxiblELRq8luI
yjF4qmkt5GY0zVlgCDnSJT96+Gk+u8qmnGZUEYfaT5EBz9UvYE4MWvgVjOSlLWq1OvcJDGYiSNuR
mU6daZz0iLNGmhACfIQ5gKDkdVYwFEaFt6FdrJK25EbfCXaYa+uo//cI2zfdtBTZqFF9VK4z7h31
kgL6bMvMNG0ts7rZPyBXDZCcah2LEQto3+INz5mI64rYERshXqo9rbaVCSrj6wwXbByJbu2woYnA
KgNmUzoekEnZJFT3QLD6XSPciokOukUeW3oUF0Ms47VIl0aECwB87GbC3VHS29cI/WT4K5lMsdbK
APLOXAGRzccWGCux9DWsY8gd+RURrGBn1/xN2zzfT+agYqUkA14Xt80qIkBZn9hjT7bjfrBHcVoE
xFU+ghPTlztaf3E/ueb1+LSfG18AiUw/3R5Am1iDnuphpAFGWsq2doqiCL910B44JzWWZ/p5OXtB
gQDfmOBxxzSdr8vI/Uh0OExA8jy5mfQa+KNauUAObOKia+APxEzZAnnvwBM3fgDSUGdHCDZgW7ga
PWtd5HdnvhMpDMqnF3UXd30AkiZNfZYzPioP7jk/3lrflvD/ctQMgCho/NgjBXkTIH8Q/ZxfqSaw
hVd/EX9MpCVUKxv4+FYp+znPOH1/9fcMzCkcchCF0JZJ0TJ1/54ZKmnAEK1zXpO8IHvn4SbVeTva
nz/qWhnC9xVA6vp4mhb1Pg1odnslPaYnczuXxWn0UznmyZ5zlE5aUHTXEnBrZQUFp5+zDmta5Q3h
/fHB8VLIrcqaog2UYRDwNKOdgVvgqT9y2APunIJ41+9juHcsutOB1mD7PZ58+6FSY3fobYmBM1W5
sMszyzuCD5Yg2bObnJhjGPVGWgIfEDSXC50+ne5qx6914lBXeI0Pw2MqWiB8XnOZ2VspJnqJDwqX
mZA1eaLVoiYjXL5dcyICu8JT8Ot6OyHvVHduMddnKqo5AbLqHGID+jug90stoA2w6GOtSHN0QbgO
sQCOtrxwfXH69DXGD3zHvDAvWB5m+zfB8uNceyi3G85s4nSPLk/EvgILp/cr/74KlF6kAB3V6GVr
9ubygS6wMmRL9M0CSv+DiJV/YHHY59BugqetWDC0oVUZBqr1NYB2CeXXzUJyagKc5NbpBbRcvY1E
bRpEaqUNrxB4VI1PfgQAg8VoYJDlMg8QSzlbdiEuTHMWPyNxF8O5w5C255PbIYd0G4zveHEbmcUR
IGMtLTliDwPH5ePUkIVjwCxn4cuAbiJJRCCT6WpoA/WrS97g1f8ncW/nR3r8VrU33PaQZIhBDiRX
3hsNDX/xSJaVcaUUVCdzoGJd7Y9Qfo3fFI3wPna8TvkNqkhhSHdM97c1/w0t6XD/SGPq35wATTlb
eDC7QH30uHxVzTjgC4ZzxxDOqmyUbbm/37Xmdd6YjESqoD1xRCV7CvX1CKjD1py7xu+QG6VzR7Dl
aKoY8rhwB+4/6WVuAOyEF0ocZwSPIydPIgcX6VXr9XlG4zUUzMEJ+i36cOjD6LhnrynXju3nzxe2
McKxs3/rrBYZM+JegBQ+DcuM4vizPNfGpubW4j21OpHnGQrtjHSDIQYHXBxBUlWRNpNdN2ilEx2o
Pb5/vEpLMUsowC0EejGdaoTdF+h3h4VuBnkgXcf9IVYBRcbz71F631vPUDtDyFp7IAwVq0Egm4v4
NU/gVg1t5c00jRKpwL9qn5GzTQSPw2YHaJHofhJIINGqaNIjlwCpbsr+ERvA+ZmAjMR+V1bs/Mtr
5YG2+t6YPSORw9zSG1hQHiT3wJbLYV4EQmecK/EcIRAewcC9rXTgqKYu0/joDUwBGFalPLSVb3sK
Lm7M0KpCTPc4C5B98NFKpIMMtDsJvHyr2B1eJPOy9G7SJqxfFkUlaUcbEqFDuGjS+oMWXJkJP6vv
+/yNlthUcMX0ifwpy4azefSWu+RRvZSt/QHgM960xickcHoNqda6wmUGMsGRBxo7nKBV6tUNkt/j
32ae9AeuIuyjUY/q9HP4gV7Z3mQeSUQ01NssfOud5hSICTXJd8VIdxfrU0c6FiA3oHi5nMsV55UK
MqfBVPvdXzHJD6aTH/PLrjzi4Le0M7MvHSrdpmKVho7yO/cvy0RIiI5q+5sPICWdoGZS2MKDbIeA
NYm0spgz9KsFhA76z7DuQF976OybKzNR1o3yuVfvhYptJ6AjOeM7vo2BIBYvK3n6yMT5DBpJfU/r
YaL/8vRvMi+R2/A/gpNkrVXvKZky2DA84dxRgElmYIrFqpFiRLRg2spci9/bPXigYfKKjd1QK2PJ
PxaGF3gM7n5spOr7iKdMtEMdk2+qqgdN/DX4W75/0RCbcBgbyAfH5J7pr5MR4XZrAEcIQnGbZaqg
PvMHoqVyKsqww/sEcq9oQNNHIvOwuLbd8JBX88Z0CtIxaHkg7kJSUQRe5LKYD6Ef7DhjnEViOSGS
i1xUnZZ8n0V8zGw+RBNmtmMMpFwblRhhtUA0T+1+1DMXJ05URGUsHlbtrHRYSu7xI/K50Oe33U00
+NIekJmRfA+82W/C3OR0nF+fHFPCV8CYQAXCxzM0Zc1Ac12uhOxnYbmxInFAW+KZeCIbjQCCJTlS
v5d71JW/uD+u8Bj0Ng5qquDNnLICq9tuh23J2rXRBse082nwWHWEsam18XZAE3i6MyEjXlkAg8gk
XNIRoew7tMKutVuhWKaz0k/H9AbRAgr5BR+8B7HREVnKldn/kZjzUE1cXKYSZmGmipjCNN72GUba
HCsZ1mrboTCAgyyKvuhAEhgWYl4phOYEhKqu8BAmAtEle66TuOm67iIf7W96elYoVFq9rEhPimOR
6QFbwhNyXarEqxZJbshsAk5kEEImRcOZGrH53q9t3LvBZiOohX09JiQb5v6yoirdG0MVVinFn9YG
/OG2aoqcsCA4yhkl418ACSp7PB3vYEHBQ7vZbEUcOatit5Q0fH+ktmAkyKqJ8zaCZRWWdEqfsYGH
vSlva8znkQVxpAeShp6kRc0uNjwxdbIcp8SYaYV1AqdiuaWtc5tsLZqmoOweJMRNrsL1mX5O/wqb
oZ4oQ/k9CaDPDHYVHiEsypUkPAVNzVPWwsdo5XgqhVR2VyWFCsTrezLWPKi3n33tHIDlfWQWQXpp
H6FrHT/umMhP40MEkHtxgm5ub8NHNOeGlLoWp2f84rhD/jzs0pG3Z2HtsQRUw1JFA1PfdNc98/WA
uNPwjsKDH8D93ukgeTGiCZU863BI3sx8IFr7e7fYDyND1an2110uzg4e/o2MYqWeS+278R86WhOV
hyiPcTDOwiCFCUQ1yoMNWmYsqcMpERgTSPgCuL4JGaKNWfjMR+sgmNIobs1Oj4kMb3sXxlCddnVd
GrtgWhq7GjBnBWu8T8LvfKHD7Q8frFpWJp51zB31KxHHKjcB6pyzc5ensoth05Cjr/miCK9yz7kz
wk2vJI3k6PnFRxEUpADJUt/MEPREcdbBKOAk5Rrkq+0Io/bWQ8CQLx2dG6w4LHdUcKMQtz8U5lXK
s+cHl/afEz/RlYWMsbsHUVJdrZjqqbetBKvErYNZMj1bLeJofhBKyNPIwiZZO+x4NieLIwuqvUbd
bzUv6B3orurw4SuZaJhtERjWtdixeOxbndWvSSJ9OwBpIrheo+fbr6DqjXAG+WJQIuyLiAuR06Gu
MJxeFuhRyG/l0Y+uwTJWKoEGH6OIDAlAEe3u9J2iN8CzNRDKxd3+oFV2WY3HOTiaRCU4jpssSpYU
l/yTul+DHnQWCsYN/Iv2zFVhFMmAM9ZfdSUA8jSOpw8CX1dfJXSmMg1Cisgn+Z0VkShvzlipnASb
IGCECAn9W3axmTYrPn88Ctiu3kgdrq+grmtjrexaXRuEOlFX9WVXaG7Mkw8R+oOLW9fxpsPyy2lK
eNDX5bYGR5A1b90EbJs9BvWaoau92eXZJwXuSNHgY8qqcudNCND3B4yk+Xwid97YKN+WfQg+fi8Y
yoVn3GxizF3AP6VvZMuf7RcLRyisH1OsCrH56ZutKXL8H66nps0rLFFcjSAudkmi5KB78ySuEjlD
Y8tJ++JWSGbqrohTpsCtjMBfCOxe/4rassH0Gkz21tOWaMZBD1zZ1BYKaWoj5H2g61n2WJWb8la3
tdP1Xyr9tI+fUVQefO8k5271e9HWx1DrJYjOSXOELlTgEwc0D85JxjwI5qcvLv8FnNuEPyqInZyl
ugIqVZmLntbNH5sseKgB+WWkDYqGcELBSsSY10SFuYZnR9Z2UbuBQOMk189HFxnBCjLlAThNOqbC
/RBLS64in8uB7o3ufb6Nas323xGaAbay6W+VCFsFQPEuhETRhH1vlT5rZkpOVNtPEVjB7RujUenL
mohVKO1IKzRVAlmOkZU5QhJPoZGyRVGD0L9eLzWyWG+lY5f3YibTDjCPwaNJgrvwSNZWs3KtPMmQ
wLALVeYAR2IPsvSOxes32cZWwTJ8Te6+oBK3D7cOTAElRLDZWNC90PVssQ5muXvVB2FtuV6OjsSN
5P9fF3q6ufzdlCjGiQg1ofbzCT+IMFRGj8L25vW+59+2UtuMWQVnOl+nRrgHEb3WsXs0tEBMnh6W
i+/JLOOKiFl9YEecENY9r01bhFvRnzJvYvXVU1buMo9g9zuUaZ8tYaXtF4FmNfxZmmFDTJKeqPNQ
45izLTqDmxyHOvF9e2hF+y4YXyY/KGWsSqkqz4O6XOz6lYBCxkOTxLoYbXwj/EEOA8mbR3TS85DB
ddBcqmEkHinZkWmXuV31nHU36MZjCCOXg+BWZJPFDTmcSGgePIhrrY+wBedisvScxRe2sXfEOsdm
+zYtUq9Z2/tJNkUwvl2iIpaKAKEcwguO90vJ5KA6kU2prRXr6DKWVKvxPY2pBYhUpDkOvUY3ShLw
i9V0osN2hEKWRZhO61vXDOWkmnSK3W6C6DQhoX4gILjzO6L/8ldqUyxAslt2S4g3G/iHYomc248r
QMaLbJ8U1Hd8PBpW4y5Rx8MiMcVI4LvhVZJJEv+jFlfmlIeazsVukj9Fkhpmt7clscy/Wr2idbVY
nfFP/IduPilnyJ3BmCKExHuEnCpRzNYeQXEIlqcRS5Pi4wuoPlSheag/4HZicDKA6cYao5BIzL2s
1UEPU7Z0gNOmGzcYIiWysha+M+6xYYLCIkiF6TSuI/Q50sRPgWK3zXlZrU6eC2rdQqlDM3uuGQ1H
Ty672i60X4XToK2Ump/mh/AsUnlAsXWnLQTKAJjbvEVmZzuWIFBLKiW1hTukfK8V8lD/UJ3pIkAC
LFwhm0LIl/5tkW7SF4hoNLLCsf8ttI/u+0MhH3sEgN21cfvr++mHDc3fFgCjxzxzn189tVbh92HL
iVKoweFtUzMN5PeT7KbnZtgAmbKBHfFpC2YK8Uhq6rWnfoa9AtPKegpdK+y6xQUxyvONiQ5L+0t5
OVUsEAiymI4Td5je1EnoJ1SIWuIZyDTMPVXeiEjuwr+J6wVdg8IL8KR9cFhSoYkfzBDfX/wodd5l
ZiphUl3+9p4RXoKQDxlKBcz9w9lIuuMSQsg3YQRQqPEPt9ICBUWNAjFzDG7s/t5FvQxGL5phjmZx
f+pZ9gXhza1ZAtr4bVr3lYKnE4KsUw5QP/K2M3Zk4ZmWutOIqeTSFUDWDmJ2sChFNj3oAikYI/mo
E+ikGePjUknG+i3DGK3HDhOCMayJLXsgMdijxSb0Qv7AtHuqwrBIzohlK0M5krAjWyrmM+rqlPQA
ydPScCVyuNYhnoiBpUok0y6UGMKEeBgWhtlNynYKPGKRX7qmF6kWEu4x5eeWHRRDCOsPtYNg73jP
U+JpNYn+AAR7yZLRSxFxgB4beyQIDU2vuw6+bqVCvItIVhMQtxYiSX90gFHyb3zFIRdXpCswGa6C
GFZp6ypM5nARx2gQCIxbIXUHazYz3whziJ7EyxDvaBvvq2oNCUKPc3Odh/jATMisj9E35q1LnJiE
bEqQRX/l+5TqIH0P0ygds+HsNF9kKhtHl+9zlCUVj9fbIQ2rqiBt2mS2g05Q+Y5UzKUazfD1xcYf
rK5+UBemnJRUJZ+I2vNT0Ggf9qqeZ8w/A+ABNX84F7xBCqNEPYVzgH5dyKLqZ+m6mKe7r9Jgo5pI
isAUrkjspG21aYQD42QB/s6U7nEqJwGlRb/1Q8rZ/tWfjtOV/wwly33YjTqeU10cBNn6eubeIWet
/NCHvUq7mzPyyGdo7FCrPrby7N/AGCqBfB3SfOTwUvvc7LFRedjGiJQ68R44BPYdWp/LnfivZy9L
CoVrQfoJaw7WlkrVihUOffP5zyEMgV5u8KhWuCpC/QtqwCBXImmb05IR9ZlWiAaPov5wGxg1XJFt
2eUGAPFr5/e3QwicnObQVbZWWOYbXdmJ5WbbzNgorFi4i13U8I2ccXqw3NR3LsVLkuMIwabUbYlg
wc+ALGDFOoxe4qoh9CMc633SbthYm7sKH5pqmbux7iUq01u6f7KNYF8Jrlrcrd4bNsxFHYhZ85mx
Y4eBClnL8cFxfbOaQtLezYEM++VB2RApK7RVrelra3JVRQeM95T5ph7KZshk/W58/N/xboOK73LK
yA9ITHdSjwf8iG+w0Qb4iq9YWmrk/B+nTLOcYnDOOiJTb3xSajBXMEcmTVyCUcFyVQECBgA4+vuX
fHFu1Wdjg43nqxGpb2aOyTDxWy8rFo5J9Ok6OlngcDedplTBXN/V/m1qCbV4I/pszAVONAKnaCwb
BO2o/LsT/V7QbS5vk+NBbAmsJWKb35EAClzn0AVt8WJV1CB10/Aop58aJwVFvBmA84OlPhP+aDbX
dqxMPHebhc00MvQeeC2WITc3eYNbilNWv2Ootq+LohqJc1OYRR+SmNfjKbzpFXdjeY0gRc6lobYg
3dwL0Ph5m+wQdb2lgLs0fflxdSxKJ4xPpfH8925HBWyz0eMDCR9JzEnZ3hzLIAShaiWYOdkVSjeZ
zb9M0Wnn5K8zGev9pe4StnOp9jhlApOCPihqbSGxQYWqXVGCr9ggifd1f+Sr8SRH6dtoLFU00Roy
E7v/tQDjirHcX+uYtyB3sSXAR6o5Tq3yRMZcGXg9lfbHpPPQB4b+fE+d56ehaKbMQpQYhB6V+UKf
gQx8icXp1icjDjx+8CBdCtQ1TPGOjWkf92HHlBQ2MrKx1PZgXdrYUBb3r2wfKQhEwgkZ56L1Q7VH
2H94tzic+WqoP2wuNE+u2f1RZQ/2bDkowmepjElFCcOq3zK585/kMJ5jYGTUSECWYcUF3wuwiA9F
xQEKiIZK3EVId2XOe3FF5h0ekt/OEN4QLhkl3vG656kQN58FFjd6iPSluYxr6+Cj5nfOsNm3Udhk
YJVNlo7W8IjlqogyEt0QBJ3GvcApqy3vmolGidByP2XbUvuBnEo5nkmt/J4d4cgg+knZQX7f/WyK
wGNGei2PgcPObNL9LuqwnsmXBjEjTOWAO8GwZODrzCQOUNfzEsuEUTHJc7A1gFYI2uwPlllgGbAf
Jnwfmrv2B8sfZlBxpa8+l+pHS2g8AvLtqYHkA8eH62gndOtB1coQqrdfdWF00X77OS2CytC+La7K
QowchJwUg4GwWmvREczkZjN5EhQpnG+ut0FwxDDRjK6agYWovHxn77Ttxe1ok9+CHx/wdIMn3fen
YYAHK/nbFZVOqf2zAIm6PjcV0DJ4gvQZh5ARwTrqIjwgPR0aaIfJL8cYI5Q+LK/Hs0rW8J5IwUTb
SUGYTeohCeMGD4wGkwWAPFg7zrOX4XkcKZi/4DnAYbyy5lGwnGPAa2MUSSvib+tN9VCRCwhaFeA8
l2o8Sogd5MZnukEvlYySlF+I7QbP+F5ecubqXyC6K96J4W4Ei2ej2CLCPS6pyyJPBHVlmSyu3r89
EpB1X18IfzdUh7KxgHeB62GpxAzTAuHIcrbp/aKlMmprhfEwdxh4HOPZZ6YwgoRfnPbkvwCEdMsg
Z/tlK87bFkUA+truybQO2EK3tJ7Fj9E6JFJvNNUvfcrFMn9csYHxIfANhQPky1aMxqY3bgfmjPqH
Vl42pDLOAfM9pdkcTX3yzxn9c6e5SUjOsz3Xb1UTT0D+YI4tAjZhJWOFcpT80x+sI4wMYWpzV9Qp
CcKkCRFx5fLwv6tzKEwVFYEFXGnTgW++qs1oOYV3k5oYCBJtzx+jpnBnVXb8leL4iwPnZu+Qo+oQ
FlSC3ws9SiXr+JrKgXdOj+XBnBHx1RWgVOOCk/EXS5Cg13ZCGUNoR3FjaHOCtGCM6rYnLQ8l6XMJ
p8IiF8KC/ZvMB/V5SYnAQ9u27+FDTFnzT7aqB2fwB+GNFDRTgsrfGwb87Nb/JnQN1w/igNq0NnEd
MH6KH9UosvxKEBXLf0aYm6UcCFtUvpp5zIW2/f/Wh32O4k3VcFgK19A10xAkZG06trl6bPZ176JZ
hB9qju+preHSjFJE4taPAaXCMPruqcJW4AzLVktXGD4cFRGP+AZnkrF8cxGg/MzD5VoX8EnfP+1c
tkXLha7idHUIx9a7TwuzaIAgx0S5yFZR04NkV5tsTWo5dc1GTgKMrSiHXk86CcIBIfloO9UySQ/d
dub55jKu7Vkc24buJVthb1A4PkIdBgqZXOmvYti+IJ8GFtaRDDPwIiHerbSMmBflSfFDc/xulWBy
H1dCIUOyDMNICQc5gNU0PjsVU5pKAYsMBZt2weUuogItt0XxBPaCAr037/n+gfX/qSwOLg6bE47d
e0XL4ePBOSQFPvd1oYm2W5c6mcUiuYWv8NZiUf1WDVqZ4qYGqWve0Y7PLvjDdNkJVCTxfEK8Y29U
iyc8GhXD4kmOakuKoLcKCUU0VhSnMhm5fueBmzw0cnrZ1D7j1yV8t/vlYugiMjyiRb3dR/iO5Qcr
KFJBM8MEz1pXT95sO+agVCAUlvTljzEAT6T9RT1PJe+7aBSQ9Yeyh9S2iI36RsDUlq/OzX6ql3+r
VhQZkMddCk/0DNarHF4b2nkBD6jwrb1xDAp3NN5uSsVqGGL1UMh8dDSWb05WMEFoPIOF7duWlmSV
qiI66R9UprEzulg8VIvOXyuL7oYtPv7eNuBUrwXDukYeYIwSLqeYZIOFsYy2qgZtc3Q/eF8UB4jP
4LsT+7UsFE5PT05YoZDJlpzlyxZF+TcWW8s8DqJCUvGDI1pUISk1AfPEQSmZWlTN2v/pcB64e1bW
eQS1vHavs1Ot4DOkU4J+KYzwkREdA4Dc/YqvH6+EsPgXKD1M28YS/VI8gnGx6lVKA3epzLD/Km6P
wFG/Gwbbu6aQYFBCtnQQ/CvBYgNIGMBeIoeXeOtsJVJIeEmhdDgQMNqjM1W5QtadjmG1+0RQ6Vp2
4Ay4n2QaTuLFB9XEJJxXTHlz7lg0gAJzSvqt/xr5Rt+8Q/j9V/ViWllgm7DUZ/02FucBXjA8ijck
zrwvhWT0pj2YyXE4cy/9lZ1OhpjREKtGEBM7Wmws7fsk6Rof42KBPOYXGtAZODkwacgldNjK0aZU
bKUNXYIj9Zwxh+Ptok5E4WKZw8zgiSYpzAvsjSm1gj9seou1iS3KP7cEoQSRurMCwg8L76d8aFXM
ZrCLxGZYpHAmik3aZH+VF6ro+yiu1P27Go8CUXkS3xKUg6QQARPTBMfK9BYCrnKyuCrSa0AvCX5+
CTIanV4O2rah2xjhgrnW+T7ClU4ee5EukEJGWACoZ26Hjo1Gy3/NI0NTU0XR5Um/1jyuGx0jyFF6
pjzkk3NEVDACvlvCrT9puMXkjrFVTfbVaQL9Kvdzy4X9l1SiTuL4O5XvPGz5Ozm2TiHO8Z/csGEe
nbK+yYkpyBfhhcA1+pUKTmSa8ZssLkA0Kzw9sOZWhzq5emnCoW25YIsw+KZjVyhaRAUQPabFqzNL
Xon+3gC9BW/Nmn8s52hVHCahoiqCyA16AwvSI8asuC3vY+Qtd//4NxBHcBYblwJZPdqkOCRbQAEC
3rrVlAYsjgnZfZuhUkQr/O9eVXc1+IBmmY15tz4oDegiJVfG6sQVCQlWMpKDBF4fpXeE1KJHePjm
Hz/0QqyX9NvO9t/ZLQABcUAiaT34Tft8WEvPaaLv6o7VGMdJpV5PSrfDAXo8rSIKG5urMQcf6NXN
QM6HpqIIgi0fWUbWWIfTBl4BlWhlxm07hVXSsFVU5kMel2a6tuAPq0EvrbN8+KF/py4p3wXxqSbg
0/fNi4fV9GTZXrSbUlOEtj63AHO00sWn5vDHtUv/jplm4QL8UI3GyyQtyxSbQJQ9Fn72zjZD5pxh
MvMOSVB9SquPqyzPr7/V96PcfK9hFeXOb8RTeyIf62z/UoGN0lOo0wjcn1RbUFcLNmVRK2iF0upi
dWk3UIdGtqMOtKuKAG95qSQNhYssW8S7YW9pW41OefHBod5/o8dGWCAocCDIRSEsdDLm18N/JB/D
Xi37FxKUiaDL6+04ZAl+W3jk7tS0bj1IeYrDem628wK2Y4/ZxevqHhq954F7BLihaDZuAcKqOoqM
/UwJHojuCewsQyJih7KZ6EPVU1dMm4VKHg3y0zW9/5qgNUzJaDyFX0f5Ey5riFfq4crOurobycxB
TQKSVvuE+UCTVvQpTjg/gf3TxWk55fwPP9CQhve+c9CcyK2XOfNnYhchPP8jd40rzbQjb3vUtkrl
jMl++LkGrd7rQf4U/6NkEAz8Rh5VDDIBvVIuKqJvis6qEWvpLPRJGdR1dt3IWkOA0E/gKW0JXXTh
p9d3tjQ+ZXPwM1MBkm+SLPV05rfHGF9XIr5hIYfCyLxzbWB7ZklksWX+6LYRur/T2H9LUhE3kYc9
zPEW9CZJP+qV/VMfKfIW+a8t56WvCS7JPog/qlkiydKiFYg5mnPPkxzD/+P74YHe0gohwB9I8gUD
GVTzA/fSiTJ80/lgvy0bVphh2PYqXIOL2hUX7zlPkafMn8i6vQ0MeLnofj9qK8eIsRmBRqFz2nZ1
1tE4tEMQjsjGVzbl01KcyoePk2t7CxfYmTUXCzoc8MYqLuaJQYxPZH07/Rce4ZduD/UkWzv30UU5
cPGdGJSBGObfldEyetK3h86q6iT0WCwdPuNtSOjQ0wsm/EmYwiR9pbnct4ZReGpkHV1PUrGkFc+j
2aX+NivNZSCi5SF193AO/dFZXbx7W/pwcJZKoSGR6grGAziv9miIzwecg04vfKi0iOlmmFcMDSrn
6u7p2Dn1H8OSB8htT2qoCx9g3u2RoygvgVUDNvBFgF6LTZKwbwr6IGXeiXKhqh5NEz9euPbE4l0g
627/PSeyenjSxVVAi0Ls9GxbIMC6t29Lf1KM419sGLZ/EgD0rJ4UpYdmm6v3i/xKpBs6mRq/Yryk
UauwWUxpuHSE90qm7iUIwzzCyttEVr7MQriNQik8SaVj5tX3+kMGnWJbb4iDQHp5XhozP7wREEla
/PNS2EVh9LLUqiWm9VSN2EarGdOU8e8Hb2cQ8Fbi7Xn3V0Yq9n2omVC+iPbkOAk/YizMRFn4crH+
VV6j4NFyLGWYRo7qAUA9nQF01+OTc2JCNKw9Gfa/DcazZjyZOPvip85bWmYIF0pnNkXLvg3l4sSd
S8QdQKkVVyTWj2cIQ/0YwJ7SKYiycUZ9Dl50m7XrfH+DnqmXs1LiX/BxgZ8IfPKgKcZZwnCGxYIb
qfPuw41Wa5BEm3iMcK6OKiWMNSSgXlPYAklxmyNLqOfSe8Yjpn6FKjRQ22IGiWje6HvFXnc6Vods
3RbEXxxKdQVrmFEUIjJrPxxscpKahsWKsaycoyaupe9ND4A/3oVp8JudVK8la2ZbDZMoDv97CgNa
EcuGqpGX68d3k7+vfmRZAObiNIfRaRTXgE8yFb6V9wVYJKiIhkFzy6esn704u8pjOkRAMdiM33zo
+BR7UHKToaNlZ6TlPpQniYrah+aUrSlViCDUvBmPCfbsto4z4LY3wqVYwyTT+J3QOmhOJPYHta1X
QZ/7Q1VpHsMbAKcRwQqNcg7fRqyqhRiqNda//oRjwcgROspomD9rVy0AUVQJXGFqQ2EewMIorGGw
gUgb5tFGCRhTjT+zllx7RevIHhzsu4wu6T1B10qArv8dxBe9+wGNUMaJkfXTcSKc2EqgjhisDCzv
LForQPtVHGAYDU69T7ETrQq7Xt90FqcbapFzhtRUyjRdOUDdc9U+opHYv0uI5Mv9/Fmv8X/3/zMm
3lTaC9CZExhxzKy+2ukG6ZKna85suE63Bt3cT8jeXBW4bM/Sm7o1FHA6oLJeMUkz1xIBtXGeWDf2
SrVrdATTSdhqEFfnoPhG9gI/Hb3SlBdPVEZ7a5EOVixcC8xxX5css090dSfbwjA6X5qqCzYcJX0t
M2JA/nfjqej9xeKPo+hjnZM+FcXX52SalxdoviYn7bniwXrJMr5crtDp4ax/pZpOwjC86CfqhVXy
j7Nld3uM8Bc4AzPjC2YoxxEJePh/fo3R7kzv5IyCj3nHZBGtBYv1uZqlnDLkR0hjmKOhxEedhPZi
0go/ngahwNXeHj5OyrVnh5vyLO01dedJcYfNIOyPlPANeghEVKdN8d+oy3TuvNz5QesAICvvQqsJ
Ux/UQqKgF19tFqQ2RiTPgnLiLTuSuHMNYMalemyIanSfnKjiSVEHu17wT7uh6nPkucDC13oQTKAY
6ZbCzlYBqxrR+LiylGoVs2jH3v9u8j7coTN6gNU+c6iVhXR1K2UHceygVX62vEr+pjv51zFWOigS
US9d0EyzQE8qLk9B4GhB02jNuSBqqnL1j0YENGfECs9rfocbJNRS/QNyzwzaY1ECDoyTECRgwhNA
MPoAp8iGn8nGRyxDYPQC3Ie2q8hs13QwkNTybFYZCJ/qD+OJ0hpHSpDNAKgqlWjPPsRgAotCExpM
5fWU2zQEcNA6fKeZtgkeNKpdeuDEivuU6Mpf07X5sd6wAZjuzQfu6kJqGked8SdkVwLd+4Gw/NfE
a+/90oKOx18B3U791rnkUaQIVjULfd1MfZqbMdJDNgsGKfgfWCLbiAZESN/BcMGEp6aeWfk3nl+w
n6CirDAzFd3Pn9dwyCou+VzMAl4rwDCqHa4ZO98QSkWTH2LfVhlfa7QNdG+9WgzqFlynKkKN4l3h
R+alP2w3aI3R/0dHqkFVyNd1x/MmtKhN0H00WiZMH1vghJRCjPyABdoXFVnQAv5S8iDeEbk1srPp
jKDXiLkyeDE7KK/eVCzDssGfh/nA4aiZCOC7rIr2zpbSTiU8AjTMttHTlmcnMsHig5zX0r7l3vsG
VO1JMvxVs2DgEmrMRag7iBwHFrly2xu8/6wwXxgo5NII7UiBKz/mV9W3N8zXf3176VdvAiW4pot3
4CBd/AzV5macNioygUMz/40+cIptoiqAkMpbtIxCRjLJSB90o8mFNQdXkg6n0/qkP0pV3KeUDTFj
ZRpEHxXiHHNeWjJOd4bTlMhgKPrAcEKQuqna2LWJvE1uyNABqZ/5cvOzAHnvK/W2mb7g51CiVCaX
pxYZdcYRmUQf8sF6VR7UocyGobRppv96nte3HMneWcHAcOmRRpsEnDC6Lz6Z5BRMVw8MxfZORGpX
kWCkNIiHDkny3xqrG5R5zevKhqpeDITAx76QWChe0PsJf6AdGpmLuKvqcvpZxwaTqVVbWJ97rnbX
Uy3H81gyWFhoWDrePu+5QSoNTl8s/H5DDxcGmDwwy0JcpR0N4udr0xv3lCQJFgwiplL0lAf1YzaS
BRX8lQavGnk+01naPi91JrOE3VB5WeewpNS++TNrsGE16ev56ZawGYO9+uo+Rh3Dq3Mpzr8U511w
69T3sctWUhKqcWBRdnPWqQGfSlApeskaWcq9it5OaP3PaSVTjSE/F2h9vYGn3/jzU5FiESCDQRGT
/U8yjguNTY/HgXbG/2Gmp69schg0M4Brs+qwfEHcOIxfLuKT8xcTqxadgUOa8UOfvyCed9T5Swct
mzYesGx/lEL6rxjem88MvPHJP78rRNcBb3EivoKFsA6zlr0d5kxskZOSTSvRuyksmTuobDd+YhWl
6IicSkd3BF1MYC0Vnxac8rRQXLjq5HRH7W4Yrc9VUhHFPyXUJk1TosnmTmc+NLISb7R2EPKrlwR8
+jzCuonwwFHL2JybS29c3v9SpMMNqTv8Dwx3U/bLew+Ow4MQdmazMbg+j3AUkI3a3AbTlQoO/Mt1
p8orHGccvBV8klgklgSprQTaGficY7AZ6UaxThfV1NaUaS87wOuCO/Qc/YbBhcPzKh+4NyTYFopE
TJAgHeITsHLU785u5xT0Db7EaZ+BT6XftTJHAXa3bX5KTu45gVk16Wk2qQu3WxURXlUphIppxOXE
VQx5j8/7C5Kso7Eu9n2v6hGmYu+LW6UiSwtco0y2SBizaao3m59lQDwnfiacfbQ18flEvioYTFG4
d5mnYsNHg5BkeJlXSdckRZFv6FI3cKpW7/+8jqXmV61N+uXYMql8I/t3hvWBxNEi7FUeWW7KSfyw
BfGQi+CTpzvpG57m31BmgWb/nTTxz4NmyI594TDZ3GIt//bUfhu6TMuPaCVQZLw6ISssQzzDaEPR
gIvHLsEJnpmgjQE8G9P1XWhTtdV7vn1wyHt0Q2Jf8ctxD/zl0Etzba2PoxhU2b4kqqSn5qFjsDTz
xYkDyq5JBo7hX9Ug5jdiIREEJ+oQ0i8oLFvbcMuYzyLHVRq0F8p08hjySrOFIEHdqTFaLycDkCf2
RT/SX33+kRntrFMD8VDPO9aHuFckbZhrFCt3Ep8tO7KoPOEW9+tdGGMaw6+NhwBrL8gwlqA20zzm
QBs5vm0XXrenbO9uE/FTI5nC5pYlUtpUt432Xs9J7eGxpck1lJbx/gm6WC1uZcmH7nD5SgkuG0nY
IZlRFElXbI+fARfJ8wzhg/8LSSVR7pwR9hkwyvgqPkU99rSPE22n8koH+bGVsDhxAexNe1u1z4FX
E9+AbQbF0YR0hKhHcPKpatVWvUNf7575eyxhRcP7vV3joxhInoR0uD+XkrtNh0guhFK2SzKM/6uF
0vNdhXKmFdtFw+qxFgcjBi2Xn5z+JKhhbdAdkQ+aWtb4J5EaaGqFGGVU2MNr5HpjEwLb2gVqXEme
PO5JP7TUD7ZgD/ybZoGDC6YnIoY7Hykev68smDEHKBOdRSIwKAlmIqhijHjTfrPvSMT1ErGM2IHw
J5mnZg7vkiAm9Bj9yFkh9Ut1DKan5KK6qxNZEGHcALz7/DtQ391nwTdA+0auiw86ADvUjRwU3mmI
79nJ0qWHaPzuaC31w4s06WrKd/0QDBVVWPBIHgVhvPp0s78KMC6vSGXKXY5tD6MoUqtT58Qr44I8
TEfW7Ditk7sPXA25mTFcV5aF5chL5sJJaoPxi2m7KFDR6aRey8vZKUp1LNEUUgpAAlZjdEhADo3D
HCM0qJkUjvNOgKzIFonDXWhVDrX08s4J//FiyMTaLHdD0ptHpi6/3y691BRbBIEYImdVTpM+OhBy
cm2c4N3Zv96ogtaMlXznOvLBcMi2qB+J3Anc6uso+6ImvMZBohse+WA9rnIS2c8yDSpSsOkwOYWN
8TPMaUau6p34eGUws+AyqmoTV5ylJZIBZTwxZi6woClmpUg1ot5SY48yn0ZOfXGvxFoemLRPr5jG
yPf82qm4VBs3PygqZv9Ez1xOvFQIqUjRvcKGnml/rXzo1LJLnRwxnyPkk0TZZRGb7lnzB10aivFs
bCgjh9+Z9scD6qmABA46vHayS2Ep/seXb2vY+gewT9ObZNjcwDXkJn0+H+mS5f4ig6RRE0mKgv9g
92ywGowXggv/04o0y/ZwJhDrTPbbuk+eZMHJdAlgFdlZx2xB6liD/ANMDakEOFQLISnNTyc3UXhE
U/ZPSHauGIMqITBIGjct57MJzUjDvSDyquWSRjVBU8m8OwDhVOQdj2r89PpHxtpzmvXxaOCVnMr/
pAdGif5HcY1PgEHn3BU1KuNqRsp9nfUISCLpKDlddQXngBPWK6dCNHdan+/tx87crVLDECwx2rJa
LewxDYs15dtoAOVq9RfXa5+mgr34ZlaFTN0GCh4JHUwb+rE8mQPwrVihc8cE8w1zH8gsebsh8iaE
Kpz99667NgvoG9y63Ypo5uJNFExnzaZ31Y6eJ/2CfszhCoyaWg+XOKE4BYR7nu8g1WT7RpVJB2Ao
ynQUhZyBs/DXRPJ+4eBiUbKxS2yYepoQBVilIdmshKvbbgTUyynPACL5PhkFBpw085hqcT/re2Xf
2kpgfA9CB3lO604AbOr0s4zQ4GCJBk5sOMG9MnLG+3Qq+tyvJf80xeg2mukIPi+QALaKJDVRMMuU
7T0CNE1ejirjOtVUG8OQG/XAvcKmQH+FB8x0XgkkrDF6USggQAtJVL5MQvsWSH5hwBKnedduILc4
0UYNFiMASicmV0KFJSh3MCWSGwZ+SwaXOTQ/xOQizxGu7rIci+XXVmgG0T+RGsN1XUL0Zf2XFVr3
gODGJjStxVPtWVFdNffxJTyoudsPJFlNOXKqZAhkjkYv4wXjLdwOy6hKZvavuUuk3Ma0jKZmoqlI
A1rsOwYv5PANQqNoBk+Ipp8ej34E4qE+nbS9/AjHfXPsDbgEjoVrD9kWnflMEfXksyhW73B8sGf9
JQrb8uCELYubnfztw6ycmfNThSLYBhprJ58IchpVnbignTs54SPYqkZ6nVVJUB8dnvdI7buHY2Eh
biyE+3h5c+GKjNEucYFP+Q3DZ4D7DpF3UetH43L+uEBxgZIiJcz7jI16zUYOiuZgDxdeGzcxhOyH
R+HWwo/ZIvBRBTd1jWume1OQql82udUFLPDIaXVIQtB5LTryS8hM4lUMpFMDD4a2dZZY9TjsfjqE
bXAMNTR7BRQ7EZmkxMly7sYc7UKvp8gW6/85iaLzYIGVloJaIr/CFWNBTYvYL7xc0H93sjACeLFo
GNrjPkRROUoxEjlNuQ6pNr19Z4IYalrPPCicnw+WHhpv+CdPUNWH+k2RTntiL2ZetNmCYKX0lJj+
Jyoii8gwcA/rhz+eyMAED2zHK3lMmlpvlQdruj5kvf//IhGZ2aGWWH6UbyUnRxusFHEm1hKJ8yO1
gYTqt1kl9vucqRiODPYh+gWFLBoRqtR7tVitR5K5TjphAVp4wx1KBupbSgY6Jkr6WNQAtVV4jOK6
vdCxgVO/ER85/aMk6BT+bR8QBCG7ZXN2LG+EKlwNHTqydBHqyuINJZl9JWj1YmNgBUbkP9fbCPNM
BWw5ce+zyjcOyO6pbfuCNHnod9NWFyzqR48mbPHyU/wkwg41NBi88IFJgu70rTvEUb3h5VwlF71n
hr9pqWQ+ApNo1m6F5idvEUK6/wNnIRtQwsQ6zmuEanMZ3nBnfYfvoPiy2j9+QulIqGEajDgVq1cN
xuRfrCOnvnJkmZ41WfFyRkLfVTwQDrxXMt8dcGPq3aEJ8gTDquxMaFlfdqtb/btBf+rkaD422Avv
kvJF3TrRepcpMydt5OHbG6HwC13XyNI1nVPfZv2u8VLR3mBLGARJGWRbFffcYeEgGHEi8AzVlOW6
PCt9J8wQ9wMEDaPzGs8ZsannBGC0kqcaXYduMCen7SiTPkL5zj57Vbk8ZvMna/nQA2MEAzGvnhV/
9tEfET/TTfXIkMDwJt/yYGYmqtYHRlSZDnnS6Mq2qmWrdD2XY7PGqDZjx4QMEbD+6hUuWu6kJJ/2
nfH96jfP955J53P1xL0XL+DZqNYS2BfVKt2WAgdvJtHXlIX0mQgWH24nbyqMmZOzjVfN7lMr0IDu
R4PfktfSjy0s1FVwSCmaap/40PrkJKzRhaQO4Lmj71sY8HhO2zWqRd5L44TSJh3B0kOssZjccqQk
m06sZX82fykvgOMNHI240nvaUHoXZqQxH0do+nlKHsImz2GX9l197gfcj3SdoVh6kL0vtkcGBAKl
9TNehVbNlAMHs76FB3HR9QtcqQqjA1HJvN/YtRVBIsQuglnvo6wnJ6PSQyZHGuvMtS3djiab+/md
rU/fZVALtKnSDaLyzgepumTI3tbfylLQ6W0Iiok/lvxlYmKOyJjeQM/w5+pfv78gKO4W+C6X0L+M
j4kJSYf2joYGLl9qh1rNadLhmUoSemjBWbCPFB+9HnUUAJnvCydpzGp8xJVkVP8NXaxAk6FRcaF3
V0Wht9ZLfzxCensnKqd7CZOZRVAV+wf0XMI3q93pTB7QPB+3ahEjzXXTeGe6UDcnmpuZ8391Jcuf
mQwhC4QTFv/q1w4ViYVG0rbFVYnP2KWwuv61xkO1ZrU1vgHUPGhDZ82ciLta2tkQkPvc+JIMFiPO
HDN6MWKRd61zTPhTzdHhgFFKqvLUyq2xgHZJo8nN52XVebhlliV1x9yZhF37PVMT80+yTd4qGFiZ
eq9lVI9mXFOJQEyYxfvwHxL92m0Y/qNQzCBaNjLmIFsbJpQYnF3M1Pavq3YgT+48Bgedk69W2CIm
ozJw287NoLUl7eZiSi2Qc8MO+d9xXxDak+v9iLLK6iKOdbbSKryCaln3Au/BK78B5gjM6xQE2ctl
gx+mtEOV4KJyolRN3dRIKiH3ssOqM0m6L5AT8Zp+G52VfsyeD8g4DcrCfApNdK9yZvsjlMqcr2Oy
wxB6lP+xvXIkQUPmzuxr47lJPToRZ8BZblFZBiFo7mUg9sWGs48C7yHMkAHUNbN5/2QczZoIJy4K
ZNYa6hxwO80IUBaz7JKn5OZd+7xcTEW0dinSuSaUdTQEMu3k6SfhxvjibotVbcr3RS7H74gWkYbR
GUk0REuMT0kVEvHvfusXxeCWml9MpsuG33qPS51fxV5Lo+KUzS9yGoInkaAgEDBQ531czBWdEXFy
2k4jF4Drfe5PYylJjYpSJQIiDPL7gW+KzbrcLdSG/0fmej433rNhCLG+bOSj9ZRJ5iP1/1y2HE6i
bJR1p9zZ3WA6qbcgewVz9i6dCsSerM0o+0itKZaXaDzyBgJnQ0VgWf+45yawDEpLLN0298/qgFn2
nhKd8FiIeCMHrPq0I7BRrGD2sr64SlcFs51u83ROn1bo0PZa9pT4zT1CcXxQk9iQlneoOucwAPG3
3kL3U+3VSOVtwig0Mz9uF08QX3WPZlfwCt34du2qye2+1R49xoSQIlwMaZzcTE8oUNmeWS0Gkj+c
VpC1eZwgEdSfu2AiFto4BCTtz0Hg7O1IXoTKaoUIR6zjowwfolq/KVY8SgWK+Y0ZuEQgZGvdxMgN
rX/Ab52ecDAnmYAVbesrMLQp/c7BSn6Iv52Wkyh/dKScGXkPjJ13YW3ZmKSc4d1mLw+FZj9YrWcb
lHSIM21aEbOeCrdwdRINQLRf05MlcFh0ZlE7vq1qQQXkCOds6gvODgx4R6fehc6BUEyq0ztFNCkB
41rjoJduX1FXHQWJGtHdm8WRLsaA6M/ZLk7F1BecZRPYk4d89OobS8kMDmOdx5oH+Qqz8PGsbB8z
kXb8gK92yqbH+d43oS5b1Vwmiq+M7qCyZkScXEPknyyZ5rzQITg2F8oMb5YI193ghIBZ7uok6C4N
YKgwjP0rDvudBdLKDfSeJAHI9t4/daAIOnzARzbQgPKEFjsajUZp3Cn0rXbWMnBM1/92U5r5jyEA
1reMQoftodBhhP2CME1CxB52SsCsRQbcogEOQVoRbDbEFAqKpQyVOGUO/CvEWzu6oXTPcOxjhshd
arkzKT0zg9L+cxZd5rCjSwT7yRVnzM6Ccf3oWILM6LC5Hh9Yv5zGN2pb/XneN4kXsvfBkStf15oV
W+egJZlMEF3K5EFWB5UROmZPJSb8kCmZl8wp9hzcdRVDEOYzcYldL8x+c7WnuGMvDfOaw7KC/FHZ
yQjNFR/38xNv3EwVYtdF9p9njE33MTYIS9CJo38lANnmUcLnBYZ6mFIhTSbnjxtyta8QkXFGPDkG
H4Eao39cqM4zbGVBYOOSlxgXj0UPHsW+8qnJhjk63RRTzTvtKnydhXxSeEmLagKM0gZ4xFfW/GEh
fP91FP8hKQrmy5hbaq9VFuglPz0lB52kzOoCUC/Jnbw+QAac8kZ4rj2uUbLeLG4LkAmOFt3+hhlN
ba9BumVIp90zCrmDFBpnRZzGnR2jSQSQ/a0RC2z9rQL1lxJXmhkEMzSMdD+aMg//7kqNUhuWUibC
AYj9X5BNumuH4qTo34SyxPrTUdbqTn6ID2mXFaiKU4jJLCM/RIEPnNLURPfwSIuq2LGWrAeyOJcH
224DqCQu1C/2SdGbthiL/OsDXwjfkqYCBxpTcPL2le3mNDrYneYy5U0dYa7Gkgi5DNaXLPxc2qlp
ioGYpWvMTAHBAdIr6fjAugKRyFYhE6/MCFl/Fz1jvYFJr3BLPc9w+r3Zby2uFMLGFBZNWbL8hfCv
z+2O1BXsRW/7upW3iW2JUGZDldFzi3XTkGx6bNdqqY9ZS9z5ihJ+x/6XsqGYGguYLljU8ZcB2bcC
r1/AxFhp9IzQ8o/DlzVOFkoM5lu91tEk0bkAmkhnCSmAx6F0BSsI3htSE/imxUV+K4mR0YybbsZh
/AsxN4FHQPZg9FkbvI9oIce+A5jOCry5GYUkSwxSnuttbnVU77bXMFJ9ppBlCUEjaw/V4RXekE2H
KAsp5/w+Xa+MC9xGjarnswGkdOuo0SfV/45ncGh+PZcMeFURvOhojrlbmSmaioQFHr6QOtiIgrpq
BZpr9fRt89vCrTyLua7VhMTEAXmffqM69N+YbTQA+hZXCAotUGwvHiEtul4O6BSTd0qDUTQ/GVen
b9KXZA+2OyEYeTZSoaZFCaZaJkoibDWeqll9GU5anwuepaMVpWaXo6D+RvXXZC3iVHo4ghepZPQm
WjMCGdHv7oatl3kqNUJCtlwuoO4uVlditQPDdYuJdvBxdHZ1ldKE7paecXW3IwxcHPoQw/ozjcym
GiWMZW07HaLcLKODIhUqQojQQ7jTaIaa8XOqaVvoefTR84uFQ9uR5IaK79D0QmAZ0hWEHcv0soyA
mRp422mvJBtC5WTDUEwnnjPqv3JAw2wvrEu3D+nvivZncjIygC9qxALPS9+WpqUrYusAO5zVQPcb
dBJbybLk4FGnrPHn0/jvM+R9PjO7xQ7P2NRHU1cR3o/ZC3gGUJiP1avZEcioc8y6CIombVjOkYQ2
xem0Mju1c9IFSDa4XSehqJZI8any4jtYIPpJ7st0xM0J/NJHWIpzuEDL3tuspa/O5N+BUUpAPg7Z
MgU2cscgu1jPsiBCAVJlvCDHpUCG7G5EGTJj8nvqLFci5iq6uHT/vorRyKL7eJu+qDnvwq3U+zzF
Bw0yut36UL26eHKjyctPX2z8rC9DOdF10XoKwGhCZRlaHf0k8sJx/2KEK1sh75d2OiVyzeVFAnPC
rfPRMlTEuQgY+RJPO9bGNh4t3bYGUCAPcAXtQ601CVfUFgsas+JNJDzMOOtczizHMqgfvVSpx2KU
NSFSb9+FaGw3pBPVXfowwkxOLFRu/xchYTvAh027t8/FI0dDI9FOa7NUckS2Y0NYQgcTzOZJfp+Z
us6q611tE3CHrWMo0+maBsuxedAQkIZGclkIEs1ZC2RtcgCdsa4vVXz7uhkOGLec/KeOFF1jbSx4
IuRiLrqXpER3UuBrXZVLpLOksInChBirmS8wbQF2Xg2hLnQufsnfjsWZDnArpLzOe3coZ7KIdcHY
5srSvTooUWEw11uTfhtauc6eRGv1dl8CMjfaGd+2HRMJZTbF6NLzFE0KrfcrHHsn9G1hYFR/ojbu
fggyQQzMcY5/xhgOEyT7w53poW3Nh+zxbSckZ1ncDKkjz/9+cLFhCEoWyPadR13g0Q6F9uDQxJ3A
MW9roV77z6FtmhBD+PWheeBTmQRFJH66bllIXShkQsk0fo3QEslFhnNytGn+ooQbl6xEySJdxCg/
Ghs8dewS+kjAsGDfZR6Gt80WdMzzKV1kTSEKuZFgOL35Q4xAExkIs0gLZj/pLA7NxSr8STpbmyU2
CquiaGi7g2leJYkkc8L6f1xbj1T4zcz2iDPD6C9Onwi2HGgtegCN7ziqe5Vk6jzY0GTzTiqZ137c
v8GiPq3RgaRA4AE6jmfJ+px9nk78HtYDi5xa/E/V2LglTzhepT+GkJkK6hOrcxUoWOel8AW7lQkA
HX6P4F94qe4i2FqnjxbNz763Ei+wwXBhi+x6qfIGzcQoG3caPUyEhZvdo+CXAbvqqi2V+qeeFh6o
rIeyozI6j3/MQnD8SqSEfZ+g4kYfj0JnjE60Hk+xodKWrprKti6zIBe+bWPBzF4ZEqck2DgGkFSR
GMbiM9kYE22W7nIX+kLbTyB/uAMhS3M9IDU7AUkFjX+es9BU4kyr7BIQ5/IC6CDR7Qk/orxAeInm
XdXelQun4UreR3UF9Ft9R2Ex1xiXbPoT+2vVQPPguuH0NIcSqPeYPjK2MK7deXHaUE1T2cXicTLW
1D1/DdqSIbjrcT7u11i2fkt6L4wzOxJoJq/bYHqkvGeduCQA/UntT8RPtB4ETV29UZ71Jd/OpGqJ
gMQceFpVln8IilnmY3Fqh2kk8A4CSUE0cA/TsFvQ68HCdj3HJwYi9AXlPLGk7R+GFMcUOUWxYEbM
ZkL8yMPsA+KU2FAAsy1z8TuPFEdp64EyAAoGH6ieyEt0V/cz1ElppduNJVa2xsC5nhpQENMe9USd
SgWAJMjt+ZqLZuMXdwb7Ag2uyMI8mCD9euQvyOXK0467yFdYoxAb/LLgaG6JVC06cTcaK+mpySaw
LJ8VP5ak3W5h7DninhbNmOLCJ4+dpFqz5n6yKqMHYMrpgzDBYoPJQe3fwi8Jv4LTHCUMrvYahnhd
7b+YO3DDLzIq3RHEOoZN5eig4lRocbfuVhTdGJ6G26Ow+RDEUAZT4yU4/RgA52iaTMhK6eDlrpOG
X3ZlizFzTnDc8I5kT1WcDTbt7KOQmNYrIXWZ9MFfGUhJCpXl3wt4/qc9t6FD+DZRNRXQjTiGBve/
DcKfXGjUg+zUvg4EPOamidkBGXmPna3JzYcGlsaUmO+ySkwX9MxR6d9yFqUPSfoTfyJZZp3NOl5p
TCz1/68D3P4IwTGUk8Mt1Vs7y8BbU/vkN54rE9SC7DT9ed0KPcsCf3LTJFY1jIuQE447UG5qOtre
KKnoF6Tc1WTiPbRcnZD1IMl96k8JfFhyqoycE12egtbA2mvJTlkTVJdoD1zT8nqwlWhWwyVAW5U8
T1dcQJGWgQO7e56TKjwYz9fkuDqJjmWYJ0YID2urQRJ+RxfP904CrMXcje2kX8Vk1uaopXXttE5Y
FFBG/+l6U9QeA6ocqa2ULNK96hw1oOtRtPHbEPf2b3pO9yBZ23kSaEXVolvufptJjcShmpi+TOe8
1d+v0NJlrIfNLwv57NI0OqGrzsS9xpEwVkX9Gn/FTIsslSwixw7TPutW5CKbWAKd/aiI8WxF5LzY
IBYfCGDZ/15QxRXHMY0nckS+mdYTlFG5k/fm73B/DMPQ7UAt7bqLk5qLrIXqTSZ7eWBvORhGmAvX
T2o8zJ5eCgkxAtdl0aAkGYI8WZyZjzR1x7Y0dBHpWHaKubw1nx2Yh2Toyo3H87L3BRVuQEHTKFCF
LJOjSaHDSax4muq/r0gPW20vSsWu3y+VVGSl+YplIlYG93h004NtSqJqF1srI+GBUjJ9dgYeVuav
VjGED1WnuRoRrZ/zYCIpRcn0Ti6UX+b93Ngy4NFNOJfpYaUSCeMwoTKVOIl0CSHcPhMVlaXb8H/T
LKf1bj1nIhq78HG7nSnL/wFASeODKDit64TNtWMHiLhNlge1bN1JerdPssJB3AZ15/7smzkXDhG8
P+ggCwtGSesXbQyBm/255NDz+ur/AkojFLHrthEoZhy4Oe3phdzxBS+ItFCrodoc1txKTmC8Oyy6
LPPe3psB48pEPoiiAWSS/QCCi1idIH2WE/bwUEus+Yn3xpdQJoEE9aPEsjubm5NuSx7eqRLOVMIk
73+2uHNxuiXlC2UXeEIfJ1zpHGDd8EqeXouyzwtjhJ4d3uJzQfZY4lBu0zBHQaYY7HRJIcHqO1/7
VCOw7ywLXcxzAEV2R/LzYN6IVnu586CI1ZJguNBLV+q0NiCZhzPO/f7mSWjsx/Xp/nufke1VoO4U
EYEBgBw0BwGwDQYOTKOVPu+O4r2482CFGmcmrp6rZzdnrAV+eN+UKs6B20Qk8gA1PgzbE3E39pyo
63q5zzLn9ehtwMJbFxKyw44BZIx/rwsvt/0E/nX1J6kK+HSt55Lr14plsEHX7+8Nie2se2jycs02
Qaol9hTM4FuuvMeHHtNSX7QzEcpMX6wIQZ2mVVV2f1q3bSllubWIznAmaYkO1D7ESeHdbm9ozUBg
ABlZfJN42y7j1W2j40yK8aNg7x6/RLnU3bwcW9M9k1rKePLJ+2SUvzBcQXM1MuD1KM/oAXuL/IMf
zr6C9jiO+s3ki+tE25KaHvYak92iDiKaEiTWfiSLXZ6pjaa1WMh4cYA64Gsfw6+LvOWGoucoy508
/lOswHTcPYbXikWXjetrhaGhlsAQ0spykaRA94Iunj1LiX4njS6q7ng2G3ee2NxbBVjsPWCa0O2/
PXO6TcbJ9nuD+mEiAUbFMDHDmUJgjM0qm0G5QT2qXCsL1GA2LEVndDg5C5zwXrNsjYUtvRbPMNxb
4Zssw2TTHfwiLNpRKqYTE1U1MgFn2vYHl5iAMuw3SJ8PltFGYunLEW7g1CoNXpi/FZqB6xADOLcv
3FK7jsrNIOInRkrXhVScdk6i/G9p/bik6fQ5SYGIR1g+2F04en3lzq/37yDxs8S5vtDNtVxNzRHw
GNbYrXheSHKQNZ1nln6q75FE2QEl8J9H+sFxrIjtBfgeQ0uw9RavrCPPYmtN5A0ir0bCMAmzHu0x
4H9HRLf9FULgSuxvPxn/koQNzx6iRERMKOYQhsC1HFgLwSlQSRMor7Wem76tDymnZbPuXYUl/dZe
hd8yoFjKvI0MnosgCx/hUhjI/5VYxKl7AHJwFY8oT0tl4OOgnzXms7qIaUuDXw5+38h+hI6yQZi5
D/rYr1LJytyhxpABMMzHsl1g+uVoane+VqiYp2TjQg+bNf5atXLeSozj02W4vgeOEFEtsFcpuo3c
Xlkzxz0+6gOJAFJKA5F6kzrdko2NZFGvUqiPdJPCVNZ4a4VfEXypzos7QANjCpRDyOxJhBwEqI9Q
n2laiUQWOxeHh2KwTdaKEcuHx+PB1anGrtT3RZUoSCYsWs89EM0T10lYLynZLphvFLnw/lyH26IZ
3fzQbw/7LmfnbrQWGspM0FL9+erTBlzrUIM0RIcIujqP39/DoPLY3e0TBYO8eLK2rHOHeoXyIVd0
gZ0UcC8xXElvyoci+bf8UvrZAYFAABAc1RbsC13fVLehdBOzP8eQ1V1kGTrDGFOBR/KtSjWFcmw0
fHZB3RXz2YmeRcURAjFrZMq6ZeMmU2rMoKVLRrT5GWrRrzvE+vbyMifytzllHsOhbiHscLgAqdfc
RBPi3ZabwuaTSWcDt3ZtIWll0yk7zJwN3cVzsuc1JuFhknZ4Huft/yG94jvjRGeaLCXkeRFUxD/P
msgeTo8kBt1PgFVJ6WU/HhrM4Jw7xaKpHFPoRvRQSBneF7oMcb/10l1e1xSstuScHDviCbIbYM3y
V0hwyebPwywvo6VZevpdn+fj7Y/CEUWVyRaHWnidUqUkLbxyuj/S07kHOJrLPDuMu2pG9ODSR+Be
LJYtQlWBRxsPXkWzdET84xfnFvEfVwCxIbhpJyu7w5DXjLtBe+0PaOm8VGPxpA8KISQKXKJUbXz2
uhON5nirMARRxObdH3bRmxKES3di3HOlmWILGCy0M/xFG2VcVwbLFInxgGK1bgUCROdOTZBw72r2
idJrI/Zg779NXo+C21igYntOhlSuKqx+3gf7p839FhT2O5EMhimtoSOFqh6oC7tj60YrLwXEcg2j
CW1FEC9gVqMZXxQ+8+mY7Gs6m+rf+xP0qW7L48D8QKH8h87D3kld49orr4gHJujYn/yONQzxkpbU
BWYf8n0r2H1cbp2TI8c4YyIFGkT8FpAiDJrshMVI0nQrUuI0CBiIxp+pC0VdnFwYyYfJg14YsIHg
SpPploFTbn/h/F+ArpF641BhmYdHDAsW3c/GDejQ65hXg1x7Blr9S0Q/EXzyFXzN/sSbLxHUgic2
5c1bH113X9tLvTsL3yKJ4ewYQfj1xuc+KrqAEXlorNL5A9dfkEXOi/W6A7OvLbelCsPWmllwC6ov
C2mUW2dTu+51N5S0YoubgyjlNs+qA3anH4z0CxnJacESJebWXmzXqbldMvzLoKHsKlWbztPrMvyd
jURf3y72oa0LSH2ALB3XvY1Dg70zgkHchF/4mjuVOHx3Hdgf5Rqsa25NLHWeIw7Jy7/AOKDggfZB
bJd0B2TJb9+Uqxhd4eLyZVdOqave7xlsd6du9xZU4e8bLZPq6KXK1qt77K5z495ApxBTcZCDOowb
sbPTIvofEKi1knTz2Rt7g1t6pl/HVPc053cQjQUF+kA4VzNbLjcE5YPyCW4fVot3SQTB6pYIr/tZ
p4reVhuiU6wGgfblI8tStwnSr3oxw6DxYDrXKdPC6aOsz795yORD6hDGpc4yngMKIqbhbdqGu/jL
jUJlqNXEHQEnH8GY2rk6jEuk+ZzAu/2RKZvDr2sre1ynA9bNnMU+Aj20Fbqt1DrIciUR/AtGL2BR
hz3TTWMPOcqYpORvBAxbbJmgouMl9SWQEkuskaMKe98DA9AWseif3YJymAoWmZFbs9EH9lLK8mmE
rscx6xptEWdUgjuZrQ6K9E6gEuTOwNowt9Szwc09anaxOrKbAJqA4Q2dCRDkbnhuubWww1ISFt9M
CrThgVVXdOPWEub0rzVyS+uQXSCT3mlPdRaIA5PvsRk+7UD5o+mfm/ssv2UdvdEteYd0gnhwqYvG
IxjaKaJp/47dpPObogVe4I/rSCRdoFPHgsbUEUbkTvlLUN9LydWFft7uZQTlIakmgBEVPX8n6Gyn
9utl285Wa1Fvky8BlqgspEkYOh3qVsWGMqd6NKB8rnOlI33Wq4EyqHdd/SeRtBW/g+kSZeGAkrNu
Xy+1SdZ1PFIUaOVgF213FwA3PB/vtbXlJCeuO7HHHqbASIoPfgPmC3D5ahhE9/fhfI3mbAFeBzvD
HlHX0BnXInjprCdYuiXR3CWdd33dr9JN0LNP02YqD33+XfMYSW21E0h9X6AIsY/60mMlqvzUXkzY
YBQbT9FObVvE5H6Kkmem0l1jvMMTX/FndFit6KKv3ASKKPKCr6HWwyYCt1qFI+VYeTSOERf0jyS2
xDieu0MbyUyyMW4anqZC6DR6eT1UpqnDS1lvu8ZhLZjQP6DwF5V0ZQ8MVsp0cGaLnU1qhTDaXGKk
JJeBdJlAULuoSd1tPMa154JEEZLh+w4Irq9RL1rlHNrSRkCa0yrZzUMpKsPp6xqsLX4rTvNg3Y8i
NNmPINTeJKBRu6it8z8GML7YXo+k+4fJKwLoYjpBiWpdoDTF/MRhXVBZEmfIELHQN7Yb60zcKE4n
nv3aj/JT01F28GWNI2Vv8kmO2qinQI7ZRCZYnojgGj8W8NHCbDn3YrXA5j1OVmwmVkZkLTaLY7/x
aWOrkKcKcRHJE1awr1RlKCy9QyKm8ZdiOUf04FPShQG7XV2fw2YABDYX0t5zuDZeGBXgtGC1X3lC
sLZ0GFOh3kKn90SSjnOKwG3jXvYwJWDfDCIvqyrMy2GTebM/m6rTtvpcbSUKvGaCCXeP/6ah5JW2
Oi1gnk9m1NS3tdlhY+T+XV4wvkZKwXaZ6UYSh8MwgIYeqEUPI94/nf3LIak/cnKYA28HXPCum0tU
ABgM9R3K1nNQDp9Wrda01ZUrN/nZ4Tl0KHULtoM6g6ahlvyTSgkO57I8NbqSaAm+TmKhWhxDkMY7
KoaJ3SspuP+Lc8VUOiNf0NN5Y0HPKCTpwGDh5yCxkOy0MrOQgrAXeNr+lBfunWEbwl8gma2GkIiN
7fP3w5Z6IcaaKvHmpcYk+LmTpg7Sh1Gg6lQbwDPGoBUkBZV8c2BZXBr4FulIBIzM4/qYqbKcEh1f
t8iqSJRaQ6VPZ8OVQRy0JQfdufPz4A4i3nkJ45CpM96eAODvEvNI1Ebr8gCrMoZ+HL9TQh/5JTsp
dwOwES1aaSu5VNJ+41ROaZ4/0MNVXaoyhDhBUjqZSWrOc56vay50A3pxV5hjTvMQ7MtoWGrgY684
WWPaZMjY09GkL4dpbjt2qEFZTFhVzyJ/dAto5r7XI27lFnilV8JF9QNj2BZI+Mkz6BaSvr2eFQN9
FpIrBkDGvbkFlEjk3uAJPM00JTi6tiJvvtXx9SSFDLfo3fw7fxom8SNSvfGtKxw16VxIMOwomNme
IvA5G/y8dRH4kO0B+2IuQ6ro7zUnY5JNAAolnNftpS03nPf+qkMA2mC90HEscXzpLgt/kc75kpxE
doqkfAuEkb2Kg5fBLRPHBO1N3AtMDy2ca5ygPyzTFbE9hZhrdjjwmrwR/FrhvuCWY2J15oI5xUzs
AgHLwqE6PL47RPeYBjxpxMkmJV+4+nVHA4k1Wb8F1WCxbDM3Kc7vBal3ytHIKd7oP6pxk8QIIodP
nK0787tfcuOy3LNeKoHqKadDneIrSUB5qEBSPgJSEyrRPGfHJOzdj6q/M9KBzxVTkc0xczqu4H0U
7JzwTEecW7qfRBH/31Xb1/ckr+wx4aA+LLF3KIf+evWGM1KZYcKBNJaOog8H34FT3ACZIV9jpJI+
MBGSz9UeS00fQdJGbRzyMxpgskK8HboKd7O1HjdOKzwPj3y79wmQAqwC4rlnOAhfeTb/ASY8S/se
viQVoyLtpQQ3TeAlCX0aboiI7myvrxyG3Xj/fsR+XpmqzmMSxxFaJiGZy+CWN57RRF/EgA0Y4qCF
bRk6WxOeG1uJdUNV2u8gjiz/L2iMKJT4DqcfC+eHb8XWG9S9ABRuPLTlnf/ffhX9KU0Z84m0lROj
nnWZaeNYQV3ku7+aRFgxe3oLuVjMefXs0YMWs7IJQJ+qtxS6v7sTe32/5X9HhZlAFQhrGV7PHgCt
nVp5DFAPzAG/e1tHk+35ZeKyQTkb7No2WRR+s5Po+n45jqvXWBDEwPFDUKpBWRWKIZPCHDtM29Q/
LqLtUtItRBB/EbfnHhRT54Pk7TRf1pgZo+b1ntnzDyeUw2BU4SgNym7h4RK+nfe8RXR+6e/aWp6d
IrBn3cGoSVXX6Yv8qQkvTMs1lD2J3EsX5XCCzMlfCDSZ1LzsW0hu9s6OHrhC8FJ5Z1e4E89ruV9H
B4MmMw9yRpYmjP2/dATakZNqrn7Eg0EjTzlO1kZegW7LigU7kqaNNDOEOS+wtns59RdyKd0+8RrJ
Q8YPKecAFu2KDT4TiXUf4S0wMosJdSQxHFwIe17FMstxirIZ40JPJV9+Ca+dxS37CoukSpZLWdf4
Ebt1LsDe4ZidQJ6s5CD/+u7GkDD5Pgv5lQoc++XEGpBfmoZd3+OspLV9t+gydKJNEtrbWCXkBLws
Q5LlPMVH+SlPyLe1bwXS1cavdH+eU7sl0lioXZlbdR7UbXm4AwNX9+NCbN3etgujNljQyZoScOs8
HmSmrKZLYnxZgma4yb3BO49tsaKCqclsTjp5FuqOj4rDonQJUD/Xb90Dgf2eTa1RNvibGxhRC03x
oh6YLs7+oOqZF0odzZtS/qiyxO9QLlZdOHemesX1HjNYz+LOZ0b55H3ZZYjmJ6We3M2b/L1Hj+PC
6qtLBH5MRWVER/pj8/29ubEBE0e2gNJNMBQo+rGa4otJMdG0SmyBfov40WvZO02vKTPSxSIGD0pv
JZwgMO7bMSQohZE4TBABKvTyHVAmjNg0m7QEWP5TUlMuPNevTdmoFkpeRDl8NrrZmXXkde+k+jj8
Hbc65M0ZcVOpUiTG9TUeMs3qGt9VnRg5EiGnO9/FXfPs4+z9BbjHkxVA+1zPH6iE1uSDBxCHhGcj
SYx9OOiqilr7gx9ROeo6R7Z6Vgbk73AZAnF9Ouz3O7yhQ8zCcEoSh1DHBxrm/yRdxpXq+1L1Lulj
9RwOvLfNslpfni2BufpLy/Iy7YuOX++fRhPUf0aE14wTaXdsXHsJZ6mW6xMfWV1YCHbvlmQI8fA3
Qla4KKVJcIyS0bxpRrCzNDzR/MNHeQPL24vhReMiiXVLE0dM8TwqBKdKeSOo1liqAY4r98m5Rrh5
fL7fDiPdvb1PNNbDVeYX2mljEJwxFbwyFasENETkV6sBt+Y/2oDuKuy2Z2VGTkB/BnmBz1YsmbjY
Oh6It72Dv+vL2Z5yNfqSHABfpt/1gx3ONswKBMT/M5MbmF8qmslfedVL5lLbqs6+uOtbu8nY+O4m
P35ufkUxm0yKrkImGWs2gnBUgZwMYcDrUFi+QDAbVR31Z2sMngwfUY4yZf68dT/hu3zSeSgR66tj
lhFIENlPFxF6NdrtI3htCBIM/HMumFzifQhn5cU70fZXE+TFANcpgPdwNgR/npkugPiEIfSW6QMw
qr1jAygxjfU5MvTXt5IF2wkWwp+tDBvCAulPBjQFw0lBgTQcMY+KCjAhaGWE8HFFFXJGuqD7N3m4
IahCFOqHhfSn2jQa+n1sbTOwwc3e7LHKdn0rPXFe2z9LHchZUlRPM3iMSwLDYRQASAYYk7dJc15r
tpiJ2yzhq+unj6tGPT5BuVdrmy//5CGY/KaqRv/hsmeACvGFAMmxXD7ZwbNATu2VtMy8nidBwoD2
QzGW1iseMOfG03janOuiYvtRzkiYxiWjqd9Apose7n52sijzLwblYmNpJBRB/yAys4oH5mi6OrGi
YBt3DUBbDjmVzwOblHUcUuTRWZ2KKEBLue+ywGJJOPii6drIGShrUuMPrYBVUiu6omJ3ufGFJhYq
4c8d/RQtzpve896i2ADs+/V6PWhtZsRGM4428dW2lODp9KfVG9FrfavQ9bvaSLAiFP7zb602WIjp
PtkefCHKT4FYYdtp2q6ImDZNgZu95+tspVkzYQaISpH/dzoSTZ2zZW5JSxtEYeyPvcj6Jre9sqsf
qVpydrb1fjRM4B78mdlf8nzj0paVeVd6nfe88BL/Gp0bf3n8k0oIGY9SrRI2DT4k4nCNWFiO020V
8BcE0lls8UECzNtTSwZ/yhIbFqvfj4rE5SirsoQpHMNd/hPRlmJfnz8qnclTG00lt2bkBkVL6F/k
xMqvbruZNw5bseSV5gQY/oP6QzqF7v0wsLALRooTpN2vKoc52Ib9pFZm0/lvK+vqPzgVLYbMMhHv
1dobeAA1VzyHnIppy5BhG8+0uVHD8Rhe7jCpYMFmq5i4wTv9D6hMNjHK9dib1X575E6RVRhe6P1S
6S7rIrHnRgUKkH9ckuiF4OGCUYLqbK4UtJ7jyNu89ygl+rfkw4tMf3+PbyjWMq535kaokcf14sz7
hI5Wx+ygWGDeinEt90BpO/Zu6eSaR60x4FSF9iZKzY1VFCdQkZaJo8gmo9AFQe/9Eh9qr02EKRGA
AMuvsL6J+83OAmz0KcFY7KJgCd8bFX0SyZ1L000s0+YOtNylLCSsAJdciZ+OyZ1JQnRdHAWu4Xg9
srwj+oqfLIE6Vn+9eiB/R3aLjRM7+Mfz3RuvHc/UXE7HdcH6rTJC6yd4KGzjqiWZQK0kS4TyMwNF
Jy+qDwQBYVnFIOr4Uj7eZ7KaRXIIqE3RgbAUX6QuqZpmUX2IszVOZaOCSEfyQwuA4vroIFH9hfrl
WwZvdGceREg3cHyyvalGp/9CLYgUNsuuK8TIWEsBLMNxiLo5gdLhZ9eyhIUmLJ4509qbg10raYTG
k6s8J4RJkTqEgt5xBIhisiTURKvV+YG48KIXf7X+BmYWNbdPRtihay+tNhE43QdGMBbAIfOw0dao
Q1/5Rz8y6LW9FE7oPfTNXvBKJ4OA+3y1Cfa7JOTPsqzzs3eA9aNh/dN2xruLZEpUXe7ppzPKvyq2
1rvLgAi//6foQc4JSMqUaG/xu2m1KjvdT3bdkmLL/xpU0s5Jw2mycMCn9FhQ3RV2KSCiC4ZhpsN2
KqJmlujfMZwm2FuOzbh+0MS9+SUkqfBqUROhUYjHZiLJKO7Pw28kaZOrUdf9vOYnjPUZeNq2gKV5
KBfBsvs+zdaVEKZ9w7HZcixw+3NGil/UAaOA7aaCzfh6CJjoxW0kFQfI5F0Mwn1uA/NUIyi1Ac+G
8WHsj8zEhz/x/N1Q66cr0RP+Pm8PixY28eNznZRfcsiH0y6MgtHRAep8iZo0a1ON7pmdPpmomfQQ
Toyn07MHsAzRGcA6yKIXUorAOwm8pEq8SehiHx+4/qIdlPkQevEJL40hbg775qDtQkdwp43UbC3S
3JuBulDpJJ+TPLuHiK0JuGHTOq9o+MdcIzWLlgYG3dwkOY6c2UupTGTrWDwLepue7yLEdYo+/I6H
f9WL/Lkp/r9C/UBQ3GTYhy/7UzlogslmOHK5+aHzj9qnU4bklxzheRLCHEgx2RtFZ4zmWxswRCaA
zIiKRi4mVIfArThSJSK603Qj+s1w+Dmk4xBsxGHTZOblQCIul2SAnB8iqVaqg1vQeQ5gUBjwlsrg
5EZky/8fM3vLJWYFHN+a0tLzmTAtTQzDLm0iUcmOmiGHVMbIYgD6L1xMLb6+I/Vgr9xrggudBrl0
B5K0X4oak90iREGggG5HgcdUI63g54Vrb+IwBuOEiUiaHH7DefdMJ5G0Jgo0uxwMxKSdhvcNmeCx
Cb3iEd60W6qfKxMD4BrIyMj5Cz4HcyNlEz7pebERgj3b1H8iH7oUU27j5GYkZCedKh/QbCkmGrrJ
EFnrfCeN6/85pyyW0VfNPKNnpZ2e4zV2gdPj5+8BWwlYR5msrHrzTn6eh5CyhIYxD1cftnPAYkAg
7MJQ7LeP2iS31NQqo5YGc4qitp3UfqysSgAta9jYs0vyVgTEmOx0WjKc9GD5rkXlSqyALvaDUGrS
8j4vVgEDKrfFgS8tDJEDCUjta7RhaTBDmhp/w70ntDi9JhZaEH7FUsbe3KwS1IC8KtN2dCMgH7Ph
PaU2c8+dxRNSI1ZDT47Wjx5k4tzJb4pMJIcwhCL/b3vk3tWWCXZgugcj18AvxLBYmUu1b59hrkDr
ALVqjIRBpB93soKUEkWKrjaVts4n2zkWXZudwF3c7fm3BVcm61QVjHA+MXeFP9O+Rcwjtx6S1skC
YTI/75HtHyCYODZDQkKvaSgFBLANcizcONLMBUccpoS8wKEs7KpIj4j3UurcINk76Yr0Z6Cxunhu
W/6ZHtd/AGrz1DNajsIA4otIXqiSBXo6cHF4u1R1BetVL5dfe93jxigAXqFRUHM717simKPFy5w/
GmCBYLfFyNpWhODWW5M+CC6Ow64vc6K+55j+sUXmLxwEoXqUBwARhVznLA8Ro0/8VbkvxMkoTNc2
2HUVo1ffPAANzJonXCUFGpwSJ8S+THm2/1WYU9En/snd0yhPTtg8akNZUu73TOGWP9Ey0gfZuAJW
LOgHesidk85uIrGWV5MzttZ5ifCtme4lGZYMwe4ypHeXz/YKJvOQsHa14pTxRQYqd5sPGRawatYu
tnro0sMD6BFRJB37ucgzJibT4Km4pfDaHT2GE2m3UvSs+5DMILC6wI3ZLtGEEw7r8XwUMm1BOZsh
W2BVU0Po1Gy7zqr+a2AwYz85u1umx+6JwmFS7PCRUU/qGBN+G9AgkZBtS2E1cqUokvAp/LDGXHfO
2ZNspxYxZqLiZkyY7vtOy2sbLvC2+7sAXSZrVgjLzfR1hlVX2XL/CoV3Bvea19tqKEAFJijc1XBC
21r1ZV8vTCly77o14YzgmReMpT1LIDfBC/19mh4YZFY2VOCxI+EOkGnzBHDe+rD4OJcQ7RL8EYJd
+23e07opzCwuVMCE59wRP/OYjOM5oUS3xg2G2NPGyropWZ03wDusUXIDONnqO4aH8L6YIVNGEjFX
2md+FkUkR8PlTKXxetTDxXxLqDPQOHc2rP+LpkcdS4JR8pxi5EAM9r1QS+RPso9nnOeafgovA46+
vW+ijBnuUJBGAkSJMyOw5/E91SSiiNhWAgyFEodj3n39jc+aFK0RLSrcTdPp9BLs7BZiDK2VrDS0
bc4flXMt/4SKoKFvrpfxI4iM8e82pN3lLtCfDJc8geh26TXQYGFtwhW5/4OeEKqdr8MQ0YO7JSPf
C+4zzL8hvLSfJ81oF8wmWoH4er+yy9OTSzPBm6K6aJfy2RMq/qwlznrnD86edgIaZdtaDT9D86d2
za1JlQhAkbPsQh4ThzfwGSD5SiC1PS5p9A2CSxC6YQq4PXDR4VejqIKdsl29my5Q0eKX8gqpi+++
DVsVmNIrkfq1uEHHRkW8e5Ys3vQPNDJ3UbAimCY/83+0NDJR10dh/FDeog1aTfVkL4U4s/+9CoT8
dD2KmNx6xSeOOi1T8/eW93wwixrrSmWWJ9Ksv+M6Bi+BTcJcX6xJ2AdUZWOMoLpywGZCFJltpKtp
ZivL9p2ErXnBESn0ZiwfxGRm3m1i+xkxIQzehA+aykFKlqSnRh4Ta840JtSNFo6rNuhWamzdIeZm
8D+lETdzYmGwIaGD1NNPb/ExuHZuRAtSH/IUZDjxk9+zJmgEeQrQkmUFClAxkV+lH3vPHJGCg7hL
HrlBH6cWHAM9Qht40vviaYKT6ywVQcMsDVKvUcoEICOiNmMON5bmdvrfHBjDK2sYQrAb4G0Sscbd
t0tE+rufA1gv9UoPxQyCj36MXKrNFNAKJyqpFelQB1s528YZ7lxsgMDvDyF6VuQXk/C39LrjeAzU
V9OP/nHx26OXAy3JNji7aCWcbe9q90DJ5TjAPEPqN9nO6efKkJWnR9L/yyAMUGC9v0jSKCac2s7l
h/RtFb4qa0rnxL732WiHWGJnRZqXS2//pf/Cih/PkYsmcQhlDkwyJYeXq64D5P3vYN7RnoYxWUH2
5GhbwblAqfOGDAFt88xi8gQFtx34mqaAYSmAazP53i1jEEMSDNU0JsljOdpXCAAnPBB6vN9D6D2k
viD+02x5CtHyGcLkc7Bw9DLUimScUGcbKxlB5CV8Zfz71COtTGMhL4BJ2Iol+dX89qONQs80lAlB
H8P2Qyo4YfOgA6RQAGnmyNjfgSOy44BB50UIa5KGzWYMEpfq3LxGCMkzfZ9M2NIXpoKXc3+JTYvA
DIZPZ34oGZagH0DM+87RDbmXSbWnDprTXV3qfWe4yMJlVPOrso6V+Q9BISDElkdU5RfSiBnOOFcT
kVrD3i4Ztx5WK4BempkyU91MKJbvSxvFdVF4QWeEMqZDLa3GIQMp1NdeJeCV/SwynTPJU6P4CchF
ztKdKeVhKYIC6rr38dEPS1QrJ2CaYPmBCmkarYBnIdu58GvmpYaJsfwDWLRta3v+q+v2VvkgjYf6
fCvZEToWT/D/HqDMstspPL9NvxjoI1vdZtYYG79Izn0BYYVNv0+060zaflUCS/XDEa6e+Lh5Vn4c
oOjVGyZsrK4UqYGbG+WKUYrJ7fwdjUtEB3+36mOD0p3WZ5NSHLsgzAmg3W9vZUi0K9O+4q/mDR2G
jkxo4EWmHvu4xNoI5qGizR6Af4r3MfOYY2PVHB1x15mi/ItfZVLUhRt1hJxn2Kjz274/mz+7uv87
hFlt7pfCmf9AgaCbtSybjBQ40JUgeD5T2ipx0ky5RuYHYXlsSCKWydJ2muxdmouW6nmMIUpvkve1
46EgoeviYY9MhqJ/vMDQY6pCxKs7Emd5QfrKE1+6tGPqzAoUMB7UZUiV+n5sS0I/2dfUOORIK4eV
27NcJeMU437DPp8v/P0Og9fjIlPkgTm+7jzYgp1RCaGtnd7NBQBbX1G8wvpK730RYELjajoEojrH
4tckcOMFstk7wT1/JzHnoJRaFvMPsm8JeKUd/TIT1XkcoUCy2TLKY1JpkOMjnSTTmg9myc658V15
m3q00paZ3QcvEkopi1q0hbiOin2td7KpFGt0kcPfRfhtzlepsue9gJJcOP3RTEsOmZD5JtBnDCoB
yGpcSKA5uIJc+S3Uuo1x5fAL3BCe2g4jAGszfoAkSGyerqOd/pH1DVR4l9NSJGUWmlEIB0teKxAR
6vhjizTAIO7g4T9wI+FhBad5ik4cwAKpj66NQzwaQ5E4Q7acfvZA714haQ0OKD20EFxlSz9K7hNV
H8NuljU0zCpA7jAwys6lKwzbVWrAGA4xd4g1P/1hHTe8qMeuLrvaCJ/5q0A55yar/zqn7I0Pw6SC
2CyLBiYqpgZpIc+KFR3c6I2ZxWdZdwZWZTEuwy9xKJDL7/cspPQuc21Ju2atUOKUlXg1990eGoqy
ZO3AnpR/pAPJrfxf8C2oO6ylRgiGamQwQFC53MSHOfVwlBvxCNlU6LA+scqeH/hqskOt0RbAdXaL
TwgNP3Vf7yf286Cij/8X2klGuxLl3XqZNg2hmtrDSNBit94HhQHWPf2HHB3Wi9i7ws2WGGd8MRRC
GerDHTZ9n6ErJ4jO4AB63wt3ENhEfoZzggZhtURtte7ZaGGGwK99iy+FUz2bJfhuaSF4bIUxDfWj
2KbYpAecEV/ek1M8ArIeeJpOWWzFVfa1vLNespQq0O1zJJ35W1qy2KE8IfRcgMaXUEX5Sr2T7ku1
6KKcH9+fMNwsbPoXgYG656YrGLtyW1+uUmkr/XDIOr4/W6RzmH82N2PAa7ktWga4BCd1AnwmEdi1
dzIBIDgdulnNM7QZOeL16fh2xqLX0cSRRtBOBNMX5rMQDhSu1IgLQ4oNny7Xw2MTBnoR/WH2z35I
vVS7DRK1YRBTAVtNwxMeZWXfjuJCyjCdCCJS1pJqM3bBDM8yywnI8/2P2G6bBPEdWhQep1E0SnGT
0Z3/k1NtSiVxFGSe80hfw+Y5ZHIMtZutLrbEKwHtLqPzbxIyKuysrv0tqrm7l7VEDYjTKUVMzMIQ
9VFVuN4zeUxm5wFYXglMX4T5aq+eT2PJkHSG15TIw3PF35TYoDGf2ME363BmI6Ml6q2Spu+WPezH
NHm28113wOn7SwFSrzj4VQWGYy+sLOb1hBDkzmDa49Wt9HTm19GrqQC+ej5QIjgX+K/NtAvHqJs8
Q8LCHV0NfboaVy9BJ7BFbwwrfMbPnIOKuWAKljTnhq0X2dCwyGjkzxAlONk+bwC0io4OsiR87Ykv
uxgielGK4KeGFkxWayyYU8UGu3c6w0Le14cs9b9uH8ziXJyjRTLl67L7RsxsDaA97AYNU9k78Y11
YW76nCO4T5kQi/KSvZhDi+IqLz/S3pU2pBCohNakYqz21iAiHiNcPEbN6kyFTF6RcPHwbiqJkzBf
vAGPeFbPNgdcCKL0iTfdO5nQANwQsO2mqtS6YM3HJtWgYSDA+MwWYXb1x4cOxnTZ9+Kkso11Nmze
BY140nAAdsSvQbYrpscuqzczlBvxZoOy/vTDKywL7apcLZgqO+G4jncip0n/4i08zSppd2QAMepm
UpUNhYXmDrf6e5cMgHRStb/WAS+E7vli8w1fHethQOBGNLpKfuv06PcJzEr7xj6OuVBLDexXIlqU
axG2tlAwNdjdrgyI8J2Yo+sp/8EtZI2Nlt2DxSml4/JxvEgLSHwS2Q/R5XjEMUTRFfVwz6AUsGZ4
tDUEhTBofMUj0ipOfoP8XkPiDLpzjnxiBzoEh+EErz0MRRYxEOwqHriyPpVr621lyT0HFkU9G9LA
1TqhrDH9AjsAiSH2mrugCHw1wTcknNk5oR7dFIia7MfTjMUnP4FhLlhJ1sk7E/3v2WULF22QbfaQ
+CltDaWu/lz/NHe+aBTHfN0riijdAqYALAnbAEO5pWE0kHuKXS986Kc+nSE7judmNB+p8myOUwit
Y5XNaqYe2VCkCqNfRExIK9yq3HtGoyV1lvs+I701cqiLGEWl1GHc6ZEb4qgmifTdWQ06r7OLt6Xy
4jDae86brlh8CQNXh0FbxFoOlJajDROJe8VttR0cy3yp+FSTfYVXivP2c2DPyRCjb+2qD9SbxCi1
1gEJoygB7EGs+/N9dLEs89yx6kKVadgRxLTN2jzkG/GyhiAxXM1351p0n+FjeFEdpjyGtb797qt3
RUkTEJ01UM9ymFh0b0V8Ik6VhHDnaYnUQEIfYEm0B5OS0MpNS/g8BxPzr2bnxtxgIHze/xIl9ZyD
CxmyNdNaoeqV51feQaafB4uKRZdAl6KfXX+omJsC/heH+hukbLPGdUImW4C2aYYbZR6jmhySfXCv
w9vHvfOd2+CWvJRfqdIn+6HpOmIIfam0GR14aQtlzjT9yID1jrGF3+c0Qq2p3zG1q1BDXmMIjWvx
vd/k4NM7yLqqrgcGH9lBhK6KKsgx0D+Vax3+FXVs6sBTf5UTxrcsSx07sgqGfIdwe/a93ox/JsnH
rc9QZLCmpRZmk8xe8Ul1TStpsAWl1vN4JF6XqOoA81p+jZkMu9Nc4zLD3MrQRQTt9SkflBjFQaHR
2IZWMEhBFUmKrG/MxUP50HLtdDdZmPSanGrjqBCeVcPVY588+sM+Sm4Sb8ZJGAqpTS/kiw4wwGYY
SvIVOUB2ZwOoJmsCNKZpy4CD7NHUR5nWOKvwVdfWLxztMD9Beg3oYLJi5zEV/ioBCdbhs7QCXBr4
W8ItYYctWHIeWZC2uYlDqZRx5eFAMqw5fXuysChjm/SIaxyyJhIvH/f2MCrckbd/qo8r7eBDPmSm
H27Vobj0yZes4RCBr4CyUquKXMV438i/t6obwJrQBEp6/JrwN1bSsFvFvBmH9UG8TiMZEsp8zPdE
ge073dQOJTOP0sZ0yc1TSg3ltWRKhuYzV0GbsNWDYKJxXe3mSBysMk4ST9coHU763oSzkp30/Cdi
hdW85b38Zg0/qSTBDADISb9SdfXVonSqJqL/uhxdZ3lN6O0P5jfvCtQm3mJgm1W80mUe6W9LTlYk
EoEo/3O/st9RX1Hoz0fuV1J4mJEl60ouj6384efbo0ty8uEaRgU03kKfQfBZBG6Ixz74TODdfnBh
DjYOBXnuTJtmZFk2hNSH9UvAZgRM4GdFFySz4SXK1j/9IFxifTZ/WKXfbajHVuq3BCm4UzlU1f58
UY2+fu0bD+DSDSUb+Jg3P/6hkXTtzPUf7vbKj5iIsg98bfGeuz8PThztXWp3OdjDzSKErOKX24vM
elx8Qjh3Ao5gDSgXErPyYorj71N4WVAnBNDYU7YNMeRD8aJROb/fKch/YhzWqth/zZNwulfE3kEI
d+BZtEeSV0gQbmWssOPiKmjCR3BdnruB0EK3oR1vUyhUYYOfVnlZlNgjOdWekZVcnTocZl0PvX9W
G5+eoPb5RbNVdAR0P0LXBwNxZMWM+g5lQ8/ohMnSW3w6qVo7xSPTodBuTMONnlh3+mGj2bB8pCv8
nnrkuFN8u0aoVV1+SPWV7crCbZPwS9jDNkE4Qgrd6Npc6u9CBxgxpTl1O16h8Sji5bLuQ0HUZwA/
QaICjaRVZHk4+NIfGEpOnOFC6HZrUaaYO4GkZQSUKiAM+QnTWnzkHTG1m2EHMeZkXbE0xQL3XapI
9kIAEd9EQa+G12X3xCZ0n7qoZnwXSH8OwWLFvqLKF7OZYtDCj5mIas18nCaWuV5hNM9vC9ikvJ2m
7tn1nnz2+cXqJZ471hEIaIwf9d+o0xg2P7Fl93fZxuICDCnnVuN5twleCOyGSblVc719LmyPQGfo
RApGo5hN2cK45LzUAhbXLSZiaHfaNUaa+a5BskGbz8BOQIgHvsp4PD0kWkdhtal9UIM5X//V6AIk
VyV95AESwvSLvmxdwIf5KyoKBiQbi/XdG1RN91ySykhahAQQg3/VIdLSIQlBl5dRUcBcuVtDBs5h
NWCxy6eaZIc7rDU+KiXBsmqPbQfl2jkpko60qPxR321z9zeUkzl88TGlJKVnv5RkDHATm/rgA7AW
p7xZnJUA5EZ16PCZ1Yg5ueXSsIj3d7sh0U5BA/841gT5eY4aRtqeqYIA2Xc+VsXVvc9AKesfrD8C
/+vBnQrLSq908OI4Vxo81yHd4AoF5UAFYTtBVJU0IoMtXYqiB6QzLwmhk2yeJUXzieuDSHbYChfH
ov8p8FYMRUa3cycpYa7xA+NeSULEUFM6tG4bzY+ch5n+qP/FW1vWopdFJkUdMmVEPOg7jPIUArHp
8pgHZ5idk1+DP8jNz1XAoOQU5fXZsHrW6yO9Pzs1gb98kPE77BWLabiL90rGRyfkxSqp6PijCLJl
PZ9XWSWBjwAUwbvkn1iCtcUDcVvnWYSHw24zL3aL18ZyCzTZlWpGeFsayGiTRGjyqARKNX1Bw342
EPYe7zCjlvYdxTtML/Zy/q9UqO6khrvFJUb5O6kYLC0QZpnJsccbGf4KVp+CT3NHnZxfF3xcjZZy
QvfxFogM/wSE4/kGP77DV0PRI+giSvql4GGav/W+UlsBsFoWith9VNRxfAdFiEkzJtU7ykqAwsY/
rONcbGTL3L9hdoOMEQ1Ztn/4jZGLINntToSz738or3uWSTH2JlfrmBtsy0D5uWPwAMhKYmoHJbkI
ep5WoQ/YU10yir+9s9gUICIBX0uBR4rt3s6VBLDSmJ8seC0p7J4cNd2vK9zWDeVGxxpj/4l0+u8J
ERU+skz2ZtgK+Jatxnj9UbDFLNFHaStRjH4PKe6HN1GHbfeBliZror/yASNGSG2avruAsC/1lHZ5
L3doXjiulcKhEBvYQ8fXK0suRgoREIqgb0ALOIsj7WDOWGed2L6KXx8+ZEvfArgBk/wAIBLNf/y/
OZ0F98GYSPLpoL4TFlkc5It+iGLXZDP/TA8mXVWA55Ldu+HtWEZ0YMGkEbgPidlQqwlWP+wyMGDv
lmziG11Ns+40hW1yfHCbR2iInytZCYbD5wwCUwzQdKp/CCYJCWq0bvLnWqRX8fHwkAOzaXxsbcr5
66HqIFrRvu/2srwWHka90RneG2zKBuGg4Eo7xSCtbTsxzZja4zcbUH6XZ/rx+nVHcFkVz4qfXpF+
EFG5h8J6UWNX1Gp8OaRnqyTewFVMqup9noSzSXUd4Alzw5eEDv6ubtlKtGwrDfeumzVBc2b9gOBP
NeJgtSsayJlYa8/LJQd4h9TrxzIhKjqIdWWZ1PaDMxhiqBOmUXjA/IQ/MDivE63vm3W0jzPAQKO7
RUpbvG9JqyO4zJQMB2M8Hd50hHQ7T/Ugr8yfeO40MyELIYoclmZhCkOj3AHitahUrnBuWdiNc0Op
4sC+iM8JkmsefiitOVhv3OmxIfj8Na21F0JZ5ps86Lj9WCX8voMTYmpAjEUNkM752f4gysXhs85u
8A14kxUTpxtB/+n2dgqoz5QUny7kNEHecJ9KrA9jOIK8M12kDFyqzSXyt+5VkY1p0dqiOsvdRdjg
VXJfZUPO504tjLYRtKhSv81/5yRqy5MozO671nOCmbb+9vNZk6oDD5911WZZ105ZXgaPm9+FpRvf
2ou2DZPJM0xEfdfo646KWtD5PMTro0IBcZEFjYh8q8B2EN8YvKnw/WHO4tFm/CKQ50kOK0W3fPS5
n2zK9JbcezUT0foeMWm3oRi5buWeE+w6XwvQxmcdfD/lcJxk3tzNX7DOWivIsa2oMy7B22rgqUBq
nzCbbknioYepkYsZG3/19ikgB4k4oO2DBvKltxIOFzHv2watWEfEFNRDCCLJyNsJ55X6wB3wWUwT
iN5L2mfAK7a1GG3loCDz34/N7/EJ4GUyiHl5U4CYAZ7wAfhLP4kSWnU1EXSQq7Aw/BCmLcpLQ7Lj
NwDFxtd5Ei4kLuvwdjfVqncM6B+g29qmdTSj6SE3iQPJwKMXHdHipWIrEEVIg85WdKV7WG3kw9O0
m2Xztam65PUW0egLNfFkSWc989I+VArb2VpbowAYCDhi1t4plbF9nkAFxvzOJ3JfI7/7KbAeR5Cf
KfrdpvqCpkIYOl6JNERnIbJ+n8B7EGofW20FhIDjsBs5riCWhr+PSAkZJJhzB600CpZiSo9pCdze
IH7VmMyDWmtdWpJ4KMa3iE1myjFEMpXK1n7JvfcaR5qQ3+GvgohYbWt8XbIn9j6RKkr6sPlJuXoy
+st6R+qj71qD2/5A05VH/T0jLyZR5NfMiSIjpGBPgh5xiOssjNfgt38rkphe4EylqrvPOkAtbpPU
g1A6/P3f9Qtu95BxlM2fmjaPesUbleLzX/UWGVLQn+QVUqCUSml0fOCOVCMWzhxsBM+U/0ZkzyAp
nuxZxmuptHVAnvVGav5mhooRPRBFeSi4fMFCVXyoK7xkrSx1WQRlGKYJyK4gi0JlFbfTP9rhUKpY
gspWergoQEKdfsNLVtnE32J2VCGdbFXyf3OY6BbwxEHw8dMbNQcubaEm/xPmMlZFzx1KhmUhmHvf
9ao/uaIfXy/5nhSzKA1YYpBKwhPAIbhSj7tDe1UNH/uYHwxViEdY1cNkyCXZ965ecpM7fK7bNbki
JPSd6ccTTipnD/PFOQ5wOJY1pBhkmt0t2D1LPjhAPPfpo4uduHNGddCFHCaWvZR1t0UxevQ5IHcD
JWGKYDzoSDnCkvPpwOE2Gz1tn3Ia69KUo7oSVIXO9vxNHryjE1fO6vKQLkRFJuYNE+EhJ/Y3jq8P
Z0jW5lmy/NO576Jrisv+Bi12mKRFluMFZLEzUSARTpO7nEhWg5higa5UVKE4ihxAlERnaCfJECR3
vQ2ikWmCz+TwqMk19NxKoORMe47nS4haCRoIgc+tflPkNKD/WvT4NVO6kc22MIUcE9hks5rYZ1K8
FU9VVr5ffKLeN8hTJOlLouFyTvIMwXq7TSJ0ddc7Gnk5Dbt4HdWe0lqb2sGrsuWbO718GfNXj1ui
eN+FXuTadBSjfti8R6sU/jB6BLXdA7QL9bJWP//ydEKHxJm7spIqYeX+6OOx5QIjN7NmJGOGEylX
Zh6mkIsV/liiVUt/ZHPVdlys/RhIfgnE1kiBcILC5eg0TUKIIH5HARjs2z1rVVWOgvfaLtbgbu66
AqfrXB1qcGN/aEnoc5NkVxw51XAzQ6C/QTmFRFeCxrnjBHpKD0Fw+amdtwLnKP0qWOaX2bxx6FjB
ZZ3Wok0L9tI6pgk7nV8zCVrPXIQVT/nrM/KaVsczTNC+HUuL/tR2sG11rRZQ0375X6qIs/b1q/ZT
7w5eQd6EoHSQaHhjf8byaN5QnuXoyR7wkCNA4LwFptFK50SJN4inf7bxdWX+rCVcH+mSqMTBuFcP
HhfUbAVMbSj36x8AkmrsOIsMuoDusGBNbNxWhPGkfsMyFbao1LBLaO/hNYXq6XTAizhJqUC3C1O9
DHPnR1irF05nkCBE8edOuQSyI6O6/fAWG+/pwU1+NJrHfZZ2bzOMuqxm6/lChD2KiiJ1ApY3vC3h
V3p6mhMyvTZ0op6NEUwz/ooaEO9UBjWkXZs5ZPLey0wmBNG80BU1lZtPVEcbmjyAXIQsxSi9lH99
+mKaGdpGT7ealdXM7vmIhmCvB2Tvkhbsm3nDTYefVq2d7CTHXY165GrydS2/BobBW1rPL3Y5CCz9
scBfmRCGzTSLwiTeiarwc/tcpfiaG4Lvpbjh25o0n+fUY7JXAx2dsihsfqA323pwQEFd8174qOJ0
PGKcgBACCqz+jDMrhgDFIsHIOjPRw1CG4AwIwAGeQT6+m6dSL0feSCfFl/oXPHpFdOp+5yLgjidF
WiUqtiLXA5fAeAaYrvpgf53hkjDvnHAaa6ics89vOvn70RN/2zwfdgOSz/6mvFz+VJYuhs17J5ir
JHPXNYBrAiXVbV0jJDIxPLILYd/HIIL3JMjVCXWzY1l9ZECl97NqltjwfDVYW6qqdiqiWdbWv0mB
ZRhIYH3lw5n+DdpexhSbOwqnOrNBIBRJypyEQ6lgACYYs9WAg/YO4uG/ez7Lhw1Zt5m5y+IBAAQv
S/avZxb/VbaktNEyA6C4tukrNR33Q1c86fWIAxjFD24/ipaDhTQEvyUw7QnyLQwHdWg0kALDhh4s
idO8WcOD8iGrG1u90WSTa9xnwQ2NBZ98I+hvehgmSh5wDTIfvjg+8TGvjUXJq5SUe6arUTgAGQWe
zWk/bciEbiAkxeuScL1D7R+Qie6B/HLw4zqDi0VG13OnPO5ai9haRU1hsMbJbWi2Wyhcr/HJVzOV
WHiROQgvmMPjkCAXvwqpScHKzZxP6ZkFDMdLk+xpW7f/izk5mTv128jFBcDdqnKY7MUZ707iJjVW
KJBxb2NRqDtmC7KdYZD640eH51onDTQeuPfpQH6TB2/rSVOB+7vS66eA0kG73pr0Gmlx7Px51jtt
6JmHxyWaBzIBLpU94Or9Ue+SGtJW0UoM9Oj0jxfT2qjxNVFCGfcVcnuIyx2osJy9dMwjCZ+zJsaB
4pi5pYC65D/KKBzTfo1JS9rap8oxUUUp78ABBXjTP5w1Xk3Hf5oWSl100rnKCQv+Z5f1szm41COd
f2mxof5NIlgJeFRWlFEIyPgdTNUSA33SvvbLPI3Uu2u9tDvXmCQvKSmAzSWQjVbn1MoxLlAM4N8f
j8FaODYMZs0/r1arXO9o+fwdAmxWGG7MRnNfyXr4VwQyjQ7HUxAnd78ML8ISEBu+r0d+vcRvzQ+7
oxaOSXRCaKUu/3/bQekVRDw9d8mm8UgCAo8AyFPTuAsCNdEqW53nb9Z0IJnX0ZS6cA76ydZbKs8n
4LfYbqMToA9aIjzXrlnOs0u14ETkAr1Zm2b6IJESDUqfi4XqocyTUbu+Y1cQK277D9mEYd5tjLDx
Y11P49bvUBlU6cBuBCiuOqTAwegpjtG9u60i0tp7eEZmMX0f3QWTNyuH47PI7SU6CTwN/lZlpzmK
Ht9lxlWrb3HgHThbe/RFFxhblxViFVM2QcF7LZ1J4Evcaa6stBdXz4FUpkF/mxXW4LnZc2T3PC/0
iQtve74moMAMXT+ACtLOmPzc7tT3TadV8r+m59v/ySM/5DjbUyI40aRib9vO/Aq1NTY/V5Lqu2Pc
AMzUPQS58KJSSRevVWgeX9pQlvuiJb1uUOjIP9DamMiM3HwHhl3vN8woWDczAFeSWmlDI5U90xHh
lNF0UUcXB/dYDGKIfU8OI/RIvnRYJ/t9TncMEAWwiMgeVbqPDfLr9Z3Pbhozgvyb9dm0i++7gMbS
JWc5u3/6dQQ5YhHXmOgBaAUdsFWWIcSN3Y2x2R+Uum86hD5E6v/cfZTg14tSZ65/CnNhoVJxLtxD
3yvfPmKuC9HeeQNeecSD9IdzNXMd1WJXJ0Vw77Y1tBn9kK3/odyZi721d2ha9bgY2iICGXS0eghX
xq3CM9jlW8jkej+OlZQHykcJfbuj5tjow8fauKetVLYw0svEBDKhXQgIP4Kl106xPSE39MVCCkLQ
KMX8b27+IWFExDE0MYoQhyZa77WzxLtQY1HNzmBaslY3VGATk6GHG4oLHWOkr6KMFmLe9SP7drfe
PQaGiJyKFOg4I8GDTWmT0bP1dbqB+OWJJZ2atpivQ9teCu4pvvHStGlycdFV0nMNdinad+F83+hP
USXCz3l9JWd9dWuTdubVvpP2UUF5XvMRw2f+8MZDGe27STydIKDwvG38tFfZfwFyTrIzmlgbRiDo
Fpz0/9j93qGD9lBOmTZDMRP68L6RnE1b5SMQ2zW0iMIhRK1bLP49rxJUtwG3bTZyXZMxLwKAFr/R
/UQoLhLkYhh3tzxEzYzFwFpentufrUDWF9y4E6od0FtZWa3kIoPsh2gkXueX/R0o3EODl0mZPCz8
BaOvnVwpKC1FnTxUah9zMqGQC+8aZtZmvx9UPla0kKBZbbDS3dwsT3Gf8xyBxnpLk7Wo8iWgfchD
wH41jnU2jJ5W81mJzOvkgBYwk2IEKfmT0YmSBpg9MlXZz5gnlDDNXAmgO3zRHiXaJZ1iUCMzUZEn
n2P6oek82FoRFaXyb1Nhyf5yp1NJu8oWT2VgfQOOjvs/+Z74SSASEsrlC5Yt52Jbb2fjOtUHo3Fe
QGoxJfQNgW7ViKj7p5T/b/YRyQ59r46tBCLmpR4xR5iMxYJOub4BNmQUTUCmyxLTuXL+rp8bjjH/
Tkb71pDwroc0Jwa9/tT7oodgbNGRQgPaUhTCe0Tfu2MN51F8fD8kNkIS/292Tk0lRbyDSS2N+8Tv
zo/+Zne0MoprwSjGGV3aLZWf+EBotJErhXVJxJckgeXdLWphIi8hJ3P+lKbnyZvS9DvpHqGdr1Eg
4QaS6ahnsyBHLh4/EcG5q/j0rWB250uecVblwwskMvqqhCm5aN8xoTI8GblUS+eM3DkExVGNOIRJ
Hb+0q1v/WfqavVnpKfkXN3N/azcXJZ/+1e1hUWsOIERGqbRIq5lur4EOeuSuCaXjWUUh9OZPLWDW
vo1VkPeuI4Ksc3py17VPR+M+r0h2scOiLIeFeDRcdxqQUsziiQu+XoFqm2lofAXbIwB/HTU10fzo
6U65AD00qvUv1yaCrUTlJCSJZ7k1qUm6hq52zNOiCW3FhsFzZFEINbcMnSKurZlt6PzAh95uCbzJ
XHNBT54jHE/JKu9zGB/xfjay4fZOTiAoaAVvao98gWNbEiQVdXUst/Z8EYtK9rIS9pP4Cf4yv6cp
xZHCI126gOXfU0vqefCIHcwdzOEVweOy1zyWleglvr8nLlRjtRe2Gkpbw4P1JpnIvfIsVhcPWc20
dO6bWdIr1Guqtc/yx7m2NkVCZZ+8KDDyRHMdBiL3eyoMyNoKi340yV5HUE5KgTu0LhbHG92NfPv4
zG+eeEKQNyq8UufBTFqk64AOovI/dcVIAJWQrG5SCNNU6U1shlHbHGjuKhptzhk0OSGEBeM+tFtv
VuzYuib6+oEBxR/o0DAKRkPKIb9eQ+T08qbOD28klMAcMq4zxvcUmdrN3iHQ9vOzk+TL7LWuMk3T
R1VFAbsLPA5gitAjbQV6YHYTsWL7+xrmaYBQRXlXL6zu+YMTFpv11jV+JgTLrS8OvphwrRp+Fdcz
3YNX3SItH3NO3PXZYXkg9aZfSuZCixagTcFTriZjqgimLpr9n/mYRlEC4Ah1axBv2yIcWWfEANqI
x2ysKqNDDFPXVsKkjeiB/g2Ysj0JL8mhAaA3FwdwqsxrX+3vYHCZy8ls5Y57tcc8/7aJ22UNxrGi
5w4auc4sv7rrn/pSpBJfdJTECzhBq8LpioPd637KRhCnuT8Itk7UjPsIHHykxzB9lxLdF0QT5x6q
7S1d7S9ksBaDCd15dWQykpb/igLKFm9mBEXYulICfRK1sGCrXiLHk0v1Eu2rmFEd1fwzJ7nz5hfC
lHG3RY6SZA6kUIAsYPHj+4QqCDQCy5T07JQXBdKahz6dEvO5MCwJ2b4+4Z5EaR8OAcI3+Gthv3+W
+zlCORpfRn1qcpVB11ep6SV1gmUjq6iFuxEJE5hg5lpM1a7fdSh39C72+S0SrzbOz+S3Y1Lg36EF
AkdPMZCfIfvyxZyFEsiYV+lHdYvktqliZSBB5PnE/93ifp5PIBq3Zp829UVD/nt+2Jn8D7yaZumY
354ssMUoczlt1BsCWcTnhxqK7tF9DmP0e9yRUrn3re4pRl3hYPmTAjyNBlEAn/S5JtjSbY+/nOl2
M1+lkuxBXSMVJGGMpnEXKiuBrDqFWkEA3hYRxwmW/1+5tgl5o1mrFiqp7mrH4TB2H4VCQogqFUWN
tM9yIu17ZefzBXNpP9tTUBzzhOYyzeJZJNNov93/cAR4/dnSYMO3no2+N/BwhZyWnm0iFF/tjOVa
2nAz3HTREZ/SJVFttC1lPYiM0+u7V2CT1v8+UdF12GbY6S3PfY5gjkw7/MBey0SiUonIexSFWl+f
NeuW94X2u5uFVGqcAhiL/D5NheirR/WEcVGJauI2zuSzLlZWN1hfCCOk2UkJUsz/8Lp1N16cwjQi
6dB8m2cQkR730p4Xfe3Scqrsb8zstsEELdy/j1rYlQRSNKfQeW6kD8x6iD+BRnVv4C22sbg1U5CE
wOrXay6xz0fMYHDlyTEAP0WKMqSzInFTCBXM/R8uvKvZvjSoAIgO97mCwlyYGQu9htwHAPTOAT21
conWzeMR8jAJOIlvAx6XRY3pJz3m9iOKv355A7CYYzolTM/esIFKE6xXDIesthoKQ+xIfKhPQ4J5
yu4EvyBVER96WDjDuyPFvzcxGlOI5pmbjF3rhSllJ2q+L0Lcfrk5CP/ph5NZorwQJb5TyYwjD/U5
Otv0plZpxmzZCpwftSzL+XAcA9vd7bVO+1KeurZ/y/fDxqHDAmBGFQ5RgnOlMVU0Olar+5hDWQXH
bIYhmrSepfPal1P6xdg7Fd2ELemBxy6ILKsaVi7ZWN1KztauPJ45drSkKAzft4kxZczh2WTAvPnl
MCpROxOazhQ3Z3sV1ntmibmYcYgdjdd2IYqndj6OF4rPNSMTPFkHa4PtkF1SrqbCVccTbfn1SVpd
gZAYD+lTl0q1UV07OhICqXW5y207ZywoqOoiJAWw2jsxzL+/QjjNc5TQEhkRzCf+LrbNmC5bz1vc
dJpx+AirorYUKXl9bCMCHXeO8j7MrSLj4ZF0YtIt7xkhOeFvt8P9GMiS7wtuHzbpy+kUMVgSuuI5
WhC/IACucfI0DdB+8CE229yUODU0V8H7nLdcsvfKXmclP4gvxt8XBcHdvxHoo+LyYVvc1TPHD2PO
hg6fgwaJ7gGSI8U5VZHBlE+0k9uRxNFbTjrNi2cbX83OZ5cix8yq9Qqr8uPHHd4E8mg4h9SqCjKI
9sTwdErcHv2PVKeWYrxoGINQOwcLkddwkM5hOt20HliHw05WaIph87ZIFUOuroecL3ZswfoVLUx7
AUl9neP2bqRuy1BCfC/LzO8s3K/kKe2i25KCanygrDQ0+tz0tXSKXrcL+i+7GLW55t7OUA5yvfKi
Ouu8SvLDJN/AY4BLHVAXy46emuCDCUF5dcc2sDW3VD1rcd2zsUqXia28C1oIYPhJ/MwldLEIHO4d
4u49tniGZMrHqYLPsPfxqDohdWkA2WVS2RQZBCgooSK+FfccbEsrS6nnl6pyQKnxx8EVefiEpiAA
QzpBVLClF2dOC2jp1LM7HMEWLDiOX0dPwe20zPv5fhOS+BaxBm+uhujiIeAXXerLHPgdEpGJWlLK
uGmaGjs2ZCV/qmk1eIcaicVmvbsxHbjwnKiBsfBbq3PehPHHWDHAf9goI+GdonrGk2utpRABDs/V
lddJriNbqssiJWgeW9VDHYjeiztQLnx7iKT+4Iq3TNdOZ5tkqnLfYzhJyXspu7hRjFTXXiAfi/lC
rfh6XcKc/xZ4+c3sKDWUZsDcPQ4nvcm+5mXNr5XkJDpfgmxXtPa3Wde2hFlfgvT7bJdAhwcMNQJN
ikrrzaufmqLc5bSuT2rjwHR9xNTfEAmHpZxr0zGJy9BUxJUa1BON4aVvFSaQQHV7tbjfDV1oLPRC
AyGKiZHm+YV2mIcZvc6ZnXFONT7wxnDZF+1zxUIKqUKgnCwK+tULR5gQ4JMgOtia5BY0a5LSXa7r
Dqisd5IkYB5KaYcNwXHDHfePjwzOZNPvXo4NyOkYHudlA3f35GDePHU737V6CKe/gET68FhbGOeP
z342XXQaxp8G+htGjM6VMZE2Nv0CcygteifuQai+JD+SHngnYStNH0ImSpdXEO8kmfffRqoRcJ0b
tV8zDg/Omm6Zbh67hcnLa001fJqSJ9/In48jCpnnwWNx70XOjD9iq+pPO4Pd/9yZ92PBoJ57tsaS
4u+AXYOHoDdm1e02c+2JJoW897AVJ96g4llX2d6sgt4D2gYy7RRdoxtnvNZdzw3qUrX2KyEhpzNN
14g6CmVFF7s6pkp+R0/9ggNIyb/aM7vI4D051Tk/b0rNEC0tzMHIJtvNbOaujbGumrdFecBPMZUb
hTQBs2g0lr1KBIV2mnxwA6BP83m5OwTS13h0Ng/1ToTAaG3vSa33wvJBu6mi05OLSqD8qp2ukWkf
WDmk8rXiQQbK0HtZi5TKkfbzogcKwCSzbjKLuY/wJFS1SuKvufdWqnZqU2pIvCNWFnrnd9pVu0Fc
SjzUcTRy4AVyfxPp1dHqB5iySAOJSZbh2rYeD8pfQM0IqiYvjXKn56QIRRfZ2gyxpUZixSy/8/kA
xkeGxD/5Zv9jWEv5klfSd9TXExtDK/v9a5n8f60jzWzbyM8ZWRg6Oj/A380B8Xc/jyZEVBsYxbpG
nAK903U0vvWGRXkzzGVmbOIBqjz4oHT/5NWy8SvD57zSDyymQjmgtoIT303swdpSr5IgFhrIi4S2
vvx+ROsYCadc2GLSP34/Kil5xgsL0HRxG/FeqckHO0Fq80slnu4wVmQY3n1Z0UBmRydNSVycHpaQ
zdoWS9B0e78xrq0lokqPdouY3AEi9iKdLQ8ySYefIxoFvvwlJW3288m5ujWRIdFaLL7prAF0D/av
XPmBEr3G0czxtZjIyZFJ5KVUjCbJWwzFfryr1BL8sY6+c1hKDZxfaDadmwdlXG3pq85pvXLL/6+G
PBf8pIokzjJVrZKIJG+Tg24s9Nc3xNSvUOwoLiCXdZQhcE+X5Lfv2nsR1G2iiEBCx9yDWqWItE/P
Iu3Ee3rDLwlxlpCkWcAN8FS1GBL0XZn7ZVB6kwSHb592IczvZLFP8HjenwLFmUiutg3oyy3sUJY2
K+/ZUwpQS52S9WIvcTXrK1owFo5wnkb+X62AlkxYuA64GIZJ1Ac5UO1OJNO/NolLKVDpPxvED4t/
8ax5aqu5K/oST5OmmlKbXrQMHcFcVmu+zzpmDIX1CGk8xs0Np1vk3zAEhyd2gN3KkTD9WbyYyQTj
B/SXQMd+Q02xsoty5pNypaaFvAwUq8TzFw4xoReoYZWW3GALUxPU0l0nCLacsxEzGYj0HG50s941
6B6HNxv9kyR+SmYxh/ysBGfVoAZKe9hRmrRfpb8ORi4q2VtcrPLbfxCG8Q546c04rxSy1FIxmlYo
rpUtx4ovMh6ND4UO89JzyX7Yx/LpJv5v+JrNoBAzQAaaRHr6Vzr1839dXLD/+lHBciQz1kVGzJD1
UJp7xSp6gi01awgLBJqRBaXIrDnGZEqpZJtUejxW8CAj+UXp4MO2b/OUKP+5LJ0uVYmnZDkhoGbI
S9n+Drfw7v/O3AJLan1UJZK+JgWjTgMRvloImOPUUAbbnukaTvEBeRis4absYf858G5GQ08BZhId
AQ85ZdXjxACGOo6FXdWvZw2bolKbffZE5lv199tAuyfOFUCs4EIFOWTiir8Mtg1+HPhkmkOAt9z9
koztKjMCbrJzltvHon81mzpmAiUqjyKm1IhkY9OCi4IJJaVicldNcMMJczvgRzPNfJooLNbXlLB2
dvf+YsP7xNUI1a9Vse+oqStV/7I8T+YGCquY5SkP+SYh4cg6+7c5fAkYqvC6crVsLCljuTQYI+d/
tyF8psDd4qahxU/FuwZcunSCcRW/Vv3uI0dgtM0thAKwvtzdz0LgO0rtSSBzv0ufwsq6fe/2SKFA
aZSZRZ8LPeCVW8erRUPvjrOdBqG4ZdbDzmd6NSQ0M2UGBHPAgT7+SVadPjIyQdD405r3OhX/Os/j
eX7bfBbGUa9XpGesaydIRN/4wYYHpPWqhqErWKyUX09bsYWwidIK/5/XSVvwiDYA7M4bHeXvV23g
GT1t8bqRMcKYAmqC8zHkiDaXO46cuMt62NNfqZjtvy+NQnE7S0Fu9BJsm8qdUI8xuX1fHllvD5WO
/Y7Z4gcmgGWvhg0ceOddWw2/vQWI+D0ggOIk/S+ll+zRYVUHhRvV1oIXy2mQ9noAn4tteubSDmj1
bChzSVqtfu+CG8Y9qM7PZhHsQtoBRBPcZIUTpG4UWQRnGXlqZWPXICgt3Zl2g+yllCADdzms4TEP
U5YEzsCqN+b8N46TyZb1yg7mBbZpm8fK1uH+JqHjIA2+hm7gxideYgAvWtLnCqaRmQe81znapjAq
z3KCLwESaehWXDVStgrVrN8WjiwbBkSgL92t1D3W7uyLSuoapzDSSsWwfdS9DG7BZFQBH8zdiErv
0aDqKanLy7sfO9/i5n92g3ZOkOOq37Uz3dXiXqN0cTHNoYkn7da2JqP+RLOhWCtzg/KX71Vp/APW
sIDs+HDoOptfN4rGONeG2d03ltQ4HyrFd1re/bdojQVL35SUlMD03IPfPkWxUGQX7KFY+iAywmWT
xK2lHyTntmffCwc5Di5GFXjBoHs1q45/82h9ytK6hrQIbSCOGc0i+JODJhKUOhUoI2e8H1Xvx6R2
/Jw53YHdDJrxCDAfVj2YQZM0jxL9n19FApBoXD5UIeElls4yVfQ1u3RU33hlVUbujQWi5RVmUS1U
32DjJAHLve1cxM97gsUMWQ3r84WoDZ54DPyPkG8taF1Tba5gKAfCyxxZoTfTkPmqyVTm/yxYM2uZ
jzKVJ3TmlhBbiihR/cUv2W2x6m07f7JpBt5iG2mPcJEirUR7vkjkvzIT1l0qa00pzDSnW7dI23Ea
Cnl3YKDHG9mKu7GPOPsT8GGtTk+hSB30j4urCAbniRoFFvT3yjvOU8F9ufdKlS/6i3w1kMGFYKz2
I+oVgj+EwhZUAuutyWXRCquvqRxfCDA80Tvd4i+pUKBNuOxccBZWLbwJRO1I7cuhPEVXW38ggeRc
RHXCSJ7uYqDkOUWBIxz/mGrXy2U5U+AZuvtx7RF3/GLBPA7rMY8Natr+85KaMO5pZ4cBrd6ShkUZ
RZcYhZEq72Ic0h8wTJEvlptd62Fv3D6SHM2jnbKDC2h4E5JXKYlG7iCbA+mOECOvamV6mq+eSiS6
ff1dSc0ilm4utz1kYttyPtqrWs7JRyFt9SErSpNO3qO0hDOfkGSwc0uxFBt5W3Rv6FyQeD35ioT7
MpyiMMsRELyb0n4k+il+wPwFET8nMwNNP9vy9fDsEaeUIU4VCdyVE5FFvkVmeQhyU/d1V8CIGUx4
adnmL8ZIZALTKiwOew2aAoBwFhvgbLzOm8WfC5I+T15FIc13bjvrh1fQT7VQjPNMhZxGDqn3NSuv
fLaml3QOZ1HX7G0aQ8S9QraJVSKY/7+zPjuIvmS3Vw/tMM2CAszxl7TBKvAkB8Mp9Qa0BQlVrupT
+lzQQ1OYDVy4m7QxBG+yZWhDNRYF7fUdxPBlk4vZ8Yl6ohc4sWg0CID/Ln7C7MprOrlL4b30pFqx
DIYhkTYI6qu1917ADEu0rfzpuc91VA5OLKQYZNu5JT5hhe3g/YAD4ErBf006xdpEJes2U6rLHCdS
FVAMpKpYKBvrWLQH5k6pi7jkDzJBYGRatG8++MQpbzwW9+6nHDobbK+37T4VdD+VMOPKLEBDgS4I
SpMPhr3Y5e63EAA002+U6C+uLFEXH0M/zmr7K2Rk/yEx3cOwlOG1ZjP5+f/xdpKlT5UQrkqzC7N9
t6bpWYQZg7iqIxwui28zkilKQUm5Tzxh7XO4P2bWDU8Gb5tVU3sIjonfUFBxQ2KR0oHio1Eeppi1
86Vm7k6KW9MgEkCRAg5d8jM7VYHlQTw5ZwklTbEMyVHz6WMlHd8oXFjX2CdTGFrJckQdjdsrgYL3
pBLik/07wGM8WyTigzpMw/SjQnLWdlniuhOlFHn7bohk2NTeX6tNWciLPbzERtTcRJkGur7Pol7L
sWCCLtBqw4VK1PmvlyIo9Q7EbAW2EGzwm2pCuSHUYXCfiIEg3hudt7kwXGwOKy44ueici0wwu/hF
PWRh1TjbBY05cMD7gMAx/gopAch4F0GtX883V116CP4alx1UrN57Mhyu+kQcPMzmfiRY3SyLNwQS
ItLOmtkzrj/sW1sZbozbey0n6KnOiK7Y2FCzmwlCC69LwnQM1ooRJCjBV72iFfp4SEp/KT9NzzSv
8G2r3oC9l5ZGHx5ms5lj7eUxEWYX2Sqzjvj3SAzG7WI1Alix93MIuqMfrFxpWyZr4Pib/SUuRfDZ
VAHl/n3PNr9xb0TMfD0Ahs38yjNwJqPS4Nk5RusOqcK0Qx8V8v0Jc8JqiJFPLcgv3HcCxCvdI/lZ
VdT+q6vB0kvDNqbd7UtKn21KxkiRPljgKOQyeUALqPrRCYFLkVhYpuTVsSHNhtUqWuM8S4gcJkQM
fiC4owAkYTXnRRaz1O95NzFCCmTA2xs0QuSIyD6jXxnTt+TXIgfGV/+8GawjcY7L+E1dgQZgGguI
nOK+ZuPiKQwjtHe5a83rfF0gbmaat52Hud8+oVQQMjvw8pmDq/OKlT+52BEMps261AkTA3QYRz1Y
AcgN0xmZ12qZksJh/e0Cf4dchALt9IObIiXG8C1JzEwHceRmrhmtGLC63angC4DbdAhnO/9/muKv
/ptd/sZNusq9o/KAg3vNH2sTjmcRf/9CuHZPNXwo3u3tCHCTY8XN4a52jpBBLG5NxeKbvnlfN50Y
1NmkEVw8gnoe3Z41KW/jXtvSfoAbIrZjSAtXsTmCaQt2wgf4U3uZrEQbcBiFz/mOlWW50olF+fkj
CnqY6B17tHtHTXWdNcAGvpcJ47/dpN9iyrymX9tioo6nXiyS19LeYCULwywuzVrniDyYu4DAPZb/
KkSSfPoN46TJHd7QaZ2UQKyxRLZIcgKa+g8Rr2HfIh2WXProYsNCxnTiEx2IMYFIkOnw7Vc4eVpn
Yu07viGNQIpkwF/0q2egRUuFIA6NDiR+/vKVxMmOlUiGJoenhe7Dq7x7Acw7hoz18kuE1KkM8Mov
1ioiYUc8rC3JZ8q1I28Ha5B7F0gr+P+BTeFdyIDrpUmy24aCLbDL4a03HNZz0ybmRg01f5uCKkKR
X+LTf/f2l05OEVu2/PDMKG08GJ18sB//wYGCO3yFQQlnRgnFABn9DbpFfS44OtwB5jKiZSM6qX1M
2Q04foVyki8lsl432kBbUhIyEf5ym+fe+ZcayBZSz3m/teg9drlpgxCvdEWHg2EzcjHcYYf60Cv2
6LjgSU851DniObcXa9qZyf879f8aC/wCfmltLzlXJzhoC7OGFMgS9M4+jcrApDdvXmQ7VKMbbIL0
FKymNRMKBUkx5v9LGOEHJyzm8prlCn/9QlpZeXT2q/8u/kol4SZX97JHp2oTRh71WVhctK8iXQio
Dd3WgApI8me/zTzsIIw+OptROQcI6eRZGyDE7EXEpo9tUeHmyiL1G9ysqe95KWYyeqchBjiKy+G5
pDC3rSTi01FZ0jeLKgtvGbFiQR5H+sLu58KRUF2o9l8Pv9Bi1Ydw/Rfq9TGgCCCoF5OJ24fT5aJk
YbBW/f/ViTce4m7na2uFpg3n+P7BsaMf6qdaXjJD1ckGagGT2F/K4DvKKMBVBDL5dT/CliNAqhBv
9QrWXQQeacanrAF2q1513RilBgczYcYXD505fh4ea2GL4M4zj2IHtTxTfB1S4pZhMqChknRgr9mH
4nSKvh7xUcTiXh03erJZzqdckYR34ln5gz9h0hyvKGureyxv/Tre5APrDFjokc3zR5Kj/MSF/OnD
Hsp7xHSJZyBcIyi70tCffGh0bBbk47sOFBTrPBPKGngcY4ZCUncp7gZGbId15Ri6eJ1Icl0RVK0+
ocKMTxAmbqBvBGfl4BTiHgSfxIPZnrO7WcvsYPa2WBJlBWFRhnmdjb1bOnDIOXsWw+P/OGJg9r/9
V62zi0ONT2l1czyNGuzZpALNQXExrV1nGVQzJ586g+U6YV9L55WfWJm7kDIUgnj0DzLkynqq+Aia
OcalV+e3oFUh8lVuNh21wMtRP1jrEG4hf10MzJWj2m02RkAczmePpWDHGy1yDWexx2hrz3TUY1Rv
NKWOZLvULn359njtcSgwooVtyF8yqZDeRbFe4UaHD5KuiaP6x8nuss8z+050PU/TKeV95RNib0Vr
+NQM4rr7Xf3UNZdrjuE4CnR/KhJPTX4ABlOiI9+WUF96p48BbelZB9VSJ/Ib4WAN/8a8QBxETcgH
HqGNWedSyAVVMtbvkq5yPWNeVvq2T/aVbhSIw0b2MOUciBGUu2GTkECyCKdrriT06jiOYkcoLMOU
8V8r8M3LZS/NAzu4ybf1tleCU7pHQdYjTWVd7gHYUWiiLvky9DX0amvIv+RoYRSbIW4te63x0Epc
vHVBx13tgAQbkJX5x9fP9mSMIuYzaTr7MNhFx/XutWqX4Pfj+fxYbONgBXXW2CH30CkBZsVbRN0w
y7YE6cEp17K2gMH1irN6J0DJOFo8cJhDLiSVnXPPkra6dnZTCfURlGC4URZe+aBg2trCxBHf4QfG
ozvxoEQaEVP6zxYmC568ok0r8RstDN9tBF0GgYKbuW9py/ISeURB/DybIlKJTNWtIbkOAOfucjjF
0AQsUDhsLhozPB0CmeVledsh/lHHVxwe+C+qZlo8ykKu5thz1Wz+SHbx9ac+WRxDptHes4DDIlGl
CW4RsOTWjkO5460tPaPTx8y1T11OBF/THIojfWvb7Tw1lQ5PzWO8Zxf/hhvraX2QJ1Vf00Z3TgZ9
+VFPrfs/fX09N3erlgB0ECnb8+P1cX1KlFggH5uRJtQRUgopbn4u1+/amck7cdHHmEHmErfhVQwm
FxDcJfetrAar6cnKFK20SRDOq37b7y1bzFVJq4oZ01mX6Xu9R3XnQJ0pPL53+klpPd2pb2ll6kI1
hWlpl9x6uSE2GX2wbPIwg0B/M10XUu7lkKkMcpZJxwVbWFsKlOizrRnxiTudhqAKx/xvop+abai5
MqgBihPgEcpmnOlktD1+vzyBfxc7xH21QhyGaQr+2lD+6gZdqhkKEOrgfeRt7XreJbJQ0AaGL40W
so4DCk8WFkDMebimuTCISc1+hnZ0NIr50sDEYdMt2ze/PjwLItrB/lU0E9Z5hgfQHDg4NSeakzfV
RqAPO8KK476JJ6jb4XnirSXHKj7jLqE0M3XXrDIUtndVFyUvFLWmMhGBXeiQE58hkuZl/ZKnZbPV
AnZP+mnTcxOAXWxnKUYBhJmQwtLuXGiTLF1BzCr/Fs5EeavrZYBQLNRgMIQlEfCoYIuwnX8Ya6Qb
EzBgPe0dkjf8pNqChBC9MS+9Bh9P+svOW7QLJyX6jyoC2dQqMrNL77IpHozOnxVuihLd6CDyG9SS
m7SvQMngq6OvhNEwTkL0YEnYHTbm2DcSLWvyN5sMcS3Y53DHIOLfXnAN0Phx8JyFV3WmjryJXs/V
Dl7pS+6OZoMrEtPXuXsnwk5Rfhf7NaZOrA5wGav8DxkuGjgFq0Sz19gi/Y3OPAl5VOd9lrb0Drz1
AOOQ76wgBG4X4vitX3+fV5LdzV/btIP+sZ9IPNSQvMDkKt4Lk+xMo51K3tVocvFAGQTTXQL60tdQ
vgNUeWSMtxbkbSWXeEUoIxqm6nVu5ssI4idBJCdmI2E52Dj8k6Hlgkd2sCPyHxXvXEiZArhtMUAA
8FK+LaGhov4a903Us4IV+oOAAV7jf/LgbsMnXC/t3oqQicQTorVPAgQGOCJTJTtBK5CyMuzOKo8P
ZAUZdf/X3MspOMd3ICz+8iPCHgIPz8E/wVyJHLEQncKmmHFHC+9DujksvgGXzGdgsjucKZ8NDzHs
BzwbY7iwN+tZRZeLhUW8JTJEDN+SCLh/+qNFjdSquHaWMZGadxNNLwHE7MoVV+CH19tifYeoKAsO
fWAL6qqNK8DGKMj2HEM14ivbUSDhwPxiemkyNsd02R9YJkpIIIao8txhbrw4ndWW5+uuPS224nO5
WkkWXQrA9vgauNMCx4/BK85E79Fxqvh+S26NiGNKba6yqjy1CwZsNsUA6LV2NSYqFjcln9zjYI4c
YcuQ8qY4wRTc6OdPzT6Gice0FCUeZOYifqeQMUp8C9pTxJjvqvvCGVrRgcpYjcY4RboaK8Saiju0
pbkdgsMwY8jdN64DL2V9wsEEvZLvwuDK7l0YYmQlb84hYoiYnMg168l7UhxTx6iO1ZH3SY9Rg9uW
NVWLXSjH+ItoLMRzSgGPMSl23dbmC8k65JkY48Ozgnk+sWDpI08k1Z1DJzANPcITTWvRRd1IBGk9
xsINOOjD7mY1fvGOHmAtw7hl7qg2/RFd3UKMJ/fjcIRhQF94OOj0j0XdFHc8iYkvlgjT1j4bNJCg
P/H6t7LJmy17boiIjJuMTVR+bDsZKypONFbdtWKvvhGB6owHJS4QDCuib8vpHkVacui2hvKQD3ZE
bgIESTuxFmcLvV4i41RVrBqhm/ZVMOCUEs0Nqdyj/+06fXhusHCjdGfj/1GtrcG9/tFWKu4G9Ulh
nEHcZB4cPuXXJtop/G+RUVyTWhqV0w2nZMnDNUz2vUZoTnFfbMZAjoGpJOo247d1LQ/AKzZRzbS1
+3aAcehDVhehAc3whUS1AivSgsnlUNoqW0syd9ovMxf4a9yEBVA06Kf94kwGh9zp7EZvPUpMIoqm
94VUHo3FbidBZ9mFcjjRS57SR3i3j3fQdlAY9wjFJyPNfvlySefcNsFja3SfHezWXhz0/TYrhNfm
/fT2V/U4wGyLzpMvOrRXj36ej3sED5o+4Y6uTHacvFc6X5PUTZfCxHuB22Q7GkWfZLX4j4zGLjbv
FHfDq1Y77BtLAniwGnfZz59ht30FjBi8Sq7smHt5VKLbpvFwi0x9kkZIlZrGUKQYGsM+79ssetVh
ErXR4y173kmEK3gjMzZhP5MGSVETlAZ4AaKS3tyuieauSpZwmqtTpwl/hc5qu/Voy1qzhzjNWXPO
0b0Jc1hvAAr/oaFEDMXwshBkpqP+K2Vm/rQuDU1KHnXk/wCtzVXBu5a6QFItbiUAlIMtuDzy+wUh
g4qWLwgza4e6dTWVqbO7laHPLBPMzphwJbU0guy3WfSnzpiH0/oCjVYIFtTdXUY1FmqzITUXIDAx
depgrXyYmO1yY1YDoReUzhTtCPUFNsHL4x1V9UUqnMNAIs7RNjEM0gmjNQWjnlzYgcjmREtozoT2
ZDn3sqCzW18kpaCLL4gwczfimIld/Ng+hcdEwwbZ2SWYNzGPOSBhV5WcyxllhzVzAdRnUWggIJc3
/SE+B0fwc02irHSuWmvZ1e9Sj7eqA8JyAbUhz40kPr3/JfN1+zbGunm4ewsNym7iVWC3S5VDUt2k
kdpy43b5OHYcieY17hE4SqdFadGDSsZmx/CkH8Novr0w2410G9OqcViAgQjZW9nq3PapP11GLAtv
E+3AVddRR2xekHTa1rGZa7osspDK48cBIojorsutGI65xSGMlDv1oEMYn6QMcoIQQvFPAcn2d7IX
KD0Z9E1af9WaWNE84xuRnumPQO/vCTTe4Pj2qVqxcOcIZxSHizozrMmy2Qjc5G66bLgG5xymckW0
Y6xm1PYsOeCusy5CCPu15GxeAYI6k9ry9Vrz8Yd2Rda6NdVJ0QI8DaFR7ohYUIaR0r3bbC1nAHWK
be+yW3J/K0vG91eWIbhaDw1u+XcuVOF0rHty2lJjl8IEEm/tjh6r/bnFt1LHymqr8gVmukcvO20g
SRrRNnOK7Sd/KC1uFnSUmLKVa/kBZknFGVjdA7m9M0KC3Ww70myLsCL6eVG+2RqWvl6Qw1Gq11lQ
cfmUCEBDTAlnHyyi84hQg+IOZ9vZP3iAVymZRtKF4F1i93FLnZchHzpgQeX+FkGHyWsAj6SaRweV
AVRnacA0r6yBS/pUoNoCq1guGXz4TlUwCbdQcLn7UFE+SWbVGdb3aXE09jHRRne1hRlQqMrhPxwm
0iHT/xfMvYZbF71Owflyf15NXWBzWmPWnGsutUV4INrpwgaVcnt7UErAR9ehVjaxQazCJ3zLltnW
oxlZARO2DPiN9z1MFsMcKTUXPBz5mb1wv4WJMrU1ld4R9THHE8KaXN4Ywl6n5rIcrO0Z1SPkHdfJ
jM/pcnbqctYb+c5Fi6cyEvWohHnICbnWKUvBHWwEW7bFJ5G8TxKvTiu8h7U4TNtH+cyuAqKV/GJW
cA5Vny48KriJu8nN+QpfdTXCHI5+AxjTrwSwqspucrAw79blOf22fwDSZqojxTFtMArI/0zK5ANf
0gqRU/5R7irvFQIr62FhfxTlNtsqLfctRkuo+MF/2h03qbAEU4vBCqEzGx4BQyQ2AH4SgjnEiJA0
wwwTBsIMV+fAOtoKVfWuD/KJjCOXrxdlDZM0kRKQgEJ/QyqIMziCKw72TUy60H0RN3uXV55E9b3j
Y7u0DEbipQEINUgQSbdwfvzpiMIKWk4uVyBtMF5INRrLwfxECum5H495jpyNHIalebj6Hh+R81nf
nHq4RD2VhtnWi1bzmQA1NV67HTAJ1MkQjZX1qL8NJnk+GZnfhicNZdx3h86M2D7OjdJ5rr+BqF39
0FN7DgpGqZEhjcQXteWROvUW9fdE1Ep3MSpZlgel6oA/04XGIO+oHkti88eKy/koNokyo0HRbPUv
8RhDIvzBEfFFJI7EDwH89DaLrN/6OeRvTDKzau00wJYA8aO07b/gxzl53xmRgR8l6PYBMqSsDCPh
YjD7iEwmZkN0mSZ1R3CDRzkCl6Zu/WIl7GnLT/4KzY7VsdLfyEdfL2PVj5WXjkowPeZPjLZHEss6
vHbRDcMmysho+6tZPlFCMNzfUOsfE/gDrJ4yp2oCzv8rb8wULwM9kid/btTvWp481s68hu3xqgP1
w9837APLyqbxsq4a6juEjDDB/7L/os0yKS8Pv6L0/P6h52fqVIn3zOm0MR7p3EYrzcA6JWRjXOIN
DdQ+GKtWuETkAaXtJV25y/mt6u8qtKhdtMQzzxjY0xPJkZa1h/YlHGnzN/nSOOVGck739tPK3o0Z
wV2OfqYB4zwmlrqjFd26hqSjMH1T/V0mLPpM/a9q8k8ENmUfPsgICPjsIHft+GTVe85HOW6s9/Di
sGhKFgfCMMxKLZ0ua+pwMekSWKpNObw7JQSI7bbzfdgA5SISK9oy2ivfolfUzB3CPcrkPAU7S9Vd
ONJ/Z8YKcHTF0ZM+3y3E10Zyun8m94gGfDI+YQSgibGejJ+Sgxqj0XWIAvkzOwtCeiOiz53BABPn
GuiAzZA9sD1XXvk+kDPNbxqbRJ5XG9QsjLMiMwF0mmpDf3HvtoVGx7l5hiDpf1XmOB1GN4weA89V
ashL90bUrqG8JAqt5GjhJneDHkocz+O/w2ooscy9j9shYwBVXkiQfl/GX4/85qN4X4rAzp11aVsL
RLI9cYtX6crNVOkGcmQXA+4+gUzGjZVzewyx3KjcxqDOZj1WhFqZC35nT37blNp71JuXGCV6YRID
Sc0yHb+6HdwuMd1a7D41fgdDexIIkVp/leSmjzTVYmwm0MrshNwVbuqDqbFO7hwEzfjMgUasY1Gv
aBjM2DL2V1XtBPRANAfyqo2TK2byy+7gpubS7bw39BIe5+LxO4lkqKuJVygjX34/tjgggXbySuUu
hFL11No2UwY6CqvWGJCK4Kd3dD5OyQqmN3DhBbdhxUOdWH8zIBM/DqlqO6WkZtpKnhUQ0n/QkeT1
rTYK6lKqYuTyo5rK2Hm9trvJxHy/7jI4x1dlo8XXZvJUn4+8jL8NVUkfh1VkpeqzzAH8+LlmGkO2
8rzO0c9K4ztPdG1WrTimDzFGjHydFb3ECGyE0WcVf+OOspNUpp7hgBAHkpDLgbSmM2aotJs+VeFq
OovQ0QuNcfID9wJI8muI06+2itppSqanoNTmW1a3DQbFSDHeeiLaB6GJrkCF2mgG31o+itIlIi8+
fOXLA4SpJna2peNrCq1PQUYfVcz8ob9DnFsBh7Vp3TS3ZgK7ylYf98lex+Pyj7zI+D0pEnMgXzP7
lSHBHOQBLeou9H8m+1MYE5ZCfa4PLHTkZ5p4YgkVRVxgo/H7zHfmYgH36Z0sP6E0sDSzqiJTvzuv
Y5hIGB1q06zozaSbU2VkMUTADvBp5CUGutv90XeEaRVgPQfMWYwxlUEOsVPdCOJrLRQbERYYzKoe
ULyVnGWi50ImhGePmvBA9UduQPP0n466FfsmFiC7OhfzJAU0WoBYeyIGsrUlv/Ar8CierD76qOwu
3nL++3ibs/PqDuQ8pxbg9AQIGuUEMZ0+aS3+4MHo7nAr+gT0yfL729XjS9UBe5okOMokqIqehstz
xCqXDdL7wecCz0tpC2J21vtY29UK9/1CaqL0wePpBEU+nYGF2CMZXMLf37V++QanUqA8SFLV7VRC
kuH0mK1B1vsqbVpC0ocT3jhQS/NRDUyszwXsnZSEfGFHmccN2xCIq7e23zjMIol8cyRWs73obLqm
o/j78KdoTuAXMIDGbxrOvgPeHkCOJa/TtHZCrgqzKf8s4Rd3cNsbbpdbvzP5pI9g05olj/FEMvxk
+aJZgNXmQjy6tNAH7rvg106NFRFPLrpFevT6Geb8B2NsjX8C+Bm6yxKjfUkxnSl6jilU6fTJEoEa
udgNtnVlM7HJE2XN68As5q74ueFfswCh3sdejWPhzSteW7vLVJrj1uYumVqOJINq0Mriv8+VwLnI
auO1TEYV7LhDQ3mnmLTLJln2Tauy3Wr7G4bQYLvlpW/KEoQJnyk0BeYrBJsecdTsCgRlpyBQ3XQ3
akx5STfe2IhesMlWurrKQqn7v7Xle3a6CUxFq7EAoYL4xy978MSm4fyT0GQoSHd9IrKGYvuCcg8W
P5ueXB93uLZXQxTnciTuznknAQjsRHHc0qI97IeYCl2iFU4PUJKM4LIv63Qk5vVSRePH3FsLmNsa
fIsbVp1+8DXbgM5U5dY8vTy5Djdut6K9rzqw8+d4y6QLJ2/6Y3+dj5jyRtAm5TUE9W+qy1sZ0lJi
x2Xx1sqIgr/0ULQ6BFTUUzqE8sCksojLGjHGttCaUZ/VTSuDz+D3NUN8qxl+JCQ7b2wdAR3OWtmM
pQYH8QjjjWIoIthO1/NKn21eExHCl4df+OLlrxLC4lywbtSOddra5JKY3KdN10A6Wul64Txhp4UR
DwVVD97xarFXBy62cmAFzOyJ5jLJmndgGIKGrQBcfo6QiOsnRFtGQ8SDFSCTKwifp5Ljp+zxyg6B
JbKvLFfdg+a/Hzn19w+KiYD4/WUOwva9HGZoQb1BlomHR2zNIaLL9cStYwLCPsLVUAQuJIWJqhgA
PymTU48F+/woNE8Xehy1hJaq8N8/cg6FLS4/Q/NxqDsWquwBwfpbS06gtxEamMLDtgLzvyr6Sd+b
iEHrGL60EjDKRSEz2YB802akzxbmr1fZoJBTbh8qYVYr5i8hZAhrr9VlFQWn5v/CCk6LZlsp0lBD
JJEAgmejOHfwuqfxu5P8dkgIr7AzrxHmvRKnRMNnI4/seX2BUGsrDIYFWjmiZq8rhZ8Y+dWRyPVb
GOk6M4aNkl1VgmW2SnOqpzokwjDc/YryoI2IGNN02p+mzrYTjfRRH9yHgiGbls0y1dwFcwzsqNIU
21TWvf/L1LCiXb/xVMOuq4nNcfqVlFjYXaM8Ozi9rsszbuRpcvU9XNNlfmIpwIV5FA9pBrRK+zEj
VzaTT/jGKClPJfkfBUwEnIFznLRQ3TZ3x6ssBILXymkC+ixPvIxmPS8XWhISV7OT9dYUCJ8waF4W
7Vdodrfu5ADXVQHfDuuDDH1qjTwNaho+3lVvNRiIl1RLmwNBFYv3qu5dCIkiCCKSY5faShJJ7M3R
R/xSnwT8xckMAp3gwwhX2bDzFNIF/D5O7ChlxPrFBXMFhLWOJr9k1axpkKGE2aLyMYvkyT0qHr2X
gdbi1/NzROotJT4RX8tX9KyFWmOgbrFor38o/RpHUDavvCCeL9e7pW8fMGtqLJ98Tc5481iciZ8V
u7kSZaPdoCuy2WvAhnk3eTwQrYNFK/MB0yDmzZGkdZMQ3bm1gnZG6eNHgdVxJMIc5i3hPkBBn8qu
NdzA0LFh1fP73h+nRn9u6etQ8oIwtJCBC/F7D855qHC0oMb4gU5WLYrpOmCrJm2fok7ce6W9o6wL
A6fMuVczEhLoYjFws1BBh218T9UL9sEBV3mVtsCp5KuXJfX4EjPTNHMUErmK+viqc3t4JMtMBDn/
0VLnDAl0gqZyq0KJE4fVOCL0I5EToGLf/DFAsRSGWwTzQciERrj0RSmDWTv+/L8RQy3WyxlpylKl
QbhjKcg4ufd+kv9rgJ1fd0fS31UQU9fe/eRpq50Lxi+4a4JPN/qOJIalZRrf+gFcye8HzM8kUyhI
bd05JgPNi93X8YIDHhRccHOp2mZEqvnbj/kedV9VE4qXk85H6ft9Dnw6I+5Z+d5/+XJlc2qLzQhM
ELg+F1bH/jReLfXMmr4ji9go3pjTV0ZeANkqkrIIjrb187QsQyFAnBgFDCe0IMIAtCtJjfNmqGCt
oURbJOJEQFsRziigF7q4vCI0cp4vvgZL9SnK3gGhQatxU6eNS6JNVwAK0fQxxwMVcuLT2+Ahn3qN
FxvcpOeJfUEG+Fyn/IpLXCmtsyTOGERNFzVJ5n/tz8pcYkI4UM62RqE29VYH+0OF1xxRFGeEHhEJ
tPDWtDiQZWY0gBQLlGJMHBM0k/y/xZg13FbDvt9JawyerLSHA3g8VChf2K63tmAnqbXKHh67EcO3
WXHV0SgtSflgB4fP+SqB5pjkmxpmDFu8u2EjxJm0H3GUOnrRbnYx+ityiawG7wBcq737wuAduVOi
rauCZzKQObqL6I8T8zn5GNJnyz5i3pPZng54JGIi1IHNWFLBfvlRfl1HDYnhOIF0KGWBCs5PbN4i
NiIKh2L+Xea6rrxFQ7m8wyhHRdWSZ4mUT+soQ/07QxuDtBPvEhHUtvXrFeaM9R4XmMiBHvyR4MFf
DVbZ7LkIGg/4g47EwnvEGRZE8k9oqHwDSgaA4lGdg1VM4WWfZJqgoFA8YcSrGXfmqYB59rBCcwF3
Vddzs0qD17TG+CXmBIcAbFj5xh71/w59/C+j4/sRt33rTgxmbG7mSvYCr5VrxIF711iSpg8X3YK8
MuAgBwQr2QFb2DkWVVhE/Mmd5C/i1FMIvTu96UEx5f5o7/BgpKE0CamNsF7CZ862RcFTvJvtT1+w
8mTj1T952IMyPsvyRQ76wYmvvZqB5GYkKGMoIIB+ANMx+PJhYmIGraB8mFf0hw+Is7Ow/NUBzMNd
NNU6bKRXQJyEserNasLMjXxC3F6RCkT8dOHZeyDaCkA03UhctqKCi96bVDvnhhc047nJbU0lzFXH
Yr9ws3rlYXZ0U6TK6UsyKshihbjbwBIDBCB2bZPG9sLsMRlbRtpmqsuJ1VNAWnjZTCOJDfSVOai6
J+Wzs/DsWsd4UY4uHAvhxjJmwUPcLw6msaJ0OAWWKj4jEOWUGzEKbEquZVnZhXTd24Q+1UZ5xPHG
tSrkjmCtZT+aiJGPbReH7IyBTKH9BoDFbzrNWQRr1V7oOotXdNrWs28EGKllFlPaKZ64tX8+f0D7
1ES8fZDrKboxxM4p4tJf4UusMM9dkVYYOHde3U34ciLZ2HNe2nimnk7rRiCMIEnGYNG99Xb+ktSC
tZnM+sTZGmqQd6yHjYQ9Wic3V3Jp7SXbM+VgFdE+wCpXSd34bXZJN8tsWPhp60RFKcimWuXMI3Ly
avg1cdX9zgAvC2BE6pZeGphdUqHtPeo5D4FvtsdnzKGlOwdsagGJeEPmiXrJTs+5daHV9DQLRR8I
mdRnab8xVaen6dn0p6ZLoBexe1JlUqMRUw21e8hoVYVgp+SNrtBeZbtL1+Lz+RA+MUydFC0qnbjG
VcrDSgsvYAiz7Z2yeyEICPoFISUOIlLe342zoYDKj5l6PXEUNqGO09xHhOr67o20WFU/PEMtcsvc
WWOdcY46tKsJ+LIb6n3pdxFgj9uBGHf1WizljT85StWPfMPnxRJehLu/ai0whKd1CBx7GAtZSkG3
T27STimfhuzgOylnPh7FXHNyJYlubG21ulKxD97iAt/zNTh/UO92XSCFwNig2UN08zkBNtWFzVyp
6BX3+L4KN6fsV5JcU5UN6tlXN0o0SxCnxReYymLDhwZIVbLY6BfL6t1ezPRCBLi/eF5Zfy7VWKK7
7gOmXBCfQgnSIU5OEwM/uobG7RlzxLil9H3rWYzUwe85m8+mmZ2uPPSAmNxI7tu3NtUqP+GXNXzV
ANy7mYeqqUylVbpWv9tAqSsUtp0TDVuhYqJW2c7bY9PTY0BWWd5nEfZWfve3Z/E7TxX795dJXaHd
7ifKZM1w+q2JqI4rWntQsWtmNdc58tJQuLzKuARG1LzR2HcxwNMJ3YF+ipYEzOS8xSucRL3y9Ib6
Q7TT52FofTGbViojAw8MBfsvhqN8B9jK/o+SjjZZM4IfT4EkoUG7SblUyhViw2sTWZE8jrE+Ahkt
9lFL/U6mGuvwHeO9H6U6dUE2kTksb6CclHqBuOe9ISGaA3esdbC9XIYJp/7AFCHTUZ8mmGuA6MkE
RX+T6ukeaUz2d4JB5BhzNGmJvHjj/g6B2cAICC8yi/WjxYnHa/63uL1cA474VIGLl/3Xxp5R46XK
zKzGuZ+lQfaqD1hTgX8k3i1ksm+bK1lSTgq8FbN/J0eEFJbpl6OkF0yQKoRzl47m5FgpRvm/DNSu
y0Q16oacygNVjQDLfLdqRdLy3HO8TCdDcjirDJ+q8r9s0wauEYofmktJbvhzzTnZJxrxRsbwLfUD
HKlnBKJGL/iMAVnbbqMAYq5lzBzsjAJpsHazs1FoLfDLxShv/9x1lS1DvJ6rTXdf5g7D7rcFGGj1
PWgiML4VqZYp0PiVeM27gF6HsIKcmZCcQR/nKa0SzympnPRTkyZWoRTZrD89u09RQ1JFadEKJdSS
Y+8D1wxcuTsfoxGjc91lWMQLk6V8Cj+FK0zsPIiF9sikhKsdA0GtqnU4anU8x20R5xhjGsGSxWfE
GwBEP4gxzOVv5y7E5QthBV7EKQfYcmZpwpp2wndZNPo5In8yWZe2NPnyCDDKjLrxYqsoolwaJPdG
ERzBE1UeqsPzn3zLsXBAhZkzwtPP044B9nwy/mno8BRjZQngFEcgU3OLjQcpl0SMBMt9oeVHFVMz
kVR4UQXhnZMvWOo0U7+MXDQ+y5bgVtHTX35086QjGNz0ZePwDyqoEOh55a7eJSvxX0qjvgvrEhtd
QQLV8dfShPHys9Jz0L0bcRuv3b5Uough/g06SnKwlfImeFNLggnELKuLJdZzev2R63xeG9zYAW93
QxzEpvitIDMNMSCNqfur9XUmL4QpEg5GEYg/gzCUqH3rxFxJC1Fa+6IQ8z766mCWiBJ69S1cxsG0
LpnonuTcdZznE8ZXWyyKdRNKrnvUQQI1GHANPTnU0SnA/g9g1fXms9kya2mXi1NYjKGITg5dU8Pj
v1S8skYisX4J3T4b/6h9TCkUXsrZeFK7+fFRMNr13OlF95FGuw+GeaYBZAaxWKKWIdRK99F4Bi2j
iW6pyzZQQFYume1F/ZRnh5i7Um8NbSN6WO8znDzR5ezMJcG9Yr4QBnVtsJG1K9rO1aflQ5OCY9ir
wjY4/l7+bKNb/RDLguS5AlT0yRr6LWmCPZBZK6FDdwp/hdu319CFgMvrTisLgCHRcvhw5iVJu8iD
sTKDuEhpIMHy6d56mEulvDzAfxe/pVqz9uW4yi7+TAq6CoZ4ez/Wu4+oNiRk0OTrEHc5etut/iSX
xsiK1QXERTJNRK9Lw9RiIOceNlzBfh+bjSKGKKPTBdsTan22A21QKeZxAf5uqvcaQY5zaNikbrNp
gkd4oIGdwi4fEXu1QB2lhnobfsfzjyUX2rAyQC3dpyWhBLXmgxuqypw6B5OZwg+sL+LS+5NISBXG
jut8DzFURfo50eGZTslA0PJx7Hflp4ESSJEk4oB8OYohcrijvYAO4K3KS3jDjrOX3u9NboGoYg8q
ItgxqKFYAKQdbINpDegheCL4WMGrHxsLHlraOciTM1S7Mzvgs9DXOpz4yN8EgZ9JwaWP0bVYcmZv
1Gc7OUPx+zPiV6ZXmevfge5sLl0vgDUQhLbM1dMfdQhasM26wBcaGJ8Gc885Yg7CjaKCLqv2qkuw
eZioTofhBARNA3SlTY6FEOhF+6FyExxzTS/anY0b13XRthUlN3W6LU8EyI5vSOQ3z5uUEwaq/vTb
G10krnVYj7wBtKsg6hTeYcgVWskRCqIWwWAf7+ERqOpjmFgXjvLcafB4SApCM7Zx9dKKPPcfBR+c
sUyOnAZlMaDxLCfHSHJdIGKsX1Wg469SgJZXuno/9DaXdXlHnfYNcgDDDV6Bci/ttl0ZKHaN3q9O
woG3ev36l3iVGuculs4+FcAelyleu6fgug7qgk2Z8RHDqheB3Cil4ENhzB66LHuww2ZDl6YIv4hb
VrcbLFYRM6o8hsEIPY5vDspPyB9y0P+lblJYSWAZbtfvBsPGCWfXNv+q0rRyvwaWD7adTKShtkoD
uFGGBbIRekvQJg+xMj43vwglNmtkDcrsjDSc9bqJCZ4afL2cKnOv79yRfaLX7gXssKleOrH+SOwo
uFrZFzASe5Afn6Rpi7azQDLDDOni8BUhEyiAHYcr5NpAbWHAo4QsKfhV0S12gMYhmjPqfFdqTV8H
beG+g5bv8FXQSEn1KUGq1pESb43zXpG+Ax/DNmvM2ZVLhYkMFLJNcUovnD3KNTWqyA/PqPcNvS6g
PylCtm0JPQdYlKzX6qj+7Nl1Ap8GpcCOtKdqR5jXcBlozcJFNXztnDhzqC8kPu1fo8OZpcyOOpB4
y5xZbIoMQKY6FHHmeGYfm9NwVRCoMJvZBfrQofAkC/4Aya/RhB7lPaCZq1x/9E7kiwFKEVLzDKmI
RN4CMwAPzwqlM4aez+6v0ujMhZNL3tZgYYPhSrgpfTG4g6K+tv/XH7pHQ+FpSqLAunJ4eWWEnkjQ
g1yTHjWbjEFnLMObUJvtiQhPFDlVijOMmdh+DvrGOCjty2Io1oWSXtbyXzKlDUD1BPHQQKh0UcaD
MYy9kOTEeL+VXdSW1ctus3Rfwn4xnEZUzF8dCTmqMx8cnAIAnYPpznnXpPM7MWL3H+0LnoBYOVBs
Kh1CPCd4mOUhjM+sYh9JknMk317VXxUULjkvSxTcU1tXl3nZk9bfI+ls0wfLXlHVMZ4zCq2Clu6P
vEtdKEJD1FCSLJKeAPe97KWufF8q+j82ckwn5kCc1WBjhJ+wsQ/nHmZfvf1DVYNOOyg596Feep0d
resDn2cRPv/mkJi9k5Hts8xeGtVu3++SYVSPYHVOtkrDpLZydQgFgkVI4zUFviA+Ma3ne2ClV2C8
N8P1Lf2xbPOaarB6V3Xb2I4TvRxWvpFI6/OyyNWt6sAO1rs1XU6oDIY1sGQ3gSia5B/tcmxeR5o1
ivyIA/DOerpLkVexYd22QMV3UUubE2iFWQHOar66CdOwcSc1a1C5hSyeY8cWDAhlrChbgGFyM/OL
zno0abeXXeqrF2yGlxxvI+M5NOqH1OUTQijCCwzJ+6iSwzVU1i/UFzbOehc/6l/lv8US0Cjqm4lC
7BtPmj+Vcd6nnEUNHExUxCTk1ngy8s7sj9paxDCwvxM4sCyHMg6jMeDo2udNE6Vd79ZUYd2B335n
ULSubUXBm/yO0jk9VwR2axzkexkfsXU1n2a1JfshmqfnjcpxurnRBYs/b0a/iy0kUa8diXGkMLVz
zZ6cvWFtqQz7dvw50bN1KE+vlpM0AGvydzh22g1AXZCTbYrrmjjKT1Wb9BzUkoh0BFqbxmobAbXh
t9aujuRqUa9DHNEEbPC7atFeymF+U44kA1YyBzrkT9h3332uIiamPrnwqyKHfTHlkciosgkOTeg+
/HI7VZ4OBIEcW2WIvmBX1RKGn1FT7eLhK8sMGiI8PmxaE9Rcrkp1jPgqC59GrJQ6M5IGWZwcSSAJ
ESCBoDNnEd00al7IDtCzYj99JcCuAhn/nWlIx6MpRGSrK+3tBGSxvis8P9/+2gLnZlWu68xqCSoo
g9HdvxTXdvIZZpQNga8yYyZkaDoYy4k+kkOrYGmF3Wye2QkNWN052nK6f/6qs4fO6rQeTLsdLIKO
IB2BX39keaYxUGCyuSwDRM1FGuvYtQeVSuojDsCA1VzV/DiQKwK1AsT77GMPB7U0tVX34WQ+u2qp
O6gq67+4GF0Gg997z4TGp/SmamQhm3T+Qh+qIR00RLP5mVw08oU1BrebnrV32cMlum0rnP/5iggX
3P3kIcEDv+a3PXxdv3hsS+QJq3nMhxN1UDCbkyuIFCJkHHBv3+ex7BPgfE4J2ifThYI/zDWVjYDr
1hRSDBqRQmcTbcDzJ01ARhTw7KJ387YCiZkUPusCSK75FI3zDRpbLMwwxCiSgRQM6CSQRGdSwWXn
9E4IVnPVibmVqijxu/gqER4/9Z2PlXOnFXUtwkSnR2jIJuY9qO7ajdmK+GSZT08urFSOzng5kFBC
rt5puwj0QID0WG1L8HJ5yIWVMAzRbOvpw0/87k0VEVyuIsQihc5ggu7hTD9Herv6hKiGws13JBs6
R4C3/o40CiF/3tv41WjBZotehppfhRjv7ONWMMR8Z6tq9CvcPg9NcwxklFtyG3Dz+SkZkx2skR2v
hd/tCXXP5y7nCnmIvXkIFvOW9HViBY5G1OVvLGxH0YwSW5iYyD/q78Y30k3y4NB8Rxj/fmluHC6y
4PLQXvn+/rcsveiAtLwvVVsaofGv3eX5+cfMK1BkWafSpfYm5mv5Dalt7Bn0kph2sAr6GWzRo+kq
RAjNzf8ALNlABHlGD4DOOp8OMs1hOHoh1BSkjIX1lT/lptOJKeveGefDNIbP9zgpWQLspZJg+V6h
j2Kexo9jmbFvr9q+dWRF0kikZtzmN1JwN+5A0zOGdlFZ0t9j6OLu5SY3W6afi3ZUFWMe6S35bjdu
cnMbMaftX5yn66nP0aZUFmUfnMN6jQ3PjxYVLWWtC7yIbTHfePuPqzT3KZtqwo1OCr8IgqADIGFJ
os1bCcraMvkej+/C30hLBiCnd8tNryGcUkFMwb21vIuKc9PfnurwKnnZX5gBsHRHlWhrx9mJJRUG
4o1bjTRQIPI8afG5BZ1QpJrfJnRzZFCOoaHTzlBKUj/0V/01dF9ZrB3JPZV6JUVamd2/DoE1ZQkk
yr46qKYaaWZyfJfk7hgKQMcEDbp4Tlagrnn2uCynE+uMSqsNiyWmVmuUxCxqJtvchj6tmc2yHq+B
OcsdFkj41Tmn8A89mVRKqo0d6RFndHhsXorw9wGqWCQMNxDceao4dIoS1kQzEa/a4k8Q+3zoE1Qo
bUSrySsikGc0AT4Zyrf9D5wJCapo41Y6xzw/flCjMRbntcCp85ATSLMRasVLGQ92//i0KVl1gaH4
19l4cbHOjCtsk5xC54p1FnL2oM9fT2BNmh9L/++4veJccVGFVSRgIiUj2AADsPuJli4enZ1n1jnE
XV0Q9qT3omppjYPJ0HWxCax8Vv7KNo6zv0Jt+umL7gLXfAZukk0U52p3y+tQbfBonu1NyNGWYKpw
KuiaLwsNgKX0IjNlKPplADTiS5Bq5mfVEnlFJwDV126SAM91gkO0qEvGyQJrWp/JzrLfxoYln/z5
HJITNsr+So4GhH8I0TuMWr7XUKc9YJgQxjiAeH27ByrUrcVU4js0ntyqNo13Mti1BzN/dBLww3ID
Mgj6BieRDhAIcwNVTaR+dOH14w55DshY7OS2HpKcK6CbLvLOHRDGxICbFceH/bmPiHXkjlK62SRD
3MQbORfBbNDorydgn9kczPz6ABYyUkUwZNPFCLvB6PqkllUh2FUCCZFXvVkAcAoQEM9cSM+uEdA2
ptPcED/B6zDdnAD2nc7Sjn+9WuBbbHaBEMCDwp0DpYkiV8sf5buhRZXHQ9510PcQOv4B4MQBrRkj
RQ4pNRJKfh5Dsw3ijYmSd9XjGRerBWe1knjXzPKgr2vxM4xE62FgKG9yu9j9Di5al3+0+HoOoJd0
QLKiubsQonu2vrIdGSkOGsFk44rEDftpnsEYn2JKiBMKeghKEufNBa86bAnHC8KRHepYDesogGKv
j12epEYynFIx4dxJMq+56UACvLQXSZtuEqovmLcqL2Efon0cl3WngXCw5+mE4tWeIbwfp8zQ+WpR
bT5TmXtpDbLdP9Gfbfy3aAqsBitHxV7hW1DoBqvLxnjuPnONjjGGXCxEh+D364vhZ3exuTJAs6W5
8eeHY0DqZHqTrYRBh4vkNjw5vfpmA+n1nMyhOnV7+6xxEM6uxHgNmHqnLrbIzbsx383mgvS3NYec
5UKAoPL+Jy3UjtiSD0ZsM+OAN4UmorqtLoYW8KSmAse8mbCN1Q9FQ3FvSLqfvq6dLjixWXX/u2Fu
ptTuJ2k4erso5l8dTiUdwLU4zcaJcBvhFnC3O9LV65EZEwlV+mbfZL21hHBCot14fEqT4Uwnx9LB
OJTBLbel/KzLr1UnFtL9JXDZtMZc6Rbk9AkrAM/wrznHcGtzM42djxanXrbJKXvPO1SP6koCwrsD
UvY0ZscFNLXGWznC61DUFOboizKEjtaVc9KgYwDMWmIcJLtQ0QhyaXIfAfS2cG0NTyPfP0Sqyb7n
OC7fq71g33tikVTlqhdL6Lx9yrk6LgMURDKRu454W2ziW7aiFI/7bJ8WGzIvgavPRMeCQg5zbPIv
8dyVQD47BBOlPKS7vd2bb72f1UH+SQQ1+U1SclwER+/JqBB644SSoSW5cmLXLHK0qJ9k982f8DzW
muYY8gU2UCdMUoEUil6dyOSB4JJY7oUZe2e9AruqbeMabhQ9Olcwr6v23XF2IWWLhbbMXAPXUPI0
e5wlOJcnPlEVtrXzkoQAepnDgd8BhizVibmiEcHygX2RA2yybtaDF3RxR2O+Y+bTCTQd1UTfQHgq
YoXYqqAw5uTEAJykcapzBVhPz7YaJGE+8NDlkyCPjCeGDZw2L5E1lh6aR37apTWXPlmrLV4h8FKd
lNm0AbYYrgrTPSfkMIGvaxUQ0QKSTZnG92QM6jZt1pTYWp5QTm+nloHbVYOjW9bffXn0w1jbG691
f/imHSDeE2H7pHfj00Ciw1jyBtSpHePFySIeBkORmbUls++sfrZurI+14a8qayTWbDSIf+eSuqbB
FkklbnNdWQ6b4fqj3GU19jJ+QZ8OEIVLB6hGEz0iztNuFw5LBQKliKpx8IhKsqDMWnz1oYJMorSY
08sMjBrAJHlDcwppWvZHJWKa2tHB2TcnDTXj3wxvE1Vm5nb8yGBvxwsjZsc5CKk7GG5IhyV5rD2s
OK6kOGIESfIEkjOIcOJA4RZX3UD8pFrDVaeI29Ogu+qoSKUEXKpbo87U4aypmChi5BDEOzSm3cY2
as1ztZlMmHggzq2rFpu2mnUlgReF4JHa7hJ9REnxaZ6DrAL0o0H0ZY7MhPMZkLuroMeeMovrvhxp
Y8olysfW/bZc6RRPqZI3qlag0PrqFTi94J9befdeHgT70mwb/3h718qCNesvTyTMv+2CEtgFwDx3
1n947VMSUuBVE5xTyE5DK2rKIx5AzTL44qA8asosyBbJh30Z2yIp0Ymjeq+3KX6TzHNW5pezeYTh
fsuMk5Sbf5WCmIsDSrtpK17yHL7g+rz+tDZv/+j1cS/fuvIkZB3u5LUQP9zlCRYYTlObN6eC7U0r
qp3yk59iYNT3oXKXBx/YNSnxC/8nW5cg9g4XC8fqZoDUlQWGvTTasUFzxWnSmxJIepMRiAyPn42X
v80kIQFirIqdYOyc0E1IjHv1HCru/CVtWShQ3f/XKUPi5NcI2KDk1ZycsY4MF3dK5+Dh/lGqq1cH
ztrbFAW/4SE3bYgSvCQIumZZ8VX7t9jh5xyDiobi8Kr7CO/h40unQWn9LKE8PlB+qj0XHdVpnyS5
k6qJvcVUcl+IT2Zq6qz9uOlnCaAoNSFNgSd5e7McOsk5luHZVkiUAJ8Hdz1NMVCHqr27jQOwXyGD
3AinAP5ApZEcB0tEVVrkBR4Matq3dyBAF4CE9PNizI6KG5FD28AUswy5uu3MrYeSfcivDSBE7oqT
u6ECooNQxa7l2qzTAccfJ15Pgn6GhN4WTYOHZc5YLUvCsaFwT+Y0K4xzLfmP8KJc8ykChhrmjsiL
XyIfOap+tiHgZiBJKlvM/aW0xfPAarWulTi1Jvp7uAbr8jpLBk+/6BnwyqmbufF4S5ejTGnQy9mD
47OzVymBToIaAl+0r0dMav4iPz26TjAzjX8Q+8Up8laR57dgiNl5uTP2q6FY5cwfXbVXAq3ZxCDR
dgQtlrLORoveR6VtbIXr2hh/pkVet6yumo98oTDmK/04stIwTJApZr4rCdQPxuxKb2T1Qa+x1EEV
dxPe2q0wMzcGes9wmLZIvMxwPkXnnfp0KaOAzCBTf8RJhwwr1K3uTD/mLdwdvDPYOTdThWcihf3k
lGYI3sJ9iO6BPtNnOkQFdYem6YiuchkkpSmtAk6S9tTOpOC8P56KFrdsdcr0xDZlXyvx+J39w7zz
fAXShmLtqdDW9qBPEi5mP4sxdWshIucu3oz22AWX1t3mKxuIQjU5604yE4SyeGYVjuq7pjnwHUzq
5+FnJxAXQvQJX7nY0AowmsF0i4Kfbb/DwZLAQCay8aUWa/qxKDVnSlcX/RCkG/Klq/b6T/Zyus9v
fnKhFfJQVh6+2U+TeuB88gn0zg03dqJvuCZDl75vUloXZakWSZa4Bx91bw+1rvQQnU/WNFvV2tqH
mYXeDKr2RhZzgjZjopJeelx3XEy+Cis0G/eXAuHN5sU5pZaisxQAE58Sgxkp96TXiGg+6PDScF3q
vsb66jrEiH9Skz3banROAyq05JqFzLlsCDN0qyoraMyehuiUmaCcXJx6tt6A9PR6y5QxP4KviEZp
IkFUn+JcaAZpRRrI4gB470XZxjqLo+kbObu4Y3jyDbeQS5QAv12aWqpPff0HZ9rHOFt/sT7eBj1i
a6IFK95NZIELWEUU1ffpm/Z1Qtzx0Sy1gZ7j3wWKS6Yxtshd8OWRTq4UDidDZxw3HqbET6AkiPeG
EqIbQBRSlSCB3qJMWxxgb4ezqSOSqlKCDqcLBKQ0grgx9xhiEJUO+SPqUwowJLKKQb1Bno4yyCRs
jOlDaBYi3Dx0oGtk6WM3HPhZIaoY0ACwYMWeUj1WV6+Lp0OWjGR0swsd5tcnbC9QIit51Ud3u5UB
o7+MYxV0WNYbWw/D5vCczeTaWKBW/DSk9gLfMxYFA/HTdIZK4yk/MazdTjJaUrpepdN/FZcHEwkX
Rsdit+7udtMyMcIW6fHr9ns7m0VrcVMhx561JNGnQWQ2VUbR4YRTT5iKvKIiNbrJbQ1mg1CRll8l
ad2u9s95qFdHpkmWmVwlH9jDijtvNvllYDlsWoKa4CEddK14Jc2damn9bbF71mdGg1DZLgq2hs7y
ZrMirVhJf8khSTroWRK8EF2I2bqVZyUXJbPirw8ZETbVfUzxBk+n6r8ctqEVzk3miZssKwXb4Rkk
ZwXCulX5a9USkgliQMkMZdTYQhIaOzQ/ydLfvvylAG1qU2DMrS8rxKcBzQ5EOhDRgD8ZudXGad32
bAN9zHn9hp1h4gSPadpgjrKsKsb3ipYrr0jK7sbgZwLIdt6URsMM2mbrvhOzmhTAXdYNBMLbrN+N
Rh5tY/VyyXMQ82qLcIooXmRsT4DMDsK60eCVsj3bTiQmakOD4Zags3pQD7M1RlWWB+oe3tBurFaZ
0MCPGcm1/f2WzoZbM/Afv2+6pdxk9VmhthXHgZy1GdJoT4f5k1+1EheYRov9YQ4qGya9HYzGn/5i
E3yyzzjBn6MaU1j8AVr+16o1t1kLll5CuRZAr3Wz4sJipF68hmZH1rQPwZoopwv8SLUhN3t2Jb2j
bplqt6yD/m+2ecpafjoTSLPyvCOK/tlvfwg0Qg2vhEhkJkzXNT2GE8DZs8im+1WJZDD0t//Uw6Gy
xxEJRFXIHKmeIZZHjINjQwJhEySr4lyKUFvlDReR245p+Zp5ypNhKMgruG7kSyWyFQ2JoeJkbavY
MODHsuA0jnM8ZW1hi1cNoHVMOQTrk07CAd2NirqHbbKHjkHTj55fIKW7vuEYm3JH8iSoj8R7J1pI
IWoMS3czmKZtjVjsr57rPKf8AfDh+u/mS7R6HQ77DqPy2fzDmDXOLQc9PWTxsctYo5qlScHppf8q
jj9vDBWh03TP6PYjjgQHfMpyf80Y7sMENycf/qcZAqTvULUlvi08GcUMBCx1KlT0TIp/4w9huSQg
OKAxFLxegSGrhkwJH+z8Y/4gs8dzHvK+hh2ngDtvjB3470/eqjSAyZlkI/sOglSINlYaWDeGXkcV
brabiDHPrx8IOmKnU0R806XICZv9m0snuDmCx62voPBDwNL1jih2wJ0e2PfLWBTWU7PNmgOFQQHP
GYumJ2rN3d1WiGYf9VuichAFnQuoiBlK3UHdydxIc+F/UKrTd8HsecKuyuOuSa0kTC0x40+2v6pI
/6O7O+ad51+XnDODKN4RQauyuzoOQgxtxoJDW+5zS9ty0cZO9wELnYCtFps2TMgG3LNZI/w9D7wc
A/Ts7gt7rlQmPz2b6ztdWA1/1xEj1JbbvQiB0w1Dx7h2EmLaKWxKrBWjD/QqWi5Pcg2y9RRBugph
xDq6WdPt0NvjDjnvdCtuVsYC92wpFVrm5Agx6iN0QeFp8rcUAYyg05AbHkG12RpeslqqGRv16CZt
kmQa+u6LE0wRyvbHoWDWjlHewBFbxbKfIlXPfBM6nBbIBrNa/dEQemjAdVCrAsq7PsWf7mtZmlym
tr/fX4YdZlUtB5RUjJ8smX1FEz5EyXwG2wU2HRwIFLHBG8KblAMPfal/DoYD1jzzRW+K5VUfVCvJ
GV0W0QeqdL8zTaxgsfPfMGbqi3Ma89F8zMuZuwVp3JEgnws5dc6eva8BPNoGOfxkzjXbmHC2QgYr
73jRw1XUrCAZowHxo/4JGg2SSBOCknk3O89IW62sSqAJW0BhtDbewx1WKHr3rx9zQe1tEyxbO7IH
wwtSN7p46sLUsTjMoFyYGo/n6FvxVBTjtuqBZmviOtOzkA/lIUpc2PAwBBbG9U67tY2ELnUZuMvh
WuAgYPsMpJBdVqtTPsGvsgAz5NsxAfH6Np4Ffiv+Dw7wVqbhd8TwIfLikYbtEDHspO0VZGnpzFZR
jU0xFBYPTW28cx6SuzFEJRRKI3vS8LZIY+XWal3bL4WHq8Og4cpyYG24vLGRailyZZfq1nggN/Yy
HcIZIqvZWm7r68DLvumazuS7+iLRKoX7hbhHDXvCWKvOAy545mfhg0w/4lEBp1Mi5aZQ2EcE+ekU
fIaPi/gVYPeNXRRboOer7ihNzoDTGVaXQMLDGGtQlGnB0GyuvNHwnKXB4aY6uuqUZ6UhDMzcT38w
M0olD1ELV2HZncc1ClBVULVB2j8ZCENQFD02ttzcLFFcJBz838kldVdu9I0MxHsLxV4ST6lZvWqQ
GzG+bENcesJVPserrTKBe0/7iIxdovYaBMvujd4YHTmnyFfSreXcKM5JHSX+j4xkHCQm5lpOnkf0
ODF6ZRtLugW6Vx4GJS1/DRJ46ZyqBFlXrVovgCFx1JFG7SAwr5A5cHZhvwgLyoumL2XhpYUyZbDf
9CJelu7eki+Hj6pdyOtdrWYQ1qn+HDePyhgYrs8Li5xzYWVD2uvh8Ta24+1Tulf6e8Nho5HseXVH
D5/FkfLvoYVvvcbsyJE2L6lanamijbi2I0UHxfHjfO1Kt8qmKiOs1TuQ1OVTdRioIz+DVkulfS/C
CnG9wnr2ddGi8rawRy2TLtpzRjxtn/DunXO3hDKFWZF0AyR3lRn23BW+aG5sVpzfpTRax1SyTm+7
BjB+Krh14G8Bs1GMyjpwj8xFGS9/9xPF2ymQsOahoUmu0cSpUMzB5GeES9xb1EnVCSOEiumbsQUk
w/fT9QaVJAXOe84FdhwI9trxpp0YH2HXlZIV44/Iuydr45m0twrCahuUGID5lf59qKVU2Dlxloug
QsD7lpLTE08x9jWN7CmpykhjspfsOw/1Pqz2/fpLMIxTsiiMdv6S7JkvFkfHD/xwgyeCSUFrO2AC
Bkg+mr+YxgEN4o9aGPmJuuIr1T2jlBHS8YmVgVBiih2E/2jl/yLl0nCJJCIoOh54gP77CBXpSuWD
pdsYIJz/YdViNhdceqCf/+X+53cCRElqxGp4YNuIafX6g+1NusWYKt3FD4CBZHMfaBeSHogWj6oy
fDFxWcQ78eBJ18IupbDkcgHtZa26nnih6sLmNGZER5fNyqbFhI+KH9ltVXfPuMsI37xcYGtyCIpv
rJbFCHdppurPmdp3A4SRXAsVSD0rafolev9ToOI/43nchYpP6iRB3NfkTePt5nadQujzpIqVIWZI
aNXm6S/NpYe6Hy5CX4sBqxDhsKPHtXcM0VI7MbvzlZ3URd35wpLAOCcH/yYohpS1NYbmTBpDrIZr
ygy1HFwyygWOwE5ZEQ3ahIpv/NQ2jiTraPYD2NMKl1XSrSOg+ca3OtwBT3DaCMNyxxV0ouA/NXvX
xVDbFlSgbOY96VkfE1YhhMtsq+sUu56a5eIIYCaeJN/SiMe4YpN5iC9enMLZ+zLVEmGKeZqSkkVJ
W/iBijLbUFt6KwaEE65oXYII9tb66B+7qwWS0ri1vXR75IMbbiWRypFZzTEACpY9mZZd4MsNPq7f
TIwSmH4dALm1LDW9TWyZW1FAcNEubs4G8O9izhqCxDIgpW0KoddgaL90TRRTnXsmSv49O54sr/rU
5guX2B2MCEuibyBacg4ChLR+sOifgThyEa35kL7w/my+/HY/SDyc47EjLWRpM+GpQ/qNQk3IjTER
lMiaFoG1J4NLq6cprMCX9KQLH5av8TkkzMWzgC6IULCYd+96a2WQDEqQHiAtYHNWGfNiJ8M0X5HE
SLNBUjZ3g0kBIOjkKj0a+7kQgFQI8LOT2ALkfplf7WJ2MWPswiWyGgk9MNYtBMckVI2CtgQqyDSa
5sktJHOd7tyis6KFe6Ug06CwguiqqovSQuhhngV1WIF+/C93QEE6DwfaUghnY6m43C0nV4bLMR9K
9IsXG9PwZZvsDkRFuP8oCiNMHEsKnaXifNYXDWCDm36TqERU/S+39Bd/3h0pnV0jFUMXtNHo6L5T
f0tJf71Ojsw1+5fh2E1wWr+QFafWaanwsE0anwHO9ctABtq1QOVAr1zrG+DAulsUGnDT5CUOw7XL
KxH1dLWNVpgJudiFhjsNlbc47Aen3RkYaMXCQQsvdGWasJ4pXM7ZlqhndvN7NVXRYQRe9oUXdlE6
pPU3gClb7qGtftWoy/d2VVDwh/ekdRQc+pn4iFgakKYaLy1UPpcaXsGsfGpA+b8HkT0Tt038N50A
ZaXW12U4JtD5OZ8yiF5Qp+VwfH1ka1J4oCXXDLnHRdb3LjYpzL6jeaMLiwMf2pXcOhNqmMUfZv2B
76m3wUBD+Rv81ZINA7UWt48ccsIgkTk12Ys45IokCY4G/2hfinHK2B0I99Fc2gPfahbmY9yEJcuI
1Q3bA6xk4MjenLX74/tR6CIRbcWecSQ30tRLuo07yc4BvsX5yegLk8rEKb9O/NZtT84D+1R0F4eA
NZz+H40+tPmgohBsmeNC5HRlOqK3lEYlx4WuTcbNfx1FbfallA32/W2F/j5IzJY3cEOLsJauFoyH
6ACZ2rHRm4+URzLzdix5pTVIxpQOVQ9RvmYlIGb8pxcwpgd20V9dLcYi7g7v7nyR3zz904WosO4C
HCBP2fbEb544orTM2i0fnZDH6o/Zij5d5WRCopIy+h1zjS+CC+TmcEEy6WG4hklI3qJ7PGf6l06e
GtbMi7EBOBJ5LMPe88Lhl967GJA8FCNYWtr+7tCPohv3WeV0TSIc8yTxt1nkthmdGWlmblomvEuX
+o7XOMjmJZBi7ZSbp5TjPd8D192o19tFMFS45gIe38h45PlMHhx40luOxKuk1FOjePZWR1Zh3yAb
sztO9UVPRdonHTRKjjbZg4pWupCZiTxHdqTWseOM95Ubj+tVz+n9x8f5Yvcds4CXZyNyU1W/N0k+
J68VJmkcmxIyVy2vQMKHhFkomIWawm1s/DebIr/ejnn4rl8sP7jcy5oxNinVA+306ziuwq6AD7TJ
zgUPOb4Hn1lWqQB8d4HL2I3yVcadE9QeuBsnirO5hi5kWgxnu1sS47qFSirxhcn2ZZRVNq4PQsMf
2ABS10BmuTFRKQi1yriq6hBVXs035+soUA1rHvg3wbGjjjJaQ4KHdVQTr4czn7fsKT31COpqqFaE
IMPI2lqbY3lPYsjVt7lhD7skIMhI7uafqpY9GfgmGHyh34rpSftsKJqYrm5vSg7YyZ1sbCzXO1ph
DH6IGTpkjh9H5zL4uSxHdvzaJ5u0R94/fji+s1at/+gi1WxHU5P8hnNM88uhHZGqOlPa/b3tSDgw
x5juxAqRoynu4xhDrJD49F1yku87JT3iw6FN1+rYQbDPYoRBChC39FibUv2tCwYXsErJXOHykn1Q
sBhu16cAhCS+pPxZk6mVZz8iac7qHq4G+zwQ+tEIbG8XOqEDR8xRe70/iPpEAKRkL6qaICFQ98CP
JjPbks30uWWZX5qHwOe5mnYDYLBXnP7wDmacPkPeqMP9DOqRHTENjqPiM7x+ooXim0EzbVDEGaef
KFBa6RdX4r1T2fMJuqGSo6v1pZfCSFrxJyx8p6a7ipo0iIUdYXr7rDPUDL5zi2/puzNZHA7giFyv
lcc9tMWIYgf9PIong32pHGKnppr2u3MLCP4Lz5YlGa8Eu62Dei0nOLkwe1QLRLntl3Cs45dUAanE
1CrgnumolvQVW2e7THH7hBl1x7EpFWsiWsebjkC/3KFlmYLgKW8I9ff7e6D9rTdBVUMcRVQhdF+T
PNgPegQMPhxwOBIwxZLn5uuytEp0Xe7zneKiCbLeEGKv5QK+wq2JGr902afIn5rM+5reIktSABFJ
7XitHnjM9tcNGqivJxktV9RMVPgNoJEjfrUj7JpPMRBGOi3PIhXK+BwL5wVQ+TN9ntKZQ1loq4sy
LtTWTfo7Ub4Vyyxul0QCnS8Ym1AFTS1d0myBqvBQmdzMqM/RZoXgQRAYF2ITBH2TZtZ40Ktr7BgF
HwYbDRgict3/2Jlo/9yD72EE8LUcfIodJGoaPkv0uI79mVbRrkSpBe/7/Cxc2k7ybmXQastgB1L/
u3yeSGlQtPyWB9Gk174NYQD3o9ZJmfS1ifPe39KomWEeRlbMh/xOCbDUMZZHa2W1vOGhA47fSxE6
uoVETMmsEJWL10pU3psTkuUGxBPxfHsDjfjNoxmoJE4JlFpptxhG3vZoIqypBxKd4FRZOSg1qU/y
0QWz+z260v7C48eFztwfDduyx72j2FO8yhASNWpqZB97vPBbJmeE1HOYIyuJ6fuMw3ARCpHelB6Q
+sI6jkOe2n3BlofOHSaz4Ith3cBLKko2BCYLkIWM3pXgQVaQEWEigF5h9u4k5jcoJMf3tXER6XAO
VJ9d7fdZygRt3M63euCUQ3oNPvWCasWXISPMaFSVOMIxl9KUgXJTc2kwlYTVd2FMacEzWC1MS/TW
46LY9P17eeCsJEnqFE9ZbZRriHvuALVIPXed+hPSeCKehph8MvEzQbIHVIhzNNuuNWEWa5zv0/P7
nvYSm0E/13w85FZfSJR45u5NBC6J+mSfV2Dwdk3taKoV1F7E9PkJC+sVl/SZPckAGRJIOB2zR7bC
qjOwCGKHulPtGOEhmUlD26FdnCwIt4ie7pw6OhvbFMjROI1oQE65gLFn62VrbLnZH0cTvmBmF+AC
XwNapy/GjR+H/PWy8+uqDspw04JyZPX7v5KkFMjr/rsGymaTelmOUERYAEK4+ggIAx43DQX25YWW
ECh+Yhd6HgBcJE5bIMJZ1uBiPSWY79vEd8M9SLjqmPa9YNJzCbeyxOCxDG3DXRGuzTdsC7W8lT/S
oAsU6c86J9rA5jR2pd5FEMEJEMi/3bLnaRsut5XiCNK3d12QoZTSDu4AHbq8LWDcXF8T1bRwBxP3
inTZwsCW++hvI29FhVyCKcBbpXA9hJKlr+KIbOdMWJ/6of/9kz48YcoyTRpp0OBlzaJzuWTKSukS
cpeBwrey1C4f7zeQ0Yghy6DtTqEb06eMkdR3qtAagAVnwOumP00vVEKemeI1qOQBUuoHpwOM26ni
P9iqWuJPSNKWeqHy69c90Q5sOj3391Z2SkCVAxLdUd8BW4sCx2YPEUia53+qHw+ogNDt2EDFMWpF
oOTi2xcQiAJqIEFCsrC7yMHpKEiSFpydqZl48w4na1v1SaJeAI7i4qfFJXcsAqr7D4y+cB0PobQP
f0lJoFtewGM9ildDspccpj/uQAxhWpRESLR9C83NFBWTcmOF19qEaHd4AchRcN/bQ4ZNX9l5m18d
lGxCBfM5OLL6gtDot/aafMV/hFAYiT7WnZSp1qkitW6oWntpRWdjQ+k5ySSDIdR92oKjm0MCsa4Y
KSZRzqsFUJEsAYEloqvD2r5EgASoy8oFcFAD88RE9OpX0v9dNZvQXSF9kZof8jJ3aY96MGy79O/2
eW3p3QyR1Qy7VZ8LIlaVisbHQQUkPNmW/FcCp0Fxsqv/ADZuex0U/JhiE0P2UEs+OrNebzfbTfC9
3v3MQ0WPk413NCoB105S3PdM3o/kHraeUrNQp9eNJ7NNvtqSw3MStacbPpTCjjnONOR4Eg00AbbP
xNjJ4W0jnH3TcuF0yAxcfqk0Q6vsT68ks8gJc3ufPD4Y27rYouWuay6Qi0MOmY14h4ciEW9s27V9
z93QIf8qfwqSmJeIPPzpO8qMx4SzbMilrab8JiVnBB0R7/yfCVr88wumpWzluAwgbVd+GFCju48w
+GQ+rOHbuQsWAOZOg2WyC4y3lJ6rsbR7ptoa8QFw2CdubCPvcEFQZ3o/5ENHmXy+pkCCXhlQ6v6y
rDVN5905zAE/XefhDrlumakUJMFnbZoTNraBFp2K79fSA1j7bY31IFmEP1Yw8ZStAv3V016M97tt
LKWW8BPCB8C7kmlF3de7mDHCwYv0ItTk02ep3IzplWKmMUcpws+k8zuy7YX72Ltr94V92ktIOXdQ
jzT34782J5DEy7XzjGS/RfbqjrMqt8eCADwa63/w6dD1BXyDlGtv5s3abnZm8idbjM2gtXsObNYZ
S0zHdzDCj5nvhATTyGAlKHKxl1EQyXDTyizXs4aiAoAJsoaLwox8k5ln5PGhr9OS2MWunEu3XpyQ
pP++/OHd3JIOQT3p87Ni9c4CCL7BtEVLZT0E6pdmL8LYT54vIPIVGN5ENtreyjCJ/ZQNN/DP60y9
TLIbxa6jNGurD5EGf5UBU8feB/NZBS7ndU9AhiS6/eSWSyVZSCI3zoewGjCP03NoQyC2gitwDadX
oXpsR+Fi9NwjH5ztrt1QTrRe0VlukQ4O60kxcCrIDWFrBN/HUHJ6Xl3M1CLap/pHp9GIebjn/7Gy
XS9hTgMKgiGbgntSCDSDzC/1rpHD2BW9jsg8uCFzD/BStGIt6C49v9CnTgiqqDquacx03VzUrpkk
CZo9mMLaJqgZ6Wk09KMZNrMmbsfmB0tmZJpjpSfE5FDHHmqbbc5ZUoXs0wXmgbFeB6ZPwDdnz5TI
7wAmQLb8FCmORHg3apZzQpgmodlRsk7xM0JN7rIpIuv9c/Ttf0XhUKaSlKVd1Ht/RNot/ADnuFpy
wvSDtT908u/Z3+kDqms+nWmR9/RUrmlxg3692Rdi6Qk+1o84SBIbTTOzeztWMsTxvPxHKqn7gX4K
H7RdqYy1X2r3tBiLcTmWmfa12idr7hb5kIugI7lo+0xxcad5l3I4PlzgFs6Yma7krAWICIMwE/y9
05ne6sapSUOwxkBcTmpPPSEexm5itTmEx8I7G0F7GbSNZAo67HlNBVN4DJi/dJtotivGLVe4cbfQ
fUMxkwz8rerM/V6ffk2xD9AL7pszE0jfrkd8m8fUVuZFFZj+eBaf6yNkhOLVlxRyy9us61LGDCr/
7LORq02VWjTEOD5i6twkBhWmboADo36krfNVDflpN9Qk2ywRPG1/G/yepgr7BDnagcKmx4ZDNaNt
4C8CbM9NbjSS+I9gtb5dyOb6c1+DRAVmdUHUdZklCPjA45rpGH8D2ZBC7FW6C3e8JhF/u/lpeLBc
8y1fzPJitUogZdYWsnng/LpAEA3NT7SY13vBKViz2DcYxrfwQ5Xkp1c13ZlamX8ewbQaVOovi7US
KHVUgMkfRQQs4JEW0S/+md8xxCuEYLoAQxHd0fmsbq6iWbrzJ62IGVc9ePMqqffaPfFfO+CGwfOE
+/8tcJ+Fwpf/8+e87sw1Ub1f/C460jrD7LL/NXWrnZugp2jEDmf/MaQWlrkCMQQAo3rnRJY2ZOuK
8D1cBd+dXJTAcjt+zh15108OQLG/8bGvEqHizmmfWjelrWNbGQG3JrLw7+v9ZWMILZWxRSv1B6m9
bs3RLvYBecK9gj/pIn5TdMZmFMG4pXLqBErOX3L2EDaMP5a+y6/Xx+bWxTXQN90Q/o4Dr2oSeUTQ
5ATFoUXsvzJ6YPpPaiMWkNKI0OpRpVpGBOst3RxIkNaDw9XR5Iq62VOztA/uGyqCgpJVnm8by7j1
chK70OL2jvjQIYhodiFOSCgH9U3+rv8HO/3fmm1D2E8EhFWW6HNOrzr13KKCrWyHra4DiwFBRdxT
DQ3hKabrncxssviVWmqjWFHR8E7yb0dPB3KdasPMpzhL/oAkeEGmo13+9PjzTeldQOvJTSITOWXu
p8CjC8gmVC6YcBurftIXNK39+G7ZEzc7iMZr0EeK6gnb4hD2m9VdwjjsFJqOlK4wXEZ2aiVWAHWh
8QoiErtHv8Hh2E/XwJ8XozG85ty3jm7pocNlB+hEJ6cj1qQtTzSXf3Q1mzrj3hblRjlWuyWLVOL3
OAq2s0rIHsh/mePdNROkEGA/Kd9rFU+iUfNq8Gu2WIOnfVS82CrK5rLSfzuaMSmB7vfHC1+6ITOJ
2wo1SZB2XXni0lR3ukHw/xYw6iC6RuyhHwvdHuBKQ6xITrnQDVsyUTnlxn1p9lGPiPQ+FawidaqH
VXG5IRBn7WSXJUmVN/qqcjRmKtmHbNG+hcG3NqTA94ZuDPH+mW1JyuBcaiIPMpa3FIC9WkXsvCw/
32ZPIZbUI2SpxEWEYMKLDbFlySOyu/NgbnnS/kCHgIzqe2RkQIK4u25c2NmqEwv7Oz3KW4AmWkBd
jjBBV/eKlCGs+9Ry28glBg/ciPKSgoAx8aIk2sJIGP1VQR1udZI/q2MrcakAOwFpNOATy++xnhSA
djXeRI3qdXJOpcpNtlGci2X3BDIsHZ7HnsF/NAyie0JWSAW+3PENssmzvbaVTgIGByNRLwSXqyNK
rUf3PRI28nE5FxTq0XzLO/2yqkAonIlsh0cCRj5tUSDfvPd4csQ1ALIeZlKYSgvIg7qnPVWy7hYM
Jm3VIZLKEDiW1wrjLB27P24HemDnediSjcjJV5zFXq5ubeIXUK3/I+43Qh9B7KGwUUpHOdYwAlRh
5/eoKo/fh2BVUywlW9d3ukRTgmhGPQ0rfWYoGHxK/I9sNDorMKIChgRuH5CAqzfLxxvCoWT5lP/o
xcRHlkLEZsEDHChKv5QPy5lVHSLsQjnm5XfW9r9R09Ptxqs35kIFhHBo3TlRk/gsLWolmXEZpRQI
bXiU3nlJwxZTe4ncqT3VSGrImHgESH6k1WI75f1DRhbgmG8xJm3aYSjgvCcs/KqkFy9gKPF6NtSv
aK4PAj2xl4ofQzpftihJQbDHZ64Yqhhu2uVRRQpZT74yWUzxVfYuvhxEUGFtEP/JToxxN9SquVTR
pb6jzScAbdRcANo/DVm11XdFIB71QFB3mzFN0U1gaYNV+7IYsZAuL4LY/1e4OXIHnHikWI9o3Hvi
57+VVzgwrzHFHa9ewU8C13FjoN1mkqXNyvf3bgPH8/dB0ZtPKL5frUZJm/2hlUZokQCc0HNmi9MM
uI/uQ9/rYb+8tOn2sP6D8R9Cjd3w8+qJmH+n4z6Wz6mO+BjA6Cxub7nMDxgSa4MBB8oTDYQ6aEO/
i5chkUNNUePjvwbGwP4ORTwpv6kbnCcS2YDaEUDwxZAqthAo2UsvcRgd5bSGUhU10bBA/1/atlq7
sDN65m87/f8qOt6WGZBjNBfiBFbQCcJyjBTsdyxPcx9iHtZslHl3BT5Mm9dbpcQdSd05+qZqzkjD
VXfAwdy1jcYOXYJI5G44oSwKVXcD/kkUkKmGFtfS7enQ0PBEetsrUYdVAB9H87qugxyycRCWX2yM
Mvg+4p2FGTDhHSWpN7S6h+Y7aLFHXb1nUhkvSWZjUfS38TQTNlB/7AYWpcPD4IJg5jiem25qDAzc
dBvCW1hGlByuPPZwFI2JxcEaygd/mjaIm3Ng4W+Gown5MChj94pmtfhePDKaWvbCiXG5nJvSGJ2J
PQySkr4hTrf2bjyxjiz4x5HACreJaP+hzXKpXuOF/c535B/JAUeCjwUrJLuUkOQK71I/nMrrpUhE
o+82rsICGXZ5SXHisMDDGQKgnFGr/dvjHjQDfHTMUsW6Rwde37ljxWaz4uw8WQPcMfq856NdUG1y
rs5oSIJqWjrISVo5wd+RL8C727U9L/qjCPJ2X556ZTvA36fzKoINsqhvDd/UGrlWxZd1f+crvhUp
B0wC8gLwnjGRSIrxphp3NsLFgCniJ0QQHwHqu1So5nLVajItuqhGe9i4T1JoJt4SCs48s5nauzxm
aJp9vHK//P9eECyxnVE/QqI14B7shsSX8LZVdceQgfOnkuNqFgXrJHKUwUjhzux5z9c6Ns5R4exA
TBl5VwEZm1hrQN5GjcIJnsDOxeI3/Q1Lh5O0eqm6Plmr0WvmbvhHkJ7Suo2TMWriYjz8fFhi8/q6
BtYwPrHdVm+yJPZXeeLEC88toaPcdE1sR9stYgrurK9kLkqilINZwtPfaiSAQi/BURVZkN6ev5Lb
Wok3ErSKweZcxZvbLqAzVnefQHoziuSpopmUhn7ShyX8KCuvFHXZDz8aGgPRKGBaWSS4zjTLyaNp
XToycAmhS9AcyE0aM+s6caiDqGohrGIzFkpddxz/f0uhlcw4RyM5vOCYB1oP1ti5YRd3alnJx3T9
sBzaj42E7Fxv1UIS4gQLM+OaV5tWsIUfVrSnhRAKlQC9U58J7Pr4CIO2+/RYEEcNzooZKLkS0Emr
YvOJEqkOsyKmvCNTvQjZU2U2BJdl7CMac59VdxC/v/KL+3OTTZgD+bitN5y+3QlNuw/M32gsljM2
3DIIQcUdeKmpY1+SpRHNCJMZXEeRa16qQ/tchg7xSLGi67ua4rGeF16RoJTQ08BgEtVizOGk1hpF
7znxHKN1Mpo5ZLucFX53HilT/De2SDyh+55SorDQKFvTqMQR/zPjDTj1b77SVpnN1qDq8Zvw0nR0
ddP4jZzNbstkUeL+7GP5FtFcix5F7xPbdpY+D+OxV+ekncVuLgVltnUFM2YvIgxPBK2IzOucU8EM
YpbLq0d/vu3AHXNMwpfOft8j8hrkFZgDCgSP1uQgSfDlwRs4CzdjETcllfMevdSKpC3bXlY52ysq
NzCm8ldONA9uZ+zOGc9aHnOvdCOnN+W2j6kR0lOjDq3vVtrjE9Qr09OqG6wjJ8chYAOmV4gWtwuy
heSRCFOSBtML/w7bdaLN5ib5UJNvfJFC5j9TUWucNdKlQrL9OD+i9jEe7zpyrqiUwIuRS2Bi7lV3
OMpqbULoX4gpj/R93UYq4Gi1iIMY1xoC2jTV7ST1X2jKtwdv3OnvXRqNtEsFWIAU9evMhqqEwZKP
UQe/qYKIymzZ+5lhNdwys/DtBh/4cMKOvPGoaoeZLcvnavAFoaQTh2YmpFDLQy35MybVaGrOy3sa
bzZlSvtxkV3Drgr+JrRFhag9QsdJGtLdNmBKPvxbXISYpzExy+2UD+tqLvq67hTW4pvl6Z+P8wGJ
hQsBa0OSFTWZN7XYY8a5AcgeCfxPr95CksXrTMbecKOpmDCUrgtwLKZyfiuL09r1AFRTNB6YEzRL
EI5RjNWIGnm2NbtZ1XqHf+jW5Q802jUh2fB31SVzu2VyfnE4HjWlj0zWbNsF1gQxw0Vx0TSBBr0g
eEd9du99C47mVkPbTke7FL7WV9dnhTAUtXWA97kfQqPSdmgBQZcyZFY4CX6CftD8dqJhOyJxYQQx
ApqXC7Nq+CuxBAfhX/FiBHG0LJHwiOxNEqva0k/zaRd3OxGyDKFGGXOQApyBHbPwL/h+abrk4OYA
dFOJQwx/321xgiHeI5innLz7++ulVitBhvKZns2hFM1LfMDkt5vHNVc3BcPVY4Qqt4bNwFqba7A2
LiEkhFYPIOdHgIPzR6y1dplsBjnt2jeFNCzdCYUPmjUC8d+VvDxmWHxzubAlQK6MFqZqwXj89D9n
fzWIrA4v5W5Z/xHeaZuNLbkCItg564y8j6oL7wMT+RW/tpxYYfFLba4vyvQ26X56j26VwnfmHCcM
7kaPpHu7kOQRWcxtNwA9pcz2OrAwgFUzuBpVwQKch3nUhS1iGoXkiLX/iTiB6DtcKvee16YfcZF1
iP7d1n/z9FA1VjxwcuupI9boNp5eQKDgDoXqF5O8q3nHVmS8rttM1H/RaDnIff0ISWoeu7YM4YM1
D+m9s4SxSZA9e2ZAMJvF27ocYX4zPNxP0NIPr2kSxThuFOAy35+bnfCf6Gd2sJyUMXM2oEJQmACH
o8fAQkT+35X2Uwxp9n7ZzHLtimKEYQjpWgzcd3FoVt1iyCWWzXbio1g32NIY9qZ8yPrYctBi7hS4
Y5fZtcdKrSsFGiWQLHrqLD1KxZxw8X+tpu/qMUO0zW8OcXFNIKbxYRS54MnyWlyEK2H9q5ZQmlpi
bv00Cz3St5wOUr7S0dKMmL0pvMGL3llO5jCA5R92Cmz0+8VbPZfNAVhW68V21fhSrHQCfHrXmMPc
jm01rSoS4RiH6EYrhpILlIwM3tkjQJKL/E97dL+TLQYbZpuz+mdlLmNhukCZ/rbfD1/JUrzi1fQY
pvXnF0zg5NW7m4p+vypoJpsoFC6R7lHRkMEhbD23hFeNRGZPR3PxK+i8eI5WB4RKzA8JYpggjB/m
vpg3FkHGVStOG3C2plyPtJQ/mQ0evOd66wloub6Y0pnIPcRWB+1niKynVwHcvJNg1dydZTUfpCpb
RWGg90JmG1TeLonhuhnHI4n/F8f/LUtXOYu69UFST/GnPMfrekAkn4PrRKuQH3WlC5Tflflrru7t
xyGqfWUWoZCdjT0nx/lTe41hXhDJxOMaJHWluTI1JyBu0+ffvwjtEr5MHuhIjirvAxd5OEfcZdj+
djFzv3PujonjKB8Prtfkq+/c9ldTQpDqWorDCG+cczBHSkAAgN1Zo6DvMy5fBUFQ1SYgtypNjspA
IFXeLctBLZC13zEKnlKiqUu1xYvTmxnuvecXw23sj0K1v711ubH8KKqvFjxiJeQU9i4j55z6Cor9
F3Mlg9gWNMAPisXYAajKbxuEb0BYCp5GkqigcwDye48SkizCiM2+Ce5LsIRW4Xqf8kdSpiE/Lvf8
TLOcfeD2v58pSTO9hxmk3eKlpr9dyDCJ0vhF0E0Evo+VNcCY1k6i9ZGnGtdceL9X5ZVXITErjj7S
VKS2BFFsFZ8Wz0MNQyn7CshaxQ7mK30RxrYIaUcA5rxHyOqg72XeKGun8ybqTih/6eJLaQsrAimj
hm0NDfni2oCAMKnwvwTFD5CTcl/m+Putqm6lzqJlB2HYX99iROWMeFTo+HAxKAhlI6ZQPwunmnSN
nShvLLhm22WBgRruTf+VOTwUEc/yBMinOiIACTPrYsXOAhiUZeUDhvtpp+wRR19Syz5QVLlPSFkt
JyHauPVbbmySd6cQ9k59vHZNTtFMc4xWlYiVWlw+UgbHd5c4Hc/3dlTS2erFYO9ouX+91VYtcF43
2ABjZnUq39dd7AMgVaCKvFyNERP3Up/R1PCFTO9E3wvey72p9hoWTFc1bDCDGMIIY5mbATHApyf0
+vG41EA9/mRaj5zJfwkOosN22U2W4zDFrSrq3pZUaZ1YTBvdsGULQPfrvXd/08xl7NFUOu6CPPRi
HsoJoEeJ8rImMQ3wojSg797pi/PkqYfsCEgOAP3bdYrXKHSzXX6gb9ZJXZ5zyFC+EPgI4HV/hVsH
zHCQKLaFZX34R6RdXKl7WYTwUGpeexZFY4ycoK0dNBKBmnP3iSyNyo2XOEGiKEyHz3xyFKwEJWy4
dqTptukrgahjuhgcobhhg9rcQKDfw+gfiq5EBcV7mMYaAIm23qk3/paPCf8lRSzT4Ixy6hr4JP0E
JPHLUBU8LOdqAHznUE3idV3ynsHoh/1PYyFtfTB7AnCccE2DuS8wBuiVCZ57cYPOyyM4epEpVO7t
Cs9a0GIDCf8PNMUHWhXfTLqdSrwo23DEwpwfd90boHJX5LpsgH1Au2lv6Iwjbetm/7WoABT6o0ES
I7u802C3PBCPY3OVseHz/1d3kiWeKPibFcRd1JJ3KhP8Jyzsxi2fTYYt3w8OF87j9lFw8uoTmHlj
QfzZx42BnqpaXrdInxTz6EIEXrR7xHgEeLegcqt4DMioY9zodXe+CCrJK+UL0IPZrG8U0ROfydet
dHufH7NIJDjQxscWIH95JbpaCSuU2Pbm6a9c/ca6gGgFafoboGEKdSnMPifZm+HcHOXibPgeahis
D4Cyt3EHJ1rcOp1UvJ7M7sMZU/DmaYAEZp5fWEMfFlyvEDM0GD3GFEc6avnJKGkCC+fcsZNKjGHX
OzvvUP6fxkAH04K+90WKm4/Ui/1wjzfKk2kDSNLcgTb3u8JUXByyF8S+uQAybWnWFEzACTQe2gRR
Oz3pOrdTJcuWAA4iqfqNtdrubfnbroK7VpAl8i8fd4ewrqtvJVWYa5fk4BCq4NaQ152pHAocoR9+
RWjfuohE//nr7s9uWs6jWwWDndaoV7InhaaoJSBuBYYowFMyOB9LxILQCSDlIDwAo338jVTAg8S8
ZUii7H7PQGKqcvPmnjfYKEUYQJL1Fc5e2pgN6U5IwvBY6sCtqeXHTTEBaJ1IrtvaiMTTVAunNlO2
AQl3/0dni1Iyawz471qJih4fiuRCUFazA/MFZan0lM64DzkhI/RPk85Y5iH01S2P2kLCTEdDFaZh
PB99QQUcMPd/K0HtmSGgAc6IP8UqmPCSWF4AX/PC3C2klLJgbHRzfCvtFsw8fjGb3VTratbcdIPn
Kf30k+LWOx+KjcOiUJ34tA4j1wPck72xQyNcl+yEu4eJgOUpix0rBgUtpihBraUCddmkjiKnUyMp
S58unak4WT7QJl8WZPr7g/zQ8HWUZxLNBQx8l12Mpy3h9GLGIZs1CdqRDZw9IwBoteb9Zs1J1fUA
Ne9N/QTfkB6avQFLC299Tjvie9rA1dqMYOrOcqrORaRvAthTM9CVdsROQ1ozQNPwMpmPupjBDiLQ
lBIZvZmG5iB6lqPRMrlBEAcNFSdvsHmgWmXuro0RNixPIasjqmV4fV2OHvJdYyRevZwz7l8t2U0X
UlytoqrlaNs6vfkfTvZx7q2SCyJH8HKxSTajPE0gtTuIjph1quBJ0SnWpKDWYSqOJDdZqYFl3oRb
Wi2oJ9kBBsWGuqPRIi/RMwlyxD4PH2LG/NdM0Lwi0BLH2x9MS3Wed+fiF1mnBCwvctbrMJ3q3QtS
eTRLsNB+PMEFQKtluLB9B9Bgeteqp43eYfoRuCJMcWinCLJfA+ib96I6Ps4D88IqoguEJuG7z95j
nRaEgAxRfh6bsVHFV0x9LlWykuWtshFVD8MJGvclGqAyV6/8sGMU4gsg7hTDfecuz5+JhXcotYVv
AXxFvX5f96tbtSN3jZlRlp7RO6/STpssRfWBs/ENqPznRv2fBTllooV5Dupd2vSAVhDxNF0Su/hs
FpCnvFvoZO8w+XJB9DJCErsXWzmOkWzGd65wFqLRwhvXaYf7Tx5nqkHSz4bA1WQtgv2sTrBeu/ry
44k5Wt28heD12YiGslnR9nkreHYKgayINSLVqjnb06AbzG1B5T+PiG+ZDb6u6ThjhKN8G+X6MCRo
BRLnNlWj0c34BKtHnNPNKFMexrce+z8J2/IOtL8yNDTHG6zyQgIML2E1/fVQOPzrjjQuKGTUS9x4
PzXayBg7HUFWoJhNKuWfKHG+gW/lYgBvpvxsb6cFLzwS7VnfWbe1o6fKfJlEjBytkWlNhquMflSq
m7HPFk/G5Jr1eA13BZjQfcdygHR9a1qa+TkCwh5iZ4NDjlhzCH1bWFy6p+fWOjtSEkPgbZiPMEwr
V2XAzEpZhQSc5kwXg0HLHienJnmAEBcYsz+HZDVVwcnUxLBeI4OBWHOSTFPOJgdUo7QgmlFpVKUW
JJSKSS1xom09oDdBVXKr0U5pewcZQLkixS21Zh8ObPgEUYWp7RbV+pBe72aBr8WS9/aPnEeZG9Hh
1RpQBpibNG+2M4VkU0hrIKOKYg+NOrxXRMF0rk1V/0WJ7XRn3BZ8qS6Gz9NKGqlPQhNoME8IRi9z
iPIIin4TeeuydxtvO+Y5OKSoi+2KBHTI4W789IzazDt8ihcTBrw+dORyr6zgZ1xyEyNrp/ooNB9I
KwWkVXN7GA1aseXZ5hpIfGY668UMIyu1Fs2sWNdS3yAsJeSXczknTBEfK419iDZbBdTW58CbZHfZ
KbW9Grt5EpUewsNiS2XvPnyi5WxZIJB3QWMIxVsHRUa2/hJqSluTFP7S330SO8AAQMLv3i4idfYH
Um/m/XbgCmm68rr0XlJd8eg2Eq+Upcmf5kCMiCIlESWLPu4Mnvm4V5f3LF1ibiGcM26MLDryNZri
tqx3W+MOKqomquoOgYkn7jVvswtL0N2OeIWxaR54jZDr1euxdvemHC5DUNXySy9PdkFs7G+0OqKa
XK3fFrF9er6aW/I+ryVqhhtUuJrHBNmxUdkytvkxDzSFLE1QLfQa0gf/j/2XQN8C0OqbgljO9u1m
PwI4O0XbS0Swhaas6bshoZBsalzTMf0yfhXgM+KLVUwLvcE/z19iwlC75q8n1f7z8MvB0WsvnLEv
HXeW12jrgea7HHo0pzMVVvvqmqN2NfOofNGWGOx1i82gYKd3SGWAE/plwLJpUIiWncJeTXgCFqm2
YoO0+zd9aySvrBMOW18CALrVfIjOFUOeDo0WO61ukfzZwaK01mD/3H3a3PfhD6pJxLrQk42GKPAv
FvZac97caGipagzcTtOS/V+bLpaqflW+r77TSovxhgfp58SnXDTKn4vyAqnFU70v12Sl0HDqlsE4
xqRIMg2PfBGt+VBSZjvsARn62uUKqpNya2pRRFPYj6Dt55jonF9gu0vWeVoh4yGN4+Y9FJwWjcC6
uS23Yf21376ug+r654QSel1WcHGrCbUL+NotD49UtyfmsdG5dfYFX5P3wlZasXnlw4P/EECAXkGO
TbyKxfNq5D+65xK+Eu+sJBzNvkC8CulSvIHvzNt1Zkyx71VaYVrQ0xEeyVuKUmSMgsl64IUmgznt
NX8xEOMzB6xX3l1lR12le4X25k/RNCkLGxzMAUjW1UNZ99OVh9Qfo6YJktRKcKp5FpM9qDCAhcrh
Z6loN9Pqc46KqZH02DYQH+Zep0sHGYivFfe1YNCUPbAXn4LuEOgwSKcgPsNbyf4TdP8uheeO666w
AYclbhyRw4/hkeOK8iyWhVj0YeJwpPqsytTg5e7ZvNiRtYjY2j8V39PJfprfKq0MEgVxG9cnvNHh
Su9JOGp44/o0VC1mTwdLGbboPAXh1n+NmZXNGCj3xDJmP5daL3HZZ9hN4h5H1AXlSgExW9LOF9c6
F9060Sgmws/HS8Anx2G0nVzJilYXgk+siCfAOF/9cOB/JkEohOdQQ+r9vUSFrtmMRTx1j9xgNub4
Sr6fwFN5l/Om2irccLo/zAUCPzrOLMbpqWLfoOAPVhnOJiM/JQSD//5tcCAHQcrvF0pHtZ1OZ8PX
ALG0uPjL5YgeZHPLFPs4fMLjiEb2/CYioOh/7m8JkvHiL53gkdDbBxAcL/txkZXZ+/pKLOq/g50A
0RkzfIPSo2XLJEQpSeqW8iSjBffQcRd70tR94z3fvdbZI7uFvP7++WuHxG8QM+Rtm6bcMEAf5P58
QcKx+XPvbYALM6MZkXiie9ojsgsH63MEmJVy+rCT4wrjETVmrNibV0831ZK1WgP/RHLNxgPe0hhX
ads5/1scE9Zk4738iR5/GqduDNjfI2asS4BoZbmp//g2bhJgncQVCbk03aInTCJ8xHhBSbk7bel7
zrnRnUJr82SPV9Bg5yvi58gi4/pI6cgGaL0QB8VdYabgX/fbPad8jzX36H0mDOakgBYUfh8PIym6
qzuLiWHyT5mNzBj4jOXBFRK2YN/hEjRn02JJlewBFOm5WMBA9CAqXMRBcD3Je5SYzITnUkMFB8IR
uXYGPpwxtyKCTkmnFoke71d0FKIRnv7uFImcpiMkkQ3SRwLCw8rS+HoXDYiOSRt41DANaHOTxnm/
SXDlfpLQ1sP8zP6VeJ9BT5ElX6sbEjb6wAYFPJ/hhHP6OaaEk1VUC+mGav0BpyeCcH5L0abTHTWf
5GLDUFMml2FcqtnNnuyX+VtWmSaoQSswKqzl1cW7uNzUQzkOb8t6aGbOD0FPeOybKp1c83fBOD0M
96YU3XotQZUcu71I8MHyIq5PvhdenEtOCd/MqzfTFAH/zPQMpdFIf8oFDSz/UQlb+VbOwQIamKTl
8CpYpRvCZdBor0FIOddnKaxwvNx3Fi0LGkbgr5EQMChWqmcJ8ByXMsFEdfFNv54I2mz9MPh0OnV1
WJLmSpqmjVPKRPKCUIhNj/CT349j6NB2Xo4WncPoUSCbBEw2Dvvzhh+zNnVcsSP0Q16aDYf87Dj/
8e9xodMcXxIrYosbtnpgQJ0H0F2nXzVqNbExjgR7ifZDzvRZUD1IrV0etFpSEj1L7JojeLGfISB/
T4JfmCn/d/E4+F+mFfjYyGb2XGK0CLnI3aduDXQUa2ywT5F4en9E/cGw8aFr9Fk953Uf4+B3uBjG
ctdCjAx/a6c2GnnsU1PkTZ+YZxMa8Ik3BQq5NJhOcDGRWSGgENCFDzKjh4YnUgeNWutvVJARbJon
6egdX/QLfzMo089tqT+aNHPzN8gnLAThdfELw8cUsUHndYMSZLuCCBv2FeOygxWI5K17IdsGr7gn
hnOTj5y/LYxRIrUDAf/njRhHssKNoZPr9qKyhYwZXeQ0iU62Zq6K+B61FVDqSRntzPc6LiU912/j
F3rNyQMRKeFjliFhu0bIZvsm1LZhWIaMQ4nATqJuhazKKtrH+6ncgdgoe20UWtKtMVE4q+ywyvcz
U+Aa9Ufe9pNbkXslnZK4fhc+By/jZYoMzfZ1AWgE/UpYFVnI3gZYdd875hDmhy1JBV54vQ5WZtRL
upFkxyVZ6u1zjhAYh4NURSHs8DbKDa9qQM3jTO5GcQEAlRVyPxqyqdj5ppKeUpE7LUAY+UfNUCEb
ons3SYoxd4xMmDczmQs23ynviJExW8MdODg4s40yBzzV11Cz0wQWKewowSthyU+xUPwoSEwvg5Ed
XukrmYju+umSRy+BeuUfPN4N9Zj2yA9snISbmFbo2KpFv/KwXoes1uYrEVMP6viu/b/ljdyz+ECZ
PAOZAJ0QmcRC3iz5SNT6xR3xbi2tvup4RRk3mYsMIk45NtabqZFNQZryIrpiZOHABEdTvkbAxvAg
PjrnxO+v1NeD2zoNXGwD1bodEUAHtc43gvcQqNB/gjP/l5A0ugkgzZBeu8GuGSVEO+Q35lwTyIpy
bBlQz0qs4dDH5ZtoK3de8h4sY/dlgCKaGXN6Vp71ionDUX44NPWLc5kyV3B0cYLSqNRceJOYkPVe
Pe7StYOFJ4ErXcEtt2aDd4zL9QTOBQTLI8SBN3dlexOn0FKtN9htX5o+xxQ8uTz/h6RXd9nVpQ4D
vIwoKrnl8gOIkFTFJxNKbHP1s9qkumdUGnbGi1NMvzrJwUVvtZFwjlSqYrV1woRmk4xXjCcUK4mb
fdmUic+DDEnEU02M1Nn8Sy4Au0zSwP5/FFd/2FZfz5VIECPGubI3R2En+XoAm2L4rlblVK37cpvU
Xf2UILJbux4OVayn3Mym347eqWujCWFgP3RhNDsHm9Z3XM7XW3w0iYkIWOsT+U+BzJuFSDjpnJ3T
Sz7dODSweLZuxxu4FYcSqUiuCDMQZprcJky5OBl3H+lXkGUBbcvpZktA9FMonRehpCUhvdZpSaN4
up5gM/moB94ijkEgWybwYfO34mss4OAhwsShjQVzVt7rmeQgivCAXMGbNtaq4TcCroLArGqVMXoG
HC/6EAsq7G5nin5VAOvfmijPt/nT4L8epBcibWa/ZlKXoXUK15M99qYGwn54TjsP3tKD0rEHKH3f
JzHJCR6H97+Fqp7RhortQlkBPvPqYlAH7VaPdaE/7M6el74kBqPMMKkwg1pPCQ785cDgHTko5XBO
tvDjdQeKaaymhsrtToX9MT2t9y/MzWHz1PZ9bmfr+54wySxrCXb7976QWw6RUE7YWp4TcIFIbEEZ
sDyS+LqBDLssvju+bXcehJE1qh+iq/05IOU4zGp5YtoByVZDUD3Lx5YXhHUrVLeTDnqeBZeTNAOx
KWGwv+92opGUBfTr1sEVqsLx/f12lZj++O4gNjleosxHWuLwsrhdPisvwSiha8rBbLdpn6x0abtq
aA93A+GnZ50SxBeJUmRV4ZZHMUiAmmSP2JTcjSGCtDxbRYTpGLX+ymE7LFc8eTVPDX3URPwr3F4O
7wkfssuh4otqnIBnv7oRuFTKf9fMFosALR4NVNTNHRSxsCACdnlvhu/Z58IuQ0ahPupTPSQ3T5Or
SYiLWT+i4ljXx5juHfYuJJQFKgetR4gHOYZerpB3IHUjbFp0wjO6ejKfaGEIRcclnmYhqFLqGmiK
RNUYHCkJ3MWaAMjvbnSDBP9tv1uonYb8HFcMkIptOEWUt67+OFIgh42XxyIV2EYYUODKgfAamvmf
qg0nWPVPeJnP9g0HurktSvhGR7aMctOSMFsoDCpDXEmnhZskr2HhzUbrRnVhfTQVkZAXXCKleEqK
+JbaT4PPhsML9ZuaPxaQi3K2G+xHTyz3uUgvJfnxckYHIEE4i5z6m+mVhu9CM3lZhLdrTJhjNTb2
78q3ODmHeYaooX+cPTsG002O9lGU+OOrqlixpUQkyDEUTTr0K79YMNtCG+do3ie0aqA1Nyi3Ernt
jj6l37Mg6a+Jer/9cLGb9+6jRX3CXCb3Hos2A/MvZl/SwxmAnFQKzoUrD+IhERYibfqPl1fe49MQ
W1Iaj/oEh67uCs34H66O0hzd0gepWzUFSPSxTVrQPZUAjxUpHchkdLsFRGobgjoF/BLvZXPYPfD8
EDmlvriaJVlHnCb1g/+PfVl5gphpQdqI/p1/IIUnXSDfesQMnW5IgInkEhR9KgHqIage3gn8RwZh
T275AnK5zGzmjRKAmfSrvTlOh5RHhbkk4QcLHSTUOYF9DF6LY4M740m2DbJbHcFi21FSNqEB1lhc
FNhF4pgTxAu3krNrFBzw7/spBl2ezG3hF8n9vVQgtWT507PBKMoD/SCT/WChm+K520pk5di2kIM6
3A1tkiUe9oEChQtkIJ4BMRljHWLnJ2Wws65y5QVoBYmHsbB24bgbVHjl1MJJ8ofyuByE9B8N8UVb
cxQ8Sp1RF8C8HNOZQyAsMbWGdxWtPiMqQJSRAsxP8CLhWsq6zLX1/HJdmRWa+GmtvSk0mYVNFSJj
lTVZf0v64t57reKGEbqwqG0Th0IrVtJfvJFdGeX5O2tJAAf0AOgyTyHKmoQBOgfkmN8gkVr/N5Hj
/HXEdnzWKNo+xeZ+Ln+BF9MmSy5dDKiRKuzSBvotAEGoyE1m8AbhU6wbfRoWh8TJE9kF59cykWA/
cFgEWFmzh7bS8GiNzyxJvYizUpwhfrhKu1EcWo8tK5wOjQSGR6XbpWKlRY9Qn/KnXi20VOTZ8TU4
8WDcmNgZrxJCKYExH6k+YiPwEKsMFME+AztIXfuljOjUm7KiUTt+DGLm60vAkCfsh2dC8rONtzWK
d8mcJw/DebTl4N9BFYqIENd1WJVPoe3NQnx25SbezlowM/R9+961aOFm8NYsGqQuzUhmF5BlIhuj
hoVTU89ukTBYvdqlDJCR6azLqqqBxVS4YxiDx0cfwipmOxJIrkOfmlVvC9ZV63JvCsiywyOBOiBM
q9f+bgzFExgwHRQoNrk3cYjMMDirG0SZ/+wYlSUUFGYBaqtQ16LFfFVF4uuDRQ9JValWfwl5mk2U
/1U1zeTNx6dGrwTRJGq52K3UkPTlVdUMDRS+2IU69ArPFZSVvyzX0gRxD5afFbFwDlrW6zF32COY
ghZ1aFQkFXPPibzRe+RxOMK/cSlWJcQi7N8DWSnJm9YnmakBebgniYOShhNFuLVdh87Ub+2weD0/
2PB4tk9FjVEmz6s1cOU2kqoXF/QoSMivXQV5ToVCIa7p322XXYshf7zBkDH7EcwmIby+njTpAS3n
jbiHZq5GjRNKPYVm1bwOf2pRO4q0jWX2MfjRbti8I3aZ6hjIKGLhs4qwyMqtL9tGq2Q0fN2iQ3nl
g9ohK2NJsopHCzSVdMxZg5OSkxJ/M6aSsUfi+Lzi3RoTp3YDguO6CcFqzAp90SjTfeGSBM0Se77/
pDgWgXWOh+xa5AxnKQXKcYvUQyD/CfJ+J7vNKhozfle3LYnWM5Y+IxPL2wfH7wTDLhrhqdE6lhar
TTVKZW9xgUUxmSU44Lxki43ZhHE7mTTi2NVoyYGfnmIg+G+Dw6ooHyaUlcBGbzSlc8cqnCfzMWi+
5g82jBaH6PUPN0Uta67IjAYxSoN//Q17vKaOXqYlD1DZavQlO6GauTX2bjwZAjDSaVaarpflJ193
aIG3oZNxgE4uoxBUS1YAiApdmtgtb+g2qGJ93ucZLUsz1Ui/zeWRIOdscsCnjL4PQnGXE7w33Eew
kD6orHE9PTesAZ6qsFD48D2/aefgPaiO/bb35dh/heWByx5hfVZziZ83CqjyNgmpJvJwS6pxHNJB
yhXiD+4dqmkteutf22+YIG4/7Ums8SA2iEMZrnnvxYkkVNjzIhSLj425/djLW6cSxsXEr27hDdl8
1xp6sCj2xUieqQe4srW3Z74DWpSY94tlkxms6I1SL9ClAV27ty0eKmHBE303V1+k1nLQwiRUhune
5I4/YirZgZkzAFWUjF+VoY/N9qSd6rK6nIoV5PbWBoZ4tfvharWNVOBQbZ4eI2ijaUh8ax0nPui8
8ULIikd7HpMqqIcBFol+mtWlVhFCq0PAnUaWHp8XCztCxwSunmZjNvbPe5xPbLMuXXqZt9wcRgz5
X5HkEEMvFAkNtiaIKcqw+JY7xgUQicAhZQX9xSfw2k/6chRHUc99FfHPKVPmPB9xi3QKW9ikV0Mv
vTuvJX1hXRrb9viPjwk+bYZcVtnBkFey110AcDl1/P+OL/Zo+Ki5rwqFjzqANCJPFJ68+dpzpFr/
W5IkZhsHwEVN6N97scL7pNPuaWxCWlK16/CevKttYdFXnQ0g9b9cC1eIjdrlgLhyh364cqRFNe4w
JQF2LHJsJfLTVokwnPmG/Wd/JYd+3QHuvbCMRlR/zOGq/WPhU2wLk/e7fBKRN4+4AzRgqaKnmovW
0qtqDtUg0KmOYRiW97rzzQNRqdyh+P4lSTYKsMw6TphL9ZwKYitDRAmR9MuomVXGZE5wffYVmuph
kcN9yFu1f1PhAhmJDZF8Orj4fqJUeNpthizrCppLQtFxF7HHS+hBcjgXdffutlI1BMn8NCdXDQQK
BBoaA46G2LLLcj/K6suxiERLG9i18qvrycPjcL2P9jZg61nYqWKppEkEqzJ6FC5XnJFcXte0a6tv
IMQJJekuNXrSXQTjy0SFmcBl1voKya4e+D/Lq7EW1eH1rDMkWXQIlUZOXj5OvHnihnIWqZYTLbfD
Gx9rHsvOfBbR0C5vdMg6/QMZrOM7Hn0eRGkIcakWz59rkAaRvkoZWaOlJs9+/94rkJm/O7Tn/01f
MZQzJIOVCSAY0dCDOfNJgEXrDkWP1Lz/pY4HYQP6RIFpsoxf8xkT8DUAJZ2PoYC5B6NtJioKZX7G
gz7WmtfmfJQZCJXgTz90a2YxTyN3omAVrSthkHpafpgBnfYnmHuibwnsO8l4O0PL5fH/nFqv40SZ
DzIkuHWCPyyR35qZEoscgsAUM8l4OpfE1ggb664ZewOYe4+W3OdYlluVfR7664zmF2vVvewavSu/
dO7C8ugED1HqgysgqCAL3YvjKVZQjVeTcvS0s9QNxs8z6uhGeS4yTgq0mZiVY2uBzp1W/yr8Mb6L
Mhfovm2WayqHMa/s58ll3VfLMl4sRLyvD2/GYb6oSFgrLxeqtqyNfzvtJJKBRRlBrtxV4w6kppgk
8uje4E5//kPV7xL89TS2izMdQ9Jxzndfehg7sscmNSrwUrKLP55/HtYlsed4diXR5POvu9dQConQ
jmiWVCV40VJ/My//oNy9xx+cD7VsTW/kws77/FXodJs8BlMl5sIyzGXHQ38fLhSephjGhqvoa03T
BdLo7mJmwW3Dr+ZmbNe9peHGvL0oxZeriY7O/noBZZ723SSu9uD5Vai7NkZ6EczmqDxmvK2HVhZx
Epa3sLMgMKnSjuakm/x14JLeXq1WqhCGB28dTXKxZhTDcmXEnwz2zdbhQcPFjmt+nXtDscvEICX5
+cmqhKI8Ag+w/9F9XLf+N1o97jK/XaGP1QMpNSpg5IbK4UiIQ0tJoaxWZk/45dCir4z6Kvh5dFZU
3o+HOs38CgY8QyL+YsHRdm4OX3gjse5xjj/j7BVOoNBJVjXz1hO+g0SaUBjaTfaasdgIcbHlFamE
DP7PWUadZA9Pl0TINhmar4diGO3OZOjxskO95E/sSX4zH2cx8wH4v6za6fOFowiGxpfELFzw0yqW
EUOCmu7gRWCRuciYXWpCq8N/Jsrvr45f0xo8IxJB4bM9QFIMojiET5twXTVnWvlIynd6ijxBKfBu
D3sZYRz6fLdaZYqDp3Kcln8EEpf2qaH1OofBBBefuB+GjTG3WyG6D3KdG2vcXqVtQ8CWsHor4/WP
JQNIMtR5efKa/zhQrcsevYUUEw/37lSflog3L1WpyTLMFjgkvpSGdhqq/8oPkGrkiLgN81J/4DHh
LGU/h0xPl12tBn58TaoSTHLs/L+mkfZ8pLeKjlpfXq1BETLgY/e8/Ii/fJkDLjCmO0yZkNMyjBcu
MA+MsbTZYSRTYtzElo3WvW9L5Sjnkm2PRKgn2U66dQ9DJAXcsPs838JsvbhMn0Gs8h+CPm9tjK7W
GXOHLP83iLT8Wg5XNG6gaTMcH2RQy43ZM5KCbGQ4V0S3IVrQZnaXo7KR9xQ+jeLbcc0T5eE3S8LM
C00RtU/qbW4eqD594+8WVZ5xUpx9l832lvxAAKsSxoB3lhyU5gcgX1VSktD2TqRhb4pzZrrlBAHL
Nv3jKYgfNvOUTAhth5owBA6191P6hRCl7lQ42jlaDpkg+IhT5ByLMu7YS39nn2sxDMfSOJaRablV
J+NpuaS3zsGtF19svluGJ/10HHDZguJA8XSUbGXrJ6hGEop0251UbP8apP1Wlg7HumQWnesO5PAm
6Ife4+1T+9X9+pSAkgGhMThKbaehcHKYTwQ2o5URIIzXTXjeZy1qz9idjjyA/emWnC63Zp71+FN+
B3Mc2UfPjSzSi18kjN3qsWrcls8kZKni+TxJiS6fyGCjbaxeMmrP43GmIu8s0L0+g6AmLpi6LJIJ
q0FQkqRFSun8iGS+LEDU12TU0/vo7c6KBGbYf3QdsF7l0AH2ReMlquLlNAliaBYwYANWMe9Du/kg
zquNpCyjTrrLXW+8WBS8+GuGuy8JF/KGhAhGM/8ggXmsXjOW1Ejl6ISS9huLTgzEYdB8dpxrV2T3
JHcqS3U3+95m0oICIdTisLivVaXAl+WetvPXbshMAUUSWPfNjQnPNDb8NZ8HgtBRjWOQh+mZCDZZ
Tra5SnVD5uUCb//7XRJj9I8WaOQHEO+YBJQDt6Jd1ZxsuhZXl/9LdSDSPl7D1foHO7P5fbfuGjR0
rrlhuleelRjRO9HlRIgcC0tN7H18soARo+yl05HHG43gk9PXmH+4CJoraZmWymDma6vXSkpEnZbc
ngTX3zN8MwhfyKUlE/vJ4BlFmo6NxE5m4toZRLrTA2C5WUa5fxdSy9rsUpUwgUqiImBrgIoszM6f
4+xsN+Lvhrd8z+BTxPCFiH0mfCKO5BTssyJYyopRz88mf4LgtbBzQ/HoerDOVZJHIiFLSqYcKs4f
vKFJNP5iLNoN4vTH191RKA0qEtcyzjN/Djmd5fHipfWLW5vvhTm4ONIChsqlJwPy2/F68YR8zfeA
IBTp9w/RoCF+u522yUzTG3bQWALTUl/yk7Ltykw+9SEJrefpgA59bJfSoqo4v8nzt83n0DjuGT61
RJjMG/eSHtZsAKEv4RKzr0G80Oq5tU4LacPiOX9SttNkoV97/8YkJIF4C2ui8FwfhEWuDXGyQbq1
vCZ3gs/9H2BavWnz6nthcw+PmNN/Ydvzql8MN1BYlXTj7jMe4jTxzFkDirI5vNs1Nrydu/SuC4ZH
Qzi4q5A52eAQHL5hHH6VPtKHbXZd31GK+iFRK6gSRxBUvNeWufuhGVjO/BUCQehwbxInbqbbegtw
PKyW/j10lZa7dMyr13cgSaQeOj9Z1wrfEL8oDLJLZQjXM+dYenSX1OW49/nDualSn3fFvdJEfMO0
f/4MpgDBkZSllCbjcmnOJdObBHBsZOZzqN+Tho3+VLNRdP60PmiM4t+B+A2p0aXD2Rf5l9op5Im1
E4gF0Iyo+6xadkqDDo/5J8eTnveRwHyj/GlrA4rV4H6xiDHdeOkar8OoxnDPr6TJJ5+1pbi3TXS2
heLweN1aQqLUnpsSk2d7dvSs7DNZi/AAn1EDKujIWP4ZwMOt2nEiMYH9nFJxfixXBHR8QCCgeBbw
Ft1VojNXpU0YbGurYoZtsKAImGs56tBCoNlLpmIh5TEJ/N3mqCn2QmKrotlPd6nbHuMu6kmFNG9N
llbIewVC2l8+WVl6c2UqijOguuQF7UgKtkd30ITMJn+gQ5jphy4Pj8oTtPlNNUta6tCCs39eLDlu
yM9wp/slcTT5fUm8LC+rp6P1dWvdpETNXUy1yM/H8BCDeBOYlOxTOFv4iZSd7MyiGePkL1LEpDr1
a3JJYresVQ9yyhTT5fA5eD1buNdJweeiaRp1Zmd4ePEuFQdoLemMMcUSQWT4n35Ia51fMSxOS+ZC
9+Q+PKiHPNaqK16J9o2q57GdGOqSo1rO0mD/QH+U2GxZ+19QzQlOjao5K013LE5Qb2G14jWBprwC
UP7DcUiCPTRYV0AU1+eFxCYQvHDV/xgTDHSTttAx+0VX20ESnCY6TgMdqiN4PUPnIOOE4qHPvNkP
Nzq4SdE+6225Oh/ixtwCDey/Mbu1saeyZ5QtMtLHV7oMkFJW7pn6d/ifmFeeYjnSV/DASrP3jdnZ
kFpnswUe4dRl/tpQzmCwMBruL/QObg5kwd8iKO9CNqHNhACxoUn6XKLgKVBx+vdmFCJIh0mz4yjM
ts63Dgbuv/xtm0W2DLDQO+F6jYNBnF5aEq29GbAoCEn8TGAkz552nMUVmlyRM1LlOStxpieZt4ZU
y4B/Hz94R1G4ncS0itblLDf4r6doFMjMgaxlQij8lKDGMwrDCYOHEKfBuI3o5gkN6pIc6awe5Gvi
9752IVOR7np/DO0kFvXyIcly77rP/VA0Swlc9zePUdq8iuBjsmPueLirj1MxRSj4/E6KzXuQD1EN
4xK2DGioRQt3XVqtZCrFz5rX0BuAzDlnrMsUkvnHsMY1Vga4nhkYqLbOmF7WqF8YvZkQMG8xZVWt
qwUPHmyuY7MrBWkhXFrKqHRh4iGHOHn2aBnfWWjNImeZJGAf/s7ktCeSGVaVW8XHA2ZXhbzCs1Gk
+S6xyZD3utV8BlUeEUiwRVF+2kmBY1GSpXAeq1rzf4j7MTesrCiqSeQlHsBZ6dj2wCyWJ0zczLAy
DQWIWnQmEpUCBZ3X93L9E3zxS7Z1sKKjgI1L43hfXGv7vJGS3mPVeIiSuGmdtS89kr5pTi64/X6d
7yTkN6lcSo+GjEUB4tXHvIgxsA7xQdwvicHKqIhK8a/pSBkR8zr8kujQmO6Ag2LrS7P0zktg7XIj
h5M8/m+GgjleVbmwoYv5TKPdK1933h2tqwpMuscTZxNLJIhRsdnAIMIM6S8XUV+6245nHWAQRvjV
KYdc4weWvMjht0IvcDLhYz6Dl5y4FbT3giD/Dm+EJBDNyvqi/9F9z4VGzDdQsCm0CYNTTjhQKxRn
lrlHUOqKvHZBqp/T/7xMFIixa2N1xjFsujPwV73oLkUlOvH0aDdjBKYBYVtmyNL9taNodfhgc6Ut
ePeSYxVKf0qyiTYFKpyMOTi+ML0Jrx2YPnh6HZGczzuwjSCVFheuIcrTbT5//VMYA6DgmqaMM+mg
Dbm5IFLTsdwHnhhylUR+4nQJnn7oRQZwAr8L0bbtknDAJI2z872E+dZhaYAmzBhqfSLp4tg+TLat
XLNfApJ854yFiMCvMzXx95/6etFxt0E+YqM4SkXevfoT2f8vHRRYUo+Vis9YjHUaJiax1sQrnJ1u
X72o8Js1QK5X+SlWawANucLtGx/EElY3M+rN/wZNA61CgYmXXmxr6gxuGdwpootYcP+eYQhTBkLq
95xq7HXzvQjiIi1gKQzMqmEd9lkDBXi0alLA4gJlPie+wclM70WIsKxlQh0/aBpLUonputUxa9Bv
YMeTxh9MVrFZ4DmJ995jiAiVioLwFuJyKaUzKkvJZOw+eSRqy6O4ksKaUIvxl85PtuUWU72Yf5Kh
evMO7ALROBfmiemU+Hg2ADvxyuXhaGf4fvKcLZdV3uu3Nk4OI3Tot+PZ5Jxarmni7IwLYi3gKKDP
vpDC3g4urvIHUXtrpjcZNpJWEF7U/e5al8BJfRrrwyS4QEONnm6ChZC52QwvsSXMebrUIYtXjcpX
oB73V0RBLiX2qJZAif9BhZl78S6aEx7vZy30tTMBDBjP/qvjLdEFMwkFTk9zg2FHzxMofJBqAFAQ
oIpZjv4MN/x0+kYIpRHHAuhm5ANt7DFA8pOGuJAWWTAWDYxPOz6al5CdrC5b8pk1zdvZsz4c1m/Q
jH4xpqdieeFfpbjDtN11fUHySKPGFjMehrb650FJIRA6VrKwZaY9v2Ob14gMgT11/uKb2Dq+0p2F
2l69uXkDXF21vk83bLOB5z0zRoEz3D2CKyVC76aQPbkJZ5Trj126ZjRwWt2NlNT8nxH5uXh0O6KZ
lfjvvo69Po8WLpK4b5EwOE66S+MYNaKYwxtaS2YuSxZH637ME65z310R4Szcun/DePTj8M0Id8yy
YZlAslVVDVtLqISrxQDBVPF1Do/80hFCV6zGCn4bNElOOl2SXd+6WZiVtXjEqC4jLsV0mvNwQU1c
yuaoqI6io/1/kahoXRnfSVekwqweloez/lECVvmTAZOSozmNBQ/ykFvfLtynZuS7syzl1OuV4xmP
Jxb0yf/K1Tb5O+6anmgDCPpEFDh84KcnFDRpictn0y0ncv3SNojmS/Qk+gGoE3NXgzjf+7aaxycd
NyADloUJ/8LSDwqrHrywLVWBcHWc1LcXeT+avUy491M6J9Ulo6Gk5cKkP5SGjqlG3eFmqZmvr4wJ
MWFhEyViFBIaOpTBz7m3Eaccoq+BJcK6vV+cXkv1X8L7CPaXAZUyrpxb7qWgdvsnpDELth2Z0ToM
CX8mFtyBk6Ga6UVIzGnuICx8Nbs3PB9YeR4cfpSYXmuELw+qflCDqQloaSZepnf1RIrtT//DBTrG
5IPQTBnb5j5DZ7/FlTAJJQa1mjEYYBQ4FN9/shm5lG+zKjydLNxwsIJoFMO6lsXDvS5o45SCl2lW
Zb2gcE9dCCViQKqkLcdmCldg0wgIzFZ13qTjoeMDC2sp0iTwbpensHJwPAIEdLIM9y3pt7xAoIux
uoiSrdZQiWa77QDxckY01I9ViXvpeo31O3EhJYTjYm7R1/5VwA5oIVf35p5YSyxOdJrM7gNX+gu6
O+D0NcsGjATFwWKfDQS5TxaDETShC+0GeMvKYXgYGBh3Y9ApUSIOBfSHcJp9oNhr34gcX3+oQg6h
CQE7L/kJdUvtgyofQZtqAGyrY9hH47xS5+GHl8FOwWUdD0++ppOMtbTLAYGLs8szeW8iLADir2DW
pJ056kRUJBI2D5xwr8QE5Cqw5vqOInnw17MPznnIR/j6oE9gEXg9UKZmXRZEz3iiA1vZM8Ax0cVL
RCorVESAqN8Bj6PTUYRvkyh1Z5WnNHx49lv4tBZwrJXil6jA8bD9ia/fT7BUbxTBrJHeHboZMbpd
1vAxiPIFUDgA2YhxT75rhVHpVisrnZm7YeGsNjZpnoU9DWWc2hN097haOpcrncThZNyIZdqe8pnh
W5sPtxHyudEYXdztygdlYJRlGGa3/UModYKPDIuKu/yqetLjb2/kuJwE7Ycm0XjOqmsVJ2p4pNf3
2KRkXiAo1hDPolwMx8pgCgMhUSbct8l5t+hHwVYVh3Evy/VBqasWbjVvhTLwBsUSIo0v5TMF+WXo
MHOXKJIFTvEQwwzrRTha8fGlA0OSDuowdEe7OuIsfOkTxXcOh/aRhYvIalOyLJGQfe30QHvhHnB6
IMuNiUTMMRaCw9cye6wfpwCj7/zWfsjO3Pz4gSHlFSCBJKg5m5FR4vxLOefUb7uUMSf97PGs1vbk
bdKbPk8NH3/HduJl8dP4JfPF8GOo0e/Ejowq0E0CD+7p4vvAe5zBfcgva+4OjQ++PypCHUeVf1r1
hs8PeT/hVBUGj/1Ixsx1/G1q8YoGkGTZLoPi2msWGimFIGkS4IDvHW4NaGxYui/9P+X91bfaatBQ
VnTDjUCfudeM9MkRtHkv2qfADrMv+YazLJw5dE9QNZTfQzT40Aqpw/QqkpWSgnVCouABTbEag9Bf
F36hp30COI6Lu4ueEPmj98hxKOuIFC7vSa8LrSKzuJqFlnwO24lfaFfwf7R/ILVGFowYpZtMx9Vj
wYIUsmVLTIrBtC52bWX60jeo9TiUt8wf/GbRXsBz43jKaYCGtIRVZX6CKG/SLTvenOuhD7JwModF
5bwWBzs+ruvNw6HhJwZ4UP5ECDIiXNVUGBMgv2PYPsqlYid6ShtZkPj0FNKd5wB7Kr53vngUluHe
YE9EoOfvjM1kN7tA2j2L/Xk84CrJGXq5kFpJ3GPM7Se+7fjgIgKMyVh+7Ua0ChutwsgjYCeQ/AQ0
FdmjsDbc/axVxwtg4Uosg8khMTqS+Mlq0UO6cQJsOV6GjuAPMh8eUkZPKUhnbBJP5MApne/wZd6W
g1MYe4776E656+ASLnar2IYGWFobSpnb55eJP6t1J62wMQQmDJzWxDS1vNed/0uKp9vtLYUm+2qq
cn3O8Exq7YYSzbOPzw4PUOilZfGx8FT0wRVbstz4XWlyTj9S6ezdoc3RHU+D+5lVnk6tjo4gEgjk
pl9J64/NXmZgMwuqBMrdjy5cK+b0xuPbbmavqSNljH1/HWUE8fUAd6E6fJyHpzt/J/kzEAfUsxEr
M25EI8cdbX474vFH1TGeYqDC0Op4Z17HNAvexXfu4U4buiH2eRiGsfJeTM0WHeZxkdXe6mIXx9YO
7QPhKeIif7J4ORuv52u7FIKeh2T/BCTkvJvUdiCXcn4afi4XaoAReZPCrdZsiyf2nHnPHJUsNtKe
3CRHmRqtC+IVAF8piLHD/UjAkC7j4v51oq++uIxlq/oKWVpB0Q3y4y3iVLvAe/1/NHxSBtaEIjDP
+RdxYA6QYgDx7/LjGEb/qUg0zaaV93vxfCNuRMLMgN8vxg7uNC6mPHjlPFFRoMe2H8L5r6fGf2/F
b8zQNhjFD3gm7bqF8LeGmaOC19E+vKEcH6FCmt87yYL8S0WhhuVAuOFEJCKn6JG2YBVdJHTNyC0D
HxCQdXJBwJH5aKhCcbazD1bClVS4CGl9AIX8gVfFAs6BSzuoyv3nVF5LY6X8UgzF4d5h/0D7Ed8B
keD7gnEBOVQ2eySN5+AspaaPJK6almo3g6U0suT76BS6JphNZpBGn0RLafZ7WTXavk1UHhqLEy9M
s7EoR23V2YAVLybBn3p0EiXjZ2RBKZNWb08wCKoX2xzFUUDOSF5K5omy7w8jS3c74kZ5AViS4GUm
fHwW8dKzpE2f468SYbwBJN8VJhQCJGpOjd3tFY1R75doEZnmOtu1IvKF43t+et/LDPN7B5ju5yN/
2RnaiOfOUhdhweANIPQ6pOwyYLv0sQ5Ur89jB15dazRs/lFIpPGzeEWUpuplOBL9ovKOZ3eWAw7K
2zrdfM6Dl1mwcfc3OI+jlKkqacj5HFRobsyRtrv9iL6yF5nPn8UPcU2GvebrLr9uDm+k1S/K66mv
YffTz1V7iaDbuYJZjSsCtsh3pMsMojRThslkAYb1tG7amVEsb3mvORUgHIqqD25bJhrYplDo4GrZ
2fGhnHqXww7a3POvPZbvhnEaxEZT40Q/R2ZOLNl+n9e44ke2cpY63icem73JleGg6gBP5wDmEKQN
Uiq3vcOpRmPbcXpccjuOI/0JB3foaqENQuOyL8uaPIhcU4lk0U8bMx7KgTM+n9sm6SSdK1kfIeVE
FCqyz3G1G6H5gtChssxQ0hupONzGUjY+5jBdJh1W/Spb0EGUFjS0ZjEkWOb8HjUZsnh2OAz31BLu
RBEln67xNKwjT6gnWamKE7QayTKuliV2WJ94FtwJNNfCxLNl3/yZxE+8NWPap8vCfwptatwTBoMi
Vj+aCZcP5W/oyPhXgM1dFBfFJamZTSfqhum2Nvw08kKULgajzy3Ssl6GrwAng3dcnGwssnmF8P4Z
68wpue/4itpwSs8nDrrKnZ0uMsri84ZrQHJVPuwXQi11q5zWriNNvLDwfT0iDF1OklFygSkoXQl9
+A/iI/BvPZK3GJ03opchBGZ/kwdwx0yMdv2adNIvvyxndM1yVBwVfdAhjiQaSfWNnsU3eVhDvOVe
EsARgCt+MzMmsHCU3MliSCx1T8Trq3nZsMN5v7FxqTIrZcSXz20Dh4ukU0q+vpvW/IzeSNqC0FBs
BJjK7McXxZQE9+3lh3DW/sRoKOEly9NGJgB8LWeELtmNdBpKwzAkDEnvirSpymme5N03BUSwItyI
AdYysw2ZWxZlP2bEV2a+5Hj1f5b1gZKYmsM35alkSxOhnak0i0Sr1jIhEGvxbuBPPipFk0KpPMF+
pHs5MTu8Vkfnu91u4pzVRFp94qcBB113aFfGIbcsnkYpGv135mVxa4XrdpBjkbGJYRd1vUCoFCoS
bll208Yx9T0vhszp3uFs5zYS9/PGskXxgeyb6Ilvqly1HPSfBRh+XY+ktsrob1hzlnv+fiEwTbJK
6qBy01g1dBO1fGI8YHiiL7HXljseCNshuFlzgLuP9u66z2ifelzhAWkBn5ueWUJ4i6nfRMnsSr4a
pHdSrwUzhcfq3i3iChRAfgLzy6A1f130VMyHHozH6pEJ91wUQFMmlS82JY2dZuvg+CEC4xXp5Zlo
mdiQ28HOU1iOgB6XtuGfNkgMHdeRQQmzv2eZ92bkOymyzEsA3vGHVEEqOnlqf7IhsrMH7AlAP0Yy
DgjmFSjAAgjUJ2fWzGhdW8687Z/oi+M9lPqQYNQAQjnsNOUeRywvNTXHIjYgaG/GgLIsmp3xpBXu
D4LYlKXGCMVv/e6RmwL7QJZ5yYthhyz5OEUPVwi+2AyE92K9x7OYGHbLnPhBTpqo4VqKPJTfJKsi
67495n/W+L+7rytLQu/tk+ekBYAdA+AP6WBDwpq9PrTIECd3R7/ZS/WO0IymUaeAmCmtFzUmcLIF
fsphuhZXT7oAh3nFix0l5Asf8y9WfZWu9d9tcyGuEI2T529s2KkDrRhGHNbmmsLA8/Zv5dYJXoYi
6uWETm/xptIWfvO0r4sNp2efd/OHIMBvlfRS2uxlMNQchYwCjiJb1VwjehyXA+gCVD3hWXPCcfWr
ERyc/hf7Xwx+REg6XZXE1LsY2G1TfXPq+Kz1Fi1VMfTj89ZFoq82bgGZiz0dmkFqhBQBtzEZ9zFz
4dp2N3SD6MfbW+1bO+rXJ+/ViZ0pqJNU5BlHTJU/IWHspHMwYgTm9JYEyJbG7iBQ8FOV3JCNzaCL
jqJ39jS6LGAIvUhxqImxSDPN1iWlqPolqXCGHtoNYzMVALu8txcW8hy0NcTGlhPP8ous2AinH80v
cKcDKxC6XLr4Klg2n18J75ErzIoeLOSrBLpE22SiDR35cZHHUDFYE3jAjaF1LWKo25w0pNPQ7gmy
jKumponSuW6n9ZfQzG4fLsmbttXc6M3RsfiW1VS/HQOJiPX0JuTOC6TNvd5YGLQO+CyE8Yl3f1FC
08qEeGPRARmPfQMC28bUESCifWYi7xRKZrRT+hjnUCLmj0vGp7GrKoIiRn4rF1Eo03XkM3AQfSVD
dNtJiWs6Wo5Y75Ei2GWF2A0GCPW35/9Ide2jvOyN81vN43WN6N++CoNP6scN6uuyZUO9/IC4FRbX
ePVMiv5yfDjAikC47bgUAinTfE/graKcfseqY3PwA2sIb3ktM1x9EnNTFxl5SorH0YoiuUzCXwSC
GEX2z6ECLCxOzTLO2qE5WY/OyJLNQU3eczTul+CNDazhHgPNa8hGQ1kJkLD7tvWOSP+HownEY2lM
hQQCtEpc+S/vhROdginAqW7dGdHaUNvw+DK2lrynS9FtOXw8pvm0+YLMrJEvr4QUUFc1pwhDVS/X
BxdF1bTfjeXbSw5MVk37bAbDK0qKYrs7nEELtAgnxEmXIkG9oBbPHIYd2QJvCuQyF407PbR7QSTB
lTotmpKzLK4pfIItE6ucnSBPrgGHrTBWpiJQkp1zCHOwLQBuAGS5wccWOHOTlwBSspM0EzZRrFgU
+O4qqMW0f5h/60YjaM7IqM7Vwx3B7Ax0EYHI1hXKY1i/fiv6IGUutwaYkAlbJTDRFoZXlbjgtr72
uaKlvYmIZGpFi4Iod8xXrm3QneklcUdYUZSebm1/E6NXmbWBVqQEiWk9xNsi87tnnwyhmfe2+BlK
NkHfMzsO9isIIBsR3+6LwnqkQXhrfKT+2AXdnxu888gmHvPwAG4DEgBEL6spaUWsMpiFcihsN6MU
PZLZu0CL7jQrBlnn4R8Xf6Fjy2WUQJOEGt6qCWyJ1WoodY85pYB/i400+kONtNwMGzlipwrrPpvU
eqhH2fP9on0AsvDzr0n/Mu43uClvWmN7LqtLDaHEO5H9p5sEiu5VT011YC6equaZgNP2IlZis874
vyY9jA+Z5lGEHIcJH6yBqCbsJvX1S+5J1jkIrQV37+0tBzKlCNPLnN2O2fp11h3qRpsYji3hI7qK
8zPdoduY82dywgQTz7j3H3mF2dnR6TKbySSE4js/XVPOD8ZU0z5eFK5JkiwV9VnYJFAce2pJQCE7
4LiKajy8TQpCZW5LnUgJsCRLlHy7gL/vDTKZ2RICbuh3rogoMXfHP/1O9ftcDsD/J14KdFF+GygE
llP5Witd9nbWZIPR5Yg0YpUd4cIjxnlFLDRfQn+R1s8hKAjr2236a5qN0llMaISY3MFFNF5wEQNW
ggjec6aMaSGhQ9xTITMp09RB9+1ytm0zMMg6HzGRJeCyDpgGIeqfrhrTfyGMZEm/U+PKlvZ365aC
bAOWo129Txi6A6oVFpj3u35F/b2iCaEgIwvQU5ihjS4rPASbO5lpKreeZV4RXD+e1rk0mhPTXgv0
qi2rwJRpEGbKWc6V7tvfns89tfSTIK6+ICkEMEz11OC5zm8dJqeMvVWCTCx2zLtHT36iXn6QrzPF
Vn/NhabjKh5hrtGnRDWWw99pBuxbdx7YN5X8/hV3zhf4WnBbFMOdZVUZvqLzaPHddUgkn3gUaLI3
ucld00kJ39DUGokcSqvVVRcDzwYJAL2+yrY5fKJQ8HzYdIXTFobwLPCerELdAKzKb2bOjmxXnVjw
yJBmmtBtSdeGBhHCNEMQit7Qe3JE31SldjRYEu7RfJtiZuwwnH6o+Oj6qawVLjrAA1gpFO5gPPks
Rn25T3G71kkLil2SupFlbz4xzggCMkUHlLnnOrkE4EqcwDQlGlXZ2oswrPIrrhddt4Z1MrgogjNb
FPJ3N11FUgd613sTKtv181KbOjYAvnIARY2Nqq1Cfl0oYezQ61X9bX/VXjMpLRHypNx3YtIh9wCE
zxyAgMoLCCTMlZT4skj6TnbTYEoar106YbxArn7XQVcviY01huihwzJgbuXjs1+dkxrqFEI2A439
w0o/wrPzTckai2/fXmQ2WfN75c7vHdn4aHCOWHErFZi1ZxZP5BLQADyoLc8wm8p1N4nXawtdOzfD
zU0NhtSUH0nwLnLfyhgIvPRWGr26wXpzr22OC5LPgeAJH2tNjrKIMqxeXIwtaTuPJ/Af3sjtGNiK
sPjHMuxq2v6LwRud63DQJox6J2E80mEBccG7AkEl+L5zHfkYwhCWDHNfAGlxlNO+xFLNQ6XG7QXH
E87Pc3dcQ0arSpkfAMS363div+J9gywQ3GWdm5hq4oMb0ausS6Yc5s47DpYS5W/ehnYX7e3dqrcT
ZmRKuGODYHdvW6K+x6m3w6EBWIzYkXyQ+e3fLARMW3p6HnltVsQoApaziR1IFP3GCwCzdh7aAULY
jNAFydSVkuSYtPuG7P4AkgFZgIpfSJlnH2qJldjaLElecSafSqk8+KvAArNbAD5xkiyxfA3wIngu
z37gmB2DLbxchHVylTsAyYyKnUubjvzdHHeVPhXgD3CEenI/sqX3mSlt1PX2ltr6ihX6/+sbFaQ8
PgY4AU9VS4gJqCV7H5N3X4W6CmYicyAyv/FYX7KoWD5Mcbt2bYrBSXPxMWOS7JHIg8oyjkJzR39t
l+0Yyumwahds3j43tOrD6F0anEE3LRr9knJ4eFqUIkQHrqPaDGXK2b0H1BmZ1VD9oAvcv2qH4ESE
bxdqsiXtzwA5YYsld1/zFk+bakyPrV8KQTVPBzsSfWOBxQh0tNz9AfR/ZsGu1QzYOiL7gY7qCoeK
8UIu7Rg+XOqhmaISeVWEjldN9mSEr6V0zVzfTnbVdy+pDw+3U6Soh95dmaOr1iDMzdArfC+2vYBh
PXywjiF/pGa0Gef9y61iQP+GuL4QH+7cn0PUZ1M72z3YXv4cPAgek2Dsc4hE7fXsV9oxLQVNxbN1
O0EMyYHB2gNBQG9r3TE0DFm4RAmoStZPiOptYsGcqB6O/DHGRSspJKjGsSSnWjCW3q9rYKQtTiP9
+qi0VW6tttZTgNf0b8WmLfYeVuOZyjuXy17AizwBsRznzJPDMqCc+N5M6TvRWg7+ehdS/otoJxUM
aY/ZZnSZLrHB0nE1TbaQ/8cGFm9YhWJyw1iP8Tz3GhGA/l3GfbynICMtHDsOhAzKCcUVsKdugBeZ
h0I5VGInCoDhWeLoSA97ffq8YkiqkpKgtLjJA3yFNrBtmt1nPlGOqebl0IIXWpj/3nRHCcqyns4+
KoPVNZH6j/LIUpOULoRT5jUGAFz/rr2xSttAPzptz4Pp4BWqHauatuCcgyUwyTllvW2RzHVeAit8
raPA+Gg13ST2geUYCmjmHyUkA/9okt7cuNBmql2kLEm96boOJLA1uTGgC419oG26Uiu5/YV6XaJx
ARHK7CvAtSov2T25GnmIp5dcAKdUqjdb2vKksN9sTCpdzIQyCuYSQY3LcSfn1j7sI4Uzeo82Dbgv
4mPxv+o+bv+NgJm83wFZaRlCrhPBsbhhDucw8FS7sFbo90WuTl8qvmODVehg6ebltWgO3mlJhzph
lTBmGV/16pEX+VGKihzafFNoNWTbZbX7HWgQY0cNiZpA4Ju1ETovyulACwnpmALHPM6eVMt5ZnzV
/3s5HY1zreCHKLy53qUTYqND509qH8KS28pJ2uBV+Y0QvB0EK/X3JH6U2hJe8KI4fTkoHvhK+NPZ
dcqRahu9LtbaetP3aY/HU84zWFf12Ldo010uyq3DcO9StLebANrAAH7uVc160tweezUbLKATu9Zy
4ptAJ4gbLzcJCPiD54oyFlibU/ufp/xevq+SVPgJzVMbcs1XSjCS6tprLMLdbYOPifZiMytDZvQx
SNPZvNCZo7SLjhMhbU0DIXurIAMmczo0K6O549YaNBG7+5XMUyG0Uf92Aj2rXP90NxYj4R/Eom8t
R4OMReo1oItdY7YGpNiaG+N6O9VZQlTjb4GpU0/++WLY+vn9Rk26ZQ6asEhzA2Yzg4aMBXGr7h9t
iZM20Q51trotWk/DZJrBAsc+wfwjU2KfatjN9CpMZJGdkfo2ZJM1P1XZrppUrXqv9Lg0aRr/FGUW
k9ifjAm+P5crkrCSsCBqg7/pI2UDrPGLDnhxag/t/0DBxDogtnC0MUVqIX8Qhs8eJXUneVBdoaAY
xG52mpVivhDM+6WAWjaPV2/w8z5LnQbn4+TQpTQblz95uUEfHVOjvb8U/Xb8ge+566pxoDhEi0I+
70TBw0bH3TRRfUUk83CNK1P4xa5/nFW9zBDBQjA+JyDy+9mSzSuC6/6s1eBJIHaZbSYPt5zDi6Z1
2Kkm2ECbKv/+VbRnuweKqmwNTxffTSkrWkHK4ikojAv0jIlR2OtbMh1ydP5e+E9uwpby8SKb4HRn
AptI5/4h1ZnRgpIgyIZyiRmKlux+6KmXCG/7LcWvht3+8JlUSsLmv/MMKyUYWOVYFKM9luuhN0B0
1aqPlEo7L5Sh4WkcxWWeNJs9pA2k2j4pZrAmVKDFlTIX0T+YwYNDsKBKG68uWHfiLRTeWNOpYlLs
CqXCPxQQAUY7B9lt2PM0ic4eo46Xl075KGEYW0x/chFgg6O+eiuOW0N0N7wl2RIPDlho2Z8JJoyW
Mjt5CerHylbcqhL55C/p7llxpo5Tqj7xnTPOZZZeixRLQp2f59sFX9OwkWROcSZ2gn74JIeuSycs
NObdlKpgzCaTCD9nZAqBZegpGHSdsiggLMNeaQTnuybMFNgeBvEmKVg7hlgdCymGpqJ/mhrqOjTv
qtWpriyCuvbVdo7dmB3gqUYdOo7HIEegi0ShEmyEd+vmQ12TyGrxLwrZxHGTFm3A3hVgA7ttosYW
D6L1qHGKQFXC9DXd/yqFfxWEQajczui0/KFaKg2S58pXveJCzU1Vv+yWcAlFjyZQ2pzNpRAKfR/P
LHnS9cnJ55APN6dNIiofLF+H8sefrKgE7FO47bxtPijuqqbCXC1R1yA1HoyFkIGJWoRbDM7UkVR2
W1g+qsN7zL+isjqVjAtSrwkdX6H96aepodpe0m/a/xH0G19yq67Sye+qVqLYp75mO7EOT7UnxQA0
qhdUH8kyJ5ExhgjoAA8WTRY3T+GbMjE+6vk288iQwwd5KLsP/VO4zt0P2ek90dSjIG+HwmIaKyL/
DAe8dqJc9e2L54wCX1+UxDPijvXzYXaTlU43gb2qSsbPvn6FVNtqQGcPs7lC31PGqphwrDvPWMWF
Nz2Si/12Pe4LLKR5NfN2mz45i0H7iI0Qc2UyTk9RtQQ9feD/pjqEyxgYGFpy05l8OIG59aC0U8Ou
Utq2cLa5yt8Cq3jSy0XcOSgi2/9khfQwaTO1tEkf6vpL18V3QsouzpnyCJ76plbfGRFwyo3L3LM8
0okheVbO7tAAwgE7brw/CHQSx6m6YqYJQPnZtGk21M67WOCDZeXnQ0FRpmHsL5A57c71KZAwCn5L
jpgu4NaEOnxuvcRng+69manviG++KzF5XjWZNVnI2kgI4refT0L4FGbiNuslOt+NkJ/842rdA0oq
PYX5Su07NZKbZSvkOc9yh91/BG4bTILh6LY8GWjl6AjQBR8SsF9qhxuMqsPB122AIsaVtkgbaVZX
yWccbk2gqdITQ/dBs3cxNcLOyPsz5YWZxe0UziFXsDPzb/2WNyxZyhbvHZ7g4PT9ZycV8LHTutr6
CmqFtadz+cirLFAxiwgZUa8iHVSV1LewYhxPupwfOZx7eaCJpJ4UJ+cKq9L7bxxjMJbYXeD28kus
X5JTG0oM2BjVvyTd/k/Twqikq0X76n0ImGdqnjOuszsga6+lcvFXzAXs47g8eMfGpFLPx3fvd0I1
y3GQ+yc4JXvtMzyf0kYgI5GMGyqvswSM1dZqgBIaIZegBgVwhMwzejPXIhteTcBYrIjgnKMHUviK
e4QyMt4qCJgVhI2k0BCzGKJ2Eun8f63fsmVZMiGq9GEzR6824sc67+IPjZGnhN2cCwQ2bVDa6uq9
L3ykgcmBAJEtksDSV4ziqufU5R6Pz+3Rn5jkOExA22GuSLBt5pHMkpLerf9C7rJovinxFPKwR2/U
I8BNqQEyL3WVt+dVEBEcUrPN+dqTkZ20nXNafq2buhBtDl36ESXa0LEkFwEXfczD623wif5M7AwH
oB8bp9N0L2GSZ5g6dVMjyHXk+Xk13UuwJV7T5vkB+tJ1Rmc/3wrleb+/qyTHc96k9XYrBo+zYykd
kEOnAFzRLkPujUorq89AQBs4MCVihNlvHzpeckdPsHQ/qIFOkt6YeppUqGC7IDCMoQUTkT8V+vQE
fnJQLHnyOtR+vJqMiZj27F+wmLKqjY5NL++bz/NYPiWNXcRNbKb4Mt1Rrv1PIHzW38RCDb5d/llh
0ZPBwHyPcRm1dOugVzKp2/bkHsxSt1zLuqbU5RVUEufHt6qnbvxMEludhs2iQbQ/jnBfe1slAkye
OuAOk9Bf3gZgBwZn336Dm55QbcDsuRqr1DOQdbvjx64QgjwZCAoO7ewMXKeY7AF7A5FimtVlmJHc
IoY6CDDVL6mAHKwkscvNmB4YRhT0EEyGQFPtliG1RoZmo4ugjKdZPtOWjV9lzaOI58YG5bPBuahf
njdlFYdbHyNcL1F0r2FdPKhmW71DPTXRETL5wI/xzFDDeZNA6vKhISrsrHakdyqlwqxSOuxkfkEF
NHjRenPMFpZdO0YfZa3pfy/dPg6XR1/JxHyUIGOx8eAO5GMFcPKB0/TrvCvtixCqa5U+5tJmbNMX
UNzN7XLRSL486yeQgavdRq7g4BKTtjc4x8ByB7w6xnuR+Y8s3W70W9G/MQU8LcLtC65LipChqIMf
U4n4zqZNzOOyl9PNmB+c6U9jsKgqYJ1uoSJ7ZqkhyDQCtlKVTnmdan2JgqjQIy/Hp98Dwai+4r+G
TUOvDwEg5JuxT/6/FcnsoZBTgV0i8d3ue1L4GLTCz/Y4jI8mloos+T5Y5bedzjwjo6I402/zIaY2
j0W4uiRTLm2iynR82eo1zMKWjf+GXk9SQwqFDPnBnhk5SzkHDuyKyquAMEVA9U/jRvGlrZ7dw28M
P6++eqMgpdFiKtIlQUk3pj4CRiraP4XYqMSoYhM76J4oj8vt8Ow88gC3/tJa/nGgKifJaq0lLTPo
DfITM+odNkpBsi5pTEjE6Fj/K9xOY3fb6q7bdXNGhyccyTFOuChV3lvAGlfpGAWaW99gBNxT74GL
YbjEzmCQXo/xhKSSMbu0igytDPUFjjHsNcE8qCv+4j8oWdCMtZeUwNh+nN/N9j3VYYlR83aCfVKW
KKvJFQgUdLpJBqGkaCtEVgHzBT97rKxyvULuVmZk2j3VLGxvvMrUiQNESSuvvTwFVevxDcr6vybx
taCby/D3u+KwSR519vYB+ASe581JqvzRN/jV96ioTreEiEzoDn10TjqNCgrA8zPmuOHOYyeTKgjW
iiROB6Hk+yzUYj7OZeDGNF2AP3bbwgt/A5CyhH70Yqa0pJUZncBSHalEV8b0X4BvwH+u/pjF6IcO
d064Jy7/F/6mucGfEGHc9ktXL620uFG9jbBkPuYPtwNu/Qti0R2L4i5WjbTJq5u7kk/wpxR+MMLD
qbOB/oalik62qFnyqNLTRkpNetyLTOhlL4TK7m4hKCD2tzN+QMQw1+bhLH6ByVtKAw0Sr5oipUcG
Bz6brHrsNM/XGj1PKa/hDDEqn2ppKSyGI2pM2t4+fpofqfIPvxWTN2QPewtRORT2ae/KKhQ9ttF6
kulQVzMH7NevKBZu226EFCDbJ6uSWRstL5umwe2XYey7PMF9FeTglnpqtSlJe45kF2SKDy6wcyh+
J3hgA9R33dpg6q9NV5UxBozpkNTwOJGSFh6dkgFCXE3CG4y3JDGTWHwtuyfBZCP5SFWixeO4lnGE
szChjMzbxaWqvDEO2hjS9qvY2ulk+3iBV8QYkNXT9yuYIDSP/XAegZpVqf52zIfsJrLrTqQ0rUa7
hGhoBuEMwAElAE5vq69jjtSzFEfZG6AHvzQutfjGJ8pSBVVzYEjjIlDL79UPC2pPwpo8LOopXCLr
8iX9johRRiVwXNDAgIIjcsczBN/SeArTZRWuGW7wxazdTjF+NyDcZ4mBeXz+ar1GOKNhlp9kcyI+
IsIDIi6BeJrC4A+kv1TLaMsQKBNCQB266nXX/onqcXfQrqC9dcu23I8FddiO9inrogpr8+LwiMzf
GK9iN0qhSTZb9omQRfqIIjPxwnV/aX4AKpniawjzEayJdpHKtjBZAw/CMWu6D3Hj8/khbK1m7aEB
mz27fXSCHlYo5Ff61gazZU5SmWOMiLCrrmEcHpAgi1gZ3LyhRJXp23bYtXz5bjS0V6XYmkI6itjo
XPDebjghS4GJJ3vKv5sEMe59trn1hYGRTo8oJGwLyhmkRJGlY857ia1Zpi3d8nKJOBPdg95ws7p9
3IOjwb/3gVQXrhPplINTBB2LTii9QFsFufHvAtPdA9ukJvvNCkwNm6lDnQBeydmlL7AoeSHkUCiB
cPJKNHGv3nDQLo/IzPpad3XF7N2qU/52OxEPbb6A/9YvA4Ku1G3ljINLckSYrMoyQXIGGinjD05A
qacwrJsAGT9t1pdwCJN8WkUUM676k2NKGLfBZsBKJVB6EpcA+5BrMExSzID+MOGxbfGYH2benA6W
sTrrk47GRuIRuH1NLmT/QF5P2AXVPHTYhmGjMNLjG9B5pBUTpL9hh4zFe0lhFB65vo2zZMGpLq+1
9HrcgZ+tzCsxv5h018loGD/Kh3bdP9D50T4yAE5A9vup8MBOBKr4yPdZXQf8oE+1WljpyAgvk5aL
9nief0Cx6sEfwGWokB5Ss5/q+QtiRpk8uPjJzGzYEy/obH+Il/OAgwcfMYq7HXpXnY2jmC9L39SN
zaqfweYcTTsl9RMwi/nzlC1fva7n9aop0+EroiSDGdgj5XnbW/61YuAdLnxqW4k7pM+TVkmXyCJV
oQzYEKnrgPPipLEklFE2phRFRNJTbTtF6z5cZGVIp9dKC/oGOBR6/eTdgh+SzVZ8TUGSpQvTcaDf
qqft/fOMm1P+qytqTPrmL59yMLuiLxdrSG9m0zhlTWLeUncUNv8Qs1ReCGJCghqzQ4mMUxKRm3Yg
3aX9kFp2mC9tTJKBPrENg/6BTtLGfbvhj4qc/DpShhuHffUe/ftAgIlz17V9MurGA5+VOB9rcvJx
MMnWapsWsTzgyWgB9EYr+A/JvL+wh4U9yQfZYSg3N/kdbIxVe45dFbEGhENUElaRrhcZnXaH9zTq
KAhBimoavLe2paYKixsSb//a/2FI99V61DiIrC8KPkszImwH+CtJ7fbwcNaInL8PbzVOZWIV6SF6
Z5OZikDzq6z47S5qB68X59eXGo0YOh3Vw+4I7nx+wgf4QHLTYkhY0L/XDg966+SB/h51DwdxgoIc
/z88f7VIX7wbnvzoHgd0HSHE/KFbzRpoOTuEfUIYJfe2Op6XQbb9tgc32kxq29svYxl/ogy8R1QM
eKog5zAcUYavoHtIDlv/k/467Id9O6ZW4kJ0fIt2zOFopE5LCLu9hHHd6iJUK+/VLD7HzE878O32
E/Z8/rfinU4zrRfanziZXqvZG5ndhrWtn2+65CEEwzIUXz/wkfL8mDtsGKqsdx+pCXEDvFNpkFcv
hsDrQILVsSSED+cUA8gxRAoGd8FpF0VK7+NQQL+HcKc8nul/r66dkAjz9krLiR3+tY7NcXv0VHdU
kCZ7H1RKOsoRbHNz1yBmVsGfD3/K6KJuCDORNgmXyge7tzJAnbDvl0hL3DXluZc93r1sthPJZyE1
Q5E+KFToy8sS6HJWgNxHAhRQz8BXzslF6GTBwLClcobmGgXcHLqZsPKq1s6UR6RZVQ/mvfYFn482
aeXbbhlIyzMuvgKBiiEI0dEVQ9okwT0rl8e4m+aFISVk9FRUZf02LB3gKhkGFGcBhXVnexyTYzlk
asZIiJ7SJu1yl3aocmEwUKbDFjz3CTj32mHpQFuJGP2LSLtNb06F6XouzmKpvREXzmRNxtkwMLmB
dCFlQ3k9pkB2ubfskTX0LlNV0E+l4Xyv9Tt5msHU9RWInzBU3YXzTmUa57edxoJRE39CG3FWrfY2
j2Gyvvy3mm5dlcR4eB2CN4R+aVwqwB7f5THiwsTn+ylnAzM7H8tXDOElXKCHOzNsvotIN1rh9sBD
oVxhsbhtZMLYRYRaLLdy/S3nAlbAkF2hi592Ixw6mCLL4/FnfDF/liKXoNuomnzgTAAN0wE/6VWi
WHRCQkP6yfA0+7T1iCnvVOkDTozukgAGucEPMNgpkJ9MKSOopTczkQwmQSRDnAwwDJ6L2Pw1ZdZj
jzdS5XcNGVpLplU51OMau8l/zEXB/HloQavOs8H+A/LtFalP8yf8M+EwEB5LWpR/YDurDLakLPnO
pa6hY4z17ZMexwIoGoM7sjmzuy6aUGRzNjG2GbKZhw9pOc01H4ePgDn2N2Qmr8W2rcK+CkMg5tq+
V9ULQpj0BEXcWxUxl0y/Wq1FTfLZK1KbtYSOZquYANsJrQqTFS7M5Pmlu0+jrmgOnGhel3JsOWQ3
jxzA9M7JWEVrQ25EaDPnaqME8Q4Q70oxwtNq/Ig3sMYwp/iWdrlSiZSfNKjHok2xFV9stLFsXGAw
Krlao1prxObafcNEFDm+MljlOWadJGPXhgzCPC89Nn7GU10zIfF02tuux8EbJPCalN/A95HgE56h
bqdjGheIBBXYmNrf7h1GHxgI0S723Dr6AuhDC1cGwldGMcNi/0MAU4iGHJzacJv+SxDjBZlDI5F3
w7PDBLyFyUaP/AZhnwlhKK/YAX3bMJUrIlOP3VwY7U29RBcP8+ewWpDsrmquxem3pJH3q23WaWdZ
oQyp3e980qEDFD9uz8jcdc72lYvZ/wqLrPl9fSCKhKdhwJhW+iYFWrQvDrK0/vt2g/Ng23JztvW9
lBmdggdAjGdnOJhHBM57dQsPeaTP5i8WT73nhMmQdO5ld3lLclj/cyf+rYPVYmRvlxlR4+kH0ha6
zw50UhtIbduiAbX5Yj1lTtlP9Vpulvx5h95trof3b8bAzbCtGdEkN1JCuMMdd8NMr4qNmUoZeH9O
PcMB1M3XXoZ5M/v7VG8SXT4/avuaLMrpRFBr5zazBZdejNpw8DHkiE1bUN8/TWzKqTbmOXVSVgnA
Lp8AQyb/k1VED6ndk2AipOk5jdb/d5SqihaVp3J7Ou2UAvjk+qJSRQn/V736K/m5R8keV8iGasIl
zHd1gbz7XkOAECThx8AN0sKT4eX+Mrptz3RBIZMDZbWb3JM94wosESeiKGWN/vQ3ikG5MhvR5dPJ
d3isyAa5Izf2uFYLvoIt1FA/77eHryVyJRrGPxQ25quUIM1GCYDIuhUHTmhcHQO4wE6NfcY6+yGy
bgIrKpw7xJi50p0i9zUeQ1jJ5m4xDSqTQGyCjt8G4bi0Sl4ZX7QKImMCKJloNgz6c2NE4DBfmYsw
UrXbsI1j0YhS8cMDyySRcBQPnbPNYqBdnRpYAWzGWCdy1/JaeMbnYIOznOEo+kcTFm7rnFGs30pq
oEtNXMewSMC/vj4A7ulW0d71kucvcbgzeAFEaFk/EEm4or30J31/1wGAD4r6ININ8Y2XuLiL1/vd
1ri1KyWjaT/fj/K+nht8jrbLqFxsKxSDwaKTOClvyBB1XW6TcQ9AZWlHK85c3L/Z8LqZVD/VZN+W
exFfaqdLUFIEFDgLanUaDupGeIlQNh8RJMceaOk+FZh8faJf+I2spHbkV+rP4siTJDRHhubiwE0Q
TMxREB3aq1jXUrih9dtMDYuEcc+/xOuObeYYTfntMivJMsYfZvVeoF6UDDzh0xCDSt/EBEdycvlL
afq6s+BweES9m0MxWwUX6zX/+bCX6E2YqZDwnWSSSDOGx7YhH04nOmpARnNumxMg0ATwFCO6t1zM
JFJmE4FkRJC1Qb3y2JClp99dgYg8ygJzFPG1oUh2lGm9NdEyvFCM8u1m/7uel9zfQHAHJqqGlOrQ
/5QQPLjRY/fBqu5Ftw3XIv9CE+Bh+LY+mjiRQXZl8pjM24zXuCB01zaBPML5j78yJWsmfEeQCzZW
dYyF/mXpdCaw3Z3yn0oOATtsxP7hR9GC3ythNKiWjLBtqkgJ6TLBAkuo+VeWR3Zs5v6HKsnm6zZW
To+Jdi8rJ75nXf7EkO7c9bLk/jW/0akJ0h19EXhmJEpvPqr34ubK7GXNyQFqPDJy+B9aiHTMTBCW
fY5xcFk34g6iaEif0eL0z4EO1NcjiVOeAjxKkZW8TVF0cCSFEWXvohl0ViWxI0sQSKHSt5PfINIG
ZmMYNu6sf5DLn8kQANgPKqF9lB9xMdCZa5FkPIMbWI/1Cajq1i3I00sbATeNsFrhZwdKX0uGUpDc
v/EPmolqBW0QzaTSSWdSsdfxq+QedKtzhjzpN5tXKCKC1axoKwCAZbcdZZ4PPfMApqWEfY0eGmua
snIDrDpCNGdnElXxDWscQsBPij6g1c/QY3qSXooPI8NdNuoakvlnhEtziuKSXr91VnZbyxPQwEhj
SJFQhQdeC2qerYozDtKXhtBhRX+bxj3QoJfJgo+eBLejFZMuwcFvTdPf1evYOAOewiVYRSqB94En
bPO9bRIMT9YJ00pV/rp7Zt2dU2SuGnZ/5OaPWY67KmBetSuJe8ZOmJsZYRQ4AWfP0bSG01cffO1U
EndtQzb6yeFTVidQUQDMttK0jio3045Dt+kMmfweecSrELOfEYoRLEhsCgNW+tf71CYmkr4tD5g9
pNqSLd87zHKdRnRpYRuPqqcRKZ5hoNqLhMQByUZVUwBh9pNCLfvQGA/+Tl8/a8W20LvK9Iw5zKjJ
3T2FDIhMfqvoW3G9CMWb6oDpYTzsESSVlobBYKOqq+hp+af2fBVZs8Ylkj5kOGGSUAAo132ZvJlE
54p/I0q9rLr76t4NrMRgcz4L2BunFTOFz2suKe4F8g2Q5qlItUyllu7skzk3R6/ijpPqZnXBRrhj
iO6XeEpYsux4t5nSb2q5i/ue33xInq1+5fQvqKDgs3tMMsvVnLsp004vwvRGHLLo+hKI/gcZVO1i
eDeR+EzyYn9npowkivntxaKaDoQ9qGp9/m3nsI7CCT5Vwky7HyfsdT6NwvHDuJEjxt8dZND+6AjB
4rmHGqQRIyZY0Wr/3QF9v+EiXgBtveMbqgoHPsQNIM70Y0leY8XmqJg25/j2Z8o/XzdFY4DTHo8b
LrT+pGxKQRCi9xQwoEg3FYRBLmO7VTuSfsrQRVazWVnrj8nUMy5+fgfDdAbu3FQVK//68Pgux120
fDaTPVL1N8M2JQS9TYIO75FS/FlCz4p5c5eSx5fUHbQb4nKbM6ODneX5EsaZUhZw5/exMKMT0kj0
rkOEGkc9XdD1XbspYtlQAsd5di3vQ5q7k/aJ1IPXjeLp/oX8xNbU8WV5wP38u3afnOGHsYRltY6e
r+YgWM9e1wylckq44WPwwEx+cZf44nU1qZb2NC35xawyt1ZyD9Z/ov+thJZwwwkRTlnx7AlhV5l/
6HR5Zap1lk5g8/IbaCm/YSBtqEUwn23Va8OPMzYZe9CjsyR2WN0ssuKtFLOdzQqqArHPx/BQbP66
YeeeGftgonnXxyidJ0+Qtbty890o9JRiLt1OGmRoHfW0fb0fHh1GKTZUZ7kBCiCqgIlJq7Ckuea2
Bmn6qIQXODMc9WqarrzGf0YxnTx/dliBJpiOObduPk9d2Z47l1syeVvAMN3MA0c9cDxUDOsZbbhJ
xqDM8BJdrhSAxaLne5W4YK3SNcUF4HxzXiy/aNIQlXZZ4NPgnR4y00PAjmqgU+AybNuQbgKdM08/
N0MMiI34a854GKOc98/eVhnj4lCbPc7UWhP2qekYczyUgfgqDIsDFe1kEsgImZwRAYr9wpgJ0ksY
oLTri/6uaGJ2CVOYDvauygZi2+eRfdN9oD1MGa1BbRyV09hUG6BOqmmn2K9V6tJhMWITbhQGAYAn
JRJq5ziXes/YYzEtAB/Lrq74EK4t0B85GrjmSZbtmCSmIbKBJBIlVZRq5oNF7xW91U1uMIz4R4Ko
ZmWeMEDDFMc4QPYQYqqAy/6MKblprf8ryt9AA6ISYRrTpSJwtdyDkBlRc/VmnaH0eL2ygISUmUqi
D8p/blqSnnL/CIXPu2wTYjL9+a5P/MQ0vRMB8orMjJMKOa6Ly0XXlOYeA+ZdIS46XW+uAstBBs7V
Oqjxo7jfbEl3lEPtUhd9cjbtkM5jUuFVWV/EQnMSih74AUYBGydXQPq4zs8npbWB7LLVLw/npyRO
HjZNZMzDaLdpzvY72Kk6EjnP84GHAxldl968ieQ8tLH5das/3j7FvsTQYE6R0HjQ5MnUj7MUR/1Y
LBtAczrz5qBO2WBql00mDuC+2vG2Hk0Oia3La7LAaw/bIGxQkQ0IXQDHaMlsolI3KaDnDATqaUwg
b33qjSTFD9ajXh1Q+HfMF625qs7IzKw7pndWnFOdL5fHOC8ZeKW+tKwyH9fNNcaK+QcIBITntf5X
U72Yp2r9/D9SUYkJJNAu1V5CxMSyjB8vUgn47nVFKy2KgbHj71lbSzN5+kMbCXjLUaJhyQZ7aRBO
mmVHt1vdszC+AfwdAJNNGSYpaFxO+Yjh+lcdV/oIGFAmYSB15jVYqQ1vpF1rBsm3XyoPJxpvquqx
IPlKcGvW4Rpm/U73UsXMDDB2TOKEqYtA9TjcJ+VjLsTux3WZxBqP8Lmm3opallpT0cdktM4sJTek
ZFl3EQLquOno/yz+24a+ERmoLI5X65CGhvH85BZrPuNmauDeYpgHOJdcPWbqrggZ1ql+a0ub9xAN
Ppv+ulwZwqQPInubjX+31zYStfVYCUTrPZHR7wft2qrbe3JKDzsNKlzDWmI4f/MYNXZLbMSoh4rh
MffWnnzCzpdT0JaNLaiHasu/Qc5atqpa7OUE7IM4aQPVuwunIrD7xd+qbQMAX1waNWPigC4RaRYO
6XxklnEIgNNdzKBxeT2rhsq3IlYmzQZFNtuh0GJDY7XmZHvnIP7bTUCxVsLQTlxytCzsHYZUM8nY
OK7tW15EnFxxmIiRcyX/p9oi2NHuYb/radLTAEeUDMPqn96bry3y/3Gc7gmNDGFNz5JLUsBSkY6v
lCjmG8nfGwkoY2pAbPfra0QP0YnsgIiLRswzw0QP1V8n7OWvfqSwh8B10f4QqcPtaaDC+umb8434
9w1IEccpKVlkS9+z2lfT5fj2KHV+NRUlIalD+TdEc5rHPNxBl9m1RjkORjmGSAk9QK/XIPdGPPli
BogyO0GbapiaG3YDmdQW4YCuoLxMyJahtkUuOUnfDIAoR2kuxGnR2ynwJO5ze0b3qy3UX7cL2fta
mgoVB3kuHsfMyOhxygyyiMCVmp80L2AszDqckGhEQuzSm/Yt2ocSv9pxG5DEHKXg2t51R+BXUUN+
E30ycx0czBkBgJMHPhLE7nUVjno0sHLiYhaK+e2fzqXygpDvqcnTL5+Q9bqFsUeqmy+bkK5cBWMK
ctF+ncxuc0hAtP8JaRjpveIS2tfFEMwjlSVTHrfs7YeIFY94aDMX5idOPsA9jiVPDIzm5gT/OdGC
W6apQLXsd6WraFftHlecXssvXBK8LGKXtQFntq+jwYAdMdxScAEowTVL0Le2jB5tB+QRc363DHWw
jY2b7UFVsWNGQItVX02mc4ME8Zcr5zBv+vBdJhVQZR1hBVs0vYCCsmBACrr6sdPfTki4wrr8D2q8
1tpyNsM/0GvmKTiVH7ro2gKfJhDZLMr3zIASzV8xNs4VgYaVoZeyW1UlkQGiosONbEm0qiXjiICp
mbI+KvKzTQOkYEb0OmmBRNStkrYHlJ/+0ky1ffulqnkWX2STkKBMgcMqQDIfzD5BQVjJZ68WHrdM
2mgn7hMjSEwFAXKnDUoisqyHWIE9Rul9DP4N5DgbyiVxfZ7n2gBJrxIauAsYBm9JjtKQF9X+LjzG
PGBYwtxjssxN89Yiiy/a6+OgYWKox1HpZz9PcgUxP3ZYb/Z9FDhOSMvW1T84Dwzw2REwXKN8W/5p
y0SZ/etDTAcv+kpOByMCvbfRHVEbreayiQVOvCrPCCX1my3salq7UcX/T74O8FtS1DydVOSI75+G
/yU7LVxMXxoPVTf4pLAqPsQYw0NmdbkMPmnuye1t03kZ8kNSRcJaFL57v9Nuq+vciwQDZcTKdIII
0f9Qdnfp1CnIYtvhCz09px+zjpx4/FqUEaT9uWwSk1haU1rKuKa+4szXw7tTolHQoCJex2KCESwB
+fpjJ17J9GM2dteIUQ6+iVAM+l30FcGQH6R/3bJk2osibv0rieSgM+p+Z2E09Chdr52EqjKFebga
ROTfspqIlY1Dvmk/jhX19y4WR0y+jNd0ZGtvW9JsKPdmY+nR5oTAkhezlr5ITIWBAf+Aoa2suHSA
9kWIGNidVQ2MjGIK2HlAWH5k5wxRnY1WR30t5sTd7r5LJmgzjT5vrpCj4ydLw/R3IgxieSJLC5iR
Uk206GN2UWicc3ftCLJRw2d1QoaRQ5M0Dl2M/vREwLDaBucyqjIN/cL9Xb4bJx5k5kOgiZ9FXZvW
utfT333JkrUqS5cOv5LgFYgnba6hPuNN/OVadHfIOeKvOmn6xHQSwU4qC2fjcQkILsOqmeLwhWID
sE+WD4xInOCIakf46uMP9r9Vcye+Yd+ED0PLQPOFLM6Ct6zj0XQvQPRSUH3IPo9lma/QRZFf/uyA
RInopCsw5CQN0iUo64nyT+/XjDu68sR9Od/j49/XaKluZBVSBgZK7vNGRd3YdiOL43wkXShsvgo/
dnoxxQl3rFJj8+KbDBa0K5syCJ53hYi3X69M+BHSecmfv4YLlKixuN2aPbi5Fr+0hcbkfBU4PkGA
rFjPD4Z/XbIdAKiVlMFNOTbG+vFoV+PBh+OjbAUGINLXL2+aPfmHH+iOVB0iBZo4DxThIbA7sm2N
kUPF5Af6AYAuH4IhSwxr4IDuXWny0wSuO5sH88Sm3BxHk4QV2FTrRkWxLrfXP5uP1gKZsytcdybR
kG2QzZiiO9Y19GwmYe/ODP1iVoz9JiHW6n1MGdkCC2RFvLvKU/IROhgI0pdPJBsdNdS8lzC+Fyn9
N4Tg24qGrjPlGFxPR0GCS7xJQPDDClBqFYYzES5XIEQYH1rqTfNkQRoqFwrvaFgNo3G3oFOQlRfB
u7zYLQZjDFZW0RdzjRH61mOCYpthpZTwxa2sP3/5EotW654h5x3SQZha8oSbpyW782IRFTEzWg1x
epdewWEQumSoNmLvZqWPe5l2duHgsOxlzJcDS3v6Qyq9sk0dEnLqt2PSZOEdweWRYqqrLscQERA2
5hrVWlos8r9jd/lCZHyq5yN1rEncy++U15dpBofiQezAbTV/i4qdTpog0FJQTI/BDMrox97T/3ho
VnBXWW0UkOBNBDMXpJhXDc9zfl0rnBkGn7vwKvmHkDANj849mIqz/Sugdb19pB7NlMtnvSd+NeNe
lHcdRENEPHRlzIfkfsMG+DH4ZPUyXDszrwneYJ5FUdE3Sla4IT6JEWYX0VuD6UARtkh6zzoOxTVJ
tIYi9s6RrW5p1PR4IUbuq/IRNk8JE9qJe82+5zqKuW8mKP8LK+imRLYIlC9licUjNJHdASFgj1FG
FwphcmVv6TYRoOTzdtw1WIZoFe8t/7IwSUUi0RtoWZb7eG7GVdLJ/sp3n1XmLC7GtdpRVQuq2cFn
9czu7Eg7kp9w+WiUqVMySGpByfmdtPCwz0apIfZwfozjx//rmO8xVou5bBJjtTLbSBPAEbGT6j41
NdLsNWhtBbETuqkaq5TfmSrJkGBC09uSWrj5e6L5keP+U23Q9+V1CSqPT7S/cfWBDSKUaw5vc1J4
YumP19hSXEkFMUIDz8m/Kmzv7qi6vJypHaFoLf9woqIc/EHdUOjLYh70vov5fYXkXFXbvxGirdtO
mHqeYT9QmriKZKrlv+zZ2Eo3DPC4A8LHRak5okWArHPFqh1m6DpE7g4ol3Hst2nlgPpP7J0CTew0
QoZDHCFX7AU9stoqBn996dfkr/2MMpWBDC7bMUmgeQ2aGKd+GOpbYJV1Hi66W2IU3b1HiC/vXCGr
i3GIpQebetf4uDAR1DELtCteAPasZ6EUco7UUvhVKRlHjyRvWMbcPURff+eBJBOgpHaU3DGT4fJR
cdrRT/OvXbMmXb4xO0l7n4nFSdAV71qxncPAx84Fs3Nsg+VZ0JNSDNMXySTKM0U4tMxHKzcd1QL5
4npMHp4LyZ9FGmmbP1WUYmva2DoQj5xle8J7gdLwYQVLh6sdODXq4WFUPf6o6GXCfSRnSK5rnvRP
/91hEE7+aH8n8mZbh5IW2u7gleRnU/ZOzWPglv7Vt2fMYG/HumAk1CZvCRC7WgNMVFI2FlVTMVkU
SBJ2YO6Yj7Ifqw0OQFT1moYbEuvw8oiPlAcnknTZ4cWXaGISXv+VyGgagV2JW97yGCjbK1g61rf8
LD6t1CZIXwsdLE7fZQ4cDZsL85/bZNFs96nx50oC9FodNBsBZcxgAF8t8pZVrzh4UQSxtoMlwusc
4JSMpQfzomNmLtrXa1FOxxnNnUebyZloDaY7PyuZuTRvcA6VZf7t6pL9YCg1b3hlTfWYt1eJGtGf
HRDVmoU6Na0pKcE3hPrvZNUiF5nlh6tuqge6695m4soBjqGGvGqWprw5+0DEH5n3HHVXqTKuvfPn
3IVR++Vdzlqm5NobrM8qLGyFlz6uktxY7tIUUG306epchYDyQQ97Ge/wCUWZ2NkJHvDlxZEg9E4K
W1pCYQibZFx76ruYKp3L1t+xLUTuxXI8zCCmb8ZdQ5V6UIr8HdkK+TnRzPOkYpJiEqyW+dzP+bbb
PpVeMMpYnwobe5lNEbZYp/UjelxfQvAYxjJh9EAwS7nBU22usxnFS3K2MMIjt8904n0cM8juQHH2
WGcD2c9y8Evy5M6fLcvEfbNXvxcVdmeyRsh9cKyFzZwI7qoa+PYnaRll34ZYhDLuJrm+sixTxnW7
CA8cteGy0alrgGwFmXAzxBlojPES0oxqLpm0NzaK+J+JRUSIjzORBWCVWQwN7s/NJICxmedp9MI2
k1EorjjDeZQpeUyCAAL5R5zKocgruLkS9A3TBixa0d9aVJgQwkTuLYOQB4edTk3AGRp6+khiNkda
WlKKO9hEuw9qTgRUP3Nzit2n8ZzTAGsz3OHkD3QOApKcLyc7UddgPJfzrdYMwIeeeptNY7i58PU/
wWFO2mnkfU9INtZdRl46i27THONWDTeZpbrYRvneanV4HL/kxq/v44ZEmfMV9wCxohPGuSTRiCEC
h96WrX6rXQrd5Gng9jLK3SfyvhReNM4Gu7q+qxQxnFm4jAtaT9xB7WH6WKlKS25h7qWL1AGDsmap
KjaIYUMa+4qFF2LuB5CVHaWs6pU0vORzuuLgjQD2hv2gslyyYK1TKVm1omlrjn/8dSqJOmjssZTJ
RxFizZagtqBJR4/9D1BZ6KkUNgbH4caltj7SIzFYD/5CECGjZ/FmKlYlTEjYXROUA6Tius6jiBgR
DjDY3NeR4fNgIWHRgUbYL1x1A5K9Is0rL5b2Xr2lCwB5AbpdWHzCjUemUIqKOGGneIkWOaZvFX3T
AZfdILmV2YRop6cXzJ/ZWT1lcOXTxHIwdQPdpgrkMCW4H/T1ry7+Yxvwpv8kYcNl7antMKSOGqJ5
VSzZzmC+i9rpN6bfURifld3fCpr1TxrBliH2xRBEKQcVeOxV++Ap1Gtr5U9CNFdmMTrGeCY3EqoX
8rA0KQluOnfeUGasskFXz9qMqyR3KdAztyVerMMei9DNeOfm42QFCylvc9Vv+UPwHmZeIXok2TaO
6u8Li7DTMuV3PH7cCfhBzX+uufDz1R8YkZ7xaYV9PwasciUTKHfyYUvpw+qUy+3TDYU8+37HAIGx
hDyQluSDW9Jh3fGJsgAaSKEruDY0waNabwawPspG5vjl9vAM5VsPJMVN+WeD0EE35bxjC5xOHLdW
56vcKPmZVEKrAQG+5Ni/104zwhsjoCa94TvjNN27MGY7qvxvdyZNizrqK2aajXNQjHzezXBTkOJH
cs8Jt0UUzphglVONeWBIJ0+niGf04XvHn5KIRNa4EX0L1klIrkYvdGAnskkAx3jN2Il5Pyfx1sDd
TIa2Ak29YiT83rfE1kgjGR5vPRyCtc6Bni+loIl7NfRwokAjLA83mMCV1KNEljmeThOwsiCNBGKF
7PYKUt1TiTL+IVrFHDq/e+tMOgr51lH1IbpLT/RaOQALYv8bmeD15y/1b64+paD6LWnc2iGfTw2O
XQZidyzOFnbuN0uavy0lxif/L95rtNfhF7uvmyXnYovF5zKaR3rewZDx3yfHnlpb+iDMJRcYvW/p
B/ZF722JhAgUKM5r3dsPkpmZn19+erPCiNFr1EjhO2vDXneDHQ6Z1AhjXcyTkLiNgv7y/ifOuIxy
nz8KSMjnCLCasFZdySEsmIHx+7pjjiH3KFPSV+osKpjtsCiHNvZgiGGA253NLqqwkgXo9RqPdbEY
oZrXAfCJE51ULO21iZurrLgpDg4DAa8x7nnJ3kyNVDVxdfz+VJKcN4/Zo7wsXDqJpBXP7ipK1ad7
iNaDtAhV8OdlOgy9L03sL5IB/Z3aOSvsDN/8DRxVAA+syCneHiLCJ9huJrr1n40ZGn8HSIjd0/Y1
GcyV/5BLbwaZ7MvUAShLhblcseMnmTrowZcPkS8RuAtB385xK8G3Zjt7bwcHdr4/1oNZDb58TaPO
OA7RhZHdTEIxSZYef1FEE5+CgafQlkbLzalTM4GOZPTRl+cczFjubwbOm8OIZkvqP0F+Y2DgTz4H
fXkcUxQVpspc711REaZJH0E9/Jb1F7aLMk3ECMJ5izmqJjq0xjcFPDYfoCAY0H6EnT5f3VPWetgN
j6STOZdKgimbFz32Mf60XPS4FFEY4FkkzVRUxFcz24SDI816FxCUTshYurAE6Ia6TYAMWXYD6AwC
4oxrjyI6sJa1tNbwMbl/ZKsyUhvhmgUUUkys8Nx+EYQGXyXw6Lp+qxhV1iPI0WrjJS4+zedgjkDP
4Mxa8+wVlAiLz85JSn02FipE5QGSZPrZBSl3lhjEi6prxJAl+JTmJJ0OpjmQL0/x0+/p8+GJHIsh
QYnYxmIHCKjxZFrqyGh6TclHmGDvyvUOfymPRD7gVw+xhlZ+AYKWLsZItlwwlshtJYof9zLTsFZA
f+jeMs+b2D8zRv/VhA5kW2E94t3z2iZURMgmbht4W7QXYqKuEj03EvxajVD1DZyZz9wj3rbYMDcL
3ObK9DaO0jHy8PhCb3HPVBx7+/wwVEEANvBrRFs2hIBu0nkJGS3BDT5c66FjEVBKl7zp+UCEUMkF
cuii2ma7AIEsc3Z4b2O3RDWpwebnzPrb4j8VYkwJgMi64iWITXN3/g7bkr23606G9mIX4QCMX6rm
LaXnrDcnaP86DcLhvaDteNJ1iOt/1Bika16zPJUpKse+SuXwo4KcYL7n8+pJj7o4a3NoSt/vlMBr
QIW3T0eStP2kX11VoCJzYqOqvUoLCPVPk2dCDu2M1HbGFGmutFIFze28SUQHDyN+f7A5Dtqp/3jx
m9QC2FpUTJ+LinCyG98LTa6XWa0hxqk53Mbjt9YKZkTGaTiTc52BOqbQct9rQ6a3msB3VHxa+ynT
nRomHe4hsz6Cf60fmnkxSyODA5OVgKllQadoWWuvNrZWhJHM74V29JBSlDgdLq4SX8OP2cN5q85Y
aROHCwU4LN79TgQCj7xLM71db44EYe6pgOYDOJcb1ZW0sOrqDuUb04MmtofcwU1a/vOmBoHH9pWW
uBczg1+93PTRV5aoURgAnWp+iMp5ZSTtmw27MxHPD7OV2yAzd/dfHVaLUtjdOLWrSziyOVIRdMVH
VmSs2UsbywyzsteJgwqCvdcckNpjtBeaL/akcbzsK49QuYWItOI8GGRtei4CsG4/an0waBhAHUzC
piuybWqqAcumV950TqVYDDQjGjwVnpGrLKJCORJBwlTwOh/+p+Xa1NbQ8Fqbj39lG2ukU1aO0wKw
ER7h8JYsxZ+cqQoAMtqeoisQCtPku88qG5t72tBI7RNQEMgtEJtClUd7F2Z4QRuvnGXyA6vL2rbM
ljWgWntY0wgmFctFzxCMhaLhr7RUTzeKKyT9kq15ua+UFAYpKomP3r2TX2K4aVVjRHxlY3VOqD+1
UBFNUPLoyjqFADR3uqumxaKr+2dBAgLw9KBExlaDPBFE1IseE2ehomG6Lc+isu+5n6sGgYwGf+pQ
VVu40DZBmJGyMAwBUbYm/Qj5jQbhpVISYqx3DswG3k8lQ9XjUtY2BN5O9utuOu2pHXBY1j46DTeJ
I5g3h8i1utydzi2BWihDPF9E9dnyYHNAG12Hb8OQsfzm6iTbW5pPEHa2e74d+jvKKWNNLfS6hovA
SWxImzvzr5BWM0RX9VCK1VnKijcT8/+JnAEmFkZU8kt/q7yIwC9U5Xvu4ARF6jzoITq7u8LHrKSW
SKXFSWK88uPBNfZxq5/8aR6GzOvNZCOvTWqVgvXwm5SeMC1nmYBUAgNm7GooSFxAd4Ifv+COQM17
SGnf/LHvxABBUrHiwy2FsWKsjrQAEOg8lxQXG+MuI3lC0tWc6cephatKg/uM8BLdxSn/THBmmiP+
Nsc1ipjw7YE4/X6NbIyDHzeA9oekTLzTLOncJRh47qTXpQdzeizsbaTHvne0167z8qvDdC89jCS0
EBIXhNP4lPbeW8J674Ew9xE+dfnWc7iqjh+fe2I3HOoYeqsErQFNG8fzftH2DLDPPHUs9fLY8Q0l
EthmzD4CDNXcwOancsv+7SIASW3WkSS8BNfFQuVMeM9Pu+OUyTNbUtbzu8qjHbpoLsodi+O0TvPB
M++vMSPXhv/XHFGaJCibcpbfDdL4ezPZ/mOaf2tQNRO7+uHf8qAhko5PSspKcfgDRaVrtOixOKAT
YPu1YnVcp178Ln0P8moq5ht1HnUF8Gxw6DlIO3/bPD8oG0nPT67Ejd91WmZtGMIisgfZVG9e32lT
gXoFXvJ0pNcwmH3T58albwu86+lJdQwv81A4Yume9Tsg7JuvYJUiZ4KJvWYWrL28ZYaRN5vCazXo
dQuyeOdKwoo3ceX2RYBl0gCZMepXZN8BgBlefdqPnypPx86Zi4KiIB/YAd184zmo5Wss68iH3NbQ
C/WMsqVcT1J5AXQZmWin9Wa912A13DIzHr5FJFiJRvJpENL3sqa3pZXV7PR28T2fjx4Xy++rMKFX
Ds3/CiYniSCqj6+Ecyqmup3hOOqkBSSSAHQ3uucKb4Zx5bqKvkHIKCGXupsrmDvs7OsTjOLa3xy/
EzFfp8U6PdIT5iMZpCftS6wcUkgxiDVVFcWCZCPpjoVVu0qZRUVuKqhYt3BHwFt4Ntbo3cGaAlOe
eWTnncmVh/yvluXk3LIhMZH7/zON6pDkTPUodPQWi5P7Prk8vOGtmNMPDheq0/WnXK4X5lE2BQ0v
9QEmNpkR0YvmOkhk60b0Nnl7f7THgCVuhtzOM4QOr96G+2dfYjBlPOZryKWzTZ6g+ShCNX/7RDZB
lECD6r2f9rpVsAv/hi5oV/+ss/LxjfEwZnShgpxSMJIw1zuei90s7CYDAxPSa3KFr58zJtKMlpYI
V1W+rcLKe80kaPKLnzpWl5BxJGQx3DaCdfNdQGSK0U4S30ToDMcqfUOskfg7QUyAdvaO94KX9J5R
voDHvu4NExv3eLkj57OhzRbtPEvl0Vyx9Qwgkg0nvDvkuslSvq4KyYZ7mbAbK65a1qi/jHchTG6u
FiT70sXcV5nR536I+QyCqoOzyOw/c5HX0cMaNPD57kEGDVhNWQ0jrnTH8SvSHkedGKaM0Q7U6Cga
0UQSynOWprv/Tsg8n95REfwW6wVXnUH5DjnMZe7yndRqWmGELO6/6HIxm6FPSmUQsCm4ES0I6Ab6
ziJFxvktp+6RttETYZQN4LVtZpxDlkVmOlGjK8PdN9hQNKb4xr64lWG1pLBc2E4dJsBsRCBhbe0u
sun9stlnmysXd90J3RkJT1GtQpwLK/9wfCm5Tys0UlELl7oQot343932g8U2LWwvPiRKq7LYu1N3
bskab2ibcl7KSxPsog5TJCUBBAYHNCubn/5YC4gu7lfxowt5SrKRpOrwUqY4GqeeBTps069WYGSB
zlBTB5uPjHCw0aEJeQpY64RqQhgt3zSZRQqY/aebh0tRm23+iA8R6Tf5/DYFSaeaJyHGphKGW/Kv
7wVnO9CC+4XCVXcDmiY3Idq2/A3QYBTxB7OaVf9NwS80bGf9of+1GYu0XVCatUfuay2G+/M/vdFk
PMbbfa9UJNxWjBAn+KyieSRhsl4PqNFwTjsVS/JKqxFrMlUTu7AfYcV1SYHoeZmk41ExSyiYMixu
7sijRxxpGhAxXkvdmIhtd6Zc/khvE6b2lnNwedQaOqxGvaCX+YQHDeSZQFjVja28ONGcGWxBn+1B
lM8BmrkJ93xqg1/AkOD+SyogOx40/6FoKVWUlnRTNPJSEd5SuoMe9GMxYxSr/ouCoDnJrRs/g2qF
MkgFOa2RHfzx3powVD9Fi2xzuC+zY4pLFIcDZNe7AHNGjGhlND+ORcjt79Xk7XY2uMT3/exaTiNw
MWmO7b83zMGzZOqB6YDfnVj+6usyQqKa7y0TkR7BUQMsEjYF/sboiOu9jqGNU06SoWhcDRJKPTgQ
djV7F0Dm/XaA/GkwAz79yLjurz7alrP+6hwhG4y2KX2NsS7for2k3NG3NPap/8Rz/FeInq/WhuA6
SI+zkrvofGfHXKsuqPE2egGSy/yz8Tp9vlZmlRSt/8nNVHHQ8TE0YvV7aTe+f9ZD2kduvd5v9gJ4
R+z/yY8jDBTx9oWu5zsoWADQcQihCgAxnnycoWcqls5j6XXAZrzOKBx/HhvmUsMTmwwff0RBjxcu
HXA/I3bxWtQC7Hq/c1BDoTOM8i8+kp5hVN979lFutN8BH0osR7/tf1nIIXIbgV0z1tHqcHCCk9gS
xYiBQ0zf75DF2J3a0aoWg5Lbsp6A/pYqvhVJEMahS8H1cQT9FUcxQSb0C9MfMZdURMZ1hAMbrC+Z
W0yqS7LaYSES7z9MuO4idT7a0ZYqHiSLUV2J9a/NhqHU+jLecliHzTAk+1we0FQGXJv/FJyWDe4w
ZNeh1wMYVW80G1hqxrveAVIoFY/hb2YDY+NGLSKFCbGEdQyGmvtBcmZacQIMWp2bcEGPaECv5owP
Pdrwp+hz2T4YDt1Dj4mHa4A9T+5ZNlo4qhLTTZ8DO+ZA+VBMiIVW3KfQ2KPOX/Xnq23Vb8NfWWAP
QfwYlibStlMRYrT2W3UGnizzuHYf1+mLVduDS6SKa8OpT7Pvw2rwypNxSZcCOP8ZY7ZLNH/L2GAU
hlSgdKKFqgyAnvhksDJaPExAFS0FEGERBrt8w7cThXvqCLYIBwMXisAsAWQBqGpGEYuVuz9LrfYY
W+aQoNoZWNyV5sLQWOiPTmfvLv5umch7yN4PsgboW70jKtMMs5jzyhE33MLno/0eeKE9kMz5y7U5
j7IJcUWpQctIMnZhL8urktZ0hrS2FotcqY6UlSYptVGHtPAK/2CCmC1aGScLhIZLHj+a6O7H91wT
DZ6+oUBMiey0p/tb3Xdd5OVRnzMC425vfEK0C6SR4g6L5tU4lO7LXaz2NlxFX4jYIGjCNPNuCGYL
OVCfaaDPzfudD54hhJRqyukcvDUdmGHXZX938g+yE/g5d65oWOGGFyDVQYcvk1Ej1vWT7lMbfXkR
jKpOiNCf4azuBUf94jUqCD2A83CTLMGCn6my7Ihy4zg6XDAOtP0qf2XWBEdLBc/41BXKnmt6lNFr
XNXB/NbbB1jlSRyov+LVehixowW4E6jvnQs/A2hGsFW7V7Y8nBFLPQjuyonvKco8Dls5msRXaCnZ
JPr+OCCWWMdg8ixFguBrtQlwZuP4uBQSRxULhC4WbSeyB8dCxcJzqJqSVBwqRV78gQIz2RaAH9sv
whkcH8cOMkHeEILPWOl9sn+zgCstn0aPcMz0BralSbMM0xT+zDPmKl3iIVhsijo6Um+JWqz08h96
VUSzZRFVN+ZVpiS2cLCdy97y/oPrtbxadgpCjoOYGyesEp9IaAwzbWG+lPtnjkG3UUGYDctsA4OZ
wwWDXXIKK/59m9qe2R10Pj9YcAUip308JEKhAnsoN3YRRqyXFaxyfByvMV+i/P9siim+uBD8pd+Q
qshDGEftokiy+VueQ6cduzfm/OxguVxkbVtAPUoTG5eBsrKewjIfyRQVoqvLSTV1I2jFWVzJBPNv
SUpp9WBxINm+2y2ys70WEk1qTh12XaPt6WhK/MhYQRCenmucfAzBYwAMrRYA180jDhPrcmFQq/Tf
SWe0nxyqnQMlKpAWpqdVe03cW/Y+NQF2FC+8rdRpGHy2aIlFEDituG7oxCsK8/0N94Md7/A8wKM3
+/axCOeRqoDkRvHpZj1hH8GjkRdh1r5IgBXKrKWvhT3usdSy0BN30BE7/wf7c3fGqgAwmNOkjvzT
M7ggm39R1CIkvifRwO6u+oOq4jBwt5eTagte1owkAxzjsvdDynwhCTd/wIERa4FbsUP1zM8mR7HX
NkgR8kSws7y3BXS5o2kqt1/90ow4Zow9evFWKkF2bu3/NeBzykRhfZOmWRE2YOIPYqtzn5UEO7hI
TWCRH41qk1pkqL5sWmOPhj3pYYqQyiSpas9ZoyRGBdaZVOS7AXHGlgmkqLxueuwronXsq3S97VxI
7rKsmeaHt7bQBG9rWTMbMvScB2W5lHHYdBhLp1QYjue9Dh7kug8eubN0QaC0iz7xrc8EuZES7wpS
DcP3/fMqx8QGUbSVjcBDvvvOorASodbPAkdpKw9PCnoqfkrmIYzqVxEv3v4isyIvPC6VuRBGxqvU
uL4yBy5TL7jxks0GgqtpI3UYWkAhIWJqrAZTrw8NTRUHkSdSrUQ5vI3JtPq4Pay3BSL6xyO1tVu/
A9h3PDjyxR8+tsQ2I3Y7LlWFz5kOnS0aqcPTNP9YXKjYK4DhiQMqWMbj272Plb9O0mson5GQj1ak
tdb71FL0FNgCNXNTZU+hcKMC5Mhc3p5sKRPiWN7IBrQd29q8SM8Oh+QCuZNfQnp5Csd3I7i8REhz
x/ycWPNiaZiE57ZV7PSkESy917J6NJwvWBTjgUsQ2woQDhlFrT9PQanoaz0YPCW8ahs6/Yfg/rXF
K+8TyrYZxw2LxUseYZ49RXCek40PoDBrUZKIRPvAIXLE+UD4dO784A9/nxLbXWkaBh/B8kGUMJPw
UArVOAOY7WX/Cgmzw7zVs4ki/rywJ7Rwi/J5AnJFT1Y8CHi9lghEvApQurwJ0HaDLuJ2RUjUAh7r
+yCK2rR4OTsujFvuOGkd0NeblnSmHm/jKTn4gn2cmseDE2zNtz2ywHExkOAAU57x46RZSzF9l07s
7YLfNnnbPmFJZKI5QK37hKEriV2QLzvYU6kPt2/EVVAzR8cI9PWva50le0BBCebfmsUSDZkmCjOP
K+CLyHCpXeJIHpk+7xg4YrSI08ZzlIueY17o0TjtNiF7K2UmY8kU4h3tHTBZit262H5NlnZMLEvc
8jbSX6CH74SyNSWOmgI7gGvUGt0ufx1qDdeNJOtIWgBw0bxvsqSJEfNtaErQLnuRMUJBoUKpIfYc
muI2D7Kqr9V9wdkp8F1cHBMdW7J2E/mjJ6lSMn4n16ma8vbyewRudu1u5wHn/XhEk60+oouHdIo1
5RGCMKlY1IH6zxyMwwrbEv0Cx0H9QI9yWVEXBDSFmxkONOvX3DU5jzNLdTAZpDtjRIzyXL+XqGZ3
IcHsjGKM7/nxzPUJzzh2GgZc8pvy3CPJWDnkRwVMi1FoH0F2ocLBaHUSvFSNr2H6bHskcH6bbq9t
1VwN/ojgvisoMy7Ca2IzMbAJCP2dhChJHwaU4W2tPJuWkEBxQxH6Wvmjn7qMO54R7U22Qd2R6tbB
Su8MTCnc3vU5wO1WADLkT2xNJbSNj/RCrRWgQBvmuUf8h0Mc7wXBQ09lyRZSzEv8z/QHn/f4Zsrd
6MkQLP/CfgxJiKh4le+ELz8nkPtp0ahpQ+iJagBm8QVJfBlXy+UYo+Id0myCaIBllX23OOK1YOgP
wU8Q8ion++9DAV9MGVv667N1tVnGMsoucBdmcd5O7MlkZF8MYHa9XS8BJULTVcu/dRWN0ngg7onm
YPE8/A6uZoUauEdYRKrTrTMPZh5+qA59noH78IBWEsDmlmcxkJIoJ+pNRqIEC690L3KG9DY40eak
sJ62Ak0SJQ5H3lHaFA9cFHdp1ni94+MyMOanll3tN7HnjgJ3kYBUuSmXErdC5x2tChrvGL+g9D6B
vjtjhUW+sNvvtpAYpfOV5pXO71enYlEg69WdojxOITMntkMi/0rL6gHWj8OUy7dkf4sXuI0WEtYL
kAshSTMOa2B+ZAClP+P41jdb0P1/HXDgajc7jOtx7DSsbXzgN/4zeagJvyjKbqOdQ/MS8a+8JQlv
rjzWIRq7ExbnO0TQb8Fhe36LJd/5KS7hLflaaS2TbnC8f5kBDbmPxpqoY+y6QHmzeqyuAKlv/x1B
+2GFnVgEdB2R9NlgDK/ryCdmOOXq6Y/R4W1mvJ7vjytfqzCdyV7KNOUJHFhVuuO9fnoTlGRu3RT8
wYIesqrAqnvg4lUN8bIM9zO2u41UrhHxlZpYpq8Olhhb4OQ//ovSrHIIGlOz6LCi6NSC2S8fvoQ1
p4t8V9R5uC5kNUXOjfEfqC3CF4aJihMS/3fmk8swboARZbHRZ12srG1VGlpsXF2RwK71ACkWiG4E
5+9HJo21yXADhb8UIY6BOQWuG+0J2Tsf4gzqH4VSj71DjsgG+YI3Hmqmq/RHDkBKT/O8cg/WiOOr
/qcrT+z7Zu/sydL2aHLqjYRwAK8ejnIp2I8ss9nwyh6P85980WfoT75nsX75JKOAbdCZEd90Y9Bu
xVLNoP/vT8NXhguipgYOZvraEgfJl4Mx/wNg9qC8rFgKyrfe2CsxEwZYCG+Alz+uZHncTPIpmD1f
W6sQWBFfEE7szzfQ8YLQcGTO1yXCoAJOg1Q0LnKTboT7gf3H2gkbUTu5+SzzqgGyMzoma+pdNj/5
4RgxOJh5fEiwp71S3hLUUGj9ey4Y4GgU9Fi7oZO7iQuI12V7uEZ6nU3BTWwTymBEUwZKtx+yTGVA
eatqOrtnTqa4t6xiyU5IWgNxmycSUhmDsIlE9I4Bi42cEf+hYoEkk9O08eTlWl2w+HRNfFWSKWhI
kJ7Ko0j5/TQsiMIH9R83mLq/OyDBP6nnPYAiRQFT9h6nhV3vuJ6wvTZd7otRoW+j85OcAd564pMC
uLYr7Rb77qQr1l8YfK1taYWt9vIYeOrYa9RW9Fhr49K7mJ0cRO06PjYWXmigpaiqFBoPZlOMtUez
S5Qp7hCPcn1Cs0e/MnNitj0i3TFWWCy+0fSVK21RLRLp78xjUupZYFAPxapfFALJR4D97mKrHvNb
AayhOkKO/MqFumnVx25NP/g32e3ZKXWArXBOX4rCTTD+TCLssR17nrsZl14JoXK2+RiLCUffmmhx
Clv8vr/Zta5BRnGsm23cw0E3H34g+/xCsxsvO2PPHcRiWMKc8bV8jHJhMEb4IF3hCRWL/r1d11ca
8c436xUgVK6+XWd48MbboQiyuM2jlg5AfoW+GSeHJjE60bbc1ml77sWtktkjg2FTdMgMX/hYCvzg
GBkpJaFKYhozTot2Zc8yRSsFW2B+iLJK1kOEPhLvaFlwApi25JnIdHPE4lrlwkBZvjcjWKvHc1pV
OiKoLx9HrBtks6jV23L/+cs+ae/CYzsTBrB5VxE6fw4YMJCVrNJJum6CcJjKAHWswen/YAzltOih
9Eased1nn/mQ0F3WnBRZXE1/P9aPP8AZVWb2BcLEuTHe1UmUH17repD/coghMlYSTjVZnDaGvf+o
Ew+PZSK3iov09HOqnCyNhebRQL+kepNr6fwDco0i9QGEDWWnk3WxIOYrY6TOSruCCWAJt8EKUJbp
YmADPo8E/5NJsAJVAsuhGycGPf22kO/VLOGRTyGA0fxlLOnqo5L9xa43qYVqYuHbw6aGnJbsbYUl
0dxHt6YspX4jM0xm8/eCF76XY4PJza35uQxJOF8mZVn+7p5adP/ukU7w23TuAmAPoo9bHsJ40uTd
Z8Sc2/mPQ00mRQt/4muScnAARcMHe17ivInx1wrouwg1xc/TaaYVTzaZ6BbzTfOzwnCJOr5MTHIb
LkJVYCr6uJADEo8wKJWPPooROWbYb1izAgi/NeAATJZ/Cpiv7w81HwXr+EpWA/c9z2rvq3dGKQYq
LJ0804kQB1NtqmvH0JSTQOtvL23XVRbKHpoOSRZGkHnR0w42Bel2Ul8DI1EuGoHl8Nr48sM/dahQ
XI8g+BcPBgUwFlf12JmIW8NLgnVFgr8gYteW4FCVF1QY/tZlpWhXfqU1Fn6gF86a8J7sqlXRIEz0
sXcX8ur6ARICERYPpd4rQ0dTPDE84zN6rJQu1xs+0A/WGNtmbe9DJflCXrw/Z4ezbKZvrq+IoI6X
mHL4cwRfxkbZLfA64U5PXe0Q+fRXZpFoGdQuyDqmi80gzC/meo2J9FI/K2dBI4yhTGWUcha4HY1F
zRpPNzmHNg6MvzX2psbGKI0HcxOsD2OD6bXeeX3J09RUWESJCOsRcafCrrDIlTykGoeYPhpRrPNh
us0H2zf5j2R6PcJQReLbqMpd0v0rSw5tcVHiTlzS3KMPC8t5mBO+R7JDu8MMev1DxzngO9av8/ZD
0WL5aYeQAyGFIFrCLy6TMDjq+uJ5OePk2ssMnOxycHrchSo2RORpUViXWcOk/NW1RLg0Lc4rZb0H
V0H4tQq+VYKPWf7yFT9OysiQlRyNuV22aPBLdS5siKRjph2rqs3HqyMc8tJavGRNU+Tkhr/uWJNh
cDw38KLlq6aNWFRZmYW98ow80M4lBvaVRxAIPix9abxBaca8p/54aGeYKfKC9UltPKHMKfbxKXoU
cFQqcyelfQ8GCVihOlah5bVYJ62zSU7vzcsSaMek7iyjBrp0Rm7tK22JMAVGaUkQfG9oTlGtvOcz
Yp63uAcTAa1Q+GUT6MqngjiuqhQ0X1lelx0iKIHq4Xm++zv1eOMdsDhH8CCNScI69fPQV7WtUIJl
pOYDUMSyO8tgDhw00QAy6/FUZUgvhtZi9WabiPaeLNucuHOSqFqLTQmNGxFAHYnwbzAum6JsbFN2
cnv07j5NkD59gqGrg0o28r3GDp8qtBE/sKuVWqrj8PyPaINA5vFTTD/chqLP/uaBK9/veCb3eln9
7zLFyChjNPUwvHAW+DkDITDB/V0WKZarrlbc3leacyvHcbC35zPT4yTlvtl7syfg04SfJ3hTOOKb
R+mmy4Azhzstw7RSxPfWAk+FkCxk5km5cLPP0dVZZzmWfxKIUNefZa6seaSsHSGL19WTcr7qBov3
cffjGiGhuUdxFe02C+DJh8K5EzcMoQCw2ScXuigiwGEzIwj1vPn3uYmiMRkq+VldjTPTsrlGNTc4
sAt4LtDQCkXm6ifbShNPfXltI/qsQ8DqmGhMOJSvOpBgJQ+mXG4lEkk7W/wfvTEJaVgapm9n4taY
la9tO6HYv2/KbifvXRafoZ9xvrU8MDSl54VDSNrXjOVlQiASvcU9eCvM/ZC0Y+JD857Wd1Dy9wjW
dPfNfW/GZO2CDQ4pvJEy1EML8c7nza81aF78GSoQzJSIIlJhgaTaeKSngVb9iLy1IWbMIoRoQcMj
vyFkdJUQKGM6zSOAnpBLQveWtkL/qhADlHEcpyl525pcPH7Ii9pqEziqL9TxKdWCDqeVsWsGIqEt
7a0qqpGJro+bZ+PtmBU205ppqV8g2Ce6XsZXeWBjpZ8DxMnmOfK5wmDWU/e0Acl4fjWcNVAjHCRp
lJ3AFqbIwYZZSk/Ya4NL3W50GaeMfsfjTtE2e00t25bJ+NIj6y7O4VI6D2Ewl4gXFeNIO/FnNfCD
3JtaPz8+nKC1EH4hhcJKzfx9eQRDyTdCnIuvjYVk5KD6zZo7zzYKA3M05wuVrp+C+LMLX7dG/nOW
rJddSj1D4r8N/1rbuKdxRlNP0B4OzHKSntSlyN1bhL1NH/b52C2LSCfeHVDgt0oOiPR7kCWcm0mG
ogN8GMWytgYe65visAM9xG1b0lUqyy08R7D/SE8pM4BQP0y9zvyYKmxKWSy5+lXEEB12ospCfIgU
VgmKDUso6/69w5GsGLqVjQPbmF87rym9Fmswnt2wE2Wm+TVAHQgpTnwI8Obn8Tu+BecQcrFEiUgs
tuk/W0PtdgxSST2Z0K8y0iejnWM+l5zsxbk/xCVwnarjxdc4bC2TX6JpCobvVLTnqkS8PD1bl7Vu
QbBc+/G5+XaClb3WNEqMJsNm8mKksazT2n+5hHlctv90yNpp97eR9JoN9w4UqIbARL0vnis6eeFw
Uw+AFk5Yp8oTMeQlYCq0bI5XOMr0UnB3UTBaBocnGV51swF9Au0PDc1wEfo55AJN4kRe4r9wfks9
G3blHQZP5kJWBxf3xb0FGsNnINYgIr/145dgs04mBrgAx5dtYaMk7lGZtEAoPqND+pDPdFUXBmNn
KZhG+H7TQN3ozfnxXHgywDkE7e4a08FDGhUpVoiuQain2MgGMgeMAF+3/7bW9rskVLOBlMbuV0ef
+8ceKR88b8wQMEZlGdAGI/bBtpbrftgnFpUZ402TgBtqHsNroq3y+gqR4DzIHSXczS5KNmAYVMhy
YXMKxwwqMnGK2WzqSijhWskn9m9Hm6Tk1CdYu/wOD6GIjY4eFnxZFmmDv2DE7onXJ1xySvsgPH/b
OM16W0jL/K0NBENTIB1gn/0wxZ8112IB0BVD2eVytpdcF3ws5jR4iEqyANdIB912Ig06XWzM7Myx
v/NMqF8fMmEiYKZS5xJBN0M+CJ2izmpFOC7fsrWxhbJhU8jVUaORztsYFamNFvkJYjSQhu5zGYOQ
w1X8pjbS81vgZ3aSCHdg0ETotXIvwXwmkXQkLE1ju4GvOSOPULMl8QwKOcGxVO3Wd0C4MQxNrSMv
tTSi+OSxouBZzGeqNf05CzGBqMBYjxt43IOpzStGMzegXYaSYV7fAzEDAy8z4Jsk//pexx3Rkflb
e1VLLA/HIz5w1aqbvVcLy5qgMTHdlwxJHSW7cn7aPP/IuryL9y7tv7bKZyf44ea03BdzLS1ZmEK/
EItsocPkqQwHYGNht1JrVMCzDWXIn9rqbTiwSBpUHvVCb40REyBhwMxDH0R5ogcVqv0Ie3crUstE
ijUju3YTQJQ8pTQRlXP7RpXsS7pAKINbX99eMVKVgQtKRuSXCyDtnjqD9bi9f0a6pUTvAIAuVgHY
Uzxxypy0eS8JE6rySD3oex3LK4jSyZWFn1RHjGqwdesnKWU8Tn8q9QraVgedtyiHIN6TsyuB1Zkm
DQepRicfP1N+8di/ZOFULgKWDb668z3B6kaZyeVxc+vIHJJWfaTwZtbDXIKOs6ZKZkS0TltCUMO9
jsx5H1wk1otSmej2x6zeuq31sZkqc6jgOZR9peusUCl1fIIx6+fseElnHcDs3Wxt+/GF885ZlBqB
Vzi1F+VUSCk2unaKVucgEHAt66zqsQ4y60ICiYhdhlJvw2OOwDOmHoMbctrXKZBC8wFBCBBgX8Mc
lGtosCE6jW0Lk0I78tntClvG9r1wtODFFcN4Tf5DK3PahYF3AZ6wJR1xtsk3+5jeUVWK/d5lzgoS
IMfEq3WmISoJFtpfI0hu6gr39oy8lhRB8mqv9fg2PhSUR1+SO9jRu6AUpGUWQ5ZF2sbDy8ZLBR21
jS/mRlxNI0Jeov2MMIZlSNXeOhsU6bC/lj3/emuLDrW4H2Bj370PaGT5bHdf0xSH4nUTMtPlK5QN
WRVUat3gVxq69ToUpodRn7AtnLHKG7aT9Evlyx8Sq48MtGigMhRFqFuOz4FzcEaYyV4zlGSFfZOJ
6uPqiT5pMgfZi1g2ST0RE7BdA3XKD12JIAgCcqGROlNjx+VaTh7F0I+8R2KL/tBmib4jDlhZIeQc
8A2xzXjqC3jtsM4TqWc9MdwhucIPntv+Bb1/O5wl/0YYUylpqK7x6NUJovibK+rTB1D2Ml317r5T
/JJU3rRiY6XFnxX4hAJXCnSWICOAZsksOHlsKn4uog1BDv4wCJpo62/rGPNZl7wCs0PijUnp3p3D
zwbHSGwNCgM6oXn4BOxSjdE31gnEMDi8FnE4WQIuf/X5XooUtdgdbdn0lnJZn26PQnIy3r5e7Wuk
WEmttbEzoEiefmkWcnO+dmQFEf012N0HDSKLayC4Jw8M4SMd56C2vhdHtKdMbIxk4MNxwwsLvF6G
rbrU3t/rixgxVcnb46il30hzgidPn05nliN5lwRbKjX/4169A/s81i7uL0lvZyK5Q3tdnHddgS6L
UtVCRjl7aR7979sSYYIbRuB7dOA/of7ePhZwaHK7d6S1dPLKCH2P9Mcmpf3Wl3XdWvNs/eiqxUGL
hobYIN+SuICDd68VmN0JJpkXCY9hUVK6iqbDFnfVv0KzYAxhxyETvvm0kbRXlrLguA2pX/LUmMSZ
6GSCrkHfL3Fw+nCqLmtoN063gsYg5fsOTzdOgX/xjm9lv/lxFI+ZeIW4Yh/hGMu5AacAywSBpkgv
0gjKa4FjtlKroMUOTmoZPmxA1CjJQkEx3o7AC4/vUpoC271LIPthf1DY+oJtXBej24RVET0s7Osv
/TrZC3NjIlFM6JM888IP3PrL2+X9GZ3rOOQOtnyE+wzLsLZPRA0fag/d2Qw+LuvT7ypGY0nClxLD
jHdOmyaRMG4oBwEt1+DXyUII1C0pcn9j68zxtH29LIZfNVycaAMd7fuDGusbPuKZ1zTxrAb6kAjE
vf1N5Ale0ni+U6K7vRy2+lx1UXAgWyVHbntmvDiQGdh/lgtOknrlE4AG1M7O+rYZZaAOw/2p1don
CB3hTmstbzMeYigBdgQN98hS4JzcTHmgQAYUKP+YXTZ6zuQJBAiql9anKUyu3YPj8sCBPfNKUDHk
I0dQY+KlYnK3EC/IlAlT6rThlyeBPOjQGCQZHmAtFKGXd4uA+FXcN5FYLGhM/nx2kwnZECIaH6tk
W0PTLkyUtOT5rd6U+sXRHeN9y6WjJgcOTbWDuH//RkxOe/WiNL315Kn3mTgC8/ZfkamcDZ8xB9KD
Eacm01KaZu8yxYI+qxvRT7XMTD8YhK6M4CncCg+h/A3+jRF2MJIhZZw/GRYBovMdS7duxEAR8LJe
hGN8BBMj+GyTF9soVZzuH3hek991Hl16P+JmNneHt8/3bJggp0shWLnpu/RzYyiQr6y61d/NohIc
7Sv5uqzmE2IZyTUVwxHqQPDvc+1fvv9Kwluv1YHJkK9Usfv/NVrrvO8Z0e2PuVOMYssEgpr6d3hQ
kZ+QoHZv9L2cZhIKFFhc6DRMl3quoflOaXKJc4EQRVsipslo9NVfeb7Wd8+5nPocSqxob0bJp0Sw
7/Ws5oUyNqiLZtasQFiFJdUoD4Mvc0xCXQZSGfqQ8kkc3b1ovRIbB46c19avOieA2bQ+nYgW1Z++
AJiOnDKsx/IN+peLh7ZqQUzTerAtL6u+5YoZ1f81dBfguXOd579thKxb2Faspqw9qZts+Q6JnTgK
B3nlIrWuIIRN0iTwP1pQgTS0TbMVQWP4yn8W0X9CUht1Xsk6hhfTfmYATrpE2DWmvhTv6jOOyeiz
w/sEfJ92lkXbXVtEyjYGsTl0b5ex0dZHoOA5jg29krz5BcFnhWC2PXEySC/yPDsRQK6sPW/JP7fa
+/CVTQtA48YzU0ebzjcA+6UVA1Y9+GuWJowReSUpATUJ0zFrz6ZxEN18pt+qQtX4vPTlMMk1ic8u
oQi84QsgEr5j5dh6aBF+Yt3MvniZvaiEylgSG9+00EnJJ43naff67cwP6qT3ysC3HIFAGpo+uaMl
BgglXJdg60ayuMTsFJzNE9u9GEQ97F6saLxWIIalttM5ZplHV1KrNaPmY6mxODJYKQ+CJuSOOtdY
r4NC6qLUsTWpX47dXPkvgnX8a7H+KErdzkKyD15OxrYuJkUyayRzbZVD5uHT3GRYw1Sbxk43HURR
1txlZzPQoSHvVKLJaWAS2tDHdwDU4CGNUU/HjMHzL5gqt4Yd0A2PODjcY0Kjq61V56ozrQcPwNks
1gHzC86j4BVT2heSoOqQ2JMddW+T3G9rI7g4QUZ2Mok3o381pVSJ4+LfbXSpSkO11drxNFH1kl4d
O59ezx2Uu6yozPk0dZ87NSicQVIk1uzInckwIXMaGA64+BHrtzgq2eLPSKnEz8V6RKkFsEr1vHyd
TSGnowv8X+kjWH+CQv2Hb9eJBYOulhtdJ0HfbjQWgETBcipH9k9aCauM8XgcwwOEWuWZxUj+5nSS
wKpm3O8FVITa3hDbH6/Oigm9HX8ADetVJdhzEYBwW5JFfDQb6EDLMQXAyWycAmDrc6DsDKzwmjbV
0I5fuLp4A10YEvYWqHM3TUFJ0pQ9qmPOyGUJpkpUklq0Y6mSo6Wk1OO31Zq4W/4mXymS9Oj/DgSl
Q4u+3+ckp1hOWuOjHO9wP9XovYjN4iHoojf0K0um//zZcvzq+ukJpYM6whF3LanclD/9Uef8eHKs
hQaTDmLSzvEh9d5k56whUOA6wSL2bKJy7Sug13/LGHjj0IBpbCdYe5tV2R6/RKlU3dVB9JKqL1d8
iZwukbqN0MCuERY26GWIAm8B+oux3ZxQP7NDSpFnYloc5ZYCQDQySpTgHTDvipg3H46c6r5vlYq9
dqEs/2CL4C/feS8RmsTp5ot7dRP3BEn/R6+7qOS6LJSVxfLyAqfRNfyJ5Tq6vSUmAwnc6BoKsyXi
bGLk+ok0LJ+E7rfqioGoNxuYiifiIdIi0IrB0tE+Qqo7Pu3QovoFGlmSEb5V1WmFhiKlDVnpKC0S
0z/IHENhfW9BRT5pWMql5lGTr8lejJNTljNKo7je+Aw7nGQbfU8QFuRgcNbXjzqNQVoe2nDvZaTC
8vysQzNNQJmtEIpZ5GXGWew6gaNzHGdmIe3TzBRhuCxHEijiuuFGpdPApwuPIegKhNuo+I43V4Pw
ayLi6JhrCfnOa8mMGCGapc23fW74ZMsfr4g++ddyUK5BK9MeTYHGRoPbcFI6GuRlTuo+Qbc/a4VN
8CFjMlXRStpyefAA4CJmm2hk3QpsPEwlJ3Y/nzkAYLDmIdOJI2aN+21Xu86bJW9yHqpruDC/qyHv
VDQLjhNIONXE3wwfht0AY+uTQKw/ZEDG7rJBuMzvlywMbW3FpkaY8DbyUhC2LqWPDcBda7rUcaHB
+WestbRRnAQPR5fw3fKbFfl9iztUKbInbWH/7CTJ9XumMnlSp25CWR2eF+MZTb0FBPhx8t50tTcp
Y1UwGohPePTReOiitS9IU9rPbPnKNogAZsN8x/Hezzfmb+MeBTHwHUs8F+YNbikio6WDyJEzecBb
b2q3cCofbr2MuljI7LMbj5i9/UKa2ckjYL6oIIN0GLF6M/rkUJPsRG3BY7EgGCgpyDkGQps5elyu
WnHmySVk76lCD2WU2HRtvDUcw4LqXk+tzn8wCiXpSI+/REVB36tDIU6HdBuHpMDqoYsVLxFi7Zeu
B8PoKsZRW4kBD0mf3k8AnSvQjNR+xOrkHWaILD2BWuEjBwk2kb6WoT54abVxZWYCo1/WOXb7tJF4
IYCkwQNvPNE1anhxApze0MsudMpqT4PJJYQI4tg7zHTs0P1nKo1dEi+Yj+k6rp7QraI6MTud4hTe
hnOSZA+BbP3YOdSF84T8OHsPVttGVtH66jXrL/bN2/Cch9QFWrX/UoT8oykvXBRr2gThrOw4lr1M
HuGsGmpmC/tu7ogcQsV3PP7DJeSvc5tG+NYL6M1TLC7p7L1w/l5Z5hsNXkSKex7k4p5Nv24uXLyw
gRihXkNM2bz5cNCgJpeFBmZhPYEqmoniMO/ogd8t31tZbZMfk77ZM94RehBdG9s+eB4ngJpshyNi
KSqKeHQhGyOhiywYnlz5T3MgKxRhgWltuYPfIWmF++dtTtAa4b03KyA9cqlXduCZDe1MIKReZ3Hp
//YlD07d0XTCCtItOB+PghRfh+T79PV6sgywalkn9SR15KYZIpnX0bA1Kn96TDEmlNSQSaPKArkH
PVgxSwqUztJ8JdB87xTZ/lP9cIcXWCPGbhs/HxuhO9C9Q9sdzogmGhfRpc7KD/OCawoZpNVpJtHi
HoKcsvq9UPUfxghtsdAGvFZnu6MOHapNhVStWpjrSSqCNFN9+GlEfWxqqhCsVZgnDF1g9giqAHkY
LIihgQTGzlt1P+P86xhyYCZr8od/3L7qTCrpjwpnG0OnfOCS6ZjImgSIiBzG5Jipx8qYWs1Ww4Ck
KX8mNkkXCuOkUjlyQ0PAKERM9NQrlnAagWHdWb0LT+hCywYSwB6a3AKxw+ThBfj6ppI2z4TUtDLJ
L/w5N2Nu2CCi/PsGGH1+/TGqhAJpeflI/KWmVppVz9yRhT0lU/Q2184kIRhnHVVsZjq5dW2/k8+7
pTswRxGYoNUjXaDNyZ6mVsZaQ0D5iCj+12Tea3TmBxZcdpYPDd5ueUcyAUgdMUA49oRsyIvykDBA
Y+HjrTyypExNWf3TMPsNYLIdfBo4Do3bRZqrYRF2yucpyrJrRoDFcMaZbUjb62e1UbZ8i5hmH/ia
/3gnQyDbZmqZqIb3GV2S11WPBxWnW+42vUxFiS1HDt0jLHLKLzghOPkwQIAdnxMR0bMHLTO5OVr3
WuDTDPwjoh1z+09aj0zk54JPwPsnd6QJrZP4yGdMe9wqSNcC4/ARecQEs5z/TALUoStzT27gXwmx
yaggoP/5hkP/jf2FzPOCcr0j/zMHBsaE+izERX3qlz79L/uOXfdJmOBx11mUt93rZPor7i6F+5XC
Rr6WWev2WfGsrAFWQivc+aOrNOt78zW053HlDt4vD80aOXAnjnechG54SDPKvZRY05f276t6Jfbf
4y1jyqvZNybKJ4pN/6jRtiJS3X7PfJLE3r+MMnjImesPpdCmQ0LB62S4bsWJ6PBc+B4OVzd3V3Go
+bxKJgVU7s/t4f1nVbTKp9lxoDG1Rq2G994G2jZOkQjfIMoPlPmBbOS9axy8kcNCnVvjbJ2yaTnA
2aIm5K9JTueVk0Q7h8g5Yf5l6cuLSJaa1g0fd+kcw7JQrA0MpC4k8U12X1/5DI2yHYriLPGjSnET
23Y0IIfi+C+Wu6M/2cYUGGN0AP5s0JUrkh1etbrwZHgtRLpvVyqYPud6ob9ZdB9132xTslobUUs1
ySIopxBFA9N9x9923y8aoOjm33c4sO5Gu4tGRSbHGVZSZ9BnfwHNSc8OJrmRiPyJ2Fx7EDJSoGYU
mhUM/wVrI0D0wTsaYpyjmHOb6VP7Xa8XBiZW9/+4iUAnK/gkIhmY1Nv4J9gQxAaAPYpsFXdhqH+t
XfZqG81xtuOggDBdLHpcTrgr9uuM5bbdCulgMQVMOWmmUdu/uKvKI3/NKY8z5/oG37oba1RxJzMl
hIUNo4bkxYM5yrzRRHrLDM3qk4oqAgSTF32dUbD2r1CD5MVD338zgJ4AdFWbq7sVeyFL+ERh7QX/
MQcay67cGOoCFgcpT1Sr6ucnUW1z/gPGHOEfk5n1UDiN5JRDyiCnBrw9Rni8/HKfkzX60xYokrRP
98mzw3+jkMQosqkDM/dRVAfZTDDERhYhibpMTyHVwwsD0cZ67QgILEixNnZSkHqq3+FRGP6fT6Ck
BzWekY4hqXtqoY1DlDLPZc9b9GowRtEGnlghwyhrvAmWJAA6cDS7bATMSloPne4llVJdzMVT7qyM
esqxWXNo1ux//V4GuL11FJdkYRfmju/EiVNq6uCfTK00Od4YTUL9MG6EPY8wTen4rFBeDBhVb4Z0
gvs0X6u615c+GBEtw6JCHWsxKe0gJCcuJssXmN9exTnqKdZstG+Omy3wXVENCCVwtjHLgFjycyIX
EhPrf4LGrx0+6s85+wEGaMbx2aHE+zIUxeWQnxYBouP6moWQ9U+nxyt4xx8sN+hiGW5JBy2yAaBf
QNml/2qe68ko7P7pvhkaU2K414HMtsI6NvuyvfERM2lGeZOrJmqXfhQg6sc4/HdX2TBtLfxSNjWG
rOyBElFqgufSFG32f2ScClqHGjP4sq0TO/v4C5lFM/IS+74ElAPaz6Mh1mJt6lAhQqE5eWSjG3hr
k04UyYpSlhKjvzwtVhcF3c3JXpzwViMzwafuqoOJke94mmQmmZR61VQGRS4J0e3NSZ6HjabNNQoV
YlMmN/4HNd7+LbHh9MXLKOw/0bfaD2OA9lUgf93eok0D5b2kZ4ckp84E+ItqzhpqGfgt9TYFzdN4
Sn8ygScYBNLYtebrNcU0GDTMx9Mv7u/in3KYNaNepursYm0pfu4duFNTbLGxw0App7VIiBqNcMhR
Kp/ja1s61ERIepzZ/OXIoU2lDoKoasasv4QBu4H7DQMapS8gKuyRM961JGRUfLaHr+RYHX/n/Kno
nKmQkaacT4vNwloKhN2wI3pwwTxpJherwfi/q2R+WoOdfXtvhbVAb6T4YI2W2KsCmPky1dBUrUml
ygnXmZYmPcX11jWf70Ub49UPKlM3rvdbXDwPeQOZQ9CW8DM2K1V4B0pjXKls6aXVwFp0ojTUXLqn
WhzveCa9EnjoqznKRa3dVnwtEzjCm6PAhqZAovGewLx47pg99ScI4Bwy8Mwq4C2aNuuxc1fIC80K
5VABo4fnnGRDGQSmfPsPjJ/rikGCW0salDF6/rV3umikvkYS4UKMq9O6tCEaAkF6uXvhtXqHJMXX
R+lqCOvRpXjYmK2a37O3in63oh7t7AqFtwWdwfisxmiKA56BoHATb/YHK/3hshogWhwpwY57PO4M
q07zIx2JZEMTY8t8k6PAFdBltoz5zxMXOCYOiDmbFQvc7ZC2L00QuQSk/ifc4JDEBs0eMlllaLTX
BerH1FMYKWj8lyyd2zBuM3BLvd88qaUHQEiHdom5KHgCPbh+X0pPFbi47OxXmRdjCQIBxQi45Hnh
4Cd78kAtkzc0JYBaqbdzHzJxIG3wLblbXOfj8nBFTZLk81S+DWZFQx3hXJzSOu5aflrnEarcPM3j
3ROEDPTPhCoahZA2nwjXz5JECNHf/bODbpmIPDfqEe2inu+FWJuaKcVBVqsmdOY32jmeDK2DEJEk
RpsPq7/DW3z25JWvWLMuzCwOF4E1qqtwXYfCv1FY9gekNJ3QF+nFtPI0Q9/+XLd8z5EEaLhmfO0I
vTsb1uj4GrFO//f8r6YO6IU/FTsvuiJ8sAzoYDHTaBYZGc5a9/OuXpA9NtlJ0ybrQQuCzKDwAvfL
78l8ETGShw6l15wu2+4Ryq1i/mRvE6+oMz50vyOwbFB/733xd1U8nWQhCCFDbGMlxZKaYl90HrIX
a3f2y/RMbYIBH3+14t8+F80EZTKx3Q7ux6BHAveukMwFGEOAgyK2We46KqlJhwMk8UMCo87HA5KX
FmoVqpJ4+4G2BnX95hFf2dF3z2n/Q0/KgrkX/Fz3dJvPEeXD02GZcGc9OlsTLOw1blVio5QDCpmz
oknsp3S0olkGCaXdUesvXt7OaiaWpwLaJpxY4dsAix50hlsTBWbuFcpRMAqs4Xxrk8GRFvDNQoVE
Oyn8fF02DU8rJ7fNj9YbU+VYdJ6gm7t8m1AXY0UOshxf9ICaDeEE/iHQGifZN6qbya66byLEFUYo
aoRfw2XiZ84/jNWh4oxI46z6RzqTLOob4fWKtRrZAg18x/eOJtGPuthA2L/1Bye9Bv0uz+ZUoktr
g5Mg6dYOyWdBdHn8qrVEHxfub1X6VBy+bTeQ+SfZHktR/hn9Vs5lMcsK3eSNp8rLiz7adwhl0d01
LodSaBpXJBm5rGf7j/dTjM/KE/vzUrJFVq2DtnullmQtJ9vSlGVMf+JcXs9Vd4I/GLpcPcj+84+c
FTw0BZxk51EhQpQTOBiDQnlVgvUt7aZGbb5G6oyXcaV4eRigoo5RF4MVgpbpV5SaGN9/9zbj/erV
is8363cEqgAK6A8fATOf8EM1P+3Cgbk3og68YSH2eRZJjkXZWDJqckjbfMQtkHdl3V8Wsk9aeake
Ja8QcaVwQ0JHk+wTfN/L4/koDS+Bpo4Y7u5QsYXDOotVR4wyZhYBwjDGM7ITM8WY6oEqcXhZKAEV
Anb8OcWnKvEVQ33Equ8UHDcJrgbHx0rPe51qiVt8P2H51Isuqm0Qb9Ysj+64mziGC2rg7oDQzYCD
CCVJT/mmSlvaNGKMUcTu/zctNG29hGMzSZwdnsaFYcwX64o+FsCn/bpUaHVo/OP07WMQgDpL41Os
GIjMAQTxOrHm2iyXf9ufZ9TWI8/2TNR4LRfN5+8yu0Xsu2msV4z7vogfUQCYYQEtXRODqLZwnNwN
vSpIjrvwjcQsIp5WksAPRE17TJYfP8uW8lip5ynkRZlPpQpWBX6KVZkFgN7ILwba57n4fsChnZzr
f/GcCVhWvCKM9VmmEHjLMINABusn6Hra6BajUybb4rcir934ZiNjsT0VZ3itomv0fV7RiyEuFPM/
iLjuoXUFKXa6QhQMeUxy7HFwHY3Qz6kIOgmACDbQKqsoZCJWgqcfKoWV5f41YpaKQak3ZcpAFAJ1
X2ziL49GKoBkJ1XW+wVnv7tU380UZPIJF4kK0jcJQk0tG8YdUdMtwVZQfees1DC3OK1zwGnG5wGJ
asOnLcg7I2mkHYJGQeK23iaoDBWix92+Kif9U5CxGDHbucprq1xZrNpjdwQjZBpOyn5VDvxdujhE
TnBsvmv82yIZqMroFTp6XNOEJOaLFP+4MQNF5TL4Xjx0NMKx2ef9FzEMDVa0nqPf0NGN+KLGq8lN
PARjU1qtBUblXBC/E4KHTk0NX9e2BTCcsWUMsj+PT6KaKNKVOj8zeaKB98FB0kHrMurswCA6tsVE
I43bj8YC/0v5O9ViyZiBCgqUCd/JrTcu9haUotZ07Cpd3YUV+CCI8fGdyYJL+rfD7sKYosme6SgW
nsrOZkeAPWmessI/Rfj2Z/TJ1R2RqrfJD2zEfvN48H4glq0RG5aL5vzi7xfUw/s8K7RXoIpNwPZL
dq5sWPl4Bdak3QkTqgWMLAibl96JaDSTLxOzDFXyq+csm/ZhaGFtdNz8PwYUbwBS6OlIWRyE/ngi
rl6/g/50gDTY4vLdH5G0/aVZ1rq7posva7lLCIflFscHelnFy+USdsZDmzpbgY9CR+eTqBGA5mv3
h9NSgmGbHsbIRuKyXEF3fXJzsJQobOiBZoTAka4YH5js3J5WNDy3cD+T5AgjHvc5WJaF/QKyoKuH
FhhXdaNplORQlzno4Gq29EZrIfO4qQP0vPAHbds9ImuiWoGtuCYxCs+j/6ECzgwI6AxZCqUk+WMV
D1usbCkHM8Y5yDinJrsKhiTSkzArFMoKF8tgxmT49MIxVelRodjoc93iUq3YLFVbLGiE1sNGp+Uo
CbE/3abNhukqrpyr1RsuyhrHPQCvwi5urKcqpteYsQdJIInY1fOlTFTm7RqQwU5LLU4xtykIm6Sm
ul8RIeFe5Kgkd9vzHFLMS1gmvI/e/Ba9qcpvr2/gU13dBM48tkKZPmKaLX6adyIc4XUlFmbBHhic
b7HCcisUy/gpnFTENRjoPwKEbwxldigt4FtXa/2jJl1SVHlY9lXWDqMWNR/dZFiH6xLPDrF+FWNx
PrZRayCvRcTGyhrCLouBYYgUo/w2jqOihtUNJoJtadrL4+4zUfonaEp1xPdHXH75kpGZelFZU3ee
hi3hwVggyEnQDUM+KlDxQWvMbXmuGlHTn/VE/TVBSMq0cmSiie3EcpwkuTFPWxo8bA97g180xZZG
abdgDrlw7kqTR2sB4oJ9++XDkzU5pUpDKVUe5s6mvkqE0cAd1OtkJkWDr/qs8d/Be+9xG9PtXhXd
+yAOMrAuoVrJ8k5OrENN6ZnD1MwVsxfsdgJQIKGwQk2PsIUYxzoxbjkBCjBAd1rCYs7tAFBB0kie
WYoHqfNh8YzXUWTot25QV9+RTWdobP5rPBRmi+LfRWxBXciAugG0E88+0EZPPEGsa2LqWUgyXmr3
Loq1Z2P2Ev0rKaDheqkrUsRLI/0jCrAHooJ3ipOJMlRHFsOBWEUyqyfCJH21THuuVgTV0XeTzt0Y
hhGAsUMA4nLMjWGl5NeEI8JHYafglleKbwetL/1Ouq206jM8M3p1UNXl/rOQEFZGECFJKhqe+xVB
1q/5ajUwkwRty+hxAZJlKi/CV85p7jJO74dTyLqUKwzsV0aYuQ8E8suVNOBD/4N/UxrQ8QRTgYlM
c5eTnLEQ4olsIyWNxLYok4ZsimMzvAoxi5Azy4swmVjfZdcdeHMNrOERfKiK1AP8crEZ6svzdbHr
iRYldazJm5b5E7yGVWtu0rLXPBQL4l6qx7gxiniqRscRq6fMe7o4QaJT2lcQqxN0ucJhzSjFoClE
2RcugbD0XAlq7hmegP2UNdJBQyorWlvZRg9l9CfBDSjhkP5SrFakINLrhD8ddvde78VZWL3BzVUA
jJtepLSk8vYlVhpnWJcLlAeuqMsrFRPzamPxkF3Xa0r7zRD1RTgX6yJ5MQciSBSodxefDptqzZla
pTNwfjP+yDKKByTx0wit6zMTP/ApiOKiInavz3EgCjnii/6+cJLgEb2si21Mj/1hfXpCiKwEFVm4
lkKaD5NBzQAfqIeQocFjlA4WKx0koeX2U6+sREBjhm4nhvQmRCLe4mJ2h1FKVWE1G2yNTyiNKGeE
d37s2Btzdc4e6Q2ONOP+mgkQ9LfIZFaIQS3qHY25FlAzo+bVC8Bw5q/m77A7JfgnVFr8MYifiJM8
YhpiD7fb+z+9vQJ2Ie+lSgqozOSOHcnIh/QfySAVM8VjM9VHUmoa5yoI0+/+gBg/Wl1y2S9PM1xQ
iCwY68Nnd5kUoRmezOkUrNc988qOQ4/pgQJdKmmnscV2xmkjOf6Qdi4FBQk2hjWcgiOqRDsps2Su
YkmLW+39vN9FiIKdqTzg3KPMkVM2Bm6WMtzRtDqUHoDleRC23Vm4+FkUf61F6a/7Pp3rVd70YadJ
S64NhBS35BpMSYdUBHKOxCqiXnJ75Vo02nhlMa8L+Kb5cpFjAqWglW6hZTQHKW1hjqFvO1GOqSdM
6IvQGRwOuJ2McnQQxv6PWQme0oNn7yDUZpZN2SEVKEq2N+Yxl4PupGITA6gmSFv248csT/OTfbtr
1o4IQyt1Va6IesvHxKB6NjSslmVxDos7b9dW0XUV8Hfw6Rb0QJwbGX1Ab9k7hMwejhIMdMyJQ9TJ
79Esd9+FdBRJGLMC6qUJEqF5ANQEt5oK7dj7ap8pjtyBTCojNOKoUVISPEgoyHgt1M3DHxttDLcs
mrumDO50FOZLwKu3oqqfN7FRT9W94J0Mm/NXPbh4rvf/d+2gycNf9RnriFfhuQ9bVj/az956JF+A
ATX0fmR57A9J2rNB1D0UITHorsiaudjOPqAWkIcYFtSqxOOBur4AfTRvhyVkvURrSclBHalOgfqH
GdkRJ/CWuFZQWAwrcWW6ZBKq8W+Nzbn38SQra/K3/WYekNKH2ndFtplK5L3+N3SLLzHXB4o+zDs8
O7QE2WZHO5Z7ejYpAYfYxGPm5DjEbKEgjiXhZ9HUBpEoiZO2aTLUPr3kK2AOablOm3WVfGB6fRTe
zro+TLM+EYagZhbI0m733nqvqBt1RKmLUlt4OHCUOEnkd/Eff2cv1uWhZyrq2PyA4jZg+6vXxAti
o2LFdbgqcCV9GdDOjp/nlB0WDQfftTDoc0SNbfQhKBAKOncgZVsiCj8yFFznecQosSUcSGVdOvH1
odrOy2oysf9CrPQdEiNwHaFKKKIn5By2inn+C0q9ld8pc6+L+cLTLKbABHsVxH+Ctumj/yhG8gov
rRUNgWD9PwJhLz0hc4etX3iUDerfsBdWWf6LE2cK8BNLTTeCGBK4L/Mt3YJxTTQg1FeZDs046NJz
kWx1Te/TaUhHWoIPVxMFSEi4AROxpi/yCckAmNWWP3qtSwnQbWCi6HL5+KEAK4mL6DlLxp9vioPZ
udlQhPHRGsaA1TFnm41Ew8JfNLOKyVm2x6A/3cyA0MV77zqKuYpam6kxgUktj3xtvHz/DNYM4qDG
vMzQogSdMM2eq+OdEq3BSnJvQ+b+NzIBrbFMlA4QdDY4JlB9HPz0VQ6Pd1MwNMmM2N2GUF5/wVbc
/mrKNyIrZLmSIcr5kNKluu/MnmsS+7Jy9tmiFucRSO/dii4pjad10bX4e5cFjgU+d5JvFev0qdIF
niVohuEYniSDva9xGnSIuAmR3AiQjsLL2kuUYwgi5TVbYWUTTYxRwKaZypuSWVNkS81/2T3ND4uH
VoTUYlSEWvqa8jaUEEmMvw35OhLkjAB+as2FtNeJd5OKAcjIawZM0GLkf5z5oXzGAhR3JN1aigoP
zeUSpKFOMtQEJrFPjhe9DqFoPEbSm3434jxXU+j0LOxPtg504BJ++qM247cscuBCjgHFSm5SowXC
6YrMZIW3M/j8thLHHoh+0geAeqFmua/WvX/j6shhXHCAt0aKhLSfRpoGH1iQahWYl9NmE7frLl4R
3CfydX4U7HD8E+g8KnAZGIuNaJvOS3xA1a0swKoFw4PAXh7AiJpVAGfCOrohj3VWy2P6V10IdUY8
3mNTD9fMKxJh+BXpKVyqBu32p2M2obTe+TI97YEeZyjCIzCLKSqmcVcOn7rEixyLRlvIvfiX/BQX
2J0QRN03SfnM//RxPilXY08xQJ5k8Pxh0Kd+y2z08LYMBec9+AJLkMse8g9RI5Z8iiP2BMNHJ5UN
Ks4dU8J50+3suuDtXccTNRpzpc6wG2qDIFi/db0qgWUw66Qqb4OMhnifOxVNMS+2VV8IpFfF+HNn
tStZLpXSxWoNB2bLsrFee9pMeNWM2xbMnbsQuRf9z/z0t/dFvOqBM8c0oHqs5EiUX9dvRxMoo8Cr
aJiVaEqQheyqBq0rY6Vh1dkfOqIbK11x3EmUHg+fYRTM8tjqELwI0/fCwBFUC3eTxqyin3eune1L
ep03G31mwdUPSRxewRTSXIm0unisYd2S3iwHfmJcVrmZeDRpCPihe4LuKnwLz7CHvsp0R+0AqSaB
wJq6+qZillI7zIh1d9V3vAfgrDbHyEfFxf7lkfI0MsfaDKNzMEkCBd/3D9HkgGlk/1GIT1jMUZpX
vneTQcNgQk8misjwm8PSmimgtClH1Fq41LLfL2mcD0+u2nhs+4xCL00yNs13DGuyj3XizpsNWBw4
lR4WBM2reG59ZZNjrz1kokzbLYX8Ui4zfVs744glSlfvdHGPUKRLzzukKJRCMmIFR/vDn7s56pg5
T61pMuLdLDyH2gqTOUlnEIcVChNWetuv2tmlLQQdfwjaj4szzGkCG0S8Hpw5D4UQQYJiM5nvtER1
yJXDfllKEvJ8WN2inArunrNDDk81KvVr5dhINFqTevOYnmaUy8jA5vUoNudJFg0Trvu6qRHjh5J6
gzUV32Zgdn/8YLJ/SBlEyr42EwM/SkK3oBNcUHVpBys8mOIHIv6/4bYU/2TPVQvNoRMvk7aaT1DU
Tn1SquxF9zHFT64h9NdX20n6PRNi6+93sO85Je8qYHtiLeE025vrkpz4oW+PXs35d2JYtkuxwKCZ
ryY1dEXG9HHW9/LJgvu0wi7SRUqcSVuW8oj7pxY0J6Lx69yv8GhRRZukyw12Xi3fsXqkdZsSyrfF
3hLZ+g0x62iAvq2pL/LhgFp5V+yPB0FCefu7VkEE1ZxK+Lp4fjDLG6Dy36EmAWS23qvlGcUaIId7
mn7PfqNaQ3616/MUjBmNPz+CSzVHy6jX9KQtLSeuE87xm4dvXBpgjYenB7bGBk+pkH1CLjOgy49a
nQi2UglxL8JfZ8dipMglIrWtofcP2DPhICDrS3FfsugsNghXuxEUGvl15OOEzxe+97E4lf4Ce2HA
yppHU5B0MkfPbIZWHQXVlB3GAiyqGlBZw0ikLb6XmpIcIN14O9GyFt2cXCFjODwXNluDl197R25j
ewp6e/5h9OVHkmTTiYMFPnWO4CL2H8sxHUBKOERr5ggPUPmuEqOfRChttZWmMJgs6B6RiowQpph2
3mwgjR/Vl1D0AZY/jNTL6xcdUv8qgdc/paCdm4gi/HdZuk3SFLsLisFtfW6pAYKY58f5Zf+C9NKI
BDS4zxdFbSasxeLlPZvsImXEwHjS2afKPW16ZDRheY7VcUW9nMWpN39raxGljVBG4exuKXEuS7fd
h962cfs3cBjtMPaqrVaIhoPaU7THCzJ++jTz65l+CgdZA/jC9/NiHSVJvGjCi2Id9RbZ1imUlfBF
a5lUjwozhMQ1Hj4pTwPlcjTpqrPmL7yUKV/XRH2lfVDp28ZnKwrtUsgmOnaHUAUI5/Fquy+78PrC
tO8pEvMI+VwISZDxPi3NJwRNbRPQhKEKunxqWn3qKm3MHVT13DtxhDbFfhLIcJPc/JgUa0htZ733
7gxDLyzwau1Tb/zbYkklefZI4P/il49TNjmm7BaM+6hoZ2drjIFkJpcrbtYKJI7SPRglu8WYi5w6
V8z1nMkWz7rRcNpaUE6KIWmeHgmJmu2behk/hTIryCnCj0zCZ6RFObN90IX35K2Y5z/aGO4tY5CW
KEb18uWcGuW4Tn3mLWcVYK/O4eMbryzWs6CtRV+o8eEA/woMgJ/ALyDhWMZjoXP0vg486XufW34Z
kZWy+VDFmPnDNdTqeAlQ0x2UW3sTRbSMDOZE4Y6NJOpjRD/K3h5XztZCJQ+QIZAqTaaCazLDFMWx
R0fssZTxwuAPIJHA3CarsNRTe4pmsOZJDMbVMgUwhrFTl8spu77RorVNrPzK2pIzXpOEX4q/ADFE
BBGzuRrktyXw+9dzqY619zkgkoNni+zbGXsfFHUFjInvOZYUNptmVh5H4jvr8fvrdxHFYwIy/bac
dIAdRN2HN4vXLi5tt1grTmc4K7ObwenSxFdXV5WRwj/IdKF9DQxAlW46VqC21qdx/te1X056KyZ1
kCjjwamQIO/eDVcIsbNy/jJNNm84qtSipxFos1l2mFP5h/PTFrQn970kHxwZPDh9/1kh3/qiz45y
F3HYUEilDYXZ0vAZPg9im1ac9B/+fTurbm5ugYzas3jdCaXhoMPVo7aG2RIh/CCJHfQ4wgxZ6y/V
HjczmDzrXmiABG3aQ8U305SPls0eFhfBqNkcP6GGtWwfW5B6Xxd14t5krTClbOI6HMNVazMO6ytU
Loa5AnXd71wsoje2OxtFPUBaQf+XhEZPctMqKyUxw59aWyRehtWkT94WiWw/a77+FnKdeSiL8CuA
9aQU6K0CIwt66yFFsPzO7EaJCB4d5cFXuGAqookTjpDp2eN4PH6A2bn9uAspijE3Ns2HOOLCrReu
rNNTHAFvtyaGY6ZcHt8j079AVQgiFSDA4G010rJWGJ0aiKUmSKq2KvH0yJiFghbxs8j8FpmMyp5w
uN4rvYCjTfHfv1e1Ub55fJbGKvRhmbtIe74wsneSsBGgn8NWCRdQtBvzS5pqx9YKm7TKiFd1MYMf
bLV1wyrzGV8lRjjd6jS9Wd4lp+OCYD2/c3MLzcwCg7Y5wdBmxE/sMh59M+0HEgetopldokutkdjX
pkZCicR0qKuk5z5yjgsyCBWsCthGPIs+8FW9jFH4RP62RB/ueAVrj4UI9DRP5fAOwhhKLewytbWW
lcqzlgCgpsZDo/2zOJQkl3p7lKMPc4SEBjh80WOzOQ0BpiVDtijGC6RpSue9Cdw3/vesit2sH4fC
bM/OLkDIGj967t7KiPikeRJMbCxP+RqrY8RGJ14STqtYF2x6tKQvalZ1v5IKFpZC1Nce575vVB3Z
riBjW0XBIDeulyuzyhlYyKdxGCwZdHV2SeSZ31IlJhG1o4EfmGmRMpA8AxcTnn3Cd2ivobkPCFmJ
TWcsgICogG+lxyA2+UyRM7GvnhCKjmBh2q3vItSihZLN+zvgfkQKY6o8P1cX19wfaDZbZoJeQg6F
jHbteqGnAvil4ZyO76iqry8Y7TDXbCpv1Suab7I4RIYIw3WJlYDU1rhA9fAoCepWSKCMb4GPfag4
M828ceqRz3CcXXCNP/uIRY4ShurkyXHKbbsk8FM47yj6WTJAtXDGzOaJd7DwDWSPZW3hU2BWQ9Fm
Oi8iI7BWeXaf6VYPvqJNZioqdNdT5k+uICH5xL16uSCthcB5AokkwlJSK9qZYHtPEM0bFiljfUrV
Sd7cbzpb6OjKHhkp4d1Y5HB6UKO0dUDtqnozyu0TcrbpMoTlaTweMWgaFTZt46jx2HurdXpCxZJx
J/bzp3Mc3c0lO5VnZB8+9kfzOHYsM8+C9XCHvVcDpIwwBszA9w/oPkCFJuMS8vSsEjhXhduYNkiF
VyDt2n4sXBUOgoaD0kESwbeT3OELrcAMaE/pVSJc6LTf2X7CQONAYYCaQONZAaZde+nVgO6Nf0Dk
STkpeprn5RGRU4hV/aBzwXxrWr4V+U5IL295HSV4BXoJemEHjqhBrn6UxV0gf5vcS2MnSfwzeGh/
LovnjSkuFeZY683Ws17l5didQ8UAR6zT3385DrNsJp0BXJFvrZ6WAVOpv2z7QzvRebqAg6Y+eotD
1zSbiCCWpx7sk/4cXjwZlPw+rK4nBtSeJalCAT5/U/U1Sma0KucvNcUomF2kmYt23V9bXWd2ARKv
JvSYBqpNrRNIgv0/Pnf/PaBjZ8UOLF7EFAB9f2U4++2bnv6hgWGzfACZ63MVk6uN/i2rcqOusZeq
kRKfnInocdnkSz5fCyEgzN25RY4f9JbcST90a+i+iZg9f8VqA6+a+nlOsDteEACVG6kRE3ritVcL
5GpDkLMeo6+I8t5o7wvWPrrRBb2troxP++7rCZmZbXbGytGAGb1SxJ7x0H+msH7s4zxEAi53pkex
Yb5ErgLLnpaM19hIBc97Zm0OVRaTQIJqMLHpgcHGNyS7l2+UW9GLSq9Tn0UnjhbAYs5LQOREVC+s
wpOqE6MbsJ4LjF07Sue5HXh6kkj53bg/RIfr6uxQWpv1zOOwsQn3ng3lXjDwgQVXu4uwPguC5J4W
zpVNBXSFxPEUc9+vT5iSUD209SrCryQmufPCmtFQxakWONOY9HYH1dZrc4DIdrlg8i1nX4rPjVCM
EMG/OMPlBUYNfF9MTKq6UXNyJEGUJERuoj/XJeHBRxooXWXRg3I7x0/ZPHELerNZwELAEaGGce/Y
HH89LMC9WiCstiFP/oe6uwb8W4gtLJeUdBs+9S52e/3+qx+25miJgRuHqqir/6Zk32CnxKV9DHu3
71gIV1KDlhX7bghoWIZKjZf37pyLuuIwktkLva+SfayUM4ekuWB8/KTe9GUwvfPfrUWHmtK8N5Es
XA0g2GIZmxBRwlj8Mlc7oXzsIyhTR1jHHUSAeCVac6C9IayCKdKzszqeOKYkOw91gpTSnmvcVsh9
5Vxj/fEaaHAlMyFzAO9tsNDNzUcY1QixH1eDO72O747AlLJJrFs+E4idMgtZNtWQ3qgiYT9uzt/t
L5DtjCgdCRoOIyxIgghxq3pBKMUdXirb5w6+keJmAYPBuPeOncGcjsD1TodkZo/81S/vrG4vp01v
Y8mrdL18uVvMDhIc7odP/XHbknutCfKcsvIz2ydkUBBxshhUB5VH/iE67QSbxX5LdcVHe0n6VSo0
1h+HpdT/cAU9n4Nyrftc8nxx+nN4njgHitEa5YkBlKI6Pg6vga2Jqeh6IpMhhRpqdV5Zs8v0HXzi
ihifSFjvLAEByduasN5+bpmQDHVAQSzzqSSgrvI3HfLXAnFySS3YdVuCktU9PMlOQEzgAD+KiVpb
eT2+6AcbkrOcQGSQiTtukOVr9rdEcZpIrMxeQVWZzBu1CYJPXM6vZjXJqs6RzlkhBbNaAYvbvnuz
P8twcE30tr0E9P7O6HolwwfP1kddYmZ9kkBLQ3gOE1ZWicMJisDtfFDDeSmOyxp3MrrcdclFEYEi
o7g8JCQnHa+WZnEBl+GJ4NDhOqfoiYUlFylL1yNV26+xRYHI1U/MkShgeCesJLAcwNwrJfFQwJjr
NpRYPL9RkDDij4rSfeFyqzx5v/vkILNSkSXUS8JmjMwnHCoiOvouHQwtNTFa7zYcIOnDaQs354F3
YbAZphK9zKKbd7jQLbZpj0HL0cdJWBo4mvD38408ryqGitb0SVVRn3TLHJ7T2FTn0QU0vq/yPkY9
gP7Un6nks7V/utY+PvW3i2jOVHYweMwO4NyQ0E08ED0pqaG3JsPz15bxBjZcvu6ktZJxdrfAbrMc
bnP/l5cRJnXZdPNuuWH0HBTrIAkYRGHdXMZqPvaC4qGyfjgviqYnRPps22Bty9il1MBIxmsrDdxs
zN0c/Zyv/ozZ8+7JBmuHFwGcJlJrGRRqf0KoSVzymF6u5u8vvrlIP1Gsw3rLjPk5YoxzktRYHqqK
JmpfW5kXdjxPHN2VMQTjHEsm1LzqnnjZqQrsOvK0ObZUU8W8yNN1Qx4qisE3S8XqdTseYOQf0bDm
RkjeSa25z/CI+JQ23PFyjPKHSvoOdLPcoZTsTprX5JIlt8oNALy50xm/UtUspELOH6m6YsI6WtJU
GlZy48XwYuOyLDDRbeeAtMlL68xMCrI5JzanUPGBk6vPOX3H9CdApvyvgGdy3gnKr31JBRYPdqjO
mtX8rxpBAKiEP+GmPHlzDaqVn8jWQ8QrPVjkUsRApBLu5vJ437iBCnXcfUXnwjlqNC6teOYE26kb
5BeS7scx9+1Nq/HUryKrKrw7Q8FYYHR17Ph5ZQGNUqPWm2utRIM90+qmPmsAMxD/y8+j4InovOrO
VNl59UaW5k0aUkd9z/m7Gk4VhtzuLIHCxya2X2XiWf8YXzCZr1HEzAfS0iDzLoRf0sEXGQ+E6KyA
+QauJeQCOGRs4rzRLY37celbTb5fsFvKE8h7as4H06cBrUZq4oXwvuq8/aaZP6ApruMKl19eQ0XG
aB4D7IoslCOA6jcRRaL0nAwX2/KlDtAtkzAH88V1k+ADgHO0kVlkzCn45ksQnEeZoKpyDvSjtaul
6Xp1L6k7TNLrgtitrPOD9rs1C0lI2r07WOWcrtcPvtFD1EfkfkXyaHHWVuYtWMqFc5icQ3HZDAFB
XSNBksO/bX25QA6otjscooxSCUloW126rG3ugCdQ2loPQBVQmjpfctupBhxTaUQL/rKz0aWlBJ11
Viy0jf8VZNkWsxVLH2rF7IkeLzsE5W2zqhqGk0OCW0pakNhRfhCmdaoEcfDEVq+qBeuJhG8o12Mb
jDTvSP6ISRwd0Wfa++wWcGbpqyEbmKvwm5h8cC+4IuK0ENQ4Gif6P06eZEXqiXJxNjLZu9pbvd93
dQKZywz3ucDeTwLnH2poKNSVhrskPjxfwgqPTVb/U5YE91oQGNGF8qW9D48cOQOmBPI3eemTcCFf
Ff4xONUkMxdY3yuQE6D5CMEDcZyFY633zoDJr7ZADcWSxlYXNtvX8HcvhawfrRPbBSAPWAkZLx9Y
t/BuL7RHjS/16pv0ZS3w+T/+x0fynfvzjSw6u5e49hTWV70rs1t6wS9xgtZFLy35JhrSC/uVM4Xw
0+F3r2kDudHOD25UvMHYw5ZNd7jSib8vtH8hf3lYuApEmB7YJtFZaL91wf+XT9h/iyrv7/vL+P+1
UXC/Qo9fWW2b9JbGg3gMt75f2m7ODp723u/34H76qGjcZHteWK4QiDZVObfChg0Z1g6lRSARAiKw
/vQABuG+23KLYlG+YMsXophmoC1n8c6UsuEygGM2w/eblNRVeONFfdNZJ0PMe7qdPDEHWBsimu/7
PqA24VnrS3ZneRyx5a71DMt4gFeDfc98ussDlnVLpYVeg5Cl7p2N3Deu0A3InHI+PYsaSFC250IG
uNiB6d/bKKg72O5r83L+Z0WJU2119igBJ4664ghY0BXgVrDLsqAnqbOyrErLY/ta+2bkiG9MTbdE
WzrjDdZ4X+B4ZSDFPZJgRVLicGRVRysGQn2xYW/aDOC0gqJxkYX+O6i43jKNyiPcbf7+JS0JGgBw
La6IUmpM4vreRMt8/84ZY12W8ELEzrrVEIHgWdJ8ANhfzpUzN0U38XHDXT/WyT/dwN4zb2uQS/6I
VkRmRo2hR4ukOx5X4u+K8FJNc+glAqmvJUZRaL2Z4Sk8DEe5yIf1Y9jG+KvOTfLTymDyNIxMB2U2
NB3qNuzKcOfibG78YuuuPU2z1kLO3zYDYTVG5bT/KEdOfc+h6E42UfaDd2pCLxCytOoXQ+0l5236
rDIumqTMW13Xw/v3aBSnFruckZWtYiSs58fyaev7WD34Ik2Rtgnlu0lPnmEEaOqDVL7dOgjkfHKc
n92W3FnNfwtMPdAMWBHdJ/Gf7AZH2O31we6Gisy/eN/k0zZ7qOvKlm/dBCUzOSAe7FWGxYoxfBP8
WFuCHd+gUQ+0L8l0i/eArUHNCqwTg5dkqXEFZd/i9S8eVgFVjcmblhB9KZynu+Y2vCyrL/XS088W
r2PVdTFVUBi+/P8j67sq8B8VEwZBhLvYE+x9JWvtQZefGPLjmZ/9RxfAvAfbd6ugQgIdkWaa+fmA
s0WYOymJn8TsEXoKCnb4ehKvn8wo4crYx32A//0iy63+3KECmCuGB+WK6L6CoQxars2YauixCNw1
Lu72gHlK1G78m7mOkd0U2SiEYEy/W3Dfmo7lRSdn+sJI1feEy9sRFB0t6uwbAEQZimdXqj5GwdWz
VohiVNFo/+RO7remA+shQf1glntozZaSQC8y6rU0RttdHu987NoDyunvu7ZbshatqwhyKF3wJlkv
PyPE86o6m66xyDT1X9iaCYT8iIDfnExuV8NN4sqxXBZO9cKwjixKIW0HTzpp07WdsLG03QsyPLVM
ozka0OJPFmcR/z/IZ83hrRpVxLCcJQNCPtsnaAtYwW+egPSSiYpIgFFItiRkbXhD3gafNgajJpgS
VpUQnJyoYher+aYdtlsOSW8+4JzeSV47jnN5jdnytRVnHLQwTg6C+5xn40Q+yFdxl/0BG1/+qDQI
Q8d27o+HVEp+jUWbWq+4KZbqSdQBWbcC2UV5Tkt+2TbZvJwhlnQp6h2xzV7Xf/pIyFW206C31IWT
TM6cw8IrszhNYwveZt1kGA4Rsry4VnMtmvobclDWDXCQmVlNgDmP7+iasOcI814BQAMMHvOM1b4Z
ma/kpNN8mAQfHb5xAOV9rWIL4sq1ct1ozeM35BbC/aS2hc7AOWWE6XkieskqeRl1FsE0LVZ+XxSl
StFEJHiiG3cF3NIdzRbns7Z35/gRbAjMpV0vUy7vVp6Q0qFkRoofMtiNM9jQy74GtdrX/Jj5ZyyE
5r6llmtExkoxYcWus4wt/0t0d0dWoYoNHhjNzD4qqLtDPabhCEd34Z4HMhzTJjAVBiozCpVDiycw
/IWeZpw7buJYMTdRZwivY91ZZl9tJkLs4JCV/YEVjcQo27zRHJ+OCte1tCKHfSIfN4k5vCp78rUA
4Qso+D7QXOq/+qFCJXP81yx81UZmD/MjIBJAPMpa1Cz/PqdoA7DG95oNvFJPAZ8DbPgGwYVTr8n4
upNqSFMwN95sM9N7B2yVCfMzU2/DWmnTch8t/chlglqUpuXq6JtK2D2D9rlu3jjL1gThmskxABa1
ZZojTNm869QPt7MQ9hhDI1F9uQiYmlFvllK2SaUYRaafF66xAakFLjcZjOtb8tf/GrzB4B6hFlJy
6WsIFn3mNTbqzPr2pHnBuN3RtAtm5LLgGw+9SH7AtG8yoYWxPFyZWCx3gX1QQbOM3eEeEpphCzsi
8wjH06qSD6UIN0PIbwyxM0lRxOjUcd9UyRQUS2uGYOK1la3OOWnll5Qywk2gVwrxIEjPoI1Kf25q
XfHHIcE8yKrHByLVPLYgQFsmPgfdM/zo2AhYnTBJG+ZNJCtM79SPa3LVDnJif1UCYuKEyG/Nu0v1
aIZO2XdOuzjQFN2PiLoRd4Lw96IWK3JKH8IbnQv6wGFOcZcEkjIVrawJ6AUr2ZtYrIvjYBBlo8R1
WHuQlhl5aKpJIVI+rq2Pn4vYsGQ9tRd7b+DI2j5lb3qsehFR70Cq3why3NP1/3cMOOHUwsfj2Wef
+jADv/HgYW0oLFrsfX8sxs8UnmpvRxsCE19xn1W4ur1+4AJmDb8nhrkDkByAuWgh0AkZO+ZlVJCU
FoR7ub5v5cbfXCjZkZXGwe3YpxtnLmNgBcqDYM9mjBAdfetM2TOBevKH4HTLXA9FyJ8jUj/ujgb2
uhxTkqWDuFV2g1aR16DvjP0ytScqT3G5SB36gT20YoiWUJTtAxGu35R8FVx5kKGLncdThQ7pttkN
8uIGSCl//yzm1F3laVXazHiI3c2kbkIOYcdm4t6LW8Dkr8rCtjry7NZ51OEIGDuvYMN2HcpwfnDZ
Lvw2+TKSexvUKqBQZED3Q1p20Uht80buegD9pktcObfNOx/2u5EL0cpm0EuEcQRgSXrecaMoaHyz
XQzh2mevbzq0ujFUX5UB+1eTonPTkjudUZtOGky2hl94h3e1TpFK2Xs/GQa8GsSidcOH/sflOn96
C+hZ/OH2YaRU9Oh4vG47ThqlbZrrayxoGZ8eo+veFhlrxQ4QtSS3HPlsqfiPsjzR/0WDXv0qypHU
Hmk6kzaTK//V0aab1O2gv//w1z48t3fCzq+lJ5EBqu/5w4UJpj6j5h3EayIY2VBr/Knhuz3QkRJ3
VaCE+08/h160R9m5ySojZczHU0c2UKpS/CmNExorxeC4/Jj97u6vrOVVe847LZvjMoSF+Fs3zTpM
3hDJsijD9Jj0zpcF5quGIkOusckSliE8Js4Y6Pz5tW0OhxSpYOy3M/k3VWFNyeNUmhArl11Gh2j/
buvERDlPSoyqchHh8YTOzNpMLhQmsli+LHSgoTDGrua2+w803ZFfS2Ob1v5hwm54cXuX3BEVaZl/
YOtrYLpfjOoAb1XFlgqUT5ZlnmO5gUN6a64iqk/tCfULkUADUe84bvHf6UPTBthSitTMLqjYqFQX
Xij1e+3YfjUNK0dSNFJTOxrPM80523vqFCB55YMQ3gXejDKmipabtGGtJhHopEA3ZOOJV6wln9TV
Ly6s0icKvYUORoB8tEbw9YvT9f1QWHcSViADfwmEUSOiuzfaBbOQUzzy/Huq142Fc+ihkZ2iKtmV
gpHMjkw9/O4rxXvQ/i2OBtXoDR3F6PlI+EaVUhil0TQEd+1uCzTxXYPanN891LDioyB/3CobjSkl
2xuyRQPh4eCrEoF016iX9Sl/MFEkCPmZHLMq7egppDqukyV/Z2jymSVorgQcmUegoG70PDiPR8e+
lmFdCUqOgHgV5GBntmfuKQ64khphvKux+Fo6MHdtog/xdfj3k3qnMpDXj44bGLOLjFJD+yR57dFN
3H9iDy/ZrkrDvHtb6vqqkIHr8x/6f76aWgXR5xzNt7pe3caXIm02CIVNsGLsMLPyI2s3zu3cml8P
X8sVsQF/oi4b7/KiV+npgItwrXH0j3iP0Vr+xuNjfqtLGnkBvxUTj42HrEFxGd3lVE7uPqjNg3iW
FeGN2m/xHEo1rFJL55Q8jMUHVx8GPLGKRSTWh1n/vT8UeVNevJkEdaUahfDPt6mvnrTrgvuz+WV1
xdUwy/L/FN0u5JbHTOCwlVamBEd6aqh4gproODVmsaNTuWrZXSwzNLp/2ZEYS5fyLrjCUi/khCPe
o0RghTZCNFh4QrAkB9iOzq7YOy3VWixkbzaROzWWZUtg/gCn6S9EVi6dnOOY7FcjSly6dR+LT4Kf
22bts6vxe8eGIyv1CtcftskSd3n2asc6onzlpucLS3rLhi9jyE7mWtVi5+kobNgBBBmLKyDZkyPX
k5yItChSN0oV+KgohD23FsCZnZu3wLIA8DjR8E7tov97KuUkKgS7vs/d8JRZ7QE0M61cfyyzH8Nf
+/8ifOJOq1wtROeo3L00aF3imP4bALCe7ulZFFR0ayBszAy1bqqdGQ44y06W23L3Ux/6TvSXhaFp
5CP8eTHrYuBTiwETcXlvKraPlfEMjyow2N/F6UmyU1m1s2naUobEfqaOjuvTaXFh2VKE0buUftmD
T0zfsBVGOB0FmGpXNqttQ3iPJO125RjbRfMmFREwS0s45z0wGXFIuLd2ngYGyNxnKRc23iY/KSml
StHKloiA+DWpCGh7ir1tbu1mgpaT8aywQB9Jrb8Np8q6vZdN+3wr5epwhpFCCDw5hUj6y2HEzZ4p
FkA2wapwe3t0WVxT4fwqIqNFcxzf7Du3UBDfUpob7QanOz6/WMsaHbmKYEeGTrIZxradciROdywm
oXFKFTSAgOfGCltbQ8RVc3U0i5JHO/OYu1xM1WAdy1YAZeJSo+vk7M2886sOUzkotWwXWtnXKQ7F
GASGKhs2z0dLu2oCbfHoD8EfVt2/WINw9tcR5fkMvFHIBcElbIuXSwnxmR6EXs94LqTmtoIZ4lyP
aRLbSWG86042wY1ZBDJlVtxVArIJNC7tBgfAGh4N7onEkycCIBvzZnqPTKEIGBDtfc7doCJqjBNd
YL/kzaoaWOXroyRFph/CgkNXEDhT9U4Ui/jvgVA/CC1KnrYLmxfNMUM1CLfS2cPXHGJZHbNAxkUP
/xbACAFK3Oc4CfoU5oYGNx5PDqh/I8aokassjb5ifCvHS4RFPfVNgX5hLC0QjPznInxECBC1UnoD
s75KY1NjBOKEGYXJHdgAuf7IPVEhnIYow23dBCRHdqkHMJUSAFOyyUC0zrOy4KF9OQrE5gSRFP7N
05EvZCvJBeCE9nNHmjTKKQCta0Xnq0z/WLai1nSuPwUOHratTWztacfWQpqSt8ok4S6YAeJD5+Im
IZ7U5RO/gfeyKfkM4KT8ILKgdNfmy+xPRdQl3bggS3W14diCtZM09evOLF8tks/coUfmcy5Uijrp
RBsewBJqT6KFjfqHL1hNu1cZQysk1LS/9kV+IvGVyT3QnE/ETRv/OATW/tLEhSz1W3mwiHzmNXn0
Hnj13pD5QD8Dxs3GvaphCz5FgNuFJylZUoG1W3GBe7c8g6nmCSbAUdSFBlPVSXNFDGxJdYL9rumb
Y4o8D+CxXl6cwMiX78PXGArgfdIQ8AFIbdnNK2aavaRpJtgZXD1nXSY96xeO9skxLd8jHAGDdb4Y
GIEcQSMxd1MTWbcPuTUxOo7bmU5KZVFUKhWRHroykbl5Pj7zaYybpr4OLX787ebw8CZwepNw9vY8
zZqlctG2OL7vUiMB6EOsXdiqWW3Cr0a/uV2scL7mdcVSNvUoy0BLuxOWXBfbZXoQ2OLmTC5cWeQ3
ZeeRRmEY2Wf44xMtF9/6FW6s24AZYS8M1dIjviX1SUBBjpU3t+UQO6k1q5ND6t22z9HjRfWOnWJS
QJrFGyN31LV1s1S3llE+4XZeeS9VtSXoCPGAwIb3/keFLUYB7P+qjl9rz6sttK8YXPEbVyQ+Cqaq
5VWd/vWpU7iyriKnUSKWCE1wS6kKbM3X5j5+VUZ9eJX0aiwlfLMsxZAXo9mUqswXsjmJL3v1l5na
0CliD4IXUhBCa7DqQ+ub5Q2TeNyvM7+5vUwsSMHXzo8AMiypigSOVhn5TIRQiPuA0dYWhwzsa9IC
EyqmRRHBL70F3KIJcZnEoUK8GPHNrbjG0/p4H0V0QPpd0RnwPcTmRJtMvlNDOOCSMPwar7spK/2w
5xTcognAp98RuNkYj6bNrCVtsus7FNeCVM5GdYJrKG+kURhdBG7aWGZMafGYhlkqIzo07zJ0oo/+
2DCYeNw+GZ7BR6ONeGlGJ57CwmBDtICZoQKKEWL40n5gi1msUUk+XxfyXGj06GYZCer4SVkuGk7Z
TJcwtAXP6Ll8O1+aShEvHZSDSg1oH2uLzL/cDGTnm9snE6wg2OJDDFtsbSTl3qpQH02EDKnys2Js
VI9MJxMYSJV+y6whLDjs2Dl4IynbbW4Q1yvI/AuU+3kri4eAT0BRVPmpbC3vgcVBGtoKkIH0uyB7
k1DNWJLZKJvJZrRzrjpILgitsc2z+eiIr/wEZ7Epe7kiaxyTBJ1uLk47RjrstjkqZZYnmi/gvDRr
f/Ff6OUhhwRHmCWaUzLxVJ2JUGm5V3oXDYl2OO+gUvSgAicyTs0PWtk+ClFrXVgWfcwI0z3cXFbT
OcDDZ2Ev+eG5OlwWFmXRjFVtPCZT8kEJQ+/SYfWPp/3JJg7hk1oFnwWxSz3xxFTrGUHIC6YbD5Eh
Ujf3nc+d0J0WXAcU0i5ckEh3qJVBEZOIIAhPlFaRLwacIrsjl3+5IN4Du32gjq/ldUTz/CuZDZ4k
hi/3ckCEDlo29Zj9nErPJ3Lbw9e5MQd8aTWUnrGiSpWSHzXlNLlep4WN0FE0EmISpHIp4UprSp7Z
4tVPw8OifjTjfMCby/gvbyLafAvKB8krl1lv46nw7P49/+1YoY+lDj2pDz90+kC9/jQxrg7dn5pK
zHAhQRXfQeOraIQFQ/nBizuPl3CkImwiDCUdJIx80iaWsftidgNAEO28Sct9G3WzAw61OlD+6Hfj
yUhRIOX2OFtC7lrmx3m3Cu69SO+lzLBII/xucfcYcnf1m7rQGYkySmmuLg+iQWwp3Ks19bUXT8Tk
8zOuLLBGc6iyeL8lzkBCFmcp7DbrMvRx9sYBv0DvJVExpFVWdMBmHbREsg4UZ28m4kg2jrW6vt74
XZJuXcYRdQhDdF7hvq298Ni/vJVNqrW3cAxWnHHzZnd8Yv9rNkGpE3/BtLrQB/6Q9YgbQ7YgN3dd
cfw1FEGXI4hjjoxD1i8Xk9Sqvpazpr/GjANnvYTGEXViGcEaUXapYFuxyKI9UEdaWaQxSzthp1K7
qG2/qLnXM8X/LSEgXMRUgGezpv5qQpR0JOQ/Rqc1UAtlMqMuX3Ai+o9Nv3wPxfeX14XTrK//NAWb
i1GHuPlWmbbHjxl33iAa5jDxzPeK7wM0BCSo+a6p1eSi1di6w97KBtb4cIIVmsSD56DdO0Gy2fZS
L5DLphW4H/K05INuhWuJbbrefT1rTaYZw/rJYMds7EUldRXG+IQ3YgtNwrvZO46+wdfrhl1cZpCj
6iTVdaz2wzQ7oDfV/qerX3xJjyhtZ5FAPIwlheYF/7Gt4oXIZJz2M6S+m/ouYwD89BHAYWJAZYjY
teWgFwmiAj4fl9+sUU5GVluiDcMDytMiThMZqLjxbEXtSdzAVEE6elNuRXxBHO/QUvOWN67Tz2Lm
xdJ7OPK3A9pdbd13/yU1YuGdV55K8uXzOHBoo+Emcek0Oi9mWjBaBQq8AYImiGyvzcEjCNfzkZJs
2yglAi0cQxMISHUCCXhwBkDHnPj4I+68m48Ad9b5s3A1tOmXFVSVpDDjVqjXGmgXFC8FoLDU1J/8
ABHyreY6y98ioF+rIqiyK09qSW8fWYHfrXWwPBNG7T6KWZn99BhDfsYt6JnlAGLywBcQEY/+K9gT
yN1qqcgvUeXWkgdE954yYt6eD4/bS22OTWhbqSZvUhGkOdD+E9fbDB+Y9F30zgnRel5kXyehye+V
6KnOjHR5/tqN/fUjk0K9wnV1qtopzIzawySCCkFLtnxLNbKM0YCC/zeXNb/t6QpmsIzyZ/W6h07k
Dyv37XtoMfc0RkAM+Abxj6xQYqRS10FLgFrw0GY7XJoGac6+sCJmlEjC1UXuxGzwJCDdcJebrIAf
Cbc4Vlw+XlRgzI4Zu2fRdvA8hlBXMVFmyE20jIElhNWIEKy6H3Mt1lTfOG+DIF5ZjO1PHJZ+LJoq
Vq2xHlBHZdXNYoIdH0BBU5QNkIQHpkgWZoDD68pweojFWXDyIro++9q5wOCuD5zMIlM5/h4parkR
uinn1QVL6jg55Omyor5IJOPWv0Wys+J2+2dOiJxHIVBqqoOD4uMNWPPFVzsfoi0KnhiqMDHZpgCN
9KywC6OjaV5BVx/TnYQv0/WbASR48igV5Ykz8FFbQdxP5KYjJ/BA5XB3AljMUEFpRX0MLx8Q7vQ9
Zn4a8XBAP6p3XaEVq6nXqofgXf8EX+IStnrQ9fhzSCmka+frklXA/8tlUPtUM/cNPY8lqdwl19A+
2xeGpHFiqpqfjbA7L1c6pZS4R6+h/oPJwlb8R8sy/1Mw1NylxlkYBQXA68KMPbsNUaTfPhrScO6T
v4Euid5sXiciAbmTggOMkogaH7bAZp74CFGWiYve1iPMRMWGlqpImlkpvqqpU9w8qkM+SO+ZPqsm
cvUoBszgI9VhcQCphZ4hbWGky9K9S7XjNDzsMNjWGZ/XR9FlmsiGL2OCybUSxUMvsZOr2q8irmkA
EhinTRLg/UaJ2GYLngOCMaR+obedTtyXgaontvdS/ij2Y4URe1QSOkzdsoElysKd+K7dSGxaLPGN
SK36+AQ/NeEBpW9pBreCMks6X70PJDwYCFhziGG76JbTtc7rGGaBqlXghJdTx74iwy1I40LtbunA
T0T5V+tUgGjY5uZau2zYfzxxw/zRcqrUCB2HldMlh/zIHHdC5nSfIKE5NTd10xnYoezcQlCRpypT
PCRElQWUbY8bPVxODCmMv4/BpfZWacoCHoTRPt2P2XnCBq79ynBbLAqKhqosP6/pjdFEDYPlfBVE
Lpf+hEsw/J6QZJdfEfIZ9SRmTOwjo9KuCKDI29iklkpJb4qRctrfCymA7Nr2+hdEM3p/BpGgsZoy
Kx4JFMXIBiO9F7yf6YgkSK+TIwEWpJn3iqF3/yiOq4auB9xYV6QDyqmwWTo6ZSot81Hmw0BppHmc
NqXjwtqwuUi7QsLMBoqaaEoJVavm7f5xcAssVSLiBY0DwrvCO2SpBRuQmJBvvqaMBU5U/wdCSDWy
TSvKVDaqZrFIIHTjRmMB2DNmN7AK7u86iXEMXmsQsKLhsO9z8kfOeqxuHiCMxX00RXfByoojivHK
5nhi4nyExMNqJkLTmpHTW7Xrj+mRnwD0weQP0m7MdzNa92/01mwojlGLEe7vxbbUfgafMpJmyA8R
+gXc1QtwVV6+TZYfi8vHCIL7Lq0I6lft9M/RmSzbnhbdM5dtavfzi6s0kMzE/pNAN+qKT23dIc8u
u5hxlWxnaizT7EteBoltjJ3jlpnPI1/QDNjhYapaZMlup85Pq2v7gPjrb6T/QT2jc8e4D8rKNO5b
eXTRhHlwCWFr9mOgerW9YWQqNLjMU3vlLRIiQh7DHBJhhkdx0Iog1EX6s5QQNLG9MRVCZcQqIwE1
4QvKtFfJZuBAnS4bHExdRYiM7wDHOBMdsNkJ+fkNULNFVBZTIhrRCnYcoDTN8I20Z9MdHJF2q12k
inYCPEIj77/zDOyalYYLR9qD36NTI04qfGjbD5wsborv2xLG+awLaTDdtLuqwhkU29wW23QMT7m/
NvP0h3zq49vqOOtAhodtOcVY0e0bu2Q0sKRQSuyK45xLvPoVRlEd1n3Fz4UP78aJF4uEI1rUcBwQ
fcbJ5fCJSD6ZaJUnS1D1CNgUwnYt5xoRV/P3F2lJlO3ARkYGRNm7K1A3qychUl0a+YqYiGHn2nU4
LNdP/07zpvhVq9o6Ww0WsTUJui3mK5chNOwPAyh3vLXoaz+9VC3zuEfBs87vlovGf1hh6qNZ2arg
y9FIIiHaSSD0NwzYxSvgD9ljVQasmPP7Yco8m/H5Ub6nym7QEz52twJfERJRN0ztHUaFSdM4zhUe
KZC/S7X830m9CDCJsMG3+AQftRsx7ec25mbVvAfnp/nzq0KVWv15eud751UNPDmjM3GnhLv51tqd
WV2N9++EwqD97GRlllIeWnXTIfmnRyJObhIuLMZfcMGo1r0mpikGM6SGCeP3DPJHFiRdxoJMNqne
0BZqKt4zRn3gkV4XJ2Wj4e8bDT+ezsnGbcREnEPg+D1sMc3H0i25F+shLpWMJ3amFV7ZDLIMaTPi
0FeNPhsQWfWHbheWIAqd4nZUfElC9eq++0BWd97qBiqsWELmqH0O0kaDA7bEIeOpyIayKutiju8p
aNnNdG+2E8dCE0lWU6WjAMms4LwLoYuoDfgLffntFs2++uxje+yAjubtQ/khXCJAX56KYOF9gYsC
f+zAC2Hf2dstOo5uxKtmH2FWU5K5lVmK67sy7YrdKYiAr9rRyAqXZ8tiMQaSfkGe7G2aQwDBaE1c
vCMSd6zpmoMADZhN5o3pGfxIJyIf8G3vWSKs1Za0Rcx6M2fm4h8+Zxz5ZmpOUjP5NE7QinWVcAFu
Lf2em4X/YnCnqFvNRQ1EtOlJ2nyzsK+w5WTC7+FrX461ItfNITJbFM9In0WHCxoLDnhsAkc7Av/m
5zrru5DwnHzKywu9c5VmeBlkCyeuJnLoxDxV3vKAwqULVnPPLIBJSJGy9EasvyA8f+nONra8DXDU
D0VIcBAAwrhj6lQG6Ht175UO9APAgGnk9djmHPYmvH7FPKsCZHbM8HTW64dOTXJgRCiCGirLbKcX
xu98M/eywgQdSJxNNcVgrhF1n55q8KZIRerYz05T+HdyhHGvqIe3AkPK+0aPpakWhVCAcmHiiIYt
bh7c7Rpiw2UCHw3QlnGB7gAQmFkymbR8KZeoEcNVytWlUXSZfmCuaqORy+QVhu+VUalLF4gc8SaH
B0A/bs1txiyZItVXv/X7qFM9DFU/6kUMSTwMVJYlk/U+9etNRXv5bCD/tXdVDEHLOCZi1s2NQ+By
Zo6rX+c17NAzAlH4CupCk5cXvOqd1BeUKdpQZHB1ApS4r+PzxD1LbAldLM20eul8V1EScztRB+kY
+xz+bqoqExraWcRbPTOviLFCr618x/ZZdbYiBrkw+gP6dVr4QzIJ24SFVlib9vtd+6M/4rDzPRJN
FN0ZT332lUZPMKSo2gDKbNTzIPUt5KhnhY3X09xeqMy66JPvNq+T8QSUXO/79LEf+VRCnS51hEOB
h96RzC7yDCL0bjjIeDFatqcSoC7fKo1u1zv1JWJOGzPYF6KG6yhZxX2fxU3nbI9/s6j4oQoYoLyb
HHluJFgQIa89PSaNhjH3phY3pDamrSMD/BgUHpVLXCGpAAwuFtYhHYDiJ4Cw/qBiwpZKLAKYRlRy
7XHhkDT2H3o6OkI1XewAx0xCppXZqqIO/1SB3PSOsByWwFRPXeWWDEHErKjYm3L/4/3qLc8ljeaB
pKMrlF4KBcoam+K2AgD0uDdZPUJBRd+sgbgDsITlZM3sNO9nq7OJ4R6LNtYYGni2oMkV7eo0TW7X
/y4Q4BPPfIujnT+eIa68cw6rpkM0sCqueqTrpUBOUfNIb/HMoMRt7m0ASX0XEV6jv7V0V77teNI5
L6zuDI3qcxgFNev7dLHvcMoCXHA7QsexMhjbiPSIqJNJ0XI7boM8F2pEhF+gYlZ6ZYlfn7VzZUsg
Tlo731EPGzOEEO3T92OInKWPWzVqOh7A9o3iH5btPBxsrGv5IPtou9IFl5Sk2tadJYwb1fQBgy9P
qSCva8PvyOvlevggXe3eWnMrAZQXczhlzPZmUv1GYs2c4MxXXGsXxtnbHNvO8fZPZIprBsvY+U+Q
wJARXwzIJdxegztzlomtdL418ADeqT0nwJZjFtrnWnIQbHtqVCcQfglL46uqZk0z1wqt0taCgmdR
Nq0K2x5YjlOy7cHbkfXeMFRe1prLDn8tDKstQ0kaDk5uJrQhoj04yw8r+SUPL7sWobVdAmuYZhSj
ibZsEfrO+LBGLaAK5Sp5l6v3sa7MJ1Mq5L8yFOayMfWuCf6Ys8NHTW1YtH/TXRIiO4W+NM0G68I/
orNQQ2a4UvpnPGptf/9cpXzBByFN8ujedPbCKkuzjM2gOliSh5fCBdDlZVDMrvGfBWQmz24rkF3L
LpMgzio+2cF8eAtOsBtbKoupYRIQTk4P7SV7RQ9XTNSYOZzc2rWMNvSJ1K7KQQFtNF2gikLJYBqJ
Rk8QGbvKOftvHyoSAiDGmr5TaxLY9XFpTsFRQwmNnTLLi46kBjQWzHzsCqtANHfXIu33WpZFeKza
5mTQz/6BYMIyS/VDPBU9FDBdMwAlOo5/dnzqxqiALUloviT2Jjxr/vIxCXpdvQSaNFVXS/aYlcrs
ivXLVGlNQJtiokAOnZ4uuCcuDuUxiGdNn8J3f3TyqmnBfiFlObGsz03WKT0gqB9tiDDy/XBdC/2E
VAhav+SFWML6hMSMaeQitYxt1NbGmBZHRnnjgW2Dd/izjd1UzM0HJi/N5pc4rs/MAkEMzriN0vhh
AlCJTtOnr+pALLAXSvNMgqdSxyom1tSOpv1yDZ0ud71PO5izN1CVCKQuAhDM5V6zYRAi6fbAEtrK
CKiHvMtNeLgqgGXOtMIQfGk9vgQ1UINf0eGFRbOjpflZ1dgUzBodUpMO5N0T4ozou12PHeWef2Ez
hkApth9dEiPWVcFrCgtNHpC6MpaqwwZrmCXzOo90UkgYXaKjYX2Dc+LDhc5JSy/PVtUuWuDh2G1i
YAvJnIhfOTcQAkZnUPTve46lfqqzfwyIvTAGS1REeOGqAGT6te85XjkpDfqAs5aphnjA/NdRMtaE
VAWyGIrCAZMkj1rB40jvFN+LhICu1hoinSfeRZdA7XtuqiyNJlQJzHxplbb1fqe1lQWJyLv5zQTd
B/KayFCWVADZq5ajGAiESB22HqHj7mIp1YU3RWhMeoubZUtVRK+HxKdjEOaUedRvnQjnfwUbAlsq
Sqop8BcxUFL3QCC4hWUXnd3/jyXtT1KnJIHhmeRpdOkybD2O+npGOA/0TkcXStxXAgxN+6UWtJGl
jAVtGDNr5GC2oebQpbGoOH/EuwHiTgLXHnD1pVd/dpkkUPihGBjPwn5A456LH/hOS8YlAL3fEzWH
sq9K8jzyQ/lcOyr4r/TKjWu+y2G2Jdg+hTauUNEb2tHJNIFPGXoE1tcIiN4BYc8ufJAUjp0QzJzr
OdUsrnreW6eLmUlMyDBRvjhiDKwBHpajUDZQGF7Sc5iRTUZAOWHV7aPbloQyn34OJ2/F2K7Gtz9C
k3gN1kfWyqfLqXR09HNvGvHzh/c+fFTsq2uuRe2m+m9YGGQ6UIpn0swba35gCxQUFB6s0LvBZmGa
QjtcYh8QUMzGpwQ13ARBjKC/+Pz67ifBK7sbzv0NZkG84x2C/zRc3COntt9NbxhGv/O3u64a5FMs
SSF80bpmQdZgCBWZfy9FNUIeEAZXRDcm4m0y5npN8pxejTXvTSqjIEY6P2h6jbgtG/vQj9MusYGz
kIQFjdTUly+efK4SZ+5rN3mrHpW2FrKoXPw/9U4eHHwWfL7d78MNfDc+wuYZoRAhpnNz4/MxH7LR
Ps+CHOa3GLV5HCaJvZafTCdBmmCsj2aquuSYP+TRGriT+YHNsOv45RqPZLoSH2LuGa2vMyj3KndF
gALMh8/2tKArUYCLYQjA9JVoZehcCax5DWYcGbsjkbweQ2OiFBmgkIsw27anFBR6XaTG1zbbyycv
nDIQh5tQWikknpeyiAmt7CNRoix+tKXUpP1TPQBVwqiHmCRVBkKUZg3BFx9G1XXAV6ARYeR1lpt2
1MF0QtrTSnIgMgv0knf2xeWMpNVWoTT6826pXjPpP8BFuQLU3qD4iS0vG1Ti7zk28+o0TSDvasKq
M+WeukKk+xMP2lGIhoW2rjubNz7IT2a8tUp5DLIhkDz860uLInUdO7xjTUy3EDT6F7SCGJDN5zXX
juLBinah3Flf8UPNSudm087R7kAodjizS8CThX7oJiCbcjgqDLOW+vXpJnEMzMgPNjFbFblGuYID
6lmRXsTli/eeto9Ol/hQA+HzbKBTPgSA3YOaEOYiQTJCBwLQsAwD6uuLUw+QFOYzReZKaURNfc6F
8HtfrmMBRYn+pAWvTqIk//xxwZ6Xt/77443Idyq/6UeFbxYQrqXD7JrmXEKSNXVvG5BQKvPygSnb
txp45XKXNBEZcdpBEnA8G15cAZ/85yRbZ6SCwNnA2bDahf7S3X/u3JdcIDsAjppLrqAEQwAwG0dV
v29UHp5InZnIAbvqZvIpnthMts7t8ShNUTDjwRdMrv8LRU/uwQPypmundPYdqR9SH/RzDsL+gFjK
SVD+KBGtHbFINqRtrtYwLqiV/UcgIkTsjehVuK4Hqnj6Hi3eZFxIXWuWfz5isz0578eAEfbrvyDg
g2ROe890yj01kWis6mmmOFNPeKDJ6gpHZSpcEdTBhHyI6mKytmMoWohNtr1Dx6Fhp/lftwqt7WbU
Ilu+FX+vEmAiNkQA3RSMaJ2Gc+7CqUC93u9j5ODj0mARAedJFbC+vnCiyafIP2mQiloFOMm4Qtzr
Iusun7S9xVUpedjc6TTsD6Ygcvdji9Dn03lixAli0c7y+GR9EDD/W1hklKQgR/SK0T1bT4QbQliR
dPlEAuaV6q0JfkLTiuzJK3lc0l6u9BvdM6Mu3pCGBcDPKwtL087ClwSj21ur3tEk/bTBE+nFaGs6
oVbJv63sGZOn5cruRe1GLy+UXT8pwkr6oFkAk0VZrxcREq7BIL7fQ5cSPkN+V5KsnwWP/76agapp
QhJm9Uhu1gi5SqEFEDWklNc1foiOe4efjQEa38c9gwJegZF2nAbuG6+wbxUH5XxMpqS/jAunJ/Wz
bOZWwAS2kdoJKwAFccVBYgojzKCUCmA//TagJeggFAJHWjtVxnhprGJYH5G7v5MNXojBX6vaOYnP
GJfAt0q1jfc1H+8KQaI37qKGMh8yGgAcrjQGlg1nrG1On9NxLLv7FwUxnY4bu/z2PozFnZZwE2dU
I6Go7wQ9l2DXmWtUbk2ekVWDekp950bMi8HPmyzxnNtkISQgMbxxIB9DpGYHzABkIPqCLi/NWdcS
mklRCpAHrqLCJdltPpVay38xL7GfzbsUmbo3p8mM2BSLdeH02W5jKJPREkY9OlPl2cPqIQncRyBk
di7zFOtaA2mj9XN5YkCyYN+R73pvlMpvoRVmHsPqFr8sd+kgBU5txBhe4ON+9alEl2wYo4dQtGni
RrbD2MOuisW30hg+CwWO+ZEtC2bpuF3lUqJzzWlAA1/aumonFMkMBYQDoHQ/QkC5RiK5pb1pprKQ
UkvTKhCq4Oa3H3WwslhRKJ6f1YcgUssUYmKLWDnxcM7W7XM2+p8ZwUz0arK6to7/D7tXVduO+dDM
Q1UmN4sO/9PvYoTJYl/KAVunu1wVaQkQ6/Exo1KvH+lJYyhONX5Tbj6vmm2f3/XsGRKqnKw0MRf3
Ry1RuYHCc+Tg85AlE1nfyBdqJ/aOlLvgsvc+0plBwJmC9tHq92Lx8E5lE926XAxdLhv8V1HAW5rx
ItNbws6wljols51TFAg6hPuot+IvV7CYhDtLBnyWHUv6D1ufjw9uj2D/RjX/dJLcKzmaiz5ydtJw
fNHFmX3us8iTTaraa1NgfHDNS9zAjYpNCDXQdlwwdKYUKDEI8e62Y6/Gh96G8Tu+gPna5s2alZVW
p+Lxxi61UStLje4FARVAbiLZvVVP7kGJPW12lxIHzfRMkUnAETTk7mhkPA+7bwvvtfrPtm8YmfQz
wDr7u99ZcZq7L6oclmfxI27mdeYIuve6nGnJQzolzcP1TvfUgWXMBOjU7wWtjbVxLOhtYfyBozXL
s4f6gqFGDTjOLDvWDmLhEu2J8sFXZhvojBsyogLgfH1Ob+8Bt7gVsXPrrs+HyacJqPwYtHd2m5LS
zW4bhjuRUpHY6XhuiL0GiJwCmHZBFLGTYPuO4A6ZY199i42RNjmbaTByjPJeh0sLss0GS+XWdD0q
ya5mUJEBluv1fRPwP4caRJhKNH57e2eD3H1sIURiEuikGrJOivGzbLbpCdASJHSXHz48lanqixHo
NR4NccgeIDArRs8dmG0eX+bbNy6U0WtEciEQhC3RupUrNc1NTo3JDFV825ga2o3zEt8VX7HTG8RT
H7OdX/0chDca5EJdlOmmpYI+U3cTn2ngPpfr/q5T9CDQnpwRLP4VHlaK/cQQCk5uymTtELn8egql
rzouWxEoLFt11yAPRhicPlvhk/AT4sr1CkQVCQISTCOBOwcMQKYXGz6q5BxWnryzpga+BHup/Jnb
Db+aQn6/GvJ95yRxDZEir4FQpGJAwcU8vr2xtYTrn4sNC0FSDquLbVDZtEPhHpuuQEooc2TjxYLF
kAgPDoPhqawLP02VQSI6QrgJecC30gctNjzkixdlZ59fU53YPxRGDeCDvM+wDr4UWj90jMG6wQJ9
W5Q4ev+oQzXGL7kING3oy1JojL9ARlegtA1xG7XgRCXjkd/UVS0qDN+CHGsVg+zLR4XUD7xNkXlu
YI1r/BoCQ8ixRAsm5ZJ262oLeP062z3BjcCJ7NKfFtesd/Fx9dcGeHakjeF34fhH3v0JvvELiUwu
hJvVpA1ydHZuEEdAEQO6pR1MyaNLjc97DigyVkkQSJp4z6+xsS2A0808OH4T8jEYJ5YbpartxLZX
qMX4WSBTKxBstbSm7Q5V4Yr/Zkn48sQKwmEVlkX0Cw6L/ox1f5H9F9CidEk/bJ16sbr6QyMLqCiN
USDWIxaufgVajTXJOAfPQrxSl92Kxboqegg5kbW/G3iG95lJU0LOLbrl8a2aZMfJpeIE77x8RIoY
YX6B/MoowsAf3FMlsmk4rWjVESVqm4rTO9vp9VDP7WRvWlT5CHhCY9ktjUPc2OeUTcPeIxz3zzzS
UlKGYS7irL2dp8bGFjBRY6sWetHXVI6vA3M/4VjpnIRT6As3DetbjzzR0nqfXL4mHTZVU0mky5c7
B3d5+mUsuP2LuTXUGOSgmhZxKa9u21SN8/NeYQVzMiEm2Lgs9NbmUgIRbONvpmM9btBqz6iyDvZo
eAbUkPvwvGUZDzfvSYL6roQS0BOzKRt+5Nmpe1Tob73WpAlF2ycjJGrrC5gXBAL/pJxDdJAnkoTT
1HxansJo58Jzp9fwIPrw9Bat2zwuM9RB3ZBblpa4onr6MdUn5TgLF56rX6rGVBSt4JC9EabAsN/A
36ohdyZGjOw4fBmoZA/vFQHMBpRqMHIVqiBCtQqjePAljif8l+Nf9ehXQTDpoSugv2eRf8qmQDqB
zduFbfMYpLe7aOnlPWHPumsdWJ5L9Y9WaplIaVpG7Ivg/J1OEKMMwaLVc//4HAzktpaSyJpGadPT
m5nIFA1nq2L7gXeIjjkIBhoz1EGXP+gmIkynzy1Rkk5OgaQH/zJIU7H9imX18p/NYQ9IS6nPOsc/
Fr3/BU3CyfnvGauE8MKNyQBpmRw4mAH1UONOClJWU3pEnNAJQ3cGrv4mi2QQvk1VnpLltXmA8RWo
bpuaBdqohms5EvcaJhWT+SdHMtXx1rZeksktR8rOMIGKO17xDDSEZDnsIYblW3l4rqJdGuHXuHr8
zuhD5gKfQPSzu4MHWteGiKaWKzFZhtZxVo1Sab4KzQffQnC7BF4FbCCYdlioynjDN7kCfHi4Nqpz
E2YvLCGKn0grLOuVrZDwd8H0wYwjLyg8wcGIb6Mmw2G3Tkutk6CX+e3j73nep/jU8u/zyMmQfHsh
84L5PAxp1dV1blGDDp3WqHFTcWH1dmlNmXA340sFXiIp5Q2EDXUTrPJEFlzZ5fSpkQ3NgaA0vpqV
G7u7z1E9isrwnKLSFhlxQ+mJvVbP135D1hMKxCa5k0WYE/9KSOO5o1mJX6tZSF8bzgPNF7VxpcF0
uHkQI68Zxe9GgmXXcj9Yl57Gl4Epm3aTe/zHGkFQVp7YCgA00k8EWY8Ey5kJR9z1Evx+a/KH43S6
kaPGrpmHKaeiqMa/Cx54Pc/rw5BxOI3Mo32O6KpMQZ0ohl+TRwxC6PlxaEca3dPEA2t+Vighi7jI
TU9bK5Hgs6+Tr+dM7sdqxxt4ofMY2FX0SyZ6QAkt+N2wZxtDOH/cT7A1qccNFv6jNi7BBScYN/uB
LJU8tvs4TmFWb6n70drXqtDTsI31SbW1n31DjlsEk5JbGBoFf93Jgzwc6PZeeVMG782FWaJBV57X
8r+KjaGEGeZxGn/sPbYgQVOfE04/g337kywqQz3my4P8vfglOqYqQvADfsKEd5o+odyguFFFXleD
CEtNHphsu1F9M9OITktNNFZGVdxS+dTeLw6r0/hjaYDq39d/UDyD3VR/pyj3dqRL6lG5ZWQaH3wV
kZXN4BK57HAA/KRPKFyhbKri9SO+rbbP0TzUAAUO5andH3zo7SQDXp1zhLOnCydNPcxIf58T0mqr
buiWQTaJESCgZGzADffdegGD0AKUuu3OTFdHd5Ag2mqeXYAB1DhY/yJ/Q09vNpFGdyWPPKA9I1O2
Rqz+DxMbPOECGXO0xrmIkDN1kX0yZXiGqeZjXbygz8a5GFTmVg6rCuUyQnz61T54H6ZevLsYlTbv
XQHwBFkc60pwCMvwY1IOaZPtG7gDYD+/3TGEGwQTenefK6LtXsdGu1PeqvjE+cguE3lq7joDZL13
WYddsqqHh5UvCQnURJsvWbUgPQ0rVGWVIX3t/0skynslnDWGQBSb2sg9DDcaYQ9ioyUQtNnll4/1
tWCAZyJOtD65cC32U0JTWd1SVFrMt5udL1PpgiLYOVGqcruIQYYmt68efxextL3tofN6lagcgWpM
pSWpHvs5GmtfLyZ/Y/RieU7MA3QUbdaNG+9q6Z5X6GbvV3r+49OTwoyQNfVztSAJuCWHWqBdQrGQ
Zhp9UBcFhf4MqkHpcWtfCavIWw6/lgc5FCKxLgNGc0uLj41lKe2bAXzR9OuS1CvlZ5iq75Md/o2m
RUA6daZ5i9xjX5bTdzCG+sNqMhVI3aF5LFtwG7QQ8WmPyc24Cu3qBmKYLKGyVuF9hXv2z9wlw8/5
kZZIqDF47Tefk3EIqiTvfNA+R9jEmWIcsvP230SspeYouTjOTwmMFqLtuVYMC/kH/H1YwwojWld8
OiJNImhYmwdBKvdzyq7Fp2EDGp/78VqYvIF5lhHEN3Ic+E1CyGpfhgr0YeNJjqNl0CLikZTL4tIh
N256u44slfcf82s+rl1Zc7jQyS++wOHrIjMHP2/QoNwvmFXbmgTU+goRwCS0vISBwmJvrOeoI/A+
xyiAzvN1mesye/nTdQBiMVqCe+QLCB9IlgAgoZneTMJKe/2RITIUWaheeW8AxMciRuqqskPmh/Ly
eGX0s4ONtk6csLKWBBlEQAlMSVW53j4e7BsVHgdVqTheyIlpLh0RnYRlh8yxUUGg032FQNEP299p
5UqB2biBvNecex10XQ16zq272/qNAHHCvDdU+3eGD8btpwkWUtqzV+t2/t1gq5Wy/ELLk4V9Is33
XbI+Z3Kd5dnjkvZ+JYjXbuBldwygat9C8ElLeg3aL92URLme/fvo9j4IkYMeS4k4l5QXBHdph+WN
vURIStWcP1TP/aZMhrmS0MVnAqfiw3BieoHm10DddsNJktfVFCJef3SzfB9cuUURIXRtwrOKEUjR
S5kV7fZ8AZtvnzUyXfj8J58vb8PsfL1QUF8AbDHH0Bs4SGyEFjA31y4KH2v0knE/zK0JdVvQj9k6
XPloSCjJ6x3NgDiEyC0vlmcIS9i138Mfrz6qipmwLC7YmVp72+z4FdaU/k04crJOFh5wHS6a0Tm6
VVaCMvdPLS1z3boGEFkwHNdQoKDE1NZDCtFy+0fCySIikCi0pkA6y93RIVYeIO1mRMzNxxu2q6g6
pptN4QL5DTYVB4yuuWicP/eVaKxh6Du8LeWdTzUDMA/R+OuZLGWm3nksaUs5G5CcIRL5r8ylV4Qx
r4T6Xxfe+4YmqHkCn/Q3gy0PbW03H9VXuwVbDO50LnmCOhCHPCsr9wsZrNJkrfMxYGCIp9FJNws/
AfC2suDWnHkoLfAuSwGZ8/oFof3BqdZmSU2C5HeD5K0vHrC2/GN2zGTaGWaZ1bLaToIcQ3D5rK84
aLppKz9UXU6Y2ONHjqSGVrPcIQpey5GajKgalELsw133qdVWwoJfnE+/1V6lqratW3ca0nEDxKPL
V2qa/doQZLqNmw+SpI4NWZ6SHQ9fDwXeYHOU31169YSukhHwsN1U5OOHku68e6jRnFQ4G/0JlVbo
PJHCRA0+O4VTEst3n82zScg99eZZZa1VUdUJ7laaauscbwOI12wHr6MvAI2MR6bX6qlrv52ajeQ/
AVMd3fFPO1wCndN+RwEl8VDk2XT27LGgOSV/gMBnQcRlGqh9KLM8YDO1J6UmJ2iKy4bUsqzzHFtw
cXWgxHwxxtXfZEvTq+ItvpgnNXuoVitlmE8vZNcAk6LCq3HpVLgMwhB/v8+8QIeHTjhS1RgcDK3C
E+HReJqgY+mYCnn+klYNFabGr+PGqC6kw2pSM9+Lm+ItD01iHkWmEiHRqwL5hfHFDNXLezem2REC
1aVyyVsJUMX9CuYF5mSuhhTIfcbttMgXzMoDA+7ASof4XVHDWFOILBHS0ysk4fZsBVIXxnx2Oral
T1D7sX/7Gqrt9ACapzIYrIIT0ymaEDxIuV4pcxw1wIcCWFvF4elfcTy5kcY2WApLSur0l1RtuJxn
HA+RXkTKRQYdag8RSpZCA3oeIie36ErZUmqTOrvbbki9xZDwIABDQh7Bf16KBANUk+tma+vc/WiZ
cRVrJohjCMf8T/d5Zx2S1FsIqa0qDkNMLAlKI3yWCJFRm/YETqbNDC935zWh1KXDlttW8UjrEiCW
DUD4l9LEBW1PBWmXAM/wux4n61DRatt4Lbf9wBOQwr+aco0Po+YVA3xFhWg+ltstl9heWR5RA6Bp
BIflimEcZetc8K+z//Y4LCWPgEdoWplHGJiDJhqZikQxAX9/p7jvEIISWEGcCqQzjpd4u+6Phewi
IZ7EjO7iOobQhrzVjEFtiNYkZMAzPfSFNpMU40ac/MxOpKcx8KhVsaTn/h2qfRtgBWACgNWHSN0q
hrrB8A8b3/sIA1OUmWZga9645pgQMdEKhjTVP1ldRhG+cnQiF8qJ8kmh0tOnP8n3KLdTVrcedYa9
ieFV5yOddEliHsjsyoyaTk5cqESyUnH7xlLA0ISZQf+pqWdkyHs9x3aqaGDqG29Fl01KRSbYxoyY
pZ6rJTfAlTEBV2CnPM8uUW0KG9wCwikg2NhVrT/wbFDOR8De1heuPy/JeCSkbFG8KrHKRFqBvRFJ
loRhs304Gu+PapnQJykckiiGoczQ5wEN6t/HN2S6nLFdxjf3QpXiGX21i64pelvQdj/pNb0g9N3A
UFRob8CSI/J2Z9nFPxEMAkXJATopG+P3Cj461pYX34LDbccE+gjo9OiDgJ+ftCLlyaMTAmsJn9Ql
yPz2EdvksH0NVlEngnDIk2kL8nLKXO2QZGQau6H1vRP8SdciW+/SWzTgEQU/MxHCdyb9JsDh04Zt
WUbeokxAJ8iDHS1RwInGwtuhpb/ViiZS3TfuMUnG0fNQ/sqFyVlkEFJy87duxkHDwMy4qj2303tM
oUkpr3+BKjqecrGOWAHrPEDVGNxLNgxpwqDzK5mbsa8D7jd3SGHVKQlrfeOR5E2ROWhzuxZIQT/e
A0WbgueCz8YzsBJaylJpsqMUcQvOZr/2qXZrYjtJVbu2Jb1MkiVvtJz594WEcf7be/DaNsPKhuXB
j48sFbJnjgoEqjVZ6Cs/MacddLvHe0bcijgAOmYuff/bIRsLuZpY5Z3N5lRe8LFkE115HcHg0/Jd
MHpDybp3azTpVGw6N+dlqpIkkCLoaBmHnitqkCC/mCwFWT8KhnZG6ZFSxvX9GFKT0bWJadtKcU0c
QDBpkguKc4YOuCobzJ/OYoFL1jwa2+BCPBhl5hndqcLdkUTcapye/qpOy0XxVdiwcgAFHG+DDAHq
5rylmPH2wjxIYOrQ3rE50jBQrHExKsedxZAjRmi4hEtcBCglHvZcoxaN6vEXtXrlMtc15OdYtvAK
ZnyfBXtUQwzjP9OJ/XU68pPN/ZX8IItuPCNz7vSRw8zumV1jw458byvcP3b+1JScTPBzYQnzaQQE
pQJzebTbzhk9zx2dyuqC28ayGquKJ9GyuSyYYmBndcdYEy6ogiINgLCZBCY4XprIuLbK2Ctbet8V
j60NseWOnih7YiME+wYKzTNf4tmdbR8CHUbWicTPDDpwJLHgdpN0CykOABoQDJ+r0CcyOhbovwFc
v3k5LhfwhFuh4tFlVNEJwjJsxXpvjV+p5z4ARA6YdQsi15AaEVHUbxbHGsXBzSW34PH/fAygNse9
uI7OfM1RrgWKrc1bt1tVR77T2nH6FUxBe8T8iB9FhHxZ6RqabNf+WyjjnnAKhbdlZpQarKLSuW7l
FziXHYYszeYVTP5PagmvlLboo9mqQknuzRORGj3d1cabNq+BI1ZkufZse7jGtxxO6ILCSbPVMGR4
iDHoXb83Pg7IGlTqwpKLdajEHGcmuEDcqF9U2VU8ckznojbcqoqOfbzDISpyMxo5ul9M8YyVwlCs
F+uU6ujjVrU2aEs9KQSnp4xuN3FHgZj8vqtURIoYHVr11lMyx47b/hnxVFV+3caosgd71DWMfLaW
WGM9VILiXRQQI2cNnd8RgPdqQ936c7KOx36zSVljP/JySAOje4CPUkkgHcpJyLeACFExaHrMW9Qc
BcwJ5OSErcCRMGIaDGC5elJ4J7HZS0p+yr3XWq0n1fRaskL0VCXscegi72BKsZg1LWLN+v3G86b5
9z0gfxCEDfYsdDbAfm2IIvNip2njU7G2z7WV/Xx5/yufpc/VwDIN6Y6IZsS42B9M2uWelt45nkKt
FpFYPoaJaQty1BZhX0Bc3kBWlnlYjcMebOG0skbirC1pY5pTG7AeqP23RaUd4ka0exZnud6M3YcQ
QMrvl7YEdBGM33WvE85VAkOCpBRt5v8/alRYTgLh0579A5+5NRdL0iLdGSYzJc9VntMdmmsy1vq2
cj7ziCgU7SdMgL8RNny6nue04mlA5Z4obmrIeV/SFXyugGuxi6Ejn2UOIPMa3/h8aMKkCuHNR4F5
S4aMLPxlR+/Pgxv+No+Vvco4ojOcaa7USHylS5faQ9csyADh2L4eVa2zP5FfF2gZY1eHad1efHdt
VLpb7EkiahXTVwKCMmoB24/nYRNMY8Zl1eQ0OdKdo5JuW10Q46hgA5d/QjULXBjGRV+iFAQd7BUQ
6IZf1x5YY92RolMRR6acHIOoE43Qq5YvG4kxl9F8qkO3gdikEtMcHu9bQN1oTgRiOHC6iXJZYIQ/
A8qrhGN0vmINSe9Kqz3BkJlWlhXJgr5I8uhtlMJdCVlQIhiI9Y7h7iPxNIna72Ub/z6F1alpoPk2
qCuefdlduRiCyQzx+Crl8UFHwWiLIZgHcvucsnWg4muo0Wzbpc3Lsc9HQbSdg8Yz+aBobJ+u2Y+5
Pbv4IQ3caqkSlHyc2t/70S9oCIudnTFFUe7+Y4X2thCwW4SvzMKFMLb6+G9kHqSnwoMufCOyozxu
JUerCNEVHCrMOfgwFu/TXKmOMZwqZhhK68kT1z5PAPf1BAwDgBEO/no7RFexR8hFJ//mF+bJGXQ6
UZr0/VKa2cQOU7dMSwfTJnIThfnJ1jVhQYJEnuIp++70iZRk703J7ub2Kazd67m8GCiYzVDtLc9G
Dh9DNV1fMq9l5ecJkXsDUs7Hz+BA6HrukXA65MH5eBOfPTiXDVoC2SbY71Y1f/BAFclV7q/UcuOE
zwx1WxF8Bxae3igjLdPqSFYmGsY7Fftg/ajkNCXdIMksXuOx4y1NyNJ92Eh6lxwSAvOCF2FtolWg
qRx3U+sj7+/G7eND9J+0+7caiGyLKcyYZTaLmGJPb/M7w6Hzf8xNFEL/8Zh/NGmE8FJrzGMHm81L
dpN68qCh60PjQxbhic68aczH04d9AWZioFDKRbh8XmtP15dEYhqz4vmb3G5CB+pMLZ9XCSnvkPdS
b08F2t3HtNt4YloJtaQZmqx8jqMNwDNiE91oW1fZN20WVFc2FVwCf/YW/8KP4NQQKiwvE4E5t7k4
XBu4ENQ40ru9JuXI0h/90XhbFeUzUt6sNYxhQEWtiN0HqLLnOQKbA+V/QksRmG7dUNVfKJQH2QpE
f9H0n3PTy6NvD3kPanvHbm2ciuvyEXhCdmwW/iMKTXxFQoF/nW4ulQmbQoa+E2u5vG3Xwvji3qOk
GRHKtf/QZuPUKN9IToQxjGqi97aj/xpZZagqxWmfe2i7URZfZTARDLQpNcxcWWNzhHOeHx+W+3An
JJY0+ZoY7b+faaOiHofzVuBL/aTTLeE1s+6cTHDecoxY9hk52pRTnQctXppeto3GBmTdq7jBfghH
9LOZX548jcB+0RtSqf5Lf+wVZQUYNYC88b7IKepUUxZgZXj5iXfA+lNFQphd64x+M9i992aDxzZx
ELhV0JmuGSnrkpSaXCFEOYEt53n21N07ZJb2e/lRZdX4VGKjpH2gK6US46dox7igM0eN+LDNsuqM
L8UAAwdZlHTjVWZJ+65qrYqx8RLZF6Zunj7BOcXZJkFBYRr3jJ7aXhWacDLQ5ZbMJTrrlyUgZc/R
drhDWS0LU7dhvM8JYJwpM6I8hlevnD8tey3NpxUMD1QGVOWssy5nOuZs7snW7qzP7ZLuZY/xgQ1A
OWfFwR/afVPBCcXgRgbM26v21+HBn0a2sjQn8cwkk3tzgXj9hyjkI+VdVn7BK2S7hq3E287xu17w
7V9MNBFwz+4Cie811ruD5jQiZXskwhNyFFm0WfiaZwqpwggvrwqh/OQ65sVM6kIHhXBs220Xit0R
MYMwSFIOgi5KZXf0MEF1Ds+ZACrsXW8CCqJtBCaagbmgbC7rwg5v1Ni9QK2sVY3+aLmh94p1DMZk
MnZNiO9gEBIe+yK+H93PIuSuq/iRyS5NT11kj6l9oSRITiBgX4wc2d0b+PB7JpsY9BmmVQyLV7Z+
OFmI9ztHlk7UDj8mkWh0jhHbvxmrt3mRgEVhEXKcOcPLk6/5eq/93HiKFTD8tK4Y5+/uKfN/mB8Q
nKFDHuBd04GqP6iU+HDtGPIS1vlUhcIyPYVwhK30QiCkJJoXs0+kxNPM3Ru7jIjW8miVgzCrA71M
tEo7HmoaEXvzmIucp2oVNB8+3yq8JgMjnGqqE+JMCXqok7sHA2aa1TSE6I5RSmnE10yftxdoR2Mn
new/fzFNbA7GvwaB/RE2nyj8tQ2ZTj6KAF4yKDV5dZWMp6RiXKCTvIfNeFfgB6pK0uOSvwkdgLku
8StMWEk0AUBTlr3ydl1x4rZndCWZyDoyCci5QTRhgb1bF+uUpWKX/rVCzWnCtfgoDi9IQRRLBE2u
I9VfKn/QTJ4CC+IUbslwJH0UnmVPd1PqcYJZSzgQlr+vuwgz6v+Wqd9vO0FraVHJCS9CuaxU1Nx2
Qq1zwHH0gJTwnw1891VgRM1tM9AoquofqoeADvJRxKI+0g9WNgLpHFfCs7mbDjZCNMwptE0gZ2fc
j4FF9SxtOJ11AB2DLgUi4UqO5aroqvY8XEDf0NWyv4w6fkme04d+awgvMa7GzbuNrXzUBQ4o/Gih
Onjs5fIl12hFbXqKyaWbPy2PComLyq8i392DwVzxIbcYt7NvV9dtlYhOUfjOI7wtfNWiqBzN1mnx
0vb4a+HNdER0X5zXtBoTfYuUhfWfJCPQs56RpyL/AoyYeE8dji/YP+xKJf60uRV7p0LHXqKR/EwR
OlkjpzVswaxLCrjmBatSb0tHhUOBC2sQpY3JhJUotIPGoOpTyPaUeveBEwYOcn5Iuo54tcyZLWbS
VCZtOLIypp+GHQwPwhjX4OCr008QBvRHUf2bzFpGf60yz0O+KAxqq7NEWhNrLjFbshzWINZpM2f9
fJUX+vRA767oJHrFr9hF9UMC8mzjUN5hmaaEHnRfyi94ayUZDXbJkGPrX0MOMDX6P8eylmxTmuWi
27wsUtmpgQ0siQzz9y5pspj4ays8+KOUUBXXV1gbuJ65wbhFBYha2FnO1pYHqAA/g0GSeSWjeDG3
Oda1PytKg9EYzIomxUg0gYFrxRBV+3qm387rnQLvIWG8WKgbx70TtNk/whYMDtSg8NE6clp7SxoN
bhcmiBbLI5NKtJPrZHR4DbIVpCCsLNFHlhtazBsT4Ny7D9VTnJDaOBFWw+Roy3jaCDzO7/+OZsrV
66Mfto3cA4ngEfW9DhntIMBAVyuCeQzD3ygJ9OeObXJeJ6Z07jOjmzVTTtU/ng3wjTuS54786ctx
myeZ99vmN415N9s05BZdGFblHt/XGtpG6psP6zgk7EMSIUkRnAi7WFgWMiuikQWXW5r5wbZy48f0
HVaTKVYeI4iHuaJxuxL593OlUSArRQ3hnfFpwXNFi5qMQVuZSoAeClTXIhMGQ8XLlF6E6GCM5sbW
RwEWyena6GOfZJcc84IhJBtraNTHW6q4qK79oeL9ftm4wbyeXWjgpH0cK5KAS5mxCZ9lJahg3Cfk
F+LLt//NqW8yvR1RJ0upqLsGcg67KqgRTMSLhucJ1DHJIwulCSfsxN8051l7K81rKM02vDFQKQb8
59sLDq2ljoOKRb98B+05Qbu+4qBrluR14lwJXE0F+i2wq0WvyGEQqvPEGtWY6m09KZGjUwafaD7G
t6IyP7EU4L/rZwPXqTUU0LjlmkytMe9SnlM/hVvo8j/lwpkGhH7DhENvPAxLP95AsIPkvcyc3L2g
HGD8TQykI+q5nhkPGsUZu76IdkMU8sdvItRYPhY3yc6Ht8n2lXzMVtrDeSSrQjgiWHc0g5PD6h8t
Rw2olaWwV0nIISsLBgmkd31UyYB1pYkcZqqbopW2z6NB5IfrEb50iO3VK2gD5TtOzmdtQI+JHYsk
DCKJC5ym7nb89WMmmnKt2nfRTFzFh+v7d0OIu6AkZkXHE6L0sGYw4ym8XYdBJc221jzghyiaistF
GlLFvy3nKn6t2t1M0Qt/aWaSL6Fwuoxi1DdEJlGDL4fE24A4Dnl1WNSe5xftzBbVbWcV2tpcKUob
bOEzhS7aVQT1jiXgiOIZTC0aoQzQdV2tlI6+YQsTInuyqPuDRAy3g4pbgLjdCpabXF269y5KrzB5
YvWAS8nwGfmErhifT116r+49bdsb72R3LwVYhT//AHQntP730rrkiFJQdjekIfS+cRAFBfld6sFf
cM1hRPVDqRnMUk3/yE4bu0xEBkXV5xMBgbRgD5/+NJxTw6XV8jWuG8anrOmJ6QCZOwsavo8r2jiZ
dyEjzOMo+z5WVZqOr9WSdmXoDo5DYtWCqIJz36rcRmtZFdSgTI2GmrCisAd3vGQr8anYsrcSv9h5
3G2vSwqZWE0CXnjMxLgGfR9NKjExkFpntjWfBp9imvwoIz3RgHZvSydZib6UCWU7mYTM0Tm7dB0R
OLV2voPIOdAFma/kp3CQQmLLLGvXRh5NeQHP4UfhShWA9uR/qGDi22XIK7iDAn5Sw7vLdiLAgOXh
k6oPVwA7TuAa1VNvcZ2f+U21sXdDMVzKMauTlPge4cdb4YMwgp7hvelV7G5Vmn9wxBPGt2yWNU9Q
sYpNP43WdZA4NjcAJIW+uUci4ToQb06uuwrgqixvuK+KUidUUbkY9xcdn1xhHmXAOGKAbSHQBEX2
r0JeTCvvwhNMiw8d2rfhMls21l0/eo13vfNl/DUEfUTKXRIyqXbbEPmwGoblDAM3sP5SsolDy6V3
9Rn+sRpOLqs2RdvDOulKCBtA1VI7VnaVM5JuOhnJ100VlR+ezlKjtgPJEoMZgzR9bmXUO3ei8L5c
/Do98g9dEBaEmKTQbPDpIc1Tn8VE6w23UtoyXan9dgJIdgF/QPP8nmVzdBWvWCexEqhhO8iIZrdn
9w4mxSeGVYUENZCxvf4gNIZXgMrp7iY8yx0/tFzSW6M2eK/+Y2Qy5Nyon1gpHhhvRBsndzVrWol6
U5NJwTfINgQm1167hVEV0ENyx6S4gay7Qkez09TKzkkpk03K95Qgwjnyd9VglOGpdR6Cm9BMWEWK
Msi+fNIEFBgUuMZHP2KtfS4Wo1eMAN1r+tu82M3Ud1yw1Lj+xbE42Fyv1aS2203DaDFXKu4mjN3H
IOgxEwtNw3sbARH5SwauXLCIFvRZ0f+yIfKZLdfQn+GFnPQzbxiYp/J25JUlYqyX8m/po/GwEO83
6QzBgxLVyaP/eF3hr5wFMAFGd59hi1zwlAA3Rdeye16tZuJlkg1/EHU7VOhRvQ+mo0EbCU0jX/k7
/72rzEyIFTksl4hINys5CFVn9INqrh39ik6Ndl9FtBgfvTzkQ5AhFe1XjLTnYde5/q1VpUD7Ve5h
2khQh5efYZwRDu1km1gdwI2/HRE01SAnT9Qb0qFxohF+TsJ/Ef4ihKacfFLDr5rAUH/W8ZnIB6lM
lb6xIZhpt5Ip3Mz350QsJ1QJsOFVr7VrnDl2sCmkUiMvJ5Yz9NTIetXNCroieG88vN+6JshJF1z3
YL35d5RyY82EZoVFI4ZBllOOwgl6S4qJHehZi92MvTqqvMZXBBchDSp7enmSfI2KaHZJMykcm0M8
49D/nx+qwOlFUFJ+BpAoaXftUUfO2imOLOUJoMFPmPbYTbZSUyxy1/qzi2t23U2S96gXP4cxMYzB
dL0CM+/s30dl8m+1+3SfvJLY3TbNICz6RXPSOzmWHjMLO8U9P0G49okvZuK48K+rEKdGsgesC7XW
/cb3zy8mxNmuxNWyW2S+9UMGVKaBs5Wk1L6QC1GQki5FVnBLYwyTp9YO9WAWWSgqNG712bKSvnwG
9uc67P3kQaXDeMWUp90hCPZlpUIDJ3dH2XMRct9LervGutiluyLpgvU2c0uchLe5IdYlfJpb65S2
g55Ot4RSVlXi+ExoTo7fQvRmM+0AjuBSxB05paIjO8AezqLZfy85QROcbrnbSUTrItpYOqykbVcj
OZQD2wQxe85mokzVTGz1WP4Lm2pij6cC8J9sirLtb2eBeV+7PU1M3Au8wdigDaaDkb2AmNXAHM65
ZtdWKwPLob+unBeioud5DivExYMqt7+6RoWc9HgQFOdiKeVherwtBugJw3uq2EA12FpqKV0xbxN/
9rshT6omXZzjrbWeL/AiDKQOezg8Y3dHIcNDIweBBH98It99XhlLk04KSxbAIeKEBW+q5CdOBuHt
8JYZnL+DPxRWQkL0v1H9zrbvXK1FWKCLFK4MK8FbuR+iscKXZVlP1/uYZSXOSkNeR4djcZASQxQ5
r7NRNHoHkuWdaaZwBihpMoAM01MNRetDaFPk+bCfmA2c6O51BH4ospjgwjFj7/KktSbGICsVuKex
zV2n2GGRJ+aXBi4AmKWKRxK3Is2c4gA1y10nXqAONUVo2otz+C8wrvKGFSoAvZRNuwlZc9mKZ+I2
MI68iWw0NYdUOdcvo4Q3PqSti043Ka+eMf5maV+9Dq7pHAxvoEsh1Xp1TIiI1bX+l0e3ztodFajx
5cjhe4yHUAnwj+LEXLtIe2LAnthTZIU+W2Lo6boTD+0vAz5Gi51Lr3ldBs1KhuQGL7aU0CmbbKd/
0T8k6mf4nEzzRQmBtd4SNK7NdAfauumb+Ot4COxaPU95E5uE2EqGmx6Jn/aGFZUKk77+1EI40vwZ
IbjkYu80tmO75D1Bhgmnl6QPRgeGrBCUcQFb6wpHBZrb22+zxN73WWFGHmfDDsXG8hwn04Ys4w9G
aV5r26ddw8855fWtgojGeZP3ltAjKoGwFIZuC3d6iI1Jiv4VwTdaGm0UleMgX9OxW+ehTk1X8mBA
SR3bg2nve32vW1X/GUlXgygoMMSmXoru5FIIU3bsAOTG2kjZauLsz2JQHtgsLM1/YViptEG55S+D
xoIBFiBILtXvkYvITXYkk9/4y2ROP5EmwuSEZQGlc50Z2xiPXPXBv8iXF6igsYGGUzO0OxHI1uIq
BFnHGxfOOHgNhCJyAx1prwFvzIZzliLWTQckjb/GoDXKsiN1WiM2sBqQcMmiXOF7JeSu/dProTiF
55gpGduIFlKem4CZZXFGVAUlE2J5qa3QRyyA9wMIkFVfEYSjseAintT+ufLgsW7Pr3LB0enOQNcr
NyA5QecU9vp+sZC3ksYV3Hj//h/V0UKCLXQw0kYXRcn++U4qGh7fTQEaDblJXNhHCSGe1dc0s0qn
q6b8n+cM2A6xVD75N33VECcNJH738O/qJf863yUXTgCR1bicoNINKUjViMDxkqWDMOd04bWJ2vzO
ci/mkjasnljmSFtvXN2fvkCNM1hg/f77cNNKx7Orye2gok/YhsDhD0TbuumbylP6UPZVolwZXLQJ
u6jiu7/YfsEk5436HMEyWfoVLgZbNn+eRqE9oiG/zMrJ7EeJqW7lE4Q7AZecbSZolhP2C4+OxyF+
jUyZ/3ukaFKR8Gt0F2BhZ0nppmF0hUgH6pTdQZ7QtyWr3JE/KvA1dk/1zVNAjsl3O4UE3YADvvR9
o6VmTiwCKXqAg5cDGidz1F5Adn6FBnZsqjk/FAjtrq/qruIZOapAV8vIjMIcoWIVXOTX3D19B92Y
dFrtH3N+U/j3MJSaOAxXHXuDyA10drODUd86+DIjWxS1by3QoHaq37LWFQ4155P6cJRtfESpbb7Y
Leb9Pe7ruNL7RghIJkBxo3xM2MG4KS3A5ceLK10HubCZKPwmoUiR9TOMtXOWIKWhAxnKG/U5kFFj
yG9mfZtxFpa6TEeCNH1WOeQWlrz6/86AfJ27jHr2CNdnbOFiD1sJ5HyQYXy0oX/R0wXGos12TlB6
PhzbTE+j0sNfyoMG1y20ioj9uuJHYK7ccLGTLpp6/Ej0ywiM+WDdFHEIJkyAkr6zHZOcObxp6qM/
sR5PS8kS4S3lK9sI/Q5JGizpIqN7MBF96jhvegl2f/eU/CKt51O9jslZ1sJGvpryB1LIXtGn3JcB
yY1LD3j3Jo8lSvekOtIjBM0ftijY+geTBrcE0zEnEo7sjINDkcskAhzNa0bq81NvX1+BpJaKKVRW
TAZJ98jUdMSEqEUTLNptOpLz30AP9EANioppI05eaGHst31ZZ1grtY4n/fDj3h0fCr/X5U7bK1ig
/l6JuBHrt2ur8M3bso57ZtiuBNQB5yEx4ixqA8yXuAYxPb1MQJIok7EHiDknKt7j19UuVlO1Tx+D
7bD5AdzavbQT2qJWXCNbbc8YTUdfAjPv1HgCkW1J4Il1d8IPy8e57hupfXmap86iYtwUma8dwnf2
n+ui3fcl56XQaKZnpzWcXAc1YMqzeiebTJgf4RINRjN2Z9iwBRm4x4KzKL9AC2FWw9gzFldKb/Ky
z1IrasXRHmcFGpvRo92w+jEtqI7p0SKqEXCK0BShnMhxMKnS0PfKuPn8HmF62QPM0ofslZviS9R1
enQ/iWWsPX4xHWNiL53Zkw457uSzTPF/W/fOL3545qT4x5oIavFS13kh+v6q8hCeGN2kTRAi4OGZ
jh+KJR5yNJVIKh+IXUW9+hZCU11GELp5/oNY7fp+s74RI7d5Y85RVMgqJX0oqTTLGGbz2ZU8/KF3
GDAmwV7a3U3W26UqCRfg1mJgbfICidI3p4vJB+nirhaCHCsxnAe9J3aMw6Bou3KYwNDPPY1sEzSB
mOvm2YbqLupNvRoYpQUX3Iw6kIX/Jj+C3uo1q5NIkcrkB7o9arsORA0lbvqmDtexdTB3dYMybEiH
RiOCT26wPZOZstMAufoGAE4BMcjbhV0EttPfSeDeve7X40BwHLLPcex/0TurRnmbw5sdHWUzccVS
dve6IyPGx4AyXvcyab97RiGCSGlpEL1CiSjbLj46rfQ1nApZGECHseJ9VInBIwodbcE92H4eeAqD
Z9IDoyIp/NZa5JfRIjPXr0KfYJ6Xuu2vsL2VOUD42cTOSqcZxrBD4ff0obyujZevP8NGmp2D7aun
13j4MHXsa2Q6FJUeNNrm3PAStwVYGkCfTHJmonOR15XY/eu45Bkl2ujAQDXLoC5Q6epussOtfXfG
7ff/+RRTstOcBk5VmZ02htW0/LFcE/VyfRhVZlJ3lha9aTaMYw1wT1EIFXoGhsfOC1VmhWdGAxUN
StAPmsI0jwdCI+Q4/7zUPyZEx7FdKHPrNxCSBtv+SMu9UhQXxy0Dgj9DnGQE/F+3b0ngUwsl/29Y
ABiKOdqdGUjNsdHk7vztRxuBB+yL5OlTsyBPOHEDy99camHK4IOTJuxvnJImHkAjSzdb6mLv/3j6
nI99g72AFWpjZJC1iSrThev9XsIbDS+1ikFSS6oUK2kigr5z4nvR45CVg3so85RoM56rGPGwIk0g
JEi+GU6dCcbRF6meViPw6aN6qQVnZ68usz+NU5Trd3v1nDvHmdkYUXVW+46llANWKOCcQoBIQL4B
FM8NiHlsHKn55gVMG0PbtKEjBLScKj5vFrKw39DFFX48vUnaoS3Spv2ENfW64ve3IRh6aB/Q/t/R
inSyu/f5fn0wvwL2DQPXQndA9wF+q7davCKhQ0w/tYlMrTJmhNdOyWX3sKhf9GY/f6ddafNvxsnQ
mhYDcLWUcK/nJjoLQC6CxdNEE2WRx2O36DNJFBljrjOVMMWVpwtfxzLTNnI0Pi8sUBpNPLd70o2o
MjLhraJ3OxVBe3TS3fBTB1TMGkI7dS5Nedw38Pi+PCl6N6rEaAq2A7NBwMlHeRMFKlok8XxvAuY4
495MBeTlQbf8gtV8gfI7Q4MBowhVGx94oxB7g9VPs0aObSMdCFEilk51LcIYQ5rLEBYrf6pXzIHh
6xOemVd7afoV6sQkv6zgCCJ08+B8dIGFAf/LOJ5CTjOuFA+iG0pk193m0TubQ6hoEqc6yjZFHTBn
/7olRj1f1ZShV73OkJ48NmL+8vA5hZUfIxZimRIjMLhDzR08DEuzQHJGqzLXhIk5i+xDj4XQzEoD
dCgi52OBHp209rnYqD8ffyluqJVcNaCw0Zid5hvXgDNqgJzwxYn2L5A4i9S+MGCZYmfm1O+IuTnB
oMMImP6ifzzt3wXlyWQZPsdxu96Y4Bm2pHYuvsXXI7yuOGLIHm1EJ6M1h3AwOQ1ayyXBwI8yk6mA
v3aincjMQNDkHwWHXQ3h5OmydL0OaxJJP8Gi9AgC/cexLtNdmoAlj3MdpZM/rcMd1d2QRNcu0svC
ZbSTHFtVTPlzJVuH6I42fY7tsPNvjDwOBozcKPrODiMdmJltj8xsQSQGyFplpWXnvD3eWhCm2aqp
ZKdBArTyimFbMqfbEl+qI45vp3D72/Uk03KpuYNgXorTmReShMR+Z/qBnk9eI1iSbbncCOVEiBkG
1y7Q4o0YMJnfVEOOwo5QCc3NCrbjEk3WbOaQhU1fxU1MGeUHkLD1Xpw5AIKeVmv+X/rJHnJXnDOJ
0j8ZA0Gs8z58prPDLYNwWspSta8CASqkwQiHh9e/JwJgeH8KBZav6fAcUgICjbOGLSzJq3mAMN8B
6fBwz46wqtpJmkQiHNsAecuKP2NDgpAHdYopgqTS2Datf4ppz/2tHMULMK7JTMUmmHskO3ChwQX6
BFRirErIgTbChV8apZTgTvo3FgQVRf33QS3IakWCe6J83kdFp31elFJdfzoqqB1a8hkMguDRp6yZ
4hP4U04cPvpXHOiSaxp1GLSdapkIEr1VlIyy9NymxLlWNHqHfGKflFOVf6ZaVBogcTerl+gpbfeV
iQhhzz5w985/+O9AnKTb7Q5yxDlDG0TQVV2S4WiXTdaBCvI6if3pRGdEoS1weXXA5krbf4nKmbo9
wOrsoZExyWZYcoW+UEcWT3oCcNkFXKwi45dXUNzNWYyAzHn9gZdUklsL5j7rVmn4q7mM0VaV9fLp
esDmUS+X0AMtZDJn283FX+e1QnfTZpw4ichPbwgMq6cnXaAVHgzTQCvF7fFILEwbO9aV3FDMC22j
9oerToP5pTsLengpUnlTfKfi+Hu4VOYpV2lmsg0/DruXRet41gJRtHvYL/TNYN1NlRUPEdTByrxs
XTpppwufjrz/YqpMddWUkc7avUmRhmMJwp8Pbz4iqacaHrv6VK2CvnN9twMMCaRlyIAkUxB/oqXG
IDpgLgfOErfTJ2VcUbPZP6FjJU6g9KPzkA/daj7tYrcrvowGUWph9HWRfhFfrx9vLqWQvitSVug6
ZvpwSD4WYk6CRqcvEf2j30k9/SpJW94LrxAiGCNMQldcs8fx8nD60eDrqCP+XQhBt3ib9n6GmwvO
dtSAczRKdSghqr566+HecLD6CXtCb29IeEGvRMF1hbw/suoKF2yAzrtmbpX7SkOyM7k3WzsJIN2H
G6NdeGoIeRELY7eTnLCUVCYwnFM+BapOXS5E4UAmyiBN48Zq0RSOfj5YPd2Ce0WqQbwKZFayd1A7
VnMvpAFjKXzz8Xdnp7MnyqDGYOVPOQLH7WbFdEMXPE2kf2rwgehuXTkfcVRm5nW4qwNhIMuQtxSH
dKBmS/nxPmOHq08SelAB13RT+yr8Md0CfPRJmEtH6RSn3pvmBm+UC7UA0YLSYlnXx32dIgnTQw2Z
TlMS0vEroHbEMbBEBBiiJreiq9u9oC8hLM9AiJkK0bbu0goistaVKPEn1hcyl5hak9uxjvAHeRa4
mPWi0tnFNgefZDUzUTUsDdTBs3C5d03/LUYJjHB3KgmtWw1nPCypq2xsbedjh3tXJMbn/qM1lmpw
s2RMlVQk5fzaPWLXb30EVIeLBBM/sS1/IQ7UgnUQbG4XfwJY64PoyMOOxLV86jpS9qB5oxTjJYJz
U08dpMh7WPqc0/wFj73ILCcb6T+FKAdBaV6NA0HRzp3mj5FDVMojD+42gJjslXKo15eYqvVTE5hU
5lr64ne4krnxtd1LpTotGhtPdoO2Z0T/VqxAOaeauQrrlDK2pwYj7pfQAtB76DG4kB+MPCzq2ODK
/xKyOc9nBQE/sPMHhdUoY6jkAaIeIxnkmoH2CW/diTUMQPBtgmWLpRPA35k548/u+3RvWNKZz0Y0
cTeHgcB//AZIym0FLEO2xNG3wiS2uqzG+x46ggbzHxcIBlDQqHaswPDoWHjRk+vSz+PKT6BoP8uD
skAOr6eeoGid4Wonq/KRI5pl4tGtfa83NFeEX2h/z6abqksBBi7fTCy2r/FeW3ZT3IfBFlQjobzf
PDQPTmtGWoU4NAMf1WZE5qpFmdoFGbwLpkNL/E4AgxuFJ78FvcCNODQRtc9/RXo1OVFQSRtUORg3
th1oe0Her9djTBR3KLIMEqlR+xTbxl9fHxrzqhCBdn9ClEUixg+Fapji0QuDGjwkpdI6xABl02kZ
pb171sumroiiOR09bWMVd4eXcnWTYUVwSKbNfA+19+5w0PDXip7NJPpD8JrXvBFyjLqzh+PSvlnR
iY6cqRDdU/KkF/3Cpar6PmkqnswHKny94nYmsEpO2Ool9GJIhD5Jy0X0xbFPR69nfio+FzyWXt1u
qWB1fZkvcrqG1JHOLh6M0/2W+64kjQXHn8ykC7pqTNqNHRP4AhmGq8W3I5K1hYL27AxeTMColaY4
3PGrlrGqlhGsabUyuXFImdbCU/zG3Qyrg7jfdHZAHNsyuTo7mZA2TNi1jthy6VjYmMhQ8sTE4FYw
FjG8TViqq/WcdnsV/K/T6vfmG2ctng+6HFF6IlA77d6KOH1YPQbEIik3l3JdhoKh76db0LjPxURU
rK0icvoDvCGrvIandDZrNpvPzMP+UZ0VnTb9KXtag0PTrm2fEVDzVfnWP9N/SdFZ1uTLCT87bqbj
etqOxDpX/Eb6xpoT6Dhxfv1neC/v2Ow1CHYpkV5CtyUqHa8EJG9HJXScToqQkbi7vjzgY5rIfoHI
4b1sXUGDYFchF4P6uZGg6TawqYyR3bwi6xRR3FPIEwbdIZh/yklqA+fAKBR44YnT+6WoY3a/Lafa
xmSbk+k9s7UbC5f9j857FrLQWRFq+8bLY/jkQDTTUT9pNnSeGQmggKYJUv5c3jR8a0vQx2jOd7UB
qpaA4F6kz6ixtQ/5zqXW2IoASmO0A2wxpoI5EDuD6BdL7jK/G8rLlVLPz9wW51mmVNmdqOjyvaKK
qorD98kP0qcXoWuZK6Dw+/mwxx4bcMfoQ9PRcKTjX63YbfVvLp/45vSSactz8Q7w81eW5iLpDSbx
vE2xN6eso+Bm8HiBILGGufxH5yS/ajNDDU963L0SLW/L7UYZYwGIVBFyZvVL2XQHf7U+0SMUSQnq
elXcADCjTwcjEb2MJTYnRLdeSEmLuhYMZ2lrCyv9EdFZwUrtFook41JuiolA+O0Umu+feECdnihA
XSP/2XwapYj2FmU1Xec4xT7WntrZ+4YIMWxxGHq2l0tVm620frt883jeDot1TVRX/43X5p7nY77k
qMd1DHxJjPgi24BiC/34Oo0mvjO+lPBxqeN5OUiPkw7n8AfhLHujyptIAtSt4f623esW9azkd6az
e9IPr/y6eNkXVhxmz95rjyaJzAus9KQbr2TQ47BnncE4cJOmOFa3BdL+XjQRYCPMBvfPMojyMYTN
k4cswwE5HqP6SnDTDpEFGT7gdZV75uG30H2GabtmTaT9hUL3M9B2NICuEqc8ZoV+4WoAoGNQGhrr
RK8aLJcDrkdSfDgFTVDs2ZN/OOUUJm0Y0vnZsLnHGO1x+dNnNmrMoEaCvt1AoyPpZ04AgXMGQ6Hx
5wJqMS8DC3aLgrXcC6aWZd82inDgLKKzcfYi+vXZdLKccjCNezPcgLH+e+siTN1FkcakjI/ggZ/i
KZs5W/IZTveBigmZNLR5iZfpwQnhZ+UfR9bnSO+tLGbXPLcx6L/AQ+TjFyBJD1xsTEn+m8MNEoEn
Uv/hX+oy41PCxU6/enbC6vtZJnCuwdXIoPPdY8AZKwp32H4Xom0lbBF5+IZ5j79VDgajCK9bycqa
NDRwB5BVTUByC38tlIvqS0g9hEXHASYzXWp2lhYZyezNns9Qi6NwOl29SnNnsMLlv6FaSeQC/N/H
aBQ/RpG5QnIkECAzCBRv89LRpdRd/nWfJiraNEzCOC7xfC15Ws4PzcoBjaFz+WZhouvobDxMXT/t
N4RwHfz7bmpTTtUm/aCCf8pnJBCSvbzww9N02Nl0xp6SeG2JTz4CNrei5Y79Hj0ZZhiEJwWwsltu
wfJks41FH3FaoHFa0YCMQ3l4cN6tWpjoGTkUU+W2vQp+aNTy1fZxsDnl2uzMEThgY6dSLGBcsz3O
Ng8it9tXyoYzVrClSQ9lpC6fnt8zESLagJprV9l8NPCOpivYbSrTViyMdbS5eSOEBAW5LTb3p4eI
++ZFvmmSW6qZX5B/qwKlW6bKVbccLGH7NWcZ6xC7jUIcwDs7NhNJtNmu3u1o9kZA4FtIH3/4G8HA
+OlAny4tDsE2VkAM0HqVGuAszR2ftfTwctSl6EicaDJPw9HwlPtx5Nmy6RnNw1f/JdEKT230W1A3
8QoW5RGjuB8StpSQKSbWN0yiXq0NX+dKbcJSFOt9W6AKdsUkR7n7DZ6ONsAZwRYY4KkGt6LxLqx0
03Z1HQNhCygFYsZuklz7JFOvc6k9kYve+OannRjvjvLU6D/a5JM8txJ6qvpaOTeKzOXCn9qUKNKL
eKwxDao4Ka3ycAhiOCRW3haxQ0h84afkDd39mltM8djlnz9XibJ+vw/8a18EFRSDKV3Qs6cYoQPl
XpfpDs4ibQqgHKQI/pxr1GE/cFX2BkkgcRQrbyKvrMZvnOpuvC3SR7OGaQhX5cXbMLlcf53D7SFi
gnYTohiQ0pbTEVjYxZJeO0hmxsIJ/MR6TBTAR1V0jlbLUhl5EnC6BBfzYMyqf3JI0kMln21WtdYT
IycLO608K001n7KMsMiUBIldSi9KaaU50N1H54grBGcqjp6pPse9KIFxOa34nDEa7V5UNvqHu96f
FHno2gItQDlFy/Vqe64mbGn2iZ6GjyxPaDHg2sDoOE7UKL+xTdAlIuGlL5rNvbjCAnGgpJDPMfW3
Wuj+Np1PtngNfVANrqxGPC01fsrdpDS3XZYjBvAZpkNFDv3uQ5Yf+YGb1366OBnzAVvsCk5USgQr
ETa4+2MlhuQJzIQSgJ7+amurkdmkcinIy5CqLZT+EYdBPUnQsC31cGDIjPTmxQOOsdWncvC8nfer
MXQfZgfcwIhPBy2hkFRLDLaY/bCnkVWEJ7YKjksIJ5kJaJJrqa8Q23gGm/WqjHI+oVLI22LRJNUO
Z2zES6cKCdm2N2XJVRGxMANCrH7myVNrMfWdDgO1/cnaXCaki+vr2Od58ZdKF0VTeSS8QIEW6t9U
hORkTo40KxbX9Y8CKLZD1X6j4yMmEuHM4ECErFqpVEfRyVCjUOIal+Nw3SFplczxQFcSZRumopb0
sYXbVA5MghptsEPmrOzZ+bKoD2dka6pI8uKGdn1MZ9q1uNoD8abM7gwFQtUHhQ1x/PVKsMpHQAje
lLyL7v4J7vSuMw5c2KkLThKWSAlOSNbFOWgWqt+HkoglCg9bCYBXgqSzxQ8gX0sundAJQXAEKyRj
BuDk+n6E2UfgOOmB1x1UPh2YeSUjuKFlvRoMhcbHcH8xfV9d33oH2D5si0ixIwudjw894wAWwjPY
YU3nodBhspdK3nd1D+J5LTPPexAyk14ZWdTp9QZib9chwYQzl86HqU9tgHGYmriMxlUZopkwdbCK
QUS6mF3Xz/0REsUqH7sTaQq/+qiFbJvkSSiZZOXBeGwrNZF71UpIFdofGN4i3Gy6e7SVBn9be8RX
3Y43kIInaHiiS3WhDa2qbzKKA6X23A2XOuRZw4L4/dO7koGaPL+ktNFoIqhc/yluZIlmmlU6rEwK
bO5OWh0WEvqjq/I/gCo7kCvBTUmdRThASYAdHrE35+Z9XFIsAtuHi2th04IIXxaTTVRsvgnT0IMi
cu9CVWM8lQiYi1QcZFUPv74byU5fy567+gXe1DUXNV3/0g4PAA9K2LxWyzgWlqmIvkegVVRu9x26
kf+uAB/09T3Q7TLdVaqcxd1EJcR/Az7vSRLIVRJK0sDN0pNyk3W1S4FYNw+2jmG9Ju/yC3Fo5Oun
U4g4aPuL7qSbcsYx/G7cseWg6lu/qFpce1tM1tCDsfk36/hndFbrogDXkeQ/5QYPh1+U6XZGwcCi
mgbZ1xDwhUCJwY3UdkJPp5xJdUzBSz4RNRN6rjMyHpFcZpgA7aAPXHXeSg8IojKFalyn6gF3sxMH
x3LblsIXtLzw45+tpiL611C/jGUfz1oJcQhd2NljbRjXllXo8JhFPejh4yaQZWFrG4lYph5J/IkJ
Tc7u9M0tQJsMOr6YbZobP2MWS82pp/2Xr2//UK0A0k1iTN+lbF7qWftcLYS4xEimS2x4O9Vyxbza
CyNPojaPqImSAE/g8Jya+no1AfU3RmLNgz9JixWp8sv0QiiBfis2+XCuaIOWO19XSPcDMfGpWfua
XnxbrIvzrmFvndOQ7wMPnmbEVTqlVxly84f8yRKDokPYE9Z9Bndr02/LT6w3BlCd3FGB2/HOBhJC
6xU0tY3dl6kURvYSHmyZC+6IRdKRw8+W5l0KjfoOzJGaVEmNDyVmQvmeIICsY9+MQdiTvRn1dxxy
OJV84Ash7pY8kHSL/0k4cEBWTC05sAbGqQzsuptUA0UIAB336sCpRTLH+OgJ/+jmEhTjQaTpXEGT
i2eZ0GmwUxPsolVOmnlmupeZmHdR46SuUJEqTYllDuXYo1WhEVEDVV37JL7LIIPKzc5cyn8i86hh
GX9hgIMmESU6kun8sGRYotoZ7MTyxIz6zdRJH3pruFVWGAlDq0kjWkr1ayT3/BE0F89gpMNtvr7Z
lxIQ/2GMZx2EKZDPvhs2/GAXBQEj+L13eLL9iXZfHCruOLEc8LEekaP+IJscE90KOBjmed6FpgFh
ncTRhTShIl3Q0c1l2t/GXRGJSMddgRQfYGsDzGhtkd/FLvb/yOA8ybjz+K6yYOLsPK6vNBYDG9Xr
pMtSflmNpYugyTbKfyQCiCiINHqk0UC2BKgJa4F7pYKiA94qHDWbN9C5fwGTxqa6CpnxFjx7Qjq/
7WHA3miQtUOgoz/qLjlSyirCw9c6TF1jSvMa9FSYSIzZci9XZiWSBTLI0K09BePIIDOPBzR1gCrw
91cCRZcq5dF0o+grqnbS/gX4UZnKBBfUaMSsASMNNn99rSgQO/JbwZHusCpK69BGyhC1Ni9PTgK2
KT+KLlClMA08u9yyAz4x/wfoHEyUEJ9Vl4CcGNpjv6vh3gDtKYVawb2b7YCR6KX0N6nt0J98dx+c
kLmCqwWa5j9R2VCxoYxUubwPmRzddYEg3O819Q0Wg0S+h7JAiMZqg1Q4OdFS4jEciCVuSEEL1A1i
kjWOpYNgWGpY51RszSSQXkdWZX5A3bqwGl7bzUpdobs3VkitNqD44TqjnoRP+gw8CRJ051hVln5r
SfzgUcedzRPPwLyarFuWlYFTUPPYS2E1dVI03beCFSq0Wu3Vd+NhNSMb+HP5bRfUhacs2cJ81uN2
Ijhe3XtxU1VTjrU+45W7KszwPMqu2PhtPBQ0B35vm00etSaEgFKpmSqQboA6KzC1BqJ/KFILpAKO
NB4OL8j6sk5lk/71sX6SkhfOcXW1Xd2+Kuwg7V+L7yH+jhZZoSsNpsNsJplhvy7S179F5NgK2XZu
BbZnDY2QhCGF5AQVSl/qJOMHCVqIO51sRGM9F15Ub/InruiUOFLy+adzgNM5mvW5RuO0UiBIhcq/
+MbpKth2nJDFJvvdgjGcRLZ/jV5dGdNSAkbCZlAo4pEOh3tEuxLmiKeH9FGrgydqPap5/OzwAtfV
VONuR0+8XemWk89P1tTrxfiSheLpLUZXgfSZXYF3fqi8wyQLQUY8xD3YRa+s4cJGTrPQ03kXCoJH
pcw5kjItZi3l5hLa+IErhgzYmhR9P5xQO2c1weOLm3GhGwu2q+XNqIZQONa9QvdJJx8XuOBbjTBi
qPgALpsVrJI8oUUsC8tYvMrbhy/u/RXttUs49Pier1rj4BDE45ZD/NtUjDW9WDIHIl4bSGoJ0+Ix
vsZa8xMqS1O19NGgEB1GAD5dMDvcncyaAFUFzSyQGYMyF+g+6pOSSVsIIYzOlCCUNXu+0fTLvIjh
N9lr7IG/s/QsxhkDgjofD+IrtcGA44eMjVb5DaFTuhXSe6seox7STHLOpQQltLJbYIfq8WSzS11E
eAXtZqvuP1emgyWp2QjcvNBMO75pRV5yihweGqfmTiiYdcNk/ZOwjVcTLVFmHWNuVHTB7vM73917
MIqNUcumuoHgicvx2WgqrM78vFnKICYqsI0F7f40Cj7sIcdo7/b8qORUlSSMl0/vc2zLMLWSH8mP
WgspH8S/MP91aTUAKzWTvzpkGmAP1bA0xYeD2waoAPwyrtS/kzsz4v+2Ro8g9GeFfYXG1rt5b7mB
L6BOZ9SeM/od6j5HFIrxbKuidDc8Hp5OVOtvIzCLro1Hq+MpR1nLjX9jB+/X8kX2SRN+QDDU+NqJ
qu099ymAugh/gaWWXpZbUvD2aLEqWfdJM1H1QfbFAuuss2NRpANC+JDNQUPZ9HDmyDclzZ0lSal5
4LvD4CWnVdtptrPUF6/m4q6RR43Ks/vB6UhbpdWuhpKP9D4mEEfvSIgSPUMOIgkGk5gRwLRzhbsf
YRArKjQwrqHgM0MZ5ReW5/oP1nJG+ImvjROnK3CrB83VohYlfGFOttgARo0DoyWLADLNS7YXlfvs
KC6yOz2ilNVy1Zvff/8KPTHkg3x/XWdwxqe3RAt+YpTr0gvMVilUqBFna0KKLrk7E9hGuJ51OW+X
dZCG/I496bzqiqyOE+t6hv9D9FfTREVUOJ5vPy19RJf5PEES8tAZ/xU1c3wEEMXA9jyDA7Iwi/e9
O8aCxNT4+yjchf0q0bz7vmOCll118S5M8/CP6F6DuyUFEeiwcnjtSBtxmSoPtwtbx+7TZWDtjVhN
9LEvXUwIiPvjp+LEz1F7veP2H5T9f4zMMzX0mku0pNo4lqfOVAjIGwxCkhBXpKLnzRwKZfTdji7c
yag8NonswTIWgexQk9SaoQ9w0nbBrQ0o1OssBj6k71gORDSNYw/9sGxfuoTB4lenY7YNMgshrcEU
GmX/mfRKZBfDBAcRofIpBbz1W4L1jOEf0e4F+3OPizPmQjYDrOhi6aeASJwGQTtfqKHyt33mKid0
oyO7smEdJ7jQDuo18XofQtd36SUWA/boVj9QvlyPksnWNUMQYNkFEIbeWH+dNjuhirxjduQNLPO/
QUo6f9FqnO6aTHiqDcx7NiVF4u3n2VqIBiXAeLPCRV/i7SrPSjsOXXL/KaphlsicGFaVFde99MAn
XewBATUsMB8pU78DWpLy8JJuS5sDdCFbhEPU4iFcISmQOkwpVVnV1Y6HDwJg+N8/g+KJAIlEqKCK
uAkM/5hSRGmeNZNA0liUojrVuKlapi/Er0wvX5fcINZHLV/mxS40G910ekp3Ecioqz3V8TqNzSHp
p2ip/JWzaP3x0dbVekp1huuOzmRppm360rhSEKk4R0ugbxVXN74prcu+l1n/GVcLHWjL60i4Wk8l
rH/hM6H98qp14HEnXX3fAx7X8nctvs4NwDVB6ybCOuKGYVRYCz5XaICvMQ/0QIdmgj4WmnzL6y2D
q1+/vd46hKU64J0X3HmYpSUEbSl4M1o0lgkh6XqeOxYXYlqoyVbqXpvWeF6pgwjfk53DCFDjTsL0
ezwKDLhtjNKpSzr2NtQmCGOLvp6DAsi43YVbICjxqM2o+EyciivBxskWgsVkGOnOVgfESZGT6CI7
Lbc9RzwEyunDyxyJwk4dpWdC3pNZmOyBIBsGMPY75UrjM5/b8mIcuK76HS+ZODCQq9foJS/mfZ10
bwpVHOaT7LL0QZxyjqdC0j9w7aHfzttCfPvj9KFPPOiJ5krddsIPW1dwnSsvM27fUOSyGh86xJIB
AtLoF9wSNoIpzg8pWBNaAeUzReKdsa57D8kbuw3hKTsYYK16EDC/2X3NUu8wiRRlYb7onloP2QDj
UMH/NMjdlbbE+3NLsMjM9y5I9YmCeGtClBYMZ62Gfr3ihEHT+RnZvj1rkUz9swiAUtaLw7LxzES1
OdWVbppxsX4vv3VnP/SAn8W3vUpjh7mNAvGe/UBN25koQcT60u7bv4Kink4qORhKlpIIfnlIdlu5
Xb5dezMfdIT1twRR8Pgf78Y9tuPR3mHuvglfj4y9slLlwTWH7fqaYXIEQ+nayJ6qMDLUvMmYJDL1
mrFpaFM18bNkNMRzahGI2T8AWsZGj1YEY8u4F8n8CZP0EIXdRInn2T6bodRhrCTP3M/sjXXUm2Ef
yuC2HCpW4czuiKVcHIvThlHpoASxE+XRSNqD6TYDOx8y+s2jO0Tj7qrAjeqYCZlVTXZKqXmWgbTO
cRShGxPudPcK1X+1qU/9CuoG/NAmJ0PHuKFm/n8DcXTdCvo9FwWZSWzuayF9Hb/fOBLYG/CmYKxf
0zNjAEBGsy70XKoW08mxvfhoY8pgi8XQGh8iLt1pLKfySEx9W/oEuYYyIgkd6hawpPl4S3JaxeDG
6eyMZ+aJL+b6x7nNEUNnDaNDzmIhvX7It6kIpcs0G6w7CGoXIJkhaZZJV+Y3NaJqmxiVAWm7hY7s
4ieOGKvL/7cOAJiZp/aW7cbM+PIh7fp7c312BuHsHp8jGUYMmzn61nukpXJRvXwRT82MJy7C/VFk
dpdkn6R5fe8JIrD7EDvu7bulcys1GcsvbD6YRzgX2j0Y5Zk9LsF5I78h0H8CTLQYWTxHg2FOE6xv
jfY7J9cNp9yU51B/V3tQQtfYImIrjRxtQC+RTnNOpHFRWiLIvZt2DMiiiq3Sc/HNEslw5Touudd3
t8Eo0NdiWNQuqzGlmeRLG38dK4vVbWjYt4jx7HOI5y8+gN1GJPl+tXAFgjxZhakT/2sAqxuXZIxX
PEc+0DJCvrbgIXkbdvTquALlLZxCwU78X4WoL0D4tUsUmCKN5SLfkYE8u4OlJxYKf7JiBiyaQ7Fz
fI5Bhwnsp3dGmTWVOiBuTozKM//Ll6KwfEZMXH0d/WF8mX0B/7021Rf5ML54uNuyKuGkdfti3SL9
jDngRqdIbyE3gcRyFy+ESAtxrbcKzmCHEvDHk4DdSlfccfM2vGdIlWTj7kirAmd0nWOLFJXhQjK1
1rZGmjsg23T8mzL+Z1YJYz9FKmDH4wCnNah6oWqshAB0rYXIp4DYWzgc5q2AHTsFBBDvpKwizt8h
7ZX6Qbk8+yE+Kybs/u0piJ2a69NoT9y37UD38ILa4ZROSw7n8dYzO6U0V8IO9QYWr5PZ87qtXXeA
Wq8SnqMZx+WWEq9Hr6K78MW+TF6gzqDV9wyoEdaCOOiN4IXPjQJVHDRXKFsMSGkhBeV9H4bKjqsi
zHBycs7WcdvflXBwd409yMChd65Ai7Tc5mMhRZ7jUiRP/MJu63B/58s/RXSKTc6T3LJiUBJKgDNv
ZM15y7bMgb3ZNnRHPR5+pyLF8nlnsBkwaoZN9qgsHVBKk7zUgA2KjjoY4ZMZTLU+ZwymVp/M0h76
emZqhA2Q04aoQofDEO04Ucgad5dw8tWScIjWbRfYdoYQHqkGlJNiamOwiUxSbzdjfH/JFgmnqnha
vVCB+2W/rhgUYyj5dXgYomzajFsg7XYYE9vs5DgtXVxaVT2Ir0FrXO2PtwKLfIafjZVbQq7nCtvE
6iaGpAX/TmZnYVxXemwFHC8m1v3h4kQK4Vo35IcRf2cWK443g16DVXo0/zhTXvbhzHFilmKAxAj2
My7GKl2Y1FbMu8Dbi0B1bxB7+4n6vIaw+bZzsX2f3Q9tVOqG49HXOjIFcIeKGhzE5sx3BLrVUnUu
pamKNfLSj1ohs+SfK2R8dxitvhyXCg4PLoj+5hiuBo/Ju0Df4cvwUmf5VvNPKmEMg6LFlArDiI5A
ICy+6Ll2zEjkE2brhv0+XHsyZ0UTmY1urSVM/EbBsGZIrVjHEUoBGBHwIIXRR15AFJSNh0c72OUZ
r4aoDGdJtUNTve+9HT8RYQK8dDVcfBfQgbfFZI/fF6tx5FeenpTT1CAtV+9i0CIJ/QqAIpKx/AUu
Knwh3L5eAg760tGbjlcoSiMs9hxIyvvyYNM3tFDRvOpns5Jenvl8rQvOXj6rVEHgllF5Ye9qsb6S
aE0gcRpDMDxeQn3D+Hqtrx+tbCMo9S/goGeQRxVukwe1Y/yMsNgF4jRp4Scm9oQhtHkab8Salo2y
fcqgJkYjHPq703vJElwximpWq0nHfNQlsL8b3tarojch8zJZhvT2oQG0AYy/ZU2G4jP7PM61dUZE
zr4OotRPv4OhbHWhFySXi4ZadtV1bPAZ7fC2MyKouzwvD6fjxEXmv+z97R6HD/gLObIUHfX4vJdW
mH0tKTJdaLQAvaLYrrjo+TRfD+BXCN3EaqOV762V89chZ7Dvi2jATnvqDnLpdSabitxT2AeAfLwS
8Qelg8s+TXPdeFv3nQN3icb0GjSbMacl3RLIpUnL7Z+f1symJhK6p3gC62fs2F6oE7pp1L7LIEZi
XWEqLNBbiOy2za4mdSGzKmxyO+O5TDxca0xutUQ3jIpFwAhoMHbT11t4gw9rtwJxjjX6JVdm1158
Hnij8+ENIHVKc6RPDsqxhGOMJzhB4BYscXqToBAoftWAMz892F9YtwQzvLanZLw5t+NWutdTVqgD
WuuSNTBtbO9+TDcWo+53UMjKCkBQYWN1+m63fRF4boYBIoAWMSdJM854Qxsfh0TUDvK+WeobnctB
kM8nUUKgJ5B5I7iYKF3zdqqYD/jjUSMWJSsw6jDdrRK+vrB8sZUsJ+D5WIh4WJ8OibnDZLXD4Qgr
yRhzm8SqVuvrQYw69qqslHxMTywpR8L8j/Wn8gaKwZBf4VJkMhWNns+hLXQQxVff74TCzg6Li2vt
4/2VSEBlDzS59JE2qMVgGaxL+DWHQiDmQ9JQng43YY/M6OM+dCr/DhYpimnlGQ2fHturGlrOpsI0
2xFBaSh1eMCSibMP1f30IEZ0wnhNbIFO+Sgnj+XDPwERuLrkS+GswYwAEalLGBMFL0x3TKrnq2fA
QkffproEW1wpbAELeayf25zm/o5uaCFNAhQ7DFoTWHpuIqJNko2X3KOcDGf3Yi04qK9P/5H+rP+O
3pOzTjcSz4dXyLCnjUDr9cY60kUzMVxhugGR3lE7mHcc1gewNRL1Oxj7pysByPTW8j4qCYs3UL9a
wL70QS141SX0RWf21LuTWou2zewPbtVKl/SjH4DPFR+FmNF6I87LZyDhHh+fg2TTNqW54CsHw0ur
Kne9LLmy4chV2Ec4Rl1z1HPGyezt4VD9JI1olnD5gMXMUPhq0jZljrx9n/9BiNX4Oym4mzY/kF5S
B3UDhfFnLWIM4w506AIURVuX69hLzqEzcJoQbm8jgGYt7KQcpMvwxUsxLpAsmYTOOG5oW3R1M+8w
JCkYrLbZQFqyMKF2vcv4DrT29dR77WcEBxX0rm9I2jKa2UA1oZaav/NZ9DfNNJ3UmI8BK7kinqfV
AqgjFVk1Q5f34aLZZpVv6eED0RWeeqpVTUKfjyRyEtKJ2K8j/JBjZzZNzE+chOwPFExBab2Z7JGY
chNQJd1CEQN3MlGDl+M4IwDeCAg/M2e9YLYkDXzzpVp5bOfjmqLW8QeDSM8W7gQLnHcBzFruGP2F
KDpUe/inqOIF8rdWQLdRahPiChrke7baXIeXDjOGXxGbS0el+a57YBBfgYF89WfppBH0T535vbpS
rgs/rcC/gTt7Xt84fbR6O7vXBDeFbuSNWcAFdZ6VuUrturv9UqWQksGz6KRcfT12+RRGJF/r8RyA
8VYvNQZluU2qWG4FIBqJTCVUrj0pBWcdDmNf1DaeseP8/XCU7SfKZYCST37hKmWPt1G/6o+d979t
Lrxs9d3EyhdgmXPjtMvAr/g1HFyBvbnXp4v8QxDw9JbKdGWUFVCIDLK5jkZNt1K6FhD89fmeO/ET
iDzsVKLFRRw29DdHmnlruWyKSgl2VPbB4T4FV9rEnRp3yTdIScv2YtvikfWwMdfXgcYRRftLbEqJ
IiLbDcO/wlqiyZc6M40wdVdSUG0DHordt4Y172nk6XpEV36+1aGoGKduSghdvycqRtUuo0gSrhAd
UYJFZ24ps6E9HZJgqiyvKWzGW9wNIZ5oqWaXy0K6Mq9zreaosSy2KZmFcteIHVyXW/5s/ABAm3Rx
6OM0BQR1Pr6z4Iwpok4+3Zm+0F+vEaSY9pYdCeqYgy7IxPaGZr6su+EZWGwlPThb82HrSiNQQ4lB
4ocEPc56vsrM5GXy7GRDZxEC+CXWarn0tX+ItmwhfdHjwbkZE3L46fB9J02VN+jcu/pLqZ3vWRYE
HDeQ2s3Tq6tIvtdjRnD2/oUNr2+BysQ/I4yyr2nryM6e49egJINDr5cf9u+IR81qC3X3nKDBYGxJ
9kQVcWvMUXDbB8iAlfiQlylFjEUpmi5d3q10GbOFH6901Zd10YHkrtHfpb/7uWkEnN8rV2oiYeTP
l98dNT1Ccbsv/hiRMZs+2ECrJah475HRb4Oc90hYugbVu4lX+VQZmGrpkVFyzGCpTEV5YERXJCK+
zHUkSQ0SHnRPDtzP1ajuoSs/8koR3IXCAqxGf8zqkDfe3pY5AIUzXk9NCypmDHeBgwoM9wxUl7MJ
EkJ4uJU3bI0pM44JXk6bYP0cVKn3dbOwsGtep2lvMFV602NUzOkOsGgtQ1D5GnXpGXh/Hqy9sB84
I/ysRdTcOqIDMHB9lQ4iiJbg88gkDl7S2skYuKpiJJOrDNtUagkHslgRm+BVzETNpsWDtKDgFoCP
kwhynnDM022zpHSAhETra35oO6ReMZIiM2giYen7kjer5kaApih7oV4+3cuSHgYiAxNhpWKeJmBl
01Jf1EMbA3L0/DCZ7m20RymMfRpm9OkWZ3U63yvG9YwqHv65sUtQXtQPmWjTnB+D/2EttdpNjCvi
hZIwW5Q8V6BUBLoMCOiDj34HpepQukQGrUyxH2YH2AvApCAEbwN3ozB7gWb0XhiUfP7+UHWxN2EJ
6+xQbW17lyuSzzdL8XpNzO7A1mnZZcSQB7r0Z3DGEaj7C/H+HuVMAQ4CBQLEALfIbN30mDHGxc3R
FQ+z5zaPqMj1gAKDdfJs+D6hxawntGC5BrN9N6Ke0dqEcxiIZk3BRBfq5Y8AgB/1Hwgaeld96x7p
G02/xe5nFFnXo3G9iGRDEHpDGH37H9A2zny0B4WqBv0UwFcNSPpXYfzlU4K8vVhI2J3zooaN5ABs
41VYP76ANcB6Xo0R15piFWcupPod91+BOqVD9dNaju/myjkE/dC4kdI91bIB31jSxJyHK8oDce+A
8R+ZSaQlqgCNa6GxZv4U5/lxBhPc8lSyxtPh3sPpdOOHkkVB6WlVkPszl/fK9meJjpsDywIL44hL
X/qiH2+6K9h2LdJB4ut86JEv1abKEdTqne0kbxHT5rWm4+bU4Ca/INR7FItX5p4k5GPdEc1gxdOP
ukYSHbquR3wPM82f3qJD60oV+lcQ2jYR7uaOQMhRF/8R+dRLWZSeGJy/7OJupA/2hwSOXMhWmlX7
3urdssSUKLUiZgKvHQf/F2CSh+gHfE5lrL025tY0qmenlT0ARienHxSvxXQmipoL8i7XSfcZYtOE
CBrVb1av6/Og7Bn/VHILzdjBAry4TlrF1/5kpD6O5Wpv9PyU4SBD/F/ULJMKs5ptsUuQYnvnqBe6
M2iZFUBhTCma06Aky7VQcndGZfIcj5kPCFGJb8xihirIm58cJoFdkTKPENlgvKNevcE1F9gF9Zk1
jfjmw+pfbu+glAP1ReN+cEGDSXaEsqzCA+Pzl42sdOVFK/AGMabVhGomUaSJ87HL+1aJajvQLJsR
MGZninFYwOaCFyFsvJtJAGLGfg+LCsoGUsqgm5tZm8fPV/RAF/UA6vnYoXQ7EVXvfOE2gc5CgM/o
5g58K30fqcWxQkZrYT73zZ4sBRKoF8dtlnEF68oizRmc3jq+fhm7/Q7oR8TH6xRD58acalcGoYdZ
54Vz++T0g3lPbPqnQLJ/25Pd2VGKxhPvEzqGkU7kKJRWXgKN81d2HmLudqjt9k6q+7g1UsedLnC0
zM4ffpylJNBuSnweTJx2peBZGXD3Gz39tCCI88sLwkMzt+aHRs8TljXqvrl/D9zPIoyfVBH6Xs8H
GtdwnXwIAMLKuDKUP1oqleWCsroIlPiNvpFnTmeMjzy0KARVzw5+idblcteKnTBS4MeTl2LRcOar
THesQIBn+6AIw6kWz0P0ZOvkdBFKmj/pbWAuLTGZKACq4JNog7xX++S8eO360Qj0/hnlP/kNDg1E
C3RojaKEY8dS0og6uZR3Unh63QhDKRaYyFIZu8dcLlc6fya0ARjuQRoF4dnFb6c5YoM2kVihooZD
2yzNWwEXu2GBVOtuWkPGhR0/OvIIEXEljOuYwCKo8piNfIygmmqytTJa6bm1IE6A3bBLhCQUUtvA
QfyZAvNF2ZJ2wCEWbE4x8Y+6uCAocwwbZovN+v9HkKnIn19tZebM5JeB2Mo47uHHEX56ycdULrbu
+vwxsYDYQL/GkRbLHaz1cRaeXqDYsVFZz5AhKmpZUHPwRVoDgXNelaqkyyUD78pFAXUun7VxolDI
/ccDOgSOXTC8gEsT4e26zErJXPMaPSwH7EewygyVsTS2P51PSaSWqeI+/4zaK/szL2SUIdVQ9ztJ
NEl+hvA6GJrHndKxpaZ4SQgGUCVFFai8HmnDPpEZh9XQzKO1K0ZrI0ezDwCp/XQaTI7OW/zQKGYT
vejBpaTIpM5vILxQPxDHa2TBk0twlBClEO1LOXXaIGAFjiUSvRZllWkm2wPgyr2f3zkNv46nNuO8
wduvryKhTYQgw369AiULPjP/aKYNv3NLGEXIGKIBiE4BpJqF5/SSgQ5ZS6BCwDU2IGmqBaeBvk08
2JcQWc6lZfU0to/MlFeQ1ecPQt6ZNAiQxVI3aFw+9vVy7aAwQtlN62MjqyLesyb8Ku6VJgXZKl+7
NzUD+oU86xSB+TTZuiUwUoCxteZ7TsWluj4e3WHXPVCXdfi7QhQobTroWFA1b1V/Fd3229jSucnb
jEe87YjnKRmylPQ5MQvC6Q0qals6affZDewZZiRhwiSdJygQXVUejbKaOU0swPeGjLxyMJj8TFtI
fHt/TvKA3Wb1Axthec0UieweCLcw5QfmfkFY7QIwMSQ32+dYy7aU/L61PyvvkCSHU5tiY7Gq4X4P
CzIHra+MmpsJo2e60aNUmip4MgvamETGx7X/MpYavbPSVuRj6cOiEvYaVWTI47pAHidRPHey8VvD
y4TCAlYxKd1aRrbv1U8hORMRmMs12NM1GQdlIas/0tXC4wYSsBREuFbG8EMrYATYz6F/Xs+H9t1Q
1Uiyer3m1P+x2/JXGRBQw8KXnmgNlYiKb13+TiFKB85HdXj2E9+gdLy6EslK9BE/JNQ39TWLvuTd
b1l1DltfnGp5kVxOVcHF7Kmxre0zDz368EvHFf9bTuXCiQ0PeLgQOtnnjKBnKcfn2CEBYzZyPrei
+4beed8eOy9jtrDGniLVtsYhsoUP4xRo/dNQBv/McEEvC74aSwKAHUtclJ7fBuDDWwDAN8MpxXVL
cTUGXQmKmHv9UonepqNCz8ZZbxmE+/jX6o/efYl1e7vR52Zxd3Wje530DuindvkRENvIGMSa8Fhn
JgXWcyGxxI4X6KIPuGh8wq4TrPszrq0Awd6bKDfO4f+99wSgWBBBGOqGIsvJLqjQw+izObgcPsJm
n39JhdkX7yD0E8F3oyjEoCN4CozyFMRAXdjS5mWE0HZaxTTRL9QwHlASKG3jBwz0q5A8qEJdJ1yG
uiAMIukCp+l3j9OD+bvf7Cr8I0UAoydWu3gmi60EOhjD/ltU/yU0n2n46Xc+mt/lt/b/lg6d72gn
Nncxdr5WHZFUBudZRQuxiI2zSL0HDG19+8NMZ39oOxXExDXPh0pH1pg1sj5uYYylV+OuxYJM+h5V
7X8dRQtoNP50xO5dH/SEliz8l0LWpzOJSeUTYjodf6Lii2Wj7E1OM61ibwha5KlgiotXN3uOsF2t
iN801sqHRgf+qVxV1AgsXIQEEaRh23blXhkDE5Ny0AtZP68W4Su3klEA6RnBTHkpvP3Bh0y62WLS
wGZIKIMgxXvwtct2+IKf1yeuYyLqoNhU7HY+4CnuHhyM4pr+mua5QG2Z9Npc5DjDcDXtB6Z0Tjf9
ZIpOfSRsmYTjZN3UywrwOwxVVkdfPbAkziV0sGKwFPNIq6WemNT0NizjiuWxK1DPSfRrZGLPoLB9
x1el7s9tbDjNWMPurmQodNfu0fs+GYx3AMSI+rf1cuCtpLZ+xYDaKwv5YF/qjjT8Ac/5vqqpUQkn
G4foywkZM3YVZGmlgqQj+0qRTCstpcpbdcMUrBnK0lD9e949yIyclk4PH6OS/eHDnwo7+GZykPj4
szbWrz7I4PPl+yLXID19iYv6POy2zi4hSYYsQq2hGf+azX3epc/xq6B02yqY2m9dnA6vKmDqYpwp
oH7J3NRnD6XXyC/C7ZJuPrAwg+wUD09+QG4/zPzqQBh9Xzcvd8XX8QvKSBWviUuEV/cuV5y6MFdP
Lnl6kk1a7RBQF0cy065QHFd2yRhi5pNgUL4Ls3k1Mzf7W75SNQe39/IWigpAXMQ2gkKN9ZMt5Y9y
ZkvU29s78KZHyVeh4hIJxc3qSTlXDPAuuoRN9UMqN8MuSWs4XEBkDQ5XRTrFMWYKatw02YNhlK2s
1FEaGoaMCBZd1A1aAJZ4DwzBpzG5PEqppNx2q30Sqkc+brMFlkoxzDwqvG9+acD8iGQdjDfBCU+I
VoynewDzYZTmTFsY050+jtRhQVFcrTMLLYXm94Bh7+OldZXpbUz/rAd+Ntqj0Rx5wZRx4uZF20fn
5lhu2bJnTneOVDPZJO3CaMF4TrfcUi4d0sKrEkozOZ7O9lnURIyB5cqYUcbSt04PhL7smDotMkiI
7FBtBF/Gf9HJ5Crqm1R7P9a5w9t786qIqBIXRbcvRCJHqNGbdxCEd5ObmoGEYLKe8Li+WNWzvX2y
Y52HxkiGUquhDQkHCzNwsOJ54nrhIDm5U58YO9KXA2xAEuPAC6/mGckpN1sOj4Cniajn9WHJV0LD
xByl7WK9HnhLwK+llQrJIB60r6eRO6HrVoPRXvjR2SR3Sq1c5nV9Btj5Ofh/tHFBtgReyTSz6/Cn
eL5DeTzqDa0kbX+3xoWFm0CluVnEfh26rWQP9yGPvwVLkwPnQ3r/wNXuZo9/atCOywwAASxd7x2s
RcrDVh9HixyWUD4gJ7Vg3k288ixd1npWNcZUA1rpyIUeFGGRkFFNcCYLEZM8SE/4PPhmxE9+189w
/PyjJyqc1Rc6uXnw1xPkqQcnZugC4XN2wUGj3wnQwSgmWEpa+0Q0qk6Kp8/RVthtHPB3D2IQzAws
xEIU3mR+Ktt04A24wTihcHhnQhep451bgw5lXSJnllfbS4J5J8pXPtuI7MH4AZ5+n4i6XkyE/Y38
qJ4cwF13lYeO2ZcHpoBomOgRHTE8hxNxYS5ldKULMMH6zfCbd9rfrMTKeBFYp4OwZ9Ztx9yovSKM
dJVp+D8aV7tWsHm3XphN+DIqb0P7CC2nAvtVt0pHyy4Ix1T7ZSfOjxEtaswy0ceJG165GdTH+pD+
MyamdrBGEffqSGaoUWbCpDEWr6ZUO/muQYbG+fe8fZu5jxSAlOHppQxu3NaNruFhbbglr3Rvft1E
oYB6FCH7uUuqLeC50b0pSUDrjUKjfiz1j4zyITUxgpekGzJbNSW5RU0g22S+1StmRf6C6WjJ4iBD
YrJtGO7/4SXXGXqO6igUrmxh+LLB4veANYnmFMMmAW9WJEtN04s9MbcADjeJEn8xmTH511Gziw4d
c74vplPLKKLodLxn85/N1M7/fAO0ItySVb1dg3Z/iDtj7bTRDRVkLF67Xf33FMONoU2kfonk3WDw
6mTou2qa+LvdHJk5MvPZyDqRbASn0j1wzVliVfRgTp7UdVTedPO2UbAmF+FVNwPFrBdzUoTlVibD
1JxQYs7ybTUtakZ+XlP5cuREHBKsTJP+WE9p8kAo0xLoCQgHWnwwf2a44fms4PDfAFwth+Z4x+3d
grQnLX/0L6lpcyVTahv+VMipo8mdFJ93HYiUMejKIg9SvEu7luet39A69VVd/0PDytkZk82xzA8v
CRIO+WxyjvLhUE/LogGsvy98UbrSf5SIMBaUy8KJnZFRHXhYOO6kjuE++A7ZSsBhhYQU1WKGFs7I
/+GhKDKR5f0tldGncKO4VYq3eOk0Bm3b6Uv1Sbky6vxGz7wX2s6FaQ6O2OWAwPUgUj0sQ2HVQBF6
XaBruTiUOW3PFCFpbioiWDNze/+3oNdsyqoNh1iQHOBeLj9WvvchG5/jhnKThBlaGK6DY5XJN1hb
7ab6elCVktap1zxR1Ai8p92U6eY6nYpjX0mrQ5TvBwOWKJX5/1pKFKxuy80uHcIxDsKJHvc4ls7l
KsJTV3GgQKDvexkMYJhzDXp6rSFAvMursxRCEgPyqSfbMCx/oyqOonb+nH2nrtj4nxHItKnpIPrJ
Lore1f96LloTRIV7k+twHCbm38ba4WzmCI3JkeIP66ah+/gIu6yD3olHTSutmiX676qHuq5VxN8d
RfgCHa3fSjgyCbBm/7H9ebPoQqO/NkYlu4lEt+uR5dvYiAx9tYqCUb7PRqOlAuNDCRtqQ2EUs9pB
EKZ+406bv6Nu61kBhpKrsG/meuu7Bdai0oZVbv0tHo0xqw1R+jyilkoSCwJZxa4PELE4Q9Qcx4aR
wAx8/yFpsbWwFOK0Pg4gsf5dIYpi8ZR+ORNGZunjaJZJxCwlcc5nxfQWTDlks1VF8JEgzpDheKXT
AWSe2+TlkWWDPP516tFd3KEOT+nnTTQ5f71PjXDHax5voFS1v+tSLtkVJXNFcxdMxYRqaP9HhdKi
2Z7VVTGJHMNt/vJOWE2THO5+QMxbUFO4c2DHZKdoiZOgV3YD6VvI8YdhNyxl64nL6UmSicq+s3G6
ADZ/ED5W6eMoaX07+2NCrXVe0KgMTxLUPQ2FBQITqWVLkbR31dg4yeyhmTYlRXW74YOtxG3Ryofp
ea5CnyPyIoGOWV2ElE8hxCFBu3mQF/Ado8QAl3LxKrCpoClZMOFSI156TzYlP+dB3xqk/x12dlVs
fX91oGTQdkTruXPT8u/BQGzcPXWHwL8ZvqPUUx/Bln6BXg0D+knyospOLxf9I+aZfF5JNBV2TRhB
SWeF90bM4q4agykqBGiuk5768MEGFjZnMPuZRyqcXF1DwIP/FQyaaNPvDUDiILwJ0T+0csflP04Z
pJHodrnrCT0Ds0EOyuh/6YJGYqACuCveVkG+Cq5frsLrsK+BYy4kUCW/1+HE7KrYTE+ZW0ItA1LM
YI/VIfibO1G5xqsbe+qsvsd124F3WWqqC/Bi1jIhtLheL1XPnMS03DDo7ilyiY0gomva9U/xqpJX
lKK5NzwMMztbDFNTQW1+a4YIE3i2ifR9OUz0CA2jOI8a5+2Tz3D8/xr4xJeQWWwa5ud9N5Pp1zcR
osrdpnT6r/hgFXPIM/Ic7BKADVKCjuepxAZSW82pQYyBYBDA15QUcRXAztFbQcuwJHHLPBu/oJQp
r0NkZ0fMJDxpIado64M4/PBR4bGqf4x8IiF8mNz6o4P4wWDB/+CzieHwPX8KpwV9p9n14BhBd8mL
vSrxNPq32nDyZweuAzS4/QeKsuouXF5E1BZemNCAIg/5oLPSvMi7CIIdEFOFYydPfr/dnIN45WmI
1h9EEkjNhJs6HmyN5Cdtufh94i9QMVTuYD77C3j0Faz5We2/mDEm7CKrFHvWqGD7TqQcdDzSqaSF
0DuOsQkfz5OKln7Wqwp13Nls0HNjRQ2q5qxHrQfV59ZwRCrC+S86/7noFeuONESun8LkTK+LjPdh
xKfWT3uPLE9Vr05ju5so5krSNiQgOt7/VWD5TQlaH/YfMxgDwlf2nt4soSmn3zj8DklV3R72TQ5D
0sg2ScM3gpf6BuYwS0b6P5C8qfrLvO+lENQYb3EwpPvu7NWyvo4rTjIun3NS8xJMDMKJWm37Wnhv
EzNWTYwKcDCfTvUdLmZhWUQe5+DDhuFYcUcBsXUHwIn0zxkAZvqkNLXyW9VWFvTHNbCImJz0Th2t
rkxyj37rrKsATWBKTTa5VLo/uVXMGVLEonfzTvVOc9e0v55lEO8k9Vc33k5NBzda3R1HCbb97mCs
FCrCPBKWbpTaYWqy840PFZWx1jAcvZPjAhnXsbPopnZy8DHjnVrlEcewrLZEMVGImjVXle6EkWSU
JKVFkCR4a9/HC02SDTfRQCrl47MXfs8EEnAfOjfabiq+idbUCqogp9Rfrn5+yiWgmEKrHCDg6Sc2
OXXTgFiCqHIsfvmRpP4Dmz6A6EwrwwDW3EXy7BaqBXRV3YULH3GvQn/i/IqLEW2zUsBetAvUBF8E
gERSsJ+GmMU89rn0OT5atQrd810LLIviPUlKWWL9bp8GZDhqvxFsJmdWp12CD4OtT3/kfh/diOn8
NnrTzF9aBtGQMGMHloNSdaf6weCApBxvr49AsY6iqWeEdtZlVtqYqGAAv939DhuX/F8iD9LF2Gsk
2hugtVwwMq9X70Aij/bmu/AGK5TF3kwFtkntjI4n5511MmWt/8UJZaSUtx+3KTrXfeYKa1AmQejO
bchldoWSZ1NPeTGpEdiqOLq6pvt0yUz0f+coZcsZns7j7ynTY7BBLS3dl37/KANoHu6O2JZ0wMLN
fIHz+wYefqrOjiWtjM/NfiI0eUPt0EdASGFr8gEQHpKHjfqBP6SZiMkZRuoKvxDB4D9nFNq5lNCF
n32HIWKxkZKQm9E2qTCRvDFmTUTEO3QQk8Aa8kgDLhjeBrZwuVXo3cHRZYdWOQtHJnumatLf3HuA
c75+bbatQ8euGLo3ejTVJXV9oe1NMCiJR/Zg/KUmtRy3F+hud7jQa2re2ZqtXdpSXLC2/M7uGHcj
6o7KIowrHTgQBFd/KsDpZ8UpaRnKHvaoxqJSP95RSpXYBtBbprLFMp8Mn5bJgf9wbcLFZGOsemQS
ViqXWaI7VorAgyHN/laRxJKfUSEwiCW8+LA/V7yZLBb7vH/Tbr3zDWMKBAJ3CQuGVBvmMAYyvll2
PnUYzDQqcIBf2CYksy0NBo18EIbF801PaH2jIMdu2ssbSgYNp6ZxH7GBGL9o16e04zDiA5ztdBGz
orcuZuXiRMOoqLVW38QhQtSXjIubR9ycmrDdJ7bJ+Pd41UVPrO/qRoYu8bY50bGYPDEERxdFg/je
e9nxxYB7c21FPt9y9htid1RDxxvh/F3ikRDmnpZ2w2+Un2vVTYSmFbv5ceYe9qSmDktwiSvtphXf
YHwOp7hNLdPsedbMISV7RtGV1Hnc9294LBe9MNObU8l5JthiLvVMyFCexzwuq2gBzUAeOuLZ8bpZ
hkjE3TIDlpsy+jiLjPnslRzYxkPtsJhTRfCKkITmSACUImibBsIwXvnSkb7DeVmwBlKebfJfBf0d
+eN8gfqdQbAR+SY3BqKlyiCGfpQX40/EOhvxcB0efvKjnHjVCCkDtEDoEuiDNN1zNZjQzp0I04DL
bthFYjqv4cfw0n+C/OzR0NQC81BubyYr5S/H9w5AM38G3hcZSbh581ebV7Wtt9PHF07nXqb8ayNb
fjJpVlCl0X6G+Vqs4GMFKzD9j6D2TZNrkSWKZIZ6oBMCKnQz/axwDNtjzlqaVTNfKWY5pHa8l0Dy
sytw7SgJLIrzx+LZr+Sw5NyRNW6+suUbykdRfctpDa1CPplFpcQfqrGif5AA3+Lz1wVS/KUJlMsC
nziGntNZ+bFAXD+y7mAo1bD5xF+RFm9Ric/opQ75lZtORqs4kx4Reb6xzkym7pDa4jreuSbI2YTo
QGGsuyto/grMJ9E1ZH+qS/GIRqZKi2CA/C+oPJNLtge+4Ab+l+Fatf257K8lJvUCeaJBw+f6+mVx
tQZIsF1e7NLeFKzYVdTkvN0D56qh1rNuxL4/WZN5X8JUnCOnFTjsCnQ+iy5Xl6Ba3tiwtCF83Ywx
I4gtE10DoT+NQieNwBuK5KzEFBozZAKNATlYxwsszjjnu4InWei1L9S4LxLJh1iHTbFZlSnSibbR
2rOUX6EsOFdjFup6YCK3QadKBT4WKin2lGl4bLlR5LI6Auk9HWXNuhYOn5JwqZVUC4ve5L2k8Eqh
FPEmw3VNw77L/xrhJMV5m913VVZcn1+VExblycRgxhnGtY7Cy/vBoWF0sCrGe+h1cV6SsBfQX/9c
ULYxfTKpnMSoQlmpgX6s6F0HTjdUSaKn7DnGJMaE/Y3lfbMO1g6uC23Nj143evx4lt0N4Gw9Lxzt
1t4otYY8aUKnDVpZTrhIB30v6GlyzrM/CHCfDIcM749Twj+2SMo311gzG35E/GBpSLvn35aaZmdK
2vkDY+HUg+Nf3FMaYSJTgzmf0ZGtnHKr1CFG/H1WsJYLbsnS5TZaosa+Rt7yymztfZ6Oj/oKTiBy
bCE4im8P5FQUwyU0Cu96J+vKsPqI6eW/t3GL6CoIn4HgXTFrw6aZvRoFxwW+6f/uWc7IXzd0yN6v
wnXlLvEMYk77ETJeAgE5/ua6pe+aA3gpCF8e7cwzwDVgXlgDHd1/k8stoGfnwDqR//toRvA6zF81
lOryBsReuUDhAFuB/ErwYJY7DgjeDnR/Qm6jT9axniX/SPe6GEmhzWiDuDd8uKhqiZ0vj830wGj3
i3tCo8/6G45h56khx0zRK77D+kYzGpumdDWLEYTB9DEWUpAu57zNWFBU1Bjr+Oj22qBI7MYBRLZ6
xqbcanGv5X09fHrqmExHa9yCiOFo+KVjTscejRzYB40huGrjHHXF6Sv5HZWzdzlrfKrKuwxgwO/F
Dixa9QCLtG7cT88Cbdq9spUJcKLSqM/bbw3xZPwHU+ziV9ND/NwuFHn2arI1RtlWxzaiAcGDGKLu
z+fE6NM0yBP9KdzaIFN1LiuEkxDj+oOp3MwTCBh0e8HFaW/f5yw2kDJCkcDb43M38j3oKdAEGR6k
akU/dwS/4BoTkmqDD0EoYLvQAdEGs6GXBVbv+2FxaKqmwUNAKhDQ357WwuoRV3GNUwvGDZFCYKLM
/gG4VZ4S7biUUs1kPuYbnk2rGyWC2sajNMTtNs/SAb6hja2nM+kajSvE0EDfFyJRt20VPU0z2G7a
M8gQ+N2k4d4cuDsgiYUsJmfiEEFZRkGQXTc/UqP803mQq0d3KOfs6wbaZA/2tDl+ZYIcTjJfnKBj
O8UDgQWaLww2/NJ7XCLtYWdh+SDoRKFM3yEuePNUM+e66x2/Ri8DIG+GgYFCcoZNCYq0zkbLCsYk
d/kFrXUHZ0D/1VI5ICIv5L1+d/ellXsOwEMwSOf0IR0H073RU/5Xqze/FnV87SUYcFzvKjvFz2Dk
GJ80pzA3PDze4dmnOOY4KbRE+BNNwQ6CnRbJ4VBpxBAeA5Ycpi7fN2CoZUXoQsNsGOh1sY+3r+dZ
Nhb4skACSDGpuo4rMUIqkri7phDhbMGgDX8IflIfFp6ePazRtdffOVeARSaFoU4X1TjtLpCrpItD
xNNSMMnCwY5Zy7ldKYjt5RHqKxCsAn2Hp4xxbeVhoLgqcXRL8yLcArxI7W9fD2D1YpWv8BzAElt4
oWPPlLYIQR9fm/o+Ld/Amo2Q/97ojH2P+iyG/wX5G/ipDCcgmb4+g/L9tiiW4TYK+2QRXj3WEhZT
Wum5bI0aSFHceVxb5uOYJGpaLj/gYsgE/29WUQqe4/Pwcj6dM+nCgiunbmwQjFAkRQVIDIFxg5+V
Xnu8T99TRlKxQGWu6CfhNKwE7Sp/cpo+aIJCGvsO/9Y0s6bkPkAz6P7MdearvcEXOWfmyoKyxH5W
mv40vrgNn9Kx5ZCKYn9U+kyLA/z7rZ37Gp7lqOGaJ+6EHN5nZTCfT1ZbVqFoeFEqxjc+zDRq9EWV
EBcGyDncg/hhyayuFAifnLKAf//Z9gu4SFzHYZntP5xjiW3jWiwLlm6Jf7ZAlPWsPMrbQldglOWV
nTr/jQBpA3F4CXcn6gWPxiPNcKWV+V4GFljzhF242hQmFhKj0seSvZ/WRo/GTU4G0PW+jcxOcxoZ
0MCaBYupTopeK49V7+LgZvIn1OXLA4kMg2/OIeOQVGhxbmvJgANOE8QC/Vu+TZ6K9zMKfphNovfU
tpSNBed/SZMhrVEpgh49UfYLjlR/CjQBlmdqeQjJlsldQaJZkDXDy7EVHoxp/ItjeG2OiB/BWemf
nOhMTwi/b82qzIzeTku4kGtsvqbHf9H4wktzPCRbLipoNnYxVj+QK2Mc9HUQq2xJmzF4gwazQLUH
lCI40suVVm3M+gJSUVIcPEaWqeju9Nw6udgFsEwp2bb6oP+DUPXtXP3rfftqzaIftiD16eOEPRiS
GbOLb/hr2m/2hmhThPT612LZj9AH7bicwfRjFf+j6ZxIQXizQNxsbdVYy52vHTPGUv8XQhCbtfK3
tHTD+ExArO3u3Vjj5pu29AzCNtaWG9zCAVvnCuzoBMgH8X3bgI9rbaz6gSEVDnHWDE+PY/Ks2TJp
OEWrLmqJ+BNxpdvE9iZaaREnKS2JZnBYfSqDjk2jafhDQjnwl55QXsCjRBYL9ZpuQNbPx+6XWff2
lVlE3UA2RT5mlUL3520/po4DBtVA6OZey9KKlNPf4/5kThiI3Y8J1wAZnBj3QaytdCxKjmrjfr95
VemcCSBAhzBg8RZyz7ZxOabIKKg3te2u7YyCrUSBERtHMkZNUtLTpmJYwg/Nc4GX95fFGR+mp51p
4jYzDL8N55BUMyr4LZug6uQcm0di5t9CRlFPbmjx2l5LeVR3IWlmDmXo+oUPerX4/L0UMdpZH+x9
M4UPXDsMIymWJvfsz3U7suEOOnSvjAU3gYH+wIff3Je/m/fT01iN9hU0lwce3WkIb7nCJsJI/6lY
geV6fUhiLIYlX0MQ/CXxey75DuCNegbuBqIWWvVbOl9YhxJnu7z+16y8Ul2ensl6zqp0O0FeiA8g
cMm7su0m92hBCH/N6cAejsZsqDxUbcenyoH8eBUcqIWhty170OjULF62sN+rHmSpZB3uTwMOqCgH
g/f0s2+2MucTb6oTWLP0nj/CEG6sgVj1ThEsf0zEffe7Ss/k4wOf/ZsC/Yko/dCuCJwyKGBBx7H8
tEO04ZWBQCuS3iXruYSykcDXHFQPjkKGd/K3y6+J2BdXkxL+tx6uYVr8NdxGDN4Vt6wRee+hQIB3
xwSvAWjvDfGpyBNewl8mZNKZIhQGu3vLFjxLdLIQtCqbmeh5PViiy0DenfKGEq3trkMzwRMVHp9p
1pv9OkXpA/FqzHsQPmjdK8SDtQHarShdPKTJ1cTMnIMadAugRkNQRrjsr/+WJ0nBCsgvMJJ0r8sX
4qkUYgrxHcMxMj3c0sIzzO2PCL96YPJIAKqcc2ZPeeulcgLsWJsnhnC5V2PHLwhghDBIw9xcUBHV
8KNApEkggYc7KBsUZ9bjyF//bbRZLTTQk5R2MpLcVImQ8YlGBhvQ4B/7C4UW9kgyu+4L2Da9Dg/c
I5gsFJ4+VFudeofZw7YSOWqG2xzAsC/GWtMmYKWCpoVJRIwq4tkUE/rXtQ9qwm7y7Y7SdX+M0aPj
RghhCx4lmY8EssA5NlaE5UbThzc2o0StkIahPgvMqDUdWlhQ3wZmLdQR6A0Aq3lPHj/EFJ9OdWLQ
YjLsQJGhSPsfREXtW3IWd+tllV5f508i4OcLzCOcJjzvG2ikAacM4Y/Nk+ftyHG3kbfSaJp65Rwe
aB/AncbZUuYJwWM5+JyvS9tu1p+u/Q1vdxCT39TcX3erk/QNmLY07wQkMzptjfHinwk5uk9UAnYh
syq/fx3zlM9FFF172BitAjItDNBJwh50p/yWadR5g+SwZbHspj41hMekOH2mFh71QXWJd6TEMD3a
Rcz7xhwvw6GOJyVrMIVo3gCrfJDFz2TfsZZCYDsy2l1eHAwYFws8wV+cZlqcbouixM1tD98g16lO
p1Z0JfSB0lr0z4CDSihd8CrZriD7RGWt55EGiiRsx+X/O9GhOPnmJmNrmBUtreEj3hAUZVrazn0L
cQLhLHWFennjI7qpk6DXaMdqsV0eTHz6JHA8sC+hZr4ISgR7iK4WKGY2I5Ifki/eBqa6WYEnjFD1
l49Bkr3IByeVtHloVBBqxrNtQ+RRM7oeuC4v7s4BwWL4BW1jCMcnkLW++uxZVFKstcD1Eu/L6A6b
UFTHB/wvuZlz6XYrmSdDXjNtOo4viq98NeRe0QDEtO1IwymMEOI15SolOX8Bg0/+Zcl87Sir62N6
t+d7AOsv1ZhF477oY7or/pM8Uu1k3H9ZOvXClOHNOi0rwnz0WOILOwnP+rsJuuOt5K0OuhUG2FAG
LiyRI2fatCICuVS9sRlfn6+pdv393/liodPUNeL8ulcIIJbP/YBQd9dh2ZldhtuYAyHuPH204QEc
sQS7oRtoUS0cJWx1ZwD5MPNrSl3f3oO34J6fad5bU30dlr3CK5+gX1sHAq+wna2VDa75oRk+0bCL
IpsSUDZ0wWxrFHQThzZHBhgR3nV7JIhI5Ulk0LrnvxkHCUlTRvedqtbcs0FUaVMpvXioxXZYJe7O
ZKRSQcqFJREKkFQT5Qo1mg5cOuOsXdah6uXoUzGqlOoAFk/zOfM/r6b4gRtFgI7tb5RVhffCQ5O3
whkhFaEwqQleAcHIbjdL1GnOMqXB9Eb8tvpefzmiXoJ147/r3co4jmzvwKvU7mAy/9s+/19gsRSu
eIYFLOoxzzMN5jobnCBKCzwa20SYFSNzuAjzHEVFDQmfOloJJLZbvuHpbqCg6OZeJxclf0o0K7AR
vwNydLEF9FaW2U82cB4RFGWPaKSiQ56QqRmLbzVC1bqJNV8Oqmhux2510GX1D6HzPJ9F6w+lolWB
aQlKrF4X8MZcyG25qF5tCh4Gf2FS6BEax8QLWTihGoGkE4FKGFFhZ0EFDOHakErCaUJpFCl8jrK3
lhWvFPIkc+AJ7UMptmnGQd9mIYavPZML99uqkCEHmfHTJ4aJl87J3QnQ8pqMfCT8+3LhcKmRmqjz
sSjoRk4/BKd85jcQEM2LCmHStbdNGdYFY03K6ZjmvvEaVusylN9XLkTc/LIqtd/sd150eQOOLSQK
i9ji5rWl58IPKp2xxbASa7Xh0Eh7MdHGO3oRhsoqPVa8g35GmqbCaa3y1GnJXDbwFUf/u45L6bKD
+jhj74zB+RDXuNSIW+Z/gY3+Ww/hWexQtxRCwLhmBGctUgIlWa+k6rq12HuauJKrcro5FdnJdi5u
+mKEK5yQ2jCjtQFrm3nthQu6aw2QlT63V4duArn3p2tggv56IaVRE5h+ERHaoLtjBeN8vxMCp/d6
IPChwzVbAALwb6CmpKPnCLLVc2y4tQIj3PrmvW1MpbeiLVMgahkJZ6yo/dJOnWVcrYhFcrOlgYT7
/4oesdOjBg/MjycAc3/GTN5uSeYb75WuGuM483wnqOECIf2mRxF7qYvGakzbsLHrnkWGLZcsa83n
NwgG/Cow51YTjwkxlfOwtZIb3yOnV0/FVLnVtAdrFBM77sNhlvMjbW1akfckEQjinDXkZq/B9TtU
MV/j5NpBOTh5wRmEQ+TjnNz2wqmjNfbURnWCNTvM4UjBLRVyvLZ0COLsnSN6JK0Mw+O8iMtne/ga
vA7bk5EeNfdbsLnedScuBPGCfLwPKF6WP7Q/Uu3hIO+xTspVF0sYtxMOIoSjFIqtcJ0gbyDf80wG
J7AuBL2gK7eEzoadQI+iPMluTSRjb8+CSOCn1fdH3LrXAtwS2iAbDXadgXWvp5fUPMdl69huKaBz
tFRbD4S91SH/tCRz+B8TzN6SpJYY7ris+I+P6gSxB3GsN8Fcn0q9CfycEi1ujepUWi/Q5Ltk8sje
WBgJuuSHuR7cJtTBv05jXeHaxqc7mFQYZCUoVu1jCsi7itPy++NTknrG/q9o90DFq8dCfIbJtJVZ
oej9ZOn+2jUv2MehToXCLr/C5hUvOe/ariJKbSL3BhRMsFpmaXH5vxUUx8pXiSaekl8W/kVXlDmn
HegnwA+T9gApyO6F3zQJx5+0MOqu8gLTtaKafra5phU5U/3ciuCJ+fefEL9k0ICqbR5hhZm/axUb
dlLT0yEKphiApCKcS7G+vCDGMaPKn1Wr2B8OSHwazdX6uewE114zdvPf6Dx+6ghtNYkmbK2y/4kL
YRxcWpTQC0H2rkllRhH/d1RyvE3ilA+33WI0cYbkvKsDcPNapOFthExPaYHx/mhzNXyWftVSCTvc
Av7GjdTD4jozK2F5qwSRb8T04bMU3PkquC8odSnOaDGJZ5h6SsmPp4x3+yEjdo+EI6t+SebonW+X
h4Q1MrivVtMLOiTm98mkUtIwm88HlE9tAEy7v1RIRoBT+ZZu4P3oZaguKVPUUg7uXzSatfvw5X72
zJ8KtHLi3Bmv8cCyiTIV9Eg1KicKFZHoeyPJbaEGh+BiJO2iez8N9zwvVmjKB/+ZQR5hc1SoS7DI
TpyfCeD4IjzJTJY3N2vjJrpVUF0fE7pv25ykyh/vcNPPg4RW4knUoDSQaftGu4cFH3jiczHUML+0
COmOMbRkeVgBUBFnw9/KRFMy06bAc7FINoSAfGF9IyL7ARZO5uDz/pIY4OtaqEuXDvgO4DvNJfIU
oQnf7iEJifRklzG8D8VIFSLuarp2vFeeS0IEZiF+IL4cZrJwvTYzUHieuqCiCH381AwhnBsWhBQR
4ADNs8v5fEBgTKLgKU49umWywJzSROoSi+BD2q+SdvFEuCchr2RbIbYjjeBUAvBuc6BRIQtuFoDq
HvjKCX4fKos27F+W/cxzNfC1T5GA/2J0cq6LEODslDGwUR7fovnXhh6bzRPteK5Lz5jhoMF0i8bq
a7ZfmcrEk9tbw3uy4cKfjDGwTykU6egfibN/Q0PQ7GbCf/49/WbOAhN7qepQx6xMOnD+4pGOaq6J
UOrMVTsuYFBf1aC+DLd9nPMXpi6Clu8MA4Y2n7wctr6CzX3sVIEDaxIc0wypqa3bE70Q5kcQHS+9
RalEgH3qn4b7Ifap/TupUJ+HJsl7SwUisdjKQhTjlNT321I6x3sAstEJeBJH2Vu3q/BexfRN9w7x
M0Lu5PrMqYkju8b+wY4b/wpFgWtBUC6j/+XBWakOREpeCokyfT9aFmOUY2Y2pSmXxuz8+FhI+SmJ
pz4UspWmFEp0zpGS6Y4HBFTUM7PTNDxkdXfh1mPBDRP39iiwFmi0oFIRDG6Zt5GURE7Tyt3rp8yg
ry673tv1eHdSwAfWHQi/nMb2RwvjcTrgXDgavZokGDqLcGe31jfR6QNbwZzN1WacetRBTfJQ8AJ8
3Nnf1BmdroZuS3Qq7PYQhzppDDCxelb8qInXS/tfhd1mpelGleM/UOz0UCoe6xMBoZciqcPfDJyF
eVmBBf/QYnBMe3qOJ/PAT+222MJehu6K0qD5JMfCJWWrXv2Zjrcvx5ZoYG8cOgR2aRpgJjGzAJ+B
5hSlJmE6nqoP7pTZ7uD6C9eQvsa37nA5eZgiqztgbNjAJ109KyIbTlXZKuyoTcm3s1IIx9N3o1/K
oobVQccmCQKyEQszuSQ6bRTdtldezHF3HLentAh6EKtRrqMlbiPWXL1dp2x8xSUryP03C/3eTAjg
jyNDhq3CzF9L4AY3AN2R9EET2H8wi+p5JefZcagoDiKRg5/w5AuKqeoXIMeQla1dgcKNPiDXxhPm
CVU2xyhDb/GzwKVo3q0wlxd49YJwfja/c4rbDm/uDLNY0vM/N2ah8NMgLn61y5XkHFPJbGlpp712
fajWuD7xLEp5uk7hxgdGlcmv1FM3oTLSda88G18bQiqTvL7ZXTlIGkUbztmH+DWqhBx7kwZ1iRZc
VF7MDYWi9O5sPeN8vw7m0Eb9xalMHoLYVtY2ECG7DZilF7rGRb7wKBpwXjJE7xAJdCUjH5YYgZ1h
wCrfYngcoqLoTeLYVaISq64mdv38RdNtqKc5aOW3szUHDV+UQJeCGmp0i8mCbG0qIrrj/mDlyFAD
QAnpE3GeoS7TUnI2MnfWtkrm7zXMzQvY4qKvEPrVkcx1ryu665oaXNQURw7arV7uGO+FB/MZRL2N
GSLPi46CSsQur2q5hPQrlYsibbLZOpd79KXjZVfCf6NOKht9VDSrt1S43ch9492Lk7nS/bqZdD3i
z2R7yuH5zd1blmI/NtVU+cYvoZTLhWhlA69h1RlyrJUcMZwWxBhu/UCluGoq7e2o25JwmFebRGI8
09+NHne0b2MktVErdkf6i+A3dRgJJiYADyqSDgTAECPCXcisasl3GAYRpT5QmSe6zgCbMPmGwms+
aGaGAkPgV2Vo2DBw1LpeItE4GIrKNRK59Nx4n7J8VdSEy4cVmoZrg01iDA4keVdG70IpGi0kveK9
Jf33r48tz8nzuMrBzbycydtflnA3Wmyk36apssYdhStl3B/u2giWepEpen+xC5hOfjIrdXLvdtPR
wuuE/oQM3t3GjSB1+yDAm92mpuCiDlnLGDQ+NCeDfoigjKgiGjlCeVuoil6z5cJU2nRNenEThZCZ
/FH0ts1SvGuYRpT8K6ikvktHAAdSmrEYR5FfM+uirDkooXfr77dmhb3f3ttbV/L7oeovGIdQn9JK
DvE7n6A1qF5GYtgIATRfbqbYCJtM8DYYXy2pyQoqvt0vPe7lZ9WfGCOn1SJubIhZxhbowltNI5GC
YrGBecEgZLaB+trlPzh0HbpthZWRL402c5ayJRYXdNJ99av7X2aKnqU2qWag8SwrqlM6tiPfuuCA
Tzt2PGBswzM4ZzLrSwrq7IZ/OGB6nc+SFZ3W5u0DTEiZY31q9BiCGHtZze7GytWxQ1QMo2r3fdKT
TNLSvd7g0x/BNMNGeasOBK0ffX2vDccdVLsIMOOat8gSGOIWVIYiOsGfHXrUw1c4X6qtpND6MHPb
dIr/tWJ7Ewgc0Uk+xutz0GL36GqlfCtBXfEGRmorXGdQ6VhdT2CKV4Jd+CQBlYZEal6eaAVLV/lW
Mub3oFiHz9c1iLhPNqSyvLD7tOXFduEetFFOWaP4E7YVm9aSPdS/pFzXvzy/MA/O8wJVCqosYRrI
gvDZhme47FvoTVAdBRxqOoAF3gUX3mKXxjCJnfUarUOun4uRkOXl8uoT/Pd9A7aA/fZ9/v/sIQYN
mHDEgMU4zV/6AABh9W8IGm+rXahE2F9k6uMOLMwKmK38zw7j6waKIi5EmUDspmYQJzKWpKJ/yLE3
Q+KtihqF2lAhYnXyBaYWXGkXN/kQ1TSwIjpkKhZpu8+J+A1i0vCzzFFt2U+e0uvybYwv9xehGnIr
Q3uv1gbahbXk265LWO0TJS+Hu4Uknm2ga+H1YnBPemaw3w6Vv1KH3EbFj3NqFoRRao1wHTKgPY7/
YSW/JFLuOUlNi/6/3kAKrP5pd88ixzIq8ICw3uNR4I7uMQVEhoJkf9gFc5uwu0iicZ24Srd7Kyho
A1yoabTJ8cSuZet6TfqzQl1qw/dE4+h3gN3HBT0cWOmPsqgmEUP8kH8sxmGI/r6mX9swsJdno8pf
euPDcaEZU0/zKG1toDiDaoMWLCD1EiBzBwa9PAjSju/KlfZlk9vFX5XV17ln0IMW4GGCGpRIGp6O
iE9AouGjjB1nxMJzmr+TPM5Y8CTBWrcOdEh6ZYUim8ZeRBDk5KZLVK/ZlXwyJdb5BvisAZQj2PV0
7wN5oX0FJgYuAWEcaSNx2wc3EZ1oSQTm1bqTV2e+ZS6ikh2PUCLtpaPkU84S88TXO7pZQL03E0YI
UDIoi3cizhIvrqyCXO3mId8GVnx+mzvRkB9IfNuAZnMny8oT8IHD8q5WSvpM8c+nUIH8oAot7gJK
JJ+Jn7s1saB85vBUsA5aQJJLbpLOWuItWXMVXXYWPTy2ee7BWL7RpGimX76XoHAaTCz0joSYpmZb
VR/61Qi/UHQNhZqChPfaSX4adaQL11GFNK+yLBHZF5ujluCaIlwRyXEyBjgaYYivqM5YGWVh3l7K
9wk9Lds65Z94/IuQLczgUVHee1ju0/LMPQy1yj0eGsp+4C8l4YyHIOxSd0IhNt1xwEQ/t0m/w4mF
d75D6fJ4dwyL/k1BXEJzA6Z0qP/1C+om8I4JJvNN4gbdhetKy0nfNgqyKMPl0L0eZtmtaXpKcLQj
OOwhquIPpIhmcd8YSODllQ2WeI9SBQKx97H6b11h9LvufuEsvLNmE4W+XEi6sqZYB2zsXk6SaNK+
4CFJ98/vV9VgeQMOxQTNVxO7GVi7CwpCgvmf+sQh8Hp9Xq1IG3SBJU380xo+8jDUBwl5kBjKweiI
/MD8ocJSmADGJfKGzAEnrU11MzP2kgjjwDYCX7LCZhDQ5wDbYy+uAdfcHKMBpVqEm4CJwvnNrWj8
oaL6ZZRAxsYVc3OY30pymQLUlvJi8uN/fm/DHWVryiUrgEEuf9bRGD14yv0Dz6KGB4xyPhrUigkZ
7BT1+3oC9z+DEGaed8Ih40VZwqYNj8Ai8H/Nk5aZ0UIO2zcMgcprlSbIUhdeT8qAhiILQEMV3STs
GSOSU+Oonm19xYjX4w6qvB4mJnPMCEgyvbH+wuNbL0Bgnp82BiTGVH7WFiJvIj9Ct3qh2R9pb/7l
eppvkIeUsVBwDRzsGtB32U2UaOId+z2PLbfuKgH6vwZANcF/sqmPkFWLdSvM/l9VTqhIpkygr784
aP6ZmUp8xptirPeObnu7QykhtG2iUiP0aDtysToh4CFtTrkjewqkpqDQLYgXhMe20IsFqvybJGQC
sSbIz34gr+8W6D+S5s/8vKn+QpsZVTqmcCQuI9pvw8TEdK+LC1SzMQQYo4CAyV6YumHZwmTsi6cJ
keJqU2QfUkMFCFsQd0PO8DSQRazjfBzcxfpcvSFxCjdfxGYMWymdCBNeL408H9b+mef8yS6Oagnd
+y9o+WWhkGkA8mz9J7GJMV27qhvCre2GLRDhVlCyxJTieyKyG4AAOC7TmzwY6dpiSlRnCcXjX+VL
MTN9L6ZW+U/HCouKxulxAxSHe9xquUKpaV+XiT672hOadtN2oPs9kSRMtiS/gV2Sza6I+sQ4xumx
m5qKM9ZlPgDZb035hKome9G3U/97HhISFrYFgJwFP+URLmMSmMTiVzCUMKGC10mA36cS7qJKgE9Y
ooKH3Nc60e1MzR2t3gN3Kt1IKM/1btZJLjfa9K96x0Vty9TOake6Q8VJA86gXqiJHVqHohDmg6UJ
AaiqmRx6ZFXOKmTsSNVL/xMvmEI7uJcpFLbFQEFgQVRSQUYoIWY14oSh5GLU6cOF/H1SOywDBf7z
geBKqoUGebPmUlxKVoWypB7ibEFFa0Oj4yB7TPpF39zCTEQEPWdPOe1ewUhXDV3HxjEQdVZdesYh
h4nGIINwXWDrku7sVdeeT2XuWzMtZIChEFfVmFp+ZhDi6QNTtJohV+KCrFwdF2NigiUjouIdMR3l
FgwUEt7VXrzTQSHv1e7HnmFsiARKhuGhh2zcZmvgi+FaVdrvSf14qGtPT8206J/xlA12I3FV7/QW
UI3VUtG0D70KqspLKlxANylCPoHFYdokignGHM3xDYSaL79whBJv+9AvuVtzR1pZRUHqScf6187j
6UbeQ3XhIeBp29Yv3mq54osolBy8xSzX3HT6j4I1bL6icd5FHSZ4oUdw3bUKTjmc4blMZd2/b8uY
SztoJdmRASN4/Vd8uoHdbEQgZS5FF9KLseJ7fA3ThTNwUnk9b2xgK3vRq7oWNhxFLKcUpDijHEQp
BE72jBvIGNaqpyl2rpmtc13Pi0l2RZy/FgnEuuOeQq+T7cc6t4IPMT38nrd6LNhpi06RowU1HjvY
5UCzmqglFhZqmGATdBoE4JH18TDmZfId96nXS9JoITecsrA+35V5G8zfx83nWlbJ0idaMfBx4ecZ
nkwaKoirPPLaQhmucrkKQgQV+7HBrrXpx84cSpl6llswbCNuZeqyu2wxoZqY8GL6L3MVGdPvu09J
Kqo1GfeU/9KLRThnILpSMo5osE5wWl90sd6fzwPIRb2T7p8i2Gq26O4xtErV0tipvVl/ZueB/R43
AY1x7FNyZu6oWYiUAW2INKCC0qFYYym6UWwChERZBDYvINy/DhJ5UXK79zkzMI0oWqwtCZ9aXs2l
01pp9luk1idnvVv1I+SyDaH9lG3RerIL023m4mK//Jbhzbiug9MpkO6JXcQDDTQra4qFOXF86Eel
BBFPnYY9y5rnJwME485c0rKOkRfhpv1ulmeAQUyYt4I40WZk42ATmiSDdtOwu9E6QicFgdFCHxnr
mJa/C+ewgdUWO5S7hCbeTysLMmqlXZlth6IqEyQ2sPZqKT7y4eAMwWYrZiri0C2a4CkgHOO9jAI/
ZdFjNYn2+EymaMyLfess4Nj1zRo5G0U4nKDcjOrwFtxIjgKbkWZphz/ncc125AzCt1pZpBarLtnJ
w/41/1UVYI1PI4C2j1RdkxUREFT1ZhQff5yAO0AQcb9/cPym/1sCagboE4g2IvnNHm755hGWWNxI
R2Z8fA1re+plilFHZcDLYnWsyafe8lwLZJigclrj0QhzImeUA9ydg6FK0qM2j51mqFqPVt/WfL3s
Ag9F6Mvq5X9kfKoi8fIRoeHsCLGlKzkTHiygecc2QQlPMJuzTP14F6cF7LltMD6pG/fSIpVbd/i7
MHRYRTHqcTTlwc5AUplgYdGoh/iKUOAllJKPVnSyR3rPCgOSWIWHMNhv7xtK1vNO3BAO3aog/DY3
MT3p+QnfmW6Wd2M6EhqcWu3D8E4qHKzB3sdh8DlvraqBxAOYkfwIT6ntCi1fqkOYZeb50Zwu2nZn
ctbW0pfuNd29ZTKy57ZxHT9BDmAUm8wtCWVyCjNihUekHtDNnRddeCesCnrdHFO7YT/3C7C6rOwe
nn6jAwiWy7KEFP23bIMaBH4/muQb2YxkiGjapGN+bmtkcedkbWIWRYipj8h33GbaGTvnXtfExdUo
ZeV/O1qWNPUxoq0gzAOwmiLWLdMqDeArqOTzutANIHGHTMSNGlJd8CPkPWlNsb2frJbSJBJUXQ0C
+SKUnzaWOp3i7ZLU7XaN0yE44uEtLIBGBPo9ZRCn+J/Btxi7wQ7V9kY1CI20wojAIm34GBKVS/Or
kuS+aq0m0/21kOhuEn/9k8NYO2ULnjWA6aNVFP5Ruo9Kg7LTDPKBwa312CjRay0VOAvmzp8MtECt
Xc5UaXeWar6npYqJmJAR2uOBZ0VaqfxXTiHwToCIi0YxFXQGWG+bNIr9/xJV2e7XB3akAvDfbA4V
L5vHf2mTsxMKQi/NuRojmf5P3eYsjOpcSnHaNDWAYXVl5hpgyf2f17ct86vKFyrJglwcAxOhRyNG
/A5ilHZdzGvbJPJf7EUUuqLovQ0uLmzMOLGiL9T6zFmmZjAMa9nFLYa71zCuIi5EJ67B9SsdNIZQ
qC//Ng+LLsHBR/bZKSOL27O3hOn/h62wHXHBjfpG+nJ0mKEoe3KzAEKY+AW3qsATfScFmfrbS1H9
DPbLWXi0zg7on4t/NgNjVanZmzo1LXdJQERQdYVH4XvlRr81ftiVzutLaLFD2037VPuFMLLrTC8J
pPcqVNJK2QNFwZNqgqGO3i7N/52zlNy2W6CfGzi/2AC+egu5H6DLMIw8gm1Kjt7s7kSwZAlhVMbz
YkMgvCBT2lwvBy1EgR18qlQlacVpZf6aoLq+IlX8gPZyAh8kjv44FI+mcWMjyzJgj64yLV7yAXE6
ni3UIK8YYyWi3gjEROH8sNwxXSZcTXEui4mOlTQDnEG96WoBf+4GzYoiElawhJitUuHraDyXhLqF
o7iaB5jgqWtE8NL3LtjLAEdbR5WGDSPWF0S5jNYDJA5cK8C5jb5gYOJgZZAWvW7JI/YsNAx51XcV
72RII5L0XT18LVGaf6Icb4TanQkGGVNZSLk3jEOMpJlRXgVOnzzzC4ScqS4sX0eKAz3PPRtENs7g
4N0TwwOpOT3FJDnsyJ9N57JwDSSVLj1/7veEPR1KmgRBGIvJp947nv4xyYTMPGe12DYpMBSblsC2
7bDuW/UclPq4cZFh/4Rxnm+1QG6utFqxis26YX9MRmeQskkU11Yz1BPPz9XF7qw9DKFHMEu8KOeP
3Hz2Y9/Vs5RWtC686TRjrM6OZuq7YnOHU+Dm6qF/itcrYFrUeouoZ5y0iNBhrtFcd+B2OlzG+oke
0zFnXy3laWUq3N6OAfwxXQVeYKuzNCXTxbLEGUWf0AKDA+efoo/UZWOF9Cb13tdlaxnQ0xArTRwj
K+PFLsiF7KU19QnFs3QV9pJRMwZB9z64Llu3yAZGnnqXtWZSflkH4RV+V0iHt9/kkd82oxp64kvv
HaO1LgUkXAWaKp8aIVEAnc2I6h0d/ghvRxam5I/sgBI09mTveKKj9Yl8j+BENCqnUZrs4ZTTcj+U
AqpZlKxJWox3vYCCtyIE/CF2uqV9yEiCrQZZSsmUib11QgT7KXRSRrWbZnN3h56hJD7oDBXNTEI8
h30GotTMRk0f0CRrFl2cBpFDa5co1V+rOw7VKlIz4N2lSN8BAedOGf903bjYZngtdBNsIiAI32Ej
qV+GJHAtlUiW9Gj+dMTAGEM1hzV4ADleAuwGeUp9MYvQzGd42dx/EcXz9TohQUaIvowMKGK+SlVm
jDKRvONa/6FX/fnG7NFFvGJLiSBBcroDo+y35qpIq7LL8EN5f6PwmNNFSLw4Xiiqi1Lvs/O6BIrw
QwNQHWxEmZXWN0O1w4nK0H7982wPGX+xFBZJxL50zp6jlP/vnQ/MDn0nq2Vh/IAUNAu9KEFezbAc
Mq04R4weFk+k4gl9MxX3K5j88HfZgG10pGcxiPcslvtpTLL5zz38pwzimuUuGz6QBmJSbXDNXPg7
1AiBWnJAAlaZ1o50OgLukVHxG2HwP0tfUQyJJaonyQlB/DVypfjKDmBpPtRRFC/DAfTCufL6hQ55
EhEZftPUsR8vCdki8vmnBql/brdndxqqZVjY1G+lppl5PYnJFsoHqNhwLPyV3NnrVLJXBZUmCvIO
xH51tyYT8pPN1r0wTCzkfcsbimsdLHPcXvV6x44esiqLwp6FbLFPmfMXL3W24jubUlqChB0NCWLJ
EJzCOWto0pD/iaG9AgpT2pQrbDf9WfoCVRNLXvIlNvE5plNv/Po44UDNQRn/tbH9S9xN7YNlqN2S
+KXrlXVBRVL8dyuI2B+Ze8VlNb7c8M0a7hRrZU2G87LATe3nFm6O41SycsU/hfLq0Ufz530WF3tw
Jg4bQ8TaWmak4SY/VZafalGM0GxuJxrnBuo3nXOgP3ktfKRlLrJWPxpqu8L+/vI2DzvTSqS+8sKF
ilHUenX50ehHEMPR5fhrxE0Wbcsxb1um4+UYvuAFBZGHNbClxmVICqOSMqo5C3K8jdDSDhCBqmlz
MsqTdXU1q96i91RScXiaWP3525zdyvUCj+eV/eQT4WCvtj0Mpgi+x1+x7dUUjD1D6vI6+elEpxoR
DTRaheSgW06CAPfRi1ZUn6Gv8y7BS01tnCy9xn1WR6P6LhceZdYoqFakwBzMCnj1AkwBcDlF72Ej
ckaxvHPHkJfnM/oK84ndKDxqVGjVEiUgXAubsyI+xUOJLxvOtfmZKbnXgfphpgv634maMr1B3SlK
6dSWGuWAJJBR7RqbvxUaexyb01eKvC4zmbG5wwypAnNEuaxeamWCx60w8ETyjjZ8hzHeKz1ALx/1
c0SCfy2YjmyPP6nQcT9Ns3jMHL3Th+f3fYdFzVA3Q5ncHOcArMlm/wBX6e8v6OIqIhUbnx/Nhut6
DOJnqmNpaDg+mSEKDwQingz5KLQMjJMWrtjVXczZrOtXIR20V+/w4KndmADvTqcTfBk4AbpfInYW
nw5qsJHoveXvuxjtEu2KupLn4p4LPwFmVjTD/gyIPwvlsHE+6igTEbo/rwFMzqkLnvVdhVIFknhB
ie12LclPmwu7Dto7cVuTl3WXpe/XIJ8AOZpa0LV5aTtk9elUQgjyiaIsc2BSj1Z0Zrfmrw/z9FGT
U8T3Jl4BhNT/C91rUp2sicfdzbPyYrFu6BqLrY+v34ma0n6O3wJDjqcIS8TIS56qFUSaZHDq43CW
upHshOX6YI5Mdm8VU65orAVnphVEj9nk8sAngH5lfM/M18t7wzDEaGim03isdE+xUVS2T5q2nTCl
8+rL8Ir2FNGpOP8D9ZpBpr1m8I5nIiq2r4m8KCpG5ebh5eXKQBS6yONDE094eYBOdpMV8lGf/nC7
tv/pK1Awyf0XApK7n5/Wl/PmKnvNRn7kG+bjkus/OE3OjLlBn/kCHMLUqlHOrnS9h9W0LRDRM1S4
2ClplGUlmmo6D0dCOx4KSAVv9bsJqnjsR0b4Db261reOcuCrMryMgTsZnhtaYx7+cgnsd6VH3C+3
u4VYo32HaSEPAeRteorp6GrGjxuQqeHNfqZvxBsJlSk4JCOnLFjcNcxmtAtI3oCjzU4ztoslw2oV
MHJKjJtePbS0uMQDA70pooSMy2Yv1tPOVei+pYOWHj62NhmVVNQw5QBCZCgssG7CQoKthXPLil2w
JVTn5JufScF5WCpSCiKuWpjK7yDWhj45Vdf989IWk9VgsICBMsuFF9HNkb0lcJ3vE8HhYXuJ0ZLn
87AkSntRX0Pf7JUXdEOoDETQxFEUx0svsiZQJLh72QMR3HIEB+tJcqRk4wi4qgttMxaXEhaioK3I
O79WC7Iqn1rFEY2WdHU8Fu7PaG1Nj7prW/nhDs7OybnYwTaokMab8vELpTEqUSCfacVEPxZH0h7X
LxfgJ3vp1rcohozo4OeURHGLCGL3QjlFDHz7BcdJH/bmFNnehYqXK+HYGZX2RuMkrY5mAfeJTZmk
8L6iHGN2EdPs8h/uk054MB8tevxno46xEaxi/AG6PDN75wXpa972dDKJ0Vt9l+lJsBiTEZRBATTE
H0apSMCyr7qTUqihWtsONJ9k6HisctBjsJ7qmM0qhJIobf60AQ4IhwtXlRJGsLnj7XPs0LZVCgJi
tPGoxjh1p8+eOVP695s5qF0NN939jcQNbwgV+9bRVHFce7jglZkDM9zROclTa+P19st2mExDQlzb
XwEYC8U0MONuV/71yxDGd/xhJYWOmqDXdCLpV3+Z+vNsIGbnTFTmBc1T6OgO53/jY+reb2Gq+pYn
y5Pw5NBMx5Xetnoh2v+CPQJrV1lKY027eXV2uVfDLsajtq3Epu0DrucwnQ6PiiWSy9TPqd43WEw4
XJudq7uDpMdfCt88PMkGY7lIvWdBtMJemJFEJ1n/TXxcbJ082IzgJOSX2QfnyHCozthe2jRvR55U
CRNzFD7+e34DLtqp2pzW/C42JVw7eaQUmZH9brOkOcZzW0gp1eFA4pRwp0bHvc5o9Xw5p+E7jjGi
VAfQ0GMFhLV/g0wk1lSX3cGlffWi0kSCDjeLYpOThmraq9Z9SraqYy74gxXxw5zAAwB8zQd0YqDl
8muPXwBlwLlLZjZIQDbXyBWWw7j6ZsOorBcY1dKBSDyUqp427BYZn6CGPAvdZXcu/xWnL2Wyp/YS
gXTWqOL4lmxezEwBSsnE2V14jC0hVaAU/wdtBOlnHQeBrM+0HJk9+Wr6ckSUUkdLWtYK5oX8p6cK
C2/kq9gG3h/cfIAd1yE/qemP1JmxK7JUouIxqmJH+Ws1En7lFnbiC0pTbC2u+mLDHuqT56MskS62
a46c+95/Tb06/gKczwdz2Qqk+2iwYamDvPp+flw07amqRRMwbPTNUO0AeV3tywu0xAZtC4RbJug5
if65yMoI/tOm9AI63IdXD9K8Q+O9Xzlp8ldD2eufLJaewJb+XmnTLNSDGjjiEN3yx02g6RUxoa7A
8KJ6zGjnM/leuBD0Yh7gG2u8FdKNisZUbdgh4xhXbzh8GpqK8TLQEOVbmYW8olZnCKKOanzzJY+h
PJ9XBXsj1Jyys/1L2VtpGe1PLikcp65G598HOIav4q4FeZZfL+jhRr+H9XIFXdd63zad+E5DvGhW
SfbO/pdMdW/4szoMoHr5fJAtPG3pb2pPkNG1g6kDtP8NQHWRHS+tYlsnU9CpmbwSNZVDGGkr47aa
sqlxjRiCibg8TN0N26ZV/IJHr1YTL3sGUzuM6sikKokBCNbAIfYiwHhWCjHY2QtCxOgz7lqjXG2r
7c5P5qE0BXB/m17CrfEL25Rs3jlF2yrthIBZWWFugbpUyPJwRH/lS7fc4dCEWiBKHXSM+9yxRwyw
SKKbrWR/Q7csvRywJodkUmy0dGx0IyAf/1Sogzo9nCLyJLENCU6r+bEf7Pgde7eZfymfisT+yddk
/7t74sAKZv/XODTgrkltVcBM9oZHTkv343qb9rtb3EIa0wqMaF1FXrWWtNTOxQl9DsTx0p/ACZXf
NtAtjO8PBN3O3D4DGM6QoVV5NE/DdPwgixyoQkOChmZYfLEGBo44AJzOWrzNSyFhp50bUJ9s50ux
5MafWDr/T5dabD3xCigqGjlBnYokk5IZUs+phhax7bQJDjD+agNkwyQV1P8sPYFGV0vr1yFr65c2
z9QmFybG7b/crw+syGDyNg81BpPRdrpOrasK70vE9IJKXvYXFnFoDxVv2mkWe+x8ZoX8H6yrMN86
/MRqsg+WuRD0rfWVDwSyYHEXC34E0VNVz7FByx3ulLW6WJop7VMHhQGSDXgDcwwP9DB0sRdgNuxX
Id3b98CLgPV1lzvpFD5TP/ixFa74vOxd1ReIUnqJuHq1ZA/3a0E8tnr3lccpYqG2dMlsjPuaWXzA
TbkfPmvWxZXCn9yjIwF3P7nZO1Lq+/86XKCfj7ikzOBWV7SCyuVw6dn5DJlpnKr49EJXv1r3Ssju
3CiM+F5q87B1K0vSxyXbDVt1PasylgCo/kWBdGeBh5HYdcSFXq4jTithezooudmrEkMKA12J10v+
tAVSPMzEoL3RyDZ9NBDaUzKCt4dzLoirOYhFzKHXOlRUIJ3PbMu9Ac5g+QwPyR4ZXclsxePg+/wn
tiBpxpPUZXdi+fFl2/pWteOSt5jEDPiGuukBUKm5LZNLN4mGVMui/K43ksRcj+dqXI5u5rhTqBeR
e3oVz1mnXuIYF0g4EtzjCObYyzucJSi2CavLOGXCVl5h7uBg4F7JoP8nvsxsi2y8fJqCfzZfL0Nq
7oaJGW597psKkD3exOglYD57q38v1q91RGflaO92jnxXGltjmt36dMOAWoUoiDCUlGNhlu3rqU4K
MTrxNSDyzNUIW1uvApUBbdLPfgJy1dZXhWEk1YGL9Mo+zYFv99+3d0HagNPaFebc4MoijKctohgK
/HJuRRAK+X+CjjtCfgLYYejpRdZBlrJrBYfQA/xbcB4hSkLfPcAuMG0WbWMajKJvGEFnXP2CVw6S
1T1kWH1Vf3Wr+PA4DHpoy8DlMuCBJCd9s0rVpp/wyDcs2/42zTZP8pxm+t18zCtugkSXajsONoZS
aSV1+TONezK3I+m1juZwKNQXN1ccOldur+RmxQGn9t8+TionEnjGBzlbAOLRk9F1Koiq2GqKbxLY
X/oEANEHhWlfuhzief8eYP62L/xs+tEZl8IITh5cgKxpoUTPAybgV3HrZwNNJWBI3qKbcYB3InTT
euJWNosIV1h2/F75e6DastZWWWntxLC+uAvoOGk721+LogB+gzEx5xQ0UxB8TucfPmjaKcJtslDT
vX+Ham8MOOauehb1eiA8xQbn8hgixm7Gctvift9mYp8Vo/IIsLspTVINw8F0DN4G91hsI5yUMGsk
p9CZ3FlrnTtk+fZVvx5vqdCZfC5ApmZgYwGyyORrH8uJUVLpHo7KPoXaJdJ/QBBu9VL0B2CwO9ys
TpTLgiRtMB04ISiX4Mb6q4I0oc5VszMOuHQMyM4pXK1g1yiB/ibdRA7ltUYOu41Q8qSMRGplM81E
1Vq032/yKKszF5Xohc4v6lFqOYp5yVpFqp5tj7BWULwp4YiliFMl4AtbnTHAvgn5T3uYpf8R+YUQ
MeEgQiaCozeDG14yc2YbMzody46e+NjkxQlrLHXZJW0/R62vkawyfnhf5GvYSJISnjnb7uk1mM/R
l1IP4grctgNtwjQU9vyn286vyTPWOMviLn87GSI68rVbEiQ3IEe6Oukb8wbAkwZ9vH94eB2OHdnk
VXS1GtNU0eJVeMZkSwM0/xv1bwIkV9uczf13mIhZt2lDE9b0efHcJfROKLhZcmKipnomKwkx/voq
cyjFgJqrMMl955X38shxh2GWxB8K5W3oCgEwBpwZ0LMAJpcdqWQmdZj2kZ+D9A9k3TqOhV/nja/4
7w4qn3VBonB9sj7ZmBIK+e5NQl+/V40yiSBWYaJqmxVouOmSAds6SWEybmjrzGM8YDtVgHkBfITi
bmi25IQSSFfMTRTCHLqyRyXb2JY70vnH95vnlyZ7N6G88IitF/B3Bpnu76b5h8r7GH/oqmhhNILp
Vtog58Kz8bjtZ+oKh0PS5e1nh3h1WFI82V1+hsnOoKxmOxDbNSFPJWlCmFT10EQgh90wMXbDXg4K
2KOFUnBwy/EMIQ1s1ifpM5QBPl/bzbbhgjP80HIt6QF9GYatrWGFIilKVzW4F36wmVAtOA/+LhOC
xUjpA3IxR4elo/X+XPlIoibvyrto662+P+hJfxx5T2xipX+Qy+fyE367ZxgVQ8Q7q7yaaEBvU17y
SFGzPrM7HSX8V/ty9QJf+x6A+NAXNB1nGfERFrraD2BRU6su0ZrCpnUnc4uzDZCzKldjS/puDl/d
ECrHDRlI920fEjYnjHlupO3Tq5OJDFz1DTKwiPHNAOkLo2lByG+ezyhsyF335lDd8WEZxIIwWqzy
PtTZtqb1CA+OcFsjYRww7QcqY5yqcrpPD3oH7klCkzvMsfUroi9lvTf4L3JA6bPeTHJZPnc1iFnl
5skdpwfWhMM0xkQKeF5Vmn857+uPEu3ST8feOQNYnvmS964w2N+UY+VjwkXY6Y6rstC75gzvEH0s
AIpBTWh1NOCC6Wdz1RKE0Ur5Qn8w/0VUjAbHxlwm/zNrDxWshA1m8nvHSUaigvlD3UNctSuvHgEO
65cX9x7eLK6IMRn2iDNeeMDBwP7r7ptfN9hcnfEd5K83xdM6dEg+MGTnHvN4DjMw/7MG7ADT9zvc
Y41DmbXd0IpL96Jvc3ZsDhDvgOUoA7qb5sUDjo+/o/eKRkuFrv7z0J0jvsNJswIxmqB78uqkAZYC
W5yu5O5SOwkcy8LaWQLeYpn67E/XfTbIohs6yHzIHbPaiPR2ZlC2L+ZgOF/rmRU1EYMWZ2UGL7ci
YOAAFu67EA+pfVpZsEQTCphQaPcX0OtARow5lcvImPFE49mUHwVBId5oUO19sXKMyxlomMxrqi4/
ds5E1Bh3kHXw0V9KGumA0bX2VEoCR0hE5ganZgaZQG5ASc8+MHkf5nhb/XcSBXoli+zpRJW35jwW
/xBz22Vj7LZp7MJtqGJruZL7clqQZ84ACncl7pGxJWvCsaT6dZKpd4Ehu+Je4CaY42Tx5QESas07
6NcLr14xzWTiuk60Tblk0Ytnh6OKZ8NUaFwpm8y1iWI52vupgrUp5rQZIFF1LfJpE0NsuCHDFbvB
FTHtDOu3ursfmGEop1dZ83pegqtpq38K/FbtvGuCjmsb5d2aJJepX73V5sDjh9sUps54OE6mGnvJ
wVIAN2ALreSejRwmie5VfvXkxtZY86AGHKyUYLkV1bgQGwLxEu5QzXxTalTeSpqr5kaIHE+lyjSj
hsiMCla1CAQRgvdVwIoBdcm//O1NBY7nN5VKT1lVQ7NIAlU2XzJuWuANKFsHsAH5CEzKHJcjJmlf
Ryv/Z/qqeJ/CVrl0a6ZlyDFF0Ld0M0zpyTgLBHsi1h3EWbPHN221OuZ7H5i8l2Ti4VGb1CmEWHZR
5Ijky0ZB2AQDr2jVstgYIsRgOuaCxdmIhfjXxy4HGtSvwv+7HkX8KQgeVfaAC47k+XdTEzhAKs2Z
MpY2RlfCpXA7xDK6xmz2W3ZiXXACrL9I26QeFfURQaSFFgR04NTiWdDiyRGI7yofbE+3WOckj29l
yaMfK8DjWKYmDjA02Tgj/ZpaGWbmjk42w6Wcktg6T9iZZJ5HUnAXostKHAy6HP4UON52qYG7a9Dw
f7YmfrERY+Lde21Hm6xAR4yaBmfKmRJ6v0uC8S4Qh8gQnWJdvOkvIGz1MposLTML8g1ngoHbOOWJ
6ruBeMTUZfZRm7GpQWjsC6S8sfmHp8npSUYHESXU8vcUWElThh7+Ae7w2rcdLIlBALIY+F0KtIWU
SXB4qeVY1cjn0BtcZSdS2id3QlhlefaKQh+nuIpdBnZrszhUXGqonjikeooACk0gZeF9mpEk37RK
qtwcATrAalRMHoX1ztypg0oqzqTjfM37riq+X0dlquh1JGPVk7GJoxQDUG0/e1e4VGdb/8jsgK1z
ASCfzz20i2bsrYCB84L4pmISvbSPJGg8QloiWWONVItjIaGUaZpQqVBdWF1c6BvGGZWzvFNETcFg
wX4NEycjzZXN9s+EwrsafyRf60am+mjMvz8lnuhjwuAWTKjCG+AkB9WUtHRVPe2g+Qr//cLmMAig
8o2RJm7sEa0Ud3bbDP8GyOoWu3hcnKASqJzL/p45mTc2hv8rfh/Pg4NeHwaID38BsD1nEI9C8FzF
KQYyo/YdQbASNLKyOaIgz2M0etLAhbbDyz6h1w0n1uv4SKPVy9iWKDoYoY9dlhmifH+3fvugla7j
GbZRcQxS9zA0f9jht7q1GWBPuoK30p1f/kjGWkGalD8XrXLbRdCJdnw96PFXs18Y4VieaCG9Tbdy
2x9r/icftSaViru8MOif1yDgmA9VUz3tshyM0oo43rYHJXz7ttCGhE36xhlYB3frojgMIXCMAsbe
vz4eYrzjaotg+sY6bVibs5xceQKAhsoY6AH1LxkFD9U3FOxSZMjOT/b7A8BiJzGMaHwuyMxxNQk6
fGrfLOatgSskUy8/EUY3Sg6q9KdfXlBkmPPMQaUX9BbouIBkw5Iffokh2JaDqFsQ+0NjaGu8GoZ5
a1Oiq3MuhGBeLG5UMPeYg1jMyrCIQ1IMHrO8ZyP+h9V4fHlEd0WA6C1fZ9K77jk7CMxD5KzfxqF3
i/fH108BkRRok4sfvgWAddQqKe0xKqHKQIJcjEiaS18amQpVwWbta/ihPMoPgF2VoVeMi4W7MR1t
yngnVpX46P/QwaWE9lOMgYWgHTdyk74eFDVVb2txoQJhF1sqwMdMVdXdXNjDVyWOgMQjxH3hMOmD
vCXVz/YHcSkg9/kWyYAxDLAtaOw+8g3UGVZT9OAfnnmkaLyYxMcNKgnfBCSSP0YvHUaOvzBghldP
8LtBG8heA2TgUJZ5nusaklTteleAEtJxarpGlO1vXIhvDJJienPIIG2WzVpLVIDKrOqroTSIjCDY
vbjBRydnW5eSAvQI/waoEP8WHJ9URYSpRjG2nf8cu/Zs1uUEL5OfJ+1sZrU8ke3lorIss5VbY2Sy
CWwFXjBBS5fAEIeaZwEO3UGqAuN3pQaG63BQWd3R7cr9SFz+NMknrMMW2FtlZvrYz/GPqAGoQwNZ
yL1Xxnbp7R0RGsVtwbSSbBk8lYiOMG/HvPUIvufhlJ4rJEwHyfSP/ujdBaG4h2SLR54WoOe+WM7w
j+SYR5nf+bZj72edY+K5fwr7Ax6Cd+gmcLC9FISrok/n1AL6q67NROpwpKK72jLC2lO9L6JWVLj4
9XMOhCuJYsJVkxJ/VLXC9kq6iyydk1dlJx9SrR4vP5lzeCyCx2urAiVdNQujYqiPLM5A2xmvDMZ0
evlo6ijQUrw1cUH9mkjoEcZuVLa3KuA6uBCEugTe5PtcnPkyvzXGqOouTFheERdSNiSEFr2G4pl4
hkAF227iN3FZsQ9l5lALWmaDfRqrnpw8O9pZP3WaPyHQq9JRVx4uBD/+0kMI0OGWfBHUHRB7Q0tG
R5kCZonuwyuO7fMQnzQX3UZHzWSvsqV23WBZvcmBVruSM2ev4HBFd7Da9swUUbYMWww2QHLLHzqY
qH2DisDI4o2m27r7Hb6gW0CHqa8CHaUum2b1UVPXohgNtIWdfqtunT7nsdM+WV+cWVJ8vRBWpkz0
V3UsIZ0q2AvlHcyXDR9DyvlxgPxLZ4I5n6FsHlxzTmHOo4DVF2Wb81rZQHlkbJu53doz3f9IN3/1
5Hhq0dQtCMOd4Y66MOEBSWthjjD3/HWfeWPEiwy0pOkfozwvOoTEjEmxybEp6aJi4SrIb5QxdLHp
xA7UywGapcThgL3D04jaNgQ4wI74mC/SjT/iUDuty40Yw5JDSOjfW3oW7c+upOtUwVmvNId57BwD
xf64XuVdyXcbBWenGH7SneyPSRA0jF/V4Gl2CSYIc3k6mTHapUIbqecUQzTTwZ0U5FyN9b+umVm2
ebJlxgZm1fSS/Tdw1OvO2BoFZWmzbyWEgh0IN4vSRXrxqGzwFgyYS17+j9FfQLgkTtVRpkBL5/BK
BQrrSUhf/TMJqCfKatfqdjz0XedI5O2K9eMplRltl/4c6pjQyB9bhH+TZy0hFgRlF7PymV11NUxX
bPe7ojsa3vMWptPQYvMtHblxx2g4F/+HIHmnpl5fq11yZmPHKdw0Y5thtw5c82cD54qgli2R2B8e
lwcPgrzMeOsxvh/YpqLI3fwi9e52zWvIWyKajDI3UhPghfhuOKEyWqa25cO1XoHQquS1nhjszp7l
uzosH7IJ75Bmw1fpIEpzMJuNPtxcj4xjkkKwURn30RwwnTuUez27zYvq+Iv3J21ADln2Fbu0dw1n
IzXV0pX6gw51LIqgZ6mEXZq2AlcDKU9x1MMOER3HdMRi/eE/90v7l5YPsi7KeVyps6QMjbsATKnT
OeaLsBTuwGprwZlVCXJ42m5s4iO9KXtErkSPHzzADjTXF3DyulFQRxbb4ZGsYCWOb4aEXzl/qIe2
MgV79z4PiQEmQv4cOorqOEox1j4K8ClfavTJtczKhYuqGT+4TuEFOgd7DYgrfZFYpFlQMeT/HE13
EmKNKX3tR0wmw8yobpGpQaV2cniDK11GjPM1mopI1IUTXkpZ4I1agNuVudARDD8a+MMjGsO6UFZp
HOgPjPxAvgbHJc4I1y68f1EoOuLUuBZeayg8sNMP29PtqFZr8AaoDghkLao37FqBxpJ1DyK5X4oc
2lHoCyBo0WUoQfHE24L5p5lv6xT6MdQv4R9M9hBF2lGX/MuuVM+ZxoQYnKBvedhUrOFsAdbmv4Ex
c9t5ZAr6InMspsxMva/1+0sN1yS886jzW+t064y8b7iMIqFc5BsCA2QM2ePnj0LKBbSJ/EQeOIPg
AbihgcfpIizTJxOrCuoAB6p8diSOkK74WU4LcYwco1g1pGaKRYdU4j3d0UiC+6cAgX+CMYeVWlKE
KO9D3sqYg+h+oyEZQuTrBD1i8Phrd+CjsGDvRb1v0XAgAJySvsnWcERqgUoZ9ZpBNwGFRbPaeLaW
731OaIu0392kBmHec3TK4ZkymrqMHGuYUt9T7rKaMbQnTNtbaKy+aPLCqxhJn7e577UDrA+nLBMH
NpBNGV52mTSGrloVkoZ+ZCeUSFOYDE8oqevt+JbuIq2HZpRIafUygyXFbJpTQXZ0Fc7TZwL+7MLX
3RovhxM6jq9hQrIRxk/R+c+Xi9Uda5JP/WgTY/U7W7VLw7TLslCFJLYWY0tPh+QE08ND9iXgzn4W
c82AQCY0ZMD/PL2JZT8ZyRqp+VYOn+T64mLX8nwDqX2SPU0xYMInrUyKVeHnxV6Wqt0GUMAjsoUB
rjuIbUDsJd3vh6MF/Is2xXfrmkelnvkzDJI1+nguubQz2hXJJ6QoOFGiW8aoqbXkoBJ0nE2BxCOw
AnTs9pBLKVyz5KslRB0oXG0ZLhWIOvBvGKUcZmr7IB0FNQqjvG/4NwMdp9+4xky9JFEUrTcQswDq
ZQRqZeS6wil4OT/VTkbB2uvVzTDdHxw7BH8Iv9ZQwjR0RTwOyJ6LmcAJ3zFfEsHzg6pDCJ5cDwOQ
55Ezm8Hw7KNJQEVfPuE8bW4Fna80t5fnGtUTQqPuhmtNYhvIgxtXYAaicjybYEMk/tuI4DRlw6kq
QiYsySONPF/+aQKqPLRZZWyMdeSrMszVkH5SsX0DD4r+7Goc89K9veN/p1g8S6r9bFn8uEz7O8Hd
w6FCKHlx66l+oMuBD7Omv0T2wGkK+DbxpAO8gBlH25HINsOQVBnAONrl0hX8NGPdYiTdg6baKeIh
smPaQo5Um6u+zQ8afbf9VgnkfQVtFhGU6yC2mCxqrab+3V7zyzCGS1cnnKrJT2CKLCAvPCzWqqlB
4KucnehHGPSDm0HS8A+5ECyWwbhOh00t4ttGXyxlhBZ247zLzwZS2cOSzSdBV3PZ2MCLhpOI/LP5
52ngAsQ2WuTMdOg8pjPaVD04bVhmSRGdRsLBzfqhRY2MHNg86YvndoDcR/JFKY2ClAwwoonvUaXm
v16YnfrBFupaP+stv9djLJJrNs0pisSP5/yYGWBaRQr0l4ZXZr9HQaR3xgmw5jlkpbG8QF0u1Nbg
JUCH3msUlgKazDf6ItPbhJpnVFDjdACoWQAoAzlNnfJgs1b0T+kNtvsd6XgtuqAohB5GGNpQ7LSP
UHmuDcpuz7TC5sCZMOw7y8nL7bdDUUty2CryOKGO1Yzzd3cjTOnxybJn7nSAzGFpOth4WVH/0Nbv
bhcO0SQeh68xqgZfq6kqq+oIhXgoRADHt+XJVp1GF3xdHBoXptqmI3cGVkqqj8882sRa81UJnwL9
QugfQ5dBGwTfj3wgFQyZEWfcAMwHOt1tlaaWeCshW7sDH9oHiRZXgDZM+g0MYLJuvIfqwAHUoe3/
5lExTAJIFJK9nWw2vBcmwHNN38pzgVpvjKTsMBen+ck5tvX1av2aup1hhkJ4Df7FcOqdgbh+P7cu
RnKVcFxaWlJ0pkTCgrIg5jl7oQurERwCWrvpMEY/Bq/m3PiFZJvPvbFWkipMwnU2uiO/1V8F47bG
9Ew3UumqDSQaq45RxsJ3ytqr+l2IrRnTAY4ZSfzGw255zyJVWJ5XTsjRTDeHcGD15PdumxDLB3c5
gHv0pOR9uo//C+GHiBS/MJ0py3q1UAmqm4nHKLQxfTgOgFlx3r8t7kHDKiJMCc9o5NWD76n1Xzc8
nVR5tHDM4pzwd2QEoRT8LVtaOS+W514DBbIcLE1QLG1B+lTr/82KjbMxMKFWT7W4RnZcggyg8ifT
XquH0GHiIW64QNgJsY+Tp7K3Wfuvvfl0oA+1QTvC8M98HywL7D4ppE7s0K5WE/Vo/wiswhRNVpPS
0tzdwbzUcubGLNRnzUp2MPQWhGNeJZm0KQwezL23I38SJZaDZO0ekB65Gae7xmCmkwDBA6AKKwK8
YeUkIX8TiQBLdOXvL32EsSY1CDrq047BTG/LONMn4NmviogScrue4uTdftbCvCrByn65dONdnlPu
kIyyBLvv3YonJXppixEtLv7NITi93QmJHqiR/YsjF36lGz/JBTLlUZYzlFV/WNXz75OaeLloLWoM
wX7+p72+XQ0nsnrvot8qFtbqgHAgyKa3lHVZH0tsuxioId39RLM1p6UsCUUtF0nslr/qWxcgTgMT
gse4m/UX92QhxAvYApcevgrikPeqfVRW6IccUdd4bjyGfY8nn2fSrUcEWp2QdUtNxPV7M7Epqk+u
+u/Cu0s6bGJTUfSln4AsaV55A3RuE0wbu6IJDTiceIBeSUWa/Yu+GC+tQnDb/LPmqXm+FrRR4HOG
sHybtdJ0zr/f105Wt8otOFAw+LAmVIaulJm7uO2j3TxtmZrr+3Ly8eGcPcaCH8H+9JJmWvN17j6p
la8yOXd2NRuCXkzZR67gonObezmMolxbZ1XDVb4CAxSb5SjVIqdIeB5tn+AHs+rQbQlDV1bRPN89
iFwgAzWDv9+9CiMKQJjJcPjHnPRgZxn7N0cA6YnbaGAnmsY0ATWDrNYWo+V7U/7Rs7WJKp+o1vLv
9828DZsj384h06tdOuSMFlWd1LpZP+JyyYUP3a0gVQyrF6weGeyF0pS1+VBqW1Tih4Ksa23hG2hi
0N/hEmRegtIiVPrF16uU1yeK0ujF6jabXwrBBwTc1ECh7HR7DBlhJDbI0Ty4aGlqVnazsEnKkm0I
ZfZ+uTBMBq1AdX35DAhEztJ1zqYUkmqQU+sKjjyIx+LzKu8bnyBFeYLsJYuG2KftGp7mctfJavJw
sCMFT2GjjaVcgpyiz+/DBTFbpsdDxlp/SrU2gTKq7KhejHVpIFSPBPxxYJIS4Vq/wEUPSX+iyHFQ
H5dCc5ZirVco5PZllz1qGP8m/frwFRmvSISxqdpg0L+s4dvveVn4fhvISHkqtzYxgU5dIPWWjSJe
qrgJZYtMnZxI7RipRc5FJMpJbOL5dLK6QKLv1nwN5mW9RvxCdglzyTuOJuT6nZo5LPdgcVTGjXpH
78sCyQXN4MRuDh6J9FOOu8qKN2ptWYY498l0PscebKCYesa3dYyXmGcrt8wZDJFyUOotN30a0BOV
fRg4at9tPuduwqnHBShfw0zBbv7l666IxK8ePFDNW77TJlcWruJRogjpwtI03ZmhC1XHjK/jfGFT
/BWKSnK1JvAy1CGm0MhPtNNKHdgVSOynvtFSSaZEXay3PZB7gSto9aCdBHsb1UvHmZgTx6SzE/CO
AKufMERVO6dR5OLq5vMJbTmjyqolPGZlZg3p5MkSbvtFhsPFCn8lrnIK26R5ZO/ipBt6kvGhZre+
wmPL4KaPXUaLyKfhUwM0cyrGZXMYFYm04hLRDz8LPkxQtQPdpq6imrLxqqfoPIbK22fe2IvfmaoZ
Ydx3dKQK++BjDS7yaZ5xzCokqiLWPOGJUNS9Jyzr9PnEeMls7InCN+Enwzu/rahuw+vCPKpgHCXL
kleTtPwRCDPUe9KOBPF12H+Uq3izdZvCFAK2n75atsB94uE/243h4eBZkgUOD7MngyQG0iW7y7jd
pKipOLrDhWr48UC8n4r7uSvFFeJoTB5VqmoKA/tlo0DrWYu+kzvYXYz9XbyMsihEckAh/R6o5bTz
evayeRX6C9vezVi+d6vQsFkzu6qkb3sM0w7B/eLV68fhofKVWoOwrFzOwl6YiJ0ASJCKVdRbKS7/
UeBZVO7kU50X9Kkx60JxzczV5l0b14Gvs2Y/pxqHnRZh4DvnfXGufoWU8DJOb/IAPd7Oo9o82fVy
S43dTJSOlDi2FO9LX9ej49DkdBYQ0J+3RF7irMWLt9OXnjfwqc0OPzttwmylie3E+zOR16H2bP1A
fN2/oZ74fmUQ1H5PjLTqiTB3Rao8gIs0I0ql76lG5P7MIyeoKXFXtE+4kbkTz3h45tFMHdRW6431
POWykTDfX6P45Ur2ENdxHJbfGiZmXwxaqObt9+YqlH9zIDKRhseENMvGlt2A1vULHCL56j7THyuV
zxUWxVmPI7z7izFAytDdWNTV1hwyfTJFuBf9Ft4/PG+qJgVnk+0UQZGOPKC8k0HzWn63TUwVOvCG
CqB+CiJJ90sglkgBsdnaAS/7BCfeMgLWpEYDxVEg/tRpWCee8X5AW98+uKNO/A+CwlQ+jRRiWx7V
kPfZh5yBbDuro007dbDGp5l2q6geqcvwA+o+3rq6n4+fdiskpIquKMCvtLBPXl6ECP5OgmSPoGGF
x7ThuXYdp7cBuIdBFhNoX5MCxMMGfLcsdJP0YE9uQRKd3MxUuQom63Z7e1GHgk+7P4xndB2LU84o
ZLk1rTL2Xvm9wQC5rLDL3n7PvbAUdg9JN0IfdcJ65ZfK+zxoUPXW2rTiWDBkeyPHWzRZTDm/hWpa
JdltRUawsixebzqNfBBrBIH+BBBn+yFF/dSV0pgNiVp4zKi+X1KUDm+1okkzR1ImEyejvg93iO2L
xgHdKFSSRps2WIlx3tG8txe92Lrx6d0u1O5LQD+H+ION35P7mPUnTwmpdsoXNokeABcSouK2Ryfd
LskMo289pm0cNVU4grUFU8wZoMB1vKN2fr6J457pXztigeXVXYj6vtMUDAwz5/cVPDkYrHlAHLfo
eH8TwRmvN+mkgb8bW6dMtB81x/DgSEFTVN6UDxtY4cvchyvMrrsFwari7vRU1vLJPjAJ0opNJkUI
aHnIUPMkxdVpnRmdt+cxujn+2XWll8zXG2wkg+zIcnxes4u+iathODM9ycq1pCnII7ZVDsu0F2im
eeerJOQyi8TO3WIl6Jb+T4SKGWjs1BgEaSKwvQqdua/c7qXFUIMwtJTXC8fzW5UxKYyqBxfETvL4
6g6QsxiHZcjxyTqL0z2bhO9B7WujwYhwAoSrxIhsdJ/tGMxT4n3L4r9s99VvUnXVVh76D4PmWoJu
7ha1HjfuZL5mf32FMj20b3+NprGvG7eZIHfw5uJaODtGHOv9Ld2Azi8aPtzTXQFhwEwjtoWx00Q2
+nwbOeJcAzu7gcOPW/tbnYC4G+0zzrVFoSw7QRKpPDAFOKZhRzA1LrSuAJlq5GliqiJjmqhuNgyV
FJy9bGTD7s2FFte0dV++P73hlrTmcrwkb7tBSDhF1ctvZmqmW/0jts+G28RuwsvQyLNZD5zMrbDX
w9eZfx1hF8a6V8qlMPxwQjuO44+7VMMyL+fMQHiMCLjtdQRjlCQOiSK5lM/MV5tiF5fIbGRwj9qC
hmhn36PrwKwv+q7KkhnVSB2x+acFPkPgnc1dXvTSXhg/U0nv5/h13OC4lgT/1Lt4ZFkHvLWBoesM
23mi47a3vPb/XFpHSMJD3MTpX3UlGx44bpUX5+z9y2pB3+FNuHoLVk2ugPHyzOMfgCzVWStCx4zp
d6xU/w/7JZJ//xyvL4k9RPJO4ntFDUCFcwbMKlBcYM4wmlBqqnXEAdRacga2c/UiMCvIYSjRrCDd
5MzbaZC7vnIjv+uJiGobJXXzrAOQk+xBWwvSGqQwKEC+y+Y81UctqGRfWc5BJi9iFggHkfS20Hm6
Lwm7PQQcafc1y+Wg8sxBAdZ5s7v3wfOB96AhXU7FqJXI+4KYYukrn9a2g35h0kxirfP0zBPn6e2u
QmZiWfwhmW7hO4SoOQBpNjuRMiG4vqI9enPOOYLVc9gHo5BfEDvQO9FXbTNp2ka8T4HceQIBQYkn
NUbJ9oizFIxXCxEqLcQUTHuUtzpM1+AHx9/qKSD84DCWZpShj730NtChCx9VmFYS54gMd9INgRB8
zwSe9fJbaUzT2TfDyLtSAcP/99LdNkwtj8zipvZZjUxWpJ5FCwEBGb29947ykU8fWNQZeiuz3g+y
EMl5/9s4LmDEpj6inHKh8lnAhV7lM9F3PSP923g31KNBWgL6VesxWtHVva//3ThUzAakcCRrDnyd
Miet0iU4kVuP9AxHsA1aV5dr9AxRmwBxeOmVL7s+swm+NSNUcRlhz1KiQ3HSoYyrHN/1ZtbUiwUr
1LcBHodu69msWyXVk7BWCs9b90NSk1z9mD3kCeairnZUAQdeThv8il6/aR/BFzaFiQvEeGwxHUuY
SBh1TUv3hWska7lwzi/FPYljmU0r4bClHMSJJP9aFa1SAbDs++HxgHlnhlu1jR/iTKBLEBJJ53Pr
+OhWHVJ/FuP6IPlUNut7FNMzc+pjw2jAhMIomxmAi5iWk2J4xpb85/6vUoCs0GYFKWPjWiCmT9WU
YzM1i/xD6l1csQMOH7AKcnQ12bO0KpmvEGI4H7nYk/VNuW2gAdk7MYPl3daegMyLVKhl0Ug4W8xR
3zdE8HvuRA1qtU2DVnr3sqWnu7af6xUcTJ+2IbJfdTFyz8eisIsGl+dE8YITVi2yELS1a1bmyClA
4ZUC9cNj/3UR0l8tMPoYQkzyu9N4uILTz/nYdvsuT5ym9DkspXOqnpnCfFXMGXVr+vhj978EngkS
2G+W0SOxVnbh5tfkpjKw5uAcsfkgaCT2TaQrKuW7U2lxyaMoTy8z5XqkHgkDqHknR8K3TNPn/4LX
1q3kY1mYhBrS8bwqLDmbo5JgaklisJ7s+Z3BTDzeyJHO4xoB8UkN3Z0L5EnjuruLWAgwabw39vqF
7xIqvNxdL8a+URwfuXwf/otKDwXsySwOnSp2l2Jziw2m1YRZDN0jFGYrqRpuy1tc3W2LpgpagsAD
cJqMu7Y5RNgWDpWn9Hg13HRbC41ITymWpK3ELZA8ENhfh3P8Q61yYmgCqV03hfOqWruF5PWKvm5i
GTT70qU/ZS+WZJb8TYO32cNyqkweW8BVKrMbjgU/Zfh9golrHYZt8dIdC+tDHbcw8udA3zXz0KnI
g5yp7vkfIE5XgEHLMI3I2i4mE/U2qkYVfug2qtsEKRB0wmci462IQaDUk0ehkM98/C3ijoVSaU5B
lNME6QWRzLC3glPVVtL6nY4aZMGDSVPEB7MHf2mmI+4iqLvnIEM63V1UA95beoHZTCtlj5Vs3Qwp
tIuJY/eHu3oqWeA+VCqN8zaim4reCVZLIi+A9/wM/n4k3GsZMvqOBPPEfa5FJEipsaIblyuvlalG
pkUsTvNRBVRwqVvfbV6+rz3/xxRIcplgwDLUs1BoF5A18aEWiSt57AI1tWShtyCWIk6wTrmicdoW
Wm/RMg3scviV+fGQiFN43or/Mm3lmmB/HCgFSvxIn5IZcqg21jTn4D9r041B12hi+UhTdVhVEd6Q
MWQEc7et3qZdTNkbg8QsoIIv/IBu2+XskljWSAmLBe68TfRtYDMqZbvzAJDMQzAxAoHOvaIki9hG
0kQz4cByJtC3qdrjRcKOBnm5vsmUODpIFbaXqDpiDMFvOcz3UdsFI2/SthJJvm5tzIJnMGWMr6uZ
bOxIYXVbfxsrZRCSEBuogGaHb0vfH+cUlqaVmdeb8u7HAmxZw9DpkQDcatxuOJS496sHtlfkIIGT
LNLynopBjQfy7I4TYkVB7IWdO223loXa1sKyDER3ocBeSJF04WAwwM+PEoEEeWNF365oNbeBV4A6
vgWl+m8KR7KwSn6IA4cQIQazDz72OKn4W8Ckn9AEWdXfODMXCt4rRZyARTwAzVnz3oFVt7xYUvmZ
WiNbuhSn9B1CYyEiOibKFqp5L6KZDo2/fG6KUNkt1ahaClLaiGKSyLlGqWx/nINEH8sMWgzglTFF
+QbIialzT2CbHy5WP7yE2tTy389qhgZZYuntxUIIGXfY2/sz/Z/F3lwpDYiyxSwlWzx9tg/QdS3I
vHDANAQHuNBYaYKWs8UJI4HrPM+2hq4+xWLZxN/OLM/IAOdLGoGVUcBjCbQP3RxSd7kQ2iB42583
oR9Eaud/SkBjUQ/YM9rZkQsRNNNCQ189luWgSJx92aPWLJCuZ0BrAimNIcr9zFp7AxYUUpcmmVZ5
PkwBQpkHSNwSNARns4mkN1Y6ZGVkS32SbV1CkS5C3YP4eWgyGCT1RqLG66YaoYKDdafyX/txBTzo
8Nw+NHDZ8GeW1azf+jiTdkxjkKG5/gtmgbxFRW8Tpn8UwMIkTi6e2YAI7rtxAf64jhIDs7yM0D+d
dafWMaKoNNIRiMrIKukmabxawlOiscOGLU3S2iMRTeVOk7qS0SibDvmW5LB0qQJexD9K6v7KEdgj
/bcNS4jxsB+6gsR9YlZGU1ZDCoW7UqdrRPUbbCs1Z/4xchZ/CvSipX684OrdyuPAq6YWK2LWUeVR
yXDVRigZh6e2XUl6zzaaL+Doy1ImhEYHwJapBgjhcKCDGDHoC1UlzKFjt5v/7rIiGJAKO2YxCDGX
VyGlROpY2XrFXajWg/tD7H8cmkxQZ2ov1ZyTiuIpJL3vDd27/irgYgSMRlSLfAQ6eQmdfKFSZ/DH
6N7G9ziVHXaW17bN1G2icoKOfUlJLv5p8q7xPbRCGry22Sl+Hc2OhRDt4EzjImp8WpJRIAs2FHzP
dumxfGir00WUqYfjhVE8UKVa4RU2E6PVm73879ReA+1sSV9WgahD5I622Lr//VPpfW0m7penYdDr
419urJ1j4onVF4vv1jVrAonuPKGEtybzHF1RNXPGIxFiaaQJtBfzjKVjhUSG/kvisZ7YObZojt8v
Yh7U8krjJRQnF/58v84bXrV1a9ig6RMkNJZSNy8UGZGtjbAzHteQxKzICLlZ1vsdpj98LNDBRxHN
PA8v8UgkJt2+xAXsDMKeDGOB6AGqhnUJpxfEQWswV70FCGY+UgwMmJzkvn6gxrx09JnIIAhW/Rx0
/tMMkOGFmSK6qIOZ+ftNFlVwqlb2nfYFugym6RnoNsbtsEyyw8FowUzE/CsTqfxOYYHijkhFRd+B
dwziHpqXC5LfquuUz3yMdtBkxCuVzZfsRwWvY422BTPyd1qPUxRdOQu+Oh8fKtfYepvk1UYhtwug
GPTs9fPQzxCVd95Ji9xWXQKDRSH6TPo5zwfqS2je44HOApSKQNqzKpFVQsd8cG3TbpXjYpqBpzOM
WKqlkK9eleLG40BRBIPfySpzwqp6apuct4y0BharGEGLfqEIOkeol3G1GvDc1BEyHKc3TJVNr1C3
F7vv3mfz57FuiIBrCwNfhUgXCWRzhVw9jBQCESNh5s6QTPygt7IdvUCWhCULNBPALF/i74IQAJg+
GeSnY4pQ6JHK3hjAEuXhUNHkPVN1vfjsCYZ0g3zf3CIXrBheBWYhr3GVR7ejk9HVWV8eBH6I6tFR
gOIp7LQlJlxo6EqHYtF9X6uLXBmdt57vOa/YHzL5VzmgUxQUm8ThrjgwxmPQuNfR+kTOEbGQszBu
sHTE5v69r8nt5vT3AJ2NCjFebWd4HajPJoHjXPcnJ/HaVjGl7KajaJxz0qa4PMg3KI5W5G8ms4QV
2h+HAoShWz5HNVDzHrhSjV2/lDNaCyDd6otC7Bo6lPUclbuI5T/cGUxSrC2o1e5pJ6lWSgQ13tTK
u0eeEYoFn3oh7vaZ2AiVezaGLvSyV/pHveQIDHAkYQJ5Au74t1sHx1wTpPCPxoowP+haXmg6Cvcj
ylYtHZpu1i+Cdj/CwhlJhQv3/wyneGkMUvswqknDWWPYgbYGGkKGR574qerCfr3sECrk8ooSpsLS
OlJa9e5fKLoE4qMoK35Yo+M11lJtlaYvIdxjg56e/k0gxFj9cwamgIqnx2rkQcBujsZ8EYYe9g0s
UHQ6/Ls839/NYzrt8SU8mnOvV/cmDfNgEOOlZPJjq/BKXnaJb9cmzMnQxIzHXszXZyUwLqoIP2ZD
zZ3fGfhUExhqGZ95CyC08T8Xqik7qBjgMpmvLhr0PFB3rITZpjQjduyIAm+1/tEAPeR9UjN+qSE+
L3dirqOGLwT2TSDw82q1p9WX3sO7+qtOy/IXBLpkgtMjaMUJsipiGxPbXrkA4gaxEVJuuxIGF9Db
GBDHLcobDOIsoqkgIUAPg88tpWwsIhsP4hDRRjUpG+aoT00rWpRIceheb05GRDZGLPD7CLydNHoU
ki388Ggd63uTvqxNWe1EDsIwixSEe1z7gZWKGwwcmIjRPIGZZcZj2Ow59dWOS/4WYFCCNls3lzgp
L3ioYEoWkDeciwVB8LXgRbIIg1UkFiAfsQUcGfN8Nic0riG+WHxLZUrncz/j8J9XFYsF/w++5RID
dUzpnIjOcUKUEPdYtGcw4108kclaHTRvete7hEHONLZVmIiveCYefaRcCPM1oVfyxs2D/ZItcjN+
xoN/u0wq/zxvgs1yUeRy0Ps4Zo/uCbyv8QdDSwyhZoWwKh3Hfprg8M0PpLHjVQVgLwBi/v9QhkHd
vbWcJN7uWPFnIy3PPJ9EtOf3MZaEx6fIRF9tF0wGSAcXAAE0g+dcDNOce2kzdRnHDK7Rv5JNY8kh
esBzZM1j2sg6AfRXyM1OqnL5KhOXmnvdNp2/GRDEWcgqn65esXvSbY3Pt5JHbc5DgJiT3/FoFEH7
4S3XuLmh7u5m1vh9QJsjgJdpd5PKb/EG6Ko4z6iXbd0a7Gloc0JOdlNb2fhF87AYM4sN9MrCl0j7
Wt2CDmZSPeoEjnY41JAQL9qecwYmhUgbn9R+CjU9nQu2aL60j8soJBu8zFWnkFYycS3hvbl7spHX
GsihG8QGOkl8yQa4mgONpEXEzqcVJVDCc05q0xW0Tefbl/ek9NcFrmuSc1ecfF3qrMOBx24kz3eV
6ycC4w8DIARGMTclJkj1wMe7bJqh9yMl36Y2hyZEwpVQrmn7Fs1Po1JgM2YqCVC+FhpE7NzVrLQN
O14yDbiSGCtZb9rUPdgZShIbMjh+lF82waXqRYQbql68kS721HmZ31hejPX1welnokYAoH6BIcre
hRQTUgB8QJhrf5TMafqdSNiBd3PNS2QF9H6Y5dTrLCUiAIFyWtNsZBkKqdX1yBDg4FBvuaqwDPee
veiH46wxiVtIE5QvF/4BCs4N/vy2d0CSkqt8gzukfvF9YbxY7IikTm+Z2/Xr9G0ehWsW8dVZ+dxd
SraP/1fItRw+1Vf9msDD4BmY9NV5JV/F38AnKzg2M7JkX1DRAou9VlH9W5tfFXKfcVNLHOoFcaU8
9u5hrcSQZuyiI2/WScx/tK3hY7KOuNtn8z1Batzh93/tMZqq5tvpHmsXlBr7htS+bys1Dzz3osQp
9geCR5IUgcC61XgOU7NhU8ZuyC4Qf6GANB+17IHTj7fxVMD55WkV3sFATK96x/GJoL3CV0NuxNTe
HzXX8QXxSEIdwNCyOYAbOCkUt19HIcsRkJK+bhBVgeiuLpOQuveFsxWkbHrlsw/Go67uK9SqWpTj
0rWR6adD4qTMWxw3ZXsrsvCchpr3mxy73DsICLlVN3SCMxzV7Q2L+iYiNFtFxJDHTuy9VZJc/ji5
6b+w5i3caooGsMSJ+lCxQoa4gmqHD4cQJi5drvowrKAD55S7C49UX+1Pfih/Z8LxtTObh+TpNT8i
plNKWLf3BAF8asluubZlz6taVye01lqixWfN6R6SjDa5ez9rNdM8G3iRssc600kpR9e6kGTsQ1U1
dFpXteS4Ccxp7BWlPBhBYx/gd0uxNWQlA5uwDhhLxCNoqTGycXSByKocLMtuITvIbN/G/Yrknd61
Yr6iURkIDhC0GXlvKEQ7imkGUtGgm5d+i67U8zQhFWcPv1EYp3NaV3PkOJEqQRFAYbqeVIxoRzU2
JaasyhI1/t7su86x02OMPUORV45T92+WBt0ukFAzezUOfCw+5NhWnJeTin8Bb9LXyH4GZFeQMPsD
EpeLsqozuSODjY1BYxqsO/L/Ovx8UpKAISwk9BeAUJSWpKlfPAghoJVFAZiaWflCM+uJSLlISy95
zvCPIEw86lZol/ubKrkqplBctUArungcZkEZYPjCEm1QAXwr42rEpstCyCJZyPmst9fWXg8ROuQj
2xFpE+59xLTLRtxHlyH4DDyoUOfS9Nvf6qjwH0rCzHjjvsiXlkmteDVDlKDSxVnMnpj0qkTsxuwu
91W5sx9+6m4li8AHSUBB/dV4tySZWX8UQ4HmQDCojUOmO6IzOmaG+Cpm6WUJVHSCxw8YNXL+/m5Y
b9ldVAeTX8308JT5J5mHID+evp0dT2JYxLw8ekgbeGwd1+RRAg/cV+VRv4Y1QL66kJ79NhlaDXk3
Y4oZ7jv5pvfW4eoO4+xVSeXCBcfPHSmjdVRU7GVjfQ+oUx797pvsEMioPdbR/uQkWCk8+AednRBP
Orlt4FQtsEYAQSBqC7pzrmxicWnT42VJgeJ0YuukhNynooI60aDWGzUInP/NbbyrzCyXbXJk/JyG
tMwlb2rXoYdXRbSzbCK2eORRf1zOmoxbZRRWMNHLytQ6Y3gnLHpajsV8u1+3mVnLxh4dBAwHrwkI
o9X2Jdx/wA8CPZwybOxIQZ1t2gpvqN5OsbazB8yB07fxnLcag8vNfNWfS5QRl1uP9eVsvoW2gWON
N7bykCRfn8AgD4TTtd2O8F3yW0Pg9Xi5mLcy5mqf8ceptO/k3cynrj3DmPa3YGOUJfRFtMrnU+WR
+W+S5wGYXzs1eoJm+MGL2LhPpzE0A6KxdscFDSQpjdFPQq13jHZGeQ/iANIgjm4y6g91iWWin0Yg
eYDHevzVm5uyAouy4jevWdChSDq8YrpZxw+s8BCFZEq6evbEi1/akTmXv0lSAok+cbdbzeQr0dnD
/Y5Mb4n/Q27fXRiMlcy5q8Auv69A7GK974gJLbtVaS99cVsc2qeGWLda32Lbu9V4X1g5ZZ0tEdm4
J0BHqxqCp38qa+yxbwK6/Q6UqnLw5ya9hE1ux2xxgo3iFyze3ZptLoEzlvqxhXA6rtrbRbk5S4zK
9LvWlx8CIfl/CgjBNUD8CveD/W/ZQX1NlC1gHyaReiIIVjYpN3A8JB1pWdAKZ0neKWvcwegrOASe
a5/mbkF2M3aIcC69xuCDDLMKFICJPd99twM8VhVm5f9ASS087j6X181GYIatwUHpREJeFIJiDifU
dgnD3B3jGEQBcrcr3GuXJoIlu2TrqYwExPrHXqn5oi6ZtbD4VZaNLsw9UZY+QLWoU/XNGQuoJ/Cb
Rk97cfweLyILCudCgEGFS7HAJ1TThinLYG8CACrTlBzszVkN9cJPZjkXrTEpTrs4xwhG3ku6JQDo
oMezi7fCCbvzhCGL9nosY9kv9Lsz+cMeGq8Dk22qv1Hby5BfLV+eSeiNhYUPrDoCk89pHd5Yp7BP
eCfltKCftGDIxvQD6bjswRmg6o1wK6/amBPCXIJ/zIZSeUDmMd8A85EnNmg8B/bMmU5T8rzujv5e
hITF9nEG/PKqaGQxCTwguQCau2AORFlXxCcKlq/Sf6TRokqbUgHDbeXgh13bcDzK0cYdUT0HNSQs
B/m8V97CJPsbeXsDdOaCiNgjeetxmpWOFzXdtxUhfITvJlcjjo495dxc6E4CrRKj7j1b0pyJLupM
Xcxj92ePRdWe50mvGYkG/AlVZJ8iUEJzWvSngcV467Cya/mkP8153MQnEnJ5BUzD7igMEE1hpDBl
2Ibti1MymCeRjQLb2Ixlem1ubr7Xa+tPrthvXVKY4xI70grMNUX0jw4f+JvImnUQU2SSwBLXcYIx
So6ARV48eDKrRzuUBU9onyn/INYsoYsWb7a3wo5AZflUgYGr/DokKTZbfcmPIryTPnuF8iAvw0FY
uIMZBU5OGiwUDJ09qY8lPTeMNbD8df12pW+J4I90L97cwJy9F/eWpgvGJezLtbC39q3SYR3MrLBS
Y1T8RZ/ZPp8r2ie6CL5qLb1SJLmy+MElfZzuMv0sWLXSj8YmZ8s5KZHXH2bEMqhtDYCvPcUazRA1
SxPGbk0vc2tPzN0vrAXmuUKgWAftM3QlPyZDNHajL68zNIWvpKA2UmuI3MgfMUAkbxbKfm0Hwftk
W+3dI4eYsli1GDy+8c7twia13dErU3ZHv9nEi4YHfnrCnc9p/beY4vO2qCDib5CvOU8APAgdRkfa
gV0vEOonoJdk4Qg0dF53Dmo3I0qeaXMAR8FKBHQ2KcO1PRl8bpBC2DL/y+d28f+WjO/qVhKFDRL5
OIf5aO20Vm15lEwHdSyvM2jtUbamGZJ2maGaSGS9hdD1lrRNwl/Mn7YL5xREDrOSTSLuBvCSQvCd
4rcypdpncyvjljrc36paaTm6AxenRAB2OuqRNnw7qfMONmf5L7othLKjMz+WXuws1osPsEP6HNtT
Isnau8X00BobSvlh5AWkTkS0RTTK7pxT0bSQkwni0/qcIZ9JRUh8dqIC3Oybp2D7bCSkmHb5YxWR
UiAHRBJPxDe+0CGa2zfVsyS3snEh6iG6NG/146AqLfg0WQYCxUJa/Hblmvqpp7WWo/G4Fa/rDjzU
d2/9dkwO2O1fC6aJlIe6NVfd6Snk34NW7GBquMToMe8AtRKTXCwjyFY499M2aAjp6SxxLRQRnkIv
EQIR9X2nryjrqOWc9yzvFBJsC9CcSca6zr3OfMCQwRMD+cEgm5OfPJldsJKH3Q3HfTOu0hMfD95N
lvRKyJVfgj234oPVdoJ0hUlx3CuLBOiLceHifKfzHL24Znnp+SRdDGe3qA47fXhLL6q+6RueH1P+
jC5vlrcNE1EhXeKJT39d+a+I7gxei3eEDgmkgdZ0lbwdJiCOZKqJXp7dJXvZs5yHhirOHl+/phl5
GkwzabzeSPNj3qpFsKdQuiFf/b32F+NZ9cu672V7fXSXDDohjPouQxQsYOsv2HWwTrQuDlsWm0pO
qMOQ2CJnYSYG8Z3ahgVfmKGgD9imJUCAmEpqMEWTVZWW5X/yXE/3eoGTJKj5gGBoZHEepKfjTqTn
PsyJZTUL4RaFqHAT1umswoBhWKZhxi7kYeBla4zMq7qbWHV9sLz8D47PXzU/CvIKowDSTQ9Izlg9
Chj/v6zKmw10eAEdCv13VnR61/hKKb9/GK1w22gI7coODgdvm2JQxcUE/aL4WuIobfT13hBQlMAV
3YOPnZp46qV/OIFoYnbmGBgZfSMkSq1UtBKsQl+HvQLbYS3iFLYedwibVeaNvITJ7gv9qmV6gqAy
/yUQE0yDjPsAMdDreA8DmJ2w62VFXl1sk8x3QBBd6B3CmdJbnAvZDZ+rjlTugjZ4iD4n9vYhwlw3
v5Q7tJQXgcZJ0qvvQXtPBPRmjhevq1I22A/dyx+mcVEn/Q2okU6/SShYUiUF9qyG4RLtFS2835Y9
qsW3czBM8BpIUThcqYiVGGOLYGdFrmOa3F172LJC2JtFyx4el4oNsct7g5f+JFBjJJ9aAEhsqJZa
Xfds3/r2S9TDr56FLGGGZmqC49/m8wabp0Cr+xivEXMZ9Mw9xj7IrNRomZBOOonLZB5N8URSzirL
+jSnMvombUYIE9E6PwW7BseAaoF43H8E10entvuGpa1dHKz4XBJ8omYqPtFFWXc/o36cAidFsG/Y
Ryar7g2iqKJlg/3J+/o+aBB6kJqip9L2k5n718yq1pNCV7+dX89nw0E8NGqdIdf2XdjwR6SHpOx1
S87mgChvuTudhmUxftf8aZRUoncRbPjncccOsCKR+Z4CM24Jpiv7XQroAxwix2qwC02MkarLU1hr
DXvwj/jUHCsOUIQx68IBAR8+Vi2OO8RKoyLD2eK3+wzVwWY773EgsxswWnqD93Cps/BOqbddVXPN
HoJAjTe8rKRMKFN8hnX1FAdBW77Wo7H6KalBn5Asvly+RbRWnR7I/impEdAUidzwoJwjzBkPyXti
efbTCz+uvAfmrZVgiYNb1huyLQ1dAsmV84MDfP34RVbNPE5rjY7yN5e0mZ3Nj+1B53ZvA0lgbi1M
3DYuMP/O4DmAviO+zDSjaqmRZ7zOcAUTy1v4LUJ+N336Zmse+Qzky/kBbTt+ZxDf2VIsBPvCuBUM
HOGY3T7+VKocJS6THwM3j3x0HSJXmclpkmVcOZN+x+cHNxaIB7TkCkwIEFN7vJ7JVN7jPUIy+qgk
xBAuEmOUM0B0PVV/VixjbCv3tOV8qDxCXOg1FdRG7Q7Wwu2t3hd7yiJqc7g3CdzAcDgt7/xBUBmL
dyIolfX9jGE9f6l0NdQ8a5UzGJR0tFwVsDXMaM4tcxPUGOeL8hU+Ug6INeIui+58zQBDc8fM1Ik6
JA0GS+sYDoRw+z/RXhFpsHfN7Bm90pO/8b5ZSmCST3hai1RVp0haVMXUgVZOHrSCOJCKWTMWZvJ1
OYmRCXMsBzQg/2rfX9HUN/zaYyd0V21zLvMk5izX5Jx9O8v0imyz8PNsIIzp7/ULIvDiZ5O876ap
2gJzyeJaeewsnO20OkhD+v37f+RUCtyxI7bkkdsWECeP4r1b4gSmdTzzxmDLkLmVGFuP0X67ArqR
0xqZGAD0qaD9MWeij6UGVRSVFwifwVGs9l5/mJDQDuUzid0CjmPGGnz07Exd9ghmwXGeSqvwPCZ2
XJJ3Y+PA3qZi6noaAnZpQxdwgmIjVSECrqgJPk0CwCxzuXX3AsbLw7GfEJYuSBKgb7NIpjDXpmZe
jbP151loVNPCMVNk66nmSoqXBnuIQW1nfpSa05xebFr+SBvt4HgPfyEZqDJKtEjO/Y3jjBTDO+dB
5dF4Cd0GwvsX+XPULVU7a1z8ZFWySoLP+QJVMqsgXJSp9v9Dzv5IfG/n23sAbUfHke1LZCsEBdox
rDFsubwFtlrbjsQ8jthVDquXTvhi4Oq2JtyYoExiNJ6WmgZcZVWcpvISfei1cdeBm97ksoPRoMAF
+OLIJ4Imk0CdUgcoPhsyBUN7tmLUUN23oknKPJ3Foec+T/HRXppk02uAVpyrMYHKe1xrxUZMYH1I
RlFj9qWXK58pnQqwO752dtLzJlHwObrlvxiVG7ds68NgmLBTnkQWiNyr+DJNRS3MDTEH3vvs/N30
rbfJZcyDvGV80nk3stGHqaCqvny+GTSoS3pF1Ed7GHJKs2EKX99SFU1Vxpl3Yi+VTDCN2bwL7/Xn
+2lOeVE/3qQKRGcPzWFuHG+Unq/xX37r0mdoT1YkOaIO97BzBcn1UWMi4hnfyx1IpbzwVYiDMMzA
npo7kVk+sASkKm8tArRIeFecJI06AEiypFIQoqqvDOA/s024d+Cnzkb1sKwy4eUR1Cszds/USXed
QfzEmYtIqkvUENQjUqNPFwisHhENcJPfJN7Fv+NhXdXKbpYRUilEpEUM+B+y9i2V4QOlUsCkgDlF
71ui6r0hrGw5bnx5W4AL46W2e2qCXM1aseujCmNJ1zaWBalkSG7zf+/U8hMk2z9hVDfylRoL9kef
QoHZew+t/HvF0C4kcUXRIbwURYJQ3N5MTIeDsyMuJyYVeQ4PZuPUN4hbHJ4AqhuR40QACdpQyo8F
H9JPuWW4YS+BIaVk0/dU80mD/pATO+alnGiRGHptpYnvXgqmeU/jqBfunqzGSc3AxMCHaFk/3vmA
c7tUpgcJdsTlMhJMxSLEtyAfijOsWuOkU827nGNY83oLAtWWyKD4JwcC2eGX6z1ViZIyplCXfvYh
H6dialjYlWuWFtzeSaRS4rAL+kV3pq8uvRg+Q/Z/NlapulmeU1nCqNlukHkyYJN6ugm8dFF7PPeP
fHyVzBdvzrXQyPPuloEK0YiV/FD20y868F7BBIU6uTdAXroi8ZlnCAWffz4XTUwP88TBjlau8VZI
Ra9OSx0Z1EziaeQT0/gEQs3IOO//hRQExj3IdyHuKY6WS8Kbb8ut17bit0AEuIfeh/mwp1gY/hDL
EOgM1AmPN6BnrHup8TOnCJgrnBNWOMHdeKNDgPMLa3fBtUu7XW+ow8rYqaxbXYUTPzRIi8Hx3JCp
dRBQERVkr7dtiWYaBQmAdpk4wEhC6HmfDjIHGne25Bhk1rX2DIoUud0hP3udTJiEubSUQ2nm0WDH
pLNrQuqQJjf+CIORFbNUFt6PVhNh7jUVzUdaxc5uinVuorBlfSeG1od79BiC7Pm9J//2dAkwqpCn
EMAO27sKtGw6zn286Al7bAMXD6IIkpMY5qH7YC5YIIEaFyTxTcoGCyEI5t9o1xwNcAmkiHFmpWwW
IcAW4SNkiZ+Arowlt0o4t4qjylGNAE5+tXrwSOlHI1zzeaFdOKqOZfKcTar/p7AY87jeXHiMbJ80
LQNfQU8oYzrQ8iyNcqpV6LOuoaGZMuD/CYtqvaoJNIBmARlRgyyXyfKOa1MoOtk8/zjS+2+T7qKC
OnJu8OqQKNmpRs5GcFkc+Ho2QOIvFY046yVrUhH0OjqxiQf821dcP6hn2M6HbMSFpqA15xVT139U
+aT1moWV9RnxtU1MYcPAZkDEYw4s6EN6euW0EC5lY4vsD89AKtUFGo2xxRTMSO/9W835Gcp7ODzL
SG1wdZog9RM6qoL03SKowzpGqyNoDRP1raNHT2YjWUa9RzzfpUU8p1t98kb0JWRjxxKI6qNlqs5N
fi353niJhfhBiLb+TF38CyUaipV6T2ucavcz8jRp+yd07LBkMNKK6Sfr0dAdbW3wl4s0lKKnVYk2
cxKimtqk5nnwm+QcQkgESeu7SBuJSpzSlZKkzMZF+3W2EL4/n3NfmHwXJNxfLu2vVGUMuHHSS2sV
+N9zVJ1KkmaNKji/ZgfEloxxCkugj57+9/h+RunPokzCOF2pZ4tK1HMFdihz7NT0eYboEEryuBoF
5e95PkG3qkIWE6/G2OyiPCx1rpYaK0G8730o7ON9u10F9H/Y10sMuDyhHNRm20SbxwyV6mp3Zcpy
6LLX7U8bOFy3PQprmB10r3oVfOp9jAgnnxpi2NjSKOU08uRh50DuPc0aAefbymJZsWEdlqDah8KS
yIRwrL9MTV+z7eF18PDh7aPJzQ269Crd4tiXQAm03utRlnEyY9B869js1i1x8MgEFAAFv8LyQj1c
z3Oy8xcXc7VnPcJNwjoAmG6JW2di4CPZdWHSq3Kc/MvIE20zL8DiLx00afpB+5y45TF0omV8o12R
gLHsM0CVtgKlDh4X+tIzQe9YLyFvrpohFDiu+Q6nwt0I5M9vsjMlIGIbfeUKpDENdUvAtlO4kUty
ts9aSQlfjex5xr/noYBQKFJmpMxBFN2DtL8hQajLWWyzGX4YoPEhmlK/IYfevysttqDs2/PdyOEF
YHtAmlEaPRtB0aqA609ZOdJ+W+9DJ3NMgCfmrOMazjM+2f8aS0Llv/s2mLBJBDR4+tAVEolTTXS7
Jb99Z+VplCVYQXPFOyVFSm/DwhcJ2QdazogRzZpAvA0D/xcKNut4ZARZSL4yZibia8SyOL4YENYs
9JdaSBmUcLhEeDwnS6iUBfIES5uJaKbwG0v+Fu3qy36XbIXgAe3XKs/7LhGlY4VAMyyLvZTZM4tt
RxxCrjx+GVwkO6adFx9jExjp1K5BSg5/m7oNklrhmWep+sX8gO4Ol7HHiAhKy9whaaWhvpncdK+i
eKnFX5MH4WptVn5zAmSPQdfROEf64T6K8kim0BtMVitbWJfnDTjDJhANjc4BrOSHuv2JiKL8g7gT
xcSuKnz7MOoSGtJV4RnXtTKEpWeeeEj6y6kl8t5lW+TGaOK+mceI4frftiqKMgNIA9/w8MXjwldX
36U6dh8g0wkamv2pAMgkjmyK9zF6PUg2al/O+7JyBGasQJyhEGYK+fgmfV4aqCKicF2XVecpTRUG
Jt3KW2FOwYmncmNAsMXs5lDj2nx5+VHDHq0sW0lADHZQn6gApZqrr6/pPWOW+cykCJ6Q2ilum52X
X5mjh1OPSeyLsGxzsEAVcGBswHeTV/48fc8XqIjFkg5UDOsUu7MzremytMWMQasHkw9Gb4BHYqxR
dwYjYytot++lj/0AjlINTXb8G6Ci7YcS/4qn2ht8FDFHf2S/xtTf7GwB+VN7tNV0/jJXe/qwGWCE
2fadpzrBAnsxfbDsJZR6EgmJNnjbWU5hYKOptJNeIAokcA2crZr712tOrFAfPbQ4218sAalRkJH2
MT+yRy4zo8BRYOppieugzNBFHfBEn5mHW8736vQQ/mEIefDyyPtykTwtnTBckBWZVjI2m9dcVK5O
8WWfGEaMnuVl99tK756RSRN6tbDSMKahE8CLEowKqi4r8Z3qmlwfuCb4eAYaDfHEK8WDZ3a1ACLu
BAVoZ8mXXcXXT+jc1CpUWLBayHzGmAp0JpQnQ/5Ye/+HiinU90A1B2Ot1YudDYKtCRaLB6B+QFQQ
XXtkKGylVTfGLI8HE6yROxP8kXt/AlXzhxQ6W2IUYROo6KY5bPRZBjO0a7TYjIuNwLubKKutYEjY
nDOSETKKNp2R7VeZ/58fPIDku+C+X1u4YDHHHAu3HTlsTQhXm9ZCvy7nTtnLb9AEYYLcBDFEtGeH
dT0un3WoUjjOXPJtHz+p3E9+BEVvG8UD7twPI6HoOnVwVI32O9YXKc+HghQMgMX75FfxACLrUFg2
+ihXsKfQUrJD1nHtmDM1bWTYDqwSsFpk2KzjkNEKeduVAbB3tbQvN4iXWojZwpu3qqRM0vd2a1CO
Au1ElPrzwigzpcHSGZ8KCbwozNxjlWHNhGhbdLdZV7kzKaCLNpA4IbRzXl7m4adaDj7B3XnvPaEv
Iruq+hFxAGtQ3PDwLngUy4d1naaantm8moX7lMnv9bs6oTvrqxZRVQIBuczKp/S59WIfVh+/S29R
6PmIyZNVfE1lhRxYALua8HM1HUyPege9mHVomL+hvCZrQrN9Ecwg88h5YA/RVZeNtPizRsU+0uFQ
Bl3zEuMN7OetS1Kxxxxoa2aVQJ1n8jZ3Pl8kt9LJVHYJBPlBV6RC9AW4aLcNSaFpPLyrPGfJQCsC
amfExLD9P+EM3voYigOonEVguxzC81LBC8SNUh+mv2q8EuewSiJDdQbACoAz8sCceqvRrrOyPYu7
6kFYnLbXtEkR1hONH699Bof24O46QEUHtMPb20BIDi5tx5+9jtx/23XFVJq1NmZ9cf5L+Q1cq4tv
3iqiRAi2Fvark9hHvmkSBFekZSzrCgLYHPRSXN++T5p0OTxu7j7NTeQn/B98XoIG/NBd5pLTLeEo
pPbsaFf0laHqBDD7KGZ/ETod1IBArhnVA7ilVwJxB/w1EmNdnKKuNiKryuaZalL/4UT91KFAQ2N9
dGIsxE4XUST+n4aA3k1aoM6RB0f3lWLBglAL5hqclMRwNrw5Bteugw9hrBFCK5X+MkJWtT1YYYyy
0hYaDnskh2TMKOZ67oAPdhaNqhqTOhvtMtS9ge6FOvC6+F8fBgs20tj9A1sOas5rj4jEs2b+DshR
wYj3tt2OviWV5PeOUTwdi5Xt/o4oBZ0HyXGiepY35jCKQMTLYNoud/rI1BO+KX2PGr3F1kty/eRO
NAFGt5THQFz4ZscgBxHfOrYAPS5lz0q3LBOMRUGeFROZJvuAMcb/ZD/ORYu3Ho7dFgV2BMXViB06
qtTPBG4Zb6X7bo+0dufHtZH54gITQy4TWr6L5A8sLtomrfBnRd5VF3rROlLwORPQOYN4mkmG5Yyg
PvLV49h1bsUKlFiriXtvqva1REkjnRQJR2FzD7P0c+O5cjsRS4vWAN+yG1DENVFso3LPGzjYB/kv
j33U/7N0ZUqoXvfyLr7hZPgoElLz4g7bB6P7mATjvE71VhCpFNaEuYJ8PzFMqqtLUebOJTphadmR
pCWaEgMBgJskTAR+cWdH3Pq9qJ1lyusxl1XI6r9R4Af3fR4aK8xh1nSXTpByjdIgmuhjp9O0F6PZ
oLnLMdZKlvGefWq7yXCNp/NL3a24sLlgRAJhA/RApWP1TBqOK1Iln4lnzWhK3g02VAwNWf6uMNyC
T81HluCy4Du7o/O81JXYJ6gNJ5KtwnZOhDVsCgrxcpxIcn8Dp1/M4ze8DAuzc5pCRI8uC1/2UWnP
4LiPPAkpl14HlFWQ7TlJQvz1MxrIGCzkiImWQaoLzQ4e5luP7tgfhUkMSz/uRATJn6UATnNN7dGs
3TEZz/bRDx/bH2Yo3Z4Fj99t82AQWp52jEbUOjKGdJOCFFwDI5EhKov5/ySFLJ6O2Yh2E7fSmhNp
B77vwnDt132dJspQ1MFe7RkgCXurKFo3gWOK8+qAEcLlxxQyZCyfEn2fhCQtUA1Ef8h5/Dtxsdp+
2Qymxjd6rA9CJahQHhyBtBZvFY3aludApgUGgdpdJ1svt+n8Z69VCAkx4KdajheyOoI6KGkZ/2rT
BXJ2clWQ9E3x/vjmagrtQyya4n8abvEz76+et/VvwGSiLB3NhEdl6j3xRbrBqtpLMnl1ApS/Lu9n
4rhRtk/SKaOa+3AcS+fBN2FN2V7L7gVRCcdu1bOKxx3WCaFvg7yBA9UFp/YRwxFpMq9aeG9kBhvg
GGUFpw9WPFK4Y0Kiz/mnLKuANkn5tc7tk4KGVVGpvYahXKxyy7VGy4pE/AUF+hZLG5ICEj7SYjgU
aGb3Eh50FoamcWrEXQiOz8PsgBUxlPkbo0GGOE45aLNsTY+MR0HJVdBslOoYJzfwzlB5eKLt8flp
wkmmi1dmD0g1/5cwAuNRryWXrPRLVOichuh5/x8O6eLTgwheIA6QqbzUbVM+noEHBI2HKfs4KYTo
Vi7lg2gz188/jQQbSwLE/t29oyykoSCV2n7tjnPnSW1k6zO60LK47e2kuxHlH0rU2MPt2VhHLb7m
NmTFvvRnNKDZDoK6dD6qoJ6JHnqzRt3/hv8K7E81sYkCJbdOdxnHu//VXZaPdtXyS6Z2QxFPFzjs
EuLrZNF6chBVRj1KLXG4SNCVcwZK4IDeDxGdKPohJf7NTvc+90zsf7rtAVSPotDm6SLNmb+hxFmk
2ZBRYUzj03F/SJ2enYC1lOpAOWICJ6RAqYTbI7SHfOGcJnT1lq1Auq/SAlxPrIQ5Dh8ADvH5Zx1T
W/EtnghDgBp4WS00vXjLuSTm2KPaxIM5ySvO+5Iz6OWKGQM1fyzX8oAkA6Dvl/qxXSpETouqvzQl
NEOnp8MjquG9yvCS/NVGQZjDqlB+HLODZcHcjvrrOU9Ndl3LNqZBmRpAb9QF3TZq5golsWuaNN1C
dVIdzlUtPWajnm6nzhL1ePM+z4tstM4+6d8V+6PNj0NTtGj5OeAKy/7KBVci+6lzx+CMgh2/m46H
R/Fi8/pph4pyv73qPUx8FQ6lzKQTete16OsZw6Tz39lJmoAKQhEKcL33gto6Eco4mZ0qxRjZMaZE
LU4B5F2E3WWPvEKDYWEmLSivh2pJZ1d3qC59JvAqmLYxh0Y953gNiDWsw9Cgm4sxMWIET2jd3qvX
ee8UPrS9b5fI/XTeUdH1I3x8a2ycVxBUxJenM01b+ayTZbCO7eoW1S2C9m/igZs6tPnw2Pbn6Nb7
MRC91bBBVaaw1RlTzuZTkXlpVrBvi2vziiIjCq3m6R3puZXu2+7s6EjqAUS5QY6Udc3XtsdgU4wp
fv1DFkDbR8snYmJGJZq/RFrKEHRVDeBcorPJqms0damKBedMEyHmZ40v1kAdAqqsyQk6huRWdGDm
EKjifcpoC6v3TDzMzgc20Yk9cEbKu1hnSX8Fb4XBl0WXzYPld4sZVgcWjE15l9ZHwwrpG11ETPeT
97f5IQt4O+E6W6VCeypX5a0CsDJjKlCPyHCIPoY6J0QdQx37qoAXs9zHDbyoaNTnL3Bg5uaJccJU
0SfwUVyNqfdQfKkHi9Ue9F3haPanj+tmdzjGvOXuUIu6O1D8haDEdEX7Z+2icRdQqT1YWIXkVbfU
vEvXshqpprpjcBk3jJNmRdAmYAkwazzQyD7y27LwODnVuV/vfHnwesODfMtDr2vYn5dGX5JyVfM3
PFOtAVxGu9c06rr05K+nVFuZ/Mex8a9nmVmqU2NQKBgsbuH3fIh9ZEdDbXWqKFX1dumjNIP9n+CV
QQDR2KkX/ELQ++kDXOsYFxUvPMbrJ+UKg4WuZcX1nzYLQh9Vn+bdFYfmoST7m9yvP00msRFjU3n5
dqRtlPhKjexy8rWGwb9Mvp1CCk5vZXSGX7caPouOOfMlFySuehrIywAC+p3yvtPlSnC1I0+0Vr4I
ARwQUw3t6pxrWl/utcfSVuj9GkL3tKwNG5Bn4N+1X7PGLCQNG1yukFal4dv+CYN6+0JjojBQzSk1
AeEOrVBE3BA0TH0EYqj1/OqYUgMw/o8BBxfyPMrKbT+sQyswH0a672liMtuFSVf8+RirbvQCGoQ0
QuMbCrnxDvjjcpAiYuamIwtDnUx47WP/ai0JoW1oQxmCYYgYjQOcP3/AbN85GhC623fU0GNgmnZJ
QP9QDYhvaozugUrlKcWzfbxbA7eOoJUPGWvlWjzk1fgwtaDPBdbzEvb8RKrHm/7VLmJiQMPYxN/J
7L1w6gKlksPDmIsGy8Jeqa0dIQk/EhSjrQAt8zglY0YGx8ZnRw77G6cKIjxXFjKw2Ib38F4NTRJd
qYyUTB9hx3hQgItErzjERUjpgVrMNQehY5i45KMxU+qmQsJBX0fWHKT3756CQ1sEiOTKBijEuVoy
NvRxnRvopVZLxCBXbv8BZhpaccvnvgNbgrwJC1O+ueDWpJYwOxEBKI9EpoxGDPLnZBAiRBiOQB+b
xivL2k/2mRdrL7qP5p/3j/AZ7QveM7YAG6K8PCzHxeNMWi7nk80L4Nb2szzlIFIfyVW7Cx7Kj2pe
LzJLnDZe6tyofle/OYGg4CoeaVciaHHxk3fmyg2JMy+/wguraG8OscF5RItOLPMy1++6WVWprzSk
7KNTXR5p1k6vDJnk3CgfJS8dUqiePwkYf4d1H8I2zkbZTzvL+mxxAgIyRXy+7LKDdzZwL4fQYrMl
q01yACZkBlXQ96e2IINtdjAeAGpGEMSZ09EoAeJy0r0tV45+ctBxAHXO326zpo243ZKM1xsz3gZ0
jMfVZAr7eWndKTrfQHdIWgCkGUb9WppoiQquVGCWjl3kAPU4LBqgGSV/uoIxU3RCxna6lc/bl6sS
CjYDwz0f7U+N0kS4+CuzB+qVO9B1S7dkkt7I0Mxai7TP40wgsJaBo4OXQL02SfC2Sl8jRqZ8g5LT
CWOIhPR400AWRh16AEl8Zo6ffrwu0/gkhWPAXjQV1xO4sRCD6MzQ76DskFF+XmRLkWtDrqUgXFRZ
bKsLYggwOguEvRz7w7tPh0E3RPJkhF5RRKNZH8crrfIsOCthF3pJ/kEIRgNuSicPL1Rc0k+9MWvV
lelFZbUz4bbYkKF/Bm3GgziLN0auOalSRxj/ZcMWP5uyc5XSHHdq1fisSmvzMOf7rSkUP+J1IYki
ymN2rHcJcp+X3cA4BzkHadB2Z0ala1R8bRxE89hS3FoFfB395gMZuvU/m64FT9PBR6KZ4Q09lFht
mpZaVtAuM4yYnXWG1atJSU+Hedo9Y219PxbuqBUPdt5khZHqGI+G+ddYu5PtkeSQJHsCKn+R9JWT
B0CM75wb6yGtzmQYMclGcg3Cybuc0Q7xvdgG+rFO6rzfsG51rnTEeD0RuzeXltufalA0/qqJtECo
PzphbUVwNotbNZLjW99naMSijEVUGi/5AcmZtbg1fdDhZUb2mzGPAdF1zQqQ90ErAgtuC2coY6bn
ZdjRJIk9ov0ujDrBMQT3JEUoMU9ByvCzV0YFkkV7fXnWtLBgdgMgB4fJ4c4J9fMBb0WAtUNRIqTU
O7UTm2+DYl6hUQbHHSxVDGkfoh2JEyb2oVsLp/0FBS/OuklQXVX4NKe+aS/s7de/BUpXrGxZqHIK
Q4uMEjAtGPvRYpVs0mhaRhkg4Bz6+D5K2NsY2WGbpo4JQeVt6djhEibRCykPPoQYpOO4+cUHs4l7
TC/HjJwVH4ZE+oKM0w4C311Xzx7fScBciBCUn0rn6PQIIuHcHxjS7o6SRF5WhtQdsON3XmswC3cd
Jx27uhn+PCf9UnMf8RFSyH1sZFRw19AyOQ5zXAjnp9k6CzQJN+sm6nJkNQLnyuR34HIU60FMbtf9
+FtgOCwOvk/ZyH9ZJPzAH20BLQxRXQ0Hm2sSoXW+p+1FDoK/he/4v8PfrUBrdOFHojrf8nUi2S+s
0rgNV7Ql9WvLP88KwUkyDeoTOhFr1OnZaeeZMV15PKZsnK2VC3D3em8KZn/W1bBB0uFi02lnKDSO
Q9OmlAZeqmuDViFa6aD3Wh3F/8MZ4GeI73CdpYqdInZ/uyeiasnUYcUhDYWH6Rj42tEl4kRkyraX
4r4h4gqW2PRQk++YgBDJcXmcSl3qcDpf4fXl9eouZ3e4qCBaLPWSo5XOaow/wjNJ+rGoK3m3ZSeO
ZqWdOM40ObAVXTYfCPTu5KGWbl7f24CdWFOvIH5FDhYb5re31vhfyQjBlXHR8m8lPte//lVZrQtV
0ueZh0CjRMU9UGzPgZGYR/unwnYRLJE8RRDVOtFOCH1SC+rD0rsqJPxCDJv8e6DhhcNrs7UwMBVK
pfAGdzfukUeVXJGnQdssbGUK61PvjsfyhVs0oDgG0bmYHZqGtBjTQklJr2LNwaXjT5TaE1MiEKI9
a0DFVsOpMRDFC2qErvfNR0M4ZsoG4zVAPReMbGB8Wg0k43p29yAXZQ7sYErv2kaPSyXwRrNsg0oG
yCJE/lkzWhHWjaEIJpF09b/M2SkHPO4JmQjgO4c/tPumlCXlAT6ss9/xK5BB9Jyx5qt5PSb5sRu1
q90OpdyWtkfUtkfqC9xBLC9aXKj1bnpx4mK9p+Fw85LnvA6GVLSiKy9Cv+ARnGEsZPbKfpwhWBLQ
Iia1Sf/PM9vgSSNKfxJ0WlUrRjnsNTDiNqeeVxfVtmMueoShu4wcb3pnKNt1GxcxqkACyt3pPYi+
ev4G1n0NKAUkQOx684bB0VrJOaiDl4ftuZff9jgot4SGb6ZQz4jXi4eJez1WLRkIsZtWjK7T6Cy3
AQwe/Rxho9Im8VU9R+8WMEvjxSxrJWclw3SRL9wOQODdj0mmzBH+Zv3m37NsYl3Gw3TF9U+wXViq
iX6/YrCkyNOvgME3rhvdaD3BHZSYtXJMOxWjVGXbl1w7fv/I32G+3OfNHIqf21OMQioPY2fUmlEk
HTf4OtU3IiTpF3ISXEOoJ8Slr5epUu5XEicHfWdaDb21xGXwDITTqQYcMYa+gtY+hZwQrcmj9x51
Doyoe3ijzXyzDXiwXsTSHBM9yA9I8j/3YSYRI7GncyBBqQWrXfaJ9KMba8K2+OG1CcujzfqIS7eT
mdZ5wX5Myn8rwJX+mqS/PlvANPhSetPjqeMf8Ibr/Ns4az7FSNGSYwS8V7gzhUeGcf3FzEKuT/Zt
Iq6Oag9QaghlMhbJrfu9eLRls6jBnY3BZ+f8sTqOAKbX70C4SRSLLK89thGQaPg4+E/kOwa9qGIf
vATO/N+4AuMUzxzo+H0Dj4czpgmQRhYQHsVb9C4KhxKnSJj2ZJ8wVnO1lv5QxTsNQrISfBiKt3qE
Oyb8bTAN7ojTkXxCJGnRfl6Inr1SGxVAo9oZKm+f8IIRkDh+K4KcOlP7B3OK2u55Q6P57AdbLzZz
373PCQwbyslawaMfG4eYlOgLQvPQnHqbtoiT5ejNUYqieQKBAFslCpqNMnZcCzpKnEQiI6mTbkDi
es6KqvPVOzcsCCyuYyPl0dplhH/svLEB6U/O/wBICR/3Az65uvMluiveqICGPHUf6JbZJSDi9Tgw
O1+gWlL3gWSNvFY5PGwMiT1zyFdGISaez2IdtXSIfzszDiY4Zkd1lgNz0VaMDi4I8wzZ7XPKG+LF
+yds8V/SbTsXv93adx0Sg2oVhJZAJwlKwiLuen8mtiUyRV7skHhb92fawDM5HcMO7ie2iNR355HI
CfSSiKtJ5jb0SSE3LwTqQEi1mUlBJ5HsNsUuOCOssn0bJlUW0SbZs/h5rOLGjN4CRvtbC4rfuShv
nRSYePC7+0npwXq/LVZStjZwxHjHESkzYS+Btrt8mVcN6C/wmOPtTDXYBEJy4lVpfigtvinGdUVe
raaNI+CXO6iQ08QDQz8NdyHN6Jwy1UdolQIjzgq0G1KwjmpjGdL3h4SvNPrlQj4JAO4ggiBHpSKF
eaRdqA7f3OPL12d/8gtS1j6biHxOIUuehyF5b0KwN0BiXVkH7b7CodOJoE8Jrbp0Oj0NPDbMLvQO
nkBmVg4xwBJk4BucdNh5OEZXYbQST6SoEKrNYssPwaZbaAExFBXcfnld0a2PQzHQzZ3RC2I4joIn
uLB/DHlLNJqyOF/x0etThPGP4QLOCbZYirAD8X0UOF4Frrx2pRzp7RVpOrmwqovv9uiXbbTl9F/B
hdxNyj70Fs6lsYg4QJVjRjVhAMZ7kjNFxVZPApIP+x0faa7G9np9nWS/OsaVLwuh2lLiX8b6oAVs
jc2kgYQZCCtLXCJ6miELLwM5aGeCJSjwHBzHVRvGFT6O2PRTaPXm+RjUEJvnakz+p+tEyi05tjDG
C74+FciTQgKn9TPeUxlrTv29CzA/WKCSlMXC1hpK+MSHB7iVvavATbcLSdT5+HSt9BBEbgsaLNCd
4EZLotjOFaq1o51jeWxROFlyToPoV+lRkLZyHtDZ8uAK7w/xwCW65nF4wi6XA+eLZWqFTFjH2ykv
DrkL1GW3x05z/hUkVGVoBMvmcVuMazGNp9j3/6TEdnGjxwFaDLh/oQUPN/gI7SC0PGoWx8jVnnxd
vf6mETWtPy9pTF61ZaNlSq4DytxBtQPfr9Rn/RCFGDEM9IqmlbVpMya0VT3BLSZ5iYd7ZKq3x1Lk
OldI3MOr3jfd0gOdkB+MHZdEIAvVnZJg3tQNC+O2HqbnIlFd8KFgi0uQAoOvlOvJIxUMc8F9Cfkd
w2iRIpeB/TjNg8qblpR5GaG9bchMnh7cWhNal75fWDeBd4yMEwuGScjvE2MGAJoHCjECvHzZ/JS/
ACZW2+9gHVybGBxJnZqpiQ0PD5zMslE/bsQEVEbfI/oXdSbQyb7TY9FW/2PKSWSLVlpaKUKAYhg5
avd92ACq8dCktYcTCJstrF9PnMQ9SsRNmL017tUI0Qte1OiO7X/hL5Wp4iPH0N+S6HFH9DZe5ESE
WZtZ6IXC5ry+FwZ9jodnU6SdEKf7KKZUhaTvfiowNH/X71qehGZt43l8zRFe9nembdsKRqme3yMN
Xw61Q9y5UM/aTSt7/INNdgKwKMrL4ailurIzCuNH16nu1dMgIixTDJp1+3S7hNOW9SynssC4iH5Y
R8Kz5HISm45KYq2+58CSzgLl54kOlp1+0ReYZCSF5hn6xQfBgZ5zrBTCJEKPWMvfJXxTLOWh4QzF
GsFCqY9Y7npVeyn2FbPJ6KEJmFjHT5c38FDCEoupT+TUorHu4HXbSTh7TC1HFBXA50F/YL/sI/No
WPYPX/V8TsRgZwdTN6k0ScR81XM82P3KeOOKiAUbzVW47qxWyDjkN0dQ+xqKmk9ccNq3TK2RcDgs
Zcn/KZRtjCiUaP5VJvdtqRKcpGcfkO3idgiLmcI6k4s/e/6Te1xvbxmPiZQhmU83tDGKelZG150+
JxO0F5XWCfN+J42jGVIh87y4hSgHRLdg9auTJXSDfn/7PPJOAVdIYXzcSvG04Wvwe75LJ88qAA7v
SOHZfAHq0IA7q6eksdOKlNiLMYKTgRaNrQXsv9QwYQLNrsoCx8M4Ades87K3c3fwimPMfuSU7+uh
u+VMKk6qsr3Lf2OQ/H9vYt8h+kiysMWG9aO+TnoYU7HrAgwOIiKHjM5IlNHA0Tpd1QGPkScjEz+6
bpHkzAOxABwVBJ0nvU1oYJQ2XubgNZpRPNiWsWtmawrV9d1lGp5YdHnD63VNy/ocDfmSdvQ56l3i
QJbTqlqsgSRZlxJnoG7cwO94oLeI4ku85ibzOO/OLKmPkdSQh7/kXsO+Xb1pM7X6wWXk7dH30z4U
/44TaSOYGVdz6QD0btUIiVs+bca//OhkPO2rHIX8HlDfY3avj54Q1AiHYeiHPC4yYM74dCXDZiNi
JXWsfvxp4SYQgF64lGkyh+zjR96LMHHGFmoCr50Q0J5NwZfWKvIt4E8MCzeYwgv0ZGtVqmlHLiOw
vFS3pZe8p96yVI0tV+iMYUnt2WZnZN/5FYdfUCm8n0wERMTYKbcu2Ej5B8NTuYguDDjhs8bvKClW
p2zksk5jP9yxILJOY1215MfF241S1bY1MagaA2sQSz6A6a6++rE+ReTmrz3dXqmhZiC9qUnW0EX/
iNR257KmwJFyBUTmu08aG3NYY9V7uge9BkMz0ASdhrbOqtv7qPoYRCcnle98ylSFdDZMRkF736gK
hnWjxDHbur/n1iKr/XYJ4i919d0NQ0ZQUmD6ylAZ+VvRIht18zD01CNNNzlBd+Yr9dKOZvUiTTD8
BbWVqhrN9bhvnSeXHfx8DcrYitCg+54/cUUKrBPkc0SgvmYk0mgy+J8uY980w99kA9RLX2LvCNib
DmohvZtDiPq0vylgnqixo/btkKzSEeGmY0lVyiPy/QVmPECpTiFTdCGpkNG/AQraLzBEL2rf3sAb
tINAA46nh7RXnJYdEaP98HZ/PBDAwOu0GB1hYKVrw2IoLNKSCUxMiwP1DoHAPm+MwFJhGHHbXWA+
xYVGQ+IwKnXzReaDEEHBuEZFz+y7w0Czj1hZYMviQ0ElLdijjgpibJescCd+uEUX+0jTKX61bJmm
SPsLlo4QC0V4AwirdTt4jt9PBSMkZBjzW/4K4UWU1i612VNbbgzmJsJ0DIGkaOVKwCLqXI4K4eD8
xxthMFedOVDlKkrpfTmeMIsZQxbMy+B52rTkOTsqsR28osz647ARgtCOBF7Ss7ig8NFDVjGUxtMo
HNvcPKjcllObRvVB39jK0HobpOLw0WJJwG4t8PT0IZgDake/hzrcITT/qrq2XsxOxf0UOmQgTZAZ
WlxCykY7RRuUcW5JN+fBw4PF1t1+gZLRJqGU+6+9IIyDTPR+RFr+R3Ix8RMkRBh6bKZUVulsXZ5F
gcTKp/oAXTvl79+3Pdw3RcU4V6k/A9WyNO3xdRCa4e71W88e8xyRGxJvBe3nROxqJZia9ZuBdoCz
9pYInyqvrIeTaAZPBEj9gMKgukgVjScHi2X4r1eNFAKCRgAYkdz0YTOGJsRP+3CFFSJ7OvlvXXhX
mnJiz9gXCc4H2vcVhHKlWyczXadhjlodpEh10qeKtAXV4S/SGlGxM8k5cfl4hU8ycka8P8t4URF8
i05FhapDobE6XgiL/Gt/98LNTKdVSXDtzEQsqz25R+wBST0gYwvKCW4ZeFttgbwvEBxDJMfnWyGO
kXPTVfX4OlAn3scKZsUFldgwQDl9JFSyGeidLAu6kTmCudNz8yLcoyOH1fcpy+HmkDq6dKE78yxz
m41DVSZZIBFfUsc77qH4chb+WhYVtfiu6zgDQTKE7m0UFMMrRP4rqyPrEkx/oqkBzI6cdVPunzZz
LsHHdaORRTBjz44AeSLdZ9rsb+cXtkUpc0ola5QOvZ5FMYa3tfuRMCYR31dqTSlieiDy5tzf4XYi
qwHoi1eukmAYG54ZXLlFPzsnfzuk4a83NkOfCBjHCiNnlZbRMFFqvPJm0UGYSlLBW+/4AtYjrYOD
WbVStj/yptXi9Ss5wPGdy8dZYV7lo/X2nuEeHoH2AClKtJ1ifF7lxDHbLQU9oJHIKg4gnGNgTNTp
JzGzi6gTcjnNorJY9vyBrxlBX00tFRAwpvv0tyqSnhK+BbJMQf8sd/Ld6oaiJ07M8ZT7uNReUX/q
gPsY4druaBOVK9yqI2XvfbxIOmuGxlL0TB4wE2XBwhvp2y0j5rYFo51xAIH01zfdf31NVH246KKk
/NPqoIIg9DylSOnQA6hU7wrVbR1u+GmE80JJh4k/YPlrhkwvA+4JcHCVx14taaFxbfcYFJ3Jr4pL
GavnFCukBWhIyRo4m2i4ySIB7iI3lUjdGLfjnUyM+A1VSiuGZk9D7HqM1gO6rvqx0pSR63vNJdkn
SHiO9O4ZROzamGl9Hh4KDaEFb6EUjyAJZH0GJWYsf/1hjbosjUz+PDoxqMuUBrLycHv3Vef75b73
qfBSzp8pu+BvZdV5Aq8+qddHtVkLu0WxxiNQmTXyEz+2g87e5ACutgzv4Xp8tv0+lfxGzxFp3URn
8rwZFAgA1UFNBR2O5sOaLWNb49vEJaMt0uFom6Wb+0XeguHkEF1mII6fSd/ju4NyC+e6G3XduR3/
Bu7Mp1dZFE2m56DVtsdq3mPjjHyA6JdUbVN2mlWuZyeQOc2hGlpM/OXSy8g1i7ulR93G/z9mrgqv
FHzvBCHVFz7glTsxFzQf2LXnqCdZeCBwgOeGgqiptI0ckMXzzBY8qZqM1waBHJYQ58ku758/VsFR
r+LkyZz8HAEQJUfoYXRkPu0lzfkU2ce1AAZeZVV6LHyBA4WapSEvFTyaBzuYA5Q7MgZXDWeCyVB/
dDWkz1KZeq8To+kUfyW2UkryFdajwzTKs2hYspb43zZ6ARpjhf8QK2lkSGg4ZJlwIHVCrEnTFNz8
kN1T5H1mi3Sa2slofSue566qiJfxm/aHzwHVnSlEUu/2I+GN87Xty77mvXKcA/5EJNjvouy4zQoJ
da4CZebMWEdXaGePceca71ZwuWd/kKouUuF0iZC8G/wOH4uhfHCVMI8EjylrdZ/bQPe+I0ZTxUn9
YNM2BiJPPuY7uIQ88f3poLH4NiUyk3ppgUdeY9qNdiupffy1jiGc0WTgac6+reeE+w1h7gb4MwmU
XkcjCRBk1RFLJfhUs07dQU5uzMyUZW66w+2Pe9ddoIz3AzRy8FHbzT4thtgfawlE1IAEpxt1QYCv
DZc9Uu1GFMgYmcPbWwHRk7q/upvHcvjxTRn3h27QN7PSXPrOIh9cJwk5aqXZ5DUBCfTUEq7Yo/Pu
lNAjkrNIQTmvPlvxcdM86Aln1Sarcn2UbCNTWSSvYCaUIuesU9rSAk1J6GW3Z41FIdo6JzHfRaWc
QVRKsHyZNMjEaxbEUzvRNSNG6NfnD49vVSFFp2kZS38CVGrJ8EZRQD6RrcPjS4VOm2F7wR4PWKsH
a2SfF8OwqBHXHM4j2542j88h2kqBzSHp7Yhfqnu+uza8I7wh09UfdRng2NlD1ZLQmJu1vibrbznJ
IVP04Jlw5uZ86h2g5HjM75lkonj1SzW4UoOsS07wwQkkrX3yq37pnjd6Y8K+WCDOzsry77kHS77l
jb6zBeQtf5ustCnpHq5IFg/PC1cCvR9za/HfNC9bvM6V7NrseZKupRvEsFNMZHQx29O+V9cFquKM
Krc3j0SkE+oTXdxGqvGBlhfGeMULbigiT0EBOehQSbsiSJLOZerWQ0JPH4d6Jmbm03V+GorRUKxh
L8lbpHukHqynTyBPvjl7AMna/1SYPddGY35LCUHYRLALufGAkSmoEiyqmY6qya6r8FgfKkCwF7sB
iV5YSdf6v/W+m16MGfDey0Q2/T9EwLgH9jaok9ZmUGr2+qV4PLzh5q7Io5DSO4RXmos6CATwvw5U
MMKM9B3d1r8ZNAX/JGq9XrP5oZYNUK8hor9vrPj18kaze90OOkRJNRP1TwthGL+3evW9xI0xyDSb
lWitYZgWM91QyHESq9eDDC+WnWxtL582FogZ2WSzrifk0D43jl6TtM1RPeCcIll6YuQoI5bJDyuu
yfHZh4yIKh/wH+lrLjDyAGiRsDZqKYwfdyyRuOy6EUgsYltHAcn+uipC/UI/RnmPdYadkqp7sAFn
gPvP4N+EYFlS2lU2xJB7IxmpMHElcGqNJV7pQvkDMWGASq1eBE8krf6ct83BFdGBBIs/krbQ73Yw
5ESwA+Tl8t3xPuVfoA6Ws7tM9QZfpwJA+5KwxaOqlALB9UrKLYckpfrYWB7Yd9E7qKoxZCvPobHK
cEMXVQOI3u4jndHyuEiqrOqeW2wuZ1+k0fJNkRM7PJrIVfaAO2IRXb+wbcsJFa5WgZgL+8P6ag+I
rpNZSLxC5LvsRcFDGu+0fx+d0202a0fnvOdhEwvZBquiJg/rjznashxc/vf/cQhQXh/SQstjD1HE
5L+bM58di82YpukOuRSCn4TQbyaoFqe7qQHQO6Ju+4wgg2AAYKFdFwiBDD8afI0hOWtgvM8PNyrw
v0y/AX3VgjJFEMEKFi72Wy8CQEzA2h3Tv6bLMY+eueVjhluashQJqOKtW3cOCXFDBOCgqlV+qxFc
nBUoSdEfWRkDCu4caS8TJUUrDB6xh1b2XUkvOZTv04sD/Ypn6ydA9sOBL2PyoWzbOTdYjCnOh3vv
dNEBNf4GcRyAxaG95GESDggg5xmMSeo/V93zT+e9e5Aaf2ShZib13Sy2qYuXqD14rD9KhSJVoKlh
aXKedn8swjpppKD+xxJbRiF763QzACfBC7gn2+D28ILSd6Ueo82/lURx+o+FgF2AoxuaA7e91Bwv
k3OkdoSt9eaLVU+NPHX8KaPRKCMrUjpNrH23cvdd4e2q06sIYvKnlnKPqW239kNT1nhH5uDQb7ci
FnrA2Ns3xy80auFhAMkmnW+DbiM9aXjJYi5VDvrAh73GUjGNAvgkHvG8aucCxpOS/ar7nJNdQnzO
S4WdWiOa6Kjaw4IkHQ3a/IC1+UMaFBAMyMTv91IbFcvUjat0sCb00xR0a/j1D2BkR3q7GilInzf2
AnXRP2HZ0rBQrUDlSGV9aPg5Ir6UeN907JHRin5jh/jvT1rUBH/bSzhtb2W7NnLz3of78uwRa95H
XZXxtiOs36ioWD8WmhArcrYo5ahmOdooTzM81zt3TnvKoVK9sQEUBhN2/v5fny9qXRk+l5rMud0H
OYE6Wn6O1jkbasBzNAvGtSA0OK3hTpb5naGK8paFacJETGwgknh9eAOBR4pfuXhalcZ6I5HM/Xa6
1X9V+6pwgskNd6L+6GmmKOXZccL4xeQ2PzpLab3Qu8rCCoTMiHdQl6LZY5u9fhoWke0ZcS4AgQuw
Osfvmd4MD0wV+XO3y06KE592AnzSE6GmNSx0rgX/xhdGi5lgYeNk3qQ34VVgmYUBoa/hDhewxFAV
gDlDzv0dIHmxxihTDKX5vI5wLKkWfmvSbFGaU8vpBB335QyG9sBoczQFhRbzvp0m94n0bbG3O+3l
IDQULH62/hHkJoQmZB1bPsMoqK4VSBvpClhbpobuTFksbHLJG/sbenDFP6jKqk80EAIhUFhkgUQP
tHa+J6PVqZ/cV+SXEvL4xfSlK0qjcsxM7+IyMqku2QxiV+JLorNu7IBWcmNFB0R3tgLCXJ8OGeCU
j1by3QA+6UV5/DqJPvQdvvnFGiosj/xr9X/p4VferEwhLz5lkTuCapQ9xpJgolLS9FSifoC6TvnF
Jbu6fhuI2XdfDQ2Cubsblj2mZ+k0MCewgbUraxb6fX6H2x2wLrsqkoHUFTPqEuOusf8Np0/LFlkL
vkeXy92ihzeRehDpmivljClDmu8AhMKQHHWDO+DePAOnXbFlBMNmjDgNpJzKn0QY8INc8uy3hLWt
htMloV0/5oLll6r3hjHFSOtBfpBLGlliJbgCm5B0KmgABC0JjnVQVU4QlRdsednaOoLTffq66h+D
gtob9pmH2hQr2IWNPx/csz9OO4j3EKGoyM0QsVhhzlXeQyMGFvk7a8vM/aeoE8lqE7CEbndr2zma
+U6YJ90uVKKn7axKluAhfeGxBnn2XhsoO1bi7uhOijsu7lTYI9j1ULkfan7IT62nuc5s8gERVHvM
jKY6jFooMm3QaS/XvgulXJu2tyteMGU/DNP6r5NZwfcI3KioCvCxK9bnzxHZVmAHQPLzOK0qFdyM
W+9lHGkVayN8LCJ04dJs+vrzxHv5J7fhisAzDyF4rPGglKTFosMP8iYbC6gm7bx2HLCjEK0z8ceV
ZkbmNDJa/jwKUxr1l2E1551Ib2ZqeOifP0MyANmiO90iqJ4GAcqm2GFQ24VoasBS1k3F3bQ4aDdE
aD1c/kjT+o3dOK0XbGQYmxVM+2ioheRuHYcQO4bphDEN9bkb+0oKOZiHPvK6c159Mj0YYCc98tXk
zdeY/3SW7u+hUz2YuDWOD+66JukovNtQVEkmXTksSUJcHazALtgtupUA92mLbkcQUFIoKdh3l/1O
gOO1tgRDK/H2yytbOyiT9mh610WwkFo7PD/GeBosxdbvdJo5F/eY05bkLQT4TWYL+66kVdE5rDOe
S4cWWwtw6p8sx/YQ7LaMX3kAn42uuTRTzdtZq3oiU0wx0TErHkOuyxOCA8EeTmeYp5Wi1RUkmNa1
IXAY5dviAUQi+hSBBzrAcLjQMq98zJDPlK+stMDgqegFkgwqlrVlrKVGmYxXS0tJgfaqhRvbsBlw
/e7uQ36FInjVjyEWxvoib9S1D9Sd8Nr3FOU8zBRuP1ND73zO1deJb+qf7otMUU/SEwWkz40BkH5I
b9cJmiEwIBDwJNPPMY+1nbbX1hNSuEeF+oW4EwNzk/tVa1tuH91LIRdTxpr0scFOewODM4dpg+tJ
yQ6mjl2SW/j8AODqzAbMBDgfCUbVF/Ehzn5GxQEicvPXszNi84jwlzA560YUKXNpUcoZYz2UCKfm
z4qraTzGPQ/iDDUxTxcLZT/H9OacRaH0XfCFrXgtn8RM0V++0DOg1P9vVrSL1eSXDA0MXWNffwOn
KH6HIYy91tgPI5uUFiEmo/c1q1s7BG4bwrxAMOTSWrWQmg4PMOEKhJkfHAYAKtaVArAxhLl0Zs5l
S90PK1kJ7fVvlZ6zWtABtH1DgGKqBtn1/pwuBKbTanI3IZbgWLSZRcCI6PzT0ry5xkHKXwwNW+BT
26XqA7T4fzctZyoq4ElSvhoUCN7VA/DPllJ/YVxcJWQ8hP2BDm79h5mT3vuG+p0tpHKZOdCiW68W
Cjay5+ZE/8evguu3Z+F0LWx5gcyl5cluD0rHHTojsAhzbLwRwQcHkevZXYC/rt6dE5v6NJ6Mbh1O
x8y/o+StKgx4AX+15UyghuZ8SOTmxUncf8SA/lNo/sFV6M7Pxn+ZbLj3gBfMZxL3GrPq99n2q7gu
rvrThmA13StWyJUD0mAhi7STllFzk5nAr/WyTqVgpbv5v6y9h1olXI1EKKcBuKv7FhvtmhhWj6AP
22E0vJY0sSBPM0uRRu8Tk/jGyemZXLBBrAEdbALH+RpeIPBXugPzLS0Rc0Di2EqxwWNpKmHrhwQc
B8w4xRBKHiB94W1KCDe40JsevIXEAC9tI6XrXsSGIvaIlcG+lKmD6mmDKhLGSxp8S/9WipdJizwK
WkjOZurN95hpNn9BECDGq/Y2gJmdLUKFkcW/1A1mU/j4c1CbSSl6WOwMDPfwyQxlmMz6FjulITJf
q1FxRyWlIAdwFhaIq7d2I+CxxY4emWGLEM3FN1lzW7IB0y9Bm5xNBneWayMk+d6jlelFICYJzs5s
GOptK3Ev4aGjOws5dYVUXIzHp/UK/9E5n6NLEKL5RDwEsXmXsZDPhkqmz0X2HS3SWMtSoPrkk8ez
3DFt8voDle9a6PxPwXxB7h6R7MEsDYN20A3f96DAVTcb/JRoDPKCKQ7NME65a8XArNGbkLpcqCJx
KJOA2FqtUdoK3GSBQnc3bCaAtFXDCmQCavt78xhZoZDyVe7wurA+kDXjATfzJUNXCbTwqoiiJjpf
4tYUMxaO6/ylroSmU4ARmEJNgqaukGiBhbQtgCnMlNCtle39nfVZoaIwzq6A1x2tCCcan4L8h6nD
5onobATh/7kxDrG9Rqi9MjSpMfHsIHybNH6zVvwMKj8DZlL/ZZZi0nV9afZbvmZwq88KXdg3JK06
dHt47rNOBvIviQ56pEkZ0oDqBKBqnd1QpzZ7Xh+tWlgzYCve9yNxpP8esEU44sRsUrsy50X9I6H0
Fb7sON+UmJpvObmsc2HE5Hltjhvf5rm/IJvdXFP4fbb1lQnOQDonLrEb3fPzyh8yFK7bmaGD74/V
hbYSjJsX17MlygXOTrrcn/loEPhxd0lsOUtWD76OaRX+4D+gul0BOjntuQRifUmUo2ZhH/y9T8qt
buZO9hiNmvYA/rTh43j522L7ewTferCqMEZljRylHmUTvLEjgR1xoW4Q7ChK3EIsNA03oDNbRXiY
VsS+R5kBO0qjXh0mKjkBZJfAdOgd+hYYwk5LaGQqukxrSmsjXlcfr9hY63WN5IVPqI5u3ASriS3j
hFjeAcQGDlES8eJUH6obAAjzfPA2vKeTNU0AD0teYI4a4+A6RYCM5OYeyda57lBL5YjbxmMCfPT1
CTNdpND37RXB3mLL8tCOeKmfX7TtUt5yPZs3ptuXyFL9rJcFfbDW9G0YsE0TkHz0UwvKZGSc9tJl
Ge2ovIyVSSiqwwZ/SHqV96EhgkJ5joPmaXkFzTHP1af92Ek/gtG6rwuuzhJ/q0ocXJieXYDqvNww
6MP27wlda/OSYAcqCsnWPTWNVKdWvZgBiaKwNSKqBzFK1lGv+lhXiDJigZ2YQdf4f34xu1B8UOfd
YwMkz0Pf3791AVAq8z8yQ/0r3Fzw+2q9wXcOeEnLBhstrAoikDOtqbKuTiMRTpQT09OgrjaDQyAH
rh4kKWO60Egr8XrrVMk1N4P8j+pitYsZxU1st9Q8C7YmVL2ZRP0DJj6mYYfhv0I1UiJ5k2KADebV
xJ4TzvhE4pgTZsYPZTNlxu0hJHDFlSYNG1JJWMG/z36Nk4Ib/Wd0XmSXnrSpp6o2EeP9/XKqSnfr
+FTc6ioH/BOQtUrsLDSK//6RPFZVpROfUvhCF9A8HaW0S1WDn155KMbW2cHiad9zBHhvdmQjorXp
suvFrw0RW8P1zPGTzlbk0i1ODweg56XsIMy2Z2TeytqOHlB46VeCPGeTwkvIiuf1UqRLwyXCIRaU
zFojYprOrDBZiP5R86UfiaIhHu4hfszxxrHr/24KtKEr+gLMAKMRzQuZHBEmy3Rm048MQR30HPet
lFE7pO5YDiQpDvcCPiuS6tSqF/2mZllvhI4V258Uyvybkgs/3+b6oNp/yg5V0eLyYzXA3rUdAdwZ
EhWqnfQisJNisOZsWILiwBEO3VwSUqao08b9BD0uFSFRArAHwtme+LB+WpI2WoG3baDT71YX6mZd
3hWj1Ni/6pUw7bkvUbFFRkx3/wf/oq0KGn8IuDw6txeMVVFfOV3vqn5x0WcRdud+A57813LEcBKi
DCcdPT1V+h4Pp3QSt5zEL8/uMdYkFfU5q/0+zaeaOv5J1+xlsDB5cNWuPSHy3V4ekdIjM+laR4v3
3xpYnmtR/ZMdmP47g5RvB3N4emdWPhTFmzmzyRKGpNAoim5jiLEQKixE6+ABzVFTDlUEcQk2Y+9R
RVEqsHjQsbbNRUnKKfxxeoXrQEAjgT2GNBXmGZ+LlTo6ErxiXPZmKXl3SVZOI0tiuvHaCDkViPb9
JbN/LI+oh+flGafvM8XOPaMj/NeIKgfOz2hgCtYmr59CWx6+Eis0wzlA+LmtYqlPyWjLrSWE7vRD
XqtLb9rANM8JU+7hRMXOlciJaFHcmEDK+tNYMlQjxzhTRmQbQRynTfjbBxyf8vD1Bm/auQOKR2S4
I16jC2+wtgTb3KTMorjxqmVr3ICkVl9Ul9bFOaZr2XVcfi3ShU47n5F7hrYHkXR+4Lnb4/Ea0TnG
TbfCHFxWZ1gf95MfDjFuTm7D6Xx3iTI2Ur1iB71K8taQQHVcjapjQlN/4NcYLIRMg8h9KPdp4a0n
GaaXLJART6ms11tE/YUTpKMh5CYfVtQT8KWq0Y+z6k36YehLvh78/dm3wKtzT7tIOeCPIPBo7NXs
mx5HUrl7qUI3PenZI9YucJswgSpA5yKCjhLM7Oj2ptGTPOCu78/xBMbA/wtNp2d3kjLYx8oiMKau
9lB6cq6VktdurYb8F/feRfiUEBnAze0hJPYmGzsjWvYrtsG3Y6iMSXRrzi03GFYqKYjXGQenfDZl
s5y6oSnSTkCYTjusWQRWotzKeH/LFVKtvNOoEOdWEvPu4FZuRq59WtsW228q+45gl7c1Rn96Ad9L
Y21u8D2eNcWlranhjlLV9s+WBG6mj3YJlheNJNxmfhrtddxix9dIfqT5RPIuUgVuO289h9YjgXr5
GAqM7EjKccXElRLI+D6M6pfubV2PicBl3Qpb1oMMJvnOMucv9+F1Y4E/DKth/FCFCCBtFF54D21v
zkxo/GHG+4+CcExlDFfL8GRCrz6BYLBprlK0aJWU7jXuIHvHUa5QJfcTYIKrTBPszQ1O8S67fTT7
JOIKoCdJT18cw1y6w37iqvcaOzBp7xL3IcAutW60PYg0f3z/WgP7oXcHGAJA9M/8IcmSFkSxHzaO
pkqzQnRTBAnebyff2nAb5z+Vz6iRU1y4mTNxXJLMUyV938udDED+I9FHMjqKt7MhbZ8yFLow7zKm
SvdWCueH85HWUJ4xjdNV8VrUrhEFXd1fSeQ+PpyaiYaklmDVi3a4rpK1nkjkRY95ozmpOSlM2qA8
Ekw5ZQMnb0ez4GUXL3nOplw6o6c2fMi/jDg4b4f6l5pJud0LV9831rWxfIywc6bLucKuA67oPUVV
qVyAY67pbkAxmpGTPwOtFyypKsn06fOIT63gQlrAQHye2ih2BQF1CfCi8gnEvZUUoZK94UKMxBRK
VjO7gg4Cn7vcvahZKSHTSr4d1c0VQGbt95gOrS/r3WwmJzoRlv3T7TTRvdgCjftJrdr1j2iQKBYm
+4PN/L2XZCPTOpCHD1pmY7LjugiqlSI3swqNcJwl57DSkCie7W8ZtHJdYjeBkAMHOrAkTL1qs4ox
zElxqo2zTr12s8M06bqXW5Xhx/+EEnqxYvTc8uNGF2QbjmogEiWlXuzfpN/hU/bcy9tXBaRqiT01
91Up0WlVT6Cl8HowAvrC3d9Js2Q+XdVSwE+21gT3xFAuGxQ9E1xA800dnoIG5V6jobeGHlcAed/p
QT2vf1Pu0SBRC+aCHrAZOSqfuisbg1F6HoyY28LDG5KbARYfe/YW//rRr35jni/kYd36kjxUi2PW
1FSpwasXCNsx2WE5kQ+ZszidW/+eLk7WJEWFMy1QNzFbjj5UKGaqXPcPPuqBr6MPN/fCXjUhlIAE
o98L6HzSvo6TENvtK2uaPyI0sAtuN9Hx4N1zZZewPiwvh2C+Bva5/RmCEI1elZwtCxcKDDI39lcK
dHfWL0n3nfLnA5W9+x0IznfMfr/kGPtriWa2qs4xoyKXliAc3XACM9bb0h2b0ydZozclMmNZSAGw
NDM8I4W4CEiHu/O3tWvGKNWIfkfB8aWid4KIOtrIfBNJW5jJCamJKluIaZkE2RhnTTO9tji0EjYl
l/SdGSQ1u/JU9ifj50LmIkLxgdaKMkXYqFUYaG4XSd7iwLTU+VEsq01R0uK9aMppMpfWx9SsvkHb
Sfi+WRPwX0QjS3demz9CNL+AUkodwUkJn5yb5/J0Hzzfc/dGB19SmTlqLPhTEYOsDwPRfF1JgMk9
XjFUv3Sb60lqGRYeKmteED15HxHWCZwA90FJ5B6Ht5EiGYCXBaZ5tgClBJHJgeJuyXCYMiezy3FO
OIGNqDXrKZmX7klic4m1lHuOMcrxQ2THOe3aQZOmcqOlV/wj6gFQEGtINDL5v6NYM1Yvz18sMIxj
EIXRYBoTT/74VSyvb0hzM8T3u1F/ZFgzVmeRLzGVSmTice8QEW4Em92Tip69W3eMRtWdzZEF1mqk
hwhOtU3jw8yCe+7BY1lTRFIBk1IG0AkjEgPwzulxnsXq0/ay/sVlQYKHgDl0POI2mhGbr56tBYuI
ZSBU+qxOb7VJI5UiDppFmyjwnfDOYZ4IihKLi4ydXHaoj/H6W3iwx9Fugh+B0QZ3Os+MIoJtHJ4O
ohpJ0rYkDgrgBDuSZEoGAFcDKTKRnPR58mHkLrUxSmuQQEli3ZWRLbpoMvyMC+MnQyWY2/IZVKfe
dGA80mQFVe0Z4jePzt5WOgm4PakCrpfYFYxoutYh7nQ30YhvyQtGxH5tRIcoO/e2xWuCfhW6eOF/
oLeRe0AkVRe/sCOTvVxwj4yvLrSh6baDyZ0ewvPphAv5EZedZn14FGyd1pJdF3S5+QEIcGFUS5PX
4j385UTKkN0OjdO5n2+9iqTDBGxLf2L5SIrOtE9c2KYUGHmOWSOShoBqMIL79bkiSIKfH62OMkUw
7soJN9kI6Z1/8zWrt5h+ms6Bvhxrh2UjaB3XfqssFNeDPJiNuJAWoHp/SYAzYWSj2GjL6m6ng1sK
FOGQnV/Qe26L/hxX95tKfITMRPBTh1mp40zWMqX5GsAP7H9Dr+abrozaP83WsC2HukOhtBw2KzXh
JT4T5EjUcjztsIC6DJJyyWU+UVw15ZtRKw2Hrvz60VqGET7Yq2S8Z8rmZmOZPjCxKtOf1gZv/lBQ
PQJ1a7/epOOzV3qxUbKOyLhaqMiKzikrBAp3gcX8XGd3ywLOzo7u/paDSw74099ra/3YaTIkypLM
2xTvM2COm7+o8z/sf0K5KxxUOt3Lc+VBtRQYzvNtnuq4VJksw/6raNUnyhby/afdMujr9ql1ALhN
nwDuGH2HQ2WC2WqL9bYxWk70kuLkBLtT/UVfmJ89JVRhOKpQ9VnZXyRnalp3agC0xGAWYOkAntyX
ndNjyZe6pAhbDKbPl0cTqmjCHefSRDDBbCZYggjzmKpSHKpTJ1rRmxuuGhLeelUiaYuWD3Zg/Nox
ekoksPOtL/CkSEkCW4nIHzBawBTeqDMarg+DqrFlYbpScXFTC17szeIvYkMid0TXTXMe1HLQ419g
NPX815q9wieLpKr2nqqOhiBk12m0uO52m8pxUeLCVP88Dta1SfsF8s8altoLPNbBC/CtWU4MRAu5
WwQc37a52Zs7D4AfjQ4QZoDY8xUKQPk/41e1FwxeInD2lDwEiz1en+ysjxu1ibxwUmaLJ2k1igFT
WJKJZt5n3mCfxiTi4JFsT9A8HgGDuenHbfc1uACeg2FYUow0ciJG/s3iMsqMceVkyQn+hdsuHFip
tduV9F+yILrU+Ulc517q6cq7NUMTzX7N95re93M01Hv74A2WiE2GKLDLhrNDHpHQN4+pTm6NtyZo
395Tx/lBZw6ZsCaH5btUEvsrLZJN6zhSXpIqVPokuXpUzRJpONUZUixfvPDLRkEisTPkanpGdtd/
QCvF5IHd28wKdraSsg0pzUxnrvy9K81DO6KqtUz0zgDCPZyd5KoNf9yLOPBftUstUKyFwbmLC6Go
yBK+iT+gwxXaVkV5AIA47s7CNY47uctCA2ZS9nrbzrvQhRY8/mqoWyXhFGFpU04cq+rV9rGuPVA9
wLZLXFHdX4q7t1kfJYaiMxiwBjeFZ9yO03yc/f0DesXz4blALS9u7SEAZnNWFC3u5O0oHUYEoRTT
aUiUqG+FoYpGR2p12uuZISAT+3igFRqIEha3ko25BGZw2zSJYz82HTWx2NWBBOZHUsT/oFtW/UPo
Is7rpFQIw3lIEYMbMXyaQDA5aeHxG0tagXPyRKTHfI69e8uxD+GLMKVPo9oYKp8Zpghk/CnJZeuN
d1+aM645gUMrEH7f+hYlDgYL/HmmVM2jN1Ud4BMrseIAV9WNeYuRiY82+8G8AG3V9GPqxgXOWt5q
d88QCbmXEbbzE1QoQqvTYw08qvfiqtbpnApJLJyRNJSNA+IF1Yh5i5uFuNw1eQZosClg9eVnKuSz
rp3eLkPJbUabUTJOyRYeadjdM+dQSF0lwI/GJRRtNj2VcB0Ya1p2j3L0sfr/0JwzkvSBPHF4OD3a
PXzpnMiRWcYhrerM4dIj/audxL3a3sS5dhlspT6Q3iowQz/vxFKQSzwyXnz5edtY+v+jGOSS2N7l
QB3lchsSKZiA5CrQkCw0Ug49OhiZ5ptPi7GCQcb3YGsrtNVQr4vYOx6nxx/fcgbDxMqtinD6zZLx
5Cum0pmX3LX9kf3RJOJkuWoX57q83UplOR0YnQB7VRrAbd9zMjYfGW0L2gw3mE+juwNhe9iDRfdB
tArItGFUN08TkT3G3AEAEEmYvkbDpgS1fHy/MZD3Qf9CsaBXAKscuA1CtyJgJy+VXgKjyrOA75iP
hlW31XI7vxcQGSXE9q6tppoww5CKZXafFnxCe4f0BjUkZ8BzYpu5rF1WJH8QbrcrJJxg4UlTT7c+
JV9+kWSSjVQBFyjSzi+unIYMS1jq/JCILRcmAME8dgxSJ/CFPRwGPnxO4xro9QTXFhybSIKRJbe9
LCAkjpPLpm6CBLFR0RFxmqcfs0iU5stIYlZfywZJu5RQ9DBe4ZS/HAew7WubFvPZ/QKqLDGx1ma6
EAA1kGn5Hx2tdikrYYl5It7Q5zw9085joIQ3LuhdmI8dDpVoMQp0R9VhtAjvz52e6v9Ejn85bUZC
TtDzjfxofP49N07vR25BQwKaZlNjrrkVu+awaHIviGNWSO5bbqd11q08BTLJKXGoF5Od8aNPzO6E
OmmDbMNXeFSwOI8E77/AY8IZxXzBK5wchFojnhUJjiRNWg4AjZ6GmvT/BvBAPMBBD/x+XBMB8i1s
vReXzWNdGkQJo08tkbvm5c2ghLuwmIXxwRhllhmbBAGNLe4Z+UbWfy6OScJOjNz140qTDf++RxP9
BECvmQnzJbfLTlMQpqeiChBJIvE1P5e9sko3Y0eOJrXVxF563Ti1M1TtGW9yFJNaBfBX5fy55fo2
JOR87N6kYA3gZqWSs1kdE1WfaDgoHK5o4zQ8T+p8U1DkW57ELdFxd55YysYVfgNZSw58zI8wvVk2
rVv7OjJLT1j+SitKrSZ9V2hkuXeite5rL5j1NvYlaDGoihZKnUt1T4o06mWDySTD5JypEGWUn5Do
leBosGEr3yrzQL2vCF0mdtRm1QBOE5dQwS9LH15kX0Mk0pZqKE4dVyfh6IdUpsphboTzUWjBdj1e
4af5FjFNWisYikuMlu+U0nqj8r8FMmqaGdTHrHws3WirqRtDb1dBK2bJdiWAsqpYGZBL9+7rRc7k
5tk14WgXfYFGwhK0VprF/8/P3j+OLO+Nrvf1pKana7RUQ6GLgNIKap3qFqDof+ynGmPZ9vVf2w+Y
o6C1R+2+xsVvfbPymSce/OJCuTfvG+CHAK+WVAE0RpqgZDu8fj/HBdf61xZ6sNeKnlozYWNZa18L
AnClvZI5XkUsPsh8WRJjcAgTVc/Ot6S7PGzn5oxE0K9vHHiHqUBy+d7PrmGoxMLwU1I5t+fRtzwW
bAzusaoXxG6ki1Ei6yBmlJeXJzGtiKvo9oAq4zk0LNBIEo5bD1JU8VO69p3o1QW7BLqBR29mbeUy
DIMexZf4/23H5NC+yDEupBDwkoZw/XTfW5uBoj+wEeGMSefnlEZdCSWDOY9p2cVISg0+eNXNbUeG
dB+1XGCyDhvmnPEAsG3o8ZFx0caixvMKkDEqs1P5LCiNFPpXRpM6KWM0kMDxyq4cDtTK5vI3XD0H
FLKhSBKgjk3Ghbm+3mrCzr73m8t9AW6dysFy68w6bmqNdJd2t4JD6fcyovjIBPI3qQ1E1/mUETc9
cEF2y60MZHUVMWrlBov3defGxY08ayTW76UKOJBmPqG5V9lQsx8HQjh265iZPnJMx37oAOEpU+ji
QMVDq7ROn+Xnljdol3Ee0Cz+2YycNPWs2Z7uWtKGldbI3wLY0Z4ejRHnhmcIJhYBsmjv/xJAKyj9
XBMCvRGXb7qkI4qkNArwG0F927wpy91lBa7kWc6mHvpOhYCYfyINgyGm4xZ0PSkDujyU6DQWMDpS
urP6wuQnz5JsxA36s1OQ6K5hJJCF4S3XIoCIKO4ixIBVswvjcD+h8aYxVfUyuD5pJLPTuEi0BdvH
QVIe+DQ4wTiHQiOIGoAlyuRoi9OZzcJc+H7lgCtGgVTKRHywKW8FKTOvoqbp6jjPWxfScLTa/vIp
sTM+T0sCgCkRszsgksqSLb4LWppkm9xyuClA/NN3ouE/nIjmSfUm9NXvADsCeYs4NC0PD05qRJ9E
lKFgRSNCt/8FbOlVg/IG8lmZwh4+fdJmpNgbwil0ICj0v2cBYX2Bdi8Zo8X+7IvxeTLaQMzEF995
wtImW5cB3F9ap81yCEtmuZo9/XoE/sNmRIJxt3slJaQek8t+XYTgaF1kz++NMjAN4w8X5uxmq5Ov
KHb+S6CNKSAVs34bInWv8AEcgFpSjOLdOxAkhr0h2mgL+coRIN8qPHBNO6lnK1135g9vZ2VUBySR
eS1v6FBe/TO6Upe1jNxPiKJP5BTzEggl1TRAMZsD5kJuyLnwFxA62I0lS8KtPZh042i42hAiV9qC
vge9MbKaoUY6LlsYmbznsNRH4IE5vbX4xjqeIC1MDYp4URY0zF1m6USRC3ymqJk++rmIrH0Eit/4
2JWKnYRljATETYySqaYWIHQM8bMo3T7LJkF2imQXF8D/CX0ytyFGdK2/Qmus/FQHUfcqYp3aKgvl
T4IcW3b056Raj6NkSTI7o9pSwyIim8FXXF3gp9iRjpQnfaWXvMKbwFtaaME1vMxQr+DEZvnypyHk
190CxJ9T8uLBo3v8Bq9zBc0nihvOFWeMcX4FykGlWZ63AtwKl3FIx+2ZE+tTeDjrGhKKVkASewm2
TWEbjWnOzScGJZMhR1/WybVBx/xK9+CueZrm19fUX3b4WKrYjDx470siu4m9qNm/QiUeyCWmXLPx
5k7wuHTb8xQBn52cs+ipJqSsSBRtSG65WQpSthh3TXWajFqHhIGa6Mkum5rfdd3rmF2G+ORx1eA2
CFFWPrLNOcc9o0e2deMbY4jBTw7LbKcpLauAZdGBV2VFzMVaRr0lL4zCkCSjMEyXUlMAiSRrqWVS
mcHAn3qw/A2KltWa5fbfvbiiW35ITBh9Z2mWhcnaY1OCyyiA9dq8RD4Q6VeX/918ggbw+4qfHcvA
FdM7aKqpL6RP5uBFvEhkkaFNZCd4e3qZ+9L3P/z1AmQw+TDMUd+2JU6Cmq4o5xh7Ww1RyBvTTc9u
TtEVh1NZM4NK57g5160DXcIrQNRqj46Xb5g5WRg1qDXwITIXTqGNynUkU4dHJn6J47/93msh8p0K
Iko8IYVc0JAwyqDPfoDU531kBrkh0GTbflbw8dDdIlrZBrqrcn2MH5daQza5ujkGvSSBXoYeNx2d
JcXu7ZqU8crEVDnfRxAMpNtGO8y6rDbEeWlh5bTm76/c2vUtHvO2dHmUyR8CC4rIhmuH2m8oSe7l
LVQzhuqMb/dCi2VQ35frxuKuKTySZz3YUiwcG5Amadh5QfOwvUawp04Wyj2j2w+F8dLcWYJvf7m/
U736RHLdzUh57/rG71YdAIQObshEdF5DXjIHpupDTaIR62AqdrpbDza6CsklM6ura+LriqHlEeRc
bsnnLNZt8DdTeRoCQru73ZAnim9SPxOFKWHE+F5X8DnzJiYIspAHlO6AYA/WoZHYUHUpI3JRksAk
TdPuiOxQ0b9JZhbgJqlahQ93MmpLoOhLIAnmaA9geaO3e5ixgNxEpd7ViGSddlJEBfgSfRa5h/ql
N+f2j6NSb75o6V1DyPnLYCuppWT5EWI4pCRCkmBmzXIqF+9uI3YvO0jQDhOoXPzXDon0oEXQ0Bdl
2zdozF4iO6uF049vc4VeOGDTnTNKCJB64J38RwiSPCzghsbfNJdNre9fgYH9mqNduC27oJt/vuk9
R18s07OXw4wElATzdz9izpVORK57dG+mPqpsoPaFM4dsNQBWq72DyWliay5hXQh15eJFf6fPUI1A
5EvlE1Wn/jOMXjqgwRNzZcy3K5UcOr4dj0oI1m7fnF1HNn2ypD7P/lQJGqbAcN5JrNC7WELlWepz
jk+w2ifbepfhZc/IHcvN5THYQWePaa/joBQ7/93TUeluv1lHtmpwYcMf8D9WGdeGH8N7VqW5Ve+p
8UYGCJkkOz8XO6Zt8clCKasWko1f3uXC+S17MWovvg5tJ9748QUhfgFU4fZNWqFh9nrgqCqMAAfg
VCmsiRZyII5/dHDG0QmJy6ke6nXU5+lDn5vpzZX7skrfDFJp8GVHIqBAZA952AQLMdhAU9GCA8qH
RfQi3NHT413+b9Zo62CnHQU7O+2KZ1PyKsMSXkp8TPOMnenl0doydbgq0RxFsd1GWCXjRQ+BnVBM
5Ppq2ZjdxvyZ4URZEMqW9KlwvDEnn7x3erBqfS6SI8pAWZvJho6D4Xno9gsgRCILm7zQToQdRR1P
vc87fp2BQ68HHjyzk2RuI9u2a30PryZrZ4+OQbk5GP7L9m2nQ1RjWNkGkbI2dIV/Ay6Svu/oIM5P
TNaKY+yQ3AD/qFvwEE9XRIfApxaZN1VNvTPmJdw2YUhrH4KEheBdAft9fXGzCrYDDjcqSt7+nsVb
4mJyeBuHYl7wIsDJP39BvuT1UE65Kw0XYRHOawe7Md9tcSUOoptjT/rSjtQP6FdkmAMqn4s5Ky8Z
XPJWVJ/hM1tagbwzOu3c5QsznpmzHpeYtFt7E8JkPVzJU0llAPBV2MmiwN1mH1HUidzcfCGEHxN6
O+vFMvA5Add4Cr82fbkjyFh4vLjCzxnYo9YYASH+uniGDBMAOLSAnWyBMZcnheKZ3fO2oJvoKsCD
VCUmSQcJOs8M/W6X2OWF8n5intVA4g3Cq9mCGu2KdEOtmiTLR1ytoTsEjXOeBoiOuiLRvPX/Xo0T
hh34HvABrXW3dZ1LHvab8+SAZkYCjwHpXGbcjK5j3LzShvXrEqOpyhfU8YxUjX01zONCZ/ZqNUY0
hOi5TF0h/mvGda2Ap8dZj8WdiOXNigQ0zZHtMYA+Y1zJUdAyWr0ckoX9wlfV+YPXGUHtQ93kGoTz
vysi7dUfl9Z0nuAZZphOF/KFj9l8LMvcEO5BU6mlZJCb1BVjKjo3/i5+Ky0OQ1UuiIU92uy808Vz
TZRf3ISrNj6bgJ2CQL7S1pfXdc1fvwyj9tkX8jlWVlDJ/5SWAoayu9z6A6SQ3Fupn36lgB1wfOML
0HN5DHe9WlobvfumIIrmlR3SLiptTdb92ImKzUlTjiSTXyj0ycOOOBX4fu+HkPpHJXA6xbE/JfRn
W2HJDXSMgHb23crsP4zQhNB/3uSZ99ZLIEUwxkMPwdxFb3cyIf8t4opT6y9cdBPWl3yBsp4fSCgq
S3pC3JgqhJhaLI45Obs/DA1yvcHrPI7SfDhyhCYJU3DdY/LbC0gj0Do8fWDsfwSumsXia8Msuw59
BRjtpZaFMBk14puhoflXs7gu6laJgVvxWIpcVo8GA55G1kIzCw7/pY9HdxBWVUwbv62wlad5SAp9
DPuAnaZ/HBoSTnKkPx+QYXgtye5HCyXlStpaCnElIGi8y/Z0UB7UQY1n6WwKNgQMvlNxkVjuublJ
ZOgQYd0yjUNJQH2gCJicTU8ItJ7Hbm76XuSxYqHbQLWlGob4kH/Wq2ZsHjQLzrjHdGwT/PQXEfaL
DgI7ow7cDeMC+yr2XIgOqOG8mX6F6CqvmjvGCyfJ0+rHUSjurfoC7OokG1vIb632aaVlgXmnVYes
RznX+Cvl++BfboV0gMXqzcscsMeGHRNEQhWl64ESj0fqK6vBbbEw5CdaJIwwJ38P+76X7+J1+jtL
d0Q9Rmo9r4YXKACHpWFYMb7KuW37QHAKKnS7Yt0b6bjC5gSQk/pIa0DneOSTczKgD5hLtYp46uhj
hU48/mm+Hr+YJH56W0qE2HJoh+d+19J/sbBQRE5b7CGpGajhdSXWX7oRO4ivFK1oGV2KnGY8LrEN
sXn3f2kPLeuL30MKDxU43dlYSIF/N2L7pJ9QWNQylDmV4Ah1m0BCkm+ZyhThZpaxZI83M53b5rXF
wSMRcei+QC/WXXaBvPlbyO/rZpElPwh3xpjVhcX/9yuQa5SSXa7jGP9rfO9lTi6kcZrOrK1UiV49
SsEJNKDp+ZSCTT6wWGM2tfc+ScOk4nRYxYNz2kF3K49yDbfaKfhuaoCGTP5srPuWk5e5zRftNO18
DNP4GUXDm69l3hk3YW6We2HIVgULi29I7Bq7mX8KpUhRplcROmSIwW1JA3LFhbvk2Ey5Ja+fYWdJ
c9eIc/hAiT/ibhaZ5T03MRRO6Vmkfl5WPFEQCQGyGVA13jxuB9jGuGEHmhzR3aWir9VU9z5NsORV
+Fp0vhJVSLiZmvysMqYp2yTqux/g3kT0GDAuZYSAKue9QWBCSRi89Wtwp+V+OnffRkpY3JGPNNx/
JgV5XhvXqP+CIIOHCTtRnM+MUFy/PGSoQFZtaIWcf8z0xr6SQhwSAPbvaPJSX3rJCJoY9xfjFy1k
HTrh1D4Efwf/O51lWmFDS/5GYAkCRqLvyk1RvlIlHU+Y+apIAbVXmjD7VP3UuByyl8J/BDvEIDwW
jKe78n0xs7ya1VBAjFyR3Tn3j+g8HhxHxYN9h2ufzC5tpHxAJWrHlLpF3cf57Uoj9iFj5UN8ILE4
bxzWSKMoT9BepHXCDcBW/kZWLRjBvn3DvUl3rXZEuUqpJPckMjK/yepYIMIm/GN6PWB8VyZq1LHk
dv0Gcu+PhNeSAg04QyraAMu3fk5Z6gPTN9xwDW4jZ8lLURG4Y8kJ+/uEtdBgXzew79JeRuMUKlMZ
ukECKIvFsIA3y1WG0e0T80ypC425oCdTY7sB6Nq3x7yMgMS0xe24Isr+f75BYXVTGUvSp5Wljjhx
OAhoWLnBrLjWO9oxUC1YfKqokbP3lZ8iDUZF1GChBunAiIRJAuA/GtUz/bQql1THvwJ4vGS8V3NZ
7lONEm47Yzs8g7OPtBTmNpww3uYGztSg6CaNETYgv0zhfAo+P+LGQP/MmkKX4b//bDsSN2t9f2el
8r2JEBMoFs9D5ylgDFZ6X1tlyLXz2HRSXcGhhfu0aw6tCeQWKbjKL/uz2wJe+kM+pL2idlqJHRxz
mgnqgabzxwlaWYIY5SR5tAk7NBP7vTf6EXml8iSsrqCCsiPddVtc94QwMoVDXOyKyajFHQQaXikx
5tv//zpjrDhhD0HTgi0emj1Q6/DS5ZiWjPb6IrDDj+nxDXN/oB937mStwL9EigFvo1Jt4fyT5VqO
m+EvXqRBp28wws1g6tAF3dpdNCtww5zHBTE7UxnBzZ7czmIat3k/MwgxrAwKRaq6ZA+g8Vz9ZsgS
AZLftOk/ZwG2hGKJeo4WPj3Pkem01iPbf8pVIO3fD9K/H/9dhuPTTxMWK2bey82w67lkfrrLnDon
pqNvy0CGo/1MoA3k0frFi8Ww09I3NcNX0ImPXbYOABXUysYBFZmXn389HT5fv/AZ81KBc+3Ker8/
Nwpwt82GnoP9f0wotiZeLn2HQhl0RJ1gh6L33M+baevWdv8QotBYiUGzqxpmUc+wTL+v1BUW4j5o
urbShVxB+LDo6ePJIje12FMQYsbLcy2XKdKB+tx7dc/BTGFJAbnkcdTvjTn6zEvJUzZwzstDbrDr
Zc9PRZVJAGbzhtoHfIRQDrzbhP3tYBVzIwx2ViYz0NFED2jHYwOgIihAwLlmSQOHVc9tJ3Qqq+mZ
gTjuPTSWi/doDu8p8vOniflHMKzGq9x7+EhcQ9X5UAYliiML6PygoBlEEme2HnNtlC/NR6V2F47H
no67NKSYWxwjvym8CrSKVmdD8StvFGTVWn2R+X7QNuQQLzYczHMVN9mC15F/8CxNS5pFdONi8khK
iPLbz3A3RlKelj/3nRR5W3kmr2Jl6pWs/UaT+se3bs9qT91afiUIGOohTjSm0OrdyiMtq+p3ip7r
miLzkWOYSCfOnG0462luhXnuMeEAqJHyc3yZnm4OqTNhIo7cVF9MPoYVAyeyLFXdsu4a5FwGxdXC
tKr9ct7fP5L6yJ/mjRyu4TwxJdiesrANNQQRXKyZiV4jMnR5uO4i1u+YlMdxBd0nZLeX6C3NmPsE
2ObXAiYWQcIy1hbit7PsRHi18EaQhNAh/EojDzg5p9cXsc/PDN80kVctiTKxLn3GzgwFQGFBajYe
Yd0KWdDsRM39x4U2hxEJeqnKGvR1Jg4EE6PQxJ/G5rCNGrO6ukw+aKJBKPe9fdcOSyOv/sm0iG0Q
B1Pm+FPAU5H6N/q/xp6Vp1NhrG0oo+9goMPdkRxP1UB7kaFn7JsV2F7gLrZsPHfUsfE9WRvP5tfY
VWVB+/xuCVBoJvQW9/fMcQG+O0aQJ6bFIM0E8cHJ8a6+VxtmAJSrtM664sFViyz5Ot7VYaf+03ZQ
cdA/EJpLQYNSunpjNiMIMZ5upTAW8+AyM/UZQ15PQyJ9uCIdk97xJ0AVZOJnbhUpeUj9hmDP833Z
Os0jfOM9C773xvHu0p5ieyc+yASc3ODFcwN8HpCnFBY3r1+6IC5ZoZH/LIcnblFBfzbbPmaBvN0e
RXY1SUbP84Fns8kADq0YyZgn0kIo4UZBES04EBIauDnGz15rQjwEBNDXGjQJI0BFG8c+aIWtKMtJ
yEfhYw0yaV2x+4508OeZbDUv80UGXfSAmbOGIPvarvDdYFkCO6CJlLr7kLcTZAd3iV7dutrFoldN
v/qTFBEMIRHVvQS08wSVN94mfip/EbryOqFKlITSI3LEnG0V344VWoTG8q4yzYO02jU/djicjAdr
qqsqE9pwJPSyiLHBv5jieGZzB0rkaKD9oV22jlz96BSqnxDqjWrHIkQvolwbt3DzSkTTRXfOhR51
/nTBVPpAaK/RJetZBa9m7zkWuWk6nWhG3ITYvbxddtb7Z9BXQ2L8rUHHi70dK7japmni1H2jGOPx
qIe3rK57S0Ug2BmN/lnPUHoLwrm4/oMnzztqsQsiKWOcb4PVN8N5QDEVv2cKEg7szeHqlWkAjipl
eTR+dw//fJzLtzP78UB7UXqfYVSl+gXVCFiGANnHUuqZgrK/xbxAKpoFGrVzV9BKf82BOl53TCu1
hOhDAwydaeSurjEv1dD5u2qbjijXNf/DAl5pMs6LSbvSUhYt+hfExJV7DQQ46hdaH0lKy1eZCANQ
8Z7lHAGOGBM9ZTJ5okmd8cJEqMkvdHJUlZh6kpBk9Ja3PoLS1NLmIfOZnTuoGLb5WJJDjh4grMC5
eToRDLJZxFwz2F6YWl32bi+4SRzOZn0Nz+8fnX/YhYhu5L+O85CjiqjHEZDMctlbUynOSDGVL48e
Q1kZZRUN9ac8xiLwRmtE9JHXNv3r7+gcWiF36nkjEAvFbesKHrvwxbKvwlFHVoTbAdTtr4NJ9OQA
YVj8WLUVwmIp5zlsoJFhnshukItlMa7qQJe4WOKh3MLCSmMKyYT2xECNyWc6MbDhpMZpc8Jcp4Rq
/RrxY1HPixJ5tkN53edrwKDJg2BtklwvRm5286U0VT5nD7Buo10DSTKq2yGw2DcL3BwFOAFcFgPl
dDfSQ66Cn3hlPOKEXOENBmoLrRJdxhANhfB9bjYx6JeJmqXmcy9gILAO43dhmgfS6Sv6ODKpMPgp
aMQadkDpmRgKaDcaLg2hozZ826ij91+5BrGgEALRiP5AWAIRkTomSVq8Dy/uPxjkm5v42oSU8KjK
Y1js04UedBzmzeKSR/X1gBtl5VCSKqkwPNrdsPcyFgfz1afjr9Y/LVfnxk1RgvyqJsimjwwICh/B
H2JGLhg9UotC0vjJDMTyuYIL8doGmO7KEpzIrWJBUNOA/qgXpWBJ2t1paEyl7e+vdatzI6HyGPRY
lHbMfHwe1WkOuC5YYHgvbexK/J9W8rYMEh2RXbcKaYyOwGzC99QjD+KDHdC33JgPiH4u8++rAWgR
7yFiR+99kxVExuP8eZy4Z4OwUho6+H7F5/ic8xlq5YvXEuW6WoBQ5DLQRO8Xb9HZ6uV43Q//iYkQ
qazv3YZfTNOsRW3O0AOWyy1GYL+KvPjRwbJk0mQpZcmDY3jJVMoswb4Nes9TnoMI0+/e77Q402Lq
FJjUs83wvutTqS/AwVSzDY2k2kZW3aBuTn/6LxI0LGfjqP6cPMq8hMA5C0r1Z3+9BTM03LqF4wtC
1BeJ8140b8lbLUtKifFIFnJiSZaOKOurmESX+MBaCoQSIvr1EUy7enG48dDtc6hRxheW1rNyz6dm
+dejScCyTHiQkhomOxeUHlEUzUgKXwzAKjC1wZmRmTCiMcbdQgm/1wbEXUB5/xr1uaIVwlxUqOWs
/ZwUJA9ix4+3a0XWSz/wwncaZ4uI+xeBwincuT5KZZfPLRlRZe/GAAdrZwEhqwq+YNHuhznrPD2S
6qpndbH1BN9mB2tS85wFv6deNQRSk6GIbtAAzfWLyGDFGwZkxBBaY/PDXXREdle2JWRds26DoHWE
2LD9JzTRvAO/+eBaH/8B4TcqFEDAsZmeAG96sjKTG+hQp56EN3zRFLFhmvroh4S3FmWtQ8xcKUIv
PfO9awhbBlPCRIkmNhAA+yJnuzy2AgrXUTsLScLfEjLVvbsjlJKt90bELX5sTyiu2Ferkllae2fB
P0DwwTszxDPx98viM2+Dmm5Frclhleff+5JdAQFCCHMOAn2uCD1ogKqDmG890nCy5yp5MhUsQxd2
d6tChJGcoKbmioaps7rvaaj0mjIRvsXBlTdSwxKznWIpFjrVv3fieSumEW70RcghBx1eMfztX4R7
va922RN0a3u3hpnPiaymS/ADx1Aj/W/oVCpJ33OiHdOS9PCC1x2jR/jNiSSvqiNWlnBozhav8LYz
wfJRmUkYLha2qtarPviWbtvETTa05lFKQ9B/2YesSk/PZe19SOqYcd31olPucysErBFwSak7mNqE
jhcAiTW1UttYEK13t5T3ftFf3LnUvRRv2hr02Hy8cnXdgA2zRIHF0StTTebFIE9nPnl/ZODuDr4L
MHLX9I5CAkRGr/imlbKJAck9g+UCUZrIvBWfdOm5LShzgpxwnhQ1WCEpPA3VuaLcfLBSsXzpw+uM
1P8ZcetCG9cEsF72VEEFlGH4JXY10TiDx94C2WCeDnKBMd+tt2GmxAzSNUMeYDslwYmhJFW3Cs1N
nSIs18nbp2f8Z91BgBrVQGroc+KycKlLy47qNp4wPiOIrS+ihY7JSUU7k0G56ua4W9lNYKnWfgYb
rLXNWH2lB7ySZe/yMpUHC0rhvO7iM8ABwDoMlofVeXpUpGZXdGrvSwIGvOZKmjfL8zIrqV96kScH
9AM34mAM98yE7BH42D+sla+q5wScsCflAg34IqjAfxIAaNLj4AHQWuNBuAMXMNYKRRau8k9HXjyZ
q0t+dN5DTUer/uZJgb03weO/WAtWHVa9Gm9MqyBX703x2amT5kpq6jjqEKPA3UpQpCKhjlgR+co6
NKFgQjhPXANR/xfII/fkVIgkBgw4KKDg6jdpdepbCQdstqHFC460TbkshB91r/PaRCQs5Yyc18fy
jZjlzRFn32F/tKv64GpMCF03OKggQEZ6GsTvL36Fm03JBoNAGuSEagqvqu42WZ8SMGfG28EwJ3uo
lcl/wzuKk5gDuv5iwi7vPpvaudqTK7P5tD66ma0psogvdBv79n9vXjCY/XG3LqPWFjU9MDxJeCVA
WncFEDcKi9n/h0UNJM5AW+oPpk7bEzsRp4C78anHYt39uq7RIW+CIDB3u5Kr7LKv/hUYaMBsZ7ld
K/2BRWGUIqxsYUvE1dXdSOVT2TceXeUJDXTdqH5xPl21e8vLY9QEjBAalwmrztZ2h6X7OJd/mIGL
2l1PH98GKwgtXCFX1/sCev/UK2NEugB/2kQbS/oboEGGVRbWx9fINXEzIPNXXVpdF7XYt479ji/r
Dilcg+erSorq3HVbcEJCKczs0jmd8b0hgd600P7u4tFmgWcH6U+d3p3LibyqDFkrTML2Jf65qSHD
imrxL1YqPT7orcOY2EYzLHEXgy9m2vm+ID05TWhOgsa8I5LQurFU7THdxt71kH0HziAnJaAZTcH5
Pu3W9W7+Uu9CeoM8D19j/AnRv03R2VEz3RsQMJBGTgFd9lSlib1xCxuDkmqgNE3hOpfk2uIbMi7k
rN/DsT8V8kN3xdcgi1/RBzwcc5J5q5YalrH7Sf6CjWFbtt04zW0wpoJvJxv8WH4nJAaWl4KxeDr6
2Kwlm8chaQvm0EE+KwsP8vCdvRo/G7rT5xCOO2FrEIuUy5MPQxrrzA0CeNaw8nOuySgwOA5mpGun
DQB+MMp+JehwnmO3kuL6dcrvf/DXKAz9tf8Zzm2ssfDBUJ5Ww4a49o+owzEWyoFPjCd1neJH9fRe
BGIUk6c48q6LWG+mrBXowCAH3WpicOrgxi6U09Zxdyt9qSnOkfO1vTh0JwAUgZmYovZWQGpd09Fm
63I8KkgxlfwU/UDWM1+6A/7rjvcxMoEwz/5AjZ9zZ0g94lkANVToxvZfhqp7CdlHPXsIpw5ZMU1b
N7zNL4iiKf2CJZymiiQjT0cLkEsEbngteLin0rhLrg/0QdJuAyxdgaBjXl7mtk+wYueTq5BWLGYJ
6y0YS2C9qnODQgd0r/5e/JurCqlp0bdQLk2Q17ccLX01rP0mMkhk0ZpXV8iZ7+xi1mlyzHSPo+IA
uPLpuiXYH3KIenXuZ8qvNY8NKHCztraD5/C5xGtnf65oim9QEd/YTrZxmus1MN4Tk+QD1v1NWayz
0jRLKePxVhgf9Bb6HEakc4bDUIdP8Ep11d2JKMEC6MMgvuv+K6fIf2roq2XYbgEmn6LkTkhJXFFI
sua3RSoC6orCd+yaQm91IT0+QgBqn7+jAcetRkedLRTZB+Iw8e0cKzP/cpj6XfN/nRKHCJ9CcJ54
06JnEZBCF9NuyFJD1Rj4ob5FTKiHyILtZ4k47gTKzXOzW/RqV+IkkatV0qgoigpEhTu+IsgqPKAT
FxAzWde9/GkWl46fB2H0n68doHyoO6zu+tunDUNSldwmkkrgILc9j+F/QkkNpy0RQrdyu1mPgR4L
IOOkv7YlkOH3yYQ8uzMdD49MMNTaXlKLZYHPHbw9ixa3Lu4C91pxhmfuR66YOf9nxZkS6bTBdjSS
q/nDMmv2MBQUjngJ8RhkdA0gx9JKN8FC/9k5/z9J0HvrPJzvBFZFZVBQL1FzfHzoQA/vdrk9B3I7
OIFPx2lsEvLfDb1fqh7A4oPAopjlGcydN+Vqq/ebjy6x5w4vh3HgMSWZTtTsCjJuapeodYkRrSIw
5ZZrFAlfdpgePFmB3UYjLrIxXdFROi8Jl3Sj+CCBpZapLQ+deMtXeJ3PtFggQWw/5ukyEpcPJ/s4
qGzL/LrsTloyQ5uRix/fd2fNdSr+YZAZ38cWckj9nzFZL4OCwoflkM8Gd22MBMHfQIS3gu4xHfAH
rdNuE3TawKr8NMuNDOa4E8CkBatgRaTuTbHm1x3LLs8yjZITHETg9gzP7wJe+1FI7aRgwGh2cwB7
zhxdfQtyp2uKoDrmcdRPf9JcHMTmqbab8NMcBJxmjmOVuCvbYVi7ByacB+wOADPpQ0PKfq9YN8sn
cjpjboLAV67vRFJ2s2k8Ku4i/BGziGRonoXYwwxa2EkhiMHNBNKxt0KBTfTRVh2T0jdffm2zZvSk
85Q4Fe9vtvWsuYRknK7GJbRiVlusb362Wi160utWPZpLXlBYG9DMkbOE2e80L/A02KIMspygwMM1
tDjbwUtIeVMLgNbho7EkBD2AxAvgsEIJT0MFYBMNlTsTftUPCG6pwZp68w61wNGd0B2CgrqQIk6T
yvPLfoOUaMu3kq75nBqTACWXcVozESeYIXogdX+etKnErji+1keNiz4QXYRTQJeB6B/9QzL6Vssb
pta/6Dl6JZCICzZWsIvk9p8OvaHbIURThzlFO86IMxyXOCUjbLZUbCa2LOC8MyaIVU+Rgco+aPeJ
3ZO6yMd7UoNeUROSKS3o+673WEbZchO+HgaEORdTjAurkL9k+uQnCXs1kFpl/GwU2XIqEy4+YYrs
iPXLoSJoy9mhpovN6Er7uyEReHx0ERfz/pIl+qQzvHikW57dlJLpPmq3ZMcdq4I9Vm+4pdIs1F/i
FaD4VC8PFuzSCQGryCjMdgNHdOBOYTp6+z6PhpEdcgOWMAcMU38Rx0C73JTQoDtbLn4N85Hp3qym
r2XjSAMr0NtQ3CnO0z+59CtXAklW43KnahLsQ34oKGdKoIP659I9qvtImdU4dqmobQyneCiztpwo
3nWnMn6tYc8O+xaaq/BQcRYyZZjff7bMdNN8QbtJ96YfLn2VOe5wL47r8ADLl6p8Zw+Hcx6JRPN8
9s+suaFnEDZYjLbV5oO4p3ORKsQbnUcGgAPe4BRto2mOVMpdoUfhljgP/AIa+8+4l+3wkR6Rx3fj
CPEG4RUhGVDfocX075IX3yZoMhqS9+Oq7jGC5RiLRxBZf1wJYYM7AQfZaRtRhocq0axApcUe1vmo
0SCqBnKioBkqnChOATrK4V5MpJ+vZVj9w6kIBGSqdvaU6Z7kyf7l8QAPygHB/URAwSzhExZg/uoH
Gc00E0btM9/NQ00D9nmPXaQU9d/y2JF1PFTZgpjYu3t4CtNSIIEPFNP1LHulejDmXjtIO9edXI/l
rCye9fWK6AQV2Kb5SnJI4WmpbGjqKRnn8RwNBf60Yh6Cnn+u8Tb3nHOCdJfQ/WMepee1pB2B0YV8
+bnnxafa4vLiBoE0G2TrH2dzkIqIfRPyxFYl1mTohH4k6pZ8GJkrHn9ligSDhzf9YXpUWxmYUZ5f
Xs5v8D23Nx89DGNuwd5/A1UfHeve1d3vISBYm4A29TdONS4eDtZ/liyfA9ump0qaiJxD4+7ljN5e
NVefHH8JPqdbzaiRmM7DJC/QL+g8wXR+6w+doGClBba3Pd/AIJeMFJ1EUeZ/yxJQgk6SOYf92wYx
UP+512fo/QhbPjbTOXAmw7h2NbR0P+tFGrKPRMsSzPjFJVvpWzlZTkbbGJUP48pXd4xEeleYtQM5
GOTCPDCxMEj6P8G3wFybOcG7gDJdrm6GI1V4c9QAhMVkVC2rIBeHXG2s0Rq/h0Bj7uogHhcV3D5K
VOdVSnziwLVKwy7XZzGVZKgf06RwV3prPZkvZg8LXr1myKsTPu2pje1BGR059rwRECsm8VKXku5x
5k2qR5UQQNy+b2riioYatfP7m5Yu/uoNrtMdmaa0e/ia3BxXZyJZk8vHDK0nPqU4HHtMh6ys5oO9
J5H0dJ0fe/Uz2gWbpPm2j0p5OdaRTWhI/swKGvbCq6hbt6vmJ12MBx8ngzB4LgHKI/GNpU1V5Rsj
OSwpBX8Goba4TamCcrBlLsoxNaSuH9EZd55vIgweb69IxQDErlNXaJ4inrxrNAsJTqwSWaUcYqxm
Jt8vGFWRs1bwzwB1Y7HMG5LuJ6Mt71i8NHl94mGcIa0L0zyU0yl/iJyfnZq/XUaeLi5aZZ22ASl/
m1mnLvfhn8DlGqyUdpxa9E2Pn09oaWahJTftQ5Gr2wRp+r7+ViFZEOM78siBdF5jzR34ASZaEO2T
jJ5U3nGPfzC9MTtqP0eewzhQh3Vvsgtdg6utsEcjGwRfd1tDJN2IfZuUC6qnvRsXpmyYnlInrwFX
dppNdKw/qCQI2eb1P2sU4YgaBeQ2bEJ+OizRtYdJWL0gsO9hubiwe5OUz7vEgxMsUM/1yObq8j+b
A4BauWhNSHa9J3oqDf9zh5w7xt4CuAxzWD7CYb3C3UFAHK9Xw+SB8by0UkWIla0URBnpLNEPjQzN
l//nr3La3m6kBqCQmwITRQTotHb1thDYt8vPvvxGY1YziORCHASBUPhE3n8I+Rw/IHIKOXp1ORJt
Dw+vzud8ki4BZL+rWUGR5I+uukW70ln6+zDBogq91pKNAGXyqMXgFadLzx+HRGfUuurdE/F1/5Sl
zb5I+dBTxGIQhy/97mrVZhJ/Joi6IaSj7IDXujg3lCfgWRqlDPe8fECmymGI62hNWXG+owru5qTd
45PfQRw8d5cPap8TqXPaWqvFQ3Jz9rh8cnJ6h23CmvQhmEXdZ6TuxaSIxsDkOrP8Kehcfp86wIzs
68FMCGsmAsCHiMEtvHqBt/VdjRtK2ENPLQys/maULfxCx6uU73DNwKzRFyRJFDiDORmOkriSkJNj
tsM6qT2IE85ZsUucqcQHlIHbRKBXGpQMzxRzFptrX50yVv0Bsw18osaKijAWPixEuD+3y9weEC66
jd5jdG9qOrd3dGlfOcEL5C1pxHXgBzQJOtSxDhAzUiF5ee8go8ELfoi79dpQ0dX3D1Nd9W9cdRYt
HjJ93kWgYfiMIdrDVmYHs/4E7EwvSsD5FYkPxalxHu+pW55bOnTicvuEMM3POjBqiyvKX1YU2juQ
vQc4rSSHwQo6F37dYrKuZZD9cGzADYmYPumGVgjMVu+LUqNIPz2t77KSSq0UaU7oiiHEVus+K6kH
1yeba66fstpRO0mzUAM0R4z94RlQAdRi6SZzyO6Nl1LazOHyjcfz8zEiBYdHuvQt7AOIe9XcA/ZE
YtWcEdUWQ0CGRZK5enW5vCg8ZKxKt7fbJVLbU0RCIY9e3+EN4D+S/S3qKykOoF1kO+BFXYkRkS1N
TGzwZVaZYzUxisE/xpU39eBLzZ5Z41YawDtE+REaZ2C1R1e3mt9jF2+9XvJTTqJK/60tEfzg+jEo
a7PYwKR/YagfD/70zv9TWPdAlAA13qlCu97DzIfjTLAry0b2vAa7dNr5k7lQtc2xJwL714DkHKUS
gXF+hbO9H+haNrFMMMKoUNXqniBJQqOGFhnw9gACxc2jli83+ozywNsviLkZO9X04CqSbZVrmpDt
6bROCO9Fjv1GRwaM9Ya/EHyXaRbKJp+yDuhMC9culbj4cpzHPQTH8prcNcajrS563xR+PPlpw11b
egJD4AfwPObTc/ikedLis+REPMtuK7meJpkLsbp+V4PO89uQ5Q0bUeWl627/ANwhkSVCvBFZpaje
mH3oVAdDdTKM1VDRhfqW9NDpde1Z70j9VrnahcnCE75Cv1yppSXy+DcU73KZqmipshfdDkU5ZYKg
xYu/m8qngUztPkM5xYSNnc+OZLHNnxYBPGLC7DSvhVOKMbR5vkmHOqko0VZsUuU7YUJv36Dh356g
enc3UEGhRay3RCfPfTI8KCWYPjKQL7D4LTQD1INRJSpgMmb4PUIv8lizPZBjs3GMoynuliBalGAQ
El1d30EmPZmG9glt1dymUhzrYz4YfJeXrOTJGuA+6QnDclIcgN3bdpXjY2w7ux/YFEOvt2+mRQPt
7heURcPKbCduT96WO2Nan0sfKwfDGaK9MLnwHJxj90EHcL/tQLEsUkLbKukqo7y0EWCfSwJelr9D
dAm+X3ZgtorwqRCnA/M2IBedgjYZQ39Ftqyo8l5jwLvzC6/ua906dlfIdGAfz81yANgdsJ2hWpOQ
zkekr0KWySaEalZ++MMnaoBGQ6i/tVXAK+IfwYAEjX88fXPtEN7IBFW0JZSzKUR7fOGVoEJH9inD
unvbpt7a4py4G2rZ5DrxRVrHUGhmuvPjnh7E53q2k65CRwIlyuFK8ro2NOJNHtNBucS9HQV8+uGU
jh/wXDBL1X0HMweozrkggv8wiODQI6BTkU+gQU1i/QV2JCT6fZoT4+Jih9R5Av/EGgremCJFS2Pe
31DOtsvfzB+jEKmd0uk6fLFUSf1LfWKZ6VopndX05VuTEwtgJEHHcTvQnw8TpszsYNeHWUUffwPc
kjIyxSSBsg8AfEqfYFfWF17heuqT8t0KHX7GK83ekKgxJ1H4bWSyJWTIrj8wDMwhy9d8hBRkvKsL
GdmlQQrSbgXsox7h+/1aAWYXrnMI0mTt77HIsOiV1SwXvwuwmGWE9exGoLBmwEqkzfZ6tZTBNIa9
eOtwzWdD9+emoeMXNotQCj5VvmmwM6eSmWoTY65xe1dCUZ9xHaSOnozUcoTqb+Va8UJx4ss6Ush5
gmrhhmUT/fOgzuNbk4qdkoXKJDmxibTZyfrdYi0TZ63Mo287dhTsCB8qfKHIj5HzbGLCHtNg9TXo
VvimAyVDf6w21K/kE+1IjJ9cBa148pAHFn3elneZYlWMb71/U9M8JsZ0EyApQK5IYojF3QFGjhT9
ZKVXo+nN4yckVs645rY3qo+iRXBG2EgvJlj8IMgVFqenn3XZWjLDRvoRgZlPD/GwHngJb9gN0+jY
5Kfpj6Zgp1+pyjkHbUsezov5CE46oILwubyRcm7ASjhDyEIL9I4cMAbmNWOz5Nnna70CHg8JJt3d
5ipUeq6BPUDS9GDPaXiP32Yt2M+kGOZnP7mWK22UQkEzZAgGvgxzgH/F8MkpLW6B7t54nD+ON5R9
lUExjfsf7hQggqN1iV2V20S2Sx8el3IFMH7G/lNGUpC7V2V3KaOdeR1xuq8ZtreT9dNDTsCnU9xt
yGmM6ZLjb3aYa1d+Z7RJ/n1WyLXw5xv5zEQ7dA91gdx5Pbdmp/1RZoPjmZuhE40jkB8tkT6cu9LT
4+MZieMvj+H+HgXtt53yApb6Ga/ngwEcGY+OMnxTb8R1mshMu2U8KXvgw7syeP43z9iWl5mxdvSb
CbvhrtEo50UrPTkQU5sRKV7lrBHhBnIJ4mXOUxV3C+3Acm6nSvt41TY2eE1zjC+SDHjRfNvlf84t
D7XXN1yFwa3yxKVzxbUzjcnzaRQQRAkCxfZm8XctCqLIoxuzTfZW3pM7tcc2t+mv7hFvxNmI1PkA
xZ8sRHx//jm4xm17y8rf1rCbZ2TmsyvrC0Eo6HfVgMSTHznqz9akMbo477HYjpOR7PNgm8FXQ8hk
xRW4K3b2YJbc9s6K5csCulkVs0V/dVD4avUqBrbYrqrleD70caJlcVzlrA9Pa+hqvADNjflVUeOL
EUDDRASRFnlAp/TkRMo5FuVGhaRiY2Hua9jf8IwkZW37eQ/b0BOJb4MbHcPVMrVrHgH/egOWEwd1
ok3soZqbGA+bP+IYg9/8YWc6JjWGuYjZxzoaIkTHrOjPv7az4CXUgMcvbYU7MvpejtY8CIxNL3Ag
HiL613DjOQdCnAq/n5kucy8duyaHtBkbj7N+LYrC/QiD0MM3a2H016U0lFdLoN7UsLAbxpQ9UH7I
n2wUhtzlMVJtX3INCPyXeDjKR6JCWSE8FCPVElavMwxKmOzs4GoV1BlypcNN4P6/J9ylSFs6LpcY
Cq/QOL7oz8L10+t9QI/iNp1KNNAluParcV3zDNtC9zO2G5X7nRCo9hfrr17sd8GEioeGrIoFXrT1
B737DE4qbfnafTYPyvIQf9gY0JHv/NIBJFjgg9FTK+K3mKijQFLmP7X9GLZo86CHhxFOI1oYkBAj
rRKpTSGJIjmtnhdBGRUM00ASDU/E0wjEtMIGDsLr6GzAFJ5sUTeX10nCqIOqhocdwCvtLljFh8FW
AJHCkOzkqgyahiPWVtyKl62fXZEv+TDp7Wko1WEX2mGcRWEE6AItoYqJkNHIOTmoJd/1H66u0rLA
+XT/1EMjYZPzppkbOQ0aUCH7iKEgXswxcYG3V2EtUM9y9fXvM6s06NYmyw9G8ApX/wyshpGMiZ8i
GrFYu5dq7z/gcTuSaHlAM+yQxPJxKxxEpN8wqE/C6a5722l8fUGswJZjVbxTmgSC8Ynk6cS63JXm
bshy/JKPMa3e67oTqYT/G5wCQxVedkSIX59eqJsTBeBevny8/WfxNAh6638NEo0//HXfnyFTQIZo
3EbjSvPj2h+8SjgfUC02Xq9Slgm4LE+PY25HtRzjYqMCHfQPuWJUvlgUhU2Yk8dEibckoVM3Mat6
idur0A3z6C8gA1IkH/Hoa+CCGQoVe2nSvk900ARskX6rJLC9/JoyPsdZD83HynwAtlMz6gc6Bj9y
jwekPSknC/41rsYVbwTYibtSm+34SLOamLBgtzb8lYx8zsPLRB6ZZMCBkDSGkFTCzvpD1+hmTksu
mquvkIbk/W2PfAh3EL7xJOBa1I4ILSRp0UrHin0HJDYQGjzMfOzHYBKIJGU4MkzNr9MdtR6I6d3d
ZbfBIq+sRzz9RQS8jEICFhL0/OL91RM4UOrQ6mdOfpFayc7IvOJtsydsXeMjckGaNZ+PC94LL4uB
LtsCnh7UTlMkl1Xnm0T2K/s1DHi4086b/wkZckc175Ac6QqH2SV7ZvwcbJTKrmqGrJIBMbm/RDCQ
ltfv7GxcCvOdIuRAhoXwj9gvKSxsEhjUlKfV78fD/FkIoXzT0xrLlWTAJhMXuWSIRHx3zlXNFmZx
o6ULw+JHzMpJeRrm61F06hzOBMTnh4bbGpdc1R/jkYbZ4sXJUrabfZX1uFqy0e2Ea1oPD0FKeO9J
lLRPzFKLlScANyjigtcTnw2vbkUxzp9McgfWnqCm0nf7gGwWAOSFbNZSsScRLpwHBsDJdPSoXyei
NYl1QjlwNjPyGzHGiDzgOvwzNxClCOZvTFHPzv001cWCsrryT4kpFlEuTJeDdDqKqBF7qqvDniNr
3dL62wt88z97sF3Ni3gVxhjSWHmKeiRIGs3qkRzPpguGiOxT9u0dlT1brR96cIlJ1nWWK6TqhPCs
8YfuwL3YqEdkGQnd6cMVrR1ErfZrwFQ1A3PYOiZJ1wFUku5q3094imWEQpFN6pOlbaFhO1PBxSez
qhIkVydtemoYkV7ezRK+9MfklJB28ehjEXk6QkjJQL6KGXQiGWzfbrdRVyFqBgQyPIuQ9V+ZeMZ3
w1nBRadh/F3ufOxc4TE268t0SG7t6FadNj54BCamnKOP1tBQW2BTrTVvEf+GZmJJ7niQzbD7bXYO
VMU+eJf886GPX9Bo57ixNMr43q1vpPUh3WkJFn8BvRJ5r9CAN3iXTPAxcxyxcnxubVptRoyVoFHX
ALHr12kfAf+EGY0v4JV+h4mGCRqaeYeR2AarHVror5ZtpWyHD2/2gGMRJEEKnPqQ/+nLID0K078m
kdhiOIOK2i0JvIPxCh4eztQpWLOp9hCVZpKCsVxaHje8nCWqSRovJsbR7e7h7yHBbpZ4d0bF02SI
cH1KvdOrWNFiwmUSlfWKnBPnImBKkUUtzIbyPlyQsWbVSVMSU5FKEpoOkIsPShZAKM6nDbY724IR
a7FJE2+lCFH66iEF3x2kII+RMYd6mPkDVeg8u44D9kEujtKDRaSq0YmwbFxNoIzJ7+0UWfNur4q0
oLYYgNL7l4IuXTYiR79ethlp2epOLUQaSJ3Ah57UCHspdZ18umu/jqjUHllamEbU0+Qtua70ZIKx
uRXnu/Kjlq1M5b4IP8hqjxbDik6ROKyBpfNYpuelJUp7s1kzua46Y/TG280+9LQeRWk5r80JwaKP
s58SdXiU9HRrwO0X1baDYtiKKcAjKIMIgSmj91RauU/yCcWJ6cBSZdwmQ5dps5DoxXPDbOM0OvfI
DbWXz3ssFgA4O1g9/81oqNCC9eVDuFdvvfS56eHRbWVQG1RfmyWoErnpJQlAwh4UwNIAxeC8BQUd
c+mmx2Kj/38/Z36s5zofHT13GB/tcuR9AURddr9tFk3UI6ZloKRaeL0XbewyFMcCqnGYKHJ6CyMT
ET8h38Ozgwd3Zk7CpDUxv2CZZ9h27HIEmKcaUkfVfo2ZvkiJnU3ZtDMiVpMVQe2JqgfjxawvboE/
sDdv9ZnSJ5apUtnpLCZrgpIr8zwJcoB+vok5jMeRk9EtJNUNyToC5QcK4mgc1vZIcxm0kG/Je3IU
6O3PbpKPzRynz+lhr/mS78eNCJ3d8bIDAKu7Ia5qyXtHPeSwbvNcOzwyHoRyxaYmw2WQaVgL35nr
dy3dKUOuYM2y2F1niyMEN5TSvR9PewL280LFvvhl6A2h3nMhjR/rI9QoXJSNlS0WlBv7qfn8+IA+
FAHiUv+nfmOkI3pW5eWUz5yo9rSsGRjOKDxL5VUuSYzpUIzbcMfGBioIXZ7umUAKrdWZGgSFm/CD
YpBuM7EUMW5FngGD1lQ511TMjlZFVcI+udfPbSeNbE7gXXb+G9LMfDezX2z6gw2PxlYauTRDly5s
TG5liqgND6Uoi+9UhD+lpl0THKIonmvhtNQO32zXDnWH2zh6nRi9NKo0zttj6Vwu4WXYVBD5oUnq
snL7KNvsAFb7Yxv+SZHe6ZkO40N/dxQ4v3SYwpKbQVOWF4KzhAwvpCO9TJO9f4mTLqd+4MM0Wl+q
TQjEEL87NMFQzQimTpiL6Ru+iy67aRl6lueQrFi9tabMWxVC+g5Uxi+OX8a78546WS2KTU2kOt0l
LImgpqDdJgg4Ih89gftNELRAyYU6YkFP9k3QR3MahP1RqLOhfv/sTAi0fu8NZdo4eArVud/Vp82u
iVLhhhA9Z/d/pDY4bnG29piaxpnBYrkftX4lPvcjwNf0u52Yanm6cGCTYgO5ENLptr5BHJIjyB6v
Nb3ekZphnNhdg7yVo318rjtGHw3RF8Y4bPVtPNoIyFdsX8GIah/vnLPpn4paAuu03ZRvb3PIdRY0
xWesWo63kL03e1JTnIK4gRq62kYff0poErRzXVilGu4b0tZfJSmGkFXQ475fLH5Mm9ufZmhjGswC
Y7lkG+wWM8/QAsBpPavmtB6Payiw1xpIADAGzudk22D429lJ2168LH/tRM1RwvG8IUB3niagVZQJ
Xm1Kee3gumKB3QP94EH8LKDw5GMeJXXQ4BYKuJ5nHeDO5tRn8tVggRHpbxx6amSDlrqAYeIK2/AW
QtulZOxkAvwvKd40DjSYnDYHZoPLyL3HvX9I3AevOHBaxgQw73NHvkuyY4+UUJ1RJZ9j7RfwA5Hh
OJx+1KeBuqbxc8NKXoKX5FrYr4GHlTHqpMtRh7hNPK9bgls2lVVRkAlajurcjQL2aAc7Hv4VMxHG
d0Bgg37/3M0Qsuce4nG+X/LwIpR4y2b14vkzEyRJMZPdVZYaLzHuGGiktNm4KjWrLgJKydY/Uxra
u2N19KCG21jg8UY5r407WWPUBBCU9QaY+y+OUqC23ceHRDLAGlfXmtrbZADCyS/xrGxBWCMoxafg
wpep8T6kEcp5k6KRSfYM/opogHlRT0eZ6OyF2WSJeJgaK4Kmbp0NPM5ZQDwgG6IkTso5/TPGHesa
p32aZrfkIXWlQfbqkiydodwtyzjLZTjNRAhxaqVr3jmPUhxAi8tmVFduk/5l1S4cKzdVITfev5U8
GJkucCMR0fUX0rCrkg0yNfFLgsFmpwV+ZOM0mBgiQj1rJQbkuXTa5e/UnMwr58ZeXJ769jskQJKz
Ujgpvdl+L/dp2Lzn7XfYKZQUTpcyGoA9/0P2x2K5wRf0Rh1wShTHCJFOtqNNTgu/JLz2FtSK22Oh
DpgVOdu0YFhapIkFqGlzo35IuIRX2iuO3wG2zyzX3Q8ZfDkeyfFQOMqN0XsY9i1DX8j+XMY5mwbo
QxCMI92u3ExKP4LE1wpRHVG6dBEteXqkz6C8MRT6BEj7BHUjJ8Y6vS+G8o+mmunHWThGDtJQrQEa
qu+rMf8COymTB/GrBRSjKSQoCK6dvlra8d7WQsq6c24frXGe2zYSXDpFCv+edMkW7+cdCAfRatb7
fxc11gxZm17qyxGzWs4QYNt34UdmMBslKnIhOpmah9KUoMD8DNtxHp07oNOxawPec/yG7xQ7a0p9
76VU2LahY71RXwghGqWOrAVmMcQ4UN8qa2DWqGMfRcwDVVM1h68MKBpi0I9dA8Ns1SS80tDJ+JDj
pRKq8YHV9hJWljmZiLof9untvgoFUXfQZcb9U6sl7w6xNCYkmtLZkbOYsa1MOsmK3z1OMcJfQu9l
il6WOMR8sAd01Pv0z95XnI+W/K4c/dlbunBXS3P1Q/HPqD/OU1XxHLeao8Jd/fpQJGrHYoH22A13
DBXdzftr8PT6Oz+gCuGWDt+uEMOO3bG5DXQR2JlW2GXqxDq8TpWNeMwJAoSuv8MXvu1UH2p03qRn
pSG0yPToCTi4wTXVoJiz6TXkZRNdJLrumqv2paBlYAX+0hgEFQmL0Ox8nvYxO13Hqc2ppxfu4n9Z
saZfzjoeVwpOETjHxig1+qAM4mQ3JE1Gt0vA3isqCLGnHm71KRWCDqtxqKpXZSJd6AMSqemTj41U
kB3i1/ho46dUT3kH4v+EedOC9925nJ2E/HY+GSXIzL2FsmUUOzoBVfkIYGq73FbBHIiVdtg1ls0M
pVzh1qT9Rxo8Z2vH+TyXYXKIwZ8lEVMO9vzQNK4+WZ+426riha/psZc8InEckUwigI3tly6mVjMw
o3MqD1gmbuAmF6aD/eDWeE9096KQWImEihAN7FNsEiSCVExTz26e5QEXGjEQh7K6XG8X2bn9buNC
qbgDbDZizLF+VoY5xzcHjdsG/4mdPATDM8FxMLNpPMEkmfZ3+i9UFYzfMdianR2+s5wMpbw8U2Eh
+IplGvK17myX8BSCe76WI3kY0Mk+Gwnx7BeouVGfFbiLVZTQea5riLbAGv1ZCFPSsOQhlB/Jjzkq
qkzzlqPeuXrzhNHjenDGS0neTpaKvLOI3U1FjfeZrO/lCSxoXmZNwV+GwQis831YaGuzYeyzfSdA
nkdh+pdOTx+buV/C5W5jMbM2D0BErKWzsZu9eEwy4vA93Qgi73WElHp3go5B+wRuIRSXsrIN9k4K
xCR5G9wcktsIm0/PS6yu8LKwAt2/wuQM5U7OifpS/sC0T7sNfYAnZ2bTVx/+H5E0mDZKIPpJGzTe
Sh0+O0mjecjuXt9NNulr2KdJCvXuuLOtTF6KqJIo7eATTwU45OXYi3Kijc2B85ZBaWEm0gdCqfA6
Y+HwFdWNjArZMhgu5d5sL6D9Pu2vL0zQLKqm9MlwSiS8AOqMHlxdWsJ1IByYKF2lyDsbY+HV5Nnq
+bC22H5ruMB9taX1iCVZmhbAYpwuJmpP+tsZiTyoqlflV4gnminC0iikL88PxC5Ci7blP/afj6Xz
3Gy0Sinjs6J+erDSmrSSXg6sWmujmk/RIlhMC2bw0PTHdLWATlMejr4+dlLlXYzWuC/EKdzKUbeq
qpqBYV8NEqSA9DI0yRu1SJ02cYqg7Xc4DxVl8as9qCgTc7GHF2EKaYlUvgmM4RAX9mhsHuutF6+p
GWTD0IaXVp0ko43fkEie6cp3OFjpk4HOnyBucY0kq3b5HB3Tm+0ZjQw6vb94CXq7aFY6HXluiwpl
RZCTpgDngBDSXX9T98/STGBPkr/gYls8gYtARuCX5bmy+86+e8O39ljDuue68ojRKMUq8Eqmvjjq
8AcBkMSnIAJR7lCF22gHHRWLyC82NKXoejhXlJ7/0HphHnCQB4E4O/FhtHxoicNORRigR3lKcLnr
7FYe3Z+j0tnPCN2ccMQ+bLPVaX7Knm96zekU7H6kmj4ftIH4X5Ue0PC4LOegx3OTXM0Fn9P+JkrQ
nrgXqQH7VGAh9geIL+XtCqpqxP9VjL0+K4t3/JjyvhZmj6/hBOINMWYerr196+5IZWE1MSkfCJLS
ZK1/mExRUyG3bsJ3ZCBwr0YfOJ2yUkkcZgfUKaWfYAaPwE4y/oWvmOTbShiX8I0TFQwealA2NqoL
ozuBgSiZlivTjCyAvLiVsRzvbbLfLZBsS6raLlyjDpJMtUAZg+GeaZ+Hjscg1zIaOfcksELEGsSd
oX3W8iD3AwjWQYn6cxPVlGL1IICSQ3Rrcxtfs9PPvTolhaktjq645VIOlvvPNE2sJ4M43TAB14aK
nrnNa8hedDcT3WzOpSRq9zYXcOXo/Hk2qIiDhu1JVfzhBrOudUTvejziLAp7ZPZMjNP2SMg1UWhG
hOU9t9JpCweCLjDcXi8zsSC1c843lZWzMm2NXW08XNbjJVClMFhuSMWB2iKBPXGw1Yb5QSZPRSlm
pEHFqu217zlBixp/CkpMwOdmG89LnLjWxLgtWSM14kU6zanA9x0UaahXzVLscjGOqWr++5p/TINZ
br/iu+36Wd1QRwaLSEIrb1dhdmuTPsMnf/15oFIwir223x8F9IM02/QM8NynvQC4GIiYTHykvEq8
Mzl2SYZsNodjU6CdcCLCJFQGQ4AeyeOAOZPC9blqGkfyoL2RvUVb927ES2nh6xZGbwYODcUg7hH/
qAM6o56zbSGB3pdeNewaMvorn1nLXd5NQ0qzkzUKv4ABdhzpmOqfpaYoduyzzL1GIyOLO5R23GHg
aymxKLy30r5GgvkousKK+Ai22GDR5S0lgMcZfqDEfEJ7GBUm+XV4QN3VhlDuww6boocdTNjgDJKu
g/0ssl64jHsOmQdyRdmeDIS/Y45MzHMej/Vn8Wtck+eNHWwXdEEbuyBRTwmRALSn3Z9xN6Rv9IHp
kaowGeIw2oGy5v/OmVn39OTUhS0vPLowhIL8+3l6r+fbUZp2LQYkMlTBiNzw7ZW858ZSK11VthE/
lT93TJ1HKzEcIRm/fkeU8GbS4Z/LQlota96UyGGGGYXksD+Zbfusbut8WJqmpHYqmxGScs9k79p2
0T8Q2N2bXkerTomVhfC/thg7M53kK3VjjOCdqG4O2G01veYA3rxyu6Q3s7tOexUxwUe6T81yz3QU
ltqqgoVM7x8CzwSztbuwCAFFeKbDPp1vHnT4JF6m0U/RjyA2+nQncp4gId+bNEcqTawgz7VnzU7v
hQVsvG9IJr/EIm6WgPBvHrH2bgXlqPYgpE2qCdXBrORslUBGtmGf4TjWP06hDBt4B0GZtSj76uaH
5EUSTcWaepen488OLT04kkz0Wc1748xrqCvz48wRcO2H40Sis0njKmNvJvggiojC5vtCvZCy6leS
L7DZjq2pYdjR8a8qGOkvKiszgSSW9IvegaGrSdzAtK/RIGnNPNIK4FnBZyITp3yjQDpu9MEbyS23
ftdMV1MR1UyUnfVsWKIOB//AL6dpEEs5JTec4cwUQmeoG0nvJeBgPQdcSrSX8hSX+odHQ8hK99A4
mn+FpidzlBrmVCQQty5DTW3EvBoKohFtjkwT3kbSuPP6rwG32gBjjMqBBeWRhELrlH6QZVdxLdnK
kwp+XzhyPnIQOnqmlC9xUjtULantogK1DeQ3mBMmKYpCHCMCGnrDNMA5KQhUtfjbXVtdFErsWYdc
iIh9iGV9QXRbM3KyeEoJJjlbeXFjH0LeBDvB3vSwi0HMWa5SVGAPF5ufSZjEA4zruJZmoc5H7mDr
BS0dOGZM1OEcnEgmh4C2SaX6liiS0sRQYeRkkQzybDjlUqMJ5mPt+2Qb0KlfSAXbZFQmlU2nb2TY
P6DogqDEju/zGFuPq7Zutr2gwg13Z/TLlaRsIeUVztq84gIISfaQ6Wj+x7Ay+J4FprPom6FH143W
RM9BExDUwf+/rn/5BOMTvsOFdQpbkT13kQ0pfjlciBPdWPzGamAvWsJv1hu73uFJxtbKDqW4SEOk
C45sL+1REr/g1V/aJOJXDGm/Wv7LdWJauiDiwFan9SCQe2ZazYiWYdTirVSJdK4kP95EO/3Ltg2h
p9knajU0u/s0jqwlLm4rTMryVmXdkhpdQPMa17j4HsOrfaa30njGFt5q65nYdVhdwaIiAK7sYoVn
v9GzBxmwjFknL+cfwoORzXlgwbR4W6TJIfoqa0a4R7fte86ODUzUA/PT6lYPIpRj3OmqSolEK8zM
acQiOTajkm/nhm89pDug+sbYij1XfBmVfgrlx7w6oShdGpH7aGfkWeAnPD6ZgV1+npzWK1N9nR+I
BMZGLlsvRuDRo/69Pkrhp9jzC71+siT1s75jh8dF4iQZDuajubMYifk/Ct+yIFkm0bon7gYuci+8
31St0n5TGMml6dqSb7OpRoay3QH3xefKRYITxltgUvE2bnMFcDR/O+QwqAj5Ds0DGerBC9HgV4ya
3dwW6QJCAUl5xghPuGckWHbngYCmKPqEnSanlHhrDhfCgaQQaHoirCrWhmhMGGgnaIPCxeasT0bI
oHjs8yFZZ/sJpijOkWRtXArf70zfHcOBi8+MF2qiUv+jlZmPNa71//y9B3QDpeXsXBUp3nPMv30T
1bKottplsS1F9BvXPUUyKHogqEZnVe/cJZVcxo1ty1jb/67uYLB5MenwaLx3UILbwXP66LZBIzjq
+nZs4L40MT+Th/YHSKjjuqOGT2T+0hUwm4ZWOLSXAUKeuGOrFgyO1s3YZpYbAWviJiB2eMSPdFc9
Zk5KSI+OQfjrqYBra635fsf5JLrOi5in6YhKsR4JadRJ4ywsyQF/0zVuUi3+AMPzr3dr3p58cB+M
eCeogvxxM39qjB6lVzJpGUA8lzIrfTLlB+yD7qEs0pToEqW8diIpMSgdMfDRXzdQUiZF8lCAkJfR
RamNAzufvYoeDvgW7LN1jrl35EqABI466Jlh3LdEsV/nj5yIRlvEDDJS6ls7xICOoE+F5I5uyHbS
0DS0OqzNKUyWsyik5SOFwplRRHziXfsWV7iu12bObfZzfNY7+7hUDZdP/qYUuzRaXrm6vFJaYD8v
RShQFM7+Hviybt3D2/uUzhQXb9iAB5HMLATWuXoFd7Ll/9cLAdzuTEV+JBGa9f4ExBEduL3YOk0H
uL2JAQ9YVi8vXrTYWwrmxkSFOc1A3P/iKLsAVdZ9ZAv2A/vSy+a1G2heuZAT9QKQ9dqNUi1m7Fpz
TWfDUGoCxpYjJ71mO8FlRhkUk3r2GDTTVnE7tRbTlGxL8EAMfJhuCuhFBbv/mf3GlR0j8OAcLNBj
0Domh7K1dG49cZKoWJdqfS4f3Y3UgreBcd+0FKddMROPGz5GsE2UvIsKmlyAVoa5C+IC4A4djhB/
rBpusmDW3qp9sdLs+YSY0tRhYxzJ7jOztUNyuXsiSg5nZPm8SjjoxQbXQ5p32e9lsHzG7eLYygva
u/m1yDXdB9DeJHwti8dA2DgSJU/+Mikeu6n6fqS+cSH4sY/nEkJKJfNqzM/ovT0gAJYOYFqHLhW7
8YHlUTldIApMrbJ0r10dNsjU4TIlLEN5lu8Y24/ci0wGEy6Ak5ep97Y1k8ekAuUicI6B+TwzZWEu
UolVqO8tmRP55t0tny8HFklBRduD/swxo/2+JY/TqlGntTp9PaLnSs/oI++/LqMzzEhOgiFlRKsG
ngAzGFaKAkWAEe18krQKbyCmKuVq7eH53/Pzu4R/35c7gUpwMCVX6BuJlS05g8dYpJ5d+Z+oboOj
ofRhV40VdeteS2e3bD6l/N0oeVTe06on42ggUVnNqRjB78C/ezFWAhHmZiPZHvWmiSm8aPhGpzsr
qxI+ICjMNcICvfyffmeB5LlXaVkYZcU5q6wevRnp4bsA87Xxhv38B1NkKSHcmw6gEw3CdhDE/Wtk
UiBoGOIUzMPaQOHTyaZ5MaJJnLsdhvIvzTGJ+Sq5VvabQosSVakYXeKHLXeZUWOAIfzwTGY0xKAN
QZjYtCtxmcOH9avLbMuCJuGUzLHcXZEj5rYhnDRb7oXaz6eHAhuqFRtY22vSMqNNtKHNoUDA2R5m
deqmnKkhVGRylryNo4HNyg5950wCWqK1ejazj1mRzEeUH3NhqFv/QjSo36SU1nxpzW2fRA+Q8o0a
x7LPi2OrQ6z3KqnSh7M2FZX5wIHWmNVnW2WqKT/q9BjH4cFExpeXVMn68LDnJZfC0wzWdtsoSLuT
Xw+7x9TRmk+CcL8rkSS5GNQp6mDRWZqywu0BetfJoEYXT4ZeAt4gE/prdpCFe4mhPlGu6APi8iwa
o54QPantQbRp1EN7xorQ48uY98XbdOHUhzFtc7UegEmd/8O1tPp+dIEhwPJ5VaePwhv++/ZxpSXw
C5pQULYgoIqsg8uxTa1My092TjXTfDRO45ohWvf13XSAszQvHwMedHZZMOO9aOcQiPS8YMtMmRm3
xRjpVZhVRyGN979Og5wqgKLyEhYksLmzRElE1aV4aSOoTptiHyX86b0zZAy9kwDFYGrrQAa6Sno0
Gu7jq6b3gcXiGhPYaCwict9hojWP2U+58LwYAqCRHupHs9iWZVill3kAH5fkuYeP1c5a8xvNln3M
tg30PV0cc6dfKmDlSptnvoKPYztUXnnTqU8+Vqj8QiWDHY4m1DTeZR2QuZZLYWbxtB7xYKMzwftS
elOxeRGJkb4UcQOQ6A9rQrs6o1q0ljQeBVzY/fov61us1sAlqvPsZ2BN1vMdqltOPKVkTatJ5854
n53ACxly4XRjTLM+Vy8rRiF18TKu27XrPGIV4GwmwMBvwvO6sDyehvYqsHQ2Mbc9iUr43JVaw8CU
M21LVq0T1+0iF3vOtS0kwiD+5pmhfCYREaSd/N78mH6Pc5o28Uu4Q4vIp/bg5bC/Ep4znm6dWUS6
E1jDQ49psigpklCsOCOa5zLa9HYqhVI41a4ESc0GoVV3q7sOLdNg4Gvti1aDT+L78WaFcW8i9hQE
iM4e/TMtrOKRGu3EroxuhwlwCDjkolJA4XOdo6tU4Q/i52UW2ooVRkFg7xNroCgvK8FbA42dCvMx
Bt/YXPyT4b31HV+1uy4IYaewEWq04yJabaxPl+LljanWingxohcColypr7wb6L0yoNzcA2H3DygZ
qlT+P4GtzNKYGY1vwsmbHEA6U+dJWxY8TlnRdtf6tpHaL06j9JKqp0iWlzTjTjgBvrFfFqAr2ubr
2bejOE/a4dyo0WpI9qry/ZxmTydDHLErCjuVj+Tk9QtdBtJE2fb07gkX2Vj1EgutHrY6zE5pXS6S
aiRbnXff43zjpa4fS6wy9g0Ntw2N4T56WGDXnyKH7mUJhs2OlEBxpIxYCKREAGqVe9IT6abGsoWl
lqDYB4bmBs3plSF+Pir4IpwfCctIOqViV/nG6MUNOwQxjBYxtmv5WJ4qIjIhMgb9KTNAhmPMn/76
RwT1KNPZlHKqtincZC27iNxv8txsuZ8IE6ALd6geRhTC3vYFYoK9ax+hnstoywJvBmLLzH2Vo5ju
ig5v7N064wuO0We9hzvA4N4egsuw17yP+BHt5nLh4XkQMmv6oZ3ydpTDosHyz4O2XQ7YN+ynzwYA
dgPrYuIy9wQTTwDnDgEPZJbd1zNBsNQs9WbvHTFhK2BIOIO9CBwM2qWoC1FsY7UndWLq8hL6SBDW
wOCluaZG9Aq7WLrPgcOSRtiW6EdO2q05h5GcrQXi1f3jS69zskALfzmlTmysSmq91jbnaFxNk4Ov
8y6KPt5bumth3V+itBRcopf6D4W+bTX/+mweI++1S2hQ0TwtCMPqKYpzIHyWzFLHxJqJWXcaBUzo
uf29jo6eP1q+Zxy7O5+VI192gTAV4JGywjnsDuLcFFGHGYsNWcc5i2E8W+d6nEybyqZXM8ZsnwdY
hE0BT0BwbDEKUMX6zMX474MvliIpbISsTINKS+lW3XcvBfe5+8nzOxmWJBsN6AI2xBPhvouI5er8
2lT2EfQ48zC217lqQMhvT6D0XugJjsEJ6FRoy/SL0J2mtq2CBRlmrykHp6a5j0WNYb2gmVXZX8bR
ksiR2HFukb+fafPBuYl1F9k34pZQM3Buhg9gro20gq3B963Kx/DCl96MxyWCTkG72ai4Muj+wr4b
pVRBC+2sZ7RbVZa2puI/37tccImNqpr1X/49aVWJkO2gxKNjN0hsnMa1IV35V90x0+rRrYZUy1CT
YOeqAjAwFozqaye7pqlOwnUMYDTQ0EaRcI7yDcrhSTy/aowIpgNe0gLntycQbhCPkKUS4ksQKUKw
S87ywwuATepboTXFNN9BehVIRr1GLtCQ2aukA5rCm2+RwPmasT0u9P3xnQYAKeKJt0ID3n8v5k6E
08JQyfHsCVIVvwQypejhv6thIJFVm8W/UkgfRWHc3W0cQzFDiJQoqlPCygsQQDFA32DP9wPMZIDJ
oy0gAcnla707oKAIarUTfltvXHnIYEkZOOrlg78rCjKhLwqiPHHfHUFlOi0/MU1Fj1Gsd4oF3Lt1
z4Wa5qjH5yapyh+S/TwHlz5M/96Q1bjCS1XOGus4rdWSX+SHgt9f1NFTk/pYCr1OCzeSrnFDaVS+
XDWOzP0yiStHm80mgZehSk7lxi01bO59R/4T2fPkwqvTKLnygykhJpoofOSytfSv+xbQKbiJ6N96
oNkY4jlhp9fOPK5BTpejLjPnQKUw0ph3vsgKnLGtbdj+7ciES6XW0+0YjmJoUnHpqlpxvWwYW6tF
Cnhge5CGEoin7S+DAHLpeLXxh6Ddnm6GpJjW9zifbFWTYbV06oFoSBfOWUXg0VCcSQ1wouhF+kgW
pIIQfx1eyWOGy2rRjCpnKdeeA9bDJYuVfo2ZsBZQeDrqkziT0KEHFSPIpHvKo4iM04NZrX6TD41i
fQbool35vsRrwNiA7I5VRotlkzdytKZIh9kE/cjZYcvTdODgPIXkzfPdR22qpxl1lCdoW+9TrXbi
imkgf808UuSr7XluebZ4jSW2yj1/NFJL+N/KtcE9+y42bEju2zBEhstLpQ4ad7gIutID5LrvJ7yp
f5HApUZor0Ca2VNaG419y0qFX5PyPmM7x8Q7mKI666ezBvlfiD6G4C0kZigeaJRcDBqpQb4tPPiF
xtsbLJBwsQguMoGbuaZ1TWz8i88uC2URn/KYuDZP65Q/acti2j8hx7P98V9aJQVYsgTJt3uYnr6q
JrHZiwHYroa7HJ3uzyTaGjIfIJAsHLrgxIfAP4udDslHP9N9yDJgE59oY9S/a6FCgEK4y93t3P5a
ZlgyuRrmV/tDWnok4W5F2Xd9Wd8buDyCmslRoxNgkXYOkQ9wwiJZRaNoURPG/vD6AcZk7hY+kkhZ
vphAV9w3V8Bpv5QMA248pSzls9iYholZCAEIU6I3PrNQT4jTBi2Tu1AEW8Ats1wemELZA2ySUDAg
t+LX2PYBXZLTtICxSx6HtIY2s111gUiij1Goyc7MDdmzxJ/IPreIj7AT8i73xUgpprglqbDZh5Q8
EhPRP3LTlwPEjY44lZmzEjdNiEv1QbuJMJnL1Qpi2FFGuhHPREb4eCsy4ocb9mZN6kvTlkUmL7Iz
d2J3nATdC6AEgF7FHlBHn1w/iQalTFZIbMDCIMt5cNFQZre7vlAwJQIUgXZvVbEzFVoJSSVPNK7l
i/5Ak+9lW2A58FLgREqYTjh4z0tDmBwOyU0l3hV+6lGqNvSXUmUHUyKqazC6MD4T1Bow/miZ2yr9
omk1oZO46GsVbTdJE1+6MOSi3I6Bzs0EfIQq8i9h5b5OsD4pnlVoGkXM8zhZKUrw09uK9ZTpp+lA
Cv73RpURgUx9aH0I0ZYOmsyYZVjMMJ1KU/ZZrjxlmUyB+KehzBgL1Vgp+BSU4YXThGKuDHFCgkGR
zXbsGf9Q/S1RrV54rb/kN6OPiLGlZ/T+QGEPrTgFbFioKgaVGoSdrmiY5uOcWX+3qLqya0gLzoQU
LYz4szKM257wfaiZsfG1xcGs8KnH9iHW01Fz6D3mDwFi1JlBMg5D9MotwiMogXrRIkt269wEcSvp
kl+MxQsxropg/OxRN74aSV9xWAKNUdQJo7aRskY/hJhvidba5/X44nz3aaKhkxSrQVSJW9DrAA5v
HSeELQB8EfVoBt/pVYQYmb0sDLjUJ/HY7bi6rLl9YetkN6/kbxvXv9ZmfQIeKN9krpplN4bvxloT
ImYkIi9s8BqmlldyN6tOcINEGHNMTsByokXiKEBHum9/HUcessFQK3T6mul3X0h/DymQ5fFm44cJ
lWxHE6vv4uWXDWuQ/PjOVl0DfxJndqvFya9YH2kvCWbHxeOkABrera9NFzZIrwHQbdhVy73kPW3P
npEt+PXLd/m9PiQVAdcwfXQew/FaBsOrndLUFePA7zv8sHjQ3xL19UbVWb72xKzJDEbwnrWRD41x
7g9E3ij8lP6OSlwJhbWd6KtXMG2CvoJ1CagflAhqMvpats/7G3JB8rFRMdgS/53ws4EGbjzy5o3M
YJ/7jGUVDLGdO16xJM2mWZRF0/SVnf07ncGTFV/b8/REe5c1RBx0HzCCU4Mq6lKFw73UtlQjIcY7
EzomzbcmHDqyae0OMgTTcggcvZkVdb9SfDiHKd9T9F5HnzsQtTZHRcW5KXc+uykTaRvcrUjo4zvW
JJvXwFS+FrEtWeIzchBr7EytarMuINPGN6qW2eSY4ufW2M4r938oIe2q7gXuEVbrfGDpkEXGTDvK
TtdyLcsHhaID5c7RVSV+aY2jVK1K5l6Um7gM6TceQQ5heUklE58/mv6ERkAd5T7R45dIfQOgUN98
n2C1+n3IofE1eBDNJDtTQkE8hEB6SmvGkP2hmZTJ1G6PsNYZpYyS95wsJA19hnAYaVoMsj+/QBbd
tyE7fj33a0b0jRRKy84xNe0Hct0K+H2qUQLu7lBexo2A1uVL6VopxV5DsK8l9jdFAIx7cNz+68Yf
68VQ+HdRQlj3btim9hFgVYvRtgKuoUwV62x+o1KUiAPHycp+ZqGHN0TTiNaqOcNBEWOelkbaNnzk
U/1AY21V6mto7RKjywVGqzjsiCzQSyd5wuyF0QqXpnm7E56gRq2uSCGtxMKCNejoXv/D2v4Ul/yf
Rtso7YPpOCe1pPMSXCLx/yMhd8VdOOBfdvkfykNRKYPkqv8npLW2wmFszQEaBnq718+aJZbacEn6
ZPU4WNopaInWYk55r0YXYcfzTNYTOHz7mDNj9hKnwx8MtsSXyzMkIgWhE/FUi6504425x0K4TjvQ
9ZXjQKCFDOZqNJMaV6ND4FVKuMfFKuSkUfh/Mad5K5gkDzoyn/jzBXEPafb7w63pMmtfkRvhUqdj
HlW9QAhokueIeehqgwKiBy3mv/iZB7VAxfBg000XQLH9wKalxYlf8mITGsQA9/U8rUszAM3ZWDxw
3FNJ+4/aUKfrakKg8z4DKevw2amBW48rZysSrSSaxDMcfSvj1/okkRoVlnB9gxFttiVeyd0ow7vp
EqR22GwjSU4iYFZglLL8WixRg6fAyyFYIGGjU6A1dJbK6Ayv9fydDcHB4h/EWKvx1rH7wr4+ofs1
19BauIXbWAq+AvfRkI6Ek+fho80WZZF7rqjoYx/pPglIJXdrKcQAvBybuf8yT45uZe43Kbwqya0N
Cm2DOn8mxyyeMWY854rPYglKUZnqfy+wq+a585BB/vKkTlSUjlU51cx4fMlSpD7hTNv7YaFZlcJ7
wI2EB1ik0uPIB1S3FfS4Alkr4DAToPYhpclePRbFLDdjqtMTiAz3nChjHR4XU8aCVK3lHTQrQNEt
ZvhN0zcRtheb7FGOOi22rGliLy8x9kPbgb60odTBQhI2CLEz6tIPaa48jyZQaEOleEqhxJydc9da
zRRcs58KOMpcaLKM5cb/2lDqOtEtb/lfShsJYf7AnSAys1EwSK1RYneWaO6++TwGfTsQneiiYO+A
FVf1id8vTpfbPH8HiobimMX9TMKu/X2kgsibWWUMbVpSBAfryK4FeD1GVoOpvwviRFHORDJ4anoi
d87RFOV5kgl2CFnjpcPHY9UG/QG3R2P4Vy0yP1GHsHucPIJD2TJKY6FZNj5gUh31s+LaAiDIOk/Q
X/ChvrqIJZVO0/hy9OUZidqBW/cEFh2HqlN4zIBd7+E4KzXz4ogsqKMDTa3y0LQUYr9fmADY+16+
V4Gh4bGmtHKrq3x5H5g25JYoWSnNxUtXak7oKjIrmuFMGP26M/riOmhvtCNjfGKRY4gynbkm6oNc
CedtD9ilmGhKjrQc9AlO7OnbZH9e96AZLYCx1t+gr3xOS1Sj+OJoztah5eOt9vr+CVgB5wKYJpl4
JZTllqogXfS7ttqJvsCDVoj6W6Aadz79ALetgUw1UoXYps5mSLUDUkzc2BIQAYa6BR9xxFijSqt0
pO06vOl9lWIvI/C6cD4q0R8qlaeMc5LQL/qANmUtcgM/vJpm5HGr7ebuZDEzQbuvzHDiiklpHRw3
jZmIT6L8q2AflciT7dpEiP+Xx2W2XE5/jLsMO7etX8BXk+bYAbWgBQu6OD1/Dyl+/ngCrOY2VpPX
KDWVKYA0jTrqoPUPCor/iGCnZaxpZIIynVeQvQjfnXwgXqNLVuEmZ/dXT3DywQ4mNI2GUBSt6zaV
Zvermu8SHr/zq0PbuuVEOv11nCLqw/RYPIlQiX3biWueqcLqiUEizLHpoRzdz7uQ5Qhx6Y6BkLaG
VwExOiph1pgEDxIvnED0kVHoooKlIejLcSO3W/HEwAKHqqwV5s/jIi4OmO50uWeR6+ZNUEKWLl0E
cvsfjc6dT/pbS0NwYsvxaIPu5wU9mNASvuwOTBGEXvYe1z5AWUb0iMFQ2+PnoKGEhFreYftYG10y
+AmPv/b8VbIb93R72KqzT4Vj9hKTauybY/OpaCajBRsMLD/nCdi7mF/aMT8UDj58CgbOHOYDAgCv
3t0rjGt8c9gctK4y0sSEc2E2eNJp9IPmRt3FTI3UadgTTH77YzrxD572hSPTqPqZvcl9JZ2NwKgs
2q+Tcan4sVV6qnAszX4sV/P2UVW8+YckkzcO5wWp03juUDylPCPQGhBmrU3o9gSM5E6dhlJ8ekRj
j2VjEf5UPsMyXA47jaDGQhZ9c7/HIYZ/6t/zBw8gk7RFUtIbK5tKgtTgrzmdSahDSDo01DXZjMs8
qQ3Yd9cDHBmXgKUBhgUgCAW5I2+ZVUofPMbnv+1jpXCd7fF9IldC5pW4z7gqzKfJqjBxYFe5zylx
lNvL0b8IdfAtLrY9T58sxGISq123vevk3rOQxZA44fqAt8wKSG3gkO1SyKPud5u0l8Lp3znD6VLA
IM2KBF4G+k8FW2n4/TlGWBQ4aNa1o3avtIZx14NB1TPwMX0EzdLE0jyW4FXOrVFM2aUmDP3KsL44
fK68VL1vEl+fxU3G7i3qYNffwQkPqxkH9WMynuNbuqIXHIhKJBpIcUCSvbGmQ/ys2sddLHCSoDu6
LzV2ksWJlT3xc4Fm45zsYiuBYg5OPWQo93Vvmda0CJTmfO1X/KxvogVKu3IeIKzY3I0DL+k98pHh
a8WGXkOppdmKyQDGmL5rJl4ZeiPfPnlqIY5r4oMxD7QXBJJyclhBkagkj2CukUJ23Ih2zS7XlOqs
CPHsNFmt7CuLHHf1f0O4vDR3sI6i1IOmim+rsB+a4x2fwdsCOyv3LycFg2Knvt7B7tSPA3s5blpT
oDO+GOVOMf1e3xLWGHROJ0Z4PTDp7FCXSx6JYBqRSLA3EAMQI5nmrU4OVuxi7IMWk5ndGyrmZNIV
tH7Kl8MnOoJ/DDxdWXlzXBnO+xoFto/WvX0/vN1AvsQ0gwjMjYbzSps95irVL7c+NZbn2sWTFvWI
4SCcBSwqKV1ervAgWSXNEmAWe/WDr7IBGdxHsgC8jl97bXXUv8Xq8G5IVSRpEuRASB6y/dgmQ7Xy
N9qEU5QFp6WTJ/aEJW9ns4UJU6l+x+tC3yV5LwUMGULtT/DTny54I3kfYcwN/pQcl1fbX2GSjyRE
Lk4xP6owikFZADx3Oa1eF7q0DB9qbIQzgH65ylew/jaRi4Kbtb3MJbm5+Qx9CjBRK+MZeTeHpkiy
tVgvzFIRYgJJTIUm12VsPZaipdYKJgH9YWTYYOAtEdnEMbgfYcfD16vek0/neQkJtFop5d0LpcGm
3y7ZKFuj4PNcB/hOpaH+RUia/sHvnTF6A0q51ORfMW2ijNBGL0UOtB3MyT95wm1ThwAiZQK8fCg+
ztW3g5LD74uqKGPFhnn5rM5A3zB+XR8KiiUWKGu2MzpBoHVxzMbrGtFowm1KpRhbCW/n83BsdpB8
cIB94wIxZVpnEOnJsTsXxpwR9op6I1FlpQlUZdb3laCn2RYGm/Etqr6dWnvtDn+dWMFHK80ZWLRN
MylSPJ2EmDeR36L9Yiu+wlLrzWg/mcoEUW3H9huGUg1/zUTb56sMN9yFMiJHEK348uwM074Bt6px
OjVOUofbjW8hUxzohuUjH+L3Ngqz15zd3PCva9UDGoxjN7GJyuIcaK4gdZ+60iW4jr79edQhhJRY
Tv9pIwQ+3ULu2xJxMVqjWqX/jKNlaMPgexUplDB5WErohdW8KoTzAgaIYeGN8G3uyZ2fDqSnq2Up
GeGObi1Mr9F7/YblMi2l31jmhEqGXaf/Xoc9WCbcnEyjHvM6y4oDsnR+geZKINtyY7nBzkQzAQKe
un7geLciEYj0hyxDyF2XFYGp1EpiePJemhkqB75PfDp01xZnxdvNish7CzBWzN5uCJC+A947HNp0
so9zStcZeduI29+pUHMf1FQ2YLO22SAE2JxKnn+sWW8q31dl9H8SLRYDfk63+OHioL7iaObtOYuU
xnhmpmMH64TfnwvD3VGAly0Bav/9JNvec9DH2QzgCRuI85WnaRVccbRFXBfsvWQgjoDHvuCLb/hV
qhgZ3RdYg7OAQ2CP20KhC+p+kOnpubPHroDRoiBEghDtyaH2ZF3w8+y1jwFpTQmPA8Ev++xR7fuu
nLsDdGL39DeHuamrUtuHtMW7wGYsMvbpFCooodaLSYl5QdhmOfCArHCUvf/GG5sHNWB/fb2TNt+f
iIGUTav3gn11sCS6r+PQKCmLyfH9x6XXNhMXSTpdIhHa6eTTkedavzNUSEy/ZMbZ/Se/kHPgABNE
ljz0Fu76zfyoUcI/ortbrISGAQae7uWUJvQEcgDeBF4AmeB/GRFIpFiClcq6F51GLB24PpYNA2s8
T5RyOdDSVadXwouWKzpvZx0QH1e0fsFg5mxHHXuhN/nXp6boHwrxyrAV7ll8LpB0kEKAgYL0i4Xg
lYhKZfs+IIO7crUUgQYQdPYvJIhGbJwig1xVrRFHK3e2BDTFAOgbFAr5p7oui6f8A2cIFXcHj5/j
9UsTE0Rz9NEQJZKKm01FfT+TaxtLw3ZCLXi2vvZqpwKNoMLdNbuWe3YxPp/ASAJIpvJ1gRSCjGpB
8gg//Qj9DAFzCoeuh2O5cfc1buUKcXI60nh9Sz7TpfhidJJwTRQYNKzXjE21S73snBuH3wAjdln6
Co+ZWj+3rDHkmigYMvMPFAJ6UEsqcQ1rmL7DOPk6vcs3Cx3aY0St0UmrzsJgsX+8brj0GiHF5xor
I27OYLQdbLni+B2Qa6KU1/4zfgEbOvDt/6S+kwR/H4tRqyAX2bzKszcQnvx/G+jjTltOmyHAijCL
qHQkAMmS3OtO9/hHWZLTtM13UQu2pAovy72WYqzcjbRSw1UyqZTa2ILn4bJ70w1LGhtUpkvhLZAm
HBcjkvx0w25dByzXMYz2OtPF7TEoOLgd4BrGiZRbN+HEK1La/ynINPxz9UrekwM0OzhnMm9pv7kZ
r1Cir+AvDI5ee3bHaAKleY43iC4jX2d7nh1HOAqVEYY/JwJgX8w+ign4RwEg/nkoofGRPtfaZ+P/
HICu+r75eSKgphOU9Sdc3nn7MCzW94EF0yOF4jPVWIlUbDu0271vRT+CJOhjstOQ84EGJaZGaQnU
k8lsfaAp8veIVrrsZD4MaMiwtypnVlL8eGIzPy0+6vWzZdrgEI156bMNYFvbUwUgWXk7RnnsCllK
gM49jTEFuh8aCLvVfWFqs5W4G+UQNtjX9d0/MljL5e66d0Ft8A8aAo2BSRdBbrQ4Fp6THu6dSWon
gLU0cPNQDgVNpmohrTCn+JqZgEZMmzPqY1R/eWYm1ETdjM5JKZJS7WKHVzDpeRfckh96ioXlXGcK
pxYVNTKVgMJzrb7T1CFyKLZrcTwa0xGRSZxd2GbfsYSIp5tlPDIUVCnzImgxz/TNFBlvNEIjmYkE
Su2/6BLV6O40javCvKIgc8MpMia9vBDpkJV8SRqCdb+ldzBYJ9f7V2SLXNK3ptf5PPVl++TrUc6N
aAWFZbev4ZonGWiKESqnWOWfsk5ThFDZib1z2+fvQuSwFBaxgRSpyR1yple0PceRpVw2zFiEPP4Y
csxV36vmlxCquRJj7ijdkC/8S7JBXVTJIn0NWykoGzLk1ui9Qx6HuOneHGjgJQyI1EU2syBFWvik
aESFFx0hpWd0TAJiz0VRIROjVSgH6JpLv97GIZbuqYBIL32254HrFsxq9DII5kJOfjX0WL19RuAj
C4FFGnsyPTIjwpShzVNI/r6bY0eulmSBMKzFsGjuLp0XFI7KmIJKJc1T02ev9bWGn1ujp3RDyfNR
eURKIN9YbUJhv8GyRSNDuX7tNg4BlPIOMm/SE75ViWibjJLIjDhFXBjitoNJXnnbyAIvl7OwGJem
AJM/aD9KZxhrx56OHm5UstS84NUIYe3VBnoN/FLOKIt8rY7NyP4toFWflkKKmi0Z9m7b06x0DfN6
7q1BT9xYjgY7TBXXh4XLcMXi7aa0NN2SW7FvzfJ3EEFfIKzn58uH+dutnEDQybjSlh4ruMggHe8M
o0zHV3ae8IoHo3+5oFbBWwMHE3pn6kMINh+VymtzBU63vvz6+PY55RDT/j0Alw70C9cjC9EFeBmR
Wqon4mFvMsXQAILRH7HC2IcJHhiHUogNibK11/Ovg0y9g+o9KozL1y/3TLjfTn4AXufjC8qLYFr6
2mCFmnFdMvs5aGFfkscTlDQGfRZOc/6hoGTtCPXd7w+Ab7XbDq4usq9Zr7qZpwwqXrP2yh+IkmQ7
m+lvPPq4IHJxdUuEVVLhLW6dxJPU70E0Oee+iqRE4rnJMdojxbc7xEZygn4+I/xHRXN8EVXsEWWv
lsfRs6UJCY74r9nn+DkVBXCx5VB511wxbyBtmxKdjbjIfe/36sSFbKsKfkPywEYeGZii8EgySv/q
NO47bE9eZg/HIB9z1BFx1SEZcbBwdC6GyNookuXs+VPHk/3JiUCmSFpnioF4D85sDOV/3bGpY1/J
aqnZi5zL539Zassiz2Fy3FTM3WCfDOAAdMeUBtqd9inIUeoOS+j65ReB8o874cAuiRgNd9PnOHbi
lWeqIVmKROVbAqSG+rQq+MwqhOBpBrQlqM70sG4rJNqAFA70fomtQrooZTijfHULynoNhlbhp6Yo
chGdEoepSIwF6BHR6VSjNd6fyRB6kOuibNBgn4v8v46kgswlU98hncRN6MYJzsxQuT8dZh+EfplJ
tHM9GAjgVDjnYxE1OvKCoup8HRBhRhkcALnnxIlLEiQGy9OC4K462tNMbnt6b3uTA/nAui84Lc4I
9TGIgPFMx6VJR0FQKbVNdCGnrUTsGwcFXxtUzWlWpSnp6TmCtvxBhqEJTAZ3bx476JtwgWfUME8o
GU9a31qkgSYNde/0pl2x27XrmgBIceFh5v1NJFxSCBHbYwjONAprl86n1KJWKk0m7LuTbE8W31Mp
P6N/ArvIYZ7S9/vyRfV30BOGovkL9gMMS5Vvkph8ux32BohQjn6bgNSJj2k6QRTwgrx9thPuuFG0
LDU5SkXZ+Ro8lA7IdpeuQ96ca8EYkYtfUQSWP2Xw8QVTxxRaQwXCVPp+N3jx3Ys4c7aFpzEIKl3k
hkCUSHCvv54o6oHGO5LaqYD3rNPbOuN60zZ1QU+FUpDrpxpHYCQFI4jhPzNb/ZjmixmTmxZy1Qpo
vqrj0mgHsn95VuUvmZfYmFf1C4uakHrAE2ODP6d3cqnnYcqyBN0ku47/XBhO/C9qkmkAJzD9DmRR
LbmmTf8SgBtWokFI2staFwMDQ7lJBqT5mQjAvV6nK3pmLd3jdjcX8FSnRiCR9jrW/Z/DSlHc/wVo
fuwSzXNGW4gIBNuQvij40J0aUbhUNrMTvGLFOelsAxexrGHKbQrvo1L879B00vDmnEZTP55hVx/q
fB1wOzJJnHhBQEbB03+d2yLwy4/iPn70vtIiBahShACmPpsoUeQdQ37HBNuYMxG5OCFXDr2SSdMB
OWwjKP7cQcQlOmm/fMX6Al/U8vZC6Sw/rnQus750HCKJIZI7ZapG0ntbayL6BdQilco6YaHdQPvx
TiR8KDCE3rUXYLFFr6KqsiiY1um7ShsNAjIsjSjQuYYgrgSvsZr8ymvh0I98ioYJp0L4nuaZ39Cn
zIMP57kef+W8M2nKCiVTOx8u1UetKxa9Nu9RGiU2wKiXhXTgwy80hogxUPdEy/mfB0itRhoNlajX
GTVTr8eBgquJPKASc+q9hfTN4spk5Cibw+qsrMHz6osY4RpAwh4FQVpz929OQb2dXvDQlxduNIjZ
wYQU+5fdbQZLknd/oQhkSQKpDJK48Oa1gPj8vFkl7DR2/VYpQyQyVqkMX+Lu0cfCHQB3Ma3Zx0UN
DoDFFYmcuvSxKNHhIKYOWagEVHRgMXQtP2/AUda5cr+2MMJAd8m3Xg0FZf44QD0kMXB+vlLIxd5+
B5Xdw/F+RxghQV3h9z+B8j2VZxM0pPYXG8PpnixOndhlqbyYomDTt1OWyZhnOwTjMHe+0DLB08ms
HbD0G0+Imson6BwtKl70xUk7FTVCLQwlNbV3ga19xcBgYVH8hvTjhZFPU8lFWZWnmGTuk/Qji7SF
BbzLFMJTJyGTT7AU/sMGxZRQNGndzr+QzOQtnzvFbvGgemzSSWB7WpW5EQnz4ffpB13yYIlQtPGj
u8+0uNhJfyFRBIkxzmBiAO+udi+x3QeV5T2DwSlhX49A2S+MTiolnUTBwmYbQtewUzLWImwSqT3y
MtHTNVctypQvIXCMsv4b+nxQyUoK+Hx7HWazOOVV78SaiXUCCSFrm6Ag/ezSS3jQXL32sZOIxD8C
puL2HXEjEKKKGl7dkLAbCGPvMneWP4hD4H4xfjhZyCsckGxz+j5V/LVTSdEiiBU0fF6JWefAAq/7
qdynNPzSwuBlk4HTxMs9NLzEwb0oVPe617T/JkWf0S9VPeO9oOGqWoen+S54UjxmYZKyRNe2umVR
IYZTMd/NAS4d9Alv0W55jhb+WWzFMT1dKLLmjTFA4L9I8785kJxNEQikFmah/v1okIsu2bWo2cMZ
Jz8ArXxSQIajhZcbgc+LXl9/G37JLfSngH4nhlkNZmKD6wXw5A6mD2Oyt1PBDWBJMhtQOpOTFwJV
6RxJPQGOVz2r6mglds69K5UBAXnV3SsSkYCM6xdqEdPMHnbhZ9n/vnDlW/ZnWI4mdq7HRnHbVMa/
Kyzp+Bv1NYtSs2oTCw8yj+A/myrXQMTcWkyxVmANRVkK6BGWQzWmNGGxso6dJrEZZ+ZYjK2y6wY2
EFtDurhiBNJ1flKeqSD4LR/IfORuKvxizPAhAg2223LKDLwX3jCAhGAfy8aSfxYvQmF+wmWjcyp6
tZzyLGA33tGeVNNHac9Pxn1DHv6D+nzc2yg6RndKjYZ5+xNESEj9MFUgw6omwWKWHrUfmWV3iuiC
0Cw2ORZBVcwc8K0rzELZE7Ouogyd4DNlxdblXIcmilWkFLwmWlJt6KIkd5sfjzCbXsf5XSEsbHBo
fv078r+pce3WjIunHSvmUsdZfpj5Hh/+K6U0fq3NruSZVfpIDOKsGZhPM4trUC7HWhRWhXjEp/zc
cVplPlcnqoVb4Egg1+ejTp3PCXWfaRAHMh4OSAf/muRrvUZkCg6tQz1CS0QOmQf3+hHYqK139/Uq
d9dRIJxHP8gxcqCuF5Z+G5l+kbjznvjKjTVtLJKu7bFezvCClHOMCcjDuBGxLrasxjED3NLh1fhX
jyoyvgqnIxN5F7KK+FYwUZ8vRiTlHHhrVVj0EepmIaMKHBJmcgGGVTUMa23rWoaVCsafZ/qYdkcY
5Lvq55+HikQZ8Ukpz7DdqqVe69iMqhJ+YzrSD7odTmSEpwyG8yzu7dzHX7iHuZ4zwqmHAUWaOZ5L
CBDtrmXhOt0Hs0AsIWPL5A5bMp54xgEEDYzWw+J00hHpoSd6Y1NtHjvbnJR7af/mQBU1GSMOn7Zd
z60X2k4qEOtJ7W4Cj/WfOMQNpKwdugZzuJEjR5oX5G6lxi9rKgLop1bf11bwLLm8tB7BEIaptInA
4pXBFo42u4VttpIBGh51OvoNJYaZgtMwt7kqw6zGrWWSEVnrZ9Id7ID7eknsZS7gwL/EiyxZEHyO
PlDBuDVbVJFJfQbBN9DKyX6+2MfQhrPyPmKXR8Q32gd3RNrLowTGxM98B80Y6wcT36R1dVPPjasN
MRvDmD4Y1/6sxwM1mZfj2MvHfzR6aWKds4puGScbY1gXDGgktC81IkjSJBFnRN1yL0qaIkgj8A+I
F8L/x6MNPjj2wOZ/uN9W9K/UPL+cTxvdtyd6F7jWXDPer8DtRPRxbjXv+IpYuaEyISFVaDE96LOT
ZD1hCfR4DAdf+WUNUcogFIRM1fYyhO508eS6x0p41uRqN48TZmli7KPmELLaKYJX+0Bdkd0He/0N
nUJAmbh/tsjJ5C3BSt1GKhKE0UbZ4Eha5/6QkUvabbKfS1OKfmnJ4PI+Itwv2bufGvB+bUYbV6XZ
Tk8J4kk9sv76qHoHN5AIvLWb9mNLSMa30XVyfxFFPwWDvWRYJtLI5o1k5pXTscADRHtZggX8v/ev
TD8wA2PsLrYQsqxrKVgygrJjgckN3+sAEtzWKjcbUwHgVPICv3jgWxgI5fFgmykhilWvPbM/7j39
BBn0uIAa78iaNv3ticKSOkA2VKv6HuSo1LeoMhq7bCCXCC/EgYtvNVuhXVC76Mii7kMAxV5teU5z
iIQJhGI1Qp65k6vIT6yk/JmdTIYodMcrBY2uDiOkABkVGfPA2VC53WECyS5jsjU7H2UWy7r/ybjB
11X7IJuNwT4IcmYWTXjPw1T6RkMrwwcFRQmnPxXOhhvEX46zRYyKfnjM44orNhYHTmI/BCLwzz+h
YwzvINAU6kP4zlsxLQP1nCHMSJRBph3xf3+wHdQ729rKzNVkk6EUmAPTuKPrjnPzQnXQo6z2gyfv
f55WzRAfgsU2y25j6wqUIOi/IRKZpwBi4rp7k61JrsmOMv2vFtlgOvuodQJLDFkM64jafHQjbx/q
D/cuRfjr1oHL5uOU2kbd7CU9BAPkJjF4jDMtP1hKLdBjSB2eTTUV/SNqbf+TVofKIJYFjkDzDxwx
Moz9n61XYzP0ztFyLbaQAcSccNBhxPo1kXuV9kenzom1Lg3U/4SGu+enqwd237hru6G6w33mdhmz
7t0g/vu1DNwJqQet2fQszaM8OsHof/nu2BZv5LifEqdYRiFrnxnAp19g+CrwWq1kg/eV5g+7Ag+D
wVC0TDCFFlMO5T3CkLC1dNLiLc1LAoolQkf1t+DQ9tcKlE+O9yUyvX8vswV8+BcUmw6S5Wy9cxsw
o9NNRsdisPrNMhzvI3Oekj/Z8OiFk+VNXsL5VF0be38h1HHwF9/ujdScaeVvKjO5ML4/wkPGhAdF
QknXleI3jo51nrjKjv9lSfR/zygC8fKAq9MV6nZXDZzN4B+zwPZHUXfRMemV/ZjUI2j9ezX34OgS
2wB/rfyPXdr2mJYlqaea2Usq/pMAXFSc/UVwgLBdTk5hMHDTwesPhbPyqRHo1+6KalTWI4/EF/Hb
NmwcSk7zCeATkES8Qet/szaUf6cVRT/jC72DCxIK90bayEsTAs+NGiUmvCV2AR5/b0ZIgD+cb4Sg
mHXX19Ui0cCeHYqJJ548JzDHhMRrl6tTGIlmj4VXczRsozHMru8CjFVrN4cCozw88hXUHXIYBqA7
rZG0uzc2e6DeK3ghqWDtHeAaWllCLoo9Rbz/rXqboa/2/0IJDpGJESNY+UaXGg1OZdv0IxsJPVFC
leI0aKIzLFN7TPjv4Td+jV7/Cfh1O226cHGFpYMDs02HgICPh4fLLdjWPoOAjB2UD0TIHn1786gb
BBkcZ/54lr4/iLmcV9nhNXMZn6LwOUSGF8rF7Mtru1cxZMDlqbdy5lufJbWlee+V1zeQuqpUB0sR
072ZfUSRQXqerDPDbJc5qRF083e/ZNSW1XL6wvjB4rPv8/P4OqnS9ZOE47Gqd8XzPhuO89hcuU9k
UNrbjbfFA6wSNQEe9rFEuFFHEp4ORH+qgmG32jv2D7qWdEKi5KOoTP0QgK01mrnYcFYtsKz082FR
eSFdzcB/LP10v12f2Ar+66FWTZbklWY8B3HExkumG6tK3LVEhvwbUMJmAgiokCJ0bt4Xf2WFwBYB
oLmkaPcVt2Ix1ydQ4xrbwyb/8MPtLX6y0AVttfP05c1hFmwvxpM+dXV8stm4C9HWY4l5e8wAIGdG
v+MLwidnybxx+qBQvSJuTAkrgwGAZB7TPn+zh4DAl3aItoMJ90xobgmSy+n8iuwAvShpqxm0ItYN
NLxNdAHTs+4jgJq2vtHb5JhDtC3MFnJ0dSv1JtIUuBIDCvwIz+5+H25vN81Oas6SmX+g3PIeWdLF
tFVcdimtn1A6eyz2eQ6AnHCruod4ztTbsnwCTX4D6GDjLq+C0xJsW9xnPNYotYIdxDi7V0kUgq2Q
oiv++2zA0PcvvWhAMNkbz6fBgZoinYa0feKJnTYhNwUfyYF6KOxTbUS9RxSZKHWUdXw2C6s0Gbsy
M3c0jekd5Uv+mCvNao0XmGHpSwXv0rRwWTCJbxUCXCLgU3FuNDfi4nnTf3OOw7gPVBzy1wJ6jCvc
rlcBv/FSsE83Y3kJNJgO0/b4h+WQgpLI9zT869nvy4+4AohXIXWDMD7qhACcEdvmAOjbJ1cAEngR
96A05KBm4t16imbljedIpLUKuafouCVEP6MbPBtZIu25SHdSr2FfQ/JYfMW8bfcMahfNFmJWBxey
i2ipDNpi9kgckat00NI7dH7BqkJ87GdQlIyvFzvvv1HLGm+NvIomS+1foeaASg/FK/d6LdlIPNNg
CSUDYaMdoCLWqXDzn4JV7c9S+cqW5ZjBilrxR61WYsCWlOgcdtT1pQ2LntYhopCq94sjVy7YxKsu
wSJEQvmsb8gOd3bfeevAB+yRcUOu4rE1sZ43WaHB0rADU9bRzxS+6ufEINYvudws64Hr1Xf7lyof
BKDJtTt6c5a8qYKaVTTcrfl1DEs1fUXB9YkhkdTk7KP5R+ECNpc7Qw4zRxaEbP7ChpbwuvrqQ6y+
b8AweKXZJY2XLntZoaDwAw3R2rBZ2MJQHe2zmvmcB/m+xXoYhlJAwjEHsKhYhK3EiKQUnwADsDEF
uhNQKyNNRdLEx+jM5mQOPCKzRKHJ/YiHC1hxfeWEYMxIOMduE6Wa3kjbW+CIrQ0PUH+L7j+9yWCl
352Wn2vU0RgKu0stituGF8NVRNT1OI0RDJftgT2ZDHb8UszZnVq59AcPj+WwB63QXg7tZbTlULP+
wLhR4tMUGFnu7kMAIjVvV3oJj+MNBZ8RDVz/pg+BIYhQP63usF/Q3/4y5htAcv37BpdIXhrqUKTW
RF1/bkThHkNmGlbgHLSH8maB+GAow7Ozyvyh7sqjALGBi6bZReIEzGyit+B/v+mPMCx5j5xa0yPa
luBharB0TWO1YmrOyKYTsotqxaS6uSW/QMEG4hB553HszyVvnKTFdhaq077jcLFtWkTI/0JE9G/C
uThwIDJSzvMnub+FB1kz3Sr06bgR5Dn/CEdnFarr2w3iiiSiTTbIJ0sUD2CbAP/IMkTT0MHhecKq
GlpzbX3RTiZb7nO9YZxaifzAOLHRXCDTQLA6y6DfJA+Uu6CVkkG/7LmndqmxWSquoAfJ/+viku+i
2hawdztnLnLZtq6ys9IBYVwg/uMhSxT3qQRflFMFEPgC/UivB9Y9xU9OGVCxj+E/vQSWafBtZM65
cm1+5gejXZ8QQOs5xXpl2YnDclAfL/DUDjB8HKDLM3j4BMcL0jjc+8oKFsKiwbqR0HGX0Rsvtv35
1UBWq/kgHiX7ILovP/3o6/RX7SRJ7pal1hqAKHHUsh4tw2GpypnpkOYuPR4n7dzQKS653SHDF1QA
sUiUQ8HUo/qOxzVdh9zvhpf745jcO9egB9rzwqJIcFNzz79qgitHO7zhPR4CRWArPnCkwCfC1/hZ
bSEBt2/ny1kZcH2kKt7GYBvPeqdzod6Ja0jUxxfVaRYcUUoKyYpF+ZQ1NpN5i6YxNGmL68Zbiut5
1m+cgAzUb3WXSl5PSVmJDPkPzvfVyTQau6QERn/I7twWGlUiXcnPnrzNC4R2jqMB+n5gv+38mXbZ
HlAh0BbvsfBySVJW+0x/YRgYzhIXTiosuY5QtdAUJelzJOqtSzbnaebeXQKWiviVnydgD0suQUDy
oiov6m5z1QO2e+qrjDZvX2ae33THDK1cl0Reu9Qt2hMz/lhfcDby5tyzRI7jXGOC2rOrAy3zvNnl
oikARZ57YL08unokKAQfZrAiLYrN5Fz2XACNg0PLR/cCjSLdkWxXaQ2FduYByyXuYc46C/9oom5L
99QCnmzRzD4RcfRTsK8A3h82YlPrj0DrngzcfvZbfuatVotbLjYLebYr2MDL026dH0tWyYBxMg00
TBA51Q1nXyl5BX7zJNwQ0h0509ijiCcfIuJBIlcZbzvNMdBmIeH8kL8xMFriT/yphFTWMWG2SYJI
iGZ4yggsnkaJU7hMAZ9NG1eRfdSD8th0iagOq6XofgELh1qs1S+Ks/QioQK6pWMh4DV8HO03BKFf
LCQwe0srckYuT+yNadhHvgMpUItJMMuaGjdtxGPxJPNKUsL83cBZr+AjFuc94cwDhfozjDNuXYVu
YZeWZhldtBW/eCNs+GudybkIdIcbWGrWiKQKz4jY8QhXffr/GXrEEoR3fEdUMwA+HZ0liG5V/jB5
w2vOVioN9YExnPfVcq/JsccEb38Z7QlCIpXh+3Tlnpgsfqk1ykHjk5RUTwvs0MeWHPFukZKfRSDD
ZOpX7DI8G2igQq218i1xvHOItydFIPB5NqHIaBT7Wf1w9L+Yl3FXzrRThuA2++MqzWwatXxBnAws
ToN16IXdN4NQpEtJ7fojm/wziLoz6KnnsvTWOGfI4Knv4ikxUVJ4CBQjqEAWayN0g3/64KBAxnI/
y3xPiXsfyYqh9ifo/R4DmfMYr5n50rD1FdOsozOShFBgI1jCclxC1aIu88EMBZaM/uxJDwgWaHPm
1JEXn/1fvMcp82mBxVmX41raGHG/5eZuwK1NojvLjuNRC5tP5aDjB8Nq9ZoFX1klOdLt71NkJ55N
w9mPd2tXvY+gesHYPT9jm15wB33e1TBxsrf1RymYFjVknC/l3YRJjtJXgYeYsYpHErIkUR0VWrYQ
nSAkZR1aEofh5Gt/vDZebta+aNbZZtooBvsSztnOlyxn7YzA2voE/zspV2gXYKkI0aLEm1x14mCe
5F7V2YyHaFteJLGPRocNwEfj8jC45lVzCM86lPSTp1PdUUKFMFbdmaEMKanXAsqRfh8sgTNBuRxa
oPk8dy2DoIdD5Dv5lrb4UhqSJ0XVP7H51HeFMinHyzBk6s28h1RpORYFfNKMcwEJd0c2gm/99Vnw
Agweb1hmWiqSffoccpKjCjivtNV8Ts7s6jY8BgRKcTn9rCnS/4OxSm6vYijSMn5phQjQGbN+J79T
4EvjfiX9KlFSUoL5uQ9yyvaPxucSOElEG8KH2u3515Mb7nSpSQ1Svdd2bXyhiZjPvt11ZKNc7Q1+
jP2UT1FbriczsSVq7PKw2872Em0RG7Mg70xMn4Ol9zpyqnAvDXM7hkD9euhCDgy7kLrGZkNtZPe+
Klt2SMqH45Dh5rJ3GJAx3xIzoG0ON+Rnb11tUvwuX38GT8j0FqbUjYHhgQNb4vxIVyd499S8w9F7
DYOGikRLLRUaB8SniAIVIaeGuLcNXZ6CbkmwBQjDRmNI4xTYEaCU/urh9SNhC0X/bK6ysom0hLoI
yWbI+aTNbeJg50hWhD6kCAl3Wj7LMWfW/r966cS4jexLB3Fgy375SuDJ1OtbK2OYqMIoaUSjIAC/
ZrbT3bQjX2KF67gW43h6vhPOaL6UGesojWh899F78+ZgzIu1MJNrT+mUKKONiQDI2CIlS9MXbXhV
st1bryrfNGtJKR6hGc48qBRu81DRd9VAYmfmw5rXH6eixXg6btIj+7ngswBqNEjncbjELbwpSzlh
0VUktTzbRkT998DqaJIvnnFl1jERCoR3rNUEGob2+EEsQhz9Rg/piPo5RNCG767tGN69Dc8fj7j3
8kSjuniKj6OdbylVjoGXO6dRYDB4ZfweerWucl4U23ESnYfWWFhd4KCcBwmVh5ApQ7bvT9DXbGc8
tuoWZv2sh/IZvFkagda6mOpnEzGaRb1EbV6d5+M6rcvjWMXlZNKRAuO8wnzZ2jdtBas7ENnyAry+
FbpecvVK7vy0SlaH4CXjkLaxq4V2AcKY0mdhaazoDFNa5AgKG4BCfRqSi1wdWlp8kyU/m4ZkW0cC
j/Kda3ZJjrdqWAYk8W+zH/5OHMwNpyrv28dGVhNd1fQERNAlzGY0/6B9UFwUlUidG/6vepQhXdHX
qBtV6KaMIo3vbbmV+YcQjgv8qka9QGqbSAyQOlgcyfSXvpqdTe4fde4IO2wZ572g7i4KSfBginvv
u8tF4WuMSFZvg+W6BWfLryGwdlbcuYqgv6+vUb6+KmIydaq6/RV1+VLU4+QzR5IvtsNkmtN5nCWa
xXZrG72CwIUuUpdSJOYIZQu67Bd7ODx/TIucUR03sVveAhuvfdMRd3MZuelt6xde00gJ8arTbuXp
4mzBJPLWPmldTjErKbpeSTfcPpWHtmvK0YNNQGT/vKk2LX9A4FwGdLZhuppLh+9Sv5bHBumzARyi
gNhFgl+uju8lLlhIpHLFkvexrbPVac3ATx9ZIdkESXqFXD1uEnb3b9SCGh3cq+CGYqPyn2b1rGx7
YE6rBF//ZM1ugq2WXfTgzGFuXXAieOU+C2c7z9bUGdxvFloB3tlPIBCA+nlWn5JMsZTEvpvRKIjH
JRWeGjMaQEeSaB1p3tJRl2JBt/WxwEBoRMM+NPyq2P7PK76C9ze/Ii4U3Zs0luoWTh8JUS8wnpgZ
3wIjE5iLdtOxdK6XPsIusGgBIMr2yZYw/5kEbGL5eJu2Ics/GbG5aavBtw6WydrErje15skV2adV
+OIcb0U9oHrYSvb9oyAnQLEFgT6sndxDvkdcuRmTC+BO9DUJtUCtTsvMuPJYwDz5EQNFTpQi+eds
siNq8bin+iQ66SFILEGBKWc6VhfQBx24XJWUtsdmJO21WTaKNzG33A0PtamQKm6aSH3GsEDEUHuy
/jRmSDmaPWC0UZ+W/7CRPCv7wf4HLVSVw+ChuEe6sqQx9m2ORQpfnhlhqTfOUVUIB/IRxu8DM2hc
ExKsQfa2QDDrdml89y8AtZuD47Q8H5o9kjeZPYO95VmRet7spzvc7tXBndH7rvfYCG/m0Mv6B2UQ
jNk6cyDHxckg8PV8UEW+l2kZ6oD0JXPVspvt0+ZJ9m2r4j8HW5/0JOWwXJzsA8lloC6tUE2lmPra
ot4ASTH9ORkHMh1QdWztM27x8IDv5GiQ1xMlaS00c6EuqVDyth9o5kX4WEgDn0YzmOjLapPtKv42
sB6vfssRFU2g8ITMkqE+ydJP3KmRK3yC12iz/iY5Kamy6ybSPFUs8GaFGfTZkxCNMgKhIFF1rnWX
c3LXk5C1S0nn5S+X25rjcoO2lIImmn7bEGkc/LNvId2xIABNtlpu6IkfwfAnjjdBjI+BOvpgKwdA
0OeRHg9Q2SLYtWTU6xcHcx6DjpnrvlMk2yJzDlHH0BeHv6tBgoKhgdBcWIPRu/yZ9DNbZDhhqvEf
w7/zyQ9+EvWh1sfB0e83uixprsdlPEikrshK3RC4QQQeTVGg3oB0RA6hyOzItew4Cl6QYg7tzw9W
qegnYvd7LJWd1Z+wIFHDLdXKrRvfMAMxh25JpioDt1/h7JNx5I7l2tjTK5Xj2xoPq8mXYKa+fwfp
VEi8yDKo7wyRcuvBLSZqIT9ZSTrAdB6pgcNjDuVcTcwmYy7PUKwKZcAcQ5FZktIy6/tOyCdAxNQV
k2AwHwfLU/0/8eJVilRj1eMTt1U9EuyhLWYLL5IR0m5VXUR/o4iWxiDQWlzpGxl/RTB/bR+XAJY6
R1wh0o5w2DFzYsd1PVA5IYO9MoJ5bz67vbnD37I/QZIKmPdeNpnevCN05YmAFiKtIsvexYZKE2lh
gGBqYGL8G+WpdpcDXRaU0U1lYOOCdPrU/ztyyJ5FqHDe8AIYZE5HquLfdhABLTD+sDE9071fRu9z
5jrrOdHPg5G8PxM//0RYzQH9V3+Qy/jeeGIGxi0TfS3EHhnflRCX1kS9gbBBMZTjpe6IsjJNHLik
VUtHt6fLdaIeYwpr0mEB0DP20cYrVhNi/AhDX2n0Vo+S2c3tkUdgSX0mwjF1prDp2gRtTfXlyZc/
1mGOb/xZQXMYO2n8E36JA63etwPw/ceAf9q4L6D3ss1m/O1jqmVs3EbEUfKIVinwkOs7b0w/L6+8
oKhJiTiPTHR48MIRtsGIfCezGZdm2BZQSxXy4tIeQEAA77BIiZpL6TfbKUMyEUZPOWLjivFmsQxA
9CiQ9plgoiT6Z4HUi0VtiY707k/AWTNkB1s5gLpPTF4W69xayED50MeuoJ7CUP/mBkmh6HqwyFxP
Yd+AiGZP5j3n01B3UmKL9zCUbykuYj4/c7qBdBpvieapB5GyI4VOSzkUJKy7C9biM4puwWLlgvwZ
GiqxTnMqXv9wcGT6wP7JPrgDoxfulr/Dlc9k3Yj/TNYjQVpAvXp5BTcL0kTQDXt65Ai8AAO3WZb1
K7HyDpUjOY7XTGtW6srDmQ/h89QCconiCLh+hsFlk2s2I5ecuuXokhCyYnK8dqRCzomcnV0UZuWh
Jw8iano8MfEMAz7Nhfmd6yJOv+x+cctsoVL8oYKlwZt5gv1KxhE4buB+ZXvbjYGWenQZ44NWoxLR
SvFA5YQdEzDm1cz4v4uskYUiU9TdtpOSgseByiaBAyZxiP4CreQBrTRd6CGcJi4rD+JRLriLXSEP
Gwn9ClZleWyvj8m4LGLWfCtv6U7JX8yz2yjdrNmYRoAWUJop+o54Kft89acrSaTjlFmhGT8u3svj
6UEkPnMR67P0tHAbBN8ADgVrTHpDWElvMTm3o9UEFG4Yk517Nt/diA9zac7DPbcMGKKFfIQkPiww
/KAx+0bGWV/YQH15CqqwFP0VIXEwemBFr/plVVqbol9vAz9dpgqE4r4XzuNohnHbaPAfcwwkxZ2E
raJ9bXTK5IVrBon9SOMwEqtcNleQbWHkeY4yxA1mpHeQ3jPnN8QZTB1TD/zophYDO3FVXQFC47ZQ
lJ38G00crvAKWqzJOEab9wX8CSVzSDEJbHBZE3b9w5oz5dRY3FDkhUzglTJXzRZZwGmJAHOeLUIk
YJbdSKKRWO4QpT77JksqM46Mv1tFOixoUMEeroKredDoRpQXIfnSqTQmbXw3Fqj3IOLlNlwOwNnO
gm/OWkb7/3AAqL4pdmaXW5d7fILZ53Xy1cIsz8qH6qNYBFir+k8bCng1cZOtPpBX4sNWUdWt8yoV
cKAr71CgjJ5XaTxGWDGaP5k93E3CLkrNwSZoNrne51PrOHEYVjNZEVCUTONOnBeqLDHMHrzLVpHk
RUD/bYdEsnHMoDHE/JNwSTrfuchuqF0DxSE/JJT++6kD727UaXwD5EvlBzTOCoFEOx5tDJgX66hR
brt+qGOxOj0s8UEYZjDdWxq6NNE8HvEsMYB8pi7BZwArJnHLOE6sM++bVcEPS3qq36O2vUfmHtV0
reCYtOaooaHEbmiTAyTgwtIXWFVDRghnC/hVygQOHgJef/CgbKkm27vwRlG5TI2/f8xE0RHVrtr2
yiyd6zf0ZS0PE7Ax2ERB02clFHJWH/6ZKPz9VocMrSkKzPgzUMS/FxfOgUc0mMQX2frtiq82LLhR
6uWt7maECJQ7Hi3H1+957U53bu6BjN5YF9RZybWxQJ7Nb7jKMThjA0x57/l7OQvBWwXNkT9c4O8S
4HOPCRAWAi1pqeuTiQRFrxqFq9JtaqUWbW2wDUTHBgIpJ+ojnMAZt/V3PLXumaRzyrG2/d0d67S7
dhWdPVnr3c919pcyiZtj/RlMHkVAnRqY7KmKvxFCqj/Qylr7fxUuyImSoLyGi5lbnB3dH7JbW7vY
MyZWLmQQxB9Acs55FgJONC6xa7Qu6FmGccJbZl8vhNkIKABXKgMy3k0EsoQF7oDM8apBpWgeY+dv
n+gfqWbeKasDxN65HMJme/xJnUQiRlerKqM4Y/CsGjl5oJ3kcq6buFX4lXzKgtE1fvs86GAmVNMX
/YC7Kc7g2q5sbSR+QlaCyViDbAvsXRsch8Lg6GqvQn8fl42p8eKBxk1Qcc/Go21KnDFUE3I6tmx4
k1brsJGzyCwdiD6vFtjb652eRkIOLm3QXN116CkrkZE/IDJcF1N8kwIPRMMYtlPFArew08Y5J7RX
ffW1Jgsg3W7igw+IN4sJEpVXin1i0yX1KPo9EtzN5of98x2yJA+iruugbgryq9y3F4LKpqNLNtEa
dhKsynQ7HaYBXmthbAXEVkKXfiDuK/CGTa6cMDyIn6f2vWlR3p2EkOyZ2QzM/CquizWuKChWx/S2
QJJ3fbK92qQkmpOr2qoT6kSGFPtdpdgZa8P5Gcp9TyQ2Murttshls3slGXvliZb3uw1ydQ/y0J8L
BwhKKuWDeaB/cvHCQatoLaIQ1YHqgSLkc6ptnfiLkNCx7U4jVWme/1zMFZqB2ysePso6SnHsVfhN
z6YgeWvzs1lU3eO3HVYIxssvbLy63bCI7ZHSsvuIgHRaNHlri5HxgiZEu8vlhkbRJTW9KvPnGIWR
MS9eXqyVaKFbJCfxijapgR2YKWJTn3DelwIugmC49HiCRRxhSGc+gNt8dr9IFyDkBU35utEgg9SX
ffDYRaNYp1f8maRjEPiyME8GmHZ2LvgunNNEL3yf0UiNPKKlQETqoFR3vGjVvlMeiPbJU+zBZBjc
YBal0tNBfYpcEdbGPJVujb/c89myyIvULAOrnwYad+ajsy1KleuTXHnAYDVmZsxAstGNVVzqHPJB
1yqPcX5sKJ2tWIqyi8+UNtatNVlHob2YO3kuRGJ8kmaJejmIjkESm98rTMx0S41MfdQ/a67rmChN
vM/g2/uNsz7IXXFVrCRSUGEvxAEyOuncb4Ba6zz7emI8m4+YC3nUn0pPhd15pfk98w/97d7LcWbk
3Wk97Y7QRsdxMmo3MAVIUwlg+E2mwE2gywp/qxWSR+YubKLgYN219eWa2H57KJ8IQkRb8SqPWt8N
zX6nCCdgt0T92AvAQBNvubzHdK0QdKskyPeRDmuXxU1KgO65U9xfP9CJBDSvfoR1MCfQ/VEKxQHP
MjqS4MX3dLbxtPQQxo1PkSJKLioNIrxSCBqWZw+E7d//kog2q4UznmO/vF+OetHha3hOzh3ty6E6
w0ZSFiKRvB8VVV4WoGCHtjX4fJjrEmJU3xqnHEIBG35rKFYNaknOWhOyXcO0fMg6iaWwMBhU0nOR
fox7kw6bd9AU4/xmdaQ3Jgz8cwr8qBBDmPe4VW25XNzCP3zeZgBq0clpt5KwPvAq7Bcq6sKLgEWa
PoVvhS08g/+y6NXaLbFtPsCKHE2YKFM7jlXJvtYnxUZ6FcV5fWlkXN4oODothq4coRfGUXSt118N
t8IYSBHp4BQVt7iFkjgKq8jNewdkJrF9fK89tvtsn7YGcM0B2vRTlxe1+9biNoIa5Zgz40qowMBK
Tim2JrxGybxrPufYSspBhXC22UWF+mgmdvmA2MWpFwtqTrE4xFyO/FnbFE+mwWE8AuDmMClbl2Xh
Jb858RL6v4jxUNu3AwSFgssuy4wDfDjVOwenxdB/KmjWLFYxcVZmS5oJg40vbIThbmhRP7veOC+0
I14cyh9KoBDvYnc6KuH5JXlBQQpJVFg4JtjjLpq6bI80IrcJaPF9aO7Lzfeertjkjboly/5mtBnQ
fEYyDHPNWQjnTRvYMlRmFj4B7nRMtOxlIeWI7tBlrD6EVWx1X0XwbyTFuiNKsPGY33Z8q6PeMolr
2W6Ls/eZWrpikg4Jd45sgh20yzZFLgPIDf1hwSEjP5fA6JqI5R+NLrKS0xGUgWQah8O9/qQhYsDp
jN1D58n0PCFGgVVqR3eSDjUgEdVm1e+4XxntwHuce4R+cOdQq+tlcuI9ZFFkn0drY+wLcsT4sdmd
lPXpEekK7unYNLqSzha4DeE6Q3Rp0J1S+StfjUJRh53f0nvUp2yfOyToK1ioMPA4QAOairRogRY5
Pm9TdV/jiywBlW4grPCkcjiNrYH2E/Zets9sP3w2KRYhCm5XrPq6bL7aFCM4F7JI1lqrSRVcSPMY
1NG+fp2xYN3wl/VKCQBtfyroZWDeNxuCn0KJ0M7gRZY+0ElklqbehMGZXmc1equHbu2Wo6nuJhIK
RZNAPb694Q/yDV5nSHXzfD2fB3XccgstXu0/PnEsBPFx56FY8dh6+DefAUM4rHKodWa8IuBgbjPr
4ToFR6XGSSmwPVBV15+ZXuSHaezD+aSmVFr57AP0w0QucNV3lfhli470rzTLp6PkZMciA/wZiYqA
qiY9ZmS+Xb5vZB/uqpWyQYbLmQPl0TPGi24bmi/oZs2yX9OvqWg2so5fco+zc++TxoX3DKeu5Htk
fWeafZmqOBf/rmL1jK4kIXrtZEVmLx3SB7pstEujUXo2TQLG71WXbkZADwNnNXVgEf94Jg/i1How
q59PGlIbBIk9Z6RpS7qGFx1j55kgDrmaHPoh+9206kHWPFG02JY2kYinxwqPYUQ1aIzs7nAyfYFm
41KelGRFEfZxyTChrC78f33A9rKJHiPo02zP/bP2p3meJGkWvpaGW+wB8rp4Abem46TIpLHL+XbP
bMcGx1ucm1RS6U+xKBeV3p7kP3OjOqiMtbhKofftem6QhYXawiOiQ3UXb3IjDDFfYNRN1Dnw2O8O
escw5PtaPvCbHN+Xv2Q6TXdqf1ri6x04PbORsIHdBem5rq6Ueys5BqEPbT1peDjOkxEG7vaqQ6Ja
n/+Ex24b0GC2HxTnV1/FftMTkZ1xCYkcdRLZp0XC7uevNpYi+8bF55TmrZa7dCU+MAoPBfv6EF/2
UHQl+zXzI2xSOS2wzkSeWBtWDsbhO6lBLUw5kVZsifmesZCL3sKLPnDbCtpSTyhMoG1xdmEmorlG
NPVoAfPM62367te/fOy15AYW0NQdekBlh+G0BHsikMLcP1i1WEYgR6ulIA/KoflsXPhkhyxy/5f/
rRnnVfrgiLDXSszIExAbalwHZOwn7NRoMxD7ET8/gpq5gA/0wmLksWuKcrHFSc0HiAx/FKIqB33a
GdMy3xghqKkeoY7fO4c8l73bGjiyrVpMZcWrqo4zka73/vPEDQSVyZG/pCJoel6hZD/2KQA3gafj
rViNxPN67sLH4Qq9F/0eBMq9eSZjrt4YH3EYYuArzd5X+ZJ4nAg1k7p6WlUg65MMTo1xaw/RdOGq
9/aoQMlvGvcLs7IImNRYtdPOBy7n9zJO93NYXGY0KJvNO00iRXG0GF4xJCkmmzB2hBAD+kzyjkVC
wlCnQ3WdiVJmFGAjyn3ZgJEykIntgz7LjXWM4GwgLUbPJndSwQy8vlOtdsyNefFEUE2xFoAmLQ5T
kDUJudCbhb6DSOglwZtKFdNpLgoW3JfdRnB22Bg3WyZH6BcHlaLmoDwhyrG973No/2Nf6+8+Kx7T
warGDX8VhUMAX0YyaYuB7RfVPEFwbAyjALvLXHG5IuZY2J1tawC9NTs6cCWylSVDRSPyHt/D+Tu0
knSBdZ3U1asD6MJKGZEI1JyaQ8eIlek1VOOPN8cBYcENVRqd6BUZZmN8BaW7ifCkFtyb+M4Z50jh
YIxhv+Qdlvx3oGn5dqzqyxJqx3ehwzZnVrqGxvRkP9bQTUvsWWbhcY9XEdaI1dBsV63nqhBbF8qs
A0ojxdLB+fjlM3dV6IZdI5aqeugP8mmqiXVNus4y4cDM91ry2JqtER41HkhFz8FGFxKjiL+2EFGC
luu5vib//r/gAO07g/m7JTB6D0pH3dJIrNn/MI1d4mzkd2BEVED5YjuTj/cXm4YVX3Y4bw/P8+KJ
weFAoLFnNyR/jPlcjLExXngj86HCqjuvGBqTRKadPhkU+x7geNFdsVT8O8hw+9dU3unstIaTaMfK
erhy7pwQnSN95hFQff4seW38LcqPmjITEWPSkPpwIKYem1BbgejMY1yOQSogB9GQsR1fUHQfp/K6
lAF8cSJ9v2uQWWESsUPutqNxWiSUAiQ6mtKNmmrSa82upHnNUM61yswOXAI7ly1BbrmvafSogdhF
lEMQqEgJKsyDvNuhHwUDNJUJOTRwjQLpkP8Xxcb+lZQMHLWjaIBgA91hjB/FGBW9O/DFH2QZrQ8L
/ySWF+gwfFmLt4fzuPlFX21H7NWZHLizI7U2bh9EfrvKwhjR/udk77e5BpWEUBmHp/EgKxdso/8H
y0t8x1RYp8+LKezJ3ko6tcl7e2y5u4f2nZwGKLp0CkzUa2S50a1yGNzhL1qeFTvKjeT2RwOY/4v7
1fOmojvpD7KSw/aQM8JpJbYhOW8G7do2Owd/gwnk5jYiliZaY5T/nwpXbT0uMgJx6S5kAGdfPjAZ
+qa8f5EAfnHeneTy6q856c59RL1FNmAqbIBZCUMAc5JkIg29w5K4ldi+4IqsMsR4aZZ8TlCGu7mf
uLCuXJVQ6C+MDZup5G9JVxvS9IRz0nNlATbdbgg9gNq+9Q+riKLoVW1wfGvJMv2Cg/sDcJjQQihQ
7D7hQTGcZ14Vobzkl4kYulQLUUJGyK0wlArPf5LfEwdhWct16/r4AYrXwa4rPC19Y5Imh57h7duI
3Iji3w6z4Xa9BdrSIJOSSEacdF/2+M1V1HKIiCs2suZzCszaPYWGHenyZAICKCvoppUA1LHcjBi5
UMklbYZYmIV1tDVrV1CoCSDydUBllTS9WyUU5excKXamTjsw0N/DsitdjZgiLdCcTRMC0s7+SXUS
PtAiCmKDYDOKoe8M9H4BRbO3Q4S1VaBJ6uFgo2nfroZcbgy09k1MUyYs4Tbh32cq/8K/ct7hM5eF
gRowc1tIQB814KBrcEHwFWUs24KmyUi3S9SS0uai0S3Ud/IXOsxLve3FqTXb7U9cG00laHgZewKU
0OaiCPKL5im4wBkI6GE56T9mCvPiKNuV5YHM/iYcFdF4owsK2Oif723N9sn5sL9x/RJU3/aV1ETz
JBH3L3poCbWLVyeFJv39b/g9iIS1MFfaqN61la0XVW+gxde4rssvy3Rfs1uTICcVPHtMhhZ7/W7C
FCI3pDnsO1dv3wu01vnf+e7i2eAyoj5/n1MXfLduOobkz5Ufb0A1ccfM+EJrg7wGKCOvmdb6lo2g
Ef9dHh+dyl4bvHelNuULFjRCB1O+/jERQMsW2nYMpllB2OsbTdDPQCSAYkXP6Kfuwp56bqHFmd1e
ms1vEsqO+URKdPNlaPl/cyLcj0YnRHtwT1qIvCsdQSz8Fp70bsiMDKvv97ufNIydoMRcsvbNnseG
TLV1NPOLj0RsI4bKFXoPDyRaZHsRKlLyeaSNX79+iJadwmM8S3Ei4YPXBTKNmzfSri6DhtAr8f1g
YFweysKKLk7MyBr+o7PwygqdVmPsfvzvL1ya67UbDr4y8n/vuVsC4FedIN0Hr9Xmy1oMiOEAQcnX
zrnYfNfNw+JLnGm3LfaPpgnfgr2onDQSys/a7l2hZArsz3SU6p/cSdUnmU4CbT5nsTMrS7bTHsOn
stxaZHXjxjiqykUognvw0krA6OXMiOx1LuGJjY+s4SG9C7X2zxLXtwwuuSldPN6VFoICCKCNEEY+
Qlm613BwWUDy+nXR8zYln6q+I765QjZxDw3h2I7bdxqg/fKIDzjqmS0RhKPx+zx5ITwcxKpRJQJe
6eJGdJsRspEtXHE1ARD1K4f5q7E3KjqXnFrV9U4WW407soaMu9PJ3ShXH9XUA99JShl501Cs8Egd
Jh7knOaK31TSt5c7vGLHUaR/5zA2LZ+hBH2nVZSKP4XZ45PE/jAPV24TboOpWha15yqiHlCGj1DL
bXCI/0W2/bAhiQBW/GwlJkR8/CczbX4uUEgGSblOjS36TzqyRDvNxGi4bIdGS+eyaf+hfKZHXKfs
U3xv1pzx5YZ9sFS1griyuQQrGiqlZFvoYJRKicwRFOTgN6NeGvVne3vZ9a/6NAmoulA9VTfztV/p
qTfZ5Fb0iu7QShn+KEDcR1H6L6qeHUdWhNanJvCtPhhZ4z8sP5WzxKt3LNPyQEplq1/cPSnain+X
ZmhhaIPPYN2goIbaNuRP/9pQmaJl59YYpdh6GFNgYu0kbpk/L5fjMyMZzefDWFCv7p4eQoxQo/Ji
0r+2khu2zrgGUO/kt6qUM3V5hCwQCUx1io7/zQ7tfT7ONK1ttaRm+ZYp3AMnXE27tD6cy/l7E226
/nj/fpZgKI2U9/eLe77gPMyJPoorChdkC0OWLJSRo7MHv6z2zCumk/TytcYUAUh+hTRtEcaMvMbJ
nWL55m/EPfsU2E0uiRec9WGFz7tk3b34oDUIyATIYRRcrGNs333SOh6EzInECFInfLDkLwt1j2YO
BT3B+UXryYlTstfRVm+kYob9/gxeNt5An5PaJA199DsmYgZcpyCkyAjNK9vAzfDSgNYCxQPmV+A5
KIye51J1hr8q+0e8CTChvRK0RMTGFJAj1YafNrfASv7rxbMoU6d5OZ6cez7ycLANHWwoCcHaJpRt
35jRqh4789DZnpDouUis/e5V/ABipyR/anxmY1j3Uu86Q13pu483yBADKM4YYSPk/JfIsbGPT7Mk
5V8lSiH9ST/elaXrXf8hX685H51R2ZhnSg6Im5b/IZKZQx1tvqcJ4+T/X1hGuQBT8uZGJzDwJDxf
gANZnspfHdL5JtTj0Bl+4lDui7a3MuQdd1U0X1xcdxs5xjgpGej/Gfh8FhgPbSvMl6i2zVSNI216
Y6lmx1QI1n+Y360ipt2ihXqcH4df3AkIGTZuBlBxjFUpw0IMBQBMQhdDftGts7x3A0f0bzYL6Gee
ps74+llWoknc4+/q9VMBWbCeIOeqC3RcDB/VJDqRnlUn6scw1MGN4K0EhjE7a9xYoeIz3us+BGwW
5Z159YF/9cNgOSlc9vXORkpokZt5v2TGCJYD+fvIgTfG5qfYD7YN8mFXa8/xQXpd8ZjPV3qa7EO4
pDyS6RPy0yHWiSHDc2xRxeVKOe4oyHBYhBAPytO4t9IzT7GWGLAuV0cdfcJG923/LPq+499EefOX
aJlz6ZHoH2LtLyPmjxZbdlVu7i5FeNHRKmL0BAgL0hVnz3E58u2gC9velYAkPtkKlzH0BzfiF5GW
KBcLxRZWYTKK3uYKhGdOrQlyD7a2tmlUIkgpOQKuqerfsBS4eV+H4NC1JIp8OxJotiNKF5nlS6Xk
f0XwPI0snNWeruT2Ilp4o3nv3RH/ccNtZr5MI7a0Casv6ZoMa1dAdfRzNIaN+NGPwBAQi0jgkmP/
Ke0Mbt2+RzeIELkIubav2CDVJFrUOESn/s9Vk2525pIrkQYf7SmGJUQP8QIJNl16ardQ4PyZhFe3
9uNwb/fNGX8X4rRPQ9iuxqfXfIPlr2gRqfhfP+ZzwG7165PpkCWxmdTC6Se4PozbdunAvAk+q55w
ZiJTOqugVduqchZSZ7QEyztdR7cKzsJQ7TBZNOdKmx/95bNvCE27VZNaFkGsqeBDXFInH+jpQWnM
OIKJDcd85/v6W+Fz19zDQnwykc5g+VRQTd+8NaOn8WimlbsyhShEMhybdVyjpQJrN00wAVHr3ZCu
BMR0xWM9aGlSBa6VzGUFjryTVILez+2BVAkspjxgI1i4DgN1ESuKlokhXxFt7LT3G3S6wK/GcPZV
2M9/InQGE7Xy1Yu1sO0b4xCCydT6WidepyajyQgzeMJDp7WarYFd7DI4mkMWhbZrAw+myK2hGPHC
D/zmc7rSndQiEjGlIcAaapvYIVzUvT9xOiLxq9LAXuZ6Fo6fu4DSjpRkDiXwFMiV6G0oKXILN99T
shNBhvQ6IAyp2Bt0e+e0kC1zi9T9ejoSrJYozVyG4aIPSa7o5+FpI1bpr1OJB6X4wOcfxVOj8uzN
6fv0CI+Ssq8xH1Dh3Ho0sp4AC6EvWi0xbJzx1CTZkrWJmJuR8JKN/OZhelwpzJm53STaDa6EycdB
zEJWRsgOqNnyuGCuSWxaaSelmBsCIOm5RjcJlcJqWVkUvrFIxvCFI0oaEX8RtKGITG6uGKgP+K51
17GCx/TYSfYb684zmDzIxpqKVFPZPrVTMbmA8AYMWz/a+qmCs4jlYQ+bnMCmMBVt3FdssSsj8zOv
2HxnRdyuC7dMjqib3MV7VJQd2A1YI4VDvVYXFJWmpsDql71dOrM8NpAjXsL0Z3nWGIY3V0TJs9EK
Wu01JiWcYvoDEkO/oAUJfnRCSMQ8hPnAObK47jaIWeoXfQwJ9I2GdeXajNiLYuCrNkV5BU75njm4
qgAEGl9UFznpmA1rwpIQQBJ2l31pnFVB2iRoz9I3kTmuczSvLU46c2WP0LKO6iWS+6HVJ08JEer3
VJBvUGiwGdBgntgaNBz+TdYkNrf/t4g0KmuhB7+XBq4jkUz3vbkeDHc2TDQ0kJXUuaFYlklFlPda
bsvubj7PhP5sLAfb1cJu/YTnBTDcaT+yyiO4aCMHlch+ShSWJZPz2tZUSOmxy+cDeclMrhb9D+Wk
n34YkvJPQp+uVgGOwbbUQR76JAAHqrK9fB8WXWXlnpM/gjE+QK8FtsGByqKDRRrB/FeoCE8dNiNX
GfzyETUe8B1jFkkVh4KMK1qjs2UZW2luzWKcf6CaU14TpnOHMicS8MJsbKR0RDlotKmkHmB2jW/i
7fTKAbjr00Ui+ic9VBSnobTzeJdg1GK9nq808B9wQF7ldi8uutuuGTUXewxSfyYkk80h6EC09q3y
kdIjtd6ifQEElaXD4sv2pEaZ29T8mZzGfMu56B3SiKcGLu5ANn6ee/hJNhJS1rtnQ6vttqvtS574
qScuq86qX5qrUFLKXla1gmXM9JtEzr9lTvVYldfcVTvGSAgNcGsHSeCGr/8DQiqCE7T6z01FRv1q
bZUEhTEdYNBGirQo6KmcrlGGBqcBY8RkmUVvo85CNhm2An0ra43fxP7UerjgYjLg6KxO0FfkET9j
qEdBmtPE42JK0tUeraiDX2y56A2eGSiqPfmD1bEIYESI3fTiqsHHllTIr6GI+qrkQbR0hFide+6W
DscZ/SEkv8vHmH9q+jAC91mI9xbaktP/HQpDDOnnsQof9TaK2RSfcxTmSgHvnUXA2qg3TVIigIIw
iEafsgzECgC7M6IpYacjll1c+ZE2OZdi1ux7pbNjt94ffalsmageOosF6YjcdUBWWrFpOZfmlJHt
Rq/zAE0OcYCosxuIzbuB38EZCaRL2yk2IfrsP1r7fX4ECuWStmd6E9V9YlBNySyXH1DnzlJgv/f7
zu61+LDfX9w+gw5vHT5icrYVDLn7ixu9j4ZH5yllhbukKfM2n3rMRahSNRC0NFcmbnbOglHuoSK+
iBQVC2Che/s3YOlbhxE5nUStL9JbDvyV/UP5RiTHcp/BlYkNH1Zd8siQ83pJH125atmoZ9bEJH8R
WDsLullOlXGY8pBbKTWg3xEuT12wdsQPYNO0sb/acHS8FwugqFrKcOVrjE8sglOQGe2XmRnccBwD
xLCRiB1HEDcwT9u+PrqA5PTB1/A9gzO5h9foqvUcve4OWNAtgpsJQMwSHnW98E8BkuPDERSABFnP
X3j11MNPBmVIQfiNSmMQcTmxwcXHIW1ViSgQKz+UHpdZ89KjD+vSGxtdsp+7IhZMDCWwOKAhadzz
TVjDP6JJqL0cejpnXXbG3BtsIkckAaPrTLBuN0A+SKS1PV6dLxV+kDLaMCDgjEm9qABsYtVLgPiu
74NAPFFlP5ePQqD3XiavZZ2jUwgv7KTN43Ldvn2CpxBqpTwgbvZl3wwy8qdyFpFZ4SHv4gfTh6NK
rjVuYFzxhvb3Wv0b0jNMatE85QNydQKiV9MR7p1i1JrfgyatVFwQSS/xeZbVvqXZOFOknxJb55dP
IMrgrFARhTXqMGkfrIf08tqbFv8KKS4KTjG/evUlm0MzSt8JWXMOT8S+CYw0PmhkrZxjPRTxhSMi
vb3LyucxyGoYN+IEtQDkSZyRzg6mR5lMJbxlNOsdX0wX3srt4bBfTKJ6CRy4uCcPKdZMxRnqcv/G
SXRHnklXrJkmGdRxPVyBEDBUL6BPejUNwXxiFw35UtguVB3Gjn7Gj086AlXivbk4yNZqSSvueZwV
wD0Sv062yQ2/R0X6uhYvuK1IeDGF0LF64WVTASUcDquW9ktS9T5qStp9fAWaC3Pce9amarGPRRTA
pbtWVZ5MpH543vhixvfieteH7qVa+cC7T6BMFHgYM+vSKQCBYwKg8ZYZwttBh0Go+pNCrYrwiKuj
j/wOkHJW2wLCIgPa7/1EnUtKSfmhYDqUK7NWQto/EQ1GvYMU4DY+l6BnsPOsIfkaaoo/SBf9R1XM
RbrkAXIz1VfSEYvmo8LWeP0Gfw7NcnLpTTi5fwfF239riOL/lo3ZYqe5eiGNCCtMbVtXpr2NXZA2
WyZr5+04O3IvoNJ98EO3nlnNwNKhVzz9qB5nd8sAIYlwKyszg0fw0OiZ3b1d3+4Phzy4XAZZKsfS
8GynJo9KebRgTmxNgxikdXMC76Ry2PCdgxXxtIW0kHoj23yXUjGB5nhWKnnaKNHiIugtQ5KtFNr0
xfKX6bCGQjDDp29b63Xo6tLz8KH8HAPFs9ZEMFthzyHW9ksFMri70l5gXdtBIzQ1nNfSHsk2RMXF
1TGqEZ6C4gsdCERpAmNIF+1QD/Cn6fHsl6e1l7QZklYq/wNuyGjRmhaMk8hD4HLWBTZE5r0pfMSs
hEW66djBb6CqPYRVrwCQCcPoQ+V3RSUF/a7C7bsuvb9w++PeSigI87GyhZ54bNcOHwaXnnL1IMK1
sTDELZ9ClV1RopaTz/HTDs5ZkSyWXFwXfpe+bwoByBESLAfQ53YzMdZgMFXZSFk8ouEHmtBHJdCy
mnG0rD/KbfSoYlIzELubLyMi3FCBxDN0j2lTWUlUc5RQbPyj3dbT/Ndegph3kYj3WaX1uxHDFLWi
LHfItvUhC8muSpcTprA+oLUrt9BwrKWJWBVGIHnAKsLNAveJ05Q+KE6NEH3HHWxnc1nE3E5dQmwN
gAlbAdEwURUJAzTbUryUK2k2V3Uuwm8RTzi993Q5tgVy1Co510T0zlSKxHiSfGh3IX40WIK6y8k5
8gJpOBnqyMA4yGfUe/HnfcFB2Cf8g1K9h72Jm0hlTzSHPGCBUL2gwyuaIxBnI2LT7/bkgozxkCx1
Vk5f2pPsqBZlpao41sJRTuuzXxI6t9lZJRe+P1kJz8Bzw9L4StErAPE67mDuhoQirpTIAGZZiL9R
FbHWRm9vcOFjN/JKyOFzN3i8MxTFIdubrgPaZDTRToKJjmofMEVzl7fvAHGhWo0HU3dooBf2LGYB
RlELQBA04RgB+zZGJrQNJwsWQmwD3Rk0WG/IbOLIaESOcKb/XWJxKTaC9UiZu3IUv9i8YveQO9fv
QHSMO/YQ1KkNxOrJYq4doFIY3lxuD03mKk0h5hiDnPx4YKdBTBu2z8QyqlYtzG0dh2qNGvGUgIr4
w8+W80s7csJKHrwZsq5qRZ+pwdzescpK+Znfx4gN1mFQmMXzDX8m7MH/TRI38TRivei//4+IiVZV
RSD9UUfu+kph20KrO+VUEDwCDLc2DDe9a3a7Jm6HK97hNP4m+Tk7fR5Q/TO9BoKHfu2zP16XkZ5U
Pg4rSyTITZbh4LDD54k/Ssqy/RGHw6m+u5LDzJuXbb4dJsAeRFg2ZxQewroJdL/oPEmw5FAV3Cbk
9QWz3Hzcdm7IQJxxMU+SSI4yQQHznH5aLmWumNpnYciYBIuStBx5X6J4zDFI3utQTOpgAgsxe6EY
N4ZQxucBAbbdifmDnQdNorEGBBV0W5VQnzGm2rNg2dcvGVtrDN38uuS3RR7CQdlYT7a6/Amwqmu1
+YhzRxWmu3dploROmKI9I814Fesw1NaK7OuKpFA7Y/kusHGsch1Wi3DkDUSR/Z0wo9ZiQxexyhBg
fow6THC/BoJAZEQRyzADqfsw/ix0HtffV9/+LzS/PoJhzukz4r8cfYN9LnOJ3LEGJXMK9I1g6EzU
CtvB0ZDmFbicrqLltOiPRWqrjewOBUdeKjWY2aX/tA0+9p/FH1mdjb0liH0R8tOdkVPyYorloyS8
lqFsOa+e4o8Uf1beCY3Yd9lBpU19EIRAdOOx43/h0q5xs1eygfQS02v8gVIBLYuRujntIJmisejy
Zvql+I7S/KUh/5E3Ou3dvwQECtWPHTLhvCuultCmwK9HGguWMXA4xDinhz7FYH5doB/p40ZTYm0X
ZH+CLEV0sHK5UIP/kyJb9n4jXuhvyaLU2ugDpL/Ypj5ITFLReOVVRn7eJEV0Up3eVavJ7CWWUVbQ
ZU16dIp/P89h1xj1nYmmralyyuuE8pAMXnN4I45i866XCvetdBIwqiF9z0wjExtee9t6TQu3OFg0
t0R7mB3vbCRLMcmjiRJVfhiJSorbUlT7l0woURnogJ5nwUSbKA1x+F6uok4TXCH+MgHw1obhBjn0
lkMWHn14w5S4vDSjxDbfiKeeqFgHlf6pZzBPRZOZDP5Cz/Y55UEqBxkKIMlnQzxPNRUVt0s4mTko
PwMHUqDrkue5N4AljmTh3MRmdR1wOQKvsK7aZ9qDXt1mRBZBas/T0wKbLDbq4X2iJQ5LeOGVwsN/
Q7WAqJoTnxwlW59GbmEOL4Za6AkmL97A7HUwjEoYccjSZVHUov84VwbbvxYMckehC8JcQ1Uu+qJF
Ygp0agfhogfrKROgANrFASm1dqetNF52zrTpT1V+KHj5cELcmHCZiLrsoYWfTFKhYqEZ6yO91/BX
a5293gNPsFUMwQszoBw2RIze0q0HIGn3l1a95VmUMhA6e4ld2Xl7eCyY0TeH8iYXG8i93fh6Owiy
EO+YCaTP8o6huElI1y80jAQCTNon1lajkkKjLAMmE3dVaBEOBh6CY5FubTiCDlPfGSYXW12Rdpn0
g8mJ7QwWkfWtipc5taFd70ZWQMtnmleyGGblz5/k5Foq7ta5cKi0nNLpTw4l5IAFBhxRQYUO8rj2
qdCqnpKx0t8EQKbQhHswiKWvUEt11/U5Ubarih69RT4P6nt4LsI6kJxhlqdHbBiqPgYOkWA6ZqHv
MG8vVcHEzQBeEplpsKzRsAkUXn5Z6rg4GztFVMhlbdOL7wQRjbNugNmIOPt1PonUsehQbs8LJ0cG
t8bNNVImvO6KdcqtXLFKoeZ+X7M71GZYv87ZKc3Onpvbuc9aHikJkYOSpYg6sXn1UxNxo2C8eRoi
YX5Gdig1msv5M4j3ffRlulqlfaMLlVyMRaTpZkS1/Yr1DVdN2+JbNYglPPhaXSxJNnhu1tKvwyJb
YmPx9EKOw8EWz2HPly+dREl6OsfVLm6G46Q01jGzjKQA585el06UcWy+widIF1GF6XMGa2hrGTZe
Exw6RStSFJmR3XpyR6dIQsCLtaLUJLboeSLDSk0JYUJQ0LBlysiLjD9Esg2Ad/JBm/Smj0MrECPD
Y9acOQfLICntcScuqw/N6erPxKdZNFGGemdhElDiWoUlKSKeZBJ+WTA9YLlGH3+tYhlPne/7NdHn
0n4OdTct2Nium9DoWp7eA4tDX4B1MO9IjBzlIFH7R0YJbrENqq7izl1hZaJUdNleu2OUPtClYQxZ
4RhvylHQzZwD9i90DRkDd9XoZdE1cjfrD1NqAlYglh3vJXhDJLw9BYmiDib10pw6juiKyX71LlzW
7ZuK23ZHL0tN+ZpLX8iUuDKo3x3pwGgFHQMGShiAkIfBTEDpJGAm09Y07mUk5mijrSESp6oWCv2i
uqhf5XuYO9Dt7MelD4h9HcQdiXxTJYZVNZNYWnWMeaMQHQ17y5dS1bokSxDpgB5cgUUNbL5e5/x8
PCmYcAc7P0e0EY7gvEFv/AfoB4vaY0SE2wiErVBueJ7ifrBYZxpvf1YhHQNJtSa9SLsYTivSxD/A
VVQd4MkUulr+6txXcx8ElOHGSTthFLMvF/jHINqn+R7Gbo/WPKbJM4N9YK/pRywo2ZmoCwPTtE6u
uZNkM9jzqYOZqOH43xKBHIKLCRUX2Bxr+Ev4dq524qEIEaanitzf9c+z+zFlf+5+opx2Gsf5NGo7
IsaCIL7xBcJ9TsmE5yDv9VmoCwENMVoH+eBofwGk1dI0BvsmOyKlcRaFv6RjnG2pTfHtDPht4RxX
d/t5vNmYFLAw4LdOLlZjcrXrbFDvYQ1K8KheG1Bw1xRnGbYU5TFTcP/C+cluAnJh8+iBVtaOX8QH
SyCKBQ1DppqcZ4FQ06ELA3tGrzjN59h6U9JC0qZ4TCOzuB+IsKh0zLewwbHsJBdr6iI6Ww57wMu7
R1V01zfd9JTMlMEsRX1oTZZLX5CqkxPJ0qf3Z3ybm3kB92dzOJdkcLv9rQzH31kJQjEf6gm0iIiu
xb55UGPjU3NZsN/IePHuVRPEXRlU4xSzMpUeJHa238TvW3Wb4tW+8oUTuMFHRD1LfQGI3EsOxZw7
8dphDEjZ6kwrpHAzuOT7Lz/v3XTdog+m/n4COkfsBRTHuXlaPysz+RPFyuXrM9hGdzq4vj3IiMHP
cCmkhPklNxQsWE5F/QUtWQ92Xd05nHk/0LYaMlM1/6MB6Mg5ynTgpcjFJyrktM8hcv3qSk0UvRLy
RN/uNwlaeJsGCjsvTiXcERRYkjLFW6TBEhJPRS1NQZqn4WOcPA6XVFhmUFbbT5j2CB/QcjTGrj8W
cmDUQwidm1T/BMmJsAhHvYpZAiJDMkstnuLqqLsT+2ZVLz7l85BAFPXrh00bob2ysR9ZI5glTUpi
OL3EBaL7cHTT0wtHwMSgit1aywZs6CPxtIHwzx2mlxMRljFJOf838OsmXRvxI8FN+n8YEjAILZcV
0wqyTKxHr+/McBBvNAeRGwyPwgIPY4l1Qq8pCQnNEfrOakn6ahAt7DbZeXFwlJwYwv51f+A4OrqH
OyE9WO8Xw/vVhEbn7zBFILAfIn1TIuaUFiNy3r2+CjW4tV2ZWqUo4U2YnVnSwt5xcv7BuoWLWb/q
qe6+P6V7auulUcKIAqBUSzcNolOcFu0VUMtD6m4RTVfePKxyMrPJkgcdYcDHDfPc1+f1LnUwYqtH
4owk1f2P72Yf3HQswZb0StNu3nmU1rIS/wN8bwtxXCIOJI8PMtq8/ltcC2hBARYvwSwXhSR9MGtB
aL2joLbSUSiZFCAKsdKsu1+H8zO3nGP9W3x4aqQ8AGLi707E0+pO9egwzlREpfKCquil9KsIV9Yw
00SC8ZjegazEhYfQeSyj1qMWPDXD3xQtiLgNgj9kg3Cy1JmhN6WsvQS1vnK8tPjHR38071YpR9+4
94NNOdZ3Ux9MrZie/5fKhuVGJ225rW9qKMzx3Twlid7bXYS/cFn3zO852gD37/qPESKLtDJ060dK
jICMIv+cw941KgxkInD7G9upDSd/MAgw4RT0HS8rXdtEiqpQqiserGqxgIuzNkHKA898tM1ydd66
G7RYdIr6s1KNVa79kWEelsP5k3f0IOtc1hrQiLa+1m9nuMuq2qByBOvRZFXXl7udPYkj8SuIqbVN
qpK9r27fu2RSUXBEl13mUOHq/0rdzF8lUDJLrzS1vaD0NeZo0UHGYuhvAYHrKEN5OuT+QhkaiSLt
keulEOUoGYNyEfmglpFyIyDNZmajnTz3DXvHloCAiyaJm/3qes2/FcFRUPJVqDkAhK4vm6N/+/PA
N2L3ReHbD+DiB9TpYsMX62Me+Pv2DAmcSBezs3bcbS5elPmcfgQ7JaQgBpCqPm2xqCj18/YhkhNc
7bJ+rOK2dlgZACSyMpDToGgY8A6Rt9vWoUdYi7+/LBwZPDBmVbiZG6mtSZcD09z6pqsfa0eaOgwW
mwyaiSMz6V+Vu98CqaTUfxZCn8hdtOVo0hQs6Wi0auRjbU0hGk06cr9VBdnogN+K/BAKO8iDoycZ
4qKb9PYcVIrxJMs6On5kcp/sYwBOS6hp8YoUo+Bbu38YrGNsT075wTE7mulk+D5IBDsEN9xRnI6Y
H7+nA5Yv86EH6CXVovzLMAk3gpy/J+zLjhbrEUV/1mTz3/JaxcfwDLWLAQPoBKwKGfIUYxfvy2zX
iXLcjfftf3ZvDVDHuPx+ymy+YPN2AlCP9PQCyLK/T7VvApc5lnWluWWXEI0P/bq8xQoJ0jmOsb6i
9Y/A8cPEZxc/oStmz8VapFxmzFU8k0udm1XBjTxXWvA5rhFy5CBiqK7mKfXcBeUqrUsBi0lI9hl7
Qkr/Sv06GQo3Sc1oinLkDODLwo2lQn5s6tLdt/b+9O0WqXfdu6wHC/VjGKorf8Rt8ES8iVEpEZRO
PNsF3fFIKsYQCXScJIAcQs/luGZg9sybPtKU/Vw6iJ9zR61c1xqwi2oOMgOedmWmHxb7kl+zjJMu
t3qW6/gypXwFBevHnI+MVNvlqGp9gSEt75t3q5VnNBtf97V2cizRCtWDBw8HFXFmfWXqna5z0BDE
t4MG5LOIcDk3fF15HKaeJzaKuf5WzT0m/fbsxghL0kLywVo89iZjS9TX9WLIMiWyZs1bWt39UcSS
N1zg2caFd4QFpefdSzFa5pwBqYv2RLgD0YjI4ciQIVgj/q8OyidkPeP6QGGkFLsl+Z8Fp4yDk6aP
FV8KhFyf2QT2dxhM7W76tmQLvN0JcaHtsY71669UA4h8neEeL6CEBsvQK3Ln1KxLhwwKdwlHXhg+
9vX2ZWUScixlRHuenENCZ8lOoFc5pfBz01+wnK1OisVdPMp6HhtegY7DSNT7ac9TYkopA7NiTbPE
46q5wYlp+rnGBQCSPdSRpWH93cAFDUvq8oQ+UarT2oB2sL/IUk5Z5s19zPCysw3IIPpVemtAs2qv
UShd2eqkR3wRhvIxA0IxkvYMvwjFZdGnc+JPan0YG9+mSo+HubkxGTj8z18NiEVcGCxlBCGHN92R
XhMFUPRNPXHA223PxB6yMQrTWSRvoGFfNxkP93+QJYhSjoV2I+YIQgc2ea9mMJRJJ9WwreVne2E9
eMEn9G8iuiu54ntKAeo9Cb4+Of2nf14g71csFsExnJIOmgL6PsYnT0uAcBgI93+njd9Gc0lD1rRT
54wXj77zT7h569AHUB7FxrQLk2plW4Grr5XPNbRzlYxj+gY2WX72xCmqrbU7CaPbKm8uxocKhtUs
VSi+CEnLibA7w6DVz5McgSd4VOimBROtgHD4ocP1C7YITfIz4xDbYMPzFiJG7SyZbthTl7zGegcH
FkEQdPmVnr9zDes/9ixaFfLy7mROjcMngggTWT7hh+ER06RnxmHL3mi8QNrv/ljX+Amzp9f5pvDU
930I+N+dQ1VgIKKARV4Uxpsp2cJjz+6DjwX/HZ3DLlIB8i7OJ/rLYpIrclWhzR3Vp3BXUKvCvVBX
cJ//W+vEdt9NYqKXaipZXdi7i0ojuIqxyQkC8CybBA04AYduTmmRf5pxLYg0U7UApvxFI11sRJiZ
LSPTzwwXSZ269ybISMXHPY/MbwERuCjWSRGTpsCT95HDhagru/VTGTYwINWlGZ1uJY2y6V8uhMGj
hbIzVI2G4xMHZVQpa0NxP+bjhlYw5Loo4MD6CMYVieUs4+KwwWsycKzPwqy2ZCA46v3jySuzoIKw
VNU7abQZiXmh85zNS3iAcpFADHLPGTX5+0kPam5Q/WdE3F2i5v4i5/WxwY3qsK/c6JExDK/Vcned
TMEC/2UwLPk0wnrkHdPrzUjsP4YEwIvyUK9odk5KEhwRZPLzqRjN0ryxz1wswj/NR2g8yba+eMBE
RboXYnW0qH169jFcwWmhHk83fix9u9cgdapwFd0TaCmqG+1hP8eaOTUk5SuFdTOM6znQjRrmRbon
NwpgG7PgULhxlKvOWs98nSAhfucreKIAEc58oDysuI8TYlzokWogKCz3i3285Nvq8ZEUOvcA8guh
hs2oEMXO6oEmfK9qTH80EXmx0XIz6ZkhaFoC8JfBG0gqWxegS7ov5oEjFWMwG5nycKSJydxpI4k/
3+k408VZi9gM+rDA5f5FoxPVMomDQ3G4xSJFhCGdLFeNwnkM63hjAORCsM2zYzpYo4O/DU2/bRiQ
zf1FwG8tY72QsX9DqwNvYHE52L0kZkn2o45PsWTFvErpW23Y76K7j1A/ifmXN3Pewziqal/qnK30
fmjMKm8UC/30dtBf8psL461piKroN3d2QxbBkVAWW5OfqAARYcQ5g+ZUGp90TgDZpT3S9tU2Hzj+
z9iwDLWlqN8L2tQCogeDHShqXGWQJdcNQhKbKJi2/fDK/Tz80G1iLAvW/gh36e8YNe9pRy89gm1Y
RC2t9YeGfBFMbsuzBMdJq71OZXQJAFtce4V56wr7ewNg8rqmQ7A0k6drB+g3q0SDNbvLrBcAd83y
EzocI1UCaOainoLPzqB4zJm8bbVxBmcvs4r9o8vd9uC7y2Ppy/nZUQzVsse1j2ad5RKYw7ORyJsN
opNBkd8ao+Dv/gARIGg/O1H0DLm0/Yq33Sil+99rOKy2N9YZvREH+V/FO5LE+tmEbTK2cvZD01Yt
G9YRHwMgJF4UyZ7NUx7qs3GTbpYzoz1qifSkqXDxMsgAJE1VXePWq8DllDx695abK+Uf7ryFn88X
mPvIfcu5t+QVDSxnkz5ZZnvejWvQNmgrDlq5EFOs7MikXPd/gck82ZtMtkOXzEhoHxxSWmTaXaq9
EMBsw5TNSEBtJYSITl8bicyp78j6kleOtTLbIZSXZ2BA0pvD5yhC3NA5FnfEnb2vjbGF7tM/Vwhj
xNGjvPh6+0VeIT316jzUmnUXv9p1AVFRkmVtICKL1Vz7QGzphy32fGtcSTrjXeSjyAMoSsyyD+zG
Nilzy9oFwmy0SOWI4Khd/xk4LZVExJWuoYbBcD8UCXB+i4o/d7Aikn1zmvjLTcmfTGpuelUannlq
L8WQw0suR7ama9kv45pomSZ0qw6sKGIt0lIdz72rikp1GoyX+KgkmQJQe/znbbzs5/5keFMOYOmp
wg6sVs04AoLV0vIwb1e6IXk8Zlsz2q8EAVFQWRhQc+rqR1FgzVPxlan3d4xOYdHYSvPvs862lqaY
WTxpzciLT2KtozaBD7adN4chLr0h0sHYT3nldvW22Ns5ym+TwIFxq871Iv5DgAJUrcr5L4SrzczC
5ONZ84hmKrKxE5R8mWvGpLcXsewbhuhvPR3e1KOLOT2qYrGTJHjE6oVXPTh1Iw82/BDVz1x/RoXy
5kFj+3mwEeEtyVHL2jke8CmpIsc2AnRMOE+m3jld/pp3m1/wCFxiNLfWaeow9REpDrpygnzmx+Sl
EPiFWaKAz1OdSiXf75WTCdD9Pxh8vdDxycv+uwJdKG45rmq7Ork9Uq8B65JyE3zMEtFcFI2zHiD+
aw9NbL2P89g57S4O5t+CvIWRDvU5bBcJ5qnN0AdY5KAKEqpWbHAviD7hG0IdjfHKQzCb9y4D3rkl
6Gu5pY/YXRkRbVzyPa2lqXbu7gc6n/6Lt1Gb0Uv5BUoS8dfG2J2A35CjohldcUKxCt/JpU5JWC+C
pyWcUo6F9HbM2Pk7Iy3lF6u/As+V7iuP7H/ay2zzp+6BDseHPa89xoP5qikrdbIqd+1SyYBn0nbY
kOg8tcvwKOXfq1C9w0Xse6L4m3onuDyPhbTxCXyYENQ1BW6ad9gPZq314RNlEHnrlTorYCzz7dpy
ZY0XAm5m0GDuqoSKIwaVUtKB7W7eEP/YFxLVH0p9zbU9jaUW1K6uvD5WEgaX/MUZytpoC0YIuJOk
nl/nsZq3Szle4Rs41astYhHGOzG6O7aelJtdJgnLcAAxMEiFxW4HZTYr2Iw12mZ9RGCUK0iuVWiZ
JPh3GNDI3fl17rCVsR/+dd0QjH0U2dve5FNXKhZzj1FuIyUktogE+46QDoYREXgdNnS4dTx9/2Ak
EjwK60B+cdLLmtQiL/bL2/i7SBmYmRA07tV/VPjZgWUIuVeQexkUEJa4aEs9yeOsJ0FHSUaNcIOk
s9sn0dDLaInJbC8YNL2Hpq1Xqv++M3LeorRRqYZ1UASF2oEnOWKsGxkqWZJgWnHy9+KCw5ZjoHcv
uxTr45XHRkr2tSLRmpo5E5JvRzScqFKkSHDNiLnkAUhxxXaXRlqo1ZLAqkWLy67Jjo/y9iuHzfZW
FiOIKR4jvaJp1TeY9D+Vq6NwqSGVyzjKF6CaRNmu2A9XWHBJpj5DZ0BFj1NohlsipNzC4bGmQFj8
yzKi8hn0eATUkU5v2+wOOB4nZzrloLKpr4jXuhb0ngUuPOv/jijF6t51sQk4JMmYNM6jiQMrLOgE
GpqLN0MK3nu1soWBLTI3zbhtsTB3zyy17VQH242iI44FbTbJMnlI80bRiJy721lR1D04xq4hlksb
KOi6xSvV1GSbLe8F7CmS7oWdZJJjUMx4H+BcPg7WuKXG+zRN4kutxTw18oJd13098zMpaj8JuUPY
MfBDcTjwDRcHTBjHyZXxhplIGXc4w5L/OVnWvzvzCp0GARJfUgd3BVhZsCjGPJv3KPR+3ZtPFpp3
2riPIGYAbRuXkBXSqRMQ3UlYb4mAGMT7rDfLqV/MV2opS3zAoGpOe0nTYY/rLQu9TCR2g5HVUQ9v
40xRf0yKyiXw0yvIRGgP73sXz3uHVhU2BqgJbjwG+4VidJ5qLPgRjW81luyuGnblis5zGF++87Hl
Vi7p6hmy6XGABrbdMy6tHvtLYWTNg9dgal0VS6WJFwoJEYbow3pyTzmw9ZF2oEhPuzsON4XXgwG8
W7r7iqvsSv/ZTxwdfayEhBJhPn6AhC3vaXPta7CiiNI2fhfy+/Y3ZL4czJpkpOOLYKNFwzR1WB7q
CaVCioGITWdlEjSS0RxCXKhz1ECllByZVClyJiayCoGsGHhkoxtJg5z81ogzk16mJqSx6bSN9Wkd
ZoagC5sZuNH9yuq3f3Sffl0QScGAvOS/oNCQLDznnS8wi+FcZbEGaja312uS4tPz3o5uH020IMsN
IC1armDus8XYvz65gTl+koftMK5WR1S1N0JrwEHwk+skyKpzJbD0qrpo3jEckZZZN5rVWkjm5uy2
YRcVpX7tjGjUDNLANz0UAZ/EfV0BYVmPhEW+ivRrocnuZycm+fSobIMOMc5riZbbTzqkT5hYZy+5
9rRpcFNHfaIwDrBtzR0Vyf0GDMDBHAAJrK5BoeB/Php9+VdJ5pAv6djlxWjv9r9TPx5jsXHi1Gz0
1/7fqoEH53JvrmLdtk0zpR3eR6XPcz9FCD6oNG85ybJ52S8XDGA0sx6mVoA64mFql8o6d+Q/SFqt
xFOn/P6eWQY16VINJgnE/EjamvIWMmUkJx6/Mxg+QQ4k63WVc24WBZ1nToRcu2AcKyI8kx5gc2oR
FJtX8XzkVREeotNRByOLBP20W9WncpL1T1O/3sQj1uvqm8ssU87JqiRKktWN9yZfZJtuOKHQjyv4
Q5EM7JuPBVsFVWdEeBXhpisM8WLRMoQdaECPg0sHOy0mvl8N0JG9P2LKfiD9O8lmXlJSZN26WpKS
swXgKYnPxdzpu5fSfPu6fcksj4K/TxZ5g5DCsRgEdt8Su1kHI79jAkUhYi+ggP6xfkHX+s3zIZo1
QUBnR7R/gvYeCTSnfmpKBHztU8tXViXUfSwOuUxpXB9CcfRUt+YKcEsRql8RZ5gVTsXw7LcXhhdG
ffiAJvrqyi0SbLM18k4NRzx15O3XbYhWyx4k1wNt0X8w+oFaZv73n5NeiBaREB8D91yE3WnvvVwH
uxXrWzjtGNrNF9olfbWEs2fbQk1Zh9TspNWpbYkAj/6pFC5u7N6NoYS9ch4pz0kQU5lA6lzm5FeA
4cMpFCXY69L0jIfieJXjUPZxGwutC0SQYV/RnLbzqkUFYVepYpYFOuxmT2949RNjIEzqXGVw5Vlh
6/PGCHTHiVdDZ2r1tbrq2e5s6sT00oWzSHLik0/9cqG+WtzbxZVByeIMfX5eYaDXIqmAlmBbGzWp
/BD8HR+YHxqUR5YjQkX7SUOLuTwe9S9fDxEGNnRCGO9KazxH40EhjqOzBV1VyraeRhc4gU+tdhex
niAVhJ6n5QV2b1pNMGoa1hT99NYB7wXdAx7kYg1Wm5dXZLxN+BRJVay+tQ4sAm5LPHIW85uC3g7i
rn10nyD4lwXAWIKyHPKBSX5cD7Pzjbm+UktK8fzzI07nHe7feBnyoMU8rxnq7EMw0PZj9TnUqDwU
XUfs8W1QN0SVpprQsjHdmDzgi29Bk05JgG7Ib1NBhhsl4FJUeoVe57M0YfnghY4B9r37uXs5q1IW
SRS4eg+ljl0FqqHEf8SB4BJlDeh2NpMuuihC5op0rtVZgAm8uMkf4UT7wnYL2Kms46m7ofxPalmF
F7KIadpeZAanaxeecS5iMyuWjxaPhpcJaRpBkZ8mlkTTChUNCZpFg96D0rJPZGqpmPWXs6TbOd98
66Q0/eUliswQ9LWWiZQUfI65+K0j1jSpevq2Y3tOSjfu5jGO/u/9iqFH/eoVLrY3hkbf6eF+X6wi
wef3c8iE3eBEjajRjNxbc3mLcCINd9pR5U78fMj9cx3iuhznMjWf1s5DOSi0GodovLF/QxOZlNug
PgpLOVOEBeQZJ9xFtLASr1APjTNQKRT7yztY1kaDinS5FJtF/HKvOmgSN9jnN43ulkGOQ3sBdW4k
5OnojPsnhy2v38k70n94rO5gnIfZIUIqKwjI4pfDdA7vUeBPe+TJplpeKxR4PWzsGqgbG+3Awlrl
+yLBYsrX5t3YFAKNRiEIUpHYNZzouqWNxGMUnHau0Pu+D4ixiXnknlmW0YVwDx9GaRXZaNyOUb7X
FIa6hYoHnGKzV0hor2o6KHc2DcAQBhmz+PWETSzy2htHYc72AC57GtAjLucQ4huReIVjrG47lggl
GiJNQHlRbDY0HMuDaYQYJE/QqaNI8AM0vcAQ9khnjRrKK2+Auu1PHzeUt1VT3YbaBmxe7Ue4WX5t
N/+98zIfzQvjrG2ria/5I3EXKlq9aLz1Is+SK806xsPmvuHQ1xhh4TgTBcQjHHqguLTrUTN41pAL
SPrc5dV+LerPHVFseszVjiDXR3AyBpprDQJclbc8c51BFr0zMAdwlw89umtgv9xk2G7iN2Zq5p19
ERG/UMIj5Mc8VP7dnjhpxQQCkCkiQ53qZTmwaSRfXOj2+twQdmQS++B2VgvPdiGCVqZqyahoRy+Y
EtD/gyWWNvo76L7rNvqQkLHHsabRsvBAmo7Hc1vKkuaYST2ahkwf9wpxEg8il9nK5nBY72TSz7xi
80Lct1FVfhW0OHk672fbAT3v1TMqtFjnpH1s+oQ9u4PrBrMC2Hpf/i7lhr1tjfKl3FPLw3iX1HjI
EWNS2v4WK30oOkBjUiJTyWYSWmo2hVAcDeUZwO5aIVEmnc+vYFcnj+W52OMsMh+Q6Bzgmn/1OCZ1
Jgr3ydhoYKnP1wrfPGp7h+16fbowWKAw2L4xEECA67tRwNs7iYo1Bzp75tKMInLuEBEV8+mhtuJc
8rUerhw9JBWwfSCHAwAWKW+gbLlh+UH4JMIfH0ljZidC1aBgbCRdVUbKoAKw1CwsobvefUTRLeeU
XagkbLzvCCikqKvStlqZnmOYmpwgxzBgfrdik++17tgbfSYVI100/xDGIa2sqllZarqUps9aPTjz
dgeTr2aw2fDsNTYZHiQ5uPQ4YmdM7mESUoCXA1Ei3EYhUafoatWmmXemEld2gShZCt8E5FQbPeCs
0w0gF1vAuto45dO6SmB3paygny/wUlEBiqqVlbOLneQrxapWUr4/ao1VDOdm3mf7e409dej8sCV5
mBGR9SN7pyc/6JvECAc+oQOkjSkTFkypgno8dXXHOW8zsm2WrJ+ENkEVWnW8OkpF75HOmHx4qbud
RwXqpqPqJVdicR6jmpmKBuDEEfzqPXJEjmx+BzdC3ZBHH1KwPx+QYZIv5Nvatdb6rHSE2kvd6I3x
dLgStRXinDBxaTJVg8qVgwWS3VAlp/XNaHXCwO4XluQ8+OR6M8ta36DFo7fTpwrJAQH7E4ON1VuO
uq7dp3wmxXN+DSD4pzGNEaWqhqCC0Rc4a3HA/DFJ5wKNM9cMeMbL9M3dSY4ruJJL/HC9yTuAtYOG
S/NradrEWxjRkRjRD1YfuSvNedPD+aFbV9E9tpbyvS0ZfFeUzVH712PdZzOftQBa8Uv+5j0Eg0KE
wl+Mgu1SY0wd6oKcDlAEiQBKUQNlNrUiwVlz4vM7dT9q5ZkenDUfAiw65AFN13ntRfiU6cm3twvh
eLtCSmShGmVGOST5KweHyQVc63NaqVURNBNIIzStiiEubwDGJPt+Uyx87SYM0DWz4A9zIFb2NNs4
gCDWBZYzuauaZuG0lX1r4sgelmngxb4w6QJZ6rlo3kfa0g5NoG1rlQKqdgIKlv5+tOW5+NyYz+lO
+YtH6jahMJ2+h6eKlkKnBTamNR7PyHKzSbg6jDBpPiRwmodHx9dFzoyDkmvuXqPGz5I55ZCZvibN
5ROYamWvCTJ5+UUF2ynVyj0bdfvMtmLLyu+y7uH9CnV2W5qkBx8S5DQuHjAKx+igHHy2Sx0x/NIz
BNqp9V9DAH3X45ef1Om0xjlvydBv2UCoGANW4ilzPtSx443QDEL1T9XmgJlky/GCeGdlP+bvMJ/q
JcX5yX4pqkEq7e0ojWILFMwTg8T0glafF+JAX5C671bSJpUBfcH8gOhmhctAsshP1pFVriUSGWuF
mcWV5U7zYj5VQBrOlZOmJ3EQutpjGOG4iUqwzhb5l7D9StCyKPTN7rS0pouKZQHoGZuzsQLYPWo6
0qdoaQq1Eyq2aSZmiiI+MLzTfeyv+QZVX/Dz4vsLVb2RHnrde66GL486LgyCY7/l6jT7ojqTNKtO
h8UC2UFX5POF4oUCvbzC1/U/gF7hppSJq6CW7E9Wtze/GYWpgFseMXe3FEkkMH9UZwrQ6geQ2ITT
iuqSjC1KW7jHTLepe9Aub5bbjSl4Fwg9iVWVGfYFWlgEB1qGMYkA8QVcCZ14JdXMKeJJ6drQ+lx3
1W+1t7BDjAWRtOypV2zNVeB4Z90ialpPr4gZmve9ulsOJIrudWO82NLQW7TIIaXag21hrAVdi1U5
1LWQsoMqBiiYmLlPBnMj5brhwFIPnFph3Q5oLh+oKV6zpRzYaQ6KGRHpTP/29pWzuEMZ/+7jwWS4
zKRwBpXrmkBb6Rth2SXnRdiXMI4f3mR8WF4ne2N1uCeTeQ6mDm+Eh8woczQ9GA+VQ9LkOZVQM82I
myMxOtchDd0VZCyBW3btnTuBc6lwmcNlwQ5hfydGUJkmgaSuFsq9AsvWPoVk7hP/sGUWgjhI4An1
EmfA1q2aM8Zpkgutd+wBbNmTiWqoccbUjQ1P4SkHjx/gZBXscxl9m5aKgtA3aOQa41x/Mf/jJb3P
pPJP4eZZzjlf1AH4cbcqLjfLL9UYxo0SzFEFmD9zZKmAJYNJ7MqcKddtzz4T4eB2Iy1UOvjfnyI9
z5j2x8+1JLTNYFqxsk176En8n9khXk6A6YVlbwVKmsjtj7qBB79kJbFpMPFKHEgXpp5EMzNWzMk8
AyY3N13Ckyb6e5jFIonCRFZVbwir2WJ3NCVw73nyk/aEOe6+ejnkJP2vnPFDuQ67eVNl+iKZcy6t
EQnRRnHoJmtCVJvXy/lb/+BeDmnioe2frkbQw7SFd6Z/eDFAkCBY6SGrz56Vz3HhXIzOO95+dz7+
Ieh4rRaOP0d6DzhKbTLRioZPaHVqKR1IIGpxQzEKtnkxCbaA8Kz0BN7jqopwS2r7lUS2M9ew62lt
AFG1pf9Wy6erN4fTtP6Py05fAlDaKKNc35XiCiXvuqvIH16EI6L2hvXoriSY1k4P6kT2P+ZDxL/B
8HdW0JhBwRrYz3CTjsIWJbJRQYeX8WW46Ayi4Me2xlEUD8Ziub2nZzQ5sumizdCDYWxpoqgC98Mf
53cc+EoM2uzp5V5yc+MEf8HeFRtyZbtbQjNRfjhENLa0nPsiHTfLbOaTh66hcGH3aXAtmbsQNO/z
keONWxFeg5RkI7u86ghBBBH/mIC7dIHSxjl1d8XfSJJzLP4K2Dvz1Fyz+yzFtqp/7+ziQVoPXBIA
nQDSHPTTA+mLFJjPg+NFTt3E0eD3erR0LrR7N5rpkw+492knwZb7qVIFloWdo7M0g97DeFAxwpDp
YI8evZUDNd4Q87G0xIDC4Hj3WMHs9fgWtFBB/rbD/OCxLbhKswgcd4i+UWFjew/gL6H8MkOtDtlB
qx9acsZduHid9ibUVslZ3GQYB0njRdAuXzUUtZbcR1+0mI03YVR2WQ2EolKRKiKcrUupJWFkT2Kl
DB1OuGpcLJJWZZSLmHOtwjfNryn6KDeEfUsQWFPt/63J9RTwcM4Bx7qVw8EFH63hBcFXvPF+lCsZ
rcSTofhx+/+Y70bUTincDeDDEE4o3HZuieutwTimwibFeVFvYOGwci3wthNK0nd+kY33DapwrpG+
5tpoMat8vsaPPYGvSptDmfKrVNm3qJPavl2UcgYhG4SviKQyldcYejpwVI1z9Ggv88tRM8xVSnC5
yeu5wDhNK60nnJXPrA+yy2R+0TEaGQhlk/4NNRABkyrt68zmBc9vHjpdgcVklDxcfLXKvLFcCbdB
mWHfmDUFZKpD4EFEdHWYJqys98G3eFJVSVyuL5kyb83blzUY6d7t3UZgLgl0CpmBQJaj0GSDIt6s
N8YdOjT0FBl7jKsmTVTGGlem9uZcFPSN/6M0UUDgqRHPimu9YrikJm+kTtkbZD4wFFUpe2fRRu0D
TbeDflEsJytjtMwHUb47ujMv6IvSwK4rDw62y8tIEhSvZb36+ONj+qEkhH94tZ8PhCHhttr4pTjZ
RtHuBMweVvO+IGbSmUhTzxxzBuIr31Xnib/+Tio91c+3yY8ba8AHC9Nl08cP7g3q1H3By2opEB4o
xlsh0kpKu/qwkgPfMmuX+Tq1qActeg3NUSaTqYzRPPzJtImuP/YnZcsadJLjIDC7QiOTKl+J6pxH
V8C1CVnekTSx0VIItZPdAgD2qVHFJUwagkaDy9TvEDHV5YArykwQASiRim37Rc3qXwBRnugD+aJJ
yy3W6iMK2l9O3vI5kM2ThpFBziioKvy8pBQgGzUcB3Ov8WhL1wPRBo7sanMdvgsOaumvwKMMvfrd
CjGOMFDBB81Vm3hbem3KwoU8G5gzgEUM9jGsO8vsHGNOTTF0edWjP5vPinZcZWuGPVk6Y3pKplAV
7egX+0RyoqELFAWw8BuCSmRFz6Vl6W4La47I67n7tBhJAYCoeeW0gWxDqm20Zss15h17ulsuFA2T
mstb5dIjy03icHknaHfGXE/qm+vNw9apsuAv8oFsQ8eTVAk8v+CVn5m1VzfCro6Ls2QZQAUk9knP
69zFd1vV579qVtAelIcHkYvgsBNIUWpwua8jHQ/6vOvU5SHU3L9pCAvkoMuJlzJgf/gENN52WZIm
RiQFoZe6WSM0tnpyzrKx1UV4lF0FJO7gJXiQRGulvhk99wHjrHv6jOi+9T+/jzmoGHhuv2ysJus8
nBImxY59fZ5kAB8+FaKAu7kLVh7BRlqnlMxZJrZJTMopU8sL9r7Rj5W8UzSKjR5uxQk+NljtKMTI
L+wBj5M/7RhdjWIoRgTCCeRkFJcf8CKMaeVoWTmnu4vap9M2eghtU9p9ukqrQHWE1DHFTnl9c4r0
+ATHctsIrzVX8/rKy2Ad5XYZOBsEkuFGn/tYLwcMVz4ueNvTGYGo/zDKt6jh38KgsC9i+fjFSWOh
pTWcb2W+ib9RgqyXEBnqNRA0TAtmsGXY0eFXIY0IQPqa4UXvB9lfGojl3w0yj6ZomiE4u2ziC7Ah
OAw8VXHU1fjUXnMgVY0RdwPEcHoRBXR3/yTqlZRY0LoSCc0jpaGnxZ6aaNaMEF6S5lBNXjI7OdvQ
aS92CvpG5iJ/KwlH3pZnYi7SJ+7vBl+VJ0d5d56VVClzOHind166MCs9fdpyXEJgLF8RBP594l22
6iMGY17wk0wvYcq2Y8etwsUPzXJF1OfjyXBc58pA5IOn08GDRGrQ43Tf8Y5R7naUWLrzHZ1k8R1B
QdVCUMBj9vPJ+oOlj9xggD6fYr68Ov17Ne0HHF1HOfiGyAIiEn76GDLdDSDFybrtrnFrHjC27zMa
6RWXAvUv15scvDI4ZOB5/3ZqPpfOJLTj+rvQUKxHyHOPV8FqOB84gO5gdnFjioczbUMCKKawWfT8
pva75/BqEvaXX4qIFwdK/Tr/lrZvS7m14E2ZsCxDEweYyVabZqVFrkiqiXir9xH1y+Cr0JIjyu4T
sPV6szUk1IqEQDWyE7V1ahgdv3eF8Y/l2Lhucf2Clowo2fzeY6qVSvbwUcX+Y4AJBGqd+ZUwulTV
6KdNdj8UKPoK7la5yTtqrlo1u0aZcG0hm2trmPlTS/VItb/xnT5nL80/Q9Wb7KyAFjl+xAORsbPR
Dl19SD95ZfWIbFG93xUu2nLknPikyQDXHi4gAk5/3+9MiBmjt4YKfCPIRzkFlGcj2rCbEVnSLxSU
A3g6zI4MGUwsuVn90w3vNxBY2Ag3DZ/VnVbTfnu4W+AGE7lVvgSpRsJw9ewKqRF9CIf96xrffu+X
1r14A/liKZtSrWk2CMtFDHGdVVrWg2o6X8b+BVeFMZ2itX3ey3anEg0kOKChUX/sXliz72TrgEC/
NeCnSj0SnHzDaX9hZgm51srukJVjqtoNeeHIoFBV+9TCkkmgv38hpSt0p1FjC+ZgoLOM9CdGS7Ig
9vjSTYmsZR8eupOTmcG7CWDSEaBLrp9GdM+DMZ4wamYtOKjKN5yzB2AWXNwmSijU1r54c60YzPCE
BXXKrltucPGYF0joqiDg8ecDaMqNwiV00k/sCQrJ5VwPligE0wS+zNzCnzhesBJ2YzKV2zQ6qQGa
yLBrf2NEZApFdhRSj90fjpTTbdZg/3mTUSZ5Izx+c/TzFq2hqTzyn8dC+F8zl17D46h+6CmHvbeK
CmIpv4KeGlzb17a/lGTGQdkHvK09zLdG7CF0A9eVAr8Z1u/Q9jTrTc4iI+N7QPxzi3NDjLMvegeb
CDPIfmHozPlygXfbjckjKtW9YYHTUR1x161jpBK7yX47VmodfWkt+2xxEGZx3zuUCx1RgLD8hsU9
iqDytMOs8PTE0Lt6raAeHyCpYKs4KUkkE8GZNg27eTBx2kZG8hUsovTUM3V/y68W9TWJZCnkQr0T
Mdwxe9xYS61RkDwYkaEbqZBusqA1DbZ6UYB63NeryRcbtaRJvYNgfvsSYGGbYrSrfsmPuG+zJbeI
3yyqK73O8Xoi9tWonJ5dE7d/jiM4tJ/jBCoZwHdbNRzkUMvXoHeR7gOOgDVGYzq7RYr2PFv+ueKH
XG7ACREjJsBmoldl7iZPZzSroJoQS0x5b3HrGm7KU6dVJsFbEaD5d6M8OnLSC8ZKMTeRQQxuszUS
mHt7RM/eJGV90y56KkXeGLyndlNBhYWCT7FTgZlBL0K++S4FOCbM81PkV0P4edkNBV0lCmSZaZ0T
xxCB979NcUHg2/I81/O0uHg8Kop1GociRQVWLGrEURINUJIcSGzBZUtUFxAn36Jqi4EAlflOtTmc
LILtWOa42lUONVgGAOff+Usa181qAR6DcV/S8+haY2b4NArrLtJECirEqXNR6lcdWCLAFJ3x6skq
QKO455Qv7ID7adQuSffLqgtp/l33KMWNJH1Sraq5BF/j3fpzEIzS4c0rN29oPvsLcEZ3ZcFQCWhE
Sn+PKWN9jeAmG+gKREnTfLAkQ1TtZ6HL3ilea0qRm15TR+4odv6xkkmoukS0yAXvt52xHJjMORzO
aW/a6/uxMzaQnxecCq90TjWYjISZzEMibGxMl2DUY0o6NCg+RBI/7qANIeE5+Ky517sVXdunNim/
YfMgPA+HWaOAXMJp+yrO0MHJH1+QL5VSuQ6AKxyCO/SW7WZNGIVDSmqVsV6FmdBtRR95pOTCtgQc
AGfFPn40eiuwSWmKQI2MhX8O/sZ+CwuCUeb6wJrMnqh1Sw/HjvrqQ7LCPr0pK8Lohi3mZ2D9DoTK
VUsTmWGojXmGh2PnHGW/xjHtESwYa0J2iHCdOJanAELraB/WQYgcriPj53D5lFWw5af+U8ok1134
7w/tMrT91o55Mbs5CaV+UUgGuDcZ+Ze20S6c0HtXvkUFvrQb5/HQAhN7FyPV0BeoG6e8loZo8qgG
//bi95UkQrE4sJ4RSgCYLETJysW5xHSLaJzcE+LpJjO2dFWl9qccqQxJrVremb1cqWpgr1yl2NYl
6G0wWpV8DZoeDzY0JSZdvrHtQrzE/rDq6F8VOPWBjFOF0x4e4y0KEyhiIoGK2wY0XRQnqqCYOpfW
u6OVx0tDwbO7/Mz5a0rhqlFqHPUVZ1+3nF+AzwxkhCf8XYmZIj5c4ihMCDKwo0hcUeHZz/Et8kt8
Y7hsz2Gmw13QZq/0vFWsW2NyJu338BJwLnO84w8/vg+kWukUsVme5QMHR/uMMAALsNJ+kNpoGq1n
p2QyOL5VLdxq83z7JrSDrz4vfcXgFV3cW0wgGSGcXcl48E3dlBtbDGrfnJH0PBmgkI1KMvPF1IJ9
QQR54pxYp9a9wfEXbflYZ7AqKmWjGKb+Agy3/9HhQV5WLhbb9HJR9JEdo5h/B0kkir6ZO6okHQsa
Ea/Fui8WaoLefLC5ug5WCGeyjg0brPxWA3odG/er+tkg5OLY/YjH1k+2y8517+QBr6TxdnW6huKX
THewyqRAeW8nXjdgsxVlBWSTgxZQ+cQWJse+y5wGE2CsiNckN1pwLHMKxloO38CDAPe6iJpqHRXo
WK2GdFe2vqJKliMfWhwa0+88WeMoS2H2gkdwyRZdads2ELnQHvHGHzcPB/tuTRd3s1ojkvW3ApUG
zd/uVlOSJvD6wr9XocnJbS1KlzMWbKwRT//2PpGdUL6ACX1zkG/Xnez/Z1dlZu6VLVaFrZA3NzHF
50BXd/RzwjaCEPT3bZofQvSTDjbEiB0QiY8AqqVjHx/lVfQ5QT1HDGN7wSHPHzICC5A7Cz3bvyHj
jFyLAJ0cav6WD7rs7hFd9jPB0JFin0YfyCEeKIoUI519tohisogixrkum9+9qQkuUqZN/NR1NX3I
HyrsiXCOKsFEsF7W0QKdpuL28UuFtD5xmazSKPoia0RDWx0ezt2sOhQAfbAiwmloF7N/qB32Sz4W
hjdkZmY1SqpYs8EDpkUSbp7HmhiZzCPp5CA91UvyOEh36qGHqNUjYGKWv4Cq7IDzujXQTQ8cjyUI
X08hTyj6sFLcT0yXwYdH0y9+ph8nqVhyvdS+alkgJf6NoFWlBr8Jh2ly9oiUCFCooGdIfWwg0YSp
Ao2kHbwhfYNVYhyE3ZHovvRVKkbYRCH46FDNh9+GWCQ+z/YItbUhoh/QJFzwJZgQoSLEHe7uokyp
CgeVVHOThtR03kZvOpLIY/c1o9jB8zkNvVMPC+D6mltWfOyf6eyu4mUaZV9seGVoubwXQI6lBisL
74B5J/O9qYThlcK1VsDtbwAB/SkFolgd6h+rq3wGwqXfoGengiT7CU1fuj6HVnyxQ5XMcrj/54GE
FPyeTtpjdvlyY5P8gRbMm73TZsW5gSbFVrmkdk1ANaEW9oubHZOUrafs2DoTlEJ4lJhVWAQn/3+X
L2XgDQ/lQl+HCt7N71vOjdj74DEp+/LyL1ehmv0NkfqJzIfgXdA/V3rD2I2mlObW0vAV9f+hAt/W
6MNqA4C+QbFiFZ8fDVqOIefA1qYbuumsCb1KsbUUCS650vRVN6XF7K4aS+aJHpTA8v+/MMTCNTuA
GeqDNnFpKrNffsuGqmbqm88AuzLp04a42T4ItLZRCzQNK4XUAVapmeSBsrlm15Rbnx9gK34FC6CO
WolEp4Z/U/K2eJ/7CbmkodkYYEKEdFjRm1J5EE/6E1aPxBNNbNaGaWEH9qNkWhn1W2XE4dHOHjLu
bFIBKeI5jh8sTS3Vq68lKCjigmiXE1SzpnwFttuowxZ7yHZUvrVY90bTFn1BhnjkJhavWM0QkbZ4
gvkAfaPMfKrDgqn2K2kPGWSKOXWzcHlniaTFoTqXTqhZh/+xlr9G4dp9pPRfswPC1VmB+pYbPIZS
fZzmpJ3HOgzhnCcAHUWdH1zV9x5MwN8Xb4Q9u5bEHIrM5hs/HeimOwYg/PjiZuRls6RH3sjZGDkv
V7cUPS2TQvx+qxqAURCB+obMRNDB8rPGbDe/agCTdGkhPunhbWaEjqBKT5EndgSLRTvtPAGd+mrM
4nXPxOl8MPEjzRnPulbKtBjZ4Jd1gBNW5skaPwDzt2cE5F8orSmozyFPEUEQ89B27PRpfCfdhXJN
j7Y2OcVHtyytvz56fWbf6eii+csbuSp7WTVCkFFYFsNHqdp8PV0c276RxnQ4ENCbsqmeVomFmGsF
KtCxG4aKAon2N26F0+oRjn+iVAT/S7L/9VgQ5rlcKEQ2AD7Gour8NDTpeyBcuN8uhFF2mkX+ZFOx
7rtxZjz1xZuCax6l3NpOS8qEBC8XZlGPXbfrZuJsij2D4m7xS5u0QiBxx+UA1BkT7lfc9TPXZLyt
YyHrSwsK4BRzt7e3lhxQ9VcVD+4DBeDx10c2iQQAO1jnd5i+MnC3PhzkXA5RsNxCOsLTGQNRm4aD
FpO3ogjFhUbUWBbadeqKZ/DW1uGokvJ87TQmaONE7u2CXp7LufD7MnQwbvRCYM8NZrx3HYwTMha8
Skkwf2/s7RVG/T/P368ZGhsZDb4Hju3p9htZCNB5G/+/xUmgf6SIVYFEp02iIdAKfjnL2JSK+FWN
nFYTaOwRTJCcqv3dgDdgEa6SCezTHmRiJk5zksQaFwOohPauVfJjtdCxIxSjkJq8yiX3SJLIxEZY
AneSxsjFBnj4z1YBld3IzhxgAhL4KtfjGFDK/qcot4uSVU9gm4GsD9M4TV5VV+C50Vf5pgoMAJSY
HgBjIQ96hF3lIMz11QvNSlt2saBON+k7JSXEStGPd8G9pkbqQzGV0i1uQ35pH+6j9bww7nGGvw7a
uO+MCGiZiYHdwD7UioAGpKUw6PAMhZw4fMSBySBZSujUgjDo+usot+pbYAeZXNesIRiziNvkRKni
TvTzPzOCdJjBs0Dq2w+syfqfVZJwB5dVK3UGYN8OSK84OUDDsQzWUWe4GW+jzsk1s5pN+FNv/nqA
L+Rk4Q2yGuEl+mUca/x9wmqh5eSyJpy5oI7amittfFTifwosqOMTOyPrEHCj4S4oXrm9mKP/6lPq
rFietMobTcLoLGqtmse9LNE2arfd98G6sFiAG6Z1G1PewYGlLkWoLXH334OQPHXAesIxJvkLy4La
IfacFXgDb9w78JldlPHJKMxYRBIe4iMhuGiiMKBC8YNatIV6xEnFx6J4GysR4B0+ARGBQhjZQ0CZ
QfEH5nWcY3nzTab3rkggNgDZ7cVbblvRoVOfpmwFbc1VmXlFkbVMXgYyd233OYJSW0cJ78WA3mSY
AybLfGGH/vPJvAx21H/z67aMM6GpmDCoFfxPyHo9cNX4HOehmjeYJqy1M4tQ2YNwwR51khI9Oewb
657bnrjyiXhB3MQwRJBAKe5cMAeK0Iu45Q/PzmalvQnJWT50loYhFfKGXaUpLlutGNjwawBm+aGs
ZIkn44Z7oFmG3qovwRtcCIhAWjmgYScDk1EcnNNcRSqrPoDsaDzx6B3kf9L4ryg+d2P4OMfIo6jQ
/h/C0nEzldqIxZpdwtlsXrlNMuyzU1uPLCJwQMyrhT1CNjAWf0HNy5yRR27CQXtYookRf3NxZCY2
dB9An96cpaUQ+bdAEK3aU1NnzBowG78PKKc211kT+f7fAuXBN8Derh/fsddA1buZJzqCWJghB5Dl
yBZhq9/zL9abMnuAYwixP06IyaSF/X+41jQFx8YcgRT/BhPuB7Nuqen3YlEz83zuMU+CGAIKGhTm
prx92u+VNAC88Sn2FmRJKM56gNnhPOMUrCuGp/i2RnS9KDFwObFX0MPGls3njbmQMCerxmOStK0/
LJmYJq3HMx5XI/pBULywUjepNgD3AogJxSjOGbEzI8YP4nGNZWnNqROJubzM2F+fmMy6cduY8yYz
6Gthgd3wZRwg7ghTMT9XIeycMkl4F+TWxrOJ6XgdnYJt7UTVHgmfbiw/weFTLRStuDC5iR8McqnZ
iTcIrFbRqymcL2wwEHyILM1C/DcIk5nVqGMA72mP6BYwmJqLcmP3PVEiFwROe/b7l1y5rw3bEYR/
Fnj/utmc3c/FCohQf16rZz1Zw1BHWKM8XbchDVPGjXVNPNVqnbblR3NpqXivWveaYsCICxycj1WG
I2w8EcVSbPjkGDIK6Bv0ipSkigiO48VEQz69OG8RUzGcbe9LobUk+DtHy46ryYdTayRn6nxXgunx
3hcwfMlmswGFG9SE/d9mNiRSoZjqBY0GjYiKtdKJsEECKxWRyfhACYNvdefOCenO5QeRIF+2sBGM
z26rnOm7yi7ePdsl3h1+t7F0PGs/tNp61tls2dKDbh4z3G6g9vgx1lChT6/JlkSFrXqvujVfrtFh
7xsLZ/MIncvszualYaTqoeyTlD4en5TnmIPgymAgNtW4Np+kiNiM/rIGblAdH5oNKMtoh5E58CDw
9TQNu0OYX4YEFT5WsdFr+AYVOgBRTLx4QrgK/tiFtu2+duVWPzqBDjmMOKg4ktwcDHFALxlMhO+i
XZpZRPXIxWS+2RicciwNAGnUTGJfRBsaSxLI5CB6hQeH2stQBqY8kckCE2RfwiVyc0+stAWw9+9n
LVsOjHPWOAxhBjBxyR7qhmenu5GwpSSEQjmPWIIk/CFNJUZi+Q+zQUFyd0Yrio860iL3YYy8AuJF
qYMQegPn1iDDdwZdNut2koQJ7c/nIOCME2QhCGK9NSjFq7Q7vQeXelnRF8vEqX0ld4qYrMz2/rhQ
rQS4x/Dsy1FUFoRGPWRWRMt8zwRxnzLGwLaU99hM8uw3461Xs5klpSkn2bqxMAllaGNslzatKYXl
ayol611rXzfsWkrAeaZDdWr77+CyTt/C0mq/KOgRU4DJ6vXxca9vFFuhfNPHRP03eJmjDyo7Wjk/
1fzy4UMQpTAH6wBxKS9k4c28P400rf5yQvMPu+g9OA4bcp2N/OM0Ns1bEiDxnKqbgQSsMXJ76mBW
doAVhTBf8JKnL/pCnZRR9Pe/3RPlwVO1Y94b6x2JNGzO7AnIBtCEzNcvWL0uP50kDKHZXmPTg5DB
VR8JMet71dZcGhCEc31IR/ofISG/NJeFT6ryac3g70EJF2jyM6gThcOJSXa9N+lE7iLoGUDJx9/U
X7zo/duwcR3A1GWzNBAEUAvUA7tBSnxn4Wr6XR/FyF40WG1Y1YHGykiXB7cW980IdVluDOzfcZFD
Idwdne8YN3NTdxWVMKds6Hjy8q1FwFYSJYJiQ79QJ1VTvrqtD0wVcSkCx5SJpCqVVsAo0kafvoAh
qCcE04bGpwzZzvWujfytVDbGxlg5gCc/xqGFIFOXVvuFP1FTTiRfqPW5tUS49RbPMPIe2BJi2iZj
fShd2Igl6TyS7pXAWVSKJk6XsivBHiQuk3Ocec3iTKuBG6MkQwVK2EKmw/RpmoTbBJnkAuY+ulJq
0019hMt5Nz98S/4TD6tNaCqRHDzX7vUzTNtsqpZNyK5p6Dua6FmQmNc5/ia0m5HLjBxOq6zu6583
n10V7wiv/JxXIvJTdFCSL7EOtP6Kh9zlkUoeaFUzBGjGqjaLiHj83K36Eq6gq/skbihrd0q0t+f3
DxJU7p1a8ENMGuKnGIYTiu7ii/9NFgNYkokbq5pxaZSnYSL99LVpGXgzQvD6ImlGpFpeOSbnYEiA
jTkxSssEPzbmrqBg8/FpRH3mORRnoKGPPyxJg6Hjr4FgiLCG0m2CbzyH9lizEzPjAZUuJM+fsxJU
51px2/fXLOmo2jhvzRSAn53K/36cxtSpnqbx5Z8YkrrlpkQi4GUFA6//TZhzEM8QI6wpYBSSpDRe
G/LkziYN3L+fNN+F6KpRvBL81gLs6I4HspAZceZXXE0TBHye8iuSjIuH2DjqCfUdJXCNiKV0ZLqk
n05A/1u9D796j7c3Y0WAIY4uzqR1yP6Bl0QnLXQ0F8kJhDRclOFXyXp375PDKBq5NVccODbur8L0
Ov7E+LwkoAE3ulH9jLUovrBEUYkvsh3kpJr4XiSXmED9KQCRosItvFtHv9jckSBz1nfscopvdSx7
zB8xv1q7XUUHkHRiHFSZLHMyDxH5HG7H5Fhq8omRgyeMPi+4vj5UQGLRBl62PBUxDXy8K8eX5zHk
NMH+tJFwJd2vKnO5ppwxJTOqCTMM550K0gbTlMOO9ESvDzDSsZvQLVty/3mnO4Np7plkkzGTKLXJ
B/w5dzlJ0Ptix06BPuXC5BWujAP9fhWp5siVM7zRUU8YLUyhti+YbT6qM9OAYv8w6Dtf28/qNxRv
ZXnMEPs+GfYJRj62+HS1S/jw6byggqkvrPhYnsN9bZwU8woUrZ2KoQa8oL7Fz9i8+oIcCsIFJeCR
b3uAMpL8DwHKSbxynfQmgLXXCAsGN8i/Uc4CA4GtKMYAEpZaZBLx6CkGtcxuUoI0x7M8BuMruuft
8VjrQ7sO39w3q4GA6CP/yDFQps/NIblPLIX6aSHs9ruiOM3cKqB8EnI+geV8BAkpPI3stsbgEqTv
tYOc+GYNe3GgeAamn3r5zmO8ifYZ1+Dv9nPNi6Y1plJdhdKK7GtWrzKltQOyvOxAm76KAPl4AJur
XAkZ5LKJgCf/rNKdh1Yz4XjSkALpYZ27rW6AxxD0clbaBetkkP7LRuqzw7NvoKr/AV80p8XEZ3Y6
x16Un8zy3rQbDkYzPyhsAdCviQH+NXorIYYqWW7ra3fOJ5AQ0yFrIXqIDPxyWi12XvhX/Fu0pCk6
35ALWVHW2GzDDfHSJFrE1ywqRGgHPKj88Jb1WwjWVDqS3IsSg6QoP8VsovG4cwCEHgxxtp4NvTNF
6jTm5M24ZEPTq7dAj23YsSaWpuMkDE+/7jwh+xWIB9vB3r96GoxxZ6OqjOh8EYhZnQNGWVdbE89P
9IpvpoyumdNgY6u9daZIznnj3MpDw+Ot0fTriKEYfYamJIkxe6tP2EtmmqQjsHG6ja2kW/D/e0+i
dlhYBxkRTG+z12QA+gT6aO9DeClemg2SHWPhnXdsfmWUaTtlXNXG8jAiWTx41thFeSTlaTBSN82+
fcSdB+GIwOj5a5hCOkXVgRfd4sNfEsQU31GvywnPWA4WxZMTs7k6xZi+hLVy5GlpuYp9GqVCad8p
wyPRhTYMmmHbuYRzIQnHJKClMzJl/fZFPnyVuwzUShWaAoB9GhS9RFa5xJpaPHs23Z3ryR4Njf1U
ebZO+af/Mszmb41Y3anVDhl/8NSHP9kH+Sz5DrH7WXFDkEFbL6kY+SQZBlRdnzhZkwUfzjko+YRM
GXlMzO5Viz5cY+8ax7jclkxsi+4m9mWLAWHO+++OvCAmT88f8S2tmW6PUAHU7/2D37P2WEqGCHr0
QkUS+Kl+hEl67vF5iNIzZI3t0lLuGRom3rvV6mJaAHd38oZ2pEHB+iYfqseSSXVG1N5/oms+JQTX
GpieKQ2wQWHpsRRwyk26FRGCAKAS5S+EP9le4G3QWQ0qAVs73lLxV3HjAvpclzwJqfTCzui/z4cj
XUm6GWkgRdz72rtnlS4yHy8dB/qnulWbd8yosS3v//oGWi2WZgrw23hD8/IcInnGo7wMqItSNVup
DEMrCES2tzS6DQZbye9uxVWPUVEXwgcDe3d6BZVFzsvDDMDk0ngdC1SemskMyBx8KDAJKsBgTkpl
Tr5PTVBrJ3apvc4ecwrYflnB42lpVlgLpHphYtqztXLP1jxuT13pBOnCfWfjO/gkkWs3tQlxzLbZ
Xw2eVoTKuplfDjJob+j29/gfOxIpYz5aUEQiec3pMPHrUlSEPPfhvzakrQ1RSppqXqzACvpN4blu
6zWDrvsGr2LvzrGKelPlnCHeqDBxfbpnHemy88cR5LHtqRKr4qLwlgRofbOmPlf5ihd/12M1E+MJ
mLMUANh0fuLITjz9/otng/MJp/xQZNMl0iBH4P6u6X7VKjTrB13hJ2Iw5MWIJAIf6sssx3TyXSsX
7Autqt4OiA+J8PA5uWmKR/7lQRA03kuY2+hUiF64Cah23ZfyZoMCz6iZXxEylPoaWAotiYPAKLOt
TH8Xl8mD7DXoH+JbsWLAn3yyB9yVNSeUAc+e4p6HPtJBUuC2OxI7ZK4CFOEazIIfhwC83a/nV+Xn
rQK9ATvowZ9oU41G8RRs9PkR/WtPBKtT5OWEL4FPSFpTHo1WuQMphPpQG2gs/WzdJTI5+B/S36m1
fbEovCOpNgUzh+u4kWddeZLzpYWmp1XYTkbmGdlRZUejhvwHZS3LpaaLVYrb2stC5kv0C3Rvm+jQ
9syNQb2WS0prrNvUWf86KbzAg8NHEze3WBwmJBg8/p6F55K5IFDHbjWrsvVUjFW2802uzUe+X0b5
c3dFOME5gCqumgcLUhBksqLthmTPu98lC2o5A52DAcJTqJhIsirqOu+6TQx87WEmCwtHICHcTnG3
AQ1Ns2Aqoj7aHj71BaJclVN2MURX67AVjeoSTfPGtrmlMPLqWVQ0GmgXz7YpEz04vGVh5oyj20KB
SMF4cJzSRFOP55NrUBUFK9FV39XX/Xl7n2ynAyLstxmQ+bEK2/k8xhEgz6shw3M/D2c2mix3Mo7g
ZFoT/Yse01Li+MCV+o5rGiBHOA8q4lhB0QcEHN3Tof5O/keZZYcdC/s8IBWNtcLqo8pI3wDuWk7r
haXPrYM7flXeRzxGxs/zw8pd+ssAuhvRW8jOgfc+ZqfG85TmxktcOHrIBbc24pG8gQDJoPrYk1Gp
PqIsDGehQJoah0xfmzRnyJHBZFZGF/3u1Zr5oJdmdMaLZEr9o36WfwhoAfl5oIPEuNilvEjw1puo
7NzbJkA9orUarJN/aPUWxkTPBPjyLmMOxEd5CQ0m4FhrNkaGEc0qdAWGJaV3cWBgaFwl9oz5/ID4
ho+TKPxl4HWM4G5RZTMbyRJ8MGImDwuq+GoFe5Tf8R7i11o9WrGLwCFbJryKwBikgYPEZ5BXzSWn
hKaaeyViQaTx6It00yD4g1bLWNb+ueTNOJIv2AXmkqzomxY5eFcOtT7kxEioHPyeC/DgVYi08cFA
10C2hbGA1+QFg6Ws6KAFi/lfAPrHWGRmXGvAdepe4xaYzuXbE4Jd20K7LY1FS5Q26o8DRMReucSk
6XgD3ZF2CQ+3dEu040qKIrlel+wXP19z3vyIlIhTKzsetGKuSfUVLUtxFbiiL/fVtL3n0knJY7rD
Wf6oAgm8SNcQApSzQR4RGKcCaEWng+zv8PGlQDQo4aPtRuQ+5Y8A3r0j9f3EjjbaACSOaholplmm
OknDivqpEckCJ8+OXmdv94BXAJsyGcqpueSTy9RTUareY1EmQJ2pHMW9a+FNzIT2cuoup6nFzn0M
fYoJn4cNZsKsANai2bRhooEXVMQHFah3PKiK7LRnKcCYfQDRNvaBLLd8pj6nu9wCNZxudaMjvn6o
Fg0lH9AuH1p+xza3wvdybacEWYDV3/UiGrTz9fBjwCq3C/5eIZ0C2VipKViXfo0b5UG53dq9mzpr
V+UQtHpYnDCNfN5cTUixl2bvfd40cmY3gm7CIoNfUqv4VLOBLUd/QSVA05DnSwces2xkeqcKArs5
PIk39ppFVfP1t15tIgzN8tKi0uWO32wJ3qzXwcPhDxcYlqO+DzvNTVHWTWgLW71hqC7ZLSzxdWS7
qUNt6uFE0mHWxgQJQ+V4L/dWArsApnlIzLCFZc9qrqQoVMLYGIQcvQFJCls2uFCu8o6kvoaPiF+8
84tppZ1m8uY/Jre4UaOmswps9p4m+FJHuSpVd9XuPc/nYNSDfTqEUfi3TOwYKfmSWGU38IICcHDI
gpNf0wyqVIe4uRQPwX1nBYCGdB18XEPMG8lQYCOYU3M9R5PhDJVG3O0przf6w45aRyqg4BR9zSsi
VxGcJuwl26W1IC5z9S8D9W7YJEozy+Iloyetyrvf7zCRg/ICZr48Xx7ysBVq5BvWipBD/YQ+LuZc
F7MciWAWfi8s3MZbiDXQjYrTrKJ6Y55lEJdqt/mYjvMYgp3lpkPwjDh2yywfzzj0Xs5hnEHNVxEG
tEBoTDw0alndjQRouQ+2218L4aCqNsL6kREcv5a9naJUVFkJJeymcT5Ktk829BGEinLCq7t1/WmW
CvymXhgd0OVFrn04fv2r69HvJH6ILK0nk3CcZxrQuRKzeqFSq1E6FKBWweLW/tFY/B8tzFZwuea1
GLViz0PuIQ2Q7cub3b9YZud12yPnYzqfYrHDJO+qFAeEz/045v5GorESuyjkcpHy99aAr1aVz7nD
qzmPczvvA93Eq7mBSYajBtqZq5ex3t9g4sv5G+a8uR2C3a4l2T/YPRNp8OoXfz6R1jZfK6EYcp4B
I6VRcynbFfnA0iXMZFl7TOW4A5m8w5Yp7++e0Ks8+01HRvKcVpE7fqHwb3rKyqTI6W+mYsnoHDiV
U5LFf4o43L5U6romtmTxEPNTtQbZx7+/tMhlEtMyS3agkGVZ3tqp8+mwRJ3tWHI2FCqkSHQ0lU0z
D1en8VldctqsffhYih1IByqiIKvRCRuukj2Z1j4zFmPXgt0qRDm/kJv6U24sajFX1vM/9iVKNJYP
GqAkl+LHJ5txgvAA0r8C/n/ZMJaywk7KHdIggeWGCDigNROZehY9y4icbZLXSLPOMIUyeZIGa/hv
B4GJnUFsFxfpp+gixymMQL4VTmyp5SVQs31ARFjKsk420Ogp+nyMegk+AmYUb2+crmJzgos3/T0Z
5kv2PoEF+gVYG19CETQ6jpQMorI5YyrRTgPy9m8Zsn/uzUHDolVF2CXZu08F7Qq3LNTJZtxgvVmq
pTRjga4uhvV0rcFE2im7lyvg3dSHiGTP30gS96KxKy5w5CKlEt0/Vr8NDU4HVqTGEZXuSm8xS+9K
+P9HSbxKzQhkDcZLJcicegsp2CXG4idIuiV0AjibjE2OrFP6bkWiTWXBSeuy7oOE0bSm3A5lwPcY
UsjTF7E2+p4ISJfmJ++ld45m7csTOtOlgW8ppTWRT3z+gEwcbnaMPRsa7oBEHyHcg3LMV5eo/j5r
nhjxLYQ7BRDh0Hy1MzdY4hIYqZr3KPc7OUakHfuWtJqIlHoTOD+z8BNTJsLFUerMa7EkospCNrte
LRcP/R9AmeXKVHGCVnC+V+EHBoA9iVgeB2ghcg9hyRaC1UxvO/GJKm0JNWTyM/QpgOYPP1HGE966
deiLYj0Xtu7qb7qvjye60hf6rF4PYU8rIoc7GPhAPgPzX9UEYcn87AwtlNAiX4nLXp6hyhLgf3Y8
TZy4FHdMB0Cn8HOamMgBeDjDPqs9SYb+hDC/3zaHy5W7p6/TS707+UEmpFxjiI+SPFX4VXUKpf5R
OQGpexF723I9bTkvodUQdjGymmFaTRkhjpAIosK0D4Fwr+c9XdkloPZRKjeTlj0VRa7dPmBhKM1d
9wxHgO58CaL6heW2UryHwb1elcDvSvJxp6aEKgwIS+IxqEWeLR6zVl5mRzy5hJZ156Q2V2SNY92+
YLkWF1Fx7fM/3Cnmv15BxmlfSTvoE/022k5ltTO4sLTXNSwagieobliq+5ESsq23QmoGEsE1VVLu
zNNIoZVNjgJ8WJ89/d95yKGew2apucQB3f6JmpG9qCrc3CuHTmYKvCtn4s5ITKOmcl2NRgYWeCfv
slCVNRucyCHQjlmVGSxmjuk5KjYNv2nVX+f4wDOxbK+EjqnjRjsZM6Kb8YUaO9pnGBIbaBA2xIUO
UMpAP2i3PCDS1lZirXwytDsFP+06bH4+I4bsuiHtjt+pyMVR0VMUIMFZgyq0/ABQ5P5lcVz0S6Pl
y+b4F4H3GSKJst49FoYuYvQxJSMaY2CCr0ppt6tCtYmSlm366N2dmHLyjp4tDbYZO2CK+Cks5eI1
wjFjEviCIR4RD645IVps0Ovw5mAqg/9+pGc0YvjRkAiX36tnqX27H7O69VXXX6kAiOgvB2VnG+ZR
cAQcsa2gcZyexTJUTBW0Zi3Lr+9biTsiQeSFFEcOkhQqDK7eumv3MckGg1tj533eh2s16iuK6rWK
F/uvpDs4IXWCdhfj6fdcnO/K9qVK7oQ3ldSnWmhDSXa6jm+419iGqGld7dLwJMNkzV2wFxqM9Ekc
fh6WxKb5gBk/58+sVK0IQEaz5D9muhXDJ9rkPhfNjH3Vjzcu8nIAaYFqxS8gXsWEBWHE2vcbLj9d
ZoQRg2P/PGeg1TFjqLCqw1raslIBJ50JGBd4No07DabFpMTIh+5MELelnTQb8u0DC7F2HEP1WCQr
uLJfnOi7yu6vS5l69IQ5IxCZ4NXE1aYC7j/W1QDfC5SyV9HXddiPbFFOYFA28kmj0jIn8aF6mLhM
Dofa9Tdrlnj82Q/QrS0IHYhU1tAg8NZfa0R3G2kt1Ru7ypVw6pkeNH12XL6sIlx4VAaXj/iZGVs+
yTi8+dq8w1ZW0g9dBU6/tZ75UunEvpDIx3QhzwvgyMYxBbZTPRS3/unL4I4t/aub/vlKUbh4fCu1
qKH6Hk+IDN1XokHJgA55AJ1ttMWR1eRx5Bih40skSBaGymQZknA1N1B+AjhqPVCgKXUfzadERL3n
O8nJhWvcBrQ22a9CiWQZVELZ0rjdCsrmfLjmnC2R1HeXJPUT+DZ9qvtjj3vQwyQaJncN28JumYtV
m9743u6ZWzr5WHXDKg45uS9MvUCLGxkYgvzC6kjcaWL5Fgt7Z/CaUFy09hKprw3VHZR0jqPIwEmI
F4vmNQhrurPGbRY+6Z2QPuB3X61qTptAuwtw97vMBfeJ1eXtys1aKz7Gf0YsfIyeHiZcPzPTDAEo
sgsfQ03cYRzsVIdIjVKtZK8lGm0iZ/nbvkZQPAPCS6s1pNbul3njoeXfu4oj/tkz/ZQwB6qzbwd9
moU5tfIBJRbtTB9hGP8J+5Am/MDF35WWBh3Qr+OACJl5UIrFrtmdT1C05ghWP/Uxm3sEdubFkPTr
d+1BBbKYx8b9EL7iM1wmwTDBuG2VIvCsE1mwV9cAu5LgyCivANF0pcojID+pBw1ew37tLjZAtv+b
k3bqjaeNxHnObFzJ/Kwi+EzEuKf/m+HLPgJDVF4blcsf0uqRHMb5S7Z8qJ1zbxH3pujieCks626W
6HcJg30itb6rGIXWh0Y9K+Nbr7Cm/P/Rol7bOjnZQAi+KX8BeJz089yrEawxF2CNq8wRXttQFIcN
zyT0FySPpAfrfn+xvqcDJ7ElrlNKNM7CV3smJiybvFH+Ro0GBKnPrN5DI53GZOPG7SldAc9NILRT
GENDD4VQpL2z7kskRgILVL7vZS6RSMFdgMujkQKde+hSbhM6M+of2jYqLbH4CvKTAHiLLUPY4khm
RsSnN4BvqQwT1r2NePVuG8G71kyD8R2tUd4q8n0N6oTbD7nSAPQ3qZNbSChQaw2ZSR+9W0lVlOFC
QWpmrXtvkbPx4z9Uc0AqRNVFkPZddo8fdycGEgljC14UhmOVNJ6uwbaWzSmibfVJPeWoqYh3mTgt
K67Q1do+3ehMNUrZMBSytLWXDb7l7Y64U1oEdd726XzFrnCx1fmXuTzMFxErRtk5s5RrcBLHr/WO
DoNlW8T06mooRubLYyEZFJyR8MJofITY357cvc5dAws5GF566FnTZa+bPglvykjzIEiRbEl9hkPP
IyBXkvKr4CeO2qTxNtMR9n5MeooAel4Uph6Uo5qXioNhW5Xzw3vu98zwLJDyYYWDjrnb0Wa85Bph
BpxpAv5FzXf1jr/cUz8fPWRgAXdtlUspuYXNNoBrmqNgLkfjoG0F5KTf3NR8io19ePMIi3GCY9i8
J3iLj/C4zkA1GJh7qmVWPYRgFZPEw3orDwVogoXct5B3kruoF7quNS0OZObdpeGqqbbQzRqBIy0o
A6TPW07nukJGypJC06aravAeY+Q840qlGijdt8XpAm3QJFlhXhnVK9eGSGr46LTvv8zLE6cbzgRE
/69Gq6O/dpYSuSOWS8UvX6qxFdEmbTwjOgPJqc5QYht+/DdolErmEdxBwryorfRbN0bUozH6spm+
yV2FRcCrzw3o9UpM1hnWwiYpe9a/zf2U+ljYE+pG3seh82m996BRG9EpE+n/sET/gNGlA6ZAVi61
hUJmVqR9DP7NGfbzRxnqmadyRdxGLxVk2O/WM99umcTqqo8H3ibsLUrlAvwziWfbu1QjtzsBOvn8
JgfY+ICb9NfZtPithDoW6BJ3Ogn1uLars5C+UGj3WVmy5WynBfKZfmblv4ilphC3TssCR+IhPO1R
6M0i417CTMt+bBAFxTm7EeM17I0gRSbWd+XXz8TZbMOihb/A2jGq0jf4qVLaX7RYaq8msVGRTX4u
Hm21PEnf1M2qaJlUAWJX4iDmwKuxlPIXUZ0vT2fdirMumxgdB7++3f+Wc1JPkAjLI2waXTTMETJN
SmxKPYOOBdx1gO/8CVpeYodnLtI4FaBR1euighkVF7di6vgyNPcfxNDxGl6X4gHUHl7Vuz7EFP9V
Oih6jlEwh1gi31VSJxsQMYl7ewmf73CQQc4aGjvC45n0OrJf8XuFdCiFbUeHPFh/b8CPE3RslB/y
stfJp2LolEvEhN7VO2DDLIX+b1W+1m849RcexL24i/ilnCIKeFlTpsaI3WYiC9P8I2XauKFFj3bY
Kq03DX0VVIqmtaUGg43PU9CJbJyz/T+ALV85PfE270GFMnYIC7+kKp2nxUrmjnLoBEs7OLJ02LHF
P3+TYjFY4KpM8zBE7WpfFFMGhI+xgb4CRhGqNAc+bjX5Tno1pZfTGdVB8BXkXxGpuWTBpU1bqZTp
et9vjXTR6UMil6BkrTguRGeRzr7ZUAK57uSP1uvlNx47/S3KU4XErfyGzddj0NJczOgQE4BR/anJ
5a7nLrItH+LsJ1cBaZFl2cDXNx7Gn65o6pQv3p8SumFwlqGW5gZ29EbIrq+UQGaV+NugKgamBkKD
bVhDuXQ/c+MHD85TlRxFaiCLzMRTaOIXptzDRvlE1xSu/ngnafsZ/xq5037d2Dpa5PnPxwGkW++O
/5UKWYHgwHzNwD0VKGn9+b1VjvZjjzc7/SCDeS6QjN4UGcGTvRs1m4Xq/vlZP28QCpEidKzCO9hb
K/9imhbcqoJKW+bJeceUlfzGXAf5hH/TSl7liGsGGo+xdYE7zSpE4M8AB/RgMl6ue5SSZMAw9By9
j3QMNUwxysRTy4JOo5+JdXNgrLO0bimwPxpI2CK4NK/QLgQftkQBUSwgiJmZM3mz3tZ1i/qn35f2
gImEFlxX5eteqvK3Sk/SrWb+tpe1u7sdHxlcB3+j6T025vOLiyZDPIL/I6aB6973fVqVC/0aFSx6
p7CpO3aC4e08XxkiBJPUowH2bTqAn5SbKGeL+8fQJHt/DtXvyp3V9gOheJXdNrTh6EUSbveGvUqn
OOsVlMVPc84HTiWjSdthYW8foAS5Xa6BuoWCT7JBN895GuVmQ01R8qCftr8IL7TqyNIcqf+xinnd
K0lU2wlXa7An7io1Osiki/q19G96K7hWfwlps7HfLF1lxUdzdUu90EKNTterf8fGoL99kFeXuF2L
NqlKwDQOPe4JyAY4SN3BRCCBieD+CrVOfWQeGP+pUEpbeH6pGVVmpM+TCTq9tjPgFb6JjtcKF81d
EZEJc3TdbZDs7+qj5nGttdXIkOcZIz8s2X8+xDjozUP7N3rKr4x22rpegQJhZReN7fqG0pAUxw2x
VWiNchPWTXl+Q2QceSOMw02f5t+jRiNSG/XfzAhrvzge7fEUeAn+NLeEEVQFVbGnvc6hxRjSrhbr
SUE+RAVXzUY+6nKsWZcKlzwBQhNLxODZ0KagFzOSB2nELFqVJP8A1tD3j9V2wBb9nUzEETyyDyFi
YyW+c3aAslJmfDnoe7fEJry7X2X17d8G1F59ColQhtu3z66H+xqKj2Btq124uACLbbdkR8i5EsND
oukGmhL1eHF68TC/O0aneWpzF7rzrXZX+bR43k1mmFoSqj71ooxEV0XI4mCKrIX1SH36QzZvX6t5
fqu8kRhM9ordwN/BaAfBKMoJsdjhfeVW4BusH1wF0nylLgmn86hS29sVYdpDFM9ebfGXyVMkETaQ
GatZdABOVMiOFeaIIMSipl8lJqc2FGQSeAmeluAFqsGNfheFbBLSD0NnV+v7cPhxKKM8ortvrA5H
HR0nvVYcLKyY724zmvEIPtsNCZiX5hJCrZ8iXw4AuXwX/0J+aH1SeNNjCLOosn0fb8LMCL2CfNiQ
iSx0CwMrgN/HNnntaHYV3W/V88FT0u4+nFwUL/3epanLO+a38IJj1NsYPgtoqJqify07Fo/o4zXj
RxUUOcelqa68k8fqipBvuGRE7hLFg18c4lFx+NSDXATjB8UxTGulSoUbo4+kUerQX5ixfloj41zG
kXJOS2DUlAEmdGs6OnCV/uVm5CUYXoUwOjfvgksw7J7DcLDyK2scgaBjwq86DjfdhUhJSLpNMCKc
ZP/6C/C7gBJZKXOqh2FIs9DEcj10Awb7bK4vjrU7qXFGlG7IwCQhQcYpb3Ly6eOI5eDHDKQp+Vk4
UALFikMAQGyA08x8+Vyk0DT45VwcYTZEsZ26nuPrX2jWyIZGyOWmo6mz82l63/ufDAUWQr8EPMJh
gjVZLTbc9VB3EmRELTjGUbqPTZEWCDwKtKhqDepjz3O3l7bkcn0oDduWbbyVXxSX+oYGketDGSM4
ihKGTtK7f+Y+ZYtoAW3Y612rrNhO1sWR7ZUrEsLeZ8otTqWIcR4+DX0BlIfMeEukq+HeIOa6Dpqt
TIl1ytIR9GkNVtMd34cemEfzAkIJ9Ga+0aTDwxuk1iFJ1XFtcGvF6c/XqUxQLR7tYGFHV4Gx4Z6G
oLbMYjBmAIHv0OVnY8FzqIi2tvNUePSJbEBtKowy8cHZddbSALjCwBSAyk7E1er5+zzKc1lTnfHy
hv8utFQu/GAVQW6E49yOjl/qxkWQbD0xBC4iUaDgvqSUME9XbLbUqpd74vDdq5HmAa5ROOrud0EA
m4eqsJIHJmfIPwPR2gFqZY2g+mhp6vQ4vwyQV1ToG4SmVoa/Mnafl/V7O+zmaVUPthxYTEMPm698
uDI4SHlmGAP0U/tXlIoL4f/kUBRFyzPPiF33YtwpbM2cVBPWNdtN30BGFIng0VIMN9w4fYO9rEH/
fpRyGVv3RRfePyg0X1Y5OfCJimvqdSStH8EARmHa3AQgbhLeRJQWTW2S46ClGfw7v7V/R8O7dW3G
VR1vaNn1G6tkgVJQukW+4iuMjLoI5hi1D9NPFdjQu2qMoJDiqe2NAP4kU2HPLzXindc+aTyVZ4zL
3tJhYtekIEMSZx2BzaD+HjiOVNl3w/V7efvqNZaXATNvDG3hEuDP2LS9zM4fjJFqJg7QjihbIgSF
PaM+bbA+lJaPvsGSES+8w7ADWzhwfXkF9t7ZCNdihRHBQWQ0++QaTSWOVRPrkTsdyDbwHtB01nyh
2FU0UEDtgLO6mgDtekrWHpW5Kumxk3AkUVq2MATw1/4CrWzadJFFiABgMs7ParmtKwSirp3aHuyt
dfY9ww41iSCpTb6UqVSymNRKgj73VpoaG5f/Zv6gsn0ET2VxERJasjTGAWSWxRUvA9L3h4snOl1y
fwzFmdQBjCa3o9DX/TD787s8+bYb6yVkwaitobMekmL1oh14+4amNb2Z5O7xYSYmvPaY0EluIj7L
0iDe8Yw/oplxlujJmSvmVsYPLcgLRY+vvQ8VL5vCa0dfXBgAzMDDvvVr3CExizWbf5sOYY4imdmM
pCPiC1qbHD+yQHhapSSaKpea7ap3j4nAx/zQ413b+KxO6+QQiRYV9+0mK7nQ1e41kTZz1uMM3UTI
fqJbCCzMRGD27zfkQHuYnwAPDbxmT0AIHgOBQa7k2rhRWt47Rn0Sy8E02k9LVjQfzOLrOmmyXBR4
N+jKm82FDjfwwE3BnaLp2KwXhWuyd4um5Kf7U95mRyOn1cwxnDM3h0pnRcyU28PbMhG8WR6+2Xiv
P8oSR4aGi6aA1i+9xsrZ3DTmnJO9vMc0Qw4esioJH8mM8xuF9iuZPYQ9DJQSRpfYVqFMSBhanmJ4
3lcxYrzZBcvpRgplDqbK8cs+rS01JaXnjGz9zWjpR7wg+0x/hoqdz6PTw9Lit0XGzNO7mhSga0Cd
aKuMV0GLMNpQcVkMkcuz3XzQ+jJyAgOvVOWqdtkLJ85BTZ5DOMd3lVW5Odwsvr5qaq2PdmCMd54I
ORft/JHMlF/lKSDQixAkUvPzNOu6PpPhNWHR3XGSBXdmNQNMsFqPExXFfM/9fwLL8YOf0YPgBa8+
oeHFGS3ceQwMECvVr3/zH76VDX2IEBcvAvsfcziuPSHDqCtSo/nAkTDopyjf4tGFNKTh+t8HA6QO
raOlF3TOfDiyxV79ML47Ouxg3LzOmwY052LFdTMxUimS568jwC49rfI3Bcp054qz6ktGivlvdUjj
xSI/Rq9KScKBSuAKuBZxwo9Imi4blYai0isxWJEszcbl4dL5Iv53yEAeROvSIrAQEDuXdJJ4rGJ2
equjBtC3gEzl89KFfGkoweB2XuChA6WOdowm5y0VUD7wNloMbewca9RdNKJfLxLiUN3qNEKp2eAn
t1UoMRGzDy61Yu4cpjmSc4RlDgqmXQc40p3U5PvxBW2QAFiX5oz6scogT9LEYvaTaXY+2e+Kmvvn
IlkG4GI89YVYro0aPfZetXZC/UFgsHLkbpZSGN2D0VXC1H+tvGsv72vrZuDpg4GVNWF2zot8dTHk
8hbdacNkLdOSHjn5TAEv6+jyTIkWM1xlbIuzKbQV+EJ2kLF2amsSOBtXzaTadY+F3zLclVNkgGzS
fU3UXWcJ1WrDeN5cWupQAh68INg+apmcmlTX7If0TGoiNeOgj5FaxO7RpkLzNuJDm9xEiYx8fpDr
RD9aOPexCkyhs7mzst+Idyy17y/kYyc8A0MI5Tgd/iNx3/VxmABB//TonVyyaYzl6CoFNqwf/3hz
NjSxiFskQtGgbLlwDARXjSbdL5+EkGCtJXT3Pax7Tbpfq4F68iodM/0q6Wgw4R3/H55tA6EfT2Qy
2823xZFIQbzgnELEGc1z/4j9iKmGW+ltFhapdVT+2jB/nvXvvQNavq4dHSAoF2ZCNl8KrcuKr3SD
NSeYudI95EN1wFjhnoXmQNkJ2yEu5A0ojcR1DsR2HL4qIeaTkrPdNJQGRhslT6EFGB0kYuCQVPpX
r3YbiC0Evelxc4j22ZCHMZmRwZd+jOkMvIj38hRGPqj9tjImohMUKW6XhgPMHP6fvteveIl/SpHj
D0oE0JkXzzuXUDWWEZ473XBW2+lavaahpjehFZ33JuwZ+WBB1vRM5DU9/qAMRuOUTglwCCry0hkj
7lOxERsK8tw112oTWhL+vOFDEAP9dsgitqI2XXtN5cA7SumvpQMteDy8a0EUfOtLsunnh+nqnJDM
yhWvcvgYSVH9gepZxJGkIbbMVx33a8r3trBF4nOcqjTiEJdHGLKlZ9bDXE4d0rs300wyrnGRi1U1
3HX2WqYrn+YJo5PNIBMpJKdVuO+VVwZj6MHthZbN6DOoyRiJJt6HWnguG3Z1HEmiEwYE8mXzw+Qa
/K/0M49CsQLNG6HmacuC7Ji5SiDfVuABj2Q6RVCZY7KNf+NF3IbDMKii0Lwye01wUQGAq3ftGaYb
phpC5AxJr993ooD3Ne/zvUlyxnQjwYTsH7BpMA6s/hnrM2my8rjfIrm08ds2tYDGqr/84mblXMCp
5xjlRMhObbCyqXl3r1JEgnioGLpCD8tPLer0Ivuh8cSWOuEvV+mQM4AdhWrTg1xYu6oIkSyJXG8x
lFJtoUMEHaUOvqpRXXKb4AldTW0MdvtvhHnwSBD/gXlyVRDYN9YDUOZYHMhRuqf8alCpPFsukGGK
iQx2mlK8PiDZ6+2re99B8LaiOY3QHGnAuNhtnYhbugLHx3ZK91yFY06EsdYyeXj9CeKZrzGKbRX6
qg/6yEHADDWhx2iyy5c66/ANpHEvkz9F24bxxyCicfb7256BfKZ7I9Ec/o+0q5adQAKC+UEEU1Gd
awuahfRcXEIhQ9KMmfGqpQolVwqvFbsAOM+1LkcIBjcsHhsUbgBjGqyL0NImA5N06Pi+WdnYE0tn
ka4W1tg3SiswmHjdqn5So1qej/oBLygvqVN2r1FkPumL7gubKXvPotKn9X7c6VAaDOdcQXvZKJ6+
QF4RllhcfcKKiZAPq15oWx6pNCViAovpHsr8lb4EzgwFA/Zc2CJLFZwG4wwVDiJYgL8vE/A90TKN
g8aDgrwHkwUGCW06RZeyCA9uWu5xbrn2QE6tdyEPCmXh+SBMHFDo40aS9FpeJX2D+X5HLh+F20wo
0O1Bc4ciTlF8GZ2SHFzTxBlvb67mI9NZ1dsU6058+21Vw1f5NEKpePtNzIQlQ6U24wcvABKOCc1I
OPMlKEQ/exf/eMEKoH3q6sJEhElG3vMrVKggd2GWpVMg50ev4G8wYOJjdJzH6+eNKe1w2DknaISW
iJv1JIW+b0pxUH7M8FQI6F366BUttdW7je8rfBG78JSTMEGi57wPfXkCwe4N5z7TkJHqx3FnhkTd
+MTB9HCSUushfroQHnytXkc4I0EOZ6H3JvX3jMZGD357+E6Dobq4epo12IMGazyanld2M1iKKG6j
EdXIVo20fWrG6rcy4FqWj667dmtYITFb+ws/Q8oLgW2A6x8mnytfC+FTWbTRnuUb9z8kaqQa0WRV
cQFNYHpEPooQMz9Go5iZ1g6YSf0zJAVHeOhl4InGye9GIFqrjYDcLDMt0W0jDFMdlXbodGPsYC/K
yCo+7bA+sZv75kmTZQh2E9Xz0EYyQ56e47y3hFwHK+33v2xMFB/B/xNOAaGFbY+Vq0rrG7qxdpoe
eIRElEETe7V6cyISa+tXhzJFkg1WWTsnEnPVAVhgNCT/jfTXqnr4ht4wCap/O6FntH0eIWeaA6MA
lQ9qGyv9CdXX0v44UkYN4/UAXPiv8VYGEhzgebqOrdyWFlCsm2xOYLK23Aww1TT6YL95pnRVbNzw
lwsBUEJRywPqfuhIW59XHUZPw8Ae6zG1Z6rgcVK4MHfUuDFmLMklL1bZ4XTTZ2htI0T3iDvVWZ0/
rKU75THCStGpFt6nO4DXZOuoKwcy2nCQzRcg3L7l2Jol5Ka1Moxf0nB8El0EXczQ8vr3PUIl9Dx1
PpOZjZ3DwCWkX6b7jPokZq32O0MXKm3lIdtPET1A4G3cZYHreiufdNT7jdWXaZwh/I9kTNdK4kBm
VtnyHE9Y7GbPdP4S8Gyi99qX+f6mMaA43/qRrU34DCd8R8lPz+VljSjLW3HHPfnrsfFdLE2AzDgf
ymfVj5LYhtqDCKF+NGrLEKvxywn4kmCfh6MjEUZWgyGbJpt+x4kbanp2rN5VKM1+T9/LcBq/+sZ9
HuMkVYqG4ieSGzpuYVWpHdCyZ1r83AMvGPlnyRkw5awuiHAuCredAbvlAdOuowfEdEECeyE6brhY
ZV15quvaSov4IIjn9Fs30MIsNlYtkW2D0LAkvsCcLN2DNoVTCYtRuXitfKXZC1pJr0cA/Jj8Ux/9
YPK/xfu0+LJuTRMz2CytHMeqx1jqIK55DeVtKKcKaRqbohMbVfSHqazoiLJ/NhFZS5yXsrf7jF3o
hEKAWt3Gs033Bxwh7btdN2gRbYZtMli/lPlbb83RVe0z3vB2EKVEVP85n33/MUlrvQO896wm7dGe
S+Fej6Xghwh67hUA5NSx9nNnkN7PGvbwZuHH36nM5/Q8nc6v7wmGeqFMF4dv+vIOiouaMl66B/K4
MRJoyAH6NSxO3SVmX3jqBvEKMTvQpxY9iR8iAwWPFf0hURLKo0IZaXpQyRdbjlW306wuzs2T51Nn
d6YU+/412qgQ6c9aiVwPFkmIByfY13eb3Uc7t6TkNSFvTocX4zK4WltPbAS0iumsRUVx5iVEsOYW
NueADkhW93VOeCctbj/xnj25rn1YenMnBXVk42S2g0c5hSm49a1qcDF7pRVewQJcBnKURDw/fqJQ
Tr6T1x+x305+CzBWl6X+uzPtAvgzOXsULfqC9UqhBNez7h+i7TazJz79uoiiVS/xzZOA7hgt8iQ2
8a6i1YnHPCHq0VNmCe3EYQ4b6i6NT+vl3USRRPp/xJV6Opjb6ugFnH3aApT3fRBksapFnRyBPNH8
tXJ++xfl/LL8E7VTpGh4PCRumIPkIHCc2OpW4LEyAXF27DL8EqObXhG+GFAHUH3AEuKngd3qZKAP
rX/HPDsOzI847x141kEGFrKo/lhlLNDxtdHJzQ5dDTvQ22p3og2C7MrX4PvEG6ARp/XpQwGztqVc
P5O85H6DGFejKNykgdbr+ekJvN4glfBzBA0SJZF1bvdNr16oXTHvbWbINRHYJAuTSDwH/nP4BAhs
WRdBo3QelfpxkBss+j+pEQaQqlTwXzWq/yAvC2TsuzRKGpSyDU7geJFpd0Uq0SXry5pppKbs4Kvc
wz0FGpMwiH+znscc9ijc16KOHwppVfnqO3/yISc+JA7X4UMeufxozFEyEaGdST+oRJIcLu8kijse
EzLSx8j4KoXZVyDkfcnkPisYweZGD2Y2ZbpshfA3OsoLan9pF3vI7orpRR2OSpwjtZOk6kyozpb4
i7pVwP83vkQslCPfDuGUaMSN7kwQWMomRz6rWyTb3DY7e+eAkUG4j5JYkCix2BPHGFyUP3HUJWBX
iMWUNyYZ8atxYeqQTi45HT3Rjir1y6FDarjlZ/aAar9lC5u2yBXtLFGBszXbgvvMznJKk2w2sn3a
qRO/MWT8oBciphcbuBBFb5g75ua7hTrrgZOP6u42Z+wVXn+u3Hii5e8ftoMJ8J0EnNalBnSl8TvQ
lNDiRA/Oiaii5el5cIpIP09LSVYGdAVvU68G23yGpG8+yXCDeCKsqOvU7jfiDKydvL3hDtgOl5SA
kILkpUpvkNvXbQHHIm5f/lvCyACEHrHAH39tdwmtnCuOkn+H/Vj4hGww6q1e8HC0L2SpVnAFWpbe
mKpNnq92zDP9twv2q6sVeXgUaewO3E8E4iP1B5Pp5yXv+mWx9DEQy0vhnfuXT99efU6rU8rxBP+i
sYbta9+qd2VztuDzxVpUV0bboNlPkYC3DEOXf3159fFmutXgyIZzaMkpl7G/IjtjOC5WQyPNb2H0
Zd4a28AaTAX3ou0vtuR/PWiqaB3rlGvfyxQ0G8tUfydP0fo31+W/GYCWHmhJOqSD9bkuwscpzD0V
aNzEtM6kHRAvtJclOicOhkIaRESTG5l8f40mm/Sn3CVJhIKr523uUafhA7s8uNamcOjKS0mj+ah4
H3LiEL6kZFUnHnhzdDXTQGaA69pC8UnvUdjlKnAsg5a9Yo3Ur73VMs/Ev8zlaHZdfqZl+CF+mXTo
FRGHBk6GBzh7uDCKSKjCjGwdr9ZJYJbucFNWO2cmHrmJf6bFGdQb5cjJdaKBccf/E+0XHNFc7HWG
2KLiFV3lV16lpP5hILiDqwDFpv/NBiiW0W2KieM0qBJMl9m7eGm7WjwMwAMXWJLfyoyKi4TQyadP
xohxxhSo5t1/zUzvp8tfxk1meL8S3lPRd74Edvol9+GhUxhk0R0PfxZcMC5yCt62XdToqkg/VdeP
eSojmujZaKIfIr6EIawe04b/j3yFzmIF87RQXWkFLRTpZTKOqOfQj1hw6uLy2I/W8cEjySniry6K
VVlM4vmqXu/jb9+inHjm9rb2ISbOoeMcPM4p9w7oEB0gJeCcrY59gehpJJycYEIxu+EPvypGNwA6
kMz+XHkOMDFsUjzU7DjjPyRk+YQKaiwTsTR3S0taaH11ZCZ8Vt+F/54UZ3JHuDyDXT0VNbBzcQPg
cB2Cwtjh4uTuFqHq3rvx4kbiVao13hU0A71yb1/hwrARu3LRfoKe+w/GRtui+PcxMC+hJizVv7sF
8vmvyz/lWG5EtipfygJTh5hMMQln5ge1oMWa+8ZjK5Vi3arG8Tl0FD3ZVOhGyRDdjIM0L5vcw2T/
1MrKEKYZxR4yc3oAgpIFCrYfp/stfUhe6vf6YaoPOrHWiEmw64SPEoyXExgTvOl9/wS+zJ3hE3WQ
QDrSr8A9U2ewtS5WPH0U6tsOYKCHmr3BMzGu57sdSYdLeQPDPgllIQ/W7c8kvWqeR5yBfn1PniBt
Mt/x7/AWjhlh5WD0evQZUungDZ8HR9QGQD0lue4euH1g7nbe8rXOtQ4y73VXu8DQPv4eV08w60IQ
ubU0B4lVVAewJe3rbOxq7/bHNnf3Akggc3HvnNjovtohe4qFjjbgGuunEGVvvj8FtTnozfLobOIm
QQ5Qoct5irllmE/85rbXLKnfcOKH8Mq/kGEO05b9FrGetPxdyYXk2OmZrJSQnAf/PUTG4NCH371+
CjwlnThc7wqpe5gaS2CLmoOSRJqErX3f6Ew1WrQfNmgMDptEt5gl7kIEnKhoX67CaZ2Xhc3Mfx1T
OAPjjDd5Cn8foM59AgXKl+rcHBaEVjSKaGAby7y2xhOWzBr+Z9fnw7I/16HF2g6ZjMrFV32OUMIk
HgI5r0WAivNZI0s3CTHsdexnDgxc8X5wuDcQWqQOgHqFdP+IjNKgCZ2Z1bo/L7N5V7hdZjll6eqi
h2HrmOFlKmPj5VtjXr4wVH31pUvF0++oBJZy2DPNHaf+HgzRvrdT3cRSkvjgpivfMVhNG3SX5wDY
1nht9OyiMxKdg38zu16kaO5SAyEMWsEGHBV2vzGDShKHcwn1PDFTknxCU9JECPc4J/+UpkLlIJUO
WFBYiuJyQfBC8e9vMtDoBgOedYgHGUEpGs41R9ViP4FU/E5eYBQzig0BtW9M4fqvbR3InTuBFDnP
SJUTSTnz7Bnr5oWwmUnjeMWWzYK5TvDLbcB3/2IQRvU7gjgVBukTdpiF0rERDl/RNzggrLI3ZZj9
XcGcGZxem6EnTb5HVNuwlu3ySRx8AQifYYrFEI11gywf37MLatQ8AtbTdltKTx6r9Z/k9Q2/LNBT
FnP6JLH/kUsNBJOaWcEzhSAN53ZGrZcp+jdKOBRiUS3oX6Xp0H+9HqrxrShSQ4dmlmh4PjKxq8N0
En+pN+UK5Gn27JcfZW518HUuKTmIdPxB6ztXSPKnVEnoa+Cw9R2zfgQMpNVJY69fdY+yDCZLfH1F
VUaNq43pS9uwLNRaM226wcMOV/qWYzH8eAHyYqpCnoQQ58LVXKDxRuBoGNw6Ae2+11UeA5Lqfcm8
IcE2Y0ZCpBoY7fEdwaswsZFczw0sDpfJhPjXdfafsUl6+lXdgBG6Hf0+1LNh+aWvA1JizDfNonFe
OGGEasTfHZ6JinVSAGPB95WTkn7JxM8QHOjVqtcmYIi01nLRmAL96Ukw2o9n9HOGXPfaiX7AtWO5
qokl/YNAGYZwClK/LKJ1uo7okCDbWM2DTzUQlZEwdiwLlAwGsbURnrvvk7HzTUyqurDtofKYRcm5
Mv2laX1Pa7RUmD91O84BqrN+5DyDX1xvWFanzo93z1SDJhaNhO2I2sceVoE/dvDhbr+7bCHxpWwx
f4P499jv6U44pcKaEYcQWURgXlZZme32xaPPLS5l1hVSnHKy5YY4M+Vi78h8sDasFqscfxMWnAng
kCQ+EOXTnCwPTCkzFFqZGUWCcToEqILYpp10r3uYJFV922GDOrLm3BxZnA/jRmhSCc4SLNaFfDb6
pUA2l4NvEF/ny2IbN5WC0+OMVLxefM8e5cS5dofGwDzg3cdEAVwm5Dulgdnr0TIwcer3jVs4bU5H
5jCuwHAsycHq3+8c1H87X86PQ3qtQwBGIzHZlz/+zmiRJvSd1QLqfYg3MhjkK/qvFagyfjt4dGxb
pWz21mFwhYYhwZr2q2oO2J1IzWmKxhklYU8TTVcJmhrmcOG/APTbPUzPpLjPxRsm4HZIZGVgfMq4
t9y5kl3/P1FkB+Fb40mFQS8jicaN9nsZLSSfDPTPV2bUTeqWtuiCdvxAswEL8v6mtFotHITQYqG3
sdlrobKTnJ8zdAqe3ZgGj/6gCdvdCjVDI2OtJ6TW9OVyNNd03Vd0TpIeRHrVIn/aXulUwxRCnD2W
SNbfWDdlFh7PSlhE0jo4aHbgBH+w267d7ikbdEYZu9xWrpVHg4bB/1yQs0lZqPCxddw2n0gr2uJl
dosPaswuK/i/TcIguEyltdbPe3Q3hOJ7pipJ3UJ7rsZGMS3hQ0gLdCx7+s3m2heuGZtgKqPwzWiL
JBX4wNpmNso2vJWFx95ELA3DfeU22o/jcOgGW363MUhCVj1ZcOF1sHNWSJHOL8qw+MpHtUNbcGMK
c0+K2xeVGgMVaJPUX4RxbAxUkDVwtqSfLPQrCQJOIFWwLzjtFqpqC1DEAzz4AOM2xKPOoz48dFyL
Hs8ewaIjs/h/tXY9C9lsCor7bHZYe6gGzYNNQGyCKRO/Ak1MzBiR4z2SSyJj9yTCDWSoV8a75iD4
AkhLfczApu05R5ix54ms0o7XPPb4wajqdEFksxlDgXWD/UawAlbpnUYLXAQcLEIeOrrHLeHoPuZr
/tj82pm6fyTwfO8+VSCMYzfaHOW8KOS4Cq6+JZNSUEQObe+rFpUlsGt++QoiEF2Q6wY8BWQESeV9
cYvK84GySK3eEp34jGGkM/gH/3flm5zrmUl5QNF213AoaGR40iQz0oezJ8sHkOGUMMtwAXCQZRYj
Vf2XxiN9AbhW4IUGbHROroJ7PPDEBBsgf5W1ERdHcYNyO9A0oDAdPNs4aKfROP9x0NJcsSoDQ3lI
lrHENzx0P2YWT7z0gliMOvE4/LWs+CDfhn2F+ni1uunb/3zgM8OBdDcBdgtoJlseMpTQvwOlYvQa
Ma+ouEHq5GPIoRgO/Gb2EnLaaEq/6UKwGOvfof+Qgz4NeWktdDXn7yj8q5+2dXic5QwIJ6p89vTO
UBa53N7nJrRFm/hTf3y43qS+gvTkrsqq6nlrpCMoBG/d5pLMjV1lvhcyoHq1lzeFddEuQlbHz2bV
hLYYnaLzQimfqj/tZuTvjzDQr9BKP/06XVigP+3r146uDLsW0SUq9Yw1xXxyu++57QzNDPkz8+me
e3h03fHiKWs0N46LyPfCkAmQbTQJ2ThaIqnC6+n81Roy8dlZFngE0QpSZeGd5hEBQA9FNhflCha4
xF3ZYUiaFF005Vlb2p4f58C9aVTyFPz37vMRqM1tvDcMVnKbL5s28uf/eB9Ke0WnPXsOkCGimiu5
f245J7NV35RDfRT0i2pMawkbaxt+rq1MYqE0H6USd/DMCB2LEABZV1Z0nXt40ggfIzwG5iiB2Pqr
YTchjFU+tCDYE17X5pOmO6k4BJCl+REqY4zUSELQufUqun9NeTEf/D5doqNUv2c0lpE1tPyxWdZu
LeTf139/Z2iwEKkMEXhnWBmbQ9Ue85jn7Yrs0JU6YqNKt4qPgupKgn5KgzGuIqFTP6IftDLwUVB3
p1GbLVyla1FOtrzD0J7i1ZW4c/Tl0vfcnLFIlcSHQk2coWhsR3hcd+Y5SMJK08AHVuQQbpihYcaR
IxRhM/x+PAcw4wirA2ecSOIoGMeriA90UzyVvpT4Z/Nl4/Srt8WcbuSd4nf5v6Z0v7LD/ZrGcMJA
swPApK2xu4k740vaoFebf9luTyGAL6zWpN8OpkwW6evwKATHEhM8Zmq5CmpnEVqwH+7cjyVJ4X48
JaHt09uAMs75N/uG0Tw3jJU5VQOlu2tebkiBkSGSsBVukkubXFjmkM3GOIqsNzYDRI0EAVxfGOUb
ec/tx5oIzaeOrfdGHBoBsRMCquUm8Yigx8UZtzXJ28ulnMeexw2rmJFAIOYrqkCl+CtuVWziDD/5
ykYNWtBvC/Jj5Vaa9JHdE/YVXH1xeWvmMVONvOEBlOaWPSCOXUK7q5vYQ++2H8QMQtGN9L31kWmy
m91yLKViOvWsc9yZHY/KDIih7r16aIvIBWeGRdtP4sJBrhHyK6nPKuvgqf8UU5D8LXA9oV4A2hPF
7lenj7LkPzJt7dSFXfNSyWdwKn5cpDH0szvQJ3mWsM7iJxRJwF6IURhnJojZGeW3ukoUuj641trQ
onbwKWucMtzvals8WFbTpvcX6ze9Bdz0Nr5ZLve5S0zRI5kT8/G28m2P6dW0UUuN0cTsrQXdDwZc
7vVSlEVUb8qqIqWBmPzBaWz2iXHlDdI9VxOj+KVXnyxX0IXZdPMbQreslHeiKbaKtsPURp/KWRLm
OCRdCZAEygz7KDP9XEJueIcVT4LhxntaSQnJTDyRdbNkoBpCxsSVENvliGNOWOGMRRV9Oa24AfEl
YByA3erUEkCw+oynOkXWOeN3gmxR8v+IrxgLs/cqNf6rGBPVYmWYAhmLBDNAF6xwcOwcGWcZsu4e
lh8RRURwyc1vu1g1XEQlsLVsCcM/pjATNU/a/ePAX4nRN80LaBHx7uRmlab33GFKHTY3lqj13oJp
m1figgCkRYAra6v2o5Y1QMppFmQPq0Yjwgx4QlFPddS4qa6mklEwZJzscR+HmT8QrQMyrYCnJvLq
2oUyqhUJK8JvGeYMSzeDay18b2ewF17yIx3n9vVIlgzqfaK+OD/uI83LvFDqkWeY1QxrC78bTMdb
w7OgLUmGosyOAFhD3DBVUS0rrlOWtE0BHHJ9wknIyYL7tSQ6JRGqOPqEYQn+U8N9bSc9n/kbr17E
WpH62AwOfa9V+l8eMEffJcdTal4BBgXH+loIaNl0lFNCUAKatOhXTylCvZDqTKqtN/8Ptrz156Lh
HSqV3jtuEe5ydAmpwYoHz65ZbMu+eFLuDAgauvKAVfBs988mh/psgwV/LqzuhKsiYb6Y7X45j+/M
2ixMpaunYGnOkZVEqRPZJWYhK7ItoIiYS0RwC2lWOXqrrzHKYAICxD5c7lWfFZ1lIRtYgjJRLJEz
WKdsTl5QQ2Zfubul5efXo7YE/zt5ZaNcMDoth+yjIAonCmp76+4PprW08AD8wwyExnMd6IOiJ6pd
aWV7UCXxYHYWZvr2MdPRdVYAF/cbZSF6kPp3FZj5A2eiqpaHvG3OfNZMYfvRU1sVXsqCa11FTy/K
y99vYaxthkwMqcBPGAbTVK3Izk8gT+XeVrzPbPlPM1FhwKcofsQ3fb2/I/B2XJsJu4yaDdnXXLlN
jXUiiH9yMYHgJfFbAK3u/gweT7j1YyegitjIm0abdS7iUhAdezX/iBF6W1O5OOeOn/pH2rzeDyak
z7seLfH5DVOL1Ca1Ks8Wz25/H9S/bBRECuJc3WdHhUaMoBalJdjjcTNRiZ/e3jZVgccO4GRLFFey
gvmIDvyhZHLtuy3ZrdhvOqB/nG1lo4SP9Yqrc02JMZLXEc1HnUKalUkfj0n6umQDuA0dXKqYgEnt
Oo4ZBoXVMteLe+7aDVNYum3YCYkFJZljjjyL3WJw+WXGPVFBEDPTUjQd/pj2nlFUw2jCGNN7TeNV
tSjY7i2FmFXmjpu6Tfw16loIw55i4udjx3OW1vdGXQ5P8GqIP9o1iBnMmFMGwPNURb3rBV3eHDUs
oSfFohb9C8GwG36+f9Nc0p8tM4udwCQk50gVoXFAaD2c9FmtRt5jwsISAKe+UT3pQeHmp9a7trgs
DV2j9fp8wdRVc9ZxHalZcEgaFcao/sf2tRmGd/xDEzzmJ36JjofAAwrBhJZ8XrZj5Gk+ST5YA9ZM
hxwhyoOqgorxwZ1OnLDqElm1A0VxKqxVV/Ri2Arvb9p74J/fiktpUSFvudaYrcRFa1xicvv1r19F
69DNI56zUfzgHI+HtdUc8B2cVNDnajCsQhHHjsvVbM+f1wBPWRrVI1A1alDEjPcR1pNK5tooKUM5
L0rytP9C2YRmOrhJbDSiBxrabXikSRBfFT9knNK8zkpaYWpNxPYefVC1INujVsMekwI1epw1xAA4
z6fLaMz8NUHhAhNG8oXIewI2FrsnYbgtkcYx9aAtB/FQNHMmzPxkbKaWh1XcF8lLc4MKu0eN5fKh
XJ1qNm7iUfwZodAHoSpXlXDbjUMR2fyQiJrSHPOOhvI3y6OOhQjwefP+9Wrm62lFy5yVyIQtoUyC
hkeN5YHw150q4mB4WLkcbhn7foaziGEMZ7CaLdUvqkz8pUDZN103ebL9ZCT07MSM8R3qrzk65/3h
Y5z/MkUWNZ9cc1SQl9GBXnRN2/EnTAFVZfrvI24woWxQz9Cm0Xl1ct3sbYX138SiguNoaqkYNTag
7q5CV7D2vXzI9lVVd5rDFdUGsmQ0jTJ5x3uNqXwF7w1OxI1H76LUM6Uya+fS0+QKu7LkfsXWHwQd
G2f1fMBX9dPHCmbVifD8beGtsbzwA27BLhbsuWJts2S0b1lv7V8Yck1C7oxGr8n0rYeuTTECTwn3
SeIhx6czO7085wrReJtVnxoAA4mp5jBy0ioyW1ndsHeoTm/HT7F9gGrQll4iJgkzEh84L1NK5eb6
lMYvCkBHPxfUJc3V7iLEGQ127OTOjdXiVeI2gDYv+Rx+Y6EQd3DKRgxrklj8eFAiGxrXsdSZTFKb
65kbSkU0c+8gB7AKIT8InhA3ZXbBidbj7yYJuagutwY/QYFxLdlTKd7DIRbSM/WvYQmJ2kFEfWk1
L4tHzSV4j0ZcPAH0qGF5e+Xv2KYWx6VdpbhS0pYwdYpU3B5ls9Cq7QAGbKCTRavf/Ock167MQePs
Fvv538srrDA6oY7CtYc7yBbrmAtzRIFpCXakOdzw1wA6flQb0m5sTj+rNu6NCIMup+MhRxlhiBIa
MNSzzmbgYRLK8Az2Z6kF98goHKRNuEM2ZSPxqLXiPZGGVE/Om1xi48yd/ofdBMXo8BPUs49GpQmP
5rvPTzB4PpqHBqO73WpANPlgn4CJ1GW9w4W/pUWot4WSuu3de6E9JWYYVnDtALyzFjGrzud1liM7
KViCT4mvRKVXg4yx3FHe2WeWBblkk/OE9FFENr9Nbp0yZO1J6JCWgjJ7EvtllYmfcmsWaFstw/Zk
rv35nD1C3bmTwBKKHP/ovUQWscgxlvTf6w6lJF21GAQWBDZVIHOlY3x6SRkpiEpobB0JVQFB2K65
IbdMqeNEVxjlErlCj/cd0AQtwyWByhqZsVJ8LQ+TlGk8C0S5d93YoVacZnZ1T9nI5D0W3DYD1mHE
neERFktjF5IScli5zhm6Guu9hhjYgdaR2mDxFlp0UWjXmVCFjBVnOeNwAjTt4HnnoFfdNTIfRqgf
D/wmipoBrhl9zwazxck+MIgiZBRshQOAJMoct9SNcWr9jVR8XRdolAaEZaWNLdS2I/p6FZusKcPY
WDyQZkTyfcjHpHnHDo07HEvJaHorSDwJYecFytRqIvxx+ykB+ufeBDdynz8lN0zT/jP2W5P999UB
8yn1x6v7S9pd/5Ntz6j5vu/PglD3D8joQZox6IykT445bvw+g5gz1XGCXnNSQotoyunyD98mtL9J
VvDpznf0XQ2lUcAswQ/1XyYY9YmSOM+upPiJYQdOkbB1Ql7vJFr+/fboa7I7ENZkSs3+R+D7NPQV
DTHWQB9xzkW3Z90WIplr+gKPdpSMuPe0xIaHx2hRHwJoIX9+Pr7GJ2OuYfY87sxvRRs/yAXoz8hb
3pnP/XYvYJi4QmtLKYpwlYgGbMf0kHnKR8ePbln/q7eCKshvdj/iXaJ6zc6vRMg4o9N43X2WIu/J
szmSj6OD/uqj9BOCIumpqEv6Pi4EAzo+eb7vDBbkjhfsZAembJmaGsVOicjWq+xK9/rPCJeMH5oU
RQ7Xr5ppeLIeq/IV7CWmMtR6UXycxeKtSOim/9Pp0OcNK73SFhokNoP1E45uqo1XqURrbEnVQS4W
hWU6WOzUtf6rCY4mPbql8psx1/hneIau8mVRMweNnDzbb3kyI//phKWErMHaZB8N//X4Q7UzGDq3
4PedlbK/10puRpDJjL1sJhZGGcBJp8pSHfWb1HVRGrpGGu7oE64sDUHcx8cpFjqm73VXCwzY1wWy
vLvM3MkvtO5NcR43sm/2K7CEf2UNB9w6xrJNhiNdhD1RFJo0da4ls6JtkKaN41g39711opY73wZa
WYRYo+8lyQWfiEhC2lxeH9l4CMNcc30VyF0oDuvXV4TTRpA0mB9KmAEY5AK9bWZgfpl60MAQw7s8
f0TRNNYPDCu+FOVs2VCBf9P68RZfXh0BR6EFMbkD0uXPb/qgOqhnd96tF0RSQJKf8geAiCsz3xqT
D7tHhaohFWw9SthMJPFhCv+3yRt3WE2ft1ooN68nwYGmvMNO8OE1UOncLmnvb6semZUncclakSGj
eaePL9hTkWzuh8VUykiGqKeOg2POVEIJCxPg9RsoF+IbXf07B0o8LhIaMH0md4yp4Ldj4y/d3FdI
zeCxTXYeUzVsSxetqGRHO7S4VRTC65PwzIT91kJmlQqAl70Wcre6ZwFhunEGrFKPEDHhvfIUULZ8
gs22/ZLKiCTn1vJntc4Eb3o4ztkr9h4hB6JLL2QdW2g3KJGMpmCcc2rvEBaRD7P7OBVYMBHoNcZ6
YwFMi+22nUGONBb8bs1qyMShsln0Dtn+vc1KcLw9CHU/VqdQQ5LuLUM76vHbZt2bIX3gj223jicm
CGujJeoEAo89UhjBh++WJwra4xaNQ/btV8z0Lv9O5Zhj9QbVJo/Y0UTq+MtB1+uIibNpgo9dU8A2
jfyCpMhN4OIJpqrIslUoaYArW4TO1DaJYdxRjZhqLZFVhriRSnn9+9eCEytryBEs6urXsh0cVSmR
ecl9xZm/vt5+zKVydI1MjHP5x44574WhCWRQ7hivTtEgaJucxhZgxtfmgypqz4EAsNvbYvXkgtpr
W882yFf/5C+6x62ORGU/KMlMe59mGUBCP/k/bSdFhCEOXIeetbliEMssQj4XjO0qFR2gA85o/ouJ
1KmoYjF46fKQOlgYksat58O3Z+DPDwlMkXg/uupdJhNYwtpMShrl1NNittqc+EQVsbIYKrVSSMI9
pLCiqkTPuzKSWC+8EAGIGhqQFXMPvwB5zypNiGWLS/w6j2P6GVmgHCHSmwuOO4JMLcrt4tp/WvPn
ruUxFWjxZ8zgbHXkXBuvF/du2Tt4ONtV6YIbmlsCUAZSdFGMph45eM9og213TLOzBjpPmMli2F+p
BcZiNT6Pz6jTcepsgrPBQmGI5MSbLU35P79y7nt2E6++sItfvjnOs2mk+5eOg0BFPKN1cHet2h3m
pi/LoXEc+2gbw/BtWnL8oBqEN4qGMSaK7pqoC4hqLPleVSN7iN5lOGmXsOKJzgR/RtBzApZkazO0
VC7DMd4ADld25CasFG3gNfu7aPtwSnu9qi5Su4soLZubatFphpFyRmMDpcEtRpwqZ/TGSx4jhfIR
iYfxmVBSoxrdop69gtFMGtpot4ZKsOmYbI0PGMRhNZoUEWWKQRNfxCmWUQdM62x4TnbBd6qbQoHM
BXswFE97NkAYuzIYrAuHreyx/+OVuAX9DCgyjsYpw/IPKKz6zDvjeGF/0R4/fXruV8dsomlMmg7s
15b6m4fb6KD3KqB7WXYp9uxSugwwvu19ptWWUO2WtIdkewVY+wWQARiiX0sreA45HZu/6KP5Kk8x
II9tt/6bZBI+UR2TrJd7rY1lle6O01ZtSsddrlmZcCEKZaSd8gJgkx8GFHf24TopG1wkXgkCZTjS
nqdkI32qBfMwGgynn5IEKs7O7Wb+i/q9m/NNndmr2kz4GJHQqoQ+zQRCCbUWyP78i1OP20hotVGA
fSvgpOyL6yqynqve3qYiRBM5HAM75DjzTW+SK3mHZ+PWoqXL20IfINenXaGDX6ZYdtFoHkYKZ54P
mvGCVYG9vOHmgiuO+xTvCcPmY9wBNiFlqxuEqAnEzhqbS2t2QA8XliFPBdkW0NNNaINVh2ufoSxb
Rf1b7fDWspXloshpIfuTtHSYxbi2M9BSascKbcm1usqMNiSfTxI4WDhKwPtBqIZgGoj0Qsv8nABs
aMDqiErHVcWtuCtajIyX/L8nwgJaYzsyin7jhwkkpwmX1YzI1J428T29+6STHhjfayF0VoLdBBCS
JcUF4p7vM1b12QfPlHIH/MgZKLGRN22iDm+AYHs0zjFZhvLqJjURqI91tLHQlKbiWG5TntwmKEMZ
Lii7I+pXIlW9ZZPbfcY/D/Ezn/ZOPMHas031YP0Bqw6WKgVCAcjADNaEm0UR8dpS85D2B6QhrQum
Jf3IWUhY3f/gTTt4/wBtchYRKunxIn99AUrYkhEVSIP0n3Nos3d4m2CbEtMycDny33Nodeozkncd
tLaMgYSrdQ1YFh7D5OaMciUA47OrfDl3ZrYDn9xOtEYfLttKQ/5hdsraq1mqWhVCMON8qjyPysLi
q8zziA+dWLLQXsqyV7EVjFJ22ZZvS53Qmg4dLeicNf5e/DlIvYo6OU9UL0Q12KdSiAZVtwtP3iFi
p5yPcOXBGShr/ETGq6YEIzfAc3rj8gSoMxlcJ6f4OW5hUJsnCExeHdIbR27nmo+RXd2vASKipbLR
yiNkMoBFqmohxLjH74pf41ilc12LfgxuKixbUiZUxsFYu7ohmmb79/CbIeEuY4byObpZluuyT3Ty
pOycJ1PbVa5lS4JX3bnUtjKGAmw1HNkyllDsiABxdwqJkmg+mVxjGjWy/SthKFt56QivH2PeB4ep
iVlnO1yqjYp7JG5Rfx0Cy50PjCWFdo8fKrwzFSL15wOXUC0qBco/4Pzxh9aDj1fBZDjh8grxbvpa
STAL8ONpr5CMuUUbNVAZWnsF6tRsXKOJCn+rwCVqqVZa+5QRC0tNtGwQ7TNNMlpRW4nOLUOtG3hM
KphLeJT6ysin2wBF7yFzWGKoQWMhMs4+9nSwAdJ/uLVPi4m6TE7ihSjeZvBCEceEV/CUdg0UqQli
iD2wZRdCKZPIVqxCrK0K6DLtj/H6OGMCO66fHa1CpX9BIAc1+xBkDG4+mMgm/DE61Sog9Ym9z0g8
Tkx2GloC85pfjqztCS8ADYxMxbzdP96lshrc71H9vsF0jSRvammGC0LfJLqH4FzEBN+rUUqK08zY
Y3XiiJLMOf3zS/sM1B41UsgyfkeAeGQCu/Pynvyf44ouL6t0270vfbQkhKkX1PzpEs+L0Lew3QS4
wTGxo98XmPBUF3iVbdsTCUWxp4JVoqYRlD4SEAITdQGaQDx1ymKBA5hDOCTBSRIJcbZtNclStXwN
rfCIRs3rLJBv4146c9l0Byyxu7eLa4wzDElMprblBh7OnJNVoc9CdqHU8prEU0uAhMiT5JVD9TBC
SQ4iI3MAoRVO4K5lxZvxHQiFRmDDJEsLPcJ6T4tsl7P8XJGnZfAL73OTYdqHnmO4AiQ7XWaxtSto
shxXZ+9UN0UAmEhpjKfl6iBkTAcm0brJVuob9DB4tdZLeR+F8Ct+QrkhMrRA2+W7CVD6kkeatAXc
/lQuVTmIScgdO8Qh2mIAWXAxtbkNOUODO6EPkKEB9rckWl2hAuU5wEVHMnKSdD9ZIw62zrmgBp3a
4zp8NMLtRY5qnmrf9ktkYnJiChYXbOD4CA2/es1Nceyi9NUeV4ZVGykcXNneY9WVBwRgBDS1yV7w
XXQe+MuBTB+mV16R7L3wmnk9YxLLQk48XtrEDA2/XxruM8V+RhQTlmjJeRzA/UqBQ98sXS5OG94M
DsG/H8ZgAyLzrg9efODfvaGGI27qlqrPgRFd0wP9/Fda7R38BcWEk+++et181XTYeNy8C6OFe5Pj
TAgA0Lmg5h8krjIjQVKquJgWoeOgE3gcLIFlw9+CSMX8w0m7MNppW6wdtyOVeTHKSplu6m9OLJ0/
i/Czkqeh7JCdCgW+k5boeMUuEIltBaLoPPS1MSyPSMHBfiO/K9Z4p6we2x5AbKRKLDSUzqGB+WKK
uXY5+R7SaNnpiQSixN0xtvLExi04ULePo5q4nbKMqro1Wg7k0bhUZx4xcJI7FFP5iP3yHCp4twgL
gmexPeoy61D6Mbw2/hV+VsRf1dlsjNTEyxyWmwHyMOu6qE4cjpSY7G0j6I3XMbP41qkPV5Ad4qtQ
4IVfTcQx4Zv0jucYGovnrtMD2btFJxa2AZL3Xx8nslKXG0+OkRSx29tDQWRne2XgtAXS3ojmba6R
LZs+NSiAhQ0/ZUCcQb9fyWx6UPJ0KAkiB6ODFjhrPtfibo1zERbhY6oVHqbKX7VZ9WAo4oVcb4JE
wp1IYhfSaiQymCnvdkMneaGPvLNQQROyWQkPx9ge1U8aufWuGdSWgkJq+X/nym7P+rFcSGvbnuMj
+Y7Or1PwjwYWqTQXwYlpZLbLjIUl/+Qyxr+2F00aTK2XdPYIvXMhLvoB4fsgtNtjSCjGykZAULsm
qwPg5cuXsg0OkZUxSk8iDiRoWFuiFvvANleW/RopBKgpNQGN+3qd47+saxtSGafqtqZGeBtsafqD
Ges0P9i7Jewfehl/nRSVoU85aYPTpxMG18zcewIPP70h5SbMFKpuFDCOVJY9Plypsnw151CDCmcL
egZYelW/IEw9QSff9k1/3q14abhyHjtmK/m2kN1POPWCqYwjyXy3xHhfuYAqXZL4sbS0SGdEUb8u
uQQQfR8MLD/sSw/ROwEZoa7jm5qdsmw8Of/5iZot5LIIUJMnwPs9qL/+7ZklSQoYUtJMUcK65IZ2
B3UJQ7/FUOv9XX4xuW3eBdXDPdHP4feC3CS7OjVQ/aEO4a+FaYkt5Zyj7QPzHu68cAvjTe4pORE9
xZHHDaSU5nG2oUwczolUR8mBXXhRDhLZqVIqmUoyQ8t+TFnP95ghT3hnaEpXV0OrQO9hQ5ZVx5Mb
/9/hM/0d12RlxfTCtaWZ13y02FVJr3Quqtqm+YHtZ9e+Uw+gvjFE7G8jnTIv08dqbAN4lwKEenNN
EJ3Z+Tuv+Al7IBf1n+5FbqvKJ5ikmGimIvAfrhxkl3V4ZW4cvwOe5ehuhpKzEl397Ty8tYVj3SQF
fXp6u+DpopPBQB+gaogl822eS0vcdH19ZUFQuZ/NNmSJsaL1RrSKlWs45YkzEFZfw7bEL+IsJZ0V
IJ2KiGVb9CgUVRbmiXoenaHoQ759qFyr6XJE6i7nIMkXjwQKtizYrKLXQx9ATwc2+Zsx8qYJvQGm
MrwoQT6CrepR8GoBhHE7d5Pomq/e6B2JWXStXm8Ppg9maW4o9QMEDcAV8sDp/iUMP+ClfQ1GK/YV
rIliQWpxxUPAG5Ky8TcPppuVijqfdRXINdlFIHPE9puXSdJnISRjnh6suxzaSRLkakj0U9w5fO6R
UVo24LpckLuJWfmYHLVnYD4clC8NFxQKUrnJHVQ/H1wl3KI7MTv/+Dm9pG29NSTubwn7Pkn/1c5H
IudFC17q35xb6OhXUB2mbAjIceEWTmvpPjAzm1DTwbCbtHWGaHrGVvu8Gemc71JGKhk68HlFqgXX
9V0F2117mJTfyz1+aFkYcWZ4ukc8DQCYBi9Veawpfzf9/tabVQMmycPZDovQIkQpWD0BkS3XhzDp
zod6VrLg/O+sIUuB9+MW96f6OKjIqg880PENdLSvh0SqmhRo/trxHaeH3DbDIZUCb35c1JUL/SQI
NNj8bWHJtEh9d1cFyAWOPENH0Eq+nJpZfc8A2uYVk9yyoZ4YIWZEnQuJCPwxQwOh7rbQsNMMk6yc
dIp4btDMWygCihQQ9a5F7F76HULu1pRnBb381BIdZwpB77SuwIpNmPR17XcSGqHnYUo6VuRKE1O6
/Hwe4uQbTOtxOD8kzpxA9EJuDeUyjsafU91pFBCUELGyFeK9sOeAPbqu3IJ2VP++w59V7S8douHd
iM8Pf7RpQhTxTyTmVieyHht4HP7CAeZS67I4SunbxrXZDrNPvrp8yetxFaQANCQQr4nzlKu/eOpJ
FH5Unajx4OEOnhRFcON+omivIQ50hImXfWhDOzNnazWkiETeSg+Tf2ya6i0qk6DXVyXo6vwcyIHb
jDPum5+Af+BU9e/9WqELMmxyBrEHxkZ6D5AM1cQ2NWYdu1o/Bc1i57YXtmo6MYJTg4fnTNz23qbY
EZhLT9VQLwk8PrJbclioeIrv+UehNyiwz7xHrDuITiPcFcKvudIANtwPgfoT0utkixjhODd8rWWB
F7CWF+V0cJzMxs4aY30e+Ty1lIFztFs3kaa+b0mzaIHnmXC+xMlKwXbm9o4H5QL6ZdyyQ/529YDh
OnB8aohrCiRQZiso1J5PSva+UrUq6bobLxh3ia/SuaYnD81sl+bBM47nZxPxwyLKgq/6CKUzWW8g
x/SWyENaPaeoPMZy9WJtdb0mNOgMPFVs8ZIfIcokMccpYAS5GSA4mqK9G6UMlhBfFzpraqD30XFT
YmQv/4DboDAzax34hmiizdqZ9w8rWoGI8njeyeN8iSfw5RPhKkrHw+HszQQ6dSLYccRZ+VX3gH2G
azRBMcksd25mxek5t3jGCpzmScHMDIZLaoMQbN4Xic6gj4jNzBOONjkpG+KnEBMxjRyRRMHHCt+v
OZipFcKkyfcGUWXLDBiUThXcN6TLmI/3gTI/wDq9D+oSYcQ+jhs9VRTObi85ZyLZd23GZiomHncO
WDOE7lCPxwuUb9ETFo6wYLLSrVpsSXjQZskSbgH2dHTC19cgRy5C/qSywSbVuFSepfDQUUFamAFz
PlHED0CsX2cIB07khjh5vbEje88TcaKm/qz2V+NcR3iKo4RBoOzCmXZG2cZPsCAqHYN+4I8wIBwU
+1iYE0QdTumiPf6ZE+gmPX9oIBPayctIxcfsBsFuZjxzGuxTS3SgZdlrIBUVGk4H7awbVgT8eU9e
UWocbG41lcnjJKJnMM3/Gww0F1VYZkzHlYZ+QdKLFbQJ+z3owEw9yjP+dxoL6/4x5EDrMi8XGQ1i
35yWZST8XJvsHqBVBB5RFl7LAenpnXY/9KvIy92KX89SHjqBiwZLQTsIRUBMD6Nga628VPxzEDst
FHo8Zgi7zbCEFaFmJcMfN3uNx5A9cO1aVUMGHeJx2oGqsBXcGNgHRjsBRuYkZ2wEYrYmN7BfYnWy
3kvNOxPwMkcMl9T/pZI17GQETCo30SwUbpfHdxb7urJW1dfwsCuoZ1leL5dC3/6mfEo677U2VoWZ
2DCvUFS8y13WsyOGmiKcx//h0dyMSK2Hvr6u3c0cb69Mr55dVbfUFp3JF5BN9/7/wB0FVOnUX74x
uQhHzW898NZCM21XpViNBFZM1rlO786y6IgkmpQcx07df5N2afFZ9TvjW1gUSN3V00DtFD/dWqHc
Jda96p+T0eBjWHjwe0X0F7Bc2TYLr87Ja1V7TcKSyUVnOQNws8EsPlIDYGQmbnXa7W8K38o43Rg9
UzT5HTWRIAPJJBKirl6VqnUGalr0pnf7NU3gVL8hqcca8nux+ypb79Tom0QMcbaEfqu0UkOpb5i+
dXzxoUdUmz16BXNFgPwmdk/x6E0Ve3eNeCrMQEQqG5YLHY6YOJtsgZNyqsrmtfKLKHnC9lUkSu8j
g7X3ADM+vrtpNpdhDf/X9s5YYeynW1p/0PBhe49SVIIAtlbn48O/b8qyXhCnU3JD8s1WXU9y8E3t
eH/hg4hrze4kJsS/PqGJWBmk2IVwljNOCzQ5InCjlowp1ux9rYjVKsclpe3+uEkc22EE+151z96F
bUjGJNKDiKXgGkRz/CLZJi5bwhUi96yuB/2NVPLGF8KIDyxclHKt8nElE6cEl7dzMH/NPWbBT+cs
927gEl3/wR+pct0JEUgoH8GuMowBSm61LkqhUNv8/x3MCwrGG6W9HQRlSzKacnnsmYL1A4e0ARWW
F75YNnB7k4DQ2fPihwFOGbsOxpqtXVCrp5tMzW8sevdpdPwGQ1NF83y89TUIlEiMNCshVVajFD+i
H/TztG9PYhILtBgV96jiTyav1CH27qSZI/Uv7iGZuFwj97z2KkjvKwH+Qtak6Wpg9nueNOS+Ei3N
5irnX0kqMUG1qG9Dk5+Igi/8p/3bwukUTN1hx9LIAz+U6XLVKERvq1MeUzPN2B4G+N0VnZ7+oiTf
9Igi9Wjvr04rEV9jJ7PcpvV7sp2YyD92qLWA0bo7sMMAmDIMVrBuyZEMfH+Se/HlvI3nnMONlVZH
GzPcwL/Q4wBSeJ7sVPxF+LE+bbOIDmDeu7Gqn74nu4D/pSz1oQfPUzHcuypXu+pFD7w+GLBo/7Sn
a2fvYx241CysUjxOJR2n7Krz4d0zY54qyiwk6KehoV6E1RxSV4BQAvmENHWsGXtEJpfQreCMmdzm
MrJrJds1lDlckvYcm6F+dmeyOpYmmQ7J8W8wlMqS0ny1COB/r7b+jAuOZKOfU6N1kcoTb62hbS0q
Y78OQSF5WHzxoPISys0D//xcKLzCdVDzfJdTyv1SXWUFUx1wT/lcIijCRIfadXZesQ3oWThqRKqY
SRSyfTwLZOT3Np2xv2q43jT0NzyeNtE8nDCgZKZ2QMOKwFEV2OAe2JLxWdDDfiWQ9zHRR+ULhyM2
KgOfSK+JRo4s4af6xbq48ZSAr1QzNNivni4l0biTZJtcwR+dG8OYu6SK5p7Xrkfg8OQe+PTYTV4R
L8GII7vtl7RbaBdz8c6zeR7qpZs1y3N2ECsLzaZnMjqPY6zXtRipIyPTwM0Ww6xYz2zkkgEBz5pd
oxgvSlBamgutiDWJ/Pr6Tq+FO/e6SZ4ZOmxstxn+a7DGfo/0Z1L9FUPULt8JEEypsY9mOWJBYWa5
xI8BlE80HJjTI0/iNyAGBhizvNXNsxabLIW5qBbpie3oEBaLHIfSGk9o1Du6yK/Wf1ESZTvHn8lp
/gFTsZREapoopnPAYtoM5IapQ31fg8sUqxUvupbMgh6xK+9iRkwUhPJnmSoRp5PR2er9URcJ953L
L8ateKIwFAUBsxYk/dqRDyUMK1iTIqWZQpaCVlOl6+0A8oeZHjl+3VW27oc6UVTr4lFpZZ9UnmWU
Ek36s2vHPZVJ6Q18LOwjEjA5xXjhpJpbar+7GhyJa9H+DEeBJbvucY4tuUyvhJ097gLFVunJCKcJ
K1aTJy/0EPyvd480tuLTXMGFhwM24Lml253gLks22UEkbMVGmKYYHgbXO1beHqLy71F/mWChCKiC
rjOFY83d+eUsOKq/vv8k2O7zysk8oDSjKZX2IHjdUoYnEEmZvoLiSjslee2wiw0bcI0gKmC5LhDJ
vJwNdindHmOUww31FFoM9cPs7Tp/3/AiDCPWcaJ058TOCeuUQ6pAffA2QD9gaIR/wyFM7qdUsyty
aRR0vUcbp2Y4Aql0FfueIpEPUMiwu61kOX2iuAta9EjyDtYTMjoFBBsQ4CJNlVO8jFjuk8dLKeEh
T7Aok96ojnLkzN4t4eXyw+52qGwQPRZs+C2IRh7f6ltd+oMg6YzoryeOsUW+03QLiIEEb6+/FUtP
tztGnA31ahPuouoorZUWOJZWz4PwSTX0uN9ckf/gkGFqWNruj9NxhkOy7veeoZEdgapNwFkFCTc5
qCvtJBUZSM/pleq9+7lYq+rhvx5l2mdq86wUzXWwB0ATT/xswyP/28O3ng+TgakqnzTexfmZAuo7
y+rRHw+E0REx0M+YLGNeQI8w368HluZlWP/7w3qeB9RrXaZzYtmzCXNI7e1mAxJ4InWGQHg0DjJd
yro03GUadfDQJ6aKZUbJEw8htj8VHp5XwJd7bUbfZYx+8cBrSbrJ49L6nmDf6huoWj+9Cj4NplnT
uktxvL1BL9XOJfVkFTCPNoBK+0eHY5eSAu/KN/U8TF6YWbGkoGcqq19DcJVO5Z/b/kVYwgBBbOE1
LXcHvtvHHY6b8kb1RUA2Dj/Ap7jd5a80P4lsR23HrvNX3NypbKCRj8cHpHZ1LxrxZYyGTUw80H36
TvwtTR7IGl3LsfMxwRmuBJ6IBU9x++m53um3fuFWgvZ+tZh9HcvTAzV0n6LCoMenyDmsxbjMDJY7
vuzXvtuex6ZPI0HwbZVMEXmYIs2DfhaN53aYvYgEAUcxQqbwI4+e6hIJgnXURL0SJ293ruxPQO+b
zXrnnHjQ9UF8E0yecVdRMBQ47N+dLnLeI8XO57GX66g1XEZEXsTVgWerYAC0gTPgVdWj1zpgVzhA
aWfIx+1eoQPq4PD+uy6olW/yJRkKLPGEYw4tTIMA+Hb8pi+z8GM1By7/5yFkSAxu2wTzA/ktjXU2
UMco5aY8+S8gaP9YqwEbKANUkKGR7bewvnEdqHo7Nm4MiuroC+JtI/jcRxgHQRslkUw/cuFaOQGf
SaoYZPoq1QuXVeqyvWlwEI1vadYWLlzEldp3zb0L2BStq018z9d7muUQe7gzO8ygw/dZ0Bc1W0jM
IBlzo4kTQD1SzS8QNNgqeww0iZafNfaQTyXUGU/ToOs91zo7YRJ+mdddQ+LDqoimGay3iYOLRUpV
ZqTQk24MsTpTMdTYQjSYgCui8JqzhaNElv7Abq4KdukzzsUqYT2iOIWEoA74Tqk/IXv5Y8ZdIC36
IJOtAAzrhe4DysQQwX5kWrPUmhFtsgz55I4UFks+/eAIAco7y42j2FT1jIPfMxhhdn7kwFqAAS+o
E/MYoWbbb+QcQTua9zgW4EfVA1hVjgs7h+5/8j5zz5hfaFuqSAu11t0Gbn/996Hw5cPm6FB6/+V0
1flgwA/qAeFIF/G8bFCn4uddF+YbEqUZTwmv5Usn7hN6Sn0W+UafN9AT0afPmP++St93FJz2CTmv
nvYCQsjd5PNd9p9qa5/MzwS57jI7wROoBEfo6vuAdpfbxgV7jt4FZG0rkbBUkX04cS+nBN6carMN
jxmGfldD/v9ZEWEpbD+5DcGCZb/8K/lK8pSgim8t1a4tBFaNjBtuwo3QAM6B8536yQF3rhBZXwhu
acGrGXRoJMWqaJhdoZYfg8kYz7k8aNBPJv6cmEmqGfSxUYpqun19kud4uk33z3Lz4pRQlv8XE9mG
y/vOxUeSWr4iDvE8svINnqqnTznjdhjncZxbLoG2olnaNrMAe18H7h6rcGGrqDdKdcCVDQMaa6UY
aQCVeMMY1TMumRUGAXT4/3y8BADDWnunEOB9dhZqOFYStnlQdhQExf+ZeZ4C4toDxig+lqk79eGB
n88vo2afdV4vZlSe7E1ZoQS1ztIkWJLgjulikx/AqjvmG1ckE82sZXaeRc8cKXn6t6I/i32HNuiC
n8yK8CSo8mSyX72r9evBdBblGQm5r38Et9cdgShaAc82flep9Go0qND2s7c3esUY/9SayyOeNNv+
cGykLwBhWTlpXKn7fM6SEo/kVDFwBtrXKHv4OinZg02cD0XqWP58Gt5QFdtmNJj+DiDjVTELGidE
oQ7kbhbb7MjJlt4dy4Q9BE1KpjlOnlwBz/bMb3p/wtei3kMbIrYw5nQgqx/yuwvFZDPVwXYtZrKo
ULcryQY4BGdwG9VMQ3tcVum5q8knsVNis5EkvIXA6XxStkAxXsj1q7sJEEvMOrDuH/e8ftATFOJr
45XX176kYRSAhsToIu4nh9pi3Yw7aboiCgRSQ+rfuXwkINhwQrCRj2aXoYPfG4GDyGIXP1Lcet7k
SSWWdOZA/Eo4S+O78sPQmb9IJ/ygD4eXfx0qv+Oql76wCd/6m/A7kMkM2G/nSzszeFC+p4N7j2fn
1aOD1MdgXsXD9pTlZVEiXHF2UCiLUOH+a46gsI+qT7LVI8NH7UAOV9sleUvy7LK6WBHgYQIwBeNi
xazD32O73xejWtIRkZfguWUIBksqAii3tqIyoK/ERaGAibMwKr4FHdbWOCQpV6xTn1NynMBdmrnF
nFwHuEmjemXGpkor/md3UAGL0XPK/H4obRvjtu47zKm3LGBlAgITfc5uVIN8FGc4p7Aj+Vpo5a6v
qCLXNrjK4F1U3UH+y/gjRvAx9DdmHpvDDcxasegVNGZBguNuNm6XUN8TF9+NWNUTXJdJBLZyop57
8r7cK+FelDESAmhKak2HQcPhPCTscA72+/Wgy9DNEaY+a9EjhJNkhIc9aOcOvdlvjg1gD7D7ihtR
ObxSWGijl+sYIFqSIuaBMHzWZ9WlfREQA4MQAzWJKUo6YX+d+gkwrfpfuW8P0+ilaJx/MoAGGhcr
Rn7sCZX4Ms0/X/M4Gfa3Rt8+gRapl8VPcvVfHrWRSZpmph8Ei6CZnybsv4H3g9OiSIx1/3N7AT5z
GdujgUKVsb5HxK3yqRcitZzhGKmmVoD43ve/0nQEg2aJs7zOOcUxo/qZb9UQhjuasuFxSKlYq+IU
c3xQzlx7m7t6rHiID7igcFDCx4ERTPZGGJbMOpA+Xg7uau41nUU8KCdWmLXBgVUoE1jdSKUOMkjh
lsjcuXoPcuf8f/H77vJYvBbwzXnIXr4w7LhdsiyjfkUqs6XjivPE1TK0tenPY66ZlejO+b8aBncF
nYVFvH7FrM9xthBuNIJewUTFWH/A62lWln9BL6sAc3ihdkcbzVjFb8nNMYFgTJxa2GDa1r6N7y4N
Px1hKVJJWqFbfE78lmEz7a9z+6sH0m0TUS/htXmE/+3stP96zclHCo7DOUvlqZikjtfwfIuuH/gm
5xnSpKTHfcs+NvAbDbIlNMO/GWyJYcvE4p6VFzoU0Xfi3U+MtTMTMyQQdYEScuy5du3nHtQDfClO
jJnj4M5YaVqOWDdcOwmKgo9k5O9/219JEKUfS9kGz+S3JNET3Aidq2QYdTWeDkn/ShTauGHH/JwA
unIsBpCGr2SNBOxodCh/btESSVVQXCy9KaiT4GHpBg7Ai1YNzQnbMW9y7B093+bjHL88FBibLAhy
Zt6CjauiBUXemVgtyZHfEwxYKOMz0FFErbtl6dM1SLtYFBcNuL4zGTHKyqMMTOpxp509gPaXuMWO
3jNrgQQ4v8qhQ2yhjj+V/KD5/8ksGuBgBqB5NVFTKZU2JPIRLcK3hfrQy/g2V88BXf0MKRTZ/iRQ
EL7N0tlDftFt1+O5ZZKmrc1eKdkWI5sgWsiOtsFgy4t5PcqekFxkRzoztfR+/DBBGl88x3tAFV6G
n9omQsUh/MBG9FVryV1jEzFgB06toQPlPLmhJxNHei4V77MDs4lCbFkUBk6ArnY2oFX3RGsdJ7r4
m7TWqR/lfI3Fn2LyQ2AAOQ437hKEw/gO7bZHuFaAB+8E6ga/dGpl3RaS1JR6a8vllbLBb4R6gvGp
VkIrkLuI+d90pwfcVMpqWrotEEeOvkMxMauUEeBU6+Hmj/UnwGQRhOtFxfNNDav5DGXIcOwzoo4d
G8MbKuNYA90es8fNDtVziwJot4hkyNddFHQjWf2B324PmiKUwgMXAj25bAZ7xssttZCttxlW+75l
YEFtOanENh/qQZ6MmFaVMPOez1xx2xo+OwE2uMlfBQXEPn2r15dmtC3Ygw/AWwxBAA7kucSr4hco
kHhLPit67LOxIjTBFVow6oG+xg04Ks9zzOnyPiHGVLczRWiNW1KJ2CeblMYt48l9qx0rJSTnZ+1R
tzBYSbzCJESJgi9zvDY/kULCVAGJb0LJT7mbnF0DwIN2ARTkVYbhd+BAq8/b3terVgBC3v1SyUgF
gc41EewEE4Tl3hI0mDebjeqRd1KK7WbHk1M2J0f/JnATUI1iTt8COoAzq965VW9PnubBeMGLqFNF
eEyoyZH5QPlcdwUIMjOe+QwSesmCVZBcZDdfbLOEMRAlLr30Us6DsS0RGqZr91asAEtyuc12IEGP
CYggG6L7r5u9HIbQUR70Xv8itshr8yNtFQMT+bRtyzVY0jIl7TwNd/bSTyqWqp3sf/E9HXW4dCl9
nyia/uNtVCbFQ+imh0ah1YGliaP/uTzAfNNjZ84xjotJsolQNncBxCTeEXfrzs7cxdaJVKaDjdT4
F0CyH0sgNoGcoazm/CCwLQB88zrGzDAgAH78pMITN6nIaqrsMJCCtIRRN0wo99VxQSbYkxSUsY5/
XHknn2vd9ewAjC7peG4nnCYCijgqwGm1xkHCcArOZJ2jkgyuSaYDV4EnuB5LmRnqMn6BFpVGZRM0
Myut7zAysl8VcDUyyeDfbzZS2Xc0uYvIbiMfArJh6UrwoeHI8LsU4FIclnyz6gM/5Xh03aPpe+bX
N7WF4bWk0nDbkHOoSkdzyV33apNMdT+L+sIN4BFZEmAnc/CXMXl7uvRr4h7zp6Xqa37rDhMx0TLG
rxz745TPzVbnt+z1ck9XF1qMa/T+unN6acClw4SXTgjGjXlvgjgBo1+gx+fKFfkgNfRHZy5OQraW
4d3TbhIEgcaXj7PoXWinOiL4FponiAL/fj3M7LtAgc20Y8AA8BYq6Yqbx7mC70SjiDMcnAKRcRqW
aNaSI4TTJiUgYSpu3qaECQ5cAXTeKWbYrO6ae6ABBwmN2unXxKH42raBnWM0q3z3HY5A2eFTCdA2
08KclP9NZY3ac8uUedp3vjLj6110mzCdivhArA0JqPOcTYjoe3F39yEjVqwxWcf/PCOfQqH5FQW+
IHCKaCcFkUn2X6suwxuaAFvYwoDoRa10WPni/CrlJmhqVNk1AT+QVgEGVFdS/xRyF9tfsqeOv4M0
8QKmeudnDXRnUpSccLJVR9AFNfBP+HeSTyBa0u3Lu6cwmuzM6DooFGMMMEmvz6Zx+SV6496/VtBV
sg8Iuc7+joSZd77oj8qHRuls3WU4ozEkMWNATTyAKDg2aYZFuoHjjEmpV9EwLp35i0T9FPt9LXgt
CCBj2p10KTruys5bPlFCXkB103Z7UwifXG3dkOv1Xu4SPMKRfyy0jrCyNmqgtATo1kjPRcsVRo88
1b0bOwxEdbbQ+AHEem8gkneksQiybomIrWq3THrCIqwJivAnIaftzU5pxQCFsg6RNLzhf7LG0fe2
0DPzMClamJy+pYNmZPZN+TPGlcaQrKf1mBbBejRviSSHZ2nsoIQBqt8v71Y7RI4+osPi60S0qPlI
+LX4CwtHEywmCEwFa9gH6ExeuQgiRWIh57djsyrT0Fm7F5kitdDVKilrkJPuGtkwTuql9Ey/EUeS
WiyZkTtTJwEhL/v+pQh8w4en8Z9Xmv378fPoT331VmkHOb+0DA5+6VnggVazLMgmfv6xT8yPZlgn
dKgRZDCpq253IKc+EovpvCdscA5U65IdMjvE2RLHNs81k+TI/tmiDH1csqRSbr5ayUQCDcPdAZXK
DkyxtreLVk4lgUg1+1qR1t5Xgk6sLmgDLHOh0jf/yWjc3ll7Acj1q2wTBmN+8asb23K56AOm514t
2/E02kPKZL//bgX/fqE0BFRIeBn4YQYUSwPJ5ILEa7Gi3huoI6gBPYuUe4nmqwXR4VV4dVFQKnXX
cw7srxOF1Sg5+oYWOtI+NYcF1sBh1H3PAaA/DXqUOGCLix+sWjIiSp0f2r3wSvWqavL6otWm3KDZ
mmT0J5u8jUWApjMcnf6uR8ee8KX+tEgrPx917CHKKqxDs4SWrK8sINE6M/iro0wX+ue6LU7oReXd
XdwIVwDDmyEcjN47P8PZ3sdPgjx5dsjGYNmsIoHcwVw1bnr0RviktunVrcBupHzWH6Da6lB+/vcH
VqHt2aHg3mmUBOmr7QE01/daj0JG57kAvAapjuuTbrm+SKwaOrTZH28c71cggaHmTJjEIlM2M9E8
HMpa6pOyeQc/UL38HqaBMVHPxMlu7PYjOTxQzq0trpoBjPRzmNGikktjut1xuzwbY/IkoRoyQ4/Q
R9Oa4mpjuFAJq1X7DLqfcgzhY8cSEHNGoW93i7DVV6usPLYkLn0w6FU68VfFHIst5rljLmNfUtp9
pYzbTBQ13sfmjZML74Ti1C3TefWKIW5uFr8IiExV3mR0UeoitrXTjNZeNuFiUYOCwes/FmUK62CP
N/kgRZDM2J8EBzSHV5gd2XP12YJWk0/SwBBBW8FWSRTGnpgM7qGoFUOEDAV43mPngWhpjgEnbeJh
sRee9Ori1wB2zBQtbtfhRwUBiJjhD8Fuqu1qAu9j6zYRSJ7rhc24/tUK1s0J8la3M9PXlv5JslhL
02robtG+6UQUhpJUwO3DljRynfQfwXCgSNpFg2vYnnTE6U8OsTg8bMjjr+vFQ8jqUFjahYMzcJRK
EpakdqRvvObLqZrz+ClEJa3nm/dxeSWuSh3nw4nVv+IsxX7gUkG9bDlMgFE2s9i1aPnUBimX+wGC
0rnlRvyoj/LJ+aAo710gYJupCowCfnNOPjKQggU2bdOX22jpjAbcixn37BAFNV/2tPA7nvcEFZ/E
cUuktrVBb+s2AbcUqvxJzczFUmkwSDQAWHzuWAiySlxvh0TUG1pZINFu8APmrNZ5i3/ZcnlyWxGb
uXph/B8yE7n96udamnIpG06sDjNlRyewg7zoY0DPhUFuC1prk367oE5//5Q0AFbmpamn19ZeCpwJ
xfm0AKZBzqo3LeDnf0IV94zm1VWpLbWKEpysdXYfJuSSmJluCWHEmqhjYtqCaAUaCn5sRNSQOz8c
bn/IiAd06bugN3RlVvV7g3QNluRwXdqggSgTTylw3EADpVs8wXWvKco8Mghx2kODLBz3JvRA0pR7
yKtIKsJieuMG549oQcExWHBmDrXLXHsqlpIWLYLI7EmSLFofMihFd6p96e67VwwQj+9Tn7NPYqt7
j68GhBMDqBudJWagn2CHvEmnBoeu5dBD0STLoqJPjBEcuGX3zxZIuOBX7ebJvMMogWmoJJkiL6tW
C7NM7pRpCnumYQLRTEZAaboAfi5J9v6hznkKFImqOWwT6gxnXyTaSNrQgHen0NkSe7qVfxycj5R0
6DQSzLjzFSwkDF9V/kzKjQyCK3GsO7KXyhZw9Bu1QPUegnCHlYCtaQwEx9KRJmdovyjmJwSzWy/e
NhroHMfdp+/tmuZXUdMOdiExLaAtLi+YwBn3vb2hlR3aLqO/N5F8SKJh+xUd4vFHiMqPd7DVRZ1Q
jLACAUw4Z9PK+JzS9Et857iUrSiCNQKO6/REY0Bcp+JIMMHVrFAowq1Iu/Xj46XNQ4gFf7E8UgKj
w8IXj3IkZ/zWdZbITXtbvTuCRIG7tCupmeGBq75J3Hfgj0fyQip2mfrGSCxe42PNQPTlG07/MnHE
dQvJFGNyku55KAlBff2nCXNDy7kqHJt8aZdnvAOwDsd8AEYP11GfG9vTOWKWN8MbaxnVCBDe2WVB
QqZZ9RDt11DTRKVW2vM+F02q46+dYEFEw6i2kyvZLIN9NcfLo/7H1mUs9YzHF3/2HH3KFO6O94hO
G2DzCpSjmGeEaa0xjmx3yr6PaEb7v9DfzKZECdKxf0Y9QR6xfCB64+3oYf6PZC5E+Z2VXAWccecm
ZWWIp9tLn/OdhcD5jCQn0hGt/nT7vxOHqXZdsb098AwQLoBIK4XhGw7Hzy3ormtDn2N9NBewVv5S
YLtKYcetHvhiXln5L/MXDnhkJD/6eItwcnaxr5wtImn7a/chhHmpW2X0BFtPh4TcjliMuxgcdSkz
twOXeLHZWRevTRftXvUqJMOzphNC5SjUKcTtpMSDFaFhmO2szH6d7XeeivMufN2644Me8wgSYZrR
CLElqL55J4A041AayaJ9E57fT47mlGoad+Tyq/ghY2SRPKa7zrnCtjOVJ8+mDrHKg6ag6ptgNSrR
rXaaQsKUcRS73v6GxLoeTQod42PWmnuKBTGwANpLqLspcJXaQaWZnNF4mGYCoUZqTdYvdDneaK7X
+Lh5Z/6kcsryL/YEkOoroHbNvd8pKcxS3D2VUYYwiJ/ubKEMcNWPK2OaUCfJOGMQ0MhILYPG64iA
4OnFRMX3xYtn9XG1dDNa7cl2Gwhs9HmdUYRtT5w17lNjD4MxWJLaJ3zk/++fpI9sjFQ/WdK9y7j3
hLp+5PTuDKCcS1pqgE+8bcmfieiS1fEc2YvO+QNWNi1J4lHtVyzQw+w4oO7rTVF6k3JMJ7zQJG5d
yquulp3PUxSe5/OFOf24IgWj/mxBL7zYTGTO8Sl7wGc8YZ4+m0vY4krnZOC8NfDkWyL4BxFCL9m7
WNeclNc5852bo2kpaDAHRtaNTBtXi9CUNi7PNKKVtpRkd5iBRCLVR6NpnejbH0yqRKYLK8Bo91jQ
S2WkO47SKCHIxwCkD4h1tC7J8fit49yhWHFF+ZS2G3j83EnSpzhbQORCrQrBCE7ZYRTokqLXddZr
MbnF2PhsYb3EuHqrDZ45/XHwo5JQISxjmSII5QFNGDVflYJbxZQae36vLS3FFR1qZb+fJtqxqtAp
RPbxRzGA5xnw3epelmqac9+WkpwCc1UeXSuixvnkxhcvI0fBJN5LevZs6VShn2sgFWzqo2pdbcex
Gd11J1viWKJ9QziHDzgS5s1VN9o2ZlbnanT/dCy3Fv+FwVBIPOzQU6F7wi8UNFulhiM/R6AgdFQV
ulLstjQExvDD9eEWuq8ufRRLf5hCn46EhTJtA8cHBm7zOZXgwDwR19y0q8NlPPOThLbOD9iP1ceE
w23AgvH0ScOjRI2kGjzP3k7fAJJLeZC9FeorC7ZjmtSH0Rbm6CImOOGcCyYEZ3e/SMNDEb2wDIxG
aHdtthxUomWgnUy6A2lyxx4nQyWEgGZ5CzpiQb//79Aelvrhhez55MdAXCdjUqHe4ltL8mtxeDFk
wCoIbcAw0RAC295PdzMYJZPo+0CCn9wv35THpbyfbr2ZFSPECWMM9ud2MTtw1YTyEfnhcd1xn1v4
a96MtdBXc6ka/VPsB3yoF+MzgE+ILcai19rV4I7/i24+eSZOL28RT1eqnglHIMvHJT9o2BoCdGtc
88wdc9bh8Rkr/1YmESg4py6qv4/xwXpYdUXEEdXdy7y0PAzH49ICYj2Hf33CLq49ygjdGHtV6TLX
wEaUrSaIxNuXkMGxhOOJWpc3W+4nS8EDgTWKk4PQn0j/CeAH3F4+hukbQp9Jkv8JmQzXXRQE+kiv
pRmh7q2W7IZE0Nz8cMHUNG3uK/YX/H05vaPIrJU0XhTT+IT2DsoK/+KIzuW4TipJ14Hk5L+AphNX
eWoIpee3A4TNc42Pzaf3GPGDMMmu050Q7AvqHgsdWMeE2796j3gTs6oOk47qT62v0r1NkbGA1CJs
UtwMZeASQNqZX+dAI25zygtR23RoPl38Qk6pv+228CuAPiLs1hJl+atiTYllnpcSFAiCRKpFORiC
dLelBqkyGngNHNkRvk1mVqB/yqZtkq+Al4BLsV+5hWCG25+eElXGOQj7nMfPoUMUyec2uWU56eR0
vOjTij4SwNpi3k9ZEuOSrj2Cn4qmFCYPfJVVsbHkpPnEZnYB8QFr4/4JWmqIyKwPv4zpzFFypkM6
mVoTr0Ta15q7f3CbPQodu0gjyjT5chAaZuwl01Vj+VtGQ4NF7YL6OGbYyiV73brlDZ/s83Hk9MYc
LR6U6w55EvTzSczNaAyanQPTasWhblLe1BNHjYuPIFPWZFoDZ/fKG5pwm8N0Czn1xQt6yZFwB7nO
W7hNeLR9koTBSyG5ym6e0WigTwUZovZQENfwyoHlEdAyVRNMoYoSBRnu8wbHk87DIrubujAHY9O4
BLX+AfXcXaQ1fdtgYXCSPwLrwFRfVP0yFm1wpeRDe1zBHOoyeCd6bddVxaOGkTcyWgIyMJR2uysW
yn2rxz62NyPsL/YLzgDFNLtQczVJNcr8//u4uSsivcvwR03myCoob66guCzgrhFNpzPViegDOdFT
JVvlAwvT3keb8TacnGfxP3R+eVzcuW31QvgIw5K1SyyTTPjB/0D9Vv84+oMqYEJJtRuvZ/gpQhSl
c19n6x02BlJFy+xro+ZMskYGsAAOv8qzlCllXSm4NUnhsIa6yqWdUB91DeflhBnHS23abp5E9SPs
VBzMbv+W42lPMyFgPC2UyTYn/N6fc4u6wFy/IaeO8HEn04F3sEdZgNiDg+R+GeO+IRcADvNyclAW
9+g7kl8L2u9nt7SFW+B6kA1Sc5+B7zVuL/vK3/tmcQEqTodYCWLKoMhTdf2kVseY/meCvKJmZ6uq
cpzN8jAYUiEc30dKTIhTb8SoFJHkZNrz/WbrSvR1vsMa54mj0P103kZUsuhegLnKpclIUWYu3ag7
b7YYgzu3O011fePo8d1Rak7oL2utx1wHIUlnJNvd4kk+pC51CoJyWL6Uk/TpcxwJtFro9xgwJHjb
V8/ucXfEuJiemroPL56wx8J2YaM4aVIIxpAtQP813KKF6UhSrBgA8Vjp8PlMkqD0R1+YXMrqTZZ0
lFB2V99MH3EI+qN3IQOGvqKbB1Vg8YSG2LajAaiFLKl1Ub/kr1xuPJshM08x3Yk6zxarTEqNB5Sv
81x3aR/bFhzakI618uYI4Luxn0mCNiPhmJtrjXDrrM2mSPAChJxU2vcnReuTHzySNwAF/20XSMyg
mWo8ywiXQ5+MwBzWdifDztufQ0mDIzXNzpTiMMgty4whdrkbb8tgSFJ1xAHXN4PRjF+9Xwv1lQda
JosAo8x0DTsynGzGd2ZlyhmPB/9a2uhhokIHfcV1ZW8h8hMKwRJxyHlqRcDx9oKntGp8TsnVOFYO
2R5MbJuL3Q3xQDG5u1szBr6RmsPB5fuBJjh4zC/drbCubvX5khBEss6lsg+6Ppwd37RxVmxhPBW8
qKp+lSEQiz4N+W+a+AXeiTDAX1zZszXTYjsdRsGwFPxdiujaBpYNe7UXHJV6VB79sMxrcg4gqPKn
T0YxPg1IdXmx4jXUojSAhXNtUxuP6e494zi+Zf9wcZ3+O6Yy4zVBl6MIz47JdpEkvwTlNDb21nlg
EKa6C6aAB78HwYW4T9ghSCzyb+ZvI3fwC4+D0hLrdh00bnwON6BN07yATSwjdq4qqS5sdQKz6Cw0
luJ+l0RhW/SLzcuu1QebEGQkSlJNZc/mOQWjgF9STqtJhSeDwinMDb/V97CquW/YGROH3V6zLx84
SLXpioV2YEL5ndkup93i9fZilaoZqGSZT5IH0KAZefG742IXLrw93mlhMolIupjDFh1JqpPFjLHc
aogQoP8ltfGOlX386H6ap0KspW3+33pJbQwVGVuIIAGg+SZvaihnlvtAxgKp7Y8BsvSG1XHzTtVK
FawShAs+0EGxwqzE6DckVoYyaZ7KSy1kJyNkCfgUlR4PYBPXG1V9Twb1jz58MeBAHV7f2oFSDuul
3I1NOwh3KzKIub4/eNJdwTlSyu/WempjuqQLwoNvqrRezjcJyq2HJ+WLHmyu8I9fJhZ3u15q4yBD
UiEWDfxAGOCpqdWuOBIVfGZHNAgOtAbPiMS2cv1ENNQXoXytI0MIt+QwKgOpeo2sN1ArX4CZs8gv
uevHCyBncKSVv5aF/R1IexwaxM23/Y6k1RFoWT405jRxZ58yzAL7oMZmyiO+m45vubSyPn2QZ4wk
ciMSXb3mxjYw2kEdY3WSOHR5ngYWgrS/1mEpYfmDjLwNU/fhYwQ7IaqpVDbguL5CQ0fX1m5D/V3Q
KSqCqTNZX6WldW3XK9dFgKkVCM05i2VAgSG8C/aQjPButLSf0K77z5pJtsV1aCAD3FP4AcTW0vRu
Dt3ms5VxiVo/7+I7xbcryka2vfuil1pxzRMDfZxmwxrhv+ufs4lVQvbpnLvHBN2caW3MdW4ag3w6
ti0DjOLPQmov+y9l4FyIq0uOeyVkB3uvZN3PGrj5LTOkaDlOXmZ9Jq3UX6MOcXkewec01Sppq4j0
SvfcLynEOEBv+2eFrLHfbs0Nf5iQohXjWnUHNGZVK+vBFCRzOlpxpguYlHvYdEGHz+zEoLIn9MVP
6C9zf1DzD9WO/YeP0nCW2H3vAbKiNflVSPvR9TBZcfalqU/NIhu6p9NLVDK7btVP4khKNRRtheDr
gWLodY1HugGRgmxPK0xwtdJaRhS6TbpiPlmEd9GV9LkV6v0MYJRX0YT38+eCffdB7JemQTIMcvlP
AhQFpPyG8zcpDfsGw5MZLekfpNegCkuoRmV5Lf16jSWi9yKYASALL+rXpS2v4PdfQzzf2TKgwbfG
kjo6pU0S5jEPV63OMX6gbsIZUnjUJG/olLYR+Fc7wjO48P6HDPV57VSXLCyQRq5YvlBJbBMD4Vix
+uQ23cnkl+C2lC5fwmo1FD0GnfaryKMQVRn2gzVSRJ1g3sfPMzCdjVyG6TDLXhz9joztZ1VY0Rxr
CYEmPyMFeVnnUio7dLsEtW/IutAXlKIXUkJIIfzZh7baknHuDx8hg5HROTR2eCea0wLQ5g6N8AYP
hK7+TaivIaVEGSAGdY/kBres+YCeGDkEG0wCRPbM7Pw6TlOg9k2HcMIFhSQZ8PWOyaB5ezRIb4VY
UBVa9w+iLspktzIztPMFM4uISPw6Rd4Vp3VZzvIBdxuaxC1u5AeGVTkynr/O3z9eF12TYPzp8Zvo
V8sFS+mJb2Usw2RgNx3IKm2yCvZU71hQKcyLBrrEunIBg4v2oKKLTP+URCN9bGwvtug3bRFe3ODp
ojcniCFhleUD4H9i/pQj4cSt1GOZKaf+g7ZCdYMBV5F69xS73y64aC1NpYIm8m3ujVTYKRorNJ8p
Gk/v5DIC8uEQblLzSSBkm6PajI/DhvBStAiWI4dw5h3mXxNKImn2zd42upki+WuCq3NO/TunJRw3
LbLfL7Dqa6/XMG+1HGq4o8M7gZ1UidOhqiV3VF1Pi+yxcc8C8airIsm6VFRZaC06/HT/xBiKK+Ue
hzo6MzVVxk9jmEG6kDp4eTnQKVckiXTM2ZmZ1F4w/SFhIT2+3G0OYl7HEAUjZIW+lCIUlSJ8P7to
m/dYqtsSFBOZ4/kfurEKFTeUTV6ZYRWIK4/ddVt9dPqe/pRWlBAO8u13zBEDr3tNxoZdr3xpzarw
dDq7X+25vmn7zPaJzZAbwXFoX3KRQVi8g2/O27i9wnKdDt6eUdl+e6j2oeKB1J7kiK8rBkmnkDoU
xufqg+T2f35mhMQNPkCPCGC4caUlo7EbQQ4E72DkN1PosK4/EsyeZ9OU8jRhqb7qdsSXDVVFPnEA
rijBRqGk4m+q0r0p6dIVTm+USToEEwpfNXIUhLnxbQoDJWI0Uvg25jhazFlbBKqnvY0mPSgR5nGo
9R+1hEOBX62Qi8giSfZupmKjQ5HM05Cx3j6YHGJPqACiuUsXx1fHwwdSAOzazwT3D79cZcioh3D+
Gr1kNeuhubMq8KyVG+zPQPr6pUlHIAjyCXkla12imfBHNZzNWNruHEsT/oHBZvc6svKwXkMc2QHP
zBh051dTGRTS3jdEJdPCZcpjgsnMVc4XHa9xEF/jOUcN/njztn3W72UOexJlmYEFpWTa8C2sD/KB
R7KkN7m0OMmVF2Ds4yxKOusMmZZiqYkUJgqNkcbs3+XY0s61kk5GkqBvGsREvOlGgS3JHhvPC3Z2
HYYVX0om0/tBE0I96YmnCLxSIxRyToUFm5I9aCWy6ZzZnkijb3Q1AiPwxZyBcrA/kHIl29kEOpWs
+ujxslC2QE87AxiIqx8AqovlYZVO3ANtXjehgzWMk3eTui/4quOGGnGnukk303RFnwvncuTRJbWV
jAR/KrpUz1BMLsj8YcXYWBbjDRaTgzfiqXltOcVLMgJ7ZjeSgf9HTdCMkMPCNcMyBQm77RR1XXaJ
Dx8orzvtAmWJaneac091w7dghNBcaVfAscynYCu1F8ziu91cYYh/PgpTVebO+OL7p33/eq007sC7
YANALEoklS/ZEpKEwqEvyXdeGLjbtYQt1QoYrLZGcBYMycRKRU2NKJxwV+xCXlDg8krzKFS7IDyM
On2GCcRyg7BHdmmuu6o1IbV1Uvxb/5STLttFcUf7MxJePLJtbBaxDuRXJvLqwGfMrhwglqRAWmQ2
u+6UAK0CkiA6wVkHRVbHHgIa2BmNwK2bmQWc1OPYvJZNNzWWGw88gHBPcybVdENZkIlyKmyJf9MA
+Gug2vyfQmbGqat9E2Q81ZAz7qz07ZQJEL0nG5jjTiqfCG49iQ5rQtqdaMlmy3HMiT9COYNY7a7l
8UzkivrqUxhuphSTn34LQ0rn+wRYrJGTCwTdta98m0BP93y+48il4Mvc2LWyzbfZiiRyMi33hMs6
IC24CsmzNiK06sYJOHvx7vItj+X1zDMU156La7lB+sQGvM25fngWjnTg8yXiv3o0fCrYyX5SQqPW
PCjUYiywlpiQeIvO/YHZCepNexY1GHz21XO2ZIjsvcf5rzM7qAn5nWY6ooR5SUT4F6w0wTCMY44c
eX20s8XKTJr9YrnEplEFhbZnsRp+qMf2yGiNT/jWAbGTyIx8INZS3qzmy4nAjfKesu/RUqpk4Dku
gOLxsB5jkEW8Wx8cndvvytS3AscnxGjgF/gIQTZlSxuEwagjIGSfYpwzv264zrhidUNc7pC/4+YK
e6CJKfUoJhc4yh60fY7hnMvxNhpQSq26TpET0oPtH/Q9kxUmLd/yw3gElVPPAfPN+xXPre6msyks
4qvucewnFr1Mk3/rTcMJw5WQtkRW+Pl/sllEG1Vzlka7rB153q5Qw4V0loKAE1cnPSc3V5rX8K6c
imX8t9GresC9pgj9oKfDUdVd95J/vQizwK4deN3YMrVkFVA/zp3vBrjN1H4h7g9wDNauOeme5ak0
1J4rbKCi4nyRDR5ZY3xemnXvynbMiDa7nam4dhjCjfc+LFWuZBrSpFzLzmLo13q+wDWo+gLjv/Vo
bnXEXVndlkQ+Lsy1sgWTUoVxQ6oojkKxa7C29HanVBBCoGoG5EYAYn9Tscvik+GSmSxBgj1mc8io
hXBJ5QAA8Wq5Lkefz+20erEwixGtwElfEK20t2j3gcnVlYkECDYBV9DNMq4DMgZOgZdOLtbKDaNq
mshHcC0NzUq8R1pGaQJpLVZXlS9xIqqYCglWoBhGECLFaZzjzvRyoY6pa4fCwHk0OxaP6/w7XQhK
sq15HH70uyqJvu4+IBo4mK4Mwfmarn6JGjUEvGMMmN6eFRM/+bY/CXbC1ISXG6OWeRmowO1IgzQd
2jME1vJVpINuW4Q5ZhMXlErP5I+uEFKSBcjqxYw0ZbEpXGAJM60OrlODmXoXXR7rSzG6Zo0RHIVQ
wz4I/XtZhqH9OpskraOmdeb3zidUU9ZFdyH5GJ6MB8cgipS/ti6iAtd2vMNgjX3L+JNxCFRywjAF
On92EAu75zFsOCwVxS4DbmOJVyXsnNmVW/jxyCbsIYl4vah3M9f63WO16idN13YMgqgqzKaJc6qf
KZCgC/WQg6ZVzIC3BMdx5quV2C/MTq36wp59VfVo1Tp7/uDsOKoM3lDFepBpyRBMEL9CtNawbpwl
Wu2WlhbiDse4/9A4gfH9d1cLFc0aULeqfgg2C0T3ByseWlQV4i/4TKkCaHKORvkBJn/J6pA7YTHU
pFMzsOC/U61ZbQ5Z/Kskgc696Y8ENYseQqI8P3DDPHv6iFNjZ6Kwip6QfSOAaNk/7VU8ZV9Kbday
LJyhVmrALdg+h3jxa3uYWZy41Cq+PLb94sXqZ6RbXf/0HUgumPFMikD9Zi3pjM2vP3ii35Wsv0C6
N0kDNzqY1oDr7fFDuU8NoI0C4MfuBfEH0lZE4kquDk/1cADME/U+nRCRlgIohdeRQ1PMv92siuuG
/Wi1qibLOk89mp8GNRbowgsrBNr82LQRpa1ZapXTfThslFCGwBqEOOGO8miz0+W7MWuu6MeH9XNh
x3G2rUjrHunh1K1yS+YYx+khSWJd1WcXuPbN41IiNMmSIfnJS5aewb1ZdfJuArUA2yoPm1U4Sj10
O7piER/p2Zh4wlQ2Rr/H/uvffqSboPpo1GSyXhwH8W7X3k8pG2euBulw9eaxcIf2fuMRLgUgNxl3
+16KSyucPTm5N1z0IUI8EClguKNEFzEB2KPutGvW3OhGwr3qp8Caf1KH9Jk8h1LGR17YcwGfL7ey
IaRIaFGxG/5oFW3bAMuDGnnL67UH+Uw92yoTGSd89nr/m93Bqje0Lu776lmyMVg8SWUsqoV8bxjE
SHcNss/BVQRgJqi4njXX+kqiTTrE2iesIut+w4OGq+O1GoMzqSALSXDcYVXQ71XphZMKf5ciOMBz
ln6fwjKFBM5Cf5YO/EALqgYQ5dAl+XVq45EH1UibA7J+s/fM8hLExFh+7F817xi+JgkHx+Xh7COu
nGhvf7uuGu/2lC7EkwD/OjO8UPb9DwqaEz63TPIBidoQTYECyEry5g5ft4///SCve+5dUIDGDnsm
TqfOkBjGgs8rYp0j4RxapNJwtXIVRRBVNiTLCVOXnE3XuEXFwi1zKGjCuRSS1ROXo9SyneRRV1QD
n/ABryRRpPylkL8jO2brvOgdCwwgqIN/my2n7zzNkHdV0U/DqJw+gksh0Cwi30fgBpJ7GA+dJts0
yKCHurUxRvHTaZ/OApQf/SJSoXf3C4UaqHiPJFXhgZEc5NJi6aza3Dt8f5qfD93bZvbhCpg7QYSR
kXp6eXtjDhZXtFxdgj/3v+mVQWcbxRmpXnfy8C76mGX08MMkUi/nftYYfQXgvB7s+zi6ogO/IBLB
VC034MX+RrA4EVR+Cyg0E59PlReOjt4WNCWj0yLWn63MZf07zy8oTnBXE7KVa1ZdjuLBFjXnHwAf
CHJ2/xKtAL8ATz+OvAbvNoyYqWmeJd/FIqVygEz//40tSJYOgo4KzwJhKLoTzSjj+P0BgNgAhbYu
uR4VcJ4bFpRvVtI5fmlbzf8vNGt9cPFyPlzVHyyu3HjJsMFDkks8j/nHmK4e1epY1mATCqDK3ywI
o/2yo5zAdItfk8X47u/sHMGrzdjF/ZdNSP3fBicMVJ+/mc9lbQNP4DlkBUPF9X7GmcLgW97uHqAR
WEU5J3ETWWzuBbwbyFIjTuUh6zU6Gf8p7FvnsBOFtxzsEfVN6uv4vuGVxpY3TO0MGDZZpOw/FkJ2
HXpR44c7Wvj0Ly1cGyKnQ8qAD79b1+FJW1o5RMl/hcEDwz5jpdZEWlszfHmvxYiTloHm4E2ubgf6
YBlkBRRHuFhN2l7aEQhIzIbmMCXWIDDpfdjZHufscr1jJhenKUgNJ3RmhJbAHYtIZT8/UZiTaszP
B2Yt9R/ZrXQPFKPSW1+zFZrdKXANPAP4zDSkhi6GlmwnWyMfTBl5kg/rYz5zhe51u8m2LuM3ONyk
O9M2qp9i+3cmyxzcoZh0RqQPXYNxzp457idzBV/eg0yQrHd2U+ngJzK81LSGK2e81c7TfpqNU+fc
Oxiq3jQHUIbh8wsGchK0aRt5bdwkRearxY0psnxZ0+ISFRW7YBBU4Q492Q9FClXQ1G4Px722/GWw
MjGnVae+xdCkE63UGa85KHkAVDAmu73d7sZQiqkg/OYMAJ5Qrr3H3IRbKqOBXv596ZUsZ18l6Eck
JNFkWsCMHkFq5if/n5nNa1eTNt+LK+Uky/UQRLYRt+AK9K8j9Dj7ZQOBJSPzs6pTuVS5q8EUirXV
HnSWHpNd5+U7Md/HO2Zix71yutoTAcCbVwgN3Qah0dSiBbADWWhQdbefPFG0T+GJC+NIAlxTDAJR
QxDV6TcF6PenPvPU8BqqSkxWCHPti9vipEFa4btFsTlkNstFX0SEdtWg4FkfbRF4l9x3o6GGZq0h
q4TFKnJ6l8GbhTJ8RalhSwIUcwt4Qzyn8an6iaSHUjEe6F7G+IFKuq3agc0hVJFPnZB4/MzuDIxT
iKdDsYYy+iRJznc8oLH+fXBawLl0s4+xPBzkzwgWgsKsnloqplOKRWbgI2jJBvvMn7wjL6t4rfjx
VPsU2vhKf8CrYJ8pbQrKHb8ivN8j4cp3z8h/Ji3QEnRmswTCnCnRQv1DNCKkQP3O7dzjw2xI7uay
XWTDdrgD+Cw3iYr2upyVbw7G81R4uBXUng1+IKwN8JLEWW2nnGUWMIzuwWWhgWeYyEQzqX46VW3E
ehuGdii5ozOvN4I51f8yXyAmya2jFcrsGWPMPTUzHsXrn8q2YALQA3J++VNBCDvGpPQJnz3bbevA
rgBHjjxsCacthT+l4HlbnqkiB1gEuzbM1IlxHvjcUEMS/BL8ZRQ1qJOfADKJaijNlBWCnM1BQRK2
36XmoQjbT7e2jw5pPEGRavfwM1S7r6ikVQkcyMOIEbTL4/7o1tzZFp4CEnAiYQsfu+ea8b6MZHft
mHyJpcttwsyEcZcyrHbqcF/lqrHlge1yT+hYu2Fy0PYA0DZR5mdHNM8NPRxH8yx8m+vH6wJfAtbG
Ao1jkPr/+STyiU/H/lw/JbSye4Ael/UTR2on7/x06I1KIpTcXzlXbN4Fp/+ghlIKRzU6QACJBIRg
N+X7NRGVqC1y1VgzFy+DvDfoIxWseuQv0kkfRQLbmIBLglhpSQb3OQtIOKZZCcUE0O/rKPiTCGPQ
2hM8HzTIThtf+f1ffOE2VvlbxSliRSGIHdTxNmBkzdprYzYeT0J7hPNgLRZSsbhWlXxVOtk6vCN2
l/NmabL0lvJJnjHe9wwKeIbqY9Si9jy4mo48eDdRczjbAg2KEpz69SCUv2wvqEnQ6I0fM/28jnjm
BWGf8jhRJpaAijDTFYRSNs6qYbFVyiIYk79cBAHwfOhmUbmrKLuIq9AYdQQQTZ+xBMGHDN4DIQOj
PCJqGVv/PHD6QhmrQ9fAsmjBOMfbz6fnzyqRqpQtBHBBGrrzNOUcGT9nubf7utIoeL1fP5vOp9W9
e0CzdnnFrL8QNWdp4Wyl22yVvN/BXKMkapNECKeL0KLF7I1nIRRSfJWmIuRJH51ucJBdzFuZMCu4
BB9i9Mo7JlyIy7rd+bs6mQbButbjHzpNMbuBFip7zpV6hGLMAiZmdnkf8Jzkxs0RhBUa2rbegr4o
+fuMYT1IDV2YLzbXqTR6V3Ls8haerIBJK1uSv5cfnkV6pPvQ4T7GbwHOZUxasRzuhkesKBMK6B3C
/PV1spNYsHR3S91quYVvbnK2tAl7ZOQvw75dlWkLMHWyvHfIH/YiVhe+7UuHzuCdK3C0vCnVTx27
ZwQyHcdVNZFc+fkxdKp2zYlQGmiP6xEUwytleZ+a0U+GlECtGoyCy0VEo5GP3teo9S5blXFEj5y9
ddMBWhPcCoCNX94g3COhGJiOpLf309uArJPw41NkicpAN/IGHSw/xVk4CxX13Kbcq37nZbVEq+Dv
DrFJTcdk+cD34RgBYa6GWwhSQTICMjKpe6HxPCy7Z78Mda5F9oT0XJc9X0NQPv8nGpF05mMHt00q
46ciZIlGLejfzUqWEpCFbqwdOSzCN0QWOUy4KKm7M7MTP25C4/hVCrhAc8ZFSjOX1Li2rX5uzEyG
6b+JW3lqjhq+Gra7jNpqdc2suC9NXZCfzzeFX27QlPJSDKArB4MMX0u2cf5rytjtNP/3eZTNFl6+
2JUJly/TlmyLpfmwSjIys3EaQKj4wkOlBI8rVht5MF5Hj+9ji5aM2fFtV+E4xNULnURNUZA473XM
pq8HyLyzyUE50WcjzwasyuNSmnUyYJJwYAigZqXmJ8FXvhW0ykh/Ib5HoHUunYQtQjQlCjJoy+Rw
kz1NpB+TvU1rC8nRm2ArB35OaNiuGlxeRd/x+oWY0CYclIpHz72T8ZpYkBQTYk0gM/GR9szXhX9y
kibvEPxNY/9OX9T+1Q9HIFHRVzWxklieJ72Dm8hawooUvYWNmltY04Z7S6LsY8NNIBljexXdIpdE
HFmiRa34kKCWWmgNtSXT5WJTHqRKZvmKKviTWQtuyxhgAjL/2FqwBHXArDknoC55qXyJ3aJRBrwb
uo7nC3uZ65HMP0yBqFKHEV/0uMWL37Yyun5dHS5jfnwsJDluVWmSMnKFDxlSGaoQ2CuD83M5qPSM
wnldCxvii65uh6fy48kuSarGwjVefFk8HR8w3B2V94kh9VSjJiKtd1gxFyok+lynke9cmcufMnjm
Xfav3EZIotGFpISxx7LZHLD/6OyPscplT/p2VzKPcZ8IeeOl/p6zJf3S099dIx4VV6OGFobAMhPI
fHVX6R9/tX0maSKtIlWN5xrCTXHMMHLTNp8eHyczv8zZCR/5rnJDMAYnqECqjnG79GZsjqWnSVqQ
FnQjbRj8+7lwtJ9YWOY3n36nzQQ0vTN8Mk1h2vS6p81RxhJ/E2/kqAqZQHwTi5S+YK1KK6mOYTE+
LzM8HCV0it6qPIBLK8ledEKzU2uXsMa84ZJlatmbGoZulhq8/ysVkIKB9OQUHWx/FUeBTdNXG4Ju
pPH0T+BwPVou23wCYUADtst2h1cZlzKuML834C8gEhvnH/9+DID6lFlNmzBq0+8l06vig8T2Fc7i
qI+qu2o7pkqPDlHbW41A05G9PqV04v38m48Pdi+7tV2bPxG2oDKqsraSerbdXBthZ7rR/PtSM3lL
RLn58glRjA2P5JxiOHdkIMlUNuCp2W6aOgd/aVswccOmyiQ/J885+B3oNVRFgOd88nQue4SIFWbH
iAGxkFqVac7VPE0ZqWnu2gUloc5XcTWqa4dgGJ/mTZjg7RlOuAGURRw5qw8zKsfDP91bCjIyG6uD
zordOI6ySzSkTo/5GbnRRLM8q759n3mXWTLFHm0bYJmGlXuBaBUOSc6vh9RpfFClnUpY+wCZU5a3
AGu1Uz0L4xFCo/mBlWW7NvVNiqIVJjYAkycIpHta4yX4l4xvvXsol8Y0OvILbzgbKxcpZs+Y715d
aP+zF2rVMcZgCFbkODkrSxAj2LzBUkgDOZCVreGGsRzNZ/O4YpCQvIUHYezKDkZD9vawYJ0QpYXJ
bqICT5BZz7zwfC+WlgjgEhHQLln+4rOYI2cMnDrkQn1Wf7dwI1tfJMiMlOP5cuv6dUSspJFF1ZnW
bMlhp2hJnY6kniAJ4pbvn9IXq4z0+a/fQw8IK7mQaWru2cMs3rAtzkgsBbmtNeMky3zRdXD4wtmQ
wiJoGCOXC83jwURgTchAuU4LG9TGtZJBByZ8Bya80dbzs1naw461FcNQGnUJedQeQHFvWwUOfYAU
RIL+o6mvdiud/GbPrEaygdIEbb/I6W4I7BAFJJWqBenCEatitxFpjQEgj6AG0tLkJJJ+2NfNiYxG
bCwlDPTtccldt44mhk4r3LWpyqq8s7EAirWFKjMs8DEZS5T9Nr5qoJWVk3rbDM/b0o1CbaQf8YN+
OBbuFr1bU0Z0cwr5QXpFbMloDG8VqMwSZfBz98V6yPM6SmocIEbZiL5jWEAejjt44ZtRNboaaMDz
Jej1BEbZNaapP+PGpL2QIAiZjGgIpCUW+coRNyk70D5vqqmXg5Iu741fV4seeK11H5E4f0PZ8nei
gU5UrU0UJ06iHWDID2w+u5HAVTo8atFbOR8olgArHx20nY9MwuWcLQhY87XpASMQXVV3cNVMKlsT
PWMA9Mqng47bJOICTMi4Ab/FX7q5oO1BYwgDGN/xNNDi7NZnefJXidmbom0yL6KXHKgn64iR5wr2
nVqLJ3f4j10hOPJesSVSPG8CchVxYgucSRWewasf+qdbo/APThWyWOizUNIlaLuIX4F+Z8kfQla/
AmV4pzufHB609Bsz5fQ3mgAnfod30OXVh2iCOci+7qo4sK7UlgpZuUBKP+eRLo8eetB25Sbbh7/a
CnI+TqhfhZ9COueLL35FtO+Om8QoTXNYlmYd+NHwxyo/P3OACAksLgdm6VNziBbR4Dhh19WScnZm
sWJ+28XEwxCg0UuTuWcTBWTVl412tVyXCDanVVXOfFpQ9WyZZ1aoOiDNMJ+p6BAlSZ7J2tMeEvl5
Ge9LpygeC2F5DRfy6+10K2/MCtY2TbkLbJ8PphR0UcBvWc+cejabVZtEZh5oV7EWzmKFTQ88KhzK
MujhIMMP77fPvMe/+1Gvfm8yqg2BFDlOXFv0uGHLEvbNBje1IUIKlV2xfaxmfC9qhBHxybbJp1Ho
kb0RyvBntqBgKCzdKiuPySE1PzTugBHsKqvb2HKNJ95mPyiUZPpNafqAyQHTWo3j1chSU7nbXL48
68U08CVEjmVPVKm000gyXS6YSb1lami3RKWtM9bqfg9fIW++9wiynFtvESJwc5O+tUFPI0bPmShO
GDmpXg20m2TJAwTD7XS3bUiAhvnapDsaS6vQo4UppM4dmuXf2/DP/70z37E1wuVE8scV0AphOCZk
j7Anqws5TxQykSwz1c7ax4r2f/NnHrfhYWVvozGv4xf+l1SJI59yQU3NplL0mZbsjtWhtKKBKgct
wjYVeyI1KCMIyYimzH/JjZMgYgVAM057dB/oPC2nuaKwDZc0mUq6nBN7EhgrMRuRiHuFZGzmDkSD
vYcnkx0PTUJDikx/mFY50DFj/Ik8P4QvQQBKGHbzT+TZCR7myfhatIthv92LPklt0lpii+uPBO3W
wkLGGR2+dzXZvrm6YKL894aVUx6WS1r6v1NBPN7CGSO40+GMl//ZYRWhBswU2YK6bJb4g0fun4H3
L3FbJCupDDQ2aCrWycgRE8Q4Hqa00ZaPuliGSHpRTfa+EbvOueVwzpl0S5X8tFsKKOjgrIa0spxm
jEYzEjYkoZHMrzKg2HkihkILyAhzBUAqsbgrpGIKZJ17a9xLZqpX/Ga7FvZQ3OzoVy8A2U3172wd
ifV7zFrcjwmgJLW4aOTuM6kGJ/ZcId09AdsbOBkU56t29IiQTP3HwNWLmHYjyv9IbCVqOEjC2Fhb
RsoPBAeJCvtBfPtt7c9kzjoAPsdbQXROjAspQ9XfaZuHz3VHWE1mFYsIiXQ1azt2Z2jIEYJrDHcm
Rinm8mASUiMKduVWGpkFhm3XYguSQLIUKN9X0NhsS3gDzUQFyPK1ROKka495Y2VwIuMKl60YrY1S
YDt3L/RGmSK/Npvsv8QWC13ZAmX0il18e6sEbHAJaZkfymV123nk6zbC5VNUMIp4Swiy1XutkShE
ww7uNPjVMl7fC3npMJ7Aonvr9ypQL6AcgxmXvi8frfQmJhDZwDabTIiMJP49Cj9qF68GNiNCWo3w
VwA6CDCf7aHRQYplWrmly9vGTM3eW+Jx2DyW8csAIYE/enDP7W1+PycEFBf76ecf0hdN25WKUZS6
ryeKFOJRST4g6npASXGI2Ch7q2/zCMLmJU88k8G7NIjNM4Ax6mjx1gdJNZkCmlhYs0ZESJuCRMPA
dki2efMvgKf3DEr3eufd1KMI26HdvGN0XcBbB0TKmVUTPHTERrMVPemKUdun1X9UsURa9Tc1oPp6
W5mK0Z8W+kyAsOsR78KPWD99YDANcQDli6OJd2X4dYgeV5MT4iQGxXPKqFG5vxuYCmWw0covHrJS
YBFLn0l10HtfSw4bt0JJeA2XIwRcZEbgrRrgzrURV8IUvR+1JOmtlNa6V1419rxye0ztvD8XIEzN
5yOASNokga2cp2jpivr85cWZb0+4M5S47hP1sMSwh2Ujy8kKQl9q1lv4N4LQvwzFJPheXFu0mze2
nWalm+44rkC25P29WOQDWPhbKw2Nc91Kk4gwn2MeQLgMNnq5sM/GlobxN0iD+qJyPaMXWHUS6mUN
MYme8YReluCv8J6sogsVHKQgFqy0eW7Zy2Ga8JEl6dgxnaezcHNhJYsR/eW7lRIowgfYSSoP0sIx
ieDsIEBGTGnAndYch28h/o9IeuHj+lbNezeUMiMLeGwf7i7dz0yPWZUjBzHBfz2XUM1cOcfzojnU
2AxXds8soILXJXYvtLTNT4xsfdNH1hw+Y8xIIcTLlvK1zh08sgRIMXPhKGm0jhdih4bu0qrHip/q
SIpzm1s2vdso4maa5qS6Wi2jyJv/IajhMgbLU/LusflzII2kzXjxy52tuJoI+q8NyHk9pdjOowws
5fVIH8lZNFDmKd5vyVgJaEI3vl2HxWu/LDz5keOsqVA/GUF3UnHmbHqo3yct/E7wfkUYciMHEj43
ef30IFFNdBqatlNTR8B0g90FEmrkQnJMvcGzpafhMTu0Khd7dHIsPDqjxkWIs3JhfcpFh9pcjU3t
39zBOK/yEOgDyFyySaM46eXFPXiQwdtJTguiqjrPdqUR+O94ry//tK8evSWuk1GujksV4MgarWsq
ypkFqme7Ptdus0tdsPLjbLXMfkJInjfOEMkU3ZMFNO9Hx+OsNm0huPR+Fw7jDvTUp8CCEKVJR9DA
bxMQ/mhYHIxNvcwgzCOMDJXp8BjHpqLy+HNT84nH5+qBdLDODat+0p0MOG4qHHH33g55++D6ROjQ
b9KDOuw6GSrO4mWN4IGPEZiNcyujd5y0oVtJiJfbM6rnHytWDG5mPKxlcivB3RGccAilS8U4symf
5ZRabHIvSf6kfBoglq9TWsbgmaDksSMiHrCsjZGI0moDjvA4cnXqdU40QN2uzok60BwPpqpCy1CX
MiiuewvhJJFrOoGiu/LjvuOa/lQajJe/k444KvlqqldzsyNToQzcQf9b9H9uE3R1S+Q76Ggk4hQO
JiiTI3Ksx6VDFPpMfHAM9VNUF+bShcgqgnN+tCIQUclkc7ccWS5XKSAAr0hW5F4wsDAbF5vQm2Xs
whk++8yFQx9scRpg9UNzQHUae2HS/6LzXIIIQftNYyyLeAPCuvp6IDBasQ3+0vOLKwtzJl0W42aF
OuG6NojoHtzi2wbFFPP4ut/MCOd8s4q7NPGA4BJN+PByHCWH7WQFQDTkMf8gx1w2LNGIVJfGxueR
dLRhHEhtIjGSdT6RYBCJG3rC7uS7red4Wj4EG54VCDIoNijSWogjrcBV4nYeg6cb9VSPnY0QOh8x
G746v3X+VfgeAfiV+ScFNa+ESf1bSpo72hh13j1UqpwDrSI53SODPAdzswCPWOvgQ0jyhU9kvq+m
ZYx0T4KMMCtfhrmfnSMGK07EM1cDls60TS15laWlw3XQJptyWWV2wh7vjt/TKlxHOh5wShffzGYI
M4+dbwayZvg6Y0t+Th5YHNS4uI0KBlniHNgcAK4SuWZtSh6XVD6+s+JcPdK3WOXEiuYzGU+JyENJ
vT+K8ifnb61Z3lNT69Dtey0YFADfl8ivy7RE02Eg4vQmXMq4AxbsPJH16p1L2EUEzk6zFpQ5go3x
xP4ysTxxlZzk7jrpvOFnVnFuzFmfv9Q/3owbGd7kpTFBBWNsIIw9LB4ytbViKyZGkDLzz3FK5BqR
YlXeElta5aN6G3+17mseHkPb3AiTgaUshNKRzmRZlp+uzQ4vvBbpU5vcdawl1t4N16fSqAJnrQra
1ndf/nFUtOBhpTchD5ZKJK+ClHr8utcC51jvMbkJ1x6BaGt2aD1kl+HaPmMd+uEvOm+2TKObt69X
5xGomLR0XtYcUTHA+Jf1mdOVpY4o8sIdaUZDoI/9LHmFbw8RYl0SjYv7kquKXPKzyqc0FoyttVjt
5B4uKGSadLFHeGNO+P98+MgjfFingKPAhQH49m0FcqGtfV9VCi8loy383wpjXOAg6xQmMNOBrJ1o
1aY3Y4b1SSeuFWWAXK++zLBsCfultLSy3XvdBRGve6/UmoR0MgSyXaAKiFWxKH7pfCK4ds0ZVev0
Lq+mzNoOYsKc9JjgWJ59nwXfQ+/qTQkTMOy1TJZrMyDf+/Q5OEsSLZKsTv6uWCj7GCHYvS2ZpJZ5
ln1vU3mjftm6ZQ8llF/pdC7M1fym6TdAqtoVjwWPQv4vMJwP595VYr1DYaRA4g5tDj0WPodyG26v
pbNVcevrkJ1QNf5Q27IoWMEix+ADJAynGUVyTFghDMw+1Eecfj+hlZWc5JZFUu1p+Uey0qxjCByf
xAyQNal+u4p0bCBjaVZcj4j1f3zkxhhPm3AsbMQ8c0t7m+IL7dE3NOJ1q6+rnYdEjJG3Fvj+yMi8
PKYR5rmI/Kigjz2ED4gyCldd7kcnuQ5ofmSrAl0QvG5hQ3HbJNunzhwKuek98O45O2dGEBaZ9kG5
9dTTHj0o0QEdJLyMGZyXGRDg11fgvSF91jtAnECoyWvUrD81qcj+OfGTAH7OglT8c3t5RrMG6+AJ
nzm03PqUwQx6med5DcQW/izjmd9oP1MQoF3CvEOmeNnNaSOvy9Ewo9nEboptftGbGrdgNdpQVSO/
LjrYI2Gqackt1mOALyombi1JNiCtHMveXG0D+P4x3TmBEbZ9wOXzh5H19nMyufrMGhzDAS4L838Q
PDSZBHTeHIMI4Kx0TDZR2j4vNA1WldIUqJaQjbj2AK5ljBxeiBO4uWsKTyJTHJe1IeIqVT3wiDpE
6LpEH1MSMPYzQkrFIKZmjerkEgXD97mniUYC3wvqYO73+oPkQ24f18a2fGcEG7CfL3vrsQKr+Flf
lrs8EQosOCDjlPqI3MnaG6UsD6KFKRmUkGUzl1PRQ3yoQ3Hotm5OlIZJa0XZskq1EH/jwuEuO7LJ
y8fmjw5jNea6My22pPQfMwIkdmdm5DzuMcZTFgXUexzqGgifb5kwEbulIHVXUedYGKElH5giNggE
cuhOVxSKwlX6X6C8pBhMat5I2VDj5IKXkad1aMRJygTolkX4YOP8pDNyQyOIrbUyr8e/eCLaeNrQ
8KuZrgBWOfnHWgXAqW2/hAZ5Q0ysJqM7/6r5J6F3vFO/1L84PJGd2UugPsQ5j91ZvVOEn0eZprJb
eN4fqlo5rwKT9r3cTyROGNfUwNepk3/+/vWvE2mkiFiNc3iAvpmht4rFdAKDxlu1i0irR4S4gtbA
Y28izCONC9iPy+zcghByhiBcBgDCQb7csBv1LQas7TNGVzcbVcSQi3cWVJft8TXX+dlw+ny+Hnz1
YaPa7FNrK4K7208pztNHP4wCu9JbvMTyAyzH8nk3+gVIIE8ZxgfFSMOlive34x/hdEChW2PawzRW
3ngYxSivPhWjZosfBWxa5UHb8YFKeF0ABLS+u47YQwNUCt6iLjR1QCWGJ2Eq3rVGMZLjmLPTPUmP
yRdv5jCoOGWMesRq0YNbgOeN4vtS+xyGgU7Zl4DISWR+Mk4BCtXmEWSP0W+Y2cwsxrS9l7ClPDXe
1Rj7I/J10M+Lvwa6MFlmz9lFi6wh10ta8BlqypUHRziHYnjBCPbWWvpqazl80cZQSy8A+0o20N6n
mS6tX3LaFQC1RE89m1vF1WRm6xY4la+MdIEeaVrl68HrRyxbiMC+gktG7iqpBnyOzBb1ZqbWPeyz
oSql17oo50srOF/f1dpTJmWokSPsP0iHBv+qUFuPIPCkWyqzyO4IlfrvQS7UachKbDGGMy7sUCgP
91KLREcYDrCILAL+xBv9/j8QqrK+JLrm4Rvj15YNmuinHgxBw+qS81qhNCNPW/OpWabVZuDNzBsX
OMTnHdGT9O8uiDRTXzbYhemCCpUWMAAeCK7vTn49BmnUIXzDDgMOeSi3FMcZLFBLc8Zk7GXNcUjl
rjqLEYUKPkfeU7nyc6YuioH5AijSkSjzFB2tXjALyTJ1lEdf1nGmtRSDLQ2pFlqgwmy13wgMcFYx
Zj1UNcjsxsSg1RTBLz13IaNTJ+jD02lNJC52KhMfyuDl55SDMWJ1sv9ZndOdXn7gU7RRRYUCJyg5
qiUZb6+kpGUklzyiAkImCiJ4AtPENZyZaVT9LVrSNUxnWN+KEmj2Y2aZ4KejzVnWRAqwymZhcNlV
WCfLw9jAlhx4b3IrLp0v2Wj1h0TGJQYd67ahM22AXmNtDcrGttn1G6IxPFiQ/00c3sfjwKtHZGtN
mqcb6E1XoWJ0tYceQAcVMdqKqoDpdFQjeAL3k0ycVAEWuWBQQSj3LFWO7kJ5tbwzDpBoSm2bHXtJ
45aWTv6ksIJOTHbZ4jBP00TH6KhfEZ+oLwDFoXDEjdIsdG+ma58hlx0r4hfMEUOska6TocEkMMWP
lZV9NdzDuFhdVXdTlrdMt9rDwgED6v7XhtvWo5AXIAva1MMBoY7i9p+RTRoZEcl8Oi8wzwQlOhU6
yaR5kVzzPuYlHryLBDFvEKWDed5N0WEtSZUPFwRtvSN0cISx9LVfnlWAyezUs2axnl8ZIhtSsMV7
q1A8+Td13e4uQtfBn5jGiNPuVcYJ0wuhydXh53YCzJjlKR4ujPMfSuWyp6wxeJOBNoznPWhFgZM2
6zjk9ufU8z5VNVgUWgPOiEEL65FJhfOmVwi1NaUuJmm1iYayAUsL53UlaxcvWlcVUjIl+0ykosws
BbWuL7Y/Bg1kbYfzMBkS4aa35BdJYkhTIyQcZAWsVKZQUSGMK4wefeb4zkJ1FLknEHjDRnXMbB/z
/2DjcxupjhSfCNaeveVuWBXA+MHIpSB/G0JPYRspbfELiOZhbHmkQeGLKxZADunQF+vXSxrU0jwh
TYG4fCcxye4KR5IZQqEaGO8XdlbWQaa8Ai+Py03QMhMfUzJL+tlufgz8oxapaoqCCOMRki13cN1v
Yw/5akfrvSX6N6oVMBYasEC0KSsFCCCJcx68rYqaLqwNKIIlzSQzEFdaby0s/xUUE8lrxcmvbYxi
XbNM5xZ7Q7e0kOTWUH2Qz7sFdZ5p+WRPWBd4uyv/0bsciP5WUThIsrxwISFrEZGb6rbgGqjIQWBs
oo674aeZMy6LWKqvZUCvvQ7i0jxwIac118lHSfM8rlYmEIwzGEqSI/qaURQk3khHMA6FRkxsFOEo
A++nI0qBgs1W7jdhBPE8fhhvBSMp9sGhWmyG6+G0CMZZnywd/yAy7pL9uEW88R2E7tpPBVR7bST1
7eI9XbGEd8wTuhOZMU9TYt21iukS0WAhsmnwCaRzCIZFbrcBzZEzBTgqZ62eNRMS2u2fU5qZ77xc
x5whp9P0WpJjXSgzZ8uxMthd+CdXr94VV0Sslc7U32THaJ5leocGlvcnQvJKCIhKDHA+XYgrk72/
AUtWPMmND6ihRw06XJ3jpCMO1nlnMT6hI+ycTTBg81WckqYfE6wyMTPF9Ksfw9r4ORjNu83BNHev
bEmdWJ2LUxL9hi3KTCtbe3167DSLHsnXfaUOi0CCnLa7uPGMEoz4eHGydu8FLpC+r7GiT7yRG6Qt
hGnRPpzEikSPsd6nWP2ZIdjkjg8w59XFWNiG2JGsHFNQaPcMUg06ZywAFuaz0KWmQ9ebXu0nb6OL
3qXuA8ZYFkUPKaFrAcL4Z7r7SR40oxxlWMDojGAIjH3UJqHL3Jf6AopauGD2Wy7S7onQ2eqKX5fv
2yYGlPDNUijIIZ85p9S9skHJrqSz/wv5P9s9yAGY8drsKY/uaYZECTBJRb6oeMlIOwpWCzyLY11a
120pxNDkYCM/mynJ7R/sWVtwDLBeLQqNUpmSErbktIb6Esdgta401gp1u7NZ6xE52RUTtTs4JM2f
dcKymdHviHuLhN0urMqkA1LLtnMdRWEL1hA82uwYsAp4dBMk78jboMeNV+zKoL/tCUD7G+t8pcnU
XrwPP2HHOyIxCd7FnWrA7OAxvQHXzSvmGnwmeJAGaz9WUk88zetUMuGslhqGRRzMq1xESApxlNx8
qU9FMJhXUgjxHnTLgML5uB3qlr7NolAtL3BQ5jggV5N7kK9vjAsKvEsWkPN0Y8rNIoKpLI6D9cVU
guwAaBPHt6pZednxYkRSbKkObCfWcSF2b6oH9nV7XmuYfi1of4gKDU2/lJORrtT8vQosQn2Eg/6o
KV1CRGEm/PTsT6jMdvLFG39Mx8nlWNkKlt3gGTL9CL/GdoqRbKEeI/b3MfDvivgrHJN721B2tth8
Zek38Z4A/Rcbx2BepM2eab7sI51SUs+WzsebDWCzHNXIdrGytvfFLGsd/VLNdD4BQHQuCyHgtc2i
mS9piaujDpT1CPXeF/dihfFNaEra9gG95gbnQaBoZPgnI7N6CKqdyuhNCyqcUQl5kHzFW9bz8c0J
Zr5Rr4PX72AiqryOU2wyuWuijOp3Q7QT/PWNyVu+MpjYVs9ZXx0b1vO3itBjY02NYAXUrNLT/nbN
T2O9ZPi6sNwaGjDheehwy+A8B6WCQd3efjR6Bu7fKgoH6jfrXv54oRA5aaD+zsa9GB7V2T/XBjVa
3axPrNyqZGuW59T60J6WnLcLF/+ZaFb/VVL21t29R/yPG1xvc2VS+JXdUDOTRkBfNFyNuyitC/uR
IRDYz0y/zAktWeHRknuC7jdx6RBXNP9pIilraARtiEgKpoGkaJYJHFUuFCOtll6pUJ2qSWw24GWm
RIPy7dTh3b8jucFJE3uVGuJz8cnW98E7sM3RHpKtj8VOKyN3hbHcDtmDvoIAdx7FOYQASQEHTRTd
GzmoundVIRhmYAHOEcHs8rfs6pb9Z18LdzA6QBBMkeAOMegdjuZyr9hA1zNwWQDvdGTx7smJbMuN
aTnEDQOamvH3lQB2GE+R79FpVyyy314fmhTVL86iIp/tjK+xJ1loJQdMtBrrGRLZ01LTsoG+hw/8
62aQ3aZBFCJgWK3BhOYFz7m3+0a3MCuAXQX9VQcCdzeAQYF6ucReQJisarpRSWJOrxvQIB8C1pC9
U4siVp1Hs7Par+UXHEnXm65wdFy1TxDdksLyWPQm1/wvrwByzchn7iWAVWgvMdmmyuPxuZm88+a/
dc6JhY4yqsEtI89gD9ugbeLop9Tb4F1Da75JUFb7fBfuGxDiiTpJJjczV6fzJ64x6qhH2Chm7BNQ
YDcO9DTVpKLFD7Il6OFSjVzwHPEBIApBChuwiAO82gEc/GEpVGqdLjvTXsYI/BmF7LqtUk6HrXa4
F8Of2BhxI74q/RjNRG6fS8dMVIDrMbOxBO6tpUk4f132DWymOcFTWojHVbgatUfL5DyPZZMur2+G
dAGxawBDMxed/jzAMk1QafZ9ImLciJEZk8ppG4GF7BhQpA1NLH8gBdDP282GCYXhEiTJOlng9eIu
o+UH0pTHTcOEZVMAVRPWe0NfsrPN2Sq/sJTtW8HwkdZi62lYcJVDAMI0kIdH10JRhQf9I4oxkjKF
5Y4sfK9nXJSm4cZUVgz1pHXnEqBYzEO/rBAUio75IKlxoX3b4C0juUOSr24rQV9Kogmpl7TUdwmc
MfXPmnpF4NIBA1LecrGpysWbpRvFBFRf0b4n220XCcseUmAcDQqTaealnUmcURvAq0mzz1iz3S+J
Rz4zE1dZauajblFO7tzHHlre9WiSGrDztqk09gxo52YX4ojtMZ6GKKvAVF/UvG9VOUoY4wAFRtZl
8snGTandH7VSSVWVKIaK6agMfnHSWmxVp/E+jOQWZ7YZ5DAaqlgJFi112XRkRQUIznVjrlK1GfF/
6KEhYcVoN3xTuhQIRqZNLIs2DTcrvhrza9xqDUlzg9NN88KMjG/t5+JfmIV4zKjoUHBXkwtGxrA5
iBPmukn36LOX1oSM8Ta2HQwNl35zK0jPnADkuOrDAsPPeWReFwyOuQFrIqG/+spC9AEqitEfIVMD
jffo0qOakdLP4Gy9qLChh2lZmG8MgZtXf7zjYMd5lVG/koVc17b35gdwcBFKL1NQ/iPzcgk1Ir8S
wXKSWJOMQDQGG4kCJsb/Z/nO4cjxZdSc1Keu+Z+cQGXJhp29aGETY9XtNQXdBxGPW+pMPaMIggwg
rdiU0zxk+bAUx5JGsUd8y3+uzYuire4r5GskZ2F33NfVfTDGzDC1lK1NF5uqePso6Nm7lC5W9KIP
1gQcDbPi5QXaLEh9vJ29ji6su5SoxSyQSGeSz9DM9tY4XAeQvViz/zx74NPaYWalNU3P0l6T8iNN
MCYAu5HFWcOSb07/+EqA7XaUveETWeOKqLcLWxtp2a7UeFRWtaEMY+jJhs5wYhYrgKYH+bu4+Xpa
BQDUbr7z+L9iunhT822Su41JPuxHxZ7W2Wtk8k0gRUa2lLN6wYJjGSnXhPqQRpK2pA2ItGtlcIM8
9ZSplJm6ne6ifmXd99R3sawJWPC7dm48eEPHRr8j/X2i+Z4TfXnQXHigo4E4A8VSBZq2gKcJiEgo
NcCaGKXGrBEmuyQvKq58a7DAhaf4T/VdzeO7CfIpqJJKmVJf16Wkzmd6N145e7v8OjxnvxGSkEM2
kaEm8CqVzzuhFlU78j+7UazaV5lQrwRinaFBXGQ7Uovkx08dqzyErWFqGgfbc7DLChtUYczXxXnQ
AmVGBHHKfheZIr3AwTwmURgYh7iCU9rXRFSsK9ub8bhrzVfRrSAwfchVaizDGLKxicu6iDVMNah9
0qTLimfriJamLBAgyxWCVb+SozOjz7VAq+n6sJlvh+Oh6reixKagD0LXdJqi3oRNUhLtdmSH42mM
N554rvTVRMDQ3GQwJmW/L1qViKjLcMTDITCI993v+powk2DGbBbi2OFisNnR9MtnHVR9FNYjDRlY
tpSTm3kf+2tBGfMAjQHfA7dnw33HitoN/Ph8wz8ivrhSLYsAoyf3oBU+jM4z0JC5K0keuUhUFU4H
JSCU9padIwyWmvlNmGcZvhfPnsaqiQgv+eYtKs5M4otWMnZGMqH5v0eeoCIjOoL8CZf7SbyXQ36b
bTDMnkEVmT3hqhtV5e8gJrYRWP8R8bPwPYH/19KdCBi0gt/XrbRy4lJCT+G1Z4LVl6tusfET6IqC
SELmM4CnwC5inzdrVO/Rnr7sNpkFzfzdxrPzEuqwpmFmCUCgn4/yE70aYDx1AYyk3rF8GziTL467
7pjDb/J4mwLdPZXZG2e3dd11+sC98nUYIaj5BpL+lFR5ZGycPYTlUWq78ohD7D3HxexZ0qk7rJWd
ylgvSmxIHwCjG/kIEbE06nVTJt+MObujWHbDUbg9mjaoLcsIdMBCRG3MbfGwQ7JmubcPJfNpYXoc
bz1l/Qr+AYqR+VwchdmfO+CYMAX5SBwUV8+3zZapkkQKPOa9IefdindUNt/N8bG6znXvJ6m4eF9a
afTa2rUkFj88zgdQEkidFMclPPOB+Y6rO9ZHc1VMWEayuqJBOIemrOPniMcHTTHqO8ahfFWQwO1N
4zGCkPdWrYpPaRn23hQ6cJhnJY9SAzlIQlW7HYlTX1nbj7hSB+qXTYjXl7XBT2Su52oikEu4HtDV
BV7znz/kipa9lwfyZDQfTL5fkNeIDqwz2mLpLra6TYf868dLA8wqhNu2ro9TWi5TXWjJGyIDLCYh
0WT2juqV6xEEg0KprpHiiqROwW9BSXn/TCzIa1mYdcXIZbYl714tNcww/Q30G0QkayWOglyohv95
Mj3JiUdiN91ahhanIq2wTt6PXV/3maNFTJdv9+mP6Vei0LJOzHgxY1+GfSpA9+B7q9yWfv9Blszv
1cTIvFv7hI+fKBss9aPaIfdqAtN3ZkUSWgXTKsPFWc+P4CbOAwsyNCXJudyNyZ6+T/+5pbi2vRzC
4TmyFfKkIL38qqibKXwIauMVBKGxqLU9gzSG/c8Z6y4tlQhIL7efv7m7g0eIx081orNBu5Yi34u3
BZ3nFk9+tk5OSYXbDmxh4tUjloe9z1e1ZCSQhv7+NMCCwRdZzU8dLQfZs+CZ57PdKx6ah8ssWStI
jss2xt1AMpI5fEr0wVenT9eQD5HpWkqtzmdyEOP7r1Y2zPQSq+3diTCN+Y19/WDl6SfMUhyX2nbV
EKTwKAz1/h8GylG1o8ZOo+j0X8PBcjRlbggrUfgsXe1urWshIiGldaoYMrQKneB2VUqK5MI1nVlg
EhuKvZksQ7r9565AtuC1f4Ffn46a/I/JMm0Bl9jorhCM3pbBak6qF38zPHkd2kVoqaMd8EBqdQtc
7CoC1KMJlEAF5dcfysISDpYGlKimgqz3yDssM5yU/PxRMoyZni/DNDABWAsP+JeYFydd/EZ6cua/
Z2TF3nZeJjMgVU8xWAqNV6fw3rLUy9J1onjiJMTQh5jF8xstwZwU04Z2iqFP0ELsM5SL8W0ma/YU
2VLEm6yd6FMcIwJJx2DFSOZfvNWLclIJ4o8gSp7MdBgDsOi0r8cm0zAUn6QmSMPhqDEkbc6qgh+j
mr43GODsOk9Yj0WKgMKvFhV93WEPcWtF+o3lF8DhV3avCxNMkSGYVawAgMhmfL9KrlBA0tS/FV/i
Q9raW3QpiQroSAHuEXbOOOrKx/cMKkdP/4rbgsAAeJe4p/FattPY93CNMhla1EblLr8O/1HSrGhW
zsTUFpZWWRzcWqQlsiGc2woGfp9jrsXfFlJeUzSFO5f5FOBD15V1r2Ct1nVtE1M9vu4FGbnnok2J
nwY978k4tTZZLnFZT/yK93wbOEZygZH6zG0qS65OhmANXr20a/0uXWSYOyLGIM/Q4xf51wwkYSSw
EFef135Vx604HBJRWEpdle5qmM12vUgRX9jb/PeuK/bPn90UlAwJmo/2BPutu8jEeNKn7U7urBT5
TQ19M8iErXRS991ZGQbH5ZT7OFVq/alL4rVCLosteWH4kQEQ1MjcrumEQ6cYmBJ0mFvx/BeedJP6
edN89//rk48cH2g9pEJA+seF99ItjsIc+ZqN/xn+RfWyuCW6WqOKFLm/EMCBgaTdQaPiNjdqj1AB
pM6zncFNxIFAkB9Gz0MJ4tNkUFrXRve3HL38Q8b8h6YcNWUstRx1BVU6RQcA0bhe1djIys3iPvO1
KwrwREJyCMBx6lXzN5xJcQdoU4yId9BOXfkgnxqPE2i4yu8lgKu2ERAqfGCpurbb7PzolSek+tzF
oW5aFe/iIbxntMSEiDEB+i0b5jcRUahuVT8ThKsWQplHKFSZ6A+Gt7L29Ld1IhX5zbYFugtsCT5J
lblXujs4dCL6Zi8CKl7Kq53o8m8le2jkXzS2W8v7E2taT7OihU3/wMAthvEu+5p4ifcChQ7V2iJg
o3yr4oFpnyCXCHOtptOFsxJB/D1tsVdzCul0Q7vQqaz1xtv2k+fOFbz3jqSTqbfqsbaKMaHwZiEp
bFt96i2SQ/GdyVloYIXM/+7rFODjCC0sIciYNhjgvd1UGSI7oAKkWQfLwPBMRWvxkElrIhHdtewZ
zl/rpsqmz+fwtNepSbi0+8neuoqGbLjgE2yvJv0vmgvEA9PyMcO26MLKanH3kU2iC/Z1wmbNRZW+
Hh3fsbJdbRYGcIOxyx+u6mEHF/jVbuFIof/n9i+YkyqQh85rF4+ze2nLzzHJZv49JxM1pZpxN+k8
OTJfFohQYm1q7A0Cn3mHnGSUsuVhhWzurGD5uPhT4Gpfj+DOKWhLqTDI9DRGXK5ipgt4TNOJywCr
hBvOeMhCsP/n5rYasKrQ9CH2h8vtRK7IF7OknfOq7MmK6BV2IgkU7qrTCjius8E1WswSg+Dz3wwn
ura8Dree4Je3Oyt8urS/ngponTycU6jMId2B7GKm8ed5TB1JS5ob+5agyIieWHflZ7A4vYx29GcS
Hgin/Qc03zr+7CiBdgQDkcJPXekcrnmqHUZa6Oosi3DoyzsEVB6msJTvTObaoNHN6Y1c071CRwYt
iEsnslKoMZw1kLuzlvRvETnVb0fJ6KfUVSRQIltuxMfIiJ/2LsOnbSWqmEj0hJa1/ix9WhP4Tfi9
EoO5QRD1x85c4ef7Jk8oGwiRQScNaR4Wjeg0h6D76Zhuz90Y5JHaG3I+uamHffBUPqANz59Uy9mg
OeSklQ1alLmuj9iDzfIwumxscUmDgoLontWJS9L73N+LJrf6zmzdmcv5dYKOWNC3xZdp45oY2Rgv
QfVZpJLbK6SGB/8JvNvQZ/An8eRcTBaWEmKWG7lr3aqum+f6SCAWKJbmc1iy7nbJOI9S6uzfFao+
Tb52ndZqVICQHdywN424hpYqdoQCGGyGLLljEN9Xx67F8e5YhtyS3WbZ69oxM2kOeHjUXju4JNy4
2NxBKgpiVoye0+e5un6tuLoKiLOzoqCKh/n3eG+5Li7kOBiEpNhXIBhkm7zTOQCQF0jYBN/G5oWJ
Wxwi/oD/dRvgUhEodzCCQcsIqGLeqMV7hwmBkTk1Fnzj1RK9hZ0VUnhs72V43ciTjTFpt7trPX6z
KcWHvlqWfYCx3sKzzdOHgePP1wSJfsT9Hr7FPs5UB73F4JKyZ4B4BxIPfhxfnHC2Kraa1RmEyrX7
FKRn3xVyamA91qkhljN7H6OM4hdcQzMIIzLsDr2kfiVU63cNDRrTqvNRzUurdV/rgtCC11CyTXvM
Fjzd7HtcUxxVTE40os4xE8WylEfhU9QXpgvnK6trchEBiZrPMXlq/rJ3/jw4YzBHmdKi9O/+eWkP
WFIBVVi4NFFC+KEu2VgaJMbYE1S2t7K84pcERBwRmqBoUTyBnMW5uZtr7JI3f4wen1Flj8/Fr19Q
JJYiUNW9va6Ldb19QLk9Hco8lQzCrKhrcis9Q049BTJx4or/QKi+Uq7jVoi0iLYjaQHdQOYxpa0Z
Vf1fY/wez0wqPI7TghdkptGbpzeeWYlu10Op+YDiITzhCThjbkioQerUbVx1OuTqyex4QqAe3VDW
fnIrnGp8koXYRgNGFcL/X9ST2xSc0ay6YZMKPgBWLxroxFKDoYvJzdL6NwYx9A2xniJrMyxTePjK
ycYn/DpyLseBZnFb1hp/6HpKmCJtdEm5nYTuYtktuJSfejav/N89QUJO3yaqftMPfA4tQhT0rAKG
3a8MBmKck4xQOEX6B2freeKeYbPFG5qJ9d2rgNZ5QgOQC//gekhqv7IYdGC8NHNq85L004BY1cKp
Z1ojDWU71BV+eOlYbbXCd4zpmdaq6QD1h00SYKb3E33NOu045yFMTGHL0DY1h+0KOTyGspQQnTEU
Wadp1XxtLyYcV5gqsKGG71ADzTJMY+FxAqE/gCS0Epllfj0YUnbclsv2qfCxWGcF40tqxnMYBGq5
8PzeNsdxdc9Inrj92VCqjg38UxmD6lBH9upxoU242TZLhnXhc7Ey3J33jGcrDM2Hbp5kpbfUPI2J
LLxK39Lq8zmDq+f/Pp4g5btcLJYjAhcviZXMKGJP6BfYOVwmQYHuYu+6tz5A5zgkJPsVlL4MGv/V
l9pAp70Q+G67gKTLoLrywjjqq2xqKuwEQJVoAK7u9Eb/Gy6FTd6AUOiaNHyCEyFBfq6U5YykOvWa
NNkACIunMR+pFzoM++OyJCZbcEhJnAOz+H7TjLoSiC58TVi6AZaUVmB7XBRu4MqjtOmTkdqI6m0F
6HfBNo2N2hkFpn92IO5tq3wvknhjUBDPxuqXjvc3sKUIG1LdpLU1IgDvwI4xpryUCR47kjSVTycH
3NfotLTSZjJGqrnRG3WuTimRvUi6An49yKvObTz55VqGIOu2BTWuezEnjV60Q7PS+ujoFa6Amp0s
nLXh2mj1bSiRQsOCO9IUVK1Y04S7ky8cXSP1JAy88yRejbvTCmFACyzRFS4908/iZZzuSp6dst6K
5UG70vGPJDJDkmayktc9wVEKW6AQ7mQSceLu0Z8OrEbTfVyTdhGhzB5nOl31kMLvN69k3eAxdw5W
w0rNeqAWY8pogcMITsQ5ftzTNQW5Nofc20ZKtBdwVKXVvtGtv+tAntNkHAU5113BmxBCNfszcxGc
G6SA0sSbeXh++2CKxu0qUCfpd6Qr/vsrP1z9gLFoaPqWwvHk/NTeuixGCnBz1Id/Njge6p8f3lk5
YHhAcpGgZ3GEp5moL5waXDzT5TlI9ACe/by6Ehfx4riqP90Vk8JTmv1rASh87c00j7tsuZw6/jA7
xQoDFa5IR57rX2Ypc9rtthGEL7EyZ1lY5FjVuqUdo17fdgTVvMHjBcul4GV4cwP/kc6djDFJYW7B
slqJAGn3JoKLyn4r4ZeyBF8oCiC01o/eew7QUdfNOtgjqJ63Tr0Sre4LZCdZrUVrzGZ0qBrYRRGV
BYhgIsmLOIpx1JlF1jgcZLUKxbTbySZM/2LkKtG6+nCPGdZEy6kzwzOjUp8hPmKKNnbpt1+i/YLh
D5JeaVNVUlvTZiMxaq8Y5g97S3oWBSrG9+n5gQUQk4dJ3h0YIZ4qrc27enVERXwmSp9DGV0yH+qy
8Q2LiOuor9iycE6lgN0CbjpCxdQYczlpVZprIakrO+u4liBYIsPNis/PJUFewJhdZ/P+aMW4t/lX
qU/dlfGUBj/zOGBszmREo4Uf4b1xmH2Us0zadpPe8k++vdnrxuWM5LKNxAdSpLRgWqrzgl30tpDB
XWL8PQfKqrSS1jC0JELZUt3dzjQe8cHE9BaJFvRBqUDQJi76TXTWF/VhrmCMaPWZeJ3cbGtlH3PS
8w8MsKy6CpsOXAwTWtrmEuOX4+KAV7W7rjy9RdhhtNT6PhOky0IaKFS0vSzcCDH/N2jFr+K35epA
ymxpwopZRr6tdJtU3j8JOdHGCxj0PzMWH572ifx9xLDGL2ahWdRR40lX1S/cg8PQDDzFPfJHoBFq
vLvXc86ECpf1bmrSjNCyqq8QHyXBVEs4mPKE8d34GEKRWJHdy8LjnNnGhaJXat+hbVwol6zm6Cev
qIG8Ow+l93JiE5T2G6VB0Ei/1FnHlJgIQcS6vUo5eQSy0PmIYLh3sfO6BLAP5EyCvK6hAas6Uw9j
OWDvc04HMev1FNgw73D11HGPKuimnTGhyRmczq/qhMuoJD80DOSxnSsKED0zK1nJ7PIes6mojFUm
Kj4Qw81Rn3fMFp99pg3EHvfhLmwYYYs5JjHWSEZUeJnHWSeAKlfVnv3gLB8/dZfe06rR0Mf0ATBa
Eya54nmrLM9tLSPgQKmwTjPuvSL9B2Axu89c6fAo6yTIqT42WpLO7r8PgpAUQehlCtsqAzkRSPRF
fgnO3BlNwo7Iu+IlQhB3LOXtd7UBK4vNzXme7JnJbyQ+M8Qrio8YMZBqujlxwSEv3XRicONvu1nr
k/2tiU/QEUoQMHs5Vs0ISFpn6Mt2H8OUgPtM6hlRvHICxvTdPLdo9lazDAaX3Anu6hiBe1hpcXoJ
3zCLjm8K8uqPHDpgIhu2554xKNNYWJ31fojP/wSoTdF0nBlJbEH74rN+HFOeZ0r9h/APFz78jJee
8iJT30uj28PFdNwYFbuHcc2fByRzAZH62qRzKse/SEx0kJ5H44CkLksDFH0PJ9rXmjS0YrpkIDcq
0Fgp2M/4bTt1vtAWaxP2d2xVq8ekEWy1/uWVb7oP8QTHQPwTPOuFZzoXhkxkxPqW5drUq3Z4dJRq
jU+kiO360cULVkLCXq51UxHPQIIozzfQNKEC6pKmfsJ44GPXnhJlZNYmte1l3DHCu+hMG1JmHN5m
yi+EAffIn6hKEsxSsw6ziCBI5/IcY4dJWDVjrwV0KwnBGTmmqh4//Jv428wqWIompi68K+9iprRg
yDucArUoJN8J5eMP9gzeEM83quHBWGTd+ZpLCnDn8cPmiXNIABWFkApj4r7KgGImsUNflIiw+8mH
CssMA4dhcVZVSt9BZY9jtoNl5jppQI3HS9TuFv9rLNYNBNNR1HqJhicZCPm+0JMb2iWNv5BP1xY4
3rbPDXGX3RBlHs+k/yLhLgPmRhE52hW5eiEQEG4M3+2UL2f+Ea1AyWSusTe4sbvq/WIW3f46iEAL
8lkx65Gx74qCJ8y9EQzOX9mWjqvW0GSkgdTeurXnUlWvwJP1257GmhgEEDaY8oV9AlNtYzEYTxYA
mUma9LFtH76OOddsZokJtniTkTNYWBCuV55YV2HgBMMjjdbAvhdZyMR9apgqEEC5/N4aw7v32Qn2
fiKm0EhG96jM4hEVn0ExmxaHCCw14pKgA3mSSXC41PSsY/oM5SSKDIxa5pQzAQ1K9OnloIiFHQpL
/8QRa5PGL+t7Shai7YCow5ZJLDcXSf55RO388D5u9A9bhQaaifW7QvrKnxMMYaJTTDkB7f/dqL5g
JcLjaFlso4iydlHiSKOlfYUXzLBAqVnUEsItH+hOv0eOvLDmQW1howncp/DODTQseLfSAk03dKfx
xeBzKIey3anjywyFHVosU5na+9GrbHcsWjMZSlt6H7h6t97llJ96pjDRPEW9QiMALfvA8g01gLYb
ZQhMvG19JZ1dZWk89x+ykT8vmyW7jXNNZMI6sof6DbKb676qBK/hLYl/aZStC4u4mNeKMrJU9I07
WxbhtwWmprMomVwqQ0YoMFE4CdBRT/icXqiigx37BeXy1q7GQWnX4txCTgrrHYMQmVKytOuR20lt
k+UyIeb4dZVQtTkGNb+yj8t2YmIZWejTQ2AQ+EH4hbvUqMc7zhtWZZNL4Lw6+FxDgwqfBAkNQf+g
0G0yWVZeZ49z6y6JjMLe1NwrZQ75S+gZB0xWI5s525SFH2aFkmR5tOM7LdelNUm6Cl5gCJ7sEICo
ZGGuF72CM6jOnbW0E4bhWCvjk7TgfHxcj6s9V9J1BxxH9Wssn7+0dHtoIxRmNkXfYjP+Hc2OHxgq
GxEZFZkjrdQkh3wzmE4ElK7MyXtf7IskpWaeKSrA/o+TVjyDlvFhug8JPWggn7+bod8RPmXzJbaD
184V1+T/19rsWThuO1bf9fTdCv13O4L3HvJJ1zw5zPe6wpqnzoHZ4tzr/23KM8FLOwyjB6n4+xay
hLkYTBw1BlxwVTaS6WIb0sJurRt8/To6lUvys1nR6Ztg9SwRAhRc6Fpl6ofzX6BeCdcnNERS/MgV
EHdfxKp7FZ8wx/7i35zMBoE0QwrbC9AUWGxT87PTPER1cSzzHJP6Xb361tPpZMzGhgeQxSZT1LsR
KtGC/Swhz/e0I45QUqg8wo5Ia53tZeuryns5kxEPpe60LwOGqNDrhQvLvFheSdGsq0L4+4FfoifM
m33c6WzlaNN+7iEr2Y2Y3N3oOT1RpIj+frR/ssqSjLLH955Hy0s8/eoEpc4AB0cOpVSWXrkNs/5C
AalxkViiN1raoZnsuWX6jFA5K6/9oWcvgJZyrCq2tcYof2GWcar1/rz3yG0XbHkFAa/tA+gU9bzJ
oX6m0gF1sIYIQciPp8U1ZPQdEwaeEYLrg8b2A6tzYgz3TOffRluCvGvmhWBP//CCpmMJcaPneA6W
fkuf2kJROf2Xte6NIsA3bqKItcCZrVfKThl/cROzreDwsRf0q0SUMwaIpaipoDKTHegnzsaJi6ij
P4Ui0ELiqYivu03DlvEilTfnCRO7zB21dFekGj5TRtBUBVJQOyYlXXKvbwqbTdqBMCvQr4BByOYa
1FOLBxu/i5NWkCaOY4KT80EcVTeswM1eGFE9+fw9r8FR9w09RLi70YaqXbP4W5vZ1b2p/z/DsZC1
KO/xeLiSVAVVJd1+Suija+QmapUwvQFQIkSICzVrcBlf769TLDXGRuUne90NKWVMUteZlDHwCfFe
ThD9tWFtk/XO2wdmP4/hiNKAWM3IlW/4bWKnLGSZQ8jUbkhc6pBpEoTFx3iJH+XbyJxq4G7XPzf+
B+sVXkVPK5H9KHcZg87slCu9qmt1LOB5S21q0Uu/LTZnELOZOJ1QZhCT/ftKcV/V7kiFtnXc9giz
WqkTC4F9T82CBlvycegZoYUE7VBkhJIGzaovx/eLKJPT7ssQUSI54NMf3Yr7CqfsWcdmDBPwObWJ
jtPou0UHIZv/gL/0G2OF66W8Cl3dDNTGmaK3lUSaDXvzAHF4Kqc7TezQOFrH97bJ6NitpuVTSGYb
Yw2flI0Wt8A2mBmVe8LvKJwoZ7Cvui5MsFwDJPhDczDg9MLf6tVFVv5nSBJq1uWVZ/pT7v9t5SJz
RXadGcAS9j4EJUVX3btDCUKu8mp20ULuBZhxeGLcFDEORdfTgpP0Cq8noMhpGUN9A6uNmREPaq3c
7kHllD9OgVkVZl+SJ0ittvfl9CM+9sXHOa7opxyVJcexvgp1KJZrPJMoPjYC4KRLVHZZj6nxH3gv
FtuBmJR/cgfYqOz7/ZZBM4qKEiAf4JHw6ZR26Quoy2V8LIEFrjmGTaN9dp/O5W/HnaYH39fqzVIQ
96CwPF0fYyTxeyOlOav++LcAKnR4U+SxNuVsFZ9N08Cq2gupbDmO6CrkG+UPa2vF2CP4vK6jhAfB
wVlxTkEgEjqKZ2i+9d0d3HtUeSlj0W72v1/BJHiVC1n+yFgJi9I7Sz702awnTomsAwP46OAeivc6
z6POg6ooIyzuYB8VATozR5nDSf3AQhwh0DrxQhUiJe1dwg87eF4rshjTHfU4/4ldmyBKFBqIQtlo
H1xSvPXBtBacmwGkWQ+PfUkWMIXXqlzhE4Y9mRdWPaqWXEUP27dTmlTgtl1GQtNVoszq0yGnS9HX
eyVo7Oy3r16S/9vWY7TPz59teKLwwuamBqZhNwD6/dYfWFuHHkCDyd591/Y+1zf9VyzXNEcURpKl
NocXRNmkWWM8YayQlL77SkPoJHrF83vBRzjteqrFzCi+o1hNf+X8KMF2enB36NWMymOMmjDYR4ed
2HK7logO8SX1GsXTu8AUl/XLgdxjA/ne8ym8tBz5u03Ake7zcbNpn5OnF6TCSATMJlwmA4aq520g
nLejAuINxNsYrnEZP3OoHdiEOJboi8GISkcadAsbCEZJEdortXMDKC/rlYirpqVo9o5tB6C97BF/
k9GC97MI9CmXVaZ0laRHuo+jYQhhK/jJFUHsZyQpeGhmW7+huk3O6cBQpYMm2uoN6m7ygoQ0p/6U
h6kTTzxh0Rlka+IyqigtZkvx3INGf5Gcd4frBFkH4WlhE1MsCzVg9wTdPh8oJHZ0loGViLYDtVSE
DFRUZb9Ya8BAD+C6xaFrbU0YIJlyn4pa5Wodmv6bEvgDHqywhz2/S0EQEm1gfWuBh9syIl3edMgk
p0bWrf6QKPALAIn/Ctu3lk4+WiOwqaEMnLXIoFqU/cu8/rYlmuaWW09FOOmf/IlChmeFwbnhglTD
Ad/7PvY2HoxAUGZ2P6TWCNjKPrb7/3bLkYcOLi2zdnpjdGl1wTsvZFbpq01QbVs1wIPnCTDv0npP
jYcsDJj7lhvJV9FFkByZhsqUZMcPTssUuzTDF4o65dQ56DyulLwDt8Y9EerncUYgXDecSYkK8is9
uqTJUapTlt0RMlx5Kul4zg+UjE5Y7610IqcthKdfsz63rdWCXar7qScibwQvFhUNsRRx+7RSoo+8
xIuGwWCFD6OVFgTlYsadvNGQo+uoAnc3SC2hrepCI0OzMTYOs25XZ+2sq9AdN4W1e2PzTN6x1LwY
0kf+Tix6UNe5jZYBNxELJp+kx/3n+hMU06Wgs3rKpCro1XUw/iALx1ONmzCx3STGKP/hJokOSha+
qkP7uHasADEZ+7MdUju1HpcNqd9rQHmyPDKzCs4eScslg4Oo/dB8cnycBlCTc41IlqUGjE8M9eEK
ZfnFPUXByiyIeh7euz7ffia6aSMNM+ZVsE0V6c5JbhS2bAktn7ybvUadl72cCcOZttno+zpbSxJT
6pc6rwTQm4UuRH5SPdcDbCsdVFRjP7+Fai/QPP/Popunn7Gu3GdtYG/XLU4rAqPEdaScvviTDSQz
uHszGF8zVpkAEQRuyB3RDlIqG3DjROU36D/KyO4miYOTrPySMS7o3MgBFuVNRbUFgDcnBHo15NDm
u9nDY14e2+WcfFLypeHhs2RtUTJhi6lW9syYQ84oiJYoylxwj9iYXuHyZlSyk2mfSPcaOy9yYPu4
khZBzQFWymq9JH+hvF983dSy3/gXXQDG0DlTO4NmjdeOLd3yfhtF93TXlIut1X4clLHcLcnWMMSo
doLEc9dmCmSA3rfPpIjQwhgwEcqNXQ/RdLjnZ/LcbAI8uMSM89tDWn5nZ/pKoCqOYfjA5/G6sGpF
Qll4f/oaw7CuIPe4QaJ6Wp586rIpp6EYB2p1Fm5OWbRRwXrTopEIgzyuB750i7OuVEKliF+YX9/R
9biLgXXBkjYVRzcA74nfh/tVUtWbMe6Eyuq7B7eHVy3sncKK9RqPkL54wxazEtJzNcmulkFF2Tnj
Oopkpff8XRvlUnJ89py2OZ0j5lpTLjFw8VyVscTCKKhb/mFq+7iXTQzMXQr9Lihkbwe+adwS9EiO
PzqPikiShNqI6BRnR5f/G3fqM7xMaale49kV0yPSRxjqAx18e+rIHu4PFM7dr/M3nDt8r0aSwFu/
QDy5+r4uK1VunMTyWrmP0SZajEgCQ4UZut1uA9TurXPrk9Eg9KAxIJyuLs3JgdTnQKGOlRZxK4uy
yp3aiOM6C3/PE7QFZy00uloYRT1zGBNmFbQUjXhztnPtc5ooY9BwiMAhJZZ3LlomElUEyv/iuR8w
uaoknNzaJAaneMCQwTST0Xt9S0Ay/Ohi9ZyCu5Ih97nUhkdBu9+gFlOyGe4DarPwHUlYcAtXHtbQ
F96ETdK74lawVNUt9+icqUOMqdVVvuVtu+AS/4jp87qbp/o10s2tb2RlppS8vq/AyL5LcUxWOHtw
63qE6UmjAFs+nfhWU5wLFmg6ggOvP4SHKyAYvyw4gMTiNYzhoIEbkd7yOeZSmep3qahOp8WtRil4
9p8qKtJ25+1JjjVZUfpj/Mdm7hylXmePS74rNvkjxvHxEC7eCw9Vg58T4z883x/jUwolYbW4FZFZ
RsSnoZOdwNTLMagz8GcJvsNqC9/BwO06/S/+cxnwhDJ5XmmxAR/K7Z9CJumGg2AG3J5JeC5uyyfY
IAxVTXWsDPTG2psOLHwK/Yj9+xVxiQebhSj4sF20CzxPbDhPrW7SCxTI51/6Jla0hYuqPM2yfXFq
kAWiu+wDTox32y4BNSUjUfhqTBbewh41+EMNGWH+lqBWUUuHK+dMhlH7ckSyqvje95UBHzD7rwZb
FZJdpjUnrngNWh6a6D457K/EUhtN24CbKPpr/5AycFkpxUYpm4wC3VfZ0e4pe+rhnBnkFAIAhOcY
1174F9r00sXbYKB3fRoeB5k/G2v5tndiu/o2FgOlgvpW1kOh9nOFLAR3P8OT9BGmw9uJMSGjHFP8
U4Ttjggx0F34y1re5mBgEB7bk+mcpPgI7SZxda0L/1kc+FAVwKqBJyDImYB2sossJ5qn27R9simi
uO1UjO27+4xAZ6uyFKGDgNBJ1QCCBL/RhWe4vwbqJobhbFamKnidpfO6pL/0v7459GyfDk6sP2xj
0MTGK8BeMsT8ewdd8LcsSDJJCBHBl8e0egMLrFnFrYKCLUOz4KeNmHV6EuStyMheFSwmDkekwGIW
6PCtkVp0C2i7/DIT17619Uluqmr5I/IeAxwZAGosn2JJ06FG5jJpQ9Q39g/ulSwFBe5YYBGN4ITf
GVFVKHiW5mYnqik45K7c5lpj+CFxtvxBh7bcXnWDG1Ggyd+aTiSckLZ4gdMN4WFqSQJRFHtyfPq6
d2iQ+eaonLZQ3fSUmwGpQaXc00/C6iL/j8eFsAz8Ne0OzsbHmyYH1bEmJdt45li5iLXx49+oCtXu
JCwxVkwRLcCTnLPGF2UERWnC5w8PYEhpy6DB8J/CfdYGjaW937roeXgt5SuENikoCEzYloBTMIKD
n151JCklmv/Ed86LtEbzi8f5raFe/CSDn29wzxrPucAiRfZ+kj/hE3toaUXeu5FGGTG6RN9HFiCF
HLZhJQPeTBw3NDJ54i/OLxRtLJmTQNGvme9895BmsyCUqJG2M/CZm3ycc4yIYvtBY+5hEGfYKEML
RbtCzeJ/QS3usH41DKtgvp7cfF8PEOwEaxwSWTIHUu/Rpe2toZYUeAKb5kUT3jh4J3uy7MZm5W0D
N4rd/YdBc6ZEVqXySjgTQr/LMG3ReCy6bmVRTem0oCt6Z1Y7l2W4Uu3N3dLS3YXUPeowsKkqBV3C
2GMthr9yjSUqIuLwtBUu1jU3fkfDP5RwXtcpBZ50FEStLzfoJs2rBI3Xa906lAtgP9fmHYtmsyrd
SiHvZRsVfd6B8z4wArb4ICfS6b95x7O3MkMAi8dWDHEYad7LskOlg4JsbLtwzNS5F/xH88mp6y2E
IAhUjFIt2b+a0x/tu8eIQSkeBw7B8kigwfT8SyX6Eg6i7hMQ1OR/+KYTvQUV9jcpKQWW5UWwiGM7
XjJOT7GoFbwwQ0uCSOyBRAOzewJQcqebpJnsVC55YRuZ/ZuHuvebBwU+g5warCIyYPT/0ogEW484
X83kkQGoG1mQFOLuYexj7QcdTZrnlR4HhRA7J5AAzAo3IM75Ao1zjOf0XxSrJUKz4toDrVZyMuwN
fORoJ2GBugAspm0x5tI2+hXRDsvhFSL5FRbTJXJq1tBEukBmpKz1S24TlFXl+xruGROxk3PvLZY1
5P6zo7KzjCyf7sYJRHlRgU//4f8sDbD4KR256iXVD4NW6oEnYs2EJhAr/eMuCf9e+4Uk0nZVrALD
OszJyTmDMAmFkhUFW4wze8oGPrxaMn0RcTvJhznoNe4wRPVUJMPc+zIkR7PvfaRSVjpLNPr7aftA
3SzXQPF2tRylS288uf7GDYgW+FyQBiw+CAGe7ligLMCW6iOeIL3+cK5gX9l0P/Oye+goMWM64CqK
kQsBJ8zay0AeagUbXnYaP3Bvd/WUjrTqOOWkpQNrSuNg6yhXE6cnsCnhK43sdQFXEmLrrK0O6C2f
b8Rb4RumMsdSWzVNvaWYd1cfdDy2WQB/s6vdnNKh0R52LQ5hVZL7gkNmIONLU5A8gEpmvGYRD0sn
FcU1zShzftFQXnKpE9MzCBMCUCm0dm/zQ5h5KWBaSeOwk1xqRJNfGD0dlPtt/Cj93Hy4zAzkIYER
rKoBmG9lkcIPS0LoHqCf5vgn7Ohr7zxvBfFy7VukaizHpVp+kjnYYCXZ0/hhXJV/PzpiDerYNg8R
OxIJCYO+zCL+I3o7p+Gwx1DEpQBgJBLYGKOr3NXw99txxqImrBKZpR8gWLBau/ZcnLvaXQqTZuDQ
WDYy2hkU8MKckecTfNv+L5OJuh25Q5+5v8EfCccPylBESADgRv1Zib4CFRfWbLSAzyWDqUiecOr0
TY+8+Yj2YwiwoFgjP5G9vnutlCSEpZk7YtYvpwpSNyXarnwaAhXkHjezpyya0wdSHsZUbCJUuIx6
0fJP270b3Zdsol4++GP69Z8NnGLfyelY2tNtn3O6lesIs1wCTCqpA5FSosgTiNf1h2xv8zLPWXJ3
YTIIEHbeHWbslU6je1VStzxJorCDp/8JFSHfGXvRuxDpMYQB+/DpHECctSUeadKeDR3O8KVuiqsz
DJaRPaz3bEusf6VEtve/dcygB/vCEaTKSsUha7tYBccUlmtBmaPLFJD68xRWobmHAeh+Ifs/APgI
AUcVTnjPqfPDmyLhcDGeT9vU5OHuEx7jKj0temqi8zbxG0jgwrq7ZHbf02NlrMFNptDWzqFP2qgT
LIEbnaNr9857/GgYMjLuIrnUKo5Q0Q037NCiCIOhPSgO6ogffEqFvbYKIwGODvOjr8KoxjUjw0CZ
7gJq7QzgC5N4YmwJHAZ/gBZZKJiDU/p+38TzbW/X+dLWHeu3cIjEGnNo7KgLtnlwkHRWqWTv2MLO
JCs+Nt9+adbVQmwXcmY1fUJMeb8sNwlxDYJLzqIr0AeWJPX7PWcmcHrxc6aVUjH1ECSRf+gihWdd
FZtFjMLN6it7QZX4zSdpl5uc+5XGx3lrnyTIN/zszLwfysw779y75qkXJjYkUiDqlT3jiSQMyqD+
qALVbSlXbX9dKB25/HsPBLLYi4scRill8ko+I6qggSy0hDaSUxYWsYXgvRqXSp/eMEUJRowIlwrT
9ODiVRC9Y9pTCAv4nTMLR+7VVhInt/7EZovGEetepJjFobsP3yBWIsYHYzaS//YW+MGAH9unRn+I
DRQza5/MsaZAhLsyGU8A/AHx+Gp5EqD1s4HJu4EuK2WDzpVuzQZt0DF3sMGqVNb0eJkAkfktBCwo
1gEFQEGBeEgts+CtVd0DniahHMXyS0UoZqzq89aZr3uHRRL8oukP9hCBP591YpiOYnD5BC0DN7r1
lWNyAHuku9URjM3VATFzi9H+66Vw5dzvR2qisrtSMG5PTceca/dddHw9IX1dApABTurHfg5J8YDL
ihXDVPcdUf8WZ/igUm2gWhzZkkbD+t9psLAPcZzBq60uGJjedYnIu9MZl4cdO0jVv9rlLWy9LBK2
nf+h0cK4NkDnrr9JtZvKS57aYSmF+v2TDhYNa4MbcK2MnBT19Hc0nflKZ5jG6dUSFTM5UqiLGCpv
AaAQ7LNKD31HTWPYF0lcoPb5PghHlApeeMgBFIjEHhZFRyV/1g6V1lqAIp46J7e2y37PGpc0+877
lO6WSO3ejTiCAP6wv8Cdp9PX5AOpKb76Tb8Y3MooLozcT12CNZHfqnIOZmpcPOldaZR6qg/mue9L
e2l3+536bqkyS0bV6p2pZm77r6CjReNsvFBLgmTMXDProHh1gzKheI8mtWuc5+C7Z6BKT7dTZflq
eNVeWCA1+dYYtuUvcpKpmec+fKMVhWrQP5ZGf8ijlSAeTTPbGAkMMemjDVx83iVn3sWHjmPrIldU
OfBSc9xsQpu8ENPGVYAJ96YQ0nM2oqTjzFGfDwrNI8f/d0ekQVlnNiVR/EqWhE0jEzGcRwsX2VzV
qhY4i5pNjcf6Fsu9n0a5J2hv4jNTKNh5CqWjum961GvvPZyYXuGrJjsr+xnbr3ta6MHhYcAhG/jO
WyotmO7caE0nxQd77FP/WhbaYGwHPfu2SWFNupw9Up1K+o06asSRRMdgUGDfnLfCY5Z5i3qw4p1V
PnTJ1YYDZnt9XNdMDVb2NJqsFn6a9VchEQb0Mkbfu1Khr6ygY6W4hKsYl5GUMdV8ZhC1FkU5Jx+O
I7dyJFNG4iAmN412KfjBBJo9NBWh57KBScwIkhwW52oSPz8c3iE6aVke4ZosN6qDLgYD86q5P5FL
PRZu18hGuwrITf4Ph7L6DWqhhWgmLdMySSKJEwFq9GC69BrJx01KBqtW/0y8kigUVZckPLGxnU+y
wLG4HI9575CdJ4zhmaWMxZGsuORw10kvpSI1zdBp7EIQU1j9IT/8HWHJU3czieG37sg4COcqQQK5
AmXiUKRKLXq8tx1zwZt21YF2mbXjbq1H6to6DxMbVO38qAlhWVRXanwQ2uK+4rEZ615v0f2NIFUW
kSY8JJOxedqJNBN6aeNr1RBexS2vHlvUP9CD4KK+/xC9pArfXgOkfkdY88L1zheIOp6QLmqmiyYT
eoGA7B1eGnoVxDdg4E5yYCR0y6inCxwhQb4TAVaLupQltbSATwCw1vDRbpAUsSya7yuQFdo0thle
JLarOacHwmiNt8FtV/mEm9m2/l6/Wy5XXA6kx/gHPS02kU+1emiThQ08uHSsSLZk6hKVr9xV1tn4
An8xRJTciBvvuGlkRY6AZbTtaeruTDro3Q6NQIsEtSCqldHcOi5hbwO2KrkvDOy/mDPA11PxGxz7
v7N8rZvOzb9qqsCtP8FUxhMWi4Ao3ZgDCBaawN0wB0OoMWDXjrOwJA8HL5/Go89DO9H/aBFfp2xN
IVgUJeFMCRnqwsRdVwkH5JczJKhs9YZ71QFc1ypMZVtWDRNpdSL26gNxDgqEr18GTHksRQ5/W/I2
DOsrfEY13cnlAhd755WXmzpbVtxwgO1fj7MW0Fh6JdmZiBTASvKcv9jB0PZ59yo0EYR83smF09Jn
QD+M9JUyz/vtSBXcpXauIIZnGEUBFIQ2J0BtCNi+Up0ZAxvd9PiL+gosy6dZEVo0L10g+gjT5OF2
ZK2XWfGJh+ML1iwRSMcmcgOdLdDG0J4fxZsBw/IuKlheR6yS9U8xEW7p4aaS0QxdBBo01TzmdppR
u1sx0CosN+daC/2NPU0oIGp+IRF1iH7d8sGWT9rMU2/avtwSgf3e1sTNd8NjC65mzmUnEf9+Mxlk
jF2EoudawFN+u9A/h4KkarWl+sxj+ApbsctxWvXTQDdQpKrBEkuABw5b8KFs7IQSy2Bt7Wx+j8As
CU9RbFWNGMApW+b8eH9GdK7HvuV2g3gvq+e6pzXmZY3YNM1xLEVu+/xPbUT79eeg2eb7SPVt7DwY
dTObOrxUMlyZqQD3D7HZXEM9ruLBRJIrmoDCqsOulNF1sVsVLy4I1tAShQk/Fp2yCa846nit3wm7
2AquU86gAN9zfl3kNe2cw2TpwjCk8eHDqeHuhZZDonZqjP27rtER0pkImivEexZ+gMLh6UA84z8o
cp33tq4MFAqXnbqvSW7mf7tXX4c2yS6lgnqkj0BBe2YvAQf7RjEj8C9bYiBVXBnjgxOd7iDWUfEX
UhO/N3uJpFZveMahqAxRgwMJVom4UD9FuHyNRm/okvhSa57DbyFxXI7NMlXX1o29nsoxCbcJ6EU9
PgBQzYCohseZQ9EZv/Vm8N86dN7ahAnZmWV1e+yfBXeHSgOryinDOscQEPcYnCnsiq6z9rNWD1C0
1aFSVVeg1qqcEXbgvMT+HEQ/MhQ+4BT3PqzQffbv19+y9ejw8tpP6OeTzResPTbjLe3ZIAjk0+WH
roLCEMHb11gzF+8vM3VVJ56qWaxoHaIX6o274WDd3/xLGUiqLrBd6xcESwoRalWe80YPAActfk4a
8q4WWZHB6HydKGpOdItAcvBJc4rH5oA9Wj3QKk7NzKUJM5bCTTE9lvfLuhfORedaImBUHbhSMyql
REpOauOU0R0yzcmm3KIjBf5OP0YtPUJ5Ez5YAPunWXWfCvwek5kAxl+q4FmKvTMdXtsVantBjTej
Ry0d/Myqv6hZaX92vVj+dELFKKFgf1ssnHWO/VjJMD8I5imUye0CmtGo9Xa8wwonXW7ynFTfwJoZ
FWRpzEfJGHrQXDGIaNlVNUaoo6qXpUBo67IqnVIoPAv3bQmDwrqeH2RLCWT745ldMC0M81CHRAey
DL1SOlFpVqE3KxR5zmGK2Wd2brI2XY0L48bUKjEUl4zbb8en1eHiPCmRgtn61hW1tSbTpMAS1NDd
ZViHk7b11feRbqnsiBUsYSp4JC+uz+d1fD+TU1bASSLV3bMrQB0yyT+/8Ax0R1FDPtGxnOeeshrS
3mqiTjPqYJWVuT1OyyqVabE/G6Kl86rYotFfWrYqqTsHiOpcFGiUqttUnQiYDalqLkq9HPgwiG6s
tDNjv2TeNrA4mRuiDoXS6EV55AwkEcAIMjxB1HVQxM0tMK3CUxm5ighueugEoqunJ7C29hLLOiLV
W6veJzOKSwoQKSkDY1CPkvY4n/OdeHomVooxNnzxeVFWtr3q5BVmAYWd40XuS0QdeKZpd5T+Unsp
xP//E8VRHXzds1SAWBldiAXaipFxuCJmWByR17hbNGFgOKZ8qD/S525//dmv+IsDPwF1F8GADTeE
dO0I9zWAhWyCXzLkDJADsVNFaYtpJvUmD0cnecC9yV2X3IsKHPMB0xsCgblWRZ9COKLTym9DN8pi
wGUZ4bHtUlhF+ACJRzo23OIOeBv9MTbESIPRaA15DCWDQl/idn9vjbW+OZEsd/CkBEF61jEJEhw+
7FvLTuuVW1Z4pE9heH7W625wwSqqXAcfO0uMuCcXJPWu0Oi399+bd+VVa+Vq2fzpDW3ISPwHsIBW
kthUvINJmj6RzTUAzBnCZJewmBkCYPHAkFLP1pDq5AWzCTwD1ILuiXxvgdPr7guJ+uJOf2af3Ej2
+sGdS/RrIriY+8hInydgtxWw3G2RlJRAgKO7RdNSp3a0dmIcA+dyNfNEkcd+AVwtWv710xZguHEI
yLlCH0jbI+EmVMRLbZTylOs2XOrkV7KXnVuTfKBpQn6ROJUvLwwIlVB+RFGlf9eG+JGwQJLlkLG1
RRgzmiJ3R6f/CTJDviK76XRY3x0j2ZKC6ndsnxfIlRJCy2GLFJNGeh6XwgAdOokgeHRchllFIOpx
PWcXeVAeMWcsDRDbpXwKFWE4+PveVJS3Y4sJ6zmi9zzSkq7fLsCIFBkSjHirgKsUtArGld/zhpZW
Mm+d3T8cM35HpEWasaHacl+5bbUGqHDiKslAhx08DvwX0P2ddIe2XGqHBCciezwasVmo93d0ilnK
TBpGwaG0Iv1hSwOH0Z91uqAa6O0lZ9vdVewJss56+Med+UIQv4C3hC7r8f4fw66Xef4psVISYZRz
YPdDZKB8UUDzZEck4pBqtRgw7vpIb/ET/GvmoR6IjbiqZ9ZDdLMPZKG0LlSJmVC9VTCAPgiD0apb
uBpR38I8yQlRVf/14W3aVLc3ekNC56sUvxmWo1qtNjcet/Y2ff5XU20E+sjlmeYWBEX771S7utYT
rHPqWaMreLkXGfKzfJvAKW15qP5L6tR8vo5A1bJGdP9FgDx6rLxh/bf1jbC2HLCNTqAi/yyimu+i
dHuyeuRt0Sgkg6YeoOTWEhCMxMAD4dUfp+OtrkkdK9yX9AAr4EnhcHOEbn5ZEiHZOzgkxjbjpz+l
i2XmCuPgZWqUvGz0elyBUQVZ5PzrvqWSo4jvdM9bFKjugMVk7+FLAuVBF58eC2+ypnLGD4lIs4p+
GF7wxYHZL01h0muX+QvxMj5VsRZndfgOBaGfqQlUtvin/BjLPpvhdA1QOhZjnswHJWawowWiav91
Gq8tq8pOOkbc3fbjJeBcbsZh75NMYd+4QzAWhJBXuO3v6XRLXGaFH8hu+3F/8lEb6CC/1B9M1eFB
mt9JzciCZKWg2A2HGiECmEjMrPO1kMDtLzl+LdMn2gYff2UmzHWrzxsJJWdDhk9V3Vg53G68d6u1
6X7SGWwfBUZX9BBZdm17XnjRHLpzTKoFi5+WwlJ7cbSF1vZBE3pZ3YmBInt0KsFS9egkYOQguKM7
2c6lUfjzXKtz3PMlxcrQD8p1CanQ6FEb7x9lOExSqUH3gqcYTOYxHWw6g900UnJANop9IAI549HP
UlPoalMee/HfVMDRx9DQb3w7bObjUTkfSJzkJ1srg9rJOXxgU4kY3ccq0W9VLbYcWmNJtKtx53VN
gjC2Gy63VCe+OnZNGnhL6fFlJULFq/CRKxLZqbtDRZqg6nGfloxia63DN7oP4rfxZ5cHuxBj4chP
M2oq6ederqMr2eeGXBLFffYuQHQxCtEwOXT7huhJ1SzME+ZhKoIFhASQBC5Z4xOJxEGjthJy7DLg
LDAsaIyfSGIknV1jtiCUIbLinoR30e+1kqmO38OVGBdUh/C5PV+0SZEiP3/t8BodzkyJ4vU25tUj
YbHBk36P57rb2E1UtLDMtvmZ/eMmy1+rHAzF3avmVkGK9u46U2AvFxeB3Q/d8CN28/gsOIw7jcMl
rgmbru1CEGyUVTOwodTBbedP4acH6JVienZ+dJHmg8Yxxn5dmPEd9Pbz6UdVzTofizsKTyc9WdSU
ix9SMkZCqgSyrhXhZMmNUv+vuEY8vZlfDez3NNtgdZFGWBo/Lfrc8vE6mszYLZ7g72kQXd0bLCQF
LwINeGbKq3pJASNCnFbTY2ScslyTTsEje2HjPTIU4p5kEnryqGpg8coFQVcWT4heKlZH37sNuGrZ
2Y/oyQbzti0/OljS0BSlyZMS2Kzn/C4GDWzOC5kKMUlmKTGg6gxytferVbOzddOglwUZIunKRFCe
yVf6D0oxEQ4V17RPDpFiwal6CKS6dQdM/g3Xk4eeOoimiJ8pvsbt1hcZDYt18ccdcdpPWL+FScQU
vP0DMx3mveBVX862JS7eBY2ZW5FEME3PxgNiu4/+6VjlX/i0o6vqQmoj4KyyqO6M/0A6XL62V5ig
CZ1aX8E0G1pbMwqbo/IePRSq37vcENbx1S4LxBLa6rYFulN+R+IoyvWy/TqMB7fBwRH4oKqs6bd/
PM+zm4snawfcLakmR6mPNAZnDk4PqX4cCK4wqFl9gHbeh51eBgo/xQUK81kKOivilAVpX8eV/s5v
wxYixO5r0BlILTIs5yZRQo46Ck3CYqVZgcSY7V2SvgKG3cnmd48TuXZwwa1uMLLUwwFjIWXFCmZE
sN0U41HRdylMbBubhLz4BnXqjIoozKa9MGgpn4Q+todrQa3T4v+vfZp4Doeu++faBBuJFMc4jizf
m41wt2oonMFwoz9quHKTyHUFuoBOv1fqHfWUvcLCRZMyOeVoSO7LHQ4KnMP1vdI+jisKQbPvrrUP
9gFf+jc8hShOKkvK3ji5DodXhj3SzSMzT0t0AyIZaIj3DTVR8M3YImvtvuaZn4FzFAHmVD1ynAFB
HJ19mg4ncwN1lr0YNAIOP9ZJPRn3STwZnLghyJS60VOH6cIvNVBFYwqzPdpIkzTkWStFGlq8HgHV
o08kFkcrAXvCgl3T0pM4CdAhtQA0ldIZEhAMvc0KXjxuH3Q+ziiFbI3JZC0aFTkqBp9cNIRmcXMs
qhHuvUcWhpEAD+mL6XPLZm0qFE2OTtf9JgXHz6Xq0jmTm7KhiyJLaIyf5hKJYZaATgwqs9NLa9xH
L/GC+N4QpOU51PMT/ovCxCRRyPChTyMjkl3HOOCVeDPJN5Hh9ZfsiNblqUQzIXYiIuKJ1wI4DJOB
RBVoizf3joobhIxgz3ex7F+jnPafQPElh0sx5hUmcfbKfLo3BFx8lj4bNbW9aXe4V0E2/DHZr9oW
5waSbaicVCGo05Ogi8gfrTZPXKD3GMeMq29mpF3d329pWMuBKp7KaySMB5HGcFu1jFoQmXNosgtT
134i+M4mdqRfCUthF92VcuEAbfktVYKfXLbwH4iZ2frXvPvAMqCEZnxu55Il76EBOXlCIk3AftUd
RYaIHlwWe9gakyDA9sCwubpPxaNMgiTmb9uns3LWdSFwShXge2IXXpTXBCGLUxq4OY57GV85aj+i
Ko0+ZIWXOlK+jWKy8Fd4K+fhNer2jnAdY9/V0J3Xw+Li8hW5+APBtwe+24iG/SlgZC2sUe0vJUab
0JLK+PYBmgVQ5xLOvNeFg1kR0zNiYOrDvrnJSvfSUCyoAWIQrBwX9Or/kI6xZ18QyyiFToixBYym
I+BxCKXdInYoEauDiSvsdTh9KTdnE/9wqRZlQarvuEzC+hKvcUJDOl4eimHJspiRAbYCZE6kyuav
CtgeOPjuf8ybE8/hAEJPxeX2FSaGg27TA8FaV6zq2ByniYelT/Lz9mz+v3Vy5ORauoGYuSHoK+Qk
sqRD/FIJhfH2lV2WQdI5hKBPnGO3QLDUkXhfEmDVgbSOAn4hT03zQy4MRC9iF1CwC1wJ/IauP26l
ApUIVCm05psKlNuIKuE+cHLsNfOCq8gAgsmAz5AKCWDW2ORopfll8MZhvyUuNhkaDuFaN8kUC8ae
lWTInT1365Xj9q56doClYeHPlhUWXcCVF2NJroEFsYnFc9DDG7+XhJebZu2QTvNxEwo11rpetbKk
XtsRQTFEFeawWDXChIFRiZJwbvIzfEYcC9hBlGFlAwtkt1WcsvJ+OdMRq/SjdzIWdaI7Ht07r+eL
CtXrccy642QPXgjNLWkydReEvl+bu/DnFKoXeCFYVhgDkQbhttiWnhjMCGTOTBpdlSFOgw8+S2bi
JElVTz+hxCV9wdkWc9AjWzDpjWWjYAfPHG6Yrr6rocsnb78QjOL6HKd+7WTdp7bgmdkGp+JT/Kw1
ks7OYqtKz8vjI45+6lJ1rI/pHDFanmYo2hc+WLGMs8LS6/juVgdtI5wr4tgp8R+g3lGtXjNf+qOB
YGRRQRQQvRAJ0QVjMtgjWwEBmCa4qHwItFGgy0CkR5o0/eKZszztgNoSxLisG0/DcgDFsRDunsTM
iw+0RR7MIoilenDJoJn0uKf3cIvurFBWIKnOwg6HQbG9sjG7LtZMipFOCIlVCdqbXhMhGlOpWmdV
8P/fdf/XueDRuvLx8BgntnRN3M/N3GyPXaMI0cE9KufWGbfWRHDPNAsXj4eyA3njNhda01QqfYIO
yRjClFXxDeX60f1yRcBjsfJDe+HvGPfPbi9nYH6e7gvZ5pzhGL+aLRq2ZHR/S+ArttmNRgfyHYc3
bOgUdnvpf4HpDSJ//BksO+i0t28gHs1HcCxduTiSzq1utlD44bVm/rIjgsVwvTpUO1nAt6go63/d
0E6OLWSB1hM0bQD/QkSkkJq/5tEmH+8JEKQTx/43jawwLXZ7+lllPCYS0i+A9bUFfTZz8hW5y7wE
zqnjLEfJAZl/DY9LDKeYo77mTaf46U/VvWvmX1NTA2U/KvcP2swmQjq3LNqf5VlLH67td3ZfGJFj
3XrDDsStiK4Rgb8IASQpcqmeul6gWdbZIx1WoP8chcrhBg3XHMtlmRsQa97xIRpLd+mF3caofOkW
zpXOvGTdsXvN66ZkUNRsOhfOsUO2DEmA5lYZu8vjfi+VoC4Hl/2DvJkGRyhQxqi78Q9RYDR5Kw89
Ry2wAbiCfVe3WBpYvr937pvJyZEC9wdnzcMTvjmat1krnDped8CCLuoNRAijspbRiPVrm3kqvdT5
4WxhWFtf/25GeF0tpZIuyE8GNHXxmlj0U7D6qj9UsZ6xVF4A72IJi4KC2JRbPwr5ZLM+/1PhQfxF
FUZQ5zQEgGLYXRhPl4SayN19zYGajv/IxUg04bUCrik6JKyP30+MtYPl4fiUWhLz3s10zPI/gGZT
Yv31SzF6K4sa8CRA6pjQykW52+UoS0xyLWw9S5jfaaUpnCcWj2GqGiUyBJDK1gGnYhJWJdw2XyOo
Sp2W0/P5KzI7OZwNBisvpn5CVsU/riaMyZRxaRW51J8EuAENmpqx0vqpH25dT3+u256YzguV0nT+
e5MyjWrQuwQqi7lZ3TO0yop5Xngh1eCKRdtwt2dAIp+IoE+2Fx4L5CvpzMcFH5C1sQHsQs3UD1XB
T/y5uWawITsP7VXd0K4hXe19ngDWjO8pzYN89FgAnhEeNZCdhawUZXVcU9CnBK5t4CxaignuTZtE
Ab+edupuPHYE+jb6lrcuSpzqD/26Dof72Z+HrRZMD+d3vqIe1NPzJP40GyaJW87zY1Z5hq2dp1bp
4naSB9gYYN0FymrReDqn+rYy6CkNQc53yQtSA/+MWhYKSs4LiESCgT26f9DW/F/S2S3taxNOUw01
LHHmM3Z0gBqDaq8GxZ6lKExus/jWpE1K9QpOSXhfZdxJJFeG1jEpwgle/6I1Caqn6yrWs2qlud55
w2KOkauL67x9WVyMi8clqtv08TZijvCNA1yAFgdjVjIyE11lQtOtcsH5+O1D38K9UES7yHowHsVK
HcPJop9IquAx2cJ68T+5/8nOebvZrhTLgrlBmaDbnROIwxNwWZyMzXpEmMMfw8w6w+jCiy8ZNaHd
9t1Ej15XKsKT31UbDQijJGNNa4cIRGWsZrw5EAprSDoASXu/RRTehZz6mXA50t7SSWAuGH+hCQdv
Emv9iGPW3JFpDsMjznCKAe6bu017CWeqKq43ZhqswX0Ad45OYN6vp17QDW2jWbaftLCxwRGFdRj3
qfUsAZaOx08douxTmCC8bRkJFXCmLsDeOHds9NGCI+sk9CK8PLOKtX3vdofqpLwaVytBDDoTK/q6
ElXbxwsEeLovFSIfI7xU8MafYVr7WFpC4fIFeEIMu1ZHbmcgLOlcKWAnVNjCjU3A1Y3+OCek0E9y
tDMck61j0IC6J/55Yq7EuVEu/jkPsxQcA9Dr0AYWoylfuqnQ/CUlUkN0xk8tzT2ikhYQ3etZYU97
7f0fo1F1KIpxy7uRMUO7e4Lu9QBCXumP63EmfExXXUN45fLKBFjK8g1/ttko61TrpXAIxo60SaAV
kdDclDP/3qOnp9qAuF/JHFveUgySxLovTlOttIIXnk9SOJrlALlw7Dg4ZOIZFUB0XL0aJkaQOqHE
IPa8AT0BkWWM5GEMEASU9UzGDvMe5hnlTq3ZWW1SLleSEGnHh+S69eFVPf8yKFvyfyHs9/xSuMaM
hGSQUgo3etIRomvuHbOdfSYHZDjpQv6m1lfpeuzjhKEwSSeAw7+j71oV5MvQk1cdgEVOH0sKaQi6
jTOtuVvK5/TuQcSKObGK4l68L5dpgHxQAGefOvLbSDBD7Sd/XltwqP/4zqgqGUNGNb9FRcrvl2x8
akmOlT26mHhWSs989n96dEWwF8/OXTagxNIpEmBhQ7lbZ9l4k7miCzQVBqHf2Z9flfeQLsJehjWR
JGSpbPctvey4xiEKNoWOTy3nOPFzlQ1yoWumwzwzBPdt4UkRtzrE7ygHMP3hYnyL9uBj9Zf6Uo/k
0Tuzvy3dRo1WW5ka5hejxd8etvLuX/e2fyQauPBQWuporVKnZQ+E3+S8h8yt4iMcf/KGCPBAScSV
IFR/UaKxKEh92djfeNW47qQuvwRMlerk1ipyVxi+wQ/MRWX9Tz4E6Bkw4IvJrT4mVIjHTStae5PZ
G7S993jjrL2aeaNh8WsBkq5224Vj/G0RDwO4pMT94GVMxfvm0kqvu3FHSfo3ufdM4K0YpEk/Jo55
59vQmU2gDXCqM/rIMpU8pcD/g/peFdqQcNyYgnqQ76M1VGnLWWShCnAWxx8neKCFfsJwwwbG77a3
uhAwXYymDPeUFU9mK+1NHCZP0g9RQGfF11XVYshKAqpF7UKB+2jpsV3wWHOPllqSu+aD5Mis+wLU
kDTRST9Xt3RfA1plfPLR2a9Q1UjdjZv7Rk87LCPxYfSMalANH/NrqRe3t9LCd0XTi5f0XyUTbXTY
3hz640pGQu+elANwn0NH42GDZUAP48wUBlYrgxiBpwhDt8XltiFXaX5/dK0ga+iEu72oT8dNWIHh
TXlhj7zWw1+GCg/bpKt2G4HKxbACqJshrGYwEZM+XoZk2seM1593z4h531WXZFNMAaiYcEQM/38t
v8O31tNnFp5CLKK/un5kpVfMGbpee2KelyacG4IljPW66eZjbOxDkNLgyqHQbt2haaRFKaL8yDoZ
K4pzf4bDoqetTFvvC3IssoEvvKT3iu4gKTmUMXU+q5Sc6ZsbZirOPeedlV2FMT78vU/yWuWj+Wzj
vHVa3/WVI9B3+FE62td1NCYjxxEAoa6RGRhS95GORrzzrm2cQOBSE5QVpmixuQvqw2prPXJ+0Daq
ur8E3/GK2VOErV6t/3zGhSZyef/TkT79StTGeIq1UJzbCa1GkzpnUnlj6zh4SOmHBYkWj38FDccb
BsXIHTrT9SywG5yVMNNBBFCEqlGiYLriPoUjzB+gwkCYKFFZFQ7F8iykdUC32a3m64/hnyPeZPdx
E2yls5+0MCdMheHjExLkybPmMboNfrsoxu0jpYfCgX5NlRnnobpkIXqAi4AjxJ9lST6zrYxqWpDV
LDfTb+54nmxxPhJIgWd4iMt+FW7Yv2v8fN8YaDYV2sxcLABQvBzlOMO1CBfIAA6Dz/DeYNfKnjYH
oof3xD9EmMDVLmm7lBO4BXIwLSfyLPd82ZMojiPjGSd23rwH9UDqz2znKdJywU/MnO19D+Xwx4Mi
xjb1sL3IE5s/V16C23UqwlNwbKrDN0KOIbCp7BP/81JvK0xaGRwxaSLbUPTP32jUcsqhDSNiqMwg
QLY1578GRc5Du2AHcLp6aRwoWNayQtsoqvBnPaALbzu+ZcZ1bWXDpF77r8/GiGKiR5GRNvN53aFc
lysG4fIcUk6D5XlS6Ajtm+TkkLIl5Hlo05J7teC5MNpKkAW+AXnrsmsPUxVCiQUsSoWKPqIP1Bzd
Y3C5+j+nP+kRS0W1z5Uwz+8CEAn0bjTY3vYKkqeD3AWBizvz9MDoEvXMwq7FHHrhBe98HveQ0Y0c
dwpno5I10q94z0XowJ/gDq8OGE3q8B/VCYH2nV90Xulxefb1L7PhbJ2NK4d1mrdG2ACR4UxhaT5+
VR+c84sNceZ6XOkyzdCiXHUK/CMa4UQ+UI0CKt4Pxg6sCaP8Ub9GBuCieJmxHqK3iJ5nk3jJhNOQ
fPF0yu5iYAwouFy2jgG6SFMalnzJiqY2v2oZNoV/UYHEOf30O1utiDGG8edE7vbG6cDllCt3A6LE
/DLtfBg/ectNPjchxro29NcYwVWWAytbVYL1gjHoj5i3Z3F+aA8dMrcjFgi33KPut8VR7c4yzn1i
qL3RMUrrenmR8KcwUG3FFKt5T8LallZ6aClMGcnwvoszln0gb+67Z0zUYNVaTuBemGVcldNIL31X
c6JOejwDzZoiBHHWXQYG2tTMdtKNjuPF6v9wXDP+S4ntMzu81Mca5vrQLKh2vtatLKaOG+w8jk6/
Pp0KVlrD22gK0kjCCepICDIe6sIdS4uWJtrguNoPtgkhy5VUjsCPIo0p8KSSFTESIdpzaj0RgVCN
O1Di1UwMQ2nme4ohHuZ8Gntjv910NH6eNjSEbQ3j3qY2msUGMJUgfdzWg69nUKGMurgDJ2cl0AHh
rwLOMjn+V28f2JtyjjNzZKu15BE/MyQVzv9JbmwGWkLe+YKyDRTgGSqbZPu0FWXoOYx7mpCII9mY
EaJjFsh0Js232e0aO5Vqq3T35g0uPjHKi2S/j6eAOPrhW/fKRpr+TTVwd7fKhYPptlgecQQi/Zix
+bg65w8lyboVV/L4DJRX8Ig3MDZ7uL7PyuscPd6TarpYyH067z03zFm4WEmigCSy2LgRAo4mUNga
7wSW8c0/lcEDodHS+x0TywUAuYzLZM0DCES46zf4RxYzugIYDqHc4LO6DCPhM8PJm4wk7w/enMw0
1+ec6objMUTG7YfKKlw+70j+SCEC1Jnixa90Vq1dEHY6yOCpMGwVlX6rOKFPkl0vkL9lgBghTR6y
3z7z0WjAbIaF9p+t3n8DxGBvgcWV66H5r7BtZExcqvRK9Boz3xJiIP6d4WtXACgOmkASbfiwWJyJ
Mxo+ez1WkasW/8Uj9QoFKO+gnTxtuOEJWM71pY2pGopyuuZk3bJOZ+1Z7KFDAISxCGFeQcRZKIAo
4U6+hMLYlk8EJDgHhK81d4fXVEtbGELktvx0H8GKKyhrkrYYCtg5m4ZxWAJsbFX9E88V4eUkObdM
tvYk94QNNGuk8FZb3n8T1hoqmi1wB18C7L81hTSTDeYtdqEyzFIXen20dr+AFqSnKF5UaYwrO/YJ
pxqbRoaMgkZ8t6rIuJM74EJOAdkE4UE2Yt5f4xH0p77sHfhQG166t7BqDj+qfRsFsPT7txJ172UY
VxyNogyb4ab33FCCXoiW1YPr+hLRDqOH5JQC4jLUfjMizMROdRGwWV2W8LMNrU73OrdwYmhQjgG9
PrIVmWdKnxbHCm9Lv25f5LMlYVX8ASUg1upjml5S8Hv62XLKVgn2yLX3b9vSHrYgsCpYqPVd6h58
ey63W96qaqEzRV5GKPEkODve3NcTsGmU+0zoE3AQPTUUks0dOqav6u5D/zdIYMcVy+fSRf3SZbCh
8gAokXL7UESe0g9wRmGwl84/y0u07A7b4qwnnNoFYhF1e67TA1mwt5axA36bEHSmT6ZU0YLHkBci
Z7YdsEl6AzW9gxfhBO2v0Z3dBP4OotoFzTXit+wUvSxms7B4VA8ffJHFp64wL5csU+fmeD+IMDZT
KNUiJjkjrl8qFzaFhW+rcKg/mt19rhPe5vBzMq7YJCZpzcBJUanfSQURfZKS6oemajPB6EigkNUH
VFoFRbLNPlhgCPmkComKIqREIy+24OxAEpwgM0etPeXx6F4eyTgXaM1KW/NmFSRqSZswDV+tfGkd
RwNSQ1BWwXYLe0qsdvAnHw1iM4C6LrcITpjZVthCikIXU2xij+1+GZaD/w/ekFUGRHCC30Z9xwF9
Y7EcfX7uuxT17fh9w1wD2yXS0QGBMP/JUHQeehD+KReANlZhfqEzUT3b8v0MIUJS0JzTob2Gnwli
cH6AJWxGfjlKnN+B4zIo8EsG3qwZ2W7ugQbZh0LDNRJDTiokO99N7/ItjuBYi+LCVXUwXQwXzs6Y
SeRbBwHkzv1Bib+BKtpA60OGcCJzQuNtWWByNIerrMDa2T9PoUzWJ+/cljqFdQghebw17Q7Yx7am
pfQKGPfeAc4YbMERGpemoNk/+V0B6oY9KThk9h1TNqs1tfKOUpSSYTesL9wa+hFOdC59mVU3r4JJ
usc1qv31xnsoatjBVWdEcKsUHMv2FhOLhfn0GQAFu9PNDkJ6WjWQZTgQtWv6Z7FPdJ8HIewUDEdG
CdYQMbGO4cqDDOOxbaE35Y98ySZzDAbsuBcpxSEzXbIvPYNffirsG26QSPUy2i2zRxQfTVBO/69r
XsTh9BmFwHdLP4on/O+Q6ToCNRjct3JKce/PyX77Q5RkRxM6LgmRsBDbGC2JXgcKf+5Ey4PIuVPx
YXgklrRFAeg0e8dcV04AktUXEzi+qj05V4wgE0K4I1vjeD9RSQkxgU66Lbl0ZXBS0qffK49hBd9G
Lz48hl6P9XgRRvaTVlIJthPwAhFtExYDbmkGY4rhB8w+g2iaPNj3GhhoP1WjAyvLuGRZr1y+zkkP
nH+pjb8Yr4ihrq4vwTsGWIDQ4n+VpKM8sck/VUB1IeKZ1G2bFjCZHb0Yq0zRh20sGESzoEDVFESV
S74+ToiY8Yj9EKEdHqlONz04yPgzAAe4A76MSL3/LTD250Vr+fqgvpwDohd3lWJTkZljd3Pwc0vk
EzuCZuGmK8mmPA6g/bfQJzZADEyxJxrYLpnNS6yFpB7IbyryhorJPf6AxmYwYRLfqXfFPaAqSq/H
6qY38hVhffxbu8KnCfi0yfResWRknTRkDatc3yORnH8rdyiYm/ui+zhz7pzJE0jSAFd4CjYhO3hh
tiXNbVGWOTFpBt3hfQwuhYt91myXc0gq6TVZIwBQ6z2xdW1JPl1p2zyks5dja/AZ+Vn0fAyp8BPc
O3MEUMQIBdE9TTH6SUhYchhpx3IRFIzXdRijg4K0NYZYyT966x5WTT0U2KQuLzH+VSgMx+Ojozpf
saYsIy7dL29EDrFP93FyJaIFSB28Sfm4Mvp+duSuG6DhkcRC/aAQ1EThcN9btbe2mCPNb9tujkor
XTsTP9zPtshMoH3ukDSkbHtyXzyUyfOJWtNuWUjg3F4f1nrhIWI7sAioCS0M/CMLiP13TG9Ihe36
YW38ZmylDJK0VmvaCWraUfF4D9A5q63JZThQx7GA7rIPwyHJmmUUnEdXdUIYJUyI2BlRVrmqJfyG
wHYRNVqMXIX8kzXWpDZZip8D+eaxaUrtdHyAt7bzutzFX5D2viIiEyY7SHFR89eYZkOY86lC8W2g
grJ8ZSEFa687xaI05AeakAknF/azflmScCt9azM2hPtAbk2RvCmozPCdYxmoGelVpQcMo9S2Kmuy
7JaDirwT0KL5ep0E1MUK20W4e80IF4J1vLNxE7I2np19zGpZX5uCibnxAPM/8wrhsvFCUAeReIo4
0KZwkx1JBjvf+vVJsc2+uv1UJ+wEXMIf5Rbp1i1WvNLDQwfjsmSCy8lQwgB2Mc8mkgEJFbskiDw+
3SfCxGQf7NBkWxIKKLcQmsX8tHBNYQKkDk/5fhYiAwb91H9VF3FH9ILTxs4geVmKQT6lltQRWBrw
NZoA+oGr7kn3RajdlbMxQqmo4AWeERCgstM4ftiNdxuF02nRTFkEsDuY5bLeAMgW1wF2ZcnEd9PF
K6b34Slryx4Irwr7qwverUCZRnVNc2dbGDelomT/4S/dQvj4nBjlsnPcrGwMywKOq83+rlmqXCr6
x7Zfilmi/Ivb3PoTYMcO1RrPel0xiFxTT/zYQmlMqFk5nTPWQ7f1/OWzY6t0tDiFH1qRDAaitLzA
ZTggCw6AilUhKNTaAHHJJNGnx2ltVPrZpNf21aMNsnIAn5camVx5DwBVLIz/l2VcbEAWc9BkFNMC
mv5Usy+VhdBQw0SmOD9HHT7+fbOH0P7HlWWuFbIDa86qc9Z3kJ4afecaBqRZg75zTIroTSt67fgy
/2wzwXYcnj1SPT4E/N/c/jmZlTnq9qpZKGGKiG1ATFG/jpED91NDPK70HCvnByz//SXXSo6PKQeD
w/TCeWTKfAgRokC0XX8NKQr6VzkFGcJ/gTQd/673mtNkbaMrQxYJVSyfvli7jx02zCVrww10cu9T
nVIpvvi/vMKB/lCdNOsge1oiTWS7IDaKWfenXkAgtoFtcsU5n9HdC6ks8khI3RCO8AfpaGrsYutp
fBWz7gLcwNE1P9QkAVukyqcSldxMiwqlLSTXtHUn4MPg69joWPZhN77e2tenqnGFvHGvJoPOv/in
EO4BBhJaU1eZNpmUrgowzGolmSlhTE3Al115dqO6ru/G71/SKEivelnDQMiliPzABkR7t8i5Nrgw
vAL1CwW+DczAjq5NYWgKWQmqN072Q+lzAXU7XNC2haBnR4AJSbYc3CU31Lh7zzsFnMnF3zX2yd+M
3gTZZmWTw4O5Y6QHs+UNvwkA9Vl07K90b2+lZq6ZmVElP9ZB+4ulzgY0hCJMOxMiVErqDHZnQc/k
+GsTPL9vqsMy9R7/8o2RFrk6rLI5X1jqYcSXDD0OHwdsMDr+uduATmXisQnIwRH+bzxg8NZhis5E
tFBakXK1pH1VfOgA/c7HXNMYVzn+TiGp8B1Pe3djtCUYv7NBySad3R1ZfxUhZW2Ww/0qXXXgT87i
tR6ZHB3yMn5kNBc5JcPq73lVs/sFbb2ebfQHMnOXv7FCk01HkRkXXl1TUmxs8D8OFOCQiOKQKEAQ
09KZSeRnGILvx/eIzedlAnrJu0m57GZc/Aaibgzvgyp4Ka/5P6+DoL/Nu51buOvnQmWLw/Tvr4GO
xZkNez0HQsoT8LPJY0+AuI2hFIb+6SwhWgMJHGIsKxdlBm9yeTJIvXy5AvuRUqKXsKIwpvXKDbuM
/0fkPpLvCBIj0gCCkc0S6t9tRELKCTIxJnPEV3VoYaXd/FJKTajQ3PS3EK+mOAjPZcGu/YvBguFw
y0ZoVx/do0nU8dn5kmeDu/+YUJk6fjOSfOixM5ALBascHqlw8vICIjQVtERyb5Vy16o+uxdrvkih
Ne1GjE0Pua2jgPkmVqzAKS/mc2310dbHd/9rWq22+Q+4SpQOEyYocpCMvc67sRxMVRCgjVIUejjM
ZbXsur8uEE4D+GPvF5RzBX29r0Uvuv1IYgF1/P0IS1muFNtbYNo1nKrSrOIy1Oo0OxH72gz64bG7
SL30wOknAsVp/USjbYuE+cOsAC3qkSu1GBRtVg4yiOUNQ62XqByOJ/MuwtFm5DgSiMF4QLMdXWYh
gIUsFrEzQSpYQ0z9cDSsLoLuQ/ox11ti7WGugQr1KsBMrV9TDLim/3IZu7CdBR5MFKFIZ0HKinvD
9bqgpbeQKmrTSJRuMjE2U4mtfpX39Egvy2IWGw2Nyd0boTaWCxwXUgENtbEd+SaBQ4GlnmDNaJ8B
kM3gwgmOxftCkLT2mnuA3DK8N+GYEKjT/O5xDTkIfzvbkCkuxX0IZrkb/NH5D4MGYgZc8yG/Ua0c
oKKOp+hNbwn/YE2DLlg6k+6411Emro/LgXcFQ0/1eOJFERKrl7d+62nJLVrX69ez1TwiVM6Ta8xl
900K2a5QpyKiqPCW51o0EHe3pa5nDAtQPENT2iZRCvPKlz4CBc8fv/sNHICcZEbn099Qv4eFklGx
RT/+zGNNzLvQsFbWn8eg6ZKJ+K6ot8U24H8FRkLe5SSiuES0gCxgjxrSjEcHuM82tjOWf3G1xR1b
r/ZB5dtSOGhk0HdB6EGdccJfP9s9T5C8myD6iwkvdP2AaduSoB5EiMWYTYppD9+yim9/ZzeuZN8v
WrzEAxWoHQmHXUVcO9/sbMxpMIkJQowJ3rBb4LurJ5brlcOpVIGgCZNwcd0OD4zMMna25/Dc91Ev
jDrt/SvFXlMGwCHft8fjzZGTI/gTf8BlQO5Sngk7La7AFMq82EEiSxf7bAnBvOVwxZEt0EX8sZrn
u017a2X9qFLW6C1gFLja1RuV+4ec9V3dheS298t7og4RxsI2UC3HpiCPr1IKNcqKkqCRpyLlEOHQ
pOoqpciGvFCg5PWhnXVAvYXoBrm2OMbnE/1y/2/6qrr5t6BIKIq3o+UyBhaeW0Ji19TSmKueHMkf
6+si5a7uYlIKS+c3aJscbmj9QhDRjic3XOJ6jVroV4dBzPbEZWSxEPYtcPcPpRB08tykkKBT5s+Q
nlRFLRjbOxdKmrdPNKXf6h/MfztkrvL0HSlvQqFWVN8T9PNJLF4emm4N9ksjWr0JjBh4xWibJA7Y
zfT8ChfR36gLymO+9oFX7+puRqU7qmROaYXX3TRu2gL5bf5tS6ta+XHvL2852Lpq1ngyNqiFm1nl
TjO+OsdKFpgIEJaALMUhDfYsw/3y03Nqdi6yLuxgdfuo3f1ygp/LMkfV7ovdsTFmmAh6kvzemgnB
kCk6osi+/ASFu5Q/Ju6I82zeoMQGeKTb6u6DtmSjlSNLruY2ysOc4k8xi2bKGZnzLXx+LMKPFBaC
lYUyPRoLuErv6FC19UNb6Z3HpukKDKuvtYK7tefJJKY1boIz8eOQ1jvyUN6q6gRu1aD94qwPXlyB
X9krb2D7JkpruYSvFmo40BZU6aPGBR2E8WN3d/60WYquUJcuCqVtHCJJmL1NFoyc2mjo3K8KEhHo
B6jUBm7b2ccedUwWizi1puJdz6yOHQWlQNe5BQt9Fh5uhlXhrmOGqsZyRuqAqV1Ng7t6aygpdlR7
JuWXEF9p/wNpkuM4DNclewwX2s0NIWOI8kBeL1CZCyKtbMBAyBKf5uQEL1i2uwny9FawGQENG4tu
nCvbY1C0ybIUB1MOJ+fBp3EvJ2dhUArzVDeuQ5RbE35mU2a7cwQ85OiKa9stjRSb+xtJunurKHT2
BiSer8Avu7ttm0u8OmDvY1XPIDgC732+qlnlz+GOqBN1IBWav1KCfHy49+51aIOiBne2Nnz8AoXL
vrgHrQPwjjzEVvnDERdazLmFb6QRco7hDSATg/52a50REFGWlXlqiFcPhQDVYhRP9WIuJ5EUk1sf
GIXGmXaReRNum1pShOelc4v7oh6ASE15/FWj6Y3wlTnvnOM6c5/LfdYA/mUrtCdP4OAMtTE2CPaI
LirruiETwWWCCgA9P8klCjqrbyqX5dPbKNUyATKVN/0F1rvHNgdijJiyXmxJ1AxLtprjr85r8+wq
RXmPox+NQV3DHlmKBUi8cAH6SKo9OrJOpIsopYb+z+3X8urtNxUKwo9+xy53bGztIsnKcPatlH0k
OkZLLufKAZ9idlr4TVah2LHwilOzIc20wkBkueOuTZd31Q6rru4E1UNe+7US7dPz7739Mw+vHX/9
mouSLynVATdV5Y0t/2M5Fb8maIQ9nzCPF1QvxqprACf9B53vchKtle3YblvvXa7OBumld2czJHQl
OKFmrjbRf/DaBPHXiaeq71bY+mpFgT2k5wCkAG0K/3j/AvcqpFhGsTwvFe1u4fG8T8qibEf2jYOW
07snXn3Z6Xl01+jogtyyRzrjYNaIiRQuv26KVz3Gc2EhpSYv+WDqmvp8/G+4tzDN9eMzzzlCXjfn
/KNIgLsMnLwjiUWwpIxkWJslixYyWJVMZFgoFk7eappHxuSGXrlYgEgLNA37XUCEM9cFZ5pLAi6p
OyExAvupc758SyPlyZgWVukf3mt4x84ZJSBURrPHq06a1PFLOf1kLw3AaUbGzMHp74eHhuxFiOPS
eKhyxSFof1Sv3m+gC2JRLYxDMAWlJiOdibyzRRMg50cgstDpO+ZNQJ+CoOG6YmVIoeQvZIHXIH0L
2FnKE+/TGRrT2bHIvS8vbuF91D8o9VBLyohg2dlAY4we0gwuGOacODkTnArI9WlgTyc8Q8OoEtmh
DgOTjA2fU3SarnV/Iumq36/yHeJ4i47Wyq50pOoGBuIS6NKwT1krbO/sdjAK6DQ7jlWqRR+s4Yem
hLIy9icQuAMFeNuAFlfQqpngf9UMbGhmHD19vuxzPU/ErO+14WobuzJ1Lq2CqTxpfomRpJnK0bTr
huCLZKY9iuLXpz3qs9/lUVK0OHcTXtg76CT7qBDCHY81c59Bj7OumKqAe3AQUGbBdHFLp+8/Mt8l
jJJyCVpY6SGvQoexlQUdOa4r6zpDik+A+FDXM8HtAg4repP9+1wUbJwPFam4LkhZl6crBl8+XNHx
qhQPQRut5hXQYl4pIOF1MB9IEJH4izwkGgmjUpI07otM3X8Xvvab3HIE83RoB/aUhO15SfymxQpd
qquvGfwS0oaLWYshdY3G5Zz4sXNP7TQ/YSwp1Z1OflZ5ukNtQQZQjawlhQy6rjE9ff6EJ48k8XqY
TDLyvjcyWELLOE0X7gA9sYGyPuFbmciWTNyJ17Zfui9YrOTUV8On33b8t+or6uuSSdGYuViiKgP9
evCV5urqnshOlgkSFwMl+y9+76FiGkIRwhJAGzaz92g7cTIiV28e/v/b6OV1HcewxLJCgehqJBYc
uNs7vTgvW9PFChL/8rToKXq95nswaAwyzeux7kUqRQGaAsl51D06jzo4gv/w/cQKDU64+1AVigk3
KaeHr0YlnjuvzWWTBK3sKUOU8COYx8the3ZdqOl7BIDQ8IZ1H+9GX4khkpqhH3os0PNW/gl3fvBs
tIT/UYXHT9KdwNVdYIEmZVRr62l5tZXo2KbDu+mJOFSssqgcDcpiVYu8Y3wTxjGmG7qliZfiRrzM
adccDiavk2DSY47Tta56H3ni7/SDMfwyg0nFmOHYGgcGQ4wMFY6+gN6U9ihhPc4N37YDHq7Z0kS0
tT/rE3I5AoEpOCfJktqnJXg2vfPdykBjtb4b+NvRNp8UuJLMu0yQo1E7h2XxMO2DgODp+5wYVcvu
8FQRVDlY7PvqkILiIyANakgIPH1HrmNrp4+HFKbeWppk+ZJWMgB69iAlxr69Nngb6wwoWmZ68ZRi
6SYZBgkGrvMVfyIYozgtQg9m6NNxvo1cDHQiFCV6k/f9zL2jkklnzV6vGozNO+qO3GVjgR5EU60i
nn2vwpIQ3btjeVbQ5CslG462EZFtWyraUK+daUXqrxGJS8cYazIuzyy8SN/Z3A/cDr4RyE+ueu8f
37ugUs9mpxqvW0BrantzjDsFD/tV/HK0h5SLtuCauolYKBRCekn/Ssoevuy/8iuIzGOoNYtGqYde
YK69i2c2anXekbnYKY1zY4R12/4TSUt7s+dOJKLqwMBx/cM0N+qDIyW82OXX5JENCA2Xt3c9hvMF
ji5epNufD8Bp8QC8rNgrSQaynDMKpGyHX1fPmbX62Q8bHKWLovNPuP5MthaLBJjHBVDf0gpEwdTN
azWF4yJdF0Vf+2hnyHrHstYuP+t0gVPJwUilzgTXyVxE1rY1bpKXcebOsPOyW963a1EYMBkE2BER
6I5B1G5ikP53xIfSA+LYaJ7fFdmPhOUe3JwSghqvReHUEk435L4V2IZ8iNw+qSlZCrkbhj2f5hDr
42VEsw2h5prwPew7vmt0lr8zNCEI4YQzdIvAUt17KSXmSKBCCvWsRYm8rTQU2XwkdP0Ksmh1ll4J
oNvVCEe4czUBvmobwpIrE0efVvE1ZGmYVm3kkXV04uOx8SB/OQRNw1ecrJbi8v2xlxHYghuRz/FA
fIp+olNZGCgnP0htWVH99gP2soAHQro9CFrVFqbvZlLqxZncUZ4fIFkIHR31uDsFhUZxhKybLYtZ
jzcOSZxRrtdpogKPCx3B8TxgzkT4c0ca947F5JAmae3n+q1lRDKMFp1xrEqEIZKoISm710gpzRSV
FG4oXZksSecKxEfJLmHSW+84TR3Ym3q14OV3dyEtCnQHPbxyU8VpZgA/3ktC0IMtke5uD0mJ62Mp
p3GahjRMP1klVoEpNlay5g+jMS7oFk4Tz2osRufoZCB0B85gom2S9iOtM/D5SmmTsIDd99t94RBO
Sqn/FRDkQ/DX6IJYViR1lQhep4Zl/4FDDzlUsJNIddlZtIV9CaDgGVO+nFYXgaPevZj+gA+6fOSE
mxxTfWWK6//ZdReFBsUWP6tNGFrPpGqKEbWIuwKY0ylPDwdrVB0l8zT62Un9q2FMu62tVebdRCPu
UIdcsoRWBdNpCEF49Bva+4jk5aCXgrwh36lAJjhDINB/kUEx/SGi0DIBfWgu3L6Wsjy3OeGV1Y6H
xD/ig+e67rgryX0VZizqMS6JfKpxwOvcLhzSzdYXfH3NqbtM+bz311dK/Mvu9QRzOZo6+vGbXyN3
BiF31qyXOFjUWXpoKN/RmwNzDijFIqVXLPnaTpvK+Qc58N1+k6benXu9haJ+h8mVZnj82WloOvxf
HH4Um4K2HT0z+n93lt1v7Gh8xm8tyXrDaE4IcH2m+Xmt/xxNPGnt7gHjl+POuXIoSr9RYJAeVeAd
OwVvy0mXuzGMp7HweijuHbhWYqt0RMZr2uIAFGLjEqbIYABhQJIuxws0dSAhacKL1Yjb77t/J356
ZwWqzX+wMXvhJhdWOYSK5bX5gUEmiV0T16pKLK2xq4iDpB/wW9uIJL9YldHZB5L25LW25v99XkR6
dYPVbFR1efvv+utFfKTixJ4Ag9LAm8HHiv30k5mEGrMceaJwbtY04xn2iqqBveI2YPIcs3zKWVZc
8uyba0gpGLm6YRbsNNmkdKEIBXh9b+LuBsegnSwrcabDiq/zxKoFJ7uxyXDP9GkRcctOebMHGGIW
/I7W1x/qnUVDixyI2Gvs8nbKtYE1EwQTh/LjbCyT6ppQN6PVIGkLi5dnS7xaksKYEqW4Aa5NDrOy
Qq8zLD5J5a2dl14tlLdmB8OzD0T5ZWKtst2vq1E5EKA+RgEZ3bSPtxNSdx/wraLi1l6Lo2noc6pf
0Mkw/7KBd6GcGZ2gAS+SlwDVeYEFjbglWqaOofECWGzVudTrXoONZ9P0wGlfQb7FDdu3c4Xq93Az
f4C2h+0n3wAaL2OAQqHdqzJQcub2ZfTr7r7wQyMClXpbA8CRhh1WEnQeBDVOwB3tkUSNe45tmttS
EwVLNh61zfp1Wj5wf7kNCaC7Sj2pHukgYnMRn5HZpLW36jrovtj6OXHWkilcUxmk8pLvfpXuUJ8b
Vvmb55qbssCS+TzWhK0HYbBNN4AMKRd9WTUQDYZolAT6bfftZVXy6VQxRrED66qN9PxSk/GOo70c
5TWoAZ3GhRp6lIaz+FunCs0JaObM71eOYNKhD2ok6PaTTgSljYUaFQtNqfcHU1jVtaj9KA/dy+Cq
2fEfVHMBJb6HDF8QkvPkVJ7YVHeAEhlEos2h/riot7fiOhsORmiAYM/l6CiBR3h+xfKjJZrNCr8U
gces+uiqR9eUGlok0Fod4SEhsJ7KQCqcZLdht61qvzmqQ/1V+0pdJnIsBtA4BCdk5C/VcuOVpVrx
P1BZ5d/koes8dcYhzq6fzyGKAwLLKDSu6qHMZ+fbtQVWAE0mG77fMwHgi4TmLl97kHRWxaAGcRtl
5kHmL8Zko0/X2sU5IQCbsDDICSPD0N6P0WGBmESvNoOa25GLOcEcWPZY+5Lzx5zmqee3adqPyLWy
V8A32I6AyMpytX4zsRYAczYteiWS2g1Di+hYtrx7YclefqSMa7vnLYm1I+91eJTnXoRFdVUbif3p
V/CWP4+KP1ODinIKVc5ZyA3NR0usz14tnJDkrED1XKjgU3Lqjj84350lh24vrqqN7ZRXz7ER2gqF
yJXpdAaEU4upj1IJV3kFTgbBvCsPvSJd+w3dpXZQbC/RUdheKYnOPCRouBzEjVj5JgWOvFBx3j6l
CrVQGfPPV8U/r0/t27M+XjbSUvvWL7QuEYhvrNHK+wN7sgFE2Jy82l1HDvxPoEkf4v148sIKkSJ0
hY3PFlQ4I0+8eGee5rKZ4LiirgVvNWuNqgF0kkLkqZ+h77xbPny//PUsCBa6DegzZVDqzyW5B4oR
fvWrq+Oo9GsoPnrVDXkeeVK9u251e8hnYuEs0MaczJBgzwy2NDRBF4tUdrzAt6JzV4DkWv0PnMh+
NWElmAujr8FnHKz5eTcz33tQsHkDr2Df6bSrd+FlnMaiOzLb6ikjwRPehmdbamkhoEgwvgHrD1Vw
GKSTuFIenoiun9nJ8DZuuDEiY/dJjmKZo+ZZLLqEc6r0eGDkUJbumGJpKGcm/cUtmR1TDi96l9cW
bqMst8zZhOhfUOD+O99XAAFdiJvCIHpd1wF7oTE1dKJPJjPoSq9Buv5GccZFX4zABmsUA9W0GZI0
Xbu3ttBhLvphON9DODMUdDvHghan+Nh69D0CZ4TgKUNwwBRR3/9NFkDQXyHusnv635mwEkMBe9Nx
BL+GXnVGizrktjk2X/sIARQTR0fj+JEssIS0GnoOSdqYFCAe+PF9gIBwgvecoWshiHNXMUed0rcu
+dSkgXHvemaXEOGzGRr+iHangPSxKTcjBkd5ohqvRLVfmly5raUExEZdpSg1JrfufBu+H04DOAI6
b6HiCwnC1Cl62rWDzzxL6Rg87likGTUAcEw8biN/D/gOK36efTZFv2/jZbIpnS7KOXki/YZEAV2L
9Ny1AxJMgPd2mnYls6TDd7HsZX5BJV9exE6z77MAUBOXOfEglFTNk0TERxZyxxY7EG3pBFWEjfsb
EqZqyNE+9G3gsDj6CLIKchT0bvnVsaets/SXFaHQ2EpWi4nCOfQcS4FfJmYHtbHdq62PU3Tp8e7/
O3N7J4TBQXD2p17jlca74Pmu4RCvcHglMeObIlQNdEWogCjSwS+GIspVbOWLVHaejQ6ZARu4I5t7
v64vcaD0j1hHemqA5Bw8IGN1IR2cpGnaBg3TdLMfXl1QG3e7VAifkUuyKnaJzEaL1/EJyjY7ssqs
PUtKaOxrMbI9AjMwTs9GlUVDK3GfOyszNYaBRyGRc+uoBkfK/l3J5RFBFhyof6knZJLOBh7flUWh
YG14BxECjlSC7jDRXO6qkNBpSjsvy8kPRBy/SdiYm2HhYw3zcGiUi3Q1KC0zVcUnEvPcrfEnGzC5
tA7Mb2VlDoBHHb76utgx6fO/9WzcKro4+Fwi5oazxExN2lYFfjy4R4lUMol+7ecV4X/cejh8lPJL
YQ/BJbzNZecQWYMIZBf9NBpqOJ4j1bhYMfsTcQT6tu6RB0prF9vc/CtNvTArJlapLRq1/r2jibkF
O8vtpH7qwX9cnjSdHjiFzJ032FiDhir1KdR46EbD4anN9ZTJ8w1Ytf03uCBkxAaGp9kKoV5F2j03
KWhW+XJDzzpHSZbyjDZ9gayhmBi1o+YbVLmw7LGjmvQtyE/p4hu3NTXCaYLpfuMnvHwR6+rAZ7s5
u6y0J0wvdckeAh0hPZLbzhP6pkKHyVHlxG3vz9ZB3hYvUpKXZhH12Q9MHC5NJE7RD2rfWIqGb7RR
KmVFNh14XrmNpsWCKawCr9D92tP0r2nrlAPFnNmAep4YJDdinIc7cJVWg0MkG11fei6sHoIt4v7t
b4cyXAD/ylfJCwmVrmB14eKz4Wb8SUA/KuTXSi+pbtCymfgT6BKUvL9noKW4/qs7Mv4Qhh+nqvDU
Y3oSyYtum5AnACcpXjb04olfHfMVaZKnGkhTtD/aIkj1Fs/4wclCxtLu3gzt5UOD6Vz1+HpH6+kQ
NTzzla8zveWzxx7Y6LbvpRpQSM5+7jC3jHZDBnD0zLD0TdZxvFPKKsC5wVliPIa2+TM/MmghqJGP
NN7yd76ChTUQqF557mlYR9Y8cVhuWmCIpXpZDRXiD3H8ecC5HQ+RIXuIP3qj0RgL1CAkx9lm9UXI
WIE7l02weZCMwaNBl4Kik+8mO0fXtWTwme6PRIUmQzb00vJ588d1ERoE6dukgW/qFemTRPdV31Qi
tpdfgrp3boFqfIYnv5CV6GqEm6RB+Kk53QOPT5bvJX4DR8KvgID7vMmEijYduftZTagP4+UxmjGF
pPWsp9N2iBgecTx8sGk7iyruuhhg9MPK8qAyeurl7ZKTWwjFkLUjqJwEKekliyiCi96bOF9qWgOk
t84ogozDK4/8bDFS18ZvSozzjlUGoXp+pfblfU2NOWGfcKkHeQ+wwbsdpe8zNLEtHM15ZyLcn6z+
WcpdbCGQi/XXgeNDftg+nxWh+klkzzPNT6hb/2s6UDOz3FaTP2NAX3/coO/Dy37/k/Yos6Uz7orS
G8xFcrkYMuC8Vrn+a1C+osCb4fqe7xF4WaIo8sMICdcw8Zfx1qYjHUduw/a9Yo2SHUiabLfVjzs7
FJKpTyC0PfNBJxCvVWJOPiXvKwUD8tSifgk3keNs7jJH2bOuiWUdrO9K9dm88f2DNTZFKlEUNzLV
a3y2JkTUmTTItULVc6Z7h9Vb+j5OicnOqjcQvIvMjsPAxECVa4bjuxT+Dk9Ln05viHUI7EIELkiG
Hkm0RsChDJh1Vc/sX7nO23u+OD+lhgSG/9zXBqOww4KiXczmG2VOsKmyk7jCDDmTaJwGlhv6lT8l
bKkhSc4brFS0DLCCKEFDycOGVDplf4Njq3TswpE6UXfhfhUvjfK6IWd8rSh774y5dEInqkLDj/VF
VlmRk2srIQm2MmjhwENXHUyQ+pHo6CHpMQnJsIma6e/AxglNfrggsssk41MYZYDeuq5+3XvlDNsS
A8R6WR+GIVtGV8eo1QSvwwzjqRxMvaPdXFaE1uadZroT6qW3myXSXaMk3M5TSmhurI6+oVw4JUqj
9qA4401u7MGB/a5wcRUg067bZD0J2EiZ2Ae2bZxfc8qMVpYyZiP0uvCalAKInih+r9gU3nVkKXJO
ExptSILCOq5faic7AkjbQLljg7NKhYBZHY8YPaS5Eoh7k4JQy9Hk1ktbzH49d3JgFdXRdSLx/Xs8
YaOPl4V2SwNRnOO58cz1fJmbqqZlnjHU+B+4xDmcnvX1OJWbRCuvpayu2A21PDkJfUmesAEVKe5p
lKooXu3ft8o309/oSZ/cfL0FnVu8ZL8CEpvlvUN73DnoWF0DFcYkl5GHZR17Ofg7Bfe9q2URE1th
iuJ7wsRP/KLjQJPiGebb7N7S8fOi4EwMiR4VyFmuRG9QlscrvekBnA/eE4aYYjlcrRxqZtZy9qlg
GreFKhtxOeyLO2wzP0uKsALtkmiRwfDEHAgz6k8z7DGqmV2+e3/Picx+I+4KAJGJQ4wjulGbSDae
RSAnRW27K2kBRkOaQv5HuVKC8e9qK1oHtaHEECtQY3gGIr6sDIOrgV3ozp9rvQg52HdM3gCv5cUp
F+rZohWLPbJD2eAND+45PDMOeU32d/JfnBWw6ZJiaRIUVGr+hR8HgOV7q03MeqxugFxV/ZCpPOMj
ES8rrea8q9ioe7uoH1N4ENjuINCACG2mQmKNU9oO1Riruu+A5/TsvJM+QIYYpMc0CWszbYC+jz6p
lYjAAJ7eGBWi7X1svxNVux4BJ0tYzQAtNJYjYYZiKAgCQ0Kh5kq7YcRm2m+C9b2BnfIQhqb4G2QJ
HLYKL1SGH5+hNT4OcactqVuiVUa17n4OZyAxRETa98vCCcxTIKDghnK+rcbkM8bo9nBwhost1V19
GxFasgoiAItSdlgrjzPiO2NwjvnOaYYTXR2fbYkHSGGXxr3gLdY3sk4bnTpBECFi65uxIigWSS4i
YnY+nEHh9WfD3Z/+uQz+Wpc/XQ6Yp3VkeW2lyMTdVmufbaAQI0+zrietfwMKcBPrv7O+ar0ubBkJ
Z9zt/qMaQGumEMRY/dEdyck60GmlcU1CbQPjLtXCyWs4KyamHNp5XKuzqeQS9jOP3pEpWsmUkrHF
luaKsgbZyD8MlshxHay3a2iRdnYd+k+GEPtKQPfrU6f7owooPbMNS2LV5tjDpVdjOouuOVWbJmxq
4HbnJxMQSCZ8z5jNOaOBLmsrYNiwSFx4QhELEr55cnP0cR6H8dTOAAqhT/W6XdmiSIVPpe7E09cT
djQ1B/CA8Nqhp/xMzmT/DvvQhhi/jrCBv+n8KGw7qfGoaGFdiqSi/Cz5D15RW22ijtVzpjTqrXP5
kWxR9QQaQO9AxxWAy9X/p8WlheKa2o+NeXrSXvVl1slAlaMyXdGp8V5JOWQaCqRCKMVc9uC5T2zM
f0QN3mC6uzgU33JRZALLKhB8MXJykU8nX/ZzWVPhmVUA4TbUBh7ZXs+mKvnoYobUOBTkPw+RMKzc
/VKLsygt5NhsV82KrJU4Z2v+K8FYuYurG4E48i7VgRAfV1e1T03hMQGgMJTOb+m2MKAtJY3w7L8q
MsOIcXHKuypkoFRNRpM2gXcxahAqLEAgoWlvZKCvru8VB8xmIKhiIU90j+fkTePW7vcdXrY6mDHB
cvbRDjWEtznQbA9HxvA434Bp72Qr2SCpR22j+Y9srrWQgndfapvNYvkNy/KeOhBBCPAXBujNt4iz
4JRAKrWjyxBYxGKlbkt0X2oeq6x8VjfeXsZWBimuLhUlpdcokOqZtMq+rJp9bIuw+2unv1sX5p59
LQEnBB0qTDl1HJSjvFtW37qyhGPIfoQ3h06u7IJwT1YkPhEVUcUOee4KKQOIcLbfRGAZjhiAYji8
y5xVJ1wpMQbRmTDGzBSBx+0+TTWn6gHHjTyK+gLkY6t5TyedOQBpCFFzRBVwBonhbxfifaxLb/GI
Wo/VOyNU7ZfIYzJKLXUAmlh14PXPrjHrxSwOfCzZZ7v4vpZb6nTZT9XFJK4M6W/9VO3YMLpHZ5Ke
PFp6Q0giZOwuk0A6se1Rz6+zHk01Lm3Y9vI2beJVk32aJMY7OmYx/a/q0NQKWUUpRwFlMY1Cq0YB
JirOdInsZyobnOVNWU0QOAjDwzMwj88VcJLCURDyYVpuEfSgcgYJHEwrV3xdPeeFFwOAgbLpd0Lh
j8X26QES30uUREf6j9PsnW+G2CZW7Fo7ho9byTUcf+AW6FCLPKDOdznv/qUmyH/HJNsxwkmkimcO
3/3LhO6OnRA8Ot3ZmwFhlesADUkgnYZLkyHvxtYkt5Tnq+oLCgUm4hzF9Y4wDbzolPOi7X/nNYny
zdLzjpLDpIQ7OoB6iTsXHKejplzEUZiQKARsmvSN2t7jPTG0Xs3bJ4resBwPBnfvCgJq2lsywlKo
tgAhz6WVdx+x3ZO6IHQsVS0RcBFioEkwPrybLP5bsTzJsa/BlNgxDJbX/AuNgXUk3Pe0G9jFWAcf
zTMdc6otfwBP3mMJ2MUzwzmq9L2jdalyH9jdABDogtU2GWSMzjU3e1QGfeCSmN+zfOzQbiD6Qns3
ynoreCriah9YgwdURBK0rn+jDfPFkH4ORspKvxWwHlJpKI/KGZuglzHNW9uzQ3/1fkgFKlO9pQCE
p1aBjZzaCZGZO5NIWo8OvTA7nqHtxtF95RPQoPOZxSloMnObje2POJSNLZV/H4mJDv6nCgUVtm4P
5kTdSV/7KHQq7W/fJOIVpUcXX2CnZzgdWpowtLMaYsSNA1gqgrwIp46FAn3yaRndhbKUv5sjyV2V
mrntBjWdXHazHgvbzDIw5HQxt2wrTUjxZM93bKhcZx9T/mnOoH92r8mCiMILQel5YdQm4jyudhmv
bZiDzncDZSkYtTvdKc782PbJdNlLvgUofNF6vF3Si8ZqsmMh2INl21QCf0InHAAo6JaCom+0aj4A
pMcUi0zWGv1kfwsAvK13iYTbNRL0c+tc7IFuftP6+/yveCQBT6OelzvI97r7BZKFRN7umdeesQlR
XdmMC3quf1BVjwhFbj/MxlgsCufuSFkeMJvlNdM2bUYkJN+gLm1cfQTUHKVGUvimHZg1wijLBeJW
DFyqoYdUU9MWtAU9PIt8nxecQj9oaG6xTp+iLVRnBbKGSvCPj1iQSmvtzrxuR5KpGqGxX1fqVYhp
buIN1t/VynC3BpGFilFtN1TQOwzJXY4FbUsiTqsUnny1IjmQyBi0WYklgzNMrbrFUexFPtSTEBCQ
PCSTO92mBtKVS4bSeIsJGU8AKcO+Zz6ZNCc2oVlPMu4c8nWxry20WJdESxPcs0GoWY90iQguPSq1
DFUWSegLXMzJ90c3eXZsGrINXGdwY3EM7xvolaNZvwQ9xq+CohUstZeLfcLec12ulGLhgfGrr2V/
oZFp5zBgudJscJJqfsWb/RUPEoFf02bU5mLs4s2NdErhSBb43XF4KC4ADSFJnW59Sa71vOfGW89R
6wnvQ2xD0NWioLn2xf3qh9cMiqjZ9tdKuHlvl2GHXFzkrMxpOX+veRDH7LTPtiqMwcXWgZ6I3jic
BP+5xozJgMPnpLmEBPe+lP6qQick3nvTSedUVG6m1zhzlRhc0ihA15IIVWp1dG7ot3dCuswKnLt0
JwsM0nfER1qLvY1lKYVwIgOHniprsjDQTjSWXPtuGLSxqWeUj09ycM/x3b0fnyqjqj1wBf1F60Cc
FrhRZF+6dVgPdq3FumPq4csKlcxHDl4uf5y5vSpbBl2lAFQPhKK6zwGcPnvMXYI8fYF86VfiYALm
QZI8GBxRZSOBaS24C6XHPXIfldshSi7wdimlkgmvhzndoTFtJZSxwKiGZWhN07hLt2tAgb/SYkr/
8TxUUZD+ddMDf/inYeYBgheF7j5i6dU0qYvFvb4og/je9YkUXb2yqNTummfpaSxCffhH2Gp+v/mX
lcaqvPUzZ0W7Tj5ZHkfIIMMbiDkINcBkWHcdWCLIjjCAjwHKUwdUvHECvndyg5XyrZNK2fXMDPN7
/0IPz1dq0wkR0vb3Llc225hk9su16HVxaxEZu/HnhyJ356nwWmngJ7jlC52UySEdY/SKQVqAiFYv
lrhrrOIZI5a0PctVjnykbF2n/UGq2zi97fvA/BajjYpw7fd7ExALLGnnSET70NPju/VuQUUMPkQo
c3UPzcbvo7FY8morgy9y9gVqtlEpHF1OqvlJZWiSejcWIQbW/DV88sirzp8x3DyXjxl2DExHu/BR
NTT4/3/P8i+mR/YxvVlBqfALCArTmcGAq2kUY926p2flq1dUwhCSpEiHBGSVxOZV+AkrLIdAvieo
+m+R12mr+68etnV8wy+5oHwZ653UPGEvFRm7pI8dTwY9Cbg6SSg4Ozx18q0UedKSwWEihDlc6aGX
tIoJ+4r5Rb8A99/X9AwUswPaa3wumNP9RCbBuM6nZS89VHOoFFkkPoE+7xbmI+m4yXSI+vqRkwa9
Wz85Ml9AbovbWrwNBIiSwjjFIUCzStbYgLLqWw0Ovz2hVtaWUztgwgZzTM3/3joV/wVgd6XDqHr3
NR5dw2DEIZZHzjmx8iHdyMXky9WekWbmH51eP3WlD+K1rTlV6QQ1vd9oVN/Mio8m4CP8hDqsOPko
F7RLMTsAei9VBlLi4b6KCnOBjeZ2buXaZ/ezb4W7eroFOtv9xSOd944MQKMifj0wUk+MBbsDm/zH
VER4+efdNoPHSsZxYlfQsOUElcJGExv0Qsw9h2ab02v77E3ST/PwQYttP9qg9n0tVNMzxllhBI0h
JCs1XQ1jt1kxPq/UZu3wVK/9zTvIFF2KOv4RrAQWlV31qTRQiuu5GqhFSb++ML/+cG8CGO3RicJd
WDTqxCujQpIUYrhy5wwwlFjOSygzfdb+IfvB6u9q1Zs2zUCuEu/0MLZ/+hYs6BpuFJLAY9KsNlfa
EEGYZ6ZXq2EgLukufo1/c68BxEyoc8KIfqSpZ9IrLL3abyM7pK4xFCPRDkjmLyNwT4JkuLinBU/U
fyMhw6+JULx2VlcH6OhSXSFIKbtjDM+zTbr7dw3wkyJpfWq9sDP0JFHQTKd/OCuhFkt2+/PZrrNB
KLZOFrbmNFLh+MhrI343c9rFTaO4nJmRoNSGQVri6dADSeJnT2d82N80MPRripMzBGHPYGujYaRP
OKyZ51wc7oK5wAO4I11oMo7ykSPF9XIdxuHRy3XfwVxtInADTpSdi7cZPWUADmnjNZX1F40NXZzp
iU8nX2BrPFCVZVUyw31tkBiQ1iPaopGhDWIkyzgbXbBEIAmuBt17vIsHGe1mRrGDxGIWimuAFKYF
6zXdMVEnzdePNeVVWZn29zS4zpqOED/scgd54/2vtdUevb+8mQFvPVQYDuZvId0XrlXOJeo43S6p
//0m9xl9Oit7yHonvEuGV8COAw7TBj7JqyEzL2p6/p/8KXyv1u845Uv5F9fRuNVidepIA+vWZTwn
gXr4Bm9l3qJ4JsLM1dfag8TvtHlQYRQjMdAlnKFa4ttHQP2MUtJf3Ah4lbnEQ4g4V3r6dPedCg9l
RkfKeE5u4Li4E7GyK923gD9gf1epE1mxYP2q2cgy8xWG4JFTJmgtG6pV0HIurpE4FMwd9kuLHYGl
l2rwIDzquo5jWIWdNsg8I6rZU0qRhpMbqzK4BYE3MYYmTCBVODbV/TeY/fwBIxUDn8+JOzKdaslC
OLaeWl8r4DZ1n16Y5IKBBGCcKzh7D20/DThG3mEuUnx/triwpSE0EGurqJXpobYsL/ovIYZSAa+g
TPXYo2rDk5nsZPlhvF5CToRbKwRLvUmsFLM/cnffK6K4AS8HcZgSq44eyZwEigSg+CLsVjxu3RTh
Khh9TxljYmtG/T1O87gPJ1WzS2wlzvxfAZc3Ifqz/ShJIvrL/X9ccSRcy6TRDkaiKE/0VJCfBGdD
DIdne4J+/pjDjdUujIZc+DKcyydOSADqPcQ5MBADmDQHdyxPec2M4a4Ez2R9NrME16ka/ILnbRvM
PM56DOYpW6VgGAVrUHD8kQ0ZMN6mjYq6zRI/G0HH9AHySBQxj7O4RH3bLkU3EzTbw0qNx9p1rL2a
Q4Qp5XzTo80QMPB5NNcncln5EDdfGHzEBCgIUvYD+Od9675Qocn/S4EGZpWn3eyQt0b7aDHlw1gO
ElyTis0OB6+NzECqKm15fGhu2fej+XhhVGivyBLea6kZniVqBaAzAUbxcWu7d6Sb8fwYJGYHRQxp
9J3x3cOzd1wNJOhkvMCd3dDFI4IuVr9q3KAQlZSI1pDxYRrhyMYaIvfCzDe/mWaLFl9BinDCsfYa
IFu/tgy2WIOcgJRvS8VA3pO6AulCu541V3xpFnK+bPLy2AcTJ+fFxoDREW2QnijsIAgdQwtHqUJ5
HSRSaC68GATlky38Nn2ygY0coY+Bry1HWmT07PyoVl3XnszHrMI46Y0BHWv2c0yUo3vQVjPnfEDh
MrVSM0V4SwjACFrkhYb+o5WJtkbqKIm+a69KxNsx8Z+8f3R+WAZZZpMXNbuPPqhDp1jb0zEiNYXP
KL1thFU6meMeVaGP7lLDJR3pbl6ut8SGm7cBBsDPk5lTkU0lZLiL4OxD0tFWGGj4qoP/X6ooA85l
DLmKgaBdLOFfuSi9eWlosM9OU3bLLP5VELQLC++AJKkC9vnOedUfUPU1mKMPErb0UU2YaKgB1GQL
pWFlVgMob7K82hO1hgE0ekldFNJMjHeBvgxCqflJsuWLAVaqn3gtziTb5WfdLaCHA98ULN0BiCig
ZeBrrdWeywy8mmOr95cp/uIuy6Wxeg8+LBzpO2toyUNL4oFxdDUjAemghGMeb0PmJj54eATV/A45
LvNYFIZAUEXi8aSt43lVY/pkB0HW0TmsUYwV7tNtj8KKVXpCSiHmZFyh3lFGrufFCq48y3+xptXC
+5zuk1C63jfqnn1D/BsIYMHF+0MHFR6RM0XwAl1dQxWswjb926m2VIefv8FZUgaPaX+koQLBAmU/
jsW6PdtAm15SDwo1bxa7R7fTNgje7QB0idii62a6uCD6WXi/qN9ki/P0oX8V7y6reriTeTgnC8hH
+LV6yKS0pjHe8610C2UDdajGCUErcseJgQ7GAnP0eEsnXAJGQLphA85/pG68UKhJFbpG0RQSfs6x
nD/CRE7uZnyd08SY0lm7pWjmN2k3YDLr4r4DlAxYtDYuFIeBBpRzW1+qfmX3iREIGmW3bzqDbK4h
ZS5tpjVulZfkwJyGumO1vXWyafq4kzbuhVfqG918O3e/ps/CtDR9V2q7GI525lAxMgUAgTuIJrCh
AvyiLFSnbFCUQ0t1mBPaVyGU2Bx9+MGF8pgz5w8bzfZJgg4dmMiyKVU1CxUnMM4XFSuDHSN8Xc5X
HCf/W3ogmblhjnD+6iJ/bzYers974NpRvseDne+SG/kzTtfVmWwx3IJXCdXapctPzYaS5jUOUl4P
VltfXzAw1Pqj8YbDFr9Gmtto1q6rhmXm4Kad5tUgeeTqhR/fyyltx3D2W6ddgwLG/g1elfm/RZVA
46eDGmrjYgbfhJ2N9dFMZilTDAGOHSEL3UcdaaEeqkNcsJWcS6gYmLUGmWkiuBJZiRxfmnV72JHq
yNb59kNcfr/0kKV5IL+wlJQxWg//IAZWzuziYz/oUBwDqsK4rYdpj/DpaFiPlr0MCmJI4aYcGRzK
zbuuQ9UY6JlLHqFRLiLVs5EZ+94DFo/G1CcS9z+5HjsfU+D/SffpvQq5+7rVXAqJ2/JlXEOgu7at
Rb9xYsWqsqkhiepa26d3tyCHf2C+C8gi46sNEW1EO7lTBiTeFkVEQw0pTvs5VW6CLtS381yhv9cV
JkpSwJQGXxJaqhKshGUfIzJMnGA4BrKzqNiKMYTjxOP0UYIswWh1uIMYHXeFchpEPetZ9P/tJFX8
2sxNVwhkOs3BBh2ncRF6gWGZe5/5g7lJ80GsaSQxD/b3nONpGI9L+aB7KryRmu8htWRc/p7qosJb
5K4ASXQO7ulJAjTNWqh5EMCT983kr1OO/a1VafUQ3UJw9DfU8OVKMyZqsQ2IJNB2+SzMi1QXnwLU
Pl5q+KsvO2x3SujD5OMpE9BaXBpB8ZgRVySnzlbbh53PakjJouhw9ec3+4VzAUkLgi2CogKIMtdn
rIY/v/RSZn89znvxv/wsXNQ+s3WmNaLMNz/9RM6W7R47hxe3HG/PjcyU5V5NMgahcbmtwiexsA6j
NmpKfd0udf+DGXNUHvPl8VQVrsjUveZetn8ge5jgsqyuYB6hufh3PjLMopgJu0uWv20ZrjDgOoiN
rann8JRAMgiVJDRq+B43ehn3SNiNnKH+yNMIVfmLTdB5PhPLlVrv+0ruthxLszJ7TqvujX4n9JX8
Ryc0kmjObvhdQyeYHjqgC1FPHhmnI8TvKDqm+U1+4PprkU0JDVYQt8WJOT8XTHesxqCshvdkKwiA
sLl/XJwN+9le9LTUnEGhUQC3GHBY0tdVaodoyJC5ZiZTlrTr/rmlQ3xyGjHi8x9ajleKCxytlyUY
Aljj2AJCWTjKtCVnXTGRDBG8DZ1vAg0G8fAbKur4J63Bv7BkkunWsAs52oDixO6OLFn6S+D9SNfs
DFisINQ8TBqziSOTQIbmeM8AKuJYqxlkCk57NNlgx2UeuW9iGI4RzfZegF9KP1SqcIMXdty26Lk0
wjSvNiiVAaCd6SxJIvdet/aJQX1s92VCVyTg6pW+NqbDB86tWpWkOLJiZnwy4K987eqX4E3y4h8v
kXzmyf1MhlUc2lKuIxdh3204a2pPTjNRbAbGESBEyBLD8DmRPctNSFrEoq8LY4r2YL7XvCij/tVB
7dmfKVgfwz584kOSWTfFIua/z6N1HSxiBiOCF88y4Mqv4P2TnORhJHAe0YeSrYNksgvki7BRYyNu
9bb/7fz0T1BxrNG6pZdq0clZkK/2Pu8mk/myphVwhNQ5aNfdIPjK4909yKhmh2XL1TDx48586c5W
ln82M/Tleuf0ZFrYsYtCGyGE6d0X01cqMxOK0nd4g6E6kRdoKz1uKycYt5Hp2ZyIqgpyqeF/9tUs
+I4DpDb4iS8noxxV+SOZAtrkAEpHzOeaUVwDaBmzkD1o09zXWrme/XkCoQ4AxX4oFV/0eEmTXTYZ
S660NH9woWoFy5vZCpRpe5jT6R3dRlDcHVWIpjOB5oFFfn4WH4uYPOjMdCe9IMJD4iEVR1+g9+EV
KbZeoiYenXP0T0Qyx8qP2hk0Plfeil/3eWra574CqaHhLsk98my2aeW/cMnV2mpUb8TN8HaHhq1T
LKLeB4tgkph/eHvtZxFHHTBOZZO6eVyE6WJXaZ4zfuBM5juwjWZXMevwU/wMiB9qCWmcDAGbDtaR
jBvyITrT1BKj1CqTP5i+dAiWrXr+W2fef4kWZUoI/Qt/LCkclHET2TEXZuerIa0puXie16R1ErHJ
KOnHLmdpSIlOnWL0duMjoHicDeSIbFRqtzZkc09v0OS1DHpOteXQZQB0RWnZhOUeVL4eh30bFEpu
X8SDdGiyRUd3t43VxeeA38nrRI7U1N8EoVEABiteT2FbQVv9p0e9G5WY0cpRVKSNA2W8TBWNXeWZ
O1qJ6hfWl8YCJNq1Dwd++cj8SCzn0Bh4SkLydk1m5jeohk2YvhUwpP4lufjA2GaqQlvOMh/0lbL6
HC2LJIUS5UXhTRCsCpfr87ecE7C76Xpj4quZhJKWU8bmpvCP3v+UV2BvPvD5K2HEgsaKKGdORHoz
FoJs6l+Yk8UAgz67lzBBOuftAlpeCz+4Z3RtXLehpaKog8b3g+sxxFZE4YOiRK0wAth0L1HSsqN9
6qAIAFXzyAR46Lkep5xFBihY4zu6QraE9CSrko0OwxvfekjR6pKiaPXX3ExiTXHFr6YZzltryHJ2
9w2nUiZP0BY93tNnEf/zKrHY4BPSDzGUxKHdgdruu+ct3XnYlWD/OKXn/txFnGsWMt0KpvZgiu7R
8H5VsB02ipN/psLPwnsKPc9elhxIYn+lXPwBM69HQ9XiaSjH0sqAFwzUmdTfmgm5s+R/buBaJjrE
8T21q3rkGD9zTQXkLGAzbBgk0rv3Y2xFWq7Gm54Ye6G3uqswWjq3JZORs6RopkyFvYyQ3VcsMnua
plRv0OZTGR9CtZ6ZmhkqgifykkrEzQ0HNIAwT8Tqhi2lcFC+UdJil1xk16x1hIpEpe/wfjguFMK1
yxqGRqT3M1jx0C6jOWpVeHOP4Rp9MAM0qzkFk17wy62NfkzclMjDqp9vIDvlF37aNO9aVdZK2lkE
f4Wvmo5TY8+L2ITn6F93nzKHP8kP5apZdA/VJ7PapITH5eG0ee3ucwfBvKBtyRe+xYjCJIMrCJmk
5LtOhUsGl/UpB0Bl+iZ6Eo38aXW2KUwa+dS5zMQu/ftcwWd6C7s4V5GSY3U8n0KzaKAS/kAiDZKF
rtWPGy7cssNptmUfQ/pzx+SD53+oi4UhNGW57qJGkFbhg+Zln2nxVwWU578A+DXp7+QZHul3WZXY
LQv0TazykL2VgD+S7NMu0/nm26kO+ivZiE4af4pme40PN5pxVD8nDj7l6XQ9ck7LSi4jTd21REGa
QYaWETgwUzmWOllx7YxEngu5DDrIRpWr3U68cKTPlw3c1wmA6con3AvKMQ9djtlbYuHS6OKEnTPk
nZ99TmF/oFlTTns+6rmcIhk1mNp2UQPjG9LfZXEnxPK3IoTrH7DG2qBRtBtnkLb2EWFNCaApQkp8
FE5lrFDT/ZoiiEfzZcp6QtipkXSHS4E3nPPAcESHBZvXZXQZ6YU0JsD6h5fPceEmB7eW5r72tr5H
UakJrygB/wZ5KihPhTsgVIXXnz+wRQuAIIxeHK+e7BPWLyQrcK8xB/3QNX/eXG1aqimgeqE02bnN
yAp4si3UB7fdKb+dlvshMLRAvF6p/2jf3M5vLhAeD8PpBHq3Pelt7ogBpl85HNf0m6Sqa/AUKx3s
EOBP39cJLkfrp0/nnk/k/GxDK7Y3z5gena/SHhiBGX+rkCktkZUmMWorZFGmVoByfxH3SNaIxxRG
yToWLXq0/noFEOlw29toij3Rz6uvcfR7maPgLGIK0jUibdxHpJZmPYhk4g00HL7sRzXMkLBqWwQs
KxrTXMYduucvYi6Asc01YN4Qg5gOSgXfWqB3wlwmKm8O1hyAFKeqG+PVSAACWI5eEu1CNejNS+iC
qy3tBj152oxCx3KQI+RgdswhJtO5eioOE4VEV0zWjlWHiVbjEYVfuj6QfxO5OrmqNQGnY3ht9o+B
f0FL4uuCKBkK8jTRozIf5M1fuGNZCt3BGPsHdOQVISz/oNcf/LYKpRQh5/QDYrKLew9ofW9K06CG
eY391ZOivNVN0GmL7fBVV3Utn8AeYZuARLsn7MEdbvJJTd94LfMhXGi62Ozm4nXuXknFw96qeJ0c
G7Aq/GOP+S0whVnYDRsjWByinidFCDp94M5U+t7+qiivMoX9dgE45UzLfR/8MHPs6kY2+EQ2z23Q
ziQsjtaoD6mezXBqcdVqHz/fxjx4URZdasaeokgP63novryI4Xi6kdnyew6dTDaBigi6GkbSOuZW
nKBBuqNCVJpvf8L8XkalKyD5WGVUduIP3duiz/HBhtufEFignHnuffv1eSonC/NdGSMTzsPawphh
IP67vbgPCmBX9Tg2gbZ+LBpGvh5WJj4Mx5vpscU18UPEIb4ZZG7YQ/EgfNP2+66PjASxGMtsAFnY
QvO6dajBBV3/wCjXKaEO8jMNbt6ylRn9DISIHpuAhnTFQjAsHp0mVQOu6JaXEXF49PWA15Y3TnUh
8y88kBfD7yPMjXtbiIxMcJ1ucCavHVfYlb5h7zlGop73U7iWUlMhrJC0sGAtRDK5zgtRUZAcF0/x
Ik3Dtc2lbsW+wtyxpfOp0yxSzEMtUY+0DAsnXWrGLL/GtEL9tfzSn2kYm3dI6bwHahQ10QK+wGqn
4ilOS2wNMEA0eEmlr81yYq87i/Klmw10jeI0Dvh0FqRMmpTjOT+DXzc8oRsFI1RKM5G0d72ThX+f
y4asLczUWlAJ62mN5bLOauMtX0oQ8pV7RTBK8tKD9GgIsUADZCpGAb1Y9btLYb3rc40eMMJ3Ub4s
76a7UnXuxUnQhm4ioVG3CDDmpVTphIFiGyg55KYmAPHmyzL52LcDH86mNVsn9m7m3NcJ+gMnzOSw
AIPScO3mLiCNG3Qoe4G4rp7l5RYlxGJHYNliDo9QTkKNy/PcJYicNDhQ7E0muhOsGIpD9T704//w
yH06RdsRuod01tZP1AghKqpG3JVOLA4axLt5ddG6nS05oE/X/FPRtkKdC18pioljxQnnRbUxKB92
J0oT7hnsnLK4HnM3bVHeRWqFshIZDPNVYJ8aISCMrckd5wFMqWLKsW40Zwstz58ZrQGdz5p/SaHo
A92aryZl6IlWSO7Iwt8Uv9MRPPJV/L/iLFDSbqQ9S7D+penRUvX5jzr9gUq747gFotaJclao98Pf
fX/CFcqLLxffMNq5rOwClNMyW6+kJyLMAGHS0O7uyDbvlBm5BlNK0FSt90jsgT2QzKz/ErXm7J22
PHLAPILibkSfhfgLvQ9u1yX+qkDmTrNgp9rLMl4vMipTmCE4JBwqh9CgWFPgUN1mzIuetVKtwiid
4a9ZcqufaIM5Bb0uKjjZ21arTeg1146FZcTSTAHfirjU0EHkdqOe6GQv2qnhJEXD04E94hjYUqTV
Mpnte+dq+5ARwSHPLEEoyzyZPGdYzHpF3mLI3qARm4woJaiyrnRw8vvcxS2ORxUnRuyAAQdeMtJ+
sKyL9WVacUD7XMzZwhVr96m0s5GiAE5F7CfsvHfakAiLgpqHU6lN4Ss7NqVMXtAsC9m1MWzGf93s
B9jJwdX7yls5rkjNdn9oOyQmKbG5IyDacFTpu1OmbiDmaKxzCZD4pu57E43+FcVGNtxkXh7talCg
giYyqGyzc5JMeIq9JXCbWlMi0VDxgI4sn08BiCozpU+K5FaaykKPWe2RX2jF+r2u/igwxMY43cLu
8JO05TMSFI9GjR5Sjtwh5x5a2FoVaiZRoiJZUJqOC8494lNpmaTSCWdnnhd7Nkg7esbAgCiqLl1W
Wh0wnP06P2rgv0OHPcQ9fnuQH1eRh9SjdVyglqY6hH+RmgDzA2DfzcNE7NK9/ZUj4Pco6nF0DlmG
uEiCEWTVAk+zeqQofNnxQSandwd/JvRPv+tpGqPyaOVMn4lzuxJj5St7pTmDIzhGZ7Q8Z/Y6KxI6
t5NwrYCHmIdLiPtgfiqiFCqFTlUgVZcOtZLf6TJjU2Usx35Tp0wEnImeDhHwxnQ/DsdQTPaQ3ZbJ
SczY1LwZwvTa2XYVxUxGZm6zEUxI/5xS/f28yauMlt0zFasZb+xvAd//Ep/U/pczXDX6QBRKwj+J
by1GCyMRadXWFp1JgB3hs1q9Q/cqRMT13LazsXykCyUkdluAjKOTyIuXlXogHIUtYwjalWBaKI9E
AG5xpKwAkr5cH1Y3fQQBdV+tHa4MD8fuPOVJM+JuVxxX1bOljBxlvp3Kc7gZbeF3hCTg4b8T0MAr
TIpZcWgZozYfc/agYFNV+aoy1YHJ+LVMbCga4QYI4Bm5SmrPq6GfsV+lGN6CXPPD5BUQ1oG0YHE5
kQBQxH+qOdPBbnk88hmELC6eplaK8+Zw4VN5ejcKoEKoqtTmbeYEIwgkrwunGawdofpGV5xOqGaF
eC42g0LoCN6x5hmTyMAgBvW7YIrNmU/GkLrlPeSCHt3mSOOtYt32VypCijWjyYfU/pBGtW9ALKxW
RCuK3AlE4nlqL2rpuzIRcpoOVfKTfY9UPCom4TF8u0AB3ZhnISFG7fdstWa5CyrW2wbvX3tomEaD
6N7YRjCASSXd7NhpG2OvXxa2fU4Z+UAcsaUPdjifIpMbkZNJukHHdEaO2I7qzD/tZy0YXOa7DVf8
iLZJ1OASGq4OlOf3N3lAJ6y4uujTi4RHUFMjt8IvVxcYysvpcbTMpOihXNgys2P0DkYgqnh6Wu8q
BpjvZxGjtZ6Wsg+PddEfDGfStFjtj2+8csRFV0j1ewCtKp20I3oZMygeAiPw9/s5laf2NqFndJgL
KgcWoNIjYWaFEX/BNOSWRoDDc6krgGDV2d8YfAOhnuwDaeTMfZpAZJ5gfcdHKKEOfJrqhJTw+m88
p1CPTCHIGLVZHrsbQkq/1kABHB5owlRG8Uz3KCZDaeYOeKorFLHy7yJYpDbO/LSaGzZJ7jboAwnH
mSwKdh2c8IkFtlR81z9SFJ3bBO81sGir4zT8JN8T4hYRiOJU8l16GGkyr2OeeMh3WKA7bL90RbJZ
Y5ZYfzLXQi4hkEMWO+r9diHgZejELefBg+0xbul8DvtDWn5HrO4B9IWQJfm/mEhzbtgz/bUNE8A0
1Q5kw+CukEHZEeCtxAznkMAkq8a5HeNtJHdVspGOoRgoDJLWJTHP0kM7wPQmcKyu5dv3y7renkuL
WGYORxJMjSnVRLxtvtV9W6/kNoT1qp3KOO9+mtLd9jNVm0D46rQj//lihuYlIiDXgelk0mxlQJlz
/nJ1etwfN2K3XX2toAJCqM2bgN6cQ7OWpfDgS4ET++eLN96kqFHSBdOIsMb6R5EH+YZKp64YJTW+
i+n6Qt29HKAMewtrW0OCUFhpryS4t+F0OfYxOgd34MVE7yyAtBoT1Lue3SHD77a8pdtCRlcmBP/a
Uo4OBUIgzO8/wESqKXOwtmUWdZOqHo8kLAhYkKALovuvZoqpHnZlhcaUm6tjyzC9rdfdLLFgwbLR
o5nBsg/+UcTI9MnwF8BhI7OY4kqnFZOZ8EX+2Nshn464JQ43bls2EdEIECKGmh/vYYFsDLt30khA
1n06TipxDB1lBBQEJQ5nC/JCLnftEeQASpXa/f74SllV67GTlXERFY9/1u9M0GM6G3yVA0ZABk1Y
XO9TxqShxleV9Wn1cfGQXwQfacCCf5l4j8zTizQuBJNQrozo6ENVGtSS006gqUSGU1rXydkKMVXN
KCBX4vjtOs+bfaAgccBI1M0N9jCQZZr6ydHwB7BpryjWlCDk9kvWT0NIZhJ4EQW1FLBZVg8/O+l3
TJqIA2y3x3J1tVhp+io6uiUBw/YvxtWHWminSaT2yocVi4o8ggRsudA/8evTrdd+Ql53vZkIUfvb
bcRCKjCoh1PWY4wHf3zJJICB+6i/TJr7SI0g9Qi7z9imrQ+He0hMOWbp73GfrkQDhUP915Surgwk
A0/5vPl9NLH68eFCz10xiMyPP1Bl4iZEjTRf934ivxdNQfN+WO/eTi6RSsZEthqd4Dz9Eifh2R1l
jUTBWoA59s+tj2WC/r04nqGiSnR5o6cULOyE2nZpVjjKqEdPbzC7igFSFOmuwWYkjT8EcC3q51TU
wALn3yIjRF/CPzURuke1X9gJ+5OmFcDiMOit2gSvLc/fcdiPCooTQ5pCi9NKca8KMV5qGSAM5jps
tKNGLvv+GDVyVz4KCVeOwTfNseKAltLUJXHnEt4zQJDbNPaxWer5LcUii1yVE0i8jwaqyKMYrFy+
vMCS7KR88T+M96InQLPjyCo/CtDhWsdio7v+psCOkbaOz7d0FxzR83ZyRFWEqgtL/sSKDUI+8VQf
czIMIO2D7wDd+cGd5DNLlZYxO/QvinRzyW/LTpd872YKYziI+WvZfdZ/RhByq+6ui8qEs1qySrwU
luYilpRVm4V9SWrz9MnTYkX45O4Y4eOw/4sJTGgjUXZgr03Ye1uXZAQya0dzEFXpBDKK9oizh8a3
2RrWt3W8OsuiB5VkKG/z+693lhA/Tbw9R5IMoo5uQLcealvNB3RrHVaKLnS9JLAAzMf6V5if+y3I
gXcNEq+oq3BEYgu7Ra4YW4/bxrpMaAuxHOeD9LY3T7fOYOWKkIO7DzlCTMsfU+ROoFrvRyZD/iuZ
KVb/MWaUZH0/sCCMzpqfnCZoUl2b0pRLcql1kxv82Hw1DtveTQG13fLpwVKPh5FTd8FSpUxHhnx8
Fi6G0s+HFG7hy08cuY32enTPO7QHWRpB2Dpakr8fqTB0O95khXXjuBtRfm2VPDjqdlCdeVgIuuV7
mbJM/4roBCi5wVmQKhbvkNz+QEwlh1HsjwprxYCmSukUKUou63Fm5yfjNvhIZhw4y9/EKfGp/z5e
Dbyda7SIooCn0iFjir7k0FAn7OtsjGOBXro5F1WLr+oSJ3isXDovWucDBjdY26hM+NPC/BV5xxQR
FVpJ5d4wiIbB4c5ZMUgJGfwhQLSa9IH75JXDFX0NlsQFuQ+oUZXELRvO6OgAEQYbXsKsSUT09Rmv
lzAQE//Wy9d5VizeBkg69XH9dl+Q+YwAHpIYcScz1hjhXxwTUnzug7va7QodZKX5DovrzF6OwF7G
cZ+DJbh37Er6GKgNdmznDINRQv1/W24ARpnFG2pCa27GtpIMOUVfvXSnnyRBtVjdciLE8e1Lkpfz
L3hqof6pmhMijff5j5KUOEAuv0LqdO8gRWKZgbRQSAhJ8w+pnarvRsKYn+yFFV705NJF9Zp29+hi
iKygXjksPGBzDSwDBIYhjkitCyiQq6+S0D3X9tlWmfeu7xdk5eAtvI/Ka9EBVTkY4cmTadAqOVE7
KxxYV1uR1xx6wFWV4haQ4vX8p4isp1aXynd4hYkfYgcp9kTo5N6ZNZuehdBVLbpidlh+dOS9PlfK
3Er2CdIqeSk+FTO2wbDqpKCCI/TLr/Nc4OGAO08NY9/jILiuzyy/7kXWRDW/lXR6/1gkCqjljqP9
dCU49MFe2+JSCYu5pByZxUH4f1IURt/ygZ4mF2ow4weYKkjbhZRw4tsitKVTFRa7EAgUNzd3V1OD
fyFK9Uoh+2FKQdJQzQ6hsMHMYd4YXnwzjmBLJrfOuckU4dLMk7WbWPfnbRgBbbHnLV6qp2faGAly
x0eajIQJnlYtJnjb/h3SBLr8kqm3Gcz/xYnKL/UxAcxyENLo6itRrQX1FLnGgFU02ObgY/vtBYrh
vnv0OzibBElqL0YdrCZwhWfRx1qkmZdEFQ/xK8n6d7pSrADSmOLLdOmBV1jR6dvE7+BoW+4Eixau
zjiLbEGCPhXHnxseyZw7LU4bm9HlcXUKqulcXG20AphYcWKVdOGIGPuhiiSeGtqIAldaiBv/dpmx
iPS62S6T6s0S+QNePKtimf/nGJ2PrgiqZLTMs0RwFo5vUMhpa0/FyM6jHn8W1kybgGTIQrV1ZrrZ
C1RBigZSU5/qECw8xyY2+jdW+uRIP6zzI+q7H3LurBTYo72KavAnlovsnT1FGPBze8e6k5Nbtnb3
9jUUjLko2UEZKJjXPIwmH13//CSJxd99aAEytCqNyOXKcd7QngeCx03UM/TW8VPYJtXXBGlxM62s
S84jhDNYF/bz8lEOonx23X3VORkBjdY4FK4fjYzJFI5WbQRk4puyF7FzkBclf9CvE6VwO1tsSz9x
LWGsFMn3WtdOCfnL5Ip1SKxw9yxfXYuygG9C2HQb5fjYjM6BICyp/OudzJl2EeknRdAMEMGBM+fp
l+lNZ+hKoMsooFMkaSto7ZWIwuKlwo0tZAJkgvxBBxtrkz1hl2U+OF94prUyQBkWFA4twvD5JoCb
hOX9ta/ve46WmYTYSPNCSOjjPJQE4fqkOjvw/odKpZM4CPNnQ8ylORLnebaR4uew5DEiIk8HCWVI
lWDZs8E3CIsLyu506Q+xlVt+JQ8XDFdxOvWjDS7J7Z9VrJBTurcP65PL40rZgzqjJDser1PMraEF
51sc1uVf0iumwwIJ9c9wysQuvNulYDCjs0Jh0F7fKg3bWjypkLycE3+593JzaiBq0kNwpSKpi30z
rZcbYxDLUJM7h+hOWNoVT+3u5ICedn5L+wt8emEIqVoOa82u7svGaWDiQl0hxUhw3ro48IF5NdQ1
aql+YxjKTY3MFZgzkvn4o/KGbtBfy4xZpUAZXVr2RkUH7ITvqlS3zGOcEx34jxyI5clnr7woRWt4
ccxx4LR8cscfPNDv6jZ7HYhqIkvCaTQcT2G10w66J+OplQAKMJ9P+GkAQ14KwBcQpb2auI4Uz/Nb
4MlVVf5aA6h66fVvPq1/cSiKwuD/RIqRjkrN8eqYJFWWvMtOtaEcUJpUPsFhVgT2ADGN2NdPeQMT
hhCZ/omnB2sGimYAS+jc78JSL1nTCBqYY25hxTNxkAWuGMv5ht12+LjjaCzn4cdTKeFDE9JIaARt
D3Q4MlqH4/U1c96Bk/ztQ5/b4NFjE7d6Ip4asuk3Q8HQ5cC9wcN1uYi8luXzhtx2gheJhNfFA1Uk
lV9qbN3cVpLS4Izrbbj7SMcqoAjGSPbSQJ6FSHDgX7GeS4ztbumYRVa3XF6PRfpI+moaOpk+90h7
DPxSY6C90nIJCcwRnGolDEZGxkDxqtdsaatIi4TlqTupUt+P1gYve7MPknfI/N+P7LdVtVxjj+9r
SYaE2QznI0Zx81vbavprg8yzFhlvKljh2E5L9JOMGcOhfAqNSNJkzgs0a2wWP9ATQ0IWrxrhI9Pf
iWNww9oZA2IOvqaVx1cxPlAoNkXn8yNMgWHQ7AtURZKH3niroD+WrfH8G0D4JT4AIT0XJuerj9X7
x8RONijEIu0th4ggDgNWb82oBcpuxH8SbBamdBFRLchYwdhHiH6EV0aSPLNkbdJLKd4no8z9/EFM
nZxgicnnsAA1YEcp0Cq5D/rrEjOap0zuDntU0V3XQU+ZLX7n/Bq0+znDILGqjfcYxHMyN7nOBwnN
qg6/lDSOgzyawkSzaK7Gt5CfKxB6T7j7/ejsQtaWaLEGvZ+10w2fQFEriX+kg9rV5iXZYfv98fLa
Dk7VO539ZCIrEQ/nTTiRRqs7WlgfnhDS/INsRlzkLQApIZBG2535WPS1s0mEhkBlNrOY7OMndbNr
sWQuOM0bDaX5T0iTKQrI5DGHljD8Ys0MbAmJQiFXprzo5rUg36iMun0S7WIW0AnLSEPVujQuXfIL
CuDa0Hj7RZolpiNO4tLI1iM1gWzgi/+biwAdeyLs9cz2dcWwQbcxp8ggvNzPKroV4mlHPjG9nAIY
4qFMPHJ9aGD8HiXkty6JpZznwPR5O34sd2EylF35BbfjgbwdkGwB60QrJNA6OnSRubdDc0mhu4Hw
KvR7w9tmRtT50TepWACgx1ROQ9HL/dIRLvMZ0WMGr8cSfq0dOiBvKcvSFg/S/gOSXL8UJFIZELyI
HUlJgi4lPNzL0ipN54X3VxMO9Tq48O2GxVDJwlIQjFHyP5HQW+3EEqpBV3X0kUeGAz9WzQDsqHQL
AekRIAAxX1BQnQVPk4nzJGZxgRkVSbu5vTICCvbwRGfCoWPx17grDUPOZej1ecfD5Tzt5DvQy4Wp
eAUyJcm/LKLE3qttV+AYHUqV9dCWbf/5Gp4ef/3AaiZ8EB8my8V8OIzFUC/vhz5mcNm1yL1Q/Aud
Y+4xwo6Jesf3islhQKY1bl9X5YXD3mkuH8B81DaFSFkmgRNcJlHg8lnntAkPSyFp5TQFJIhnph/M
FzPgVWwBFMMOD2bR1MhoU2Wn1Czx8mbg4IbAgTfyvmw8AuivKLwq9/ZFjTGyMeIdfxJVXf5KFYic
x2crKvFjswJFuRK6EoUQEx39vQAQ4WdFt5iW061BVRRud/zeBKtSXV9TKak8OmxxGyeikJrr7lZk
hs1GM3MV4Fa5jDH0XP4s1hc7Cwh/qwJ4Nj6RUXyuZABpJ2GYm+Kn57VnQ/W+c2DR2WuvfrZZcwUX
zrv7oQ3lwPVOo4H2pVc/VjKtaiwrbHVsG0YwoOtX5vUr83q9G7zL9gEYFQjwn0d6kRI11v1Ajt/f
U1VkQnUB4as2j043l+dS3onmhVWz+SFV9o7tkY04hCIZokRWj3EHORaVEJu7HJ7wLbAKs3FJeEn0
ZAVpJT6VATGZ4YmKFSJc+uN27uqtzNA5M5rtG2ZNqa0DWRb5Psu0OuwXRsOX9DPN8lw2av8QBUIq
1juka4+0t4lGB48yBKwjGykw6YWzfM5uXz82CIdqQEPLMrBn6xDRMd1IspX+wuw02empqWcpDPDl
VU3LqBo1pC1Ub7rM6XhkLL0EcIbsJ3LKPfeEIoMfaoB2cxXkLaxydPvuPyl3pfkUNVMit5X8PpE/
cyU88cX9f2mpNyZA0+JCGqYfjP3pfkUTFBFgtCx3A5OrPWV2cXg8JFcz1qKDQTlwaPlilM6W4C/P
KFbk8Ei+n2i0Nftckm6L7rGOjfox+8UOiNLEix0RW9JdFu8MwCaV44ghPSqvhq2gAev2Y8dNNCHu
Wyd1nsLXpSuTvxH0mQVK2OwhD3ozchsxUsbJPMsDPaT7W6X4ZNsipFDIrxA2SqwhESyLOdfOoFxW
5iXlRaQkjQndXcS/GdSNzJo844sLaI1sP2wGKfW7N05VJL3LVsyaRidEv98KuOaepmZJ2C+75VE5
xqbMbzSe6UCl8PGrEB+cYugoPmQ/Dq6nzbPAxxSFH9MphQ/fNVvDm6XbR4JwgIfCI7uCfZi6ZUjE
Wb1588FVeeT3Gwo5wqqMCmSQY27NrtOvuy1GqpOx8YbGg9mCHmoKXgb8aKgdAprGIdIjPPoq3pzP
+5vbPWMUPVH4IZg+AniFOj7LQogDvw9254xn4wMcncvct8CKTDHhsxPwH6Jalfawk/9TmKoS/1vH
PuCcILzZgIIvy4/jPZD52Nz1ViX1elCLxs/DE6VYKAkQEawVWH+UM1PxeGwvcirEqoGHPEKo8sWB
NVeITJPxyAkOIL1XXIRavYOCXZHrgTHjwyNXR95o0EpjZByS7opO+VI+Zj+50au4dZbCujcqVL0y
v5lKDbRj+zjE4d+v+8pAyZhFQIEMD/tq6NlAgMNv7iu1K2cRdNccYPklHMZRmNuQLiaWNX85dI6Q
xUWBj0yupHGe5foKdoo9D283nnwowe3aHm8gN+LbVgoRNynHUTgoddkQNGKuwnoQPq2Br6XT+P/W
1gdd2KbBY90E/55iLpb5C8uXWXYGSX6dIsCx1/pVhbjCbTxR4NZ3DPvDiooFAqoaGLl5zTS0q+D2
IcAtPE1pUMVlFIT6fQNiu3SQxtSxjpMXEKFl3yvA7YPXicFyIBWoH8PD2VMt6NN3XZDIsVMsy4dO
z2rS1vxZ8JqA8anuLbwMspQ8o2WIu7voTn5RerthX+2gVM0MgS8eKPr/ZCklNKRPFeJJV/jZnsxf
KAizvxnesekHAZutSCLqnvKhQTrlq3r4yv5q+aUDHiLeJTKWhxwnsr8bXRSGP7oNDL9ZTTgzbb6D
jmrhmUufOZM0l31PotjAeznPgsaiaGpsag9+tjuxlPYylP+0CICyN1CMuq2lOHEPq4fl+wc0Kn7U
UUNOk959CltTsk2944YR3KCpqyKj8jJR5GWyAoccvdjB9Lk6LFgSN7nfLx5ZjmZVRRpP5O82GPXi
JEEg7Xe3JZtDLb9W+e9ksi3UIwudiG7I7o8M+voMdlo//M1OgTBlaQZV24Xvu5dvxDU+PMrft6vb
anRcOX8xr6wgayDbhZCq+8PHACQUasW3sIehI5ScAaKxYWO3hsrZLQmuW4mpt/dxIqJyYpULx4Tj
hEbxg6u+zKGGtIMgndLgRQPY+JSD4jFuTKCemNsjweNBtfKU+Qep22f5coUjYNFP1lSO/4gPAZPn
2XYpARjEgclErElE/CdFPjZurCbYxGjJ0xiexN8BhtYpA5Kn7pyW58eEQzw1UK7P/V/ygtNmi5Y8
Kn0sZOWzFc/YRYEr854lpacIdldalR52GvtI5+CPIm+wB8k2oGHf/ruie5FYnvd+drTeCj3BvoLX
l0M8dsdUBG45+k9B2nPRrznR+8U1Bvi33TQmo5GvWf0XLRK8MTLZNe8erQ2KMI57Wk0SORrYXLH6
ApkaSojo6NtPvQReCNWl/lOyfJmFPZHwvljvCv6T653GdsB2brtXfiYvi+iLTNrmHCPpAVKPc0K1
8iwlasvb0Xe1mCOi/2SNgcCONVAsMj5/XLm1o1hTrz4sPk29CS4atPqbS5sR+wyAZrHH2PVsMr7E
844/Oc00GbS9DuRDzA3PaYOOsmSO42ymAEWg/0orO0OiaLkghpsenVMEvS7nJV+gbsIPqwI6Fxgz
ffakqrbzpYbz6aOaHF8VmTomKw5SVuPG2BBMpPzgs4p0uubYAzt2TzzkT66QchyxovM0YZL8YbAI
rhLmYYfW4r1RAgsKlLCo2ReHCBwjNIRzN7HgqcgDPODdg9RVXfRX7mJa4xMByOawESebMEheIpLr
lYgcsZ0SzgapSHInU6Uuzx58WJ7EzVHi/sSyBC12V8QfedCUeqDhu1oz79X7ckRKJ/cHOy0kcJhL
qJ/WbR5rc58w+5YzgIAObaxV9ajCdxT74aJhSfxri9+hEdxx96m4kwWKh91iDdPyhQsruUa5VY5T
X0QevGjqrJi7XCs1ulSZYFxrxq4fiGQphWHACmiVY7GiwK/99nDi+g5k1IT/Tdq7HdqdUGQlWkwI
hYzEVm4fe1h9SkHRejYf7HPThdt+lihdDdM6RfGD/H8k+0OQZV8/H3xofz4zy9pVIUA9ISmn/3tR
set/T/cSxIYiFEuXV4so3w+VUtuECOqmw30wQBbFdPfXO7WF78nrYnQy5JbhrQNgkfqg3neXDk1I
4V3DqvemWtBB0pvSCLrkJfGt5g3kLT8gr16mlG67e7V/i1hh6JtZIjwrT49BEaKNjQHLB3QSY/bP
1jG/RCLXddJrWJmHeKOUNlhItHPkOL1pGlhmCXLB2mU+xSaeCopZAn+pRcr8GGeW9fzk7jOvHZzz
MLdFgrfItzdJhLLBqN2mcc+bOZ92jo1s0DS5YOLtklSWhFQNxMoErdrRVhmldqqLvCe7kd1BvKtY
LTzMzEkqxhmpr7uTh9KNDeMMxxjpkaxHi6jfimxoMktlKFJCsGWvHglBqEY/nVvnHJy6P7Leadaw
+9mEd+ocHMhtNBUjBA6MYwunruadWvrPHWMUbKgWNgT/k+VE8fYdfXdsiYrixnxpR1ae+u6LWdS8
VwkV1OqygEQDQvvShWzE/FNAUaRs+zHC/JbRKnTlJg/BfXyWIMgbXD6YzUy1tV/Huonme55JrQqd
DF/CMYS66/OqIwplpD1hWrY/suKt9RWvh8+oyPjalhwD3Zo8J8486hVCG4QJuCOkgergoMhJ21XG
+BuZ0H4dU5DEGSx2uavhvZrk7cnPpH0ccRoCoYmEleixJQpSlS0RcEWOYi7gjlvL9MjMmyYDhsQK
/uD5lHDjpZdQb+9/S5pn6QKWyfv+Am3uVcP4jw7zaFdijythUnr+OeaxgNT/B/6wNeBSeKGxiItS
D6Nf1XdC5Deyj/94gUwwGPaGdZiCGPi5yMRAZ9k5PJLqQydRlIelVfr3Mtzzd4UCBw2sZetqbs3k
qVroXUKsCyvx9RiOtrE9t1rcODsijBUwcaKghqODEU4XA+Jk6mBpuApqzOp8XhYnfryOKW8M6nSP
2TVSHEyqezeAQKNVld0Ln7n15jrs/DS/J0Smi+PA9r93HWAq/ep+Uppms18/LDgtK7ZAiK9fXmbA
K/Zp2J8G8jje96+s5Yqk+oDARGfNYBvocSS9GO8Cn7WTr/8W5YB16k/Bi2ZnBbQ2eIePKklhfxLq
+13WSh86DD/2od2yMblzX/aR3bgjRpurkz3KWVqLVKK4TZjJMxDHancygEF8X3VUNLbYaxzVU8+Z
LqaK3Mpm1jNx/lH9waiZwbObannfKVn21V+pD9lyqU3vU8L0Q8l+ocHaZum22xmtm9q37k56cAM+
pPQa7eAjmODuyenLR8BVfJccaD1rsdXfXn9CvSzS9nemvLBQQfhEDnaDRxe6qLhSEJqhd/AWb1K0
mEuj0VvipPxUW9u+YwCrH+4FjMPWsm5S2sy2a35I+UnyskUOZQwkJc/+/hA9BP3EVWT7YNIZ3xPc
OYxndCmt4ywmReP+kdCaZ4nQM3oCstz2BZAx9joXiTXlZ3+HpONzzX7zafFudjb1Q7pMkl6gCqrA
jS/i3kBSH+6WXLfHI5W80Zgwz+BdfrNw/W5rxqRM7WPl3pJAfwW8lMFtN9f13dkyAkSe5HQePDWV
N4zhAH9PQul0uhAL3vnsI+Fh8YDS9hh+vD7P5c35CM0rIcapXe7MpCcdHhnadJVM8yBN8O2bBB1s
3epV09iLhj54zQ6+iFkzBU8chq6LkbSuQEzx9x17RpAKChqPhXWvvG2C5yiUusePN8oms/erbUim
FH8NZSA/V0cDLKVUrKZlMmhM7bbs+qfqm6CBjumRRShDVW2fesgEqBMxZovM13c0pW/ZIDqdt8Se
z5mfcuBIEQuy6H3I+9wEGOy/d04/7PEY2nSs7KXh5w6T2BRTFCGWLODRKCs9g4+DKFuWzmSpvpmq
fn083hYC4cBlkXyiSGexISq5RWHke90Bml9ZF8cKCVX68sDlM0HntbQq5vTqEvxZgnbpCbn6WDh/
8S34ROhFLuSS7TnZAM9we1l98UzjBXhvCPkyvM9BhOVuKNiWisK0dYKfGUrYf+yJQLCJSKBqS2yE
xUEUz6xA+n/DW7zHPxBoBQn8obQItAzwAUOpkgLWIiOVBnyCQmP4opNrnW9PDNd/QtGRgVvy8pRE
QWAp4pZHOiRKTg4y8mrpRrpjo6VwxmTvMX0jCfeZQmXXSZaj3D4sCJEuCIpOBg9HgYkfvThrVR0K
E4Dvjybo7bk771REQv2SxoJukbUcaib0RzOmUHbGDYzVnwr1TFoyg21tEcPZ5Qw9//QLjKWa/LU6
DeAHwyUS6tnY0yoORBOuPi+zkRklS9S8EBlwWcFlLU++4DIApEqVFVPrsHhZ8yoodhNZQNnN5Mzl
6+JVxEqkCuyi6XtAdPPRBji246nd7A18AsT5PUbPyRORoSCqTfMULMfnY2u8cfZ2hUQEKGPjj1LE
o7czZJ4R7PJa+Kq+1GXiNVyrFnw7PHXw3QlSiZW23JSQTMsi8hHh2zHFC8Rdjd3JYAm1Bam5lNah
xX1C17B5y8mZoWL6C4BwuopE9PgNy1+ng/u2mRKOKMjhY2QD02mxYjabZJn7f8MJ/u5/VwG5Z+LF
oL7FtKgqz6UDM5Gg3B8yHyaNH+Ui2/EKZsSRMlxzKx4jM4uljPQgwP94P1LOBC202AzmAKoQ4ybT
+ohPyDrLSE0f/PwU3l7dZHw52Q63kzR9q00JZLAetZwSSO1bjrXO1VthV6NcNnK58XUCAt0yGhWB
zXaJQD8JOdLbkAYNern0yUTE5Pi79cqg2yWs/7TLXFJbrcN3ppQ5NKXGcrT72oOZE9mMGvPrMKzO
KKzDEUzsD5+yFtVXRWBe6myt8NZ7MLF2TVSYP99p7YcEzizDuo/BzuSTA+ZmliF6EdW2zSnLJm+/
0dN0KnhDJqzMNEV9bB413dIFtHQCOO+fpH4jWdi0pELnD4A6F1Gov/mT6+T4uwbFtYV+IfEyl1sv
8JDyV2XpjnxSXfj6hHTC9sod0MQW37vdU0E1JfkEivU25MDw0Pf8OzoOScnXDX7uMDxO8h1zXWFN
pBhqAhGLefzKohdOfmMU8B8YSbWTcgmX1i1S262CmcrMz2RCAGv7sk49iiUDoxDA4DoV54yvNXWm
utDm+CaAmtPrOiNkOoJuxTinRSC1O1wqivsw9A6fltSkk/GRz3TzYv61otHCwqdCdHAu5dHDBFv1
yh9bFZLNqlUsojgSHHfx5pMKQ7FXop8eMRt+kjtexjrrVEbXVxPN7WQTTb2OXoHUXcWdpJASfO0x
XKWvKfmULRPJg5UjefsEjMecEJbjayzmWl0DG+meXqHCx+0zgYe4dcowERHk+tDrNniXhf6XJYcj
aLLZ5k4JrLGEpKfu6+qir9NH3KWF9qABXKR2wUAES89Y4vjOPjp5cCntob4U09LTOaukgjeVSHBY
PIqOezhXmR2VvfEPC2k9/HbkdBM2g6rY6k6WVvU03TRVD76STO6x+tQWzfhq6v0LTrZAbuUj8T7p
gHEyCYLf2Pmw/LTAwi+c/9L06d24X0FWT9E3ImU4TflVjxJACm+ZNT/YRIPPISQ0j89lPw8d6h3X
/wUvwmgby4F50UMAOtasLbWpiTUwrYGoFsz0IT2REIBDln0CT9Gr8Zt4QI7ANA4imdPhhSiqaYTG
gp/FqUJfyMWTbAFt9T7p7Ovg0xV6mT4exnM/tuHRgES1Te8avjbhp3Hb4E/vwp3gESvtUItUuiYA
DwS3Mta/N0YfOD0aseCiL/TPa7qX13uGAfQykIja3xVqRkdE7bj2kl+JFYvBqCqUb5usUT7fWZWE
7Hqnmuan/f6mEb6V0Zd6iVfHSgCBcCYJ33SX8/lq3Dm9bT4QzOrV6xIzteiUqMqqrVUDvKsbzv1z
yZHmucQeot2J0l75MTvub2eMsGBhA9VW+A6bN/2/dTCO3gwgyBMPE6GNdphMovVOoKP24Bwxh+H9
hrGkwO6uwls8GIq3yT1hgfqU055RI/c+SB6HdUbRxb11WhAZY2xZb01lVPiDz+udkWV+MchQl1XY
IyGN5q63LLxi3tKemqtiy2k2wR1KtNeCFABuIIAkhyWQu6gtUObma8nD6RMcLGiYocjvnbjpvIzC
3zA3UWzCpr+NaB6MpHHy9f9WeikHnsmzNTHV5eF/vOtd3LkGXLZQz3M29JnzgcLsGov2YS5JJ8hi
IZcasQwzmw8KVt/vWSdYfz1KtxJS9qsiDpCDnkZGKerM7mxxxdrHDuf8Sdca7HdOSzSntxg1g4Uo
XyFt9zVhd9ucNyw5EIBKj2RMvzDxQydTFq8al5oMMCvsM4XRWyd3VWqzGXr1JVGXp64IpKCNRcQA
ensl91n8RVK51Oa2XOWh7eSs8Ry6Fi7XaJNQVPAdyzc1mL5uqmYIxVoyjkkZHcu5dTZS/5+5lpjx
QW0BlFMKdbjSJdQNS5bAz3ko8iSF8DBjiZJC4bAeHIiTwk5266s/Rs/RbnJrSepoQLuqCZlWGuwY
gqo9ana8yObjvOhlIKiTCJ6pdBmjvZqDZJoaWbJ1psJEPDP6nEBYaJuw8AArvn0gQlcqNjw/WrE7
rACH7/iGXEh5SPZefpaMoUxWYON1ZH8cPopqrm2sZniCa2AxguQbUSU+N9E7H5O3G0J2Gw8Za94g
l1VopZg9DyDabd8d3OmsjY3h/kl4JvrL3KayR/LkMjJ69Dm/dG27EOmDtaPMdEml2FZr/Ma/D1b5
MrYAvp2rX6O8+b7uvvZLidf+rQ5xWwmDJzvEJYj+0mltWnJ2NXcpm0fjnd0DxiCcuGg4es2YQPiU
W7TzUIwRPRgs52eomhjvPH4Pk3DIOnbZJhVCPWa7SYpWPhL1sKSfMzxsGfmK03fyQAustftph7l2
+Weq/dXjSf9ovYs/BnMh4ETZaoCfHNB5dWsZf0IAk9Muca5uGF9V1P0soOAqtu6D0REe8oEK5IaC
/rNW1+Jwhh+btrmDAaRxGkO+CR6M27PUxXclOMlWbdNmV0jdxDDXrutYelWnr/DYfbMCqlzf6RWe
Nc3vij6RJazk8gLJuhAvuifFOL31nMfkOJrt/cPq+8ftOLTXppYP9Cw3dl4NRcidj25gWSJOVHy4
EsFe7X9ga4mvrT4kS7yFQ1PF46AO2OvQomCMk+1YNL1itxp11ZcWkqNjALPOqF0PXNHj1++1E42O
jXy65fmi8Sd7aUie+cOC1VqLU63UjgUU90X51FtOIfu+nwH8ciXmuJ+9smPuM9EeOh8TzY8jTNWD
t3A1QDShXxIazDu+mL69LFTd0dT7MwolNGadiBmp/eOyKVZxfNUAocBH4bY2jjFpku3FvoeI6Erm
WV5nVhypC0Dio5cDZtYUJ0jFsGI/y1wM2yZrctYKm8+QNvYEjJED87nUsJONL0gm0acqkJRTzZDv
6qJIASvVlJCPd0VjrzgYN3gK/j9KCIIixdbr4k9+o89+3EfSU/EIESUY6fn1EDYJOttzrrCjDXS9
68/G3f/haSTqKNSJbuuFGHvKAX7qJ3jT2+bNgSTw6xjzmYddMsseO6H4SyIOhdPe0u/xdhLactmt
lTXz3X6O9yPb2HXm6i+g+RIXwEnlIurrVSyVnrNNtRd2M5sQdOZFKIxGboIwVkYfRRatA3qQh83g
T5VLThFFl65jtrkORs4GQQe4CxET41eDNdr94BaX/HwVo3ChmLvxEV0142UOXaVcK8WVF7I0iBbu
qZoE9YWTo+92zhecmdWsyHg4X62VddsVtTSk9j1RemdcDX0R/0hDYIFbiGgETLd24fv+vHZXfeIZ
sEqxe9IMyWUa1YQu880av3hEf49EexI2Tkp7LqasMT7qyRddMLMTTbD9qM0e5sPRcYI3IkC2bSuO
9m3/dv69RCiXALlJXxB3gL25m3u+JuNwjPXrjCFa1b37c2KnnQ1vshAIwvmX9P8c1EuxZqeS6jF5
/sCEx10IHzFeTdqcQXgq2/Y9Q06l2hnOcw2Hd8RMttJx3r9fCzGbWANt9C0rhOwNVv4QiEV9Uu1a
dLaJNqUbxa9umstCoWWSaK5/614JCUFNjQXab6TfSazGiZD74XBkawKWii7cd7Fh5NWqB4m/iBm7
y3R+/1rmJ5NOmsX++NyHTxbXbW7ey+mOwDY+vVT5BAoc7wL7cPFXxRKyw+2e/YQBZX22wYDjsSsr
ycFtkeTWfrALDckw2NudEDfPA+o3xsTBoVM2eH9u1l30tFBQsA54J/Zj/p0agnxPeq4ng/eMCLeT
niNYFVGUB3j4qJiRLbozfUNB7upnNkjxE70YawLpzExRMKz79s+Tg7b9dPFqhNxMx5Ab2nECznFF
2QOoO0337BqnL+/A8plyVCIqURU6dcDh0QHWfDF/i4PiU+XjpqyCkynsUaTCifC0uLfWeU5zqb1U
3FRnx6UGcQuYZfepYtlAyG4unJa2lnYoSFXNnuU+mYAPQgeZk42fYx0P0a0o196AIDcdFaPQ/s6S
4CJr0XfY8zs1FbNiB9UcTMxRl6xHEwIN3C+mM8bRqIrqnNDYVbz0fbcI5A8uIP7ZJPfGV0+g4VfF
bUe+TtlLIvf0WCXIZ+3i7E9TLidNUFDj9F4HJGd6Nv9R0BwHIBTH0OWHPr42/pcOpxpSG3gn3GQ5
xIEMQrTHDVMkITVU5EKRsEdHM5cii7l90YBarNIm/FPJPugAHFGE9EkIbqpd9LXk4QB+w5cfCOVI
Lekp75+6lepcJofChbq1fIEQ/jKXeBHZ0MH0EqjJf0a2YIjk5smrqxMZPZMvpf7Zut0pzFeAJsia
tk6HsVgzhCGPnrzNDym4qurNhBr4Ldy3tMzhyuRZS9Mv/+o1VsqY50jtSNGEv5EiwQovLpdR6shr
t4pECJyeX76qNw5NzV2c6caho5ZTD/C0YozO6NcjxY3LEuGzIz1CwKMphiHmmcfmynrjqN9VWuqS
8PUbhBfl+lZ632wuO3lvukKzbnSUZKz7YP5+ZKFlK5HueIW90ZpavP+InrlLLat8WI5j6ZTb0pq0
KkNEL2yNL0WzmLShX/uKZQJYOQzcAGH451avV5Y8qL7AH3iLWA4FalU1fHv47aPfzH6kJ5cyhzNe
Aa1cY+umlRXJlZabEcbUvi2/Ik+wXpBT9h2G7ERj4tQpUq5hJY8iUh6HskUiz23g73NQKIMtUaX1
sjQctySj3hamcihQg7NUEkT8F/sQrPHNlCKDk9Y1RnRhe8RDgLUejsZYtM75Pba3C36ZZX581Hfk
IU7+gsu2cqn0xpXo4J1cVl/d8DjVG/jYdKxf/tOm7O3zBGj88rMcQQxuKUEofb4Wd5TiFqkGIqVr
MSShmgjR3/4FxGsMJAQMQXV5pK2RMsm89xsZBS5IrtqNBiyuvd3LDWvqLok0mtq2fziKnyJii6VK
Q+mSn7ij8FuuWpDn5GqAN9jYZsZmqKPbD/4VhpnWrikGUSDpOXbVLE9hti1oS9MgrL4Ho6yWQwjM
S+nabeajuX9vv2rVdQn/XQbuT7B58W5q46tH3celUAvfwaKKLqx+wWyAmq24t+bZYRo/rfCUI3/a
qZDd0QY/9tXheKvM+hA6c3Np0cgBKstHB6mE6HZd2KYm7FVRuNAOL5lJlBAZ/dsdgZj+D8aaiA4r
NZ+s4UTgagV3UgCCIM7uGcIy6wqkrkqp9InqjYJoly86YVfh83p1RCOrFzxBx2XKBvOto/szz0In
fGKINXv0AxCOLDpy5lAE1/xr4ycZvOFqZCHYLozns7h5pk4PCU6WbnrtS9s27oulxtF8pe65VC4o
jtMyDvSp2tC4vpvLGo9kqr5JaodqmIElDCSCNkYOvf3b+c/aiHlC1dJWUTcmcg0K4LcaqqNTEOmt
ONOm+W/lq76r7+bxGIB4ud/GPdr8mreDumDcfkwDMWGL6+TTU+Ucx0aLwDkjN2k2Bja+d21J5oOZ
Wv6ViOf/Y2Bdg5otpYymh4wNzEzfFFKxfi0cmeDYEQUfijkYXKVLCXHX/GWaHJTe982dnxd5uI4t
lGN8zrZ6v2P2xwLEUZ/ZN4b95x6f/+j1FMONiBRY3OHdJz6nP2xI14+Ger+BYZwDJuiRKQNfQC41
OV4WOWLi49Agz5Hvo7Gg1Tvge2dbf31qsiZcgCNgn4lNz0ThU6PWIKgSs5H/gPnWvq69g9fFqm/2
EthhNbh6DChMpErK7fILwu6u9iqDoXCgUBob01G/9zpN0AScN3H3esXWi7zFKHR44Zxh5piuNgqX
L9/gJaHb8+p78s+oksVNcxKrKJEfDXoYM9n9OVzXPUXK7rEuwYR9d4bbL5SdQn1jHL3c30L1rKN/
3zrAuBSbbMjBS0sP2QzWPdydH5PADO1k8e98Xi0lTbDhNK0emQbrPz7ofplFDvBgkISJfk5QQ6il
AwRuFmZwMB958DnTsB9gQxH4LxrZqZ61wbE1wn8ZzDzNaU59UlWxwqdn/WkEWldFUnIpkLyLD4JK
U7hrJYRvUTkCm8yuKBPsx4eXePEWQxxYn/x22vYuSe2m6/D8G+aYl5rqiUab0XUDssE/23xq1aPL
h2JG/9D6VYhsY9R9xjWa3BbTJr+4CSyChTODEwCUq7xRZ8VDB12yRZkjBqRCD5hiD/kV+uPWkYjz
Tlqp3M9f+wyypmY0kE/VNMX+rSy8e42GjSeOcFqXftmj7xckQXmDV1CYqDV5FKqo/hWUO52cmvua
rZuaPLjpFsB84y7h+8PwLjI4GRGc3A9hZIyRe3FLCBIn+ENF+T0pkGAbif13sORN3sJNEdGBC70T
el+JeKDnd67a0BDDsQ5ixgmqyIt9bT3yalq+X5ODY56FwEfMXmsxSN9BcH/+DzttvIlBcz+os+Bg
mE5pi71uRR8u/wBix7rj7xx7yR0OMJZ1v33ogFRD0Uq+jmGd5CNULMUJguxVmlCTvruRP3vVv51a
5Owxd7axFeR3dYzMlLbvsbm5ewU5+IaeVxpEvLFxQvQyECOIOPLQDNAOn2WN+HT6lRi7k3xJ1afr
PtlsiLkQkGJ629v4er5XbEN6bc7I9HK1uMU8Tpa7i/3z1WzzBXH3+n61KI/m3YztGgGlz6k+zR2B
HWIN3HidAKk2XfnFP2NJc1TrIBayJPQw5ELsYTBX/e5G6AwZvePnMsUB2lDxq6i/1J5CvohMQLNP
erCaml9fBAkBr4WYXlAtcVHn1Q07Z8qh1vBf7jO09wnwBDujsYNRGPzww45xk9Uze7+53KLx7Esy
M1TkNq1plOpYkSedXWzyo7KCb8OESVZGBiNQFmNAO1c2VfizdvroM61fLZUH0f3q06OaiJ4SMNn9
KVrE2A5/OPNZJc56txVAoVswbR6/QPIZGBLT3X9LwA+v7PcGS/qGAV/NLhOl+hl7jb8HNOH2XACT
OZh2+hqHJnBuxrLuncT87t7o02O1NtBiSSgwP4u+4FsIP2Z/2rCfJH3wTAIcj1mzeRr+Ij0JQhPj
wWOGLIsL42tvsn6UB/N4RpX4vGMX8THxu0XO/EqYEoUgrureqprPUd6C890kOuyImHRwVus25pRk
wArOrqs3IBaT44RW1INxrc1r6EhyxMNPwzT74EncQkoJLCkA4MhL5VFRSbQjENY5o1oKLsXRwB7O
rSN1EeO4c5Yb0uD3PHKcsc4U4oWj5v23XTuoTz28QbdpVpJy46AFEDek14JQ+wOZG63MabBWB0vL
rU7RUb5DwF9M+nbjvi+cOjTmVW/mvgCAX4/Ro/bZZ8NpRc7zwB7ckktTLpl7+blPtSjCoRxS7WPP
ERJFCKI/Oqv/SoQJfX8B68pJN8Q5pHe4J8cnpxM0/7rpMrdOzRozBdm/SxuJhZnEsXSQzDVLjjvJ
Gh6dCQaN7eq9cVoMVXgrkQFi9Yy+EMObrCgLCi9PfvKydU8akTrB2KveoFiS8elL/bSY+IWLPCUb
td0E3JCwarEd6cOiuzldyZBQsxMLxW02gTIGIaQ2sQKNR3Mj2qjM8EyKhSqhFwCYYlkD8ewqZmCr
NfAZGSlQh3VJje1ozfg7Q6+aTZtc6JYMt+eD3GiNj/oyMMwebbHhEIOFCgWK2TrAw3j7h7rcTrtP
tF2MtD+zInbr7PlDIGxkAOW+ozZHwy2IvN04It+u7KaQT9Dv3I3o3w7C9d3vgdWLfVm/MY01Q4dz
mc18eqnqkS9BJdHEzGyPc41ztRzF2AqSRztescuVG4TTfF7zSod7BLx02jiMQ4NMf4P263EyYLQw
4cAB4iIJA8lOfZRZJk3mNF+8byvcMh6lHvSVAD81FJGA90pgL1bgY3kIKJYA5eZ5t2SuZu+kA7b6
ejUgNFKSBCih67yfRtGbnEWyxxsIkCFY00zL3mlI5b1FptpPk1hmtGwbAz603yrRX54vk8nsMwyj
pLVgL3beQhLJRY2smCGY71xtsaNfnrTwbwWCy6qYKgTjAOm25UpjUeZMGO9tVeJAE18mJOhytGCC
1ZMZtZ6/56VxnN1Q/tv+HFhDTrR4GQbkcW4jebrUgU3aQQCONZ0PRbfB8ObQDRVW2JoEXQ/RWa8P
Sxn9vm5zj9mo/sBgVJuBQMAwdGXvEkwte17hBWfPvDQOBKMkHD/4DCZ55gt7XaBJJ+kluoSmjCqS
ViaVxZPDYByfKNo3SoOAzvDQ3PpwbpIHeQqXeSi5CCj49608gT8h+B0Bnrv8DSDpNM0l3QqZpwlC
tb2j5lRWHnk2CLgxZbazGelwcBq+EGGlf3SGw0xrVmMltrzp4xY+zN3rQ+N9f6Mm8L++TMppUgxl
Epemy+661sMHtTNouJds11+X5+xCFRZWeLcYC1jelHivLwdlmhIQVzDPwJQw+xIzjoP5aDLj1+WL
/2cbT95jzUks3y9n59Iahwt/lNEkMZne2Q5VnJzUZNN31DH6Rw3sKOYf1/5SJimim3qrweh1XTir
hcGMjKX8fVAzUUjWNCQ2GJ1Ia3Fa33fh6+fjlMbk9yDFGl7CIil45Twj3tfY9NoE93WWPKSKCktr
mdzJyJxyoW7rSPCrazqT+K0yv+OWdWPpmrY5e9ASUlI0i8qikmkKuIGuMQ0O2rkcdQtvJDLG/Qgc
gfvV/8555HNZeNNdMnu9rjO4SQ3S4h52jDJaxYNvYtszIKyMTKreeoc6wg0+NlsF1oRktPESQVmG
vZU6edm/EVs2ypgLh0Csfm3OAKuYcpRkq2ceVzTwsREMUGmi1mISVLBrWyn0hoqqGdtedbtdQZKm
epv/E6I6qUwIUSUJy9XLvX6/3HvlXvPNdkaZzeEWDPa5JyZdFdxnYsmFdR4D2UFIRwh/Q72eLMTz
Fi4AVmvSFm3FPC7cl+vLQ/pJ4PjUgaVg1PV0pSur5q8eoTBAeWmQDYkHKeujOjKZs5u8B/sKtYse
eF7zCZp13iaTHnTmjJrFveN/iJfqtCHjE08D+9E0l/i3qAfwF97Mz81q4aPisQOmbKuT0hdOf0je
Yu7bcsBYLq6F89Tm/qbKfQysXSU1nEddY+xcQOO8J3ms3Hce/aydltPy3wvqlFoV/H1BdwL5dnPq
oMz5Fdem4HqVls1J+xtK02tZyB1s3acl5eUMl0ZeIS7KfHLTaZjyKyalJc9xQVNGkXa0fqp2F5It
TCuae7AXabNcAwiTdJZSdu+UAU6DEH+TpaIJAkxgsIJz7Db0iqNcEgp2j8lGytUjNYnDcwl031go
VRhcrheDyKBwOCtIW+iY+n4ZnpvgfnqpMQalxD+6NOpF4dT3t8Rvb273chlZz4nso1+V156puOzw
QtrB1UJEFfsleDPk1JQbGq9BY2O8g76X49doXEirIxBrAfzIEuAst/2R/ITqFs05Q2UNib3A20Hv
8m/M/ZZ7L+ZHdkBzF+2+k6CUutiVEBUPFbyVOSkOOM8SvNP6icI3bh3pIYyaPOxJeuNWgH3ljcR4
gvUcZaX+AjfJ7/yioCjdvOS93D7Z+rZGiY11tUFEmYkG1qCcsD0PiduXzDivb5lb3mlcyfKTeQkr
QFBOKYTzm9N39ckUz/PeSoFjXaCVsoaC3dO124r/1wF+Bf4fsDQyb9ZdrJfnqOpihQvDJty1b4Mr
q9Lpo0+mtAaGEssazZftZzzJSAFe9QJN4ZIOWcZp0fWD3M4NFppuKETAoRajRSVyJCFFBLJBfiQt
Ov3H3lzG2iGHvqiTNnEerUdbSqFqtaDCv+j+kmSgDqRgQEho68uIWqw9ONq7DxduaoT97jSZWz1j
rbXwxG/UInQs5xtn+razxYQ5to74EMNMDTAg75Dcgus7FDn2HnX3YMvREgC6P//D4jkrlXyAFHwK
KGf/ArE4BZSpMAMVpApsIk4aTN+EBoD4Xw5n0mxgE2y38BtnvrSQAdKPx641Wuk3UfDXzTtJ2XRS
FxVB/Cksb+fzgpm/ipFwpOeuKWi6NHux/5o18pzvW9HGu8uPr5k2hxV4ZExMcnPXyPwWqW8kV9kR
Y4VE8VQazzDW2AIwzADJhwQ9zwwAwra7u8NXBuKctlkUrFkhz9QIHcVxCG6iXzJ5ftwW4jEUR+wb
LavJA3AKkh8YDU4wEhIJSdw0S3GsC4K7zD0eckEnjh5MLEUP6evacrka8AbAIgwYh/Qj8DsbhGOp
rNAePWxkapz9GbajHgULdUwDqTkUeKSewlUfYz6zrWl0Cgv8+6CFAjbc6lj+36wWUsdtkcKAlZLF
6PU10i8pMqotdBgxVnwlepVaJEGpijFfquDl7GUFialOv484n0InQdS1QO23XHDDzTV74B3XoFms
4Fagdq+EIdhqbf4/g5x8V44LLIVMuys1H+lRYG2C0HCadpdS8l6TY8LNzy3rWGlqPxzlfNvfpQh4
SSi+6WvsWssM09jsDbynNkYUyxQ/3ekM8kaUxDl/6VI38DNPGCzA7QN4JX659g6ispU2RSzgvpsn
BOPjvJkyvUW1WXQAoKLZKkNYBMGAXPFnOHAuYTNBVXa2gEahMntvY2ryRWrvLdlz9ru3XNr+7lgz
9Yd47t1yf0WE6CApiemr3azizlUq5AyBOqjBqCWYoI8Fg+UebJkiMZjEjV+EYAhdNvWt/fQxHJzd
uwSwOTOc78pCS6U5zxyWJF1C7hTgVARRjDrJVltljdykulggheGPVGWNBCZFg9LQveCGA+zGToBU
QLdgORre+oWk+ZDBMSnr2UaXFv+y06yerHkK850zzMphxEp+WZpNd1ELsf2gVxujedRAzuxhi8Hk
m9gkEcYm4aBR+r8/PUA7jJCWYTvJqxChW8xB8w+2BeYNC7llUFSRNB31KTZ1g1K57hDT+Zo/R0g0
DXCIxmOKdekWKQOxHuF9KjjzvZBbV+pieMW3CFGJIrdGoocW3ysk3C7F0nRsBrZjQXfP8clMAqa7
3kt97e59BPJRIDJTbKCO3NDmWu+HtL4Jk2VQ4BK+d6lOegURj7sDh493j1cr+6DnZBix0xUlpQln
e8IXF3aGNpwyonQ3tFkfK822OOiwPWTKAOSOdB9L+4C5sl0w3RVwYYb+79QB0l/Xp2pccIyYpdT+
wo4AqXm6moG4zFchYh6JbikUxFMCn+7tYMqu8rqvVsRIhwHTu52yDmthhEZdQRc79kWorUJFkAw6
bm/NiPpBPNZRRQULykqHUOgk328ea/rjp8ZtbKBI8/4atdSr5iiIfvhu7olUJ/YhnJBj2jRsNBYS
xk0iSXQkjUg2nJv8LKvm+3+W1rQRRUToF9YrM5X7MEEKRt9JYxkqQs0Vw8FZyf9llmOJ2T/XryR+
jQIjYbvNS/83Z652/qOj8wu+VtJeY45El+fJP9+ZoLljtRUNX460Fe6YwZCUbDWpUy6Uzp1jWooC
k0P1vg8P0X6dTDFP1Usl/BDMPLSOblUVd875EKQ+3rea6b/DW29UN3W5CZ8lUCDPeGON7xIAzQ9y
PC1X8PigbQ5KOZBnBN1V3GhITTTsyVRrAvzkKPGTjqdBEzjiE2ZSqHPYpDiRL8XJFHx1NDCb5QZH
KrI+OTU8L+dU3yT9CEnycL0u/V6oJpN0Gb2jW1Jy8onhbGpI0HpvB3juPn+Icqmxm9vyBRJ+w30J
vFlmXXjqsnf1ftjrVymYvJPGzP30fhjfDsC3HK19Wcvqb6DeV+CQjxpt9cs5N7Yp2+i5S8TPJw3p
IQ5Wdv3ItvGV9bMbAg11+F/L6sCO0NkQNZ0f0vzXtSFizcuwKUzOyrIyevB3dbz//bbwl0F7jfI6
+vPe3w4xTlbGoqE6Ubkf5ZzwAL5FH8Q09okUy4xpcvv12kO6MGlY1yElNQk9yFpv4P9oCzkZMh1j
1YdEXOFDbVIt+aUDxr57ZtwZdbNcUQUXsAWsw1G4n6ZRExqxPFRxdrfMz08G9IgxlnuX/J6FRZLX
a0hJh71euCDtuu1Wd6KaQCiCI0/blJ1xkmw6CCkVWOlstj4zRtwzykc46ygFo1KX04xyA2ov7uk3
tw08g9lnmmJWaPW4g5mLyIsoESkAanq0qsRwPyZp2BXrEGWP9OCVCVOD2p/8fJxui3mw/65P/hpt
/EcQkqywtLmIBrv3uiAIq7t4cR198dKDQMGnqY80PaVKYLKM7o2K7VRgOBLvaole9edjNia399f/
sl9Y8xPm+Qru0RssbpMsrI+RhspnkIMcIXnu+t5KvoM60ih/l5R/zq1Jbd4T9vxqbqIVN+s3TLPz
vQDaYUPAj5det8wbFWeRc8ZI17CtgJcFnZ1a2lG7vVFEP3+EVGPOLIlddKKmGsqdiCjbDSSzM+B+
CLCfAa+IvbGIerMgYfv3oN6ngU/NOAGHJmeZxNc7HAdy7pg/jSWBbRKf94sZCx4KwuR6RL7ke9mF
3mRkJmKKA8WAmTC+Q/oq26iRCLYrLY1Vf8SSmkA/aQVxihVlhWJqdhfTr6kB4Q1sS+9VI3isdTW2
hZ14IwxuVlRihQfKpKdabLvjTYNGoNkitESDtj+zzcMVbHWsM3cybqYWR1M0wu0McUiBiu99jJZo
8gswU7yU9UaaBqashN8ai3Pir95s0wEZasWAsaQe7XW8FI1s+vLuoSbeaaFYVF4TWUVeN20raqFx
FgJvv83BguDTJJKto+ZVCMyzryExkBeNGnpLJU+DiYpZ35Za/PPszl06HPPLJioi29HtBlbFfNeh
stm+I6WB5WyhGLEzxCaR8MRkXU5eiQKoGHQJ53k6JriPp3Ks7oFRo2v3waCu3pUI1iObIeFt3OMj
M7ScBVp+vdjPxdUg4N3KYbUeLDHZS2O71eIofXCAqHMZqZWCWXzT298SFyiizGitSjs3jCfAPBE5
Gg9Q6sLINmyLFc8Aj7E5KiqLxwTgHavvv8kBM9UqC+fPRKHtLwRQaLuJgqwARCR4f2asvSx3znKP
J/O2f6vE8mw3G0LM6yrygOAHUlCDHCwkLqh/+k40xAapcivjtDm+lWCDPrsT8dgHApP0nMce/Ult
UX5ea8Htm+A8UgW7rOARFLXlvDSUnaaiMsFn0SAonS0L4kx3sihsKA5WMolcupkjmmKrG2S6S9yI
L+jC56GpWFW2qKTX3VG4B3j3NEZGzUFJuJjU1GndFCYG3MfROfYjad7b2hhdgzgIZYDx2f0vUz2e
nzeXT22vL2hWbUzf3dY25Hhfy0GQXWm7dmqnQGUohmIYicrPL2AWXo+YgvsMBt8aThk00axPgFKr
vd2BoP93fd9P3Q7lt5R8Ci0MTvR28gHIynFmizhiyk15TtnmfJ7m2qhulvuOhRlrVyuXbCwXsYyS
XQfrODV/RxnggibDGefD+6EMGaCfRnMfBwut9xYxzTiqoEBqpUmMZFFj+kTweaGlpJyiSWfYCOAA
8pKkiiWSU6umn/3WFhfJQj9/pv0dVCrMnrNDsDYzfTrsQZQGQwumacwjDDRvzANFQF4UAFbB01/X
E2BBJVlSYRB4JX/xCFMKjqeAOnjUrKbiOuCWAfGz3scWTlo+66/hUSphkTWy1UQuAWl1WH760YJS
i6rY2rE5tIewDMX1HxHqTndIWCYj4w52We1IfBGbcLQJ8ti7+CL0+VoysIge8Y9Juby4+6A55Cvp
X/cPvZJpnfyIiYih+5uovtttdGl9hLChM+7v6SprfTuntz+Vqj49YcLP9yEET4qYdTXA8ENFceuF
ieLzcrBsyhZUeLYl/o9uslLFMYkkWSdMtc0a1vtSTfnKlN3gd6NqZSNUQbM+s5sLyi9n7S0bFmL3
6hFDyymEmM9Tj33URt7DGW/9DTE8en44Eut5bwQiEgph3iLoRmdANJS8JOrXw4kgUhuU7NcTysQx
P4rvOG3Ciq3IHHZt1sXqN75ebGfrNVzIBkXdpf38cVFBrO39c1O+0j6T287U1f+XDFvfxHk6qoM0
3iu3iAXKNF223HUOG81WI3A8Iaxwthy5AIDM1+fzqlYQmuUxZfL3t7lOZfk3tlxJ9SYFZDG66O0J
OmM9j2IlKIfkcI6x1OVzr2COIyw7nZ5ObuLlsXVGfMPjT457m1jM5KQYx3++qulvwkz+6MBLWsHz
ySEbhnzTymEIpsCuSHkWjXAu7TF8equWJTuu+kz9v2zMtRDju+98zdYtmSKsT7jKBb89g5vTsVjQ
K/7bzUmKNNz34BGabOvz8EgeNvb4FRJgIn008iJPOVi66vHRIz5Ao5kBhtCm+AoZuWIful0LiVfy
RjrrxZQrkI3uQbLcVmrSqgywPTpORoDaEJoeHm+pRq1sIZCEz36O4E2ll20pKjjBA/ETKmOK+vjJ
q4JkZL0HXsU4KG0yBFIahZ9xOmZ+orBzW+wo4ktsyyO1g8rhgEQ7xz1Ra+mBKgIxLTk3uiZ4/YUM
UT7+2eqp4xPtFW30ju5JbF8ZERLWz0FHLCKouzIha6jDv3KhswnQXbXO6Ay5mbkOZgltPQrfzKKQ
EIJ8GKgL9GevpT30qkDQI6RQMHr0bCsVqr5VwFC7DN8tMaatMIUFrVVM2/qvTUyDs3fzGA6ZYIqu
EYCPGjZa4wzYogrRgDneOiPPdxDFzkP10tJx9YcXzCDiuGX+4lTyn/3YQT6v9zPUxY1OP16i2JpI
AClTMYS32r8tkXduxolsnfKDFXvgiDaUsMk3Sz9WKT2VZsvUfgqOf74pur8VsMPmugijfpvA/giY
hQoXHxqk7UF5FNVagYtqyBHYKuR8xymmH5x4USH4L7tcdhIMTiU8QKjwM2Z5dtQNEoV8phDi1VO8
F4oRfXokJEEyuFUVRb6hwo77lFR0VXyJxtRlNQONbw8j5ttTHtOr6s/4sqPC+za7oS4KGMDAbMSL
IXU0zOSGI6vxgpXu1ecrLQhk1y9KUD3NdFMswonTSktkvZ3K1QXbEkktir06cFnCFl8RhAXmgAbH
/kbj36Am0kuhn+7dkYFGC58Gg77AFHsqrj6fwtIf/Awiw9muRRlj3FVyYqwf0apd8qrjANBv9DQE
h+IkMghXsn9sAo+/QC2Vr5RBYKnesDb4vszcVFF3FQ5pxZdzpBiMpkVDfOfcg8XBqfPqkLKEQO3C
tIuTnkNEU/gcmGK5KbJAlpgbDXoAjdY5hMiX+rTy/phaX0hErYzYa+dgzfv4QPSdbKhEpLrXRt99
Z5KPrAUa2hoyylABdpfSAq9PNlRfCdnrPjxSLc2GSB8UXcRWUimTGAW9EWsXWiUjorbBPEXnJuuB
45cwhXjZ7u7Bfg2zAMdFQaNpC29nq4eoTjnua2WSr/h5C6qA4n3XF/e7Ynop9KsJhweMXkvPMxvr
t4Ap56DDKUWbynVeztTcTpGTqp6DJB3sDAztglwXN2aXXp2F7pE/tgscqtHZpXMT157vQweu3fHp
6RJ2Sm2WpDbJ+pPZytigEpCEhxXNrP+eSDGPlH/bdOJrzmLSNaQ3QldxzIvKAOOiBToD65GaVSzC
JNGGSAqc0hWdgrX12U1brVxXkEXXxhOJ4fvHuuqRWKPpAuLarHprH3So6AlRSwFBd8KPaNTNCyyO
wm8jqJYL4lthCFEiFwaFml+6za+9nQBLMDdgOurdN3NdMOl58iU83qketB0MN4ng4lSp3W3ROUia
OKm3c99rSZdu/5q3iSygTj25f/xsGesh6rq5WFMt6PvFj/tP+qxJdn3zMMzEyaXWNeiahHvVuHIo
6nGkeKNCC5/WGl7pR78hnskpBVPUblxN7r7yQr+I8RNzVdKFTERJjCiDkgV4O4PCEdwcc57MKBAw
QpRnfch8cG5Hbh1X55jJMyZ3EpINMms+WMCqlohyeXjnRaY9bcfztJL8qxV3hD20tDwpZHlw8kft
2WRzbNWvki1+MnqTB9hCpxUekcFd48Y5n8AZlIkzpCuLEKD8044jHP68j7Zw0NTXEc9X7XlW+ai5
CgLwYKIvAZOASu4Zl17QaTE215biRojey0SDHJlIOnWTWje2W2+vH0eLY/BSitqNugGTYtSyZf62
QTmZ1UXI7z3R3xw+9wdk8J15jWAUUd4BXr6qgMln6CtRdJgv1GEseMj5xIj+8+OY6AmRyJ2br71t
/haZUPLphVE11B3BWf9se7qz116hXkDh38+SN7JU0knRNZKveJ9r3Da35r+5h22KlAkPHLdxQvSZ
f1j6KuVmTpR6eSKJ8tvbIkzjM4pDIWO9Z+MZkXbU0vyDhLhbTWaIgvYW05FTALBj+EhDqPcNTmzP
u2mUJjubhvhKIjvwsPFBY5TPKqIXqknWZiJUY6VXoLhm37cEMbQE7tTA1HymHOAil46KuMppBGAj
bjmE1d4VtjhSxQ03cF/0ESvkoUXdGQwBqkFwrrgc3pEgawN6wnSYOUirlVDNNwL2TYAbwhiKE/oD
GSruxWGnadwko5iUPihnW1Bjx+mnCHwPT8dgoKHBFQv4gC+bCrBippDyhgBw8Ad9WxbKK85vkJ2l
kpG1t+WyBSuohL/Q/29qpydR3mr1HVgi0H93dhsf9sQjtpMD0Y9DyNVXTsitC6kcUjTik3dO7pm5
PwH/hj3toTKKAjkJ1BcEmDi+2ZOBZgEBeiaKgwWAAzTXMXBqxgxtuDJdOJwvbWiQ7tRjVBOZIwMJ
MOOCcRNLQs5iesalmlwi4Coq04bWEv/UqJD27BQC9BoRhLioNefdQGhe6o2SkLEHbMk766Lnl72e
JUU2JEQNNIVPZbi3PMwQKi2NKJHgF8zzllgVfcGAHfdyDtX6K8sPhmv6ogLDyNm5dVzZ4WuF/nKm
OQQuabBtjnXh8p4VU1hWvKQapxlGOIxYUOMCW+ODWFQxvQL+4oO0j5Yi02cn0qVKV2e9NIZ05Gne
f1spl7vMvThbFssQPj8E9WmiaPPfDgX2IirDv6howyB31KaNlvXCxepBUsdEaYHw4Hnjn77yN0TG
T2qi3Y3HnuRgs56WSW31QDKXoUEF5Tl8T1ptqU52/3NcAJ5FbfpwFRyRueHR6ZUsxd1IksdiehD4
mM4RyFnxSDE05Xy0V/jKfi8tHhSE3xdFZqtCHjBhLhXPlJSKyaSK5dI+Lg+4l6LHzdsR5HOtQyOr
JWlD8FsOTZjBuquJCM4oPfnRa8Ll0gjvfcTT/AG0TiDb8ydDaWE7hQwC7UxBAY6FRmgnTfYudLiA
fPhsuytfern9hgetsjWPI6no92h0VAwzDMuZBdjjj50h9YEJlFNEuE0KBA/QfbsjHGUmLTntdUiW
SUjQH8XoLEIJxT0P62YS+ryxGI4INND5c9WHa69x+mYD2L3lGnCrilR2KdrQ2el/BiUoz1s5H5GJ
rHGa9NW89ghcGsOMN6MFdILsm4HfZm0s0DUn4xYRS8XZAYmJcGalC/en6z+9C5flN1mnpRpeW+iw
8DZOQQvLFuqVxuZ8PnqWpbGIMJVQClUtG/64sjeqykcll4jr5Cs68YsQgSZZZghEG5gs3BJnNQ3D
isstc5suVyToStqbGxIW8+zhLnbfYrpmlTgMcG+aCWLrvFoVHeTFXkAsUT2BGSZz25FUi9csGfGn
moB7DauP9P8D5MGuvJV3s2yMWwrbbGXAPnr+G95FVsdK3w67wZb/x0bTqVUuBgiRKcBdXZKhKWku
nkD1wctsFSVo9YpgbBRq6akutxkpOfsLqTp//Rie5eGMytX09yup+ODhHWFlel3a/YQczvCxjB4+
elGeMNmpVEQQFb1aLX4DPx1yIYXepunsVmH0nXbK3NXiiuavtE0fDASheulglkA+SfZB9seFzYTn
Oto2SYE5XWLBBAf/v20WrzPfD3hvB3DxsanlLZPbLioIhH1t165RxDJwC+ZQJ10nS+ZkKDM+36es
JH9ifUN/RK7+dFN2drG6lZ36unHq/kOTs5u+/UKO6XZzY1Tndq+a1UyOlV7WnUsLnjKjjbRDgnIj
m5I44S2x/rs5IGdyoxVLYJwtlAPXvGPVpUASXah1nM/63TvzjiWjACvSxJW8TWksKD5NGC1V/scz
NPX6RcILNh8R6DdWq20RioBEI3L70wIsdpwmBXLrkv0kTo3cQXKJVfAZoi3aiiTUk9iLFcIr6/if
hIX0YHPWFvz48WSR4LrscvbnZwTRs48rRouO5h2SFbrcSjBrdIgNeLccLh8bOosCHF5F07DMwGE2
vLnquWQyhY3vvjgDAIHUvcDFhsraSAV+R1OG7sAoH2GqbTFs0/aSlo1wvDWmhKG4VWCbuT5hBPhW
nmfsec9ntsy/QiX/gOGmXCIAkzQr7onv+OOHY3+3tt+plPylvWdghnOlhxYgQzPORv+f2hwUCff9
cXTcgHgT95U1/Rhl/5qHnLvIfP0wFQ/x94NwXAOJKOYo7k4igc8L77euaf7h12aeKNwtsE0DRIGn
in8XuGqdByHiLnT+bABmpwIsVRzRi98iJ/8OZ1mRhJturHtxjAo0dMG8nZ7mx8rhXHqqbBTqnaeK
CxVrorIsOhvRK1qalwV7BNf51+spDIYy5fRZaiXFP4iS2XvXVDXMvbiRzt/w93DcWe0vtqVAI7Ek
4iLT4Rck+TMyLRe//wDIa/aSUlQo4Re54syXzkhsdrw+AQloQh18UDMmLPIYVlr8lrZ5NvCd+1W+
F5LuYAcHEN5awhd93cAL87tKQIqWhlt2TRoRtg3yRV7zFGviCImggKMRBgwjrqy7twZxZCAGw9e6
BVas1J4yCTPyrXRfYk6fCOYgUDb0aAOobxHpM2qbNRMwBP2vFZfCG9lVd0jBhxpqd74oUB7Eo6rD
cCBGUPZ05tLgzWunBSmCmmCTs/no6g2KUcQYWI5hKeSG7Z6+U+qxKQaoiaiBduGi6Gi9Son/0W0u
MeFGFCtcNA8LCYp4bBI09VMa4X36lRJD0kMQnEcnrmF35+K4W6i3gLKR+HRuPNj3moxrN7qu0JjG
5sxN+jSEup28Z1LEgCwGdJ/0DvxpN5QO8hr+CtRH22mN94fCIjenW/pezcK4G/EIUAkhkIF9HTfS
zpOEy/zdupzRdODjphZhzItVg06bRHqDZIxRrfDTSXpYs831QnFEtc3gI/AQRLLg/MwmczzPlffW
BtX98HK+1YaFn8hTDe+BqYUnjGMenpRq2QSkYQSN4wIg/k9SL5BaQi8CZBCyGequj7wkOTQia6gZ
HqLWlR8zWtWbBU4719DDyDcNscvSYx7uOZoeB1edeXQT/MsbIPLxxLE0Z79f5PgWS4f724045Qpv
ox/vo+QqA9V8G/uwNZVyrzGnCxXG0P/L0T+UZU97kd6Qh3Xo+K5eiA1oNwqVJMWt2KjP0wP820A8
f1Sf/T3vVwpWeIcY0bfYkQ7vUb9HYkC0rcy5XN49N/jlgRvbWGpfd/WrIEvYiBS3J/Iflye5OAG6
B6tSZaR28D4e0iTp0SuYhuHPGS7K98eW0/qtYsZDS5tLigDqJDQC5rY0afAgHO1FnZL8mYRgojSo
Y/A7A1Sj76LXUnyP8nLQJkvIx11V2/Bd9MzXJm/uH7aWbzomhB70Ra3DmUrvynNaMbnej/8hSBtc
BUl/zNenbon114ugX+CXlePo0iwFlJ42+ILido5MEvi+mSgjeq84erJE40Fiyc+H+/otnr86XIxG
GIadawEyOR41i7AQrKcmQoEJm/zobTHf81Pkt+2eGogLEn1vrqtoagqyhNaPFfZkLQPqcX7hSuZ5
cB9Ak8Ud9PJTS6Jqgq9lnNM9Atkg8y08SWyjjmJ4tO5tNs9dKcDSA51EzdSg+bqU6plqZVzV/EZ7
o7SPyvJ9JR5mGiXQ1hjGCBvB2bx6e7HbMFQNfy7Ow+eSo+kyXSi+rP59R/kFwZTY+uGjyTdaH9ey
UUHNPMjTMHI/tx32x4itUYEfUDWpeyDO5jz7wngAAXvxILKIasysLecf4Rg/gJAG6tqezzuruPrV
FI5aAzmoeuV0DicRxsK+aLluOww7g11YOI2TNvoiKIB1RHHb0o0FP2V8u/Bb0ycBAntq0Lpi8DlC
cTa3jM1bJ8yNL/rp5X5dyo/hnvwj83dOu8X1cNICAEGYr4GUQKnbwPE0X8pUJSXCanuuPPhs3VzH
r4kVbvprICFPFZ8UqNA8lrcf8hID4mQUL+HF2OMmS8LLrOJ3x49MzKZ66cvP0zzCiT/IbQcr8lvZ
4/cMzZ92h9RJ54szLyFwcniwxg+6G7dOBsvWgN+nF3idXSRCDMRBiPUJWtRI/ls3FNRgT7tdw6mi
EH2bjXgx8MzwsUaFx8KD9jSVwY5aPGcXqgV8qD0la8h9phVY+9PXnjzEByqr4BJUn5hcpRqgKpk2
yPbah5Veik6cKw/dTZgUMOjfNSu38U7pC4WmmqWnZYMr3IKuNh78EFPSE+A2OuE2i5OqkP9Qnrmx
GqRTwn1Ngg6nJYFsrA43k04qxzEZ/vHa4StXjBikTywCWDsK4oQ6aWYO0rUpN7urPuSGOG3uixps
Pvq5lGCnL0LTtQuf23dwC2PwrABwcQ1DpsdLo25gmZnGbQ1X9B1nAwGcfxw0czbNtaPjSf07Hsnn
q0p+cbrr01SdjyGCfnbISZeSOXkiJL2D1jOg8Xtfxdg3xKUH8ZHkZsACJDKcbT/xOOjj8CxAwZX7
jT52L7qo8y7sukpg04UjjtIHYT/KtifHoVW9QkFHDhID89IV5N5sNbmlmlEfNwhfANPxlJetYRcc
DI36v8JMu8yzdPhAQsqg/5ZNuC7r2VSQJwOnny4g7SN/1fSte1FrL37fbz6ILTrGpYOFUF7yp328
DRfVHODARCbSpPppX1BSjh+BZgjvzOjD89FSsuC9mqO+8s7Bz2nxDZSK5HEhGeKr6nPpA7BKiKX8
qxjseNH0U5bAHmXrWV+Xs09TP74dBFyUR2uKBD8oY9FHoJHol8ZMAi1QDcFnb5Quan2u1V7K2xjm
l93Y7vK3lR8m3XjO4vB28l4RvnUZYrNJuGWmweUzk68oV3aGL3s1B8y9uuQfAAhn28aUvFloqkpn
CevarEbA8mLhA3vDi3GVisjCXtEDS+0s5h1tJuBkhLXHQTx1i8W4vCo6WJpCwfnYiXfllCmh4Es9
k2cARFoYNjKaczVj366qeb3I0N6rJQfnJJXmp/VmlBH4lRvWQRemQwrYWh9ii8awDPD58wvGuue1
YBY5m7mwLv2I9WjtycZNadFpjyHO7jdx984mCK3U0jmss0PgkVYcBFWRP34UypK56ab6u9La87Fs
gk6HDyWGOEKhwKcZrOsyoWeuIJQEnVnWkuDUkVhxfd00BjA+IuXveh9MG+TANn6O4Q4/V98XqQQ7
L5grdi8pySGkeDvknxQmr51tkjVKwc2caj/0HYJn68yzyRc8MEGtrFu/wRV87MjwbX3G9z+SBLbd
YOrhuZeuY7QNig5DC7IHfollH4BFONd79aB3BPSgg8EZM8LSy5yWaX1MBz33mzw4YDmblqqInn6w
l1RPc7qSlgSOlKp6phKdx80pS0s0EJoiLmy8VKcvfibhEuhp5eCC0oZ4IcRukh32P2uheGPkpe7G
KUwZXWWg0K++/LJVFLXa594/d+mc1vdVfX21juuPDQOOY01FCnpzzyUTNzcrgy5MgLneWi159cM3
RDx5FLNiHDdq9yYe1Qpd/CodL1qJpFlmTOJ2sGUG3ShT3b0RpI6daTZSDEQ0G9+k9iJqyK1HsSzr
jN/DjL0kflHtmGVdFAON/J+63E18Q1BIyYp+fqAuqgR703gQVIYBFoR8QwAntRl5/Gb2ruRH65XX
/FFj+PjuW/AR6j87GcM8cv2/ERsB1yivpChOBciVL/pRiJroS/nnW4MYcdv6BzIlvWiIJwo+0+Xx
MreoDncMHT2a7vRd7VSmueoCQ5wdjv1GlxKkfxydVBT5h/JnaheY0U7IO8eZsNJ0VC12y5LhK0NB
wd73cSARQieVQ+zyIHUTxeS59BItk8yWyeia35XCGpNCf7LgUOEmmz/PDbK/AxmsjT0fyVJyRU5N
fztigT28v4+xhDHCjp4xT5zjHWb3/Vfk2252n6TEWrvinZjHsLOyOyLyRzu1dKUhyu1pUfT5h0Im
e4A3xnqpxLqJN8uzcPTWoLBEF3EhMKxgkoeYiSJsv3TJD3E58xAYkbblnLnStqEEJb6eDNWqdeQd
hmTBQPKmlo1pE8JbH909OCkkjcDMfux+IgUpmz6yySZ/T4Ae0/Dd7lmfQsIHgQICEo3xcChiyQ5/
lqURjEHvZpLRiYlXIJVys/Ksy368ktW5R21l28CVj3UOc0jl6A8p22rsmuiAgZGSFHQnFL6Jhj7t
FfVLUTqhKhdezwBYxYxBmeRIb/gC1n0YubU/NE9Z1Dip2oGkm2aqc5Arbm2oCDnLDnOXJgkA8/IU
rO/i5PCbiTJj3tLL552c0iRGktXaX/fVRmpXaIi8MWJ3SelnVem9VGSTlok+qUrQqmW25G9Zh57T
OJNTiHGIUQxw63yk1M2t/sXOJRQj1HOmhyMpJ3LMv9BDhtiRgqTsKKSwxl/tDjTwwPwXzZ9KIzRo
WzL0WhSOFNIFEHadF8lw4CvxWddsBxwepTEUcCeN+B/swsfQ2CdAIJyudC3WVzUFgNCF2UHS9U6Z
uPZDxyK0VKnlgurr/iJpI96naGo3eyKWZmlPJJ6KDTo9PJ39FqFhC9UYqsLL7fiqu/xUin/a4vWq
5GI9pE9Sdid4UX+V3d8I1dYju2EwVDQWNLvius4x6SdS/HKfhwyCqMzNF6LoDW5I6eTxcpfMfMwM
4fvQYixpXV2EOv5PyPJPG685jntik2X3q3pJxSDWRZgy6C/HHzhLW2UMvFgO9R/T03zg9HhSgy4D
KQBTI+WcoP2DKrO6E6fojtOaAduzcE6v5rq7rWxkvqC0eYhNKc0E1/83QEipUN6jyD7ZZUF3wxKq
AOEq6Jt7MEwMLQ4+I+5N6vjZlL9fpFRrBhZLh86pHHtN7ikkjsPddpqtiClXCbvOObEJ+QVFnMVx
VuNcfd4t8ucTynSjHjHkdf+KVtfMev0/LHh6XslPVF54y0REAN9yulPgGM5e7Yj4UfKMdLtAoaZn
J+YJYxMMSxJWGEY3DDpPv2hrOBLKrJ7r/GU78bDg8TO9QWwAOiE9NOBbsI0vxCk1s4gL1DtHt9qF
0YbjstJ/ydMZLqxc7yjo20n8aEtI5v88nsiAogO78YzWBH/VlaWoDKfe8gCAExvBhxTgs/3roJeA
3DScb6ftaW7B8rf46UYrKXg5k8cchOvjedjq7M0uTAg+D0Ao++t5criiDRgcDAN64UpDtzw+AHWn
GdTT3DluHDjGVs//0ZroOv0SIHxtbsFAC4n7+3WYWtJ4SaQe7I6irhaJ9bo3H+/IqvYoOtyVlcTf
IFExwmPGHA2ZS0n45qSEz9bbyciMIsGMVGsR/zf8O79YSA0jVeRR5CAc3c7CLX0jVVhs/F1/oo+u
HFAz4aTiEETj9l2EI17zxk1Q8IgG5Ec6EJdu1KIgU/yNoEwOw5s/v9xoxTypbHcEn3xJGrG+Eki5
f+N7y7Mc10vO8PGW5V1NOkuKL22NZUwI81Wl6wTxZ5sCcwPNE6b+bOlQnIwaVkmXbqqS4T4AyIMb
28EdcjBRA/ZzzcuDd+j5Vyo114kXBs+aLhlOR1l+kPocYiNYrfeMkJXam+RvAJP7kTYJt41IMPm8
zJimSWAHn+OlJZnDSmZbGTPk/I4Fuhu6SY3xYp1Bht0qAQhhimlIdMUU7r2oBIYIJuiJ2tn+tqEn
3iWVAD+tL2KoEtv4EvSHxWVcMk0RpUzqYTPVwy/mNfcJffDbjwpCJQrh0UryznMGQAInA0STek3y
fG2gCQRvoHJ+V4Gjy0zlnQJtd+ou8CZyakDdC43KTbfY9rzQOEO69rAeqanFKxqgOcJo90hTtS1z
UbM6vrXHz00S2IC7Nxj3dZucm9re0Hu7vCiGo3c6KDgyWsCyJzMLlZ0Y2Im9JlRwjYIphPD8Cj5r
0chM9etyZ+/zmI0VbOO4qJaZJxvJdC3mo6IAoV13CoN1f0f9Cnq24aFzYt14QBe+cJP7dMGxpJof
BgUWEh/pAzGJvS0WRfh3eQZcaaIMz5U33bXvCVKmhxp9eUl5LNfbCpgVW0zvsGpI5plSWxmjrLAE
hGpfOV7vW/vwIAyTNOAskSuuS13B6yRrcl7/Fk/lNvB4Xt4OU+RDHTLsi90m7GChbVhEvFs03Rjf
KlSCrYqS/vhzqjZ/fXCmVBD0eQtInkKehraRcBOeU/7WLYuwafYi7+pBB0gWv6lPcJmN2O2eO72j
cqul6NKMQCk+cicLnoMKy8of2Q8bJdsOOdcF1j5VM7ZMN0bcaeKIAdfqLWbVbO/M5EbEceSdUVut
e/KUhtdw5qPC7A17UOUAwY5nkayx/HehxLEazBb5v8YFQsO4bDKWwgZOZsTgvnwAY6cDw5G5WlZf
dpWZeC4MKRZz6Tp8S30+bjK+zDEHRaSwvcRr1jbIwHdVx9fiOB9OlnMLmuZiW+SmEBTRmUDMZF8j
/T83GxQOR2YNLSDtHqkfxGYFOvshsk9UYzF5ukiuvc+SHApD41ZjpfZ6gA5A19Zr54t1e8gRX054
PzKkkhqDQMGKy3FYFYWHPk0PUvWfJfVrLns4F0CyE6RyXfxZ3g0Ffwsx73I0KZFF6G83LdtDotxf
0nW3cA7A6ng65rKSie0AcHAot3ZxB0O+8MV4bf1UnpcfEfsqgrwixxS5+zIAB+j8AXNCjtzltqB8
L0wizz8S0dIuwMT036IOjJ/oR1slqesMBK0srtL768U2rdzESHSqv1WW7hSWry0EaaGMYx9TVMKq
hBuIYa5COYtxVuEb5f5KayfcjLCSuQQPLdYkuAX/wKIHCWvQyVzIERTdp4dMtmts7k6r1LZD0HJt
f7DRRhauHkLJ2L/scxQtljmpJF5pup1IF86ULWyRrIWbmNsEMInDGzoS+wBKwFqnl8wQQfkb6zTA
oGCkP0lE1toK36GwLcNbg899iLdDWifrbGClB+vvOfH04s7Lzx/HFCBbp4pWo1tWbkNcwzqmCfYV
e71Nvb7ElcpQTXm3QbCmiL+j0JBsSqDt5nL/8/XqW55c498Xyb27c0XpDANugXkjlkGUgMbxdhOL
2wcoR/zvYDVIB2cfCedUfb9vzkk16buJxfx+vraFYbgf9kwBNcoVLU+0M1tFS9yLRCpQqNsaJpKk
tPVWbxbfgPDhVYvhJjFNnwZ2B7JhOfTZe548XECKvN3I1dzIQBR15H3GE2lgmy4TOupOZ2IZ7XoL
yVYkYmg8VS86h4T7Zu2J9fasIn3SZAUK8CCPeT2yYefo9G0xfcW3qbLZvS0/nlkNH80itRBF2tM1
pyDe1NNlAIFcCnWC1Mga42Njc8vBIRDVPyxERigXg/dra+wUtvJkdwuwDWxQZ3CWpmv5ZEgk0V5u
g/b1WpYNf5tEKWRdEHY0OYydwsmK7LXGEDeMUIXmXWI1XRwDKGEe5LUwNDoQw+vIm/7QwP9GYWQm
qO4PEcKlg64LxIQWwA6ix0PNiv+88Zps+hA7J1OszK3fKJDFXIkoesXIizs/wwXndo0ZX3pEsimp
pTIE7+2eyxkrv3LVENaG/0ZLiB+8Q5HtWYAHpILgGSpNxGtoYWr/Spd+Yqsg6HGxVkTCZ1W3gi0I
hMiFiS5M436FoFYcBkEXkfejMxfH3XfqmUGsDKM53h76Pby+zEoCPABm4L+XKc1nogIQaZSpR1Lb
LqRFB4IsJy7xHBEc2nnKWKkOaERKUWI9k1lNCkH+MySZ0xKo3nJMk7F87QCH1Quoj6KFgfMYVJlQ
Zb23XYIZdXvU2HPoY70v9y8ckfiZb9TjLL6sOw9jVIh5ttFRnF//BG+YTR++SyuEz7CZ5JkdxaX7
NOdQG6SjoiHgL4bRCUrIPskyr1HNbccl/cBDzXCGiZYuAGCtP4EPkw/jt4MJV+270azbCd7KXtQ8
8Yde/7cw3yGFweZcekoyrUoDCQsIfvhatlpY6aP33zmvG9SOyBuH8bKwdios/PFwMQ2LgCLEXmx9
71PIpOqV6NJGezp37RM6m9w86H2M3HfhvQup/Pw/vuVZLHeV6dFXGl+NYknViwX/nXvdmkFk9VmR
Sww0V/7dPvCOGvqWDYbuF6ge8b17V983T9FTxkWhGjOH34lv322fQF6l5jQJNwgMN6QlF1P9dipe
qwY4SaTIvg5bMgodGjkSaUsX/Qhm7w8Czgti7aZv0LlZVT2zGomAf9mGKZVDkWmB1S6jX09rFpt/
rRnevrC/cgpekhgLGrT3MkhLyULZvkHQQitD+KpkSU/LF8jfI+Z+Usy7QA12GgCXkFdFq8018O0E
ENaX+J5rSwyAp/lWPWW8XBv5yGMRkkmcSEDqi1pbOWIOK+0eXzHZTnkViVQKMyMBwPkrwV6uQrMp
xhZoKSq5e1HomLqMmfG91SD6+eSGmaj3nsjj+p1rXG4knwmWy1Y/pr5jIiTL+cHQm/T1fuWcl5tz
/qa8z9qtQSsBttZmKkL84a4bVbbjsMnGZLTkgPvT/tRp5X9csDEqD+gcm3E9RPSgAPejSNIODJlj
/vjwgBR8yyn9FVvKylGqzWSKlKfCsol6Y6ZActbyhYLg5g9Jn53MD0IAkxFIXK4KCLXsYnP5ZFgO
nXgB90X6BDyDL+va6bBn+PF1qHNTT4sZWDc8rcQexGk1ar1rKHLWciaQFzpRcl3UgTk3nyVRX1Yy
eWy7ZVG7snDCRxq/oC2gZtOuK65FT+H1NObGjWUFx/Y7/hEowPeq1GU4WikTvM93Sdgzn4UcG26u
rvgIl3E4glnBdFizuS35ozEPH9bWAGKEmWjdxJXLxX9SUjuWLbCyGZeacz86hV2btMJ3AdbfXlWI
wXeVHCfbgeaf+QQNbNUpNvanpnQsUoB5n86M9z7Br6XMAtf/pjLovwq38GpPcVhmR5gS/5fJVWr6
cpVQhstSWzHr2Bst4cqRraikvybUgtouiUC6PROSDF8QiTts5ZduaBauO9TDi4KYLXa0N5hy7Srs
2Np4DQ3UK1tDrMYD7GLqvuQ2dcJgKPtywu0ETtEXNhw8oIZZUujXw10uTPH2YXR718GDOVjiSq18
HMNOp3WR1EgRYew7tK78teoh7Nn7aWL46PB3I6qhXCvpNi8Pteo+skj5B2Nqzqt+i/xqMNMBnwGg
QLE5HzqRlC7ZqoTA4yICmWtFbR4QPKax24HjVQX2Fgqab7Lj9OhVns2L1Cyf9BpTOdWsNSYJfWFL
EqVbXSpro34WJE2v8topTmn+1WEYNXR4qo7GUZnZjgryuzJ877/5RYhGdsCiRHgY/gYEJlyGEsdI
u0Q7yWact6EMmudszJHFjsWZv7e4U/hoorSTE3+KJICsabfRp9UyxQIYlIXAS107ryhm0UWG9k2m
H2N7Nynx/JNx9r7RDOlLSAw2a/J4F/hvUcOKGzV+zQImw3VXSgqBDzJA0c9Ow9Nppf4GTNy/NB/w
VPNsS21S/n8/G+PddD3D+/ysC96LbvQawhe4iQKXZDXLZoQc2SoVhpSXuqX2k8F1YeuZ00L7nOII
AwHJMOweEsC7P9Mr/5imxmFfBZ9Djee6jSbuUAWFRA/To1FNVEDkqyJJG/qRzZjksdcnH2x++Np2
3WSNddqSMLWgYQB7nOWUCmVTAVADmNRkDZxUujBvnIZRZYykvE5K7u/fr50MXrmvTp7CzO2JRCpS
vzL2MkZi0L15X0d6yFznfXU8hnh5R9S5dcwl/E66WR3AzxAl8T96mP9OLSxSlCciqGGjvnP6i79F
Azwxx3vJT0QipRSv0pNbBf6Px+sF641qVC0ZFOuqWMjVOSKE42Rjkf76fGMTO+2B0MYM5LuFhhuH
In6MC5GJ5zAK/A1rRgNpyb4BchMUIKbUKrsbwgTZd2I4S130hLtcq6JD+YYjAQLdhtm5ZCAu+lOF
J3orM8PQpQqHUVcD39+38D7myCcDNLTlkATe952oKazXzZ8s7odXXao0LLO/ltpODWEOszvbJ5Tf
bV39c5m0t7Si79JL+HT3a04VCkhlSawKXHNNz94AeNKQdgOOakFYw4dahjDtU+JEr9wduBjlqJkv
K6xfBHDyBkDPBeCNqw3a3M1c/cpzd2aCcgxWXP9X1K+Q17RF9/yv2+6K6NVbkR4nUDKEJDlQBnTy
6En15iY0qxUfOUsvsA0bfeI7nYD8VMP0uXFF57VhyOOJcf5LWycuAU9ZMb3W8yp7n8XwVflyx4+r
BdJZ5EZiq8IrE8Qm4G//caB6RCAkSYqBDhnkhyIWTV7X6JGCwF2ahhjRSdwujOqqHIgsvp+ffx08
QdL1eiuDhd0YbJajqOk/uxQVLXOcwi1KtKy8zVf+idRKXmBh8OwCE0/rzBghekX55Zb4FRMsTsOY
aS2QgmtoNM7xwRP3fepEitqd5TEbuLO/L6rt2unXuUH9ny1e7Tp6asdlhpe2LM/PB9b0b4bh0jVc
wC1wdrGQRavLAhCkfkv8KPO6MGacnu0dJaHxbCc4ifjz9SQdjqCj1XQYkTThwgDOt2Nfbaft+q0e
Jjm8u9OkqLhUVD2fSaIW/+f60sH7RQe6BPk6cs7ZffKO4PrgJlypzCa+4HGTPetVrDRnro7DFPNx
j+0fLY5wSD0l4RsL6UZcafXUq0H/cz4xL9YEwxcfGMxuqqnEUVqsniM21bsJUDOti3vwuwdNhonj
LVBKr4GBsKOucJgg2ItQvwJV1A9v8edpIcxAKPjDxYGWN3GSRyblwzqGmLhuKljy+GmLJNgiR9+Y
vIaFFz4LHZ6zxt5N4TYjqt+4oXanmj4akIvPG66RYiseYyZfoQLiziBQMwQQXMotqb13lLosjmGF
qU5DODCPoEzGWyz4pkYUWy3iDy89gJpitGjNtb7zykHaWbg+RFXiprsv07DpL4L9rRXggq9V+4yr
sdwwqolhNJwmz1Ir1QsWgiMIxQd3SwfopzmEtF6+N6K9Yo+ctwsAgRrHVxKJjA0SPca3PHtjy0TD
iPrqoeQK7k7KXc/IHau2bpXVA52KA8joKjc8jzWJaE9g4pW08uY0pQJ6dw7kRI82XyvAq+jyiC9e
BFJq+KNzQzBc9lvd0++uN6xKi0gw4AebsWeqs4HPCj1I5EPv5jhjsu3uVqd3K9RQlP+F53hHhBuB
kkmXUZJs4RkOKpF1S0DSrnNm8JqweTtPNnfWGLGkQPb5fMZZRzdlxh7LLpsi0OfCwYpWTX9VEmsw
1DOTNaXyUzl2nX4MwhuKOfCL8csTFTPi9ELE/Xd1nNQQwnO0x0nu8fM8UVnd5+r29bf4UqM0QPjB
JVHVhoHRNVhwtSKpBF3wht6g6cMjJZnNK1g/dSXzj3hMp+jx1VB5s2GCmZhCNRqB0fwYTl26Adtq
/ar0HJo78hvAv46WiTnc/BK+ZXfr8u+RA/WmK1nX/1bNxdL9+U4dpL6DB8sqz9RymnXsjobG3mKk
FwcJ3WAV0eiteZBJdvhtgqum9bWU/EckbWRc6w3yX8HDmxF8F5FvwL00RDrUoC7Sv9BGcgYaS0HB
WnWPnvMLyGHcpqiUylaTfU6rD9IyBisUCPPsg/H+OLqytqWlGMsEmjN5LWkui5NAUeCLzSR70Wzl
Lke8d3U38bEdvYCMR6icA0GOYadL/X88pxsV97D0on2BFgIdBBC52Qjbw7IFNmkHwBe7Cpzvh97R
aOQt7Ncbz6TL6TEL2kJ6XIr6WC0LlcB+JSBuBF52/bMRHybMKQjyD3f/PyGMK176RgUKw+Ct1kUe
69Zozlpxkqmd6WlySZ5x4npv/li/BQ1lfMMaoY2riug4O/T9QwguyAkrihhpEGBf1LsBAvwrGbTv
ZkKfz9LJJX239BYNj/8P+KN1lfyk1c9xaVuiVggnf/7xX+/NQgJPuD7Etjy7NcBER6POmBvWBr5H
6a307Ss4ofe2eZjszyot1zseNdwDkkee71kUIZG6QWAPkT3GQ+PbUspE3zDJk0UOIUodXmLfTK88
fSpaDYT9tfyBjbI0+HRmx8aoQdCxc1vfRWzrHMaTtYM2qn7jDm7BIhAvfYewtXb88suXZlapQ5XJ
MFUuFZVObUSEiYan2M3CaBHvFx0LEpvw2nImNwUGMTmgvn4yc7H5hcd2g+UaNIumRKFY0vqMR9L3
o9yPB/AWe5hNBH2FznOzsFrApCRjZvdiCXxZOiwZUK0AeDua1hl+Vg0y5e2sFYxdbwjiT9VuOa5W
7Jqkx/cghC6jyCCscjT+3GJrTCYCTSSeAH+FjabvmiN7Pr9AhyLUTqRDZpJmqC6BT6hOMFLMc6Q2
v/2uvlE7cZZMqJycC0oDgWHr+nFYxJCZRVNVQIc7lihKMLpUbRJGS0XSXtzQF+y3CrIUCWPB7IoG
AnylAW0g6+t1iPys0oQ2/cFnljmKPnSqqM+mjNk4y8BHSlECmhkwJGlkieSjIaKEmMS50cxQMti5
T+FaO8zvhpuhYJzDwgVcAIGeDUferX12AiVeeyy5hOfw9IYw31v44Xn1CNWN1/d6v5UrDt991gvG
7FJL7F2I3KHJ4yugSLNPVamY8z0yBDgVNgTGoyEcwuT4ixvY+NRXMBV8mM3zyuQpMxMMsVGNcthY
Fad4/QY8GkC1qUsuH68s40Uz+KBAJG6TxG2JQ4OiCDxHSP6Od8iXG5LCJjhiOdCaiXSgvLFv3ikg
giE5Ub+psI3m+RVAyhpV6zr/DpmWr9kfnlVdzpPTriGGCFdTGaDD2GlK+XjM2+IDull9aqiD7ufQ
kfw7TW3rfO7lKGg9CVscJKV8OLLBuVotQfY8qFBRVrzc4B7PaAJoN3TYBmBGtBkFPEPtUloJA661
54iH5e/fS84Gs+xf+r9/aTVm53SkQRU9tbngvuW1lyK/J4z5REa/DSPIz3fKhum0L5QPRkDhNfLQ
fhXcF9o1hCTaOkVHL2MQ2XMjGTZZRcKGihEpVf4/hfPHcaYRgFH4DArUUg2/3+dl+P+CKIe6eumX
vDxECz6uO8XItG9od0QXbk9TfmUm5bZ5+DaHFnWpphdh6iL/GS2TVcIeQe8Dk9waDMga1i+oNtX2
HZX0qiMYZwwiKItMKEYdZZzVXR6tYNkZNPTj2tSrDIKPji4VqjE9Z3S+Rbv9QtQ3xMKJmSSWMub1
tNgq0VYlU+TzsswgdzhPvCt4ZfgjTLs6fxIf5HU8Il9D7keycOui0N/nufZWg3gcqGpNl98qSTCg
ITTm5Lqwj/B6thmHvCQzgqEQqha/2Sc8iJ8BnucmVIpBEzrwBijkfPeskMCJYHmKm3RbYINLqyOZ
a3XNj/3OCk0nBH870oYb8fh23N8BonX0/iV1k4EOXPr7owdGRKq5XvUEsQzIhSzrque+doCPKDI6
tPHO8gXfMJkrj/lIBwg9EO9yna4vrSS+RFwthx67jsilJPVeU6Cm9vC3e8IINXfLZcUDyPsCuumV
MC9h8cMxfBWIzkj4lELZ6ACBY7w+5jM4RJJRQ9S6pdNp4s7Y4APeXdD0oDsfdLC8jiuvqFurceBJ
6aJK7G9IvdBnsO+LXurtIEwQvC0y9h81ENBJ2bdZp+XyVobVRbM+fw7pma88iqasbE/pczdMB0iY
ZpFOhD7BJRBABGGmKwHm33gsJ5rtu8c6jytR83waaET0gnvjoeirWaYJTvfpkpo+I014O7UKZSS/
1aToehnjVsfnyZoLTwm9JAu06GCoyD3pX2fI6VfoZ1n1vwMvdt3ROOWa7qJvaBPmh++HGoN0hIsI
z2KeBOPsSarhuuupL2GYyWSmPL8MlJhZhSYLf1Wyss1m+4r2SChoQH9EfRqITrw5g0KxmS4/NDfC
pHFEdFXq8apiJ2U+xfW7t5AZ9U2fuyx71DbVlVJtKeZyWovnxgnCiI3HOyP0/NleqhElb1R3szKe
CYr76BDZiXPtncLyuTbBWqdbpmjSAelXJ20sX+5jEjbZFb4qRrxzjOazoVS0jHxtg2O8V70uLQTB
mAPv4p2LvH8wYOpaDDwt8fS64ZJys91mJc02i6S1Ek6UNxR9iPrk4oysHY/sOZ2MB/jrSVZKQ1+X
fwxwYTJ7vUgckbcyoWDzWAy1wUD2z5hretQmJbkv4vPLAAi/CFiWAGUHN52HoYikl5yJML95H1CV
mTeTUq9XLFaXd/uXCB3Ws78p7+nyKiY5pHACTKd4tW+MVmtVbmTzvRPA4izpVsaEOtLdWqmxEkh9
Q3HblQ+V7MbijTohm2krmqT/W0z5cUHtzL93xd+7kuCq2X5mi9RbkGFPAouJ+sV7x3sH4N4bGWXN
zk5SkfsY9yX5361yMzKf7qekt9dodiwZh0DMgDfhcQIJJ5kmCZX/OMJMQOLkCf41mMzNLGzSauzQ
rno3s9SmZMDRP6eTmfTN+QVIJNRQHH5s2qlLsZCbbgQI4tSAFd+bZ/wlncMnnK3A0shNwJq3uZ+R
L6FH/hk8hrjlELoOh09zZKvjjuUxZS2mosTSx7/P8qdCgUQeLVVBa1NuFPaxS8j2+pZz5EG89tEG
OIOgvQ6wlotn+ozxFvwKKgmSvCxY6ZKUKVm0eULl9pmYzBldvSTfJU8jcAC63ENL05R8jNtqwUqU
JYaj7wJSTqD9/lWCfbWJUPYz1a0mFgyGehQ8dPIo0GBtIJiuLQ76yvEL/yLhywvwIPnVTrNP8P8T
K/Io/5IipGA0FsOERmFyXgkG2jAOVggId0u50wQpv288MoADg2J2X7CXXP0yarZeDvfl/z1SUjTm
suPPK8IMBfGWTdMtluI1wCttj/iHVahE/BBamRKSKzOPTD8A79vO8epImhxgd8K0EOZZh8CW7O9X
dD7E81/rabDAPoSwaMs81+HYhbZLX8twWZJ9rIPPbZBmEAov5+HFKsmVjNix33IN4iL8F+SjUyts
M9Ea4Y8jzJFBdFtAtZaTHK5nwIx8Y0eUojQU3tf5dI6Gaft38w72gtDapuIVA5DIa3i9pLS4S7M6
97xXgyVihp3SNpXOzYp6AMo4Uo1d2dKp1lchY5fXfAd6uLjNsRunLzJ7i/a/7wxdXQFSrPQy4U34
0j9qqae3g8JOFMiOdJbGA+FzUAcQha7MuSbVsUdUc3YbqzgJ8azSyfxqf0tCLkvaE1uqIPqxLbQR
OXfHp9GD8R7fUDziiv6abSpCphY3yhUxUl/Qy+lOC2gCQWqoSlmY2Y6OBE9sRnb74To9ZezgW6Lj
nEwZDSaMQD8gm/BWOG6NpvOTz6FEEK3khzIjpw9iNl0JhgTdU8Q/I/FWbz/KmwWDRwjA9LeWwI8T
D3xX4GhPLBiUG1EQi3SRW4xV8RLd+6QuzKoTFNayI07HrFE+AEan90gclaQvPoURv/uZ8m1r7HAH
4Ej3it2h4nmw/r7NvydBUSh542E86gmSo+nRQ5SUGyhaj97ym5DrSzmDBsuutcM3wdCtukriJgxO
oIULu4nxauh7NPQfUaS+tGNuSROv+IoHA0fPS1A4MKAkQIjsyBgD3FPyNrFnheeCCysrRp6tB+K9
BKZ2ALb8+OezSg+ad8XaQUOQmF6Wd0RbKSGB2rmerAijOOZBaGnq57OaD5vOCqgPzXVqDU9S1e6w
zJAwmNT7PWc5aH80qpaTP6dr50BYxavrroAub6ApiCp43mSJ5yh14Nrpi3y1b9j7HbBR4wu8cIb9
gY6WWIkQbrau7GRjwmxKpjJgj5CC9imsU8hX8FUGBU0OxsVUBaCZrfdC3jpqBMh6R1CwFqHUSDhV
ZbCNfmm20lYNy6rBhQS7oCdlkZ1dWgn5Coej9+OzCON+pBbIgBhNRB8FYWQg4yDVuOfTW+ko0TUY
kzggzhcP/WO54PAfyMkkjLlt/26sBEcokbOr25t4r/bhk54FFUV6yONiLdhJx4U0+pC/5LPB9Njw
vzDthDxdmxSJervV+52dP2iVtLc1iirY3Hg5qkanC1TaE80rKdHO0k0TRuuCedQRBCyr8fy/6i2/
zIBTWrwrASWTyM2E8ecDonrH6jmpr8HS9jLREvatmSKP9ur60BKKjCe/sC2nF9SWFkoJokLvbpzy
5DFaDzt+pc7Xkq6QQEMeRNUx/uCES6tl88mA/FMbN2iJ/GoJ1WoUchBxqHH+X+fZ/ZwnzJ+h2AU7
nhh1pptGO9bJIu+9YG5VbPWvnvHi2VWb0Qk8TBkbuvEEvMwpk++n7bRu23tBLkzwlQjkkMrubmM1
XgXSaCuYmrjY0i6LFj4V5qk8e2K0I7ks6T+cnroTT+T4RKc3+YuR5p+kjrK+cLY0urnw5QMIJONn
TXFQok9zYRTQawFW2EBOmYbGHqaKa8nLVRZQ2M4zH6PGMCNnKiUKUYl9VU4z/9LVxBP6Ak3z73mN
JDN5iLxcEo0x/qd+gHm8CLvkW6a2NReSj3GgKvV9koPScRnYcYf3VTf3qby9d0ewiwRp1dMW/G05
5i+dCoAitcpY9QLfhzAhVBo+WMQKgN5a9KVb889z4l16390Fi7524uor1nJZRAXmwrc46jZ9lzaH
LL8nPandNHYhg7iEguSQxOrGH/kGGmnh2mg2vsBjz85epwwM/HVF4QDhNxLaM5LbfsSbjK6MdrMj
y7p63yG1KDN6YskdFVrwnGE/ubDaQcFtMmlZKXsqnVfdlWasAOWgJ/FWBc8IK8B8tUqz5pKJGGTL
zPXlTushMzi5rc7U36K8P3WCftl35boby/TQCdT5TlqdhkExkWmX5MpaLTsDnjD9YnoPMGZFniOY
hU4BJggwBn2TL9VZzKORuV5d6arrOxw1GWaJ9o9gvgnWzVtrG/CQsEVWLLqZa0+2/MbGX66iknAA
XyxrOQYQxn7OUtllVOuJGiVTOv5JNXOHL4awKLl5BF3zaGwVb0v/Oj/jsC9RLzJ99ZDjVgKRRnPl
gj271bZ+Giv5cvjF3z0gs+7Cg7+e3gAozetgm/H1m8syVrIzSqP8YtgFf2oOb0M2or8WAVs6wqE/
k3XBdEzU25Bv86F1sjPWSnQcGtOq1On5ld32iBr03WnN3TocHY/OGm58Mv7/a5usz1MCEr2s02Dp
jJas5acc9mN4BPpqvlAK8wXBioefxCh3DXYDXrF5ev3cHk7qmiByfzARnzKv6h8k727ktWd0By0h
tJl2ORP32gobpDwlBR+rn+7QP+Gi0ZfvG4VM5oxVg/7daHHz9UdqGTDELCHGEKCyE7UjEDqG2PJT
hPBqya4HpThmrXI5SU5n7LyxPbZjDJUDHB7fCkHMZk/UqLoXyRpUW05ZVoH66avEFYUEe2CvQZdk
ICjl5bk5lpLB87g0oSYGoqiQr0n1DAXwDt7vkzudtwDm4t9mh1m9eE7aoULIL87mM5EhwPxitLV6
88scpOmN3SNt0kkW6uWf9ljn6OvE7ZqI02HG/AjBIyTaMwKE6LqN5afqfGLTCZAbUO6TzxhXEOM+
uRUSYj1G+E4nWj3PxTUsGk2iY/6ZHD+/jC4gLmtsO2z15OeHXlw9UWd0BNlm8QQ/gD6tNrH28997
2UG0r7rXMENpqUAljKwhLP0qQ0FrXlIolsRduGKegZjSIjNsdnqjFukL6PKeuupaFXgyJElRYdAR
4xIDyRfTR5CPsN1UA7gMcIyMwC15lmY9paNDFZrDyUhBO0fFd0sqTI8NzaGkZOYSelc+skjM/IsT
ruNwhR5T15eunpxzFU71yAn9j+Sa1kpesqxoYi4ycdy9QWJtZ7Tup6/94RlKv6SVwZBQV+2lkIwK
f3C1tBnCYKAUKopyhjegV9hDiCvsqd9HE0NPIAq/zmPObxwOYU424BUVDDBkAYDIeO7wjG9XKe30
zf5Egr3gPvY+C/AOwqIlqa5gWCWdFKHIcP5UOzl6S+1M+TZ85BaEF+j8XUc7BMn3vKY0QZ0Flwhi
40anZbfDlybxekLp5Ujf1DYpkZvT90dvhE0tdaVCQkPApNbvrqmtezbdtg44BBsJ0ZKMr6z0YKMn
DACu0yvlOxZS1FeabhhjUzj9gjxFBOg/jUGc0YC2Bd+IW4NpuFdanQEj9EDS2EXFtMqfaNO4UdB+
Wd9Ut0ELmKXbXMt2xI62M9lmIjiYQzSSK6wruyzW1UHkN5GcmeOfZF8te5zIaY/X3bHo3LHWy3/k
HNPB5WP5F8kiFYZQo7x6h5SPwN0Bf7FoKKgkwKIljG4DsvLBAWvHJPr+6v5HXYwzDz8HgAtO2+/T
QNwqedSHCfVkOTfwBtJ2dN9nhT4nVE4jA/hzjb/aj4SMYnRxPhGGLQwma3lUkX/cbOzqZOqlwRci
fF/QnTLKbrC2hdcQZ1N1YTHRUb6xGh/RNsQMZi5VL1GCQ3AwBoIcFweDpZ7EyxkeJpZjKceuht7l
xRjvmDgur/re4tgGzlhxKg22ygYcLgCt6y1oxVuPaCr8ySG0GJoEz6+IzM5tzNiSTvYosXCHrEvt
YNlaF/xP77MS3ZF6RDhmqrx2BQoc6l8uz7YLtBFhvmBdBV5bI1owYs2OzP39HybGqQNbu/2NGamV
TjfLM513UT5nsMS7B3rLARdnWVnvrqSiHKQrJ8qGNPsHnSsyZuyMhZRtHeHf9+IE3DKgp9vUXsk1
nnmEWIjQ9/AGiVLWOMS37qb6qH+4SOhefMI5ozgtGkd4AqL9ZSQUcSvRnSoYavQs9sWpz8RHo2zp
yRd6ahKYhjhHJC06fPc/fCVliakE85D8KTw7EIWWc22e3Gp+nQluUWjYiIraW8Kz7+n1X8or28PA
Xbgy9v2ZtYl/Xr6jH02ESyUdCpkT4KtRyO2TJYFqkO+GODFB58VJlbLy0315Aie/rFBShybE7pS+
nCH6trmsGiWDvLlCTCNJOlPvRGDLBcEFSjy8XHi5ZB7ATa9LMwZyPkcYGcOG03JSk12SLx5UkekW
FOylnY5RmAQus1IZqkYr07FFJ6oYr+JvqkgZ9Oj5zEGLm/WjaVA/r/2rYIlCdV2cAJ4cAO/kVgy/
b5NA0hVJPiAhuhw1hZOTDBpbkkdaqfrJMePmmg447DtppxD7ZDbQVc8EAxDxs6Bz8ESRnvUdySgQ
og4Bry1u2UaceFpPEZOm0YPI3qWm7DfCgFFSwKi/5GG9XY4o9jXYLzIseU4CEwZV4KN/Edk0ax23
I4kELLWU42sYfqz2MAsEbAIKiuApC2TMkAgSc3bxoKO+kRtSYa4gJwkaYPY9m+14LnRyKtHGzENL
SXRZTwcfYTr4BMKzb0FJ67IgvIx0hv55oZwxHKx290v1/TIs0jU36mZGZEG58WNPhPd9cT5xiMbC
nKcKQ0/8ScipViDZZ3rFyotBk1Axc8nUSimSfEwnAXMzYmN9qp65WMGltaYRewoqKgSPf2o7LgpB
EgQA7EABV9BheDO1LFUxTh5846kxCP8jg5vTw4J6rjBPoLCL3mS0T2gxOrJO59ugjlDm0Jke3aG0
LtQUvsIAFykc6+SiGZnpXhTbzSiv8RGoqDs+1ed+n/VhaHphzXPsMaY5ndqnzqrlisJVVwuZ440I
8ILn29l68BmpEpqcu6KMu7QxOlxdaRdPeDOjvsFp9y9c8eg0N4xoDp8n3+bJ+OsrgN1g8X0S2zLt
V5kCyB8VDSQACVFr1oi8qdPtYjWm0g44C0XAVysJwtH6TWKKYXUR3eQpOQ5tit9k6gAjAskrsE8a
M61ZAcV5w1JZPTuvtjEUKuClkh1l/t4qmlzpueaHBZvNB91InJWUJ4vh/3CURIgNgnMxtyNAI2xY
ar9c1OOaqEMAwxaMY7cxHQTKZLX3+MZaqFLkLHi8Ic2Vzx3TdtjmZfDztCcrUT/IIp1wr7DF0m9H
EYSKrNOPgsiupHzEz51bEjfQhRmHPpCaO7eEjF1/ktktFHIGLgzJ/+ZPVm+CAg0hVeKoorK7iyid
Y9FQySLJsESP9AKEmeJFIAtSywTfLGEMrYFaXq1iKaXalqe9pcWmCe1PY4ZIzvzj63Cpu+zvQ/o+
+uAAW1pDMaIwLaLgVSZFbHlmH08VU64FX0ARHN+lMInqsDgKlrX6p55AyC+dVmIQsziQ5dHbkihJ
aGULmk+dDxk0zT42hXfTjRL51EPY9d3wOyD0RU6+EF9haha5OaT0EJaVjOHsqGID0Z/FMAmqG2z1
n84UVeJzqgQ9KVn49znhLL+R1QVEpA/Rm+RjBodSvT81Bs56VDsOa77qqHg+Jm/xV9B6QVQF+kw5
X5LwOY4eDVzkE8IPShl2bjHK9LEYAgnMtHwe7E5UCTTVmFM5UiI1DKOredHxcVeRR3GL1Aug5/z4
V7m/u1Gj+DfYB5hKxijEYjLkkj1AjiLDcbivASabxdChe90jzam23VOZPcSDQc9Zo9okzBaX0mRn
VvfernOMLVGZ7d4O0bHcVkAH20UPdbOWtG09xuHn8yeD2URK5wxCsHHKXBBkGq6sHm70XbbAw0LV
x+xebtQyV9u0jyNWEglqtdVaiCUct0T8SSKgrH5biCwC/OnvxMLOc4edEfBFzBgb6TR52/pSzeIC
uWVIrrnghc3g/O8gyJ6mBAXYzxDqlbKYvvfMlBac8xEVAGJ8RCt2B0XTsP9fRygR9gQzlHm2UC7Y
m0oj7BELOtELSIUMLbVgZkJjPQsgGosSxd6FU56OXudfDUoLvBlKvjnVkiyegh6P9HTdH9wzYtTj
2TduTptoh8WnVwI5At5j/D6qPwLQa07rGKjfIcSKh2yOG/ukfo1G2i5dxYVlYVa/FUx6MsGEfVb3
bDn7deRbCTXkjPbjlEYKaKHcAvko9mON27LVG9nsB8M6IcidnMERVsksGF9vKmJxlqC/qtSLsI8M
i+HY1PibeluUazVVyBOfNVyziWLgIxMf9/18aQ33ACfuJZw1zNOkOfoHFfx2DEQfKoqGEpdTrGWL
Wt0nl2phOD326yrTcmiCadOPhXGI/vdFmiGkNcopGVBuzjQIs2IG9TDsop8R46dgEHYcJcbLZvaN
i31p7nvNhYMJxxlFUx0ZHxOYhpUjaQ3Tpz/7efr/ZxUQZLmbomtLSNlI8fjubJl8fOnPaY22YH8d
Z39MlvaS1+R6EPWdSVbbCMWuPhj2X3lrsNGJnDebMTN+qEM9BMEtc0jF+iutP4VmPGeoGmpdxtxo
RpsvAkILqWAzRNPfZuTNTFJPe7J5dxj5r533yWE9tvoSEkXo7ddIklzaKFvKn5QjyhozjoHOE4PL
I6bbHtHNhm65pojfupefSH7Y2QP8sFgWpQAxJfNGiaNPFkqz9WJmei9QDnlnLbD5UiOxhWQdc9cI
reJSY0aJr9fNzkfZ1s4OJV/sBdo21Rpxjegf+KhYpyeyOmumxAnZDgciUmCdJztP9aZav4kDaLXa
w3xP5kVH9ZP/UfP1+pab3WC6Mty91QaiiPPBRR0GG12o6SNFyGgt2Z6ttlFf9wScIPaNvoLXVUXM
U7yqMbGgXIEoe0tLMpaYjo/D4zb1CGgMuRjmT10Rs12xIKcan2EyRw0wCgVARa8xD4VDOh07Y+ih
E+/ZA2aXSK7MerJ6L7bwT4rjQSdWOLp2Ohds0QhAfmD8ipf+uWQEHFOfKMqO38DKPaX9wAMKAAl8
xHL66fCtdmOhPOc36s3ShPMWONioNfcy8l6fItwGsUfyvnrYhZgjYYSUR5oZwKx6SrGndZTOD/6N
QkU+9PC7wIBIwbA6PnGObg8VN1XA959aZzkVognThMhRMh7v1N4e4T3TxuF59qARtZa0fht+p/76
fdMLCKsaoiOutZqYmZcow3/2UUTFBUb66iZhM12Rlb5BTVEKhQqM5RIojgWse+i4tQTS1eJcthzh
US5uTzZ7v5iknYFgtemdfCV2p4vgpx3yMALaWe6DOlKeT2vRzlZXXR0Xl4cScN5jSe05RZr5FLuQ
BkK5rAcS8ndXCkU2GCniOELH4e+d6I+sjvhc0KAYXBAepFp1cuQODN8P0N/mnuWyay1urQLY4O8R
4oTWUhNEP5u6hqHjRlkweU+QyMMwCbUIXds3vrLGBw2zYno42QjzBePXucCXRhkc6QKBsEhTd0Jz
fEepxw/2175cTptyOWoFqkbXKpW2Deo15PRw+/IulhsKneoG4uMcpOeR8WRbmOH6IDwaSsTDDsxZ
v8fCErxXkFzXSNzq1beOsQAzl1N0LBENYMZcFCs8pxYVcn1SVC63DQlJuCgtpi5MCS2QAM6dS8Tf
n0AxYXjbCiH4LtnSHSRp3Nb3r//iD+ujWVOUaM8wo5ZawcDEH+UReHTn1EpMqHhPe/OQsroBcy+4
bDXEqxRXHy/hUu8+S3ajZqysbWWr1+gL1YoQLqOkzBUkCATNp/w/PANQOp0Cntep0QPSVBFtMFjY
RsobVqtZ7m16mRwvkvrdZcpAlWUpB7FuRgqUvx4naR06PATs8nsJEmvyDQ0jkhvrQTkjJxvWQX8n
Gg6OqylS/5YfyZpTrBhA3kzju8nHfsbS36UnHORvyZomW7LKooqfgTrDgJxnIdnzzlqxoYQU7wKa
c2CYdTus87zKZfT38SyVnUezbx+wZeSewEvcN6KxwVacPKQiSCbztWCtqKMAulsyi8eSxluk7RRC
QMpvs3nNgMcCUd/TPuZwaS51j3pD6ATD96F0/2vTqHazB/mjjiLTlbDkus4BrwKgJla64Pjbq7yx
4HFKZIIBuQ0YZZSNXFvHS+Rbez6/Oag3kiAXlKI3wzB5Zo9HlJmAQKGrnA7fcRsjWK993c7m8o2K
L9IWVLOy/Ab0I8bKNZAHyaZkz2plmFLy+6OWyZ/uCSLnYNBUr7Uw8zRG6ZiGkuF3BGAIs5Aj+DVV
alrVmYNutMSV4GggV61mlSokb4UlMBXf+91/BEs0iDQRsYxwTzLyjMwqxlhHrW+uI/E7vYG1LnUk
oN+Xf1YPXF4jUV7A8OyNFk27J9NLWUXj1DSD3jVVB4Y/383k/XTOLw4E+o6EUzyjSowmOUqdCuYS
L8AGqCQCLD4Sm4zjrQpWItslAmF/t8NmfSpVcvg1Oma19Jg73It9dyHQh6lBr0ZpQT435i3HPTDc
4AZXcTfP0yjdUWu1fEoMvu81qEE7ukT0vq9nkRUSz5kQ+fi4RWsfVFlcgaB2z5NZzCSc/o5LgfCW
3OltGfyHFMIBK3TnSvshcFrz3fuHSI29wyP+n5pE3h3xLEVniD9Po/Rp3175+ody6cuZs+x1hFHU
JiLXJVtOZQM7ctg04stwrqBJfFwawKlC4iRFP20CA0g3Rd18TlvTxsMA2dD6tzWyIeN9FwHiKUzA
TX3GVkwnwFDOoLgQGgKwkPOXmtaUmo8CIK7VeeFT5bJmD5KZBoEj6BWSWDv5SNmfG5xTaDHuWnOI
6EH4MxR/ALBveI4uWuWbqpy/1X73JxXBN8lxIzn1TprEbDCQPR5eKtCu3w/xHFpLC1VbkHavpBuV
/wAIkoOL9TCtzApL8ctUOW/lHApTx+L/Z5IX7Wj4L2mO95wDQrYAbX7WLsxxks0hrIXGX/cp7+z2
bRBAMgVrqEkOfaiAgW8nRujJDO4VIX4Fm598JM+G9fJsaJdxKA9QvEviX90OGMmUQAxNn2gzDzlM
F4kFwDiQOZVW8bNdR+QC2DXhqhW1p+LGyGxESFbj5AVwqbb1G3luGsVO6ytXFXjIaeiYwgrQv9PA
het0LOO14FLvN8z+A1GsCWZEp4cXDnQRzWvTUYExNcnoOtFanOzOvGdBIYJ66buiUeDZoGYHY7jt
4pWEDxmN87WzAiPb9VpB9FhfNaYX8FKJhLseWVgoEae8V1yxdiB3en25dvJcsnty6r95CMLhrJjK
Ui2dpwsyUuM+SVSf19hQvL3yeJX55rrkGLIxxpm7WW1oziG9ybVhNqN8HvbIikChTajZzUel31NF
XWPwZNokLUpmg4OPlBiX+/I+3XoAZ/bk7A/QjEocld5KCuJtMRZfX+nUyBsOBsTg125OBKKzFAq/
5FjN1u6BrFfmxQJeD3Tqd8yTFCmgiV0fOJqH9g4o7lsvgAWiQJ1f53qe93dth3DeNOdJyPLQxr+Y
RszGkcdZvC1O7edfBbdxV37MAhtILt47QD4ERZOZSu3zX1526AmaKQsbMCNHgft1ww1KoXOXUJCH
sAnpcfTGdOwgUtHVBEe/Nhj5zRzuo6w55W+xxDSBtiItIVunZAxi4XzRR2EUhbZXhiAj1jUIl1Ku
OiTWeGpupN7gZ0bwTB9sezLTEwDRLCPnvOKyx/2nYu7kzIgJVpYvb9WOIBUBhx3e/RAN7jm10dYO
J1XpqGhvVhl8OnbTuoVINKHZTclj1t9KZnIrxj+ELwY68hFgRIHE7VYo4FjUyZ1U7ua5xkmrLJcK
FH/qI+kpvGhGtmgXab6PeptIl93dEgACTz8qeN3QvRx3qFKsr389JT1kB3pr+mVPcmgJabK8tgGi
ebSHH0JWsUwKdqSCPK09QnjTspirKUyyx1G+/ffAML7Zd2ZZhvuXx4QYuzSdbhtdiS1MpF06Z8oG
zJPgjjitKM3cevF8AQxZTW5tGKbKgjVs8+0BIPkIwaal53ItHJpKOQP5dzzcESmnSv8F67JmClib
R7uOdwRxig//klg41mGjSn8oguzADzdRoVWc830DwA6vhF1lIG1NP7nlzc5sdthyX20VJ9389Wk7
U4W2mmDyx7qD8ZjZ+a8UnvztvjBBt/Iw1rsig4j6QS0Mw/jmM7L1Ve67Lewbt+f2q/18cq4D/VUm
PKC63BozE9spqSFq9vE8oJUSNf2k9hlgNN3jw6QH4HbXZtC1/MjYqbI2U+XU7Q7AZRfmHxMz/8NV
8o3ZsKuijO4vw52HfH1TXMdoCNP6Xkesy5sMI4gYJBmRmniQ52j6Uw075dF/Dc3Dj87py6oH6+xA
AvP3xr9CXJF617EAQQ55/XX4ziaQ2xyHWyTfidl6lTHhr7dU86qBmJO6lJPkz321Az32jWIzq4g9
C3m0hxnJDjDcSHo2emQmBkkOW8vl+TTljOQMkzxQl75rbu4UHP4+amC93tMixRo19MMjYsA6CHse
uGvLbO8Ce2QgWhGteg5Q4Ng2zsiVVw3URCNw/Mpfm6tan9/+7g0IhMocPtOUj241F8mr95jhvyJQ
zgBF3RXwevnyI+dx1Y36rDpY5HOImbLIxMFXAScmePU5NgOOimJW4KrGjTvfp36nRGdgqdr2ICV/
9ZQGgHMcYyCI0hssU9zybwLy+zFPhxl3juPtF1wRZc8CnTvqTbe3DtPaVURXkazFAw4kcEm/llGg
Xkz3L6M6fwl4s4fcxHme+7snGUucgsLj96eyz3xSIYnh4i7k0iBeWFWp3plpktLZZ4IUoXjmnWDu
pmVEm5hEYdGmGC6Uc9zQ6k7qqxySRaNWVg+AUKbA9mLt5rK6R6hMJ2Y8Fea2hC+w6yJGLFgLmxWT
c+UoxEiu+Nr1qtoUBwTmiw6STNRHheGkciAjI6zzMRBND1LMZxP/nVn/IS739jP51xf39VJ5qBlw
8aX9kLclqYgQq8Jy76KaeBJ0H5hsk1ul9msH9uus/4bXAwzh+Rw8vTvwq+fp91sJMsaYbmzecoR/
O6/vX5XKI7O7gM3hMXASSeuci0WRGBToFmGrb49UXzfo9h3WzBH1EQ9bvReYJr8tJQMIJidCYV1t
/IoEahOBycYBwnWUaWbiOBHG4IEiPB7zqELdbesL3Vqe1YbaMh2RTCShZpGxGdw1mQPbqc/ACC+q
qxoNMxW1ni8TfRJPwwh4ggxARqJ2N75v/o9ryCuPebsxmNnKFjUZVFkr1VtXSkfTKwVsNXj5JJKE
KRbrr+4Q6QAdqn6ibaNTJ+25kBnc33Awx1715sYe+8UyGvdD8n81tuPqQhCLsJKyHhc+1bDeYchd
MTc6CaO5VNWqy+aQhqSGHS99w4iicNFNYL9G962MDmc5yvb7Qtoe75JrZ3J7ci/DpOH2eqnr+Klu
uvrMv5oqCssCz0IZne62qQk+y2S5f4EBVw/ZL34kVaAzOZ06W2dlKJPJznRGmlDqvLqeBQ98eUax
SGeh/OddpvjtgJqIaM0C6ExGBeXZCoWhGx8fWetRAk6w1R8DaAJysHp3XnKmu9LrzbCLoKrX248g
elmmlyIS9gx+Mfo3lTjqHkH1RQfdnWO3wEFRFYAXNCYYrFzaFMF/n4jBvF/q2LCqI8lXNDNsWeE7
RH8P7jnWR+loBBfDxqbouCEcP2BCCFuztp26kNTtL+Wb9M5G01/PFXS355MIOiDmAHTjmsmbVIN7
Kyanz05bqjxLdXrTdmFHWEYWL9wXXLjSoA0gEkqNwx391z7795gU4iDlc5J4XjSoIxCDTTNFDtAp
kVibO3LGNG3rof7PT0N+kEFEvrCg07nSlVqZanK+8Gtt3oh5ogylkyD/m06QlcvmjbOJfb/0NTrw
vD6t8HHkSDIJmeR65+mcMusKuSCDY43Fqfqzxl4lJfUCDZc0Nz4hPPJA5l/3hmQDb1GlwF4LH1Ds
YoxJkWYJiCyLAPopBKHsDr36+mW5+F2Tfqa0TrSISAS0wSf5rN40BVWpTcocKOkMMJuwewW9VyZv
lFBM9RPIG5EZyuR25VNv2Bx8bNVw0qdtSYebXhkU/fSnBl0u3739t0b6hGzSDGHKhomhawjMUDWJ
Fo85C6OMJJjjRExC7JRNnTHSUdFbjaiw8pdoyyaIE0K6DASGMfgFgjZprmUjhGHBSc3+gCi5LT6t
51RK3Mg+wpkoJ3IDWfZZSCvmeNqn8eCGnateEXhPeFke64/s1Y84lOi8H1Fdt2gNn/unc991ofzj
Zf+nx4DhilOqoSBKaT6sUIS3D1LnC4RxvXRVV41RtM+eBJanwgUAKsodEYQBbsiaEgn/yNRaReFQ
SW8pC4YkZhKF2WHV+CplR9UQVr5Jz4RVUPIEGD3VqjK8BUFalwnmNwnfLzb0da6qSwmX44uXbL2w
UFhKlDhhX5+kHcjXTOVTygb1CK8eY93bBhVGzyk1FUheeWd6WkuViD8dtsEO3rOmPjOanxaOJLcc
DK+YNXCp80V3AwDkTBU8IJzNnouLjxb6KPLfv535CRcKm+unGq30HTbwOqOaGvo07Hums7FZ+B8/
1SHgMfVLJ8IViiFzD1j03jiZlTL3W/lL7dgSBmGSeZVJa7cYzIJg+lGvXe+us7PNF4Ok0ZJW7bvm
gkFN3kcPplrtm60HgdjwAkzT36tuVATghQwIGbYnwd5t59TfbJGCNf2GUyxXBJ2kjBufwi7J7E0+
kvf3lefx97dpI8fCBGg8vyglsdmbz0XqBWNwO9eT6TcqyQH/c/EAP27XgP1a4EGZ8XJ8fcLcusal
lqiY32FT3cS/2BDbUn3TMBgTxlco3Fs8KEyiNI63pkPFAhLBbP5mj5pjVwdTog5MF+mm+xMMKZhh
+cvutNVTmEL5OBxg1AFF51x0LdBFrJP1Ysjsme306IILfc1Rvo6zIfPtOwTTOONQ4255V+8uQ4E1
81bzGjOed0dQ8KV20do8I0HFpOwl0Q/C4mnDFlCy5C5NwBeUYZN76fnTLwBei3GPJGMgy+ttb8Re
ygNSTLZhpuyCW7OPqSAb4BEB0qEH12GbNlfs5KbYy5/QBTYqVRLD5PfIqFPpfcBA7K+fknRe7xj4
0ednDSkjYbQdulyP03EdSxChaOtMF3RsAgaL8PvH7ylUtoqVIWvknRU+twiUQC/E3kHqJ48gwKp+
Aghj86FQGfrLKmLmjdaYoe1gSXsSL2N/2fM22e95e6J0WnAglee8CtxZIXIy2ayg3tXmmSlL1dxF
p2oTB9ZtK9m+3/OCw7SdfjARVojUDaqNevsMw2yh2KFC1DmvKSn3Fsg+J+mCQ/z6N0Rcv/H746yP
lpq0kZINffu0C2Ddyr73VX9v1FeitGahNvYmbXQZ/sE/SymwGaNV9FbVO60ucho3HFpRiXk6PYWv
PT6SAa/NKx3oUha6CyXXujYDB7tSaZsEAZHgk0OWye7wC1n/CIlQ+0FPBMkHyqlKHE7DsbeIE2B6
WJnyPIqJuFbMnkiFAm1rmtngUliKLPTAZGqDdwN6YGE7mqeO1NtfJUKgP8v9xalu3wsxXBb6eSj0
QKZdyZliKmvfoVfEuLFpVmyiaPsGfWwqIEX/p2gMgpIZXwHhJEjYDj6hLbN7mDT4PxsxmrrvdoNS
gz4jIcktIBxKb+tXn5rwqc8Fk1pxxl9bPSJNdsRwyJXQ5YvkTYbq5uFpC4wa3OPKxXvZIl2dcjhQ
5B8dZ7VLS0rvkfJSj21tbiLAc60mMyuYMuqXf7BG0KRPR9fm46yUQmKAc98aCeWJ+Qn3r7qVNSDq
hIlJn+YMBXaRECF8zlrx0ifmepi6DClRpJ9bsWMF6lCSykwwz3GyZhNsq9n1K1wQMetRiEYpJ11P
0wJy+U6ISb1dMRI+dieBVjwQtaGohxM4ug1tfapMNvyK/BpNDJWreF5Jw5T2/7AsHfttk2+vr5Kr
1Rxz2f1tO/6pNR8/HoV5T2WJeF7Lw7tGOvxr5vuTfLFrn1IO0jVEUahPWbfeB8tjF2VKABQfoHC3
eDz7Wrn06A2CoWjaPsM+RpeqBSFt0Z4wQOszZpb3yyJeLK1bAXcBPbHUQ66rHT+gmNyr8Iok/43D
2hiPf5jo8QqlBTkw2LIAw0OgTQFl+4r07YMydbZPc4GfXTxD7ie0VcaaRpglV+giZnTubHt6QFMd
zERBA6yYQoANMna9uLUOmrdVBs49TA4eb2T6YPIbpPJ9479rok5Jja5Nf0pwKvE/mOHaBwzfO9ux
yqKf84ZlqUzVWxXJN64145praZKyoFRWzNH5wJQjmSrnLlObAxUSKghmVGW3lAf1rSKEpPCBoerh
wggIdPsuk8wA1B0gLEWEiGgl8MEqJpEWnMmro8URXC0tfSWWG26IvyPT6NEFqRyQ2OzQUzqpdCBu
3t2U/1Df8fu0a59dNGkxBUJOxZr9o4p6oCB96WNgg7P9EcL9eq9vfQup1NjuJutC3ahV3ZUGYfMr
mdsNsyQ3M9+R3jksBR3amDKlnhdUvwB9o0EV/h4q9sImYjIa6coOmYnXFCu7NRpoiPEbBXIRKqf6
u0U6AlnM9/seUUEgyoMkSiOULkxK5DlZL4B3jhC8EJ4oelfcQiX67InCUp1+tDSw9qU2SysRW1Nu
GmN7Nf8qqnenjPOXYrgpQWK0P82ohCtejvHsCD+kFnzyF7zHgpU/URTVgYIogCLw4PIazFXw/3kv
tnSbWotbXBCZfm+CTjJ6cpVXSv2hDifDTMk2kuNaFLG3K/64xbEXPOQ4d/b0fqZ+2V8pPeBxDgwK
1Mu2jtZw2nIRR2ML1CUW2UVwpn3kkVwOT2P+6H/K7LFMyXh81wAShecY2ECq9erKdENEO2yx3+En
KAjzhfjwm93A4sAXNAymKtJOvW21kRRImDdK0NXnHtA4Y3k6tO4QCLaCZAuXTVx2Ne7qpN7V+Exn
zAkH1oAq3W7LjXtlTlD31x88jyKQL7sscIR1EK1F3Mx4QLzSkf20CK1psyIbogae90prf8S0COHy
2I/xZeBo71sC70zozmtJ44mf6RQD3e6m/6j1Z7NJJcFL9FIDO1wRYWfn6DZWWI3sdScVsqABf0nZ
XCUR8rjZT3QMAH8vcx7w2xmMV4Tl1fNz2LTIwgPhwq3QMTIGk7ZXHVOCuel5xMZBFXtUbMSutmZf
NykWWo2JEiAlysVtdsZvuU4X5Rqt+/9S2yjwTXpkefc701YYxkyC1wahOx6x0zvxB7JZK6VTsY7a
R6vRX5Jxih5Z9ROQu9QnGWK4DwAc+kdtGEzYW4gpa0+plLmrQdSwfxplIvNXivz5bNiVsKI5Ozna
HdZ9XjCLyLi/n5FqCZ4WJwS01qtUUCL9Q4c41G3oFVk5Cciid3C2r4Ocj+RTPs9VMWFZnIExFxPx
M1nqrWYLFsdAgHAq8DrFgE7N8ThNvR15Z1vCXWVIAhKvTQn3OWtQB3HBclYgnnfiMo9rj7Ua+pAv
H11By5REkcizH5Gcl52Z+oIKnQrzawsnHGtkrcPYMdy+Qj8irWlxn4HcCKqTUM7fAhn5m+3j51jY
PPdZjzefTqGHvYctHWN6vQ+FbucR4Sav3W5cMb9BAcfOP4VoNnFNv7dLfJ0Q7Xq7CPIYGulIpaeV
CCwGaXblCXqrplRMHi8KhdelzzM4D1jADUUpIOkSKfEpvH4pcexI9AT3/wFV0wIKC7C47LMZDfSn
kvGtwJ0Zpv7SzcVURqgVnG5Rowq5RFDQCtjZkfSqX73IsoD9mXUpU6CAsMwQfToWb2if91CkeWSD
5ygheZUzoAxaT9O7e7WAeHxJwAOgvzvguw4qt80BQNbeacrnxU8GpdhRoE5ZXLhirG8syNnzR+3R
B5icX/ySyFrmSUlfUxWkKMHzM/CpNjRXHbkOXwRKa1aMTN8/OTgBto5DoBjHKZ79aIWXBg4k2mxN
6puqZ0KlKVdSTSW/KH2F3WHsWQEKBOuPjZiUAiwvgLFDZnydq7Ksh7ajPT1ngoelhScf7p6/Tx4K
wWHV4qGWfx1XjJiecR/P1mJsSnHKMcXdQXmiEuE3RTA673bOUuEx4uzhD3x4bro9XmEkQRBDlCcQ
0/hgzpi3HPqddm9fk8f7H0YUP3CitUvSLhI/dfmpQ26Xa5VkLQjJAcq74WJAFQajk/pupMlGJX8Q
mN7TM3YmRzlafiXjxlsk0UqFuiwBROuVZyYquw/KALXiRcbPAQHrm+yMDqjxnxA6Gf93VikbNmdD
o1o4SiOgp8ngdPo1HC415+8/+zCzQNUpyhktCW+/VmbUcw0TqI23hYLrZ0KamVi7ueaCfpzybagR
t7KZ7YVb+aoBecj/hvuhjq+DChJ2HsmZsW5jFUUGbXxWpfnC/LLSgSGODWGZvWfbpAnsoFLtLiMy
6jVgcV6xozVG9NfJAXHvZbDanj6UYSItaADcwEzoZ7ypeE/VWeqBZCuLtQeqYcy7ceqBVMVZVZJy
XSXrmXMefTOiY6Oj8dJn3zGk8O43zFIqX+G+9RSJvkXNpw4WPekWIuqOtuNXGhZIeBl49EDyRSV1
29pXfcOHU7Ts2xkWAB2JyLOxdxtDeypCyoTQXMjVdfrgs7AdHFeKDKY2B1E58C8crOfRFmel9h3a
piB+LmbJ9XGMU2OkwA==

`protect end_protected

