��/  ��Q(���]G%�B�C��G�1�*�$�^�Z��%�������[�Wq�~`�	v�.@s�Yꥱ��+[q�~�����h\x�W�f��O�盁G{b�]���i {����~.q}<�	���`�� �)���(�c�,��e�طɍq�޳n���6�����������HZڠ�I��Ƃ�b�_��c�hd��N��q�f�M����t9���཮�l�rF�$E���`sQ��<#��:��嶺&$��pwe���bcz4���@ 0�]�@�u���˛�-���D�_�j�C�ba�dߕ��Ori���yE�fU����{\�e��g&=0�ܝ��#hU:�ȗ���C~��@�Y��I=�'S�#ԑ�ݿ_tĠ�ai��5��C�!�,܈�Û���tW�҇�T}@�~ˏ�Q������ͅ����3�'`PW ���w/we�W���+@3���u����\��YD�їR��ȡ����U��)�f�sg�U�G�G���rE~���
����˪��ϰT"�mH \]ÝB�L�D ���#Xq���D���0ObǿPh���#I�ֳ(CȪ��#N��kE�+�i���*ʧ�_ap;A^�\�Y�^5Cg^0�����yԐ]/���l�,jzJR"��7p��ٮT�wm{�as\1	
Yl�J�꫏���;˟�N �9/w�햼�g?"��9)�n���@e;���e
a/0A����!�~ʎ�T�ߋ  V`�p���|^Jl��P����x�n\��\Ljg�]�G�&.]�W�.�o�� >S���_,�hH7@xGe��D#�a�y�� ���
F}�R9R�H�fџ�Va��$3O&�]���b9�5Ǝ�q���Q`�ʔ���p���qbZN� ��PhBnyl�J(c�m}���]L��)���M�x����Mk��Y-�[�ֳ�}������D��a��nN�i?���~	��}Z�����V�\\��Z�tN�:h<|wY[:R.�
�I0/�XmU�*����MR,P��8@�o�=��n�*�h�t����~�;��$"�����{t�ũ��/�Ă� ����1��=%�Lr%�BO��	nn����XζD���}W��]M/����F��u>�b8jy��ɇK@���`2Ҩr���A���1n����.J��~a}�k!���+�%uEQv1��Z�̊�/Y���LX+�j�����bx��Gڠ�]=\�5���΄r�m�����j�<o���vs���FPG[�7�K��\�R%�t+:����Z��k�sq	1'5S�)}9�l��A�����Џ� ����JpX����p��8��_'��{9`;D��(����0;X"�j@�1���e�)��c�۷t�E�HԦ
"��=&��	moX1"7�������Co��S�|24�������\�T�
����lv�N��Ɲ���VS8OI���%�02(�t�q�P����L���x=(lԔDi�Y���]�R��P}"�I\�C���/m����%B}�_�C47U[{;��U�!�	M�¿0�s�V�hr�����(���p��_xC�o�=i^(+��a��·��<��hI�伿ע���v����z%jb���2��m4H�z�E,eTßv�e�s�W�b,N惪xx�W���x&��
t��d+HA	���-&��|��m��]j�
��]�����ɦȐ���r�%QX�I�����3���;��>���E��=,"���̦�.S�x��x"c��~�}��@�1vhjI��R�9L�C'���Q�l��+��>�$lR^D�P�V`��L������b�~]�#'/O�h�Q���*����e�\�_��]��� 06��>��%��v�����nT\�?J��2�j���p�8�CK��S����dZa��e��D�
�]��ޞ#I%�	ʯ�a�"/����9��m�"+ ��ա9IX+��_o��{򶷂$�+�@lJ�֋"�q?�����f;r�%yS�t�V���`d\��2Et��pqjLC�i�p�׃X��}$	�SLY��m�;6��+5A5N��.�c�ņ!	L����˜z�rA/+w4��*9�K'�����7K����XD�\.[&�Óx|Rep��.�,g_�3�è�Xnf7�_�Ҫ
2�D���]�t����C�N�f��/����e*����9��I�+=ֆV *~��l�.V����P��rA ��a�{dD�,e��&j.��s����B�D��5m�3�
�60�͌�j�[bC*�☬� �������+�"�>�R�)R��v|�>���y`��V���h��b��y�&��fF��8��U��p��܀����1|�D�f���+]��a���.�`]�JN5t��\zk7N��@)@da��u�"��������Xu����+�{\��+J9&Xr���]SN$,}�r�Q�w�����9p����'��"�j&�1*�z./���Q����vP�U'���J�8Gվ0fS��{#��r�ãun0������ ͸�<N�@иl�O�C�z���C&�G���>P:�p��xdٷˤ�0Q�sm&�.�AH_��{�z�O4�c7��Ⱦ�nҌ��:Y�c�����)�y�R�n��O���j'n��r2I�El;E�YB��#[�H&��=��Ht�"�p��)y��.�o��p��D�e�C!���H�y�yv�.b@������$�iW�i#kS�0����T��pO�xF�>JNCz鄡�nFZ�ý�E�#^�df��+���}�S4�:O�w3���V,�J�x���[�9�e]�>�Ӧ�MVs�<�� �!�^hNpC��eް�u�R�SA�\�V>g�����Sxi��KY�St���~�j�+���^E��'0\���~���g�R�.?S�� �ʣ-�fK+\ ^��G�.��kA�{�GZ��n&8x���0�;=��[��^r�Ey�vc��?qD���|7M�LςW�Ϫt�oF��7j�J��K���]yM˧6,�t�DVw�x��@ YC��,K�:7h��^7���2O-�w�#������';��(?��rqpi����L�/��j�gz��G�z}q=�zc-ח�5�� ,r���iH$*V����K��i��r:!��R��΀$�a1��!�
����Z�&~5��B�'� 0��@B�|;���-�J&e&u�	R1.v�����f��+�.�U�kc��^zQ| ]��rO�h�@?Q�l&��1kb� ^�����`�<)<�t���Y�d��h�p��1%�Y:^�l�[��ٶ�5����l-~���cM*�$-y�~@��DS(��L\!z��o�­��8N�~�Ղ�ڦ�47���CvYjeN�{�)� �X�Ϡ4-8G◟�@��������͢�
����G�3��ع�X�^�⯃t�{�IZ�k��cc���BN��s ��:�o���=_�NEg��#�P���-��n~kP�̩�,��뙕���>[0���Z�7Vु�jN=a��PYKK"��R��/򯦠�X��O[�V�B~��IF�k�f}d7�x�ϛ? $��g��!�y�z:�]) �r�z+ 
�C��v��)kT�w�4�h}}%s���<�I�AlY�(A��D���I.���݌��5���!T� �����ep����X�71�ͱ��^o��B
.��M��G�@*�Vzqff��c�9z�K$��a�7p�5:��9ɺ5(��͢��]�F%5�����������F��D��LD�^�:kR媺���_T3�����nva�$���E�ږw\d�љ�'آq��������}��0�Ϩ���\�'�3
� �SD�vm�i~�MԑV���բ�I�� ����2�~�o���fQ��ẵ�)�Ce��9�6sRU�����yҹ�U�_�9j>��E�	�L~�K�%���IHѽo�]�]�%�g�� c8�A	��VL�(
��A4���Z�)�*������v�4��e�%5�<R�[#�Ϣ�lEXY~w�KH�����#�6�5sL�A�!U@
 Cl�N���ip5\0ԓl��p�t��H��������<4��)O"�0?y_N ��x�8��3�<P��>���Zc�qqK��j�<C	!e-?CA.��m�1֩�Ap�d_��Χ�Y�J7�"��H���Vq�����+�tn�?&�C�Ҽ3~���,k=�+X*	��W�6��	L��r��M[Li���
��W��6��@�IIɳo��`���w�N%����̶�uhJT·ԇ0v�Up��۹�`֍�*+9|;SCO,Ws>�f��fa����d�� ����"u����@�|�d�أ�U��7����h+ē�v(Թ��&;Ah&2mם���<��������v�+i��V��{��M�Q��[���]fcAT)��'��$���U�<����e�͎��C�1��z�z�г3���ZS�����G0t�,j�B.�o�aI��c,I��I���yJ��g��׮-��ME�����HJ@<�gG�e ��wN�n�l�ۻ  ��~�LZ$�Ja��y5�[�%N���
����I�Y��W[^�b�)�0ʕ��N���#�a�W¾�s���M�cao��53��qb-(A[��z�;�]�������e�5�C�Qz@�W��rb�>���2��k��IYi]L��[�ai/�G6W\����y��\���:���(fFНc��-�`-? )�my�Bn�"MKC9I!~��P=�y7�`�{bdL ;P\��)$�������9�K�$�2u3���8�8��E��ҫ�'��@:k��M�̪�	Eq�҅:C�8	��4� ���Td���:_^�~VJ"t۲E�C��}���S�Pg,�)@�`���.�l3Y>�#/V��8>o\l?\^��+�|�����j�)��`0ʔ!����(ԅ��k���*VBNG���?��8�$x�Y�=߉[/�o��>U�������a� �]���ë�F���a%�,���f�������|�p�9�3�/��y�'ڲ����ȥ���c�$��.:s(:���l�*�4�W֢�O�4~�-
����d^���yW\��hx��~�8񓔈�A��e�'[���u?r!)9�]�#���4�d�gv5�{�j����u��p�N�I�V����0�,��:�&{�G$QE�k8��.cS��r>�F�W�h{#�{��r8��Y]Dj�3�
ڶ�=3�"09�>��9��"�f�!�#�S�E�>� ��E�s�,J�%^["�:[R�f��U���'��-�!���ُ��ͳc	��/R`��ЋprV�5�Hc�5�a���c�Ռ)�h-����@@aVP�~=oiq�6w�x�m~�W��(�k�G�3�O���>���La�V�2�>G"�[�Nes<#Α[�4nX¸k�u:�mz-cH�\��sDv���u��@���w1�&�?I=��쨗z�f5���[7��rj�1�%�v�Z ���8p:��-��!�9L��Kk���'K"�a���q�.>[��q��/nk��b���2�.�r���gp_lT��i���Y�C���yH�|�n��:�=*7�n+��3ƒ��m��
�8��{���h��rq���Ci��s\W��C鑋#6՝�:����p���ġ�(����OE��z��CB���R3�^.1÷�.��ڛ��W7j`�8g��5]�j|���^5�-oY�Re���'���]��|�sK��^�"Ȗ�/���U��L]o��8Iy���t�n�/�E���2I ��%Z�b
�*��{��G��}�L����|�ۘ�j���Pb;:v����ލ>/y�"}�k��}_(|8~�u5G폒�Oz����l|b\T�	/H*L�R#��~���Cj �Xw��S�|ƐZ�NV(տ��J��;cl(��P"<C�=�f��P�����d��Հ0���}2�Uih��h���7ā/��T���X�n�i�z��]27r��]��-3�|4,�l�Gǲ�ۤ8��[�t��>f�����^B�>-#$WІ �e�,�O�������j��}��z9���*^�ׂ#dB��\L�j'C�J����f���:�P+�DP���Dl�?УM[����+%�fD��� �;��3��?kkݺ���D~,[K�墱��D���#W?�՞��� ��7L��!	eG#�o"��zj����"&(��J W�K|���yγ'
�o��{�>�� ѭ�8Ҳ�=F_�ط�3o���Ə�K�dt��2�l���BZ��-f���  ø��#r͍w�*{I�`���	!����z�՛���X/�i[lۧ��c�)�,Q�I��F[,(��p��g�Իx���.;GH��?j��K���W�.�L�'c�y���>�1�B+w '���3��n����-pN�@i!�/��L��H������h�w~_����-wqZe���P �XKs��:~D?�+��HO�u� ����8�ҳ��j�ƣ�R̖;�0a#�z�no�I��Y�|?���"����b}�_�0Iϒ<)�����W\�Z��kx״=�T>#�>0��{4��vg|���[�Q39�����q	�XY�����}V1�_�������{ע`�=����pG��*�j����Xn�^ſX����������#��H���֘{�M�aSpo�-#O����1�c4q���Q�dA>�xC�Nn�� Z΢:�|��:A[H��CB靑�3ο��Iu�j>a�/�V�y7�[9���$�
�k؋ބ���D��F���X�w�"�P�X���^Ts@R!�t���,�Ε��}�O�8�cY�ijk�)oY3�ڥQ�f���y�ܬw������FV��ҳ������B�/4}����@����Lܡ�)�3c��u�O�j�Ӟ+�����h�?'���\�qm�@�e�9#�"%����l��n��X6F4����s�T���F���o1%�bwW��3��9��4d*{5}��]�%?������4G�ܖb��t�]����u�s��4���&�J�ib��m`h�\B�+��|k�63$ԌD����ޯ�������n�z5��������·0F�V��М��rx���ں����#t�	O�p�:�qHZ�dS?~%��A���,�-w�:�膒I�F.�lG5�}H�t��:Ɂ��tz���j[�
�'��ȕ��� ���l{��m��Va�ڱ��b��S�d�e��:]"��B�I=R�<�`F&I'I�˷�p^�+bJG�b���
�k¹r�I)~��LLxL-��c�;

�IKyH����3�w�C�̾�{�n����KDu�@]�K`�K���3��'0�e����Lj��%�`H��-H�p���&��(a���W#�[�{r��
����JR��HLZ�]ؼgP�:���a0���L`��J<-;a���{�s��y�����U�>|FS4����>r���,'��qN8{�ӓp�C:�}� P�w��(����9�R��`0�9�����P@���\F}8��o
�?�*l���Ƨ�c��O�m�!��3����n�Ȼ�j�clkPO'�IҊ�[p�8�����N�gr�	([�pYX=���f���GR Z��H�1�=X��:%- 	�H���gL�e�,��a>�,�6Ig�� T8�!���8L�8x �]�a�M�jv��� �ޛ���
E��҈�ؘF)���f-�r��!	�"݇pZ|�H9�w�x�
ޒ�26�КAt^
�Q��'q���Mv4O���w��I��݈����Q�s�O�q,�P_5Hk`�TC��:�;ٟQI_|;����g�@��5]��R8OA2�Z4���������f���[|�ᾣ0u!��g`kL)·0�/�ବ���zf��̂*W������Bv}R�(�߼x��TS]�5h�$�nvU��孺�:&��� ,m!<�i���w������廯�p�� [�R�XS����Щ{��,�ɕ[��A�f�c%(y
Mb��ˑ��_82�ۃ�2�*�����i(�%����Һ��7��u!�I7���{%j� �oK��Քy7-er\e$�1W��-�مxo��ID�`H�L����X��W�~�5�
=�͕p7t��z6̌��I�����!�x��U�u� ��i뽜�q�o��P�K81�����[�7�|�j}��X@�c�p��d�2�7���8�<ʃjT��n��sl����mᆜ��#
w��j��a����-"���5�%�v	O���ґ��eP���_�َ%}�T�VM�� �޴\�%�#���=IJHX�;$�_���4�VkOM^�ό�|�W�fc,Zְg9{�r���s<�n�]o�VzA�lZS���=�iC	�'��)b����v�h;[���͇�q�N���Z�Ƭ��dbl���NĠbӟ�ʂ*<k;���g�W�n=D�Y��d����b�U�ԶyW��"����tr�Te1�k�{.a3{S�Ҳx�R=�� ���"��7	�^U.zT�=-Vu�D��e��?����,����,�����Б��`���J�
�W��w�T3�[� h\߸R1-�]ݭ�^4(�E�I�:�Zd�}d��^B���ƫ�7i9zו�BI&c�]�aܢ@;��c��Xr��V����ȿ3�����5�2|y�!�G���-�c�����*��HZ��ij�3]�A����eL��c0LU
p!&����_M��S���Y��kެ�i��{�4�L��^��G����.|��7)n�����H�I�O��S�Q� �\p�Wj^�Co�5xY�*�x�W@��`���v���EzW
U��&���pώD4��x��̌v'��2`"AE�9B�cq�7�8/����j.vvK�Q��9��r�Ŕ7�l����'YNمh��-Z%��H{�1�b�+�Xn�D�(+s�����{��/,D����.9�1O'꿌c�S�N�&ؚ�X��D�:h7�bm�	8!ŷ��lF�r�!4�`L헪��tB�<�di�V�r�]�`�]��L2T{vJ�F�����<?�-�����{]8�����:t�w|�mֺ; =��͋�6��pa��j ��9�O#p6tA�Ô��i:(�dE�2Bu\�+ϨA �\���7����&�H���zx����+J�`6��n>���^��褃���W�/�pۡ��5��ϛ�Ԉ�����lZj��[�Wj���w���!��gq
S���O- M .���..,<��Zֹ"w?-]�eԍJ�(}#���������1�ʀ9뒰z��y/k���فi��u�M�+�$*�!F
y����I1�4���] "��N:��ֵ|g�'}I�m�\W��=I��0��}��}�������n�y�2"w�!� 2zh�^8ژ����W�b+�X���!�ٶ"Q���hJ�fU��,{|�<~�|"�/��t�9;�bTf�	�sV��s���e��l����%�l��5uo��R'�x7-a`8��䑅�S��n;����O�|�����<��=�D��\G��n�o��Dg���Ѯ���tz��SD~2Aw��~7�� ����+z��ʁ^38`��:�H��)juc����WS9w"kW����2��B��U��~Ո�as�O�2����c��h��2=�sb��/��Wʈ�f��ݤ5q7!�靺�)|h.�_��'滱�G����߇�nmQ�`���{ &�}6���G5��e,�j ���i�٬'IK,�yN^m��j���N*��t����9uоw�G�rE�ԥ������5�7��9ס��H�l_��ɮC��n��2	 <5���x�r\�#�1f5�~��jk�{�[9���s"�ԑ4���י5��4ʞ�ŝ�@S��!a ��nsA�z7��,�c9r��ǙU�l0-=�,�4�O�?���]L!��`Y�lt�kW��W���xa��v�/��gL=�%d�s�9Ik@j
='����l3�B
�s�F$�O�^�m��Ds�.�|!�_�ʋ=�m��������!b�Ww�U0�1?��_+��3K���$�=�)
̸P=X���� ��vM~�;_�s����8>L.Z���!�����E�\턟R�񑑒�Q�D�W�H���D��|2�u�c�a��ͪ�j_�#�V��f��'���=��>Lެ�r��?Ƚg�1��O���~�����5'�����lu���B;K?u����{!�������I�θ��B�u�)��ǱL�O�.�X#U�f�
�w�����H���q�9�E'C��c��r� ~B�����:PR�#r*��p�Eh�0���u;.��
��5nJ���-ZLi��)��wi> �a�L��J+����Nrn��l ^rL��?�w���]�ONO#�[<P���f�m�����"�Z�?5���K-�;�{�O���+>����{zI�;���:��-�'g��o��9�u;G��z��x�@���=|��t�y_tl��b(ԭ��0�,�����X��d^F���!�}��GkzN�6g���E6Jm������&�1�V;�h&�F��eT!�#��L?��������@�V��:6ڋt&j�Ԃ
U�#���MT2�@�b�f�W�c�� Y݇�������f1�ӛ��)���{L�)��G-�aDY��j����r����6�=�S?ce@�n�.t �J#����)��n\�J[3�<AQ
��Wv�����XMІh��8�'��_Oz��1ԅ �p��[�P�������U([����_�S	�}�x��տ�����̔ː񠍼D�]��I	��>�%�8��[<��ݶ��P0k�:�F�@X���2Y�4܄K�����"����q6Xx�[�4m�Cxȋ".JPi �)A�F�	f���njGV�?A��[���ld#�ސJ�p
����9>l�S
�~����!�z&����T�~L��1���΅a������< ~z�k����>�3��x3.a��H<��{d"8'�
��Qh���"d�Ms��%r��y�8m*�aS��h��I��y�{L����ɞ�2�K|��k�=�����&|�����5����*�پ�3�L���B�K'���@ �V����!?%͙��/A��_N���a0�D`���+j��}�fl��R����v�����6�&6���]"�@��t��1
�.پo������2�-�TkX]����i�z����5�'U�	�D�"�@�xػ������������
j�-�I��I�,���f��)�t��I����I�{a�p@�(�A���"���t�{nf�gg����Ŋ ~G�ݼ�
�n�n1����U����]&���$�^��l]�C�ܐ��V\�B�����*���W�\(8��/~��$����
�%�v�=�}��K����#/��v����/���x�};�M�巛&x�O�M�ԧ��u�m?[�@0ƭj�׏p7+����q��f�*���hH=CJ�����/<Vj�Mp�X����1a��.�
 �N�$�V*ɃW�L�ffD�X��dRf����M�N��B�9df~���F�}'dX��� ����qȟ�g;��2n �8�5���S��m�:':
�C�,�D&5���_�y��L�o|u�?Ж��`�_�倂�,���=o[²��x����Лg�Ty.��c��~��= ���x�m�!Y5�U���x\�A�ʔ�o�0�D������qzq�X)��
�h��`�g*IM3$�1��m���vS1p��4y����1F-7,">U��\��D�E��J�Y�Q�%Ӛ�<���.��ت�5� w�M�h��;j
C��b���C��e�iWu���U�1![����{��;`B�.>��o��1��w��`3}@��f���Q�q��,txC��f�i�\5��@�f�⟝HU�ͭ8l`�>H#�c�&�ҰV�
c�٣2����PC�fU���a򫚹��ӫ� H��M����1#�<vM-��Y��*�.mb:�T�&�����.�����i������:ٮO}��P�ў���!���,�~����vn��K��^�VD��3���O�N���/~���oJ��P��AO���1�'�U)���N��a+\YE\��&��L��h+s��ݜOW�n�!r�F�r�V̛�Tǔ�����3�q�"��o�S)�^Z�?�㕒��џq�M�,MӁh�M��x[N��	\7�_9ѴS�ǟ�J�[z��"�[���J$g�^�J���Z�A�P�=\�n�ʆ���>�>���s�"����6r�l��Me;�d��+t%n�~ʥ0C� 5��[�\r/�Zg���k����V��*�n�nl{v�o��$H���G��O�ӈvo����� J�6z�gM$�Y�`/LLv�>w^z	����q����;����A���Kඖ��$�ߝ� غ�͟�z�1�{ԯ
�� �M�Mm�̗n�qAxN��rMi�Y�j��I�5�5)�8���ꡞI����ٟ�D�����>�Vo�$J{�a�\�b��7�fb�!b[�JJ7k��=�c�ͦs����uy�DYL�_I%��5��:7������+�u�γ�/Pk�DdNW:'%�E��.bu�^�e�+��j���]AI:�b�	�33-#�uѹ��R	������g��'�d�Y0c���g���&��Δ±hH�N��#W���|է�Gl�͔��-��m^�ȳ;c�ܦ6�LS#'O7�*�Uɾ�)��߷F��3ק�ې�Z?��ǜ؉��%�4X(���.�C�����\����@�b7r2��>�{�k|���[���=J�<Ȗ*�H�I��y��֞���!F^���zH���z׏g�^X���myʑ���� ���!_�lZE�9��e�~�`�Ѐ�2]��&���ܽ��P9�9@}t�PA�α�e<xʽO̐	�zy[B��v'��ۆm��]���>�����<��i��tr�R��������lOv�beyq�<�_��|bp��|�r�V;@W	��Z �ć��C6q�v�����ݕ�U�l�@�B�%�p] ���P;��<��.�pgnu[��o5C=76����Sc��2\\j��ш%1M��9���b*P�.`n����&4� ��J��^|��0�G�4c�����0���1D��H#nvtJ:�~�H~�n��tw�����t�Y���R��֩��}5O)ε]��XB;�=)��S���Q�̊������F)���Ѽ��lz�g�D	>˙đn�-���,q�f���>>���n�WY]p[&'+�z���J��R>z�e���
���Z�?¶�A����^y���D��f�b�v�.|~�r�A̎�	����x>�*�r��#��{E�h�R�#�����S�ՇO����!H�t�ړ.��Rh����,���D��L�Uc�a7XE��ֆwMZ�^���h��]�)�U�`���n�����җ+7��L�w����� >��e<�9	��R%�[�&�&�D���ŀ�y��h�O�������NUl���Q�a�3�h��2T����+1����6b�;��e��}� � ����(����c�-��ÙS����H���ؘqt�T^�¯�rV$�
���dO,��j�mI��4߭!ӌ���g�Z���]iK�+����ڰ0 ��
��ֿ����(D�oN����fR'뛯�θr6�c�P��Zf;j<��e+ℊ�8��RH[4�;���џz"AR���W&����4+���N���t�4���,��}�!8�K�8�$����R��e7鰴$���-�QQ���yUg!�L^�Ҝ�wT������	��6�T�Ao���զ�W�
ҥ^�w�A�j��A�.^o�d���p*��
Z���f:ح1�"�US��;��k�6���wV��;z�v�7����?�!�s��x+7	�����G�)�(���xҪ*��]ɍw�ٕsE�'��,:Iv{��7T�ã��,�b@���
60P&Q#�4�K�]��!r� �f�Z��E[��W���0b���،h������[2d�rV��rX�;����A�����wKi~�B��y�l7���s����U���r{w�{�7�{�HJ�M�פ� =�3�xd^�b����#=�����AjZE�lb�<3�M�D>}Cg����|%[<&G���1>YL�bB�MC�f����2�h9�q�)�qɺ��+��SDB���ȸؤ����Cޘ�����!K�-g]7T�Lc�qm��6�w]ZC'-���u��Աp�B�G�1jo٤5��"e��E�H���ߧyxC}�R���c''��Rk�!8�HʬQY)(W�cg�Ry�^���A�F�9�d:/���ܡ��]��H"��h%��f����3$?H5�/�(�&B���@��pF��Ҏ�����^���G>�I|��d�i������p��6$t���7��j&��^n�#���hn�e�Ù�P�:޾V�ݢ���/A�O�b���QH>�L��NZw��O4Z��|\EŸut����>2},�]�eJ���	M��Rڲ_l�8 [� f�vN(h~c$�.�w+��7h�lP�t�ݴ�?�\�)9���LOaFUk�����&�mI`וd�ų��:܊�B�6���?$^�pu�н=�PZKU\����t�fp�:ųٖ���I�����������x��V�G��0��F�TU�������p�Y�Aʡ@1�'��r"��K�� ��-aA��u,��]:�)6�tJ���֔D�1K{���������܇_��b6b�L��Px��EmL�-�X���@F2�jEn���M.��B��d����r�{�O�m�	��KL�/0��;��.w!@l8jcd�O^�^�l�cg�P!������(��:m=��3��k��OM8��-^�����9"�݆�G	���(ݞS�ht�������Bu��q��sdu9_�˳�j8��|#�a�uC�ܙd�$�/����(`\L���.����ʆd�s�2cP^�0�2c�9:ԭ�<a3>h�IS�-�?@s-����]��w��̀��!�*t]S�?�-��N�z����ىKKZ��\����=��O#�%������wI����Ykһ&I��:�TX��f��/ ����jو�Bڷ�n9M�9d��Kv��]9���S�q&�d��4�;ݵN��rӮ�yf�Z���m��Q/��G�\��2��@�T�K+. �H��q�߃J���Kr�_�yQK���~�`��<�s�����<S+�>����������i��b,h@A��b��"����O����
T������Ր'r��l�v�KU��"���~��iU�,��tAf����9���>�Ԉ~�"�ʹk㻥���w�U#��hI�e�C��hfb(��y��%�!�c:¿&M��lN���ۮ?n
2�KV����o����v�}����4ǭFWe-R���ϕ��;h�s_� vp���)e���Zi:��O5n6,�=�*�[�(�Q"�/��	_��D錺� �3�J��D����aԬF��/�c�S���c
V.P����n� ��,Q�y�����R�Q���#��1ꚹ�F0o�(&'�(�	q�	^h��C����9�,����!��$���ew��ЊR�w)+AQ�|aK�0c��L3�M�s�R���lV�
�d���pg:5���md/#�|OG����#� `�Cc!�x��Xw\�qR�o�o7\�o5z?@ ��8�������Ѷi��r X\"����\�}!�|i^�'	�ã���P:�#9D�p��ʹ5�氜�bz0�C7v����Ȗ��\��4� ��Ò����dd���nVK F�,FG�,*ء|�!�� 8����:���"�����x��?���[5k_l3֮�6�Dƃef�}���l� �.))��9�_0͍�R��y�]߈=Rg��=�gN�����dt"-^�/9g�� Hc����0��?^k]�;���>텷�״1o��@���Wq|D�%�6�$e5:
��j(�J�	�P�֎��O����-���Q4��i���hn3�|��-��ԅ7�e���x��1��g%~;��?�_{YJ�^�p]>�X��nR�m��-k	S\�wU<��5f��CY$a��Y��EZ�w��ë�'6�9�DW[~+�E1O%��f5_� ¬g/p�[��]�r,P�e�7�Y��>��}0�%A�6���y��B�-c�a�e�]�|YS�N0DK��_v�<�g�-�NaB�mQC� h��e��u=p����2�z��F$|�hׄ��u�E�<Lu'H�k�y�o���L�|��g���d���߷h��.��O[V�n9��	,DkV@�"�m`�	�g$��<O�ɡ!z�z����Q��+WkN�� �_��an���:����lh/3Uk!��^(#7���8�t5K�8�1��-��*}؀L��o���*x=��J��0w��1<j��O�-�~�[��?Ror��f��������&��K�C��Jf
�\��Z
���0�vϿ)�nˍ��x
��x���p(�"����x�+�`5K�ct�fX�ᄇ��V#�������ђ�tuWBU<��߷�8�|�ܡ�����^+��^�O�'�:JT�' 6LV�I�!�;�A70���`�-��_:e�{0�:������.���"H�:�!���+��7=��"� �Z!xs�D�˪,u	�<�4��?�w�QP�T.~X�?�Q��ZÕ��=@c��Y=G��X5�3�"	�EE�H���%��/���yr!��x-���գ9g7)Y�Uޮ���.���Ց�h˳����+�C��p2�*[[��@8�>�GD?+��˭�v���T?#���|"����5���f<I�@�>3؍��	<�4ձڹsQ�n��F.j4��$ ��~���=xu���Bx8/A\<���}���J����Y�J�@����+.�J���\*�I��������nt�#�L�;B�4�N��r�c�O��'�9 ե�.�ٖ 0���b!%i`��t�]�ўLa���M9�l���59 ,\&����V_]�0+S9t� �$ΡyS�˅n�`t�\�mE�� ��d��8���f�B�����tYK�4F-��*�n�PT�}<!��-��]�%t�3F��ŧe��p��r�ҥܗv�6o��f�ƨ6���z� p��idfC�xh<FR;A�{�{o?���������RqP	5�e�0��8#wx���1���o��g�w��}Tj��h`m.ϐMM:M�����
*D��
��0�����F���e1�HYP�w��JW���$Z��W&�M��:����0 f+�w���z�_S�n�1��R��-��Z�o��m>9�lI悥��z�M=�0�����R����A.>c�}W������M@�>㒕(��2�'@e�j<8x�w���.�K<ߟ�(��5�a�~애�k�XpwwʦzS���xL����l��e͂W÷9U��f$�f\�=�S�pâj��]$����"B��-E����'.�X�T���d�#ջ���H	Sub�Ѭ��������߷�X4�+B>hH�g���\�ݖ��@|�Ltd�?�m�\ݾ��XEg��6P{9�Eϧ�C�jYZ .�ڬ����'�>aclT�4���1Ϥ�[ź��z�C_���Oa�i�4��=8�^�6�H����7�ު���Ie�Ϳ=�E�I�Btyyj��x�@5h+O�~t���YM�,o��pc���e����������r�(�Je��{Y� �/�ė|��o���E�vT��BA�Ő�4��8ׂ,��h'��7a�O(�p��[W��S4�� �qEH����&kռ̱a\�):$[�S��eM��܀Ӂ�X��>h@�L���A�GLk[z��j�oH�?�{ϯ���m!��X�a������c�Y0̮m����²���DD5�Ĭ�6o�`!���]#��DH2�\z������&�$��rܳ't6�Υ���Q�
dK��ߤ��,q`���[���x�S����"@5��ۤy�_I�F�a���	-Q.� � ��8�� �yr���EU���s@R-�TZ�Et�ԇ�v��~,�h����^�%<�q�1C�C�C�� uG��᠃&�C/�l�i�+�M����k���
��;���P�o�1����v��-P�5����bx��`9Z�sy}�v� ��V59�8%�����i�d(���ޢy�>�wt�q	�	�=I�uV؈��C4Sq��y;�,3�R �Sw�O>���P��Ef2��i5�Mӈ�t0\�
	���=�_B5c\G��j��=Ơ^e&��>��<�Pى��eXfN���w�4έ��)`!7��=��y�c��=��v������{1���?���Q�6�72����1���ۚ%7�pjg,=0�] (��{a��ָ�x�$�i+�=�mק@Ģ��k���ٛ���H�h�ģ���{��,����Wk�ߛ�mhę�6�p�zL��˝w����,��F�ҽA��j7�u7yn��`��9��cL?�Ml���1�}bp�d���P�G�/�qРu���-|B���(����b���}�=��ʔ;̟���9 �j��c��1�y�.תcQ�.��*f�t�2��$.�F�rP�3�<UNi�S���M��b���,��Z�݂�dm̤��L"enZz��;�����ͭ�mF�1��]����	 ���{J3��~}f�	���q_e���F�aҮ�B���	_�Ǟ\%���ZK!E����
��8��|k;~�BX��L��y&��PZp%���l4h���21�a]fݗx
��IYu)/��p��r	h�jT;���b��Ȗ��<?L��x|�=I~8%ĕ ����U�a�`��O� "ŉI�14\(��	��~�i퟉j���C~��{�m~�T�3�P�P���7s�?2�����bY6�ƍdL�F�A ���i��;P���+\(;WS��'bB���[�j��K���_��J��8�hdmq��qB�Y��<uŻq�n�
�u��,�	�ѱq�&X>Pi􊧦�%�F�cA�6Q7�ړ7y�0]��|��e�@\1-H�?/���Kz��@�jo�9���V�h�<�HL���a����u�yO>�o>��R[Z������C��S��h��r��(���=2�9	���7��8�EWǊ�ZU�j�A���/7���t��F�|?�K1�h�v'��v������e�����Fv��<\oQ��v�eɈ�`U2'�?���zQhzѱ��Ϲ�'��ͺ�6ŕ�k%�;��/�,,�n���S�J�3����C�����A8dG8��i��|В�O�<{���:��̶�E�G�=|�mA�Ȝ{ky��s35,%2��we�$�
g�����LT8I*P+�?�y�"X[��1W�em�D�qP�`bŞ)X=�[�5��&��3у�(�x+�xՕ�^��$ǳy�@�ߓy8zd�.����h�p�Lh.��C?Cj��2�b���- ׭Q�,�.��df��P�J%:�%���R����Ϲ�7��Ogx�	�-��"��Z4G��"���\
Ʌ�E�Bӈ�6� ��3P?9D�G���X˶�[P�f���W�����N��
�`�.�ָp���Je[�g����Wa��ӥ�²y�5<��	�����-��D���$�ٔu��uu��f���kpQ�5"K�}z������PO���E�	הx^�q���S����gB)Y#5>�B]�]	����u���m�r��z��Ò2Ɯ�r�J�J{#v�1�.�v��>�gc/��=��̂#�(Q%ɲ����W��w%=}Cp'���4nJ8eeG��I
��ަ�6���1V������]�oZ�
�ߣ?4�|�
T'Yȩzg^�Y�3��a�[��N�0уO�L�	��~G����
���S�Eٲ��y��,@�MA�
���Op���^8o(��:���Ԁ�5K��0��UbK�Y�;7����u��m���t��J��O����rKNZJ߫�@��;Ls��sʪ�����b ��@P�Bˆn�3��i�6(��'[@���XT���I�[s��xEH�Ώ�	=Lz/���1>0� ���t�tv��K��{�׈�%r���B����pJ3+�F�#%r�)���7�̀@R%��`�[q����v��<@g ���\H���_C��@�>^1��E��G��(�z�'?��Dxu����� no�����=R�ok�c�$U�&=����df�U��<�M&P`x �̈�����y*�m#�fN��f�2��m�����.��`֠xC$l���{gF���T7�>"���]��0'� �QT�uF��:,��EC��n�@�-�F*.���vE����㈥��m�߳�쐇T1��Ki�7�ζ����|���]�փ\J��B0(�7�D�
a�#�f���n��WE�|��X�v�?���-�A��4�8�/��eBd����9A0�E��$�篋�È�sb���@��b�׷Is$�#2�Ǟ�l߀ )�k�u�ft��
��"��[�rT8u���J�3��A���I{r�Wi>��J7����|��T8�F1g�uy`�h�_�"R��x<]�q3�w���6+���v]�Pʃ_S���-S6�,�v�|�%����>��TS��ͯ�m���i�ײַ�\���0�)[t�W��Sc�#P}P8RU�ћ�b�}=k��a����j埅�Eoh5��h�íg+|��<>���Hcc��FVV � ��M\ECz�U��I%d�:��o���=`Ic��VY��F�WN�?�
Նr��c���k��|�\#�j�;Bg���7��6{9B��\�EB��>L��"��l�m��%1�"`�1>�7��}R͌)���-�P�-�B���	�ϪA�f~�7��xF�1i*�;��OɿM薘�?�8(2�4��=j:G�OZ���bmZW�"ZY�T�����1⦐B_�qz³�1�e�P�(���wF%c��/�i^E��� 4�Є�&� E �|X��wNRNE�ݲ�t"����!4gV|d�������yO��k�m��Hiۇ��fa���ϋj�6�)"�Q#��
Ҭ�ro.�r������0�s�DNAl���a3��:�����K6#����Gǹ6��3��9	#���L��d�~�,��T/���_��.��#M�w�5��6��><�K���ջ9�N0E�Ks��	b���y�����s�D�
Ag�g@�N^&�(���`Xt�w�7�d�r����wx�6(�}cVN?�U��ʩ��ך��=��M�)��5�� @�]���{l���Y���
�o b�Ӓ��?dl��t>s@��O�9��t��e���h�j#C��y�^;��;x�w�J^?{��`@���x����s9��X:��3P��Iˤ�S�'�/q��>���� ���<��Fm~�Tw_�vĵ�*�H����{X�= $��^4@�q�aDC��~gm��	����[�.3R֮�R�k�|��?�צzc�]p�Y�q,��������#���Mk#JA�P
gfO�6�-���O���2���Q�@�||p-���'���M!p4"d�~��e1��{����.�����k�?&���dHf�E<_�����e�-���?(�����d���RJ�b\mq���@y��+��
_�j�H�!��D�OMi�d�j�i�z�G�̵��0}P(2�[ �;j��z޻7�����x'%�ԫ� J�co�nf�zD��� �ͪ���֘@E7�\��ۑ�m�����1��H�'52EޒL��5��6缪�<�:*s?@�h���t��������ugz{�D�<�P���)}߆ ���km$��B��nH���fr�`�,O*��'(#��
��Z�hQ(b��y�q�䒖,���UԾN����=����rL��	Cx;�+��.�ƙ�B��&�\�.yƩ�%)�����ir/�.^�w�i:�"�K,R	�(Q��cO��������fm �5�U�"K=W���&C� ���ݰ� �s/��"Ufw|�%�;�>+Da��Э�x�=�<�Vj�����$�Ό��d�3����H��2ܡ�a64�'�JR.x�q�җ2d�J]�ړ�j�$�s]�J��a�f2� �)���`��A�O�P����80�K�O�}�b��#R��u���9<��%<��>�_s�w�(o|/��A(��ޯ0�Dw��_��v��o���)����#�nHܧ;6
���|��}>F�M\�!���}ܲ��Y޷+�T�k�N'=�����֮�W���D����ً߯���4�����v���'����cl)�z4٩�r�H��
<q�g���N��H����PU���zݓ�3�k<K�Xc`��c-GާV�W���o��mL_3�ε���"�u�h�!e��c��ւ��:h�%}�����1��s��B�_r�'P�M��B�h� f���C��_�6�@#�ZS���`>��y�W�\e�q���y&��T��s ����[��B) ��8�֭\���Y5�Dd�Y�F�B���D�
�D�>�SXm*�����F�U���/ � &u��l�!�J`3�C�����y��R_�<�*���o?���Γ@s޷��NO�曤b��'H��(�6N���
$6�6 ��VM֫s؄1x�a��}�z�]��:kEu��ky�%�U������,��2�P��w\^�w��w�/�.Z��^�����S	����92J���0��{��|��Ċp��)�a�J�@&��<�"���O|�0��?D�ҋ���ƹ#�w�+UL�����B�k��H肺��Wu�(j���6����K���̫Z9���d�7{��u�	x,H��l�z7Q���U!YԎ��J���j�+�iav�b�꿣�G���uo@X7���"
�яq��Vni萓�|����AS�e	/[L��ь��b��)iV��݇����3��S�OcW�Y�����p�*�{� [	a�k;n�$?�n>�1b?��!j@�enb���&�<��H,�G�Z�)�����	P�H�a@�Ou{8X�E�ď"�lۃ�|���Hmm��ω�U�?0o#}u�<�I�xK8hh��1`e��d1^>�Ԯ���=[L5%Oۙ<{"Ҁe���?�i١e\��^򱉰"���`h��8k�����G	���wD˨�=�hH肕�_�Zݙ���Ӏ̍�?7+Z�_�:�c��[�����r����4ZK�Ϭ�V�Mk�'��ڏ�`(̅
6-:�}������l�������GT��A�E�%O��8=�l?�Ԁ���:��'fߩP�RX n>��+����U{>�T[vF�71�Z��v����`�-��|q&��K}�ΡW�i%��;}S��V\�i)���_�D0U�� ��XKD	�߂���	S:�Z�{p9��N�)�L0P2����{Z�w���4�"/'��0��VT�Va���,:p�t�C\����;����#��jg;Ņ2 lv?���q�'#r�
B����T汽y�H>7xomt+@�".#һ����jdɍyy�s-�E����0����3Vb�	Ǡ`�L�ڷ�)v3M�i?�)�����Ezi3H�;1�h�ٳ0ƼB�EZ�##9��oThhU�'/}�dgu}��cw�
x�y�c]Z�u�2@�~�5�<��$�X�ղV�wk�:<g��� ��lMH��J�zL�D���8H��ǻ>�͸Bj�}�=�� ̕ZM,~E��n+����^�K�x)|�����g��~o[�V��HqA
��B¼��].ZrS�%eʔ�8�0u�0�>�"^Sĺ�UT �"�Yh�j���b&��"���n��[c.�u�8�� ����N>�=��>쑼b1�2Ƞb d��u޽R6+Ў;g2䱠��1fԬ�(U}�
��<���8���c���+����Ɍ|s+�^��bN�+gB�� ڮ�nx����9�a�G�*��/��W��V�j��6�w�f�PrJ��K1E+3h����}���� ��<:�T�t>q�hp�8�����^��!�4�q2��+�9��� Z������$���W�X���(�+��Eqtt�S����>������w#D��>M�Cy��A<�����6���T>����"Xl6�	�ۧl�`��ϵ7����|'i�g������͆��N�I*�ߌ�?�FS��kd��0��gJ��1O"7�d�f�Ƌ�`1M�r�q�@)�E��#;)㲯��3i������?t�R���
�2�_5���
%J�A�i���<Iz��f�b+��&v��b�l�]wN�0���P9䲣N�e�dFPJ3�Cܕ1�(��f�d��9��V��q�NF6�4��*w��O���~	���!\�"�M7��}��w�-��dҿfi/�Ϧ0BNdp$�.�/��Ս=�#�x���=��C�+H�_:�]���۳y�T�ت"�J�$��t�$a�h�~j���k�������Ώ_V/��9�S���z�s�d��w-z]�8����ʑ��謎|<�T1��@fEs��ul7om1{��.�98�Ƃ�N@�7�$7is���2PT��j�+v���\��ݛ�D<�T�,���R\�q���G���������ְ5�a�D�м�f~,&e�R��	i'gx�b�A��vT��C��¡�^Qb���RZ�j���7c
ۏlA���6Yɏ%c)	iz�A�������B�j��<�H;J�-�B�4���*�!������Vo4x���8����o�y���0L8PZ\x�:}CG?iG�R� O��<�ih�V��	�]뮾�U���G^c��jr���?V�@����*Xx�剷D�%J�xn.}��_��e�o ��������S'D�<��-$���7����te[B�z�@�ʉ!��	�C�i3�q֏��-�<��ʑ,|Oy*�Z�q��G�����@�����}L�X5Sqo\�/�x��LS���qS朤{g�s��:����/�ڏn+F���E�b��F��� �X�.�;��Q��9"��I�}*~�Î�����p�����g�f���qb5|�?z7e|iҏA�3P�������m�߮z����@�C`�sB�7?��Q$���<���:Xi�;�^�t���d;�>�e�H��w�0`�:�`EP�ƨ²EuȂ��8���x�h"_����@#Y��tŽx)a��ο��׺Яy?Um����2���P;���<����m �N'�܋<q�AE��t�D�cUӊ�;xK�i�q_4,��N�2X	��*Έ4��k%g)N���c>�{����1��R6�'����!൦�����L���¨C2BNzb� ��~c��>w�����kB�[��@|�r8�B'%�P�a��?�������NZ$H��R�������NiQ����+cb�>m,M���aA&��+h�$������\;	���\1GevUf�#�%l�!7�Ae(޲���b;S�`I���*w�,�9��KI� �0��]4(݋����%�G�,��V�3���DxUVJ����9j���wxE��h9۵@խ� D���U���b����tچ�^�Em?ʟ\2��J�yG�]�À��JDXv0 6J��h�l-���n1�$sv���k��_��Me��nB}|>����#��b$K��7A���v߻���Ķ1���g�~�Fd4l��|���$N�:ߦ�{M��3{ú�?�b����Z�#2��
��⨊jqV�m�t<���Kq/���(9�~e:�vtہ�h���dC!������ۢ3w��?��r0�����O��k)���ER�o����R�'Elxp��Ƃ�.V.�eQʒsX�<\�EB�څ;=؇EYSǢ_:�S0�J<jsw�xj6����>Z�tJ���pBg�atG��r�L[Zw(�JW��?{�P�{�'�i 55�|�e n3�í�a������WE*-@�E���u��gd��g�B�^}��'�'�q�U������'<"�)Oӈn��)�{���
��x�����7"�雽p0���ߝ�����˅���;���{�� �b�����m�GZ՗���q�q�. ���Q�����J'|�dÐ'Ƥ���(	�m�՛$ꃿ�!Vjp����h�a��w^���)�D1��
��P/ο�h�Ȉ�4�PJ,nG�5Y,�֏/z��[�������5�NiW�����S���S�2s�7d+���9�'��`��OP�������WN_��Q��� ��\�{ �rF��)o�ttF�WV���+��G�z>-�u��y���OTXP��}�OE��O/BA�>��n�~jɴ9ͱ�И̼f�6|)ǈ-������zSc�� ��{�h�#�K�o����u�q�(#jàHp/[��0!Q�E�;�@���M9�>>)��.zٌ�wm�T��h'��A���=GGX�G�^G��%z{p�DxN�tY�����q_.x��췽P��9����C�P�yl�k�U�a{�Rb�����$��M3.�T�M����}K�a�z�f��g�K�9���}��f�P��p�}gW�s�8!f�I�M�R8E�C�2V��A9�,nC����]F|ᥚGێU�׳SEK���T�>i����l+��7���$�_1����H/�K�/�d�ym���w��������pT�ܚ6XL���)�L�L<n�@n��%���	�;%51��&jYe�Y�0�V12D�lw�l��@Y����`jY6|-��^>�'��^�r����3Js 7c��W����t�X�ҡH����p�;8��z����b�Y�`���!��Wg�p P%���q�~_� \���C���c��~��+��@�y؟ j�H=�=0oU���یO�S�����՞��ɩ">�yo�������F�Dp��� �3J||��ZB/�6N��]�գ�M�}!*����߷�Z]�0\͘�y��4L����`S��I���±
!�:)�@����d��J�6Y��W�E*��� �L��_���/�w��9K-uU�<�����':+�6�	x"*9��q]	��)�ͺ��������P@�ξ����G��*�sk��k�aL�q?怎�l;b�4��,���!�0=1>Wb�tw�[�p2:ń�=b-w\��46Z��B̃�~	�$����h�(�Z�b��y>�tk���k��>���s��C	p|n��:?w^���^U/���fG��\])�*�1���)���N��V�5�4�8�)���r�������ޥ��*�P��*����q�ǵ�N`�0��ʲv��d�J�8��V�S#I��]!F�r낺c�1>1j�Ĥ)!j�K���S�[n3dphM�+�!Q>��<�Qn׉�Ҭ��D��ߎY��	j����}�	(���8ǘ�ҩ��qQ�@H��fh�#���5�
k�\o_'P��4��j0�l�#L�M��QEut�3R��~L9�Dc���3 Vv��e�k��˫+�����d��Aa��M����l7��V6�iIz��j"��)���|�u8���-??:HaJ �����6t9�N�wݩ��O $���(5�D�%��4��e&���6jQ��K�����_�cZ`�/�[ͬrR(W�t�:Y���G����*��(ƶJq��%T �M�+�� _N�wA�S-��	�&�t�b����i�UTV��%���K�b�M��}�ӎ&��k�hu��M����5�V,��v$��K�c�D���Z�S*���M5����k�������6���k���^$ڙq*I}��a�}�_�Z(7�w���H�*z:�k
��IƲ�w>C𢽵����C��K]�(��Y,��v>�t���j~8VL�� p��QYagj���53�����kTơw�#����22T��8'vQ��><��W1W��`e��wr�M5bA�V�o[��A=��uu�lEtZt�4xR|�/�� ���s��KӮ~�L�)�2�c�S��+elu��e�Ҝ�1����!9,1Т�f�Ϭ��lS�;4��i?<�8x[�LSP�F/.���}[�!5�uK䷮�+���9�ڌ9˼h�H~3���_�u �(�'pF��39#��6�8����l�
,a�y�ﳾ�Yr��4y��`p;���>�|�|�+�:�/U��5-�X;A-,�q��l��5�i�_��E��, 7H��I�[�����fE��v�m�D���adϲΥr�Us��&/�C����.��]�wn�T>�6L�={uQA��x*|�l��rϒ���&�
��_@��`�,���l&�)�^3��mZ+�d��`�$��ɉ�X�;�.�5Tk�9����@�X�
؃�j�wKi��`n3��p~#U���g?V~�!�n�x(�Ʋ��|��V���S�	�c[�F�)��~�L�|Y	�)	j�2<�b7��CDf�/��B��s�l�U+L�'�J����G��l���a��n��,TV��m�fl�5�yD}�,:��Dc�
�q..�"��E#�����:]�:V��/F�FT[̼�bUt�]��>�TH��&��~3�[0d��҇��Q�q��޽��\tm�/ҊTեx�i߽��JM% *L���(���?J{���޴�-��sr��+�p8��z�TMz7��ш���(�m�OpHE���v	�v�7,�R�9�>$�U 0s�|���ŵg�_�����h[����/Gx �!R�G]��K^`�� m�/N�k��>����)��~?Ǟ:P�T�>���M�4@���;�K{�R-��d�Ҡځz�L����\m'F5�����{�$=sĻ���i0X�%%|��F[?V&��M<_���l0���� �&�+V�+7���]��b��c���r75
ߣn����LchEG��]�ƀ���_��"�0S���?�"4�y����I��,wQs$����ܹ.���
���ȱ`�����|�w4UJ�|?&y>X������\&��nc2�R y!Qޑ{fF�l���}�Ʈ�&�M��$����9�J`�� :R��h�|?�,D����M�u�&b�Skm4�N��[���Y�$�����x=������V͝ZO��?�=��&j����JΡ��1�ɞ�ݘ�Ʀ`�ʡ+��:�%F��4�i����uaKSK.;V˒��3Pbm��R�A�\�*B�b��gK���.���ɷ�	m��o{�۩��ԡ����
�X��@G�����"�<����`G\Z��+�;,�eȴ���p ����G���E��<�&�G��z�aN���S�p(f7�R���ƾ���0!�,�Ђ��!������ȟ���p~�l��8e�Ҙ�y'��܈�8L��U�Lx@�/�1Vl6@�͏�pu��f�:�p�F�m� z�� bb�0�yew��c�`s�p�*ƛ����.��V�f�>��aE����!T���"�e�1�`4O.���/�z�����{`���u��e�n%���f�>!��p+-�+-7.����j���#��U�����ȑ|����xM5���	S�%��������?�]R~��K�f"܇h����ý����jq���x�2����6�����_��6��A�= "��9�p�T'�� ����#��QjW<��K)$;�Y#�	}�{{z�=GKO�JDG��'���c��]G�[���M��S_k>�ؤ^,b�ܽ��3(� >]�EZ��	����]S�"��(��b�O�V`�G7D	�Y��(����)��*b��.��4!�Fsݩw�Zj�R	Y�%����:�D�c�������RƜ�ʢ�~*��q���G���Ҽ���%�E����8bJ���PlΧ�ȠE`u��ݠ-$ϛӫZ��]]v�~�2���关E��چ���׭�.�s��A�!��h�ݔ�p�y�K���P8w�΁����q"y$�������s���o�hbDl[fמ������c�-!Z)�
Q:�
�� �%���8�W����4�xD�b���`�c�@^��_�l#<� ~<P���2�Z��g�� �*R���0K]ؖ��VY`�<ߏw(�j���H<>�tk)��q�������eJ7��#e������W����Wt<�B���Q��Ӡ���#M����:02����VC�f}z��aQU,��0l5$"�;;��"Z�P���W�oN�$�x�Ֆ�>
~�;N��b�'��6�a�Ƥ,uPpImGCl��;�)o\�,�����Ye����d�C��TY���%S�go@<�։�7�����#܇Y������+�W�mU�;�X��:���Ŋ�D����������X�{$=8W7�:����-����5b��ۜw���/"����rV��YQ�lyPV�yw�hC��p�֓�Rbɉ�4 �&{�1����|� ��	��,r���<C�o�*���(�0��@��6�o�-�.��զ��sl��^{�?�޺����8~h@)�UO87�C�	=�Q2�YKH����.8��&�����j�
!4������`���T�g�BqQ==E$�՜f�d�~�w�����\�ؾ�Kt�v~Oe̓��~pM��Cϲ�^{ߒa�m�"H��1���\FeL��	Ѯ�y/Z�BX;!jD�!����o|E�Hv�/B��N���90�.�V�=�i�F	�Ѹd��;�q�Q��קb'�����DM�!��n9��(�p�CO''�eI��_B�ǉh*YX�1���_S��Wز�r�����#=%K�_}�e+j�B� V��O��$��Dhp��'3}jȤ���)6���e:��W)j�B�©���p��=��W� �{�'&@,�&�f������1�zL�6�aZ_ 7j����Ӗ���2�$�x">&�0�Taˀ�1���X)�ńWɣ�+~��Wck��Z�U��_�h�"Z�D�^���ǐ(�������Ұ��l��$4[���]I��FL#��r�����ΙǗ����12���.���4 �\�	������=M8��M��J`HeX�-�_]�"�a�����&�1�/�F�,p^@�Naֺ���@��0��QVu<��F�� �
���`�rX�?�R�ħ����C��{ay���$���OvU�=�沠,��`.�Z"��,�\5RU�$���9Hje���f,~�Z^T���4.t����ʭ�ap�L���L7�w�d	Q�+�m��-uVh������ q��V׾w��Z�"�C~��]�) ��j��<�����a*����g�Kj��	Ȗ�����s	|��x��~aEH��F��y'��2M�K'�� �[�m��Ъ1�Okv�|e�����/�0�QeDFQ�1$�G�,"��Ψ�eQ`�E6<x}"z�.���p��KR����%�qs7g�d���L������!xP�}+�+4���-�iޟI��(ŉ-nܼ/��j�-%��O/�7��iJ����ը��N�x��U7�4��4���p�jMy��K�C��7�a��}JH�3��Bi#o��t6�/���vF��P��&���}�͚�i�G�Sj�s'��`=��|�?������� �Wp�T����1X�bqC�eX�d�E����iݿW��,:��`���zcYLk���
32XL5��F�& ��0	Q�Y��\�}�gb�+l��K�8�8�B�"d�}���c�!��#���I*+[Ti&�CW;IQ��f#��͜�[͛���VŢد�|���@�����8����u�feT�E�$��㜲2�>>�j�0�6������f2y���>�HOٺ:9���OK�} �s�q�'�p�gU�0X�V��';���%n,˜�j+d�րB�ii����pjPjT�J�$�c@=��)f,e����W�,�|�E���M�׃I6��i���|��1(���2��!�!����w��H�k).'}�uV�j�;�&�X��3t��d����\�^��O�h��S��/0��R�:/��F?u���X�a����o[�rI9�ق��A��{!Aտǳ�b�bv����F�VU$���m�Ą?j�#���ވ�4n�<3�����`��8�>�(�d�i�tMN�B�{sH�\�z;!5���>�9��j��d6�w
7�'�p��w�mӆɜ{|���
Ri�<��/\u��+�?���}�5x��u^%�� ���=[�u���D*���|�5����Ȼ�"�1��+z�H��^�����tϐޕ�7N0)�P�3��Hz��Ά�R�7v3'_��.߮ۥg�"�p�I>��Z���b��
O ���r OW/�V�۾�ת��x@�I$���`s�P�oO	�b=I�?��~�~�� ��I�~�Qi{j8��]C.8�L� >J��2��kD��Zߞ>�ߜ�J5n�\��FL+��Yc[�ί5�C��D������"�� S!rbśU���~z*�:����l48����aF�]��%�d���rN�*�6�y��a��O��5R��0r��EA���E��0(��H�A�Z�T�xXpD�2�5�J�0'�˯� �5j����oCc�tϜc�|%�^��RլֹX^͙u同vH���A�Lm�?�4iR5��ԫ|��ϴ�w:x�'�Q}ç�%�؃����3AI�
ny�5}BmW��=�쉈�>�C��%�ZFf�qcj�ǵ�u$[2�����3�����v�ϸ.R�s��ѐ�����U&����|4������2z����׼��	���>�Ӿ�����)Q����k������:"�t=��lU�f��$� ���h��Mz�����V�l�7��+��:Z���#�kvGE�?�#`�j�N�8��1T	��Ґ�`�a5����v��z�hZd�=�Y��Z� Q��W۶̙�uw��{�T�,�ܭ|/]$��[f�#
_��Q����g���p�l�}����n!\���I����UyU#�86��}��6�(�i�e�@:���<	�d��ŝG�f0P=�!�'�0b�gm��v��R8�˼g���5ڊ���vb"�:9UQx�Q�L�/.% �������S�d�����7�X�������w?�R�E���M??��9,y�T��V�Gn���؊��w����|��I�B~���@Ժ�~�EB.�kiH;Xni�9Sn3|w���\��_֌��8q�\g��'B2����=�ۊ��%9$��,�@��Kߘ���'A?C��9��;V��uD�PN��%�M�G/�H����UE��zؕ)o��&�}�:�[c5ڲ�"ip�1O-��q���z�R�R>Ͱe����J2�/kDM���[�6���7=UD)��<�~��hf=��,�L��;���Ӝ�:�����<�!y%�8���5�����q���נ�/�Q������?�]�\..�ڰ|0�"��:��m�ɟ�E�k��Z��"b��HɄ�/�ٝ	5����3w�n�4<�oR2� =���7���d��~�}>���*\皱H��!�g����%�����~��O���EU�{U��肪. ���i��"�*fy��1���/o$߹�@�`���i
;$�w�=�_�1��n);�bü�qN̢_+څ��c�D.=�!}7�-�
(6b� ��o�Ȋ��2qSH�����~Y�<y*�=�eڪq�D��{��m+�$�xFS��O`���U�p\���?�Ĥ���T��
!5�����Z�l�m;E>��u�@�*7'L }�|�d��ڣh��A�D��(�%Ž�D�7v�5�Aj��\2��^�┸I��B��5�����FM�����s�6=m�|������^��oQ'ڬ��J�
��s�;�kor��Is�m�2�͖�'�͚�ܯ����tq���wH�q����lXڕ��O��,�z|��7� 8B�U�Yt�ò3�'@�$ۜX9A[�^��93[s���|����3��{�'���{TR�^Q��(_5Q4��Z�֡��=��a�,Y�{�8K�en���%Y���8&΍��LM~��Pn��F�YA��K뻐<��f����;qp]%��׶K�[��3�2�9��8m�vqr�y>Q�)�^Q�}� D��N�O+PV�!6q�?��ķ7syIap�AsF���ͪ2���a��ߙ��n���Ť��F�q�	8��q]�h�O�3�N9^ϯCz�|����&{�j#T���Ghuq�Iv�g�/r�b���Z.Ȳ�1�ݹ����Z�o�{B�*�I�"f�s\"OK
�h�7ue�b��k�옉�Yt����?v�� �T��+9������6��������U*�y��[��n�,3Z�Y:��p���x̕�ݬ�Z�e"�.��-��Y9��k*�ɖ�n���'p_*�9���U���mq�>�Pf����u���6��<��;��dp9?�3�����mF�-�Nc���^�@�2�[�J犵��jJ��DkOMU�&���p�+����N���[��y�aX��;�r
"B-�����HC�?��;�??ߋ�t)T��ۤn�P�C=�u�]^��|���_���E$��6��ֲ&�l�����q�����t1��5PPQ2ͮ,��re���N4n���U$���P7���m�#�h��,.i~$�C9���]������"GwXF�xZe(�Y5���f�����{Ak G3��o���2"��~s;[�B�L���No@����s#�����go��/:�m5�ǅ�
|���%��:g�q3��	�H��9����r��"���j� ;�Y�{���(� �v{4b.�PwK�w�\{w�ٕz�␜�!�Z���6��y�R��E��\���JaEc$�7Y���p�\U��!Q#��/�Bqid��S�y�9�4�K�LV��h�Ǣ�O�.h�\��K���"Nk�d�����NJ����O���zc?�(/�*�R:��И����}zmj��p�՚� sݰ���|?�
ώ�S�A �<wEX���E��s����Qº���F�/�o���OP��Ѯf���}!ApT��iIp�x�pƞ��������OX�z�Z������!���v,].��D]|W���j��PֿI�%*ZY;#�la�̎�@����ȕP���-���Ic�Y{��M99���.�o�l��Ċ�[��>�=�+m�4�iM��C�=ik61\o�CX��>;P/�x�z p��ݫ���3��C�F?���Ƙ���T���ٿ+Ө�8����~3���	���Wb� ˅I@w�����Y�ѿ�rc�iɢkҙd]Ӷ����cy��q�p�g�dR^���F��K�uR'_
f.d�Y��&�3�⪐S�ut��+.*�V�� ���>�����a���%�o(9j�g��o ���!�)OҺ��c��h�>�s���(�v4
>L�3�f6eܥӢ�9 ��4&���X�A�eȕ󒪚���Tn�>����ϭ�����Ґ(9��П�Y�� x3Z�����K�	�0�b�e�I�0�l��k�p�t=��r�\
[de��`�1.X�T_6^ZI8~�x��jJ���Q�k E�ßck��=v�����V����S*Ӧ�#�	0��~���io�:��3�����0����&��性:��5�(?�@�s8E���Y5D1��9���ټ�2�+�z&���$�4Vf��53�ڻO'n��Ǒǔ>��_i""���DV<�ɂ��V7a�lUz�!��荷|Y��t��(jQ�´��k]�+��>N�B�V��<L���x�bx	'Kw�� �G� Ze�/#Vh�/:�1.��70��.�����(/^�[�=�i5I�\���G�Aͳ5��U�D�~ ��rU@޼���V��4?K��AՋ�~��U��[觵���t[þ��?�A�m���Ug��]��G�w�9������yv�_X�X�z�r�-� �����P3Ѫ�a�p>(�u��,Ũ��-���>�����f�bkb���p��M?ޥ!�	#�F�O��ݦ �����\�m�����9�q�m����;N,:GQ;c��rz�ƧO�Ц����1y��L��i$�_b�;��4N�j�pp��̥��s�uɦ����I�jC���yx��W_V-�p;��/ϵ~�u�3��~����Aɴ�{���[�b��>�0�ѲS�#Y��c�����`���&�[�G2�$tj��_G[@�	ΜQ�V��/�4@W�Q1��Â�-�Et�n�gq��8�{�:iGy�7��J!~Z�p���2܈�l��Oz��Ŵ b-�sڀJ�a��N�
2��܏y�N���<���eԴid�[{Y�ҕN{��mG^�?{���w�W�I��!��O���pp��X�>A+�҉H3�hؿ��X���օ,���+5�\S��i�ٯ@��V��f�"�=x��������+#�T��"-C��_�S`~6ذl%@���D�x-8&ޗh�;rD:|��s��U����:�����s���i(���*��ݘ�DU�cfq7��"7��'\�<�PF`B�
�gd�l�����A�m�v�4y��pt���7�e:��RLh�4O��`�]��j
��Og�͖�[��nEi�x�`C���x�L֑2>��8���J�"��l�A;I�[�9�L~{��Z(��c�D�7NʫM�?
��z��X�I�Fe	(�$Q���2xVb��]U�8 ~Ӧ�N\��(QO�8�������
�8"�,(���I)�F>K1��^�B�h�^U��
x���a_����	ω�ؿ�a�ʳ)TS,?R.�a�	��2t����c�F07�M����#-�"��;���8Ԓ[��4n��̷�R�i.�8�tTg+��$0C�l�D]�.xM*d{�O!á)(�O� P��� �;�I��|?�`mie��]W������U�_��c�.���{­9žuJ/���I)j�G��$*1*5ju��VJ��K~_�Kn�{���h\�J�k�����̕1T�b�5�b�M����j�F&?Ō�Ug0���J$x���3�y���^�R�~Ѵ�Y)�Z��l�;�1'�Đ��v��I`��E'�2���k����p��ۻ�Ӗyiڬ	a�]�귪�Ƅ1g�}O�W��^�o� 1)ȇf���T�3�5�M�{�n�քb����5��+�~�E5��L������,�V�r�~�L#n�͉3��%?�����W�AI�sB�v�����j> [`cB0�0���x2l��/���݉�QC>��	ӳF���U���Nޞ���Bj�_�>��}�
"Үg�/⢳�fD�)��*ߓd|cJ�Jp΁��P�j1#�O�UZ��U{õ`]�Ëul� ѧ$9��Dw��t�W�ߖ���B��~)��y�[G�(�KI܌��k���沐���2�����۞Sb�w:&�CّR��_��g����FjOcsf�����6����_���g����P!*`�D�E�k!D�7㕏���Ř�rP���]scW�b�k�=)il��U��K/#��ؖ��7����]+�!�V�D�.� ��ش4��P��Q�S�f��=�#�E� �|Ķ_K0#�>>'��B�y�'���+���He�<�$�X�Nk,㪜TB(�-���sr�B]÷q_�w�}�T����
�s gn91��K�Qұ� T�M]�*�6v<�)�Oe�0�
�|���Cu�{��lVK� �z<=X��C{#��'�Anad�1�7&C���*����e�"`C��2��'�ރ=��yC����\��GW:/��o1X=��'�q���Q�-��:큲�c^��'��Lh��8x�I}�7{��Qh{i�و��m}>r��?�$\�r]�+��	S�
7C�x*� �	��)��;���B�П��%�sן������s�SeE$m���q�PAQ+���D�r>}���x��O�\FxT>O��0q}'! E�-�0#��Z��S��y+\O�\�|#u�"�>C���b�$�[ڌYt���hd�@A�+9�5�*�*|R�� H|p��{�C��0�<f��GbK�����Zr%��1o�(>7�Y�~�(H=]��8J9Tv�r�wX0bi��8�c���I N6�C��9;@?|�S��..��������!�ɂ����X���4ܧ9�K�@���%��J�ـn�������9bC�Ȩ/�T�cƭ�L��а�'�5g��{�`�Zs:�b{����~ �'6���J������l��ױ��>㱷�<�
�)~Q'F�<�����#W��&�U�dt�#��I�p�9���e�ǋ�V�b>ì~����7����\�K�O[�y^,�\ifH��S1�h���wm%G���3�W���k�p�=�v������ĳ\Vʢ���G؇�SN��r�i��t���7��1�،�g�Y񿄞�?���_�����"������ �a�#71ҳh��oj��>��.x�	T�0��:����V��ۢ okCB���E1N�Y$���-�dDR�)>u�Ԧ��S{G������� �l�0��
���աE����`B�@	Fo��{%[��v/��@� �N"�B��[i���Rd�!��0���f�u��a�(�����fZ�t��+��m}H�W]���gNȐEP$Ȱx�}�o��F�WHF�Rm0�+���)e��ۡ�%��2r�Б����k��nO䄑�B����6��'m�耇�7�b]�,r~��5�B�6J��e8Ϭ�y�N'R�T+�w��v7�]�����5'cUV`��9���"��D��OJ=�#�M=��2͗0�X��nݯXP�~l��pw+>���6H�?����!���r�nL܇4"����Yh7mq%z7I��wk���T�W���,�Ծ���9��L;��-��t��*(���t�(> �{�����A ���z�;�Y�S�Քq�N�to�ғ�n]0ɷ����k#k��Y,�Mq���}�!��營 �]w��;����:U��{��D�}q�͡���y�֮�bs���Å,���A�nb�}�[��}A�� u��D>n^��Jg��Fk��NwU=�P�6��8Z�QI`шEjr�܉x8�	4K�6�R�Cҳj<c�i�ِ_����"�8�|�ԟ���?�k"H�&W!��)��a"8��0�sB�ۜQ����Twgr���j� �̧(L�:م��l��'xs?e�&�������Ӱ������O��4
���W�����uU~o�d�sov�9 ���;�q�s�!R�"�/Q��Dj��kz]���M��&6R�tN�e�yk������\WF)9��q��S�����NJ���Z�葛X�X�^����_� Ȼ"��K��:;���w_�b��9�B��jI� ��z�/9�A�xN��
k���qϮ��s�� S�����??�=�\���#PG�J��4�>����OtNu���,�WQT#�^/��$��-�(L+a?����ٞ����/��̹�[]6�A�6�D(GK ��}��
!�Bߢ��Ј� ��+�Dax[(�2��>�_܊C�D܅�n�ׄ�fۢ�E�#"Ek���ˋB\_��`vV�N�ꍪ�/�Py=Vޝ:�E�3��管1h�g��B��y�Ц7Z��%T����������U�ʴ3裦�F���H��t�H�??�d���ib2�����<�����ɋ���U���%��Ԣ<��J�k~�'�\�4k���?ܙ�֛���`-�d�ݻ���W}c4�%�"?\`�}�����LAW?�@r:k���ڢ���������h�`}��@|=�. ��a]����U6�ɸ���l+��L���Vr
K�\A���;WV�8�>�omh��ߦd�����Ld&N��^[���l���R��CE��Ҩ�� �gZ�ޢ�����b�iI찝��B���Fl�.�S�}0 ,�標5�JE6��kIo�
ZiPrjM�s�jY�`����zB��90��p�G�P;�Ç��������T�ÃrC\�4\"O�̏{�ER~��`Rŉ����8�l��b�&���~��@�i��xŕ��|�X�O���J��j��p"�?`(� �-�'��G����k�j�t[C�s1����/HJ��`J���y��5g���n�춙�o�'-���@��Q+�a�۬�n"z�\rry0�Sk�&�fE�����b��
����.�@����W��%F������u��]�������<�@����^ w�!��s#��_@qra�@ր#�G^�H}��A����a���.��̗$�=�W��W���}���2�`�p�6�-ľ��;R	�Q�_�#�ۼ�z7��f��u�;pb�+��sz�(l�+OR ���<��
����s��ЙN��{�e�K�ol���X4�s4���Po��`)]!��t�c���l*�ʥހr�kV�����M4�,�q��&{�ARR$G��r����̴��������S�^�<R1�%�C�����s��,�Q�Q&W���M��I|n�9!��ϲ8�/l(Y5xx*:�e���BMU��\�\2��M��v�{�i��$��b΋�J���F�n8�|�+8�D'�}�7b�\~�sZ�֟lx%:. ��6�9IfK6�Qj[Aq��p�x��w$t����f��t��2QC�.���bj�y	�Wrz�Ժ�ff
m`+�-�o��[}�dלA�V
*�$9'����!СB����XH�-,[�y�  �	q�����L��xrSbu+-�� ��*���Z�;5�`qX��k�K3�/��A�5��B���o�Nd[��֨R|���Z�L[�d��~I�_q`�����9 ^���&�VRR��y}_[��g�}�,&D���x�}����m�-����O���&�&7�G�6�� |����lfKb�&_�h"�m}Ȕ2�� �������|��@.����<_�$?�A|��kx.��|�ͅ`[�˨����=��K�C�:�u�Y��y�W��@�~��g��b@%���D�l4~��L��0��v4h�ghQ8zz��,`�q,�j������k���4���� �M7��,˭���+�rP��w�uN�ܓ�YU�2cJЁ#y��GT��Z�
���'����1���X��⏫�$,~~�$� ������
>�V4{��?K$�o��(����!�9��g(y+>�)"��ύ�VD^�� �-��R*15*C)&k�d-���k��,5-�����W0��G9�ƅ�����÷��j�2�x��(}�F�Y���S)���*G+��s��Wj$���%- ^����<�'�i�J�y<�CP��E$<N�e��;UJ�6��
�-��u`��K�6��u"у�i%�m�UU{�X +˹>u��gW^�j|�!���풠�����)�6�,d,���X�b[��߮�S��ß	gu��x������/P�l��:��y�*�S�,��
G`����bO`y'��(4������'�K�$h˱�\>z<M�A�1h}�佳�I&���ŷlt��00XRw�*1>;F|�..n�/W���(�P�!@n6j5I�����3�/�$m��Z%��Ǝ7s���MC�q�*��
="U���U�&�!�����v�о���h�/�D�dx�+踛3e����j.�>�v�f��u?���J(�Tg+Q�_D~�ǋx�]�c7E=	���
�vG�Ǖ���v�-s�4ַCĐd��q��cZv��*<v�>V	mu��jl�
V4i�:Nt�P4p��C�<�u��x���6�/�Ɲ��DC�+�ce&��T����2�Y���Mk`�����:蓳���F~i�{XYe`V�3�OCa����g����hi�+lj3)K
�����C/ۍ�@*ԝ��<f���c
�'UO.��mB5i���y����z�w�Z��Y�Zx��s�ĸӒg��T���O�Q���ehl����Qܿ� ,�bE����ݡ�|��H]��:��9�\%m���յ�xSv�g'Z��s��/���!]|�hIu-�Q��W?��F4�x�9���&��Y	mM	85肌����~�>����P��)�/4c������^"3��ۭK&T&��}G�~ȵG}e�;a;�J)Eֻ}l�=,�����g
Y%)u��gC�$?Ns�����W�-o�+��+�ԝ~����r<��S�b�I|X&i.�z�5זj�Ӟ�\cD"����J�Q��x:�BR��#�(�z���W7�$~tv�)���:[���F	-PH���Bs��4�W��\e�s����k^��m�X&$4�G7�٧ҧ���} ���!R�>��=hP���D�ŵb���ч��k2=l-�mz��e��bm"������ S.�T}DǮCo\��.Y�3��c1�ŧn��[_����S2�%�:i\Iڵ�iҡ�ۗ��}�$�gj�0(��#Ə�u��k��$S!��4F�XQ��;�|}o��J1��[xK��H�NY$��HͿ�(� ]=媋���"�LN0Y,��;�8���Eq�O�V���
7/�4\��&�"�� O�I�@��tI*���t�j8vu��5Y�:����*�B`䞠�����*�|�ta��D���I�&G��"T�;#����[��H�H���HH��{�� ��SY
�#��ì.`x0�R�Ľ\=P2�4f�׌��00ъ�g��LB��������¶"��Lq�S?��[��C0��}+��9W:.#@
} ~��&�h�mwA(���D�g�C�sϤ�2E�Ŗ0(�&��%#O����o�֛e�U��u��o�Vg7	06�lbp|���h�����B�噳�Im�Mb�Qv"���cN��'US��r)�#��Wb�,F�� d�[���J�ş��ѓ��VA8L۟!�)A���&. ��Iy&2���F�/�t��ۓ؅%����i�|��N������@j{ <��jܞ�J�4r}��i��q�:�z�2>�x�+�Cs��y��8ѕ%��A�*��;��.w�����o�d�. y�3Ĺ�E�b6*M�3NY�o!bY�$��������_���J߬�~�#�b�Vޘ�4>����r�M�L��;�����fy.�ˮ�pI��$��g��P
����31-�)b�j��u_����J�C��
��wP�]��m쟣ɽ۶w�|v*>�+��7�T�%L�;L���~)qꯡ�� �|�	�o8�[RX��h����< `@̑���Kԙ~��|�����8;,��>�{��kr�#���D߬�V|B6��D�ٳv1���gQ��k���G��+A����>�a�I{��S�G||�6?	�aoe	1�2ʎn��f8��P��'���p��A���׌if�R�����F|V��7���|8A	�Q��"�EZjU�d�� GD�S�9�{��ώC�L��J�3λ���q]��_.�q.�T�<Y��Mጶ.���hX
��(ߟ�����{o}@��C���V�p�w���@�r����ɮǐ8b�����j�Z#��N�c���p�^�2SqS5}�w	�ԓ��Ӵ��fo?�j��Q`'��⦪�;Ix^�@l�����O�p�����D�$7 ��3l?ll��x��vǟC�I:=G���Q�X;n/��'YտI��\ގ�p�UoF)o��^����䐬EH	2���hҼR�����M<E��NI𰋉��Z2R�o�	-�e �Ǝ����*+�:P�f�I�~�[�/���afY�+o�����E���2��ֆ��2����p���~����(�{O`����?�lH��������M�Q�bg�P7��
I�>�s�ࠒ�������^� ϴ�G�v)�MO�|�r��b04(�v��?����SN jV�ƟE��P�AJf���Ц�z��"�	19�2[7��w����eԋ���,��GK�8�\̅�:P�R�Z�{��)���O3���A��HM��A����Ǌ��R����Y�Ϛ����DU(8�q���A1�D�84(�fZIN���[�+��߿jw�D�2J&Ee������o�[�e�nn�K�4G�V�\�O!%��sWΠIG����/$+[��ML>��aZ09��˪�[[]�����Z�>�F��l��~ۤL��ǒ�j}�pʺ�K�O�ɨ��@�����<�u7�Q<�@�Fzo�v�wg�����Qgm�"ƍ�@�($k�{�؟sf�H��o/�M�%�*�YJ�����f�z��ߦZ�bm$ ����<�dA�����u����:z��0��cᕑh�l� ��i$�ڹLOәZX�O�]$TFQ�*z�O/�b�t�����ֽ��§'�S����Ùfcv�.�f��w�ZW�Y���	l�]G�+#��.�*��G�m��UeW����(������tBYk=�")+^��C�� �~��*Bp3[rZ�˥�>�b>81�P��T|�9Y�zy���m���@C�{|h�N��wvae��#;�n^��p��q��#�oN@3��[f�L�R�GMZ$5���Ǎ�BS����F&�%�H�5z������P0��F���y2~�����5١�������0@Bΐ7��$����^��)(�	�r�[�^| P� �;�`s��M�@Z��!i��/Ë��T|�t*�ϡIl�B	����c����RkU�ʆa�uַ)_�%�ws�s��("9N��"A)<_�e�RkTD��|����6�JLp�b�g�����Gٲ,a)ًH?���az��V8ᡮJ��!��I������3V���iG��!�Jbru7�Ρ�������A���!D��	D4��;\��WRܝ8tc,����
�� �"���	i�g�e�@ٙ�"6��^Џ�̒�_���!ν<�0yo�WX�YuT9#X��g�e�d{0D�76��1NhΣ�./�	�;:m8��t�rn5�ٮ*4�ɦt!?񢌴D{�U��s�Q˱��s�P�$H8(���Ms#��Co=*�]�"�fSM�V�+=B㯽$T������t��n�������/�rey�R�4iN%�Y�)�R�$��0/�#K�*I?��d���z��t�2�h �˪��z>`)�T�������bpݠ#BK4��_9�n`��P��'��ė#�z�@(��)ю�꒨-xꁠ�b?{Gՠ�J��ۭVݏʒ��GZP��f㤭g2 d,���73�@$��6˃��JWX�C�
��GvH�}hd�W��e����g	�˹E*s'T\户�I�ܤex�����ޯ�� �M�iF>tT����/�]�'�Hz�+����Â���V�Vѹ�/��'�&v1�xϭ��q=����N8��H�� �#�'��P���/zy�8~��8�����8�/�����b^v��K9L�s@gp����^�@eF�^�|*�#j�!�h�$>��nh��g�Ό���)��!w�]�9�aC���5
�Q�p�)�Mz�t���JEI�A7�#!Ԥ+!�;�H[�/��w�R!`M�$i+�f@,�0ݦ�1$'I��� \�w�CMǃG���9R|M	 �7�����c��|���0%ʀ\��-�mϭ����ڗ����(W��V�Kc$]����XQH\�>�iQJP2:�<j���c�ҭ��D-O���Uq̒��E�,��O����Un[�k}�Y��������J�h?Y���fԑJ���ݒC��|v�u��1,�����n�R��q��;�f�d*���p���b>�����f�$���J��Pc���ZLPCk�	��͑���Ҭ
swP�#���*�z����e�Dtd��0�� uz�� LT������@��w�EY|��b�E��+������'�l>��1a�Mϡ���{
�$�߽�\�@m�B����I��;�t�o��Nfy�O��m添��q�A���5d�{a�+f�(˄���w<Ty �s��+�E�Cpv5�����ċ�i�e%>k���H.���������vj���f����s�[РÛ�u�Q�*�T��[�3��۹ĕw�H�gmK ������"�ɉ&rbwj�� M��@M�#�O8<Q!O�Dղ�Pˤ�����YW�鳥�%��-���۝a�`���w��7���\��L�yv�{`aք�0y�-P��sNX�~6��d��O��ގb��5���]<:��U�h	ΐ(�u�,� ����j�x��l"�U[��Tﬄ{��k/av$��D��[C
��40�sxeHD��^"��3��s�6���Hhܗr�a���6`���wi�=O;�Ư:iU�&������L��5�鄁E܀�l��{O������G�F{�{.����hh����OL���2��t�w^�͗5���y%t�$r��a�"���*��䷈R٩��YG6Om����"��^{Y�"�6�����W�V��EpUn��9>v���I}/�� ����[�ٶ5���i�7͞HNm�[\^�P��CA�Ϲ6�>����p�I�.������έ����x@�~$<Z��`c�!�v}�%ʻ6��(Zܖ�a�%����I�Lm����F�7�b	����d|m. f:�r�큸��|ĸ8��NUl%��$N��>�j��5y��_��`���+cW�Yn�%0��Fg�Ž>��l��O����-�=���bC�9���������x����v�x��RB-�{���J��x�=�꛽ -"�!���i܆�bp��W!8�Y�* Q���aP�H��kܷOK�A� �"�-� �P����%^Պ1���i@ %��A�+�1'������� 4�\�XVHR�l^��gVF�-�ֲ�CL��{ϗ�i�xO�����X�)o&_����Hn�P#M#�VB���[���S��z1�����?��յ�U��鉇b�c�5��c�O A�_��_�"/MK�=�G�N�Cn*I�a�L�"p�U;[�M�[?L�65�T��µ���)���_H��\��D=����	o��:����f黋�:`�3's�3$#S�-*�)�m���p���p3� ����/��ZEh9��u%��9`!����N5�<�x5��C]Q�婆ٸV�v/7���S�c��	�րD;����,+�&�|8�Z���'��M���v_��tE�.�����X᪼�73�"�5�8b�+kE��L�Wf�����+=��[e�ݻ���8���9xv�0��/��!�'�:O��vR�����.W0��{�
�)���E`�����D0nX���LQ�yi��>c�K�0W�Ao>��e��}ᎃ&V�W��D��?7��_��~磑�Q��y�ݯ�������=	���)���@<�õ"�lS�<[��l��̧�O~�_\�hE�9�"g�#g�͕�?�1)��W��;]�x����j�deGF��M5a��^om�o%��U�EA��U�����I!���B��$���A�K����FQ����>�_�@#�{(4�5��l2TG�[�Y�H&�{V�Ag�\��e�������v$��Ց��`ԟ�ۏ�E�bH���M�6�Z�P�/I�r�yϕ#F�vF����[]Ǿ�j�`�kU� ����eɉ��6���K�.���&�w���D�Jk�{��J<B�x�����ep�lM��%u)�w �S6`_f� Q��)
���]7H��4��O3Y,�����^	�D#2"MU+�0>V>=�����O�zk��Ӑ'Y��޼�br#�J�jx@���Ķ�O����D�nv?��_�:��()��3QRy��d���)�W��9��G?� �0M�AM�Jj�Y���oZ»݁��Mu�`�>��L�kEîp�x$��X^�O]W��Au4.��|����0��p!V�5�Ю���_�Y9�X���`���0���|.륰`1n� ]�Ef�p�Gԧ>�*k���w�QX+��l�}\����\�l��ܔ)�����DW��o>�i�H�,�},%����ऩ�_�:�[!+W�W�e�>g�Ӧ>P_�B�X��f�w�e���i�]"s���bb�$�A�4�W>O�f���xt�K���,����Ń�.�|F�vm�T�K��"H%��F?`­y,HS�x�1����MLǆ��73�P�S���FRԘuJ�'���@9�cI���§_�&m��~�R�K��܎m>KD���4���C*%�������(��6
Fv��O����'@H�E�~ ��G�!��������[�*�j�5��q�FՃ�¾@�����~#`IH�� �T1�DJ�N���Q׺q��5Wj�I���p2�1YW@ϧM9��)��d��>��=��$w�Q�Q8��m�nl�s�Yf���YT-���i�O��cΦ0dƨ�cwT� ��O��	��`��ϝ�_ޢڶG��$
�����@�\,%�0?���zP�v��ac^��6	p��2OD0>�Np<��Ѱ� ���4�
��Z	��*��"���Еѹ4�՗�W����|ЙO�Dw��F�St,����w��=�Y�m[� >b*]fsAn�����8#�o+��������#z����c��+�O�E4.�C�l��w����@}��d�Y�&Zأ���j���j��8�3��-e�*��nm�ThHy4`]�ݎ~�{H��D�f��j��v����\n�u���	/�-�A�A��@�[�Uɤb�<Mk_��1N��ģbma|#T\��/d�`�y!���7� ^9!���W�-r�st��c,}S`���'=/�U�'ȼՉU�Ng(�%U�'J9�A[H(I��+��buh�>b~W���7���wŻ����X�
��M?Ҫu7bϷW_��ar�@G�A����h[�F𐐥y��cU�@ݎ&~��^	|1�x�Ք(?�R�H �b�b82�ND~��/��0`w�_�^�Bd�W��8�9���ϋ�YC����Fw��)L�&�F�T5�*�n�|�����p���A��#l}YHP�b���Ӥä���T_Im�e�����6��i~�hĿM�ڴ$��J��:=�v��$�'��Οѹ�&&G�Z�4��XsCh���ݒ�N��*,g���o���Ki�e�1��WL1'�g�v��#xAo�� f�o(`*�GP�����'��'�Ld��k�	#�u� W-���[�]�8�N5[fn#~s��H�t�Ge�J7�����kTc(�#6��aܢ��W�t���\�7��p�X�{i��bR{�i��3�Nh;]�.Ҟ���}T�@&���.i���h}6<����Hp*��Tc7�I�P�����(ջiDT��z	.�YGT��/>#Q������L㰬��\�G,Hdr�򶳘S�vƘ���K�[����K�Ir���^�a(�\s0�ZU���v� ���)>,�	��5��}ep������:\-���ǯ�t�{N]�Frr���5���[�3��W�̑�\2�:oq�n�-</x�Iʭ���O��&��@�Jq��EM�jMX�2���>Eɐ��Lo}��=�_I?���o켴��?�$�)��8��O�q0�_�M�>������ߪ��z�G��]btM����v�%�c�����S��8��I����{��A�@v6�������[��'���Yu�X���6x�|
X�ś+q���_F��T��S��g�Z��I�6��n����@7����@'��˜y1LM׎�,�Ñ�P��tK������<�Z��)�Ȍ��0���F�`��]����8�ّ@>RyM�ɉ�іE�\�|s����̩�(�֚�g��^�Q�����cD�|��}�O�S��P8V����j6�,	_�c-��&�Mȿ����F��2e�c� h�V���զk��;�}�i^�/�"��'���HF��p�#�K\��Ua�*������g�ZR>ܪ^Z���"��E#�=0ǎ��x�-��B�U_b�>H���Yyw��%ئ]�"���%I6$:P�j8�Gފ����SG��B%�Q�I��M�`8KLl�f�-�m�����p�K��W�=ݓm;�T_��h��`[��7Hn���Yz	�ߑ��� ��H�2�%�N@Q)Τz\6��Ń��:|@������A��~�p(
X������\x�=G����q!�e��2@����a�^���lX-=�qٖP��fϽ�McyL�f�t�!v�Fe/�D��ޟ"{ �}
�yJ;��t:3I1FJ���I;R�gЅ����܇=3�=id;
7ܓ7���}��T����,�A�
WQ!H�!D����r��3_.w���C�y_J%0�>iU������ ����&D/���5���N�E�	Hh�F�;�UJWLl�,����J��n�9ѝ�Pn�M9����Ƀ�O�?e��@~��W9)������r�dCf3q[��v��^%:v5�f"��}4=��������bi>Κq�	�(~��󛨮^�M-� ��5� e
��0nh�&@�²��a޶ğ?�q���ʢ��~��Dy� oS�q�1�bc����$'q&�O�_������R>̤1���`O��hh^�������*��l��?�9L��T� ���S١�"F�����Y��X�a0TCz5�ra���ڕ�-�_rƷ�E8���Ɯ���d?�u	��(���y� b�<(h��B��4 l*�O3���"��#�Kz�J�W�Z�O�"�y��cuF��}�7|����6��d�&̆�j7D�y?Q�å;8"<�6<�M��ׄ��К"r)��%l�J�8Dl3%�k��v�3�JǋC�aq���o/�Ψ�K���6�����	k�ӤM{{��?�ߑ�[㤻��W S��N������C�����g���`��Vl��2��>���_�-j�\�^QCbX�%�M�W&"q����/"�د!�W�� ���]�ձ(T��}�J��q��Á4�m�0=O��Q.�d,�@��D-4����J �SG�r����{�w�c4~����
XeHjc�Q�#5�G������I���=�fXrn�8Ɋ	��x�N�6�/FF8'����i|��l���Sm����h�#:up~�u�jB�u4�=B�H���C�s08+'�)0]��|!ϩ�etk���)��,������k�ckF����.*G��y4�fS�UZfX��h���ؼ��O�l�뇆�6F��CI����ҟ� h3��@�:"54�@C��|E�H�Q+�^3���.p�������:.��}��_�)��T�х�yl�����@�Yp�A�����Ř��7��N�A&t����\G1>�6Ѯ��X5�K=;3�,�8:Ȝ k�'4�l�R�A0�X�J>	�ߌ8J[����tL}�>��]�����ͦ�/��)�1�{��P�[q���ٗ� SC�CBI >#ɿ�t����n|-y�w�KƳC��L�QD?�d�0�Z�@���J�y�xJeeӂw��$
¨P��޵��?+�q�2���n��ꠛ�+o(�)�w�쭟��3A~1�I�OL��־}?TR��p�`9�o
+�U��z���(�����ȵƆ-����aF>�ct�Kb
���>������Ӗ5��W"�\C��̀�V}7��GB�=y�B_���S����(�J��|P��=�fH@��U�#n�9��!����	�(;$��f���hM�������dIB$�\�%+)z��N�$�ډUA/$��r[�r�$	$�{:��e��z	(v6P	 s��<	۔�7@����\���oD��p������} .A��\F�K�i7����Q�^6C7)��"$c�	���7�6ݷ�pQ���%�<|n[�潌ޣ����Z;!�2�%�}�qt�L��d%�t*�U���ߞė�m����T9*6!E��@TbҞ�|���O/'�ʌ#�+,H"p�$�~���P��빡�l`����v�P��-P s�b)_O���B=ϩ�N�C�<�� :�'%�,O/-�7�R�6/��� ����a���՘��}d,��x�2<��!m1��DӼ(U�=�i�(�&7f���i��_yƄ�
�KKh��S��R � ?��j|DÍ�o���v4� �/Ћu����!W�����-q�!���k>|q�!g������ǵ��2Z�P/4�Y���֎�����;�.�雯i���tD�#عS]f��jV?��ъ%fO�e�E�իdK��
	 z�/�p$��0�)�����L9х��B=�cm��b!���]H���{H�ɬ9`~H��$xw��ءC�\Y@}(�6*��	����#��b_i��Y�d��6<J�*�v���/?9�Ό{��<��q������V*x�0jg��K�n���WhR7
:�4��A<4D��3|]���X �&a����d���>�R�+|N�I����!���T��4��B�ZS,.j�xq��.+����*�?����|���z7m�#�t�#��5e���2�(Kϊ�-�M��jÙ��Hܗ�*IZ�f@;�b�qs7[Qq��@9l�=�v� 2�.�P����i��.��\�����;�2ETX�˘9`�\;E�ד�O�s1��v�؀j�=;�I�
e��R��,���-F:��rqR�N��͆�i	Tc1Xg{��jh8��תs��=n�2����Rqr�U��q�R�i�����]o�X����v������X�|��~S�6�:�u]�V_�<�T���nX�-���
#ޒ���E�L�
 ��N��D�_�nTГ��a����y��y�2!�Tv>H���:ͫx	��3�s|J�/�m�9�3�ا�\Q=:�_&�rH��\�D�O?F��'�~o�q./�>��&�-�<@�M+��A&�:�p!�M�b�w6%o��J[=���h0AG�rL�0�9��k�B2�ZЖ�4��w(��q��G�!Y�l���y��_���ć�������>t��;�it)Zh�W��zѻj�������;\� ]-�9�������En�u���lq,���#�$��$�Z\0_���u;^��HO]=�,���{��EL���,��`'(�v�ýJܫ��K"F���z���1@O�YtW�m���~�Vy?�kGQB�֊�=���S��wՓ���s ѹJ�"m��>��%�FY��
�T&,�����S'�T�~I��V��߄Z1h9��~�#�r��C�Sy ��#gԮa�u>���������yh1�#�H2��Շ<��F��s!��ۖ�%륅���_��Z~7���ϊ8p�8f�D�T*���P�?��'���k�?ђg	��*e^C��+:����b�\}d���3�h� 1�A~�3��G��4�{E���,uW��0w�b���}vƹ9��9�l]�D�'��x��Z.0=��7�*7�����MG�i����\�ߧ�n6U��N5>L�IB���5�j��`,��J·�t�s2ј�^O�nD��%!Ú,½��f��u
�oI��O�R�V�q|�Yk���d��F~+>酃�@�b晏l
�.�,��E��< �>�'l��J��*�k��>'i���6p�ʸe2�s��;��0�QD��� x��8�$�>{����*H��{�	��8��dm&T�\��tKA��}�Q/q~���N׫�]~7������֋Ăle���+mi��RC	�n��1&����x/vY��<iUέ*H����	F�K��,f�sW~#[d�_�_�Y��n�Wr*	�LȤ�)��$��n]���,换~��j�����AZzڈ�Eͪ�򏵃��!�jI�i��%9�@�n���q�"x�O�;dQ�5��5�6+�v�ֺORk(I�@%0�~]��Y�M�Gx,��RQ!���\�??�)*t��S��w4s\)� 2�̿��I�aY'�h���n	��Ja���;�z:�~jB
R�w��Ck3�j�F�׻ר~8�Yw�<pLl�tK3v#3餮�a͌t�V��Y���;�P���s��g��j쏻��9��6��]X��UƩ����΅Q���0�7�%p�n	!���l(	�G�)¸w_��E[?O���nt�l��(�pX�&�\����V�_H����پu��_����&��u�������cٟ�>���3��R��i�=G��TYk~���6��%�9	há�n2��"���<�D�9�����~<�t��y͠��jW��ݤ��D+������g��G
> [?�܌��Ҝ�j��d1�᚜���wr�+��Ne��U>Y�D@���r}9����x'�6�b�0����U��l^���F�@����[P�-xZ�<��W��$��s-�=�/���)����g�ӓ�3$��0��N�?�Ҝ��;��v�m�2sh�+�#�4��D��9P��/<ǁo�]��m�QN��{�}�gv�^��V��1oֹ�8��oI)v<v��-&��>)��w�!�1=q�T�~A�{�Q�H�2��)(Y�+� ��Z(�~��q>�k%i�zS��v����$&�S��{���(hV� �#�}���+�NQ�z��(�U�/�M=���*��Xä7djS��hda�f���C�UH2m�y2��[��o���"Ttr�˖��EO]H�3�ڝ�ߞd/TV����;�TQ�>`��QCj_�~h��7x�����!㓂ق�������̗z�5T��|S�P)�;�(ՕuG���Um���Ә�X�T�� �C�=���RƑ�F����$�6�p�>�#gt&�B
L{����H7�]�φ���t�j�Ckj�#嫂�&�e8³(���?�	�y��MV�A�6\��(8��m3��)��=J>]�<��=���q�ITZ�x��H,����C��G��V�j�ge�[v�U͋�ɂKZ5�Pt2�v�f���ѰHq�Ϋ�B$c���s{@Z��Un\�mӾ��rm�+̼Wnz��m��JBی$���I�z�p��Oo�S�v��I��Wtase������T��/fi}��`T�S���K�xV���x�".! �ZS1��7�y��\��hX�I�"�s�)F?�8^e�O�S�۷�q�>}ZUaN1s��	W�6f�p�iIeW��-��D<`�����y���v���p	��p48�d�'������:T�tP_y�8¨?^��K��/�gx�M��td���m�/3�����;nR�Ɛ��LX�6�G����gDD���t1@���0�;A�f������a��}Ѻ�+^*�P�;�fGmꭃZ���Q��)�g1N�R��j?�v|Jۥ�����z��]�UE�"�B�=k,�ܷ�ceL���X~tT�C���X��9DMN��p�f=c���]9����k��}:f�����8+���O�l�,�dm?�]&�<!uN���	d����<.��BM �b��k6�!�>�lo�4���n���I�]e���H�ܕ���V~�^ Y�ں�:�@3��h�u�5q<��&���9�O�`�y3�C�V���'�iT�����jH*t����Grtd�(Ģa�ȫ�O`P��o2�Lsk?�»��U\Pږ�?���O���p1���p)�_�">�35W7��	&���ɼۍ�JtL�
�f�~�:�+��=СZ$��0����|�">T&C�p�m�|�s�Z9=�o�����B�v	��ɣM�T�h1�6Hw��ҹ�~R��ȫػ��&��(��O��j@
Ӆ�Io�A�s�����A�X���~�7K%��$7�9�g{Z�F��
���@ԝK�$6�k!u���"�1&z�Z:*C�$��RH��q�H!������L�|(t�!�c�?�� �<����R��r�:4lJa �l�� �P��{Mv�[ƒT��rd;M�+"���ǘ�1BU��=m皉z���Pz��^����?�A'�t���&^��������+�Oc�^�QB�5�3K)m���ֹr' ǁ⥓E�	"lsG#|���+��{��@�X�  4�a�7v�J��n����Tķa�*M��_զ�!79+��j)'��]�2�w�:Kz�+^^*u�� ��~�ik���܂��j��p�NV��7�k� U���<�y�e�,��i�z��"30%�*׻�~��y�L`����\�`J׉jW~^�� ������w9��)vG�ܙ*���?�Jf���(|kK_5����Z�q������ŋjNՐ�J����5�����& ;LI��{�4�8=T�1Ǩq��H��%T��Ȫ[$'�ϼyp��������W�.*dC����}�t��Co Yr�Q�y^�����{(|2pJb�/�R%�
:��xD��5��|���Cz����� xۅ�I�_��̍3�3�v��u'�*T
��F�����T=��� ��n�.��:�	�K����I�����<LoŶ���]�3S��Z�*�(3G"w��|�rq+j�=�d���6��zp[ 4h+А���3��M7 H��b
_��I(���*d��z�z��팎�Zפ5:�j�d�@-&T)H/��\I����H�%��Z>��>�C�7{�"�%+�D��0W �jԇ(����u��Y�F-����5�n��@?�cP#�j�_���T�ӊ�ϡ����5�q=I�7"������ʹ�>�h�%�K�4
"�f1�Zm> W���x�ʕ k؂"r� 0����þ��_�p��ۗ Z��l)�mlF'�9v��t�����+��ڏF�\��{���	�ebU�T���M<v��\R.��Ú�LV��������k2ׇ��	���.��Ka���}s�e�_+�� �/��h�[ЧH�a�U�?���f���=K>�h��2��l/���}T���4�Ó��B�d3���v�yn,[�A	x��fG�0�˧���L��3��:��A_a�n�"�P�-��5�Kl�� ?YAK����L׼�s&AY7��Lt�������r�2�ü=�w<\'�|�Q��М	-\a�k�lCẶ�'�屖S�x��8���G�B�S�ٹ�n�@��i��ۂo��h{�Cr�2���X���d��b��蘣f<�|�c�PH3�n���=����jDr��)���~Oq �-D��.6̵�9���c[A@r�n�mYi%-�m=�����o��7O�z/0:j\�"�ȳ�)�w#i��u��Bg�Bo���И�p��U���,���%��B{0G
��Eň�>=����ץ9)���iM��r^�Ë�|j�G$��Xn!�$0�5L��s�!O,:��{*TT�����O*!��>:���H�U�ܷ�R|L3���*҉ȹϰD�a$�hb���3ю. Vu�7=J�2HoA�|D�! \�i��K,׉yc�s+��r=\+�m��g�����R��]���# ��-V��b������\[~C�Ǘ<r�wjvm}��Fp� ��=/��1p4#��j}s~�@�<��q��[07����d�-?՜գ��"(}n��I]ظAO�FJ���KhҊo|M���rQ�룍TR��2���aI��00>�v<�B6[����`�.%��'���86s'���=�D���FO>�ۤZwL1�/�Wᔙ�Q����wv�4��:��g����6@�\���m7t�?��P h�#�{_N)R:R�q(!2��?�M/N���� B�QCF�Cm#L�@���d
��v�	ǡ�Db�7XD�mW�O=��m���Jӧj*��O��
�;��=��3ب|��dW���<�nޞ~�I��P���쑕���B�[{�!��ɠa�#M��926�t��b�d��m`H���&�����6ö��� ��
W�T��-w��"����[��f3��(��5�s��o8��~��a�L��<ï�Om��EN��<f�uǉ�e�|{��C���֫ӈ�Ƅ� �2��,�9�0���hI�$2�ɼpH˚Yl�<�m��|��d6kV�0��eJ�i.�P �J$ab7*��F�;0n3�y�+�ߌ� ɘ�n�E��;�s�5��C��� 4M\��>��Q͍g^��1�{eğE�����7�X���~X��"Wԋ��F�3��h]mSuu}��Q�z��
� l'���~-�}:E�
'�
���le��iu8	�ѯx����0'��=�n7��	�$�!��f�3��"�G}VfX:�� \��@�zf5	W;�ā	���Ԏ� ՀԹ^8�S|:'�q�����c�v �!	p�Jt�U4Q�����pS]��8��YtRNT�{�j���g֣x/3<+�{=����U�G*)0��\�/Tʩ�kx���|�J��A��8�-�*a�G@��S�[��R����E,؄�������twV�����8��-R?hL$U�:c��:Z���}�o4C�x�����ݢ�����/5Q���"�ϙ����1#�kM�a͘>n�2���]��� �;p����&�ulE�*L���̙B:>�V��c��N)ީ_�����c��@	�#!�In}�
��/�\�N�ȉz;���'ǂ�ь���}b����R9�l>ڸ&qx4������Y���rf�^��mkq~u��"�FЍ*U�2هz"��l����Q�<M�Z��?/�8��/�r������s�)�bS��o;j�T5UB��Q�ʻW�S��d�Ds~��,�濾�50$�F�}P�1� f�9ul�zY]�^>,G����dnO�"PD�8y,����)�\��V�'vW¦�Ϻ��K��0���)��=�G<����p���7LTB�swX["�*����6�g�^!uB��ٽ
X$��4�x�&e#m�	v�����.��n:�Rqb��rY!���)4�b媏��'�� -�X��!fi��?43�"�俰ܿp��;w��y^ڥ��Q�<�3�ܟ�oM�PdG8=~壍�ճ�w\�jQ�����ڼ�ƼZC��k%�L�Ǡ �E���Ѹ��������FMo��	��N,{0�)n��m
ep>
C�{��)r?<%y�:�χIoQ$Ϋ3�=0�-Sޭ�	��)*}9��L�rhɐ��
������oU�\/b���=ʗ�]f;�`h�䧉�� �mА���&m�@8���*9��0��h�b8{]�b��U7���&[x��쮊c�Ե�nHA�����Z��tPi��&�bs1�c	_W�Q��������9�AW;��V���I��UId���ʗ-�\�g%���/E������޹����B�+���>�eVJD�݋���������k���s��M�|͉Fܒ�D3e�{OyJ�,մ��՜�%[h�J]�����3��r���E`�ˡ��0��?�zh��GޖrU�e�ԁ��D����E�b������d��/_�t�ۑ�qc���1w6��& -�:����u��{�:��hܰd4���xX�c���P����01���'�u8�P����ۓ��'>�/:׌����8���Č� ϴ�|��Ot�V$�f����<J�b�l�5�ãm���7����E?�x�'Ϲc��]�ocH䧧��i��a<���ݡ\EA�����5"�ߛ� �+���L��H&%��׹&@�.}m����h�Q�*�ih<��PW��}-=�F���S�ٳ=�x ��$��:���F��̈�e��๭�*�1�3GlY�O�=g�F�zi��4�M[)�pj�
m��:hg3R��]e�OiGh+*�G�,�3��gi桷�'f?�)�:��}oE>pceꊴ'Ł���b߆�SD��;Q+�0�f�K@e��X7�o���VV��sR�a:h���(�{ ����޸���-�>���޳����6��j��C�������M���vD����>� �*$:���l:)�I�?�V��3��ԄwdW-�~��1�s���7���0AIf�����F��*?{)�ޫ8����?�{*�D��n��,aڤ#9|3��o����m͹]���U;�Ͽ7����S�Z+��+��K_�W#d���n�B���ߙ��H�hm���C�/tL�OȐݞO�����9fFWc~#�S��}0����i�2������$/����� d��*(L�/0v���aꊁ���`�n	�Uo���ظ�B���7��*�@Y�bX��ϐ���-�i�tO�[��:�j�li0���h��H/ /�l��F~�Le���/������U��mϘ'(�L��Oea�9���P��{��c��5DD�1�<ޝ(�K��%p���hoq�[\���"�>���$w�:3�e��'�Lr0���� #�6���HOs�����v�l�~�"����36�+mbZ�$RnL�E˜�&�@_3uA2ݼ�������*�Dݥ1gD
��mf�k���Fzɼ��^0�}[���g�oˌ��9�*JW��?%��bS�y����w6U�U�������έE��_���6si�Eg	MQ���<iYo�v��B(�4���rJF7�ȏ���y_���.��u3~RD^(��^"����Ij���8�Jׅ≵yV�N�a�Q��|�n�H���`�y�+afN�R��+!Թ05p$��ao�w�ݭf��2a5����F�_\{]���q�;Ur�Mr�>�OgpK.4R�'ӶF\���5��	{)�F��` �UΪ���U�\��)󘐺*���Y8�[�:$�� �@��wrK�Yjƪ[vwC�ˑ7j�d�9����n�M7O�w�0�m@��c4CD�*���?X�N��S��T�G�:79A���I�]��AV��qM�����(��j;�� oN�@����S;�y']�r����M3��]? �q���7�F����a���h���6�L��ҀK�I�����5�z{VYp���"9��O�}����]R4C:d����=��N�z>�]��jc���'0�Ys>d�F��5�녨�w�v�ẹʽU��(�I3I���[�X���X�hLd�&�|�F#�p�Uw��J�-�6���m�H�+_�!ю��n0�k��m`!���a��ܻ��X[n����/���%�np׻�40�.��i(M�q�
m��X��0�����mQd':X�*=�9��d�d�~�M�	�"���S9��e_��p�ѿ����P��A)W)n�m\A/T��T���J�0�����M�m¤�Xs���r��/C�o�� ��@n����b��װ5�}��n�P��0��¾�Ȉȍ*�s�[P�m��U3BD�,�����������������(�r�k<�����VW'��3�,s�LV�ڳ����=0�j� ����0LUW�&��VK��r�ը\K��fjT���aS�j#L�V9�&��o���er>�l9x]0�(��_1c����4S5����L5���0O����%��YXַ���.8S�C�J�b�����%��L�BuA�<�6X��U�A����� �vvB��_�J[���o��a"p�#��R�H���ߣ{}�q��h��o�+lk���P��[�vU!�&��!~��!��~�-���޿ayen,ڎI�W�Z�o�7����3��LzA����=��"�� :����
���pj�<���ttbH��c�wE^�2��6����n�,03��i|>��Ϫ����apM�)�2�3���V]��3t���s��<�6�,1�V6�K�o�?4֏�ii��"��H�6cKA��%L�3Y�C��?�޶w@e�#З ���vu��WN�Ȫ[��d�������� ��:�/?FQ∌����z�<5�K���8u��&l��� ��|j����Ŕ�����}�$�Z�w��ٞ�x�#�p��pd�������Կ�������h�E��צq�*e����)�-@h�u0�����5F�;�cq��1,�,j��5�-�ܳ�^��<KuȾ��;߄Y�r�r@�=#,�6��ߕ��@q�#�M�k.*���.�G���i���8uD��֮%�,)m����g�{�6�3��~���]*B[B�	�2]-�+P<%����k�Mz���`>F@ �;�q���8������������1�!K� ����KR	9e���Q~0~=�V|���������)���^e��Q�	71�wCYЪ��1�|
�-�L{0��"�q�Q���K����;�J���1��oy��H�{�$�Y[����W�s�P�������.3��h�ۗt��bG�	�~G�o��5Ϩ����mP89-/_GU�ʪٓMp;U������l�� TGy%����"cc7c˔��;�!�j�w��/C�K��<��Gn��9�׷H�|'�r�u�P�)��T*a'EsԜ�y�|8c�$��o�S1��1s�^/�v!�D��u٭9{��5�f�1(ҵ�?t�+�q�o�ڙFJ�MK�����o��u�GF�k�5*�E�A�W���/�V�χDJl��B���C���h�	�M�!�>�����z;8�E���Ҹ���y<^%�e��J	_��O%dq��)}C��Ͻ�������w��7�5v#R��B���Z��:8���נv-pzA��U��A+Qq<��0g��U�O.����m��J�N,B
櫲��	���=1�ΔZ۪���s~�jx+�A��5+vW�v]�9�i5> K�'f�������΋�$�"�E�ۃp�
�$�(���i��@2��7Tw1��B�v"�3��3�h�d��Ԩ�������KjG_j�C� -݇,$LPOB�/ڥVi�몏6�}'�/6�RC.A����� ���Ga��Ǐ�F�� Wk@8A�*����޶q�V,�`�l�bU�����C�k6�Bg�ƪ�d����wE�*�9����g�i!`��>����*9����T���	�u{,���=���>�;:-�d ٍ���wWGȓ7�|ܔ8^3��`��T�jSɾj�'�zy�@yˉ|8e�;����g���l�_�.B(Ë�/ۄ�g�q�Rk/D� �0�LF��H�ܠ�介�����:�.F��G�˔�;�W:s���e33���:����V`�a�0�/�c��d��:��N������Fz�)�ws��e�uC��P,^�Ͳ�Nl2�P#RP�Dw�~�#���R����u3�t'�x%�yB1v^-Ę��,�S�uz;,�g/7��HcK*�%Y�^XYPv�����,=��!���ƧY��E5�CU�8|�1�n��Mk�J8mo~��0O�nK2�������o��:a���x�7"C	��41���m�5fҁ�!��P�x�Z�
�c�Dkz�W�(���%���d�3�P,�!�ORC��tyG������Rې�����g�m������RHΈbM�jݼ��!�Y�?k �Ԅ���BO��W�!0ǃ���u1�R݅S_M��a��Y�P�:O�I6�K�wLf�����y����dr��M��Iw��\C��b��~��"]��s@��K.
=]�B>�W���v�>'���?l�9�k|j�bH��f�����ЮP&��F�MS�5��Ye��mBfS��&�'��U��y�������I�&��a���\�T�n�O�9�� �z�T��b3����t�B�[0q1�*��j�V���ϯv�[�CdfL6�e��u'�EȂ:?EQ�U��'��N`k�� �f-��|��'ik�n��� ��\<Z�E
=�?h�E�"���޵ip'��'��ZT�F�\!]�3ߩ�<y��58|w2��q:lKb�?+�����i&���A�\J�"���D�[#���s>l�/�;E5�.�ѳ�qʗ����e�l��[����@UUӝ����(Ÿ)�2��j�0��ύ�ˑ����TF�Ya�Ŝ��?��.Y'��'�Ͻ���@T]��lEU�N�joV�\zmM�N�oJ��qH,��)�Ķ��5	Wz󊎽�/�s��[��̚ʫ.̔�1*R���Z�`9��4���>���l22�H�'�ǘ�Ъ��05X��=={^��!����1/�%��ܝ�l�nSlpQ;�q����c�^���m�`,��E����|� ���
"�W�3.��$8�V�L;\��HD���e�X+���Yı[��)�r;���I�.�W%e��3��(�3�D�#̆��OsC-ő���E��\^C�K���aOqʿ׫����󳪽��KqQ�������[K����/
S���h��ta��WE�q(�i�B�GX�?R��w�#�h���r��a@.	�ҜW�y�ORR��e?=mV#k�$=;Ӻn�/�vW���A�4Y�hHHk�|=Pq��fî @ZAU紛z]��C/�<�\?�NkGO�uހ�����a,���?�r0\�v�q�rC�[����t6�B����Ù�;����v��h�wy�C���5.����Ule�,�s�>B[ܱ���MC���5y�{7��g�"C7j�+W�SL��l���H�w���ԽĒQ�xc.?O��NFY6�L�d�r�K#�;$�aʛ�d.���9`��t\~P�|Y�]V�L��i5^P�_* ����+�3���!SVl}w��S�>��W��(kL�����3��ӓ���.�����w�#�lB@>��`��v��^��t��rx�:�i�x?��A|ٲ܄.	��͛˭��|��e�9�����t������T_c>������8��QG*�Xٜ>�0��Uˍr!�'K}|�nWc�\�+�&�w���?!�y#qȢ�x���Z�|8��7�اr0r��d���{�g?b�TΠ�Q����I�����Z�I��V�p����֌��`n�$���+U�Bd�ph �)ů��۷~С��y�&K���A^}j 8����4��Ӗ�C��E5�^.�%�R%/V-�4�M��&����0/#{��_� �~�<�Wr~�C���&*���h!�~��Ep��If�����U��X ��X�L�{xL,G&f��`r��sONZZv9|[�1��3�v�����-�K�����2���sŻm��Q�J�^_�r��EW��4�%�p�61�ܸ��XXV�A�V�ML/u��oh�0�Bأ+;gH�->z�ί�'{.�x�o���9ջ���M��,iyp
�����9q6�a��֠�*�X�ߋ�Pd,�$fY���S�*��t�MN�!�$	S#�=6݈�@��UMY��7"�eV�I�<�/�cAI��J�sed���W-)m����/3���0gLAi�Ih���-fKإ�x��RbIy��V^\Z3�`̛/:�h`aA�6N&�W�Ξ���q���C	א�hOj��q��Y��2��J.Z��0��a�G��6�ږBy�}S��X�pHiO�&C�tV�:����OB�fg��,̪���%�ç#���c���H~�����֩c���� �,���D���I���2�hOꐉWAE�j`�3������r����ZP���r)��|��v-i�9F������5�ظ�@���|�GW�N�*�XY���`hQ���L,kdq����oER�/N���P:F/�qХ~���b���Ƿ) .HH���A˕)H�Q�ik�*�$�%󾷭���E�!���ْ]��Ve�l��<E���!�O�gk����
�=��6Hl e�ҠK��>��@���_���SGZ5Q�}'�x�������l�A0��Κ�K�d쬝��C��GH�l
�E�f�sv_�����R�
��(��l�y�3�:,Z�d��*:�����`�š;e�'�[h�:�l����q
�}�JzP�;���b�Wx���(��DZ�З�1S@����;���ҚW�"	����][�QH��F�R���s�6�cRK��Pmaiz�����K��/�ssT;�S�5xֿ|rt���s��<�\s�ʿ,3mBωH.P����-�ݬ��)4�zC�d�����KS#��<�t3���Z��a���6;����>�ѳ�Gp�d!,XT��B���[d�gwX�,=�/��k�W��a�UϑSz�.���
r�A��w��l	�Q!-0w����TNĢ��ھ�Dx	<�IX��䙪4e����3��k`]�^�б�߁�R�X�y���Z)��I4;�^��	��e���X��̏��h�rQ�N �gU!�G0Z�s^������\�b�=��l��2M��Rɐ�+��1��rvg�4-l$ƩfdA3���A��vp��SZt�X����̱~K��)ȏϚ*��.~0��	!�qz)O����U[$���tX�����򕙌��%*���J��z�m�H����;�Rj��B,.�j�J9��PF���4{<�'
t��QJag�hy;}�5�G*�MƩힵ|246}`>u.Ku��ş�^m��)��%k<6$��J��Q$��_������#]�N"	5,�L�8��,�|���K����#�u�gIbܤ�c�1F�[�L�i�,��Q���d��Y��T��&�/����u���0a9��"�e�J�b?]0*��f=��~ƨR��f�����xV�]`f���h�֙!��ťݻ6�177N%$�M6f*��t��Mg�ac0X|b4�M>}n�D*y	�9	ӡD����2�P
9M+����X���
z(�z�n-��z�zMJ�3��Raĩ�3���.xd���GzD��	��V��w�c�,��H�Tu�niot�?[��������/�Ͼ�ܿ �[�l�l��vX�)���xr
�i�<b�*�bH���h����SUp����>��˝����1[֐��G�e�*L�+tQ�t�ۏ�<�KZ�Ơ
E��m���Z�%&ð����f��;�����#`�"P��}kt��6.�e�T�N����
��-�ʸ�È��XsJh[nѢ��;}����m�t<n*���|5����o,�O��01gİ��C�f n[D����LI<�m��_Sx��G�-5!+�KV���'��b0"�O�̼ww���9���u���z1�'a��*�cl�x��w�ڠ�n�����xqT��w���=Z�:M{�{�8����RU=}8�X���?���ߑ|?aI��}~퍒�u4��F%�������:�HZ�1wgf�`Fڻ%����J����o�q�X� "SL��[�7h���$��z��{$F8� ո�����Q������;������ݟ��!@D5�z��T��ߐ^p�bꎾ�3d�	N��^cJ<�B��uZQ�p��2b�?��c�qQ�ƽ\Ƙb�B�*'zH�0L8�L�T�Ӧ��*�5��`���`K}^�v�xbVd��q�hەD\RiZE6I��O����d������rE2��INOl��c��\T�b�B�N9��5����Uvg�K�<���@��Ƴ� �G3���q����u<r�����w����!��r8k=�@'�n�~Ya�Z��� �H����B@�	#DB�&]����K�a:2|� �pJ�&�q2� A�W�}>�]Y$O�|2ܹ��`��k����Zjd��xM��_�o��T��w9U8�����ṳ׹}�kD e��A��]�V��CI�.�r�����x�qm�5�'�x P�Hǿ�Y�+Ў���ŔA@���D�5��J�?��n�/o�f��I�p�[��@���6��<:-�,������������Iͯ6�V��E���D�IO~ng�_�mȻn�^�Dy1౦��J�N�/ix�j4R Y6�e'{��O�GeǙ«,�P�ހ��@��Kۘy�%76"�8�� D��`��pf��On\���&Ğ��ӻ���En�|4����i�RPP�>�&1 P&��pz�4�+�����`<ͥ�n_�?�]�!�N�u��P���6���
戂�.��D.x쏡'�:�ڑǊO`(���8��2�|KeY~�dw1'�x��bg&52Ɯ?ϻ��6Iʷ�E��D��3R{����$m:�*H�������n2��)u�ǈ��4N߳�P6�N�����m�U��
�� �y�H���֋6���p�Zw���I�t����3��J+0�RO{'�a��V���k��Syԁ~���I&����d-?�С(M@�"��M{}�h�~s�A�����I�b{>tȴ���n�pO��q/n��o��j�B-:�Pԩ�2k:���K�Q:��$W��`kFX��I���Z����4)�k�"V�w�J��+[4�2 ȕ~E���d�E���|B8p��>E�ͮ���l'����ވ
�2�X���)�y7;���IK=5�2)/��u�����B{�&*[�/!�\:xY��F@ϕHfӣ�͟I�KTv��]\Z
fq7��_<���]�Q��y3y)� .��>oA	� |aJ���\ng�_ss��o��p�x vG�W!cV��,��:���l�/��::Yx��(c�����Ċ��	�ʺ��1����x����w�l�a�O��`U�~�V�T��MP���i�#*�f��
#~�0����a��?31h�7�g�����T�<&#kEl&-��s����c,K-��1\$��4���Fz�G�?�jNs�0"���NH�0��c�3!c��iQkm)ޑ�q����kl�#IVx!��mKD�&�?
�I*�ֽ�%r�����<��°��$�gp�<Fh�.��T�~��"Vs����\�d��������|�(����#`���QD�Y�G6F��FJ�g��N�'"���u�r2ٵ��
EB��p;�)��u�˦i�|��/a��
�3=y��,2-�O���r��z�� ��C�,�+�<f��ӵ�^������V�VeD҆ڌ��gDS�.-�6���ܛ��[��㤠�f!���¹K� �;z�'t�����h")G �HAfW?M�nȉ"o�he�Հ��[�ζ��F�ԗ'���V�ĺL+�`}o���~$���!���`�}��q,���Y�/�㧗ڌ���X�S�����!;��<�/������VJ��9-A|L��;B�I�6c�>�a#Ң^�����_ys��:c=ͤ�el��*����g�w|B�
�i"��3�
���
n	��V�8��'iA��2�u�(���5,��Š��1Eml������s?�z�ӽ�ߧXۥ\�S����;�`=f���J=�n�d��Ҋ1�����e������޴Qi���Oog-F}ob��Š�fM�<2�NEvt�๸�y���z	k�9��a��3�n�=����oA��'(��@�40��%V��
��6z9EB��0c�?	9N�n��D��S	�5����0 8�|Db	K�o�>���μmM����e�IO/��;R�����Cd�f�w�Qk�Z��5�= 7X�+�n���+�BQ�e�@�{ik`��OY��6�F����[�U%�~�n�P��d#�0q�i2��|�T?h�T����Q�AK�?�QCrt�}�_�p����-rB��J�ǧ	�K�e
��� M�U��Ʊ��� ��MtPqT�#���N�r�O�8:��8�"κ�����,�w�����Z�ל�$�����ٗ5-��[А�a���#����2�Eׄw�]�֪��zz;c�0V�݃ϓ�n�=��w��_���.%��2RQj�<���V�����m@A#��g�Dr��19�����"�,L1���}E>VN
D̚�_��Wv��/����#3��>�x�.�x�OP5�t��=ڽ��d�`��Kl{���k���8'4&���SU���P��xn\|�����˽��*��M*HaAFpg������)�����v��[�pD��o�95�c��Q-AQ_�X'{言�ݬw��������vʐ�7`����N{ ��6���S�J��)���f�Te}1���ell�%���9iF�ӂ�'��1�aР1���>DH���R�i�)���1�oh6qZ������>O���S�r|�X�@�)K���ق�y���c&F�Q��+�qY�J�F��ꦫ�[�����D?��B�(�� a�j���x�]x䉩�Uf<E�~eG	No�ON�D�Y�˚�!�����,L-�|K��g.�<O�������_�lm�T��}g���U3=������>b��Z�����`�;nc����IO�Bx��{3��pSf���xK95G�RU�Ix^���'���1ց���K�[�*�6��gAu7����p���4���^���T]��xR��'���f��"��l�	K�2�	��h��c��5�O�A&,�$Zǋ\,l��E�^V�	�.�4�=��m��H�����4!kEi��ܹ�� 0�M�]\Key���F����Qb	�w�``���H���'�@-����lЕ��ՙ��^��FrR_���o�<�R����Qn�!�CAe��k�tq�2q��Ikah�Z����pG��ۣ@�3��}Cϑ-�J�(��Sj6[]0yMu'��(:T��wx���<)Q�.�M@�����z��3͈�I6ډ����5���2�!���m.d�uL팝���w��XO�����fV�����x"ʻ�k<<����Mo��!��I��~	^OM+H�k���� �4�P�3�۰�1p��$�P�n*\k��y6}�K�3(�����k�����.�%��[Ϋ(Do>�I�O�¡|3Vu����S!4h�bh��绺dmZ�����<_�Dq��D���b|b@��������'�)��� #:�T�ˡ�/�� t�8x�\�7\F*g��\Lf��XF�I���!��v�d��綼B�8�2CK�*�I�m92mb
��#k��FC��ќڑ��m�}L��b��'Lt]�^sT+���Ǝ��UPƜ\�Y,}AT ВL�o8$�m]��I���˹���!��5=UEsI�_�js%��x.x���ހ�i:�ml�L��U�qC��U��,kL��KR}�*�W�rȚ�@u���})�����>A�h8���?� 0
j\��݊30��2���=�	��ǋ������ ����Mm|���عڪ}nF����޻rϫ�\��G�]�7� %����n���z�J�ц)\�����T	]�Ϭ�h�!ܘ���&D��S���J�>��o��|׷$��a���E������.�Ic�ͼ�9�Ґ'$0�Ozpv�,u�#{Hb�U�׻K�$�c6r����D�� !_n�Y���#���C�I�nΙ����f�6�I�1>�C�[����|q;^2�*�u4f��Yi�|�$WH�nr21�&^W�Q	U+�X��Z�ۈ�����\�%J�����#�~40�,D�;��x����\L2/! k����3q=nЬ���[��o�u,c�W�`��J�q_�	˴h��<�nM��Uvyl�06"�����W��L�g�t��+b�3�����I�Yz폔8j(�䝥�� �C�#�H� ���i��ѵ�E:|��}Xe�����'��򣫫��v%{bL�v�DZ�s�ZW�PܤN�wU�䵚�[�ُ�\�[Z���0�w����X����E[��&gz�����
��o�f�z���_W������Y�x�b|*�I����	vH�E���1���q���]#��uP�+,�c���[��эk�T�$�b��	�v�(��wE��+,@��:t�b7�6(�넖�ܪ���d���
Sl����K=}炂1V-	ЧNt�/���;>�ѣ�;�����%q�
!ah�'{ܞ�n��q�~�"�Ds� L���m�C<�~�ՙ	�N`	!�&<�n{��h��@���Xu�@�󂞜{��\���-H��ln���Q�L�;?f�9z����W��n4��*C�ɕUFb> z�6,ʗ��?���B�4��f�S��O6*9$B��O��VN�����;�R�F%���|�P8L�hIȏҾ�/&�3d�J�՛�h����=߆����̇�۷Y�E1�R���<΁�Q�p�>�YLW���������n�x�1R��v����)w��RO�����%��0��O޵F��LJ�<ukn�N��[YF��\���m�� |�v�k��bě9�sjroMʢ�_���P�We���wu��d=	������1�^���[���y��cZ������q���.-�Uia.p#�Wc�R]�׼��B�fV�vS2���nx���� ��9|
�o���M�B!ڶĢ�0��5?��HKD����b:m��T���|��4?])*X��O�_ۊ���G����ziw�I�g��K��A��4��*�R
W�i�� ��s�v��厕��Kyo��vd���f�h��\�HN@לO���A��5�_+�ܿ�1�툵���:�C����*-@P'"��'�k��<A�����*:�KR�*D��4��#�S�TG���"�[@�nYJ�fb�"*�&5�,���9���y}^ 9F9cM�yfS9i�;eh��" *�x���kzf��oK�6�=��qc�*;f�-�~n�:��.�	���M�>P�G)�!��&=����|�tN*M��q�K��5�<ߗ^�0PM��IK�.��6�3d���I�+�H#r^�L�����(��Y=SO��ta䓛YOn>\�\Hf����3���������D$w����A�i �1K^��:z6���Q~�c��{�u��Dbt�]�J�����e3���ĕZ���U�J�>��x�A��}��D�e�����@�B��u�����Xh�)��6��������}���p�r��bn �@�@�I�
$<��~PX�2\�k4�e�l�W��%�n��$��G�H6[�o�lr�Y�g�[�E�9�T�����4�� �^z�M4�^�5��JmP: &o��j��o�u�#�퀣����$�����W�Z#H����V8�'�� #\$|�	��݃<!����	�L[����@�Т�{��i��֐��L�*��j��7��B�s슜UO]�8(�5p?���80gC�VWn<�у��S�����,����jĮ���|�9���/�Ch0	A�:�SΒ�d��!����6+����dj�u%W(�9v�v�&���m����������Z��80��yc:�ZƢ�:�}���7�:�If���I|���$�����e���t ƺ�S�9U��,+,������D%���JȚ�Q؈l�ŀ���]�8�Ic��.�DY\9��ZX��E�ײ"-y�Ϭ;���Q% }�J]��h���Nr�BA�W�)�W�]���ӑsD%�٤A򣿳͆�8�w�7P��*�4����l�"-�BNg����� ��QGO%0h�6d_����?��x�u���G^�:��j�x[g"Z' V��8�׷�	���Ѽ'�"g���B�^��9�И8�ܜ�i�8�.���p����h�!u�D��YMX��,��~�-5 n����	����'l�UA�G�Pxd�+��n���+�H!���~$B�F�g��h��aKh��&8HU�K�1�?��A���7����'��� {R=p�5l�}�fN� ɾ{����N�&9���}�C����������\�f+o���[�"j�<��o�5�4�Ug�# ����`��`�ꌻ������p���
7�9��V�	J��:�!a�D��#�+cp:��Uđ��0�P���m�G���v�0/F+�LC�� �$���{��ϼ����W�4xՋ7*"�����Ag$�Y��Y3���,@bx����b:X��u19*�zQc�i�Z�	��#�9:���ĥ�R����Sۧ��Ϟ��c�H�N豺����&Ir3i�*D<WW��Qy�$g.@��p��o9���z�Q�Ǝ!i(�C��D��pr�Nd�r��btɔD��Dw�L!�^�����US�յ~D�C��[YҰ�<�sa��%�=���k�!bv}h�	T5O��������2K['8�\:[��7����=���gO�*�0�%#�kO9�~Lg<N~��񇖴'�=̈)!���/�(�J�So΄�ܭ�g�^&�����0��7��V��>�,����G.�>�M��D=iMEE[�s@Ѧ�M���W=��`iL� u���N�����h���eIx���d�ˁu�ݯO�Ȃ�V�0Ϸ��V��M:�x�*�;���;kv�^��,� U�>������P_E2�ߍ�b�b���ny$m��e纗�˩t��٬��ǧ��샭�9g3լO�a۸��^�'<�������������R�;3�(#`�'��B�[�?I�W�툰',Mp��� 'O2�Z��뒱|_A.��KF!�o`�fe�� T˜�̷�/����Z�V�����o;&�{�Z3{d+#�i�:f��/�,������~�'�c�24�D(���,N5���8:oPO\�Z���� yT�0����}���nV$��u�g3�� �����E�����~�L
x/;чe� o�Ց���d��R���O���:��AN�p��ȶFD��F��^
6��^�I7%
^`���>�����`���F��b��D�NK�c��Y�ZU�i��x�V���~�6�L�T���K�.g��c)�����ͼ����~u���ߠs?br�bTz�"dr���C܎-H`���]CѺ	e^�3~v�Ϥ����>c
�^ѥ�b���q���+�r��$?�7ӷ�U���j������x�
K��/2���N�q0˂ĺ��f��ǡp��]2=#���|���@�=��ͤ��OJ�A��g1�(�G ���6�~��D��xl�"ټ:�O��Y�h��`N+��_d�vJ�]��9��B�Ť���`��R�
��I��ex;�yR2��g���]^JIܿ6Niw����Kԗ;{`K�ay�%A�9���<�A�F�#���3'HB�,�|�rMg�{���m�;�`����b�y0/�:�[��|��0C'}){d�����q���c:��d��j��^�*��}����j8b �Z8�\/X��T�+��y�#�M��C'��V�(�V��eK�آ������WUl#�b{D�Q�Ss�`L�:��5�����k,�P��ñY牮O��*��`������r��=��TM��ݩ����D�zz'ʌ����7��a&�UZH��X��!]z{s~I[տ3݌�fL���Z��[��� |u�G`ѷ^��Cj�G!"Xe�7�nEbDR�}�xm��T�U�*�e�F &k��%�<iӸ&]߼��d�_٦�r��i�!��F�w����hu�d��d��4�1w���
7��/	.�4��iQM�h��v�Nܪ`٩}BE�0Lu!=�����P�ϭd+��a�p ��-B�0R����{��[@v�,w<��&:KL���e�L�6"���u-٘�+��u��'�3H^;�?���⠘��=hgL�j�~x�m�	� !c��ل�n+JoZ)(I�t!Ƌ�޽DV��BVȰ.���a0�c�q��V�MŻ��2�`��K4w��6y�����DGmgj���s�ԅ�X%g�r
X]^'Frd1�*�zh�$ wI�����]<��rg������ \��Rz@ى?����ϗ�W�F;A��U�r�љy�ݬ�����������0	��p0�a  ��T��;��NO�6d�<T_FUj!C�î_�7촞�|C{��!���;V����_���C:`�jH�B ^rX�����:; �uiҁ�ˠ����AH�r��4@k�����ߍ�8�ņ�;��yj/����@j���'O�ߐ���|x/�yZ�r��#����l���'�m�(��o�8��}�Ī﹈�9����'�֦ �/�s���!�A.��-v]A�;݁���rM���4�����H��8A��q?n�q��p-���Zw� /,����eM��mA�3MH��ض;ܱ�Z��F�`w��t�םR5+�=�(���DeZ(d��|rc�:?�q�)�ì
]�>��Q��KXn��j^"��Ed$��7�,�B`%'������:���|Lu{S�0�֩,�kwB�T��K��?��}�H���k�l��+�ǘ���(����xj��n�S�p��^F��ڶ�ثX!���׌��)�����Z�x�,�؍��m�:�ḔC��B�&E���q�J��I�@ ���H�P �K,��7�u��8�ʭ�cqr�aWa �ŔcPWP �9��|F�k��T��^N���:z��K�A�r��ǋ~�iM)o��N�kX���iGaă\A��U��nm���kQ6�k�p�����k�Z�^�4�����M骨Nn�C�C���!�&T���f��I�Z�U�C>����Sª��}�*/�4+�,�D�QQ��p{���i�8�H�x
A��ƍ+5��%�qQ���"@e[(�U1I�h^
c��6m#����ж�肾��O�I2#1�"����r���L����F%��8i�BJ	a�iJMo�Z�d�v�w4B"k�>m��cѵ����3��ߓ��y�˥dޢ~�O
�\0nr��Zקm�X���5�uPXP��}�l���l���]�{�k_A(�r��2\~O�U*�5�gL�#'��/�d\�2KaRq]���X�2�?v8���c���הA1pH�����JR�b+�;�ޡ`&��e'0�R���&j~���?h����a�C���d�9T���9�9K�R�U�^��!UbB�a��DHl$J6�`��c������?��C<�����&l��2�O(�v��{eq�j)��T,i���|��P���ǯ��ʻ�c�c���h�Md�yV<�y;��bxM��t���Q/�!�p���hu�jIW�*��1N��8}�st�Ѐ̫�De�m]�i�[�SK��vCI7WOFTZ�����ñ'�W��+u�w�)�O$>���\��-�j"�Qr_}����ց�3;�"��۸���"{��͞�hU��P�!M����	��KiSI���Ea�(��z+9�'x�-I�ٴޥ��ڛ�ſp8���[β��7���h%�TE/�=Tϸ��ѵZ��B�O������A)ΰ߆m.P*p@N���8M2wn��u��ܯ?^	��?��7��^n�p��ǯ�W� �up3�Ӵ(� p\�Ŋ���^7~���/M��Q������UX�r��CraV��f�[�[.��9X���n��@��I�4���[��u!+)>w{��rτ��=A%�.��ki�����՘	�[ ]�VG�v�Zx����^t<�|�@�o���^��$x<|���y��ʊ�����{�(ǟ��]/
;=f`ı^	ڴf�����~'+_����"����?ykK�z�cC�,�&��ޥ�di�Z���F6þk\�>Gω(��*�eXg�N%�������a??��j�\wog�`�n�@����BS�Ƭp3�(^��u=�7秙��\D�
ǆ=N�R�Zy�~�֋�Qf$�Vt�0s�\9nn��m���k�U󬓧�k[���"(c�C:EkZ{��<�v�.ۧ���Wm��zͧ2ҧ>���3��3a����/��_��l�%�&I����N�d�����ݫ��Re�� ����V��U���0��٬����?q�%�2t��2�έ`�m�x��)$ $�(�J�yU� E��D���Pp�4�p��zA�y;��SA�nFl_IT�LY]?�7X"@�[w�F(�#� q�e�@�Q�p)r�bD��n�c�Ȫ9�	��ߤ~���c�Zb��0`�����͹��7���������+�5!��p��_�~�Hi���H�9�[��*��<~z(3Uu�́zc�R�G�����g迌Z�r��~�U/��'y�@Lq�����k�_M���fW�mPI����-ugB�~�̯�;����b2|���Z�)�q֥�R<�������y���� ��K�B�
*C�Vil{�n �0��{=L�ޯ��ة#�AT��%ȕ�k���&×� {�\܊;7x5��9��������9�\���!z5��Ub�`-t�WC&o�lt�*|&G�x��+��W��.V�n!�>�D�W~g񄀮����4���$;տO�e�݂�1�y��}�!1��@?����\~�\U�9����g"%�s��Q��J�����*$�Ť�Y9w�YZ���c �(IW^��_\��$Qkc{��A����û��S�C��]w&�ʾ0dD^��Gw˞������n�«y ��&�k�Zᦂp^�t��=e|�*����9���$�xx�p%���I���d'��O��2RA����院,#�����ת:-�Hx�\�4�[��T?TJ`�\b�3E���&�g�u�a�~��H����+�ͦ�U�(��xJ�sZ�V*6b8���uQ
�(���q�����)�$h�Y����<���|�RO@��U�_���ҌY+�1�����I��0�G�w��.1R���2i14���)��Q�>����z.(�i�o/���4��t�;���kNd\�U������	��+?�X�Vix�m-#w�xڋN�T&������:N�	�%<͔�O�h�+��Ԟ�m�Y�i7�]��ұ�&�s��Ҥ*�L����]Ոo;�/3H�J9�`3�<�}��qH����
7���v{�����0���d4�!�*5Q#pp��'0�q?�R珥�-%V2
�7�@R�S���n��2���2�7�n�Ɲ�[)X�Kۓ���&��Ho�r�{�ً��Tl#�XNL�X?T�sōC�[��7���_�\���!ԡ^�\���Ls�5E)���("�>.��|l6'�#Ay t�Q;�2'��J�\��r�ZN+�yևͼ���T�콜��1	&�N��ʜ�]b��x�Z͌���"����n�:c��+�R�[>lms���Rt�e���f���h�W7D}���}vz��H����$����2 �#�5ޮ*yr�Ӗ�k�#�#f������$��J|��W�7�HKi�~���)���eo�C|ԥ�(;���e-�5܏gS�4*���Bg��Sv��a���}�8N4`�g��A��S�ct�O[����7EY��OV����T9��̸k�&v�\�R^�_)� :�)�`��ɿf�G��������.[p���6���+d��-x�Qj'�brH��,�:�K�1$h��d&��겳�/
"c�wQ�X�3�=?^9�@�ǎ�~u��=T�o�B��g���BL
�LI&'����#�6��Q�^&W����{��Vl'g	;A�j�C�1v :��5�?��R��t����*7��$7$P:��6R� =+;�����%';>TR8�QL[l@��`s�8� �6%0430�,�"�j"���&�:6)�A�xp����P���݈���OF+�$�L1�׀q����Ys��l�!�-"�cOo?���A`CJ�]i��m���Q���k��,��o�9C�Q�AX@���v�o�I�]B\Ԥ$.����Y���VA���F:�B���KD zU`K,,�Lڬ�a{����El��N ��H�l��Z�������Y�Y+P��i���$.����v��v����w� 0w�����d�Ԥ�i?N?�E���kw�仄Q� ��Xm��/OK�#ޚ��TT$��g���0A��>4��A���v"�yw���R��/��1ˋ���I5CT�Lt���N��l*���&M��)2�JG�b��#�����y>*;��x�]�#?=��O靇O�9����WW��މ���Ć��V!��}�5�����?Rl!JF��,���m;'Ϧ���C�v���Y=|I�%�Ě��gX�T�K����s]}��(Ʈ`z׎ߑ֐n����m�I���O��7jĵ�|��@b�I�6fƐ��}���A����Sc���u�*O>�o6�鵢��;T�h�|��f��`�5� C��ބ�v�o��XT���=��@�}S�3�)��N�]��!�2z ��d�?Ԁ����u4��-��c��1ia�
t�MJ��������V�1pH�Q�Ƣ���$Tڴ�LǪ(���\R��?���O����~��.`���$#�˵��u:�(��?t\51K�_���ٺ�G��w��0�AfϽ@	��Y�/��>e��162 ��ij�]C�qI���>����m'e-�Y���R��̂{$����F����˘�J�Y����Ț~��DF��[Fc�0��o�31�꓍��=�=�W��f鎮���\���������;-�?�WR�sNrp�[�x��2��"��#����%�1l7uFN���,'���4V|��Bb�ܮ{�x��Jǋd�:N�ZgQr9Wk9�_�]S����|dT-����v�Њ1bCr���`�N>k��z����I�L��Z��S�
�6ɡj��y[��H8h�2@��>�B��2ޥ�ObW6��?E�O��h�Cfl/:W*�a%��ȃL:�;'�F_��&d;'a�"/�3����5�J5��om����ײ��}�T�n��8�ZW,ĵ`�̕�mWmFF�.[�X!�Ut�B�������c+9��:�3>Iϩ����pn?vh�s\V�)6����͟?��miȑ��b���?��,8:��pʽ����
����BD��'��cKA`��1ȅ�����q�(��[=jЏe�b�,qf��tpk�9Wѷr�W $���^��t�峒��SFE����iW&s<L�M�hd�=��a�t�v#�N9�T��R�p4�L�z��#*��5ً7���*_B!����c���Yb	:���_��r�p�8�k,�6���b��*!dj*�����Zx$ �k�,��9ψ�
� �`�>X�r�N4�648��_xG���7f*��Jm�\��k�m��l���4����J,�mu:�A�:��O3��;��6܅˶��#U����2E��bƊ�^�����gE�L�;�HD�wU���P݃k/$�L�@�4�v���9~| �c ��zտgF��X�>{b��&�Fw�F�t��M�v3��s�>i_�����-��+�,T�	WY�ɗ�����i����4�))g��BV!2σL$��������*XE����"���KZU��u��>s B#x�i;Y��/W9(2ON���+�w|s$<-�Ϩ���\����0�9n"ӝs�T�e�Ch���τ�B����x�Q#nVȤs6ڇ��(6G$��B��K�a��w����w)q/?���1�h��B�����I�m[uT�\��רP����:@�ٟ�3J4�zBP$��,䞙�S"La��B���aͫx?к_5͈��)��#�h��ަqw[;�گ�>6�D�n����.+���0׽���'ikW�2���:ĕ񸬄�)�	��Y[`�T��{qQ�$��y�*�|�E�J,ڹ��@#�T�yxl`�������;��������@:���\N��u�n���
�4��,?�O͓�QЮ
��O��;���0 VT\l� ���l�%Db2��2.5��cvG�� �������%=T�C��[j��:��𰳃�&�0nrD��W��1����YY�T�e�{���&�z��o=z��1��%�d�;Y[��c�&�߻֔�Y"�������U%|.̙Y�cxv�!�I�劻���y��-\�y!��}�k8nLswU�Z�t$djj��?l`nFZxy�Ec0+�}7~�P�"Y�#�c������X��K��ê97�T�P�ֆg
4A��g��hr�=�ȑ�l�s���q*=�}��}�?s�G���h$�0P����fJ?�����|�d���|�s�;4���D�U�`�M@g!r)����I�8���1z��8�J���s~A9"�	Ug�xpZ�e#�7k\�p�5i�Yq��%�1.��{#S���kKS��-|�Qu�oL"�7@��l>��1lts8X�^(O��GQ�j�dC��.������;U�a��Y�=O��}{L_]Lw;�F�l
�IC���#;e2��w= U:z��눔#aj�/E�	��"�G	�}W�4lbu��-����W�����e6:XQ
°8i��c�2����k�eH���Z����>��g[��
c��E���i̒VM
;�9��q�='H�&��TI@��Sp�#zFk�~`��w�P�K@������숲��V��s�H��8>�7���v�X����x�˦����\6O8�������M;��q�J��������$ŠY�A���PG\")����b�*�uF`M1Ի>�*��G(A,5��M�-V���y������9��p����a1Ebh6{�����0Lm���"�;g���U��� N)�i��F�*B0�:α��
g}r-O8.vSfT�u��[l�^������m�����o {����H�x�Vc�S9x4���ź�}�Fz鎰'$,F�6D��,�$�r~��
�����}&l������Q�u�=Z�3�Q�ۮ"z5���C����(7gW?�(Al�:��{p�&;ۖ��֌j��!$�KQ�n��>���d�����&��A�!u�����߬�Wk��~�͸Dؿ�/�%��^���1��,s����jG�ՇH��`?.�5�c��t͈^�����gnl���̶k�\B����V�p��m��ǧ��/hW���@���z���7Ҩ-Q��F@������I�3#�&@#`^�;���Q�)����!޴��&��J��q��/���a�u}���`�W��#ƈtL0��#�H`�쌃����ҏ��D�+[���� �w���{�\�⡕g[8�R�RG��d4������`M����<K�#��$mROS��r�!d�*���=�����C��7���q47��J8#K	Oa��� !7�W[��H�5͙{�}4:��=�Z�i\fh9����V����6��2��J�f9�<,|����#���M���U?�5����H�2��˙^U�}3�=7��ZXE����ᙰF�Đ��MW�(�}��\$�ޑ2���O�g>Ȇ���e/|�<�w�ɇ���n�Adi���d�.ݧ�I}�6z�,��uQZf߹~�X5?���E��֩��7J����6��.u��� 
�ƹ-�h�(+Ď�׺�CeqA@,_��6]�RZ�[Q��j��lӮ"�j�po���c�*����6��Z��gv��[�'x�������uIc�e�J�����F_�
T��L�ݸ ,=�:;��̞�@]o�#jR`8E!� ��[�ߊ��oҾJ~�����Aa����(���[Y�/��-��sZ) �RG�R
�7�b-J58H{}ڼ� ����Y�b�A�r0!rT�დ%ժ�
�W�*_N.�`V�0�TR����O�}O��9!U}�w
Hs�+�J�E'W׻uuT������2�_��w�E���ͥZ���1ʸ��%�Uz���2��Z���a�_t	�#�:M��!�I�ް�p�$?q�/�o2����<�r�]�=�!<f-P9!N�x@�e��'�����oc5�#c�s �*���a�� �͈�����#�Y�	�LW'/}A��[����P-rH|��Ç;��T�[Hk�c_�"HW�ȼ�#X��H5��ns*ZqG�R �@�h� �� �|6�-�Jd��6|�3���#wv	]���jͪ�C�_b����̯�_���	�EM��I��,�}�O��hsK�s��~IY��װW��5	5{dY ���?��W��z�5arN���7�Y0bk��9l,�����^��3����S���`�ܱs;c;�2EQ�@?[� �Q���(��b���m�ߍ��-����zl2+�-8ힹ��XEy�k��lb���<��!��)Og�;_�yA�h�E��=��2��i�g{=ߛz��џ�xH�RS*t�F@����+�+�&�Ip��:=�-f�*�[dҺX���ו)*GK��65�I�5�r�L���������6���+��}�v�J�5�3�t|Q>
P?�(�����v�Z	���&IǇ���(��'��#�^8����b!�
	����+Q���>��7��Oŕ��cO�i7�<�X�Q�$o��a���Q1<�Q���kr�m�2��De!�-���:|񓸏ī�;�AG+Zw�~�@m�l�	-�ν�F�4k5�͕�����c'�-�ОEn�����Kn��Ξ/3f�]3��<G��a������*��X2���d���v^j%�'VJM�?M�T}g"��gkZQRW^�t�`)��K��Ce���ď�xң�0n����]��,������R߄.�"����ۙ_|S?@�X���+]ٱ�}Xi�kzig�����g(H������s��'h��6�JVm�D~�Tqa|�rWb�����q�_�
*��ru�����s��b%�KT�~\\dWEc
��I��I��
��-�]�%��M��X� K�N�gR�[��7�t��$���#҈l������������{C�j�~+@ڨ���1#���� �7�7�P�J?n����ԃ���c^H�{���;G2�g�!�	����h��>�YX.0��Z�M~=-W�:��꒢� R ��A�/��r2D�ؒ3���J�g��k��B��)�'�Hm�8����O1պN[�FM��t?�=�/������~��[������őu�뱨^��|ۈO��82�`YO�߬T�8�����(��ί�<FP�HSn^����7M�ͅ����Y���$�u�u��%���Aq��"�	��(h������>�D����^H���w�*	�wF���JMYpT��xmm��b�߉���n���l����4��%���K�e��LUV��(oy��k+k���# q��)���N�K�LZz�+�6C�Ej;IڶY�����LU�&�6������zR��������B� u;�U�<�]=�Ǉ�dX�o�|˹��,��篾��v�Pn*֏ؚ}1"4��{Tۘ��J�*x��5��.��t3�tU">r�"�?e4��y�:��$�g��1���N���d�Ľ@��`� ����Ҵ�y:���P�KB>��c��.��Bp�@VN�����q���|�؅������l>uќ�\���S:.��6��8�>;v�Z����$���L�Z��O�0Iz��!��TVx��rMZ�z&
8�)t�#�꾸���Cg,��28����`B^�˹��j �	��~ӱ������}���Y�S��j'�ATCʶ�nw<gc� X|�F샕{d³��zU\���G��Y�'P�/�E8t����Zp]�8���E;��K�h}9n�d1�����T�n�ݫ�V�6����+��x��>H�ͤ��.���J�����a*�	1�����V:�a0�Y�%"���h-����_��(�Uw��������%�	�o��
�C�|w�ﾭ���K�0�̶���.s/*�nQ�xY���ԾǵGӑ��S��XPuT��+�a�x�����m9�`9��=ϗ��ٝ7#f�QdP\��ʏaZ)^�ɭ>ε��_�/z��勤{,~���Ӫ[+�J9��`)�w��Vlv�ђ�.���Aq��w����$/��t
�{	�$(�SSLs%2��ܞu���P�WޚF"S�9���wrkoQ<��Ќ�9��Z�ֵG���4Z9��	q}Hg7�G��R������L��ج	��n�F����{l��&DHR����4΀�BnTB�Gq��p��
+C2���Ru�}�Xvz�p�쌻�N�� r�j̄�+�ؿC��%��n҂m0/��,}I$+DI~����o^���G��!q9YV.��q˨|��<(A�?�j� ,WG���m�t�K�l�4z����X'�*�����+��l����\� ɿ�������}k@�����T_���ڥA2m�=%3�o��`�@�M�ך#Lh�pA���)�y�X�ޣ�8�s��Ӏ���6/�f�!�����x���e{��α5�O����!n�m��Q*VJ-HC���~|��МW����;̭�s`{��Λ��Ȕ���:[�p�LX4(7��C��������g�l�G���[�Θ+�{n�,�~-Q�[����u��ہ�G�D�����b�z��V�[[��0����{*/�B=�BP��A���ԏ�k�V~�W�B.��a ��-J�qn���ǡ�{��\4�4u�>0X�Uo���N?V�����(��C#�8/j��7H�ZP����Kg�Y�x2�Ө��LP�i�z���]�pz>�������l�jw/T���^?S^Ϻ�.#��6��{�FKbP��0�~ʌ;�D���_�*po��r}�2? g2�'m���T�=F؞5���K�����"Aě���%��q"����){Rel�G_M�T�@��T����-yb�>�o����h�~���q)��ľ�)��Cs�bU9��M�Uf�X�9 �Etp���<�P?��Vv'E�;.	����rj���[�o�Lz�j��5z'���/��{v����U<�q���7��]O���&��ٳn��wTYPq�O(ы��li�e5Ѷ"q
S:#f-���Uxk��-3�-�1��lPv����phlkX���j��u�^�/ �
V����l;�e:�=�6R��S������Z_����Qe`�9<6�����߾&�#iՔ �6�r�ͨR� �m��/�Ŵ[��m��S$�rA���]Va��вhU����6�i �>�B�Na��-S��Qg��*��`��b�r����j�]�Tؓ?J��O�7e��u
�$�{XE�eI!Z;2��!���$b^qzУ�L�Z��E Ʋ��D���og���k��ki�Fkj �( �n��U΋��/�8���Vz�T�D��&q3~�)�4��c�����-q��b�xgʟ!�{��54��ڣ�P�kݵ>��Iq�R�!/;h�|1�����C�}4� ;Q6�p�-C��[��:.5�_�='(w�bal�[�B�	Qç��r@h?���\I,�؉��J�	N������3c_,0�|K�.�-Y �Nh�"����)����v
v:�IH����}��O�m&��Ə�SЊ��0-�n�{��K���Yk�� �m���ҋ%2?�1^͌U0��DQ(�'O�5s�0��<�z�Յ�4�C�M�#��rY-���_4
�'�B��Yi�M�����N���\� ��Ag������r'@!2�)6�5}����<���U%ډ,v�P���.'�Fܺ���E<�.ԁ��1�:�.��7���:��%�v&�#������M
��.q�:�U���_\�����q��6�Y1�<Ȝ��@l���R��r�C�&t�%~[:.^���@_�q�Ԩ6?����>i��y��ޖby75��D�]�Ne��R�0TDn���<3�������>���]y�����p��X?�����/y���^�����mm{�G��,��Y|{j6�X�RB��Y��BxǷΟVf�����aO��,���ɝvg�f%����Sb�G�
0 �+����%d�庠�nQ`��M  ��$��	̡M}eX��*���t��}�K5�x��%	�_I��)q0^}rj�鲸����2���/����x�d���H{�� �[8�v+�c���>�0=�휥�N�����tOb�$�W|�}�Cyp[awS�3����w=��Z#-t#|�'z;i��{���� �._k��Rd��̞0�Z������##�E����hF���&3�;.)<���\�(F���;K�gc�V9�4�f��6p/�`T־u{0:l˲v1#r�z)e<pV�p�b�h�����!c~c���f`Ԃ�*��@�?�א��bH!���2�F@���io7J=7�]4��Ë���*�f��-���]E#N����qG��f�������H<�$�&���P�+M	�1]JA�H:ܺ�[�]��^��%��=��<'	 <��	~�ҲRHM���&�	�K?���lL`&�z�x\�E����>w���N��$.z�j�]Jĕ)_V^D^$�ك�r���e��;K��c3��IӫE�p�d����Z��9�^�I��r�8Y1ڧ��jњ��ɮ���L��
��T����G�� �8:p��ܗI���[��56�)=���*��N#�������.o=�-�	�K�v�vRVG$(����u���b���3��f�2�i�i��� ���&��D�aHҍ� �8]�#�2��w�s����I�/����o�1*$q	q���@}<W��`ѻ#�&B�K:��/�ȋ�A��-�����YІ]�?A�s/�ɕ�ˇdX��b��<#n&��X	 �r�C|V�T�acGG�A�߰��sз�D�%������k/��5��59<f���EPM�=�`�G} *��Jn8�?q�f/	�<v��]~FA2���23r�51�N�&�N�W�zk�r����@�?ɭ��7 wv*�^w�')J�+"%���M+���rU�n<�πi9-�f�A�?���	��[+�p��`�VY������\N�%
�\wym.v�ՀcM'����N�7��G�k�[�)3��h!�2�t_A@��h	8�65b���ϷJ#�)��oǆ�!�\|���*%	9�_J����<�;��H�7Ev�?�x	�G�s���9��Z��,Fw�E��D�1E��'⨄���[]dV�B�/�r����k��|�E@��k�*	/�\cU�۷�M��%�L)(�TZ i��X1`��H(�q�E\�\u�����V���<aHAl�cjy��9�B:���k����ܨ̶�:%�o�_�u��(����OY�]�3�&�Im��A2���qO��,u�]�g��)�O�e��y`�y�Ԍ*���l�b�)&�]������K՟�g4Ʉ��~�<���ަo�zB��ث �ĎC;�V*DP�����󪸬>���2��P�D�X�H�+�`�-��LE�Cآ���>,L>��~.j;q��QPdx0��ݞ���?7��Fu
M�k|WV������w巚8�	�P�f[�������D
��b��22 ��.@7��X�!�i���l6x#�K�M�x���Νr��A�R�ۑu�nb;qa�
�zR����y��.ln ?��N�D�s�bS�=!pZ�������4E�s7ǵ:*Ӷ�c�7���/�22�zy�|ڵ�ô^�4t�9y��t�_j�BWb�2��8��+��t��E:�0����}�K>ocPt'�Ca��H�E�n<ۃ/O/
,)��,;/�q	
)8�+����?�T���7}j�Zϗ}D�u�a��xJq�q��nҨlB��#UTa6�0>����p�8%	oRk�Rvj$Z��n�I��{S���@��W2i�Z���5���M�:v�F5��`�+Ns�qa�\V4��PN�Bȅ����B*K,�[���\��[c;���B0D;��2��G��rf3�*.����}����4�<����8nܤf��4 ��P;ƅ���������^�g%��۽q����DE�}24��ˎ4'�c��9Cl�jy)3l]@fK�
`�]��^;��(�� ������h? �����JI:�Y�0R�y�
��nXM��YJԧ��H?����E��m��m �R��J֩��t���[�i#N�wNa����|0{8	�E�Q 4-�:+ +z7���-�����"M�[J��?�hH�F��]����uG�W!�:�ccQ����<t�+<���C�*r��^��FӁ@PrRuIH/��J��*x��b2V0iͭy�k`#M/���o�^�(�ll�}�C�1� �L5�.#]�H=$�h~MXV՚.�R��l҄�qg^�9��<��\q*A��fτ��������5��6�t�i-�'�ٜC�P�a��)�Q�l�W^ʰ��xI�'aݮ$��������h]\�.��Cu-*��� ��h���[�dH�4f5A���I��=.|O��⤴���Q�R3 ��W���F����#K~
a"Cij����CV!,}�k�I��ɪ��L9�d���V[[�,��Τ�t��"S+`~�I?���I���<��ʋPS�%S�񝓃W��^)�e�v�+}~����㊞ƪAGD��F�wN߬��#G�ϵ�R�����P��O��)�;ǡt���~V�ƶ��>�3�v8񛢨:��:����%��� (وÿ��b�c��������[� �Š����mj^G���є���y�m��]��z�PT]V�׃��@_҈^��Ż}qc�N�\���(BX	�@7U�U;��0 e�������Y�m�4:��U��^�u �Q�'3NA~l�n;�fq��Q!���B����#�{96���*����c�IK���-[�w���n�VQC�tF5�X tE-��=-]&	3��Z��S��a��rŽ��`5��ɘ�%�B5�]�K�'�NA˵���*���b���sӷ�m/�#6@���m9B�l���ɱ���N��c͡���tzZ� ���*�K����T��L�f��B�;��K2��R-_sz<�U!�R�G�M'���GS��H"['|�d���eYi�P5�����)�V�j�XD������r䤼�x��Y]w�ء��ێ���]�l�6�����r��#���5��������EdQ�t� ���_M>~5q�K��."�
�K���-�V�gPy9�P�R$�����z�����_�d����S���v��ao�A�ѭ
~X2�@�B���=#�/�����>K��������e��f�AFM��t�*���cKwE��B+7��Fʦ̫k����#��P�֊+�����ٍ7ڶ�@
��X~G���*�,��LJ�x�~Ah�ɴ���?�7���o'ɁX�Bߞc���P��^k�����奟?-��@\��5���MHs3��K)���<��'*d��<�^��KxC��>c�Pޡ'iX��Nz�3���[.�D���_���PE<	�=�k^"���|�/eF���;��i����.��r؍�:J�@.��/0i�5H��R�d��OXXP���{�J}SDM�O���~��`й��g&4���-�x\Rǅ��:}��D���3L�~�;�N&��EH�l����Hb}�}oЫ�|�Ё���7���)� .՗�'���e0�$b���jϢ�Vǯ����_�_��(�L�3�����{]0���j�QC`���l<GGc�6+7�B�%�&��j��,"z%23��+��2����a��d>	��f����e5@���z5X򓄍Nk^�X�-���=��uy��%ZZj�i�ԕh}pI�]B9W#��.+S�)�zOz9`�U=Y~�NeL���8K"j�Һ��F[���YD�3#��	���F�Ӂ�o��[��-�dW��0��	u|�9���Đ4�L�#A""f�lN�m-OƝ�
�ʪ�_#8��j��G��
�A����і�~0����-z@dN�Ez"�A�Yŏ>�|���i�䠚�]�b.."�U!:�t��KB���n�0��Ĺf��%�Qtb�3	P8D�K�
&��F����`b��*	ٛ�"^����>��<s�o�#��L�
w\D�1XIfXGHí�<�$I�߷����(��NK�"[�h/o���i��f!@~��w�/x$IѴ@m*w�0�y9.��٢�'��<��ϟ� �)P�gE�HW�X�Q��&��.S.fs`�yU�6��Ý"�����F2�cS\/&����'@���潁~?27+(���7د�9l�+@�����J�4� ����<�[l�8�!ft��A�����!tb�xȽ����фT��v�=�ԣ�_���y��B]#��):{w�:M��P`�,
�͏����˷�^���6�%�u�	!_o\+x]C�En��ǰ%�_7]�s�o���y]�[99�6�������B3����+aW�%�n&^��L�N��k��C��꾭c
e�����Hѥ���W��p��N_���>�|��iS*͈8�d�.��¿�F�H?ͥG|�͞`k��Όa�q-����|v.��:�2r���c�3@@�d11�n0@r��Lm^�$&��0�W��j�f�.���ne����,-q�k��ހ�~dN�")�?�MD����oVDO� �Z��E��<��Bu�~v_w�ߡ��%[�?����J���d���e��	
�Wo�4#����DOpҞ�cSPH��Q�m�==&	f�
GtR�'
���:���L�9���.gi��ZpG�z�h�)��$=�u�k����v�c�0k�;qǹ�s����E zg|m�Zyᇂ�څ�s���iӰ��)-rt��� ;�NL�jK�T�k������4.��aoD0R`� � 'ؔ�����A5�v��d<�Y��ȸ�������U:q����	��Y�:�M2��d�I,YCUf������r�cz�]_A��O��a��e�@i��D�'K[y��ZY}�3%��;DC��i����2C\�����'ȵ�f��v��v����726�#��Ё<�������˥E��wU�#<Rgyx��e3&�\M�����l�x�����;wZL@����-���ڤ(G!�=8y��uG=�5�)`-��_�ڪwa$؜�ŒB�~֥�-b��B�S�~��dJ�/I��`9�󈋹�����Z[ڱ����2��[��Pm�0���>G������f�
��5J4�K(�[���Y8L?�Δ�ؓ��y�h����a̠�/K�l�9S��PC�^%��Β����-QH�1>�f](�+���@����wfl����X�L.wNc;�,"F}i�6�\~��U�l�g3@XO���=�Yd��6�B�#��zi���S{��{����Dާ�V�2�s�n�d�畱:��G��<iA�P��aߝ����:?�g��#�����~�<���<�����mg���R���sk�P���Ψ���0��0C�� %�"�D!A]��-�Y���R�LF6ٚ�}硬A�W̢��(�����F��&I/��Jʫ؞��qҎsK��]>���-&$,��J��?B��K�
���DZP8�"|��(J�x��a���Oٟ���Y�tz�P?\�����~�v�=˖ɭMG�h�4��d��2]Af�p��0x4!�S�|�Kߨ�XYs��!�͈�\��l��])��K@ո׵נ���.�ɉC���a�ޤ�jm��(�F(Dp�_ѧ��R�v�۽Q73��J���P������du� ^+���9��4����䦃��$HS�ہ1z0���'�E����4����+��������	K�hw��\4���N,�������F� �e;�4�{��4w��}�W'������%~Fҙ��v夊���ϔ_)&���PF\
��+��LO������|>�5)IE(ֿ�]AL�>��.ͅM�5���3���?�˂`�f�j���_�R�墉��ĝ�7@yc�B6gН�cr<8��b���Ǹ� �r��2(�o3
���-A`{�֪�vp�3nڊo]!x�^�5��^0Y� M�bwG��Ė���n�*}~>.�B�����A���9$��7?l�fRf��>�m���ǁ�.l���R���%<.��߽��PG��\C�w@΢����װ��3�3�i'���M3QhS��v��ڼ���$F�7����6�M	_�v��	�̺�µr]�����R�e+��7b�D}6��W[�"�95\��V�h���w�J��d"�2T�V
"D���<�h�$��;�N���p�f��:��`[�c��Ұ+'Ftzv�L6�2t�m�������3���hk�}��>7� WRϏ�B�J6�����O^��������#�|ր��W�$��@_lBE;�n���Az}��E8c�u��u�3Lfr]L�<)wC��.�T�6�]����<0�Ű�=����8;B��J���R�"�Kt4��x�H����8. ��a�T]�vA)Ȅ!�'�؝�����L?�!FB -��,v�b������ h���@��)@�� HvH�J���L�F��ۃ�����<���v����}��S�����	ڎ=�}�ۂL�ǹǇM��f��N��d"��ٸ�r�6��j̼}<+4r+��4�H�����c6�iFq��K����W��O�̂Pi�*"�ξ��Ynt����}H�XR�E$�hH5g>�)?��[>�:��`74S/��@�*��(&p�{ѺV]�{���y��e#�kKut˾ţ�� �*_wE����f��D����xo�"2�h��T��ʡ�S[�hTm?y�zbXqJ<�$~k+L}8�N��cg�����|Hw�Q�W�t��p����+�����_�lޣ"�J|���'�H�z�[l&��u�SIq;�;��'��t]�$�)1@i@E�mpp#�5�� ��֓"��UU�������N�kM`b��'2@�M X��Tȶ�t\�YV�&X�5���ߟ���q�;g��Ɩ��h�)NYe�O�[�?�1�F]���hW� X�`ˌ!pf�y�L��Y��%ڠ�5So܎0�Kl��-�W��&a_�U��v��x{r�4A��GY��@�����1Z:Z��
�>(��j}�u:͆����c0��r�,�|.���U�_ӱJ�����
��q�To%i���1����.QM��5p�'JkX��)y]_ux��L�nAQ)�i.�	=�.����p#����ѢLK�zϮ`h
ܣ`UT"�D�׳k��H|?@J�J�тU;}��dI۲i�䀅?
c�Ѿy�W�mPj($x�Ǿ�s�#6��Ȣ�cJi����J��h[-��-p�>s �"T���J����)ϻU��:��\���="��y8��Ā�Gۀ3�5��^�h���̔�-�<��mV��n]=�֜����t�af�{����%�@�0��m�6f�K�� z�}�|�A���@�*��ZV�a�r_���h.d#Z�j[#�U��F����%������V�\�H��mo۲���ۓP*���-ѿ
�S�'њ��s�
03���_���ߨ��Z^Z���FFo� ����=@Z������q#��F>��%fMe��<k4~x% '��Į��[ˢ� ����j6|��W�j�A��0�x�ċQ�f�,�kXi�n�Y������ѪvǎXTW�#��2����2&�v��������(�`���ڀbkd�'�fK�Q^R���Ŏ!��&��ʧ����,�(^��j=�����u=yoқ�9��u!�▬�-�KR�Mh^��H���8�J�-���A-�:_ƎBb����I�$�A��V�C��02ƸmQh M[aLK���~�u��N��t�;��� �]W'�]��8��ί�Fz��?�#���z��6�r�OX��$0f���������?:�н���.?�'x�gb���C��;0T����w�u��I]ˤ��5��њ��<vڳ��9��: *J��,1�f�j�Qγ�����厈1Ԧ�I�����N�i��Yy�X���h��M�9�3��.5S�y.���W�;ߓ��,B���,>�R��2��藂���Roq�i���L��4��R���� E�uos�!;�0�A�a��:�]��kn��$���͎��M?����G���j%�,%y�f���z�Λ,H������Tl(�y�[u�pL�8<vk��J��"Я'�|�""t�Њ�����f��d �p�a�su���4�ܡ��[�:7?t�J
sw�E���8d����I���᠌���FZs�U��`|����{��J?DK�#Ѽ�_O
ѝ�!�����y�`�	�=�����}]z_f澸�Jב����<G��5j�Je$��ZY�ġ��5���5l���(L"���8'_���h@GE���9<~ֳ8ZӐ@k�B?��keK�Y��xQ�p5�W	M(�_�!�U�:싚X-��-���
)��H�@��N�V��/��р���D���ܵj*��wuǞ�:%��=� ���
��2P���w������7�K�߮�~C4L���c����˨W��5$0i���-b0E=1b�h�j����iAX���}����5{\�I/�.!<�u�����nT$��L�Z�������9P�aRX_*�u?��:j��>������GvԾ���/���{9aYRk�ؑй�������T�Ѓ�#�oq�tQ:5\����d�Eਛ�V����9�f*4��r��$b��F;/�k;C��\���Lل �照<���}  ).C}~S�W�$�@ǃ 4^��2$g:wZ47/�j��C�?�u�F?%�@����m�]�S���%r���@b'8�L^Fю;YP2*��2��HL��}���-)�=7�����*�v�v��}�A�}ğ����ʜ��V���O2!T�aR^~��bwBF�t��G�F���O�;d�GM�U��0w�q@]����L�o��m��~���N/�|��m%3?M�<3ZZuO���y�� ��0�����=���O�ןs�K��nD���5�`FM��1�s=��JQPꨘ3�����wb;�����N^vvJ#���'���i���t[�YX�aMY.�����M�V�끁�癦�7I�Y�5��5A�����-:ߎ&/��ْS{�*��&�Zt0G��〯*GGkk����i�7n��܅8~V�r�cL�R�l�m!*��n-X�x9e^�n�?�YA`��`.-��ކ����T�-,O*��=���Џ& /��{��b
3���!���E�r+
�k�"W0�4�3V�!%I"��p��C����UbS��(�=C�Ӭ'�����{�ߺ,$��=Y�Wn�ޒ�~�]�K�����\��9�����W�0��wN��z	�P�U�f�Pe���o���_��P����:3�ʠ}w' �6�G�r�65�$S�(f%g�[R�0����/��PՃ�QU']d͈�O0P(1�� %q=�'#YRڄ�FYgt<Ow|	ci3�8cq�>6�Le�į>?r�X��r��y7�J�Z�N��L����yi$dh��@�2�T����J?UN	Cuj�
��M��������r��/��@q�$U���T>��o���~WT.ϤjG�y ��ޭ�u�߯��}+�9�]� �Kcp@�"�v��3�1l��E.$�,&dQ"F'" �`(Ϙ�9�90f�4��Wu��	}_��^��9�,�O�E����D���pkF�-\[;5�����	
˴�[��NR��eP�-����n�F{�+�b%�S���[`�g�q���������bT$>tA`�T����O�Q���}�Ï]j�f�/�%��0��~�%�Z�{���/{�/��uG��@��8\up.n�)�<�kS��	��������
���!{b���ZsV�~��X�AaU�e]�q	9e���u	s�=�8�}�b���rIPJٕ���h=Lx�b��Fm�a�23����q�o������Y������Y D��0ə�-�(J5�N����na�@�>���a��ׁ�sQ�$�ٽk��@��D�B��	�]5��^�L�q�q�-�Y��Υ�8�y�Pd��.RX�J<���>c��;`y�v���<��~�<3�����@AV�bp�y��Iv��E��q�X��L�S�V*k��~� �� ��^��"�%Z-�RRb���B�Oo���삦s!�Wll��dW�lM�-���&s����O����'�~mY�WL��j	��mc�к��Jc!u��"�.n��=�/��~��V�\�?�����NxzeŻsbL魫��)i�*J�e����Tl�������1O��Jݧ>\{���R��u�<<�y�.z o��F L{�h<Ξ�>}2�L�����U#��C)���}��_�x���~�= �k����`1�%�8&�39>�g���y�w]���M=8bf3y|�" Iu�q�)jW��X~�SN���1T
�۵XRcC�j��P����T�!H������.Nҗ��P�A����K�������ny�~�r%�s�Q����?�Ѧ[���=��֐tȟ�<����,g�@'��74Ѡ�j�:8����=y��꾐���<�U�jQ��.xOk�I� #F���Hi�3{=P���/���Y���B$>�D|Ԝ�����3c�<�&�-;����J
]}��1�,��
�iN�TZ��ռ�#�g���ӎ�]{�(��:Ƒ'���F�+&��#���P�8���5���k��%�[�tt8�y���+�_��~�YV
�|�4^�]�gi���ukF�qйG,��W<�a6��>g�iY���K8�Ӈ�Pn[S/r}g$M	�L�7ӯ�<K�:�d� Z�t�!�`���O�x����L����䍈>��'<VGn/ �(��GݙMf�v�:��>����C��%�x5��Pi'������pd�:�5Y�eF7V�"�BP�<�؝5�T�2S/c�b�/�g�J���6ҹHҒ0a�l1� ��vº��r1o����]T�ɨ6��P��E�r�7�l�"2x�_��)��)H��k�[�H��DP�}�QagUj���.�O_�}�h��q��T'��.�S'�!�3�c���v,.(��'ȕQ<Q<0i팈s�o2.~�D������6ռ�sL����ǖ��u#�b0�{�R���0�2�I���dnE]�T@O�t&
�Nt�.C�Q �b���ea�U�-�L<L���������9�-Xs�)���55��^F���C���hA@��G�`�*��m�Fw�Xi�%�]�$�z	��.��3��j/�����D�y*��ŞBG��۩���B3�Y�ژ�[�l<��<e'�R#A� ?'R�NN�;��lN���EOL�rxMT�d�(�WX��!�F��+>��� �j&�5�2����y*�����{��IԒ2�)RЯ}�FW״���t�o�d1M�b)-A�����y���9b>����7�JOu�{kyW�.M���������F���]ˬ��{Q9Qެ�>�i�����?]��-����W'[�t�с2�q�����R
��y�l�L{�x��2''@� ��`q�Tt�_�<��ვϟ��(Č��ۯeW(�N�}�4;鍮��RE�>$��^�~��;[��B�K�TBX��X
���H��rba��܎��x�
�o��b{�b�<Q0�V�>��Z�*�Xs)�>!
�_[$i�B�n�����z�ۄ\��^!���6����J�7�@�}�nR�l
ń��g"~l ��1�x!	��:��)T�_�]=~ߧ�PKE~h�	� ����^�[-��-�ղuG94�����0�y��)�)����!|H�5��u���8JM�U��p|;�~{iN*�t5@�Z�װ�v�"\������2tA��V��?h>t�T�Qd�^Y��V�E�=J���:�ﾖ���-ޖL�Om�RE����n�B�	�X7�����rN՘.R���Q��	��hYkJ�N�t,6����(�=Շ��\e}�Fx,wd�S:y��0k5���G��-��b�3���������+,�A]��� �g�����K'�!�B�q�� O��_��F>�U�ˬ���v�(~~�ck0.ӀQ�
x-@?m�7 %ϒ�_��)�#�k]N��!�Ua��v8��F��͝sasPA�[)iA��G���MQQ��X���@�N0P���f1�ÊC�,�S,��WP`w!;�a��v7��|L[�VI(Ԯ��5�n
|Ӟ-�ڦ.���U��L����P����㋌1K���Y�%��x�����|�"0�� �ʧy�I� E�AoMV2��� ȽZZ����-��� W��� �de�l�:a�ϝD��*��u�7�Pj��d���!�h�������r^H/^�@$mh��C ���
�h�y�U���NCVe��LA!V�?�,���.����y7��{>{��)�� ��R+��反7���胭����{�GGǭB�Mδ�Г�Uʋ�G4j%1��eG��<��Or`�k#P��Tg�ZfI�e~�<�6x4�G�i�.p�JBn`hD�s���=~��,ȧՄ��=rxO���[�����T�'d�Vj[�BF���$��Lq��x�x���7��4as�p51CB� �RO�^NlGIf"ZP9t���ɲs�����vM�!P,_zb��0�e���Xb�����)s/��e�ݎGݥ�#l��Ťk����n�|`A�ʸ�AYJ�{Ţ=z��d��A�|1��:6Y&�-j��<4c�7L�(G�>\ugtk*�,*܃ZJ�U�L-/[��L�Qܱ�B�	z@�v�P�X���7�h%�O������"�)`Ф��'�$ؘ��Xl�t��������d-	��icP�ͫȟA�-��/����2��(�B��-�R��F5:Z��&h��8����;%�U,P�S#�{/�r�[p�ɍ��eŲG�ׂ�|J�	��^*W�&�n�H�H�ד�nirVa�`V֟����N��DH$'(~�������� F����������d��!éǮx�lPv��r0[e���d��V�mr��ՂP(LL�2�wMX&�B�&��d�!&� ���:
<!�"�lB4�N��T�Ν��G������eO��O�i��|>��5���~��F��Y��Ik�ħDr�PSq4:
��)�$�P(���Q#Mh��1$rmb�C�=�hc�}�K�(�P�4����O��t���-ܹ�k�F�\[���8�~��������:���C�%}�?�R]_�Dwr��w$"$�1�3�Iʎ����k��U��$n&���W@&�J�Au{v h�!F$'ֳ�90��Ŧ�m6/.m��4�Lr�wY��7�ٲ����O0(�֢����_IN���P��-�yC�ё��Mv�^�_qurOӒ���`m�_Qq(eʟ��x�z��盅�h
m�ӡG�ɛW8&��P��5�-%�k����s۬�R*&��^w� �� C$!�U(F����_���+��'���4��,�PLB�iN��jJ��%StBQO��Ɂ�'�&<�����'��$����
����f^�Hx����`�%�M�M�3�8ѡX�
�W����yxS9� ���\�ȁ���v4����ʵA(�ܠ��ƼL���v��x63����(���Pe}��tv*CU*�n7�P��^|vl��)D�ˇ'�+�6|*�o��o~9}��ԏ�f��U��3�ـ	J���P/�|Y2�3�3�|�ŉy:�+$e~���d�n��R'��ƕ�u�
/)+V�Z��o�"��@!}�����>�3I�rҁk�]�}6���8���U{��/�or��l��Wm"(n:��L���v��V䄉��G�g� Y��C���v�Ɔ<bV��-�.��l�k�[I�C-;�;���'}�+F���l��)�_F���X���S�&��*�s��1
!��M�O����%��1� ������uRU���U�q�ݠ���e	�b����;51����{}&G"����`SGb7��[9ҵ��O����/�P&���o��8� �~G` �Kk���,��L��0f�Sc���3(	�˗v��)TS�D8dib�BXiS�0l鿑�j��J�4P��뷲�U�����P�����/g�q2Ů4�u��I'y�Fhm:�j�ŉ���H����˄���^���6z;���]MV�(�� !	���1�L-����\�a�J&qz-,~)�sv����E���Q/����5�>���S5�dZL>m�d`�Ï:ƛI{n����c�Hh󇭌f�F���(\n*p$�zl������'9�Ø�C�L���z���>���BTK@���V��	�Bw�DH6.x���L�i��8!��9<�#��ghv�'�M���΃Wo ���3y�}��j)*GxX�!M/��%�fW�5������]�t
�� Rv����U�ᮉ� �yj�%����_m��9�0d�HCtV��U�"z��-�/Y&��g�&���X��WK�ւ?�l?�,=V�h�J>0"����}�Fv����yYz�#� u�+�-��'���6w�^*I��mW��b����åw�QyA ��f��'�h~8�G���CY�U�`]�D�g,?)�cl�E��i3!��9����\��_.@
sM��t��-*VA'܆�kԎ��`Pٲ��M�/�}�dQe's�8ˆEa=5�P�m�O٪�`=��q�JM��q��{:P�g�G�ɫh�����0��� ���h'�'p�d�n�qo�E���{�wl�"���Ú��:�q.���Fš���˄�B�ˈ��n��*��BqHW2�����K���TQ���{Q-2Wڴ��������NZ��N�;��v	�?4D�P4G��&�RLw�L���ul�Z��VƗ�wQ�g
��xb�S���51�`�6~�X�ik����@
���PS��馥��WC�4���q��0ػ%	��9?_BX�'��ֹ�r˗��-��le����x��7=d_Ou��pM�f^�{�G�����h7m�4[�1��䠧A"<�I|ܭ�.��Q��xE���!.0P�^�0�W�Bp���H^�7��袂t�|�?�^
"��`~)�/u3��I0��NCz�U�u0�ى"MD�vUj*�J�k��� {]kL��
qW�u�2څ3x<,�b5�&8ʱJ� �pU/�Z���D$��+V;I_h��[1���}]�U4�?��w=J���ǐ��AL�y6���͵����2�2�1�W$����w���-�q���w����#�����-��@����j?3�9���Q��d��9lX��Y��� ��&��7�#KѬ�8z��˞OOelu4;������l_� du�G+F~%44OzW�[:-��ndN�J�3(EE�B/�ɯHnuX�wO
 �-\�_.[��eҜt2��-���9���ޤ��y����n��MI+�`��2G���n������-�����U�H�p�D��	��(����\/��][�Ş�P��6(ۊ���M�2��ٿp7�r���4�~�I�&o��������9�>�F�k��1X���R/��|��	�"��z�zS��=e���U�b��J/�_+��@1αVMȆV�8���%M����u��P��w���_���	�>�1�(D����cE;�p2�^I`�9�8�
[��ba
�
ߟ�fJ3©!���U�=W�]���L�#�@��%x%�ܭY��	�|�	��^�vw�@�g���c:lߢ����tZ�2�'���r��S^�nӍ����� 7�{c�H���,��|�+�x�:�		 �ؾEl*���k��=ظÕ��t5iϘ�j�!D�#30(�����ݰ�%���κ�yd�9A�X5��S�T�؁�at}�(�p:��헪���M��79�]zVh7*�P@�k���~����Z6K���)e�Q���I���!_�۔�b�?��\[���$�v�/�6� �o �i�g���p`\���#��!�tPX����e[W��ch޽��^BC�3���N>�1��ph]�?�?��;_��MFi�O^���d�!���\�u�7粣x�י�c �]�q.@3��KE��q��;-�6�2�҉�����ά]�����G��P��Ws�b.^��L��,)��ܦ� !��W���9#-�b�O+�̱����%;ȝ�v�;�y��'��a�y�捍u6��)�Z����	 �l���ն���gW�쨘X�|��w1(jR]dc�A���W��U����Y�#P�NJO@m[m�t��ڰ����ȼS�Ӱ�ͪ�/�k��P{k���vA�0Ƀ�T�����2(y|�u��I�<��\u�1�c�e9�n�}6�{�QEd���tdd{��g��ДG��K�,<�C�M��pY�{a�	��Yk`<��LX��Zv-�Sؒ�����&��5*fZ朝�
�I2j�:Q�=�	����z �I������vþ�5��vIˇ�T��B�����4fM��?���Q�5�F�(��Uo=<rB�ΰ�]��'o�����f��{���sB��,S���l�-Ʉ���v�׍��k����
�&۟�{����^�i�J��&�XN@t� �&�u)�½M�W�v����̌sP��v=�:����蹄�a�7��:$�UP\��P,W>��L���߶­�|�wC*���N/t�f�`�X�9r�0n("1t�KHy�ڥG%Z,���H&��৬�<~`�.��������z��0K��*�d��}n��$ j;q����_�!�	)j�);G.c��0�r��j�uc�a��S̥y�k��UL1��4x�_����łW\O��b��ē�]V�p$?o3�	�d6�Y��0��j�H}3cT�5p�t]���l����}����=��N[��f�-�|�qç<Z���=�D�:�Iр���30ќ6N`f��\g�����:'q��&���~O���U��01Q�_i�+�0`�,F0r2w�X=* ���N9~e�C���@��/E5.D���f�ʒ����f�T�I��QQQN��D��=C���#T�ec0{�^A^D���%S"�^��JK\������qx�uL��`��|��.|�u���.�����Kw��ľ1�O�Gǽ�E/�v���K<���S�.��z֏!�� �Q�(؏��#���T�׼��Q�����0d�V�x�w�O�<ظ�d����2�P�f�b����kѦ���V���g룒�:%Ӳ���dp���T�Zn�'���T��7;'Hࢢ��%��(X��vG����J>�n�:�u��_�v�c�t���صL2��-��\�������&�ji��f�Ls��VD�nW�C�͚�ņ��������v�у)�^�*m�t�m�� �	a���/�h$I;mB�u���J	��C}P䢫F�*�<I*q�Kn�y�[&�����\j�YC��U������3
l���p=��;ҡv�����G���x#Ue&�m���&�c�=߈�V�^5��٠�\}ݮ�[t���ό�u����y����
�i�پ]��D ރg�c�1�a�D@4=��Ɉ�i�(�M�vr؇��#5�<[�'ê���S@�0����(d�ܸ��
��ɹa-Z�L�Լ���h6��s^���M�An ��s2��O�%���k>�7J���[D�]\�N���R�0�3��B@� 1�|��Rodo_Ώ����0A�� �у֦*� ��؁D�X�_�4U�cY`#\�e8�%E�{��3&#�*&x&��B���~�(~�?�G�KJ?�O��qY�C�8g�r���JNBr�-0����b��;�����1�@9RV�;)��+���C*��o��1G�J������|ǽ�f[i�}��¯տ�k�����xHݡ�5�{G$�_�f��pd�1MHp/�_�</l�r�G
��u�����$i��v��mV�C�HYr�5=t'�(�KW�*Һ��N�H�0�0z�g,�#��*o�a)랤H����(fh���3��w�V�72�.��q¸��9#�Ec��NO������p�$>C�̥0	��mR�{��V�q�����i��'�^~k�Lyd���kul�,_ж��{��CSg�G<��H�Ur��/�mM�R�G�Z�>�w5�@��k07 �M�3�4���\#\�a�����x�1%<Ew#����;1/�qO�m�"z�t��5���[�z��\r&��M�}5�塞|(=*����e�lq;�k�/�K��CU�	p���� U���|���C����Y"�i9�|`�)`cb(�%���W�^
�!��C4߹�b��	�N��q�!�A~$��=cjeѩ-�g!/"��ͽ�v�]-o~f^��n�΄L��[�DP|-$��9��̛q�Kf������jpwU�LG��Lg&��,2�^!��X��R�^�*�����>Q�DH�����c`N~9X�B�vg�T�IU�˃V�S����Cl�m�v���,�k?��3}y��֘���۹�#���\'AW�+Hw�zW�c��G����D���֗��_�4ޝ��,;K�?,���P]��N���/�}م0���>�I��k��m��ȴ,"��,�%"��lj?W3�Ϙ��%k��2��ݾ���R{��I��,a��Z��hV2E�5Zo�	��*�-�4�w�DU*e���BY����u)6�1I��@or�.�B*R4Yĳ�J�ϖ�(���vu��Tެ*��>��:��r*���}5DѪ�4��\u!��I
�݈��ǯ� ��?�qJy�yŝóR���R�C�A=���4�8��m�mhFP�Q+��y
�;#�É���-���ZR6�{�po��K��A'�'�r�y�4��qF��+i��tE��U�vڍ�)¦�J�,Օ,�>���a(��:z�-Y�E���R��~��0l�Ƙ�$
����i�(ұ�A�Ҵ'A|�{�ab�����(Y����q_h��̊�철T�q̻�����G�)��JX���K�h���B�x�ݝ��(o��eZ��Q*z�"�E�Y'v��ݪn.���U͑�.�x���B���i��y��x;Z��Uh�SY�����{=����#a �1��9m)t+��v1[-m6p;����"�]4 ����#N�C^�5��yN��J𸸸�Q�@�r W³9F_��p���?��NQ���Ӂ<��`��-m�k�[w-&T.�Pظ����3TҠ���k�X��w]bÁcю�x�0e7�t�XNбC˹�k|�ir�A�0Т�Y��`Ky��y��8
[�c�ئ�ZT|�f0�?�p C
�a�����^e�ȧr=5���&����%Y?	�e�\|��`n��q�y�=�=��.�����$؍A`��f@3ġ�E�H���V�y�0�6gpqm�R��scT�|�|��W����BѸ�I0�&ˑ���¬��?k��Y'uvgjF��,O��h�o��I��@�ٽt��p���(�aI�;�ۋ��e��ㅡ2R<~�c|�Y����\���3|]�#q㧮f�B���{i;C-�b�GB�#�s����oӶ�x������4�zM��y�GA�Ĕ�*ġV�\�����F�/���moZaA���C�5V녉���뗪�4�oNr�5�܄����Dw�j	���oX�.���ɵ .w��B�Ar:���n��,k�v������֫Rw�E4�̴j����,rVUס��pf�����DC?��#([�)5��1q��W[��*Ս0㶫 >� n�	Rz�t���I�a�l��5!T��Uo	2�%�+�%|�%�!ql�x���u��=U���d���vջ ���_%"�^	��+5'�q�b�{t�ˌ�}D ~�ԣ�����6�s��5��l��!�� {�1�{�z��������B�4B����T�ހ� �H�B��G��-�i{�=��G�$f
oR���j$��G�jEr�i��ȃoJ�����pe�#$�5P[.-�K�(�x"�ff��HA�g�vM�7H�5��bm��7��s���u�"�\~�a4yf��2وL����gf�3�?��߄bs�
��|�����g~�+�k�������vQ&���$�Ol3�H+Nvi��3�x�4W3�25$�ܫ�r��W�#w�z����K�l���j�m'r�i!1?��K\{Eo�$mfB�ؿ��H+7��<���j�JN+�P���/��[<Tô���qS�v/?V�z��n�`e�AS\��'���C�&�B��)�D�����뇩�6��$��ڀ�7�����~�cZ�b�˟�;X���g��b=�
}ˇ�5�h")��<��W��	�9 t�V�閡����p���� ���ݯH[
�T<�/�~�1rU	��DF���=�&���\�9ZG|w�P"q+�_�K+0Z3��p�3�#f�� ad:�E������?��6��gl@vHwP|�;uC܁*�U����>�oT��MW��-��0�S�^p�;��m!&��8V����J�2��4����
�����d�#b�m�����Iu�!m)VH�K���88���y0d?���]^R�u��gb�@q�ބd;���g�����.�T�_r;�h:Q���� !p@B�@��)���ԡ���I9 H^��x�.L�&V������M�2�@
�9ߍ�3-9�@�>3E!�2]�E,����-��%1NZ�K4r��z��؉���~l�b����<�)�ś�,V꫄�_�`�a>��@=��"w���l��O�j3�gڏ=�c56ъnrq��!"� ����EF��3����o1�Bf����i��QzVzii&NEi"�_NMT�\�~c�a�f`m���;�f�T�uJ�izn�kȹ���a�%�)�A�[S7z�
4����9� (b��8J�`�f�_W�nӇ�!�'���D�I�0��lݎ{�f9�+r�{��B��r˺p�Yā�~��x��L�,|}9z!*�8JI������^ػޯN`h�)@��R��/�+�T&�uγ8��C�K�����c?������_�#�d���zd�&A��Ji$\�K?�7��߹s�׻��BtDzҙ������k��`��X��w�W�w;\ޟ��RD���B���79�&6d�!���C���;��Ӱ�و�w��](v}�1D��ťʮ�w�)����%�����'G{����lbN�Xܻڣb�u��Ͷ�-[	��x��X�7�}(
3��B���[�'^��:�d�P��VtO�ɬ{�m*͌Ƭ]�"Ek�>x@
a�G��uS�=�뭈��M=@i���2d-meyTle��*���5��˶x��[!���]�ċN ��z���_wv^�C��c�0���
�Z�'��ފ�Z���`��t�3�˵)5�sX���@�4��Qp��g׸w�}]��Ԕ6�ޠ^��5���[6�Y%z4����t!ġ��Z����gOtO0�ԏ��t�����3�"|`�!���}$T@4x��Ò��YڹL{�Qu�Z��6n�O疼�f�ZZvd�YpKٹqX�4�=����0$�gDx�W���9}6j��u��.�xI@��`�!
ڕ�%Q�xr��#É'��P��"Ym�j���;UZ���|A�u��sA׵^e�����%�f	M~9����K4��0�$�N�W�S��'�����gM�D�!s�\���h�՗Թ2�s`"I�s}����xJ��r�-��O�o��w���q	�6�Lc�bϕ!웃8�ºS�W�,�!�G���fw��%��lSB;�01�+E=�33���I{��������(5Ȑ�O��t?�!��/��T��j~�[1+yC�D�aK��v��G�A��ru�Zݑ���a Z��o׳�)ʟBA�]�ܒ�h���m�\��K7��=��)L��"�j��>K����z'����2*��؏I�a���Rz��ƭ�S�̹��y����g� ��]JY�ߊO,�C2�m�b��&𩢬�W܄����.A5�/�L������v�v˪r�nw=8俲?ʎ���*�+A�r���<�غ;�ͿW/.�˴EN�ꑐ1���-5��+5t?T�cQ��� )>M�K��~X6����3?�=yT�m5�`�W�϶d@K'��%��!������Խ������S�9�� ��l�����g��j	��}#)E��B����\�r��:�CU�D�+B�1�9�:CGx0n0�%��2[�T_o�%Ę¡tR�Q�F�M�AǮF�L ����^*?D���p�V��B�Qk�� \��!�5x���QLZw���?��u��R��l�$���Gƃu�'(y���D��dE\��/9�������n6=;5=~(�����`P��N*�o��h�4ЉCH��9h,��~�U�i:}fX��~�"Z�,�f��F�Q��@^8ݍ3L�ʱ��������7ێ̯��m��;	�J��;^}̉���P�G{$ ;�L)0H����E�P���iΙ(k�2�.�&t��b�^�J�������b���b�eߵS��P������T�KP��Y���Q�����R��G�fb���h��U֡��Yw��_q�l�Š)Vˬ1�1�y�W��%�플3:��k�|���&����,�r�3ant���+ڮ����a$�#�=kA����u8hχ�J��Ĩ`�v!%B]l���)�Ď�k&0yjqƃx{�݀E��\�v�؄��d��׸8!�7X��Y]#����	:K�\�@��o	XB���&�&��e��}�s��>�֗��4��ĳ���G{瀂u�M�r��t��cZ�,R�JN��Y
�)K���а:����j�$��g�&+l�)���l�����>/t{P�Sq�sy%�5��H���u��:�BЀ�t}\҅Y9`@~�E]�'^�/�@BB���?�މ4������p����9���y�9\~擺�Ȉ��)Vr������iO�b_�G����a�S�'�t��@wG"�!D(�E�E6�3h�%�X�a���c���H�ɜ<�&���?ã}�`�~k� �F��4\�̕�O��M�=QK?f��e ����>sq-,&�SRz�"���F4W�N�[$v~g.CR� H�� xZ�!R�o��>���	A4���Ц|o�����(���<W��IMz-��OL�Syza�����p�����҇T�;��&1�z��G,4�G-��/�W�6�����g�5C�J�o;UN�f���2s���A]}���wu���c,�t=]e>���${��V~��.i��ңؕ� Da-S���I�l׼��T"�	d���lY��<����&F���v��=�
�+I� ��ӱ=�s���`�oz��� ��M}ԫA�y@�M��	����H��@J�ѐi]��Z���+����gQYj��U~/TRp8�sr/��(�Xٻ2�F�+`6����l/,Y0Z_p�Ȭ �c�UUg6C����}�P* ���}H�*���K<���=���0&s'�������}��c"��q���n  �. "s��X\� �^�1��ۘT�%8�ET�^�L'e��$ub73��d�Ż� ��A��y�G�Wz^��vDd�&����ވ_� )�,ѾǷ
�Uq9�,�@�=��hg��6��RKU-ω��v�������t�b�_��9^�b�5�Y��9�φ���ǅYq�Bl�ެ<ݕX���� b=���$<��{@��4�EE��6z��`��S�u�p���-�]�$u擻ӫ(�q���ůq�� �� � �i�~U%	s��,����|���,�P�E����|]XX �?�l?y.(R��}�%��N�5J<�A^����i�E���$�#�!���W�����z1��̳�q�hH�V�����"g��rJN��)��/���g�[�e;4�aj%\k�
�`&]�x�!���5V2o���R����B-�HJ�&�ؑ�Vۅѹ�DK�K���LLv>��ƍ��Mw��q��xz����n����c� �/T�MW��]7t���o�n}��B�����ϿС�ur�㧙ꝔSbj���m��A�����O��L��ܡ'��5�:�
�������V�j|�����#����/���{����h,�*s�T�b?j,h|����C�����k�e����c��3wk>� ��9e���k��Dx�f�G��L؁�� T���3I�v��}ס�~�%�@[6��p�D~��ƕ�m�&��uíR����b���g��������O�pzz-�þ�� 7c\�^��RK:	�qL�be��<�-∕���'_�`9��<�o�]�A'F�麺� a�ܬ����*`O1E(��C޷�­�jo؎�DHБ��	W�g���)���X� �%��iQC�[Ɠ�pա�s��;�`�)O��n��_ɺ��xeZ^3|�h�(�_��,�0����������;ic��I��?�*\�/��u���L�����
�f΀�T����r�!.�)9f@i�`�>h�ٖ8�X�)���� �VD���O�T�1��x-�w��~�HR���-�n=�*w�Ě�.�٧����:�QO�Ɯ=�<ĒJAA��p�h�b��t��B�~;s-�3U߯x8SR \I?KG�F�-i�$�]��d����\�^Q&�~�Ϳ�L�T�B��&����8�����=s�e�Q�`�Y��;���K7|L�{N�-��۳�G��pGy�����KϢ{$��R3S�ݳ�ٞ#�q0�ծZ
�,��"�Ɲ�t����%tP�����+y*%du'�skC����m��g>�%]k嫱���̭��4XB�v�۵#��X�vKPE P�D����E�����+�;$gu\`R����vB\�=��!yl�<� �7�N�r�;8���D%��O������������B=�M�x���B�6�O�4L�/����ߟs�Z��ӎ�?�'��s�w9?z�7f"��Ӱa�K{,��𵀣kq@��<>��ڪ+^{��$q��pr�VӂJ�q�BP�� Ф�=x��^�mbM�(��wJ���9�m,{��fʐu���ʜ�Kb4�Lw9,����@9��⵭M�A�.��fN��0 M��C�q�ϳeg��.0�w_��_�7b]B)����zY�u�D����Z2�C��2�6�e���ܼ���%.t��Q��'y9W�z��
�Kob��='�e:'6D󤒐{�Ǜ�N3���+Иٖo1W��#�����DAvae=%(7���_����kGx;���u�䚕1�Ҭh��5��$���M`?'�X�ƽ�΢~��!W[]��ek�^�
�Ax�H����:Z�`�W��U�K�H�lVXo"I>XG "��lP��v�y��r�F=[�����P$s��`��&{sij<�(�%���c����=�V�����\J5�ܞ&�T�h~?�ͮ��Ԉ�y���$RK�j�Ǣ�70�H�9�+����ޫ#8����X����|��=|,IJ�H��*�U�P�rIf�t2K�-�ỵ>S��I�q@��խ�y�Ӕt���&ne����f�Ju��r�Ũ��9s��m؛�+⢵j��r�IO�� bQ�?;5��[_V�ʥ<~
��|s��*7���2R��-�G4������E�L��L��`1^�9�S?b+�,�펿M�gE���r`Î��a�'%dq���U�f�|U?7�g2mRJ�q���H��g�C�RK�`��ݞ8��:ņ:Xq�x�����xM�>/=P�a����?W�!��x��G�k/�^%��)� �f������MZ�z|�}����l%W����/�24����	�Ak�%$xw��|��S>P�o��a�T�P�r6�!p�{wW!����0��&F�0"���F�jDA�~0'��`�CBz�/�&�6,�^�3��ӑ������Ȃ|BC���O���\u��*f��c��
co��%1�3���v��#ɞK���BPF���I�Ó'D���j�,�PNJP[�.�馘�k2��tv��<�IM.Pd�h�һ��x����'q?��_[�����^b���p��)&X�a��Ee�n�9�Un+5��s	3��l�K�$g�[�څ;�:D�(SM5-%�/�*E;��;Wg'x��0l�|M�/~wo�w � �N�����p;����~g|�:)�c!o��Cxo�-�W3�:D,��3NQ=D4f�,�()�$gh���Q��ԓ��$o��A>9{��W}��)!��\��3���}�N�ŴeI���a����m
�4ѧqv$xu�d�sF��)**�����~2��ͧ��9_�lBT�x��V�/�qK�9��b�5,�z�G�m�[t���Z���S�XP.����
H���4p)�iv�j.]g��0K]0�SZY���������筦1��E�w�7�Y�Y��4V�g��Y���u�$z�y�.1ص����(D�jW��ڞ���v?�S��0:FX2	n�_�\��Z7pa���ڪ�(vSU�o�Q)�f��i����O"�{
J����� ��x�+��+��X Uk�sE�&bJ���wl�4�(�����^��q��<J��Qx�J�tڔm�dK��(�B^�B�}pv�=�Ӝ0�e~T�I������9�W�Xf�X�5��G~������3$жH��t= ���ЪI����f]y���T�mh� z(=�d��� gPW�(�xD��e犣*8��2
�]WȢ��[��k��ͯq^�%��7�W��f��xgv�W�M�6�\3�\���p�$�"��f>�8�`]�H7�_)�"�V��k��>��Y]8�%���X2����C�Gt-K�s�h�"�"�է'�]��g־�ޤ����4��՜�ap����NJ;��V��V��d���7&�Q�5��;j��֡pG�`/Ә�קs#��=���2i?K����d�y /6�A�g���bl3w�7or�9����D6�����k���~0J�@���TוV�����P���3�����?��0裩����|.��y6�*��׽�͵�42N�"h`���Fs�m6vߡ���~6�I�k��c�^*�(*bS��@�/�uK�e�V ]���T���Kz���}*�և=t��7�㚀f�Xu����Sʺ2¿-h1j*��Rĥ�w�D|/� �!��&]Z�ê)��h����9]��t�&Ц�ۖuG,`$�=T�L��a�JkX��4�E���M�c
 N|�|S5��:��3�M6u&Q��!&<m�u���յ��ϥ3�K��Z�B���db"�+���s���3��F�z&�t7ӈ�@��|�b+����+LW*�F�jB2��X��5�S���c�	����!�Lb,8b-á��3��a&���!u���EI�f=�[�Mr���"�~Ʋ�o��B��a�H����#M�����%�p��T�39�^���(��i���~MTٞi3�k~��3��.b%��.�g������͐�k��|p[���Ә�Q�_��ZD���qO� \|�I�r#�Vy����['�v��}]�J'<5O���XKY��c��}"Γi����}��$8�Sc]�4��38B)R�����M�����<dpI��:���cy[�E'U������)��d���k��LT��Q�~0g��ݕk=K���@�W��WA~��)��Y�V��d�<���f�|� ��}9s��x#���W����Eg}A�d`�R�0��1�J;R����r=R	�e�ES��l��K~\�PNG�� x���#�h"�y�t�R=q*�\y�`�|������ֱ
2�"3�;&��l�8��gU�����i����+Ν,�N61�=�V_�*�jEC�z �ti1
��@��k�O�\3��}ǃ���l���M�ۮּ�b
��ߤ�:���g���ל��y�)R��hz��J��>���R�綻�@�Cjb��|�iyZ�a�\jS/�l=cX	F�K0���)yhu�
����b�^��ˇ��,�%�����������~*���)����h�&�!B��on'�-�#�<*(Qm�h�����䤀]�j��5:$��=�0�~\\p�ޥgq؜�3�W�
zۭ~,��W�S</�:�O�*h�>_\�L���N�����9������UB�1י�֡rP��1�	a_����M��{D�n�����2�h�r$�)+x?��(�ٶc=E�Z�)��Ӯeq��@��F�2+a�Q�W���E���%�'¯�Dtz��*6�y,8�(�;]� ����m���(��rKO��ig�?3�0�P!��0��̈́Ѐ�4����2g�����@D�ю���5�"6Z���iz�µ!i�?�d�)%�Sw�y��'}��DjU�#�.�� ה�
���
P狴�	������N�����	:Y2_@4�PCf��o
�L�&n� Ӧ�hM��6���ű�^���Œ���������8X?0������@n�+�͞�O��O�P�|�p% �t��G���'o��H��s�~�?a-�ͅPlg�#HU@\�S 44��z]��s��}�i=N�!����A�LE��J���R��}ҷ�O:�G�F�0�q���*ހ���'�3��?fLA{�U}���Q�\��q+۩��̠�fze�59��4]�S�	vIK�CB=Ŧw�(�j˵�sm��k���Z �f����1/Pi������k�TIћ�U0�g��v��ɑU
DC�"��A�[�a�ŵ�L&�!��~R0������_`t����OK�w�a1CO��w�Tɗr��	&vNQ4c�|��j̇�w��� �0���_X3h����2�MD�46����N^6�5�f$3(�Z���ǅ㧹f?C4鱱Qu"CI�p}Ա���DhP�H"��
2I|��fQi���{ؘa�ξ�(����5��&0����Ŕ�2dG|N Z����Wc)g�����G�ݖP\g���M��k@�\��E))�:���@D�h\�=iG���!tbu3�_�G�῱VM�����$����u�$g翂}�4:	�"�' 3�0�����H�pc2w�2;�
�Na��
�`r1��vՒ|_�3B�}�=A��<9����W�H�x�0М�=Q�N��'��R6��7o��~V��@���F�N-�H��o���Ƨ�S�+�Z���'����>*;!Z
���F���l�m3�*�(�^4�NL,}���$���R�8��0�	s�
��ZavU�4!f��#�a�s��V>sV�!�)���� �fN��J�2e�r�(Y�68��P}1#	�,����	�D)�M�A��X��=u_M�`� !RY8+���$����t��yI����DƽY��sY/�X�4ђ'����P/��t�W>c��V�6��4s��cڏy�b(���`f�I� ���EM8B�'���Q�`O��HX��Oo�d]P��;�Wy�I����Ɋ=�:\<�)�PC��oW�Y����ʡ���Q:�U3UH�����*�&4�#s/@�����~�r v��0�ƌ�b��8��`QV,��f�ȫj�����x��>��A������DkfJ;�]/F������N/χ7��1�vT����l��k5����'�u�Pfdnw���Q�s*@K�������zrt
�*�ÎrA�k�A��
�����r���.�z­pf澱z���@��)��K�Hʪ���o01�W���E�W�XD"��%(�{{�O3 �CZ���)�?�4��z"�Z��A���?�H�!�������-n-��ޝ(�7(���:1�8��(�Q��<�.��ܭiO��D��g@l$�v)�v���=1��l�5�c�L:�q���%K�sULh4�d��L(ۮ��ZS���E6�-��$괂���
βzo�$��S]H[1�	�ւ)�^�0,n��"o6#�V��8p&�D��7R�0f:ĉHԾXg��["V�D�ԣ-a�� �N>�P��Rtw��C�d�<�VY�����'��,*���M[?k �wJ`]i8�N��F�Y���s�T�]�F��H��[�p�O��R�)�� \��<F/��˹$��5h�u^�9�z|�0)ȅʈj�iߖ��Ԓ��ؠc����U���c�]/0
��[���(FI����|������E�on�'�9�`	e5t��a���	�X��� ������:ژ{��[JO����?Pm�,��5�b]�I�n09X����7��+���S��8[�w{D��~U�Ѓ9�׸,&�� ���0ɪU��JG�?)�%��ɘ�<�*�_�НA���4�Aq o��K�9ʟ>��w��aq�K�����:?j^H�*YpQ엿�|v�ʎQ��*v>�a��7"��<����O ��b�nJn������un'�M[��3��#i%���u-��t�)�}��>��LM�o�9�l_Ha�����A�F��5��ԩ��O�� �h�R8��4D�d��,�G���1��Q(�#���)�r%��ݔE`+�l���!��Oi�<LG�˱��`�{�|���~��ǞT'��:ޠ�|��& �,o	oV^�S��b�(c\� ���R/����Zo�a�����%%��־�:3�7�H�O���Ə��w�&���߷	��L6��(,���'�KbX���.ޣ�/�V=���
q�(�X�Jc�q4����)���?F�''��.7��܂�&�����ܥ�8MZ�������-)Q��⭍�\��4~�)����.�oJ���v݌a�]+�b�-Fe�Yg;���lW)��P˸����R��Ы\���w�u�����9�!�+J��&sAZ��Kk�_�����D�-�$wBS0`��������u��ܐ�)����0V3�Nh8�s������r+Uy�ٞ0D�Q(n�&����ɛ'��k����;7��O)�o�[��(.1�r3e#mZ��W$5 �	r�g�k�����kSX�5�p��'�{�+� ����
����V-�����b{�4�mHpB�vD=}u;�(��El��~2B��W��]b��7���##��Y��,'�n�Dk�וOn�E�:�i�\Gw�|~�ٶ��M{�+���ә���Z�H�i>�<���%%���I�=hNq�d.��iF0��bĽf���\%�%���)�_פ��Q)�-� z�kU뱅����v��t8µپ��נĬ�LP���Q��F+۾Ý��JA)���p3H���R��`ӛ� bLV��=�m2Kӽ[�d�^�%�I��x5�n�����?�[Xs&��a���!��ҜH�z�Z��PH��z{T���b�g�0��>��<���"T]]�`i�C!�Zd�	�PjgX�R�ϳ�@�֯0I`HX��Y�@��S��%2�z�Z���b����n$:��4gI���L�7�w9�L�!*�GԎ�?"��43?1H�+�v�a�$>�}N��$VJ��][���	x��E�G�;L��Ʀª
�3��h��S~26�tp���5���t��G`~��u����x�:  ��#P��.Z�O�ᚮh�v��L�LA\&�Z�hg����ɮ��@{�6�zϲ����o)$�~���XurЬ��
���&#k������'�Uy���s����[������o<�͂�4M\�y�nkεN)�X��V=��m���Z�����N�e^&�/Hՠ!"��~8���0<XZ�!:'\�_h���d� �v��~<k�Ɨ����oV�?�7�,�^/���r�,+�vY	�Q S��D`Ƈ6���8~�ss�!���N�>�_٩<��$��Gk����#)Ќ%��#oN-a*�ܲ������}|hy*�TQ�ߍ���H�5(�9V�,ԃ0`9��꿀d�A8�p�(]}��;��{&�{bIz�5^0X�f��yr}���#�����b�ވq<W.ǖ����g���r[+���Z�y�c7p�ڧ9p'W��zsF�l��:ڎ�l�o�����/U<wf��[ّ݋)}��ZN�n@���L�Q�-���Xj���fN6ϽE����Z�g����Tn�4�u�M"���{^,
m����a;�_,�.���OG7��U��c��Y�o-��
 �;I�c)��ҔD��Dd��f8��-��;c%�[��n��9D��I�h:�
�\߶_eI�Lk���,N[W2;��[������U��AX^hpNN)NZ�*'eÎ~�wQ_�x��J��+�+�!��q�[V����%��Ɋ$V1��|$����.[A�àlI�*ջ�Vxe��V�]b�b���@�}�Mh��z�S�������t�Ha��pS;�Ec�6���|>$�Z�<?��)�iʴ̶�iJ���!R�X��G��_-�ź���"��`�[����n�v6�}+��u�="����w��]��P���I�A���5�q�̏%��헝�ѐ��D���f%�=�2qw��tƞ �ݯ>�Q�� q 0�+��&����C��w�
�F��ㄘ����]%�*�7���[BxS��]�(�w��a��v����h���]���c
���H�*��&]	r�1���eM��o>����ڄ���U�i�I4�Y��%�Ae�Ro��ϻ8:��7���a7v�t��O����I�ؔ.�`޷l3���
�������ނ�|e.d�E7"����%��fw ��V5Wse��h���Ծ�1�o�-l��R}����*�ш��9���ߜ�X�5¿&T�b�._?)�1^~��Z��#�({ %��!�x�-��s�n�~����,��ݛ�R1U�Ux2��ݻcpsJ�e�f��A�l���=��#w��p�<�����ѯ~��>�C�yj�5?���x���ׄr+ߟX�@�W��N�0���I~��wKgPf[bHD����&���\W�}���]��a����YQ/�7�B6�X�A��/��<0.�z�U׮	�R��	�>i��4n�on�cv�f�"U�2HT�!A��&��Hg��7�/|�3��!e��R�Rԁ�C������<�����1�����V.EN�@�yqz�^g�LDn��]���'2M榦Z���>�冸�,|w:n\bA�����F�[�����m�ى�q����?p�l�-ÂVE����'H�����*9�������:����'��;dڹ�T�,^D��J���%�6�~>�J��L9^�xINu�Sa�s�-�)�]j����i�q�^�?9�4�r� ��� ��D{S8휖^��&X)�-
��A�ALD�sݮ�r���F�\f���������v.�ޘx�� �$�)�"pq��H�s<Y�$��*
�=�l0��Q���E0p��8��ݰ�3�mA��gF��C�ZV[�јu<8,��k�tΣw�����<r}���ɵ����S����X�:a���OK]���_#�{�2�(�Sxh4��`�7�x�JDG�>#��C��fW�}�U~�L�-_b�M�g}jq����h(d �2�����3�x�͌�����uH�H���7�;�Q�4�=��*����q����+hʜL������s%����g���%���d�܌��o��Pz*h�������3�.��ZLq���h��(��$�����u���#x�/c�iPOz�B�ls�����{��-/��w��r���x�ݽ����3������M��W1U�K����c�37��7-uJq�B�#7�7?\�ְ���1�X!t^݈�Q��{
��>��=B::$�6�֠�=�!qy��1q�ٵWS��<˦�{�C{;��囦 �!�y>�9��)|���}���t��;d����Oҝ� D1m���#��A�B'b�����;����Ї��ϭ�D�;5O��!�L�T:/�6N(�C�yBeZ���"�g��K��Y�i;%[����FƬP��y��B��c��Ɗ�恠���e;�7*.���[�eY��L��'�`aI�_�?����A�̹Y��t9��)�^a�{�ۦMC2�f�ƶP����s��q�&��e!��mF0�de�儘��l��,�
'B"��1D��$Q��)�A_߲��B�����V�WX����!��fa�^�ւ�,B�����kH%,��]��|,�58i�S���5���r`Ӹ&������y����1-�:�t7.�_��v��$�LPCo&�\����\��O5=+����>^~R�����;����*�揩���	��g�~-B�JAn焏0*��U-�}����q65u���z��a��&����b���9��K��9�9ca��W�i~��0���I�*�&`hjy��5 �o�b��Ylʶ�>�I���:��e����_�M~�̤�[v��B�6�L�7�E@��p��&6��;	�>�u�,���)��p����n<�<!mX���b�������߄}پ�|�����}��pe������Wֲ?��nU:m���^J����-$k��.]J	&U!��~�.<�#!G����;#[��#�<�0��n_�H@j�Y���h�0/��dז��Xݐټ����W�f�ꈸi\��B����IuT�v��n�2hW6�p�F�����ƻ2#zGW��k�R5��]f��N%�r�
½Q��Ro�Ƥz���I�+]c����Wj�7D�R��(
��;o��)��pIX��f���z՚��;~f=	�1�IѪ^�ϖ�Z�qܩ�[�N)R��}���a\ʦ�:�4�ȵ���~��
�Kf��/�R!u�8��ъ�p���nӑ �W6� Fd���O
�1{&ٔ�����K�NH�2O�}�����!}4:������U�Nk�D;˫���y�*����O��^0*��������7j6*�3Д�����k杲J�ʅ��86�	",�G0��/������nT�5�c�'XP�g㙺0��|��b���2�.Ul/^�����ՠ4V̂�_��Т��-�Sl~� J_:���F�_�Ud�zz���ӷ$����.��-��uRL�ڒ@��H@B}�zn��(����R�磹�U�����΍��\zG��?���$��y�m�.@��1�p�]�ii�Sh�'T�P�f�.���|���\gx-щ�i����X��JYB��wӅ�d	�����#epW�-����0�i�IC%���a���$3�/h;�P�Nt��`���8�+��%������nstK�k��LŇ��&X��@�>"��O�C���j=�!�}��jGWyfBag��;��%����B����A�O�1�-��:�ᛸ&����_�Ɯ:��`c�5	?M�C�Kke��iF�4]��\�^�/�o�͢v�9�H�,�R�.��c��tu���"EJ���F�Y�
)^�_�h�Ü�����al�Z�嶯�w^}���l���QOr�k
�v��
�i4�p�L��`>�����ͥ�ڬ?��UU�!��HЬA�@j0�?��~/Q�c�G����b���ua(��]�'�r!J^];föiU܋�YSd?\�?�7� l�a8����q�� ����p�"g|͛�"�U����V�$�3����L�
'"L<��u�"���6%�Wh��e$�F�)n�1��zZ3)�(;aH�͆�ӝG�V��߈'͛��x��ݛ��/J�?�_��֮�>��4��ۻ:~L�����:1z��?�i�L����VV����W�~���&���qXB�'-0Rt��y���V����dѳ^	�N�3�*N;|��i�m�7{�?<�R�To��̔A���{A��zI�7i
uKIr��'�;�$`�Ӆ�[ܟ�B�ff�.7�/bD�O�j�LgP8�Q���^��b���S�'�AkR�w�"�e�^��E}�9,:�ǳ)\Kp��~��t���l�b�Ή3#qvo��[$�S���K;EH�|�,l,��Ɲz��i�)�$��2�������%���%*܇��7V��*��	�Fg(*�X�Y?�/�:�����Jx8��2�<x���u�N�S+}ۯ�*\� ,w��"��zu@U}�.٘y��/z����ٮ�k�ǻ�%�����)��t]�Yh)J�,Äު�ǤD��������1!�{�=�Qî��^.��7�ѺI��_ģ�*~i�v{��}�V�u�������]��4��Қ�pV�]��>��*��~{ghȆ��4+YųA�w}���A9Z�����k<v�^��~�b�O�`,�U��&7g�3�~5/c4%�"f��a����X\��o+̲��^�A��\��f�Iᐵ�m/n��;HR�έ�T��/d�}�B����Gxo�wa9�َh���@��G�F��[�Փ�[h|�a{��y��!*v�B6�I�6k&����DgQ�Stu���hܻ�����(�����.瀅Ě�Y�}�niE���k��Q�Ř������OnY��W��|
�,8��k_byc�K�:�&�乏����^���}�&Uu+{��!2����^#08�h�r�[5"��,Au�Z)ШG������׮H�O������>l?qo���?����m�3�c���K�x��1��6�ֺ{gt<ʒV�x?����c�9)�e��lSP�יH���n8�k譋x|�q�Cvol)�!.�R�u�Ӌt�"da�I�R�=|CY�<��n(*Ss�����w�y������C��YF�ߏ!Y&�W�,�f������K*� �u����(���A'�O=8Ֆ$mڅ2���Y	v��Ȳ�$��ˇ<�v��.��pͤ���fS[�U�V�!�YH������������js�J����$�hnvRo�-/�:OĤ87VL�c��O�5�{J��hp��_��ق�]��K�J�xb��?S(���XN����X�Z2_��o�X�
J۴���䏄�;�%֙A��?2݈��B	���E�l{��=�21���4b�D���FY[|��!VI���^���I,2��&3Ա�q�Lm=��0�8�����08}6!3*v�V�D���ו2ρ#�`c��5���M��_%��e�N�M$��ǵZ@�-j�,��4�ϚnߠwYB�0�-ة)��6s��xv�{����$�:���l	����s)~xi):OHB��|h�[X���K�(�.A���jj�ΥB*��O$2�;�B%Q����4eb�ݏK6+���-2�|8�����Q�9�!�^u�f�#N�\�q������a)��%��u&�1��΁��iP^�k&h� ��m���+a v��I�+a0����s©�hy����+K��4.�e]�N���6��*�̠�iՃD�
e)�_�Z��5�qfW]`j�(`��ĴsB��L�-��3���}/V�Z3\v�A�_E��O�>�i���Y�/l�-t�I^�$8��H	DD���Ɔi5�
*�Ju�c>`��e)�a��EPP�]��8��ֆ�S��c����%3����n��[�I���9H�s�L@Eb�x�0Ս��rç����r�V�*:?���G�8;]@���b�}R�Wo�+�y�Y'�
ȿn���aq�y���%Y=2����o�	2F�����p8¯G����h�y�w��q���Rq]e�$+�c>fi|�r��@R���}��_h#a��F�9F�Kt6<P�4��l���ֺ+����Mv�Լ���3��9]��O��۾g�T�0��xu�t�=���t6�d�W���[jvi�?�d3�T0x0=��'4��>g�Z!�Rж9��{��1Ke�8�34��-��U�\�������D����b,��,�l�.XMu,}����6��d�h�$�'�dv��t�h�U�&�A�;3��b�7��N�?Vre(�@	�ot�r:���^V"g7p�� �~-2�5�W�u�	U�G��d����
:r���&�u[}�[lJ����� �hc�p�Ur�ē�D���� ]� ����ZzB���6�25�9�&�ЩH8��Nn�@�r�2��߅~-��늀�
D��"��Hh�tQ�v4��+�_�m�U��yf��Ƥkc����٩��_�3���.�Ȋ�|"��	 e#�j��jе��`�#�1�!&�l�q����J���CrZW[D9�j��roh-z+��w�]b�1�\��̔� JF�P�	�Kk��_R��� ��M"�z�q�&W��F�Y(�^.E$��NF���¨��l����w
vG��K��u�'@�ӛ֣�Ĉ�#�O�z��x��8p`��Pc�֗G�-�<*��E�ߨ^Ac�%�b0M�~Y�U���%�=��՜c�6�cop�HcD%xlf�I�
L���fL�>��>@�������X�Z:mš��d����nq�1�9���,da��_�|mL�1��G(�p�f����`����^���ٷa�U+���4#\�|&�H�#z0Y�O�ʶ�1Si%y�ϯy��Ut(3�ԣ�����R�p�wΓ���iEcs{f�����H���B�0�J��tIe+�b���&U��T�ωܟ?1��4�[�0����	�.���Ճ+���ΖKz'�5�د�V1L҃�����Ҭtx
��'w){A��a��pB	o{����=�&&�Ĵ�U����y���s�7�9�}���)�#h.���4��.��#*�f�W�!9)y�v���vt�C})�s����q�%)�+�����{{��J�!*��T�g-��z2���ʣ�H,f�D!�w�����U%�#<�3W/ɒZ�7��9V���K� �Jq���-b���s-��I4o�r�}@Ds����8[yoa
� ���<A �!J.d����:����	�>�)eM�`�C�}��k���~��20�K�OJ��]g���N�h��H�3q��X&aO.M�:��1�ѫXQ�#B��EQq�#E���o�lE�u��VS0�1�;�ݵ�c�>�5?p/ӱ�p$D���+KCG9)�R;V�����X�`��myS_�*�_z�	�h#�9B����4~Cҟ0�{���Ƣ��<m$�-K�����ê�����s�b)�����z��v9�c�ŕ��	�������m�k����|�h��u�#7:B�In�� �<�U���<�u#O���:�����f��n��ލ�p���^�nM�=u��Bs|]����;����['0Ć�(ޠo�fG�v��W�,MP=
�}M�!�M���;���AЊ�FB���o�y����&�ad�7��«�Y���'Iг��Q�]�A���""�:�q�ߌhx5��uN��7�����(O�j� e�����,DvW1���|�v����(<6��TH^G��G��/�[��C|��(ߟO6�EN�Y�$��Z|�憡vi�ʛ� �s6��#Ҁ���J
���
Fz"�^4��$�n��iym�]�t��ƂL��j�J.���sZ��>�%T��?�kw�w� V����n	C' � >;;�6;~~-��V�������UM\c��A	�_���!�I�"�ϒ�R�/= ��	:3��^��ڟ�?˝# C�y�E���8�ZV���T#SKcmd��Z�7�M�phέD����H+��%A�	ťVR��R~��~�%�o�+=��������g%na)��|U4C��8xh�RP`�i5����[��lС�
��d7��5�8��%�A%ꊧ��,�����v�i����u���lǘ��C�P�W��M�UE��A|^5ԙ�T��)�0�h�
�(�/��Y�i��F
Aj��w
$�a��1A�jє�Zf�"��Y>������al#�8J�hq�Cn�evJzIS�Zc�п8s�_-Ǜ˔�]��u��ܰ�S�"�{;�@i=4�aa�F舃���Z^y�pz�.7�^pS�+N��)�m��9Mw��Np
����`�ϲB�H����۳=��,`�^���3�Di(ʿ�R�h��Ռ�)�5$P����z�X�?�oO��Ҙ����c?C8�Y���������q�^��"����A��[qu������nnre�j6�۠������Kޣ��0�A����I��Ep��]y`��}���Ȑ���b{>� �0]*B�v_t5��[����)Փ��_!���j���Ä��2���#��Ͽ���� �%	��]�vQ��5��Cn��>���@�e��	XJ~�B}��ṱ!��)���f5��m�2då�I���ǚ#Ÿ.�	�o���Xod��5������R�[���e.����_������կ���g��-�&ҳ��[�o�`"q��b���mG���;/�����Q9jvMs�a���0���V�/W��������n}�� �/�}��[ڢ�I�ɣ��Ӽ�|�I#��.���]@[���w2�qU�"�s߂�����݊Ildfj_Zv�7�������/��J �8��`&�4�šX!a���wj~u\��l�U���a�_�Q|Ĺ�?R]b,;y��X��~;rxkw'�TzV�$D�4��EH���닜�&f�\�>G��,�Om܎���V�
�ǐs��߰���F��w}�@�N������t>Te�W�t}���S+:|q��3�N7��Q�2�G�7�X�4����!�qk�S&��8}�|����՞N�];B	�^�3il��,5���o���a��W_����7Ƒ��C8ڦ�?�| &_�6�.!����5T��nη�j��|������|8~��A��c3=
c�;C�̋:��g�x{0��f�Bb�Ev��3����wҜ5����{��Bf=#���ʝj�g<��>��b�'�����S/pn��I[���]�ۥj�8�����!�m�*/����xJ(�@��ń"X����UF���p���y��[t��8I^Պ��S�(1�6�_*�f$?τ���w��=P�����Y�q�`���r�5J����K����rI�� �Yq�A��b�|׮����]+��V�x�j��˯�0Ŀ���{�Ӕ	13��N��S�p7��Y��R%I���N��$�A1�5|CmT�T�˃y�lLt]�OTT~�Y��gV�$S4��,�|��2<g��X�U��`SP��1�k;}`m���C��NS�R���i�p17D�i��ʎ��#��tJ�RJ��Uk�"��'�i���?n)���i��3�#�d?ٴ;�b��3L�HܤtH}9��2������%��*6�z4^o"�T;��,e<v}0!��,��E�H��.�	3׸�ٚI�pW��<ţI!E}.�zp�궢v�����)�<����#�*�U&aCK��x1C
�4H�k�
%������R���0#�̩�@��u	�&>�h��A4��ó����]���$ b\S���,���?��'ҙY��G�'Yv<�7ހH�wk:�^��J�;�'�V�,K�b ���{��A����ax�~d��H|w��Ű�*vN�����m�'�r�$�3��x"`϶tZ���b��(���}��lO��������:���}.s�
��9.}�q�Rv����z2D��s�`��p[���Q���� ^�,l=�B9���o:�+!-��R���0j�c�s75����\=	���^;��fW7�Q��xn�T����A2�u�([巚]�d��#9!}�5�����yN���NJ�������'q��a�=�C6w+�A_��l��="џ��E��ٓYȀi'?�9��ٽ�.u{uI弶$�ʏ�pv�ɱ	���>S�$�S��O�?��&H�u�=��h�:�w����k�zS��	����������z,�
��o�xI������-�i��ѹ�6s��[�E�M�Bk�M���<��{F�Q3&��$�xF���� �������`�eI�y�50Ov���_��\�}���Y�bb�w�����j*8{rM�l�٧��a��w��ys���������P'���=(�������^�.T��mcۚn��j��okˣ(ac�%�`�E���1ű�84��L���~v���m�h�x���^%v�`��Te���ELݨ4ϲX�e`+��(L����S#yg�H�6Ʈ��a�w|.aq���?[ѣ=*��Y#^'_鞙�I����h�QW^)�����6�~�T��x�8ݥi�2s�W�y-�;H��r��i�	�J��}5IɝQpէܞH��.Sϫ�c��Y�J&n���4���Y�#v��h�1}�_����%��U���~��d�4w�n����Ӥ���sKY��j	��]3����:�+����&�m[;l9{F8���,���~L��U���\O�kF������(�a+eL���5U����m��9�+�*ʖf�0�
T���=��ڶs�ҁ����h�v�H������@���v﫭�s��3��0C$���C���Y�pj�����R��b�����J�Ʃ��g+��L˄S�,��M|�`�B|�M#�t�X�+D�akk�	9��8im�n���YGRۏeY�7�貍�[�Js�$�F���'A����L��ASBbRx���}lڡ�E��A��yT�F�M��o�FɥE�^kr�QI�@��m#�u����d�K��,?�*�m/E�@���_a�X2=F�Us	��m��z��uh�v��L�c��_�+��śC�헬p��t�ztu���)B秈�5k>�>m�b���R�"Ɓ��a���	%�h���S+�O��B��6����\�d��	�h��W]�н1zW��"��H%����(��1<W�,��K�������tΓU���r��T�ۛ�(���(.�*C��7��kx����acU:��}�"�7\kJ�P�d�|�Z��R���s�TLQ6s��ٕb�=���J�ިy��)����39�H����W�	Kg������@
�;@u�lz��J]*��Rrr*ȟu�#s�\�N=�{�i�9�i݁���WE4�5�'��靡�0�Ү�-_.�������|�L!������9�:�6S�p杹�ܨ�;�+P���qm�������#��8oظ�	�����8�1����a�0�c�P��6��Zh0(6R����4�㥘���|Hw]�����X�9��j������\ud`�sQ<)���9L���;��k�ܥ2q�$x��!�0�JP��4��7��4h�פO�����7��gj�0()=��3��[�0�w��i�o��{�H0,��1��
�5�rQd��iP�?��>~�-��i.���h�+����'M�kd7�������7�~�|�覂�Ð�)׾�{.{�� ������2�?>)��PJ�Fy�vU�ߖMy�rky�B^¿C��#�cmA�D�'ѱE#pO��8e�v�On��~���Z��<��B܆t����@�p�v�[���	>���s����i�C��(�XG3�+U ��=Z6�	��|�u2(^N���F����.qR|����$���!�&�8<?�:�CNg&$
)�O��@�Ȝ��W�Vҷ;����	p\n�i�P)���㇈"�H�uS����Z���y�.�)�dDn�'H�ѱGH�.��iO ![<���,�F[	e���Ɇ��Kl�bɖX�$�F_�y���PC�qޮ�;=�����@h�i�������ۣ��~ƈu�q<����?����v���l��V,/�Ld[7�\�n�|�mC�^���)��Bi�f+p��.
�1�A�4S������,΃i�|��)'�A�Q��n�#�5�T�j֫���:ۧG�-p�8�eel'�#eF#�]�8;.<�\.+��,l"�2�W�=S�-o�SٷNBжu7��4���yR�e�������)���6b��P�����kΈ-���c���OV�����ai3�-'w]Ї�s��qhRi���q��d5a�wȞ��p.�3&�n��^ hm����@w$ouL"�i�4d\�[�fw�[@��d�)`#v�|���} ��m�փ���fOK���	G"Q�am����+�O��ۏ`�`&O��,�[fX��92+�� �+a�Ѷ�����21��g�b�Z�L��;au8%iw��:�+�0��C6��u���0�Yl�����l2��.�d����N�6����!�i����3�p32�P��I�8��z2t�*���g���m�ݘ��[ZCYB�x~�]ޠc�G���oxVZR�,�hL��4w~Zq'Ǵ���[�=!:�+
��s����iȷ����g��8�f�x@B��N˛[bi���n��ީR&�N��, �����-��!�F�򝾥�20��Cd�5��8>Fɜ��������br��,��0D��@ ��[���(e��x�+�B	]��/��($����k��ɘ�B���ج�5Q�	Ͱ7鹆�c��f�?�FΨp�޸gF1W�\@~��C���Y��}V��Sz���F �j,��X� �� �� ?KBI�����>B֑B��IN��)�'�ٔ�;d�0�ʄ�I4z�D��g���\�Xj��[;�X�"�t��(�B��uf>���M�ٕ�\c�;2���o�l���Q_�΅��`������C�T1 tѱy*Ʉ�
��0�1VE�H%��晌K��]GX�Uq&�א��(_,�̥ ������;T@/W"$�Zl��f����i�����|W�4�y�2_3��:0)h]N2ř���ʲ���w��M� �AX2.�Fx"g)��nN\���wk*��F�^"<6ֵ�s��=NF|�S��;:�ӆ������#o�i�4X&@T@��MK>A�,z �L�Z��_�Z�Z��i����?��ȲL7�U.���P��X�A;6�E��/�J?���w�(q�	�ų���;S��!2�UF���ڼ��"�m����qgL��i�mc����ՃFJr��ˉ�%,�
q�t�1?�^��?>�UB���|_'M�Q��;��J�2��C֥:w�s�.?t��ڞ鸩e�=����J���o᥼�����S��H�ԪD�P2����E� ��>��Vf�|��yxI$�qD�+�3��;��DT�]D�\��
�����8}��#?;j�&;�xް�:����>��.����00�G�>[Cd����2����Q�@�ЍZ5�U*Bg����_�3�ٱ9���=���zÐ	�$����% O��g�H���B�y�}�j���5��\G��(��Z��>�m��,��&�06�k���y�;�,Mz�RL�Ś�la�fYG�؞��V`�\���wD��N_�%5 &L�1��
���4��b���laש����纴��1ب���ƎBҪz&���
�&'?�t�"?��ߨd�^�S�\G�=�	� ����ǉᘚ�O]I ���PP�0%�n���#����,
Ln?�_��!���c��}t��FA��OƲ�Ml?�G"+���=7o魄 p[N' ��9��bs[�� �����K���\�mi�S0FGѴ/�$�2ԍ�Io^i3����O≋p ��42��/��C��|<��ܭ�ʭ�Q:h��a�LR�kU7b�J�լ'�@�u�N�f�` �!��������������ԧ��J�Ƕ��J���~1v0��I��k^�q�G��h[�"?+m�imB����Y�lQ~�Rc��MK�7���
 ���&vq
 r>�W�����VrڡW���"�����c�EW������y��/J��+�7�Lr� �[Z"�+�Jl�c9|b�9'�1g��6�)T��5��e�vIp)��ns�#i6~�U0�l���7�R7+��aE�(�-aii�:�X��(�1U�����ף�?f��wki|K�02d�Z�נ#�E!���Z`��
;i8��h["����3��uK�+\�}h��ʖr��r���}�n��-O^�<�O���Q������QR	ΐT֬�[�\}�!��hOn6I�sx[ gҹ�ڱ��U��'}8�6�����ה�Srշc�����W
�k�M#l���Y�i��s^UB�m���_!Cd�5ع̅��<�wHT]U��[�-�M�Y��~Q� �E�j6�s���ިWxB[9�Ɛx:��6ñ^<Y�p@�+����[TB,j��$�RT�^�>��X�����śb��� �C�d�����}C: S1�IDh���jD`#��`L :��ů�5�1�+��^m�<�3�~�#F�|�?�W��1�+E�|j�s��#Ҭ��2l�mp�~Va������d6ȣd�c^4<�ݭ(4��)��E�p`<�"Z�D;�S;o��6s/z�p��=xh/�j	횊�W�nK�r���u�*��l���T��0iK䏉�j����+?��(�6�Q�t����T�޹'A�~����e�lV�-�jʐM�ᑑ����+�Vʖ���Ȑ�į<F�߽�D)�I��Ox6P����KO8j�nI(޾��F:�X��J��8�����f��YM�ݴ�ɉ*�v{�`"�Q|l=�k����O���\b��H;|7�LǱ�ם����aVrIܦ���qkUu����E�'��f�˫!Q��g�_�G�7ڠ�F{Xh�
��L�˒+�[QsH˓�hKn��ǒ�PΧ��D�2M�g�w?ʟ��,°��+(��v�Eg��x@�O.���ޫ���ǌ���m`����ڟ�w'��5�5�����įA��Q#ۜm"�$�>ȱV����6��f�^�UQ^�L]g6����ƠM6�2H����-���T��	��������]�=�X{��n_1ӄԁgv�D�\0�Ѐw>*S��݁��֗�l�EX*�mU���J���_lj@f��6!���)U`�j�"�/�%�Jr5ޢ�F�cb��l�E.��9C9(
����6#O�\~;�<d��R���V5�I��1�mԣ�2[�����1
u�]�}�bXC�	�f��E��\�,���~b$�ڈ��ѽq��g�~��[��	G��YO�d'X���j~�먽��������͵���h*+�W���}w��x����aM��W$x���W��!70�2�g�~�IY#��]/$v@<�N[�R`����lg=_HF���=�}Ǧ�$��T��r�����#���"@JȵĂ�s����0wXt�~�b,�8�lji��;�ߛuS�%�,�!X)�y�`�c�ps���@�Ò.��ܻ0r������~a��R{sS2O�O���� Y��* 2�������b^ْ�]�"�����g�س>�O8�YYm{h�t�Xts���V�I�IrfQ^���o�8ηzO���X}aT��M�\�pX����l9	�V���?H�����R�n��o���F��0X)����S+U�ڗ��g�0qO����q��������b�[x����Ӝ�!�fNC\���:��tb(�����x���Tc���\��v\@aj"Tt�,�+|���U@�][�ʇ�d�YÉ��	c�	$�œ^�����C]B�<�qB��6�Gj��-,M�q0�F3q���;?��㺫V��P��{<s�"�W��r����O,�corǹvc�ۼbJ�M�n��� �`Q�`擒p ������ҕ�9v��9l�q�*�ڴ���UNF
��i��j�Ui�,Z'_7_�I��?���w�"��cK���UE%�;*�t��'�p����+i'9� xIwI�yfԣ����n�߮x;��G'�$l������9���BV�Lm��꟤auޔU��
��s�K2�����$��F$�عq�"v}#��B�z�H�B=��c�*@�vU4
��UЪ���e��N=-�]���C-��&NV$��n�lC��ŮW����ߑk��L@�_��2
8�f�CH('x�w˒��F�l�Ӽ{bY�x���R�m7}&�r�X�J~^�5,�d�N������p�z�Օ�eS֛j�cr����dd����0�A躟S�^*�'k�O1�����iHL�����Mi{�����1[г�
�$�T>.����Ψh��p/���T�}:�2��#:��AN�����T�)0������<R���uWn��#'v�{g5Low��O�����QP�n
w6�X�,,�����m�څ����Nb 6"���O��\\_$eRWI�e���tzh`s����v-���hk�xn�,�%�O��?���Kno'*��/Ie�\8E�8�=�W�w����qy�N��b�$ho�����Jz�y�Z ���_��Cn�v�S��H�>���pB��'z�P�{��X��^W������g��k�B�<@��Q5ɂ?��EiR���s�t�T孜M,�`��?ǰ;��0k.� 9㶌��φ�@.�qe����g��+�C�y��܋��o��GWWN��
׏g[�p9`o½v�P�sM_�k��ðt#��+��1	��s��>����֑p"f��̸-Z���)7!�'a܋��0��a����ed� ��o����,�*��t��d�0ӮO�\�~_�ELΉ���,�Z��c>r�Ʌ~i@B�O���Y̫P�Q�Q�R�>����@.�ik`
�.�&ې� ��)�>�g��r�V�_��m����P�f�I =��J �[��*�qq���ɾ~�ߔ���F=X"�@�.���B�` v0qJ� �Xv��n���J�o[���SH��f$���;���N��.��i�+�i�[���\�ա>)6/�o�
A�F��2jt5~i��EB��{.Z�=�CKk�\y1�}L�b�H�d,}E�ľD�ϰ� e=�S���d�u�9)V˿�W�͛lo�}\B�܌��Y��V��,!�Qx?&��%�jgOr�?��;���p+�u2��I�s�>�M�4i�K�+_}[K#[��%]0�ht@�a��BQLgя�{�@	rִ�������_� �!�$t��s�����w���6�F9&ɦF��#X5W'�6�v<����D��ֺ�x��$����J��;��n#Qe��<{�K������'3�ODا��B^eN_�,\���:ˇ�Kd�5Y{��e/H�+��Ϭ���P�B�B�ޗyr�=l��a��Q	��N�2]�jf�AfB���������>B�e&��u}������s(_w��_�X�ytĮ��/x�B��`�[d���w<����י��d�M<�^�U�e��Ǆ����Ք�1!������*+�C,g4P�o�o/rg���W���H%P"	��j�ҟ������A�n<р)�������g�W+l�.�����hJ� ��큺�+��qy��=��r��� �t\��^��*����U��f���{r����sr/,�g�gt���b��8a�yLd��5���?�/�D �����BF]ґ�pj�A8�c>�KVث�Lh��v@��,�Rz@Rj�l��eA"����W(/ߥqF�<�I�.�#�� ����@�R�T`����k�e�bdY۶ʳ2���n�t/aҒ��./�.#�X~Z�?�r=@8!G�-���z.�Z��Q��mC�W��1Z��빒�����'ȿU���H����k�7���#�����me�1V���j�0�����f n�T�`��/���q�����M�fKPBs/�E0/}Ml�Ȳ_)}C)��u.T�� G	�b�C��g{��zf<��Pm֏L��s|>⻱���R�|�G���v[��ۺi�i1��|dԸЌ�Q��/�*J_U;�M�dL��t17!Q�r��Y[��o�o�z\a��oܿ"|�SblM~(�Z�������KZ;��=��Ek��;�N�[�8�O(��P��xi��K_�0���k�ia��iz��L^"0-����1�a�t��~:JPi��VTF33��?�/��һ�͋?≝>���R-.q�~��8���s�ͯ���]wS��A�6;��?0��,H0H0 �˕���i�G�{������T�k��ֱm|���t��/�<x��3%����5�E�D�SX�/$��i�D�u��_�~�h�lҖ���6���.}u.
���q�&"=w����m��>�b7Q�	7������t�L����d����(��'��_|������/�BF`HGñ�����
3�2�'{_TнE[���o:�� �ۄ���6�Yb�2��-.ߨ�,��Ҏ�ȑl* ���e®�HSk��{>X����g[<o�^~�#*��Fp��N[�&����T�b�#k��g	���y��<�����U�~�Βq�-�&!�������Ð��&�~T-�C,ԌM$#D��.ķc�JA�)�c�!��fꬾ������3��h���~,I�m��R��ŭ~�,A�P�A;��+c���ͺ��^���}��V� M�{���5z���#l}��`�*}�L⤻/GԼ�>�RI�������� ���|#r��	Q���l30����6&��	J��W ze �7Y�Ƅ�+�Y�n#n�ߟBjczq��Y ��i=Uf�2�E�����d�\��L����qА*�p�`Dٙ��c��`��bo�y(w��D� ��MM�b�gHn�^R3S	*"��6b`�N�eB�>!��бcp	�L�_��7���*pRi$�X��7��9E�[Eߺ���ʠ�g��#4y(&X�P�K,"�F���m���2\ܨ�T�-���^#�M
p*���xJ�HT�^O`��9�o���y1� t�[��\j�U�]9d?�*��?�ȍF��{9�8��f����<L�繉t֟@hrہeQ6����pW'u�ɢ;-�l��(i4�8�0��-K
*Q�"�L����J\~�@����A�A}����xW�IDa
�
i��m����I�2�y�r=�!C��N'�˄�I�]�x�eL4��g_���e����Z�Z4웺��Gn7���5�rX<os3��ދ ����ϬCyɦԈ�R	������j�.bi?(�p���1�Nu��G������[���0�*#O`��
ҤSNGW�� ŀ[<A�
���a\̘�dz�����0,�~� �f�F@F �}�3t410��/���:��O�.�cƆ���Y�ڹL���1�λ�PG
��{I��c��8��e4l��gޓN��5i��>3-ח�}ɹ��/N�����!R�1��ﴩ���be��M$����� ��☏��h��Ci�#�;{$ke�l\�;�])��;��ܜEg���xŴ��+�n,�?������׃J9 Q�2�[Ov��/�_�wy����v,�t���ij|C�7l������%g�e��7�k�1kY��<p�Z�Z;�M�JP����L:&�ZK�ָ*̬�R�0*�4�S��t��şx�%�}J�cU~""*3�߮�u���*�'5�~9�l�g��?"�*���K�����A×]�{r�g���F�o7���dXj�aC���DL��W��0��i�>��BK���=:�d���}�Wս����I쥽�+{� ��B	?�u��7%��-��x2�Ǹ4Ya��p@4�e�Osz9���|$|*�R �����^��t���SM�/FvZ�@[�U��+@�0x6����v!�c�y9]��vS�\`�ݟ���"ż����������>����Byh��獟��<����'�>��LG>����3�Ӡ�n
�n �J͞��K��:^Ӽ�>O�l8R�jp�<\1�,�-e�QoU��o`�������~�"���`�ғ�9Af��u��`ar/F=���w67�K��v����ʧqAлbLν1�Z�������ݎ�ٟ���#ev_�^�M�(�TIY�"��/��"P~�dtU�F6�,\>vao�Y9<�t[B �( l�c�c�$�_܁4�v��d|~?/�(���<�e��&$l����J��A�%#(��9��gC�j�W�,�/Z���[ŽF���&�*Z@A$�m"�X�D��Wݖ��j9e����B���8�k{f	�1ԣ��8�$�򖰳 alJ���/(�	�rIa��s��ڡ.�����T?�پ�y��d�q�n{�uA�`SC#"�HPT��
��-�"J@� �:���h�	se����:�v�_AQ�IS�hc<u��0�HVZ���c�Z�d��b�q�ˡ�J�X6P��-�?��vj ���#��Hԫ��f��?�L�]��C��,4�~��~�F*���D�ҏҦ؏d���|��fS�(��[�"���
U'���">vy�{,S�Kr����evR�흘z� E8g�^� ����o��/�q�.�T �A��l��k����Ty����G�N���aF$I�0�/o歬ذS����N�c��r����*E"�ׂ�G!�+Ú*��.~Nt��G(-v*�c�Gf�?�ZՌ/����Z8�g֢$��$����d�A��}��6̦�@у�7]Q��(5Zl�v�[�Ҭڣ��GTN�1�I؈!�`����1�
��a`�]�gŜ �����A������ ���B�1�,���B�3/�L*���pĪ��T$�L�e~���`Nc��Jkp��{ݮ��k�Q%�%ls$6��WmF����N[�pi���kx9�t����1� Զ�Fѝ��'.�� ��z#���n�@��br�ƉT��͐:dd�P�;�g�t��-1�0����ю7��+U,y%�i��	&�8�!Sj:1- y�4�%C�[S�Q��>N�B{��������k�zi"�<qx>V�2���t�eBts�֕}��lt���u�C(s�`+���k�=�vn�)�q�2�D��'n�:$s���۞�S�]�d�BZ�����6ӝ�jUSΉ���1��(>U��<���C�	j���Bn�c q�t��KzcU�"e��o7�i��f�-oĤ�����캽^��r�I��A!�LI�)�R��fY.�)-�H�X���ߗ��<�c}$�x_��1�����t¤K�ΛE�:}ԮD�;3ߪ$�v���G �f!Ye�~���?CT8��Df򧣌���a��xj2/�]� �368Q+��m���Py�7��q}��ŏ���)����t�S;�bCV�
����^
���w�\Wd��Ӳrl��7�Zt$�ޞ����(}�wM�b��8����,�Ҕ��w�_yp�(=�W���m��t|����<Z�<�j�۾�o�Z��[nRy��)Dڐ�Y��q\��6���؝����z;1?�~Li����u��3ɐFpSpᬁ�ɾ����~DF;���ݏ<� �aIf�xGg���C��7V�%(%�t��Yaՠ�1sޏ�	���i���9=AaݙB�%�M�� ���l��3/���}��v��%�ƥFq��Ӎ�A��H�C9&��Fܸ�������S �0/����������[�7��G����}9�T9*2�����&*Ţg�����G[���:�6;S�j��2��	a�����փ���8e��ʐX�˹3t8��XH�x�k���2��0�d1,�
h}�b�� `�POya=�{�����	�4>8˅Y�3��_lK�l_c��ޞ�9�i�Eh� NmX�Y�"�Dv�!�x#B�э��ː�ߘ�֞��(d\��}���*�{ q��)?��(�i����X�Ʉ���TZ�E����?��O4��,)s����T�✠��d8�*�Z�1�*�K��|��s�[� ��Ad�j�uZ�H������g�4
�R!�@1��pt��.��k��*p)e�M�|�n*d�i��U�	�y��&,����A	��{�R#;toG��B��*gz�����c���s�����m��ǅ�9P>!��G{���#��\�A���]��#9=��wk\��e�1��}����px���׃A�G~��ӑ��~�d��.*������['Z�B�To(ҹ(
zT޻E�V#I�[�E����	�[�e��JB��??�C�F�'j��4�@��[-u�������:�!no6=rW��jᦤEⵥ���9������Eժ��;���1�D(�ճ]p�b�Ju
D(�,�9����PL?�/���-��{�*ʕek���h~�N�̅��H�~��潁��o �?���������y-��~4�q'>�u�Q�t�L�N����֡�#H~�?�QS��q�I��3��f|j��ڇ$Lo5̔��\���]��0�o?b���?Zj�:1@w�PHW�1�q���6nX��=�1�JV���p`���m�K�ϼ��\D	p�DS`��	�P�t���r�r�[&Adw濧!�T۶��_Ӣ�an���at������g���wcRuse?gn?-`W�p�̈�����rΜ����@��~Be��1�R��h��[�\ﭏ�D.ڷ�� T9��k7�gG	i	i��kKv����l��3�EnWXt�-��cG����A�̈́I_��E�\���K�CG�Q�7Fe�m�W_߅���H`X!h�(�D������!W�"U��a� S�j�r��D�y�v]�FCu�u�*Q�
E��nyY���sD�|3Z�ZU���A+m�-vs��	���Y�������Jd���!s��/���1�ۛ)�2��u"�����5uإ�?�(����a��_E�����>��E����Cy�/�u�.X^f���q���t���7�"��37�d���Ԫ'Po2�2��LK*��O�E�r�����q:Ĕ9��V�u�1�1�kOlR�AX�@$���&�̷-��G���\7`�%g�]�-��U�ǚ6A:��Z��3d&�(�-��0��P䠪�YO�h ��LC�n�}l֚E��>�7�E�-�T/����K��������d��,���g\�TM����H��D��+��^9N񑣆jK-��2?���O1�Pz2�4�]���B|��:ʜv�����������S�ɄhN��H����^��^]��F��2�j�:��*n��ae(\t�	悞u�M� $�M�=�J�tXnW0�ݜ%������9�a��E~>{���c.E3������ڼ�cZ���^<��a������k� }:��۪�|��~KP�Cm�:H!νP��j�.]Aث4B�51���c��=�w���L�j�|/S��Pq��
�S1��6�A�Ͳ����XE	Q
�?�b׍.������-��,���X�/������?,lz�T���9�O[��9c��?>;�pi���#�v�i�,û'1�
xqq[�sIr���X;��>�u��ί8��{N��0z�Y\6�;��x�g�z�Ψj���c����N�������@w��ςd�K�3�FZp��B���q��0!_�,ƀQ��M��"�3�����������9I�ƋL��N��zkM����G�!��7�5�m��M���5_�~3��*W��*��(*������J�Z��`08�*���5� Zl;�2=�7z1EQ`���_K��?yI�JY�<�U�:g��W.�I���A��V�G��/�p�+���z���툘�A��ef��½Z��K[��1v޺�����)֒w���=�i�)�uC/B���ų��T�ۧ�q��AsE`�����/��O3F �*AO�ΡS�@�i\Q�����'���#2���s�E}�{ �5��C���J4_>�bS�/W�}(��H�b���m����?h[bV8>40�h�S^�qŋ�d��k��}��R锑י�A��0z�+�ՠ/��>�d<U^�K�k�(f#��
qf,`ۡ�x�R���v,p���v�C��L���{ IP�dka�fk}>�h+����|�D,�tG�K��ӆA|�Y�ͽ)���+M��ˌM��EG��'��HğOy.�IzM �Z̾��{J]��7�����Ee`���jt�֯��w>[A��ld�g<G��ՄB��D6�RJHS��jEi=�JeR��)��ߖr�v?�:<��s_7��X}j�2`���E+��0���ҽ�*�gG�I8�7� �lon�E�7SiӃ���
���>&�P@��.��.SP��wLJ�����k)��]��67��"�FG�9};�R�*���w&~Z�lו@Ч��w����p��-�Wދh/̂?�pݐ'�)s�(�0�E�����_�$M��=�0���|�
_h}fž�)�.N�(�xP�cR�ݖ�>���lM�fӄ&���$�>��+�n���F��0�~\�ד�А�6�x�j�/l�A�,�j��Wc��ھt�NM�� ��]$�4���L��2��OL���c�/\?�������jfGa#���k�'�>� �N@��i������5���R�K��fg[�+d{s���G���g�n�t�|�����������Ze��D��7u�3������"AN��M���k�k��"�>,�L��Rf撛��)�p_����X���0ؤ�Xc�  ��r��}��I��{�S��� $�1+M�����y��0�T#,i�1z����W�A� ��B��W��B�;�vG9!l�4QެEM���ȷ;7D���z��n�.�aO�����+ �."����	4��n�]^�t��*2m=_�ax¶X۲�$�`q	ͭyJP�exk1�O�o��P7���>0)�ek'�6*¶<��m�G���2\�E{�e��� ����~�7�"�/��PvG�G19$j�Ղ�i^�f��V��V��ף�]1��o�I�4�1����wXaF����ȱ����J����kȗB�h���3k��say�y�K�0�CÛ�Y��~pb�k�kܪj��_���]Z���7��1�gM�1�Ҹ����,ZsdO.�H�!�t����d��ߔ�8�4�۴$&>v��z忉r��s�V�(�1*O*9���e-S�#�����S<�T[�\�(��Q.�zywLty���7���*79�b4�QSK�8X�Ʃ��ϯ_�^xB�gN���DQ�m��
a����L�x�%��ѿ�Ů.~��Q�� �20�m0�Q��Ԝѥ$j����tL=�o�	�X�4�s4�l��Rމ�Nʺ�ܼ�X��U����/�c3��q���V���xl��$��bC�y�T�ҋ�ڱ�b�y�x�Qy��%�T�9�ѡ��;3gT^A��i]�E�����1#�PQ��%sex�sʷU#�9N�!����g�FDceb0No%��♉�s��6J~l��2��'���W" �F
$rh�|��M���E��l�F�Ȫ����Ͼ��:�u�YAC�"��M��{�Y/hM[so�K'�憭0"�� ��A;ShIv���ꄫ-�) �d��x�:�M� ��cO���N>#qM%����r�X��%�
4�z��¥i��6P$��{�O���+�q�a���'hS���������i`5c���î���?E��C���&��ɬ�#�t�o\o�X��g�a=���A��n?�nH|�@f��dM<�/�`m]�ω��2�5�8�&�d�w��|�墶��:} w�	�T#B�܌�؇O�P!�����g��nW{	=e�CT6���+��|ޓv�G+l�4�X�-�#�	,���z�O1��֛\�3񧏄�|�?]o8�;��FKRi�S�y �#�2���{�R�R�l4�5�>q]L�A��,������2�]�tz�$�������x��L@��q~��I<Eћ��A>�E�&DB��͏!��E�f���C���x�r�˄��L��Z�&��-��ǒ�b�_��䉨�q��$;��&�ɕ���6W��ɯ�|5qu���]�.0ZF�dd����mh��^� �3�,?6ڐ|G���9Q��=q�#�OM����;ui_�$��xC:i|��E��O�d��@�r�&s>����D%��^
x<fK�����(Ϡ5�Aw�V-HhEW2?&�������j�w�J���/�GJ�M�y����=�@5��]�Mj��<�KM��px��d�ަ�ڗ��E�qz�ݯ��#2�n����K�]�P׆,�N���/Wx'2�q����R����b��{��^�\[����ݦ �
�TO�M��3
5&�L&�1�ywx�0T��������|]�9���(Z9GmlM'��蹯zҋ0�{Y],�j��|���Ӫ�A���*~�&�l��n���&>�O�<낆���jt�+'�*rd㢧�2�i�>9�0��ܰd4
�ٗx뱋�9�s��-��-s�8��kѱĢ��y
-����
��L�m��E��Q�ϸ�S�s� .H
(!�[�������(�o_����m���x��gm����?����Q�M����*a܀}��l67�{��01 ��ݫ�2��|Z�#��jS�+}ҋ�깚g�ŀ��~���K3�H-���<@|�)��#Ě�i���V��ΰp6�M�ޒ,�m��G��$й����@���Aq���O����?�ӂ/S�/���}Ed�w}S�Dv���	˽u�-����9���1�`s{H�W 3SL�qS�������/�&}�6|���y[ �ܝ0-���j����m��YF��>ˮ ��#^�.+l	�#ɺ���Ml��'Wv����^�]�ߢ�66�D��߽Y�5L����\HE��]�#�鿴��\��]��;K�YO�Pc�j��� OLr4ɝ���M��v��:Os��1�K������F�&�)�k�����Uu��b�AH��F����(B�v
�t�����#j��"Pi1{������q�?42�h꺤x|�*qܱގ�-o�n�E<?�Q�����M/�@c������('�%���T�v�ժ9�o%�J�p���'v���9��/7�nk��
���H�Co���T"�+<)n�{%,-N�N�1 0�x]�<t!^����W���	A*�MT���ɒŎ��E-Zm{RJ��#��<�!Ƒ~'7 �6"�:���ǔ��6�B�#�f����5�&�{����
�$��Q���b��F�b�苣$\z�뱃:�_L��D\8Tj���@o+�i�uP�3R��Ŗ�ym<eubQ�Bܮ�n2	#�k�� �;ͰҖ#���5�����L)�rk f=6c�BW��o�1v�eM"������D�`�c5|r�r}9��ê2���J�k2�%�r�aLK��kt5��5�j.�S�ߦp���]c��-!G��pU�G��`�Ĭ�o�DPn�Ш-�ze �*K-�=fJG�mg�rq7��s�@?�����c�b+��לּ>��u�|�@QE�������:Ӛ���ʑ�0�)�߱'H�OD�m,��nB* ��=J��Y�ٔ|����H4%%j�|iѵ���m<�v(`$��'T}�z����iϭg�!�>)c��aZ�y�Q&��)#6�X��� �n�A�+�4c�kn:�{G�.�+#���G�ǄeI��p���O4�MH=_�czh`!I���Dr�����㿠�niW���>t������eKlA1QS�KȞx���a;$	���@�����]��լ���}L����]�(4���『�����' ��gbwuxAZ$\0R����w����$���	%K$�$^���sc�8�tu~�?d��9X�#��I�Z�sgg�%�ݣ��ؽd�ƘkI�8�G�I=���*U�L���v�Y=�{+�m�)����0P�hD9Yʾ9�Q�c����0�.�dMDR٥?$�g��2f���'�/��iiL�	ud,d���n��C�p�$��ZB���#���[��6b˨�9IV�6��`M7�^�@\���z[���3�A!�b��/��T�%�;��h���L�#�S�uC=^%Х��K��-�/�_���P��.?���mu�Xr����yaT��Z;�?Y�쪐o�z�/��$��z�PC^r�����}x��G�k������$>_-<\F�{N�q��:@ �2��ٽt�J�]�&���u�Q� ��ͯ�_2Q�N���)�_9��&��j�i#³�Z��x_���O0d�-ACY	N��Y��y�X�^�"��얕�Z�'�A����Gj-dJ�oF�6�٩%g@�7�Y�$��$^�ˎ�RNB�-u��ڝk�K�y/�.��F����W[H.{w��Ve1�?U��M#'e�1��ߌ�y���{��ys�S���l4��r?T�v����ΐG�Xb���P����m��ﻘ�#�U���}�:%��f��V����	��	�Q�Y��`qN�K�x�������$h��䰭|�qb�I��2�v��j4���{Z� '�?��3��-M�+HD\�Op�2o��Ԫ��Y>ؘF���_�����i�I !۬�H��Q� �Zu�4�ξw1 �=	�����a�hN�Q���p\V%������������b��g���f@�[�����2�J��P58f2n#�PL0j�2�چA�P�X�y��\R�֭[v�#����cX26�e��G>>Z=��"��|�zQ�����:�C�����9�(2X���F����%���l��AQ�G����́����2}�?�	��kt^�CK	eS@��>ͬ��
�Y�L�ek�g 0����.h���b��쎊r�y�\eN�2���[��c�n�FiB. p:�JP�Լ�Fί�)H'���k����Kfaz x�
�z���E]��a�6�k�ķ�Bn����[1I�v����O�%泸�xn���!� AE9O����(&�p�k�ps��BK@"q?���ð�����^N�UX��������:#�i�oןϟ�� A���l���7��F�g�� �.^�N`��"u@�6F�ৌ��U"��� ����T!����,����8�1��s��iF�;Q�U�y��&�̄�dCa�ʼ�~]�o�x��hJ&zxN���	���w��B#��IQ�$9ڰ~���7
��pH:wv�9]+�FX�:��p�Z�x�+$�,C�f	����3}{Np�Κ׳���(���C�=�Y��7��e�ltb�,��@0*��d�Yh�	�&i/k��-4��Tq��k��Q6�����3��`
�e�cZԀ :������^J6w�U�c)����bt3k�*�=��h�ֻ^��p��eͺ�|)j+
�е�V&)��#3Fcye?��Z�䛃����JAcB��L�~��9���7�-m�/�v��jP����ܹ�W��~l�e?�H�V@R�a�/�@�֗q��-QIRc��
��4NhL����Oձ�i����=��n�i�����T5�ǲO��P�A�թ#k��]�t 7C� 
�˔bS��㰷�8�x��(֠(.�.��K;6�5R�T��j������]�<�#6�����m/��� /Ѻۑ:�,],Z�|�R>����\��硶�_,�1J���$_Z��Ǘ��N�y� Kd]��!��JuT����VO3�</����
��X�s̚��lxr����� ���(�f ��)ܸ�b�fe�c�u]%���\
�����O��,�:��~������������*;_��t�X]Xx�����;2�tT?�<|��:�QA
b*Bkp�����ԸBP�
U3耲��b�F$���� �4*i%F�� �mk�ƥ�)��6)c����%��a��M4ɡ���Ҕ�vi�]�~i�	�؃Ԉ���?��\IE_��(Ci �3�x�4�U�� X��U�px��ƊJ��/0�a��KO3_I[A����׼���XV�:�X�,�s�}=��ڜ���N"�:Y!�Xڨ��Y9���1ҴFoX\��WC rXOy
d�������J]nwМ�	��i5�ay�ٜ7��Y�b�OJ	�I��)+%wiɨ<_j$������!\��0Z2��"i��đt��y`�
@�G��1�oO�ă)�EF��M�	�Z�?xN`t♒�Ϻ���b�L�!L�=�zO՚�M��^	�=�#�Wu�Tv������>_E>�����j��2ca,�냐|�S|񒔣�Nb��T�C����i�񃜆[�o �5�����!�`�P�M\�S�D�I���b�W8ɲP�܎����!�(��N��%��ox���M��B���F��36eN���+��c�]Rص邛Y��*5��ł���~?����#�F�m�V]�!���>S��	u	������!%�q����>���!��u���g-�9�֔���MD�p۲z@�$j�2������hs��[�����}�P4M:Z���������_�D��	�1�
���`fJ�d�s�%\�
9�#|(,)���Ǟ�ۃ8ik��N��l�ӊ�>V��s��@�@��p��t�r�=�6��ː��͢k�1�}�}���k�YA 
�}]*�%�)�B��p7���|;m�=�.DѭTy�+5L��o���g����aѼ�:�S�-&�0R�����g�����2ݟ�B+I�`E�%G'���r��]>k������z�SܑdN�`Q��v�ȑpԽL4l�çO�ؠw���p�RO6Мת����ċ���;aC��k���)�֟�{S�iZ���V1 I��t���ױ���p<���S��\�=-(��#�O�훃0���le���\���k�-�M�� �ݩ�<H�\�n8+��ӆ慠�64 ��cC*=G����ĝH`�a�V�,��ƲzV��󳻭����5M�U�4�`����1�<H-���ɹC9�S# �3��uY�S7�0���>�)"��
l/܀y��s�������+4��3W����"|L�'���ǍՖ�ykډ�) '֖��/�p�U���^G[a���"�"/m~�U3������m�@ҿ�Wm��B��!�R(0ֲnpI�<k�W��Ln�
�4�rY-	=ߦ9�3��!��E .T���i���ť��MXi��дQ�p�HA��i���WB�UJtΖ�z�HBY�Z҇GOs��N��0X(�
Ue�\V�-p�&]%��SK@8�A�t����,:�"�-�?�%�~\d�7�3E8���@V�+В��6�/[C$ORrh����~碧�v���;#����ü��ؠ?��C+�x⨰�<�[�I����3qB	G� ��<���*3�).I�5�:)�`����c�7��:�k�W���}w���<�y )]���yBrC!�bF~����Sq
�ν&��XH~�6�m$�B����q��@b��ϵ�mzT��b�oo��a�$���KLy�:�2�1.����f�d*�]p�C9Bz �ā�ֶ]B'J1d7N�����B,��R0�T�$����l�K�i��㠗�E�?trz�NىI�*� �å��z�|�:S8��ڼkc2-	ho�p�]�Y9���^*.����1|qG#-ao�*3غ詗;w�
�R���W���X�I�>�a�#����_e���ݡFAȩ)4���nA�,/+�)6˵�K�\hV�����G_R�"����?�Z�R}���w�i�/fT�n�.V<�����寠(�qP���Q�u��WX�I��<M[��t���1	�5 ��ZÊ�d��AgBZ����/�s��"F�7�!�t.��w�l����_"��/A赘!۴n���|�Ӹ�B�եkH����Wk���r��څAI�+8q�#	�DP0�s��v2>�ݼHD��ڋ!� ��=%+��8,�"U�n�yWPPd�,>l��'5����1M��T���Q��Hr ��%�L'1~�B��g	|�L#�=��+<�E��߷1�fc�ɦVN����y�>C�e���#��-��ƺ�K��e�q�hĲ�*������bt�M'��w�7��ty2�+?R苊��N!����!s��.��I3d���g-�U���!@�F4L��Z��X�`�Bj9usW�������0�fZb�[��c��|��-��v�%��1��0�|I�$q�nS��o�3�"�ٵ�
��?P�B6���P�܋#|uq�o>���� ���B����E1T��B�ܱWk�$q�����,���eG�_�<6�V3l��b�	��$��j�^(�Z������h��%��ur�1������D)(e�p�m�L
b��Y)"��c��F%��p�.Xϴd��:�a�����#C�mm�~��i�o�D�%���̅_��2�i}nwj�B���:g�d���3�vC����c7u����2r������萞 ���!�	�+��L�}L�� ��닿��"x�蝝$Sڴ1�=��c���8�n��=@ܻ�DkY��с�J�FW#�U�P�b�g@ý�V����r�{���.�>*�&�O�r��ͪ-��	�(���L͂�lY���E)w����B�P"d71�X>g�[�����s����>� ��ǰ���&���HS�䶨ENC�K�������C��(X���s�\�p����k���ùY��m�?�~k�(4������L`�}o���_��%G�@�Z�X5¼��C3�/�{Ӹ�۳|+��G͐�όP"�_P�*d���*�t]rX0���>�!��8}�Z��J-4��&�~�e��e)��yC�k%#�e٠HzU&|�xlc�U���y�J�厑s�X�੍j���3��w�S�{��x���N��8J5�:b������u5�~��[��Gzx��r��}wA�uHf��Q�z���W�w���:*���ODۦ}�r�z�4���$P�,�h��#��J�4���Z�=1�L7���:�i&����^�fj�"%����/�ܻ�9!!���ܳ�Z�����'�z��rT_�P�@<#����2���qx�/�込Jr�\"��=��ƹo��f�䚩�ΑƏ�7#�߄W&D��s��w-�w��|��2��4�1(E��p�'a��%;\����$�ßv��� uH��=9U}�'%�1hA�Ʃ�I$QH�L����MW����&#��$q�wɠ"���	�5ey������$�b��̮���[��K���p�ҁ�=|�����ɂ&W�b���o�XN��Z��K[Ŋ�N3!����!T[1ڿ;zE]=�f���E'J�����i�=��q�ʵ(]��e|PNm��KCJ���YS,P�>�S�����G�2��7�D������Y'0z,���Le�H=-ɺ�<�̙��)J���ԟ�Vi^�P�>�;{��J�rЈ�5:�nQ�(�k  vi���0y�,<�*'�������\3;�D���9�5����
�Y�r���P�㼺�V{����ߥ�$G!���M�xކ�U,�iQ@*��X�&�4v߀��\S����eih�čH�p�)$O�oo�Fw������*m9�:��
ʭ#xK�\��AdDqӖ�{�^�$���[� ����.]2!��#�I��0�4/Q��;�E���:�R�Hڔ�;��X��Q;�J���ڌP��'��3	�Gx��g������"�B�r%"'D^�b���j��ܷ�sS^y��ɨ .X"#r%�>T�#�Q��m�c�X��w�d0��A�=�������TwŚ�w��	;7*K,JR5����>�a��i����~LIq~"��^61�䧙��:=.pR*žf�p�Md"<˷��f��	M�?�]~wY#��3�l.�v1���@������s;��xEX�_�|
s�	F%�� 8:���u�[� C�$F�Hb���(.7�U)'�q��^$!�8���χ�f��Jq�����f�(�'�<~��g�-��Z�e���
�K����4�d��I{G8�tc�|'��r�;/��G���P��4,</��A��7�Gf-�#�\w�
$����۴g�#��_�(�v��<+��9o�h%-O�ԩ���S�Pť�Mc���"����X�~���ӑ���eG�g��3�@gsG��2|�;r@�.�0����)$H�!7ӕ^B�K2��)NJub���v����(��CqIu����~�ΪN����I��J��8�n}��佀���j�Vr:T�C�fyY^=�+0x�Y�I���=�ִR��@
�j�<�KL�C�����8��`J��ea�G�m�2�d*�a�`$6c�雈z_�=�n���2��sC�1E��� _�%~�G��s �1'+���:�BT!�*�Y�'��/l�f+�u���ABz$L�m��:9,-J��O�.��~Ǯ? ���P��6o�Q:�XJ ���g��ݕ��'�>�Kq��IMG.�Ȗ5��q����]���T��1�]r�����f/dl���� H}��]��\�|�:�q�G��c(�{���� �%'�`��g!g�N��*�@z��E����Ԧ�;!��CN��ߌ>������^c���ȟ��A���\�@"h�=AO3;����6��XL�@�m�.F���:�J�_�Aᧃ~�3A�Ϝ{��o����Bj��ɸ����AҔO��{��y��g��8��,���<��Q%��=A�4x��iux���dz@J�R����K�n<&�΋v���2�����k�b%����ܷ�a������E�y�-x�mb˯�h�3q���L�"�P��->��(H�tk��Tm4����S�o�K�"hq�2Cp�jK���p�0�+�o�Gxj}��?p���h ������:��8?`�mj�*�ʁ+�s����R�KEШɗ�]v����_�2���H�����p�=5=8Ţ���}���K
�'�D��t�8v�!$x;y[���b��
�N:�YVē%��6z�<�����W��s75B�6O�K�z�Vô��Z�N�4���m���G?
f���6O�Ϳ?�ZJE��b�!�\l���%@����7=�;�5}jm�����X@3f
%�����"Bˍ�S7��2�n����hJZ���*�mkِ�P��՛�Q�*�=N!B]3*����'*G����э%�����)�� �Ԅ!�D�2Ɉi�8��S�b�p�A������b��O��"D���~��a¦֮�/9�����7���e�aER`E��[ �3��m�gy�@w��:0�'`x s$<����jJ�����ά�y�ovnނC�.-�.f��X��{��)%�dʙ�v��I��G�S�[^��y⬪�^@vĊ>��\��"�A9)������`��R|e'+T�����c��\Lb����02�'�<������b(�%��������������?���Z[}��������^U��|���d���w�l��'x訒���� g���&J�.5U�7���~/6�&����^����u�@�EpU�w�Z�}!��!����;6���ʑ�'D|�m���x,�XC�!�u(n��Ԯ��X�'������G�&�c�4d:!᩺��>[�ɔ���?�k�rQ�Lo�S���ݱK��q������
ғ�q�o�js���C`e�*kZ�x}���]�a2�~��:e~?�T�{�5$V>�V���cj:���=�N�Ř�IW�O����d��rZ�@�H<0��=��M���'�<�*��P9F\�{�]�E�׺�4�ª�h�7��)3\}�g `  ��RI�T�O��^C�\F�XHH�i�G���x��=;���oat�w�`妒>�t\����d#�a�"�S��Q���e
2������)`SZ��B��s��Z�W���}�D������M��JxI�=�-!�\���^t� %/�0��%4>6�?N�Z��H��b{Ҥ|�*��+����O���z�M�ɼ�M��􍆮No�7u �L+������ID}GZ��g���tx����YLݪ���I����(:e��%{��0ݱ���qdB���lLmZ;�^�v�����_ %kHE�ma�~l�M�I���iC�B��F��8ܲ�1TOYYM8�����ǩ<�yo,��\���{�Z�*��K��Ϋ����f�p�6�	Z����m��;u_�*�gd��s��,�К�⹙�h3]�=��� =BDR`�t~�!�-���U	5�ӭ.�&��)r��(sE��~$i�F�'��?�c��@S\�w� �)P�K�8�����<�o2y��f�)�"���O����':�-��)�&����?�]�i0*Nr*��ѴwǨ�x������V�`�q����ME��)h9�7î/Q�[���cO�t���b�8�ֶ
VJpj���a�X�\.��
���G�񄨏S��H���-M���/[c�
��(���Un�*���+l��*2A:��M��w�,6�yn�'kͶz�5����mkW�e�t�]�#?
�׸'J9�_f�Q�۸\N���Üᚺl���X�,Ěr�p��R}Ě>�t���my������+]��$\�����u߱�f�O�nV����@L��1�?��v�9V��n�_6ҏ[�N=�f��'R�v�1㷩�ɮs6�8�S�L�gx�14�> ��Y�I��,:��%�^u��i���Y�z
q��}$�*R.}�O[���/f.�U]�Z`��f��,� ���)�%Ʈ\]�ڜ$k6"�n�4���<O�=x������*��%�:��?�mcBXߜ��[���z�Gт|��p�Rn��{�e��e�%�%H��B"Xv��Y�
3��=�0��t�<��tdB�r�1��8R0���Dv.
��<�ߞ{�V�oX���k�X�t�����4]��ح�b��W�t�n sKs�B�g͊��ؽ
��=L]XG��_�|��zo	��Z��Y�,��G	L�\Lb=��sW��s�L�銚���jt�� �8ݜb��Ŵ8���+�sM����D�������|��M���W�G6M�T�<��΋DMԃ��Ac�s�~3��c`1zј��\����#�>�NLU�JZ2�ݽ!�����Eы�A<S�'�1�tpU��U��������� m�1�o���-Ϳ�~�nqU�Y���Tf-���+�XdU�2���5����ل�4�$Y�cy��Fo1ߋr �Ik�[l���ң�j��;v���%D�V.�d�^TL��R��A�$�q5)�Y�=��=�Ҫ� i#��4X^��!�I�Hnn����Hu�/�ĭ!J����:��ō&4!�݃�0�cw��okwp�օ�0S9���`=��������a�#�{[ATp8���"��A��.b�u�Ϲ��}�S�d�K�ZyDy#�~�;zglK���x>!0�	�3q(�E�8@�����Ջ|� �׺��ٴN
\(�-����^ʃU�"���!��}o)@���c�i1џ�n(:5^g=�ݘ\�٦F�����7��K��?L�g��J�1tԥ*���6��x�R�t3j��0 [�)�hL���=~3����=�!�33����?�X($}�K���ZM�	��ѷo�Ho0���˺S�W���2�O�u�&��K�7�ɕ�
���ݟ��Wp���WU��*ȹ���;�ax��H0��&u�H����=}v��ΐʅ!��ӊb`5�rNAV���Q�͕�K;c�Ҝ�K�x ��+xc�*�4�pJ�����Om��n;�_���D�
-P��C��d�^$�Mncb(.U*�z�� 4�_5a� I��{���&WW}����`l�GP�lFI2��~<f� {1�Ytr|t���>O�7)�uW(�\6��(�'(%��z����@��I�c�z�Tu/ڲ�K��28��v�b�A���eu�&��nz�M��b������q&���*u?T�V)��v=�`�%'� K(�^t��3n�V^��K��A�[ƧLhg�[s��KL߉#W�T�<��U��� :O�U��'�|��s�;��S\�s��{՟*�kjO�5p�P�4L�c���"߸�L����}�!�>�b�[�� q,��2BM���?*��Q��mD�Z��Q�~6��Z'i��ia�e9NJLi ` ��잤�FWy�"�0�<�&-��$���RA��#,���7�+����_a�iJ��_фB��V'p��<��KNM?��RP�zk<���f����q���`ik4*"Q�խ8ޢ�w�ϟ��K�����V���2Cv�~��xc�A���.�|g(�I[�o�a 6���f�puT�:�D[,+c���xG3{V�@���`�#2iT~q��s%3U0�y����9��"����r��G���J�d��7�umT:���NZ�p3�0i�\K�<����P���M�3tʜ>d�f��K��x�)[(�g/n�A"d��]����v�#ݳ�E@��*3^�������.z���9�]p����,Q�='7۪�|�	�|
�����yC�����$��!�!�K�38�v�R����n�{��o��@('L��34�#9a�%�h͍�$m���&i;j��=�Z�7rm#���m'�5���Q���7��w�L�����JҰ�V����U#o�ڜ��B{/[�C��d�)�g�`q&�#jʓ'�)	ZZ���Ifv�a���)�W�ۚ�yX�+@��Ǧ�j�<cL��Z@j������q殑vfz���$U႟�W�qY���E�e�;[3ݞ��;	��@��Ce�9;��N�d;.�7 r���C�z��Ҭ�S�͞ȞF��^LȎ]��[�"�	��.Z�D#���sX�g�R��a��]����k���������=H�J�I?R����D �ʕ��$S��p��MNfD��A$	?�{ȷ�6�C6�l�Rb����0��|U"#R���*N����@�]C�:aW��K�d؋[��H��;��9߁��N�t =j�!~���EP�Br���������+{�[�@(�������wB}t������ӏj$�u�X�嬳�w[8dsz�
�~����[���m'��496kڳ��P�
�["A%���j�~u��K����L
���ܘ=�	�Η���\�<���䙐���A���[(@��Ү�19������R��.��!�d����pK�y�B[�Wj�"e��>�MCs68�-Mp� Pm:!g�i�˶�4u��*M'�O�k<�[�Ž�1�o�Rv�h<ޙ8�sl��3��Qv��q�6���5��A^� LG�n�W1�&n�t��,�&�Пl�.r�b�#�^�3�a�WѺ�Y8Z�ڽ��~p�"c������i�w_�0�0VQE��k��Rb��f�t���\g.^�]�u�~��&���0�OB��σ�����K�n����`�[8�����_6^�K"���~�q"�'=k����D�Z+Q��њ��J(�`*��j^D�y��良5tP��SŮ�����������r;���&��V��:�ɿ�27 ȓ2m?�Ik{!���}�|����pN��2�?��!���N����9a�s�e�#
vyT,Z�����7�`���m�2tA���cV�*ʡ�9L��k&��7?����,3<}��'���݋��/�Q;7�BK�Ks�A��du���Ĵ�^3o���ш�*����ܪ$�<]yE�d4\�I��*���1�&zc>7·��y��j��ZU�Ȭ۠I��ys%��o������)Ό~���!��A���Vمe��ݖV
te Ƨ�!>�b<�ԺJ�֊_ ��[p��f�py�4Էv�7�8;?�6�.�� p1�n=z�B�-,i�eЙ��Pp���ASa,*�rN�&Ov����0�rYf��'���2K���{�>W�\cZ|��M�MIz�b��1?x�B�I�j�p%+Y;*
o��A�VNBƑ@���8�`ح<�s�e�-�+�g��4������-%.�t�v�<|�I����|� �|�TjZ��x����S䜫z�@�b�I������04(T�V�vî`�}U7>�*�C&�.������6�k�W��0�kN�"f �%!�ޏ��]h��[$��32;�pj��G���%�̲<b�S�l���=�l.p�p,��1�32���`�)O��$TM�$�Kp�K��^K�{���Жya�pm��Gc`��Q�Q�Ӿ�	}�?N�9��8m�Q��D�Ne��L��/� z�k��t�+/L���<��Zp�\�,}��ͮ��pW/�ڬ�
�^j\&/%Q�F�P��w��S�ｸ���DX$sV�C�(�!YQ(���>cℶ��ϒ_�
�?���𰧇W^gX�nC'�HXVvO��IIdo@:�k�ʽ�!�V��a�DSÝ<��f�W*	'��W��[(?��:�<v��*�I���@Œ�Q+j�{#�sO��@h���0�F	�||���>zƤ��O�> 6K.�E3,jZ��*�Љ?S&M<���ǏD�D��"�ʺ�a���=�s$���籛�:Aڝ熈��xcn�،�A�����*ݕFG����ϣ�Kq'.�h�tGK���'Q.�G��?ݱfZ�XFx�,[��"
Gx�9��_�'�h��v��VAeF>� 7����NJ��|��u�m8�@���V
�̚p�&�`lԁAi�!?t0�&��`w�q�%�ջ�0�6�>�VH�&��s�N����^��u�ꬂ�W9�f��4У�{���q��!����gj���X���=`�;Q�(fys�z����ji������"�.&��Q%�����,�fOݙp���a�G�?�y�C�=�q�ȝ�;������;"�⾚�$"����2����Y�4��R]�o�B[��ęoHVS ��a��i̠����{�]r�ՙ/���oqF<�a�4�V�6\�ז7u}�&��Lon�
� �
�'�����PE1�-��8�[�wY ]�:�,�N���ظK2��v��!�qV[K^�P��a�<�
����Ѥ�,8�ƒVI��, koD�Y�iL$(=� '�q�И��]�b:��^�UZ��~��h�y���u���&[x̎�갔{��G�)��#��˘�R��$_&�|SJ�KI��u5�oWڽ_��-�1P� �jO-��IK�9�.�ⷒY��!D����i�H�&҆�Ȏ�yآ�)ݨ"���얈�9��@ڻq὆�ߡRL�/ 7��
��Z��u�V����N������~%~6H|S�qh�x��fR^� �B	!F�M�)$w�9[�ai ���周�N��?�����~;8�F��:��}g���I��
���,���ԃq	�\�K1�;�n���IP���4��[��	t�������s�����v
W��1I�NT����h��o�Nn�g (���E�vqf�9^�M����]���M�,���ah��E3��sLN:�h+~o��W��qwIȉ��U����=�J�*YTP�ֹ�;�>��P���o^2D�G�q��_�]s��7+�����˨q�YhV]�Cf�_B��&J����	S�F���Ԡ�<htc�ȼ��n��p���t�?���,E��ԟ,�U��9LL8��.^��u��n�1Z?��~B������e�`E�����a��ƌ���4g:���R��������@�U����y�J�+�S��D��z]�(��Ľ��nmFW��;�N��^d�����B/a��ZZ�t i�qC��\�{��n���y��o�� �-�������gU���I��8����It�.OT+9���*e�M��M���Hy�)�]�!�,��^�����R�(6�_��H�?^��/e��[��Zs�d�`�駰��Cw��t���,{N^^=��a�QܦYT���������:�m�)D/�>��֕�F�\���}���48����Z|�x���^?[�>=����ݯ��$�px�o�χ�_p#|M�s�;�S�I�ׇ3�n2Y���3
:%��8��º�NW`p����,
����ۑ$VݛU�1��m��):��3g��*9�Ѡ`Zע8I��77s�~kC⓽޺�!��Q�ߍ��T�)�>/$����?@���{m�q��ѩ/��z
�����ai���ii�*�f	���O��K�ƃO)��8�V�RJ1�����{�C�EW���.�[���&�uD[��~����{W⮬��<�����2���5/�3e!��T�h��%���.q8ѹ���5k~��s�!8�G-�����^���yc��f���:9�]�Zɐc3�_���m�&�T��y�0N�'��9�w�W(���	���uCV���L�6$N ��hn��K}��⛾v�wz�ʮ�V�;]��������?_��m�q~�
�
3�#$�����K�7�3@��#:j���Ӳ����I��n�s��92>{"���Q<�bm�$vr�D�~��%F5޽���Ãb�r�b�-��0�e�b3=�0��Sz|If���y�(�0��' �M�u��8�!�j<q%̽�}�Qi�UU��\��L:"h}����g>�I�Ӑ��ڑ�B���i$�̖����"�ںw���FP���p��t�"����AJ�i5O�]cwN��Mc/P��iq��>$E�6�E�.�0��Yw"s�S�'����;2TG^�Ҁ�/P�e�,���c?7?�Ij��t��ZL��0U(4/�����4�ٙ���x���EE��/��\�o�9���I�x�}�����[��c����J]}�Oݍ�N�S׆Q�2Ć�`��r�Ŋ��o�@�1�RlY@oc鏧��!m�4M��Tɧd���W�Y�7O3��f��R�8=��$3)@C�{'�O����x��۱c�Y��
�ť���E@31Nw�faW��^�j�~�����f����sP
7��o�yg=Ϥ�{���=��n�vM�0��p\|W�a ?���<���7��-���l��b���P����؛��r.�n��o<�	����Y�P���^���6��gj���PGs�U��9l������sǀ�7�RE�cKI�KX�@.����U�>��Ē܅�s�Q�IB��H�0kc�R�7M
N�a�4��p��4���/ό�˰�o@��a���o��������+�-�9���_� y��I�pyb��)��VF/Ie�6�̳Z�֓rbPZ��^�2��1�Y���Y��*���yǉ��B^Uu���*f'1�͞Q�d���(sr���W�]����3L�@e�yB4:���0��`׏��I��n�䨧^/yc���jmʟ팵����U��a����6)�@�Q�ջr8�����m�[�7��=Z�/��Q�o�vՔ��c^�B�v�kK?p`�͆���ޑTzK�f��4�;��f@�Ut�V�,�1�%a����4z�J�IY։MCd�b�N�!�m�$��x^�oU>fl�:s����!�s)V	�����i��bQ��v$&�~�2b�	 ��24^<���#����܌+�������b;T���J�I����C�;)X5��u��}J��t�tC&�[��ټ�sOc��� ����pjP3���.V��DÓ��s/��S��/�p���]�ֻx�����)��ژ����Ǥ�a`��؜�촥ʱ�aY�/�)�6\P�DW�R3Fk��S��֦��(��ɏ����T�ݓ�ou:���FeA"�_�M�� �0+��1�r${��C�E�L>��V�|$LC������73O��Fby�f �.�z
3���j�DJW�ձ�
���ŷ�r��,r.*��ʒdNƫ��n�<�c|�����:j��8���*�#���hT�'�N Z!dG��k�V]��j��u��it�BoEK��!�W���4��/?�H(�rݾl�!�'�s
{��x�.�K�*l�����žZܳ��*X}�tB%�'�Y����{&�.Rm9>���������Q��I� h ��~a�wt��St�,�&Χ*G��%v�~1~����^�{��?ݸ��5z�"�Zȯ&�u��ߺF�˻�m������_A�%![�����|��磦��,u{�Tgq��?�4
Ŀu�:����槆a���şT����62gL:�<�΁ڌ>����`C�&��J�Ԇ�,���SEY�b��>��Ksx.�؛$�����XY� ?�~	X}�|7b�P����$!)i�z��W���A��j�+���i8��oSI؃"��v[��C�)�O�=o��3{�⮻wMnW�~w��LKA6-�,�Z��-�4���u(3�|�Z�Muze���Z���8��DO��w�I�d%�F4x��4��Wr��9�M�L9rV*���$9�c�ӳ�[�B�b?IL�����>
�N�/�r:K�#�I,荆�6tW��D�"���oZЉ�mS�7��}>���r���
���_5��̲�W�X���%I�˶<�J1�=PM�^l}�r̼w�5@���6���PL߾�'��[ec���q�8�N�d�# �˴���h⍋ŬR��� z���{���W�[}�����A�|�>�L�ir��?��1�:��Nr"�s��w����m�RD�u���y�l-S�ՙ�i:b���砨6���>�,v��:�R����U�P�Q��-4�ӥb�w�Bu�,RB�2K]_�h��Hθ48A&�<�&8Y��q?�P<_��2��O�l�׭ٙ�=�d�a�5d�5h=�#�YѴ��odjpV��n�tP���2X�ߜ��xp�Q�z�K��	FY�(<���kW�Ԏ���R��t{g�4���{L��t��þ_m�������;�;�'�sH)UT��>��-OZaf<׶x\�';.�ւ���Y�w������<�ލ�͝{��܇;=��9ro��'����T�'b�0jB��m`�~�߹�G�qeqj����3<��,��~F�ր	cQ�>b���/�iV7�x\�:pء�������fiK��A�	��˰޲�睭��s&��p��ݙ��n���Z�֘�0�en����7��T�8,D�J~s��q�tQ��zY�����$�Qm8��O)A���-~!����Υ���`u��sg�J,�0�,�|�s8�y�a�`Cd��؋u��C���B�l�
�S}���"{	�:�Iw����C��9T6x��J.�ά[����3$�K�U��dڬ��M��>���uBA1�6Ǉ��(H��-��}�;l����GOe�7N�j�."�� 6^��}b&�-��a�A�w�!}�]q=�U� ]K0�����J|2)t���%t�׻?u���D�!H�Ń��;W�.��c	Ű�鑓��I�;�Bo�?�@�A�|� _=O%��n�-�����p���[��,�O�ft��VV(����r(�C�d���{ץ�r[7F��Dћ̏�yr����O��7=&��LuMyI��3�B��m|=N�X�����]5Oщ$�%È���u#�0?��暱���L���+��~���0�kI��F�y��e�A��p�M����Dd�T>���	%1?.3�D�I����.E���I9s�C����1���%�@�_����0�:�
7%BJ��&�(�kwPgI-�S��n�P{�-t!�U�T^@� vY��b;9o�~�5����v��`�r>����U�Xl�A��%m��/`	A�<.�W�34����Gn��o�y�Z�8��B�������km�j^��S_Cq����P"^D�7���`="4���-�7�Gt��ـb�'�C�X�Ok<�GNtф/�Z$Lܩou)3Ir|�w3���fFt�i�/tU�&t��x3�c�=�/��X��:�޷&�qb���EE�J5����9�V^Vө�t'�b����jpt`�r�Bb��4Ub!�I������O^ׅ���E
CW:pV>�x1��b�$�o�n����%GLW��v���2�"�J��M8�yfT�\���iR�h�{�jP��:���3��<3�B�����9��/�i�s�UY�jXAk���X�3xs�~족�U����N��&��䝅��g5�Sٷ��σ��;-��Za���
�߯�߇�qfɿX�;��K_�O>��`�+��k���~���G@�Wz/$ù��&+e'�X�x�阰�A5;ۯP�u���A� κM���c�3K��yBp-(�yP�~Ġ,�|��5��O�u&��l����P�W�-�Jgb�pӓ�j9�B�ĻK$z�;#R,v#�����V
�)/H�ftQ4�T��tcyg�F�L[w>�,��7�A5ڽ~���6����8)K߲9��Ck��Qd���BN�4�\�Wֈ����.q��#0B�f$� �Tv -Ͳ�0�2UePK�rб���2Ӳ�A��W�f����	a���Ea� �)�&䔈o�?,�bZWk�;����@byc�~W�8���H��f$;�X�$ ����#���}t�AVejYj�2���-I���v��*��9@h���G�V↭0^��1oIX�n�cT� �E��1&�u�`�t �����]ä9燆S��r{�b3Z�&�T�m>-��$����F��N9R>_(��zTXbX|�䑹�Z�`���ш���z���̕��:Wl2���.l����%l�r���$vb��L�l�9�1.mn�6�I����b�1��)(�����NW��3��d��=�H�D0G���dW�c�L���-��$�b	aa-L�f`����Z|��	/���!��T'��,�X��E�߮9F':`3���W�盷���i9%<��о�1���a�PK(���|���k�Oa�;)����V�QO�:�Wϲ�[��f�o�o��x���䐮`Ж;�Qg1�2C�� 7%�m��~CE#�~EnX��5֟n(?�aF��|�T�v!�W4����C^�!;��<���=-Sm�X��oB��&�s1�_�Zj�x��n j������(�д�-�4e��Vu�Eg����oj(T�ԅ{đ�����&Ì�?�(Nm.��8���]W��_�L��lP�<jM��u�$9R��^j�����V�⦆���"����WT#�%@�&~�^B��%��Ź�F�e�m�*˄�x�������Nx�
��LL3?�|���#/O\���|XP ̂��E>�y��إ?@���"V'��w�2�P5!��R�L
���6�&F�z �L��'��W;��,��e�s�~a�|k�cu8��d��~��8����[�) 
��f;�CVW|�p�w%����i�rV�UVelM���fLc��������u05���y8��p�_vbc��͠�|��˃F�g��� �.#>�"}�OV�Z�ЬC���9��ֻ�s*�������M	�6㐿20v��hdrs2U��.I�����.�̴�<·lR2L5G����>�:���
����򩢱�צ�U�-��٪�}�3�M��<�JZ;K�}q�F.�f$�s���@��EjN�w";���ʁ��ʃ�(�W�+�l��ٸ���9�pͻ�_�oFu�|��yV]1��]��V`� ꦣ��������,�{��R��_����r8��1��c3U�U���q$'�usB�yz�0/�ɧ�ڻ��$�Sc�B����t�f"{�(]��єF�08�b�bu�!:+k������ֽR�V1+�je�sW9vT����^{�cN4�ju	�u^Z�sH�n�,io��)#A7��
r~�dYG-TC�9���m��ԙ�̚s��4"�s�f��R���2��,t��d�����I�w�;�o�l{�hS����9|{��:Z��FW/@��h�<�@p�mim2[6��u)5j~��<��.�O�.L� ����9�`>��s�iU�@Š�?�M�Y��i�L���u[��/k��_�H
�0��aׯ��z�(7�A�v@�j��n9���WفHcàH`%��l-�	ar�$��u�yA�/�塩��63U�?��-elH�10-�����Ϊ/-����À��N0�C:��/FV��f�}��x��+����w��1�?�����X����Y��[ĝ��*�3e��>�'9%6ktUY�w.�����0� E!	�+�+�����!�?����j֬�O3ǜS	��=A�!T����M��Tk����YA���C�[�T�3k�i��Dn�1��&��휃.N5�H�H��z������6��B��P�YZ�J�9⠨��Ԁ�mʗf��j��k"B0D��b+j���<�9naOp� �T��+d�Y[��Q�v�b��k�����g���˓Q�9�.bj�I�k��E1~�8?=���^�䌎b�[l�Pk}�馻X��bc�����5�������w�X�6r����`�i��د���IG��u�A9��ռ2�%���U��cI@� �3�*.��T�!��;<�=��0�LZ���0��hݹ�_�j� �����5�?�L��:N�g��ӴV�G�9w�V߆&DQKh�	��P��EĤ<����
��o�55o(@��B��A�����5	�)����c9^������ǂ� ��T�$A��[0����Y�_�M�gI��%2������	a��R/���pq��rM'��(I� )�O2�M`q4�iPU����	ҩ��[��5�=k+��J����gя�Y��Ԣ��A�
|��ʫj9�y�'0*Z��FS#J�a	a�"�x.K��.�j�]	�=K�5)�*3n�>u&���^aEP�`�]= ܱ@?�kP��2@v6�K�Ҟ�v�Ӛ�_�hX:�E0��>�S�%<zE�5H��P����a��>�(/a�-	�Ub�a�Sz5�����(�L������ݏ�0[:����_�c	[�ӿ`�����(|�	S��U� ��ە��j��8� r�w9k���u���fZZl����˼o��1􃄸~0=J�t��+�j��[�����'ʰ[Bz�
"�0l1bY���0rT�A;��rNXwc�\B��y�T��|�D/�Kry��'�a�B�����Q)��)��:��b0�<�46���ʵ/2�F��j�*�7%�	�_W</�i
򒵬S��q�Ɔ���h������}:��4߉VZ�ܦ�@���o�5'��j%�j�C��H2G;�����t�,yx�C��/��x�۫5J�?�r��Pgy>ߟd�nkx�������Q�V�*8�v�a�rƢ�:=�7}l���6��&��-.��w�"*���T6�բ銁��c=�0�F��ɣ+���œ<;�¶ί|gk��1�/�_ad��D i������xdё+�R���V���H{�?���@bvo�7=�R�f0��i��J
�$��+�K�DaNx����d�Ũ�������h7v`�/�|Jfs}f��jr���R��/����c�6�8-���S^:x8����s�Ε�g�N���:E&	�0��i�H��C�ȻQ�3+���4�6cGӒ�6��$�;�<ɵF���/fK�`G��p�jhg���3r��v�W)���7O����r�И�E&J��w:��o��o3-�%�k��d����m�Z6�P�["��O���|���F�AE���0!0�o�l��J Ǣ���:xAi��lk9�HfO0�:R���my�x8��zn��Ǭ�}���B���WY�QIކ�GxG�%d�=�*��C�r�Tx� W������`0��yA|����̑���G*4�p"��d�l�����3��c>3ѩ�w��<�!	@��.�za
��}?Hrdk�iI�ؖI1OǼ���fZ�� �gs!]�d���NЏ�V��q���i��Eo���h�wƁ�^G�Ǻj�`s܄t�Z�i�*�R��Ə֜����6�_��I��o��bC$�$�£"I��K�m�V��:wU��5� �n���3�3��B痫��T6#Kb3��%� ���A�5��a'�%+Z���B�$���4[�{����O�n�eH���*)K���m^�\�O�w�$�cb�� �����MO�x�>r�!Yq�'<�ζ<-c��8xJGR��ڐ�	zqa�@��,\$�߹�����Lܳh0/ã7C�A���^.�	,��0�m��5l�゘�V�\��^��#��G�����ų|������B��T����N0���l�P�̃W���3�]�Y*F�[<B|������wÛ�,z������@��n�%�h�!+�'+T��[�V��[�7�G��i���a��Ys��J�=_қ�Q����|��]C#��o�YC��j[�>a7���[N��Bwˏ ���!	[��s�c�Ⱥ>7��HAH������߇�����[�~�^͘�l����3�S����\���s�8�� ���X}��X�:���ձAfxxښ�z_�����jf�o�5�2�3�!ՇϏ����	�;����/����K9�_�E�y)�A��������e����B�������l��Y����&�ҟ�F
GR�Z���!��Ա6W��b��ֲ׆���'��T�~�m��z�*-C��ܢ�<B�n���3Ֆ��;N���Efh:�O��'u7czg�U�]�ULBb�X����=����J�8|���7��A\���-�v�e�S����ҁ6ţ����-�n����X�d��$j?�v9�1�����l5je�~94p^B!���5�K�������q��1)=�"�,��f滔��,���IT5���r��j�x�u�+#�[�WyV��n97[X�����k$m�3�h���N�#�lD�y�����w�l�	"٣?D� LC����.�I��kYz����$�=�B71���⮗�75�T�֣�S��>�g����A"�K�����>nɓq���!�@i✤��8�|?�ϿU$D��)G�4��c��i��R���ڡ9_�AL/bH��ګj�O+����F2�i��g���h����XG"�WnU*�v���Dy�#����L0�����JY�>M�-I+K�I�����R���Nj�e�"3��3ӊ�7t��Q�|r�u��J�Vf�2{�S���(��r���`��,q#!�tVK�����=��\����,i��Ԉ���9
���G`j��S�Z��=��}���j�.�R⒭�\��^�g���e���Α����+A(E���a����<T�^M\��%��B}����Ʊ�4�Z��;9�u�kJ�xBM�⯩��	�X�H�O[�H��9w��N�l��x!n� �*	 �ŀ! ��GX�8�0����9N9�E��� 7����A���}��9F1+�@��QE|�J�}9M���N��]�ݛ�����D�o5� �^.\u'C�6�6]Hhq�M���W����[��$�O��-����1)��F���͝��E�t�sG��9�
� _ȵ���=e� v�����3��g�E/Y	K��'�Ҩ��>}A���;W���J�X4{i�0�6�[��2s��a�>Z��́&���1TO��>��1��$�]C	];��6��d�V��m�>���ߔC�_lW�����Ȑ�Nї��~l��u�Y�1�b���\���/��G^��M���Zb�a����oi�y���
�Ȉ7a�i�܍�q͊IG*亁�Z��W��a>͍���L��X<V��޽����&���2�+���l�ND*"q/v �"��oޠУ��8�k��� ��Rx%}�5�;�B��1H7�c5��ԝ��H��b2}�5�chp3(ES�hB_�Y��A��tI�����p�G�Z�CU�+x�5` �` 0~���η#�u���2t�X���!͂�C��^s .>-�eΎ���=����9����{�]�ϔPs(L�;��7���gf[��v��
io��B�#(u�����{���Ҫ_�f �������U�b�ln���;/[����N���S�����H�@����Do5���.U>
�$ʹv7$d�0�:P��6F��b�-N�����8�psV3I^���k�$h��̏� [�� r���q�g]��^��9'2���ܖ|4�{ն~j�CҬ�����L#�X\;x/��!]a�C��?uo�����gj�=������W��	�H%�-l�q< !8d��͓��R`T�Fg�农 ����9yP��ie����C�<!zo),�	��&�I�cM!�>�3�'c�:e���@$`i���AÒ�5��||qT�l��4��/�����Tȍŧ�@f��"�N�	��F_ԚEJ_��	�u����Ue
���ٿϓ c<��5WZ��
p(COq�y�փ��%��dI]�y�)W�m�{:i ��{`׾�8���Zy��Ђ�D	E)Z'�y�č����AUD�v�gH��J��s<���[�B�������!�`���[����94���j�}��[�W��Vz�Ʌd@H���wʉUΨ��Wv��/�yv��0�/�]�u-狳���_�v@�Fz���Y&){e�c!U��"���W"�
��'_e�S��`��v�Z�N߉��1Ȋ[k����4�BXMȜ�����n�Y���-ާ�e�-�'M}��=��R=���r~YEW��5�@���cM�栓�Px��~B����Fc ��#ux���ڕ�M�������g,�u�fb�ݴV,Me����b1����IÚ=o�J��U�P�.<GY���a����\�f���K:'󮹰�N�l{D#���Z(^a!e���&�|�����!9�n�������N޽���ڋ�Z����ӏG��^6%!���p���>(�ۡ����	?Ն�*T��b��]=$�7i����k_�������e	�@�[ �܉���Ӥ�&e�O���_nWEM���8�#ݽ�!o��v[�۴G~xz���Kd!`[���k�E��0����󹆁������P̪Ů-�)CР�Y't���u<m��KU��"����g��X8~�&30?�m�����\1�v��ᖶ�p��%}�$��J�� ��˔�YS�94���Я(3b���9��L���O�8���SuD}Ɛ�q!���V8N6}�>����	���0q���7Y1�����/:�ey�M���࿯B�ى��ɣ@:�N��L��2��L#��mZ���IuD7�)'���a���M����GoM# �j���o"����c�wy�A���ȗ���aƶ�N�-�ې�9rͷ�v����rsL���;	���!�ޞ��g�ބ�n����۶#*-&@\�Nץ�c~�VXd�g�΀g��]H�L7w�������<�%�o�9���w���)�2��gmCһ��|�W�j��A����[����w���c��-(�(zd�d>s p�H���:�Ö}���eQ�;����b&�M��DT���գ�aO>�	c�A�rf����y���/��UTZ<�ƪ��b��f��?"�1똖��W)��v�������d�OdS�[���&>?�K�%c��,4`޼N1��喝dEJfB��.)��Ի��Ks�&K��4��$YK�$��I}.�I�;vx�t;�<D��6���\�1)]T�j�F_��� �O��3�p���:}����@��K���w�x, X�9�L�0�Y���~����nYX��el�S��zm�wm�\�y�dy�u�`�L��w"z|��Fކ����&��?o�'3is���#W�Ѽ\V1�����.K%�!��P��	H�?����8"��������mͪ����9���{e�
�`��o��w^�Xгgtl�n0���2�U)ҍ�����x8�kA@�Y�K�-�)����%m3�&��d�T�P�I�r�Z�5�}񆩨Crt�.�	�Ãl���-�� 3��JG�$�\N�jz���+��Ϡ�������I�^Q��	��R�X��p�+난O�VP�!�2LV/�1?z���Q-v�dzWX?���a܋ �x�\h���P�l���h�j��qv��$=�oi�Aw/-����º,��{=��,~_�w�{�Y�M��>�su����;�M~b��=��刎�_&�$޽���f2�\��EL�/�P,�_�ǗT|d)N֘�fjwי�C{��{Xl~�I�@=�|1wd����?2!LK`���%tG��	�>�Ӈ����z���ԱZ��i�����_P�&��Xlk����(4���*�������n�@�r�*�"��{^��E�������X��dѮL���x���D/₁����w�}P�>Aj Ir���+�u�I����0A��I*�e�M�Z^|X�ˎ)q�o3e-U������a��3^�a�B`������6^D��*}6b��1ҡ���G�^��f9���y5�`s�Va�ע*d�Y�x�=Cwl�l����Y�� �*��J'|&��?�I�����������w�.?c�tAM���`���CH@��Տƌ��XM?� ������r:^ײ���
�|��m;�t��:�ӎ=7@d0����1A�
WwJe I�`_ܨ��Y��"+�lU:?�>���r � ��SK��#�q�i�5ّ2��<�zm�Gԝ^�n,l~�eY�m@Z����X��#���_�L���pK����-ح��J+��( �$c=���T��^���˔݇I�8��\���� ~n�^.D���Z�I��vGz�#av�n&W��IT�#����u1�2�(�g1�'��@axo�%���4e'�b�>P�Hۻ���
��=8h���zo/�6G -�4��lՋL���h�L�(�/�3�\�ߛ0d��Ktl���I�-̓}���{dy��k]�C��`��O(!�<����-Ŭ��d朗R>I�{�]�i1�"a���
����Hq��P֟"W4Ӆ�P��Z`�����6E�~�w�bi����~P�*�[����Boq��*������w[���t�Ra�D�֟yp/;p�n�?�@�HtZ�0V\7p��c-K��޼�ӗh갪�|YPݱ,	�|N1����^(��*�o�F?����x���� Cj`���r؆�/78?	�4�r�B��dH?��0���������RJ�I���0�K��4�}ث����T|�͏h�z+�K�4Z���\`Ҟw��to�<cǩ�2Z�{�P$/j��=m�r� DJefj4eO�)�3������Z���=%gFH��0�s�u��;�Հ�z�i'�I��U�u��Mi"�k`�6`b�AK��"G��ۙpIR����y�c!Ջ!+T�]�/�6�.<OZ�K2cVA,塕ɧĬ"=:g��'����g�ja̋U?�(�}�\��?n9����>�b*�}���Q������%F��Vl�\;��@|�R����ej+�6� ��I��'l�����=�_��,r�C�~�!Z���G��J�`E^�gAr������>�_�!oO	Զ�U���@���.�>�#��q�I,D�����՛��.1�=������������y��L�鑇D�a}���a(^����*)�ď�M�=�v��
/
�O�r��
#̳��(	۷B�����`�S�PN���)34��TY���%,��F3�s�i� �"�{׎#��L{lٲ�M+���7%&�������9�3SI�|�������0�L,l��ź�mo�q/�/5�4�3�QFojƿ�/�-Ⴡ%��P� U���qB���e�h�"8#��^N0Y4"6��UR6o�G�Վ���dTS/����Yv�|�0ʳ�H�L�)ܻ�́G�ǳ��j�6[߶�,�É��L4.ZG�/)B��à�3Qv�#b]�=����?<N&��?�����a�]�ݢP�&*�[��i�xD��jwLj�c,E4�vR>\Ǉ1q��1Prw��1Ә�����]�U��g�V$�O.JÑ����s��=����ީ��FVNSZ��e���e1���`t�4�,�}���cw���/�n��c�
M�a�;*8��<-y;�~���곀����X�ta��آ��S�mfȾ�[ME�[����ef���(�C��̦]�������u���Î)�ck�vM�oө/�єr��v��r��&��?D�	҂�{R�Z��,B��3o�TK���@d`��_�s��br[s��!�&�s�|���\�_w����降0 ̐�p�LFt�`/}\N�����*'c�1a`�ȑ�ݜ�񒩕h�).w}R��:� ���?��N�?�޼?}�d��9S�[Bo�L�?�{�YN���/����?�Mh5&W�%�T���H٨��X���=�۔�6Ύ�#�� Xu!@��Rb�64��]��t������%o�B!���;5�J���9�4+|�(	li7	"׺h^h�O�0�DB'���� �~	������������	�2�!/�/���	���k����/jm��+��� ��j�D�^}d��e=����~���t�b�e�� �(<�.�(qJ
���,�=r|V�t����>z���q��H��V���p��M����$�s�l6I���F�qL����j�.�# �NܗF�=��G�2R�cM&Z�<z�y����)�|�@$��Uq��F���Q=��u��c�M� '��Ө<h�;WGYo���G��tJ3K���;�������O�l�A�&�1pΏLp��S��N�6�Dk�}�%���������m�4XC8j�l�եD��6�/^�����g��E��j]cp����A�T_<Zɹl���h�Q���Q8��� ,�����i6�νmdyZ@�g%jSXk��ŕj[���d��o��0~�QBm�9��U
y��J�9L���0Q$]��6�)_�L\'A}l5M�Q�"h�Kq%T�o�{�aV2�.�8ppD�C
F�խ޼��P���#���L��?əS�l`�щ��}������ ~,*S�;#��<�rKI�;������2q��>{R5�!����!�͕V��%b4=!�o�X/f��X�d+��h�ʽԞ䂲��G��+|�WZl� ��B.�0�O �y|b=�N��}R��2ݧ��ph����Ӳ�Q�cu����1��S��A�^���pD�]:m���Cx��q1p�$0bM�m��]Y�ӭ���4�F[5�g����.��Q����B@ωl·{�?�^���򁽘�Bn�2,��G�V��/��{�7�C���I��L,P'Tz~�6��$�8)E���v$��Kq��B7h4���]-�ǫ
�;��\�d���ͨL&~��S�Q[휬��g`�o
�QMj?��E��mip`�^f��{�o����K��j����٢Ch�p�� ]���\HѬ  t��q�'|�S�fZ��&_��M^}X��� ǡ�i�l�a���k�9��h�E�_�f�W@JS1%�!�(���ظ[SM02�V6�;<��+< (&|�Ŧ7���CλEƽ`�W���Xu�&���0.^�y��)�����t��eĹ��kM�����ޙǚ/�^N�������g�,�������.�5��wZ2�'nc#�Ø�【�w��<�| ����n�y6���(��xi@?��<u_���X*y��"��p�Q��� ��@:�ءQ��j�leߑ�Vcp��&z*�re6��f��˴�l�q<0f�ajM� ������s"�,��7��j����wƑ̲kl������`��Q�3�2�=��*��o3;��6��j�]P��[D�V} ��рG�|���Sp#@�1E�"ѵ8�IDNmݭ�E"}�S����d�>�a���oĐh7�v��Ls����xzQ_�U�u�i�/���P$"7J���_/ 7E�ˑA�f�5+g�%I�ɐ���^�qPNՕ���/!keMLf�t��>�В�򀯫�`���	V\��E����Թ��ծZy�u�ve5�jz�ü:�~�"�AQJo����{��*L��'#��:��Y�=I$���u�_�� �TW�j��\T���%W:~G��'�6=ʻ�l�ei)��K?����S��.]�^α����`�Sݔ�d�[^+��޳�^�e+�Ez*ae?#u:W�+���.g�4��V9D�*���[�Ёr�!-���>;�E�1�z*}��Er��1�_f0H�p�Zd �X�k��H�y�8[�R��./�����F_��ZwD`"(����9���:'E�����pW���o~�Q��o�ɤDǁ$�c�b�.&l�q�(Z�*����ʹ���ԂL)�[�6�9�7�8n��|�s�(�s��*������ϵ�>�)ʺ�$��M9�pȓ��H�Mu8����g�A�v���l2+�]�������NYcj�+m�$C��YkǷ��t2���SgjW貍2���ּ	~E2!I)�ts���� �E��)��Cƺ<s~�a�yIBQOX����$
s��)F���4&�t�K�҂�}�.*���.՟��^Mx��df*"4�vg�h������f|��`���|��r��F����M�Dq�}���r�����!"�H2�����a�]���/��>a�爅�d��	�Do+4;� �>rCʟ�F�86&[��CR����`�?osk�(l�z�����&����PN�j�FmR�<xҜW,w�C��%�;�o
�X��"`%8�����n���������M�;����R|�}�!��s/��B�<��h��}W��,P��,Lq�Ug�ؐ�k�̺Y�Ϣ��µXnlNx������A�h;4�p����b(]�FQH�����'�N��!3�l��Y~* �I�tV]DN���MV��lzk�P�R���Ïe�9,�>���F��y|z]��
���ឭv47+*��Z�a��n�]A����A&�V?����{R�Pᔵ��曥�2�hX��!W:f����DE̶U�WTS}�O(o؆*3lu���cלwTD�-�K����r[B�B��.�,���̱"����-滁D��8Е��`!���`6���h$�1�W,����i�u�mB�\�DU�?��b�=n��t�����?�eE'!~���>II�72�������5{�C��ϊ�SD�2��� 9��ع�D���ءwB��3�/U*���vi@��8�E%S������x9@�::(ΛO�p�6Ԥ�(J̆�M���B3���T,�e\<��0%����7↬���Q�(�ı�v:h��OT/�ۓc��oAf
	q\|�����/�)�l����`��V`(���ʦޑ'�KM6�Vp7y|M���w�QU�J6�ST��p9�r��E}_�E�v�f�?�� j���B�/�xpm��Ǿ*f�C?.`��e͒n����ilAؚ
o*d<1�^ y<"ؘ��-Z�����*u�"�*�`��B��\CURP���pxK�#G_�[h���X�`a"�S�q8��$�8��\�(T2�L!ױ�v��L�V�:�tX¡�M
���%�<W_��tڬ��%g����t,F�0m�4;�#P�E���]�F���X�Y:�Rʨ�7�%t[�3JeЮ��RE�ݲ�c��?ʨ����1m$���~�$�W�	?iu.���靕!O�i��G����_��o�����|��Ͱ$d=��@��D�Ty[e��&��"b�46}�h�H�٥x�/�����Q���8o��^ҦEB��dnh�:l���+�Q��
��`�l����4&'z���I�(�)��Bư��뙎0pk������6���Y����v&C��fB�.TKSӲ�
�C2��� �[tw���q$^�3�ʺ(��sH4�P��qT�;��G�$�t3LG�]���RĻ!�{eX��!ih:4�Ǔ�r}W���/4	S�������`�О?Gj���
���,��b��Z��ʤ
<�a� ���]���}Į���;-�R��V���,ԥ2x��.��A�(Ot���3Gn����+篃V�*M+�F�*��*#����Xزj԰�CJ�p���$0�W��3���m�wAݗ���r����i�Pz���<#�i�xR�8�����M�gxn����j({�&�Ηe�M��g/l�l兀l�˗��"�,�p��"X:m�}Ԁj�y��Ô#z��������^�aJ�
�����+Ky��}R�/#ְ���?�֑�?�g񴕩���J�����d�B�L(��k��r�eOH�K�kj���	�^�e��â�ԈZx�a���L�Ͼ�_b� Nf��a�����)xO�iH:�Ox<����E29I:#��hC,���Zь����9�Q�nb(~��}D/W^��
�H#.ʯ��@�}
9S��<���>!�D�(���vY�����R��y'��K�L��/)rI Tj9�v�zM-Q:���D�� ��R��zڷ��'X鬘#��R�P)(�5:�X��ӂ��N�ź������Ӛ�)��Z.?���vce�{�mmA�n���&ϻa)��= ��& `,X���.����C���/S~��祐�9V��轭�.ȟ5:{��4>��u�����Rּ�W	������Zm��}]�_��2RT�Z�����l��	�bX`W�$�M�;�P�k�,ÕC�`���y׷�V%0ޡ,�Ԍ#�G�����P�S�[vяСK<Ƃ��mȉ$=$�dS�O��S�b����Ԙq�ӵl?���`	�֏��\�L���.�w
y���\o�sdT������4>�R̪X���^��(��(�T��X|v�:�:�-kL��2p���r�K����K�;-ݾ�bU�wΪ��]oq����.b1ϡ��h�=]�?�
�y|�>���?�^�F �Q����?࠳��i������L�Șy������� h"F4n��įc)PF&�����f���6,_�|�6=&��p ��̙c��	~�VP�ߡN�a�@�L������>��Q�m�bMՂ���yp�� �ji������R��M�
'E��S���6puQ���q/��u�2���G5�!��ENW֒�/ujh�G��2����T9�L�٩�x���֏���܃��G��m ���j���� �Rc����N�D�f!�!�Q]Kj���W���mz�,7�u�1D���`a�����)�1D�'�����1�B��`�w��W�<�0!*�1�
rύ�X�Iכ�Ln�XJ#�����^*�L؂6�%[�$�?Y������8V��F�A����a&\��e����xe����.W���B߬����$c�k�BBP�
�_� D�nHp�n�,�#���f�D_�x��G��в%�$s@��^k&'�X�O�So�-��NA����m�|iCIH���Ul�d�A���}����.��ˋ�i~W���zX�{-�̡��Os<��j�0��B�A��
h��\��d�<�u�n�c]��C���trZ08@}�Y�]b���7rya����
U��A%�����˟��Ε�WU��r�yrO�0�AV��azI�������)l�d#��h���V�ԇ)�X25�S܋���/���=�.-�r*��\�a�I��в�Bůg&� ��I{=��}��0�i��Mz���H�s&&����ΰ��}�>؈�ULa���疻F���nܮ�����p��}>�Y�Y�=8xH5$U��u}�J�;(�͒Ĉ�K/[��5e�$�̶1=}�e�������6�Z�Ʉ(2c��s�P��ED߃p(�ӕB5c����}�'l &���e�P��`$��UX��� M^ZDl��o�<�����r����\�H�GY��E��i�`�Q����\߿�|�ԉ��I���v��/26��g��t�����B��B}G�P�OO�v����;�%Xy���w*=����>�k���%���3O\S��)Q_Yy��Ѳ��-��'��c����Olw`v��
}�<��s{l����W�˿ŜH���úG��p�L�5gX%�o$L��;e��Yk`rdc(���KW�zR�(YTTU�84z�`4yPr6��
3��������eĬ����olѥC����Ջ����k݄�ݚ�;������n�P3u(HР	H��J�h��e�[���}K	�e�w�R���z�DW�<�2��7��}����a��p�\��%Ŷm�3�V!*^���n���o^�big"'o�b�Cn���͕�Q� ��Q�k�.������c{�T�#Cgn�w�jO^z��`s����5_^N� 5��m��|����<�%kZr�t�%`����D�����˝�O]A�A��I�ɏk�Q`����\i��t$N�f:���g�j?��Ζ����y&��~}�p����]�ȝY�3]ɩ7�,�x�AR*��d=QUvt�h�cP/
�xQJG�0��8}_EJ�N��+K��g5�9�yk�Z���(I�/']����E>�����?�8ac�a�X�)�gY��5J����2������NX5ؙb���p��˗��ɞ�Zv�#���G�{+�8��PVC�XW��c沀d�t�R���%w��b�]�۹�~%'���
ւU<ܺp.��e8� ���Y�{������rJ�S������v���㹶i��"�Ft�G"=J����,c�'�æ�r;��\�F_GK���x���fw\�v�٫�%�T3�tg�y���p��,�#*W{g���:�i�٣O�Г�ߛ��]~Ciz��l�0��߅�*k�՛��@w;�~Gq���31�=M���d]����1ǋP�$4�f�}��X$,:��j������.��A���j�L�5��p���D�)���ʸQ���"���5��Ƣ�Ν
d��Rb�5������c�2)��
��B!²�E���:e��ӛ\����\^?�"��r ��?x^)R\ڎt,�M��v̕���������$Z4 �bfw:��@ޯL�G6+ﭳ�kPL*�mQ�&�y��W.�6�9�1��$]�	��%S{~j���/�ŷ�w�A�ћ�����3 �K��[�>��z
H~�n�o�m���pE'����`�e) ���]�W9dX��R� ��!d-�'C	f��U�Ud`b��Nx���x���/��0~�K�kV!x�.X��� F<���x{y�CMM�~�!��[K���r�MH��+A��� �7#�N���NR95�]����$�]�6	�z�$�V�){��w
�0��W?��S�tu�c��4��B`<�3��ا1:N��y��/�������垮{H�C��	��[����=���T �:h1��(� 8�H,�~C��{�u�0�i�e��M�M�������� ��2�m��q�zZwDL�n\��j��z��B�,�>.�ɭ��\��6=��U%�ώ�dx�1�_���qn�����T�
Ǔ�)�h���z�(�;c=\c�զ��Aݢ��/����_ic�>���^>�W]O��v�E���>�B�Ց�yP:V�Ɛ�{Xfg���0��:��C5\;�����ψ�d�1V�ܔ//g���x�	����sXf�\/[̒����x�Ճ��I�mKm3'�n���a��C_��I �/\<��2���P��h._������]"�~9pM}��L�,] �C�淙Obg���#�����6���X׼A.��c�N��z�\	.��L5G"*�'�����KŮ�]3����M��}{�ϓ�
7[����j)�!��|�y�F�H�C�AY���-�.���T������^f�^Bh�o�K����Z{�O�v�J�CƕKO�����6�M
f�0Y�2�� k���=��3��Yu8�=�����`�ń8raC���h:&6u!p�~�l�9<��_+TnX91�D��ϓ��<��^g�`�����D�<�v*�k4k�z� �9�	��У"��U�V�����Mw@��0杒���6x�ۣEg�
�HI�Uۣ�@ڞ��GQS��@%����Ƃ��n�u�(�$1P6����v�k��dK���5V8x��8���,�ƃ�]a4G
����Y�5R"n�|^�|*n/�T	�{�@D��\nX�C�_��	�la�r�p7�s�T�B�j�������T��.3=(+�p�;͋�;���Ym9��.��k�&�l�.7���¯�A���� ��_�L��J���� �̳�y xm���8��ܣ��|#�SLg�a)����X�G�S�B�:���׷}[�t��;���I�>�L2��\�)�v���r�k6(���Q+'��
�=Bo����Sb�#���ګ4��.T��=���:�CN
Xa`�$�L�r�c���!�g S��(LO�_�S@�P�Ԅ^{��̩�DzK��K�˩yz���HU<��j�蚹�����-8_·�������M�o���[�?�%���>��3��֐��W8��Ø��=ɇ��׌�8ܬ��PҞ��	�`��&0D=>��X]��%b��cH]Z~��a��F��sH�*=&ʳ�%M�� �B�g�����c�Ek	��>����@MTxi��!�߉CIE,�:��rx���g_�,�7$���kॾ�h ֬+�y�3����q���\�Aп/�$�r�ٛ;���i�b�^ʅ:��;=��
�p@�s>6����)z���EWVf�dbs�j�-��F�,��1<J�pS�z.#�ݷr�9h���G�sᥥR3Yέ�q{TP��Y�u_	lk'φ��ͦ�na��{*�em�~e�mo���'3vޣg��7���ȶ�:���E�p�|��-{��(A���δ��[�ح�T0�P��\J(Bn���
����	������B#�=�(es�Kf狨6��z,��
eQX%�jj�m�9d|�y5x�W�h��"�	3{9��g���i���9��t��w��#����
_b%K��E]ʘ����.�Țގ�dg�� ���g���߼��پX�Ѓ����P�:*�d;I��<���\�Ǌv'5]ԏ���#b�^6}ǵ���ǃ��T́ȑ��n���)�Z�AY�|�i�y< �/�{v�&M&o�n�����~�l�����R���.�{e㯝+'��<&3�ڢǟ\:�?0���S�gKoҷm� w9��c��lK_ �h��c}Y\�}��%´�-h�Qe���5hw���Qig��|H�9�2Y5xQD�����o[8X^�h\�6)�.��e7�Vjɕ�����`�ͽZO�������y~.f�j��، qf�}8P$/W<��x����X�k+3��o˴J���w�gbs��Fv�&R�b��&7�1'��X�4iܻ`!R�"�am�<��G�N�^!:z�ʽS�_ꩁC_AѕM���
�/I>��H1��H�b�Y���F��D���qL3�2ܿ��k��S�T\��eq�0�C��c �+��.2�b)���q7Ȫln9L�6�קE�	->s��q���1�a;��w�E���C̿̇'FTGG��?��	#WCy��@���@��D}�� �GY��̻�,�vE�U0��q�u4�)�I��!ߛ��=
�M��K��V>1n�d+l�Yݺ��1��-�y��o��62�M�D��QfQʅ��G-�˲�V��Ȭ#<���!\QO�?8&bqG�Z!���q����>�m��aP�3����aÓ6�E�b���,)$�f#l�t�]$b֚x����΁��)l#�A@m����v���g00�<�����4\�4Iؖ�O�mFp!Ō�"�G��w��?��cg~m�v�������G�?�85q��y��pm�q/��s�Z,M�\Ʉ����c�c�Q~Ȼ.;g��S�d��Ta�u]UX�%����)��z�2촄�^AbE�_-���Vg�s��j�1�q���u�A����(���`s��߯��cfj�tV��nj��ܧ�N�;s�����S�m��}75���W����3����'^����h��bOM=�@���=��<����F��;^��5���@%:"��뽅{K�Ӭ�ubt*�]�+����Zx���P�j�vz?E(����Ѕ�$~�����Tn+g�=����4\�w��'�j�&�"���D��"�r_��M�BtTM`�

�U2��Rt,��S�VK9i+W5�����G�o����\y�o�M[����ܰ�4�� ps�a�MyL�0�����>� J���U���ힳ���{I^le\��_��H���|0��A}rt_��k�/�(�+qG�f���TƳ�]K���~ܡ* �}�]2��.��د~6��w9��sn�;��˓ҥ^����	 �YbmQ�`sQ
�!��pN�8Azl578���`��A����ƿ��G#�*e��m�E����d�LD�pjb�CW��E՗8���Ս�c���ȟ��G�|N�*���ƍz*J�4���y����т�����$��X�}�P���Ҷ�b���*�R�L =3&@H�wt�Ǳs�ս�@�Y�p��{�Y��,���U<,#.�;%��:���k�"����8b,_<�������c��co��^�l��;U���Լ;)����,q>WQ��'���o
f�ډ׉j����C�+1(g`�B��/�q_��M�(��=�����3���>��d�S}��y�d��"F���3r,8H`U ��+p���}���� �/e�:��?���s�M��w?'��Y�Z�����*
T�e%}��hU�^�2�'Od�=�#�y�]T+�7W�`�[�JK��8�����ʖ����%A��,���$^�`fʢz�&EJ�㺴���!.�8Օ���YgbU#�����ԫ�I2�[I�JU�����&���wb����{ �iy��� ��f���#���{��+D�5��У=5K���.��8�8Q�)0�������8�?Dh��YɊ
V 4��O6�0/B�s���j�^�2���\Y7��Z0���H�� j '�ؒ?b��{`�GN�H�]W�9��B!�+"$�N�*�{Ε?����B/*`fɔ.YOw7]�WY�
��j���k�S�#.����O����N�������=8{���	���с�,�0��m��:������URF�4�z#t�*)��?g���:��N��:��/Q��L��ҒG�E-N渏��U�[@��c�w�BX�~��
~�6���~�7�x�OvLF�?1�};4���k����F�%t����Sk�P-�J?�����m�J��ce��gT�&v
��ng����O���w�$�����]0`2=<���Մi�1��b�`���Ë&¿#��!i�}�c��H ׺ć��M�2�'���)��8B'�Y�u��y�<j)��M^Pjv5"�2W����fD�b/j�8!C�}����yhg�s8��c����8��lw��B5�@�+:֏?z��_���3\8f��Co{�,�����1�ke��.�̥t��v'�ԧt��/& FFR��%���ǦO��{_�P2ʝ���m�w`W�{�WT`�L��������Ho�4U?�7��d�؂9L��(����_� \����jR6t�v C!�:�����~�Y9�w�������ioy�2fX^�rV�G�FPM�;Hf5;i�K������'}:`��R׭}��O��$�R
��n����g���:(��4?Y��g�q*s�
1��6f3���G��Lht�*	�~��{�����Ɋ	���i�*�ޙ��-Wf}@i烺��S���E����g5�U=��,I�4��9'��u��.i*F7ִGL鄹�PFK�ڈ'LǠhs��ZE���	\>�:& �X�E���/vt&^�qQ�Hz-����u��)��d�������#���>�"�3U�?B�6t���>�y�5�ž�U�է:]�I�Mr���/L����KM �h4=V?�Z,Q|y�a������P̕�pޟ����,����kMʽV�����uOW{��`i��|~�)���uq��-7Uk,^���{H��d�tɗ�2p��SSsiD�}U�Ut�		 ���-ĺ-�62p�72���Qi��c�r�mk��g�Je��j:��b6)I+�ʭ�-����&���A�%�A�6�w�+�A�-`'�䗫�6��3��/���,��L�Wddj?���'�� ���)����ȅ�W�'��d�%���"�͋��d�����@Nu�Ŵ7Z�u����Q�R�1�`���s�Z+�nK<@�l<�_���B޻�q���ڦ2��������[T-HM�R��'v�=�'�C���ܲ���e�GS;>�h�#d�Ǻ-�ȡS+͞^z�y7D��#K�k�?�A��,� �1�"�< ���0�S)巅��������lk�k}�m�\�U� s&m������+S��Lg�4�M�F�+�/]�s��<��d���� t�]F2r���V��fse	�[q�k��n���<:k�����{�'V�߰��!x������xpA�:>ƗϾ��t3%A|N�9�#�SP	���\4C�Be�\�H��T�#�+c�֖+�Z�A�N���������}U�|1����[Hۜo@�u��������$)R�T�Ǯ�Y�� �Ε��<)=�;�N�qA���Q�2�Uq:�\�y(_�$/����Cn4����e<�ȳ��x�ԼI����\�Q��%qHUB�N��;���d�m�^gm��U�����g�����~�N��U������z�B�M�HG�鎣*Z�
�f+�K���� ��P,u�$���H�~�4�.���|���R+S*3oOʛ�4Czc�pVe�(ʅ<���>7�D�l����e�E3L'��*L�;*[}߁�Q>�T.ں&)6|\���,��� Э��]�P�D�r�`hI�_����`���A��E�H��7{Pn�/�\J��[\�cl�m�0�pP���.�&Ot7�����Qni<}Yն� ��R=��S��pĝ���0QZ��F8�Qy&��y�x�~����<�p��~@q�����)�DMWU����F�>!�I����x\�lؔ�h:a��++$Y�R[b!B�����Eg@�5r2���p����~��٫��8n�λ
D��Q|ɱS΅����\������%<�G�u���I����l���B��9���%}��2ٛ��U��Pnq��#� p��d�U3��:[�t*�����Y��[�5S�=
��rn��z�/��z��䓈=\������JE���(�h(Д���j���3���V����-�_�X�m��,�h�+�����;l����-�D��$�����n�d�9??Ԥj):R����x������Ѽ�qϩ ׽��Z����Ź��Fȭ;�RF(4Ku�����޶����.��YС�n������fQ�U$uC뎭SL��S�����κ�
t�d(��*K.�T�rv'`�G�_	N�k磢î����ud�a��cn�g��&}��o�㏙9A5�Ih�J%�gm�y��C��O�������PT��:a����U(�n�<�I����NE�+�+Q�O�|���z,�[ˡ���Vם/^ҢֺH[h0��pNR�
rl/��xG�.@m���Dp8�2eږԣ�K��be������pG�\j�5d�qkȧ�f/�C�=�%S$:.��A��Lk�}��s��{�z�Ҟ�e嶦�M3#@���҃W����S�UJ(Uh�t�,��E�6W��xA�-M�.z�5^����z��_x /�kDT�!�ư�15<O_�H��FT���e�H
"f �1 �j�_N�I^�Й���)�n�aT��V�e��.��u�0�p����<�-�6o0b���	ˤ�K���J�)]k��09�0��>��/��U����3>e?H;�:���fs�0���w^2�H[�E����KazT�
OM�.W����[T.`����.B6�)�뜓�:V��i�w=p��@ʹ���m�cZ�>�6���jWne 7Vj��^H"��:�P/#w�;%|���1.�;m���'Sl�p��wvE��aO&�f]�����UYg�W������HJ{�T�2� �J��'�� ��]���Շ�E���K�IU�:�b�K/(B@_ʓe�d�5����C�#�i��8� �wLD蹈p��h�%+2�W�mD��N����gtowe����o���j��W�C3�%<< ��ߣ���w�7��ͽt#oQsLQ���0��+��у\ot�UM)�M�+���%䆐��{�&���Y��rL�k,�o���T'�S3M������P}+�.�o�	6�0<ޓ[���B�Dһ����~��>����/Z�n-v��>,��(�yG 6y��F�G��k1���žp�����8�G�-<�3�� �A]n�d�5b��u)��3!R:1��쒗���G|٣�?`P�7��:�y�L� �zP�v��o�����-�ir��:n��ϑԷA�$;?E˒7ښ� ������ո���R"%��9��魃j(�� ��q��D8��2� @��K��N����=n?����H�8���&����R�v�:9�V���ӓ��,��Qnm�.׏�`T���Xu*:y��_I�ZE����\��~O��AV��g�ޢ�6�b�qGߘG�'d��;�rМ �u��!���#�\����Z3Нmm�����1��Wk�5p�q�OK	r�L'�)X���ɷu�&æ�O�m�ĕ�j�o�}�Iꍸr��D>\��M��Aј��E2��N}D$�LRڴ�rL�,�h�gȀ"i�������e��R��@c@+0e�|�����e�h2=l����A�����)��fI�7,l"J��
+}e�Z��������)��A��u�����X�q�V[��!�:w'&u�}y{v��Hhj�D����io��b�Ɨ�C�ޮM3�6R+����g3'��H�..^�UA	`���i2yr��Tq|P�L]�����~��z�z�DɅj�^�؝%C��4��O��]�`K�u���R/�R��k��SC̽,��,͛8� ���]=;��?w6�s��}A��6��WA�~fɏ1���I�'�T ��ܡT��C76L������(|�irj����ߝ܌)��{����E�8�iB�k�RO��@���;Ht��� /𲘊͈���X���|-j����s�\rl����3y����հ�TÏ����J�7#����#���*�	�}��
�}���`��� H��pKw�l�����P��]�f@��g^l�M�?�������n�? ��A�"�v3[e�
m����/�,7G=��Q�f��4�u���^���_��9' E��1;��M�5�)�� �$���r ���rkb��I}P��%T�@�<��z^�Z�~�Q�M���ɧW���犚,�U@X)C�%]RI�nI7F?*�7��XZ��%u
�̄X��X�����B�q��#5]�ӹ�����]T�ذ�*�l�Xl"!�V�y~�!�R��_r�͘�UTr�P�A6$�����"{������R&'�3�f��P?�~�Y��ʨ	h��09j���|#.S�`���f� ���HL-�o�am��N��3��0DF� ��2Bt���+R�L��/���b�o	N�08������_ze���)%cG��	p���Ld�W�m4<�7���0�؁wԮ���dJ���q5�).	ņ�Z�ҡ��澤�4��u�~vEW��9{�gQs���"���+F��:r�����o��8N��6FFDM�ˌ�sFNKɻ��"���ױ9.�R�eWƢ�U���X������
��N���U�J�տ�9
��
n��?^�!�.���x�C��A�R�:�}A�~�"6����yq��'o����z� BBjXy'��/)L ��諒�PA׎�+��n�Z(�F�}� 
">q�1m-펁����v_L��8��7;���$��K��L�0:
�����;��b�+�j�B��$ÿ)�����68�6��&޴��A*B�M��w���P��;�w���S�^×a�Î����u=)�e2��lI�Q�˕S����5�h/�".@�Z:���l��ͮ3�$_dV�\�=X�-%�T+��M����	jL�h��'9�Ҩ��!IP�ˢwRرKվ���-�(ѨC
w*Q��R��ϊ�/�~iG�(�"�^�vl��� 3��9�Yz�J��ݨ� 8�_�����A�C%�x=O����Ae?�ܤ<��Z��J�ɗ��Z�H����D����ڎ�&�xI�B�-�;?��zKY���tƀ���#����/����i�I����x.����J�bx��Ь��a�k�Q���Ey�ܼm��X&���B�!n/���"��8�O,��R�x�_��$p�#���y.͗X7���l����4����]XO�
�gA{T2}zF�\��;��~�0�=d��ԃ�C�F�jy�8#��=S���P�!ִ��~��3�,B�y�Bp�V��̣3��%����Oe�T���l�1L`��G�u��W�i.w<�Q(�k�<[

 �	���̛z����WZ��B�V5"����):O9��G�ɕ?T2���k�#�|EP,)��y��g�vH.M�~�(��%����>}f��c�i��B1���"���Q��#�Ha�0�w�_#C
uRή�i���26]F�JK��$�wXAo��ls���D�y�9���0�4$cu.�P>��]��a�q{�Cg�&�"��&{� ��)���3s[�����ŝ�a��z'�X!gq�G�`:�A�H��'��*~�@�'�3d?;���
�-�g}#���e!����Cwq��P!O��2��pH��+�J�;�u�6�_�I�D�"���U��e������Hc��4s�/TF�LfC|��ypC�0AN��?RO<��i�Z�b��V踠1����MB��+!"gsr�����M�k�?1���ȉ�����:�D�|Z�D�7���D��� #]�a_4[g��IvP+��G�F��a�hd�'���'��%#z��M<o#��,���eo��@I� �ȏ*6�i��t��Ȕ�I4�Ƶ7��u�;<*bT�������&�/��v��<�K�}�6�u�i�eT.��o5��v(:v���L�.��V��is��~��Q�������Y��]�7�8��[�5u(vdW���Mk�O�(y��gN�K���NmTg�
#w�6���J��̒{yg�XO��)z�+�-5�H�kR���í��̇v�t·hzd��W�^B�q��,�\���!�:��"��,���Z��B�J{_��w��gZ>�$����f����+�O��K����^�1�,C7ӥ����ڳ���)����mqS["Xi����;@��_Z���2˶���q��$9|�$s�=���Z�|w%���h���}3��"�����n��!��Z��g+7;�0�w�~�u���ƙ�m ���>1���I�!wZ�[����̰��l�DZ%o���H�;��4��<���Y$��3!��O��Ȋ�$]=u� ��?)/�5=�)��r�1��>Z����K�u S@�D�z�+迪��Q?�h�w� �������\o�;�:u��&[r[C��R�E��H�6���FG� g��[���V��o�Q��'ڝ�5���C�W�ЈEPl�9y%1\���ϖo�@Y����ȁ�F���c�c��
b��e�!�j��iM�B���"J����ԪN�{T8%��z��vݒ����i5h�2�.���;�y\�7��|k�!��&A!��d̈́�
�*��
����-��ǯو��!�9�����\��*�[�j��vP[@�+�4`��0��~�>R��&G��ܫ�o�ء����ٞh8E���}Ȧ�A�x?	�e�D��M���sX��2�\y����Q�lq�;s���0������T������*F �_-S]����'S	�E�&ˣ��mE��i�Ǩ+�
�`G�S�4u�@��*�����u�Rc��Ǔh�!w�K���t�Lh%��?��
L�Г#��n��!7AbE�X��`	B��@���9c_��PO.��y�'�H��n8�w}�ê��rF��W���EIi����t6�	c0���J2��W�-8�g��_)�GIQ�{0�IN:B�������,��U��` ]J&������k %��RЌpksZ�⤻%�������l��9<Qt����Q\s������ �y� ��Z���	�����o�U�`M���*��F��^��aU�i6:1�5岚����R1H�nq���r �b��ڍq��SK��,M"� ~a9Y+�0��̩H�ƥ<v�q�%ʙ�ʩǩLy٫ύI>�L>���;��"�}V��j�j�Z��t%_S�:^��.��\��$���a�T�,���w�,��Yư�~s������$�xof�րR��QU�\KJ����`O�]xk�]��u�^�G~�ѭk�$��و��ן,(��_�, �*,����}�XN�˔Ob���G��S)��f��� 9��]��'��p9Y��V7�Dd+P��_�`Z���Ъ|B͑$�u�4k4��:�n���G��|=AY��d���tL�#�Q���J����;ڇ�;�2��9
���Ň>)�rOx�ԣ�6'��f��Od�t�8EH��D��l)	�vIB�`ߐ@��]�&eQM'�`(��@wa鯜��w0h���{GJ��j�-�$�ܱ�7��k�D,�r��
��0c�#IO�O��C��j�$������ �lu ��~g0?�1'��Wb�ƢE�E�I�#�ǯ�.C2wM=d�m}�L%��YM�L��r�1������UCY�����.?�����|��E�	�0���nl��k�X �ں5iI?�T3Vo�B���D�߷����s'�䗔�5q�n3Qe/�>Qүl��M]1xYd���Mp���0d��#
l�5̬E��LJ\WU% ���p20@���H!%��@������������3�C�$��Zy)���0!B)��{�����H���p�ʥ&"	]�w�p�d{|tz��)� ��;�MN��R����o��H5$0���Q㵁��T���5p��FϹe��x��:�T��nʚzQ�|4W�2�MLN��)aM�uF$%����!�B�m�E���v.�Q��Z�r�ϖ����#���**G��S��c �,I��r���8�׭.
�6��ލ£�DT&Jƒd�dCKW�$a�خ!�����%-%�V��:��_^�@�౐K���uO�C��t�B���V\�)��Ha���`��#�Se-���_�\���h�ƫ�g�{�06K􊖋!�R������U�U�<__��`����} #��I�
��ڞg�Yח��U���N}���-�!��(%����;���GJQB�	�07��d�ncEJ!s��Jڀb�[J��Y>�AD}Z�b%Gً�D���LQwMV�����k�����e���j��w,j�����z�%����F�2��w�v(G���Ѫz�n��_�Iک��Q��;��h0�kw�y�����܁t�;|�E}`X�Q�^��6��#�b0N۷cJ����\^�-Η6��b=O�)�Y�;x326&6�O��JJ��N� ��p��
��ΛjB; s�=]��燅��[���i����]���U��P=N��o��W�3�%�i���I��43���'o*�_|춑�[�HJ�O<���9$臕���O��`�J�K2���]ٞ�	�ڭ�3�ʂ�����h�1�V�iB�>�u������l�I�^�@ȇ�����ɣ;LD�-K�u}0Ei,O2\V��4�[A���uXdi�K�*ס�Z�xΙ9Ɋ,������B�ss�^3���*��t�����1�#���v�W��Pm�0�Me7�i m 9�)�]��3��B�׹df{�:���<)6����l��Y͓�C�#ah/��fF����1�ôa�@y��5�4�*��.�'�0�5�V���ja��m�g��{:� �/�u�!BR.�XL�=�Qc?,r�mrn����Nc��X{@���(��? Ps���.��KPʆo���%嘗�������>�.l}sb�\8�_rd�R1lM��%9�_}5�w��_��(�� h�yE������h�"�V���4 �_�9#�ѿ4b$^���3Zp�D�Կr��6�����ƪr/vk�y����tY��/}���`�%�a����&�Fl�^$����<�k�P�=�V�~��vdOW��աQ�xilNDw�z��w�:���z�0=$�c�fx�1�Ƨ���ŋ��=%'���w�J+�ԓw#_#6�sq������@J¹�y���׋ c$ݡ����H�H� �!�Z��Y��g�\�8��������#�1��V����<3;z�S�����	<�M������&m)���#x���S��l���@ߕ��\�,�)F.z�_��� ��^�����AFT�M��`�G�J�?(��(���Zi� ڝ�W2��C��O:fU|DlA{�^7�=�1w�/@�^���n̹�'���%Ϙ�gb�@�Q=��x9奺(�M�{��_�%���m�]	���S� ���w���ZRE��G2l�VQ��+��&�H4:qm�����A��e�K2�z�U6��8���J��2�n�5F%\�\������r���n��4��ma��SF7wf��#*,��y�	ܰ��Ӻ~NF�S��{��B��W�U�)LDօ~�L�E~?[t�T�W3��
��˺��yԃ���X�����_��ݓ��sa�G�� �H� U�tԱ;�0Ok#}�xD���u��p�`�g���*r�W\d:�����}'N�)�Γ�|��#=�W�����x���X(�Z7���l:���BJ�F��i�@��A��9��C���?d�N3w�"aw��
�MB���g-N췯�\ӌ�{���=z�4��jS�
�˒H�.�5)t�跕q	/S�y��D���"�LÙ�1c��)�#�'o�+
.$�;�n��g�i=�$<��B�+�>�.��车�+�����z�40�b�ú}����O���=�O�����e�`�n���'��ZK�Ux���WV�h�?�
Q��s�^~RJ��;Fwj1,,��_�7q *E�_�ҊB���{��,��ΜY�E��>�t�)țe�
��Yy����a��A��?��&�Sa5�ss!��<�h�sf\n7;�5��A��}�TmtW�8й�wtV�t�P�%RN-O�5KJ޴ӫ���c4�B�x1�}����L��m�`-S���BΑ�}71����T��n\�>�^�v"ߺ���M]ٓ���_��`Ҋ}���ӟ%�V<ո��9u��R��v�\������il���GA��ߛ�ݎ*�˓kQ�aBB����'_����@�6"��o���N,U1���֎��rD0}Ȅ�*wW��ժY�Y��mʿ�p���B����2[��u��^]�|�a�=�u���q���u��@�y|z{n3�]�G6�J�T�@D7T�M��� ��`h��TQ��O-=n����BH���e/��Y�"F*��*@�|`����n��s����ei8,;	����`B�t�ZK��� ?◅��,��(^����x'��đQ^:3�q����>{��p!�%��5p�r��56{
�To����Ŏ3%���}�K*�C#E���s)Ξ����&*�A9���p�}�`�����U�)8�0��*�e�����![�7>�Tw�g"|Y��!��
��C�#��o�* ���
�Qb��V�YP��c�u֛�D� �	�m׈�3e{��`.yǨtm��k�C�|_C��a^�'��O�G��6`˼n|�5�b^�Vf�����n�s���~={�Kʭw#_Zz��>Zg���%w�����m���{tn_��1�-(~��5rkr׽�%D�) ����}��net0-�hTx���G-���]���J��\9\J�ae�r�[?7ֻe�3�	(����s�GaAu�w,PI��ś�Mg}�UR��d���W��v�ԓ� �Z,K�"���%��d��o뇼DM�3B:x��������^�� �Wjb�@0]�_Q��m���C�\K׵G��M�Hh��1"����A5B56\8G1R�,_$��0�R����Y��h��F�vx�I���2�^�NP����Тþ�,�H�<��w5�e�Ԣ�i`�)8g�I��0)�Zͦ��b$��_�eO�Z�V�[�B�Dh�)#�|��[{��	4�N��S=j��![wet�e�s[AĻ�*V ��@��oЉ"t׆�*�\*� �H���a��)RBT�E��N�vJ�wb�8�dGq�<hUY�W��/��
�&���O�w:����: r�U�"f�a�x���?�A�ڛ��m��3Ŋ�v%�)��hU+]���}��:�p@�Uc�P�X����F_�|�Ajf���g�ɼec6� �_��H�:�p��ͭ�;r{�tL�=D���Ȏ#N��f]w�gJ�',��o3'����Z9S5�0��*ҌV�f���5&�4�lrG���q��׋�lln-B��a��t�*?�_��L<ۨ�06�E�	SM.�Q'�愡��qā�7!��Q�ډ��§��8����T���?���U�¢���RC�xG.��{;}�h�t��-��q>�2�V�`�t���Nq����6�<R(�?	����H+����)��w�'N����t� _jS���h=�,��O�	a
P��f���DRt�C�a�y�%B^�<�˺������Mr�Sa�mZnjE�3�}��_�A��G��7�ث�-;�«t��ڎ�:4��+f���N1>�-����7z�a�ΐ� �؎bb��bCI�݊H�Џs��?6�f6��{`�.]U��YI���p7J�zq��)��o?��w�Vʮ$�J�kl����� �X��v�BP'��R��|l5�߼��C��1�b�d���o��:������sǐy�8�(���n(��
�]0iyԩ2�ɜ�����T��"{���id��
���<;D܀�?;�ݦ�!hd���$�J��C��v('T�R|(�l���&"'����޻��ku�%Us)�s��3�ج�����"��7�P"тy����vZoꠦ�=?nH9?	�n�"�'��p�����	�>V��p��F+�y���|�b�
�ù-=����&�SӃd+rU��:���x>����~@�2�:����-mg;����/L'��=�b"<����7�{ӳ\�Y��j�t���F��1�k����idJ+��D�j������5f���[>�D�Lj�i���Z]�rW�H3�Z!h6BN}� e������cҰ�>D3_A�l�� ����7H+,��-�`�F�ٞ L����G�E�\�� ՞ڄG�<Khd�2@4���?���S�Ҏ5�#���G^�:�?-@��m����]qP����lX���U�I"Q@:�E�E[N1�FROG�F��6o�'�v̚�訽�� Ј����{='�k�/�a��}F�g�$�h�xN�;)-�,u!!�M�$?e6%HN_k�D��hI�dsԓ�'ԑ���w����h�X�h�n��-�L%OSO�-z�i�����I�-\�E���J�q�ޓ��[W�|��4Hl��_�O��V��ԩ��C2�UDG,>�Ϟ]s$�l)c�����_���{�@"{�����3f5)�	�ډ/�W*]kj��5�"���̗��743����!{���N��� R��w��M�6���t���\������g���Zs;����.�]Ak
� ~�r���P4N,����2R̞7��Ʀ�بS��I���YC��D�����}P���ح<����b"y1�c��!�ν�],Ax8��2���~�������ir��pD��u��󱻴��'�-�1˫��\>�d��iO'�W�Q5��W�e�caV)gl#Q�:��E(qG�AMӳΏ�|��������'�����ʧ��4�"Y��tH?d��ø�̄!Sg�a�^ڹ<����k9�q�8ou���`����*�W�|����e��B�#��� j��@����K��W�׳�J���U�j5�s
a{�y�0@���g�"\S�{�$��xL�&W"Ow��\��Q��>j8F��᳈��(�p��A���6Hɶ�l�V�46�5[�WLC����6lM�k�P��Af�*��c�q�փ'����
a���f�1��S�4+9���CQ���`�o6����]\�R�>�B�)���E)��,�'զA�-�|c,��X���l�!���i�`�)�v�m���j���q�90+��궳��SuC��?���|ö�z��{,S�7�B�[Ӫ�f�\[�Y���,n�#U{G�qO�}~���ò��K��>( ��V��jUɳ܁!���`������-(�"�w�./O@����8�oarC�J�����~t���1�*���X�Nʱ�Ӄ��WnE sL�vHq��+�q�����o�Q���Ua�5��P`��"�[ܦ�n���eb�w%���[�m����`����mX3���hF�����g����WݿB��dO3���)Z9έ_��a��gU��b~�/���~��>ds���v��7R�L.�v�k�+g����黷�}r��`��U@R����Ƈ�^?pV/��DuL�V��� ���Ϥ����3���	�y����,Gh�i( ��9�R���5�J�%� N^�!�eU���"�����s1^,` `񂡤l=e�� lY�J�j���z�G�Q�G�( �T/&�i=�r4Q�%|>S��#�_q eh�ܓ��i����6��"��~�4�I��ˆ�3��i��`�[!ٖ�p��NY���-��\*x��W�ڋ4��;%����$�z3�	�����i!�Vc�B�n��"�t����Ő��D>g^Ru�ou��ף9k0�\Aʷ~�n0a}���n�^�zw��k�p�;�F��΋����@_�!1A�B6��<�:�k����(�G��d[D�W�_��[�A���A�K�XLk����2oO�K�����kE<��,/�>��y^Oh�m�����u\?�#Ӎ2�<T�b�G�%~x��.���\��G6�:9�&w]���NRj��>�^'��U�&�͈q�[Z�k	���Gs-&�;���Fk�4���&ԓ�����gS�������q!�5x}����٢
�t�D��uѼ�\ o-�ek��e�2Q[�Y�r*�:���]IÜ����`S2�Mv,�*����{MY��i��mf-'�z����J;WX���퍒*�,$e[#����D�]�I�n{<�sX2�����GQ��u��8����7'�DZ�:�z�i�w*�h�`
�W��Gu�+��{�/HX���L�f�T��N�X���3�;NF�����\܆��j��+d��B8�}]�|�����u�R �.����"Z�����E?���܍,�ݙ�g��v�׿\���:��9�֞@�<�J����� ��Ќ��Β�E��MJ:��ŦU�P�� +A����˹.����7��cQ�ACHP{�"��=�=4�-��@��4o3H��<+
��G6�c�/;>��G�t}�i"��wN7�q C��Tb��;7�D_�.�|f�Ô�r�>(�QA�����$"��)�ڬ�y۷y���f�8����DXG�\b�Gts�����d��E-D.
[�Azj���_qa�	��]�[�(y�NpHdW0�n�c��G��b3:#�׭��3fZ_�τ�6��k�=�LpZ"�dL��[�1{���jm�H>�"`�C����r�5�+7�n��Y�d���0h>���k�"ނ&Y]-���ܖi�D����j�l��"+(��޾��B�2�j�/����FX� ��Ytj.-8B���,IrF�?I?�؈	���&�n?J�헀X>�Z��m��zh��y�䄕m]+-
H_W�4�)7^�h7��`����d>f �����Zȍ.E���I�m�^n'�W�����-��b�^X溇��N�/*8n%��E~/�\�����R�Y`l��fE&�p�ቺ�q�jg���t��Wज�;Mq
��\������S��yJ�z���A�ݤ��0d�<p��V�=�ܛ~DψHG��6�nM�o
�#sMbX�!f�7Ο���m��b��A\̷��9�E�8q�i}I��
�D�0#7�aq�A�w*�rț!+4l���A;��O���)�!�䗓ߕ��Je;s.5s5���Gw`v��̞�{���5�N���-�,YH,9�}
]Z�z�Bgt�3o���
ఖIO`V�E�%?��=�,�pA�""�<�/ӥ������W�/��n
f��#y>�ۃ�$�_� ��aa������Nr�N:�Pt�ԕb`/��22Q�-oZ �ޙ�.ͱ��d)��ͼ�uK�C����G}?-=�҆*������8"�gӯ����P�&l��l�z�22ʩ��/� �҈Z���+U��=y[�6~s7*k�Iv���6����B�v�Ա���8���PN	�ާ��h2��
�������iv4�sί&Y(��8��lŀ؃����E�@�9�y�̯q�����+�w�Pt�(��Bş�ӕD�o{�/��|���Q�9.������������&����Te�1��\��i�b�</a��p��N�28����/����&ܖ��S1A��P�Cd������Cu�G�E�Uu�v�L�w����lo���)�3�濥u3����s�`�S����`�����)A�TA�uh�#�"]�s���KzU*#C�soU�3�b
�X~5�Bn�f�n$EN�ͧ�'�N�85��s����>MA�c참$A��&�}�2����X�ݛBE(�~�_R"q�	��m �`��9M.z13��ى$��S�[�f?��}C9T% ��tO�G=��w�4n��bi�O.
^�n�П=���=�b⢔��ݧ���w�_��Zq���Ϡn�=��b���e��#HE�����P{ǂջ߀�H-��M��	��kn��b�A!a� t�1����^)��V6���FHb�wS���C��T*���)Е�����^�+�?Sl�hs�UxD:��}�I�C���9�{��s93~oQ]֐�I�%�!;�]�VZ~8Y�d@�T�A=��F��v���� m~�\�?���FHK&���5?��1�0�����_!��C�O�`1�<<)sA���XEX �q �o�����x%��ô�9�eZ��@kp_�j� [���U���w(���4�Z�-�u	B�1Z�\5�u��#y�?���GU>X���Y=�+ab�g�P}��SBl6���k��EY�iղQE )���V)�S�t.����7��G7�?8�Q�4xX�_�O��
Ab�ԜŲ`t˚eCt�Թ���Zi�W`�S�ߘ�ū3a��c�/��ϣE}��!�y�Ȟ|�]�>�t�.DY��Nw��2x*:3K��2�Q��B��������v2�.��.>ώ+4:Jj-ݠ$�����,������ *�@;T^�o��۾�n���V�]�EvG÷�����H%a�,��H���fB�W�x�q����ً#�R�L����{]7%[Fy*�!(W�A\���k�8���˔s�w�8���=|gRk����aqՔ�_��N+�^��.c��JV�tO��n*��B<-	�����};,fE'/mN#�pem��@��dl�'����FsG ��=�Ƙ|�����ӹ0�t��Xa�r���u��4��k�\��*�c*)<K0m:�))��\��1	��zF���g�d+;�|qd��N�`�08nw{���Bd��=��̕�����ܣ*S����S���%y�JaB+�
��Ya���
��01`��
�Pk���G��tCOձ2/	�����N� �r��r��Oϔ�b���M����M��\���=�M�L#.�n������p��\Fҟ�ƥ����|O��Q%�oMz7�P
��|Kl1�Q2vզS��p��I�iB���?H�P�hH8�'�5 ��� �3�ˊw'�A��`H��/>�����X��On�j�wZ�'"�q?�Z��ĊKY�U��nJ��_��Pb�F���=�E�PJ�$+v>��-l��\
n��w5=��p�m:o,Eux,�����ᇖAN�t�����"9��nJ�nH��6-�;L��%�*��28�=��&���{Ī=���d�[��^.�5d��ऻ��l�Tg��[�8��o��P�E{���aǭ����Iv�	�r��`���ġ�:zx��rg8��5���%�)��,7d��Ă��,��t����<iWy��닸믥z���
�1@,����^��0�R����`�;۽5�]f�����-�&���D/�����k<Msx#�m=�W� nK���+��0�R�g$��Yg�l3�K[�L�����\�f(��/��5�5z<���~#�_�޼,�j���o2�Њ	�<���R��7Vώ�^�������x�M�⣫����3�,�猑/'%U�<���M*�5R���^�a$������0xAn.�_������L�T8��e`�g<p;�_�~��*��cm���=��u`-�H�S��1��	�{�S�c�A.�'�@�r�5'g�G;�W�S"|�!����^�����V��e��ޮ�#��xk?�\̼Y/vY_�{���,S��|43��H��L�m�G��D����¼�g-e�$�J��ѱ�%{V����u6��f$OԌEx�,k�<�ׄ��_w�E"ۿ�C���w�'�!���	����b�("�FJ�ԆH�r"r]��L�n���).���ԋ�nA)����3oc�Ƅ�D{;���
�����\i0&|�$�e>�2g�L�SH��R���5���h ��� >�1A^x���|g��]�����Ú�8�%c�e&���F�����ݜ��&L2���̇sŐ0�֞�q�o��%�Z�B�xt
%_�8��)̷~+�iS��q����w'E�!*(�R�n�B�ˀگ+<�"�j�f�vUG;3�8ذ�'�B�/���W�j����������EI æFg��
�o������C�.�q��k�*�]V�K�|�s9]�UN=��'���/�c�G�(`,�� �V�l�1<����[\ć(��d� �|G�<�x��F�>��M���-��3 hѣ�����e����K�5Ut˗�1��R����b-�e�1t�����m��y8*ryT7/*d��e�^�mn�f)�J��j�vC��m &��A��&.b���v�K��2B��Ҿ�Ȳ���c����E��O�U.8�AAL��I'�J?5+� ڨ�F W$�N?i�ҿ~���A=�#w�Ux���e�z[k�۾�X7��A�{�5��QZ��s}&�{��Q��(�]u��b� �v�"g��g��*޳��"L��%�8��j=�Gg�%p��4�S���SB�!�A���FT�p���ʕӁ��ž����!�I8-�lxQ��jI�;Hsܬx�C���</�-�	��5�-i��+�����C\XC�4�(�շDw��խ���n�	�Y�{�+RiP�a�g�AY�6�J�v�c�V]�m�`��DdzD��z�C���)�:,���W�	��a���D�������2�I3�u�*���%4S��(��G�D ĎK5So��c�@�X�>:{����A�Bա�DgH�q�u�����j�f4#}�G��s"�qi/s|#�����u�������X�zܝe���S"�B)����cNC��T�b�ހ�!�B�-m����z�3�@�?�O�ZH3����}GK%�N"��Q��[%]���{Ze�Nثh=�9ko
���D�4���8t�݂Y&�3�,��24�0疣���Mw�V����E�>{� 8�!iQ���X�$֤+���g�O㒽ă$��>����!_llqkAw��P���"u��ӂ�!	j��9������}g=��q�I�gW�VXѨH; ������3Iʹ�J骪^�y@���nΫP���_(h�OD���~�d�)�NB�!����l�2*l�~�=H7�
����:��|�V�6�f�`��F�̈y~Q��x��%Q�y��e�C �e8Bȷ�>�+���o�qm��S5�S<��d�'Z���ٌa��88(y�e{eg��:�k@6�F��Yw~���⼨�)�6��W�M���P;�U����;���GA�Ί�Z�4~�1
ȽN4%��>�Hb0�v�8w��:�<>亀�ONC�C�(Q$�t���"��]�3���Q�[@Ρ�o�q�lI(��ϻ�+x-	vL/�M ĺ�Gƽ?O�R�P�'^.+^�P���B�)�����f�M`L�R�PX&���	�� IPSj95g�N��2ˌ��-�d��PM��Uu��*����{b�W�dd� �~������Q�Р�Ox��է�J�e�-��˖4'�0��B�8$��4�4���B&�Ei�]���8��B��*�z��M���2����zw����G+��jcT��6�@��g���d��R����dWt̝u�h�o�9��4���$�zP��ª/�OVg�.�fM���%ƉCh�t�n��~<��0���H�"7�b�,�Bb�J9�j�F��ǎLs]*x���,�n��$>iӕ�?�72��7�U�Y�����z9��Q��?�-S�XA��+�N�0���Go��ә%t��i��Z�ިq��@i�2L͡��P�OkU�['�HNk�ٺ�i�TN�nvz�5�d�S+g����m�ē�o0�YJ㴵~~Aiɯ|&�r�:�b��?E,��a�!;�'�6y�|U����P�Ca�Q��� �N��,���!���\��eUh��= �Z���i*H�<Μ4��.�}g�\��A7/X3x���1�T��~�&��"���nK�4-UGE҈��Mm�Ӈ�u:�i��	��-	@�Dٞ�t��v��E����ڊ�\b�k��{^�5�DI��T�4)�sL�be�4��i����IN��g���H�,�mBݏj�܍M�/��P���� ?NvR��b�^���"L�*]����u=I�@����h�ܦ�6t���a���O�.#CV5.��g}+��|�6~��۱���
u0��&xD���:�c^
nB!�;ֺ��)	|�>��g��!� F�����Ҁ5WE8��"�r����=�������]�P⡐f�p��׉}vT�>"D*�v���/�֋񗦅�s�;hf�x�U�s�5�A��M�Y࢜�աz���(���H#�7��%ƋU��q��BgT�$���j�R���|ӗ�q!��:g�Y�*A�._�툆�8*d��n8����!�4e����g��P`�P��7'�H2��nx��>݁��Q����I�lx�[�$h�k���� :	���
|.���	2���T�X_oƥ�����_��v��B1���U���m�a�vϼa`�����.a�-�ޤ�py�Y�4xL���3[2ԞBr�Ve��g�QH��cHKjЮ�Z1�㦞���i�Y����;����Ն��)��Z���⋠��$i \��8�E��BN�54@}݈i�.cr(�+g��!j�o����0Q$�hM���t�L���L[��@���@F�(?�yW�9[I�w,��������@���)"�0�Ϥ��Nh"ߩ!˞�[J��^U��ض�ѫ%Y��Bv��6��Y#��EJ��M@��Ę[�ш�����%�"Ů>�nyCR
�a��R{���E�4[��|�� ����d#<ٿ���ys��J�?���5��"Ȭ��0���~(=�L6_V��u�Ip���KEBV��ZVcZ�Pyh��Rz�'���Μ������Nʂ
�+�5�`�*%Fϻ�q�,��1��F��F���ﴧF�ֲ��Aiѧ�Ӄt8�7u�
Lu���J�9����3i�Xn�}���(Y�)ZX���mq[��Q�����Ь�Ѹ�u��Es���}N�R=��^ �Sˀ��l�*G~&>E�/� �5�U�(ŵ���T8�"L�F�W�%�a|�J�@���	(]���d�Q^Q�ʼ���U��r�⫝̸YE��q<6XH�|s�a�s�+�/��� F/�B���/h#�P��NoR²���a�7m�����Nd�KSṬG4�ɱs���51\�rE��#/@6d���\l΅�A΄0�<Q�s�Yz�M��M���Ӷ	�m�T+Ã/'�|��E�u�a]��J���O���\�A7�I�L�TM��;����iy�-C�3�Ut8:+jٴZ����|�!����֦1�fb�'_0���Xp� �X�=���,3��4,=�VJ�[`�8_A
��-U��uv������g�+�r(�(|�y$�.�o�����2�`fz�9��������N��u
���"u�jU�s_p#S�7y4Ha1?�e��g=�3��X��z,��9
��]��� ���l9��{�s�l̛��gO�͵w�@KU���]E��Y?�&zاrc6�n�X2���s�� ��P�����W$�/ц����$3�!��tj��Y��$�u"�h��'	[�����g���)��č�:B�ϵ�6[��I.;�^��1�8�߅O-�F+�?�	֟%�M�4nO�����і�R!E�lX9Q#�m�Z��kr�̒�R8B��x�����S�XfQ��u��,���[r���
`��KѝI�_��t�ô��z���p�y�ݎ5C�)=og{Ș�z�����&s&�:��7�	ei4V(�z��Iݿ[מ��mҺ~�0P"
q}ls��5I�K�l�3���c^���T��9�iba<�A,Щ���*����rdւ�S[:0#]�B��)��ɷ:���pb,�M�L�m�d>�o� ���N@?��Iy���	{�DZ��JQ&F#~��_���%�J��d���:J��P���@T��j5a�[�D����%�z���]���[�R��?�Y��9� t���9����0.���"A��T����Q"��Լ}�c��iw�u�6�G`���*�x]BCc��~�1̅�P^����)T�Lר���c�(� #���c�������]��􍷂����`k1�NCt���|�	���_�Xj�O��OM��4��װx�����W*B�a�I��Q7�İ�j���.<I�;X̲��!dZ�2����v�u�Eq8Ƥ&�:WA��1���[�f�ά�ܸ��ٱc�g����fل����]������:J��M�8��e� {�t�bDi����J,6X�Ҝ�jo7����L���;���/>�ۖ�I��[�z����v�b8������g��B�`(����� �������D�ri�%�z��ك���c��"z:ϭr�w9�0	��u�4�a�T�rh�`�����f/�?#%(q+t	��Nî���	��c#��>g��(�W��ģ3K�f��b/~�*}
p��mxJ�rdﰭ����'0�����d ��7�Y|ĕ��b/��p���&0�:.���J��"^ע��Hq�S�W�¬O;��@Z��&��5=jI�X����I���%_7e�נ�w��!p��,��!X����|fZ���ϋ�Tv�>�ଗ�KA4�mʐ|� ��R5(KT)R�f5'�K��b?������Q�5��IV���2@/��_�~�HNy���G���x��C�^nꠜ]:Xg����`) �)���҅��
l�i��M��#�.dix���o��0�*N�0n��2�9:�.�����6��
��%�k��IHEE>}v��G����T0��~���~�qL�2�"��7_�b�=R_\'����x�����3|��f�S��L5^�M �eX�^�7�h�R�~�Ҭ����`��e���dW/����>���=�[r;fJ�.��f}$1o�h��k$�9��M>�v�[���e&��!Z�9��#�N��2��\��'|BJR���<L��}�/����K��Ӑ��s���L5W�W��>~�c���吘�d����Sͦ��f� Q��)]@-���y��Cm���v�դi#�(-����@�Q�G��E��@��A36y���i_A���D�&�<u��?�b/��羰$�{d���J;
��GDd/�
�(��w�������oPO%ѿ�-��I�ѥ�H�7�T ��s('��TE*evG<�0c�Feq"�>]+3x�o�/LYH)�/~w��Jz�C<^Ezޅ����/�F�8�(S�n#��^+7�S<�H5�P��!(�9�b��p���3W�"��5_T$�����U^�����"Kp�ɠ~B����܆��r�>���[�/����K�v���ha�۬�lϸ�f���2�J,�\]/��|N�O_<�[�N���^xA��қqs���Á�N�1A3bS�.`�}$�	3�F���<sW�W(;�6�1�՘�� pf����jN$_/鳵�T�k�ȐX9��N%a�wXei,��$H���5hYN0���Y*M>�}�e��}is/��Gm�Eо:V=�$6��e�V=�L�C	2k�>�zLX�Y�3 ��H����2����+�)�`�G�ݐ��M�8K$�/aY7*�7Q�,���T>�.�VP�i��?���%�e��cVʺޞGmѳK��ț�ᨋC��9C.�"�9�؁.��O,_��5N�����^r���%�>�'��&�(0�?��!ȼ�w�#R�
Y�s�؁��Φ*�o�2/`{{"y�B2�)T�nlAZ0������ ́��9��@
@Wؾ��=�ȕ�)�M^?� �,<��Y"Px=�{��$��s.�S��$O;�
������!ۯ���5o�z(��F�C�<S_�t���1����Ol3H�|�~�/�?��9�G6
N(�r�j� ����yݕ��������iL���,~Q]��<������P��?9��݋	��N��#�J/ �m+�a���#�=6����Fh,Q�	h�NK�8_E�2��ƭ�=v�z�P�E'��p��$V�@��23F�{&�*�t@�x׳@ESF;�]R���2&�,��-�$o�|_:�}��>Kc��*c�4��KqL�G���X~����2��s��V�pD��#����Ȉm��;�iW�#��;#���>6L�#��u��N�cO"k�>����)��R����c0�Bjqa�߂��ԭ#������"��?��Zt�L<X�心�Z��كR��7���D۶=rV�{��kQ x�9d8���������W��
�g�oNߌ؀ 0H���%[Ѻ�S_��/�)�Vjv7���+����Jm�Z�s�9�'�����t�?﷏�̪�A�kB�j?2"X���(����L�ck�)�k�CP�o�~񰦸,pu ٲT��:�fN�.�إ�F
s�^0�Q)9KTI�`�{u�)k��͍���;5�݅��e�ԪX������Y��]�DU�	�k�u�1I,g���7��Wd����軝�md�e��ҹ���y��8���a�Ҙ7��}�/H���M����R�B-�h�j�j����6�_ApY�:��kWeA�����m8����$�I�o8��R��5�\$H6��KG�jt�դq5uպ�G�ͯR�9�WXl
Lƹ���7��m�L�.�
D�dÅ`}�����N�����A����}�?C_�!��,4�N���YN�ZUY��MP�.����f|��O@-C)H*�n�]�ѿ�~9c������o/u#���F�m��b]�;^�Xڷ�eB��]�M �W�q�k�l���a��=��EO���"���j+���Ȝx��a�
�`�g�.C�˒�9s/��<�j7d���$f��aN�kl1��Y����w���?�*�/�n��ˍoq�y��N�cY-��S|[#� �7֓��v�3lbp���%u�҈�k��5X�e⍫WiL�_�$ʦ:�&�'W�PiA�v^�s�1�H��O!���/X(�^�}��B�1�Eā7�	g��E�h��6=%�Z�`Q���~c��Ӣ��R��������,�/��AΝW`w�O9�&��J5��ʵ� ����9$K�Z%h^uA1��F
8}��zKWv�BG��W�Y�$R,j���[��t�Sbh٥�;s�Z��,I�x&��K:Pݦ�h�z��]�:2mmlV)�G+S$�iA�6+|�dM�/��al�WH��U!���QyE�����t�f�Ԥ\E�a� �W`j�:|Z7]9����/Vk����J�I�YR��%���V�Y��R�ĞkU�壴A���&U�������x����� �°'�6%6��r#���4����e�d��L�9� @� �ٹ)O͈ia�?O_���>,	�^�|�����o��D��b�h_��ٻ��٥�k�����ΤD7w��2�G=8������y�����y��-�ٰi�L���n)��d�Uy�%��������14Y5L]f����|TX,��K��f������>\zK�HE�f �+�|�5��j!Qv�6jX�z����� �l�9�o>�U$�kR�v�����q�K��%���*�sA?�m��W�$�Q
K��Gw�K��'���W�/�5�V�[�(@ }��d16�=�Wރ3�<���p����Φ�6����f=��M�Z�J�d8|��c��NoM��Pv��J�Y5�<]Â��8�*�u����c����@4}A?CW����-��Ʃ��$���
"-��裻�������58��[�M\iPb�4���F9@�9���	�kP�j�;�Y�Z�͉������)}�5�ֆ�~� <A�z���'�DLbt����^D$�;\�^�÷���Y�;��b�>���b�6Iyl����8�C=R���.��M�.�c]��{�Zp��!2��) Ùf���L3�sl@L�O+��d���,�'̊�K�|z�n��Rn�`�/�Ё��<��3�ãHq��� x�­/ �in:#����F/�9y�[�+�����9ͮ��u�k
�Z��d���l�3V�'�@�O��b����U�kݗ��Gd±�\�z$<pX�Nb�p��p@B�-�%)�$��ꢬ�n����^#۰U8�"�!�&q3k��I��%YǕ#0=j��E��!� �.�Q��#x��w�YM���8�zs"q*K�YEB��9�X������Cǝ�m�ȁ�K ���,BcAW�G��"`P��z|���Yq��L�M�ns��t�+Gǐ5��1n�)���2m�T	W+���pZlM��G�V�$D	Rt��g� t��"��p��"Զ�z�R�ψo�P��gҕ���A��3$4�ePrٙ����]C�	���+P䰗M=�wNtqw�<Dk�K�����ljQ��	h��ܷ�ɻ�hYu�}i�(��I"�|���
0Yx-�$tȆ�i&x��>��9��3��[�+J6νji���G� �	�$r�[��ހ)���9�e(?��fEn���"�r�'?@i)#t?[�b+xz�i͐��*�;��"꺃�&S$8d�sq뷅�� ���o��5f�}"����D��QFN��9��z:��zZ�@�Ȉ%a�3Uޘ���� q�bܭ�����;���ڂ
�������*��si�H�������]o�Qz՝ؾ��:������GV�O��/9�Ҩ��8��;�>ߡ $�w�;�n�#��:���9��Eۅ�p�M��/b�ܱdD�C�<S	i.�zJ���ilV�Sy�jH4�h����GbV%q̳�jV��:����J�#�������q/;�Z��G~@{Kp��#�%a�9Ȼ�p�P�/h���=�{JB�%�H�;��焾��zy�\�7Eq�x]X���H���PyG	���g�~rJ��Z����7��=�yz �_S��)"X�m�E�A���K#�{5����"֛��>b�-fǑ�������>' ���Aת�(�X�n;�M���4���~���y��w��fv\s���T�Xu���O�i�}#�����Ə��1�Z�����H�����x �d���Hd�YPn���ή�g�I����lϜfS߰0�x��E6�k�@��5�@��~�.�dz��q�R ^�t��\f��7�H5bH��RFZI;�,�~=������F3G�.J�=wc��]���dL���q�Aop��yH+�U��$���hm�h�QҀd������V卟MSA��6�S��h�}�/lݶo��[J{��l��073d����C`r�q��\>��{6�N�qm�󀺿.?���ٟFI=2���,�i�q�������շK�Q5``�2����b�4��R�!-���gml?7ג��ZP�I�f:)!���q��S�;y��SY��/��Vd$O�����&�j��i����.�#)p�s4/� ����S�e�~S��y~�.�y�Py䜄����b2�z���ŰR`��C�Z
��;��սO,-�8]�k���BM���k/��wE!M[x���˓��H������#�E?-詰T�Y��b�c@��S��Wވv����g��{Γ���)�n�S/e��0�c��<�/}��G�M�C�����1��%��W|���� 9/�i�Ϧ��M����}��/:��)I��?wn�(:�?ʱW�:��qY����g��e5Y+����T�X
��;�|�rD?� l kl]���W�q���-c��y�;�����&���}��c�
C\)�p;S��~��R�R�f�X�R��������c��@�=@t�K
A9��Kٻb��E<���#�"�$��V� ����*��=���V!��#�"�RT���ֲ�o9�UF����=W�k��8�
3�a�!�^uS��	�fuXMC�C����9�Tz�lg�H���=��31{�ف!��u"���*��z`j��y	1�xW%P�)�U���cM[����&4+|=�.R�.>�0�rd�C�|+�.��.,^K5��6�ޕ��l�E�3raW����/s�L�#O�ʘ�m�_wܢ(%�I�պ� ,*���C���@�sKP)�@�/n��8��$X,��f(d	�I���T1��[��t�3������h)4�P_W��tp嶝<M�h�G�`��7˷i� �\
q�V��:D��/��JX��c^�J��?�$V�=�#��T9p��xt��z���Ŭ@p�Q{��Rx�V�����sG^���y���!{���7��)d~��N�W����X�j�m:��X��{��ӈ��>ۨf�.��}�<X񫣢u���s�|w�~�f�g��]�1���X�D�|�H4y><�_vtL	���J���ǎ,��iYc�9��S�8��+a ������T$��O�h����R,R��RzFײ:��ԮZ�w�a#=&s�P1��o�B�Qe�X���d�������L��u��i�.��t�r�?����?/�eC���V�+c��F�H��(��D�͑'�9�i�?]j�.k�;��I��c���oHع�D�l�z�v��ec6t:4�����RFn '�%��xA��U���$�� �W�R�Lt[��`92E���}�-��^��%�x�>Q�qiV&}���D�I�|�Rep!Q�ݡ�3����ʳ/3�\�=���t�<c���[�l��6�������4 g�6�M:flS�yJ�,Q���ڻ�6�>�^���d�`R�6^�^\���Dɛ�u�$�~een�@Uvȅ��X&@}�|?�J$�� �����qB�"2�(wlD�� TV�F�~c�~�x�^g@	Zr�?d��f��-�$�[�&N��:s-9Ɉ ��t0�b���N�_���l��.Q��!j��ڸ�t &.��M/�`4�};s�'�"V���%��|v�TO'�B��(���Q,���~T��$��ļ.w~��}UF�,P[����^�����K��D��sړ�Qy����+�`<E��O����s�niq&.���f���o���L�'﯑@ŧ�@��4p�\��:b!�^����_�h+�/��
wgh)Ƴ`a�v\`��7N&�k�q�y񼎆��WE/��B����� 3R��j)���:*E���!��]��5��#'[�YL]�m}گo��V�^�X~|�N�v\K���Z��-��T�sD� ���?���P�p�F�T�B4wOa�9Uw	[߱���u[~x��.����{����tS��i���69'H��+CFcm�l���ӈ�7|����v��>�����S!���͑�_��4��R���=D.�-��i �-e�
�[M�� ����UP��FE����AR�����$8+]��;��~gc)>TK�]S`�+k�4�Ul��06R�j+OE���G�ղ{�^3x��5�����ʎ�����B��W΀�7� ��K+6���R�ե(�cn���9p%�=�X9B���7 �፩��{�l�A�p�n�u�)Mn���jw��3����U��K�,=�&ci���Վ�ʅLjc�+�M�%o'��J��"x�3�O�z�	F��Ч,/3��K,�����HX"(�`(�;��Fk������bo�R��%�8RC��ާSzK;R�ip�6W�Ií
�� D��{3%��T���������M_�*�^uO2�H���I!�siu눛�Ks��"���B�#��^D���A^�n���*��!	��ir��d�j��l��~�D\/���z�X�G�ϭ��5�� �;��H]eX԰�~:�����?��u��Y`�9�syndj��Kj���N��&|�l�q�
[��g�?E%\��#Cԅ��dwt{�Ș��k���������hT'�&4*
����L��J�e��j'-��َ�_�T��G�x��]�l���l>��h�]�Y�zT�!? ]Pw,�-�/vB�4a��O����PO�*�4F�&��!J�z�a�z���V:����yyϩX�:��ܩ�zf컺P�7ː�6�+Ү��/R*Ӑ�����Tu��I�zv�Ek8-�i�L�n��r���f;U��
8<H�[�(�2oM��D��C�ʑw`�����j��8~�!��c�ʅ�܍�	6.�8�@��ؑeCL�R��3]���r�'v�
���k�C=+d .N���N�RO�s"�ƕ(͢rQ�w�������ѧz�$��W)l`ї�rݍ����N�ăR�K���U{w��;.H����dȼ�\y�۽��k��N�O�aZ��D�Һ��{
��eY&���=,xw�y{Z�  r��8$��,������=S�VA-�Ƨ�շs��
���Sm-ڶ�:����Ϛ�m��|<a�P���K�<hO�^y�x�����6���H��DZ�r�-K9]��[lvdg�0�{@�>rB�&�4B�~�Q|?Ҟ`փ=$���(���~G�(CDe��������*��I{W����?�����f���ł�E:�J/8���g"^�\�b�'���"nb�O� �G��`W�H���K���AɁCDAq����y�D�h#�ʄ�4&BIE}�)�r�@��業�N�eP̪�Kg�����\K��oz�>��d��1�4n�7@�!&�M��v� ��V�$����KS3��$9���^�[�<���qQ�r2�u�YN��2_P"W7!�A3��v�>���?�C��N���ڮ8�`ZIä��97 �^��BRHH#�֚6�@�dr�P'�����&Y��,Y`��!�M>]���;����;���m�(L��b��3:����ɘ0r�\�F�:�!C��{G��va�x���VM��P�P'�~vƗ5��@������SŽdH�їXfZ��Ǆ���j��yx ~zn��Ǌ1�&H� 1�*�������C
�_���`��Ђ�+�7��JXӁ��d'���H�Ȧ2�+���A�z����v���@V�/��79��8N�Át��z6]L:�:�;�_Q|�ʧMޭ��5��x��䬷.GneϷ^�)�mՙ>�������j�&��R�6��'���#%��9��L�f1�B�f��[j���Iq���3�v�;��"��a���+�*���Y7F�R�k�3V�l' (�r��&�I_Pt�~�`���sy�C��w5�||�m�|e5nE�id3��˵�9nC6L��c��ހ����TN�;��#}���ʖ�E�i�"�c�銫�V��~e#�c��8�������b�DiǹV��kL������O�d.�]	�yy��������d���;9�p�O�Bx|S��K[���x���ئ:�SA��[��ҿ�0Q%2��2�_�`��f�!�ؼ�o]ڐ��B����&U��f�	�^��̝6a���'%.�KJ��7Fj�m�3K��.��ۖ�ZTۗ�|�ޏZ�/U#�"XŔ<�����U�D��t''KBٮ>��T�e	R��z�B��5z���~^�3�ȳ�:]��.���Oz0�Yh�}�^�\�)-�2�z�"Nx�e�q�Eq��7�	}�g��6u�-�l����vm)�fo*�S�n�W"[�"���,^���Lɓ�չ|qc�i�0ɟ��6�q��	T:V�Ҩ6����禁�yҤtp��8�*b��3�\�xњ�����՝z��wp���?R�e\/}P�CW�A@k�"w .H�zQ�۹��;�Q+-�@�W@d�J��eZu�-)'^o���^3QY���ˉѬ��{�13�x"Xa�]A�H�
�-_����sK���1�!��ͦ�
�N��
a���7)��G���QD���R���vXMne!4��D�qw[�Q�1����+�y���	��lb]���|�kD\�Kb����z4�]t'�Z��t!��.A䳯��^���,ВT6T����q�+$'�N���W�,����j����>|���%�v,�Z�.9>�h}D^Gk0�ńg�Xk�Р8X�;�B X:ǣ�4l��M�vv.U�fi��&n�*���#\G�S䡝���a��]
�f�NPB34y��U�K6'E�t�\C�oέ-��=�S���,����8�b��GFsRXK&q�P8��?2���������n(�� C�𺪨/��)�@\Vrc@���Dl�Fd��-�͂��`-�w��L�ws ����������v �����`�����'���@!a\w�漂� �{��Ҫ�5�hEL	�'jYdDZ��p��q�����ɦ�Pfz�v!_���<o�b����9>�P���7Vv�'�����"LFr`U��Ƌ5���r&����zjnb���?��6`��^����0f����139��D��n}��5�%7��7�曏 �۴�c�<�mi|��/`5=m<,+��Ov�!؋ȅ�W��d_3Q����-��,i�"��Stٵgq�% a=}��3��uG.�����ðp�`�B}#�Ih���א��I���	/��4ፂ�>w�~2��4!]ʌ
�n�E�Y�[��ۏ�dM��s�2��y��	����&=�]¬��FEM��~����?�4O�̴���b�P��O��]i������U��L> i~��P>M��Х���B�\gM6�7B��l���w	�j
ެ��Vz���R]��6Fxƥ�M��{5���+�3���ܾ�p��9�߼ۡ_g�2d�U��D�ب��6�PLI7�_���N�%��y��m�ţ	��|ݞcz5�;�������:���ޔ�ҬهF�%��ʧ��}���d@�XFo"	�l�B�pn$�c����_�_Mht�J�wE��������?W������#;�A��xm*�.�~�oJ��U4gE?2蒻YE�Vf�i^�¶:� �}_�T=�>C���B?9v��p]vB�N��Ѿ53�J�3������%	��7J�������Y%��%N���S�����3ڏ�9��0���lGݮp�]Owݴ��ο���E�!�,��CG!)�/Z�h#���X�U��^�vo��C��ڳf#h�1�\Y����N��O�R���k�m��r�h�׵��(T�Q)Q�����8�im�M_�NpO���#�����1�d���x��N�VT�P�5~���`�9��|��������?z��\�o[PW���X5�v��7'����%��-�� 3N��݇9O.XX��9�j��d��,�bAy�v�.)%�%C���Jjт5*!��|��q�D1,���ɿD{�V-��i�Q�8��^�Y�C���F�M�`C�q����R�2����c�]g_����wJ6����,�I�+1�B��q0�2'~dc�J��}�ı��0Mn�S�%ߝ�`��F�) �yS֘!�y�Gh�|z����3Z@�͠�^��nxGA�����T"�)�����&O�FK��<g��)f���+��r�jd�����ҿ ?�렞�ybr���֏�q�Io�ϓrs֮� �9M��J�9�<�V��OW.B �x�o�'�@g�'~T�,���M�{��7�򓩘�]�p�m�1掦�?��}}�pׇq!o��X���R�����vR�R=�H�!�@p��o=T�W����/�jI}��ij:җ��-�,��!ܹ�S�L��?į�1�K�>���ʊ�!�ݝ�Jŀ�>-U�po�a�Č�!%���m4�!P�V��M�z��n�����ݓ�E�US�:lw���u?C 8��y�2M�Ma�F�7%���׫�vo`tu�D��-2�J�$3V�v��709�VP�?�ٖ�T�@'L|�����x�J��b�G�jyW��&�Y>r��L�j򁀣1���"�����R8ֈ�������zE�p	�n��x��O;M�����jckPB�S���7;�T��u6-�1�/T�s�?�Ա��]`ޕ<���9G&�RnW�a0�>�xD��^͂�؍�HS�����#Ѩ�&�DY#4�hI�b�u�
:ѱ�/b5�ms��/�7 ��S%�_`IIu�gdr��[�&;�ά���&�6P¨*�YH8u���ߐ�;ǻ���"l ���J��2	�Y����F��<��� RU<���R�o�.Qc�)����z1FI?��>r}���C��#�(��-M��]!)J��q]����8��d6����7����}�s�˻t8�����edt�%swj��[5K���_3̅���"�Y��j��8�o˥s���N]f �3�����P�Ժ�A.
�A�O�I3�����歇Dڎ�Lt6��e�$��,hR��%�Iڌ�I乳dj2��d�ʢ5����	���.K���2�6ܕ<�EP��;خ�~�[`ΰ'�PT%�3Y,q���S�Hu����t;��a��(�8>ա\wV��O�w�������¡�f]E5X�$<������"���5�̆���nxL��:�����qV7��s����������=?�:-X���0�j�A�+�<�2y�z�C�E��M|j�'8�=���(ZAu3���@�Jt��}��)��:��1��3`�����A@���%>�*�u�:+����Ive��D�*=�X�B����G��R��N��F�#:DU9o���#��H�����6E:�NƮ|�/�iw#-�/��A�Gj��u=�V2��ҢyJ����V�L�/[�Q�"��[yT��<ʢų�!�74�
~�������f�l^Qş�� l�ɲ,�PUҮ�íPu��a7���o=3�'鴞3,�+�\�\ݩ�p�b(|/ts�R݁���1^�B�̿&�j��O����0�U�{�� ��O�� �*P�����S�(��5���$A���M�e����
>�Ԛ�I,>v�.i..����E�oxa|���oê�}`�P=Q��I߈��_F�{בY�=]�D�1�����mcR�����k���\yD�Dh7��`t$�s�[�.Ef�{�5X=����P( ��P��`�:^:l�Hk�5
bMJvl)1*@�[����舺9¨�a��/؞MK_��t!jl��ȗP�G�@�F#"t��`�Ԩ@>W ��f��3ߑ���8����ё`�b����o'�.@a�Lˌ!��\���@+��Ԍ��n��!\2�p�����\��Z����)m�绒�G'Y����p>F���B"�˼�I����A$%��a��[���aa�O=�*f�y��zb�Ǽ����:נM*�U�D���ܐ��⊱ؾOP.�#�9��xAt�x�ΈN�����%Ӵ$�N�2t!���c|���]�*{�#@#��J&�} Lr���#�{����dLn'ĥN�|�GQ�ö�F�Ă��JCA:g~�{�3�=�3BhR���$��%1��"���O�)Z������L�4.��:�e����(�-�:i�6�+��0��:��BX��*��N�L+�V�g��=���6t����<��qp^���b ��� ���q�ʯG���-��R�ճ�$�4r^>��l�b)ղ��$u��Z�#������A�Å��mF�MCZ,�Ԇ��,�ϐQ�������R"ngT��&7M
ÊG�*1�Kd��M�Q��V �E
3CϓL������"*�0����qaQ�i���C���u6���m(Uw({K��+H$��Z�A�/�o���F^^&��1�/��=Qt`<W�Dp-S��h����B^9�
i��_iȕ�yp���T��@��=H`Q�gsI;~Բ-�X��q�09�y�D��W~��n둽�L�J��Ģ5����d)G�O���5D���Ϣu�����"L$��"��MUj�7��Ɖi��* ���!�Z�����%��'�X d`�����ѵ����>�$�K��>xk�U����'��]CŅ�Um}M�7�|Q�8J�-q���d��Ӳ�%��٩�qH����jN�e�}�ܷk��ub�SƌS �?�L���E�+���_��`��� /�we�4wu ��|��/��@ށ���:�x��X�m�H�*RH�'Y�u78�x���$.U��:e�˂�#!���{��W;b?��PIP���ؓ�c����$�l��mn��_0�k�z'!��{��G9���� �w�P�ʵ�ȚN����Y�oOr��8z(@����T�T۞(WR��?v�����k�r5q'·�!����XS�wfy�X�-�C�ԩ�PA�eAg�x�
F*�^@��E$ �"����X�4��(��~]vX�E��G�/Z�;���ƎѰz�CNǡ�ho>���շL:j����*�+��?��P���vy}ͳm >���X0_EȘK�5����Xr�b���`�^<��ȑ�z`���,�ta��R�~�hyJmIUYZ��k��i i*m	�0t\���,�0�B	��7-�q���3ːoE���z���t0&����ό�*���5�ri%�����zycdPͺDC������3�܄�o��+��?�.AOW䣿��i�H��l�1M)�0�l���}�������6�۰�ł����Ɵ�4O���y���������k}��I�3�WOH S��ڢ�9�[jx�H ���N�HǺ�D��S��!1R�����]ŉgU�n`��\�����^���+ikW5�:Zt�������Jn�}e��|�C�5cV�&�`�?ݳo��phL�;wѹ�C~��{`#@�E5�ҒjƀɿG��o^a��D��Xp�#�2�����6ܘZ��0K[,�71�}��c�GP��H�0E(��RxN={�v<}��l�������$K4�k�&���d���<�N2�)Z9�8|�
bt �C�|I��
�@:t*#�9���9��7��%W�ʲA� ��T|��a��~�րZzK���t�"�˖�
ѣ
����ض�6�̥��fƣ�.=S�`2��
a*碓���'��<c��]P����2Ѩ�1
���#E&f��o��}��\׺jtE��I�P�`��1h�p&�����}�'��X���=zn�"ps���,�B}9�ҫ�C�'=��bX5r��*�/M�8OD��@��ق	����UU&TS/����T�Ic����Y_v׃` ���	�$�E��@�ed�U]T�����Qh�m�/�h��|
mׄ���U`k����;���	���{�c�	R��l'��L�v
Wa��s(.�76���]X����O���ZZ0mV��(��N�Ϸ����M�gݙ���&��UX0]�D��d��G��lHɔZ����u��B���'4��k�Da��-[�xH��ڋ���&�AkŌ#�4���<rBE
�4�z)�hj�|����%;-^ڍ��ĒЗ��VRhW�Щ~
�`@���I�G0��WP�ZC�F�����#AF��{�%���8.R$���}��5v�d�@9�Z�q�� S(�I?�$"܃q &b�<�q,_��������~b�nv�X�(�ط�C?	x�*�IM����-!�i���w1K���DM>��£͈z&:�z8���Pf��s�h����t�Qb�J�<�N��mϩ���MI0h��}>~KpE_�������a��R�,l���8��������0�&�����ݺ��i>޵�/��#u�(�	��UY��r��k���l�����A�O�@ty��O��P!�-ӑ�y`���	�jp�'L�HI�1K�=�]���^��BH��|����,%0i�}B״��y�՜J0*ķ6t�y#�m>ܐ��V��b�W�>C�dy��:
���s��X��~�����?�Xj'�:��M����mW�T!�nYu瀶��a�
6k�%���1��vF �&���E��Ε�3����5[�d�B�o��T���PX��L/����d�PV@� Y�jXI����w�J����ܞvFeZ���-�?М�N��;{nJ�,ύ���z�A)Dgh��������b��RG\V@�X�3��Y���،����w��V����^�L���S�DpZ��deiG/�XJ3Z����6Z��.��ԡQ�*�LaE��IV��,�mV]W#L��Kr�-���c����p��0��HP0%z;��mJ���w��/Y�M��$�K=�)3�4��
샏���g�������9�c��O���c�G�|�5zOc�oLZ�$����S���������x.�_��^ބ ��fHBe����g�(��@Cq�4��p�{$�F)gy"�zwM��Z���פ�u��}jg[� 	h�9g�R0KPӈ��5�wc=�x<��q����}Q����H\e2���j��Yy_��9�}5�}e� �w�E%��"3I�����L���6��*�7�q���w�tf�	e�3飼|� ����(R`�
+�����p�"
)�����Q,#++���\}
�8ޣ>��U�!����-R���[I�n��p��c�]':E�"5�l��������8ΣX0I��	�mr���9��� �a��Paf8��|�tӘj�~����@ ��#s�9[���}Wߊ`�+,9��r�!!�R'vu�ٔlmH�������1�`�-����gՒt����S���(Q�!0m(C�E��vg�<���|���[7l�.v��g�wɢ�a��6VAMD���/
��{O������n�p�ԇ/��TP�t�_ �K��]��Oc���g�ǽRt�ō�ׯ�%]f�A�y+���@n��%�Yv��I�[8��7�PT�M��&wO�b��3TZ��1e*`m�\�:Z1C>�,�"	��
s�:�vu�K�k�`�g���1����:�.��^�#Q�l��� ���/���bC&��Qit�H,�>��x�K~&�4c�#P��s��7L�f�7%ܸ|��C�S�pT7�t:�?�c�^.�ogWs{�(�ݯ��6�B`�&&����(v����\dH���N��أ�ܛ1j���0��ډ����s�VDb!������j�{���M#�}��teg�*C�9� /k_�ی�_LC6L<b/2�'}lK�P/A��4�눜�Es%��©��R�~�eG�S�+`�Bimjp�,ov����C�{�R����?�V���.% ��/K����_�[����]��>�G��C�ճ��h^��xGȥ�����b��>:
no>r럨�n�\��-�;Iv�ק�t�V�Z�ˌ��]�\R�YTݵ�p9E[ûgYg�A��[�7�7� �;�J��U�&�z=�>�/��J"+��ӳ�6G��WȱC#֡"��u�uq�n�����1s9�a�|�f[�:��sK�v>WM����pZ(Q8g
S�j��X�&��R��,�6�n����ii����Y�%C�Р�T-��� 2�ya������HխSQ�#le�#�Y�6Y���?9Zm�;4սm���nF����"��d����Ԓ�_Џ�,7�X�M[�-��ݙ���{�@�R�����.ȭʟ���I��:�C�>}��9Ie'��x-��`��w�b�Tq�o��yB[��;�N�g�:���e�6Q)���v�
�4��.�WO�7��j�؟�P`hmArg�\@�S����q�ϑv9��1$Sz��U��t�i�ʑ1&(qR�����"b����ҵe��z��{��giy����k��&��]\�Ҹ�җ�	�-q'��ˢ �p]�)���- �2���~\�6�(.Za`�z�V�Ȑ�Ix�R/w����y�\��K��D&��2�{:=�ѝ !�����4g��خ��r�Z��J��|�{,fB��)Q��UB��v�H��r-bdɶ�:宑��`��.��)����s�s���+�K% �?R�vq�����4��E�g�R�@��s�&�����޽�.�W\-�c�ن�!D��,t.���Y@Z)Rx�97��ΓbFcA�vD�>�5mA0���$�/}įj����M���~�n�@��R\oje������ZO�e�;�����o�V����pцV�>*Ξtd���Ke\p��ΰ���ڳ�F�D�|�?�Je�˅��z��?u�g3m���jE��A�o��ƭ���uqp\"{���&�fm�����`Pi�gA��s0'0爮�>��� F��.s��ة�)��h	��D��s������qn���_�m<�*�X
��=2h��u�!�ք� ��3x"����c�;��{ߦ4���O���5҃�>���w����pA3�]��ݲ^/@
]�=�(�7�e���o��VjU���&����+��$w�xiڜ���G���w:���U�g�^��V�4 ��.(`)
<��H�_���U�泚!��(��_�����2ד������"�������^�~�}��\t��30^�Rl;���������:g��O�����֢��]n񶄿.��o�������k����fB��Z��M�,�B�V����Ռ&��G��hb�0�+#�?�|��ڒ���0eIw�&Vq���9�~����3��z튃�w�s�75��'��!���|saJlL*��6B�twY��l�	�b����zX)��Nj�0	:x�)|�xb�����	�a]r�4�H�Gq纆��V�gDi9�^rƓ�������T�E����Xտ9ƶ�*��������d9!�V�K��HDvr�����JL�T d�\�^׌^�db��@���dO�G���!��R)��O�!K��K��ϗSo�������]�s>X\�	v�G%��8��^�󈦍�
ɋa#ڣ�<G҇32�==�v)���σ�	�AEr�� K�%�2<�G�"L�%Gu�i$5,eȧp��^E����|q��C��w}���~�e�q e��s0�G^J���zn��1�|j�-�Â�I��VоiF8ˁ�j[�jOd�Qv<�I��v~a���+\���z�uw=e�$G��⍈4�1,�Η��1�>Z���NLNP�Lí}WѤ����,r)�>��:�$���v���c����:my?��fl�g��2s#��"���x�m��0�M��uY"�K�ࠂs�^E�Jx�4X(7�}�mڹ>y��B}l_I�m���we���4A�ЗM�lIO�%r��B�3�ssc$��R��Z�4���uy����L0����[�rn�I�?� W��ԙ��'���g�� j����э�!*t�v�"��9��v�b�: �6o��{�gt��z�L�B�Z�wQ]�@-�Q�AՈX���\���FY����[a,�31�B�u��>+��򪠑PNh��e��0坧%>Gx(�qq��bW�E������P!/�{��u�>�:E0k��Qj�m�M�Ԝ�I��x�_	���o�,σ�M���8�����pO����2"�-'�Y�k��.�vM@@C��
�
��?��X-0F�ǥ��ey�$<z�Mw�;�*��fP3 �Z�K�G����7F�P��}g/����������C^\�dy�u�k�1tQ��WI�`�Ѝ�|2%ߝ(I���/�<aC�>�iOi�IyL���o���N#~��8R���T���<ܒi�� �
A6<(_�"��1���+�*��GP�#����<�l��bJ��- �=r#���B�+�S�_��U%Z�nc���>;��6��*���-n�j/���G岒0`ws�T�}^;E�}'�Z��Nfb��z�Bo#�<��OY�3��b�pu�UIַ��=H �a���CS�� �H��m��~_a#�"�J����3�tc�+����"5�8�K,h	u�x7�G\%�W����6�1��,�����8r�&�U6{�G8%-+�gt�z��E�䨏�q�&�_YD\�5_3�g��lo<8e��8�0;��4�9���e�Ri�h��3f�&�$����z�RLm�>b�f&�ǸT��iO�j��
�~�8�,���'��djA|�V�����r7�L��t	��n�fz��:�����%dy3s|&N��Ýy��%KP�'��4%��5��ޡ,���U�L�$�A�)6�9�M��;�xt�G+s���z���8d�ԟu��-1g<�WM��_Z4��_'�ޡ��%=�r.L� Hr���+!O������qTI����Ž�Q��j5:�r@�9��X���]�F�\%#��� �BɎL�_�=�#T�5?�]I�'�ߟX�V~�`mAQ\닉����8�wFE��/i7
�¦vV��Y?�[�[è;?~[��fmcq��5��F79ސ��*��^����������}p�~S�0��Q"�<�62k�O:"
#;�FE����X�0Z��NX�1G �0��i�d�d�XnK����^uCdh�YŰ�7'H���)��f�e*��I�h�ǲ2���.��X�_Խ֮�ش�+�p�
:Q`V%�G�*�[oy�j������T4��JKJ��k5m��D�P��A=�?�q \�D�L!��۸͢�o�Y���	��7����~n��k���?kI���D]�Yl����NP0�&<ٝ�\Ձ�N�-sr�e���a9�$�d$(F�����Z�=�t�WH@�m��D�ɺ*�q.��v N�ˊݗzS�(�H��*:Kn�q�r[m܆Lq��p�a�H�94�n��'�)�S~��ʥ�3�")T����� �e�[@9�����˜�ʋä]�H�;U�D�n|���Q�@��QP���A��2�v7�/�ǽ)S�;��kP	�
��s�� ��6u��l(ʘ�$J���]�Y�Du뚷M)��pF����-��L	U �md�\����S�p`9
]�L7�lww,>:�FƉ�R�yo؄�5���*�3�Y�c�la^\^��^ك�Mf	=��N�`N��(��w��7�1��\U1�bl��ٰ&�v�����dۇ�L���8g�jLe�ZܳǴ��;�t6<x8W"�&���Q���2�Z`� �9�5Y�P��#9t�;�{ݘ�AvZ豓hY�gr�3��W�0^-&���A16�]�v%re��ِ�8!u�j�jݯ�Z�n����d/�����j%�-)��x�o���oϑ`��	k�E����M9�E=Q����b�ģ��Ť�oU�~y�:}N����{�y���x�V��<��f�k�<r�����(���ޤbҽ�&3I��2�����נ��+s�&�UK�\��f6��)���ɩr>�	���:���Q͢S�Q�cT���)pq�G�����o`��d����w���J�jߣ�I� �˺���n�ANtW#��}�1u�d��BO��1P���s�^{_(g^I�n�B�Ey�b��& y����	OЭΤ筕+N�|fP�Y��!�5$����ٌ9[�d�����&�ke���CK�*�X6>�W�~AL!�}��j�4d����vQ_����zw�,]u ?��#�V�r���t��uZ�Av,5�k��e�͛�=����V��,��-�9�V��ק,��6�*cx�}kŝ�'��[� �&v�O����ߙS�c"+b��b��wlR����=?�Eb'���HP��>��^�_�(B�n�4堾�P�*�� �p�y��MG4����':�3��x���C@,�,3�q��(�SU>���lѳ
�uOz릎!��6(�*A�=�}��1��!���3h��s�BD�6����/H�4�N���ʣ�s����S,R��A�f���%'�hW>�J���5	W�(>+,m���1���eE223���趔�fۢ�x\:��x�������q[#��=F�v�v��L�%�T"�*�	´"��Ы"����x��w�P;j��+`��𣺝�����S{m��i���^�k�8�-�n �¬���ޓ���j�����1�t��nX��g��Om���oe�?텠|n.V��\q��KL /037cZ��MWǙ�{D�J��c�.��ߞy�]'�|{��5��>5���P�Gfjc|�����1s��v�aNy�����`�ȗ vR�ƚ�Qi~��������C��RY
�ϕ�Fu�S{5h!c��v<˔�_�T7䪎��y�輅%F���L�|�J]<;e�B��Rd��R�x�-O�+f������:l�z��+<��d�gi�F㾙	94��0�����r��������v`5 ����mP+/��(� u�=+��`����d'�Mp��)�:����S|�θ$�SN�+�ZR��|O/ɾ( #�_���]��Ɔ]F�i!�X��� -�F(�[W/d��%GX3玖e�]@|av�(�P-UH�A]�~ꌉ��:|,E;���5���|��YqqH)%L5�eT��m}f*��P����q}�	R7-,w�J����$/�s�6�D��	�s.�M+���6r%��j͕���t�-U�������Q^����(Dބ�����-5ْP;n�����5qH�~%_�3� �	.��d�^�^%~M)&�m������%�:+C�Sb�h�=+�����s.h��Xg/XIWe�jk����ډE J{"؏��׬�C�l�;��+��[�&*���Fy���0So�;�(K���;O,�d%�9�;Õ�<R6�e�^9z�\��bS>�IS� Ն��`KE<�uw�tV�Ѽ��+�i�d.��՞������#=����s�3�lI���}�i}�P�U��M��#�1�,z�j&��Z�`���Q�U<�K�b:��0�9I-��Y{g؜�D���`�FA<D9� �S�LtB0����O�����1b�Fᙉ��� ���Q���{����[m�u1 Ko�d�q�ۆY��t}y�H�JWꘚQ��g a6��Z��s>@iC���൙߁�2ؒTC]1k����Cc@��+4#��K�չ��y�'8�<�f�#%���p�r��!$��~NL)��j�h��u��6�I�x����8ϧI )Y�C�Diihu�z���c[���˥����7j�#TH�Q˻s����B���Ll���^u���lϺ�m}�k�n�X�n���&L��qD�zL��Ft���69��4�����@zN��|��n������2я�Wp���y��5v3����,Tv.��#�#�B��f�W�!����BK&z��қ:=��B�$F�oҹ�96����aik�0]���O*;?�����=T3^�Ʒ���j,��
̸����t�����F�R�x��F�����H�n���,�N���</H_܌��e��D��`��Ib��Sdl򚶨8��ڑͮ�AIӇ񥌰uZ��K��7@�h��k.��nj����.�#Y�3�ܢ�/@�v.2�^�P��S�2���|l�o�  �g���zG,�)z�|�ӜY|�##��0z�a3'-�,������1�5���x4�!�\��B�=Ɂ8�6�d�4	nbl�E�)��L�Ýc����uA��g�}������O]�Vt��g��n[k�=!�+��~�X7u"T�J��GZЁ/��U����YA��c�}.�)J��<v�����B����:��;��gr� F���Y�"ԓs)���h����/>H�Hֈb�2�s;zC3��<�'�Zv Z4���?5�r<�kl������q!6�m�+��[��2D�/���z��ai�{�\3��mI�ێ_�e�L�Az���.ǝ9�=���ފ+�����2���U��;���S��"�	�1A�8��.�@;��R��n�44�u$�k�>���J.�B��iؤ������S �
1w�.�{���h&�ꩉӶI۬H|�@c�̥���������pQD�#��0*�/�o�_��;�����|�9�b�!&	Ab+��N���b�;��Z��6UL��t�4���j�;����|*��vv���7�eۮQ(#�!c^��i�R�W�'�Ü+���*��F1z"�x�9]��5�'�<�}r!����^j}���Ο����xvU@߷Ux�q?S�j�#�A��8t����DE�������N8�ŏbƄ���f���tvA�Ђ=�7+���-�����YK����I�(�{�R�Rǌ�u$�͟s}��Q�"OR�u}����-��)0^+d��'�6���AԛL�"#��x��I�ۜ�-�U����80u��ߩD�eZ!$#�M�7{�������Nv�2ʪ��_Ζa2�,���d���HW&_�Ņn$
�ފ�W_B �_8^�~v��h�=E+���.aΈ�/�xt=��bX����R��G�ƕq}G�2#���N�z//B�=��ے��$n��tr��#f���Q'&��n�����|���q�P#�J��>��)�o���睴0���<���ɨQ�)`wh
�.��n"�Z����}�H��x�-��a���\1ww��(rd��l�=��f��<Z�=:��Sf'.��pR�eD�àc��P^6�肢n���z�N�L7x��4s����k�+�j�6\���2���ϧ��L�rc�9��	��z�q�7�o ��9X�͕�*qQ_��<nه�X��;���o��-��Am��jtc�l��oI*��c�1�����k/�Un����Io�t�������آ��I=�*{��z�]^2ZG�a�5�7ʑ�����q��U����fx����h7o���0��	<o�_�7�{�����Zrg\@�/�v�E:Ƃڣtډ��[�U���X��܋����|�7�o9�K�c��٩�=�����ݫ��+�xX�}9��|�s\�KO� W	 !�b�$ɻ��	�m3m<}�.���PBh�.�	��9�Y\�%�Q2�d�T::��Oz��� �(�|��v�����dڒG���94��iغu�V�<^�H����'xa�вHܰ��@�a���ݑޘo��	�-i��KNc|/���ډ�ە�[ MJh�.k_l�g�pj#ԃ��jnגъ?];�� ���w޲��>D������� \2q��Z��-�5&N�-������c�M�]����U��[\>fo�s�ns0?�F���s��|K�ɸz�E8�k�>�{Ѝ���Sh'M�3��t�'O��=�Dq=��d�������l�S�.u��^�t�*CC8����� �JO�yz�Q����<�T8�#c+���ҷ�����#V��i��ф��n�,�}�j�gj�g�H��<_[��K��Df�qh�v��h�QX=dҬ��7 A���
l����m|��7<kV˳�b������4$	 ���w��_ߦټ̉���J$�~�c$�\�mct��t�[����|�GJ���K��a�N� n��m�l�����,?��P�A��I����>7���#���Wɑ��V���Q7ð�a��	M?��6T]K���Nb	�(p�~
�PQ3�b,��~"�d�c8ǲ2#�ql�꽅�I��T٪�n#�e�o;Gt6?��Oe�4�H�E ��Ը&�Qi$�n�:���1�HfN�+�I��I�����=�#��-dԽ�ۈ�����=�+i���WUN"�W�%����� �Q�FgF�$U<f�a
���
�b��U��{L�X[q��T����E�9.b�CA&^��r'�����N��YXS�/����"��]t�@G�Nu���\�Q��|���$`F�1�����[(��-���y7�S������.���MR/Am�@�3���7��\��\���dkЍ�\kJB+�g��k�Y�"�a+�b�6_��aB�6����Iy�C[�5���  >6˻]��@��f`�S{2��vр���-}���iM#�{���_��QfN]��KhIĻ��$9}ej�U��ݩS�YV�r��m,���U{KU�X�Y���\�L_и�G��b��K�D�d0 ��ն�1��U��r1V:�#j�'��t��FJ+3�q�Q[�V�zMQ� �e{7̸CG��A1�Y�MC���`�q�GbP��ݪO�i�H�H��>;�Rj��F�|z�X�q2�i���A��6&��p�@9~�O�q���7-�I0�K�(�������¨��>v���4ZFl�`�"II��6�5�U�@��yTY�f23�b�ӜʜkG��:d���q6��W�KK8�`S�|3��+4�/�<��:�g!�F,)���S<���T(����pG�9�H�܌���(y�B�cM&|=�w,�<sa����x����yΛ˩�w0Ҭ�4p���s`���(��� o(.	\_/|s�A�/;I%�(�5)9~��G�1�.o� p�FDo��i���k4e��y?�����r�kS쏡褳�V�꼋 ��a�nd�K�SR��`���� ��Q�X�L�JMFB�c7� ���j��9�"��iX+��R��23�4�#�-�T(�(�,��,-������甝h2O|�@Mo+��
����_�+uU9���B-g�D�т���Q�1��N��Ds��AP�9�8�^U�A�k�:³XIp����p�������`iC�[�tx�V���}e�������i*W_�7L�����>?�_�i�H�Na�3
L� �7��fA�h�:��o��g:��TE5�
��έ��	+����^�J\�J�QWč�	@�����_�^'6�������j�N�:ѿ
��������x��#M������}��È��a���x���B=1U^,�[./���N�`"�Q�<��UC��N�{����2��C%��6~w�XI��3z��͞]Ybu�'v�r@�/Y��w�㠑T�?Y=9�����u�G������5rR۠K-��N�@њATr$
03Ǥ[�q8�ѣl�L�d]^`x��|���ԾC��֟9�l}�����Qz����qQ� d�l�Z�m�֒=ߗ[�?�zW�ۛG�'y�J�wSb��/���ǽ��[���ؚ�g�K�s��(�|B���=���ꟶ�4��`�t��u!p}�ځ�GKJ���ڋ�C.)(�Q�@	��v������́ā����>S���	�Y�.]Mh	{�C	ٰt���5o���t3̕� 7����1y��U���>2/��W�VgS�tL��"�R���9�NpI��D,�b�EF�е���8Y�pFAM�84~,	)?���
�p�;O�N�$�
�a�
L9��:(�Bh�V���^��^�;�8�v�}�o�N���o�W��G>�z���'��'�e=.ŋ�Trr���ZZ�H��XB@)� �����PluP�,�5�|�~�s���t_��V��}�����G��~an�$ozG��&�;��r5����\�kf�7{��.�+W"8Y��|�M��Q�ȍdVP@�
�����}*[��2d��'ˉ�RVԴx���*H�W	�mo���g�l2WGW9æ!-�#T�Q��^ \�>���t��N�=����dd��&�w�*+BWۘ��i)�'���(�+�ھ|��^��ޏJ^J`�p� )���/,W?X�FS�WP�b���&����S:1Qq܉��)7F�Kk)|���s��3�>mZ��p��£؇��5�i杷��g�O�{�Zf�CsCK8$1�/�z������?��X�_WOe\���d��$�I.�F��dA��}���/ߓ��/۫��B"�f�_ڬ�G�7�I�)�?zl+|~��v���p��1�s�hB�ѐZ�y�~|�Z~�a��#�5��*����G!(������g�����Qy˸���е},�Z��P�RL���[�}���p��}΂Ӗ�E���'AI���"I�3f����W%L�si�����0�o5X ]�':`�&i��@Ejp�Sˢ4S�����p2��h�'��:#�yź��9� ߐ0x3��Ք�ϯו � C"g�ÇF���g �L� N�z$��ۏ���Np��t{;e�l����^�������9L�m6]��z��pI뛬�t
 2����������~	v̬3���*�)�v'�CS�g�Ŀ����6@�U�t�ccz3.�R��XmS���,T��@�]W���w:��6z7C2�6�<���\O�gᩗ�-s̯�⼘Dmݱ�d8ޟ�N�.����)�-�ӆ]v��S�[>�BZ��q���j5�H��`R$���p�JksX���5�s�nH�4;�֐$ � K����_y�������9�զ�%_����\��+	�ή(�5�/�����d��+�u�nne����5��W+`�9��頬�bd�?���k�N���.۹�Q�$|ai#����|�WT��|��t�w�aR��B�uU60�Xĩ�6�N��S{J�v|���6��stW����D~�h�s�no�uђ�!7g���(�!]{p΀���Da�$�Kx���wW�zr�s0;B�zl�ƕL�Ȉ�=���rtK���>�lʸ�8��B�q,A�[d O	T���̥{f8���A�� �(���]��#�0O�E��*8��$����{�y���m�;Ɵ\���l{T�5�̤uV�&@����pC�w���q����~Ԓ���Yn�z�=x��Є�zE��%P{E����B	����O�)!����6t8�����5�2t������ov΢* ���%�� ����Q�v=��;�ך���𐄙P�����V���| SR�����;T���� �`�48�4cd��$�Ӥ��Nⴥy�=�%�_td��q����>�oa�֒NceR,���ݛ�X��=�fMe7:i�Q�τ�*|�'�!E�<��9^^�S�t����ҋ� ߇�0�$��"$���R���p�
ܹ���*TA��d	�0�K AG���%���bU�>� ����	Ʀ�.�!���M ݨ���S�Cv��B�򡡑���}�3J�+���֟`�M[�
m+ET��>�h�R�H�=�� �A�9䃤�)��~ذ��@�8�w⍕M%O�{Z�~� Ԫ!��-g=�%��O�Z�;��E�F�f��%�<|6�0���B���D�J���	�?�h�b=���,�@ܩ�.6�X3�c,���0YJ��kV�O#��_,���_��:�-��9 ���+�>6[��}%���T������Q.Ks���������gՍW-�i�3��B��#\N��k��51	a���P��旱-PEc �6����)Jt��eQL3��h�C^��n�/���g&ԁ�Frx�������LT@�y�M43�$ �������{�*!���xJ����\��L�4�B�֞���ɋ���X�ቑ/'N��F	�0b��{d~��/?&��@�#�E�ၤ<������ӂ.rO��x�+���3vF��M�d�� as��b.¡�O��vuF��pV6O ����\�|���cqޔ䯼{������ 7�Sa�a���-�G-��l�/o�͙W���+���bc.z��Ć�_t�6��<&myR'M�8��C�Sn�ݖ��Trb
�Bu�z=Jĭό�jKj��	�ɹ��Z�\]���5Kf�u��n<1��Os8H��9ނ�P�|�$�o������s%�猏�,�R6�H��q��Oz`�6�sf<��97�#�!Q�<t���>Z�«V�!�ſq�P�y��r��j��Y:A�{>�����O,�{�l��6&���s���{Hx�����g����p�al^Ŷ�u1-Մ�^?�/L>��z�,�z!���MMi��$�Y�=���}(�*M��]���6TW���%�dN������~�X����C��1x��a��?j��}u��i�Z�7��ffw�H�A�
p���V�̊�I�s�+هӳ�J��F�F�4҈�X�b\{�=�JA�w~�b=��b�\Q�G
7���ȏ�F��Zw�M��FSǵ<�oTO���1��eG����A�ox"J����?�R�i��Ȉ	  rܸ�7�?-�ˮ��al:m'��{� �����)\��w2� ��d<�U�kL@l}y4sٱ�[{��p�\xe��Q�?���~V�m�s��k�ީ���)R�"���Qb�ξ��ą��VE;AV���%�6�>�|�OI.�!J��Vy`���lx"��px��9C�	��g��dR<y���K�U�{݌�H��qͻ53�m�	iF���1!��g��Uq=j���qr����Q)�92��S����!&v�dAM�c�p�J�^pF�?ǈHui��+gZ�E/K����1s>c��w*��"Zb��}�^�D@�y�Y���ېҷB�_�l$��,�a������ �>��paX���ք9��<��+y�x���$���s[���U�p7T����,
�����;<��߈Uԏf�-6a��>Kz���r5y�#aˀ?F����kN����^K���z�Ɣ"s�l��hϳ�S��Ln�g��XL-��X����!:{�k���8$��їc���؇�Нa ����ɔ��Y�Ywg�{Q��A�2]�X߃���f�ӝ��]I�]�=��Tz1���4��K<��V�0�s!�Ybl�a�u����6Q��	��;�&0+軖2/����g��R��^?Y�N$�9��䅣%i�D���ƿ�iC*]k#(��g�E�lv�t�fh{E���maT
^��>N�%����{�y]�P�s �nאǫ�v��d��`������Fn���_E�A�>��W��K%J?&S�[�n�q��OF�㣉�MYWzZ�?���o��܉��g� ��ϐ?�D�<P�ʈO�-������KʐQ����a����o*�2}�'�� X��g�0�LZW�AC�W��������&�w�m�J��v�ڲ"u#���'�"�
ąZ���-�Π�5i��;�;FO�4�dZpQQ���[DMv�/b�N��
����oN:��t��Q����`��#��y?N��o:�yld��0x�����!G3�G�s�J��2�]t�7� Q��"K2��Xw�L�;4�[5�t#t�����i��lЊ�*��}�_�N�|�fc���6�� {]�h,w���3���gP����^�qOŽ�Y/��M�c��wЇ]��y�z���b�����N���`���*:p0VJdro�֓�.�yA����ؤ�U�ܷߢ�I1/�M��?�aS`Fl�2��r�+1�9�or��2|�D[��%"����~S L��1�3�)P�+=�zv��[CM6�Zꬓ|.��V�i�
P���[>?��q�`N,�IaË���M�P��O.-����_"��_5q� b��>�L�n���:�]q&��d���S|�2�r��i���f�uF�����h*��w	�))�f���`Q�����6�/��t��D�0f���@mN���<���6��$=x`�����i��]>�eI��W��(LH`��â���pG*	UuM����� )f�(��]��RZ9�(��%�3�55ǷAu��*�8t�ö���L�_쳯ĥ���iMm�su+_%�}��O)�@h���)!�(��s 	�C�������XnY���|�,�P/.n|T�ū��1^���z��>dn%rO�����"I���QS����'o�A��C ���t�gj�4�P�M�1��f����_L:w�3�����r�u�kD+���kLX{2s�s�L��T��>�o�i����*�B��V7lD[7gZ��)AɅ�!0�5��KQ�T�xxlכ�xߤd�'vǩ���6n[���Zq��|�%}a{����d@t�X�ِ��2�.�U����H_�s9���:"S�U�p��ysR�-���j��*iu�t@�F�np������osm�d�Ȓf#|��,3cY���G؀��E�KvDe�%0�<u�-$�y�\�^n��'.b}�T4�j%����߫�0�m<@Ul��c�rF��ݍ�)�Z�ig�'0�}������ ���h����UǙ��ϥL����G5�]�w�=�t�ɫ��et�*������
�b�-P	*��T��<��>��� �rZ� �qV�-�_��"$�͈�0=�C,�j�H�	�0偍q��
p�[���Đ.>h���� )�s��,���N@偄�Q������z�+�3�H%H	�Ĵ񓋸��]�=�Q�"��վ1�����������B3����(LE���EltX����䜵~G��A��`�p��&LHt��ko-z����]����G��$�^n5Ef���u��1���;���y�t'�
;�P��bi�0����![�D�)���;�^�C^CDލ�="\l��0�`���@`�
l:��36�H�Ǩl֛�����Ѽ�8Z��V8#}�J��R^5n�v�ϯò\9��R.�m�����22Z��J-�Oζc�$���n��*I��TI�{ߒ!%��G�N�A<��<O$t +��?��p��p�}KC��gq��g������Lg�JrR��HGs�u��u� ]��������V<����G���D� j�)�G�ݻc�Ұ6�����&{�Bibï.Ӯ�H�1N'�#�x�r��Q�ܥ:��/a�R[�G8���}+�ռ��J~���z
L���M%���D�>�7H���^��_��ȱ��	�����e��M�^�{���w��ߩ����O��%��p;�p��������9��p9 ��t��N��%�p]X{1��0ACb�7{@M��2��-7u�~ҶbV����"�=/ٲ-����2E�m�&� Ȏ��*r�"�X��r�N4b����hp�
\ȧ�!�b�������i.��J9ע������ʠt��%�6�s��zm�V↣���
�Q�,�^+�dq߇<@�C=����r���(ȡi\I��V�g����!H����$����1�$���Ñ�S+5�v[����x7���p���١eq&X�G
�A�^6��F3��FE��4c�������R��hg�.�V?��!�_OLNt����h�.6�>���C��z6j?%ut��� �V�1��8�H��Ѹ4�Y�\;]x�O��^�"m�6��v���ޢv��ʉ�&~&�D
熰���Jңg��3ג;NW- <	����&%�����p�m��rC���I1Je�����|K�I@Z��Q�b����7mV�+�Fu�x����K�Y��֏�|�=��CW�/�Ģ̈́P�p^K�w�ȣ�M�=�ćja<���gp�lS#�pYۤ�ۙ�8=Υуj�����k�#j�V]qZQ5p�ƅ4*D�I��������{G��t�u��i9�~[��)�D���-����u�چ���d]z�b0�P"�k��B�j�	��A�Ct�;)�H�T�}����P���;�z�?������丸S_r��C��
U\���-�	g���L��x��K�s�8�Ҫ��#M���>�0��*��fg]*wa�E� -��W��(�K��@�F�	u�c*r ����J?����4�!�Z�^@���DD�����Sy$샔�sx����Y(��4�����]�m먟�&���"��f
���-�I�R]I�/�.|�����N��	�V���ќo��mH�+���S������i�5���d�a��XB�ei<�bG��L�'TeR��}����3��/gɂE/p-������Tc�l��6��՜NK����`ܛ�m��\%7`�񳔻Ë�� �#������$�_�~��&k�0k�[|����G�?%t����P�5ad8�W����� ��v|�|n>�	�j�qE�����x�=����o@��k.�lW��4f&�����B�wl=��}�&�O��M1ʄ�L�3��?g��G��p���`sȎת�z�[P�s.�ϙ�؟I�@��np���e��³i:d����N��vl�8'.Q5��{QvL�{T�n����8�,����#�\�:�-ߧ=G�??t��%%̶K*�~9(��r!�j�������y�R�w��DЋ����W$je=򩞮���g�2��t3T�	;�R��������k=�����h� �ί󳍴@xsf��������! ���8�	��@�8�x'���:�DdY6�^愗��%7N�]�&/A�"F���^x;�٣�3����9�?��H!iKb-H���<�8/��vg�"/wR�c2���fc��!6^ Ku��ˤ���1haش��_�Z�w���ٷdWiV;S��Yi��7���vN����8��h��Jqc]��������-�~7<�{�$a�?b�$�6���pт6����ę��w�Z�{n'Lj���6"��{����,@����L��)rF�e\[x|�98�=;��2����Uv�?0�@�{`���eo	{���z��g��ϸ�o�i!{z�^D��Z o !Q�����A����u�]�F�օ%�Ĳcڊ"SY-k�1����R#���Ϋ��|Z��>!�G�?7�y���˚�|XU�����OB���
h��!�:��ឯ7��Vk/cnrdK�4�+�k�_E&���aA��5R\	n�c��#j�&����(���s�§ky�\��?���}�B����lXI=>~���Τ�ҵ�M����q�V����58�ޤ��$��ߘ�*kя�=uP�cQ9�ϒ�����׷ ��_�������1Q
z(���S�����	;ę�V�"��7Ո�\ʟ�䥁�b:P'��`�2뙂���ΰ��Nڱ&�˭Qr�uou�F{�Nva8���m"���;��!�x'l����e����w6��w�*~g���=@l���ؿRt����2��K�HbV��~��������ob�(�{�}���y։��Av�¤G�88Qc��x�,rJ=y�#O�!F����Pv����LY��7k�L�퍀p����	+]�����Bp�ԅ�	��@ޘ����O����X��{���������[ƞ�������c#��L����qSrl��q�!-�GC$k�!(��Io��,\͋�9��y�yfg_BKYz�eԯ	��p��Fi���`��@�R�^��[�u��9�+5��]\�<�1��ڭ��y�^���ך�@��k�o�I��ӪWG��<=�jZ:�SnOOQ>����3��w�ݔ	m:�S����Θ�2�(��8y坲�Z}��"�g���&�o7+"f����ժ�T����*`��u).�L��g�g�-�������8&���np|���G��9�f�~�-�h�#�-S�s69p�w��x���U�?�_i� )������ 8��H�
T�&E�Id�Ra�W�~�#�5��;�rم�Ͼ���][������ַ��=�_�,�S�Y�k�0M�ܖ@����~.�b6JA�2^?��䫨Ye
A)T'�Xӎ���ٕJrY���r�>�䌌������ڝ��}ٰ�Y̬T�?�����6��!��l�$[���,$�r�a��l<��)*�VO[$`��LQ�~�(����2�̐���{��(ʐ�F􋳝����e�e��������+&9#���#G�,IMzd���em���Λ���v�}��	��J� g:�������L1���A�?0����8	��|�b��x28
&se)$1���r#!�-g����Q�<J|ś&�d�сT`N��r-�Y�z�r���u}�����o�\8#úJ_���-�`<�kQA�1Zmz�vs���Wf�K7M���)=���?^hs@��2.�1![h>&#2���ʉ��!F7w������^��:�2���6��t%̡6�v���B�����`�6z�MY�mZ�j�l����6qK����R�V搰�m$��J �G��ڋC�`;@�6�T���ۀ�F[�f��)�SfK����گt�g�䆲"z]q�k�$d\#�E���u&� �^|s�G����z�/��IM�T^���/�}�]<@M| �㉟�.���SN�j��7��4�|3�6*L�+izƸ=E�n�Ś�m��8���Z��#>W_&��� ��ȝ3��?� ��+R���T`V�Ko���F���|�,��)�ә/nML�&�02���������}�I��R��5��<p�3.
\3t	���H0�^�n�Zj�le��@V�z(�u� 8�|�O�N���n����o�˱�a.��a�9��D�,��wJ�??�����@\	���~��\�DAa
����4�"~G��˔	��II���e��b) �G��BVa�����w�jd����=��/އ�����~�iHx��MZ􍖿0���h��:��}r�R���|:�=��ε��~u��uW~k�����jԌ]I���%��#4�T��L�a�p_��'�Q���p]6��#M�-�hx���[u��,et#Kl2�|�h�m� \I�bf
�k�`%��+��Q�KT��$lG�E�?�-/�D;O}�e"�!}�&�������u��<��IB$6瀠�y�}��u�j��p����7�B�dpC@�4:o&.�HИR�p�iǖ�C�����O��n�Zy�Ha_��������(5���
ܼ���+��)�	<0�زE�uK5*�Z��[b� ��g��PX�X$c�� �󏿕 q�:Ɖf�+!o���d��K�%��/!}�#��6z�zMm�<���@���ܵ�2� K��@�B���hkQ�j�Qib��#��"�q��Z��Z��!kq��|w�+?z���9�Z�ŀˏ��X�kqij�j{3:^��I�&Y*G��l>�t�A�4 1.Qʸt�Xڜ+�ȗQ֬<ƶt��/^QG�Z��
2�G=���&RC!�Z
�&� �b�����W��BָN�v!% 0`/�L/Ξ���So���~��r�t_�v�B xqŅ��Rm^�T1&���Z�j��@�C�&�17�ด�7�k	�cJh�N��_Ҙ�+1B@dRK�	Z���bf �U'����dna
5-{��(��-���>��O�j��s�[����3�Y#��:\o�V�T;�|���㘂6(�\����P\HT�Tܑ�&����H�v�r<-�XI��|�� c�R$�L""�H��]�A?�U[��'�87pɍ,�� �v��L 2U�R�P�Tƚ�����,|P~h��|cn3�w-�%A��(����r�����Z���ANXk��tL5�Ȩ�+<I��Ri:Пab=���\]D�A7H��mm��L���Ђ�h;E}:bq�h�ŉ]���'+��ۋT��y�<��;jÞ�G��5i/fP�Ft� Ҿ���O4KH�O���(��׵�:`����w�,ȃh�<{��Ұ�(�D��V�#��9�B]Fs&���t�Z����ƨ��#�W�D��a%J��3ft�T6,V�|=�z��y12(�)�圾ٔXT��R��>���ıa뢷1_1���J�]�<�Ľ=R<5�[��A񜒝��RL�m�b}�̵�_D��P%��'��/�����izQ5�7e����pw~}�#5�]��oӚT����
j�:Q�}N�<v���bg'�'xpˑQa�R"�v�G+0¢�&�:�jN~8�Ữ��q��%v�{r�)'�-���d]�+����T��݀����� ���c?��ZH�c����8�h\A ������q~u�[2�ZJ�S�{���q 4����Fkjo�3�+ލ@6��>���N�<̧�~��a"��1Χ/+w�� _ў���C8/u.3��CO7�R��4��t{n�v�������Q]'͢=1瀔���Xɫ�ɋ�[(�mK�v�qo�H��A�?�m�-l@(�C/ŉ7���K�(d1�l���غ�2ezcߨq*!�����И��b�:����R��z��TP�J�N?��22H`���b[�Q�`��T�X���\_�O?O���YF�s�CS��q�;+��|�/g~9�l���ԁwd�9w�ս=�Š�"�V�q�T�1�u%Z��0Lj��Z�c�����m�����J�����sj+J�~�����vs�����;t�;���5���f/��qv7��gRG��[�ֶ������{z2P���ލ�Y��@�J�`���8庐�
�����1�f{&�әioC�����1�������  {W��ٵp��m\��[�,��[(� [���<���� 	�(2ȁlN�����`lc�_ʧ8S�X������m��EM1	�Цv���l����ي%�l;���<�{(����m����䣒���i��kH_�Y��P��40
?��U"$�ޙܻ0�-b�Th�هM��j�6�}�B '��e�aO<`a�3Lk4�:��월v�38r��w8ĺu���i�4srLN���iuQ���_�����V�˺KH���v�T޷e�9�ٰd0�dL�N��P-�4�V"TuT����B�o�SdbM���xfe��g.Ξo'7� 	4D_e��Q&�N�H*�:�&`лa��H��r�b�4�#a�4W�C$MxT!0�V2(̞H���Nk]p;#9KCA[�?�MD�4�Vl8�
;'�ߵK���k@T@KGt�xRn�s�%���3_�A�`1P1M�s�Q%���|��Vҷ�t�{s�IPȬ�����}мd\��{������K �;>��=�1�KUTz���3��l;�"�(%���5����:��́�Pgg��G#����h�p��x���_ƾ�|Mf�� %��o"�ُs��1>x!W�D�ǥC��m>���@��ˊe�����l�<�	(�lR0&1j�Yr�����\�:�C{�1d�
��7��S��;f3|h�]�WŻ�ZaDN`�v/�tRx?�z�����br��������+~����PĢ)I�k#�����='�U)W�¾f���<�!A<��*,��Gz����>�j���4���y`��Ar���)I^��ւ�I�ݿE��sK�^�G _���@���WLJ���lV�%.	&so[���k���>[r�݅��� �`�Q�6U��D�<�2�a�V���� �Dy�ӎ���qW��d<�f�ե3�|� P�=t�;�4ۛ.��l�V�E>mz�~�fG��:���N���b|�xq��V� ��I�.#b��K�n�B���Ȋq�bc���i�?OPKr<깭��ϸ�{�LY,~�=+_HIu��?=㓰"��/�YZ�B]���0������Ϻ�V}?b[�־t���[-��֞��7�@_��@-Y�r��0�@gpgSY�aq{<b�W+/xp��LC*
�&�[i�Ď���w��>��Ø����ݦE��l(��[��g��m
���]D٫=R��S���'Ovu��Q�c�ݽ���kd�2[�r)2oac��
��zU]�Q�G;�Qy��}�:�O��%�3��^ȯAn��������VZR�Z�۝�cᬘ���s�:1͚��W�Б�<9���F�B-��+��ˆ+n����-��ybHʋШ{��!�!a����E�^��}{�M�p�PYmmTntW"�Ȝ�{c���~�-q�s	��4��E�?���o�vU�,���O�����p}�@���n4m�{�������ֵ���8�K�Q�X�Ol���B��3:��x.����(��)?�!UYXm�j�I�{�i���������66���ə[= ��� ��.4�����B�9�`�	X���e����b����J��;�O�B�zg�)6P|�e_�0T;��k�y�h�p��1��.�o<�Y��S��ɴR��"��+(��+E��l &�J��7X�a2���}�e ����T�C�Bʤ
%5���^m�x�15��h�P�=��^���`�i
�w��wR�	j��M�>r�m��d�Q��ol�-,�R�=餚܋�^�2XɖL�@��Xt��ş�J�Mۄ���Z����Y����i2eh�d!��8�j�)���ar����o��w�n�O����\&�,3����#!�lny8%B�����-����v��~������@�#�RB�$E�j|~����7��x�{:m##!E&��6�d����ܜM�/����Qk0�����:�n�2�y�ime����I��^��{1����2�f|Ֆm�������>��ʡyG,؇0c<X�]7Χߌζ/�4��[+��{�v��U�G��W,�=�����H+�b�!!�vK��`�!NZ�@/5�F�Tg�':����l�6�'$��"JR�l��V�.� M��5Z�q���&��[b���+��ꄠ<�V����ؚ��
̋0n��1�*(.��r�v�<`&׬P�O�dV�'l��v��Ӫ��[҇X�a��K��>�:<����a(���J`�Od�g��;�+�c9��M:�M�a�N�~X�-�=�����d��Vɋ��z5(��;��_m{���+!e�zg��0��&��5�$qB�V�� v�*t�d�!E�R،����b���HA�ld�of����ޘ�*�I�c��p��\����Kr-�G$��-��Ґ�N���~�D*�X>O|��9s��0� ,��3��'�h ̹xl�	A}C|m�u����ฌ,a|���Em���dn@�q�A���?�R���z��f&]P��^8M4��`���눋yU]A�hX��mz]��D�\�9�=X>T���uL�!M�B�b��g�'s�T�pՑ�K�N�[��������&��q2��6|=Z�(���aK��ֵ��_'�����"��|����2g0r�p��1�cHHQu[�c�ݎ}q�p�����빫�����ޫ+R�c)q����j���j(@�@ⓐ>�"X]d�Y�Z�����/�L��z����� R��;�bЪ���NZ���{�4s�9�U����JLL�Y�Q����>���"M�e��NL�5C�	?Y�
�,� :���Њ9XJ�ߕt!-�1C.���Q���ްzݫ�����=tC��}L����z�D�eC`����T��4{f7�V�y�.>_~��GLW���H!;`��.,�N��3Љj"���ʧD?���G��Ư/�*�K�u1�y��3�W��qf�N��p��������x:��VTJx��d~?��������sE����`)���i�;�a}a�k�o�c)}�B�Vm#�B*�"�~����E���- �]g��l/?�"?R�@�<$NRu�s浓F$y��F�č}��+�6�[BV�U�± 0%Q"����+�DTQ���e��2�<eA`�=�M_�@ͧ�IL??�������.�V�L��1������%V	��'2�H�h�>t��h��#f�_��?1tB�~'�\��gO>�D�
�3o��S��j��X��߱�j����=1�+�B�R�����O��d��P9�vq��P���x�
b�.lT�7L�%� )�P�Js�t)��^JR:I��`J���A�?vi�����_��'#o���8�ˀg2r�Ou�}�;��L���h��5&��Cey҂W:�7;�O�vn<���k�+"��K��#h�U��߸!oNl�i�ΙT�H���?���)T#v��;�O�9z@��7�1���,L:pb�?�`Ţw�L��]�~��R2ک"�*sQ8Qgm$��+��{��3y���)~)��Y:�,9�؀�"Z��J3�`����Z�=�s.a�XO�5"�J��M�y���即�}����&�c�����M (h� k1��x����qƢr�<�{)O�o.R�Wo9Wq+S|m?<�Ʌ�Ƒ"��ʿ��4$m�wG���B���y����8�9��΢uj�����-�3܌��U�c/I��:Μ�9���mH�m{AS:�ϹO ��Cx�G"c�b�m� ��Z�W��!�`ܹ�b�[M2�$0��g���7٦�J��
�އ��� �6I��?P��{[�_��t��fŝ[����&����nA�a�i�^x��5� �~ 7�>���<Z����`���Xzvb!^WV\
�`l=H��'�m%t��Natz347�u&Pg��
a������g<PbX�m�'o1�0���(dZ{�\O8�+d��@)~=2}R{���`	s3m����*J��,�U�������\�
~2 u}��{?�5 �-�^>ֵ>h����Z�|@.&w��	be���Η�_�Zv��e+_q�S�ە�u�ϋ*í+��M�Z�5�y�l.��'#�-R ����qu�lD�W���?\n���nX��)������gk݉ʨ'�TW���
HlQ_M-��	�隆��!tJ��ܲE���Az�iz1��3��6�'WW1c�܅���x�X��h��4����P�%YnB�ϔ ��M<~��M���g�|����IN�Ѣ�����2��W�Q�o!q���F��^*GS�S��W�p�bH�I���Z��ȱn��:m�3�pd��2���
u|V��O8#/�u����W,���J�M��!ؓ��eX�q�_�+<8?��< �f�<NQ�]fZ>[#��1KY_��s�������ě;�"-���\P�b3��x��<��u�0j_�;o#!����S,/:��z�Y"ޢ�k�6�TР��� �{S?6���>b?yly"u�5m:ڈ��Y�5?(X��S�j"�e��G繕9��
ip6h��,&�dZ��.	��x�=\�� �']�t	�MN$A�%�(��� �fO�Ee��m�Dn�y�\��=�����m�����|B��Õ!=F���݇�mR@���O����}I�rt���=��%���.�J�6>/�Z�g2�}�V��/f�H[�Zb�㫦0�U��e�Z�\����4*�#�9MO���hf'7�:=�>���� ���C;[a�#H~�s�i��}�J����T�30v�졛*�����5� ^G�r�~G�E�=-�L���a���딊�&G�r�7�{��k�Z�$���S$���=w'=��58��$�T�U�W����o��P��Pq3Hp܁��{�ﵝe�*BA��I�`sg�?һ� �M�ڜW�5��41Qɢ�@ܜ�� ^�T1�~l+�ÿ�%��i�X��� =6I#MC�w�s�J	���ϖt���wu)�5�V�����(i>}.��j��$nQeM�ic��F^WCL��m+��h��[�\���^�X�E�\KCcG xEVn���ne]a���?�Y%U�ꔈ�m������K������xV�艻����O&��=�;*�|�\�s.rA�M��	���g�c��O,s�r�XD�� 4[�$Y714sY��M�����*m����#�m��<Q���;Q73M��P�<�v�͂�9��ޠ̢��lszX�f��L���X w��0��!���C�Q�(��F�mHl�b\�0<g���h��>ޚf�i���%i�)4��+�>�[ȧ� �Ey���H����-�!���}}?.��Φ�vJ��g�w%�ƻb�K���IӖI�����cN�V����A;*��N�pϙ�МP@- ����m�c_a���:�з#���̝42}e�p��>�7T=���"�9�qA����hq=��GEKXH_⒓rc3��8Ek8�83`���/�!�rg�5�I�N9^��1�IDw��`/��]�"�w�jtA�ś��QM%"/�:H
�nd����:,��Ά	.��7@�w2�9�U7���w3\E�@�|y��W������ߤ֧=��i]k��M�{8D�_�����j��}t.	���g!����	%-R
�` ҹ>q�f-���þ�,Ĩ)���v�=�B��ן��Q����_JC���pK]������l]ܥ#r�rI�%�^��@�O�ǴV�_{�n�NH���}~��,�f��-�y�c��>7�����t�b�� �Ԇ���"�N�c��a_�/�
g�7��_n_w`F=��h�+�O��Ig7��q��:�aֳ+�ǳ��F���Dj���З�r�K3��brۃ�O_��ޗ�M.َ�y��8*0�$���'���W����j�)(�j����e*[���~�-lʔ���#i2/��+��p^�Ò,HMi�>��I�j���,9��]��ڿ�|��M�.�^Z����zO�04:��we��A6h
#�� �"�Ͷ`�%=��7��K9�6�V$Y֤�!qHO�1$�r�"L���u���X�zh��{Q�F~x�VyOB>}�L��yGw=�4[ƭ$��5�X]�����T�+�BR�/����d^�ƣ��"ՓMo�ߨfz������e������9�|��0�AU	7�����KC ���5��d�q@���2
.����/��V�wѥy�H7�BX�8��ڛ�zߑ�����Zh譏��L&X���� ��8���=�m�Iv��L�F1/E��f��~����$�89&�˽���@�٨q���O}��T�/e̛�T�u��7y�]��I�%�m�i�g��pJ�"Wע9�LyswF��.�M�4{�gUQa!��|C��S6��m���8�fq��q�3���o�aƀކ�s�^<Qx����,.����KmYl'
�y�P���?%����U\2��`��CWaDs�O(+�@��@�o~)��3��ܳ�F�W�*,����%�0�r�E��t�'�|WѳǼ�(�%�S�Km;�����3u��Կ%�_�N]�}�I'?O��1�B��eom��j{���d**�M������dOL�'�����A	��ͮ��G�H��ܧY�g����q�bwn{�A瓈����B����}�������@�vh�3��!����#j��V����2�/�����?|�sX_4�d&Z�癹F�]�t�U}�%l8�n�O��ɾz�Sw6�3�����H��%/r��Q^]�x��D]��s����Ipj7�~�Ҹ(�<20����s=EH�Qt;׸kOՙ#�V7���F�3��)�I1��.@��~����?jKg)T_h�.L�A8���+�uG��Թf۰R���p1#,���{�M�e�R�j΂ܡU
�u�x�!V���uð�).T������ '?lN.)���scK=h3-A������K'�C��br�(�
O�o�NP/��ީEtZS��_�?����-�2ve7u��=��� ��̄�
é�N���)�,�{Ο�m�X��P���bۿ|�^��Y����(��9Z�[�5�8��Ѥ�FXW>�[A)��ɵ���� �~��ٺA�n���ꠛki�A��x�a�u+ �i4���3]49#-[�+{�J'HWc�~|�+B�\�n���Zr<��U%~GǤ�<{��t���PF���R���M6K8΁��z`��@�������m�&��}�r��>0��e6�8�\r����/��œ$jR�­7��3����b�찳����W�TK�j�#̞l����� {ؙ�y� �U�g�Jp��15�D14.6g^ 4Ùރv&7S �L�I~��{����*BY^�k��0���0#������(�Y6�45;^>i
6�t��P�{IШm21U�.$g2����B�O�Y1/��p2vU6�}�W���#��&IF�|$��)���V-V��Z��Ώ���8�c�|!�:mΖ>>~�i�2%W�7{�z�$��!V��sּ�V�0��
-cA���@0�qbA#ӺD����H�,�ʀ���1N�3kx�b��C��O6�A��q�/l�c,���q���ijٞ*�u�Sڦwq�r&��F,$`�q�r� L���e���VT�_ԉ�(���F�5�(`�B�B�&H����@1��
�f7qx3��D�4+4���֒�!¬.�ݺ6���r+L��u唸 ��//V&�����M�����'�Ա�<f¯6K>"o�13�<{�8%�r6�k�2+`���d#�r}�\���y�a�����d�x�CfA[A(7��b�w��ؾ�����MUw���}J@�*`�K	܍ŏ��]C���Usk��8ml��U�c�����8c6�ߴ�QS�N
��m�`_µ�V]�s1���g�4a�H�h�r��k���!'��W�0+Ť��ۊ��[<�`Զ�JA!U�V�̮Y}�O��F�r�=).��wUЛ�lg!\z��T#��_Ã�eitÉϥ;�i!��X�W��!������Q�Z�'�3���A�y\����4α&�O�+�%cm����46�O �<onr¢~�U/�o�j{L}��,A����Q3��V=�&w�U��=e��~�0ץl_���O� �lq���'K͔��Hc�`/z�:^1�ۇ �ך";k���("��&��_G�x�u�=c����
z�ق����`�����B��h ����?��Yi����ц�Ouqf�el���M��j^]0Y]�[rば�l�	\��/t�S��~pUL6��=��2��D���[���:;�\������B�MX���0N� bX|V\>�m���l�%M9ș���J�p��u�>�����6��Û�ܴM�B�il��W8a?fW�tyL���4=�`�C��**�=x9ƚ�!��S�QM���cc� �2R�"�)��;M��-m�����V_&ɷ�>�F!u�=YU�.�tڱ��}~�=,l����v=kk��F��)���Xt���3@ڮ��ŉ�G䥪*&Ǡ��E��mLaA2����^y�g�������{��2f��4b�H:{vw��#���h"��"e�!EIx�����bP��i$ڙ���Ct�Jn�|�,	��Oh���uYnl��;��5ڢ1���k�zϳ]�>K���ޜ
mn�ӵ��1���������Y���~��x�߸>f��JEb�C�W��\s,+r��?e���ҶC�f[�l2!�v"���[�^%��e੅���!J��n{۟���q��d�ٌȋ?�6���]m���-�b�$�̨����V}�ᾃA�~s70�k�)!x��,��ɻ���5���I�����r�4�V���_ eS O�Vk.x-����^�$P��٘��T0h��&R���~8�3={����+3d.��.�l�P
Z���s�e�κ׷x7Y(Ќ<��։���H�k-e����$å)W/pm}]ȓ��@����98�Iʴ�A�۱������(`T)LAF�~�**�`iq ��Wy�5�x�7�G�Ĺ�cR,��`���zJ�����n\U������a�{V��٫U��Zp��ڢ�; 	��#����3�}&n��9E���q�{/c֋��WP��eH��&Qj��6������[�p�z�^�D�9�/�ׅ���0^�	�Ʉu�)2���y�y�@���Eu�[)�z������)�j��P7�hB�z��ŷNR;�����f��`M�.�5i����^?�6���M���6�	�f=�F���u&����S���4���Rx�J���G��_�o��uTj[-bigv
l��&&�So�^��	q��J�-����uf;���^kj1H/[::H��4��� 61L���gC�2�-)-ºё�`��x�ҥa٤D��K���LSL�����	`$�������<��,`F�φcL"��&S��.�I�G�U��A?���HH���8\�z�̯��UV��3lyt�@z�8k�r��?�yP=5fYqߥ�$�0��v<��=�� U�_��[Ǖ�Gn�x����� �m�rzܫ��D�xc�`�V�.����?����@��{��xW�%�gJ�X��'Jִ����[=l�!�eo�|�+��P�S�+[<�B�Y��"�pDX��
B+�&�%�dA�d�x�b�\���~P�G��9��oc �b��u 2�X$Ĉ5��_��E&;��v���D�d��&w��}O����3��4evͪ���ӊ����m��`��Yq���Pal�v��Ө���wL ]�������B|��h�g�K-T>�+����`^Ý߾0���	�n�:0=�Ëc�Q�����x`hh�O���h��<ݚ�_��;S�8��ߜ͡?O���'��;~���
�ѥ��7W�Ӣ�k�����S
V!_�\��ߺm5 NC�R��	b�fi7 D/�67��. 0�j�s7��b?-C�cŭ��d2"��u�ML`%Th���H����� T"�4Uf��ēcfuG���3�&ԏ�X�z���e0�^X�5�M�9g��dn^;"?Ut���Y�!Y"�V©�M Gn�+�����\M����q�`��RK�
!�G�:�r �O"rGT/�n��޿
U�A&Ն�:(UZ3��uܾ��w���:̐��-��y�i����h����M50�J�a���^� 'қ�Cvb#����>�<X&
��ը!Ԗ�_��P����0�'� �����H���>��3r��^|�4U��3b� �D%�f9���g!��lKnS^�,f���-+���]�vA��� ��	wY>��O���g��/�&�[$~���ʨJ���f6[��1�lOp��M7(^��^���qRoX�"�g��	[fg��sH�h/��uNm�{�ܹW���=�F>־s~����~x�|�d'�d��0*"���r 2� ����ʄ-YleQ�v��c����E-�������X_�Z��РC�^�՜�;5�ᤈ3ׯ������.W�7Gcl+E��3hT�n�c��p�w��}F�?tD���'���&�s�Z��2U�=?��Z{�?�觑��2�p���h,V����LI���tb«�E��A����G|������A��E�����:�p���IU��Dr^��N[�]2:�b��=�U�M��
���*�-��a����Y]�/��dG���������h������Q�,+�����:d!�@�F�v�ȝϘ�d�e��M��PЉa�Ik��[�󧼹il��8!�&��_0+�� �^{n���N҇[(x���s <�x��f���׉(�H����mB[mL(���
�|�5Tg�h�:�b��=�F������)�q��U�!n�����:�f*�ja�Qs���A�#wn�[��|g��p�7w{я��7��$����%�'4$n斮�p��8~!U�e.D)�SR\�r������|zk�B�F\2�l)�����vBQ��!b i�N��V�|ǈ�Hj��>��~�cnd�(!��+�%([���|�AQ����q�gYy6�� �u�A;���r|�K,r���a�16�D%ޘ!�9r��$��}փkr�t���V����低�T�n���zfWL�0 g(e�Й�~H��jP`�~�բY���u������N�R�@g�F�r\�H�_�C�Ǉ����oί{{�I�����\x\'FM��p%j�H��:4X���w��������������((ec��0�ɏ%V�T6�(.3m[�rcZ��������G�X98�'�A�pZ������h�,��*A�3�_�]bM��R��C�:0t�k����A9��	K�Z�.O _G�ޥ�Q>���uy�:H��絠3��wRc{~�u�P���`�|	c�b�
E�-0ȑyP��29������a+�҄��./a�He�R��$�/O�P`�aEc,���B�Y���N����:��˄P[�y�Hؑ��-�|}h�/�4��6�f��B�e%���|�r��Ë��ңsD�+ّտ�j���X�gܼ=�z�xe�<�X"�-pȨ������X.��zP?�9�xI$�Py�=iP��n������@y����_�~����<�n��p�͉ӝL0��]�xo��d7?���9�s���N�R�������<,���Q�����u>��{X|��}�����C�7���k-P�~���?�wE�ޡl]�ς�7��p�pƻ���&!�8צ�`�fe�i�M!$M�Z�!nA0�%a����Ss�-~`=��#��T��	3lb�P�$$�D�R�v�Wĺ�5�H̟x�x��t�g^%�������m�5!�{�����7[o��.�`�e΁�B�?f�Q@�o@H�U�LAw�T�	ٰ�J�T	���u�>2�c���@H� |����
 o��b�N_��卻@��y�^%"��NM)N� ��T2�{4B�G)O=k��9Le�W�X�R�H��ww�~`fT}�j��J�T���`@��,��t��&�Gi^�ve���E.	ܙY� ��V�OƖ�ţ/�gd�g�������=E��XE�~�;�n3e��9h�����`qB7��ޣN�&m���[��4�~�V����9[	 +�Ǧ��-]��$����42Y�H��,����f���Zt!A,�NC`㰲%��#��qn�X=tQ�D��}��1V�`�ؔ�q�Y5r)к{Y%)��T�0H�pX�2�f��oƣ��T
/SB�WnТkL1�����Gh�,��#�ȏp��Z����c�+6�I!;A�#��d]
�u͇`p{���Y�`.�ي���A��B
6��c��$Bo��:�fJ
�Ui�O6���;��p��P�������5�q��Q#�E�7I�R�[7O%�t���q������/�yA�Po�dz/�W�>ϲ��:��Sq&4�]U���
e�2F�%��V[t�k�eF�-�9`�24�����\����X�>)FF���+��^nC�gO$�'RE`A�^�ze�gOwu�zO��JpKU��BrR&Ճ{�}�:w�A�G�tG�,
�;�e�Ua��S䭙��BxvH�N�X����i?]�>goγ��d���T�=ƾ�T��Jۨ�zu$�o,%�#ls�5���Zck��B��崡	�3����LX�?��nR�\�1��v���R9Fas�i�E$�m�]?ҍQb��T:_�].�@�(a��LS�R2U�������ď�߬���˼���e����i�5c	.*MlT��/�� {���#L��/��\�N���ɇ�=tb�sG���O��8Սm\���D���-�u����ʐ��T[t�5:�ҼKWJjO�k�]���s��� =�����e)�H�,�g=~�/� HVǒ���Q�H��M�ݦz�8ؔ��Ĺ���V_j֊�1 ]ֻ����g�� ˊ/j�(y�h��(u|�${�V�x�0�Bk��h��Eqq���^v�G�O��%aS��)���zo��ж��Le�%�~y���b��i�0�ĵ��T�W�?�pʣ:݁I�]�Y���<fg�=����Ķx�N?�Ng���X�S��0�<jhң��8�G��Z��B,G�� r�ș�'�r����6H�����^!U�b):y�/���=�E���j���on��{�B4�u-���Q��vL��"Nr=�@"jG.x[���,�R�nk�@89�������O3Cu�4�>eW"���H�w�z%�c�;�y�+����>�v<���1�:څ3�YĴ�Ŕ��dTiE�Z(��1�IGY�Y�+H��B��X�Foi^���3x�	9��%d�jc��#m9����⨴᷐���L��S��h!��u�]L�	��}�VmU��(䵼V��h��ӛr��M��7LSk�Fm�a���)G ."�T¨�J��>�Ս���m�O2�n��@�R�^r�������Ŋ�N�~J N�-J���F�z�X[�Tp�	����m[���D�=�W��j�k�`��tj<��'%����>g���� �4\B�S����>��0U���$���#�,�&�A�8@>�C��WT(�F��*����0�P����;/���͸ZՌl:$;�~D[�uv�?�nn����c��|Y���)�A. ފ��s����jS#�UBCI�{�Y�ë����O�<�KdlT��C݌�H������E�"�y�y!���jKHd�r�c�r^��T"�ջp�Ą���k�6�`ćQ��5�;2* ���w���ɧ���;�c/������X�(���
�#q׹Tr��\��*1 �A��z�a-��%�vH�.W�C>{x�̬3P��OڵA0[��M�)�V���?�Tʜ�̅Q��CSӝ��:��_�2��b��wI��m��k���ݭ��5��p(V����|N�C����Np}L+�ᷯ�
2����<Z��\>UZ�Ꝭ
}&zk�Cqm ت�bZ[ �u��������z�������2g�g���Q����E�y>&�w�����G�Y� 7ڡ�mӗC@Ɠ��çL�̤�`3�
\�!b!F����l�8��M9[���W4�B$�!�F��J�����K�< T$_}�y�s���@]���*OP\0�}��z�ۀ����ɽ.pi�u -�I�k��?&(�����kKCj]��-�%5Ͳ��iP�m1<Wȷ�P*��q���Rh�Zȑ�ո�Ȁ<���/�N���rFo����Ȁ�OM�1c�֦�TT�W���D��^��2S�(^�$b8f��KV;��B՝K1J��b��M<A��,�hf4(��[O�bз	{�A��^���g��:��H�����L�;]� ;���x �7��>�t~���19�Wn�M��H��\�󡔢�'�**w�(x���G(�M��5R_��'L�nМ;�m*�����'�k����U3������=o�ڏWv���!�va�O��JB���/��c��)����w5�Z�IS�M|nE����R�b��O��Q�����Y0�C#�8�2N�1����ح�
���YZ������	�_�d[,��w�.�)F��3�j0]K?3(��9��.v_�M��;�&�E��rI��Q߃��B�@�,z��x��B����l��B;���M�U�O�vTOV/�������3ݹ��0��NZ��z�J�(A��ˋ��R��e��L��~X��O"O�N���R�a�+��?�h2΅���u��ᨵ�0�'�]HK�0����x���ƅ�TA��3�{�㋑��mEx`�;h�i�'�{Y�<~�,�!v��RK�:U�'���@}�yQ=R�Z�^�sз�z��m��ڝ0y��L�Ҷ�!G�?la�3I�.ie��j����^ɼ��O�����L�,b�%�_���j�;](e�F�R���a���ձ�r�DhF��g��)��b+��P��/%�^0lό4��qM�<*�B��4�a�oU�� B]�`�Q_��:^?v+͙o�W�p�|UC��y�6�%�4[��m7�n;ʟ0�5;lז�1T�B����/b�)x\�vhA�Mmq� �d�Շq�,sE��	9�:h�3|��"Z�OZT���8~���P+p���A���6�S�ʆ뛉!��즡0���Ե�`���]��2������zB��(?���˛�r٢�\	����FQR �`��Hѱ��R�`7 �s�y(�ǲ�Sj4����埴�C��{�xɳbXg
B���b�th�uQߪ���n���ᙰc��Hwx��`[xh�Đ�6�*��`�k�7EL@êV�;��b��FB���X�i�!�)p��
3���'!��a�E+��r���¯�X��T�S��h21����嵺���yх���A'�8�WY?��g!���-�@�-&��4>>�8.�����%yj��h��($ֿ'�x��L��\j�piƏѸ@��]������&�����3����)�}��bZ6I��c�����s�j�zt{.��{^3<�C�\���ru��#��h!MI��d+d���
W#�8�i$D�pH#D���J�cەq��իq�����	� ��HjG���7������_��w����cȜ�716ܢ��K�̮��8��ZL���
̻X�{[AΆ}j3e5�9��5�7���PA�G#w�?�����^e�%8@�;�Î��g�A�V|�RqD�f�A<i{��F}�?��"��>����a��{��Ǳ��Ʉܯ���g�D����&�a�:>�B�3#�ƪ����د��k���7�>"��B���GUii�1��ݪ\�](	�;��T���<@û]��G؜q@:�GeaY@�A��53���K
�h!,�w��9�j�+�0�`΀��Q���k^�Xi�o�lN���Zсf#!����%���}:e�O�K�nѢ�N�m���Ft6� o�.�c��.���:�⨘��p��5���2��tK(g�P-����?�,��z'�U�/�ytf#��Y�B�B`�]����H�ɱ�i������F'�.��u ,S^��ݒ[ϊ�<	f�bn��N�ꀘ�@���>��~Dlu�2���=�n�n�/�ߚ�<b����/����tS�TCZ	ln�dA�bF�Q��7�T�dw{Τod-X��l���ܼXR��wT�eUM̳�R��i 1U�@uN	@�2z>�C�dx����~�
�L~�q�pM�Z��j����E	���+j�U�*U���P��'Wu�������!��ލ��G����i�g�<��%��o�Ͽ�*#~Zh�u�.�*T T��n�~����ͧ�˗�t���,gTI�h��O�@�z؁�u7�0�8�~p���
r}g�dX���"�>�e2a[ݚ�c?�紃�w�@�.xqua�w�|�r❀`��XY�*׳}����*_�F7Ĉxr�jg�*��m �0IO��:ϕû#)�T�A��_�<ԁ�Ⱥ��A�j��j���jYt}�JIr�o��}Z|̼V��<����X?�Tݛ�,�b�7ഹ��Dt���T���B�љ�R�eVإ�3��|��>F<-�ցe�b �V��&-�{)��<��]�Ch�+��K�x��]��W�6��cn�1"�+�S<�������zN��*�_��*P���������X�����X^;���X�g���DlL�r�L�h�0=���u8n2ay��IY~�"A�1#��Q���K��	���)�����A��ek��޽�p6G�����w�T��^��̲����9���&�hPRR-"��(��[9��vܲ����s[��o��F�/F��\��F��.X���7�z�%��l�Ήi�������'Q@�A�����-
�FW9.^�M�8n��]����*���TV+��r�.�Hvb�}��
�V% �
/���S�Ad����d��Mr\��{��羗ۣ7�{z�]�ѥQL�\,9�I|�m/h�e?�+?��7(+��?�&r�c\�����]�j�Uub���Ώ#"����^���MF=s%r��o�X1<���A�͍ ?���<O�x�*LQ�l��J��C�r#iE^���&�P�(P�����{�Z���2�
DD�d���Y�|�:z�<F�?�Z<�Ku�"W�0�F��O���/Nf\{�4���5�������b	R�#���7��X~\ǝ���^�eIm	shM΀�b�|T@`��6H���h)�a���%�(X��ߙ�f=gu�Q�	f��Q�|4�\]O�U�ԣ�iy,f��˪nb^����D�=۔|r�i��sJK8�𩸫��% ��o�.nu��}��n�����\�H���u����8�c��?X��l��������Fj0%��|���tRA��a����� �o�X�l8 �����p�����Q4�mQ�:���$b"2�����P�\�G�-D9f�����W��F�r�P!5Mk3��0�՞ܖ46���3�����rY~�y�r�KF�0�?��r ��:Le��l�t~*~�5��Z@[�lG�P�s�<�Oq��w�a}�;	<^}�.�~���%�NV�C<�nIq=����t�?�g��&�/(��ϕ��v��`8ֱ0;���ز�Ab�W�T��}A��W�����rꍥ��3U�0�5��=YyDbĿ=ã��V���;�G�l��JD�
��� ��=��X�����SS�m:3�v,�{�������N��^�b��X�5��8���&�K�>Z�I#��Ymc�h�d�U�1�_��h�������_y�t`����m�q8��~1�;��t1-�@�`�j������J�T��O�w��\��?��~͋G��P:�x�e��"��۶�q �xh�0o.�u=�㑓e���V�������O�Y��`�"�x,�h��!Q�L6Q��x�X/�w�����t�m:A�W���eO<ov��ҖF>,"�J�h(؈�꯫��T�>1�f�v������}2(�{}��V��l����I.��n�&��q��gT�[,��8W^�X@ݡ�> ��V/��t`�"��j����oe��Dw������L�U|Q	�s��qO"�cIHn�
�s����I�⾷�8���q��%�:X�����z���Bd1��R���PQGw��)	b?Z���}�H��ESK���"=�o,����!*�@���+�U�f���#x�Ǡi	!�'�����u45�wЬ�(C��qQ��M�R%������,΃Rɵ�FfJ�F'/(��߭�7��t�!��n�ڝ�xݿ�>��Z�����ܨ�Z��֐���� ���,�+,�p�{hqU��ԏ�}��Z�ˮrEa�@�_����d֦=�B�j��a�~�5C/�5�(T�5d4qP�ެ����Mb����5���\y��;E��P�ꔘ��爈�q�U��,�3I��R�^a2�e`ڸC������K�o�?�R�6N�Y՚���T�d^Z�ʓ����|��:h��|NBЉ|J>q_bG/(B�u�P<���NTl�h���O���6����.����:{5�C�i�D|�@T�S��(
g��B���E5͒$p��;:?(����0o5~��lb�` e��qr�e 3�C�(�i��|O]�|��9����o� U|t�ƴo�0q�a����+d����jYG��8�/Tȵ���ݺ�I�B]ȭ��*�>�[gyY�C9�?c��c.͏�����/�R&��RF�����j���`��~"1�xd,`N�Cy;�[u�"�j�3��SO���!W�jW;S���|�M7d�֎Z��t�����E�8�� T�)�u�ql]�eB��x?�0.�Qmդ)��v*Ĥ
�ϋ����ۛ��E�Z��ө��MN���Zc`��2-s�I_��J�B~��<���:�V�֛�s9�]�GlA�Ŷo�fXt?j�kE�S�h&@�2�J����f*q����؅���b�z] o�{�L���E�h���kq�F�J�GNu+��!�=�]���H�+��+�{3�p��ȭ�BEkP��^K�SjT��[Df[,*s��P�L���\爒�r�ԅP.����*�:��ڏǥ�h�Q��z,�)�����Თ��?�
2����`kna��2�'��/�Z~"��v��cl�\̏����}D���:cߗ�5�S��4��.�,Ҟ�4I_�*7����䒗�~mg�*�5�L����|�S����^��̶�����gY��:@;7�ʽM�u�t����1	�u�Z�̛'LN�g�+��������?}DW��}�p����2���b��mM�
L*��t�x^�HA)�4��{��@k�M���(��b����{E�z��kW�aZ�g������O}02p�Bk,�z����}�gQ@@�
稢aRޥ�ɐ��r�Ix�7Y��
��g���_���j�ʠܤ=c�K��[��M�!��8^:-_�gWC��̍>A�Ds�����V�qTh��z _��ʸ��[MsN��h�tX%��J�{�~���g�����d콧]�3�_v"lk��$�$*vRz�43M�j��NR���&�n���Ɣ�pX[E@-��ͦ�=��!��L!�$���(��R�	j��%���uY�!�*4�J&�LEՀ�Ǥ[k�ɟзc�S'h�����:�l��@0#Xk�δA��Kv��|榱eOVg(�F���������5׋�r�:E�Z��t��?��~��z���Q�yF��h
�}���5�a����5�B��M��m�����Ԉ�r�U��q&����
	1y*늾�
 �\F�K���l!$�:��^&���s��𘨳���_�(ȸO�sB�#���=�+I��%�۷y��z�R$��ύ[$H���!��o���f�!���f�i���Sz����� �a�2W��:;Z�ݮ���cnXy�-����7"���}�7�i͸��71Nr�Po��f`
~ATۇdj���r����)��1Q�g��ꉌ2��qh��
v��5����S�r6�\芀�H���/�D���[�*�"$��ۤR��.��e��ڦF0u�Չ���J�qgf��0H3Ԩ���I�.ʁ��;�T:(��g���-}��u�������°�����5h AQ���G�(×�R.��i��˲����m�Wx�����s�82���^�
� �d�~��O�D�JV�.Q���;�*6��&	sK6�q:������>[7 /�����<K\ԩ��4��K{v�sw���P��٠D�% ������<�0�v�l�͸��X/m�`l�*l����%����~����1��QޕtF��̍G��'�O�4��t�*�x �J��!RK����+���������ߦ�Rʨ�����=L>��%X
����t��r�G���
Z*�U?^%65��x,�Ek�����)��`���H3�@:���l��8�h�g�ϻJ��Q6`�i*���t���E�?��o�+�iF�Bj�wN�L�$x��g���
Շ��4L�B>8JhE�)&y����QZ���e�S��/uYG:`�M�S���MX
j��N��i�<���p��1���af4,��E9{ۼ+XL��?�\R�0�������Z}��w������.�z`a� �2$/��hϿ�m&4�?"�6��6@���j&�R��(	���*���!�f�R����!��M/�Ľs���A�	M��*�r|�=2���j�����?�0�V��gg!��;~ԗ�d�D�n���b�lܽ����?C;*xo���ӆ���XHOܴ ��~��������eJ�j��N#>g��`R��Bg4"��6��1�����u��#-I�dw�Oyز�5���IC� �k�U����!���e!��������>w�$�{�'T�Fѧw�-JB�Ǉ��� �%ϱ��A�$�p�;pֽ�lB�v�}g��,�qB�KE���QXŐ�G�!ƅNyH3Ά�US�! ��1��9�񳁳q.#u���r��ʿV٭��`�~���J]=tjI��Y�̭b���W�]M^��֩�<��z���͑������?I�`	S�6{�}N|䘵z͜�UGKxI��9��=��OL4A�R�9�E�k��}�#bh7*� ��Υ�������~��)�9I�Ӣ6Bd�G�l�[B�����=~N�W��~0�����b���!�J@� l4����r���ܠh��L�[��Ks�����BG�/:d���;��X���fϻt<���@a@�y��Eعj��S��#�l�w�y��N2luǦ�3~I�W<���o��e�~����ro�Cd3ڈ�)��L�����c"����I��x����3~��N�k�t�UI,p
�x�Ε�y��}N����_ypRs~t��[�?�_�]��)�8�k�K����g	,w����T��V�jZ�����H��d"y���S��C��[jMJ� 65Q�{.�q���m�,_7��`vx[�c%�Z��v"4��$��=U�To�b�P�6��zQ��p����.Q��j�l'ۤ���A�K�����������v�?�̷ӿnV�s2�\�[I�J�f#��p�.W��B����st��$L��L휜BZ�A������\�}��y)]��j+ޢ�J;�h�l7�o�/-�۴' 1��!�$���$7F�V7�R�/��!�㿃v��%�E�'=x��gL��=���*) 5޲M��X�XaGJ�ݮ[Ƃk�����h�O}�Lf�!���㺃J��
'�(�ѻb���}T�����B�+o�!�+U�Ŷnԝc�����t�6L���̓e��d���W;[	*}05�P��h/Ð��}�2v��Ĵ[��A�Ǘ��|a��._�0���%8Rp�>P��+$����l_!��l�/ɱnkf�m�7u�0O�o�r)�R�f۳�Q䍮F��jT�D�[��1��T�N��o&����O��įʤ�~Ȝ����NuC!	��D��d��d���O��~��;��+�i8�O�T�58�B<�ƾI������� :�R/�õ���%'=.S5�<XA~p���w|��6�3c�{�XĐ:c�H�r���'�O[�8��JZ?R1CЁ'��0��;.{=}�������=���D��Z\"y��~O�p�GZ���½��M��KQ�%.Iz�|��@HF�60]3�TU�:�dg�Kx�`�b���>#1m��R���Ci�=�x���w��4�H�G��a��r�C[�*��o��S�j�ՌM1YY�N��B��ҖW9��'�8b����~����scOC�.A.U)�9�0%eU��#�H�00 t�b᱿xs1��X���E�įg�'%_�V_HTJ$�@ ���n�`1�F��k�����:���`����=�L�I�FSo��y�� '~_O4`�x�������y7���1��\/lP�:��0R�3ޢ�>0ѩ��>��Ч�'�b�&d��?�Q-R;�lb���y��)D-]s�"�ls����~����BC15,���Í�� C0���Eqz�o�Kq��&OIp}�5"��*\1��u�@���{��Ë��0�,�Wj�J�������YR<���-�	7:@;���(�ĪQJ�gK�B��U=��mh�ft�rNY+��XZ5dWj�~��H6�ի�������������
�Ù����wb���(�N O�~�"�ñ��9LڟX�.h �yqvZz�v�N2.�Z��]�I��y��fn�SQ�Q°�m�	�YQD����V��1�[�I�O�.*�q�}��x�զ�ZK�3�8���`�a���V'��$�r�{��ru2ݘe	}h�J���{5[,�ܚ,���wgJ{#�g�q=Ĵ }�Z����J<Bj�ޏ۝��Y�WmO_)}�5���=��}�a��)���\���'��ѻ
W���Ŷ`�@^V"R�d}V~�KYJpާT�������K�����J[P&�*�mS�<BL7� �K��2�ݪ�NѤ�ߗ)"/zC��\ ���u!�.��#�K�O?�������5(<U�NZ(��c�%�6V�L�3[6��`λ��*M,W0&~���%�C�O������^�W�|�=V���bv|~���z�e��N�1�p�*�i�� B�w[����MI��Rtw��ԁ�j	U�>���������nP���	�*���܋sS֪o�.��z��e�f�o�}�Z7��I42v���'��gm{���f3q
�5C"���E���d�!U�Ͱ]Z���Y�-���ݽ�f(S���˞���D�m���e�����H*hb�y�Μ�ƪ|�Y�>Ű������F �ʀ5�I`C���h�?�w�+��Y�-��=�sS�n|�Ge����zZ �]'�D�FDf��Z�����f��wd��XdlzjS�u~����Ǖ|ف#�G��L�<�Y;���d�^EVA u J[<~
����������BoIa�}+
�	o1RO�Y�J�u0#^mh�\�Sn�|ɓ�X�ƍHVR��r}��'��\k+l��j0�!�gD�`�H,���)��g�	(,AT�S����K�a��+%�yY�.�E~O\���uaKl[Y� �1����\��D���O���:2#l��jw�[��˥�d����jU9���1�>
�_�@�+�y�`��VO	1zu{AE�%�1 ��z4B�a�����i�5R9��J��Z`j-v8|δ ���m��F�}��:�Z�!iҮ��1�;�\�
�?�w��[<�u9b󤿪T�yP�DA>�*3	�c��\�W�^M����h (��9�Dnq �\�x��)ƔA�0���C&�f��<�����=���^����}�M�;�b	T�d��3�Ùu��R��ǎ�~p��+�����=�(�^��-��n��8k�X��W$�="V&��.x�X��iU�}�݁}�-���ط�eO���,�S5�d����aF�3��&&���֘ZO��<�\S\��lJ�J���Y�z�IC��o]���ڎ��y':���p0~6�D� +�k�H��]��]`�7oG�t�GP%k<	��[����خ���P�e��r� ����*�����	X�r��6* �Ƅ<����CNiP&oi�����M��Q�g��#eC4�j�ք�����N�~�h6>��͙N���ХK��8�(1��P�L�_)��M-!��sj>{t~�"�g���;1��GC&���R��zV�I�IG`������:�R��<q�6�����0� ��`閌��q�'4����*6��[������`uuD��'Uz*�W���RZ�� z�T�M:)�/�'2��U���E?=.��˃�a��cH��R�-W ��e|̕V��c׍�큢����^�
�X�":�ʼ�Jg��,x��,�O �����i2t^�����J]2O~�s_����
AK��������j�]	����):��g��@TkӁ�W��l�AK�|̷�z�N��,���U�	�W�q�]9�~���*���
!�Վ�Qχҥ�g���2k)�۵�|jg��,	�[]�yaL����sL�)�9~�KGJ~x,ݶ@�@��n�j�b��_Z�#��$�٘f�qv�-����I�ȁ�\]��4���ȱ�bCP+��v.�m����s�Q�7��I���pS&0�}�!�,��l�sM"4��':0���1��:��OC�v"\�d��F�9�|�vI`���XJ{�ȭ�	��-��TC��T���`W׻�(�����}Ū�sC�r�o����ጻ��s����o6��"�5A�v�/7��ڎ�JE���e�PD��E������FK΂�kט�
�UG���$��R�c� \,>3��ѰJ�%��_�?�/�8#��9�j���h�}�n{%�R�`�܉⣀�F!�����+���i[�����B��\@?#�0����[D̈ߐ�]�����8��`��{�Pv���Q���-9kFMb:0;Ov�[8��'Ҍ�'�ԗC>ҫ�e`���%`+�:C"���[Qr� o7����0�{~���)�v��׵�hMP����e�څV��_��gy����*�&��K2��f�w�	�F�U]��x��
9�ל�G��^ז>� G����kX��&Ee[*��A�8v��#��'�s �����>vD��O8�c��s�&u�a�џ�m�����JDx#+i{R����*�O)�P�o��#��6��rI;�4,�H��f�\9�ڷ�Q��Ҋ�8j�9=F�ED"ۮ������\�a�%�41T�������9�w������~��u�J/���fY`��%��@⎎�1���4&���G[�F�<��S�$�K���ya`$�@�2�6�ydw3e	�=1���ׂ�|Eˡaǲ]�0���Ȧ��]���k�����1XK��}���s�_��&l��=Ƭ	ͬ�⧽��Y�72"J
q�K��Ѯ2�X��;�L0y�KnZ��B�vvDf��+I2��4W�@ɾt����T��)6�	���R����8���QYw>�7���Pu��)���3�-�"�W3Io�нY�|�W�4c~�t���avȌ��D 1�����*3��G����F\p'=������9���z@���I����<k�7�Ae��'<�>,`S���y��I$Zg� ����p+o�8DQC�'W��L��7d4�����5nzGo��rL=7뫛{�{_�E���4W�?�~���al5��I��Q��K���Ep-�j,˒�Q����n���?�ľ������O��w/l���ɹ��K���x:=��po�X"۰�AB� _{����������\J�?�E�o��kry�vEz=%0"��5�P�, �=fF��

�"p���	�vm90�=G	��MU2|�ͧ�zse��#��N��z�1�NM ��kch��ɰ�ޒ��'�v�7K��Sl��e� ���9H{Q�8�M!�mR�m��{�fmj��D&:��8�a�t�5n��h����g_���#�m$��	���=���4�$فɑ���=Y~=k�_/	L¨���v�\�4���Edxx�m����ۃ�(�x*.�t6o�y�T���c�
S|��Jr�p�������U�1)��@�N���]�� ���+X�"xp�Q����_��@�+N����A�>c���V�A��ß�'�&���$eŉ���!L�|Ᏹ�e'0GW�����g�p��`�K?W<3�	����D�p��{8y(0^��mb2r&X`�W<�k�_o:���C��/?�}�4�a���tU�,p�%I�OO���*ڌ��o�j�	1C���Y��3�����zamp�37�}&��A�Ĩ�H�	�#nXg`2슔�����z}�e�i`x,�:>7&cL)��1d���0�;.�P��@V�4��������;�9L$�`��bz!k����(�aeɍ���xi0�1K\A����1r5wn5#NA��/w�|����v��[�1^�+��C�]��/��R�לj�a�)A	�����Y��W����7	�8�J4���C�H����#_��|_��/��e����O�kP4���"�Zǔ�%� ����3��Mh�
�l&0[�C����,����߱�7X��~������+�(�F���IWb�%�����C��at�lt�>�OS)�(J��u�QK�%�G��hL3`A�qN5�BRV��?�Z�>�sqy.f�=��1���7'Cr���}�2��w����BRMh��]a��ɢ�L�Z6L�^l �mO����� ����Y�Wm�H�f>�p��꤇��y������Tkꏟ�!o\�Џa4(Gv��u|n� "n��M��*����{Z������ZV���%�ı��k������DmyY�RN(���Ā��+X����5Z\���]���C= ��{��Y��R#}뤠��<<1�F/�U� zm�����?G��ĳ���1�&�-0�݌[ó�s=�ԼW:�&�� ����Z�[������R�d
� }�V �C�	Y������Ņ��Ų;�npR�"����D�zF� a�Y8T��̠+	�;D�׬o��q�X�qUN�7�OJ2y��9�����sH��p�v�����U���8��;�����������6�J-�=�^��h\<n^"]��8`��oL�p��fm�XM��W�|�:���1;mJ[�h�	Fg��+WK�8���� 5�~-6���:���%��8V&=����^>�k#�ڟ����GΡ _�����Y�d^�QH�W@����ܫg�91;%����up��Z���^�c &1y՝Q�1��`%�sO*�E����HE��A�Bg�Iw<d6`D�-Z�}�]�
K�~��;їq�1&��7�nW+�N%
��طj4w[n.(�1a�a�:Ȯ��%�	l~	��d$��R}G�8���KO��Xi��]J8���Lg&��w*F�YY�<�<���R�*j(xV��kZ�.E�������M[T��#j��>���
4�"��4���,��xh�׎��X�P����j�.ބ\�L�r������R3`��p9��yƭ2r������	���|�[�իhy��焾dz̕`�|�nW��������|���-�#���F:y�z����"�@���a��،����A5I�Ld�:2u*]v�K�f��U��0����cίS&V������k�9B��8N�k.0� w�M~<@�Q�N��\P4L=���x���}ф*,>b���;p�3�r��J�:߭�<zܡ���ƴ��(@Gָz������(�y����Jp��wu�a�_o}��+�dP�j��Qm����\�z����d������ ��x�2j���F�M����J��\ ��pʿJmߴT�Ǻ�M����GQI�����[��>-�v�� 2qx�qB�F��s�}Y-f���*�5I4ҧ�!k�Ϻƍ���G�4롉������*�����O�;/�%��
R�IO!
�M�$����ָ>�P쥜���+f�	>����[�7NV���Q#e�?dIa��.������&@����
F�%���\��t,cԢY׳
c�B�h��Rݔ�$�> �@@�[6��q��fnAY2��(YCn'~�Q:�޾P������rr�ϟkW?ZcdwA:*��X��#/h��Xs6�X��Z�B��6�r���oA�D�giԢ�n�؟�2�g�r�S�bD����Vuu1yA�&��������d\�n�t�sH�ؼ�S�ϰ�������	+��e��Ug�d}Wخ������,�?l��S엸�*D��EOD�J�oV}��p�n��@?�E����\Q+��"���ᠾ7V��-�aH���j�3�l�o����zv���L��h����u��M$A����~��X�����\����ŝt�0 ]�ݖHH;Ͼn�b�e}TQћӅi'E��$��ȑU��[�7d_:�}K�,iޤ���!�JG�.���@��{���bF5����1B�y�KD���}��E�b=t��;� ��O��Ҡ�ˊ�֙�9?x��X�̩	
3���@M��T���D!�s�;7������U�l-�c�ˁ9��8���p�N�o(�&"p�Cv�����B�/" #1Q/�jC�� �+�Y+�����߂����ܞ��ʮ���s����Q��4��)��H����0")`.D����
⣘m!*z#򺌬��h�cCL�ׄm�6S�!g�U�� I=Vݤ����)��/���]v�u�E+tW���<�2=�1���VnQQa����8"�J�7�ɗ*Us�]��K�1^�T��.�s�X��@�
��T��i,^ێg��{����[Mᤞ�P��:�� �D�l�K$TbS��&��*���珰�����=�fHDI�:��Ǿ�*x&j���Ԝ�?G�r¿���r�i��\��̒02ԓ'�0�h�{�gm����U��~�m�Ζ���������}~8��(J��G�}���ZEa�M�U0C��3�D%o�a�>8���n:�&܇Z$� �ݟ��i�i��)<�W�;2�s���i=�P��T��&�ܲW�ͷ�����_�r^5ʃr�:�D��Ia�0 |���,�:(�i�pR�`�Q��;D�Qr����UA�~�Z����O�?��}��;�ݼ��s����u�b:���S7��+��赫�F<��,)]�o�e2�� �u�F�"u�b}�Ǣ��;מ����{����͖Xn�.�C��$@�M��絲��%�C�G4Y]�<�eY�7`��AN���?~WkUh�;�a�6��`v��g�e*PAC�+�2����*l�<�۵-�i�PT5�Z5K(V]l�F��E�0��˖2�F�`�	�rM�Av1��(W��QU����H/%����x�WҕaY���}�-���,a4�%*B
h��2�1�ߞѸ<ݦ}�+D]M�;���Uʨ�ifN2�)��[����;*r�Y屈�)���T�F�B�Qw�M6ڒ���0Lu24X��{<�%QYH�1�#�WR�A���UCmV�X]�ޠ�<8s�{s�޺?92�V�ay�����8=��1�W�����!�������fa��1�p�$"�)\��~����Q͏�f�+B���lÉ�5)w���/+5�.G�������:h��n>'�*l�l�f�^�|�a�5�]��l)}T��P����6a
iZ����5X<�^^|�~e�,�4�h�/��:A��p�EU��7�Ҹ�.F'����F� ��5c��߉q\k�h��Q� ���\Ʒ���Ԫ}�������"�.q�*nb����uRjH7N�����{1}TK���v!d�*1ˀG�2�ؙ��%<u>ʽ���H��ϘΥ�e�3k�״��t�H]m���C���Pw'���
���������&<��3�\z5�D�Z�4�-�m��X��m�i9h$���B�r!����=�dz�!T�aJ^Nz�~[�CjBbq��H*����VҖQ���F�]k�_�ʍ��iT���l�V9p��š�{�#smj0r�#7�p;�A}:ZW��0m6��θ6��ږ)�;��hR�5�l
Uʙ�뾮ȓW��r�J#��W��d�-�V0{>�0��r��[��X�-r:�R(����Fn5�� ���Uq�Y'ƧK��Ԅl��%0�m�>RoܲXj�s��B" Jg&���r�`F��	x�x�xѵH��:׺��X7�0:��^��)�?Wɹ��E��a�6 �=�)e��C��+���$7A�|o��R����2����m!@��8FzpSTA��"q-�7>�ǣc���8��%���8`����|�Ē�N�|M�a�!!�y{[�G���[��A�ڃ��p
�j9�5|�
)�(?�v���8w�gh/C��&��KO
�D"�a��<���<�}E9K�xb��
w�_(��	8�=��*hΩJ�s���!_�fȘ����#K�0BP�'<Xl�1o��܏�%�h�~��n,j;n�I~8�oV���*��#�T��ެQG+�C���쓓I!@e,�y)6k�`���'�v�i��Įz��I�o�V��H�P[�J�Pƙ�P���ғ��/���#���TWIV[��p?��2u�?W�Y�,Ms�
�KJu��Fo�?�������g>���]dϲ�[P�$�|i�&�m1V�G�(e�gh�j��	Y�П�Ј�r!���Q�}i�@ܠ$�1���Vs��:�)�/N'O�T�J�����Kɖ�**(܃�{��6E;1'T]�Q��.p|i��HAH���k����Ϙ��4 6_;C�xz
xZB-��?7�ң�ʔ�s����,>%�B���}+4��A�|(����)a��\r�����?����A�%HurP���\�f�}�Z�E:6H�Ð���
�*��%+
9b��W[�'zg4�d.�R�㚺1��`�e��])+[5���	2�H�E  2-�h�	�p��~���=`���i��-��4�D�>~@aosK���\��i~�E��f��]���#�`d̩v�����&n�~mj�'$j*�V�d��[KzP<�|����?�2޺�e�tio�障�0��������'��S�~ݼx�*Z��GnԜu^���sw}��򶞿��:�t�1�$���y�Fs$�w�t�e��3S�*��L�������Ex�
�v7O�?���.���Ur���H��)#5u��my$x#"N-y̗�(�~�:4����"7�U�#"�C�R�s�F��ec�� �;h��b�@jp��:ȵo�ȝ8z���
����yлp7����s��a;c,�=1��;.��mW��Ńfz	V
�!�i��JwSa�ؼ�y�ꃍߴ����^�e/�Ab��g�x,�Q#/���B:��j�3���F"?��ο<�T���,����`wq��,�֕������
��C���)��g��w1����񪹜�:�B�.`v���0���L�ªO>b��2,�����i�
0y���)PCH��[��@����&NE�<�o���H��Ν�uG�1)�+	̓�"����
͓���~e#���'5��ݏd+����f�@���ł03�zC�gD��`�1�oYfo����C��O���Pl�/Y�'��v��� hvT�y!d���)E�7)�������Z���ڑIM�.Kw�).pŽMs�q$���6��a�`(&����$�O���O��K~�e
-���D=I#U���C4�Q�g�5��?I�6䢧�P}�I�����w��?m�7����ƫ"e�t��Z��I7� *��͢&�P��H�k�3��"��!���b<#�*u�y�À���̘tjzEm���Q���R�k�L�$C8�c�'�ؕ;w����v�|E��z�rX��2�͵�ih#�Hs�	x��h0�T����c��r�T1E���59Ve�0�zvq�8O- ��6u�8��(�ZgښA+y�ZY&	4�6߷�=W�Jf��10:�ؘ��V��|]/^��tr�ش�q�=-}��Sr��3��}b�Dϊ"���ܭ�w�&۰�)�0pe%
�;��#8p�t�Vй���A5�iuO��^N�
��Y���m�^��[���H�.$��YZ���o����=��7�U��u>��b`�!m�2���ö����_�9sZ�F�u��^\O,��37��s�L=`��PbJg���I�*:h$���u"><7��!�# ���l��qJlvчd����Q���u��$���f�ε0�jvɋJ��!�F�?m(�9����ş�	��<��(L�vRA"���rCDh�i����^�1�Z�8�H�aL4]��fV�N���j ��pO)yHRA���]"tr_v�As�EMK7p�L�KJ1`]���?�qbb>;�
1H�+�A9u"��Ɲ���or	e�h$L<����|���tI��n���K�O�čs#sc�i#RBWB��H�?u��Y(4��˨:�bpvgk]@7;��@�<�����|Ķ��k�)��/�Wdݶ�@�S�z�T�l�4����ڠJ���;]��Q��o�1���(�ߩ��[�k�C#e�r�uPԨ�X�\�X	��cz;� �Y�c	�wC�u��tg.=BN5����/�2f)�n�f�.��NzT�T��t&aGjWZb�!�m�7���^�Y�R:�:�R��� B��ݐ8�h=4��^� 7��ҵ��]ղ���7��	�
�+���V ������ n\���o�E&�5|��gK�E�E���B���1hza-2���CX�2g?	"۴"RJ����ٯ�G�R�8K�;PjӠ]sSN"n%r��,�(!��J��X�]sS��(�5�]� I
{*]��(�}�=:=��A&XC��B�$g˳ ��1
h8�t�+80z�����H�=ŧ����}`��� ])�H���/���%T	����(e?[f��*�7�ұL g��$��>^0�0��-1�$C�_������G�jc�ʶ�H���&��,8��c�nr����LS����?��㈲�
���v�u�#���D܌�i�8���*���%�N��8C�8�s���@x�\Q��+J5�~�]c�d��gR�ҒR�#�Z�����m������E���^ � ŵ����E���Y�eTf�Z�e��}/�Y5�q'��n�o�x i=�x1?����L��e�$�q��^p�Yv��'=��j�v��[�G��>�8e��=�᧶���.�=�zQ��$��1�Z,"�"�;@�η�I���*4q��?�6�j�l�T�Qj-]����V�K,=��o0������^U�A(T7� ���Hg1�-%���"2����}z�_C����^	����ZL��%������LϢ�l����	Bf9��Qη��D_��1�1դ���L��ӵ��U��i.�E�-;\��Ll��O�]��e��ry��_��0M��X����P���
\�[� �J@��e	@�E�>��GL�\u�O�O�{wn+$Lۘ�|W|PSd��[2�=���&8��UB�����m�ڋ|R�D���#I
J'!�Y�}�a��U�ߍ�� �H8���	���(��o'�?z�DV��ӺQ�J繡��GM���6Z��8��������Ђ��r��K��x�򁛂~�S9U-�Ν6=�K 1/C�JN�Ò�tH�>d�(mH,�6�f�w�G '��.B,��{�'�����r�0��1���!T�g�)!h&����� �~��|�����k�j`�QW�)��c֠!E�H�%�8W�I���=�{�2B�!#i��!%���X!#Z�Ǩ�[0 Ɯ#�jⁱ�@АQ�����`�o�|0DMg,�ƴġ5�k�>�cE��)у��e�\�k�W��{a9�8lM9��DR�,=,��ha�w�Mg�y!]{�����Xw�ڔ����,ׅ�jPn������	ٵ���۷�������0�:����Wy�}x��3��ޖ-I���d�p?�ٱ._\D�Ct����R���i�������P"4��}�D�fT�y�]��)*r��Q&�Eg'Zo���_\���y�\��P��Hџ��DZ ʫF�S�{\Z�|Oe����%�4��k�b��J�h��%)n:8k�J�;ό��0�Aw~�f󧯔@{*;��NzV,��{�F/A�)$I�d/b�g�\È#i5H��}�ð�C �v�D��ƨ��=፟�Ƈ�\���_6�wp
ًz�(���Q3ȋ)���������)%&���)i�fF��ϻ���c�
M!�{sbI��9��9�P�X�^. �[_A�grWg���$�;(��a�����N�P���[�8��H����:����us�݊���`�8��,k�1	[���N�l���6!�⩯$:2��-��Y!:��&�&����6��B#������u�F5yW��T�H 
��K���i�g����Rfg��x��[�ˏ�lw�깆�e8�w���7q�|.����6�ҏ��x�7�(�*�	fP��]J�cdk;�͵��GP�oA�Ubd��:���8��!�����W�/mt!�F�{�eX-���Ҡ|��֙�l	�D"1��h8ɪ�����tR�E�;����w#m�-a���;�z�DF���a���ݧۥA�*��s����ٰ0�Q�U���B$$���.��o(�b�EH|�����$��_ n����<�8Je�e��ז�������i?
��^���/n��53���;�YO/5wg� Pr�w�����?*Է�҃�B͔�!���qo�x�Dab�[׈���T?!ui���^ڈ�7��M�n�a�ѕk��� ��Bi�m)�N�?V7h_6֗1�,���C'ls��.�)5=d؊J����r��L�+���Dǀw��P$o�\W��?�/n�@l��U;˥�~�mhZ̸rb��b�����ʺ �%I'��k�Z�de�`A�v�q}�����Vy�$#����zg&�C�i=��f�̒�aL�9ī��.��)D.Ba�GAeЍ�B�E8�6ei�PFB�s����Ւ��f���&�п����I�[���W�^��!2�-ҟ��5x*w�#�Q�i�'�2"%K[7���7&���򺧓H��������sv����1�W���@�9�
�7�ܐz$�Sai�_ϰ�CL�A[������˧(�3�U���4�t�'
�2�$S�=�Q��$�cSiw��iX����z�U�{b���si�8���U���ۭ���_�(��'k�?# �JN�l�N����|:�x����(vVTL���nR(Db=Ҵ��lW�y���Ÿe����������s�e"`��_j�O��tZ#�y{�f0dc7A��{Z�}�ߪ1�a6Y�;-Ɨ^��3X�eHٌG�{'���DV��e[���,���f �N�*�������Yծ9	�z-�� )��[2}���F��o�Wl�1�� c�$����W�<����Z��C���H@���#5�UU�GV��t��j��x'�`�Ӊ��8���� ����n$���Qչ���y���4wF]��~�"e^p\�����V�R���	��Q���0�:���@sH~@�� 
�Յ��w��'iY�V}�ƫ�S{w����sՃ�?:��Fˎc�Wt�m�Xqd�����z�43P�D*%_[�f�t�1�����]ǎ��0+�'���+	PJ˫d�,p}�U���B �ab���*���t.�4$�ѽ +<�HDV�7�f*m��}�;x��&�� $�KK������s��!N���.��Ѱ���(0��n���U�1r�^Yd���xD@@@�����l��◟B4��0�Yn�T�uy�	��KZ�o-*�T�龑G&F�����F:�q	ta��9�����P���A�&�a@2����(M��7�Ɲ?s��¾HF9�V���d��?�:;������B4 � ��:�E}��0�U1�ĨwI+OV, b� ~�b3��2���O�*D�p��AnbԦ�C<�|35G�4���d>3���j�/ �Y�V~�lvEb �=E��Y%!w;5AP`�w+�� �vjZ���/���6P���Q��/�����1�]s���A;�W�)Q��B!�n��o�w@�:7���kl�n]w!���QEb:"{��I��y��θ_� �	�G��Fob�Gr���UoBj���At��'7��ߨ�m�L�{�ZW?��݊���-QN�qt������+�_��h����&���];�M����N�����T6e[��A��<��8�f���\M���NV"��B�߂0/�({|g�x�
�$�h����2:�t���.�� ��ED�]�C�51C���'`-�%�-:��bND�'A�g%h,��|�r��}��Ƥ�~��^l��\<�F z4^���!�q������
��^mb6E�i�xb�Կ�|DU�Q�Ա��0���U�IM�$�v��B�`�CS4�Wv�9ۇ��y��''�s>�Z���`ÇJXug��O0p�B�p�9gUU頿1t���Nwz�ͺ�J�󥝅1�8]	Z�9.����j��^Y����zG�:ܳJ�,�sƐ%��
Y���x�LK����EOhd�����9��.�vzc�/�;��N[�WF��7(J�<{�oY��Ѧ����^�]d��K\�����-ݶ�1۠r�!�%9�(���l�ݭ-�Tuu�]Ά�#���\CW�~z}����f�����5� ޷2֜���o��o(6�N�����6�FǶ�|?H��o�'�@oȿ9V'�7{3vW "�����y�-�x��*�)*�\�l��(U� ơ���cɊ/�$ l~�V(�����4O�*��ꜟJ�"F�a8ݼ#d��@U�uD��#.�6�b� ��x\-x�u*݉��P��H��Pk��v��IX� 3%���+lC����kN�Q��2	�����x����� c_��`e�Y���S�!p��w���u�slrI1���{2'�v�P9`B�7�O���|���|
X��*S q�8�����QwK�_�z��q}aCKj;m�y)R<�6�g���G�;dT������k9�PC*y��]�Ԑ�/��)�BĥT���wA`3$fA�:#��
ٺjvi+��T�N�D�F'�|7��[����NI�8��Mn��J�{�6~�lo���U:��U��$\�
{a�3����Q�Ά�) O:�i,9#!��e���eX2�kzk|`���M�)����I�o_�D������G�r�y�L^@�OL-; �a�$���-�ۥ/����2�#���{�|��2�+���QN��	=bvثx��]m4��-�Y_2J��*;�3MwՍ���u�Nd��u��_�:��wB��gӊךϒ�BW~�?�g�f+�)�̛8J1<�=���ke�Ro��)�`��א/������w:&A}�vSA^����t}c{��,ټ�R ȤQ�Q��f��h3�1^M2ۍMrǬڹ���B�����"p:C��ͤ�V�����vq+>A�ʸ������8'�ߎ}��L�:�o��-��<(_��8/�[�[�kЇ�����N�����\{�[��e�R�)>���`��5�@Ϛ�@�z/Bo,	T�%w%���l+���a�jd{�̽���(��!�b��I�A���L�4s�]��7PN%�3�����ţ��|!d�ɯ���0�����;��P��랧F�ԵW��ڤN%?��z�����''�#&���[�����9�x5��<�~A����X�R`(~W7F`UTx�����O킄Pz�U�I���cv��$V;�:rr�yy�\%�-��H*X8":��mg;TW���1��G�Nr�n$>	�E��HAB�Tv�A��Ξ�j?�Z柯޺t	�l��U7�p�]Eғ��2v��KD�f���u9_N�F���q�6�c�a���B�)�9���&Y|�[��Ĺ��B�N#�6U�W�	j���C��q"v��c�h���r���-VIX���!8�D �+֩�Ɉθ���wN�^�:��;@�^t��ӗ�^�GsBq�p>���Y<���#Q��~�n/�,�zz�ը�����Ⓚu���˔>�M_��8y�Z�3�e�N2�Sd��� cS��n?�Hˉ�����>��9兗�LoN��昱ے�4���#[�? � �r,M���B�H ,��ub��.��!1������TqY�Y����n��0�f�,������oC��	L!�vʧ��2��#ϿG�rY�>&�M��1J�����H�x��I�tr�Nc��B�G(��m��I�G��,>�mD6��������P���C;�@�y���L��3����Gl��$v,��"5������۴?Q�H�&���`�x6�+~�%�l���?]v�ћ�EB͡l���;��I�V��m��?!���'J���1|"�˞�ԭ�$6
��/�B�<,��`8k���e���u�.t7�w�,���@���<��b�l��4O�P�H�oP��qpQݫ���Ɵ�U��|�blU�h�u�(:~1����{���;��Z�9k��/����g��+)���u�K �
���GZ�����*�Ǝ�|&�!��T��I�5�5N��55��&{�/���6�e����s�Q��,;�C��D�mcE�8$��z��tJ���C�8�����R��>=�0��g��=)%Ap�HҮ.{���^�h��I�i�,("1��?gͻ $���B۸%l�G<���'�sy`��M�.6�w�,;��ؒ}�*>�$��09pv
�U�.�����L�b�C�S��@�70����8'���e�/-�68kG=����.�g:9�����U$���OŇ�f{������1O����]B��f���� ��o=�\��io�t�5�'�e�}���H0qs�0~�� �2NTdFo�v�ֳ����C��n��X�� ���8�:]Y�ٷ��Ѧ.������}�h��_᛾��D��z7��>�{�|���Z�A��L���wUA�5�d�[�J��:q��Z�Pxj^��.>M��J��5��ma(E`ŠHq,1��Nf��n�D�e�ľ4�lf����I�lS(8 ��R�S�qۦ�Hο�ij�:�[��<�x�/�Dx1	����+�OG��ƥ�>{K��!	�8���oV���H���Q2*��o��&��7�7y�ǭ!�_k�)}_bZJ�4��K��&wJT��7�]6�G,8n�Hj����X�#�7I�ň��r|.k]lZ��;o�Lf��
 a��k��$rNP���po*E�J�X_��Q��z��+��y��u:H+u"��1��p.L�9F�{��-	�>tDz��x[|Y��4�m�qhXrO�9ჲ���G��32�s��L
��S����d@D�1h�b� ��4ܻ:�\a��H�ȑ��к�f 
7�;�k�*�K��.D��RX#+���u(x���wpdþ�V�h��;��o+j$rwy�8$�&� �����[��?�T��M8���5��6;W%���CIN��Rċ�0�ZY�]za_��g/A�����7�H���r�?�&g�W0��SYҊ�GۉO��`�/�NU�jh.���K�o&�v�ä��Y^�<�����rs.���`�\��@2j����@,�1�7!h!yב�%�Dj(-����8�)��+!��5�� ة��xe�g�"�V����QZ��.`�՘��8�?Hۧ��.j����qJ��A�>�
�p�9�����(Yc��x��d�St��^nv� +�+p��#Z�FwsWV��A4� ������c�(c�j
B�Qa���1��j@�awqO��뎄�1�s��^'���5�Ws�M-�Ϫ�PSСX�'��Q��ܪg ��W�[�S&FA��n�����ݓ��gCk��;Hd4!��� hs�� C:�E��_�J�`<`�o]P�}㎕a���a	c�0��t�H���������:e���8qyu�YŰp�>�K&�_�!�:-⚉�.������:�ydم�%*vK�r�<B=�����"+/5��>�h����C��B(�,�1�v��7y�B��K�ǀ�]��&�,kA�Nl�SYq0*;�Y���_��$�Y���#y�d��Z
�5u���LeX��g�zrQ�2�sa8�0�A�|w}	��=k#�)�e1'� G���]�hyw��������SQd���[�}b��foI���G\�]��H�ԫˣ��(��=��V�=�!�nw�{�ˇ���x@������Mųu}ӭV5@���}N�r�"��L�?c(�;|Y`����F���p�("��z�O,R�������?ʮ�IӇSRN�5Q�I?O���<�%�s�]S=6��\(�D��y��
��I~�K2���㴗i<)Y��R)��yby�8���G�qi
��A��c^�(����Q�3��G7-�IB"��� Ŧ$�o@Q(V�W�0N	k��Yq�1yc���.�*��L���)��ъ�mI;µ���͝�V�4�R��r�ޚ��z�
z+�Zc��
%dI�sx������,ŏ��4�A��5�8I��Y{z1
0��3�'���Ⱥ(ڭ3U�Z'Q��`�=0�GS�|��O,���g�1\�t�lS��\m�L��v�ܓ{�i�Ļ�C�1<&P��綣�*2I�h��묡�Q�?����Rr(��L0�1���D����WM>V�5���Z���A���H�ޛ�:#e9X ��&Ֆ�c���V���@���̸�� �{�%'X�?�,a�M%��[v�m��u�����|��"��������y8O�7�7��֝�_=�]ZZ�*�!���r���CR��;@�̓z!o&Q�j�t��#��E�(`�g��R�c"i�R N9S/3��O<�(zy퐐^{>݄_f	��JD)��J�Y���(���J���D���Aw=Z�َ�$׺��:��g:�i=��@�v�j�%N5���̴��fu�G�C��aJ���Y�C�Sk��F��L�yy�B�h%C��N6�vaK�K����F<2]�!��s��PaH�9�Wv�AK�[7����n!��	,'��o�a��|����2���$:?ܠ����G.����)�ʟ�V������u:���05hHmU��_����[f8��<=\ר܇��y�«4������Tx�Z\:J7�l ZO%攮���;��d[���O���gљ�A�;��- �����X�
`y��GK'�1��!3�&�ax'\�
5"����h���Jx��9����R�c���[(�֐�.eK��l䷈3�0������;�j9#a��v*��؉y�~��ߣ<w���C��i#��ug�����ж�9F��i����h�@|Y����������E�s��$�$]P��j�F���.^�2i��g���X����0�7C[�\������rܡڽB��y* ���TK�?���JmiC�.._�|\��3;�w��[�����Y
��~����ƭ,�״���3Aʊ;���u���;��s��J�S!۵G�}��r��`�b0�fҮ��}�*�:o˕=c2��*x���V��S������\/��5�r��Jn._m���[hbkR5_�[���	J��j���UZ*ي,8��M��j�&��ɫJd������E���A'p+�N�w'Ðx*'��"�Z�����ir+�����M8t�?��6	�"2�RQ����z��w}�;��b�%[��rzC�,b��w���I%�PjQ��	��A�0Q�TV�s�Ó`-3)�ԯ�3��Lw�����T�)C�f����Ds2oF�d?���%!��_�hP�~D��  �>՜8j[�:[e�粚<TK?����-�H9�� |d����ɩ�e̻���i������q���e��M*����z�v���)����\gL
`�)A�o�zg�]o1�<RЏd"X�Q�p�09��S���O�<����Vn��$���r��J�����%аq�����&=�R&�C�F��Wj��6G��|�T�O��h_`�	^��x��=�tS��B�4ą�i�s��K8ns:�M|�=@rʆN۽Nf��j���v!g�#��8-�A.�}Ϝ�phL��w.O�v`�&lT�\�U{sa�J>>j�9�,��1�^���9%��J r!��IYw�Yb5��6�.kF��؏j�i��!"K�i�@ީqE�y�΅��
���U�����0��U���x�������8�#�R�����R����υc�5�ҝ��]��Y�	��^�J�*O�y��_�X�}���ɶe6�D�5sT�^:b������W���Pd��ʪ��3�F9G���~�B2��G�,�O���a��ـ�{�g�n�8��\�4�ǥj3��Gn0��w�[�{�K&G�C/!��us��P<\ss�>�:�Fp��x��Ǳ%�L�=lª�x.�'��Ƞ�?� %/�U��}Kٗ{F+�8 pI�E���
@'Ȭ�Z��6c��i�d������;��S��V�y��w�b����g�g��*vԫ�)ag�*�WwI@Y��bŜ�	n:=S'�G��ɋ[��#�3��R��.o���o<c������JwĤ�#��zV�ڼH"[�^��/�:r/hz�~�,��j*�����ْ���
���ɋ�HENz:Ɋ�C0���	I]��`��s�_�;�!7y��ze:�z��лe���}��\�_�<��� ��e��9�Ń�T�Oꢉ����� `m�}�C�<�u>Q�O#E*g=aN������u8UV�.���x՘9}pW�s��@�܉Fه�dޜ�Ա W��G�e]�ޢ)ʨ��)�S�n�؛OÕ9-�5�0�I@s������Y������!ߟ^�,�m�Z~/�C��S�ۜ"�n*:*�2�E��p�r�L�P��p!�'�	M'��Pvb	s���g�9s���˴�Y4�L�%,�Y���2�4֠�awh��R���Q.[#�$R(�Y\�õ�sy�(ݗ���6��j�*���<�T�Us
�(�w�����P��(���7��� ��'��c�
��:v���`��m��m�|W�5�.ԚH"8d��[WA�S�N�O��Xش�&������9����}N�.}��{�K΢Rr������h#p+�]tov��I͋�KEnS�����\y�0w��y�8~���͓���;$^������B'����j.�9k��α��� �K������o�:��a��]����gyn�@�r�i���-�\�[�uJk�k�P��<7������Y��y��e�UQ��1B�&�B�q}���#�c���Ȥ=s�
ԭŰ"�����G�iV*��������oy0�I˴�����s���OcQx_��2��Ӭ�$�+с�c�u�;aO��g�2����H����߫=��.���|���".Op6Nm�DtG���qa'�o�?*wb�F�t�n*<*�DbJF	��{q��pVl=�v�(�V)`V(e�+�bs)��a��d�/M �X��7��L������S��G[&�� ̋0[v��m���-�W���Ք�. �H3D֔q"�m���di�|D?�5}�j�a�_A�W��p�|�(0�M����xЯ[�=п�m�- Z�z�YM\���S��8R�Y,���׹*����}�q�:�>���E��6��Z���{K�I��W?M����x"k�CO�y�!�)�9��}*#��>+;�9h����4m�[.
�e��$�M�5�HC���ܶS[��Pvu��-�"Yn�������ϐz�H"���H��F}MG[�en3��$���j���}�C��f���8AF����z9�����?S����p����GHo鷤�Da%7�L<?h�Vv���1W�N���A���G,�C� �����Y���6.	5-wL5}.�����X8�e��B8-�w��P�Q��>����և4�<U᯾o����������� �1e�ȇ����)?M�E�k`�uI>qt���\�'��u����]��Le9�S����p�G�8ܝ|^�Jg/�<���%�׳}�A�n��rv���wu�hҼ��kD\�����Ǻ�2�Aŧt1��-C�:n� ?+���쭛�@�X���7�S��{��+��l�P1��4��޲;��
�K�G�Z�ݒ��	�-yk�G"#�&�P���a��\��*��+�%{A��s��<�
 0n�[?3�e�u56f���c�@x� �Q	Y�)Q%'x�l�V�OB�I�HdB��/Bw�%砛��V]&���!�z���!<�%՛���f�er;1D�:��it��M����x��h��x����X+�����[�=�J�ucOu!�oP)b�L�J-�~�|�2����*�Ve�|@��c�vͷ�e��aJ1A�5��B�Yܼ~Qn������cw�2�$�DXfH�rp
a>;�4���-[�%��h��+<2��>�Zm����K9Zy�)��5,<z-"�!��xjAJK�պ:}�ds�~]CV��!A`1���+ؿ�"�5z2����̃�f+����S�#�l3e���Z���~�x�.����Xی���`�И,RumT���=�5V����7&^�^��z#�)�o~���P�����.�vM�Q$�?���zfO�0ԅ�g�� ��*����|�i{�n #��w�[��U�Ѯ�[��2�������f��kN��1"#H;��&_IN��Y�����V����V���v��'m���l 3�G���H���3D��%AZ�!+�������� Zgm��]����J�{��������E����ϑ��^�Îȇ�^�._<۹�̞h��G�|���7E<7O��|ɄǖX�뇐����#��J�s觧��E�10���/骮�tK����?e�ܬ���� ��9W�=v�>y�vC9.�1��+�0���,\ħ����Q�P�-�>�o��+`�IMn	7��R	ׁ,�=��?�m)��A��=�4���
�z("36i�çț��z���$b��M��(�����-CER3+��.��Cc�5��P&���48����z��,ʷ�2⷏�Yc5i�A*�I�����߷N�o��l�0�[U}�UFEv�JY��q���`V����cT^���R�.>r�� %�C���t͎ �����"E���:��%�S����	\�"<r���[R|%��(� ����D�֑��٦#_��o��}Y�u���$�04�9�J.z(f�xK�J�u�s�Z�[�kѲV����5����jw�O��gw���ϝ�WB��h�b���w}~*y�����g��)���!ZMA��%]�u>���jNj�]�Ӣ'�j�o�6L����w�,tݒS�~���bOІ� ��~<X�̣�z�A�T�a�\���]��h,�h�T������6�diش�U^�~�K\���1+�m����n�\�Tm���f5�m�ь�Z�X��X��+�����qm��SS�ZCG�8}o49��D��˳�E-�Js2N3S��G�u��,�mlN`}Ps��k����Y���Ó�J y������L�z9O�����T�$+!��G�5*	��W�Wa%���	�G�J��̭6o�j?�b���7�C�/��f�4m��w)ؘ*��Q1�z�l��CU�!�!�0���Vw�"Km�.�M{�\S*]h �詙��X`��t���Q����%�N�S�|�w�$<�1M�+�X�F��Z�X����0ǣQ�j��_�.lA�q�M��k��Γ 4k|���4�s�jо�p�+�@��%��މ��M|*~�`�X�n"�l��<�IT�ٷ>^����l[��~��6�RM���s��E�p�IJK{"�]��e;��h��*�j|��X]�� _������KD���S�p^�d�4��i���Wfí�xVT4��d��Z�Z6�$��R7��==S�l��˸}?��q2T��g8H2�����չ�Jf1:�iu��D��`��&�-�/bo���J� r�^� JJA��D�Z�X����O/�˙U�����Q�Q�3�[�H�D��΀w5�)�����8�` 7�����VEFP����z9�z��^���ql�px1Z�d�sJ)Ɖ��w���Bt5b��	�FPI7b�����h{��#���z~H6����aQ�x׸�K�z��SHg�\���ˌQ���8���y�"K#�1���Ζ�!qZ
�)�G����>��J�-�fX0�M�9��Y"F�	�i���Ǽ�覽FO�R @�����i*�%���9^+z�I{�D�#$�v��q�uw�)K��tq�.��D��@UR����#l-�k����f�@c�Px|�]��=�,��)�m���[�V9s��9kuX��{���F�vs���
4�JMxh���c��c!9W�e%P�'-�p?���Pކ!�5���;^�b��e	+d6�D.��Ȗ��zl�kj1+N3tm��l�r��N������h��T)�2����l�H�$�As@�`�e ��.��Nͷ���ns����EpuA�O�94����Q3�Xi�qUӗ�$y��/u$�&�R�m���-�k�n$E���\�N��w��3ލ\�-y7\�����~<��\ag0C$A- C�Y�oY�2�]}�A�|W�����O����XM�+���f�#�#��*����j��4T��-��X�D2��p�A���z��A5K�E�e膹���_�k���� �pr"U� qQ��f�$#_��?�^Z�'���Z�>�#j�p'EW>�)��|��|O���e#Zf(��S3��RB�w���SAG���b��m��S��-��D�&U����
��z��5�zJ<u6��+�����p�^�Ši��`�y�q��S�:���{4�y�������0cO8��E>ԡ!j��qͬO�!Վ.B+�� w9Gg,)�r@���o����OQh���+wh���qT�8ʬb]�:]0�泼��;=~�a#�B��0�s��!5H��K�R�M�e�^B����+��@��+����fF�|����~�QW���Ũ`D4!��~Na���W��q�m�U�ͅr�6����;Y�~�~c��wO�m�/��]�3O�nvd�UՖG�н�b������a�|I.��"��w���|s��l+ⵂ7jB�:����x��u�P�|����^yLt�*�[�TOkQ[��p��80ռ�d6r�|G��.�ډ3}zaC��¦S/I�r��/^p�*��2��-��Ҿ��0h7�O����u7+ wdՑ��)��A;���.�
tY�(�T�B�rW�:V�rh�~��C�|���<�~Vg?�_:�уQ�۳ �?#�Qv�e�A�+��˘Z.���
{����\�y��fpE�5*������F˲X�ZZO����$ ��$��m��'��L:��4P[� �D����^I_�{Ek��[���Qp,Q�4��-~�Z޷yT�e'��V�8����1���� L��5�|Q �M[0����\��@�9��c�����K�v�CO�	��,�����r3�d�
)�����n�Xuz���ߚ2[�&�ˍM�� ^Bhe��&J�!�u'3�~�a<�P"��Q+� �1���d |�����Y,<ID��ha=�}�Jl+�H�!�6j�6U�Ju�!űM��h琚�r(༆m0�U�C	ް�z����b[�A����Y{t�ږ�|�e�N�j�(�i�vo��?�/F�1�@���C(�����	���������u���UB��o!D��4y�?<���(�ԿŐ�̏]�1�J9�4������=��/�DpM ׷.��ɀA9kO`łnc����z	��6`��}��fs8Q�C0i`���ī�^E6��u
/Dӥ�6J�G#U���_���0i�d \�Tu�d!�v��L��'��c�p�(��V�V7R��/c̉1cT����g��.	r�Mn���,�hD"����.��s�cw�}m�6-I.�iH�]��b�U��j<�0߶����'����$�E_�T��u�@w7���v\҈�Aպ2R�3h���+<��<q�̃�8�<�+T�K�V�����lkۈ����<�p�p>D\i�X��[���e��`d ��B�r� ���ёr�I}Oğ�h�ф&��@HOq�+�sp��7��MӶ7u�9��܃�Q����e�@��#����C�!��v!������Y���u��x~�US�9��桄[q���o��%/�U��A��\S�G5 �ςL��7�`��?$��|��H���G�`���+��{;�($��2���\����YϗpQF��1��=J�{��"�'��A<�=��2������g�Q�k�h�C���֘0��j��������o"L�ú{s��CK��8�;�;E�z
U�P�����~_A[_;6؇^iJ�&}Iz������c��Yg�`xy�p&����R̘cUɸ(՛����x���{$ߕ&��C��.!�y.��O�ѓ��rk$$[2�C�n���^|�{�v�v~�		�(Q��R�k����rr����DYo��#U(A���F9���~�EsD�f�cH��g�V>F�6�Q��1�9b�r�a�b9�V�#ӆ�?�9P`@�K�!'��At
e}��:�C�$�_�_�	���[a���< B���*j8��4%&��*�	X#�;UT��ѳ*�U)�+Rg�9e����\�;����RGf�����\����vzV����z,�O�s5��i�^6��m���M�4��j�I-d,��xXW���m1��x=y+������&H�+�LLL�l�ZV;�YE.��JL���O����!�@/\�5�@}u��A@��N��/��q}�d�b-x�z�l����kp����e?=�@��s�dy]�9c��0�>�%�$�B.
�r�6�x�f��a�a�j��� 2s<$2=fn�oÑ��Qx��t�Q^%3�ϲz7р����u�/��,f��a�{��,��	�)��Pv����R�ٺ�%q-�<v�l�S3���#�v�;���?��7B,�AMjΏ���!N��eՅ���C��a��+��R��)�^,�����G�o2w¿3u��0MO�4Z�:)=���Z��"C3WJߕ&rxmo���.�!h�}�m�%�L,�N)rZx"�s ���+�g�^V���K�a�bI���9n� a�[9����+i��b�5�z�Q>Ae7��{b�%~�G֚����|e�)�pΣ9��iЊd��;�.Z��`��Ja[�]L�������2��`6�9xhvcr���o��#��5;����1���K�Ū#�A�M+Ú�P��љے� }fN�A��s��\�9���B�p����N���8���u��ͼ� �&���&jJ�o�#b�2��'|k�c���l����ڳg�9.���h#K���'�8�g��M�hM�
آ���9�sb�T�_,I#3��'h��C9��W;4�yDE7#"� ���Xp���uƷ���d�[�����f�mϐa��g(2H�?�X���F<��k�x1+��*���d���6����Q�D?��v���u�(�[vc�Ai�����r��<�V*ŷ�a��|��{��\"(� �����]6*����18�J)"��Ə୛��s$�h�$@P�Z\R� �[3����ąQ�
k�p{9�����������+�j� ��뀱����e�o(6���*Ԁ*i�ʚz�J��Ǝ���nt��0�f���ۼ�:a��C���A����-Z@m\W�8du7��;G�#�L�| T�2'n�X�5-#���r�#1P��S����R߄fO�4��nV�w
�~�ͅ�M�!��)�+:s�i��0��<3�T	%���Ï �u�t�j�Q(+.Zr�l�-�%�a��a.h��~�Z�gr���O��}�Ħ�����Bބ7�
D5i����C;uc{*0U���e���s�4Rֻ�{��=�[�9W�YFG�c��֌��咡�BPD&�Qp�ن�Y �.t(s�Z��͡g2&���͓�e�s�����Q��|����UQF�SNN�{�:L�6U[�����x�A3�B��t�X��}�C_7�����SC��oA��jk&@����Z�S[�.?Q"�@��B�n&ӫ�\xTK<g�~������Mf�8���e���2͢��@�Bc��^�C�Ÿ?XF�ql<� )�]@��<�#�[�au��Waď�e�x�����>�_���}�̦���]��� ��V�{'��t�G�)�ݧ\��w��	�G]M�b������3$c�d.[$�y���ߍ0i���5"�;��CZ��Z��+ѧ-Ն�:ڛ	�a��tPo�����)��vA�T���Ү������g�w[NL��K�Xs�3��Ct��g,{2�S)L�4hsr��Ł�����"�&��f,lmj�G��Lx{���ZCPx�#��Ove��O��qH}�L+�c2�7�0���^���җcS����$�V}ix�2��Ү@"h&2;� �e����`�$f�1��z���[g����"�8=�X�.��_tg�T�9� ��>�A��h��!�6�m��zށg��G M���-r 
Qw� .ӂ4sP���1st�H2�܎�Jsm�]a&��%3����M#w�U�M��ڛ��w1��Q;���X�=�G]]c%�}܉x�>T�� K��o�%�.>�>��ic�.�\юs`�T
q�Y�
��7��i�	M�'u�@Q��G�{�j�+xp���w�co�LX�ّQb�k��`,�*O����${N��o{wA�M������ x-��r-�.	epv�b5!�$e�^�c��0C�����>���B�v�#�02zܴU��B��X�Y�i������Y��'rH>t�Bc
�]��$'�b�+F���A)M2��e
DԹ�v@��i�X'.�ߑ*��j�U���N$�ݎ����m��QĬ��)�Y��<{Q�TW\�*�.��P�b^�2�q�����D	�[H�8��Hx1�bŭ�J5mY�{Nw�;��u4 8����YN�m2��=�$���j$��w����IP|z)��QCz������tO�Ձ�T�{<�����3�h�
[���9�ʇ�Wױj��$Se��
'Y)!����F�*��*�/%���դ�;��C-���ݴ8k)B�&�!h�kri����Ag8/k��8�JrJQ������0�R+���>�8�.�5�s���3��^J��US����A��?�����G�Q�v���wRn(�$uY���N{>_&��$�[�,��IJ��d�mvdA�~��r�D�6}[�cxJ�Z��9b��������w�Q���0`��lʡ���������QÃ߉�ރ�I}���1HR�v�=H�Q���Y#s�,Nѹ̷��~.�Y�F������0�)Ϫ�ؠRy����=��
���Q���m�V��*3%fa~䱱f�~�l���+�u�6��r^� �ǽ�صb����E��tm0�e��@�Ӆr���J�?�8��܇hc�ڏ�7��[�� G_.i��{���G{����nj)���Ύe�+<e�j��8,��=�<��A�'��S�f�јMz��+��2-��@B�&�[Vm���k|���--M	6r4�7��W�F��[�F��֗y�1U5�-5�h�S��ZxRQ�"!��N1��a?8���'SM)����'.� �_���m�l��
�%�(�h|���Ϲ�"2���:��{� ����GG ��G���I�XQwlԪ	0���O5��VWkk�^d�:;e.=����]hLX�&�����'!��ZZ��b�ی���p�fsFUkK� ������5B�J���溴�8���+������.w�W�=�;߿K�����Il{�a>��0�`�z���Y��(��"���Z�^Gt�
��asѤ�Ф�$R\��T�s�jf2+΢��\��pm���׹��*�j3���^�ԟ$H�����L=�眅g+Gi��}�aN޲�1�bih��қM�@�(.�g��E�?�py\:�Ӄ��k]0 �����Kq������OA���j�6x�f`�P�0Hd�)�q��A�� ���{���P�Ut�z��8�5�Ʈ?l�s����U�6��0b�p�t�L>������5(,�ĕ��0d����cD!���p����$�:��D���J�d0ӊ�<�͈Z�"|�I�-�,q�4�=�Y�\dx9�/! 8��^�2���XC�o��ߦ^�!���W�;s������c�]O?����~� �"��x*�c���@<5= h���ǠP�u����&k�������c64��Y�򜁇�<y���7Fi��~&v�C��4��<��mO0^���'_���DR`�����z�L����rt��������ޢ&�Kco���y�yj�L�Ǻ�MHڍ}��Io˱ɔe�F�-P&��~�7f��w���z���a�c�:���:�#�*Љ?��)eY�+�W�qF]Y�,>�yK ¹սd��V���i���;�� �U7��lJt����ͅC� @p��)�8�u҂Εt�Sª:�2��y�߮�87i:H�i� ���Կ�(���y�L�j{�p���vϫ��:� J�e��Mo�Z�tZ�3 �ӱFO����}�� �?y�dȃ��]�>M�S2E�܍���0O�`&���\���OD�?�QE)Y��c�y�Zc�;t=�U�?�j֧��Tg\o���ڴ8��Q�Xyf]0����>�TM��{z2��|��eE~ާt���j~���]ڹX�̉a�^fV�N�qe�'�@�a��Vԏ������A7�M�gھ3�}f(͆0$�|��Jg`�E9���j^գb���WʘP�
qN�&}U�7�>��Х�����V��6���b+�[�`�k?yP�E$�Ĳ�R֊)~���7l�F�����*w1%��-�E�Z}���%��P&Ƅ���/���sA�7�/Q"3)�d�q���d�VO��~�ƴ:��~b\��	{sdfy$�O�"�U1��QC�:��'X1�p�!���b����6Z1�V���qW�����G�� ����]O�����9ƽ��Y��ae��H@��ۊ�D �6�H
�Ι��C��`5u��-�yk�R
z�萑�ыG_a}G��D-5�W#����~���ۣ9�
��I�<,����ٛ4*B3��(:��*��g59��:2̐>�{����.�GK��2O�3@�3,�Y��)d�mUG��UN*�	�*g�q��߰|�ˡ���{Ep��T5�9����a�|��?@��֮�#���w�m1�v�@��b�m�D�3[�~
�P�~�P���P�������w�r����Ϡ0d�����*7I��D�LPn-yG&�����E��/� ��Ep��Ӹnj��S�n�N�1ŎՖ�=��|��h����[S�D��n���u�h������J+&%����p�C���L�R�1,�.�襂/�u/pi�!�L�w�SQa�VCpr��Z�ԇ{V���������h���-|/?"l���?� S�A�x�1���&[h{a�|�kj'>k{A�&�D�s'V���L�T}�
��
��7�T5*��&�U�@R<\�is#�>9����\���oQ�� ��A�����)"���+wM�LH�8)�*ݓ��}HAf��ӝm���wE�D�0��f�0Y:I�.�5��|�0a׎��1��lBc�o�ϙ���A�2���@�^�pe��U),�9�QƮ8 ^�j+$���[��##Q��Sy�P|�j�Њ�lyg�I��V���� ���c�!�cW����J�f�a2
<����%����:�����S�Q�S�����y��h����͛�Z�����+X:8����KҪ��٦�|x_� 	r�sZ�W��6���Vr���,h�N@�V�=� �;͗�� qM�N^N�4ZČ/��H�di#c���e��U,"��~~g�_�X��nV�4���V7�@$,˂u����m�� �d����v۞�h"w��'�;�
γ��<�"!�$2�ca2,�w�Wޔ'���:]=d�Z���n�z�ע��U\E�U檟=c�d�����[�A�I-��;�(})����H�,܅�@�)��=�d$�!+�w����"Ͱ�+4�=�k�l���_� �"�xY���9�Tp��F�*D�]�_"�\B�Ǫf�Q��]0�Z���y#Qzb�&�A�~"I�T��b[���Ke�pN���L��%j~w*t�)2�co@R�c3�s<B�)Z�]qg��y��M7w]�
� �:
<o�!:���t�+�j���J52>����1��[OP�b�D&�̗�:\��\y�E���؄�e$����Qn"�v�wy�l�^Q������%X��2��&T^��Q)rŢ��l1�m=�.�7@�@��� �<��������>�U�6�׎!���;�;����aDii�4�&��*<44@EÓ����qAڂ��c�y��-��t;��?���Y$q6���˗��H����%�X ��˷W]�m��n#�����$�i�KO�l��֑j�W:��f������j�rd� ��1�bݗ)��X/΍U	o��4HI����n��I���ݦ���*�P��N�HE)��1'cٶ����b�9���ߘ��D|�i4�8N���GM���AFe�;@2����Gf��S6Ԕ�}<�s%���G����~]�� a�,Ed��8�W��s���<�p5��#m!�N�q&��V����R��'�(y�2��|��y�e��	{y�����t��J��*���DAe2�R��k�@��`v���M��"vM�!��@��5&׽�p��^*$�B�0Z�K�ж�3�̘����� �	�������fN���+X�JO*di�<Ϸ�J�&�%\�R�t �7F����� �*�.��d�bc?���wx5 �Yz�1l$7%Z	i�m�b_�/�p���*�5���{�a�h)_�⪓���С'u$�ϫ�0�����T���B��_����f�;�3�/n/�, �6YR-��w���ۅ�5k[�񜀳Q��#9�<>V��B1����OD�r�5��ℤ�������6�ȦS�kSN���+Sp~}��
0,�<��"���&OT��=Ԏ��8�U�.���ؐ�*�r �<U���v#k_�o�Ŭ�|�Vt�g�+�8�`�$ ʠ�f�Գ a����7�h� TߡM��vm��ď�����6��W�����v���,8a��
t�>1xq��r1�q _�@N9�}j�����w<�0d��#��!-�ի���V$�cA�^2��|*����x� ����)�h3���o�~���9_YV���6�S�*@x���,�.Se6ξ�c�;`;~��ϩ"z�vط��ǆ�ESF�v+���h�/Mp��!^�l�D;>SX~}�T�<hA˻��ծ-�n�T��B舟^�� ��܎<�'�x�xb����"aQi&��qC�w����Z��d"�����^�v�Y�\�e�`dB[��9hs@2���g���M!�n[�~�M԰��_6��xl���������s��.��\��7�\,��͕r��%(��oj�2]����LW^Zۥ[ =�K�\�l��>f� /���u���?��Ti����6"8T��g?�ߕ��:��q�����k� ����@�0
]�V!B�S&���xh���$�	/!=l�̸: N�!GV�ywu�0��mO��4F���Jˬ���p��s(��U7K�&�C��X�;k1���i��uv����Э�+:���-��(�{j�:���7K}��nbt`��hO���*J\TL5���jf��/tb�������ε��)>.��$�>#��������I���z��=Z��%_"H���'��Ǻȥtv���M���G��<�L9�P�R�sB��h_%% ;��F�#�P����"���є��	ՎDo��c�{3*����H񀦾�G�o ��)e����.����m��
������vf��S��M��	�����6k��|D�+��"2�@FJn��ίi��Ց��4PF��,A3+��	%��U��/_�n���/�h�;^�<Ŋ"^hY�W�a�9�|Q�2�U'��z�9��)WjZ��D�lմzs�	F/a�Ҡ�w��}�����Ľ���>���p�����P<Я�
{E�sU�|��D(��@��`�S9�Kנܪ�E�7�5E�i�����������W����+c��&�,ͿnUKu��Sΰ=�4Թ�� lf����B_`T������y[^�w���\���
ё���_�č��[Jc1���%�I�؁����G��"82gfHJ���g���i �B�o��ǔ���_������̐�lQ�:��[��+�D{�k�v7f{٬&Dx5�aҞ�@��:�)�"x6iH��!��o��>cc1fO���9K��> I��e�3�9�Nk����r����u<e ��<�!M����|q��:0�x�E{ȏ�i�N��׍(�V�3u$�<_2)G�K��J��Ϊ�Ɉ2S�]<^�z��kT&y}Ƹp)�}J�^^zH��^���"�����<�7θW:
�i��-;/DM��8e��FMTĂt3~���]{�v+��Ԗ?�V��4\AbL3桽\���V���;�Ɠ��&��Ё?�M�c���do��bВ6m����%�Qr�u/��IDD��)��M��� �[�e���ޤr����$��^^EH��n��O��;0���?#Q8���B������c��z��3C��B�BD5k
M����!��$|�b�5O��	�_Ss��4�T�D���F�2��
֦�ڴ��k���Ͳ|��;$�=*���yhZ{��Tg�?I��#U9J�v��°ff�� ���2�`�������:/�]��^D4Mg�qe"�5P��`~�܂�<���a�r�Z�����"�h��-�$ĵK!�xfA�eT�M+F������|���9u�U���x��Ҽ���y��.��56��Ԣ�8�8����ZN�iH�}#�8':syb�o�̨]Q�AVǺ|�o�6��v�� #�*���Hx�e2q��7�E'X��\KhuKF���A>\�5"EQ��rGQaTT���K�hVP=>+�B��5*���s���GXZ}\Q�ˢS��y�O���Ii>.�3�uӣw��9��q��7b����:[������/���mI��W��t��e�m�q��v>uEo����&�)ٯI�Y���l�d��5И�LPZi�+�M� �Z2������l�E$�OdL�l�l5���I��0ieκƷKOC����2��Y~���h�7�u&ѡ(�,cw��&�����Q� ���^`C���^�>�_sL������w�H�������A��*�	)�T��w�����)���G�wOĄS'��/`�h5��q����s&��`($�;�'��*h�@�1���b������;���$Q�S!SE�{� �P���� a�c�F��IW/��x������5)��O��a����=$= ��Π���|�V�Bt~J��Sj� d/!-e�²�I�D�������2%�6�;	��é�����k�`�$�n9v,K�������7Aqs���2$֝��R�2�_��u�uZ��g�Ռ���������I��+.��1 ��[�	­9�]K@�j�+�Ϡ@���5�t�7<��]jcwz�Q�lx�tV�w�5�VuJ�G!C�-J4y5���FfwǪl��L���q	M�\���R���3���H�:�_����^���or�W��C\�����&,��`l�i7�yq;x�
��Y��-�u���{Z�m������勉bX��;|��ȶA��}߄���5-)��s��w�x
f�\�&l Al�l7۟̚���.omw��{|�y��u�'_$>֌�iM�΀{��۸Jj�r�R>�3���>ϸ9=
!��]vO`1A\�cs����@���,Q��5�g����j�`м-O�x�IL�1���^â�!��q/�Aײ�K�Ւ�1������_���U�O🯽����u|���t�:ai��M�\o��E~ĵ��N@�fA��i�Q�aJ雛5��@��^���TAl�\���"�`:/�ǮK���j��?c�������z��Ig��'���1���>$�{�'ب�&��ěln�L���#�#/�	8�i��Gva���@* s.�q¶Fel{�h_�w�ߣT��,n�p�"�f�*��7)�5*o��|��
�w�!�:�H >ǘƝ�87*Yl�O��*!b�?_��-������S�d�ҚB�f�\;_ M�t҆%t���:\��m4�[.l�#���!L̕>�M>���
t1���������p2ʌ�%����10wϮ'��}u6��Hm�%������+�=X�<g2��7��n��^@FUrTӂ����#�P���\&WΖ��w�����G�����#����R�;<
���1l|u:U���}(ʸa�Ed�>|�y�C�`C�Vyh��!^d�p�ϝb=ݽ�)��:��̑�Oㇿz�Jh��{W��-���7�
.�+�����~.Q�]MP�	Z�'�	�I�.51l�|��<e�zq�G�U��[n���Zg K��Wr~c�'_[~xx�����>=ͧy���^$��!�UxM.|�X/ŊEFw����\bN���k˒��]�M���[�I�������s�7�VZ�RK����c�;����XL�K%�蝖�pu�83:�:�]�;��z��?D�4�q/齡�8���O�7��[۶�
0��v�_������HXeB�AK���C� �{x�b7U���@W�s�V��X{���>А��U��������r�.�@V�k���B-�/�qڔ����&��cM7>��=F�]�l�.������Lַ�M�l�æ��pV�<@��ds*rg+j���q �0񱴑p:�����O��T
��䌢�z�塚
7'^��E3?�KU�# ��R��5
0 ꍿ+w`���\�4��泾*�M�^�B
�$&A����K�_{���V+;�
��
�<�?�5;��}M?!�1� _�&p!�>�Ջ�e��L�<��uR,�ҳw����5�m��ؼ�yQ�Ҡ##�j�;}�]���
�4��^�<X`ú���@�z�a�=3�6}��|��#���s��.�!��68�Z�7n�.P?=��M�^�}z�O&��Owl�46KUt֕�W�}�;�R"Bs�~4�J�s���ʌC��<G�=1,ڴj`|�^Yq��)u`������R��P��l��"JR����J��D���U9~,U:�3�q�#����n�e��ﻌ��u�(���.���G�De5KL
nPP�J}���~��Fqx��"��:c�v"n�L�qDb�l�M�^��X��uD�C�~!��T��QA�SCc\��r�Y~���ћ]3c�hMЌ�d�'^?��X����8bb���|J.�Ɋfcb[�.O���Ľ�b� ��E{e�P���'�����+d�lܦ��=B��t�B�\.��V���%����Iѻd��;n8�Ek>>X�=T�E�<[hu�t�Wz���s���\1ӕ2#�l��^�Q#-iv	�������du���J�K^a�{�5K{A���0��J��i��Vg�;ل���0��eY`=�(�'j���o��u���)we���(�ubl�
�-�/$��]���� ɨD,�%_<�dx��s�T�'�++���^����ƞZ��\�Ħg�����q�;��j؝�})��ʃc��`�9��Z��0E�O>Ăvq߿���jK�7
�u�n��>���3�9.kn����<�Ͳ�Y��E�|��i��8��Sݠ���� �|��G	ɕ���P膑/B���?�W�F$�zz[j��mx\��/3��`�GG.�!(Ld��I.>�|�A�H����F�KDP2v.�j�0Z����ۘ�0&t�ٗ��h3"3	��ّm�Z-�<Jv;|*4��r���|u�U.Ns*M&X�DŌp_C��
�����R�jĕ
K�H{�ǻ�2q��h��j'����3�O�*��S �	M�v٦a�3I�0���=�m�����[�dr�oEL��s��	�P�=!s�3��¬�7n�=29ŀL�z��0̵�m�?�����p���EO��`Q����(|m�}�/�ˎ��y:;i���8���
���FV`Ā�}Gn�8D�R<4pBǁ���$��G�����%��}�B�jB��]Z[����W{S�VX����=��^�"�@�V�A�%�!���t�h�5꙳���},|vS�'~���a���4���f0zc?>9�*�&���K\�);ӄ�v�c��A��E�Q[�o4}X��UgK#���z��[{چ�w����o��$����n�*|���Y�=�:E��H��V�������,���4���Sߴ9��l/=��9P���7�X6	�x�{��k@��mU�A�-��
��5�*�ݟ���{߬�jZ@��1e��tčǭ5h�U6���~�Μ@���#���ʷ�m���n�G�t����ԙ�V>-c����h*��׉ǋ��z�-�	��sj�@���Y� ���5Z
s�U��ϸ�m���9�:P� {WT"��2^X���'z�퐟�4|cK&8�՞�d��A8:Oe;��b�e����G���ҧ`�<�����i/����Ŝs�!�"��&�N��rի!ÆB����a,�Ino_(�9K��!'�ѿK�n�J�Lz�i�@M��Ŷ6d��?l9fl�e=Q}elT%��[�:�W����(��~I�����Ln2���j�|���-4�6h-E҄�������`�3��Eo"�^�A���U�tl��d��49�3�3:���s<�����T�m��nrH�UJ�@�F1��}���p� )ln�0w��0�W��;C@LaV��{R�'�����Y��s��fk�0n]�\i7��v���TZ+�R ���}��Lh��ўe��#bn�˚!��&�,����ǻ�\ ����̱M�S����t���:)֔�"�7	��}��e�Ӣ�	[����~�M�*12V0���B�Fl���	`��{�Mx�W1��5W��Y���`�!����W+�)A��Z*���}6�	_>�*5K��?����_m
oA�	�E�uegj�_@M� �#ZG*���τ�Z��l��y=da|�{sχ)4���5�*���Uߤ��>�k���9E��T��,�O�g�^����8����M>�WV{� ����q� ��x��eA�h5Z�m�l2�{�0>�ZLt��ۃwާ�e?�V�@�PwPRlN�C:N�ه�,�-#�;?�r@ἷɖ"�;���FD�W�g(5/ЩQd`ޅ�^���2��BA�I�ʞY�{b�ݖs��{���]*��*���E[21���z��ы��0p��*!HՋR�kx�讀T��W�nH�o�Bf�p�ę-��pm��zM}��� D<�n�G��|&p}�ը!c��"�Y��ch�'@��?�U�,�v�X��|��8!l^.������I�o��Q���I��Y�e���yu����!7��TV�UN/�f�숩!҃꟮�'�{?]V�A!�FU<.�x$M,�7#������8��I ������"�H��D�B�D�:��oH
���2�MK�rY�sͨFǲ���d�~Η�XgÛ�^T9X�D.*�w�bZf�:끴4x���d�=MuZ?l�NG��$���+��U�sSB�r�8E�D+�2�����/Bi��mX�5A`(H�8����a�������/a+��^q�c�����8�{"%��:p��,+�Q�n)T�������,�/��Iڤ8�7.7K�"p�j��^Jݰed�d�M�����K*�H0vjMQU�k���@���2�3آ�6OS���o��1�y�-k:�.WjEp��ߠAgA8ߦ�K��C��=4ɞ6�X(g,���>�$V��v>ir�˫���^c7���vl��U��I�E]��Z���s	�������G�ŉ��2�'D�Z�?;�����:�c���$V�8E�i1%
V-r����^\��E�5��@g^�2W<�� ����y��LZ��:w����
6i��_��QV��H�]!��`�4-ڽ,��mg�'}�0H�1g/ǧ%�N�Ko�U���p����ʹVQa��l^����lj�yi��m�x
�V7� ��	^�3���������5k�� QW�0R0��v����t�qRlk�wƏ���9~5�K�Y��Q����K�	�6Ͼ�b�OԓY�������N*t�O��1�+m��Wg�ƺ
�7�?�V��"��_q9&��׏�C��4Y	]=K��F��n1fe�'��	�����p�Mb����/x�y�ҪY�	�ǒ��'�Y����E�C3Q⣬\ٳO�)î�ងa��uV�0!;�r��.F�����/,,>�ڟ[�����_���@kp��iC|�D$}6�q1���7 �f�xL�(��n"�ᵸH?y�,�rV�özm�	ݴ��V�W˰�.�J�r�i�\�(W�m�d@��p!}���{^��M���b�,|w�c�H�r&�)^��+-$�^.���
��-y�~����g<Yy���.d����Rb�`�ф�
fx3F���k9�=hO݉���E9�A�q1ctoeS�M=�)���I�a����k�~K��e9�*p��X������k<D��;��w�"��]��
DB�x�*��^!8�<ra<0R�W6��f\��8C�V۰4:��Y$� p�+Th���|��Ӧ�KyW	b-���K�5��~`0>��zae虶L�k,�ꁔ��q<�858:"ڪhV�����+`
O}X��2�f�w���{���SB�)���x6�PT,�z=n͏!�����y�.C�t���D�ي@I�=�!/F�&�tA8�*e%�n����{��2�;�?!����T�d0{�+]�烍ج0Գ >�Ɖ�[��V��4���y�xl��{"�������q�O�x�x�y���u�ճ{b@}�ȫV����-�*ݚM���	�R��.?�������Z���Y�h��^2�g�Q��MpI4�ͨ�Ⱥw\�`��H@�"�h����!s����bV�W���B��)S3f�ʢVi���Rx�f㭇ӭ�h�'���fH%=�D�8�d4�sG�#Q��� XH��Ӌ�������ha�a����2��1%1�)�F�o�ـ�pے�q?���AA�_�����l�1�ݷ�N"�1� �L�*Њ��s��}/�wP�þ$g6�0ؙ�8mHY�G��n�@�12$�=���[��&yK����7\>^��s�b����x�ԫ�1�	���	a�����K�]_1�jῳ�6�<I�W�O��U�Xb'�ѹY�	`�����9�X��CY�{QM�+8.�����D{ O4�h@����AE�o�1|�*�����x��fHy�+��;�/s0V��Ë��I��UJ���6-���񝜘�7�|�(�ߗ���<�#��,wrۀ������zb	�$w��s#��0�G�Np�@��
���mߦ-�8�IK{{U�5�(��χ΅^��ђ?��4{��_iW��;	h��iX�i��:�Ȥ\���]��&��Î ����w:vz��]	�xEh��.���I��1�s�3����LL9W��1Y��̐�庀�� W.0@�P���?(�ؚ]1����2Q��^��H�k⥟&�9�/�9ϲ�.��~)�5*}hqE4n���5gՅ��o������FC���s���1mGH����ܥ}O����/�bF����t)�i;תƘ篗N<�R�.�]Ac���-'��dfhT9�65�
#�����Z�K��b�ֺ�3���*���M���F¹W�ت��j:��n�K!B�=p��l|�3��	<~��)�Վ��W�%�kT��q>n�A�Ln6�o7�����T`6zz8&�"z�8�� ��Pa���F�����jc���1�nܮ�|�����I����=o��\D�<��eC��^�ں��cIЖ(c��6h��N*(���X܄���s��V; ��đ��eN놔Q����#a�rADTǴMy� �dXܒZ7}� _2�TA�e��!�����]�*@c����:��a'�d[٩����|O,��M�z�H?�����0,�1<�2�H���H i�xn��>�	<��F�׈��9]�ي��:&�Q��?�u#K������q1����J����y��P$�OLa����uo���Nq�l�\���eu
��X�f��Kl|V��[�>��L?��*���g���-�F���a	U�hy}�5�g�����4]�}ҿ�U�+o��Nre�㎴�$�L$܅�e��ך^���3�%�*�L�]�v b���o��W�۩1JɈ���c��*�-��a޼UCh3D�c^4��r/()�F�N�k��C\�D��@��:Ɗ�`��N����6�su�+���պ���(�'�%�D������`ή�-���=َ��Hx&i�F]q9ga<]��2�	MG��l8���-�5X��� o>�&�8˹H	[UӔ�x蟍�W@����~�HC���5\���R�vJ���LO�(��<:�����\.z��X�lB��,�w��Mc�s*����NT�Zs�=���/3���,fo�S0_��GM��(?j}��i`(_�Q����pq ���ƜՑ@-)�J���4h�C��_5�؇�;�0��y-2��nסȒk\I��Ӓ� "�f�^�&K��L���N��όQf���j
���d�����S����Զew�>Q�������zv�:�(�XB˶�6I�L�����~D��:�&w��W����M�T�9��b-mx��y9��L&Uh�Vr,�a��K]��є�:��|qw0��΁L�]��˜ iE����'k�?�=0=�}?Wh���o);���]?`��bu�C<e�7F�S�&�4���'�� gB![�؊>
q�K�H>��0*���긳q���4�M���}a%���W�@z#g+����`bï 岉�ioQJ���4��!�	��q'~�+v�,,�A�p^�\�f�խ4i�S���Jx
�P���ݯ�����Io���O�3 EFDpd��#�Y/��ku�K.�D΄ʘ8> L&�#}l�C��1�6�Wn�&,\H���˭@���#%P�X����6V��01k!<"vqH��v�]���4��p�Mt�;�kx,�� gr����{��6ɻ��i5�[GNH���hb~(�#�J��?}��q�!�����}���1����>�I'GSTYKr��R���~]���� ���rg�]��³���D����}�c{�p����h0\�� 1u>}�I��i`<h��\D/�)�����8,�)e@C�k� ���)#\T��������8��F{�*���W)B'��+�	0�m:y�t��Z��ܙbPϴ*upу�=ǈ�%�Hy��٦8Y���K����&�*�Cq�9����W���}ǌ��c�֊��x(���8����/y�Y� �`��7����G�轣[^HjÞ>�ّ�� In-O��
Q��\�[�b����Է.������йɈ��Ԛk)?�7�����@?\@$*��E��_6��V#[(�J�'.D���2}���V�Aba���K0�ܱ�n�b�|�<�BJظRP�3ED�t�xq�2�j�3��ڠcG 5��́��%��v�hf^uh!��%��H���|��ЫL"�2�G{y:��3"����*��6b�G�jV�ky�rB��Ţ�Hbf�sZ�ؿ�r���y"��(���,��u�G f����$C��4�3�*ٹ�A{��B5���B�K9�"gGH
�]��*fr����Nɒ/)��*!���Qʯ��h�8**���*�1��~�7�Dh��i:4	��XyNi;����MQ +W+�G��)DХa��t�����ڈ~�V�f��Y�D����5�����&�ۏ�B2,�E]%��d�ؙ����嚟�M�1�������
?� ��*\N��M���'d�6��(�
F��Fb����?�Xn���eg\�����J�9ȴ�t�G}X����ew�h����J����j]����)К�����(1�Q?Ug�[m{`���n?	��y�t����H\�g?i�R�tb���T�4Kx,�H7+ּ��T39���ͷ>���H�{�����U&2��%	E�E����)bt�NΧ�7C�Z�xmO�F�-�|Ð�[�<���뇴{���++X%>���Н��ƞDϨ�:�<��"-S��X�#YA�K��HS�gYI0Z��FEg�[�Z�>�{�3�#�x@!��N���Oy�d��U��ж�3�9�x���1G�m���e-�U��oDw�"\�y�j���=?pQ�@�J���@*G�v���'��&o��F��4�]�xQ���w&��d	DY���r�>'�EҋL��<
Dæ��dwe�����n�oZ�h�Pg��7����̮+��5�޴�&e[:�~�gPF��d4��>(�Kk�A�ZU�-=a��9�+ߎ����R�z����t;^g���KEZ#ܨ��(j�2i�n��G�	;
u|6i�-sbo��OR���į��
����`�D�1�E�C���^p����4�c6!p8C���f�(�͍*�\w���n�(�U8�]��Ͻڝ�i���]ɀL`z���J�B&�����������3��σ~�_��e�ۚ� *F��_�b˶z�	S�3/�M��_��jx�T���d4��B$������,���su����k��ү��B~Q͏!��Z�8��6����x�')���M���M��r��m��'?��ڿ�X�Ջa�	�����i�=6���%����#�	���t@(�Us��穲����y[mJQE���977n�=Ҳ7�E���2Y��j?����l�w�2y�GĎ&Z�6=��4�yDc��i�K����>zӓ��P��]�� D�6��&��V��?�
�{�x�]/�%aͻu�&b��<]�Y�>쓠�~�#�xwd���'d6�$��l���;����.L�J��X,��5�-U%�v���������K�۴����4�I2)�y�Tur��J����A}_����"n�F�G�J�;��t�H�L�����O pӸ{��8�t3gf��8A���M��ܝ4�	m�K��|kճ~���ߨV>$I0B��:U�����e;ׯ|���i�=���?}]��� ��в9\�L�gȚP���|���b9�O*�0J��AY%�<��G����6�]�ġ�On���m�
���ǵI������*P��;���J�;l���ξ1��M���㢰*�J��K�'=P��`vB�/�c(�� .�%�<N 7[�,�^��`&M�.�J���̱�Y�RiӚ��ʪ�IW㾞��e�j=� �Cs>�Mt���§ْ��S���"���K����R����9�P����K�Θ!�y�Ҏ��ʻ.�水��z��r�!��`*��|H�2�+���zdz3(D�! ��ه
̨�!�u�]?�H)z�Eg�?O�ݞ�T�uj[�!Ct�Yr�c�pUś�
atR��4�`=�j���]��U�R�.�F��t?��~	�|[�[�a���V����3�[쪱o� }�2�9H�"��� �ޘ��n$RB�Ԫ��)����޴��J�!�?�6���ﷱ28g�ط���ux�g�F�9�W{Ig�#��B/��&�r������ǰc��!�}�C�S󵪨���ӏD��2��[[y��!�x5-��%EZ΍���u}k׏n3�y��_�v!���&��� �b������'��S�Dkղo�|&�mR�=��g��l���u�`�@#�&�(�P�F{�X$i����ӁX>o��/�o97W�Lу���˗�
QY�~�v�!A1�#F�H~��I�Е������pA[��p��O�Ke����xn������S���z.�lO��L�F�3<@?�f��S��#��L)p/&�z�ObE�1�]�p�>�ܟӏ��V�1��zw����������i6=�Wzr�f~��g�aK���$����zz��"PF�y�q�c(潼`�iMp�R�q@��)˜��Z%�oŰfB��̈́�g�7���Ge% 0��|���9�M�G�1<�5��]�J 9w�C��O��u]
t��|�(V��%d�g]m�!�Ͼ\�>[���L2l�W�)�seQ���%=����Er����FW)��R0��a��n����������k�� ��T��iO���ϡ�V�fy�:��:`m�D��3������Y���R�`¶QN~䟌��D�p�����o�к��:� D�M��?�+�u�bP�^���>����tK���6#ʉ�|���7�0s�B�Է肚�?5P�<�}W����G�T��ٸxU�b���)�9�*�}�*�W�]U�>z�OϫG6i���d���������5�(���?�8�P�=�]��*+7�*�G����د/�Kl��s��������Y]�!�������d^~U�١$?y��L�.8�`�b�n\�eٕ����,zT︢\3��U������0e\ ^j��JM�埃����JP��_�c�B��P+�V����5HS㙘���eI����̦�&j~�#l�
C�z�QL�l`�X�w�,7=��@wr��@,�X���!�L/���p��w�m����q+$�B����>����	q���[،|�'i���H�7��	2���F6�N�J$<�ť��& �'8gTA1�!R�棽��).��w����I�g�u�o��vF��Dr~s�T��(�����˱�ү.�TdE�;�����\��ļ	��|�Y&��8�~��	�`G@(�1^ZzNq
��	EY�-���6qչq�ao�pL�r��N�!Hb��G`��n��S��&ɷ䔮gsX���D/B�R<�̤�k#��Hx�
��fCr��6�h,�PJGW11�WM���m�k��kл�ުN�����
�zc�E�IX���W�X��u�>(��R�x}�w�A: ��Ty}�4��s��`H�?���87���Y��J��y(�^���Y�/(�L��gΨ]S#�j� y=g�����ev��Lpu�νJ��!^Ut�̃­��-7yNT�ݩ	p"��ˌ��Y��y�s1.�E�1}�b��m�'���T����	ϪA��l�U�}C5�;���5`haO�n@#(|[\��J����\�g������v��ыXZ�jAZF���R�U{o�vNn�$�o̻'(�z!4(>���}����ɗ���܏���M��k2e����Ke Pt}�[�<֌R�
h���A8�8ߪ��i�H2H�M�B�9_Y<}���t���?ٟ��,�B؞�C�!�����潍9T��CZ�O�r�ի��<�w��;7���2�ޒ�$�ˊ��<,�&W�.J#R7ͦ�a���D=�������@	�\�{lG�Ć��X��-��iv�:OP�P`l\K;ɳ$�B3T�ӵ���YTώr�
�L�5	�m�+ԥ�J׶���7�����	f����L#�� o!u��Z��������X��jnj�V�7��}�l��+7�h���q��P�À���M0��fF�O�x�Her�^�d	�I�0�$�| ������� �]��Dj��K�}c��'9�����(U��B�b� ��㳚��(�67��6�îR��{�
9/8��:�ܮw��,h�*�W�n���a,����J�����Z���%�KN�>��هI�h��K�\�C�O��Dsmݦ�辅>��8��.M�_#�`�3��";C�x�����G�@��Dי�ᵕ٬�!������BG��
G����^U���U�P�#�U02����{q�r��L>�LL=��!6���{x1cq�� ��{q���J�����N^�j�ǆK5�%`��:As�f������Q䔕��\�]�8> `�g�����w��e��֚6FoӘ�����/���t�!�1�kc]��2��әHa�$:x�Y����!��]�e��Й}���Cx�_fs>�N��L�e�m��n��ɚ����.�t1�Ȏ�t"(vW�giȏ����Et�����̪���RB�����^4��G�T�f�Xԅg{i�؅��L	��o۝r]��y|YuM� �/��%�ޟŀ��"tu0��'`�q��1(���m|dN���f��j��<�>@E��rEՙ�w5��>�V��bK�����f>���i���a�z�����O�5��HNH	#��n��8}�Pil)9�J�9~�z'Z��һZ�v�9	G[c̯}�P3&x�C^�7�\fz��������.L����@�m;��Αq{��8-W*�'쑃ok+�21�T_e�U�<����&[z�*8������֧��$�o|+��Y�A�}�����QRfd�~�*�颽�+t�����tx巧/����D\�*�p:ʃo$�Z�;���d����h��P �mowp�9��T�hc�gh7�-�T���W��W��ίvr5S��R�AQ8��+�u�I�U�k�q8��{(��}N
#��t8��Zp����6��=�hB��3�(Y������)m�μ��W�ь1Cd����rCԓW|z�wF���{���M�k�q�nҦ��\�����j����斳��BF��=�i�ܔlBvLiRˡ}�E�̧?�~k
���<���VsH�̤H�3¬L��J��������G����c靏Y��O��wq�_����Vm�C���Hn[�E9V�7?n�N��T$��|�:�&�ao�6L_����c��4lΘ1KikO���b	c��f�غ��f�V���.<���߿-+�d��6��h��P1��\��9B��$�����1 U���a�C�aV��67��6$(F���n�ݶ�������Q0ϗ,y������Z��(�|n�fN��M�1D%��BL�N��K�����T��2��T��j����:�pw�~
󷖣\������Z6S
�d����Qb�Ϣ��%�)��|�v���՞+����0I驷؟g�1c=���� u�o�'�}PW���f��|X�1m����T�m��3�t�7 b��l��⑱;f;�ҋv�8��!�ZNB�fSgeyS Or	P��V�#��1:��ghf$l�O�d�744k&��~m�� ,1��P����;4�!4�(x�ȏ�Re�IP�E�x�ƨ�����;����*�e�s�]�v�EG�Jl��JI@� �!E��A[?���P7;��7�6�_M��!��j���1�m��ِ��@a$6?u�<T��K�p�4�vI�A�c�gD�����JE�Cγ�[�6�st�ko�3d�7C�T�ӊ�j��­�	����Z�`m�~K�Dp��޹����_��+��cA���eLum j��w���&ʝ��� bw�B��/{����h@Ҹ�K>����w��w����m�k\CZ��p������G�d�����|�/�EӁDL�qxO����<쬍u�}	Hi.cp�Z���=�u9f���]�g7t�;���j�5B��V41�����{�SW���G� CD򶪾���,s��kr�~�?pR9~#~�ا��!q����c���*r����0=�iG�?��8�)�p����B]}�3_�1�Xq��� �r8�n?�^޾m+J�$�7Ґ��c�n�1��]^�
�n({2E�ǡ�Oib��\=1�5F���@&�(�0��?���l�Cl�������1�)}�R�p)+��m���T�[��N�0%�h-����.�B����9[�t0*r�e^l�MsO��6J@錕2H�1�M���  ��y
�2o�tS�"�`�K�n��8t�93Xޝ�|��}:q�x�ʝ��J�#/l�'ݻ#j6�fN���ǋٕf��?;13��)�������O��{�wC�h��t@a�Gyz��B[]!��%}�C!�aLf���b#�@��1�?��1�n�{�־݈[hWw�N�Y��֋E��Su�a�h�iŁ�&z|���+�N���Hd��(�qX�P��2ѯ�A�~��D����ǴhS�����2D�tH]tw
a\����נQ�6�>,^�Nɏ�|+8��J��ѥ�&�V�H�L�	ֹ�ᴪ�s��	�k(����0໣�9�/��rA�Js��v:q0S�&;�.q[��݁ ����§�'��џޟ��C|�[R�)��ݤLĝ]��;���҄<�r)�I6��{8]�\��c�%�T�BQ�^K@�K� ��l躞�J�#��~'����f��*un�y����󰲀�J�x�ά`�d�Jxɲ�N�����ֱ��Bq�{�>"S3@�'���ҋ�;�@/E>�l���ᶮ��<�|C4p�i�h��n|�T[���X�g"���j������D�'��ت�w/Ux�Le����R��z��uɦ�/o�*�.��
��~J\9G[��ǚ��K���H�R~�V��^mxn�m��sI���C�b�hAa�jF,�XY'�R��S27RBi��rV���S��h�VZU?l@���q�	e}��z��JW٪	������(�����Y�/��y��<�Q>
�Z:��3�S�V��V�����0�9��Է���AT�E 1���3G�QZ��0Bs<�uUw�oؼ�/��t�~�m\AN_	�6[���@�Iv���+s�_�iӥ|iF��۷E���(��E�5�w�u���X�dvv�[��EԈ�Bn�O�m_G=%�+V5��@��4�z�_�ۣ�����,"���֣ӏ��N<#`�*�Df/jE�'s�I�b{�u���_���P�j_*Y��!�2�p�r����o��d�t�������� �O�b��͑��W�����$�ل����B�U�ڶ��cB.�ڄ[_��w�u���D$�"e�g�(+e�J��K{r�ۦ�V��X�z��G�Ӥ
3�]ܯwnW����
�i������<�'���C�bۤ���A<+X�T -�ɦ��}�;E5�>�i�'Vi J��#��3���(�����c�ё��o\�w9�
��j��P��'? q6�cVjB�K�9�,�hb�mì
I��1o�u�XM@s��hZ���:���l�$Q���%w;`^"[�����ttR�Ǽ�\��b�-R���T�A���棨��W�-om�HC}����Kn���n|��8���q�|�����К�0��p�v���:q�Zmg!�Сgѳ��
^ܮ�T�?�5�����py�_�i
K���x:�
Te�	�=[�c��b��s�-����f���l[��{�K�
�L\��/[��/��J���V�K)/�kMI�r���<��'�uC��Ή�V���z�x����������z}Q�������i<Jl� �m,(aV�;�B�o�N���U'��M�vXO����3������ނh,����R.��_�Ɋ��t$o��ND�`�=�ځp���}щڱt����jPn�N�ou��) ��0�`����.�M,k@I�^��^��T���Iu�e'�^�	��ń�@��+�)�6��kq�~�Ƴ)C�)y��0�i,��Ժ��%�X5]�Nʡ�o0�u?�1c
Tr>(Nq*s,|Ⱥ�b�������̊�LMD��$�#�V�5*�j�X�G�j.��~�W�����3�1�Y|z+��g��V��I��HQ���}Y�feyL9��iV[���g�0�d�@�<.?��ʨp�=��p���>�\@���(ţ�*���}_fQ����o>���)��Ze�M��qo��VM�3\���'���s�_�U���Fף�Vľ�3c�V[�hLG��f
�Ͽ�G�rm����S����HP�YC�$(���@,~f��!!1��z͝"5'��������8須�rύ�.x;��N��	3�۸���U�)��C��F0�@�Dx�zj:e�_�W$,q��s\�. 4}�\�'�����|�Y__NfЭ�e�Ut~g�%£. S��=���ݤ��Sp]�&��E�����b�����A�ҝ��	g��x4�����}��B��b�Շ%� �<�?�W�F7��)����$�����U�M�~G���MQ�}p�`��6扠>8���f�.��:� Ɓ�c������L�F$����k&pr�/;�(�\.�:���IO�ͷ�!	�mG����4 #��6BO��.�x�D�~)��ygO߉��0�&$�bs4�5��l%q|��:!�PF|6����.�{J����$��+&�b����-9���4���%7�V�i�IR��Ѡ&��@��Mr�5��[��	����ً���L�ȹ��W���ZY�C�I��G�I]�A3pB m�J�MN �r�������	V�c�|dU;@Oƍ�R�,��o����]:̎���S��4`�^�i��[|,0�ɥ�f� �3��>��`���>�`%�x%A{�5C���"�ˉ���zmƉ����u��~ԤNl�JP]i:�$�mp��Y:Ɖ������;��x'���ʦE����� i�)�T��kTr�F﨏���\����p� ��7�����6��7�S�Ʈ'G�[�{�o�>��/M��U75\h$)}�&uyq�#������E�l7=�l�9̾<�"T���YA��?�?B,Yw\����=��r,�C�K�9�y̢0*v�n�AFx_���i�K�ݽF���н����C�P�vcP��޵d�$iW�RE^��_~�_� �����\-G<u!�ܚ=��ʹ��,(M@@�P�&移�)�j1�hK-6�]'?S�v����g����:�i�d�獂��=�h�WA�<G_����ě5�L���Y�P�$�Tf�؀�ࢮ�k��1*��Z"*�%�؇���4� q� ��w�B�C�$q� B?�K֯*{*��?Ws���m��ƺ���u�kX�YNk���@�uh~�E>�*c%1j��ϧg�Y��-w��$�����b<�շz3���]|�5$
�������%D�SP�yV
4e��t�k��sZ{׍����+�YD4DD@��� Z���a���x�������,��6q��}{�n�Q=A����s̿�G�'�N[���l:ڏ�B�F/X��a���?�����:�@F��9��BW.\3D�-曍r"9Yb$�D���uK��Hs�=;���3<�C�g�ޠ��� ��JT��x�?��WA�#÷�s��T�)�#F!�l���$aBh����"��s|�)h��=h��s�e�qpn8Nٮy*���� �bw�h�E�R� �?�����f���'����ɘ��l᷃���O\Ѭ+��/�)[���e������>9�if=���P#��i��$Y�a�y�@Uk�b�>�fV�:)��OF��aԂѰ���6P��)�"�l<Q�\������EPlʱ�؃�#�/$���:&uV5����hkI����Ţ���s{����&F��uHYuA������Ǥ�?y��U:�>��-
[1�����X���Q� �lԍ���C�� ��y�7��Gx�#��E�����߸2F��8��м�퀯4�"�u�(�&��}�j���ǹ\f��E>�9i�_������y/�V��ت���ׁu��hp�\�t��L͆H���G������$���\��,�T�:�kޣ�c�ӻE��H��R�Dmm�ei�'i�[�3WM_H଒�s��қ��H��f/R��7���M�i�xZQ�k(�͢
]r����#���H1i����ujL(4��Bط�~	4e�+�������ST�E����e�Bm/��}�G�$��"��ښ�A����+��V�d�\���8=����ͰЏ�$�)��&H��a#��[4A�'9m#�К&l�o$+��;��]I�	=�=.V���8��1����������7(ַڣ7����t��xV�/�N5�e6�-� �&��@�8�!d>�(.���4�V�7���(!/	j�^M��X�@���BPWp�?R���bk��!�de�o���o�������A�01��L-�-K°۽R�n�ua�iV�
�%�ٌ������C�B�Xw�|*��܅�G���7�śIKva�J��/_�}�փ�/��*�u��J�ҟC����5(QSt����<��CJ������c<_��<�=�Lr��lm���܂�������l&4r�vB6�L�fa��yz�өR`�:���Li�C�iو�����
:޻l�X�9�Z�lQj0�3^'7	16�!Ѯ�s��c��@��oc��5�¨���	�7�D���|�=�Z1�'���o� .��B�����X��,�K�Q�q�g�xu�\����2bq��xP/;�3s�����øJ7�Ș��tY�Gr��|�HX_��y�>>C�}ly��;.���C
!օ�o�=�=�%�0֕�C�\�x�VJu_���ȅ�7�zLb��5�X#� �9����X�!�D脫I���,LN��k���J�,�O�h����H�,ζO�*W��L6�&K�Ւ�!�Qk�!q�j�k2��(�t�n�t������ǛdMr�҇�����b�*��}�3�:����,��� ip�7]�����4ǀ�ϛ템%	'�ܖ�TΆ���4&�j��ƻ��u:9�������[�3�'� ͙�%>��O��9�����F)��)?�a��2W>Amm vy�,'P�[
ك���k8�5ߺ��N%~�.������!l;�^,��A�mG�H���6jS�l�ˆ�Q������W�-���ظ�(�B��K����v�/����\͗��L�C �aڳ��v߶)���( X���ĜL4�r��VY���I4y��oV�m'D�����:�~�q����yk�9�+�����k��	b
8P��}���]��y�-{���J��'�Ph�����Oo�H� O��=IZ˭�+���بSI�5�%d=&�;�+}ݮ�}�b�S�����ړ��Wb�vƏ���Vq=[
�'���0�&�7Q�[�I�ڭ�[��j{�<�|��y�c�@�N�[#({ɞ������f�?ss:5o�-:� Nڴ�щ��(	mh��0���[�UQخ����`�4SsH�~���5���.�R5C�˜q������-O#��fw�BY�u����=��z�z����M%ZY=(��Wr����y��z3�c�FN?�LE�SK3�p��n�˝�0�v��V��7WE��k86�r%G�'�-�}�a�1:�j�G��?a±]�q|��7�+��3ANv	$W�BaxD���ʒ����ᔸ�96|��ayH��!_=��{x4���� ��o���\�x(����f�/���Μ#>�.\��j۞®=֊j8Hx �X��(n�Pη��\e8:�-�eR�7`�\�s7M��`���V7c*޳p���3��l�tA�8�MG-Qn̖�ڬ#�j�%2.>K�����B$��mԫQ��_���	�g_���[ӋM��s�!r���J������\����x��RR�h���KXeI��^��VI����6k��7�D������[�'�7��=��k��,���
1�m�	0A�*s&�!�;���~f�27�@�gB�dqT5Z�JߥN�e�U8?c���u��/?\�y����YzQ��3����	aok�����P��m!\���1�S�/����KTwvC��4�%�0T��U���qMQs���־d�;��ǭ��+�\�%��	�n����}��x����a���E�VX�5	Zb��"��Xo���.x�E��`�PbH9�5�m�8xM��ڇ�.�x�1�-"�L�����D�4�ׅ����J���.�B��"���{�K�Ё����Z#G������:��P�pN?��ID)dN`�Ĳ�����XʾFl;� �ĞN۸��I*:>:8m�cc�/+L� �~i���a���Ow�)�(c�a��)�h��l�BI�ɒR-vR!�Z�Z��4 1y͕�q���<upf�Q)����d�w��mf�E0�����.���8Hb�J7�,���N�\Ťy�[5Ze�[��5��C�Z�^�%��������i��q �*bo��R���7� ��p; T�ץw�/�!��Ε>Q��>3%Cgf�Sۢ�K�Τ�S{��À��Wc���c:3�7���O��7���5�CKMgǴ;q�v���k���k�jڸ켖�Yҝf89�>y��T*'���_�B�Ȑ�����2Z�᨝6�����Ԏ����]�*�	�I⹈���Xɿ��Ps��ح�X�S;<�0-;���n��0r���(����Ξ�@^P/rp�UBU⧲����_���h�+(4n4�跆���?��J��R�����H��Ig74=����L��g��
�����}.:E���-�ϛg��Z"��$>�.�G^�Y�`�E���u6��_���N2J��H��Rk���>���>[�x{!�/�W<�m��%��?�D԰��<�D7�.0Q��{��B�r�ݥ�ɡ��fF��)��D�n��0?`�� �����.ZH�3��+��E��T �?�=�e�s�\FI�=w��2��9|��ml9b���8njf����hQ0C*=���B1bOۛ/�;M-�|0P
;�%a˰i�7�GM����� X4�Fl0�o7 ��tpA�y�;�û���qo]8���K��7M�/���:����C�Md9Jg��6��L,���D1��#�Af�~m��vk7Gv]ʏ�Ma]ş�:�;gv�ï�B~�t��f��{#�+�B��k�R![%��AVC�DC�#dմ�1]X�!��H���I����`)K�P��*�gL' �=+�NI�%M��)�I�����	i�mGyH�z��a��`��d���
��M��G��2�5�7����a)�M�a��wGb�[e�T�\
�ֵ�����'<�*F��W�
�
��ԌX�윆	������V,�F�:/��p��]���\Lb�:�`�7���Y1<��8eqVS��-7w���Yxwa��,͡�@���\��0��p��etJ#�)OH�u�HM�ï-�}�6q�(�b�M�@&�-��4�����\��eGB�	.B�w�i!�����V�fv�$6�c9��0�Ti�2Gt�f��|��K0���gw�x[��oc�_����s܍��\�����,Ȃ�U�1�	w�4I���F����m���&�EcH�~�g$�����ݸ9J��W}G�f�
���T{x�$�<�	h?��Sh����N��Ug��
�%n�,mg��N!D.���f�iy���i=^��7�Y�h�׸K�r�*t��)g�&M���IHY�]P��{K�� ��p�d����i�Ӂ�m���$Y?M
M�ф��mR�Kǃ�^r���3�����F5�bՉh��ψ7�.�t����閜����~���"�y���k�s/�P-\͇B�E�Pۧ��+�FU��SB���H�[�W2���6ӄ^���c���~�����ղ����<p�&u��y�W�x�^m*![<[�� ��;����ˈR���%�]x����w��_/�JVf�`�y)�8#Y?Gy�*�I�ӫr��S �|�R�Gl�_ Rq1r^����>T,���w��MH�]�g��u:j	�A��B�&����ak]�?OU�J�RA�1cS�5�p3h��3J�+F=42Ne'���u@���O�5�����U�o��H��f%���	� G���̮���N�dFe��"�l�\�����΋���f��oˌg=��V�ϙM�R4�����A��="�����THaNlZ�
f����J��lpg��\^��6���HI��̚$�C�\����㞽���9�d�s	+���d%uw]���|���ۙ8T�QY�!�g�>
#�c�D�pk�R�}a�|�{X�c�S�W���~䩉������q����N��X�VB!�!sT4"�.��k#�K�[S)�u|Z�P���v����/��^#��B��C�����ࣜ���Z���\������q(����
�UVcɣ��R�>6y�>��h���և vf��I�Y���zM1��Ob�:=X�[�5����D.��N9C�QPn�t���:�?|��+&�i���i��6��)Omn�^��|m#�h�Š�)<�^t�4�5�꩸�w��s�����B�x�����a��Zx�)����%ݥG��]տ~�����L}1٧�I}�jf�pj�.N��
vVJ���%��j�-�uo�;;B:�w�H�9�ʚE��?u�T��S��l��XMT_����&0�K����V��q
#{�0�cG�_P�R�~���a�q5f}�u�8mF�c�`[7�ݘ?�U��q�Ôt�9)�C�~vQ��#p�&�"]+-ܮ3���)5qAXx[n?6r��rE� ���Vu����V�s`#@$Y�uV�(vU��5ţ#"���4wFT���<0���F}MR�����WG��q��㾤:Iش�@f�G��.U���j~+ֵ�o��J�� �o���|�JΚ3I��tG ���3y��T4�6��s_eʠ%k�3z�?%W^P��w�'�|7c�Ӫ�l�3��fL=�S��Cͮd�t7��N9]�d�Qkc�F�$�f��8�q^��j�T��/�?�v}�G�`����y6�ArU�MYl�N���r�g[5�\�&jۊ��x�]�s������L�?���l�Z5��F���lL͖G�`�E�����5A��$�]�l+j����.�l�?���t��a��=|c�D������;��im�lB�K���r�![I�u�|:��.LZRUݲ�Q�Q�;5�WՐa���f����Ï�}��}'q�F������ը=���0ĴL��$��!�Q����R>z���{8X3����E�P40D���^��������3��'=^Ӧ��M�ɍ9�V�\�%���k���t��-�N_2S��i20��S��B߫�����*�kTb�6�l`���fޱ"糢yRA�}�/�}}~�bҹ����@x[�j�^��E#ʅ��A~�b�.FJ�9*L��A�WXǄ����͓E�{(�>�Ԇ]�kk�Ǌ(@���P�G��赘1�ܹú�����y��V S'�ms�,�TdK�T5���f���lVy�IglG�N-]�J��!�Й�q�z]=;u��Oj���%�ߕ�WH�`5��A�ʏ�~��W0	��w���;
�-� 7_������%���R�@��q&S��XO���%�Sq���p�[�G�����C8����)BA�ѵ�tX�R� ����J�Ԉ���g3@�p�C�d��%~=9d��ɕƷ���Ts����!޵��nF�i;y
#K~6��¾�\�9���D%}4T��2W=�G7.wlUC��5IEܸj����X1�NhN���V�������|7�$��ꛯa�
��������,(d����w{�MH�@!��=�~�2���3��UU-LrW	��}
�YQ�٨*���Gj>��,�`{Vc&|�c3ٚ�$��ӱ²�9�������Nb7Xu�����N�|TDBH��C���_���L��Q��d���cK��GiYi&�hҥv�Dkܾ�>h�`A(I�� ]ke-m��e��v�m`|�)
+Fl)sd>��D_-��ˤ��!.K[���+r�µ*��Ϙm���P���H~�|��z���N�H�CJF���la>���2D�����E8"�[.���:p��C+�d^�9%�ŗ�V�!;�_�#�O{��؎۫�1���K!��jB��z<�|�|ÝrY�d9�T�S����^~4���R��1!�V��̄J��� C̗�&�|%֖(nڱ4�g���
�J��=_j��l�p��g���@��z��On���yQ���)"�#q_���8��]hW�n�� �(RM#��-���S�|qǉעM����� ��'�K`?Q��>��!����AO�%�φ�^9^��r�Tzq���O�x�����N2lf��2t���`�{� Y��D9x�dG�:���W�6g\♮��B:X͟T��z*w	�d�$j�3�D,ޗāE�JcBCs���	L���axϴ4ꊅ�M<��EU9[��тZN�8���Wzˮ�z��h�=h���#��K���6�vr`� ����I-�a�B|���<</��XpD�=�cq�r&n�\��ͣ^�M�3��2�b��DD����2�,·�u���w�$ ���1r�ڱ�T��J�>��f��˓k�����u����*+��YMع��YX��:�<�Εa�5���s����F2�B��_�a�&ed�;�5��X"s(}�`txu�k@ּn��O��Vj�vv�em�RgM������~�]���_�+���4�ݺ��{�$�T��Ԣ�l�ҕbH�a��D#B.::HgaX0�3�;"��>5D(�W���/��=˷,0�!cKg�x�߸�����k��y��@�N|��Qs��w�S/�虎�}���fL�qt%���jȗ�T�D�9���	��(<��=�U��r��-�z�*�#	�M�}p�pZ?��1�o
WtNHf<ē�=���o����[�밺B!�8�ON���Q��K���ݞ�uq?_�����.;3���D�~<�P� Ih�q-��bL,Ce�����mq��Ii�Lv��1���{M*w+z�SDR�ʏ�O�=�m�D���Ef>�j�+����@,���\���zA�߹zkf�;�eHL�9�b%�pz6�Bb�v+�'p��HrXL��oEк����{bR�����vX6������"�b�TZ=�m<1�c&������}H�6(%8��	�`\��~����L��4m�:^��4��(�qj�L���?pr�w��=` �A�G�J�'�QN�k
��41C����_ F��I
��VT�R���WݵH�քͬ��|��c��\�^��3\�2�,j�q[�O�0s�A~!R�VAӠ���+��P��ŏ^�*\�-�w�uNijD��HЛ1.�'#PM�߿-\Au����Ӌ�k��M�����\�[U�*�0��Z�RD�[�a�	��������2�9�ct�O�9�e~��Uy��D�7��8���n�%7+?-<�L9�W�0���E��kH~aߒD�(.?	��/���4����/��P+�6�J?:�u�����;@�ݽ蘀���~MW)N&�����X�yc�S��;�j��_��0��d�9M��P0;�<��!H��xKR���<�"n�-�\�q�n��H����i��e&k�ߟ|V���aa\5B��V}�Gݞ��f�{>4����{��ߑMd��������L��X�b,�^�B��y�m�m!n���ݶ�l?"4	��w_�����[*D�����d���˾J3p��⯂��A�����O-��z�6"�6�H���ԈA�h�$�����S�q�Q��ٕ�٥���f|��℉��t�UV��V[~������6��P�:E�8Q��~���Τ�P����	�}2}H�wZ%�5"]+)]N�Da��cB��W��~�M�QW��S=9y7gM�ch('�Cu}fF�C��R�}���}�o!w�v��%�jBx��ʊ	lx��b0�*�+���i]L��R�Q�o�Xk���Ji�Gy�L�=1�`GvR����M� �)k7���bp��ݫ-�Ɠ��B	:*5;.�s�����`�a�9�X�p�8G���)ѓ�/��xV_'M�h�G�j�oՎl�����:�Rd�J���Ck�y��q�:���c�Л�<A ��u(���ȩ��:[��㬺_��0�mL�֔"QR�0t3�T���˰U��-��s:d�W�6��Ϫ�2��D���_:(ypt䣬�,�^�e���U�\b0���S1�l%��۪��7ķ����)W8"i�'Y�Y���[J��!�^ᖟ�tV+Jot�K�U�~�G-��;	̼<��c�98��pQc���	�S����wI�4�D���w}�z�3��:����*9��D��c��]B�*��=EO�����Tԁ-��Ϋ@��ȉ&�`9U���ʑ�+Y�>�]�
�,�����݊{te#�k���qa)k|�P�A�h�x��������u#�FO��]�����u`�������X%dYِ��
3��1�X�ـ� ���C���R�Nu�9�+-��_��u�.�פ�L���]E�Xa������O���"RvL�
��֍@Q%�'|�+xZ��J��6��*�+0by�������i�����V��3�*������[�Ev�o���s_}��4�z	k�����ѹ���Ģ��M�� D>R�o�M�$���j0n������	dQ��i�M��Bƌ�=-
p�H؄���|`����),�дD�O�؃���ȡ�� i��.N}���V+f��63�����PXޤ��$ꔲ� �H�Ū��E!c�}h%��0��֖3L�J��q	���lDj�y����S\0�-�.��	��cxzôUc����3�Fj8=��>�v�/�U4�3�y��,&�|��x���6c��g��Qİ>V����)��{����Jī3\0\���#Ŋq��	������ ˆ��>��m�Π��㾵gv�����:2�z��#2￯�ړrY� �*{���t8:�|As�
Z��RQ�1�37�YkJ򅫃@��{��y�R�d߷��w�u����|���g�:��+|(n����P��_����5X�O��Ԇϳ]BM$��{=�(�}Z'�;�a���Y7*Qn��D���V�j��&��c��cj���;���E�tn9h�`ݕ�8���jr�ȟ��j,	@q����(I��WN o���T|@�2����	p�x��~I�&�u4��Z�жU��A�c���������ɋ~<��7
����Na@4|A)�'w�M~k��j�J5�c,A�%��"`�o��o��;�A�ԯd"����$�:=�$/G��~$�O��<`�
�F{݆W�+��4F`A!^�r�I,��>��_MN�
e*gwʹ�+yn�P�^���'|���-dfݙ{�{��a/�!h5�';�O^n��~�����$1�[�"���"�!fO�KRc@ v��,�t]d��0.s�� ��*�T߶������W�g��!(nݦӎ9��9VIP�<��W��	]9����&=�c�d�6 #od��?�GgX\�[����F#�j۲š������å���W��\�L�1��z]4�R���N�Mo��Ƴ��=�`��9dw��t��C�
���-�w��t@�,�;��s!_�X}�[*�.��T/�a���P��[�"6����a;	�`�����86}�W��Pª5|�l�
2���e�ɬ��[�W�;Ӳ�O�ʽ6�p�D���.�sP�վښ���"����7�>��,p'_��R��WdnB�/�^o�$X���F=�ߢ���s�9.3��n�f�m��`gg�v21MV�a�$�R�}7�R�Zʱ�� �NCs�ȴ1�-	S�g�5�W�AÁP��x��lnP?�"7�
(�*�ϥ��Tj#4y]��s���.eCR�Ƹ�BvI�X��H.���� n�ڄ���~�X�;��-�*N����5RV�J�_�rh &���)�1���z����S���{C��Y�|(�Q҅�=5����p�؃b�3#���?�P��~�� %�,{�x���7khS�ϯ��T����i=	�C�@��Nt��m�J�7�0sM@�/��IZ��Z��1/�<=��o;��t�b�
�� �j�/�+=̺`���a��]��7XR�����@�F���v�p#�k�y��U�s�����%]/�2��[�� \�a�g�y�E$�,�����z�R^���d{�:�Y�Yo�=�Z��	�}��<K~��\!z�N���l_X�m���H�}�{���Ț�����mv���R9���Fr�"\�twӡ��0�!3q�>eb�g�EoX������<kV���ъr��W2��q3���:�܏l[Bo�,�{����KD��C��ц\��I��g�ѽxyp�~3�������9�:F�!˸C�dҝF����L�+4�Qg*��mkl�h��&Tk�	����5;egr$�|
�O}���?���i���t��8ϭ���E���Mޒ�����;R_�E�p��$�����Lc�ι>n&����`��Z��g!�o�ҟ�����W�����kS��,���)���\Jn*�	��I�I���D0�V�8��<�S�S�vE�Z�< �X8�@zF�WT�$"TE��Z���){}M��RG��>�;\�����V��"�w���
.A87�[��������*�a�/�����Z��	��5��Or���F��7��z�A�Iʄ)
������g[)|��>�`1�6�u�5%�6W"�:�gW�XD��J�z��O��\���~��P����ܡl��ĺ�Qg����s�N�M,d�D�xuʟ}
`R� U�\��
�R��u�|퐻��*��7������Į�f$�WG��޻�� �cd�Z�q���>��\��Q��푴y/�V�y�J:_B���0��tO��O������t���O$�o�!:�i��0{�˸w�i �i�.��o���7Ƴ⏾��bs�G���Q��и�L��7�6�0X�`ȱ�j�~���0�d���UDU���h�_�C2o��O�6��9̐��@N*���������]�x�B�|� ����^�,�SL�ȼ�p�0j/C�#��kԦ���y�n�GC����� zi*���Q�f��5��	�n�d��#H:+)l��uP	7�6�omB������('�E�v�7��7�	��1� ���%lA�1ԫ���I��#'��&:Y����l"�E�a}ΩY�����R�� k����*�ݡ�
ڑpX#��M?mӺ�
$�O�V=��.�m�
7��n3��z�z�/G g�)�u[�qZ��_ؤ)Si�� ����%�p#b��'�N�?~�Տ#>����x{��Ij��6Z��e�vDA~�I�5:jm^B������+���6���n���L7����G��0�fe:�n����S��ޘ���� #���Q
I�%p��Dj-pF�g��J#_�b%!��pI2~�֎���jp7�8`�"�Fa�V��1�W;��c~��3z�P/C��~�Lhm�e↠�:����b_rT�?U��eFT�!��"q�:J�S�XcR��1T�#ze�����Q�g.	ujhjǢcs��Ȋ�=��	�E$�u�D}�KҧDm���c�G���a��I
'	�=���r��+e	���荨M�:f�DW�W/��'J>q��D������<e&�ܳ<.f�8��%+ە^'���H��肮:��/��Y��%PG�:*R$.��h�^\����dX~1��Y��J������3�B����+��~�)79��j������qr�/����s�d�����bJ�bf^��ES��Ǘ28;��j߈����i,�]�(�;��ӎ쥭�c̻���/�Y��f�e|��(5�y9������畖I�t��v)���X�ǌ�"w#��r�u��j2L��.�=Eð]�ɣ�P֪�r��6!�j=kr�A���;�ؒ��d�.�5���,[×�8�lϱ�X|9_Ab\���:�`��ƞ�Z���T��Q�:�US^��6�S�Y?m�k'�x�*8��F�R|�y�Y��"��Z��j�:v��K�t��|UN 2ѽZ@v{qk�A�#5��)q�N�+�Ol��f%꟢7K0�4	��:I�������U0!͆�.;�D����٩݁��?���a�/���Krе���=K�Y��t���M�Z̃Yze'<�M��SO��$��ݝm¨͝��i^���(�̻�+t�Z(�-�@p1@!,j+}��f�a[k��ɏe��2V���C�$�U�����#*��P�%�Q}�h`$�Sbi��7�Й���r���;w�� t�:��ǩ>X/�g��	{&�JG���"H��y���k$É�N�{8N�[ߟ�t��"m,t[d!,^[�0� a�O
fM���0{�}���2�Y�+�$�0�vV�v�����<���3����?�����˘����@u.��,�﷣�q�S0����>��j��0��Y�����;.T�����Þ�lJ�C�����xuO��%��@���u�`��|~Y���]��@'W�	y�<�A�#�D1l9[m7�J���r-O�I挘>�*�9'��F�b�'	Lsh� �Y�AD�����(�u��0��UY�y��<H�3�\������l�By�<S���L_&�̲���5��~��/V 0P_�]�E1!�4��lAMn�=jZ'܋'K�U��k^�ݴ�H��{�r�o�A��ךtRm�.��se��);�������N�3w���&{:;�����\�D�RV}�\���]ѝpZt��6n=
/ ����.cͨ �~�A[�3�!��>c��21�X��ZԶy��v�a!���\�Qc���)�hu��Y�iH- �=��H��@�λ6aՅ��Z����񸽺㙷,���"��p#��BF��V���A`whI�{~�|��[n/)/
2{>���UG7=)���u���CӍKҢ=h��oM�a<xB0���i���C��D^�(�y�Z����zlm�^��/�3 ����:�c
��>/-z�����<�|�V���y_�b�r�� xT��?�}�A�Y����#�)�����ࢷlĮ*�6�Ǟ�		��%f��h���GM�����%/ci����ٟ�(��̵��o5.ŏ�PH�iM+�y\\�鎓���H���M�����[�9~?�� �I�e-��%>�B�J��av;��E����E��R��B���]�݁F
��νѝ�сeT�p��ҝ�\hN*�T�@O���}s�+�g#� ��G�8E���qӱ��gx��EL!�'���ӂ�|m�r8TNZ�?p^-���}�cl���N�J�`�C����8�k�.-��/�#Ҧ��� Ns��3쑳�#��J1���Y����t��?AY��>��2���l�J��[�(��S���F��l�`O��iW����D><�� �i��M-7G��(�ʷa�W��/$�W;�OB�Xe��ԋU��ńy��S. ƀ̝R����9I�{���n�����Q{��n!��n؄�.I�Պ�-r�M֜_�-$��iH!F_D�������N��)p\�lp��N�h�O�4W���=̜���r�D����)�q�.���iѪ�W\�!���&��
2���O�I�J�S;���}4�����m�o$�����5���M�R{�Y�<���I��� ��z�Ca<rW�]��j�6q���~�j���+�ZԵu2�zVb	��"�j�T<5��y�Ę��Φv�1����5��b�#��*����=P�K�/Cqkz9T6��q���V[0\��B񛔨�S��w���1�=wVTsz�*{�'�T��Le��f�B���zfJ6T~�-QGp�1�o+}� �2y%�pl{����8����#��X�rzr�:2۝�rA�ۘ�X�%��K�� 4w�5��̣�A��6@��P���Q�z��d�,rW�'���'+�kj�c��˞ m:*��3�Uű��\�`g2�8������:#UR~���RǌN�>�����^L���O<�LZxt��!x`W1�.�B؊>V��
AT��"j�7�SO6�JE�)��G	�]�e\�1���C�VlO�ʭ(��[O\���9U{�K���A�{Nx��(�V� "����������쨯�d(.���u�2��:Lh1$��4Y}�o�߀�Mb��+D���qng"�d�4Ԇ��\|��Pj+�`.��.F���@�P�;�^ځ��e��;�?�6{�_'1�!�zK��q4�+�b���S- ��s��]�ƍ��ˈ;�.�,)\��aX�'�3n*���٭�m~K�Z����*;e�\�S9����K� s����5�C,U`g�< ~��i�y6CTg�]]`d��Y�����l��*sݵL�&��"0X7t�"�n��el,{� �"n�^��ׇ=��ħL�Gʣv��G�c�Y`-�	���I��x���b�k^�M�^���fˬaꈀ�0����a	hI޴[+���������Vٷy����R�)��R����CEߍ��
�a��0��2�#�ߑC�G��r��H%�ÊYty��@8�C�CK��dDY��;g
��A+W��u��;3�Ge?# u�W)�n�J��y�\Ƞ���=xu�#�UO[�>������%�f&㟞&:�Лw��9�\�6 =?"b��yӒyX��}5P�snLѭn����{2�kSe�(���^"@�˵���8����
��(�°�Hu�p��L���ÞK^ @c<}�L��W��{b��Yo� U��x�y�����#�E%�O1�m#.��
#;�S�����]rs��)rs�i�`�����a��>(P~�x�M�j4 G�;M�8�aۖ����ݪb��>���K�aw8?)g�7\������GO�n��ۚ�~c��	EA% ���d
�4Q�z�v�^+/<;�U��R�b���O�x��L�1O�u̕�
���UY'��fm�53j�X�$����[%�#6���t���J*���^	0��,���IbnP�!郓���w;/�
��v�\{��q9�
"/X�(#+m��(�7z����ֽ,�U̫�!\a��r�H�Ha����\<�'Z�Z,W#x=h�I�bs"I���q��>�o�?,^5��Pz��)k��j������T�}�%���M��r��Ȳ�$���~w`����a��hO�� �X���~T�LR��p���=�P����Qf�ةށ1���_��zA<0BcG^;2pT�H�莐�J8��[�����iC���;T�\���T2��}8O� �����ǽ��_�o[���e����"��o�g��~�82��	��'�1��igv'U�Ѐ8�
MV���B�3�%�23�ષ�<Q�7�ù�̢��h��͚����L9�I;�*�[�);����P!�@�ͤ����+��$����2knU�H����{!61f1<�C���s���P��Fo0N�sDȖ�y����XcGh8˪�E�+�H0w�e�����U�V}z�9ڥ;6�}��K��PbG��!����<����ze�v`?�Ղ0���Q��J��f�*2��h��Xó�ϫ�_�"^�Ϝ:K1�D�I�m�"��Ղ:��=(��[�Օ�?�Y�8��Q�[Q��i{OG+���B��k{ѷ՚l ��!?��.:$��Y�L�"#�}��%ֿʹ��o�X)�"���YR<!���|��Tq��X��r�zH%��������/�H�?���ܥp���[�b�Y�Kʘ�vR�F�@^WbP���Q�l��l���C@	�g�e��C�$�@�m����<9q1����g�,��M�J��cR*%�����o�W�Nt(��� �u��IzE &'�5�������(�/O �.�I������Ĕ#.ܮ68�0�C���y���l� ��@'r?FF��b��BKJɐu�q�/",&��;o�p�zߊ�D�k�1�a�:�I�ڎn��d�M�FSܑ���Ȭ�4~���yd�r?C)�9A�V��-�w�����n/��sٖV�Y#T�����=���<��uc��_���T�N���dx�$���w��5e�ˈ����͍៬!��3>"��F�ds�^�\^�,�M5fh�����Y�Ӳiܧ���l��8�>��nx*~S�i5��OWh�� /�}a��&�y�� GU�nmˢ"�n3f�Q�'��5��u��x�	4R*i8�!�PM�>��;�M��Eάe��z���.mmGOt�rg:�G�����N���4��/��D�C�/۱����JXC=�����;y����[��?`#[Ս�]H�|� �O�dz#v=���_���2�0%�@Q~�'���e��g�y��,��Kp����~�:���n^s65�"�9M�F>@��	�hQ�[1oS��4�l�cts�;RR�S-��U.���ވ�{o��w�������mۤ3�ͳIFy�L��'�z�&���ɢځ1dɧ���F�J�6DS�������nh��4�Ld��Z��K��RD�M��j)D�`���8���ݹ
�9���C'��N �#�2}	F�9)z��hdURTmv0�&�����~�����MkN��&�d�"��<f7\J��?:��&������?g����������d����	n�ϫn��_z<�$,S���XD��M7`|z�MI7p���	�>�b�W�z�1��H��Ģ�e�w
e�I?k��A2u}�`�}5m��_ng���k��Km���w
h(���5�N�J��;���TSGi|�bHᥡ+`�$�v��Sl�k�X5i�w��||54ja�����pc���+F;Eugj���%ٓݦ)n.�_�]q�|4�==�75�uӹ����S�}�+d�Hf-
�lP�;�'�f�K�j:u�����ʵ��q+}�i��6}��.&4H:��W�I����Z��bO��P��t)��X�ס�������M���u��R�?<-�\JA�"L�VY�WP��?������>��6��+��O�X�f�G���j^ZI�)�^�����s�#̒k�.&�������q�p ܵ���C,���B�evn�(~E1=Gŝ�Tje^z��J�*8~�e$�/��@q����.�����cpX^��gă�j��r���w��L�cլS��U=���}!9�U���V����c~�F�?��R8�'�^�{�;���D<��l]�}�3�_��Smb'8`��Q�x�TNq��n����:�\�\h����)�g�k�-:�(U�Q|[�pmF-��?�gs��Z�7"��mOfג�ۜϦl�{��Ȍ�JE�È��,rd�{�Ho�|�#i:A
���>2�tL�mZ-���X� @s�NB}��!4f�RQj��U�uD�Zn���r)��F���]j��=�A���:�֟;��%���*W(�'��}�H���g������w���[�짩EU���B ��	B�9}����t�yՓ���ȷU�_�4��!"�?�$Tqj�*�2^p����Z�s����އ+İ?�)�8>��S����/"F2�NV:��I������D��<^7gǧ��W��j�9���&�-��~�mwr���U��7��w�U�>�cPR���}eJp��Sl������O�߉-�%����,���<t�!��j�1��>3*�jTv%���	&s��FƮ���v(�����I��|�/p��{c���Y�V�-�yzv�D	���v��|�N�˽U�l�DY]d���/�q~�J)�}��H���u��ET��V��������ߖ�r���!�j1qW�@v؉[��/�a}0~k��Dz�%�y�O��4�t��;��m�j՝/�Ե����7�����b��_���.�pÓ����%�1��z�;Q�@� ��Ed�@����6b�^�L�3[�4���V[�42�n/�x0Rc>�e_ZM!A��d��� 2b�!�􏭲"�×;s�3X���}�����[�m��@nw��'[�y�ì�w���tֻ����V&� �YQ���_~J�W\��H�QI�q���d��,�����aX��j���f�G\Xҵk��x�aS�� R�;��Ԡ�h�q�;�������K����!��@R���\7��ilK�}i4*�YNJa��f}o�a"M�!R]��G�/���R�q�ٔS����?�OhJ'����ڼ .Ai�6�֒(#�I+G�AUn?��K~vE���?�0JD���}�����Vs�k�30�R�Q���f�<O��JĐ�u��Ft/�G��a��ٕ��H�1eA�G1~^�{&��k<����l��Q�p 3�r�J�}ʈ�ExcG�O�ܨx�����7����א6_v<,׋/Hi�`̝lH���H/�% MUrd̑���ʇ����]�G�V�����J}$���{a�غEp�#i0#UU���+��ꀐ䫍�I����/!��%�LX��$/� �����c�`6�H��i�X�ɝ�� OA�'�����T�k!���˻P��)�@^���܆=MQ���9���1`ˀ�Zx9���p71���*{�s�[�Z����,g� ��$t��[^��g&f�|�1�L����? V�>��-��ڿ�??tcy:JG�D*�k�hv5x��3�9M�۟�FB��y���w"�q{r����Xy�<�(M��j����b�s��ѕ���/��n:̘�g��n`H!Le7�c��O0F���v���L�k)}lX�w��j�ֵ+o��2@�D������w#s^��D�I��9u�_��j\�?��-�"Xk#��+Z��A�rsާ�ȳ�ڤ�>1�7k���C1ͩP=_+8.���TT��J��k�:\t��ZZ�Ŗ����m���W��r�
�/�q��M��ҋCL��g�b��G��.M��� ����{�{�o�.�����l��]KY|*p
G:q*�Y-oK'-/C��ԃ�[��1�`<5��
_C�b�Nj�x�G�п� ��U�╻�'�����V��KE��}x_*g�fb�
����G]�0�m�k5�ʴ,|�ԝk��j�$ֺ�k�Rf�1�МA��
é���EY"��	�R5������h�����?*Mp���z9��+��gR��Z�μČǉ����r����V���%i와OT/��4�s���.��K���+5�2�I�S�i���_)\*e` �s��,��
 �k���-��oJ3��FLPfj�T�Rz��M����w��{��jk�\����ys��!�������gա��
<�fL�_+_Қ���{a6 ���j�wH�U�8��X���������^�4Kt�UD����� ��X��}�f�He�}ͳ��u�����$	"->�N�DV\D��{��w�Z-g����X�Z�#���˺���U�4a�����:�
is)���a��:��k��}9<d��>�;q	떏%��ܠA�#��/����>�0�j߇���g�O�oa~���a@S�5�'&��ca����^B��\�(0}�?��+�֩�a�_�*��b*��-<I1��)z��W!�te�o��k�޺��_*��Lg����Ӏ}趸u�+�u�q�b�>���;ΡԼڸlX�}�Uq��)H�k$8L&+�o���b5<�~�D��d@�~X/S���^�g�0��HMd��9 �D����(:B�`b!�47+�	��W%�ѐ<79�A^*��aT����I�@ ;�-����,��o�i[�d��Į��9�)>�9����=��㭲v}v�A�Ωz)����b�P�u&T*\d�-�}(ʊGaB�n�q�J��'z��Y���������,��n�pi>e-��$k/#i<D��N̸�����
;w
��B����Y���a�B�\a,�4˼�Q���zLj����{o]h+�萶h��,���N�G�	�a�|v�2��1!>��������-^������F��
�a��3[���+�Js��KNwW-��]{h�!�ēr����n�dz+�0G6w���o2,��^�}k�ɥx]���1P�|	%|͢;Nv=�eW�ųW�D���[e\� ��3UCMM\-+/���hA.����2n"�,��>Ɵ��o��}אַ'QPx�2>)o�9ި�C
H���.ʀ���f�*�n��X�&�Y�,�j�H�z�g/*2����[Ė��9U#\%<5�W�&Iv��7n O
�'���c�Br	�*�0�X&|�-�xy�V��+�]C�����9���8�����������|��v��?](��W�ٷ�T݀�1C@��cq�?nլ�Uo��[*��
<j�׍+�3��¸�\e.��7ʦoZy��w��:�1K�����v�U�	�M��R��-��_r�;�Z�NY�]�O^Kn*��+z�g��	��!d����*ټ]w�Sfo�s�B��#Pً֗����Y��80�9��&��X���^yauA��LkW�5hV�y}F)��`^M�a踟�߅�cW�5�sV���hp�K����`im*���������h�7�<ziF��0b~M���4Xt�3����T��2���S���Je�]�c�{_���;N7�
[W�q����i��wј���!��X���s+U"S�`s'/�x����*��I����!�F�DA�����s�D�Rr�,g�x�<�y	�La����"8�����ke��Ķ9�la)����Y �Wś��`��8��v�z� �k�ԇZ��a?jJ.(����� ��y�?�iO����a8��s�X�D*q~���6nS��!��hY��Y��7��U��k_!�k�U8�K-���/%����M4eYҢ�T�P;�~�sa^���g�/ӝ��6��K��^�&�8Q��<�ؘR�bߒ>bH@ū,�e}��v	e P�� �u�֚��I��k9@b@�;g��[ҋ��U��98����<�F�5�we C��4�PU��|��bR����d��䄆��s��SM�8s�Ϸ̜	4D�(�Br�J���9"�W.��B���)Ln���3	�v賦㍘8���+��k u�͙������d���	�S�%U��S�L�^ߣ��D��d;`nT��E��A��f���О��I#Q�w��ʻL�޼殍)��&�QX�2��������{L֕�5�D�\��HI5���_c`�����1c�R��rSʇv�p,�ѣȍd��p���8-#Q��D�m|������F�ȣ+�ɶ��9x�R�R��5�s�v��"�K|G+Nh �8ة�;�j=�MK\��$��*r��/WH.� �]��y�x6q��_h�`�a'q2���l�6 ��SX0@T<�j�D(�?]`�= UP�qͱ�B�N�Q��:x�l�L��
�#�+�X �M"����~���:��2:-����(ڎo�G���6��o0l����$��J�C��V��ó�n��#km�}�@���z6��iB�X�7�P�ў?+�[E|��K6����J�dV�5:�n��k��r��5cЃ�֘o�i #D6�1SW ǒ���?l��:��!��#�Ѝ��I��ه���ފ�$>p߆��0�[�}lv��R ��v��*v��tJh�+�T5�� y�#$j�Pt�m�\�M�9v�Wy �H	IKɻ{w�W�vj��!������J
��Ry`ɼ����������9��ڈU���V����=�|Aq#cki�,eam����Y��-8Ӄ�5���qq��r����P=�ʩi��!�q��c����^�Qc������Z;]�j$��Uȧ+Ό���$�I��؍�B/ &{�P�����A���ɋO���v
1�;_�%M�'dWA:IL&ހ�24�4��1�K+�c�)M��	߱]ߐ����
�_�]�����(ӄ�7�E�w;�3�Ar~_H�+-Zr���`%��ʻ}�������|���7���X���C����hZ�[�m�H�UNu�=���4�Eٍ�4X��YA��D>�M೓�-'�~�@U��*;�weM5�ǔ*:<�Bb���H_H�ͫ�Ɠ�r�[��"��_K�+�謳k�����z�6�R`�C"oF>�k�>P|[7� �wJ�2b�=������-J@�D�L�UwG����a�fؿ�ph2�t��Օ�����9D�S�}X��v1���$�[vs�fW��}��p��s�[�GO
f=/׾����Fh���L���W�YG�P��iR$L'�����]e����+3P8�X��D\4�z}߾����2ܧ=1�uJ�TK]x��+ɩ��.�2��sR6B��cޝ�<�*�����[>�6/��_g�!���i��1>S�L�l�XbI��2D��a���E�7�W��4W���瑹�_d ���T�7��jHSYK��>Y�B�+x�х(�Q'B��0-.~��5j�f�ʖ�Ʒo��f���5�Xͻ`���xG�&�ϡ���Fd���C!���ai��z��}V�f
��̱Т���|��|�Жl�3,�Ygʉ�(��;�!���!��>�/��BDK[ske��,�
F��ކ#Fd���!�8������X�����-��m_N��eF�� j�!1�A��`"+&P��+����-�Te�>��WD���'���|�I��ڲ�#4$����:.�Aa����9q��osϲ{��M�	��=����7#CV`��<�$�}��z�F�[�:m#��(XO���Cq����至~��&�yw5By�N���Ր�p���	�B��e�54
�#C�6j����ތ�_�O�7����p7�Y��)t�	�T�\�.[���w�V��Y�٤%��2�TC�gk��B�_��)���M��zB\x�+��[# �4�vm=��F\��W(��)��$R���+:g'�v<rLLw��YTu������$k�ϐ��3N����A��a�,�L�^�2�7�{c:|&᪜��3mЦz:�������D^ͻ|y��׫�H\�>�b��a�m12)�*�����#4�\y���
MD2�N��wC�ڤi4��>��oR�'��/�1�Ĭ�QD�XE7��]?�.���||��
��6CZ��/�Ns�ʷ�bV�jn-��ʋ	�*E���l���N����A<�-��4|���~%�������k�o��,:��P��G9QB}�Au�Q骦)�#s��Z�@|����;@���U�W�s�+�%Ʉ���v�b�n���V�r�L�, I}kX�G�Ԩ����T@��1��h,=���0`�k��(���&�t���ԏ1}�{���� �#���E�@®�'��5$!�̸�fd��ȭ��'�A$��Ɍw��C�U1R��[�yi���_����t���K���קxL���S�n$����r[�T�
��͚ź�����?˛��0p/	b��fdP���W&�$��͝����<�W	��y��VV`l��_���~��?	@�B <w����6�O�=\�i;�Y�!�.!<	 '}<x�5A�,G�|*��s��Bؓ*��'�!��0@Yx��;$@F�7	"������㎬͌����Np�$Q�Yv�Ni��@K&�hz�`l����ݫ�tYA�V/lV�0��w�`;�����}>ݞ��3nف��S�i�Mw �A�0�`E��IB��=����(��+�d��K�˔��pch7�h��(�zg����~$c{Y�#�,k�s
SMO7[���z-ZD�O����U)���($H��A������q���/�j���g�	�M\���2��yR��c"�Ċ3��I/7T~k�5i��0զ�����U��*�z����1����TO�@7���j�QD{���=�Gq��EQ�R�0��C&k�1�S>N$M��n`֣� ���GK� P:I+�����pPYk7<'�?��3(yz4�Jl W���t�R�<����I jϠ�������J�xA�NX�n�k?ݠ{�ɏ쒓�w�#A�RB���l� \���[gP����4�*��q�x���ⳁ�LD��娝�j0k�֛7�RM�;׳����Cym伯�؅�~�9Sʃ�W��k�&	�C�iZC͏���ǊJT�a0�ݦ2���X#3�U����J&��j_j�֎>���I#'���g�m38+�$_���b
V{�!'#k:����\��������\ul���H���,tI�Gl��� ӏ��|>^uw`-��q�g�[�@C~J`��$h<�(K:���a���z�hv9i�J�UH��p�g�ݛ"R�駽�
����\x�%Lv��ت��!��T�i�9�|k�n�=���Q��F:g�i��)F�
f�/O��3}`b���G�^�$�U'��>�����5T�<�_����RM{��&����'3��\ɚ2����c�k��ʌ�n�*���)�7\J��]�'g���N�F�L�:���b�bJI#�]`����ei�����*{s��5i������^U�Q��]Ǝ����L��C�sC��{^"�s���I��.�Iך�&��Z�B�i�1o��v�9�8!ZS���0�m��]*�C�,�SWVD:d,����j�M}��[yg�����ۑz�چ�^�Q�Ziԝ�|�~2o�}A)F�q��,��wv+#ߙ�����5��c�Q�?����^m;�x z����5�ڄ�d�#��?�E�����G����Ԯ�Q�&�������f�~�����{1�ߣ1g�y��5�U�:]d���
^�z��J����ҋ;!��L�����Yd�]�Q{z��WOH�M�����(��Ab�G������Ȇ
�1�OZNkd(��k�,mnI�ۈ�-���4Tv�*<����7��(Bh	J�wv�n�C�N�/�km�"} Og���2�d�&�&/&P�f�x�ȷ�Z��[�����]4�f9;�Y��-lZ%g�T6l���Z����e3�����w�Y1k��gB��+�zd��
g�3׸{�)�c��_my	i�6����$��O�n�\�{BYNN�gV/qB WO}����]���*p�vF��%����x�h�^檈l�j˧:���:�*X��OK�y����>�3�Il?��-�	9��sB��:���ݛld�o�&��|p�8�>�� �0�@�t��$�j��NMQ���N���Sif9���1σy�����j��8F[�v��c�fԮ���o���)
�����IԜ)x ���\ç�!��4r�6+Nǈ����rٰYC�MIק���l�qq\K�gH\�i���Ձt�[p5�5Z��/W��^}��*M�g���"X0j�%a��������ku+Jx���l���{�=oH��
clH_u�ڒ6R�gĉ��L�g~	Ϧ���Չ*x�;�W#��Y��+��w�U���յ��ā�E� �����)���v�?���e'�:�r.T�qg����������������^e+��肰{6�6�TrhfGXRl�ָ�,;j�؜qn>Y�
��_�Ls5]�h
hhH�8v5EQ�W-w*�Q���B:L\�upo �ە��.�hE?)QS�k�`�t9�PU�� �����.�o�� <�:'��x��Ⱥ�6]��V���i��2�+���9q��UKP�v�2���L�����y#�q�%��0;)�ֽ���q�#��@�yD�|e8���3(+n�4����{ab�ל��.��`��Q�~�tK���d�;�5��B�.�ʉ���S�o��Uė�]	+�H8���~���!,1J.�*�8�)�N0;$��_u{���S�$�X�uc$ߣ�Z�`$�^�8�4�>c�
d��ʶ/tr�C�pec�#^	��s$��v熤�b��d(�{��>�kd�G�`�{Ǒ���\ҏ��ߨ�$O��I5��i�>��d���
5&���G��,���e��8�	P�a^W�J�
�*.���R��pa��8фo��yb�}���**��̢�_�U`��7J|�Q[*��*DX�w o��}9ҽMhʀ��F�������ǘ�	��xY�	���XO���b���o���3!)
�=@�Ƕ\T3H�Sw���P��@��\���)(HY�Ĕ#!�
h�4\��	��Ǎ��� ~��>%���u��~��EGC���7V�w` �@%�����Y����Ơ	w��_n��'�ei��S�!"N
y�	����+��JAiMS)-���"H߅�X����I���9f�*Cr��N��%<��^�/^:сh�#8��s�ѤU�h�?]8�Ʀ�����f�����X5?���A)iI���Z��A�&r��$.k]"4�;iX-����Z0���c��Di#�q3Q�e�@�e�����;�<���wdc�ƙ\P�߽�F"�j�L��;���#����!Y5�v��@�^�����h�� �e��i����R4�^�n�3���¦̇\�:3yfb������zL�U���se��2�-Ϧ1�z6�<�<5�@ں��	�₎ۑێz&(������a��!����g��+0�����h�5|���qU��O�Ϫ�o��E�k�� ���h�trF ��cĘH�cgV�e;��'�=��tU/(I�U���F��/����1@^Gy��OO�X*cB��'U�vqTd-L�gK����᫇���e����ݐ.@��c/��ɝ;�������%K�s%�rs��v?�%k��?�1
�'"��P�G͌]ʚ���O������~v��h٦ό�h:ב)�zG�Aw��	�=�+ؑ�Ο�ϫE4b��X�[v�i�L3%b�������ӏHMsYL�g�6[YY^!�����Y���|���d��.n'J���w�5��t=\��8+�R%M����}&f�<�L��=}�qMz��#m�4�W�bX����
$�/��G�/o�ь��:��2A�u{��19��K�>��U��\��<���3V0�l����0��9�!��Zk�{�`�3�<N⑺����H�� K�`�&�2�ꢁ�&���x��(9}����}��}_>�m��=k����H�N��yV`>ӌ�D?{���H��2�� ��1��~9�$�t�FU��m�s�15�+�A�O}���F�������w�oJ�2�!���k��i]���3�ø�I��Ԁ��ٕDK.V�X���^M��#wˏ�bߥ�54�?�^�"p|ًޛ�7�"[xyM���������懺�%��=��X��zU7rE��U��
�I��A�p� 53����3�e$����I��5d6lh5�3��ʀ�J"p]�cAfA2�~%����(��?!�(��Ua�p/Z�}�||ǭ����Y���w�,A㲰����<���1C��m�d����� K3��v����Df��X��ɾ�Y8�F��J�P�����Ae�r�����
�yA�;���9�����p�п&��*�����N��+��C��S�H�2�z	9���/��F�rN�cwy�~��wB-���	�u������ݍ<m���{��K�0J��A5T_��vnC����hmc�^%]p��-,�uإ�v�o�'5�dPd*G�8w[+g&�3��2���g��|
ԣ��3}�ۻhΕ�ho��+9�4���oBqo�aj:�՜�0o_��	M��xB8X����}�rӅ�sD��,��r�I���r���`
��Lք	�9���duٙ��`�v!��~�X6��-
���4��}� �F�	3�DvN�MJ�����<��b�ΓV�;�ِ��������%Ǯ^��Ğ�t�:���<,xG�6�Ġ<�!%�X�-�f�j����J��^}�������@60�#@���&4�B䉫AgQ��%P{�o�e�f��x���5��[})Ȧ�����W)g��	�tq):�S��,��{d�竈��6�ya�\��Qem�h3���i�72UG$̖�cT6bv�����}�p�KD����ć�,rhx�ְ_�����v���l��Q6�}˷Q��L�'t3�"+d`6�k�B����]o����ӔD�l�\��^�i�>�ޖ��Z@i���&N�����R�mv���@M�£Q�ش��uX�ap8,�(�}�"����̘����#I��0����P�����2���6Zi&8C�C�=%1=J�6Ͱe�0;���ݫ4vΒ�n�H��;k��oh��K�7�����9�d|���@��	��$V��^��M��X�W#{jR_�.�X�Z���6l6�;���� �jv}���0[�>����
���mrW3d#�;��!�Ɗ�P-�n�]]n�ݧ��YD��1�v��~D�	z9�����?��BoCG�[�G�mB̾߅_��u4��v��m"6�yq3�Xj���'�{�}���� =&aXG�Ę<:a~&�@uP����X5�"�����弴u�q�̡g%s"��Sە ���#��_<����G�-�� Y�0�6^�W�I�Ա�!.%�@1 �'�9��e���K�������f�{:�o�&�E=�����U�|�a����t���@A��A�a�B;EH�|��$-���L_Fk��|97<��LO	������?O��n���M���o*�OC��؅�&ܝ����X��_ܾ;F���e� ���)�YZ�M�,�9��oK]������3t�3Ȏ��P^K�ԣFȂ:MYn�p��,'�$�����3�D4�P���!Ml�P�E5�\{�@�
�^���&������1 	��*������r�BKh��C�����J��g�v��������v��]u�*��%�7���0��}�S��9��趎�j������7��I��(���9��F8rdJd����/�U�s&��JT���svc����L,��k�`�_�oJ�s�����}D'@C�>x�oc>��Kx"�z�6�N�����W�g���C�bI꜡+l��H�Q�����,w������Eyay�0����*\��K��������ZMJr|�6�u�8ᅵ�ғ��>M���b5e�,z�@���8x��)~d�~���
�5:��g����\�J�qnDf�hd������b����E���W��Dh"�|Rq%7�� KņZ.Gɼg��|��Y����Ľ��ݳ`>��/��	���M����k
�ĭ�ȄAv��>�Vnfu�l����,��c_��^w(_H����\sͪ؀�}�LOF���|Z*�D�T=H�mA[�
1A�0s�Y�8�fes�[k�M�Z�$Z�Sߊ�o2qbۖ;EMQRr.K@@*������A�p|�U˜jЪP�7BJ/�~~"�<E氃bt�t8
�3>G*j
'���V <!�.���,���'�(�:�`���� `ͧ���D��2�+��CoI��ٗU���9+W�*�>ô�\��}I��D>����u��J�C��Y��1Ab���L5��8�3����� )�R���B��9�_��/?�wTl�� �Zr�R���A��v=��C�5��2�5B�+A3��u&��,�_Q
z���N>aJ�h�����������S�Ӗ�EXoV��/���,PۑORh�*:> �]�Rҧ��tڛ�� P�1W�,^�?����q~�>g �|Q�/��p�k=��G)�`7��wJΡ��<����,�Bk��N����b,PX��C�W*T��7� ��]J\f#�Md �,�+��F�4�I�?����r 	 �>����Ruà�'F��g�mf���q6�Rw�&�H�(�!Pm"�c���p`D�g!����0�cat҃�r�D�z�%���.��&���ќc�~��{��9�(�CAE[��#X[��)�b���p�D�C�G���PD�r�{���Q.���D����O�G�f�^z�H�3M�#�*8�ޚ����%>y��rwj��2�FW� ��R��S�5�ډ�9-���=���\2y]���&o/m\2��a��Gn�X.V��,�����s�ӓ�C�^���t�1����M��G1»*3#�~��Cw;¡׊������I�Z�/�^Y�E���K�4"�o�
o}*�QWK��(�򹚺Hc�9B�Y��L�	�fA��>�*|�G�c����w�+eXg�m8�ٛE�
��╫����t{Q"b9(��A[n6���]�����-�t����# �]���yN��殑�,����)�;�,uh��a������G��3x)�*�\	7r�;��oh۩���}����jm��L�E�=�M�Uoظxk�$�c{	�����!���m�8�RN6��D65u�Q�������K��v��'`.��엃'�6�]3w��<OS�-��;�֝��L�X@�ѧ�:�-��<�w(����`Fl��"���z��ӝˈ���dF�x�pM�E�\"bp`��;�xoe��ރ 3|�Zǃ�a�H�[��O��[�j��Y�|>'a�7��V?6ݾ�/�g�;�^l�>�����p�=�4�rҢ�-D�1��_N#nTr�2*;���,��$4�]�`�i�^Pa�A��"L�a���?j�w���IR�Q��rE�a�,�A'��f��:eU G�4�nIv� h�?e��|�������5KA��r���˻0�����a�U��#ؼBM���	�18S��e������Z9|k��^!��w����8r�Ty��i:!Q*��>����!�p�I9S	��t�xv�ݩ2�fnh_�������Xu3�i�(��u ��̽4��D�z�<������ņOa�d�n/��J�$�G��]u������8���-��Vg�!���h�]��.��� ��doW������R�h`1h<�C�M�
�I�6� ~�ᶆ�߃�4%�I4�� ����������YUs�M���L&�#:;�j�̘�"�g�Yur��D��l�֕���*v����Z��.u��ksI�8[��ג�9ϭ���u_������K��l�0S�{��!І�Js���/t��<L�_�]8
xI)�����O�D`�&�Sc�y+ͷbPsO�z袺����C���ۚ���l��$>�Yכ��'��|�u�����N_�S�d�����Т����	Q�:c��X�+�,�S+%�K���F�8S�<�Oמ�<ܤ�YOGtǶ z\y���3��4m��^�b-V��"s#�jxj�C��'�m���$�1�T��XJו��{d|24��� �/�����n$��v"��7�{4�fanZ\��Q�,��4�5,hAD�1�C�|�~�l���+��W��x��:;�ot~ԃv����wo�]C�H�h�a��C��SM-��������g�c������X��;���B�g��f������<V�ؚ���U��@��8��A����
fB��ihE�#����ň<�����I �;�ڨ�j�OS*�o�]�ZR9V�ܙ(E��iX�!�#s��?vw�m`�?LpI�m���B��^�A"mQ�.��h�:Ϳ*o�6:�ܴ��y�,�x���'��5KD�d��"1�o�s��;[C0�s��k6B!NgBB�����JS�T�~Ϟ��@̯�O�6�[�IE��BO��z`��z�}Rv�ز���Qy���?N���O@�q��:��n��|��?�M�)�^"_��� �P���7$x�ÕV�]��g��@(E�p3�t��˩ψ�	�����o �u��X����>8� 2W��9�j�4v�2��޸�W%>$��E��&i [1N�~�5|��]��^�m�c������T(16��8�r�񪹾D6i��P�?���R�ZZ1F]*%�D"�e-þF8���I�p����a:J�����H�Mxƚ��s���4l+S��k!%�أD��7@�u�,�e�2$�01�IJ%���r���Ͳw����#�u] �n��S=i�'!M�ڮh�ڏ�uIu�p�uyHI��:���i�k�hV�Սv��-���c޻i����n�JBI-�7˓���婚l7x��he�@�:F���(�X�hɐA�͞{M���V�դ��#XS�����v6�כ���;�����G�C5���&r̀�S2�����z�w��6�N'�
_� ���Ҁ�#������&Z-1?nLy���f�/9;����Q��'&fe�� ��{��q��)�s�T�K�磁f#�5_d��y������1Տ&�P��_E�Cʤ�3������
N��(���ָp��t�j~-���p��( �ϫ�
:��$~�+zvbI��l� Vj�'fc�;���¥Uԝ�]S�Y�����n���rvʪ�����R�b�	�!V��uf��]����4��'4f2�q���l����=�h��pc=R���U#�*ܼ����A�
���Fb{[���JVF��7�\b(g�13��H rv`�C�$U��=kCHm@�}�`B?�v\��t{��4�7������P�H�K(��Z��ݜ�}����&%�x�g+B��(4W�P�it9mphB?�K���y��w�y�K�!���ZnP�a���U�s ��:Ҿ�u�>6D�H 5�T*��*�!�����˙�l��Rk�N%L�2wi(~��G����	�y�e���X��T��Q�&IQ���չ4����[?>/���W~D��:w�)�Q����J'_R��3�H���bq �N�9�p�����B�5��/���-#��b��Ǚ ��V6�V�-��L�G=�!�`�E_��&�UP{�!�be��I{�����@Uf�\�O<��ے��7�>���ME֘��a+� ��u�#�ID� N)��n/z=@4��n�ť�8��>Ps!+����;�u�׎�S���0#��,cgEۡ�z��3ޫ��i>w�?6�Z_*C�����
N��};��;���u憂}�������=�r���2�h K!�N�ֺUr�2?�]N���Ɋ�SA���`�/+��3pl�[G�^ cF۔l���F=�|.�5��|�2���,"����A��](C���OɠÀY��,�4~���M���P&0+r^��ɳ��������B�2��l�U45ų�ͷ�u0��n>���k)�1U�Tc%����`� XL���v�t��Y����:�>�z�!<�<�(��W�e��	V��G�����P��#G�p�rrV�lT�6�o7H:ŐY����`�s�&f��77Pv�b��� <Q����6$ƛ-�l����� �P*���qL_�ʌz=b����� T9ak5����������d'5��4*��f���Ň�ש
��$��縜K^2� �; �:���\YE�/`�����O>,l�����Nƪh\pS��f�z����Ɲ��T\�ҋҵgӏeJ�7�� q��v
�?��xM�Z�r7)0,�h7�;��ȑ��qv��V�(ԋF�"3Qf��Vt�A��Db�)�y�{T!�T�6�l�I��
h>�4�?�1���<T�O��ל��y*�}*z�����G]�?�.�BX0Jx������s8���$�,��LD� ��ɌD}X���@v�L�U0xl�b��+
0l�yT���2c����P��ġ��(����_��o.G��5n���F���@D����fz]�O+���x��uZ�l���o�1/��?%���%}:�J����Q��]��l���R!�xv8�f5���CR�&�Ij {�<���?�x�8���Z�!��ftF�$.�=���w���]ce1.��v��W�x�q'��>� :W'�
hD�|�;�SB���T��X;NNi�6��[�F�8��D���bFͯf~��:
�)�W�%����5�:��^���WK�"@T���qh:���|��*���%	߬�ꂾ
>z��\�BG�U{���i��M���3d	���B��3���s���D�����1�Ʉ�ƪx�b�2��v��F�=��*���TϾ�^�i�9*�3��[2!�J�^K)�/�����+;C$����]�
p�4�z�W?P���i�|�h��YZQ���>���P�/�H�@{�_��}�L��!�8�� 徼�KE/9(�ͶǾ������g��8�dM����+�jQ!���>CH����b�+>r��;�7��C.Iݚ}X)9>�����/5������A{�~}�R�����+��n�I��JZ۳P0Nh\�%�L�Gay�BC�0��8�K�.�������S%��hYGk~t�nIWY���6��Q������
K,\�&,D��[����������M�����6�횻{�@``�-������]���H�+��e{�S�#���.�!`1��:�"w��F?К���4.8b ke	���i[�(r%�sf���}5FKj� �#�����>i��R&�P&?���;�Y�
���0sB�vc���m��u���)ym����	Ӈ��E<���S�-0q1����^�j�-q��Ҁ�,�����f�&���=,�Sd2��ؓP�癒�h��3�\��ޓ�Ft��~X��)ʴ!4H����zg>VF�$c:-�8si�7n W'�Q6��jn���on���_��d�����
�x5�Z���J{)�>��g�~U��' 5��A}Y���J:�U���=0&cj˃��l��O�P'*úM����p����v: �0����$�J�?�^o��K���hpj��|����|܆N�%Ċ��A��A�u��kqN�{_�ZP��{�A���'Z��0VW��b�O�Nݲi��ǩQg�iVGV�(�\�?d�����kY��c ����J�G{���o�1	͑��r�P�!A����y�J�g�d�ʏ8{�
�
Wkԋ���gB."&$�ag�=S�����f1�����䌉5�@٩cA��)���>�L+*K�n��3��'9��ךh����E���+��a
��c��4��hJ� ��S�L���뚂���\�0�w:Ex�SD�`�����Bh:�>#3�}��0�
�履!M��f���w�tj�������>*}�'zId�t`�	)^D�F�y���������=#����`��D�N��:�]#i+��D\a���S���l��3��u�A�O���܀
՝�+R{�ܸ��/M� U �!n �E�g�&ǽ�g�|/�:��f��<ܽNE$�03ʔ5M�k�O9���U�������R:O_D.��r����zQk}ًR��>`��hLRMBM�m|
�G�`�1햔�!�3��b�`����E���C�./�	ro��Q����'h�x��俴�kcAER�+ Df|6X�'�o	~�B4V\�ݒj�1_�B���p?�|�a��넒D[���H.�n�Z���P&�E��V��1��\�Վ��@dE6Ec^�TΤaEP/ƽ���Qrx�p��%���E�)��?�M��C����O�!U�˘�g�@'���@�b�8�G��V3�4Fi�N�0M���et�����A�}A�[�s.U�_�&Ǯ/��9IcM���_�N�钫sx޶�l�� )2AZܯ���;	*�b�dZ�������3�^�7s��e��ݚ�zEyi	��unJ�`�S�9yK��@�~��C��Mm�4�,m<�͛��ޣ8���UՍ�t�+��GZ�9����X����m~]'����n���� v�"��v����&4��wLf�7?�0S�(L�3����F�T�|��QmQB�_��x-�	�Ӵȏ�})*�r�sOtC��mIZ�+��!qj���f�7^M��x$z����k��,�`2���A�<�~r���:����G������v-�Xt<r׎�O-�<�w9A�*���`�bJ�Y���C������(�r���(Gt�yа�����I@�Ð^#(E���@w�ٳ�{�N��a����s��T�f�G���)�L��Kk�%�TS�^���j��C���QŪ�v#�ƛ�{<���v�X?���5w��{�hƢv/�tٴ����0�k�Bג��EV܍^�������?��S���گ|�r�������:\32%k�����$ �	j��Σ�?)v*�qD<_ѴJ�5�w�>5��)��g������a���*$��g=��5-<�uR	��%���(;�lp}�cי�{՚��J�~�E
�Bw�P�&��W�!jw��Z���°ɷ{c00�R��}�c=����+�RX���f�(�%s�P:dQ?�K+%ip���6$#��0����D���]��~D�5��UP�6d�`tl/<f�rR���8�	yM��Xc'?�糁n�6e�ݟ(���H�M���7 �W��4��r���FQ�����#�š�)f���"W������m�Mg�B�U�#Ig���%i���f�W~����}����X�>�9���7��Y�]���Q�5���1��Xcն�ʘQH��_UX.x,��\��/
W�� ��ݖ�?T)����5j̭�O�[�i$O-=�k��LA�Z�����:�H�Ed���E���l��H7�� f��!4���ŧ��Z���2�G2Q��y�ȱGs�s�Hyj/�5v�B����n
c�a0��(|M���~��?��	�,�X�cb��id7�����/�ԅ�c�O[Y;��BM���31�c��n+���BtՏ�6���A���g�Szg���p�f�#���QtJ��b��#_}�1�Jnk�/��lS��?KH��-bBYpŀ��ar�-U��R�ʗZ��0xV��LI����N~�Z?���$���$��̩(�Slq��Nq{2j���*�� ����eC�����aSxc�{�V �4�(B4�P�_n�_��:^\���s7<�Ja�,�9q;�Z_�AC2c@E|���D�,LI��L�6�9�!�bay����,W���z�����Y.�S�Ɲ��BX-e��_�a�E������A�LA����ʇhx�g�ߦ�������+h_�^-�%�{�ɶ���蠹P���Z��z/ ֠�����PQt_��j��ȵT�j3:9	�QFjw�W�bZ������rh�D�A�S��PԸ���O7�M=v�ă��v]9֧���g�v^s@�����X���V6�j�ۚiJ���EY����T5L�#�.P�ZLm2R��%"~�B�+2�%:1�,�
z��t4v~_ݫsI2�-Be�t���|_�?I(<t��j+ѽ ��D��ʤ"���}��]��Ev�儒0ѧ����3e����(�HZr��������35�9�-ep��5��Lt�o����,��#�P��8��\c��8K%s��hn�yxe=�f��`��?�u�c��(Լ����[%����p��N��T�F�=���i���ΰ�f��z������}��W\�!�����W��"]|;�!�R[�fH���R���@�S��n| �"~G��8'�y�^QdQ^_�`��ok��#)BJ>kh�?���Q&�?�� �=��SS���AFCO���*��4$���?7��q�;+�|���ey�����l�sNz�����&u�<n���Mպ���J�D ,ߍ��1,z�z�}����̇p/�%zxN�������\rk�I���hK�}�'���{���f9�.l�8�^Ԅ�n�s3y���y�>� rb��ֳ�7U�Bҽ�&��#b�<_�f�<��S�v'�ҳ��pz�e�c�Jtw�B�c��-����Z�ZӸ�Wł��E�	!�hZ�81mͼ��4%#�h�z���Dځ����&$��4��k~!����������_6�.3Ɣ�b���	a��B�W/���x{���E8�+���\���Gт|�h���a�������.^Ri�{�B,It�\@f��0}'nK'F���m���S~�KeޫG�h�s�F��?�d�dq�w���T3���"��%�?U�k��>���s�@z�Ύ����f�.%S�����*Bxo׉y��S��{J)�X��I��|�f�$����ʻ���#�U5�>�SyK������mv�P�/���Fuh��2C{�J7���t�(1���!��2�t������@,E�m�4L�Os.]��]<�Q$�&�6�������@�C���	U(�/s�-�h��07-ʪ����gX���bW�[R�Y�]�A��;:3B���	SN��ƴ�'���%�&�4�:Q��L3��/^�@�o���;�-g�R{�{�����_�CK'�׳fuC5	����T��7>?Ֆ��3d��<b
��
u��h�@3a�����]�p1o�Zg�X��}N�]x��J"�ײ�k�Q��Qٱ�6�,��D�c�-F�r�����g���; в:B�\4����8�I+e�zB�/i1�CS��an�g	� ��V�SU�(���g��NDC��o� r[�1>9�CxC�{�:+���`r�] �m
���O�?�~�/�<�,Jm_'X��H��twH�(<��y#�X��r��O0rX�x��(�'�5��:�?����&����8ik/R�')5�h�,/ғ��o^������(B��8_�0	��"\���#^��e�C>���升�p���*�0@�!��y
��,�����d�_6���Q��t���>(��Sc�D$�`�&�䑷�j�� yS�G��>$o��A�@-�*����y��%��4�,��v�*ZЎ��2��[3���C$c�ćN��HMt��̮��C�m��#�@�acx[o��qS�I�N4��I�q��1���|�\���fZ5�[�@r�B��e�u��d� u;�����p�aʸ`�������ʬ��Q�|��t�!'[�6t��"S�MU�M��w�G�A��O����O�-w���}%�{�$iXEU����R�d:��m���+�@����H��.w�l�%���#t�2�l�n��O�n Y85W����b��T�l�Ҹ��:j]��N?�S��S:��A(Up�t��y@��`{n�o����k�E�[lUx�c����_���Q���PJ\!G�����O�.dk���Ql��z�,.d��~�qz��$���OЧja���Dѻ��GS4u��Ŕ�����M�;���un/��}�2F����JH�Q���վ�����lʠV��w�P�Ҍe4�R9L}&+yN����E���z5l��fC>�ArK]UC�&9ґB��RW��Nנ'�5��h���`�����vNڿγR�XBG�q�j�"���^�_��� JL{�l�W=�e\Ѱ��2y����+�1"ۜ&���i�=/I�G�� �9����<�S�$�J�� �j@�ɴ!��d�j8��F@�V���g�l���ܶ�aD�[nX�$|{�=f�m�e�Y�D�t�a��~jW z0��ju1�Ah���<g�*��8&�����������Z�M��q7���o*켊&*�X�����Sv��"�g�A�P�Ru�r-�s�nir�]1�S�T�w��A�������@��=�Do��ޠBF�N##���Ϟ�����*y�ԇD�,,x7o�����ש��!Ȑ��'���}��b�t�{���>���v���Tm"۰g$�m)`� ��8վ@T�]�+!�
rb���X��+�'<��_�Ĉ� ֌|�����diڵ���w꼪)�Z���|�se��*��Ffx���I�8"&� �yg��eϺ��w_4�\\E�Q�����E<��
Y��@̂�<��d����vIwC��0�nѰ$!�%�RH�R͏��jsJ�K��x5jK����=�-��$oC�ȠGv��%�{.u�+�0�a�,R����!<y�.�Y�ߣ��P����=szd,Pk���3��<ݶ��9]�a��N��<c���<�%tw�(�;����⺻�1��0:y��^xI����)��Y�A�u���yK��=K�7�:�Vx�7�����"
-����F�@/��o��]�6���!���������{���?�����5�����Ni�S�Ȼ�QHƟ��μ�Z�{����N3O#��9�5I9��{ڋ����"�X=&��\_�}gWGlށ{_�Z�H��I�o}��f�<Z�ݓ�(�y�~}���Ѕ3��D���*@ҰN)� � ���m;����d\%�Ϫ�4$w�X�ϑ#K02�����i�B�5}|�����Z�"��X�}.��Q���0e��������(�Nb�k�L���PG��OXC���W�x���n���ǿD`����$�IA�<_��j~���ވ5�	������ɨl>�1�ȵ�s:�4������d�����X�P= P�1V@("��/�A;�B,D�/�P%"Lڳ����o�&�BI䔘��h"�I��[Br�8
�����J~�0+��"o��2;vÖOd=��D�j%�6�؅�XKz�����ڪd-�0B6a����b�97��w���d}�m��������m�c�jNN�w(�L��l|�{ �I�9:x��4��P���21�r�p�j�.)+�qm�*��&�{(\��u�1��g��u��Ǔf?�[G��z���N�:�C��m_�*n�&"��oo�|�|H��J
��V����<��Ad��E��a&B�l�	/�(4��<'"�������1�w�a��<{F�Inȣ$L�L8\�精@��_�����s+�r؃�,��-o�A�I���iF_p��`�=�1�v�o�1����,�|<SV�-dcM>�g^���]r��xͽ�%��������;�����7xB�ev��ݟ@ޅ�2?#�gi����W{�c���ܝ=���S[���fz���6���ҫ�
:G����O�ֹ��c������k�/����	/մ"��<�(���+W�| �1|���Z�:�ߪQ��%�P���V#6��_5���'L���H���^1sJ���j����~� �x����|�^;i��H�@�,�nq�z��G���cƻ�|��Badk�kwI��ҳ�����,��߼��H&��V�������K+}a Ee��G]1��d�-�p�$}�$Vo��'`�6�k�V��<]r�|�1��d`�c8��:�^���B��>�/$"y��A���n����F�^y��ah�A!��;2AA��`�M�HG&)?�����̣^oò]c�S��T�霜��H�ƶ����Tru�^�a=Q��8ӧu�#�j�WU�� h�
��W���㎇�Q4]�μ�nU��ґ���~���":Kpfͬ���H�o���o.�b����JE���7C�@��I���<^2f}��t�n�-5Q	$�C�rTu��'�Ϻ��Uč��m$o�u�����70x�R��|�yA�J7�{�L� �͕�|�^E�����ƬzB�)�N �~Mw�SK�	)a��gI[�n.�gY�{}x k �s֝�Lm�(��7J���ڣ�?B����A�v4��q��q6��z��PR�)VP}>
�gݦQ�O�c����z���� ����W�v9� �ArC11�`���/�g(�\��f�C�}M@��z'A6v3�&��4j��~��Y�}b���p��� @���&�l�;t� ���u�*De}��c�~G`(��.�Ĵ���2i�)j-�"��Co��G'�U����L�s	��c2��TO,ע�u�Yhu�K�"�Z�x&r�ۺ����P��e�'f(����IjX7����ĉ�_{Ε����
�#�Zm�In�l)roA��.�߸}(�{�n{�TMp�k��� -3x�(���B�g�5 �p��)�F�ΏX��MPO�R�1�%��!lJr�2 ph�k@�"6pn�+��5�d�GD%��Ȕ�-*j3���(:��L�^X���ɘ536��w�׏M4�5�)�̈#�%-���M��V��m��ɦ����SX�"�������6�]���w���!����v|���Mq1�h�A�{�����<�#�/���� )?c��[�rc,���G��c��Ƨ���7�A��ۮ�{ֵ/�5&q��Pp�����f��}NW,PJ]�2�.Z���n�w�cj�8�	5�p��w���	7鵺!������I�\��f��B�x�*�Ӧ�;�L����� ��+��nג+��r�Q�k!1��.ks^|	�O��y�Ƈ��!�46&�k�<Yڅ%�u��~�z��	�ww����k;��Ah�?����4��L����֛o��唦��~%���R?�?�F3#�2ɴD�5`ž����N�,�qx�<Pk���j�3k�����h*� �K^ϺD�~m�R[Q��N�SF�>q$}���`Y��q%�H��.��]Â0d'�g�>@�d���zb7=^�~�s�0�D�E�ЁC�Uӊ�WxbHt�t��hf��d��'@�ق�#��*���J�	@7dZ������ ��t���Q�9��=�V���Uޗ
�Mu�"��~8��+�h�������j���gi�?N��۸;Rv��]��j�]���f^�+慻��]MN���n�q����%(^��1	6
fLWL�7�����o*S!s6����zU���@"{׊^��'��P��I�Z�D\r�O�)�k�$�/��(�ߵ���}���s�kZ��QfF��b���B�k�b1Q����,��O�\����k0�;y�tK��2���IqG�j��T��u�n�3{���0��B��Oa�M?�H��ô��c(�������2�0.���m��͍�Z\}u�t_�]��(�����Na�<�<m-e��w��	AO�I�/��4�^���~�*��D>`��R�������,�AT9U��%0֓�x֦��p'
���5�����rOY.��滰Z<����{����_KC�W!�@�J��5�w��^��~��[�{��m�x=���e��4JX��5��\����ˉV�
2i.�,{���ƫ砥���hդ���O��`F�>�;�]�y����*;>������R��]�e�`?��F+5�՜��4�=]r72?dI@	o��[���1��wL��_>ٛd�o#W���xVVJ�=sGa�K��`�Q�$���%��^ `��8�l�G݅D��d��y~�Xf
��
N`�K��d���>��$�Ϋ��pζ}�)�{zYҏ�#�!k��bVv�v ��\����}�,���:� ��Gn5-�]T'�"��mҼg�ꋒ��,��d}�P@�ܠgRݯ��֜K@��ܕ4;1��t��u�b�P��=��	����AC>��~7��pg� �S��|W]kh����_%���\51d�k��o�,Q�7Ӯ�+�����7S-4�Q֯���=�<�Ԡ����Y{���!����FY��z2�*�>��]��rP�D耷a�" 5���ԛ��#ב�O<� ��щ�h�#.�CI֨�����$Yhahn��	E��~�:WA(�t�#v�݁6k���䨭���r[r�_���xQ�fC���H {?#L6�{vkfOS>�����<b���7^�w��	�1}�k%��\��$���G#�Y?`�7\�*�F�&�^�~a�ϳ��=�$�Md9,=h��w�J[����4��F�D��n�"F�>���`�=�T��gl+-�g�|^�H���孁�N��e|�b��F�5~���q�f����U���œ�}�V�{\E��Ԣ��D~���*%���[�ާ��Y�'jdC�����a�ZӮr��S�X�x#����v���^�����%�����*��� �8��S�E����A�T��r��fs�r�~���(����DA�G��5q�茝�n�ʬz�9"o�����R�
���T�0:��xYC�=�x�o��H��1�$�gY�?)��3)K���'?��zʢV�	��N �0bЮ��=�1���V����U-	��Yvx�ɹ*��J�p��z������,L;L�� sfs�ԝ����xݯ�\Ξ��q��pE詒S�t�N�=� 9h� ���Iʓ�Tc :�B�y'6�{9Ň��$�fW�	gA�l�I�w?oZ��{�c�)�Z���7ȧհ�J�!?���t:�7���~���4'�����C_���]�jw�+�T!H1�/�,��b[o
N.�Ǝw1�]"����L���FF�u0"��Fu��AR$�t��#����n�t�T����B���5#_�Ie���ϫTHN]ei.�=�cF��	�yJ�JNF��c޹��똈Zms�Y>)r��z����R(9��r����I�6����P�V�#���d� YU�����$ �P�4 �&�w�ۯ5~�Ak h1���f��G�/��w;<=�ab(l7I~	Y$������C���'U��[H�I����
U��8!k�C��ah�`S#���1e�(�ctA�
�>�j���M�7&�	����u �ՙ���>ܕ�ζ rZ�=�^��Dڰ�����)7�:*s��W���"e��#׈��^����#2�_^��`-�?�r~iW��>�_�o	����i��xw�#_�`�ґ�6���(�}���2�/D����B����������F:�"�}ڢ�[���Æ*�c���O�q/��3�xR0���p��������
�ֳ��ޢ�\0ɇ�`��~)f�6Gb�ɹ:u�AHdM&^)]�@$�G�Y�~�.9S�/��U�n$�l�#}�BNfI/��1��o9�f%�|�O��JY���Y4���EǞ�q�/�e3)�m*aR��s<t��e)�����S����<��%���J�B�AG&;^?��4Q� t*��l@�Uh��x8n�F������)�h�W`,j�bB-�M�w�խH5� �l�{R$��'Z ���|籘����#��·e��EW���-��@@�L1
���':y��9�DF8��1(�
�=Ebְ#x3$-�> �eKI ��'�^�UsS�|���k$P�+���hņ2K�LXǕ���̄�7�,�ĭ��Ol�x�����Բ�r�T{G�A{�F��)���#J�;z�-�Fw�KqM����&(Y=oYu$Xk���_�_c�t��].Hσ��
_0n�bpƊ�iO�^�D�a���������Mf{�H�w�|��ê3���q��X�l�6*���(��5�2����6���'9j8��B����pD��<�j��o�d��9{��!�$mz�d<����r��B�o+:_9��b�S|�������L'��[҉��Ա��ҝ�ߌ'f�7����\�!&MeL_8��x������3�H�Y]��h��c���'~V����M;
�G���o���]��:�����^�rEW�Rc~7E���'!4Z�c�ӧ;D�Jv(�s�/�d��%�(9�ӈ����dl:����:`&��<>8EQ�4'-*��X�!~;�i@j��YJT�_�ic��}�j}���n:=Mu� �q���ĨVBj�(f=����:��h'A�(
�C�b߲��e띹����Ӭ���[0}>�p� �{)j��	D��RV!�>�Q��e�%�gA6��g:d���TERZ��G�[�奎Hb��Mu�����%R��_<ĩXh�}�?�o�E4C���>�\Tq�:�%�>��N6�k�U��X+��3u�m��4D_����"D�ݭL''�5�T�я<���uKs�),�����׀�`ޢ�"#A$ȇ,t���	�)m�m�sY,�"$�;��EI�A�|h$Y��~!ڨ*���loq���c=����h.�I����=~Ru�bm�tH.���k.C�C`�؎�� ��WP��X�dބ�"�r���礪���E4���
|ضk��w.�(˶���$L�/AA`�����I��Z�^R7#�-d�w���-HP��'UߡY^���X�����P
�T,�6f��N�,��p��<� ٮ���ąĖ���FD8F6�.��mpK��n���Cn��z�������1bi:O�\�F3�(���Љu}�B���p�����������3�L�nf�
z��t��SI�p	�����VJ����H��>
E*t�u<����\H�2��� {�O�Vxxg��g�	j�9�D	�K�K��]572��}�����I�Q��4|�]y``Æ6�����R¡���4h;���XJ��@ڛ\-�m%�ӆ�C^!��W��jy�f8��'0!a&���z饘���@�r'�����D�S2k����<b����-�aƕj�z3Ҋ�T�`*!V�ԓ�xN'~*<�I�����З�y&�yX�+
T%��^ܭPœ{)I���uQ�H �}HKz�m�0��κ�sy^���$Ȯ�E�I�ۃ7�/I�t ޳�V|t�e�'VUN}Ǔq]�.�,���Y-~�b��ru�g�FS�^ԥ���b�����ω�6��7���-ً�k>��s=�#r�|Z��:sj8oܙ���	�d0qJ�����⻽�VtR�_�z"��V˲	$��=	��jg�����)���lOF�#Zq���3ނ�H�@�f$�[�����q{f��c7?b��t=!����/<Ł><w�]q
kJ��m���1�6d$�J!�]���@����Ec�\�'�����8�
v/_�pS��2���"_bBEn�X.���I���U��4��%v=�b#'� rHz�Ɗ5�y�`Y�r
�D%2H��):}^f��I��Ļj����%�j��[�f0�OJ��,)4b�a�G�P���_	穔?�2���%Z(�9V_�,���E�fb\�+���6��^}A�����ޡcr$�����;Ƞ�q��P2p�O���03W�[�X�E�#�N�6�~��X�Hp���,YYLq3��J3��ž_�Đ˯jv�#Ηd�uؗ̒nmƂ�f��\G���G#R�J$��!rS�j���~�56mֿ���"lmjF�:A1�	|L�rϯk���m���_!�_��=�g���E�����G�� }�q4TK��Z�|���ʁ-4���Ҧ�S�|F�TD��8z�����l�ɝ�(S��6��fK��UX�CN7	�NTr��0a���ݼ�	�%��#�T{�[�G��Que�=��"��Ž���������>�[9��y��8��uܔ�����=���G�G�ϵr0o���Rk�BL��u�C"�1�]_��=ƐW�j��m���h��]�[BA���D�F����衄I��A�͏����.�^��GE�Ė�w�����s��&�jWp�>�G%���r��)�Å��T\�`fE�I���˛k��#��.D�1�`$��|#��N�w��n�.\D�>K����KĎOl'�~���5쏜�dB�q����{)�ˬ�N���v�q�4�a��h1�R~��S��s�Ԝ�~\W8�|q._z���^��Q�E��ٛAz`�3��$�$Ҕc��m.f�����p�N����"&oկ ���E�cnV2s�z]*�	/�tJyt8N����h+�j��ŔY/&sۜO�ҙ�q�^���g{jIT[�)���c�Qq��������%J������dя��y�1����΄��әI풊jNRSC�[m#07p<_滒[� i�?/��u�(�B���}#�W���-�sͯ6�0�	G�+�ՊoJT�����Ӄ�4Yaݨ�k���I��I�m%������\���TWN����'
7�6k@2]��Qe��$x�M��S%�HK�9��%)e�L��R��jȆ��]�:acՃg&�ه�Ċeƙݠ{4WO�aI#�lq����Y�$�d��6ʂ:�<,���!��&m��< �bfl�~^
K�n�J4 ��dG��Pb��ʇK��9�{>����2��5m*c��2p�/I�}�+�W,� �_kǘ[r�b�%�u�C�(���gV\�8�1��ES`���6!̳�z���j�����U�؆�G�Hl�=?8K��Y���㆙�?&G&m�X/�z�ʿ�f�d.����>�Sz�;�Ҧ�ɽjg�1�>_L/y���ēA� p�.ւ.�*͜1T 	�jfL�L_�ا�ͼ�K^��B��z@����X����.8l.�!)��E���"G��쐐�I֌ c7��ԕ��GB�?�R�]\��=N��ͦ����_�{�9�<=R���߿&W�����ٓ׳�z���G�|ٖ��JO�!q�)\t��S�*�Tzp�U���mKB-x��Ú>g��RF�զ!�G��;]CF�Ω� 뢰�7D���2.H���߮ʆ����a.~�?���d2NC4h��{��b��Ǆ!�����[�-%�����w�,Q�9g���.-="�#g��ף��DJ��ɕ�����Z�vl\�"щ>t�Re��*�%�4�	d+����`��6X-Y*�5��oi�a%i4
�[��wJ�'�i����;�)�`������/o�pm���8|�8X a�S�| q��z��%.���y��ô�U.�0,�79�2^�:L��ص0]�U�:��x ���(|1�ߔ�Yj� MB�3bM��P�ƽ�@�%=jk�:�Y�W�xzNHd��Ln��RG~3��w/�=5��@��yR� ��[N���w*�1�	��ɟ����	��=�K�O	˵�]�E�@���P ���4� Zc��2G��#'�YA��T�U)����~{���^1YoL�p/�Ͽ3B�[�X����<���X��I���-ٲ"x�=���х���M���O�ѿ2���t`WNjd����ۭ�$�3�O����ay'
��	�uqǓ��U�@熆�gnO��3&E�����,H[7�����ʁtI"K��L�4�!.�⃡�{Ь���\i&�����J9�w�@#�B6��xyʆ X�cZЬ����E
�0��"��ٳE2�c;_&���7 Ӄ
*�7E�JSK�駹��T�,{F6���7�q;a d��7ЬY8�ۑD/C�z3l�V�_�2�~�T��=�ܛt�D�i�p��2�B�w�Hg�߮�h��LȔy]�v����5�!�FfGō�&��"b�gc#��1��#����-�~��ڵ�'f�o���&=@bC׆_���S��6�$)D�#[���������3Ë>f���Z���
?���O��âUi��}��]�P�	�,��=�)L���f��z������W�7\�C�ˉW��,b �[�bV��tz��˧"�(�FgZ�'�r�;q<w�������v'!^s6m�Y&���w�9-z#�/�����+B��Z�� Si��8 ky�i,- Sd�4`e��� \�8C*Q��AF!5H�"TR����ݨ�׮]g�c*��@�P�y3���o�,|�9?��ds<Bw˚���!Fp�A��R��(Hu1`X>��K��ީs����C�:�sѩҒ5��d��Zs��d�@�J�4=#5��>F?N����w2�����(V��o�%����/��D�F���"��쬬U�`�U��G�&\).��dA��#��=SϦ���z�M��p��!#���Ə�B{��$�d��%�n��c*ɫ}��֜^�[Y {kH�V��xR�/���J�����x,{�YC��k�}J[=��ٝa��F9��~���^2��ص����?�Y��eQ��D(y�d{�/�3Y	 D���^�� ���ڀ��s�(\��pöx�G&k�.�L�45�;����.P�j�ͷ�f�o��ɟ�wЧ6���d��X���}V�V&���Opʎ���T�a�d���n���{���_$]�?����Ђ�X�7R���p���p4���W\Jd�S?��9�:�#$y�@ͦ^��/c�]A��;�Eח�WۋG�,�)=�.�ہ�6�� |���U( ̏���9z��9 �Z�E�	�ܰ�d��x�2�+�� >��rPɭ,���F>�Ϻ�V���5*���+<��'0G��J|A{Q��)�Q.>y�y�o"��B}���0oCA�JBE�ɵ��a]�y�,�RZ"yK�)�����ڨ}�#æ����&�C�Sy�bsn����F�(�2��<�������%��']��(1��	�%�d�����0 �.���x� !����X0�7_M5,��i�$���8R����fuL�������w�hi���� ��Y�ù����:؎M^���$ ]w4�ĕHwB6B����Ѿf]�����X�ӱ�a���监�!�g_;����'�Y"�aD����ٮ��Эt0����g���/̕�׆$n�ۀ}%?m՞��cDT��Mפ��.�e���fc��Ӝ'�����XQ+��t+o�|!�3�(��5��"1�\&���z}�3�܇O6儺 s�|s�����܀|�` ����'�f[/�:��Ӏ�䉮t)�Y�drq|<Ux�cC�{��`nM��U�����Qg;I���������K�ˇՌ������td��⚜�9hK\+��?.^��(Ŕ��$ 鐲h������M!f>�T<ht��I��q�������z�����wk�g0X�V���*8�����xn�˱I��mޠ��y+��a��(�17	A��k���q� �TK� eR/C�)8��	���A!tO'�^�
sA8�dr|�;��#��nG�5���Y8���dW��w�C`�W��ߺ��%�F+�X��K�Nب9:��pc��'�P������_IS���	!|�}I��W��2�s��m��I��V6��0Sm���a��9�FK�)Bb��1��2!jE�wn�̩�����uĻ��%�֋�*vS������CȢ	����ۼշ�6�1�\恤ل�)��K��ʓ����"���u���,k�kl۩ޖ>V��B㝂bK�Ǎ���`T�N�\��믏�M�������+)a��O�~��^� D$7B'��nic��/��Fm�'���L�Q��a�`���.���4�;�%�I88���+J��/�?2̼�m)<.poK��.�Xrk�)�3N:ܠ�Ⱥe��S� ���\�����t���"�U���"�
7%إv���?�M�:DC�/H�gx%�/�;����'}n�~��i�-X+����HΘ����H.�'(�������M�I?[��V4���(����;�1Qc�ud%;��P`�
�%0�1Ns8  d]9.ʆd�t���Q2I�T�
"�6P��xD$�.�����;$t%Y��I'��QC�n�e�4��	���%hu����]�?�?P}0Ǭ�jDJf��^0.�r9hKV�[FO%ƺ�n??��=���šz{i�RS4�"�I��V��T�E��ȍ�F���ui��r��KчT�G���6[W�x���e��/��݉��=���7[��Fd�Z�W��<���n���^����2$�'�jPq,"�n�
Bx�D�pys�.��;�y�;uү��C�{2S�Y��Kx:�����4 (>��
HN�d�����GV�Нk�xE��^�J4���c�D�6���(�ʄ؍�@���O�����#���_��b=H��R��VRݶ�q�%����M�F	K�3#�ë��e��>�چ�# �+W���5�0�񱐃N��_�j0ر���mI!k�ͩF�M��D�2�?��k^�$������oCើK��(��]!�m�ghR/"ё<��A!�َ�{�R�r_�;��ɖ\�-h�e������㟟�����Y�+I��oљ���|'�|���U�*�{�Kgw�w'���Ovs۵i�8��x�)��m��p14���ծ�Z���LC��J�N��q����n���_��n����-�w<�o�C{���ބ+�w�O�	.r	}���s$���@ţ)����������G8�g{����+��}Q@_��)s��K�w�2���n��L����{p�v
.|���$4=ݿ�NZv)�̉rl2i���2�B�9�ix��� ˶�7�m*�²\FJK�ȇ���(&B.�V�+�E�ەv�8�g�+�H��ӣ���6/��H����[���0�u��5n�h��A�� ��fg*�HMI��Ƭ\���4ٶW������)Q<j `�R��fz�f�����t��1��X�w�&����JQ��K����Y2�d?@;�jh͢��u�-� 8#��"Ε�jw�����(���PD$�R"��@	�E՛���:o�Z�Z�:�P/c	��S쬏��2�^��1��dos����.����C(L�}W�������@��o>�$DY����(5*g�Ss0�hؓav�@@ �!��4x�*��d�nڝ����4��ﺱҙq;�{mb�]R#١��$�A���
W��Y��R�w�7���XMiEaca��dL��{*�dޫ�GMe��2�~��������c��G�Z��j�6D�S�Y�h�%0?��;E��<��A���%%����}��9�j�5Khh�XJf���=�bIl��D��:�W0A�o�U/��-W�f5sn�˖����:���\�Y6%7�� 韧��;�m�k5���h�S�`��EX�-���N�y�#���a"��^�{�����(s�]CE	;p�2��-r7I^�В�h�00�Zѿ|YK��Qx7���!��:�ByW��8ydZ�L������1���Ƀ�P��5ոƆ$����p��g��75��懆0�	)$�����}� 	n�i9�kL�q� �F]	f|���{.��d)��/�t�K0n�$�Ѻsn�k�ƴ�Y!ͷ9���ŠSD+�G�����] ���P�Uy�55��:�£�^vE�D���(����ft��?�W���5�P��uz��EMW�`g0�?7�mG.Ը���4�����P��F7.�E��Z#�=�*A����q���h:-���$!\Vط�V��C�i:�C�0^¡��|4��u�bF���C��_�Z(_'�@��ᄳ�SI��e�y�.�P{��+�(��.�����T`�ɍՆOaWG���9Lƃ�����o���Wo��f1)�Ԏ�7���;[}�Zgj��y�%��oe)��J����H�\h4��~����Mt՘r��!����1KQ�֣�� 
=󺼟�o���U
���I���(F��al�^|0]q�Zm��Yau���P�	\�a�Ds�S/����8��]e��󓲫xg�8�/T�`!�_q�jv̀
 �S������9]Y��A8�Rl�|�����=5Xx��2��8Vj���v��F��B���������J��ǭ�v�wt�,�Qߘ(�!�7i�{};;�[L��6\�O�Y,J��)�h�g�K�٘��h7���Wi�Wn~����V��h�Z�N�d���>�"N�yI��g�YV�xK%�������%�������tů��wDsi_��S���į��3�����Old��?��GN�(6ަ�o3���v��e�jwlI֖��v�
����2W�J�hS�b8��fHۘ%� z2j�в|���F�j�x�����F+G�?��1e\j�T���u;��#��k�4`��N�,��n_�=��|���;�<E�����ޞ���<�N��f����Y�~�J��ʡ������e`׻JM]�Ƥ`�~�8�@�ޣ�	���Q{{���p������:l��l<I�'l�Z�}FG���ДFt������gD�]�tHN��������}7��s����~o����"���)���3��CT65:N)�)���N�2-�]J�bn'+�!�������j�R���l��_ ��'���]�C,�&���Q?;Q�����5۫����r'L57����q��i|h��h��=�G�M���X�f{ց�O��?u����9ZSxn�$	�K;��Sq63����_:#4�s�s�Fc�F���A1/R�S&����,znr�Tb��ב����
M��E��u�AA2g�gic�X���}�9"h%2�/����ى~G�KZ�w�9���|ߚ�?N������n��Z>����50.���dOM����*�����-� ^LIR��F��$G����_��R�|k��k�l���2�I�-'���Ꭱr��+v3�%�3+�Q��&V�s�%����Ҷ[��p�N�+�le�[�'pL��f���� %�W����ĕ�8�+�[�C��ḄBނ�B�����v�:��9�S���'=�,\b�����-��q����&POS�P=�6g{�\79(q��Ƣ�}����k���C�r�D�E��Ui��h����~KBMی�:�j�b�Ne,������"Z� ��2&��p\>�gx�`��u�D9�N���x��c�w��]#���'Nu�ݝ�@&�c6�\���l},FTN��ǰ��:Md�ߡ�4I`�����nB�w.j̋���F��w�*l_!���sQs�B��n�,^lV��J��*����Y�ͽ�c�2�V��`3�cb����� g��c�;�+�����Yza'��{ޚ���?#�n��︙�Qo 3��Z��U��/]��`����7q��gծb�N�<���U/C3��4�)ܥ���m���h(?w�Sm��`MJkd�~r���cU��u�p�?�WL�����x7��[A���p�-���[9 b�=��eA��lK��'Zj�qI���1A�z�#�z��\�=����������p����Ae[x�o�.�t�s��7���]A�m=q���E�d�j�T�7wYY��@,~ղ���<�+�{��;g�����/O(&!�����'r���T�h;
��~\��%��hp+\:w���k��x�^;���Y^��S�Ǥ��lюTDB*�i@L�1ԓ8����[������Ê�&�+�U.I)���`�����x��K�K� مps����tP��|��'+��� ����zN�N_����2MF�{ش��N��I���(֙h<�F��(|�'�!V&���BXt�%�{Iܣ��G��-��Lw��i� s��C��kNI�Q����S�M����h�+� �<KO�"���ՇK�2�]py��1�X2� l��#!@*���SRO>m�"¥�F�O�Ⱦ��?e���:��D" C�1�xį;��i8��)�?��z@�M^��=)�t�	85�v

���b��-�-�@׊�qj���(�%�*�Oe��v��ю��j�]�Y�`w~-e�.,'�Tt�\��gV���R�`+�G�g�P�i��3�d"�{o/"���i����d�\Z��e\'�l����.�$,^/=�������̎�.k4FIv��O��qd�g�<+�bVcV�į�)��%��2N7c�uSU��xA�<G4���3�D����c{���=��YT��d�;+�*�������6�mڿ���<d.1K��,�v��//�UXXxT��k3^ҥ4�H��g6}�w%���We��ߊ�ّM˶�@�z�
f�B�T���	�"	��g-R�Ҋp>���,-��7�8ɊA!�8��<��m�������rR��Z�~����T��R>����]x2�c�.ſx��K�s�Y�{��5- ���~*.�\�U�FD��P�D+N2lbgy�Z��9����1sԭ8������fI�����I>���%YC���7/���@g����g4��,�u5���� QBF͟�ij�`C]�@Jm�L%�r;�7��U���ɕg�6��]�w|�9�i�uU�Y���̗P�(X�S;��%�l\�BS�$Iʜ�E��������U�p�o3�j�3�!#��I�a�0�a���d�7u���`����A�X�qrG����:"Q:���5��pH��v*L:���X?��B�^�H�<���G�J,�j|/|�`)H亨���{�Q�C-�4�'>�!^����|ed����b�Ixh�n4O�;�P�V�	�n�6z�EN.����Kub)\���΍q�U�����$�k��zp��7���S�`�WS�pJ��$]����^&�&�2"��:H��Un�ֶ~ <B|��8�W�R�7J�6K�Ѻ]����:��L�"��+I�%��FF�f�2��H�L_� �������?������-�����ۑ�,Qw����$�H�Z^���P�@��"mD/UƝ����9GC�)��P��,��_?��Ν�12�?f�1;;<qP��'��IS�l����K?���'���T1� ��f��� iٴ$��Xƴ��7^��L��}��m�G�T|*ԏ�Xp��M#��fU�^����S���`�nM��W!Ӱ+�&1Oƒe��5�@\Z­z��ZގTD�IX�����ϩ�jb����l�5a�sdO� pY14�f�z��%n���FA����ܭ�6X-�|�o�n�@!�ay�!�L�)�y:{`1;�N*���s��NP��{�6�@��u�$����ںk�6�����[�R�O(��7�'˻��Pm_���p�c�� ��N��آ2l�fKjOo��c�Br3�HI�z9����M�⛊�S9�c��	<�D���^�V��w�,S��Y�5�&�����54��w��#�4���鄎����W&��fV]#b�{�s��3'�!��#�-�_'��J���d	I+Z�q��8AP��N����X�>�+��8�.�&=�W���!�4y�;BTQ!#�H,� D��'&���ha�Y<~��ئ���lu��x1 [~�'�0Y��e4D=�mqIR�����E	r��|��(u�{
].m
�����億�t(������#���`�1�@�ȴ���kQ,I�<�`tU����g��եI���V��"z�}Os6���k7����{�Q�6b�q�[�i|  ��2/��*֝���h�������I��a������A>`�>�ɰUΞ�OZ�X!ad��B+�W>��		�bш�^�[Q<L�������t����ʲ��D��2gU�>h+�r���� �-�����]M,�X��ܖ�����@�+L�Y�/h19idĖME�����\�Q̉�f�O��#��RG���Z�چ���=zZu�pn*�RT e߃FG���)���-yX��3�y�㋙��Y5�XF��}t������ST9<�2�%�\ǛW���<`?!`��j��9�^-ܠ�I�;3Ma����J�aS�'�L	��i#!���uD�P�����u�AD�E?�bA_�+���_n��Ws�b�g�]�n��@��~H��C�&>*{x}
��"Ű�i��*@�s���*,�%?;��~��ߚ*x��s�ܝ�l��o/�?�,"��eƸohD�r�@b�SL)?[��`1(U-��q�د�}x��4����:��(��]f��0��U_��7R�[Ȇ���GΟR�HW�E�CN�ג�?�Z�`:�_�78��Fӑ�	��z�d�$o�)h�[*���f噏��m���C�3�b��}��Z�y�HB����T;,�qT=���!��R�#�QaE&M�+m�o|њ���{�?�P�^�P[ruh��G�CP*�|%����7��+��|:�{�J��!S�	S@��_��IG�HC��V�-�z��9�R?K��]/hgu�σ����ٌNZi��*�;��i.�_z��38�V��1�t��"Mn��;^2| 3���������/-+���Rė�83�{4�	*�ߞu~]2���[[�|C<x��X�/k�D�U��g�\�gF��řC��b�oFF��QM[���`r�ێ��7Sվt�i�����B��e�"��)p1'1h����߲ ȗ�u�#�ڥ����y��I� d�9��@��0Z�)�	[�Yw������vnZ��v�'��TZ�/��H�O�ϔ��ٗ	�J)�Dy�ꁌ�|�xP���G)|�0�t���nH�4kg�I�]�8$O�
=�,^�ޥl���\W2%yN���)��u
u+�.�J�"	��(�-K6��9�
&�~_P�%�i�+c�M�ڻ��XC����<��智3�o�3�[�ɬ��@Mx��c�2��_�H3��B�����C�:Mm������km�݇O|_)�ކt�u��/%��W`C��ǫ�i�T��	H��Kq��!O��&0��������]-������CR<lv�XPM�g)��d$�oз�1mH�o�i��L��l.���p-��$|x����,�X3�����K���&9s8 =l�2���eP��0Y���K�d�͠=����Ȣ��D~���'F�K�a��a�,C���\J�U~���׌&�8H�z�&ʄ�t��\֧sP�\�XcO����!�1�����p�ܛ�l��x�4\?[�sT������C�* �96QD3�a���-�}��X�(�z�u���7�򢠐B���dجr��J��Go<ǈL>�x2#���"W@|���P���u�'���N!��$Y�n.�z�xl#���w��s�9"�//@�h3w�=��sŧ���[蒪��X�a�N�e:��R�y�c0J_u���Ȱ��ʧ�q����|/�ѻ����KO�~��i�&�{��_A�q_�(�M�/���8�������s;����s�?+�����zw̍���a�hp@��g�	7�e�-m�u�w�TAT�?3?�^�}�il�K�b��yYύl�[�iyϧ���)��m�*y�(H;B�#+�3��F�HXFe�Z��(�߮����D�=)(j��w�P�o��E�ލp?�y��6�U��@N�g�z� �@����c���M�"F�(����$Q����nz�Ԕ@�:q�k��&S6�4���Iq��+E�`��u"~��Ŭ܇�q g�X�$L�);O&�B�S1Y�$��R�?�,��Ve�o��o��﫜�����5'�(��1�S���"�(�{s�TW�~Ķ��.TB���c�%��(8>l�����
�G�p|�ߑ��Eeؼ�p��pi��i�r	�l��kdot�4{���rC���?�p�v2huH�,G���}���L�SH����X�3���PO�6q������C��1Y��Z�.��$0c�X%����w^�u���l ��=
��x@��i9Fz��(��5�u�G>"1�S���F�������'�
u��L�EÑz)�B��L#���2`ˣ|rJ��/�~��|}�	%浀�ȯ�����a�����c�v5�Ow"&&D���xUp�( B`�i#Z���m��X��3u�dҼk�<��6;�xvޛ�zB��}�,`"�X
�8k񕄤_����U��B�ъ]���t� �e�hoΚ�� gaP�a���P׹��t`�����Y��#ɨ���{�s�1=T�R��Q�5�99�'r����M��n�!�{��A����8{9�z�6�W�)9��^��E�M)�	1�2p��B!��Gܨ�#zr�����E3G��:5���Bx)���:�z�S��8=���c�@�v�<�����z���Dv�@y�p<\��O#���J�P��<z�S,����G�H��y&��Ov�Lh=��+��]a�?(!@��󶜟�+8$�3#vHZ�5��_�J��%�֞8�m�r�}�?�i�=�|��
�r�P�Um~�>�'�)ٮ�
�GV>0ޥ{ʍt�ۧt�D��mlOȳ��#�^�������,[S��d�7*�3�ޝ�	XX�Ԫ���^JM�ݞ���W�@���\��l�o����._-s��[����E�����-Bh֗�h�����a���fc�o1���!<����ds�݄�}`|�"i��{D �*}id�x�	)
\S���@�E�����U��QC�F�Q'd�d��jg�f.�����^���Yg7ZrG��G��Ŝgjn�mG��.����)�L�V��^�=y����Pt�S.���la�E�v-���>�H��ngݕ�&��V��r�GS�&��>_Z�N���6}��t5H&��K>��@���|�|*���{�Hmx[Y0�m"oW��rr�h�� qs�����ǖ(�^�@��^i��ǩGM՘���߮�Ud�Rᵲ�OMHҸ˖��h�n����b0hJ��^�$ozz��R��z^�h�%��� ����R���Y�K3��(~f���Z�Z��'=��w�%��ˊ�}���}"֜�� -��ޅ6�g]���h$%�GWͩ����Ro��t#��ͨ��T�,�\F���R���5��um�9Ѿa��
�̼�{��#������j��\ aN���k(�'�Dx��7��{�b��2��@���ʖ �d(��.��_a�٢c+�oz���3�i�
��^�[pS��d���"���wM\�c#�h2b�, ��@��Gl���ʉvtQf����4�rXQG��0 �g�L\�;zB�a�>��$���v����Y��Kz9PI��m۹YN<q�R$�2�O0�����h��+����j��pS���z���w�|5浺/k�[��Z�����|"��%&#��2���N,�'����:�CzZw��-U�ؚ��ü>����30-#�^�UQ��|�΋GE2|��yN�iK)�!�r0��uZ��c�9>��ɻ�,����O�2�(�܈ s�},�շYB�^-�hpO'v�ٞK���r�4CK��e '߬��h����=�t�[ISY�6خ�Bv&M��=͡���Bn,rB��b�R�^,)w1�'z-�
@B� Asu#Y�B�k_nY
ω�Oq�}{�7�g�gR��%��^%�?�����`�;E�^j$=��;K7(Ps{��<֊��4����ն����!x.��
I	��D�2c�������:�
{��~�!�sU��q�Ğ�pl�7�ߋ�{n f� U�CTsB�1j�)>�9�k��.�;���y������=ϩ5��Mm��^j� ��v�.�4'��ˊp�=0$��<��thO֤��l�y��lC:4�a�"��}ro�rn�_���(z�����k�e���lDP�Y��rֵ�q��. q1��y<;x�����-T�k��XSk���m:��}����>���	D� ����ZN�t�M�Z��J�H�DS��#V6��	{b7�]�_Y{w"����S�ç�ȓ��Z/�
5��\�������(0��a�E✿�O��Ī��0�B ���U;.:�~e��b8����@y�*�~4�&�����,^��W�RW��ę}-o�<��{n�ͥ�RE��C6��:E	�\��Gg�r�Um`�����'���˵���j�a7���x}�~�ڀi�&0&�q��4�r�"�_o��%�1)l�Շ)��h5�%y.��������dHT�Ϩ=�@gn�*K���17�^����W��䃂�(�X�V^��U���<(�շ����z���Y����d� �RϚb�o�
g�*
^�lo[���"�)�Y��H�4 4��=���M����:��`���G>+�h�q��)o��Me~�$!�n����CSg�Pw�����t���'��~V1��:r�ۻ��:�,�8m"�Ok`*�H�BsC��v���=�QE�{K�XK��j'�·�@(���Ƒч�_�-�Ez_�5/��l����V��P�
؄i૰V^�n�Z��Sd��IS��:<w�y�f���P��?X�8x��\8_EjVb�%SS��H���<�ڴ#�;z'�癆�ߍ{z��[�9���MT��W��;���8n�l# �B��e��/�Z^�oOE;��u� 
��4��QÖ�^Y2�(s��\�5���:�B����T8� G�?���P�WZ��>|/��#W��a�����m�� ��M	�^�I�А>�{��k^�̥fL`g~|���MSt�X୬��쒒���!U�}	�a���"<+�a�8b-\i�p`�iU��I�Ӷ>�B�8��ۂ8�☒r�R�ٓ�O#��V^�}��f'}���k���]�l���B�Ol+�m�ʲ��{��yu�I�RY^��� ,��4%:�mb���a2g��8�|���"ÿ��^�5Y�P��VHĉ�۳��g�]���*?O!���y�8�
U"@�[��w�b��:̏s ���-h��ccC��}K��QjY�x�?j}��$������TP��؞�U��:�ܒM1\�,!�df���^8�	?9��OK�\��0��7�'�Aj��<`�^��R�I�@p"Z�FĊ�����K!R��9��*��rQb6�n Զb�Ț���V����bۍm�!Q�����`���/�W��/!�tMޏ����s��M�n�G�gh,L{<SgZ �@jE��zd*�n���������N�v����&8�W�'�}ÐY�/Z~0�) �D_D��s�KЭ^F%3E�)�h	�W3�����D=��Eg�C�����{���D�21)����mP�t!���|��oW'"Y�/� ���ˋ�9������G	��2$$2��d��P+4q�I\��<p��I�N�zzY��l�'�->mY���モ�wm��"��������Jp�ot������(�éf3�b�7�Xc0����<�v`�m�G�h+�����>� ����`�Wd�c� �`Qt��x���&�٦w�;��%��ku� O��XȺ�GO��b������*��;9d4S*_�Ѕ�n�_�������3'X�[�\����q�Cp?�6�l��M�	�<�?QXj9��2��ն�2a�(��ѐT�Wښ�5�C��pCC�g~��RU.��	�>��L`u� [rE�r�2��j��p�e
W��!%�`��d���gX��{-:a���$?�Ϟ��m­�՘�jXI�ǐt���R<�!]�\%@�\R��mOa���Z�����I8P�����b?�S )�nMPU��aw̅�S撩ĩ�����L��h�D`Ӫ�8��/P}�+�S�3�Y+������ǧ�߄���6;�kL�98��&���&jP5ٵ{c��qe�������RC�L��{V,kFS1����j�CB��F����I�5�f�2@"�'!�s�҆����[eg�)�zE�iԻ��(�sQ��B9�o�:2|I娍R���� ���i��G'a���2�\@�V���ȸh]���Wl�m�:�(�3�gحϩT�����y�?��n��!0�{��,֘�5�����`k�8���g��d�:�RaY-�V_J����`�3��L_��� ��{�����1Y�FՐ2��ff@k�m(�T�,Z.����_���|��/~�h�{�Г{B�7�Wu�W<T�kO�n[@/���PVCC�f�&���=�DQhvԗ�moݔ���� {F�J�Y|v����BB�M�F@m(Q�'�d_n�W�(�&����^h�a��VAq
��
8R�XY-�i��C����+����F�e�Vo.�]�N�vX/�$B�{�q+}�Ϥ��Ph�&[��<��h�(�pSv��_X� �I��7�8s�Ќ�}>�J�_Q5��݁���l��{�����e�7́����2��
S��H/�&uV�����"�pztz���Sl�aȯk��h|B1x����t�Z�����.��n��+_Z1���!h�Xf���R??�~�Ԅ�R���s�3$X@((MZ��)��ߝ0W
6�H���`�$�����+��3�!O�f������O�br���
�5�%mq\}��vV��A��7�����|�K�V�����3s�0q����A��9�cyDx5&�X�`�}2bF��W%j��2�7Z��/�{pƩ}?��f9Y�sJ
=获7����V�Y�{	z܂-*X�G��U%e%�������g����Ve�n��LB&�k��U�`;~)_��I!-��i��=`��ߠʍ.[�!w) �,呥w��I�o���<d��W
������c���Sd:��5��ZbN1G0�/�M���n�W�A�eV\���Ϩ1�K�{g���sM���YHϾr_����қ%��B#p<r�ٻ+	>6��+�>�
'�NR���y�!�; �[ڟ}f/y�n�ch
��FTjE�ep�mì�ܕ"e����f�	�sl�^y��X�d�Uh�Upu:�)M�p���hP�e�����[��.*1�����NR�XI�Uk>����|��{�`�I���,&@�L�I<����>]�'������5VV���p�:f��P�?������Z�0��
&�o�@>=I�aS^�����<�g��;����	J�l� ���q!�Y�6Oa�9��ʿ,��[�*I��/|�=�?\�Q�As�����PMr��pat���	���������_'���쾵����<�u��+���W��q4���x�k�D\;o2�0�*<(�v�F��������̧�1��m��G���	�SGo�[&J��f�%������ީ����L�X̗1�C{�K���C�߫�V*`�-c������KC�	��nY�]���[�Hy�L���_g- Z��k>�_-�C.4.Sw �����d�aJ^�.�5G���#��~��{��O�(W�5�5�*���ī|#�����Ɵr�ۄX�ߵG�)��0�eX2P������r/��\�H�O��Шm=�0`��6D��z��"��M
w�jW繷0%��=<�5ژ�'��`���Ў'$������x�;(�f׊�Rc���˘�s.��Ƥ*�v-��X��#0�_���k���!Ц�-<6B�K?埤#zj�����V�g�ͳ��[����1� ��W�^� �n����v6�R�U�-G����ۖ��($"�W�wFG3�� U��)ц4��� bg�F����v���0��K�
�A})�B��]z���y�#Y �;Ѳ��1�ɄŔ(M���y�,.B��i"N�|'�[T��	<��_yx����C�7��g�����k�����I�8)���Cfxyfe�N�ͬ6�����ި�F;�\�x��Y$C�@�	��0C�G�~		 _�d?{ybYF�'K ��w����~cƊb9\B�ل�RR�u���g�7p��C9����<5gu���+��ABƑ���[�!b[�}r>����L��A�Ww[{���C8�Nu�7�qw��g����xu�?({���(Ƀ�o�@ѹj��h��DIF�,�Y�W���c�ͳBb�I$�c��i=S~��8��x�/���zr X�5(�!/�5� z]?4d�~�Z�ٵL�6g�����4�]�+��/F��h��\ļ��#%_�]�WY�UA(#�ȭ=��P;՘�z�Q(�
��S�0Q�=�{��tð�Ҋ��4O`��GŽ�ȿfQU$��K�f��S՟�om|�9�����?�t�sW�x.F�a5e�Zʻ�}=~)��>LV��#��� ޿�G��\�˪�A�,N�ჶ�\�|�ٞv�J|~D�e�l˭ƽ�}��V�զ�� W� �2�C�%i��$cg��(mCc�����sXHY���M� ��_\�)\:��u�{˾|x'�筥\b;�YV�9�M���"��=Fom�<�>�I��q�*��N��WYf��~@}{����m�'[�C~5_9C����]Z!�9�tN����)��2R�Nܵ����g�r�:�Aw���s0]r����ެ53@.���*P�6D\����ؠ����Bb�����?9��8��\f�B�0'�	�ԑ�+�O��S��M�,hւ9�7��4��ʮ��@��u�j���{�q��~��Yر5�ȈhZ�jqf�DN\�G�[Vi�X� &j��Q�i˒o�q��Q�E`�L���ē��ʽ�Bi�d|ǌ����\ƍ��{��v�ᎉ�}�须��=I5���p{ߥ� Y�P�ȅj�w78�F����V��}?��H���d�����8f��RG�� '����f��(��7��?����c$ɲ�Ehƾ#x%�<`���
hΦk��ԟ��U�Gs�y���t7(��^��۫*�w�x��s�Cm�zS�k�`�Z��zN�(E�>0a+�����N�L;ă�2��f,ܪ�C���?���ϟ���]���֦��tK�"��G��j��'���>9w���/�����^
?��4���X�z	��$'*YA� Q_�3��S������E���Y0����(��ʏ[�B,wF�)�8��E�J'[�do��1��܅���I���g��>(WN�zr	j(+p�ݻ|��ά�>\�MJ��c�����X{jz����5�^8/Q~snXZ�Ff��E(c�g��>ᯎ�[-�o#6U�0<S�ǵϔ)M]�I�7+1���|��(}�p�N���%/�T�ie�������(l����Cg8�� ?.�d]�*T�21����-?{���|(�T���^�dz��'��!�8�ηn�����5����c��m#�)��5=i���L�n1��x��QF��wRJR�=vo�?��vU(�}K1��R���v���;��jrL�����p��!��b7q!<���d�o�������Y��Vf�&Q鴁�l�6yz�ߋ%��t_��9H�f���تB�yQ�d��5|�zS�U۷^������dg}t�Cf),MVux���<���>�o!3���Dyx(VҪ;^&H���\�Ym�]��1Bq�������f���1%��
���4Zm0b0um�Ѿ��ӽ�'�M܌��p:_K0Y��J�CO��KyG::ͦ*��7W�
FA��k������Y�sm��d~��A���/2_�����vii�}n���������v���Sfథ�M ![�Ӧ�G�� �W�s�<�}��IS���x�OM����K��S
�pG-J4�a�Z&��q�&�%�x&�Ճ:P�����+N-"pE�.�S�G�M��g�o)1UV҆�^`���:?,��TD�`A˙`nW�z��=%���%d���Lrg溹V[h5�-xp;.���}�T�=����B}M⤄�7��@���D�e��ٽ5��J>������k�Q��D���7Ng��.|�cd�{�QW�����f�#�|A�Z��#�����*��T���j�E1����<n�56$ ��'�1�|�5�z�f��Z�[U݇.�����֮�}Gs��ױ��>�i�̉�����+v�v��u��O���
��s��|�<+�q6>�t{,a �N	�EU"���u��0�JaԀ/ʲ����r�~��2Ђ�[
̋��!&���a�ND��=i%�\8���(���7�P���HI.��U��V9�9����Y��Ҵ�Z�)��4��|��T%�iH�"%��I��aj�1��x}��3�<9��z�j1y��?P?1bE�[���Mc]b�jD/o�a��@��;�)l��$���X<��\�70��������5`�f�C��LR݀��:�2�͜5 ���pq����o��3,YlEJ����׈�xDu�d2��9Z��$��I�9�Ψ�F��ڃ���_�h��}���\q�p=��1v~��O^/�e���߀�ǲ��~�6��C�o\�3��-��He+��X��/�z�m'�'��V����幬���.D�/U|��\T	KH ��w��m>�TG[�T�<�k��]���-�o�F�īE�ns�O�9B�tN�����+E5_�x�hѸV�!P浔`�D�(B���{�$0,/�>�����׽��O�O<�K��dB�����V�k��dԏ~̣�?�-�n����Ov����-���}�V֞���ru7���-�V
�����tΩgQ�ҫC3��J.1��a�&�oj�-��EP�@����;釜�O�_~��'��Y]b9�ė��\��\3��.#O��\��@]zn:1�L����w���W��2f,:s��J�<�����"	�������()�=��xYU�@�	�mN�0��,x\���Ys�����!N�E���Lar5�c�	�R�$���e���?����S>XJ��-����tS�����>�LxΩ�/6v;��Üh]��m�h�l�@�>�F�n�I�9R67�&�-�a�j��C�&7j�H9��t肐��	���8mS�A�
��*�u��ztN������nR�H]yOaR��@�.y�W��M��1��X�\�v�q�"Y��q�(	�e0��\F�m�e��Ņ�	��!$�2Gdv<T.�)v��;)�4ˤ9�[���Lns*O<�������\��X���z%�y��Z|5�����LD�� 2;jS=D[��j3�n�`�klWC��+��
��R9�^;-���}�P�Ј{���TA���>����I�	�Xh��'k�Un�r��=�\ۈ�Z%c-�e��6{��'hLsw 8Q$X�lpAO߹�U�O�2fW�_#W�C>A�E�DP�߻����-����^9�v�1P��j�0�EL;ވPo,� ��'eF�
PV�eeq�����%�t���/��@F\Ũ�~e�Q��z�2�{e�b�p�!�Ww4'��缰��a��W�擌S���'���4�n|w��9�uy�9��}���8��w�f��R�Q?�i����o����2�\}P@���������I�!I���q�R��G9���X�Q=�F�K��Բ��j�����׌>��N���a�h�t	h"���v�ZH=���i�V���M�c��㊸�$d
ָ���J�lB�	��u���(,��[2�r�2!�!'k�U��cBK�b4�`l�h<��J�z�
I��>������v:U5��`#�_qb��7
�=��R�^ܪ��P�����[�T�n+����ǉ��Y��M�d��G��ܱd5�ڧ��F��_����15�Jl�����k�k%�9y�8£�KN��x�N0�l�TV�樽�`����6Ϣ�5�� �N��hV�i�[���u�X�º��ˆ�|/��ٽ鯄��<��O�C#�Qڞ�E4�Ba��?�y �
��M�%�9�(���'~�%,Աw0��M�ΨS-H$ћ�!?�7T�~�$��>��
��S���y�4�9��M�ƀ�ʕS�؆_��|bM*�x;��Y�\/3W1��Ll�hΓ��#���-\�bɹ2aV�� �����NNxu0�$J���A���6Ք�>� ��q;ܼ�鯠0�ЈPvtˋ�P�S]Fڕ� �
y�`�5~6f����?�ج��:��0�:��?U[:�ˈ�^��V5;5�-_x�>?�����vl���I��˟F�,�W.���4�AQ|�j(X��\N��{.X�M"�����lɍ���!������F��ū'��l�g2�D�2�Qn�IQ��bz&�J�&��3����g]R��=�9���7��FB4Z����a
=B+ڿ$*
�V���G"v��4�k�U�vxUGf3��$�j3���{�
UY�I6�r�o_���b4���?ؔ��?zV�q���l䊎��Up���3~��d�2���ؘ��mꏋ�U+�z���9�,��]:<�l	R�3lBrϗ$�ZI��	Ձx�lc�OM,|��"��Nk�2���a�x1������Z�9JD<0̌�מ��&!F(DeU�XeF��H%S0�S[U�c��4����א�s^ɘ	���C�H��z����Y|�ʇ`�&O��,.w���^V1v�7�'1���u#���̴�AGp�!6m>-�Խ�$�1�q������.!+Dke֩Ȓj̢T�s���@v$���_���dWϑ����i�?�[�|q�	ӹ,�rUh��9m5��_�́�*T0�jm�X���SQ�Q����L�ÅP�GlI;s��蟞��3�c��pA�~t5�E��J�C���$��î����]B�υ�2��t�*@N.�#�>hA��-���4$��ǽo������|:e�;u�5�'-?uU����OcS�%�z�ӥ�4KY�"$XQ)gE�����I*M��<2��ĭD�P�ܤ��Flq,�3���������m]�*A�a���~���&k�;�������A'O�HƊp%(f�؝�Gᚰ v
wX���)��O�֛��EƮ%�"J'kO�`�H��ݒ���ȈY��m eD
6b��s�#y �c?��o���F��p�!�'�Gf+,Zu����]�f�ԭ~N��Lh���M ��LG!��wO��2�ν� �y�+������Wz*,�14���:�o�Z}��$;�݉�KmO�H�cd`��:�c��]�dc�� ���P�����9�t��蚘��yُ��Sr�Y�.�����&@�f�n3��-�i��y��b��������*�	D!rx��S���$8˾�p�9JT�2?#���D�~�M%��(]��O���)�gy��7<+��l�.=�t-P~���$��b$5Ϗ�¥.��2A�C.t��ݷ��S�&�q�3���0���H����Z��T���p"O�r�6z�j����?T�',�;7��{w�p�DN@���r��ˇ���U���49�
53�>_ދ��|KR�A�w��Ӣ�}p���:W}�"�m��������`[x[N�9����_bJ2re������U�C'BVU�b�����5��M�G5Y ����SI����R ,���h���P�/��`�����r�&�B�m�o��1��ڳW$s�����3�����6�:��L�DTˎV�Q8��A@.���Ol�*)ɰ_���ӏ�Vk��)}�hiԱ뉸DYr,��6|W��Dm�<z��� ����4i� 0�Ql�SE�e��!�"�F tk8�KE/BfJrY�i���'M��Ey�o>+�h���^.�~I[,Ws�HDZT{z����yG�)e�1�)�~hU�Rg8aO�j	3�F�˟h7�\N
�ݷŰ��v�/�����[���QY��["�ёT;��xY",��P���&�m�N$����׻����g��9�Bd��b�Л�^���]�����p�!�iwo4���M��d�.��+�
�����������)S���㍨=����MS�Y����� k��x������@q���s�w��u2�������k�d+ù�L^�I=�M�0��1�l_;��rK������_���X���$C����ˁ(�;ۼz�4j�O�ɰ-��?���>�tLwG>��NЧ��i���iX��$RI?b�}O�Z��.����t0��_*��j?��ng��Ǯ�2f�|�
�X���͙0�����e���Y_�ˈlg�w-�n�]X�r��l|��ܭ��hp����Td�'ư!����e���$La^�Cy6����K<��q}ZF;q��{m��uQ����|{�Ť��H�s�����L��cP6ȓ�Y�6}������T�>	7��n<9��C6�čU���[�&sl���	N�{L�(N�����҅�J�v�:fq-{��9���uE�Ց�]�����,�n�����r�uFp����nG���l�x
_��
x�*ɲ��'��_�*آ܆���%9�#w�2a �PAj�� �6�\��
�L=E���vX�-����=7AQ�xs�}c>М�/u�L,�+$�P�?pw��4*��K�G�(�~�e(�G�r#���u\4��Y�����0r<"70nv�'ũ.̰��3�����%8�(���TIq���i���e޹M%�}��z'��M `���A�������h�햙X��.f��i�ewO��f�q�h{:��b:ji���]�mzlw�`r`�g�eab6n�,�H�B`���J�<��m�os��4?9��-�MrX������d�Z�`؟�j�R�h���"��_�S�J�U@�cj�´&,(��3�P3=j��19�R��Cw6�4�OԸX�?F��Ƨ���LG]����9
���]��G�؛Bi
O�8��*|���ݙ��YK&~���2x +I�B`mvk��%I;��a����o�[9lip�@�hp�A�e�^,��M1��]�o%&I��=�t!9�k�8�fOp�X�A�����f�!�&����Yɐ8��$"�꾒�o��
B�`rjlw�'7����OɲxZߝ�"�d2��-���;��.cO4�Bp�/d��v��Kt
��ǉy1
 �w`O�l�h��b3#7 ���"�H���Q��t��@Ȣ���C�qF5,!��>�����.�I������ү���"~!��-������h&��T��>A��!t8=dW�뺢�%/����6G�+{��:&E�"�3��DH�I���Ѭc�Sj�9)G�L�	��	�J���d��T%�#��_r����T�pC�o��5|����I���>��:w�_%M-��Q;lid�qX�vKb���U_b��;VS������ýk��2�QK��G
~���vd�y��Ac����$j�=����Q�DZ;���)�[rW�` �x��i�n���.�I7�����[1X=��yj�J�=��F�.`��c\Kڗ�9�sV/<L��$��	!8Ab?/Y�nݔ�Q4Y`E�9��D�N?uHW�r�4�$ED�#]%*��0V����2(�Yt���A�\�v>���_n�F��l���I�����q�x���8�rYA���P�j37�Dc,.)U���K%1�i���t���k�E��.EI����Ԧ.	�Y,(pc��'�N$��(�W*��hP٭�ٷN}:h8��9�GS)�/���?��E�\)jq6ܹڤM#��k��!A]`��ںb���@,m�SV�9me��k�UU�Ŭaگ$4�_E���R>=�|}���P��$��=�8_��rp#��%URc�&Z8a�J�C@�ԪL�t�K�>��w
CzG�W+�-��d�ܝ`�]%�@{�! �C������"r���&B�^�����9vq����!������1XG���>y�9q��ݮ����k�}!ˁ��c���mR����X�n= r�u1��}M��@��յ�ޚY�5���i4ڀ!�S@�T�ل�7NĹ(�%��y	��zGS����2��f�f9�~�uvm���z�f',O�8G�ut��ME��_���q��=51�8Zn�G+R���� P�Vo��0�u� k`#)�E������#�Nupd�y��M8I=5�Z�G��������@J.AQj�@gә�T�������0��+/�'[����~��
=�D���u�{��㙞�7���	�w���z�A$R��q#xyެQ:���7���e�+��c�=��L�&wk�%���5	.�cّ	����9>�"�&�)8����I����"����mN(B�>\Ũ�$�6�q����#����5H!�bN)�Eߴ	C��TƟ�����6�7Ce�Y��t����J;X^5�F���jX$�rO|�ä�	`���u�[��F��7	jm΃��"���2�5h1ӵ���^����Zk�(��T� ��Ug�$�&<�����y��M`N��(A�Z��1U#<ѳj���Q�$>��d��kC_{�lU�q M�IX;N��A��&��F�qш��#�Yx��iɖ��`��o����/D�V�AE�89�c��ް���@� ��9Q�zl?�ɿ�Ω��z�x�����=��Q�^lM�d�2�~�F��h[�Z�jj*��Dh�ЌR�&��6a���+�~���'u&�쵅�@K��{�U���e��LK5���r�Rww�
��(p�=���$�iJmF���vl�p��<��G��|)����#��Z)�m�D^��3�,;��z�y��zH��@���,>Fc������\�,1���s��O<���F�~�⑵'ޛ������'�~��Խn���W`�#���� ���Y�ss�5F(	�>fgmܹ�̟T�rW�C2���ǨE?��#g�ҭ�\����I�6v�P̟�t$��u�p@;��*�5Y+��F��vW����)�K�HwS]� B�2o�g��8�DDe���$��s�� ������ɋ��-���l��~?N�o���
I^*Q$b{�c�5k�2�a8Re��F�����R���Co:IRq�w���>2y���0�-�U�ۀH�J�w��K��Ô����`%��]�U��)<�ÌU�60htR�l/���u�im/~:Ё��ɚS�c��>7y�c�~7���HJ8�˳e r����C�Dw_2���x!����RcB�t���͞n ���z�[I
׿F�3�����x�#G��s In��f�4���JV�� ·�2��L�<���[5�)�@����2n5��K)����+�v�z$m�$�*���1�F���#��$�4O�%M���+ZS�o�.��B:��5�b�N�jޝ��kHβL�QL'-� ,v?�+�Tn����)w!#����{2%Ms�]�_�ovIN���@�������h=�Ow;uH����L�j����t�~�� ����iѬ����p�O�����Ś�0�0����-ڇ�XZ77u�X���Ky����ae ��X��s��6��k]+a�z�|u����l�\��k�z���!�:�����kjⷦ��nT냌���R�s��}_�坑u6�n))������W������i&ur��9,ꊍ��~�� �~ed�
A�f�ٷul���	���F
�7���n��d{Wj?ݑ�f#���r�%����#��m0[�حケw@?�8&��`gHU_�]�+��:��xMP#��rx�yr��S�����P���눹��{4&C2#���>	��6��9}�����S1F/��l�^�
�{�/Ȥ��*/�T�7i�	�jn��d����g;�u�a�]L����C�S��^d|x�a���jE�ʡf!O�*?��Q��5��{xpOT�_IQ{î�}Y)5�B\Kǭ8:���_��{|m���=w�ʳ%�P���,�R�����
�+�h[�zh{&P���#�����/j��[ӣ t���{�U��#A��FS7��K7�H���@`]������*j�r���c�������P�K�-�RsD��1�0}����{�9LJ�/щ���M�f��(d��q���벤��e\D��t�M��
+슺�݅Zl�Khԉ|�i�_Xq��Q5�M��]zm�ˢ���!@SI^-��8��;���h(�`�������CT��hȘ^����u*��훖�XLd���3�#�*C+~�+�{8&�D���_�J��{���Є�@��/�`�_qy��L�+���᪋L��1톰L@�מ	�Ԉ�h{��yZ�^�ܫ8�d)z@)>�(��>/�ъ�eV8Zjh���N ّ}ʟT�nh�v'\�|{�Ӗ�K��/��/�ܓ��]1,����8�������`
1��a�JK��ᵐ����-�2�u���_���Q��t&���j�ŶV�UK��[�9� ga���00�_�4RtuV�]����R��~�?�H���X׹\�U�M���9=��8'�Q4t7�@;f&}�3�<�`�%��q�-��;mc�X������B���ܾ��!� ��N�\�յOuK��K���ˀ|�do�A�n�B0�*�+�M���+#G�`�U���s��FUdkw~��J�IaE�v;�q��gzϾD티�z��AG��J�?�o�`�b��H,����������/�<���a��"O9H����OL�z�W�T��Ayf�����1��﵌����=8�b�tj��Kgu��@Y�p�!%�H��ɛ*�?�e��<������R�6�CU�$�Hy�]�fO�A~�W|�(�����]�ΰ�˛\"}
@^(U��"�b��h���op��\]l��bJi��ZX9�{���ӊ��ͽ�l@�
fw}��'#Z?�Ό("��z$	P'�V��w�/�O�N?�{k�.	��X?��#��B�:ǰ-�p;��ƿ�;���4�6�]����-�����ˏV����~�b��;r�"�����]p��[�&���M�ju�3�)DMQ���pT]uq���d���~o/�H��\� ns�!�5�Q~�tu����*Y8����܊������iϓv�e'4�����̫ǽC]��'bݛl"�C�2$R���Ȏy����O�>��Suȉ��?+Rhaҝw��h��kT'G1e���)	۾�����.v?�,֧`��)�����O>;���Y�T:�FΞ$��έ���7i���0��P��-n�}K��ȶ���蓸����/=^K��Y�\?E��/�F�y�Kڸ��5��D�X�̛4����	�Jp�9.��;39�I*��{�C��v�@�k��� "�����k ��\�����ş����ch�ZQ M��������������F�E�~�'qH��u�y�a�X-<��w��ҧTRik�y;&9f��V��tVQ*<�>������8Js��cP�I��T�X��Bg_�x5IU7l�Ll�5�h���@�S����������9Z'��mҎ��Ħ!*Cy��g�nv\��Yk&�tAz �&@(P���$��R	��������z�U����T�t5��)� �,c�lVU&�)�-<�ifov��we�;C��
9oD4e�CϠ��T�y~H�F�v�|(�\"���m�q ��A��1�gA��ҿ�M��_qEs�U[8��{���&�\���)��.�$�3{4������\��*/�i���I�E�7oNb�jTUԾ!cV��6�cFt+�v�R�1ܹ�HG���-v'�e��i�V��ꭧ�/��8�85z!uѠ��T��Or�[�Z��&"���/~c��� 2q�;ЊA����a�ٳý��7]:�C1�+��Pn���欓`۸d]Eah`�6�W�Ԗl8�J(�����#�"`��l����3��0�X6��R�-�!� ��@+��h��������m� ��ր�!��nY��r��E��������sO֞.��B��̏��[���=aʃ�^������\d��`�񓠣�T�v�j�����u�Qh�κo���� ����EK���BF�t�sj����C2�tr�#f�&�+,d��ZG[P�`�E��W�@ &�b�*s!U����+
bڅ��z�V���n[`��[����0Ko�z}/���𹅀U�Q�s��mf�Q�3 w���]Tz�ԡ�7��&e]d{D\�t7��L��)���$h2b�Of���;FP�U�$��L��J����q�����K�P�fbq�5�׺ڥ�ǎ�
�j<�mZ�v�� �n.ŵ��F�f�):J�A&ƞ&��z��c����x���K,W2���r7���z�5Ή�as�xK�Oo��(����\�~׮L��i)�xt��,�0Lo�>����ݳk�����^=SM�b�s1�p0��-�oYC�~�Ua��N���ҕJHr�EO���p��]�zE\E�4�C^L\;����r�7gTD�e��~	��#%qa,~w��bR���#[��Kګ
����Śj��2�TǺ��`_H ��dc�>p���+�Ϟ
^(qW��O/-�Ĭ�N�
%-��ӻK�,1��F��bj��!����~����AEM�ꪟ���7ܲY��`GO�o;6���ϗ���� +ʪ��/���x��j�c�B�M��.t�:��"W��\������3B��||G��׬>�;*�oetC�U�)q���I1UL7��\R�mx�6`F���D48�)1�ژO��2����GB�hZEW<�O^R&��\ZR�s��|*���e(�9�o�f�OP@�H_���?��}�H�Ď�B�x��_~V��� �q45�_�ۦ���"m���f�M1*z�>ޝ��j��G�6�A�.�/#ey�T�ް�/&aX�ʝ�?޲�~Y�@y?�.��U�0)�����5�0�́�UY����Z��m��ʑ��ڰ�����̘r^�gz�4����O �y�&�n\
��M�d���'>�U����낮��p�^ѣH��%�P���M���� l"����8�ޗ(�FC`
挷2��ej��71>�ׅ��K7�ɚ �{�����f��o�1y�l�P���]�$�&�dph�Zf;qփ�V���z�3
�VeW�_w@��vwNY�\��$���5��=�A�U]w�4��R4x1�cȮ)��>�@Ơ�:d��Ŋ�N5����#������u�r3��5ؙzJ��w����Y�,�.�2!:S�r�X�8�tg�T/�'���t��7��/xC���C�3�d(>J������ZO�P�?m$�v1��jv��v�&��!��S�Ȅ6�=�|U \D2�.Q*�3�
s?dS������.;����� ����O��R�����bDK�
����/��d�$h�JdIr��59K��vl9��fF���DJ<�f+A�&K���3̷h�y1�$P��=���d����	Bn���\>��~�V�BBC���.��[�'��&/�K�k(��ﱀ��m�w~��Ȓ�BtFTCR������{����	�(T�` �8MD��@��^rI�M�ui�*�8ג�*�C;#���3\�K��\�r��(��c�� �������8��$��ZN"� 3����F��Hū��������_�/�dŲ'#-]���g�9� �7Wȶ�y�M��~-���WvGhn	|�]l�FAK�)P����Ej�lB;�j��Ӊn]�*���z�b��eP��	���lA	��!�W�Q�Y}�4n�b �b�>�m2]�xI5CWUXq"��:�sn������ivk�!{�WY��K�ۻޕ��tۻ�􇀗3��]�V�6۠XV��>�s<2�/�R���#ӌNj� �:]%꓁����,*غKg��专䘲�*���M�q��j\O	��:c�$������!��yԟ�)rлr��c����hOg�\ ������"9�&YuA��v%RU��w�ON���8Հ��T�����<In�)-�9q�Z{�ڨ�ȿ5��@Q*�B�d�9���|�t�΄��l+�K�&��/K95�W�y�hG��gp(zDYU�y�W��/��yK�m7��X�}B�)���㾙���ϠU�����`�B�p�W��T\�=_��U���G��Z�v���!+�PT�gF�]�[��¹<~w�_�T7����)qۣi�Myd���	)�Z���)��EDz��`4X	��Ќ�B6H,7����,��x�|�k�t�!�?��!7P0ll�������/ه�ך���g:���$TU�8+�?�r��D��R�[ 8�5n���?�]E6��IE�,�O�cic̌'Rw�M�t"��3>�>�b7���I����Ƈ�}냲�Q�Ah����1���%;�V���'�t8p�Ys�l-T�u0�;;c�n�1�r�%���H���K��O"Oj�� bZ=�[)��F/�dk#���F� f/�`�Đ��8��Ơ���}.�l�-xi�{�
'��[sh
_f��"9�0�Q�Z�Lv�?��W��者Zm%$ �.�� K�{�}
RXZ!%\|9EԜ��X.a[�����-�u��#\�ʍ�[�SϹU��7�I�f8>d=I�o.�O!d(��{��2���-��3�yM���@ðY5@p���
��ůXlP9\3FV	��h��Zs�;�hÊ&�K��Vi��z�˖�HQ���i�Y���-4�PxJ4�^1��5p@�����'c��h�u��M���K�ޜ�Ya�X��񒻮�����Z��
ࠂ`4X[t��L"��j3u��r��Z�β.��v:��$��s��$Q���C��V{�Q�L!l�i��G��w1���R�Z��m0�2��<���]7>���b�k,k�۹BJ�~�qd}�r�K���d<�L���ܹA���J��R	Y����D ,�?�<���8_�����U�P�r
ا�!	�.OU�"'B���+>�q�]N�!
xǿ��)@N�-<ٺ���ݑDKR1t>�b��i n^@Xk���C��rr����V�br��N�LΔu�����L���n]D�{��=Z��
�}I�A�:u#��)�}i9�ae5�K�M}*�򄐐 v �@1�GX�d����@ �&ה�U7����κ��֦B�ɜ�m�h���(9�/��39�ԹUd:�T�0DfFj����!zy�R���pP=�-eSL�]e;9�&4�Lk2ɷE�;pS�D�����'��4m:��4�������)�I�;�DN��gym*�5��ea�-�]e�5�,s�v��QVc�n��XC)�Cfٙ ^�g��>��� /�~&���H�ƹk"%?9�y�&.#���a��c���\E"�H6C� a�l2z����6���(�Gj���&ùQ���7�L���K-�<!���N�;^�z/M0n�'�@&&�g�_�%u�>��/M�������]�FRjh�:�����G���^ot�۫�)��<俅����A�9!��e;��ƹp/XT}�(A��	Ɓ<q���<qZF ��yX�S$�kVd�KZ���ۨ|����Ρ���H�rF��S��	��d�3F���l�Fˁ/=�g��3cD�,|~�6{�����OޗĦj��X83�6�i֕++�l�rp�|D	Y���J����.o���r-��z���E�h�Tt#rd��jް�б��;�N���&D�S�ǅ5�Iw�&��ו�i�3J~RH9�y�:Jj1���%�@c籀���u��xK���!��;��K^��F�Cⅎ�	L��f�vA��s-ml]N����~Z�"�$�;�I�9�V(���d�2���5���|�fL��S�#S�+�?��(��x���A5�x�`qvRI&c�I\���IwӬð�&�5:�^f�v��0Vps�����#f|�r���Ũ�8s�[�(�_���Kf���"�l~�����.)^�.���~����߲΁Q��ZAq�B>�9lF��r����{�����؀+����q?�]���Zt?`QJ^|r�,��͛G]�i$�Րַk
���*���{��9��10^��R�9p_�$q��
X��Lrz�T߻�K�^㢙Gfl)pF"~�H���	��[F��E=����n��s�p5'P����_��cÒ�	��*���d�3��Se0�%�6�Hb3=���G�����=�Kh��G�umd�-�]-�� �{���vv������k���8<D)����P��K%x�/�;�������]���+�i5�5`��7q���o���Tc��=yu�yð
_��N^��Xе3-�r�ν��,��nË�z�}3�(;�J*����$�tz��	F��Z%�iku��b����-p����k��ڦ4���?��h��g
�2s�B�591"���P�a,����'�LQCq��:��7�����%�wjT`�mZŷ_�icf1iUC'�.��FkPSh������{k��<o��7D���m�Zɝ��ǘ��,�N�׺d�B��]1���"%m�"P��g��k�#F*y���7���|���4EJ8�Ls9 ����J.� ���	��ENC������(|Hj<4�$�5s��S�ܡ#\}�W��uhD�����j\���_���N���ˈp�l�N�������6˿kL��n`q��#��LJ�a�ɡ\��/��OK����j�.������҇���"
T�è	���<����؇X�oW����^4Y����5����v��)J�:�;��̸�զ��vi!�,��iCR%����C����Q�3�6Ø�� ��������z�6桪���b)�OQ��w�,��D����g^ ���8�p��8z��ZjxW�����ުז�D�I.�8�̪J;+k<�#ְUN1�/��JV�@�����1V�����ស��6����}�A�l"��b�B+���T�?C�;`k�7QΊ�$ ��a�i�k��z���������[��Jb ��|h�#$��d� �\�II�U���SGIFaM��v��`��#V"z����n�@�ا{� h�>�.l&[�H�H���հ�EH���>��1z�G�O1;��oZ�(�@�ΗM�"�L�������cP�;�`�b���Σ,�B�	�0���ނ���a+����hI�^\�� 2�����5�x�#Q?U�~�Ļ�d��[�t=2�k�뎖I`��R�����9�'n�-����1�~�^�a䶉p�`~rF�sP_*�=�w�{���S���i.gT�~��Ḗ	�6�$!a�{m�Є���$��v���N��a�����Zolh.
Z�OhK<䄰t���3c���:�Q��4CV���4E��HR��i��
����)�����q�e����� ���ap���#b�{ ���F�&|${�8+����9�K�@i��q�*����J���"�{"_��i���7���YG�e��)c���O����P�%�ufr˙,���O�Nv饗m��<N�K �����h�@�v�{��t�J����T�.)EI+��Y�����Pp
��.нN� ;ʢ����E`+�bô�KT�q�&ª����RE������Z�}.���-�1�h��B��&p�vZ��.�N�|p�S���
�`j�J��c@�|�%p�w'ҋ�;�V��;�\$��-0��ۜTqt��~���6
��Hήv��Ͳ����,6����e�j�x��ߙ�BRm"a�YԿΑ�s���T�*W%ۘcB�!{R���K�k��I�	,f:mT6Nm��Y���𴇝K'"qs�V�� �[��Lk��OP�Z�~6�W�h���Conn�]�N��X�P�W��z��f�W��N��Qa��8�]�=����R��Y=H�w�1���	�Y�_]
sOf�������Oi�/��cD�'6�>~����^h�!(G��>��h�k��H���H?�M;k�,t�T䤻�4lA�<�����U��>T��/����t�&��-Z|�9.�o;�2�f�6U�){��������l��Fy&b�8<��f�\�[!,l�i{�u�����l\N>�{����G��h�����.�~j�X���$kV�� �$�["�s�x'��d����Fs�ͩo�ց���)@�����z�6�!l��\����4��ԭVWe�qB'��:��[Dƴ�K� ^!����l� ��w�)��X��Q-_.��p���|�^�Ր6�s#<[�R���.��jԏtm<�k[����,��Y٭��w9��fH��/L��.�>���4�x͕�4{#�WG㊦��H�>֜[
`�*�Ŵ��<����an�y�y�n���(.�*��ى!u;%䆩W�[��UD�������i+4ADݠlC������'��#a�P����[��QG~Bn��c�&���B����B'��}��K����-�(u�+�>�G��C"�'�h�\�O�/%Z)l81�������ܞm�(�p4�ktwՕ�}�����II�Ɖ�zL�Uj5Ǚ�"/���XҺ�0����L� ]��`�f�$�u�>��G��;����ü�b*gSq.�*��˻߈��,��!s�P*���S�u����2vn�/��~��,�7�aC��3�a���y�HkE��*b�qˬ8N!�B�vk5�T͑�AE�:I�K�=r<��̫�?��؝�?��!�
�6åy��q��6���7��E�ht��􏮫�P�?e�SMo���v�n��\	�ccKe�;}�?�N���>����mX�Ϧt���{�[����5��VE�� (��3�MC���l����ɢb�	UjiLkSRU�~��1�.D�e�t��¤ccGt�����@��c#�p��q��N�j?�*K�U�Q�>��h��c�r�}G�Lw�8���?M>��r�[A�~�U�?Hֲ�f�7w���v��!��8�o[��LU]���G��)�[z������L�i���Z_�lij�β!BJ������3��q{�7CRUI�K*W�j��`h�����ǌ�,�ʠ5�\q�o%4��j�[Tkg.hk��!q�lf̙�r�Sq.и' E��:H�3��2�!��5	�V1e��y0^�湘D�i,�� F_�66�20��B�$�A��v1�[& )<aT� W��a(��i��n�mvJdGx,ȹ���������N8C����_�j� �=% ͳ��*���J��?d�Z�P�B����J�X6/�@�J�n��;)F�a'��$�1zM��P�#�F���Fy5�֍�.���N���r��G�@k��1üg0Lj��SKf܀��*�iwb�i�@'Fk4~�y�qH�7\Y'QW�w���懊7rS�BD��U:�C9֥;R�[ e"W��h�^�$ds*�;���}�)l���,}��ͺW%��Vb[��b9�>�\�)�L�~[ ;��)�R|���E�]"�x\s,��Ѹ���g��08�C��u@y<;Hf��Q�)��� �DWpX�����4?��Tw��V�C��z_UJQ����qU����낭kA_P�����b�1�sɼ\�ly�������a�c�`gs�G=Vq���VC�~��I��G�M5�-]�j;����@%C��H>i�X�����l�>��i��޿<d|UB������rl�1q
O�����;���xJP��M��칄1x�״4mF�a���~��<b(he�U�@�h�?�)�r!�h�-f�*�98V���Ƙ@��g^�rS�#�R�X���f~��-ܖ�T����(�Sëܗ��������۠z��A�F[$��E�	�X��!�Dj�kD���5f(s�Z�j�������a��
$�`d��S���_	���1�]Ж��ֿ�,�I��9`����@�>\a��Ͱ������Υ�m��z���݊�Q��%�7L���M�=M����j��3�d#?���_�[. +(`g���yt�y6g��2�A��r6ۡ4F?\�eJ�Q?�U� �t��M��9�ݥ|��d^���,3���о���R���م�Dܜ}�!3���2�0�?��ܽ>"��y����4��r�B:�˩t�?"��ܷz�U��ecq;���m067�kK���r�h��'��� b�Y��Փ<3�1�)�'.J��Һ��%�!T��W�W�& �{*�"2 ���j� 6�ݡY/��$���C����vy��e�w��-��ȷ��?�{/kԤ3i�s+:�����b�� &f�R�فh���-��}�.v��Aé�P�W'T#�r�VTЉ��pJ3��, ����`���5�����$f�7 T�U�Œ�>��"�P([�'9 z�Z��j�Цih����tUMl0���h\���p�d�fr�ݢ�g�L��>mTB��ډ�`�~Zj�N𵀛J�(���"��$�GgԶ��<���#_S1����X&PẤ�͢���ΖB��LH*u+���f�)u{?~�Me��&[�?e]��������;��jfd��|1Q�-�P�X�K��p?�Il�(c���y����#gV!�\��퐝�
��+%Y�z��ക+1�2
4�&�X�Iz�{��х��*!'�[$!~Bmπ6��ܶb�U�o~I�51D#v{�O�c�|�y'Y0C��+��:�
_��^j�Y+K. �7D:�A#��4�N��q��k�>t>��� �jƕr��'S�S��H��O ��ɦ6���J߱.M�����u��Ho��gm�S@I+zA�Z��pM+�G��LVv��Ma���J�/���?�%�P
B�>�?;Z�J����u�oH�7��-fp� ʭ�����ތ�}��E�`R�!���!p��s��aj��׹�G��F�g�y,�-2��S�h\�Fp>Q(]rD�U!��r;N7��1v�Fj.;W�h���r�l���ka��A�&�dn�-��ݖK nI�QS1f�!�x!�bu� �2�q���Ɗi�y�TJe,�Ĩ�F��9z��C�?����1חF"�w���$�E8�T��6Ԅ�;��|�:��u�� �fN�A��{P���E��[�	�Z����zj֪-���+�����eEUP`#H��$D������}2�ч�59��ڹ[x0�����(� �]���6��)���P�\ʫbU����-)X�)�հ,��_��7P.e�����2�U���v�S):�q���Z3 �v)2�ͣMgP7|��dfL����x2��4�F���{/�D��͏u���S8��\&H>�=���PΡT��n��{�_�d;����y���u�@�D��j6 �ͦ~c�=hY]]|U~�Ǐ��|\��D;-kFk$ʌ��=��j�@�(	)`=���F��qh�Way��Z�*�k���ycU{���hJ둊�����.�K!&J;hP�%Xn�^zB������Ɯ�ĭ��>e������Qn�^|��=���.�b2(fP�b(i�q��6 D1%~Q�h��j�B�����c�2t[0�4R(�nɩ�X$H;�El�T�g#N�DD�GTzHQ���+�D������x	�����u�\�w��~�<�c��f�1H��7�/\�+���`)���U���K�ٟ7�QH'}og�gu��ܘ���
�#O�U�1�A�V�=H�h�N�o�o�;O�w��t~d'�h�=v^�}���q"���?�!Z���z��5�Oo��ڢ��O�Mq�kд��M�M.Ob��_"-��t��W?����e������CI����!̯�,_Ҟ�On&��$.���PWu�j�P2�����������$��Z_�P���B_T}����nD���m�h_@&�ZR��)��Ȑ.�mS�a֟:�-�����+
[�������b�<�yS�C�Ss��PJNt�I��&�-�Z&t{]9�d�Ǩ����[ %ǘ�1��.@����Y�������9v�2\O�X ����nţ�ay�Qҽm��Ԙ
Q��ѡ��r˴F-E{��t��3E)~= �Ӻe��y.���/jN�G�KS�����A�&���V����^�Q�s�.���Le��շy�7��r����be��g�O���&Pj>�L���=)�m�xlTtx����|��!r�U�+9V��Qp=C^#94ʝ�r,��d%݅�9OK�O��Y�-�q�ex�~.3�@���~�9�'�J�74��4���h++kϦp����b����o��qoo�9�	lM�����=D����� 2s�L �f`��J�zZ��̅뮏IYפ7�U��%�Sp��M�0`�~��ѽh
پØm�(%�����SGz`D�H�������ɝ��[ӆ�-��|Ҹ�"-N|a���xㄜ�vP`��	Uk+�}3Ē]r�)�iN��d7��J-���{�5 p�I�kS�d+5�:����)���tn���[��M{`a�ѓ�9W�@��b?�E�:�;ٲ,eq���/,E��"��%��/!^k��5	do�m'�`dJyk�#��J"Al���ءkW�
�}��l\�DI��h�-���&���Y�Du.|��Y�a:k7���I����,i�I��;�9������+���'r�� ���Y�,���0�#������),1�g]�.�o������Y���lSB���G�p�(:�=�d����3�U�����.��ډ�R��l�*��}q2c&k=�d�7�t-�Ц'�����WŁ���{������ͦ��,�����0�R����5*����8z�7Q ����O�\{�Ȋ��ptq�"����������Sp�aC_� /�qX��,#^�����oz�)#�&��0��]�`��������m�k�P>>T;�-�C�)�� �hr琭�M�w��L��t��_Mټc�Φ����%�C�C6k�rd������+�ΨṎ=�\��dw�H���-�Rk2�0ږUܚ��5{ٔ��7�,N���M)�Ϧ`��0F<7�MWk�JA�Fa�4��5r�_J��l�Yp��wT��A��%�D
:�Fl��h)��A�����������`�A+���R�����_jƊ��f��WElݛ�Ru��<l�䗠zI�h��^���M
eT:�5��Z���&,4,����^��r[�~��??����p<s\����H��Pwtd�n9��}D�V��I+�s�a��C%�(a����'�
�)�Y�;�MS����!�W�hf��pO2�틀���8J�"ݑ��p�+jٵRU��*6g5:_��m<�ʫO�����+�=��,z�ꒈ1t=�$W�eLF��f���_�I0���[j$��x�*�cܫ��N�z�G~'�O�	\��v����$z~�Ґ�\9O��2�"���13���b�K�_\13�%���ݧ���I-��ͮ�z��H�2A^4�q���SϺ�y��2������Ʀ�d��dZq�VI_9,Q���QlExޙ�ҋXOK)O
�KT��'N��уCL`�*�/���J����mV�����ς��1�)Zzw�v�)؂GZ��J������}�y�Yķ�&%��}Y��ک9Ud
����|a�Yޮ�<�R{��H�1��$c��5SJ�'/�#LA]� �ؼA�`[\�O��	N+�����p��v�^Ecl33���A>�b�-h?)Q�Es7�����E�suǜ�����J��-��_���e�#;vz�2�q�痣�¡D"�Y&~�)�7w�QD|W�^��~��9W��9C��>�c�����2��� V���&sf�.A-�>p`�V�<sث�y:�:���2ל#��:j*Ҭ��DƖ��j�E��?����F�5���Ņd�i��+U����x��9����� F�sf�acf�_O_ܡ���i�S�΢�G�����
�.���Z�q�h��p5��Fghg�g%]}L�w�G��S�;�S�b�馏/Y�ề��\7a��7uhK������0���.�F)�A&��~��c�A[�\REE�n��=e܇K�i�b��!^_�6�)>a�)���t_�i�u�ב8ȝ4
=�H[ly~<KYy��7�"O�x����|G�ar�Qk�]�!��|��Y���=�&@��=Vu�xj���I4+�Y�X����傪�-��AA��&�dJky�е���I�d��I;�	G� �;U�`�y�#�ʂՋ��,:��ww��>u��x{��mb�4�!����H�|��Z��ò/?�����NM`�g�E����b��;�]8���ݓ��_�<Qa=�ϼ~�|�����<���B��5Jr�SR��=,�<�wؗ�(3����{���1�/�i�c)<Ԇ��1�'v`��Ȫ�~sV�)ȉ�|Xo��s5Ѣu�x�Д�7��DRxϱ�UM���-,2�J�i�y�hP���o������'RK*G�5{x���.3om0��N��A]ǯ�d�8��Ujt�2�E�g4#�V4k��j=4r{ۍ.�f�׶�����M�YDpa!�Ft Ҳ>������-���&��͹0J"2NK�0��N/��f��Ύ�>}�A,�?�vډ�
����"swO�%}�&�*�2��tFY��s�P#3dbKk���sz��5T��Qmi���w��Aj�z,�v;���#&>���a�z|����v�����
H�?��@�N�.)��/,�E�8�[ύ~�kA��:~�Pia�_�#&�}�PK� P*�o*�j�����=��k���R����n���	�"��Cx�Q�4���Ɠ�â��.h�c>���՞d�,I�,��6bk�-�D�C�1
�Ҟ��sTa\�ꮷ����ͨ�VK�����o!r_��ne�!ԚB�3��H@�@%Qn'�8�m���o&Rp�Lq-�P�������`9h��z������/o�{j���p�δ��|D��ו��ޜ�6uQ����Nf�L*nd��C@��A�[b�1�M�3I.��Ha�����ʠ����d�Df���z��R�U����=��t�O-{0�͆��� -^F�����|#�:�M�+ԍT����T��h��9���xj2�Sn�,�4Yv�s ��]1>eA6�N���c�d��4|�ݬXVɸB��Ea nOn.=�����~�+�	���r�i=���\�d�^�����X�U*E�.�*���C�^�Sxr:e�V��;Ջ|�՚����`��������R��¶)
Kz�x���:�f�O�Oi��E��2���ߊ(�0@�
<_��7�ڳ�o9
y��qLN$YC�X|�ݚ6j�L����+0B�["���τFSzv����m�˃�y����h��[�fM�-N}����7h����3�Ȑjd�K��_֤H�Pb�Q-�ਓ+�N�NL�q&j[7�٭1�G�zpqM.ʺ��A{3D���4��e��@Y����o�Κ1w���g"�`%_�\��r/���4�I�hi�5�^;�I��*.�&p|� 7X�
l2��PF�P�e3�]���=
�h���Z��f��i
�|Ƭ�e�٥��_�q�W��ě-��-��U�����׺��-����.�lLVz��܄�ieKF�g���/�/!yC/j�#3�~��nQ"թ9��|�wC�&�!�D<�a�6N��I3Q�h�04��N�w�daK�Rya+���%�'`Q��ȷ!��S�o^kX���(�L��qѬ3�^��9�[�-�`���Zi�N����ew��#���3!��k�f�$�4���̪Ѫ
g�3��GA���7�X<��i�S$d������O H��s����&��TK�u�F�𸓵��V��CA�9�)��Yj(^<��\�0Y��s�\���$ wZT��R<�Ԓ�ޘƤsP:��{7"�6*�`0�D �r����6�XtH��$���}M��"$�3b�|�Oj��tՉ����b?�Z6�(א���,��n������X1!����# h߅�&{%�p}�A:����!��v]bR��lq2-IV��q�җw�������OU��;���> ߿`;�g�[��r�rp��!LY�R�L�8�uü	���K93�u,ૼ=���s�O[�V[�!8Y����&��Fȁ�~�/f��S��Z*[b��O��ȫʕ@�1����yq`���NT�!�o�Y��p<Ȯ�.��t׃�ER�v�;����D$���e-+Nǟ���P��԰c�����;��@t�7���1|ʳV;�cpѲiz���
�� �U0E��1�>	#g��?�zR�yk{�cP?�W�S��襨��:�<D�J��&��Č�X/3o=���\ֱ��6�-����	��T�PE&�1o«�89�S�yt��ŀr3��	"�����R�	�rx*)�p��>�o<��k�HI��\�C唐�l���Ry?A�I��A���`�
���Ю��'Xz��
�M��HQ���=�i�Wn�q���S���UL�U%�4��zޡ���BP'��{��͂��?����A�Cy�{��h'��*`�$NKW(�h]%�(����2�n��vF�O�j)~H\B0˩
�P\p
%���t���x�;	�;v��ɗ�#���7U�����=������*���1�(�3�����F���c����K@ �c����e%&���$T.ZE^��뵦���~��KF,+��J��oU��e��_��tf�� [p�n�\Ęaܫ��ߠ�mK��qN��L����9X�+Ei�?��u{P�+4��}0G�&*M��=�09��b�c"��/
���C]�6�-=
\2¬��U����ܢ�=��!�qɱ����{��r�3���w1 �;�J́��uB�(y5�����P�>�]Y��P�E�hY���D,ks���]�����DȶF�_��(?-s!n�jM��'���˰;!����/[-�m?vd�Wԛ::F����as���������H����]�� ��&:"���\����hd!���]\���1d����ՠ�}����@�sm�1_� S6Ӊ��G"0��g�	K%�߿
��/vڝlz�m�Jo��8��#���;���Yq#ig�ae�4��F�CY>5z���~*�MGT��|;ܻ��d���(T��87Z�h�,����x�Vϑ�����->��qy�D�]���%
�r`���CI�"�U.s*f�øڦb��4
��_x���=iH�u�>F�'DY�*_8tA���rM��#�K���t�h�:��תd_`C�^L�\YL��Y�f�����ęi�{\�VK��jv�����t]��zB�zgS�q��UCn%����9�,9��S<e�CL��(^�Lw��ߺ�B�T�"�*M��ɸ�TAn��ܘ#cH��v$�ň&h;~ j�� #f�z����#��@�<w���q�đÈd]�fh���2ɍ�X->׭=�-P�0�QN���"�����Xp	��Ċ�
�۵���릓�"7L��Af-�N�V��V���?ˠ�����]Eз6l`/��	/":��\���(�q��,�W��ۤ��_���!�Zi��r(]�6��v���e�m�>��Auc�S��A�h,ĊX.�}�i1�۞��B��W1ϘᇠC��֩k$q��㋐�����)/�Ӓ8�GE$�Ҟ��`�o�Ip&�vp�6L��{��$��`���K�x>�;�z����l	�O���y��J�p��i]���Jiz���uX��j%��4��g�Ĩ�է4:��F������L���h�b9����Ψ1� ��F��V§�R����S$>��q%��|G�O��CaX�KZl�r~��u����&���:�K'�_����t7�^�&E�[`�Js�J[UI����L�7��AW�]��{�hA�NP*]R��h(J}��惢�}'j��&�������W3Kp!�~��.�#R����o��-g�y8���G'(>�'H�1�Ʋ*T.�NDuT�2�_�R�1��n:��i��yskG�!��D�H��I�T�*Q�����7+�#��H�nM�0�9^҅�,��-t d��&���WF6�������_I K� ����G�	5^���Qr��ȚtR��F!W®��H!�FJFУ�o�*Z�n3DB��&��o�G0�nH���am�������$$��H��'q�(�C�S�ynI���d���kGr�f?�6� GG�3���u����`�CW�Q��%��ȃF�Qy��T�%�=ۊF��K��=mHH�9�N��@�N|�rۡƂ@��%yY; +ʻ\�Φ�`ϓRr�������w{u~�^��}�ɘw����o�T�ޫ��b>��7��]�fvmFg�nd>w�A���9�;]x&uKP��Q��D���[�5�� 3���Ltz���oB6Q�t��""\�?9�AV�`Pp�Sm�rt��0h�,�_�v�1X�m&���ӴV$�X�����@/���{�w!c�c
� ��x���<���t��m=v�N�<S)�k9}�G��)=�~��%#��ā�Y!��o�e��B�%���}s^vK$w��>X��G�WX�T�ԨZ�̋W}f�VWd{l"���-�Pm��}'A�'�]w�-J"^�3q����_��L�|S��"Q���\���Bp=t�d���͹2�;��=��U1�c��tŜ�I�mh�����o"�;����$�䙋�~iy !��'lS���~Ty⪾̠�J�p���?�)������R��U�k�_c�M�#Jw!1��mɦ�/ y�;�.^�w�3�޶/Sw���4�-ęD�1+_2k����ʏU&J�����m$~ �R�߀�_�`�E`���/qZq8�vV�ly�mj��-��[o�q&�B���ۙ��W�K�?\~�?Rc��/^��[���v��|~�� �s0aw�Mo�]�c�1 s:�mՀGO`׽�B��)F�z����f�I��5�C�iR`�ۥl蜧h�x��:��p�U$0>�R��U�`�{�p�9!-��P?U�K}Y�2�Gw,M>a>��E�KR���������L#ǁ������!�b�OB�1ΰ�����<ܿ��Z>�Q�_��4W[ �u�U.%����D����Wz�f}�(���2|��ĉ1��͵Z��/G�)�����P{��z[�>���*�Ŝ�>�&����ϱ`�<��T;�t��F�mzm�\d�������{v�Z�É'�k-���Z,)n��r�+��X��QDW��AO=������s��v)���xHJ*���@����1�}�r�"���9�/|�=�cbg0�'�⋪񅏕�'x� y=�,�q���ڲym[3p_
�Ո؆,��M�K��Z��%A�i|EZ��:Qޘ\��� l���
���a(�]���&Z��Oh٪��C�=Kx9�JQJr8�H+�\#��8�r�&j�I������9��U̳�vRYsx�<$�J�W��p��Nx��R9 �����x�نW���W
|��>yk�y<�
�A:�����g�b�9ԟ�)��>
X����f*7�vt[�ү�m�k�+^�{l�쎖�F��h:�'/��nh폿H-J=��Y����?�ߗ�+z
��/�g�O��S��>c��4�Kt<)X�BWK��X-��7j���*�q��ſ`5E�B/ı�#/��xW�Z��yڂY���&; �����Z�cn.%-kN�GQ\����K�+EMp�JD\Tp����eUq:��,7�>�m�zL'F^�y4l�Nހr� ط�6(����]����ť~_#@����k���^��`�.�)T޵	 �-��F�@驵:1��5i�A/V���N�di�Xܢ+�9S�e�V(=1�P��I!�`�B�w�M9��w�ב�8��~�+H){���A����$[Kp�GV\��]�*�F�@q��bU픙ǅ�L��9~ R�R��~�He
q�,�	Q�Z��S3�J���m�2�P��?���Q� �T����Q��2B�'{����C��܍&*>���ܒ������{�v�r`@�.k����-����T��T�Wd% ���a�p���W��s$��U�֔k֎%����Bs�C��Zf�6Q�l6I�f
�~�)����I�T��&EL�	~HH݈z� ��G���3���D(��t�Wv<}�hU3�$����J�^��u:�� <#!c�!c�����Pq�����T���H����T���3?�Y��ՁLD��B��|�\F.�ڱ ���"��Zpz�kϣ�)Z�y���j��f��&��a�V;�.r������Z�*mL?!��Z�Z�kE� � x�+I۴&� #R |���!ѳ�β�~�2�UUa�2��	B�����@�M��ף�F�i�C�}����\6�d����,s0]�""/�pSQ4N��~g�n����
b��q�B�1��Qǉ�M�缬MI�t�����hSIwr���1K${���8�U�@������G0�/��	�@d{�Y[�1Z/۹;�r�ˋM+���I������ed0ҩш�?�g����P��ΟX�\ܜ�*���գ�t��V�DP�=&����.l�uH�*yeU�򕛓��"�n��-S�r �R�e[.��b��ϸ+R[�E)�h�r h���L���\[m4�s������ZOR7+�n>Q�Ŧ1 o�`˂aACV���(HFe������Fӥ�$�7�w�#֙
Ի7�'���9��آaSOO+�P��TMr�D�&�/(uq�bʏ[�����(�S����⥯j��N�}�S��a�ʍݸtB8��pM��I�K8�JM�$��:��bCk~=뀇��gR���r��aUl��N��fwe�!+�
=Xa��U~p����.a���Eau�$g�#+�=�(�� `�^9 ������B ѼJM�{#yT8���G|:q�!����#��G�j�聰��͖'�Z�?�$��X�N�$���#��$W�wm���"�!�*����Z,$���6pIǷK�}Շ ����V�#�z��H;Mbr�d��B���4CC�7�0�?�߫_��2��mK[5j��9b�)��ev%� �G��_u�6����O�4��V�܄�fjb@�š{�"ݕ*��+9��|J���S�<�>N�W�a�V���+�D�>R���wn��c�����n��L�~u�zl쵞��q��g�^����d��%���5÷YE�Zˀ�`�̲h�'��ឳ(aj������Y�׿�t�Ƙ);���c��ɑ�Hzʳy]VISi��,�S,�
,��HE?�,�nH�/�!�2�J:J�]	��~��.�n�[��?��u��1�1��c��k<�z�W���ˍ�h1(�}D���G�����x �����e�/�
���[(O��C&A�6k������h���\#�r�{ǘO�����p�D���;�o�;�M��`�^$��覽]@�ƛ��IFj��@���$��������1����l��uY��8� ���w�����T�H�B
tr��)zn4w�j�Xɟ{�uW$.��qǖE	k�y��8A�b��k���,��W��eXn�Mݮ������	��y��F���)����'�󰵙����ͺ�Ik�;��������&�X�A�f��@i,��!���:m_�w��G�g,C��`@���El��r�Q�`� S�ΔY%�{������Վ�����_
X�Hh�]O "�Z�ء�f�a�E�l�_��r�F����<�T�a�.,�����%d�kF���5s�t��^� !H�����)�9!F��4�&�M:\�>]uuP���~�$q��Ï����t��C���.F�x�?�ni3$�'��m�Օa/V�+)��Ym��B��Ý�x�V�K'>�i;媰��D�Z֪�����Q�/uG-M�I�7�Z<����k }ע)�����C�^?!SӪY����!?��1'�K�|Pty�dQ�J����l�����2�5�U��4�	(%^��b`#P
�Y����U��y�K��f��F�'�(Β���z#�]�p�m��@:��,���S��S8X�&�
y����&��hI��G1i�@m�U���BY�����ab��t����K���$����n�f�R{�
y]�Y>�ӱK|x����8ڃ�Q���cP-�8=��ki�I���س�ce�-*Xd���/��=Bp5��t�:RQ�i�Y�h2e�=�H�%M��ZL�ך�ǨE<{��Kh��#���c�����W���gg���em6���u
7��ӵ=����ϑ���]{��҃^a��+�]�G�@���l
!�ԫ����"�0�֜>=)^w� �/9���+&�b��re5/� ��%�З'E:,�ScL&V҉��G�H~#�F������6� ��[�@lxB
&�sGA<�ڜ���*J��aII��~C��Da���F�oj��}rz҈��1k|?m�`n݃'��6���H�9T�}����G��ѧ���P���梙�~ �H�n��)�"�s��؎�e�O�I������@�ι_��7��X̓^#�q���d�.7�Tȿ�\'�������|h��9�S8}�`��8%k��S<��ׂı��o��R�1��u�5�.o���I�&Uȏ;��A��V�`�F�6��.T2\��"��.4Y�����%��ө��4�vl� �p�(#��O��J\�5���Fw�ki ���D�J��WDS%�������Z���z ��$b���Uz�D�`���|�Ҏ�_�ZCƿDD�\�vX�b> ������X��6�/bK��.�A�tF��t�j(�nζ|#�UQ�J���?�'W\�@@i��0_LD��fI��$v���	n֮=L���c�9,<{P��R�Ju��k�V�gm�nLU�DN۩����c�(5Kvֲz _�4xխŲ��p�:��K�|���o�"�jc��IQ�^�x`�|/ ��?�;V$&�0*=��1�م��?4&����g��	X(�_V�Yr1?砾����:5 FW҆Y��u�4�/I�p�h�Wb~W��A��4
�C2��t(�H�!�p�`�{�CA�A0�8u��]��;�TM��;���MD���{�����[P_�)�n>IL�ӛ"٦=P��ʨ)��pN<�iQ7�)��)E\�	
����t�N܉�MO�:���
Y��B���Xb�z>ڡ�����k�#j�D.~�`��L���:�܆�l`/b�})7�K@)ӏFv�o�ok܁v\(H(�J��"�K�H$˼�l�Rl��w��*6�q�+D �A฻����S�Sw��*�f�x��oa<�3�&Q f�����:O�J�
v��u��.�h� y� ]oeօK<I��1Oj��#�V�q*q�i)ڣ�9��ݶ#�Cz�ϔ�2?����+�d�v�����6qz'{y�{Cˡ�l4q5_ܪ�԰�m��}r��rY���Wgd�v�Z1/��B"o0לp�x�	YU3��e�,˻��k#9���Y�o<�.eK�@�ǖ
�M~{���%��^��Dn)��<�b`��N�;3��{���4�K�C�4Wu?���u��IY	�W������h4G�j7XPQ�ŜLfGz���Y�˰Lֺa>��Ō����#�����Q�H6,����8�G��O:�V%=��>�'�C֒px/�����K��e͍bL\�U���W�r�_�6�X�'�|nZ�*������Lk����
�ht$��bݘ��QbN��r{��9�E�Q����{3��ь$^y+��2��U�ǁ�����9�x�4A%pE�����:^���w���z��)*���,��n����.����ax'��ߖ�|��)��8�FR��=,dM��|��U�`��K��OM#�z��*i%���HV�?K�����6��bx.#ֽ(��J���u^��S��{�:�k=��|�;d�^��X}a0�����9�����	��˨�R�L��k�/��eK׭(��	��ӈ�: Սc:�U�~wҝ�u�i-��/�����>���>����l���Z��)�wf��TA1�zO���b�b�@H�j�L�<��fh�Ų�^G('��l�t��۵f�(I a=l)��K���4�o�,\K;٥N�|P5|��,�,9霧����~i��xO�c�
͈e�a&m���a^��R��fe �@��J��x\`\�L�b/R]ٚ���ݽN�LS�}n���t�����9Q!P��Rk!��W�����7­�����<��cYD�d`ض��4L���ľ�oPD�����"r^V�,1����,�"*��U���S��E����kV[�7ۻ8~!�^:38Cw��{���8��<��*T���a�G~!�%A;ͷ�њ	�oy���M�P�-��8��X5�$�L�{9qt�@O1��;=�`��038b|s�$6$���a6';)_�{	=P/Lm�K���(�W�8��i*�s�"y�]��9�NF�U��zڳ����hC��f?O��XF;rU�� �[���<p�7q��o�[�j�2K>1���»�d3�l��(]�4F����
N�MnKˬ
�`��Y1
���9�Q�Lx��
��ΎSĝ0���ڄ����`��oެ��QU����� X���}��n�����p�%t��h�(�G*z5@�rŃ�˙���Oc'�0F�c\��Zfw �	�$�ه���04t����ʝ̱���Ւ%��y�{4T�B�fy����ʜŁ����*�n<ig]�]�����x�nC�.��q��Ziq)F	�:��������S��E�o���Qy.ӼǙ~�`OVi���6ԓ&iov�p��Գ�R_0�8���I�c��aY�'zFށf2��|�)}ս�1�,�NyB��*�ㅊ)�C�E�m���Z�FQn#I9(��Q	�����h���U���@	�_$�\�g�dTC"�J[� u+fK p���=�:��{2�?z�}�-��6�r��J�x+C;��\�!?n48>�>�nHZ㳬#iӅ�/���3d@"=ƨ+�%rǞ�ks6�W���w=\�p?n���g{�����Q���Q�X�7>�����O���'Y�<� �D�/���"��z����t>W�Y��
w+ZD���1K/'�H: ��۔�4MѢ�T?��lU���	��I�K� �U�\���y#�Vv�PL�a$5���Ä��&b��O�q���mĄ!4��S�������X�Ժw����pA�!$�:�y�m�)��-��?#OΚ������7�M���ͷ�>�r򟍢I'���k����R�L1����b~}b����u�>b�G��@!ZB�,��7��%�-�m���Mz�Q�~G����@ճU�:�g0a�?&�M�������~dH �z�uq�<qEWx@A+���c�JCη��[ћ3*���
�Ǆ�9d��,�`���b����W_�t1
��w{"E$��@����@�V#X�g�	�o
l�i���#��)�}�����+,���z:�7Ke��S3�u;<%�D����8|{�Z���oxM�-\HмҊQ����M�Sg��H�x�Y��3n�<<��L��bU�K�t�)�'�U�H���o�l��]���������Hp�n���ǯ`�Y�����GH&���9�N���Eެ���K�[�=� �����U#8�����,d��[�eqsG����1y��w���9�1��Y���)ܐO�B�Y��D�(<�R��CɊr�e�L���@�ꛯ�����Z0d��J��C�@8sR��x��.�4A��P�Q�i^���C�ްI��J`߱�ԲށUg7񔘥�L�������w�������Wb�������#\02�� ����ӽB���v��v�F(ߴxm
x��id���H���/V\6"����293#���`���ZW=�������0S�#؋������?\��ݴU�q�%�@�K�V�栦|f�����-�j���hU=���d�����{���,(��zu&�����Eu����Q���.>�Әj���7��.��D�(��s�B�%0�b�&dTcEՊp�>���5}�HD�;U���i�5�k��`℈_j���1����Jt3��cĆ۬8�v@V~VÆWa�n*�1�o�
h0X�j���̭�:~���)K����1�F,cV������1�}�տy�kOPLW�?iHq���%�Y������m,Mz �`T _od�7�}w���$h\�=�rb :�߿�p�#∖�R}
�ֈf�v�v���T�ZG)\�[��n7�k��D�%#��cF>5^07�Y�:��k����P�y��� z�Ԣ{3�,��%J�j���k�L��"E<��[�N�+��r�匑F}
��#�ŝ��,Z�$���.|��/��1�U�6�"[����#uQ�� މ,O�����ܝُBR]�'k�;�F C=+��2�o��2��׊8��:�k�plE���N1Y}��>�}��6�M�kgH{���IL���{�rI�?�K�>��h@|pl7| �q����u2@"L`2��
����Ba��OUW^�IG�p�� ����E�N#��^�ˁ�����Α������LH�I�!#�C:E�@1�Y)��)o� 	IA��𪟲�
��)��\_�bvd	C���EZw�R���>|*��4���8&�����s�,���ْ."N,/I8����9�#<����f[1�5� ���~�^��\{N� ���tdn�~T_�<ݽz�6� vɬ�D-ha�� �r"�n� �97�m/��2�P&f��dF[Q�5O�*|�Z<i<�pt�e��
l��=�Zc�	l�F���	nU�1.�C�J�7F:V|(|jj<-�.MR\"ʋ���O�9H�2	5f��vvvIB5�xT���?>~XQ�mFT����sчQ�ơ�+���^i����X�����h�nI\��rp,l{�?^���N�t���^&NQ�ӈժ{ ������;'��}��yzݗ�z	�����w��I
3A4je��MGBX2<��nAw�H��a_�X[xŚ�����?��13@;'}u��%��y��h-�j:!�̳1:_�:��z���<b�I}��[h9�hmd�Α�+�h����7A���d@���f�?f�n�i~�j;lQ0�E��w����]W��Tk����D/�ϨV��	��ifA�<��uE?R�Bl�ܔ�=�x��M�)S��ii�G� �%I�І@�J��2��6D��G����!�Ĝz�s�����z�\�ut��uU���s����E0���)-ч�y���C��Y]B�钊�6�e�Jv!_4�EV����{�2��C�;���f�1;a�F�U0G�$�U ̓�:To1�����9�I�S7����]8{�`�k�&���ȃ�G�Y�OIj���K�}�������9�fiA�_�W��N��`��*Ȼ���1�n�5 d��Q蘨��&Gd(|�Ja ��`��Qb��g>��!��:Y帜l�c�٢��O����A��-�|;��ᷩ�{�_��t�IG6�?����]b�#��)�
<�4����0$�>5�����a��DPd
��e�O����a3{��gu�|��s���*��w��j�ِ ���s� H޲X�"�!9��TF]i�T���0y3V_Ӯ�9�M?N�qG+�����f�x�w;�(=��ؙ��|by:�L8��!꾍��q���1c٩�+���^"��d��)^JT�!^xm*1�cU�NT0,�o3���Inߥ5���`�`�&zD����2�����I��I{�2��e�a}��-kņ�{1j�zN�F����_Q����}w�� 6ؿ,˅;�|�9���@�Q1B�;�\�����ͼ�cw�w��^�۵	㑣T�L�	�6����تZ��ޜ1�N�KW�y�Q=���w�h�W�	�rP'}5�Ej�>5hd��zڹ�sj�-@o��B�i].83h��*	Lh�a;`
���L��/����d�̽r�nfz�3d)���@�x3��Ֆ�"���)Uˢ��	+���h��F&�ȑ�C'BL=�݄x嵖G]%^͆L�#D�Վ�u8�U>U�Ń���y����w�X�m��*\l�8�`�����K�s� `v�&���9���<�8TQ���[҉패���f��T��J����J?Ñ9,�4Z�x[�"���N�[j��>���u�iB[҈ v��"�`���0н��ޞY�}gĄ7���i��X�e>B��H����Z}cU��4�,��_c�Q���ތ�[��Y�C�����'��Ѕ2�Y3�g�I�T�K6���-��wȴ�E���ayT���H�gR&�P����M��n�*�ءq~�D(I �����]�R5����ǀ���'L.g�.X��1L0�<q��e	5R�Ʃ�(����k_<J�f�����:^
Ϫ��iU.���A�����i�	#�vTݓsyu�m�Y�8}���E�x�>!��6o��c��NK�r޶��8�9��=�i���D������o���͸�$�ӐM��)�� 8�+�N���aX~r�#nI��s�,���jmt��Hd���kb[%�)�G�nA���f�-��.����dckj�,�)�Df̔�-�;�$9e�q~ˡp��#5�"`��atD�*��8��U�SӜ�����ʴEmc��D�=r*��`߽hf���Q^+��P�ݟ8њ
��Q�8����<�]*�ȸJ��I���So�D�<��������-]rE����a?��+8��.����9<�f������h��P����U���o�	�0dZZ4��b�%!�'�>~8�"�r!9�tcE��
_:�ؚ��w�
�]&���ŋ��M��'���]�P �'o��8��>�w�Q�~�)�&�p�/�91q_�j	���]j��b'�
1�[~�0	�����13�˯�x\<��_Ԧ�$�5���Ī��/Ҵ��ٱY����'r�'�5�Hk1r�vBND~�c�����Ö���I�����9¨/�X���c:Y�W�ine�����/(�K�CLx����Q��_Վ1ݜ�_��!�d�1W��:�n�u�14��F0V>\m�ޤk�Xq��nBAj{=s�l뽾i+�������(�ER������f+�j�z[;.�/���H����J(�N��S�]Z{t�zl{��v���m<!�I���ru�Q��x̙9Q��x8$�	(�N��}�%LƩ�fvOť�|m�$��j����3�*_��Z���x���*��}���5��e%�*�����H8���.���(�}j�|+��_H@��5��%�z;�M9�ۆ�;��P�(1˰&ߊP��~�_Ҍ߻���ܞxT������dlk\
w���F�^܍�k�;����N^����8s�^�V8��_�A�}���du�P2FA��N�MVO�"uٰn�
��{(=zN�q2��Β�o*��d$�����UQϐ�*��$<z�rM[����萳�U�!?˫����U絖�]���s?5"E��2������ʄ�qd"7:��Q½�QL�~��졓xy�~A�"]��*�!5l�n(�?�}?�2�����OI��Q���M>^�#w�����퐐p�to�tt�g�1Id\�,aO��:�t��/��s��{�+����v#�Y56-DFa��h$3����	����wy2 v���l���?P�Q��W��ZPB�7L<���V�Y�^�-Wo�S��w�M5�Z��Zʗ�DTh)d�,�AL��WO���k"��Q1�D5IQl7�	�62�#��Շ�V=Lf�N����X+���$e�-yx�Ѱ��gQ�)�3+�~J��%�uy��$��X�P�����?�V��(r#��DD�'����N[ML�X� ��`���~��^�EJ�ѧ=�]WC��d�μ�y2|�>gy��S��*�ن�L\��&�z_!����3�.�H0ȿ>�T�&����r^V���`Ym�x�]WM�(* `��3����g ��I�O��A[�#�*���;HnW'�V�z@Օ�����CP��|��WUQ�b�����z�t���	��/���.�S#4��ĕ��L�0+���#��Hm�
V���,(�$��'�`�ywt�Νx�D,�s~&�� ��@�)���u\�32�0;��Br��9�#���i��ozDJ��O�ۊ�%�U�a�FR�ذv&<��LŘ��KB��2^����Aء"�=�VTb;��e?�*5���U15_��L������>8��<�q&�)~�C��Z��� �����  *��Q�<c�H9��,�~0�4�y�?�ı�=�~˺��.iN2����a���̬x[�����yV��}G�|V�������p Ea���'��y��zsX�w0޸����ۺ�"�Vq3iw�h��87�ht�b^��x2H�Lc�g��{k�B���0!�gq�l��s��������{��\��q����R���;ו�e���w�n�@�ّPM��@-M^����\L�������
��,�ʤ7bV��ܩ�Pgm���� ��J�5��g OΎ}f���I�ۓ�>�H���a6�n��o�u{ �Dуx�GQ��В���L2f�}N�uC�OU�>7�>�W��;u��tK={��81l'�#X[۾�[сj�_~���SC���G4�mW��Q�w��Y��@�R��An��D�3[�O3n��t}�T��E萖x��M>�ɐ�z��ڒ��yvvK�	@D�"�Hk������^��ֿKد��Qu�n��?V��,JY���Pu���&�{fñ���EQ'j��\��H9k.�`�+���]J=���(� wЎ�㋷?,!���5�<�a$X|B�^\�jG��̹1��٤�.ϡBke�>(�/a^(u�H&F@���d@9�D������l�7��J��Q���L_d�;�j4�o�&���;r.��h��N!p���h��Y W?U�ǍGڕ̔��qg���z��ZZlsl���P�/����|�5u4��W�^��)P`H��#�(�=�ܦ�H�\��d(�_�+T�?�������\�u,q����u����x�߬y�ƻ3���(��8"�Ye�%�)�F�6�Si�JE�����+
&��Z��� =�� �Jp��@���];PL�@��u�*Td�p��ڥ�g8,KN��L���f9$�n��}�?��� �u\�TF�C���d���B)� �1SD�ϝ�nH8T\۸Ip�����]cR)�`!��G�v+J������ /@# ���@��VUU�)�ּ�#$ Q]c�f'��Mph���&��0J�Y�)�Q��d��x�B$<���E�$`Ͳ�:���W{yQ�\�a���7���4�p��,�ǜ���ZaGKh^�����Q��%�H;u*����܍�޵�jK���{�396p���#[��1;����"�L8��XU߳���L����G�)!�"M��\�U[��,#J��K���_���!H"�p��1��w��cbk��E�ZhL5� ��*;�w'��O���$5�dx�7�ʄa�&,�U�X�̱`c :T���NV{��[�9�6�H���	p� ��f嘋�m�D����t�V�uTC�� �\w�۞l~�jZ�<�1�^3���1^�"�/�S�IVĞ^����[U�0W��T���Ļ�+u�\>�����.�6	K�a�,K]����˴������PA$�.=!�)fh�-		��--��yE���6�R["9h�s�V`�����au?%�*$�I�[���(���(�mk(33������*
�~��)��o�=�܁����q��_Z= u-{2���%�wIؑ![�B��n���-��]4*��L��<;��"�*I\�g��w.S`�g����:o��ט�/q��cV����~K|o����c�	h ?A^*���-9]t��;���&��F4������`wοK��X{L�x&�@�(�+y)�xV��v㽾y0���O,U	d?Z���!������h�&���}Kd�rk��dtz[�Cn����N]����uzv�������ё�_Ow�R��:v~�@[*Q3{3AKk��؁(h&}�ArU��E���^')�T��E������4�΋q���B=g^fYɬ$	l����Fu��Bf�O(�U����d{h�DBi�2�6xhZ��1��>���ye�����[Ǭ��	ǣ���S��2�h�r%1��?���!==:�����z'Rl��MQN���ӊ&��_�6@��/�ةWͽ'���NE	�C﹦X������|�GsȪ��
d�������g=�ג��;�fߨvj��4�ZWo
�x�B~��Q<4l��9��<���cG9ֈx���0R�	�K�� }���ȧ�ץzG�"�*L�/��2H��3�`�<�R���@d�P��sO:�^�aĵӷ��j=_��Q;|<�W]�2E�EY�v�G�_{x���'���v�`퓋:(�eb3�ku�q�Ѿp�Y��J^*wT����`Mn�Πn>n�gV&T'C��ͪ�떍&ܰ֡�$��W�@	W����/�N���Ч3Ic#��������._����h�{�[$}�*�͇
�mE)������d~�S���ǮQ�\���]L�W�OZO�^3Ǽ��U���	��ߏ�$G ��i>�$�e뗟��zQ�7�Y�br+�o
q����U�D�V`p�![tvm냻Z��k�Z>�.MV��&N��Q
Df�\.@��$#�bv^F ��N�j��Ϳ,L"tb���I�7����t���Q����.�ZJ/��f^[F����NT;~�L<t��պ ��U�HcKepp,���`�������P�����0+���]�u@Z�dߍ�4�!Lۓ�a�����+8����&�5�P����$k��y����g�D��:S�:���uƳ��x%����M�� ������p޹�|w!k�r�}������!���̔�7�L��퓾'��& @��`�|��`��"V"0:��]� /��@Q�w�����^?�������R�C۽^.hg7!�#�t t�9�ޱ���20�3ϓ�{'͓�d�XhV�H`두��?p�^#�j�z0��"�5�t`��@DHWL�_��G�����l���
��Ո�b�|9��Z�\Z�[���
��5SeAy:�1L�Ew�\0��� �����"r��e�ca��w�[ O���&ĸc:K:^��f�g���B{X���]o�p��S�w��Up�ڝ��:CM�ރ�w�wu�����Ĺ���v���z��(v4<`�?�e�A�t��}~���L�,"20x���E28&(I�j�Ѓ������ب�Ā�����%��L��	{�+�qY$����������g����7��Q�O� ��Q�4�f����;�� q��|-Т�fb�=\�j��A��D�U����sz�a͜K1��"\Ҝ��O��F3��1�<��|�`������H(�x���-���{��劏fah�#f��#"nV���^iN��[��\W��,�&-�������]
�p��j��K��s���*��n%׮mKF)ܤ���.�2�(V3�lSJ�f���Nmf ��L��V>ř��B��u�E��8���j
��-#�?F�Ӗ!�՜,���dj:����I�H�wp�H��co2��*a�K�;MҲ�7na2BS4��M�X�#�aEUs�>���hMF�M�a����:[�"�Uf1_����04�o�-!_x9��e���Bn�^N�([TSs�����s�8a�	�Qt&��/D������F5��A~�E������n���t�R]��6��n��&Y��f���|ia����*?kD���q����0<?��IXǣp�(d���y�#��*��%�#���ظ���>Ʊ��t��ȭ=�1�E8~���Bm^Sw@�0�)sq�����&��[�l�''�<�?�v��A���7��t_���$kY4�	�f:<�Pq-y|�us.�/���W_7,�6��0�+�LH���������ʑ��K��x�;w�ܹ�p��,���cJv�%Na������$���1)�G��	��h�>rt-!|����s�%����F��K���ԃ[S��M`�͍��ݐ�C�p��6d��M�~6�#������(aۙ��$�Գ��N;�ZGr�f௘O�����ρ��c�Xk>aB� ]�����x~���!���J�1gM� ��R-�ě�J%��h��v��T�H]O�E}��: ��Ԅb���Q�X�^Wmٚ���3|���&+ g	`͢w1��bS��Y��n�f�XtX`5�� �<X�(S�c����wP����Xx4d=4�/8��e�]H���Է���E)̣�ݯ�(��C$�e��6t�����=���Ϡ�)q�)$�* �dA�l0���%�%�mu��I�)"H�/�T+���������f� �~e7+��o4#�덍ݩ��k�ć����/��}V2�1�R�Wci��2�U� M�
l�:0/�N@)o�m�u1fu-�*���������e-I5�����Z�-	=U���=�`��*E�\���ɱ�mKA�:����=,��.(�%�C��n_e���#i9��{!�v�
V�ϱ�C�+R����Q'vnW 8eIL�Bz�@m���]�R�10ڏ�U	6?���9'�!{�A�wm,�N�֡`�6�픃QO(���M�~/�� ��UM�'�]��a��i�
.Ü�nL&��ejM."c6@�L@0׺!i+<�<��Oa������ݘކ+s�s��G��~��<1�M�n&d��S�e�jS`�O����ȧ:��w#�VR�궳e},��2W���lD�����vEMS�Qv�,�X�~��y�"�=�:��ӟ6����.��Oh��׈��9���Gb]r�M��u�	k����X�/��P�|�"�_)я��s�f����I�M�,h]n�[�L��I�X���'}�D�����ڄ6toƓX�,c9��{\�S!�鋦�M��;ģg����f�=z�����:�m��ev�lE���Ҵ����M�%����R�W�f��)&��2�7�ͬa(Oi���M�g�p2I�CdŤ�#MF��ƧL�Y�(&Kv$`�Ļi�R����g��*�V��CR��7d}��;c
��^Pe�+f�A��We' ]\il4� ��ּ��H+Z�ޯ��a�������yK�������[���b�-Y�B�e@{2�I�	A��!ʷ�5Z�l�ն_e���i1^4�;#��~ ��A���4u��0��8��,�����h�WE7񣮶{H��C�(o�T��P�j��@��{\ɫ�.�7����ܬ�se$@	@��s�O)�ݬ7Ί+��^�va�p�%���U�<��A�^�����L����Z����A���O��)��(M�ڬ�>�	<��'����%q�g{��6pCc��0D�U"�k�]�F���H ��(|��HD�K��ǁ=ϣŹ�E�c���g�y�1|�e.�/���E��cEe�渴[*�U���RC0�;�>�B�W�9G�SO�/{�壻.x��
e<��T=l�/�cZ�J����dgB��-���`؞������v͌�p@ΰgfz3�=h<�ruk�>T����t�R�;�T@�6��4�1���O���ع���_q&�6�in�n5�4,h�5?ϭ	w�e��ǩ�:�~�3~��Z�O�2���Y�k����"m̕C�!܁n��D��o��#2i�'��]܂��� չ�)F��V�kP1[MA��%�ڕ�r"��B�䥪�ْ�U���|�0��
��,�G���2���5@����lK�@/n�L��=龎�y�z�u����x�� ���<ӧ��.��J����%�K�ޫ9H�"xWe��m�(�&H4�Wv���BBbt�,h�ډW��W
3V��p��$j&���)^~�j{��e�s���8����P�i���T�8@/;� la`�\�E�f:��N���t���D0��V)��H�4*NRʌG����Xd�R
�kB�d�f�.��%a�b�p��Ȕ@C��i�ʙ�5eK�� غ���\k�����C�1(�����g�4��������vkmz�X��Ȣ���Xk#�N��&�]�%6�Rd`�$���s>��@��
���lZ;^�I���}�*�d����	��q��ʕ32*�#4�[3����������08_i�o�!�z^J(;�tl�bY�rk���#��!��Ժ@�N����(�"��E��e�@��)��;6q���U�g|Gһ:�4���^[�'��0��	<M���ڙ�	��n�
B�Nͷк����ɲ�jU0�%����,�W��+)����dE��?�� {��Eެ��5g�2~~�zV�K�=�tMѓr��T�­Y��� +������ʚ����
^�k���,k�e�V����޸o�w�a)�53b�3v�����.3���N��G~��|��'�����,����5�~��Z
ޏ�\�!�H�,I����s�]kE(�A��lYë����H�8�+6ї�Y�'Vj�@p�����}7�%�![��x�/p4��F&���w/m�p/�,��R��3P7s�n�̡�kx��Sw keP).�.�X�G8���=L_Y�d��*�%�E?H���#�7`��AI�g@y���R���1ʋ��Gc�j�~���Eg��8O����o�7�P�*����!1�H$Bք�a?��.r�.״m{⟷[���� �KYYR/��Xk��t Bk<1(�Kќ'�zo���!�]�7�.(6 -��W��ۗJ��h[�@��ǎ`���:H��C�[���lS]M��j|�\�ȅΗJڟZ酃a }�4Rh�Gzk-��\;`.����g��.���2�_��S�Mva
��h�L0��D�_��V� �W�m��8�⹏�۴&���k��Q�ü7��}#�di��c>�0�gD*\6�lw ����H!o�.�ȍ_�"��tyN.�Z��IY��,)�$TӬk�Lr���(�I �܆��s]�F4޹[��$�V$d�
�8~�r�S˪b� '�`���)�x��f,�R�v��H\E�'h�G/+��#�V�y:հ6�T��Os�s-+:��������jy��!�ք�'����a����RnG"�/�����IFg�5q2��NS�n�͌���K!�)��y]{��
��}k'�h��)LD�=��k�nC]��&r� �U��7"���R�ĜZ�w���jVɕ�V<\�A$}/����IE��̻� .̝�j���b�M�ꑫ���@9w& ��Q�к����v$�7�D�_t����du��ޔ��{Db<���]�x����ߓ����K��##l٨��OU����$��߯w��K��5����%J�J�L�Wi%q�r�}5��ߚ+��A���t4G,MwZ����Yq3O��,�bS�����K)��z�п~Rx����b�
b����.lƿ2��0�1V2-d��D�/����ѹ�qk�jDo�������N�r���Ply��ր���Q�&�v��g��Σ�=j`
x�$��E�"I��;�q'���%�lQ	kȖ��1����9iE���LJp���(�-���D16��S@�{KO�f��P�#�t[!�iQ�OK%iﴤV�_��q?܂���nF;�Y�����V$#� Ȍ/F΋�
YW4]�תa_��қ�����ߩZ��JB�a�� �⊾�����)��V�"�
��yY�|�Z��$� �x���c����柠{XP	@W~ܰ�1��$Yl���x*��~c�oޜ&���Nr��p��f�37��
I𤄼���.���������x;)8<moT�3�w-)��㿨�����9͖iSy�w���xvBͲI�J��^���x�#���	�N~˧n�
R=)4�v�S�343�ٔ?11ܛ3ݍL���W�k��M�x �-��4��H2�6�++�}�uyl�� ����[�����e�A�Pn?D_��~��,
t"hG�ʢ/��-�r\Y{,���U|NP�V���uP6��"���M�1�y�W8j�9I%iP�0�;�J�Yh��f��R���j��K�4�G c�
�k�m�('�n"����~?	�����q�ɫJ�deC��{���6�'�F��&��k�C�\�<�̟�:?<8��(C�p������2kL�j%�	Ni\><d����{1ɋ}����k�ThN��wrv寗�+-�q�@��&�����<�q+��߯,��ld� �7 f�k�hʼ�;���Ԛo��u��-?D�q���I�*⇷$}��T4\$A�z�,'4�*in�O2�M��7�B��>Iˢ��s���-D,F�	�}�h�\�˗4Fm�@�M����~�s��m<ayM�rA)DX���'|�=��E=ԟ������=� /��2���S9(���G�R93G�C���|?�������0MΌ�5țC@ �` �01�Xu���K;�� �"`&�[ݼs�ZJ.Uz�����p����8iOI�O	ldh��{ ��>I[-V�u��{9$��-4�[����β��j5A�b�j؂���� C!�4���gS)�� d�J_�y1(Ȩh�Q�[ʦ�T�� ��P�i/{�N4��H��	�;^�{oH�
�#��L�|�q�]@�a2y~�+ߟ�9�h:���oCp�m����v��o��� �����Z=Ke���ʙ)S�ѝ����~�������G<�%VSЂ�a<*j��^��U�yU�p|�j:�O0
1{N	AL����0}H�Ir��1'l7<��oH!p�¬$�z�7�?q�@�K���,���!%��]�Vѣ�1 ��=�DǾ�a6�I�v�
o~|4##z�!��
��|�:`�Z���M&-��4��?��Ê֗Y#��싆�)Ď����/�eJ!��TƟ�������c�u������7o�~� �M��L2���n��@�⥼��-*݃x��*�"K��&A�:�@� �q��5#�8��D��h���n��ޗi瓰�*=�,��"���+����N;1u��<��^ɛ���a텭	���������ѳ���
�D%B�2
5��O��oj���~ W����<S|)�6�7	�<x ���{�ٽ�~��s��v�{�E�8��<uy�E��鎨8B'�V��o�d�Q�y���B��_�W7oT��ݹc��^3o8{� �^�P�vy��$|�=b��i3v��ǧ�wcg%0n%^��yj�_����[F��ZG%� M��v5�&�X	�����Z*I�0�
���JFC;K���F�Q�`�U�A|�D�Ͽf̬�Ya[D��悫R���[`�Ռ�_�����o�;nw���]g�Q���\.�u)��a(*��ߓ�Ʉ�7f�ƅ��M,�z-�a����e.�:��n�Hx���M]e6h[��ϣ��=��(���Dv8���%�Z�6��\ñ�̖�$*�>�#o;�`����j��%�a���j����;/M�i����&� `���ݢj~�O�R�(����F� {_��� �8�︌������T�M@�{�{;h8'�QZ�4�����d0)4���_�hB��Z��w��fՉ�Ǒ���C1Π���՞@���Jy�~��'Ը�:c5�=��ʥL���b�F�AD��m.�T�K ��k��!�Ȁ#��ϹI�����J�;�e����������'/� �
ɪ��j/��kA�0"�
Z+�g��IR��Sp���o� ���|m:�*��ݐ�O���S��ߥ)���D�YX���Nn�+�[���3��'#�Ut�!X�v� ř�s�W �u�2	�,��a?���zᢾ��4���
�Q�}���
�����bRV��FO��u8��)��c��	�H7�=�#����i�e�.i>�I��$ ����?��Lw��y6�@88��׻T�XI�Lдˊ�)c�Ш�^	���OLdH\LF�hA�0��Q��n&pkA��a|�6R�d���ho�L��-*�IS�����R�X!POz��-Sp��gX�z ��RT�k��m��d�2��Hp��E�#��%��6�~<u�'�ElVڰ*~m@���$�M*��˵��|���'�iXV�� ��|�"|���*[�4V���|��/����|��r�,$���BB�EFw���}�Q�lf�:�l���5��K3�^���Tp46��<ֺ����7�|m?yipxI�}��������%��y�J.�'_kC�1�����7C������4F��i��(Pz �0�HM@QP�����.$?	�B.��}Sn�o�@��}�G5��z|�3�MU�6�a�M�,I����~���6�{�@*���%<IUr�	�����XI���K}nvF�~g�IV\HhB���f�[-�-�������4O�����\�k���|�����B�HWG��հUN ��~w��9��6��+1	� ~jD�zƋ�j��Mv���'}� �f��,}Q,%�!�䖉�	Y�,��wq�S�#��H�h���� 3&�����o�����2�����)���:j��Pp�K��c����I�_9�&_Ed^�G�8�F��s��q W�*U+�'��r>�ʰ��$C���:�wP�Nq;�ϙ�w�K���[S29&������瞬$'6�Է�(PBx��X���/��*n��ucN.��V�CF2�7[�`�m0�E�8h�]��N��	O���c�d����k�&�܊|�W2���O��s0ώ�k&��v'���y���į���Y���s1�\�E��4c������XS�ub�Q�+o�����zmM=�e��d�eU��c+�t�ݵ�x���ENSe){9K� ���̜��dEGe��a_�(��7��'I�`��A�m�N"�6��%ۙ�r4�M]��ܷZо �Y�_�<���oO��El��&�6�&��y�B�T��.zvc�PQLy�0�ޯ
��� �$������;�P��N��\��@����5,eq�0X���$��o�^ܫ����/7d�j��*3sK8�a��$�W׉Pݒ6�2e"��o�	C�qo�ǜ�O%�Zj/��/'^j���J��b^N����Tk�p)$�@�9��x�	.Q�n��k
K)�euJ���}��]��aS�_�S��c�o֝bӲ���c����7�P/��65ȁù?���'���S�K=#n��%��H�>��-#�y�:Ma���I���,0� z��6F.O`�Yq�[�X�~؃���Yq����P��P�XZ��D �>OG�P������L��#��!d���N�s8fB��vq�VAԁ�W?�C��}����B��R��X��Ȭ1<��
n��G^���K�s��>�J���It�W���K8x�5�cĨ�5����|p�uJ�-Ǉ�����AB���Iڒ^����fn�(RR���;@�	�Ǣ�bl	�� ������*��]ԟ�H�ش���Yc����)�',���C'��[�\o�!o6*��?4izh$*��=�����u��� ,wF�,�X�v���xG+}%��8�t2� ��M��퓫�/p����Z���u��}M���� ����$�#@��g��� �����)(�`��[}�Ńo�c��@�[N;�d��իGK߁���6�������y���-ĳ�r��.կ�.�O�9��"�ˠGN^�!��~��X� ����I{L�&����S^G��4�З�-���
2�'2x�w[��
j�]~ϋ	�_Xi���١��ov��;�{Ír��,ۡ����Td=��+��ӛl-8�c8�[!���4O��}�[�m��LgS��^M����o�����6K�}�k�8��5�Eu��) �yn�!���dR�"�A�<��kpJ,K2� m��#���{ >�:H��~ ���Ɩ�\ dʒ��⬫��P����J�&0-�ɡ䡽n�����ꋔ��@��  Nd �D�1L�ApV'��y��L	z6��?��}9�?��
�T-�K�I�@����g�	��[�Kb������L��eݜHx�iԨ�ܽ��w�BG��9�l"W�"�Z����Uk�FX�O�f }�x�E<�f��^{Z������<#�]쳹������x��'Y�ȅw	o�$�;�:�"��"�#Ҳ�=9��|:���<�
L7dp�3�C��F�ޑ��a����@�6e%�E���t�E�#�HsE��7)'�Gͅ���b��%�oC���"U�iB���t�#o�GC����@a����6K@���#&�,�uҿ�"~�x$.{� m%��G����?��~,�Lϭ�:��aؖ��\qo�+�)�w�҈v�iA̼JK6���f�5�*�H�f|�G���8SEyq�;��g������"����כe5[��΢��R
;%��C��* o��<�Ɯa3��<Z|Ʉ�g��V�%�c"k1�6�U�u_�����^+��WPa�l��o��n�;�D({��'������]�y��n)��0�ȩe���� �ܻ��:��*}o�0��1�lG�����)�)b2ǩ�K��*�i�DYj�Xm\Q(gm��4��`^Ժ6���Us����i��֪�n-���\�0�]cV2�7�u�&H����޲2�r�\�c'z���ɋƛ�P�;;=���* �A|��[c�i_;��zH�h7���Yn�@C�����R��Ėd�ab�!".TQ��e�؛|@����T��p�ݍT�s ��#��#�iXz\u��@O��Wd�+��Յ
{~��R��f~����M�|
�,��kk���1$q��ӌ3�*�b��C�!1G51���J��p猦թ/%���=\h*���7�=\v�(��o�'���TD�0����ϔ�� ��L�X��\6
8�U�O��s>=27Vّ'�Xk�?]�Q�*2�N�]p�^�L2S�������yA#,0p߷F�*)�O���Ź{&�7��y6��quJ�"U�z2S���W�Q�!q��v�.��tkb�A�l�ؠVn-�8kej(���Yx��R�9c�7X��X6`��6z���N�L3��_��%R$[mi��Ck^)��{��j�|���8L �^�K�\SQ�؃z�B�d4=X�7�g�p������;G����Qwl̋�$�ȡm�J/��F��yX5��\�����;Y�K�sY�Ye	H�0��H��<��X"���a4����<�[9D{����ll��D�rނ��/���k"2����* ��X�<�?G`����� ��B���K�ԗj,+͘����}�IK�cko\~L����3���6}s���Ĺz�M�t��via�������a������U�����p!�=�T��%����o&�d�V ��@����"vuf�x=w>2�X�2�0�-�~� N���i%���f��0mȽY�А��%�+D� ]Vor#���(4%����^�cnG>��&�HhK{o}��T�u$����4�e��$nd����;�p�A��|.�X�d�J}�p��*>\�9ܥ�R 8љ�S7�[B�-�e�;��]��0ɔz����T1)�'2g��]ME}o�1���L�����S_/;;��u�T���1Wm�n83Ӧ~���-�%N����!Hk7r��,.T/ߡ��\7d�ܢ���pC�C�©t|�;8�#�;T�t�������}�bŁlˢL���~rn��$0��&��B4�����ځ�G��������x�IL��BF�nq����j���Z�q���Z�Q�dźj��~�_;���(���F��7Aͫ>���g^0��?���N��rsui��up�zi�@�Ձ!�,Δ1�w
��ut�=p�x��_��hw��9Kl����7!��9��5*4�y>�&��'}s��T�KkJ�J<5�	Ըl�9�~N�q��bW�\�
�T�u]D�2%�wE�N���wk]\]t�D�'h?�;��*`U����I�A&�6d��~[7��o��RQ��C�M�o	���v�I�qx��>V���$rȒ`0�ʅc}����<�a�n���u;�a�B$.���D%��!�6*��2|���|e�z���Xڰ����(��sw3�Ȁ�-���E�_����>�����A��(��n�SK,��Ҝ����s�[��P1�[��q����F`T$���@YВ�>�$eu�B��|9Y��{�w��4 z
���Y����uɦ|�V|"L�,C	��J����R�~��,z���B�Z�c_"3�:�]�>��_���!�m� x�@1$�X�0���eg�YJ�������^�0��[B�Z1/g���O/R!^n����A(�n����O�?���������h���4?�����pe�=�6u��݆�T��UǏwk	Mʍi�e�V����8�ü�v�Kԧh��giI��]f��2�� �?�-<���������{}쾡�֨b�sث>��՟:Ke�h�H����&\g����Գ��`���BW��U��g/��*�۩�H�F��~���q���ef�o�2sR�@��d�rK)����upt6� +������Cj����R�M�|����_�5�`�m�z�� m�����"+i�`�]���ǫ�����	�D��G�3��U`h���r�1 ��>�	Y󋡞[���Ni�J;@Z��3u��.�r&�O��IK��I�E�fS��|��p�`�Q�j<�)��$k�~t�e��[�T�c�^����M�Z�n���F��FP��9�O����T��Aʗ(��r��3���F>�nz��U�.�����}�[��
r� ����P=�܏oP�#*p��h%E\�i�7!j��nfmq,}�4
͕V̂���rC(/A0gm�Bup� �q��r�x�����5vw'�J2���ޱ���.�J�:�'��_�s����OG�pi��ӧ�8uz7+ۯYS��l^�C"��2����p'�y;v�VDت��yƲ�M�[�P�w�/�ׇ�T�y9hq���#��āfG�4���}�n�Y�˳�3����6��0�D`[$h���A9�ߞ%Zd�!OC�#���3T�a� ]�H��fG���ku͇�NlP��L0� �?;�*���>�.U={>˂7@\�v���n�H=��D����*�:��
��3��\���A��O�!�밻��B��-b	#����uѸr�,� �|!*�Vq��ӑ�ͷ�7��?�$�R���w��&��3���-�P����B8d�h��&�+l�Y��0t��`��Y�A��o �7��^��F�A�b�,@���8P�;��ܽR[����kD�Z�H�� n;��(�$+��ܸ���3$=�k~#��/$=���AȐi�
5Bk��6��<i�k��Ʊo�4��5פ~>ı=+���9���x<SiZ��Ri0��yM=1&B�C��a��Z������w�$�ƚ�I��X[����_GE�ԏ-�{�Z�RY�Pȋ��!�q�Ic��P�]��ҥ7i���U˷��j��$iN���ͭJfn�d���w-�m��
:�/��V$�>WB�{nz��X�۹ȳ�D0������\ǟh�r6!���L$� �l�CoQ��?q|��>^-��A�i6��ǂ����b.�~���t��� ��AD���s���P�M�9�<�%_��ҩW�F%���B��׫#RN��1n������H���|��h�z�H�<&�#MӐ��tx�>�m��ٌT�wRr��r�S���zqz�`���9Nm�(G&�n]�;���\�fa�<�4����zi��9و�Y.(�&�G���,��M�gE�Y�*��E~(�ꪁ���z��a#Vؚ�Ub�=�L[�Mw	4A�C�YE�#̈��A�>w$����6Lg�����ft/)�F~���o$m�
3��#l6��6�ȉ��ϥ�Y� hd�,����f��_mg���G;���x0|�xNOY׀3��T�8�ω���OP�"h�m��r��2���[�o΍�$�!U�䬓��?}��}�݂��;���wҀM�LP����@iV�i��Z�)�F�����_sF4�g���D7��3y�͹���,ki����(�ƛ�b��T9Q�	 Y�=���ysN��K�CzR�f��t~*q�I���1ɓ�󸓣[�9���1yXe쎆��q:[�^�,�~,�.0b��Z&�m�1QlG�K��@v���̊�F�
���o����F�_F� p��据�]�[[��8+���]�x�ً�[a;h�����v���T4��Q"F5��>�'�#S���,%�PŃ"���f����&yR�;�W̀�lL� rϽ�����R�7���{>�Vǟ�\��[��?�D`�Ԗ�d>͌�|{&��R�w�VX��,6�IUl̇�/�,:��I&�ێcD�� �iH�׍U\�F&O�����P���.��*��ƙ��Z���hw�4�M�5��O�1��9�Ij�I`����k����%˲h�_��_B�A�� �u���-�B2]�P��,���$�ϳ����]�,��B��
H/9/=��T�9���i�oP�\�8�}P����ds�+b�R�	�m��]�T�#�SA~D�̗�����-:�Š�=�8��J��~Zd���TU����e��D����B�51�#�8ix�T�a�D�m�z>VJ�D4��Ts7�U��ʲ������}C~�����RX�8�P��E�R����x����P�ky��sU���(Z��f�g��\��?4���k?���gV_���k���rqa�����=2ԏF>]��]�d���s�9��ǎ|-h����鈫�A�׆9	{�R�,Z�"����5����H���.�k�O%(�6q�މ���=����KE2�؜�²̦�i��2D3�D6��O��W;�߄^-�ԇb�ٓwZ7	Rʦ�8!��	�$H�,�� N#[�����P�gϴj���2 -�.� �#
{n�ߚ�i��Mk��}�`�<d��U�IM�=���L��<ZNB�)��ވ����Y?I��D^T���fyZ�<΢�w��@'���z�7]��+�Q� U������rƅ�BZ麾���A!��pe1n�ƃ�d��j��/o��o�~+b;��c����v^�]� ��۰2Z��#�s��$�45�p��^JM+���0�9�B6+��������N��� -)ޥ)y �ڞ�B�˺�:�9��dl�;}���2x���c��g#��?��N��.h��*�:�P4�N'k��ѡ�=,}}��#��*[�X��b/�h��h�M����h}Ƶ��6}ժ�[��Ey0W ���Nޚ��RNw��C�͟c,FYP^�i�6<�R$��!5&#m���+���5���xs�<6�m�s��m��4e�M�)�e��dɘ�{dz2I)\⒲���n�R<����/%SnK!�ja��*�l�B���U�jk��g6�`eUN<~;e�=�f˂�9^p���Jh��S�P��!�9
Շ$y&��6nLBb�wN�(�㹞�w1�EW������F���wn�G�g�o�DfڀR�����s�_қ��72�>e֎bfS��JF��{�����j�&��@M!ԇN�2��r^��(��ݴ.��}�syp��0�V\R���]�y�"����*�aؼ�<f�:�����F��|�xU%��i��J�
�[�'0,�Aǌ��p5S����	E���	�@�I�����>W*�t�����+e` ����q�nEin�B3���q�}��v��}��zP[u�h
 ���6:V���)EJ9&���~��*C.GQX��'�9	i�έ��'�ޑ��iO��zP��Y����&���{�Z���/2�Γ.���s��5#���8�Ԓ�.�:g>.��
�p�N"�y�75b|oh�#��DxBX@��?ZiFT���n��+��Ҭ*s���E�$` sB�U�)?���Z��"�
�!$%�4<�<�I�O�Y�r��̣)NT�>��mB�1�B�EQA�ﶝY���^��7*A�C��Į��%�P��s^��ݛ��t��:+�~씄��8�j�d���w~w��A巿����4s��f'�g��c�;��Uj������)"�;l�<\�j��n�d�<������Ǖ*'z!DБ�����U�D{�Qh�^���ĭ$��b�L��Of �f�/�$�Ґ�+�`F��
uR6�C��8v�6��5���`%�K�{=u�DK~�䦁��R�.%4(������2<V͉�8��M�VQr�2z��V�Ծ_�E�.c��F��d �|an_�Q�}� �J����Vt )�1��.2�Î��Ƈ�c�os���rkH#�Z��"q�V�=5|,��_�����a�PBn��I��o5�ݏg2�ڑH�4�����ú��}ҝ������	+��Ɗ�K/��(\3n�.�Ɖ��1J���b3�E<OkJ���ȷ�)��DK��<�͓);�m�3@�j�xw*�`?~t�uf�S�Xp2q硄�%�u���c~ܶ�okr���W�i9Z`wW(���X�Ҽwkv7��Msp,o�F�8�-,����⊄�����k���u�xH�i�9���H*^P���$m/�����S�Fhγ�9�� @?����]��7�*�;��&<��$�� ���W`�*�u�G���q�/�D��\�M���`1DfO{�]�T9]c�n��p�0���_n�9>j�v�?#Y}�o`��*��an�O.�&�F�����^JO���%�UHLW��/Ut��Fu�#�:��D;�~�f�5=��R�S��ǎx�H0��ʘ�<�Čn%l`c��詋p\\�M������E�.��,��)�O�$lܦ3Bu_;}�s`���_��<�\��]�>,��d� 9X����t�]O�'Z8���i�1ֶ)^�,�Al�r��sW��t�����gX��/�c�YsA���# ���Ԍ/���U�Y�R ܠ�ɬˎ� ��S�@oF=]�P�¥�����W�&��/���|�7"�@�"��0i��.F�R�8�0�W��_�)];]��Q����c&�4���	�<�w�$����ʛ��˸-W��['@eRJ8�k�C��fk�>&���6�8�;�=M%{3�0N��3b�����:�_���wpD6��-Y��"����>Y~x��y(�~i.�U�(8�����X�{�,A ��K*�/�h\s05��|��8?X�����[$�R��ͮ�z4fnp/?4���5-�LQ���Y���e�LV3�I<��'����U��;b�zR�aϾ`�FI[J��"��f�FM����\4��8��cU����&��u�[���>�v���78�/Ư����z�ݳ9mh4��ͳZ~��ݟѺ��`����V��K5X�J�Ņ�^�i'3&Vg�_K�*	(2�^SJ���2��H�H#�c����� �'��e\.�B-�����?���c��6���� �Z3����d8�p�����������Y���I�]W��{�!�_��ѥ2�njMq�bRٝ�Qr;`RG8e����(�1�ֶ4{1�����д���İ_��OE��vu1s>�h#�o�0����fU�\s� r��S�;,�ۖn?>�K�����S�@Y}�"�S6'����>�#-���D����E�%gz�ϵ{�_�`�.���c��_-���sg,f�r�9EuZ���{��uw$�������^w�W0E� ]\p�Y�݀�;���t70t�;�'vBge�尓y{ڠF8�s�O���K��%�PE\��\�;��+<c�]S��+��b���`,�}��K������ҹ��bӱ�ZK���hk�aX!
?V6ɝ�gs�!X�(%!_ｻ�Rq�ހ���w��k5�w�x��ov2%���[���!�
�6`ˤ�����(�s0&��{o�7�zc��>mu���O�)�HeU"�-p�>�Ǩ��a=	�KTU���E�v��9]�4G��*#%>���~6I^�*;K@sE�5F�ϣ��)i�0�y�%�^�(���33���XZ1ݖ P�^��t '���~��ha����>>�M���ȅ���j�׼Eg ��
��J�P��:HI�LC���m�Pذ��vv��1T̵k�M]W͐|j'Y��B��?@�;"����0��u�BI��x��a���N~j�vev$�a��p�$�)D��}Dd��a򁳁b]ѹ[�v��P�	����I���g@E>p��{W��u��?�X���%5e���ITU~��ܶ�%���Ea����T��V�I<�2����fFln�8%�gwıS�w��\��=�6&^�3-�jpm����3m�(k�O�F��<�Z���<�������(@�d\U-a�wI���Pqn}��̫���8���^�D5�V�Wg"/JU� ���S@$�K��^�%��y��W1�"�R3��	�!&���JJ�4С�AS������a��% �-������
����ȸezc��_4$�VbHFo����h��ژ� �|GA@+C��S�&{R2�Uӕ�0��ؗ��ym>������V^H*�����%�,� �n�-��l�y��-�3�G�wڂ�j�P�X�j�9jM(������q��,�Ɗcz�]�a�������`U��X����������%ް`��E���Q�Z����f\�@��^@˷U�H��}�	:� s��G��R�|��uZ{�`d|8�ı�@�w��戅�7�O�#G�X�ŬĠfp�8s�K� �υ�߅�iεT�G�5�����kd�sz۟��B\z��;D�8+����J
�;����V>gP�!��t�Z�AT���J>��e��W�U�E?�L��K�Sᅠ���d�C2&���y��<|�D[|��Rz\��hΖ��bm�.���P�b��+�qz�π�t�4F4#�Q��q>���Yu�	v�W�ǅ��[�YB9g����2��D��$=�ךt�nٴA����� h����\RhXN'.Z��@sQx*pLg �16�*K�L'#�����rh�Q�2�SW� w���F��Mc9���Og�|Q���Ֆ�y��G�V�b�No��o�ҧo�@�nCc~&��?�"s�9�Q�k`n�b���H�2uJ��k�ߓ��������:������r�5L
l���,��ڳ��"�<P�ݛ���Ɲ[>\�+�Z�5��Kq�('j���cA&��j4u ����e�m���F��e��W����V����n?'�ɔ\`�Z��J?R[F̧��Q�"6�CEq��㫒����V]Q������YDJ��+�d� ��D�B�ٕ1�j�N�f㪶=ɟN��X��#-95�Pw��`r�<U.���zJ!snT�y���Bg�i����'a���V%mq�����l{\T�i�?�$C�Y{㇕$l��I�y�I�Uxk����;G�u�6Tk��r��_�h�F&�C:�5_���a�)Ͷ�O�LS�YPK	�5�4�ʇz�R�׭���X��
V��F�t'���{�a�J�Kn띑��Yݞ���e����(ȧ�dk.d_CcJ�~��7Q���hw�n��Vb����L�v� 5{��Y�8Ź�������~�YCq)+�Y����>�o�@8c�T5z�ɛ�j�I�Y.& P�$���y�hZG�?Ȍ�� ayn7m'��%�f������}5���3�%���6���cq,��Ɓb�'����$[C��`7}LI{ȋ�����d�L��	�1.E���$�k��Mܽ蕖N������˘�����W�Z�F�� %�6����so[��c~qSpt��?��؉������?������@��i�>4�����(j�|����4s�&�.?1y�ǰ�$qi�!H7?��U�&ns��H�)�3/��J_W��"?�W&�/d{��=�ݪ�����k�y�-Xt��7���ԣų	�/�]���!ۧ,��t�(^i�M��U� ��^(�	A}����!D8K�'���MW����ӷK��)έB�Z��%�T��"�)�'��2?�1��dO�r�Z��Z�u��k"Iʡ����5�{���Ô1� G��b7�o�;�D�f���Q���I���v2��j>�]Iv��LK\�d�jE:5	�|�ҽ�/:)�]�+5#q������+)\e/��V4��lI�����>�qdb��V�"8�����L��캀0���FRO"�v� R�r8�2�P�heE��X�Z6';� Ǚ�����8���:m������k�ڡ!6g{�0J������D��:��7l){�VW'�*0��x���9�F��r �q�k*i���fbH�d�Od���u��\[�6�,�e�\�X��f�y��+z�Wa��;j�k�8�B���!���:���"Y�УKK!�n*�%ۉ�<-39M�3�n�1eݚ��^]Z�
��,��l�S�:���n��{�pei3i�{���BmLz�A�\.Q���ET��_Ғ���AO2�&V'ي�]Q�������<� �C"y�y��Ew�՚�����j�����^W�z��}��<k�[��=�r�WR�MSަ�l�	M����G�>�Ւ�}_K��qE��4�ӑ��N3��w4r~r��o�Q�D�	U�Č������Ԫ>#ˁ@�w��i]M-��<i�f�R�	�;y���5yO	�����!���ȲE�"+����\ҡ�Դ�n�~�S�J��E�1e-��ݾ&�����箊ۘ@B9B;��\a�:�s?{�I�&�(oo7.�uȔ�\<���Ԍ��������/e"t�8�R�L���=]��@~��P(�N���󘪦Zw䟳tx�s�I�V�w�h��B$\t�.X]s�3L�YN@�^���}u�M�i��" LM��b>4��P:���"�'m\����9>�b���G��*�M��܌!770%qíh���whtB��fXQ����X��/�����Ѩ��",~
r\�?鴯�ߐF������k��ߣ�=����&,y�BN���B޶����=v�<��1��m�Pc#h,��b�N�����:�qقw�����)�4�y��7���f�X./'	����*��8��&S/|�M����f࠴������GUJ㓙�x�(sQzk����}���W�fuv
`tU�/l�(P�Z�ս�)N5���d|�$O�#7*�'�?���W�A�:�V�,�$(ȟ7�4/#�����͞0��c�F|$߷˔2R  l�D�Q����{¬��3kP�#>�bx��@ƚ��5� ��R-���(6���˪�ƾ��"`��A�2����]�縂x	�f�G�_��S6�l(*��8�h�����.��@�8�����(�-�+mL}
LN���t|�Ȇ��y�}�+������_(�>��RHT�������/{t]K�5��zM ��=?����Y��k�v�az2^:��
��*?;�v��ÚN����n�o�����X��38m��V��v�ڱ	��+'��~5�`7�a��X#�n�x�:�wެ��!8 Ӗ�^�"�'3��[�C9�|����c��t�X��CǻO��1V���nsF�C.Q��Ɇ���T&^�S�<�n�4k��?�γ$y�z;��y^�_p�՗��#�p!A1�'w Ǐ�_���a�l��?�k���>�w�*�h�o7�0��W�xR�l����aiw�^��XP�P�ɲ���������ص�K�ƞH�]��܃?��x����͏nT냷F#a����s䱽� X��>%��V�Z�����4��"7�q1ո��ɂ�(��c	Ȥr�0>��`�X2�u�\�n�`Ía��S]z�D�7�-����[D�C��@�M������=:M�����[U��m^��-�5�.���(0��#���ׇѭ|hlt\����^ ���}۬���!>8[s����w�}�e�w"�cɱ-S��Ke� �#a��`r&2��pB���-���Y��.�RE3uk�|���L��r�Y�>Gd9��D=�ݍ2�Ä�{j)׍��e)�G�h�T����̰�~��S
~D����	��Epø�S�u
��r3����Nc1�&xU���^��!�!���m��!�V21���q�"��v��|.tj[V5�Nj��U�P�_�r^P@�+�V=���:43�߰�TX�e��Z[4�R�I(tfy�q�͉Y��_6��5z��qۃ����<��<'����[���V ĩ��z�e�O�+f�0r2I���ExbT�~�7(�w�Y�&����<��n���f;[n!M�ߪm�1l�}EَOa��@�j�C��i���~ET���~��a.�KaJI�+������~�|�:[��v��:���a�V��:��*�� z��:����m��ڥ{�FSRDc煉�l�� zl׈���oe#���_p1���L��Mi����?&4��hI�/�$->�t�g6�4C?#. TR���-�68J�������W�P���K�g�dJ-�ZiHr��muXXV�
�6�)=��D,�����*���'����R��
hk,�p�����e������- xzP���hŭ<(ԍXʹ쀶Q���m�ֹ��|��i��N#g�Ni,y�>*� ���}"������y!jG��ݯ%:,��kMe�J�d�Z�7%e̞��"�P�G�8n���.��T^��r��`��^��i���b�{�ʰ*8V�(� 9�m��Rá�<\I����7YRd�@u�����"�Q�͞/��3��=-����)4��HD����/����j<��n�j5:=
q���ҌY�ŝ"($��Ff �+�s�.?�}u�;�l( ��⮮�Ӱ���5��n�� ����F��H͛ED��Q�B����N�\��.�d0�X��c�������a��!�
�a�HW�3P8*��3�*O%�Y���(i������	��eH�"p��|�h#�,$N��nn�����
H���N�6.��ƒpn9*	�z��*�q*�`�y�ɣ�y�ӻ���rX�1r�Q��h��B����j��[������+����S)�n�r���SCc+�\�	$�mP̾A���i?�/<�#�L���H�h	���4xaNA�c�P�DB�q=E�,N��b�ުz� �]W��O�e^݃/&p"}zH��Y�(КJ�V>��hV�	� B���V K��#{���m?�G��C���_�=~�R�(>l~���'�gT�b����]���>�%Z��Y�����yL`�8s�~OJ�27���b�{#]���kIY��.	۞�8�*F�#�(Z՞F'�
�-����y �2��֜,7����$$҄�M����
؟=$����x�*:Pg�����t�����]:Sᝒ-�"9'�V��|u\C�힌�#?Ӷ�ŭ�������E�@�Z�B�P����3pK o�2�te-��y�1m�%$�V|�o������E��ϻ��8�͚��A�ї%�B��]/������z��O����

Ucؠ�`|"E��A��Jv���Я���#�a\�"�T>LCp�ɛ�.O0<����2�S�W{��(�3����h�i���l0�fxoC��h�!m�j��h�q���ʃ�AFaх���kP}7�Qx��`��ժw=�="
���&�z��ڞ�n�V�a�l�j���6�g1F~�U����A�iťp�DԂ;�9~6�47
>�&i��5���)G [MwhN l�x��{U��k�����'ؐ�W�K�o8���\�%w�c~ӟ��@�b���濫���i�`�̢%�p�:�����"a��1��V-�������-O�9{�f��g"��%,�F�d{�O;���B�>���@���yVA�d;r�����9ɨ�k���D��\ԕ>p��H!�i�>�f�3�솖���Y1���8j��|F�d�:ob1hp^�O��t&�*g��y�]G-ir"�U���Bl��`�s��gA�� J�s]Zk����^0gi=i��Y�q��̡Y�vw��l��(�>�9�]7f;�ν�[.-�F�/b�'��;Ks�I�c\��L���g�e���;��iԧ��ޒ�܎Q�l qHH@{H���/�z~c\4��ǅn]-W瀔ژ%�!�H����D�� �Z/|b�����&�js��r��?i��)�D�o�¹ڗ�ӧ��#�O� ׳@4r#4+7��f°I�P���rS�`� ��q j����R������vș�s�g��<d�遦�Q[�(І�艞������d�FO3@w�������2q��q�\��RD���n��O���m�3B"�u6p{����}L�{yqQ#~�`�l-�#G� t����JUR�]!�X9Z͇^��?\lx
cn�Z�ϖ�V&� �u)P�hY#��.�����O���@�e��r:��+߬����̎�D��z��Vnu��t�/�����$�R^�������7d��_�����ݗ!�F,��_EmP�l���4Q�X���Q�4;Y���*���n�Klv�`���Z�i��$'��3���$��4x'��L�󲛘
VX�:]����V��̣m�jH� ��S	�D�r��rc�L�-�G\��XwZ�4�.;-�\j{]q����֡a%tE�M�oS�|��\B]�c�Y��2��k��v�R H�������o=8�/��J�N�Jf�Z��)0��E��X��4aU�z'���GC�{��#���5�T��L���#|0�#pQ�<]����v7
@�<����\D�n��G<�ո���p�^<���tB���kh�������d��9c�`�o�m"���v�)\+��?hq�KBآ~m��n�a�vwz��j
�Y���R$�g��,����2��]�_�>I�H9|��	pGSD���VR�qkь�Ycn���R4�!�fg����S��btq!"�A�o<���O���^:����Tpd�����(�����:�L��ݖ7Ml)������QC�-}��,��#P�.kj�Lެ�+^��f�ȟ5+�J�C� ��ͳ=E�몹����N=�m����+5a�_\���?���.E �8�h1�G��jN�w��NX�w���Z:�M�Z��	��F3�嚟f�=�T��ت�)���PDH�(�`�I��H���c�bm����+�s���F ,������ڋ�0B�.'���4�"2q�r!��P*i��lY���
�	���&��2�lr�%�|X�
@d��Wa˕l�Y�(�΅�Zq�+h�iQ��+5>�z�
��\t`G���sh�Y'�|�*/��1]��v�H�M[C�T"-��}.jI(Tv"� n�C'~�Z�ț�_ݟM��AN��T����c�9��T(Y�:q�[B���Ŵ;�I�m�����`,W���Tr��-���$[(˩ߪn*�ٮ����q?5����R������Dh���+��;�\��3*օ�� D7e`r�e��ۧ��1�}�͒�{IG�������/�y�έu�Q��~W�V�!���u�}�
B��)�|��	US9$��N�9+/�%��"k��?��̸TE�|�U%ZS\��,�Sf�(����NMq��$�uQ�^h@�SQ+j�U*��A3r^����&ý��냉��������Yf-7�[���]~�OK�p��F�}}�}�F�;�io
Bw��x�eϓ&��q+s�j��y�� �q��a�����Q]J�9上����>�9�N�[t�桻�/�.���!a����F�F��_�2q�^6�ڨ�gA�1�8+���yD�uac��|�#��Xv���c�G	P��X�A�����On�_�~���}�;`��8{a��-X�B،˒\�G�,�jx�h�N�O�рu���OL��G�u�L�z�y|l�%�dG���L*�8:�(�����${�b�%�����O'�Q�Y&�\{c�$j�7��ܽoT7m���{#]�T�#L|��G��	�E��O��a��bȰD�:_�a�z����7(5r����2���:��]�)Do����k#!��:gH�}�ُ:��_���A�*�#�V)��
ij����b5��?#�<������AJ���T�0�s;_fkP_�衈���9r����5�FG)G�t]r�z��8%���*�V1���9DtNt�����\��,ݚ�n�ScR�[j��7�[j�Y�^U�1Y�9)����W~O��f��<��5����g��	b��0Nncg1(�5���k�M��k�b�:w�pM���������Z� c��3�s��R�	ul�1%�	n�@w�F���s�7QO6�:��|G�/gR3{���xڟ��� ����}��3�6����"���X��}h�c<�� }������F�-���;��z�� �ªcc��Y�6�+�?3٩�r1��{�4�Q���m�q?ۻ�oܺb�a~tP8�9<�������R�W���8�E}AT�,q�~x�3�(7�����f�Ix0P���P��F�o� ���dl�*	���Q=�Ae����qT���(��|T���o��G8�s�jhn��"-�jϒ!+"�������������h��U���z	���R�LWT�ݽpm����9�-�@��o���p���Q
��U�`���+
�Nt�ȳ���%�/����ņqJ^ +;��i��O�$��z�o_�#T���p�� ֗EI'�v�I��5�R�(��r����T��XG��I�!`Q��1d�|��U��u��zS3��7� ީ�ʿ�ms��S��\OβO>�4ڼ5�� �A���8�!4�;>E��D�`�����_�|�x���i������D����>��j:��Z�"=v�=�"�D��h�
ʪ�g�\��e�[ĨģX�yN�3��~�7�`|8Y�G��h��0���r_F����t�s�w�t���@;�D�ISY��>�������t��c�\�4U:54�J{�Ѱdi$�����^�_���#������ߠ��el���s�ܤ�jnڹΏ�w�+���8y������+rr��~�1N�қ���ˬ�U`�%v��/gΎQK"ڴ-Ca+8?�.5
WM	mEC�����ߴ�"s���Sf�W��*m	3mXs2	�㮬k�ʊ�
G#a�RL+➕UUV�X 2��|[�a�{�Tt�[�q�����m�h�Ӗ5Ez�*�rc�o5���!~>jY��
"�C:Z��O=Q?���kXF�C��G�)ZgYO��J5�"w�� D�{�џ�b	uȘ���"��X�k% �gv�n[��e�>I�l��3��Č������k��^DO
5KOn�Q�K��`C�5�?�N#ͳ���S�I�V|�p��\/Z�Fl�ѕ4���|!#�"�ԒswP�`���EQ����E��-^�iC��l��/�e��<;I��_W��`z���{�Z�܄���E���4�Ȱ���bf��	*H���<I>�' /�EQx^攑�8

�����*|�&-�K�`?��$�:�1�+'%/E��R�(�7�K5 k�(�K�' ��P )�zѦ»C2��ߑlȦ���Y�o�O�Gv��4��}�=�xzٔ!k���P��|�s�4���?�-b��ļ.6[�ԧ%�w�� \�@<�M���#��qЮb9���Ag��eV'Dn0d	�����=�X]&T.�XgO�������|K#��7�lg`�=$�5 �/-��y𡟋��'!�ݦ��H���_��!���U��#��(�P�e8�]j�s�1�f���*��eC'���Y���V<-�/��v�)�?��t���M�0��ڀ%ٖoÝX���(��I*�W$(�H� Y�8��Ս��R<	����jܞ
���~^Q�h��]��/��|��Z���R����ܵT�%�k��S ���"�c��_K�:��J�\gz��f�]Mm�mYy`�|�{,�L��iP�h�I�8���XFǅ�"��>ׄ�F��m��a1w�]�-���ҽG������� ��P�8���l�I`�{#[�O^V�y��U�&E���n���� 4��L�[���y�&��NqK�)�jM���2b�&H���Z�S��q�$����)��;>����m{�И�
n��,��7����ߘ@�Wr[�Am��bSo,?J����~k{#(͉�Z昇� �\��ꮨ��%k�����蔢��Q1�[`ڜ��5Q�Vy��F��a��ctrMx��A�:u7/��?W0z	��d�s��X&!hX���2E��F�d�G6͌�Z�Ҭ��V[ݼ��%��A���/����Dk��&�p2-Z���DZ@�L9w�{�U��UEb�;_^�V�M:��c�<���FqznЄD���f̯K� ��u�����kY�����Lٖ�(� D��}���<��VNRd��_��9	�a>ķ���ҥ��HC�'9Q��WulA@��OJ�ء_�"�ϗ�Ý���m�������Q�j�jX^M�Sg���$%���O�:�Lﮧ��y&&���M_��I,��4�C�%JT+8��=��U��KT���"�Fn����#ÇY�)\�������"���*��ҵJ�ti�'I���״~�v�n_ìK��KÏ=��kª�-�o�ې|�!�[
Д����ǡ^��<���r����d�;����z��()�\j�T��|4��g�	��.�_��@	2�)Oܗ=�����Ŷ�N�!`N��Ux��ۊJˆ��W��0��-A4�o ��1�q���Tb�{��!i���/:c�*�|?�d�`�6�[�@d{�N@5��ӷm1���� ~7���2������@�BCw_�#[pgP+�4v�@�0v�;�	�^a�����������Is��o�p�Er��)m.�VFi?z9�Q-��)�OO�h��b+QC�Pߊx4h�cex�bPM)auF*�A2Ӛ���bv�xHq���N�����I,�OϜ�+䡋���,�M��3�I#ʤe�����Mp�Sѕ�Lg���M����ch��AtU����!dM⹰,�N��!�'�jz�0TCB�fp.]v�jm�0Rg� ?�	��DV�I-���K}�P~s���X	Ү���V*�MU��O��gG�Z3o~R&���j�!Y�ӡ&�Z�I���>(��A��Lj���͵���f	B��Zg�aҺ�5�i�2?<��U�bT���� �0�g?'-���%�g�����W�	o�د�Y\8���[���QO:p�f��<��Ox�uemcs3�D�>�P��&���F��5d��Ӿ����e�`���}L����a9�5��m��z3pi"�u,�YR���l�2���)4R+~hg�-9����OZV��&�m�i�Q���~h�2���ț¯a��a�q�rBY�i!Di$���VN��zj�c�k}?���<�1��%%�cK���-�j7|�"�d����֠��Q���SӦ�����Ƴ�*�T۫X�ߏ��猪�,�>��4��8ɖ�ؤ���MH^<z��9c`ҙ/�hOa�aZ)�k:��+� �$}��|&�i1��C�h��m�@̈GK�)Cf/��g�;�5R[u���E~�����P���vD��_���X$��TӴ���#S,��H2�e�~�h�:|B��� �d���=
z����Ϗ�N�\̨�:�6�`j��5�BH�st���[
d�f?�*�vҌ&ÿt08|�1�����(�2����d(�CZ��7��eb%�; ���3�'���qQ���-D}���B�y[���3��?ض[p�������
�sN��?J�sdA����堽���*9W��T�	Q�#��z�em���s�ͽSi�� m�'��M������ ����]b��tkoIV��-1�O��ts�v������!/�pH>�6�UL)=�l2�"�
��>�\
���!�Ġ?�P#e#yV]���I[�4�4�0h����m#/�m$q�/>��=���=�{��n��q+�[tO@�q@�\�����%�!�����e�F��֊����8l��>��pn�+�c��<�KJ~�B`C�3\��Vi����m�
��v��9�g��ʈ�':Օ��"�4�D���q�}>��$��iԡ�	լ�i���lؖ]ƆA#[b�~��ƛ�C�(���HU��!\��K#�9�@J�RV����Nfe�+�a��K��3�1�v�(���c�-�֬��H�q�S[�o�.~���
�����=E^�q�T�<j G��<��R`�����9��|�wf���C� O�������$���AX֥20��Υ����Ha����ٲJ�&�ۤ0G`�ŧ��(.D�@�E/�6({4�VT�Rq�%o�L�7�}��\u��}@Fn���u|��n��p�Z�6T�N��2Lp#�mO�)����T��7�e@/�"~M{z���omĻ*��贶��R$�kO��s)<����2T�V�f(5��'+6�<0���?u)�6äG�A��d�6�;y��^R���$5�X{���>���z�%�<�ݴ�Jy����]�Zj�2���$w��.-�鬷��{c��s �8����f��ς�7�nИ"ME��j�҉YT�����y�LQ2GԠ���9��J3)m.�4�DMVT�P,iAC��傹��vR���z�t����g�>�V�"#"�A<ޚ��~x��� ~�� ������YF��o�f�US��܈��x%��7V����!�fv[zx;�� ����ẍ́1XRD˰_�ã'�YRXX�32���! �H}��e��|�d�΋X4�j;Ŷ�b��U)S?4b�k�=�i�C�m=_��7�����Y�N��Q"�KNh�%�@�	]�V6�E�7��b������}��u��]�OR�z�Q��5�~���:�k�z� ���v��>s%�.�-���d}��7�F��SF��f.���7.�	��k�2ON�mp�qc�D�S(e�P&}w�{����wzH���Z�S_��>-߭��ECz_�)�6��
})��y��L�l��&c�Y?.M�#�n�{(�C
�e~�i��I*���19cSw��k&2ѳ�W���*��3��MsL2̏�����@5�����0�c������a��;U6'$���M�kt~XIGyn^���C3�ޟ��*o���+䊐��=���n�JX��vFi����� ����- ���[S�g���ӫ5#>M��v3Ȋ#iĆ��Ƽ,N?���ǔ||԰���^��Af�gm�滤�!���Į~�!Zk�c!x]�U��3ߘ��3{�[7(3�Ÿ�)�oh	a��bw��~��Fu����.k���X��*,����E/�!�b��2wr��PDh�h���nkr���������R�6a0�'uY�N��#o��9��D~θ��k tBn/�2T2;׊�� ��,��h����&�g��Vpd�r��������"?PzX	|Q�F�ahi�X;��N����D�x���O�AL�gl�r�����O�B�aj��̐҇�8�?	��9@�[J�N��r��hO�9���e8�
1u��f�b����Y��~<���!h� *�W/��6�n3�#�ԝ��Gf/C�q���SI&�����F
�C�}_	��ζ���f��µ``��-�
 X�Z���fߓɸ�Z�ex�����o�H�l�����/��ѓ�k!�g��A�C`̀�@;���Dn�<s�Ex۶RN,��>�A�X���K�߈+L콞�cr�a�S�FQׁkҜuw���5�r-�Q����MJ�n^h� �!��%���{�%� }��
����вP-�	��r^�0S�(Y��u�tЩne(�O�O|�=Vxh��>!�i�{���o�a�OD�#��e�����r��֤ڷ�4F]4�7gн"g���SC<Jg�O�N���O��&u { 2��<eo]ѻ.�>^��a���kU31 �
["=�֤�l�\�`�������b��|��Cy���`�ѕ/9����*�Z�V�,�_0t�,�2q״�gKHnG/���'5�y:ҿ�b�vr���;��)-�Ig���7fV?�-�W�<��L���O��g�4͉xS��" 4a�lHȐ�C���9�'��=��F�U��U|;��'�o��h�p�F�T��a?O��� rK:��d���ve�"HB�b�x����t��t͝��U���/EH�б�U��-<k�R�I���
��������&P���Yq�� X�੕MG��(�>��`
5�j[7����b�����)�~��h(ШG�{"�}����'�[f�K2�4~%��'�&���d��oL�R�{_F0�s��u�\��IY��]�jIQrޕ��di��e�L�L���B �TF�x,H�ÇVN4_�E���0�V�˻"��d�E,=ܓiӔm�E	���fc�FJ7 cv��#I&��5��AM�Z���#����)2��op�4��K,]\$�@$�>~*<Ͼ�&y�e���q׽X�x7��j]�%[�2ߥ�"h�ṅ��ۍ���}��a<ߙN20���=��Q���"���M��[���[0�}��\\���	4Y��Z;�7���+b.}��=Q
������e��4�S��@�v���r6ٙ��A1S���MDȫL[���jp*�ř��D`lN���k�\�l��T�s�	���ϣ~���gj���=�EU)���[�(Q��ȨŢۤu-�����s�d��A��5w��O)'���	+2�)��
�bA���X�-�b��;s�Ԝ�k��Ū�'�$��~[	�(����"�1�e\�΃]x}׊A��E��ĆF%�%���~d�k��˵���:T�%Xz���x��r �"�Ua���z"Cߵ�h�
��7�-)�*s��l���e�_�o��ADP
V�ź��hE��KG]$��#"��a�����cJIi�YʬV��[�i$~��HL��F�e6����`��J&�V�!ӭ:Η��(e��xB�:2��S-PO�y��Q MeDZ��-^�O3Ł����;R���6-=%!���e���(0���s�����qD~������G��o�_�����@���*%e6v�+~���P�"�g�8��,E�u��%��!�D��$�ҋk��y�4,Wm����X�Gs��:g@�Vo+Y���s���¿�'��Wb�.+Pw����$o��6߽P���%	Te�8����G�v`$)jɄ�+���kL7�v�ۻZ}8��B^��_��lK�lS�Ҙ/8Km�4I��7�D������:�00h%���/���C�2P�/����;���ARn9��;�>A��f	����	k>�D�tl�G�}�a��Z3�F<�Kp|����6�N��p�i�g�����Z���iL��BC��	�ȗx��JCҙ��
��ud��p7l"h~���N���N$v/�8&�|�W�9��G��`N�T͜ѣS���Z���)�(�T�o���uz�)1!ES	�:�`�Y��v=k�-Z Ԁ7�I�v�m�)�DF
V�5�Za��\�5��R�]�/��f�J���Vqj����\��i�5�i���^��1��WMn�S~�s�!�^�����VcVs����`����=������Ak�+�\�?��C������>B"a{�Z1.��)3�:�'W"��z�w��+Dr��o��Q:���@%����� !u���ښ��ӓ�~=�%�*8�H�Lբ��U?��$}��XS���;>����І�
t�V`��������YJ�]�w��i�g��4��xS5��s}N��h��_��tP��c���y�R���Y�v	(@:���6y�	 �pD�E�(�U�m������q���S�̨c�֣���8�l�E����fQEYXM9��S�w{��5`y掂���ø�2L� T���DA����Z���D��GRs7&�c�k�������)i��㧾念�6O�+���+�$��k�
C�HR�ĭ�s��F;+��Aн5�s~P�A���]��֗���ל�����/��)��3�����p��?ݻ8��:g_�?#|Q�DdiD�r!n��bWNF�Dx;��\$��hn�)���T��%�A/oӳ���Fꗅ�^�+ܡ���|�s~�������uP��4�'��=��;�0�Ț�<R�p�kб�#��N�L-��.�c1�bfE��=�C��Mh�����8 ����J�#6[~�Dcz5�/0��2����M�b�y,l� �C:��G�G�����25O�	�H$�~�INPy�6DKdS^$���q�K,��&KSJ]��:�=�ή�X%��	�����o��o,�MQ�MO�~D\=t��6ɼ;�	>_�?�gҞ1\o��%�&) ^Lb{���H䢽�ߐ������{��C�YbH�#�k7�K7� �p������~�D������ǂ�jk\?����z2����O�7x�g��QH�� 9�~�{G�i�,t@�n�ok�L�`��w�U K\���渮J�ׁ�5�zAܰ���6�"�����$Ǉ#>�h7:�g�0t���_
kSLtE?ŐeTo��M�E�)�h�~��S���Z��CJ�&� �%�w�ɤ�B?X&2���(n"�z����)qU���p���6M�3��vc�WT��P���1��w5O���f���{�#M���cs��b�qqHPpޕ���c�R8����:�h\�'bD6:Jhcw|j�w�%��	ς�o�BN�$����M�Bu"�AMB��+��F��]͌���� Jb��2��HJ5+.B�����%�g2e�y�qu�C��0ͯ�^�o�6n��P%���F�N:.<
�+�Vph����q���	��E��y(���z�WJ�f=�IL/�dtoa�����I&O�#��	I
i��˖�1��3Z��
+�q*>6�;4��� Էn�÷�#�w[F$�͡��pt9d �a��Q�N�4(������j���̿��N���ͪ�?�1X {�~c9���;����;��$��*�>�T�&*K�3(sZ�ż���=���W��ӓ�L�σ��W�]���D\�m2����4�g��@n��Le�$�U��b�-+
06�Ƹ�l5T[uw�|q�g�.G2��B�W�5�U��ڧR�4(�)5�ً��7�ј��PKR�)����1����k!�ޞ]B�+���RI7��3S^y�֌��	J'X�fQ�n��(�2U��=�XRgok==��.����V$����zC	�������W4���m�ݟ��`0-�eo�*IbAw�r��ܽ��G5����ߤ[�͑B�:�kf�Ks���>�c,f��4�\,Ȟ�>��ތ����o&?7��eevxFi�����;��&�����ٵ���(���D��2Ȏ���#o����0��TSfU�;���xv9w��W0�MNb�_�6!���d�����N�.�V!Ia\2D*�wd�Ķ�8*"��ni:�,����? _���pI^�y#��W '&TJ��gZ<�tR6k�/j1��f�<�*�g"����x��X�:n���y7 ���s� �r�E�ᕱvC�����;6�NRh]ܤCv�Ww�'��klK)��PC���_�����ي��PC�<H�v�i<�t�j��g(��T��ox1؅J 5<*���`sv|�qH�T���FH�c7��#~��Sd�X���X�JbJ G���3�2��~&J�wC��@7�G����eU�`�I�r�Vy4{:�B��:��$O�i��ov3�V�{U��XA!�BA'��J�olw|�R��e?'7�C��4���_�Is�^x�Ӫt�/*,
�_���ƴ�{W��f|\~��U�EU,𷦕��T7�߿쌞_p�}��Y7��+��Fy!�u��Β~��D7�[8Z�4����a6�UJ1j*��[ U=�&��j����|���Y��Q /�^颫����᫛yM�����fC_]33��67�3&�.0@�������g� #vO5�g���Y�J��#��{�Ta��_�D��T��+i�0���E\�/V�"@��d����܂v�w�p�G�`3�,�@������s{��}U��V�G��,Uw$1�O�Ʋ�<�I])I�c~>�WE�C@����}u^� P�P+�N���}���5�L7�'���}T�`ڦt3})x�ۢ[��q�ԑ\0Sz�Lب�p,*s�\:p�-&�\�S�K���>�-Ү��d��]3]N�����&�{�,{u��rގ!$ފ~��jF��L���"PT�3�&#S�*�!��P����!��}~i �Bv08�E�������J:&�H����r���{��QB����c�uв%�w��ҷ�&ʆ��
�*��'�`:�>#֢Me���"k��EX�}�)���S-0��C-�}];�������[�@���e�-+!�!��J�R�p�k����! ���ױ�����T���/!��t|��Oq�����Z�"X_�u{okL&,*+l�MY����6�j�A�-T�=km�>c�f�:i�r��|�A����A���EΘ(���I� ��%C�	�5,H�s��^�E�<��H�8����71��_+O��ކ�H�C$4�>�;��q@�%����# 3P	G�R��=����b@GJ������s=���F����x�M��g8�-���.���yR+��}��h�[�։*�q�a�#)f/��`��۾��󵮡Y0_��q��R( ֎�������U�^t�lt�d�K��|��%�x��ʤu��1Ѭ%=\��J-����K��3�,��w�$͙�Oz]���PmbW�\�T�.T���8b��8d�x bY �؆��������0�B����_�J´�X�-��Ҥ�GUyQс����Sܖ��wJ�^��4$�,U��s;P�d/��?��R1�ݭK7|���G_/v:���JK���n��U��V��YS?�V8�K������ʹ ���
�ERdZg�a�sP(�8�G�;fG�%�ۏ��X�=x�AW.��_5���C�2�Ю�0��{e/�`/�~i����{�J�>�Rn�jw�	e���X�z��[v]�1���f��a��v "�Ӷ��]A��.�`�ơ�U�4�K�3���yŴ.H���6�f�h+��I�r~�zlW�E��(1�{J

m�oު�7���"�ɋ2E�.�#�����*�~ �Z<_D5bZȵ04���Fp��t+D�13 @6��BR�D�a	
brzH�I��'����Z<�y[]�]l��3�"�U֊b�y���$S��Boʢ����:�$����
}���x�3E�/K�%���X*D������q�T��甡3|G#{�T�7�cD�;,�;���SIy��\���M�\���H��l<���É���;q�%*��B
���RN�n��h�JEG�U8�Fѡ���8ܲG���_�kh�?y2���8�!)Ö�Wt|֜ٯ9&˚�eN�A�"�F����=��]���Q>+&�<UBa�@�#0g���I���|��_�-��.�$[�:��1?>���W��P�R�isb�{�
�e�)�y�A/5�@S[� ���,��êU��������YND�2��Ǹ�fKN�cVr.��ˤ�,A�L�5����魊�%( �O�N��U#��]��?�*OEeXD6�M�t �ߟ�ݱ���8�m���xvT3_l��vxs�[�Ӫ�,�_�U��"]Ez��J����߸6�r_�������0�	 v mwo�?��u�W�r��[�66��>C�Q3s�| ����5�?EZ�x5U�ak�x�g2�K.�<�a���ѧ�ғ���%�Qdf*^c	����s�E*��0����������'Jb���'��?�&���(� #�<�1�T��;���/����X^G����V}F� N���ϗ���ի���<��4Ť���T��(��ZI�^P�oݲ������zU6?���]�B�*5	Ԧ�x�֬Ĝx���*��2�RR����w�^���`9�1DL����U�1��_ ȿ�(揰. ?;��av�I�h�1W?9�"�Z�m��=7{q�|km�ިF&n�+$�������^�Jm�H�c��F���6\g[h�B���ϺBf�&�x��r�Om�Qs�K�B�g�&��<��c����09*X
�ew\��q��Vk���}|��e-�z����7IO\��ƟA����$�Htc�O<se���V�j>���t�@��Hbp��D;��d�����M2�M���(k4Z����@G�:n�ī}�����+���e�ڨf:h[%c��w�ɋ����/�T�W^�U�W�F2}{�{�3Pp�ǅ��JE����z[�3���4L�}�Pv��c[� Ҩ�s����
?Y��g��U��\"G��pIdD�A��0������X1�H��ws@�i:c1����sX�Y2��e�D���U�Yp�T[G��p�;�������»0G����N���=�%����1/鲔�-)�n�Lӳ�N'N'Υ�h���fI��״(��M�J��MLG%K����hi�j��C|�B{`�kS����b�_"#۫Z������l����:�����{��w�=Vf�}Z.@��>��ݵe�ǥ�����lX���he��XQ�����`/9��oYŴ���z(��4�1��Ϊ��a��g�j��}j�Y���>9�l�����Lp_����cľ�ď�4u����bW���1@0��hpZ���)D 3���{{�\-�����EU�M�񔱔��Vfjt��r�VC�]!{�!��(��RPs�c`I������z
��f��q^7�v�G҈z�:K��+��h�����҈a��3�ʺ���%���|�ˠ~R�Z�� ���A(M%2�`q!�4�ܤG0���J\�YL7<7c���!�*T�_��)�	b���C�wJ��;����y�A��^�ȥN4�v����3u��e~ڲ�~s���'�/��v?�82��*����g�B����A?CkĆO�G|�o�Ry�
	�xZ^�5��`[�Ě/f���}Z=�p�
����|_�o�e�|�p�-e�����6���O�E'ۃ��B��{\��92m2<�&7�,��b���$��֌��Ը$W��`;S(�~9��7���!L�qоc�nq��&��d�&@��k�i��v��O3\���m�i�s�
�~��%tM�Lkg3��'��E�g;����L�'�$��"9�W!�b�m��/e�c������C3�;�l�q�qC@�QD��mG3�-2�����>G�	��!p7��k��>s,Uj�j�� �Kr�������z�w ���h>Ѿ�|�ۡ�Q���lV��)��S�~КiА�SzW���3���y�磒pJ3�>��g��� ��ȝ��HtH�W���=΋<�C��*�&C���ٙ܉�S��W�WD(��b������j.L*�v逇��S"��(��c�h���᫢�����%���s��㿡��eIxҋ�/���ٛ���� ���.��=���W��Y�%Z����h&��<��6�RMɸdUw@�G�b�y�w����t�.-m���������Yz��(0cY5tC9g��@�"���D�:h�i�앾��w���|�B�2�+����b�M�k��KB�jɛ�BF���.G5v�vڋȕ@a����2�j{�f�ִm�Sms�P��r��P�m�5x�L���$�?,�m1��98�#��V�W�vl����!4�|�9�wJ\S�,p�y��P9����%��\������H衸�	��d`8UM�ΐ���,
D�]W�9�5�g�>��� d��go�wv��2��;�����S:&�^J�V�껅�s�4F���<@�D�P�L���=Risq	.&K�|y���G~1���*@ֆd/iH�9U{?�1���B*k�|�����I3C�Cs8�U�>n�E	Κ\�(K�6t2�ײ���&��m�wH�'�e��^Zy�(@Zs:�!�Z�.q��}_d��!�EB���獚8�o����,\2��F�0x)
q]���ҝ��d����_<���t�Je�R����ʇ� �ݽ�gn�Z�b;��A~gJ�#LV���F�-}����@ON��a	��X� �����h�0�[��NZ����_8?�m�v�����jE8�l[< ƴ���e�6����|��bU�1Ȣf���"��nj��\N�o�l�su[j5��<�s�s�n0�W}DgSꇡ-����73%����]�]2�0,�r�?٣�ت5cd��w'�j ]�� LX]�j5�������C�]PJ��Q�ȥ�ˍ�=�f�ȥZ���Q��E�d���뀘M|�xZ��3�8�i�����>?��
�A��5%[9���1��O�=yw'�нt�5�>�@}ڔó�"(�NC��hLߛ�P�&.��E��Ol�+��<��
V�) pj�D> ߴ</�j�LHg�M������:>�w���<Y�穀K[A49h_���q#��dY���Au
�mp�lW �3����`�������
R��bF�8���&ڔ��ʑl�X�WP�1��Ƽ\�d�0���|^����]ҽFL��-��.��:�#������h�0$����T��doy�&qqdM� �T��0_��q�.���l��`�X�O��u�p��D���灄��#u�@χ�C���ϐ8t
-N�C�	�xx�	���".f�V�>s�0�8"V����h<׉�`v����I�Rf<��Ĝ�@�-׮�@<3�q�2��u�T�.�02F�j���k�j,��f��da�@oD���1���3?�H����3�Gq��M�R�1���.�
�,7U�鲦Ӷ��.�b�'K��w��d%jݯ!�x��~19vIv�ْ�-M#/�G��+���E|g���|8����< ��S�F��&��>[��w_:~��	��o�iڍk�/��H���J��w(��,q�@r�~U��� 3�$$F:ap�>:��.�֍�J�h����)�u���g�Ӂ<�_�fa�����c����/���dQ��� ���n�ۧ�e���h�<���x� ����X���פ��2�]ʠΣ;�)��%R����2O���)3�[6�1���Ѣn��C�<���a���hQ|1��x��Ww�������O�E���]�빀K��賙�a�V��Ǳ:��2+������A��r�N)_H ���^ƹ][^E>4[��D���u����A�&�H�ЫVH��]�G��l��SM�R�E�v2�U}�	�j��p5N0ˡکǈ'O�����͂Ƒ��<�����3�=7|���+�u	�+G8����p�c��|��*��!i:}/t�*��KW�.�g,��=�飣��Uĳ{�%jQ���ܨ�۰� ~�2�I�x�K��pP沾��,�������2�l*?Ґ�^MF�i#���1�*P��8\�ڇ����Z��!(���,��ԁ���E�Z\h�#3r*��ʱd�����B���O6���F{����M/�Є."�����J�B-?ev��Dt&���XF�X�~bx���`=�ٺW�V�u���g�J��DڛF��QV3�'�[4	�p�YN�`>%�r3:0k,C��{^�4b�H��/�Y�dw�v����\����!d�>-*�d~�j���5]=c׿���"R���K�l���-fh���G�,A" �d��K��S�	u��$,�XSS�=��QŅ�힉%h=^��e�,��q�f���)�������f���{ٵ�?���$ݡhd	��0�3]RK�6�N��>}�z�\��K���kC����jy7�=@Bn�Ԍ�V�{-:�
*��^:.�#�����NU�|��=�:�rn�\�E�|�g[V���cf�3����aO�^�tb�d�6�:���B}&��$?�3�{)���x)t��7WH � ��q	>vƔ5:�䆲Y�n2ъ�G�_��B� �8�j��1�Ly�I��]���H�~��R�Ǘe�Y�Ӯ��6E%��B�F���ڭ�<��r�p������VI�l�������i_x*��������_+L�(���li���5Y��){K'�K�{3�dy8QaB��#g�Ϝ�b�gxJHǌ��;�{T�z���"���奉=�#�t	���#��&p�=Q�J�i��q�5K�$�'`Źau&9����7){�wI�8$r 
�Sn�������G�&�qt�i�/��_���[���}J25��6�!�����u����Ob��|z�g�E8;B�B[_'����ϼS�����Ɓ��m���Z��?Ř��2�(�-���(����U�aN|i�Fi��]������� C��Tn�@�v� ԫ���iOX�G%�'N�����^����[ykm`N+73�7h2��7L/\e����RI�äV�"ziA�)3L�K�%�i�@c���4n���yt+Ln{��oS��\s o��c��-Z3�,��7�S��W��
Ff�#�����
�4ݜTW8/#�NKl���%{,�0ǂږ0.�e�6��t,A�)[*�58�ƀ�`��OO*�8{O��[���������rs��o�H�u�s�,�0G�_	�|���S�t좎��P�\��n����մ#��F��Ӓ���3�a�+�k�|�}����m��a5$�L^�_ў �O�I#���nQ�Sq}����Z��2x`��A8k�r�Nj5���HR۸z�X%��C��M4�$�Ff[���e�p=�-1�2�z�\U'�=[%���k����ͺu�b�p�"ݵ��l9ea�w}�O�0~����ĭ����T2���1e����/L_T�jEE���;�S,�:���;Vs�L3�ң;3`Y=���'�$�P�� @�9�Dr,�����+&34,���u(hT���(cc��R��U��#��폭���d!��cY�zZ8ȧ���&�!�m�U�5ge3f���!)��P���ֳfV���)"!(�$�&������d]u,%F��'u�M��Od�8��a�T�b�do���w�D�Ĉ�C8ڀ�IS?t�4�!=|�%w��eL	�ѲJC�5k�nwJ�Y�� ���,�\�k{dja���X=�q�Ae-D�Õ��s(��"*C�hoB~���|7�~��@U���%i	�js!}�i�zw�U�b�aJ�!z)�j�V����V�7��G�$*�;�|ѥ�������]W�ڶFXG"�%�{��O#-�%w9u8���ɝ����������	����Ui�xrm���A�'�w�U	�p���\C�FW�n�+�����%DZ��O�����u'�$��XkA[�sG_!���,�e�9����>|!�gu6���ġf���6��$�sP��az��tv�(!Rs��:O�m3�x�RC�Uy��첹�|6�ܘ%��U��|��zk3�����2; }���ɺ��o����&�V,m�;���س ��N�[/�Lz���w��Ui�&ԕj�x	�ͻE�4��!&�� ��B��$�b�[|F����!`��������/>�F��lr���j
�g"m�����N�uO���ֽD��H�F�ѐ�3���9�q��w�]�]"_К��Pp>�jrV��:��(#��  ��(���9y9����x�7~����U峸��x�簘�&�&Y���Ѵa� ��co�kR�e/��g�9�v�����#K휲��o�) ��Z6���������qǻ�4?�fʴq����T�'g��V:n#�}�ե:��s:������sr���zN?쾾��[������4�3����_�r�)��]�N;/⽂��°��c�a!|_�/����J�o�V�XfORZ��k�S���5J��/�d[��2�������q�y^	��`co-^'G
i|�y����Lq�[Qt�����l�q��"�1�[h��z����.Cr�6!�*�ĎA��`mϦ[�'��4h� ����Ǿ�+�v�"B7��z��,����2�G��y ��麛�7���M�"93۽ޖ+�X�f�N��Q�~_,	\L�p����r/v�83��BF\�O5�K-xi%�xq��~�p!�n���R,��%�Gf��˥f����07>K�t��<��)_E�?"X���P3=���$h���Q���V�Q�d��?��.��<`0L�Aaצ�$c(���Y3^��I���[�?�d"�����n^����g�����r��9��SpJ�W�`��Z�-b�F]�A�'YJƵw��bw[tI3Ĩ���TB�V�Sk�ݧ:���ك>�vU0��\3$�E���H�7���[����W��h�&��)i��B�����c7�mP�߫A��?��>e��<��#T`г��V����E��nm�l!�JAl���8�\a�ç�Q���c�a�Ų��m��8�#�^Uvc�|�}~���V�~�λū���u�aA�_#)�oKm�c������TI�(ߚW�a���P��*�(�!�7Gr��ŊS��x��U]�|]Mv��O��R��z��;��%ږ�/�?}��+�M1��:��onRer́�(,���9�T�Hi��D雳�T��q$���V[�T3r���Y��5u��0�,�6����9��b��5�&*�p��D��3D��K,aȋ��#��?�}�������u�9A��� ��ޮg�����j§�ij6�f��e�.�&�%��z�4h�rY{�:�P��H�!Na?j�#��2��B(t��G�@O��NB�I"	�d����9���܏��"R����Yq�f�S�OＡ;���I�t���,�uR��ݚ]� ��V �bd{���6�\�Cd�2&R�������U�^�ϸ��7Yd0��t-��Nfp�rg�	@�T��0���Q���n�/��λw1���L��u���ȮYD�%j@���&�w��}@�%�h\���s�W��k#s[U����s��Xp �N���d]��Fz)��v`+� G|�tS�<���E�bO�qs�H}�H�?)�D�0)���c�1",�H���s	���Z5)�Z�!B*�jȆ�sy��f��x6_�	�LE"ڛd@U	a�S^7̚��L���(�DM5�(�q�����j��uj(O�Ç�	'%�BGstF<u�4֢����={���a��5@�l����	E���{�9x���F����3�E�qI�Ժ��@��q-��Qǰ�yj��+��\,]��˽d��dZ�7��6$Z��@>V*��}��Gؼ�Ք�`���HQ�ӱ`����v.A^*"��K����u1Vv��E���q�u����� �v�5��#�!�HC{�Ϳ�!��Y��Љ?*�7ER��&�$]�K���A�c��q|;"w��I$�j�d8�V�N|�z#�hǥ-[���_��'M�S����b�/�R@���2@ ³IW�l,'�wQhf�\����ב���	���2�5�(ܺ��O��]Z��Z����WH��nM���2`ɏt�S�����YH\ވ �ڈ\)}��#��w[�~<�
������x�q1qp���q�����%��S�'MZ���ǘb�A,��
�9 GD��Z)Tv(���S�2�B���	����"~666d�XGUl`Q�	�r��d�Up��'r��X��B^$�|���1���?>���`ͣ�7/eۺ�91�Y�U�Ug�f߯i>)�g_9�̕�X�4����ѧ{C3 �Ux�th� >!�;d /ԏ�P����{Ζ�wη�{C�y�N��K09H�-;�o�S�Kn�5-���MT��}J�����ͯu�%3Ɍ�/�0%	���n�&�خ��������-��={Y���Ok�û� ���k�	ESN7���a��Ħ�YR\��e��k 9U��p�^��@QF���R���,7�S''-��Mk���1u+,��F��J�x!�+�)�c��y����Q�C���ЬF ��|�Z�ȭ;�3�ݯ� z�$T�N�ot�m,�6ۆlE��$�o���wI	�Eh�FG��}(Mhs����r��
��W��9�<oEv�P*�@��^[v���<G�S�����r��=X|�m�����>[��E����U�������>\��IŢz�/��� @��e��}@���(�Ь���>��_����'�0�Uځ;�L;j�|�v�X�,�����_�:��F��
V}r�|e	p��-�6R#@�!��鑀'��!Q2�brN[��ȑ�J�
�����ϛM���D
�N����64gҌ�l ��mKcw�RSsy���n98�6%�'q��ϭ렪�c�"����;o���2��5�\Cq�Q,4ft�PQ��J!��a�KOUU���Fgέw��q�=AmR�s��t=&���Y�S�+�jm�{�6G����!M֠�0�˩��1�ѽ�Б7MOa�4G�n���f#N��]kuG/C���Ϙ̎j\�:�3��9fH��iϼ�?8����F�[^L����s�ED��T�k�1G��^�$�*�����#��'�Ab���`�T+��EͻiE�E�W`v�%��?@I�n3fg�������`�"e"�����ԥ�i�x֭Ar��������αr����`�3N�5;§Sc�$�X>lA-�(��U�Zy�j�3�Ĺ̃�s��2.����f�����]�gn���	ю��l9���,���!��\�b��680�$+�$���Ő�͋�v�赙=P���Z��f�`���H�e�5����= �֝��xj�A��`̙ʿ��\�{��m';/ߖ�ğ*)4�\��_���}� f��?M'4�U��p2��ǿh}�W�1�^�	�jrͲl~~��W�|���-�6���feU��xS�x���:} T`3�����T�7[~׭۪Y�q��d?ȑ�Y q3M��N4�Ӱ,�=��'аJ���i���bGЧ ���\�|'ɈC�h�a�@{�Iן����e� �R���o���-�2��U$^��=����T_���(���q��$����L��i<���3���A��,�5;_@E���3Ae�*(�0N��&D�A�^_��B@!�5�*��J*�-��P��t��0���`z���^�N���{뱶��nd�����\��7�UC<K�g_���V���B)�qݿ6N#���~���~E���)��1��ټ�N��Ui~�9)U@�zA���'�xHB8�c�r�gS����~"���S�/<�d煌����/���]��T�gP����B�%�HqX�?����BD ���̜�6N��fa5y.�f!�r��"A�&�[��V����$��sOύ����wĲJ�O�А@���mz[t>5�=������E�+�:F%�μNuzΡ+m�a�lxZk���v��6lK]~\�p�o5��Z�8��;Tl���'c���
��Os�p7��Q��H�e*��Dѥ*wp�©E���6�*�2s�O�(V�P�)6Hð-���t1���j�Q�L�F��P������v��,1�5$a���d�S�-]��9,�[���k�B��|�}��hR-@�P��!�S�@�%�vm�*U@R��ce>�,ĠKkA�6��Ia���{1q����aFW�9̳޸'�i]��UNl�$$C2�[�+�h۳.9��
�+�7�`�5�ď�#�k�V�x�ς�'4�d�~�q4�T���C�5]��R	���t����./ �J��{��*�s\lk�T�tj�4�����/�l�s�xuw�'�C�(X�o�R�8LHK�"���y�"82+H���4�Z�>���"�z9�������4��ْ)�������i���3Q�}PF�̬F2���$�XЦ���{Km黡Y��A�W����Ta��k�1#�4A^F�����o����Mhl�=�|,2�F��`k2��p�F��R�So��~��`���h�[�-��/�%��*�ӵ�=��
g�Va�`���CuxSǢ����)�JQ�����^�S=�:`�趞hZ��V��� `b����-�}�$ȥ��Jw~]nۑ�S���&����v���6FRQ��O( �E����.A.Ia�e��d\d1�E,Ʃ��}`�����`�ɐR3��LcY=���	��Gi���͊QY)u�.�}�iif���_��ǥ!�����8�U��=�_�eZ$�t;%�aF�u��������8��k+�ƃ��˲`:/#�m�:px��[܏a�|b+�c9���:����f�v[��H��\���!@��ֹ�A��35�8"�͉���� ]�K�P�bBo%&b�o2Xnkh��:�;2o���w��\�UEÅ�0g�he��ٶ��a.�Xj2&��x�x�7?���=��zغf��b\�,���=_��Ӵ��(��?�]|�]�6�M�Ϯ�(�$���VFѨg�K������r��N(�Ǻ�m�OT;ivv�'�$�ڿ0�<�^/�l$\�ԺaC��z�Lt �N��j^��TM�<��4��t�0�I�05Q^%���ǐ0�`Z�ٶ���g ���9��yct��7�@f��3yD��UҒe߳K߁6�0=�KX��iф����@�Hꍐ7�ͥ\��{�P�*�wK�b9���Wf�̳EG���g1 �,p���]6 ]����9r�̕~,�'އ�&s�+?Q>B]WM���+j�\����Th�׾��Ք"���|�=	���z��Сt�tZ�N����t_/��ϳU����j���֍̡�F�!6�0r���V��b�7��[�Th
x�r{�u���Nk��P�֤������זr���K!��7��ky�qB+�^�*��x������W:FC��̶cɊV��h��$�n�R�[��J��d�J����~Z(q횮�.V٭R�K�|{ �������L�5Xh���n�����/�E�������oX���i�rA�B����	ъ���Σ��[:�I3i�%�:��@��E@�?x/��W����E~���+O��{�g\���1��]C����'�����.���py�| "��<���lz�%n� R�%��|�r�@�����Y5[ҿDp�r�~�X�~�Ҁ�r#�j�&k^���l�+���[��y� ��,�=!�����*�-�6�������sY�$S͖��3��3Z��U���ۿj³��;��)�,����{�D�T�Q��aAG::h��ϊ�|Q��(m�����=CV<�e5# }���"�����y�,7�:	�S�ÿ���گ_���fx�5Jo�m<�OH*UY���vl=���>�o��*����~�4qdw��6T
݀��o*�齣�x��g&�t��n�-�W43��h���XL����Ρ�p?x��CPҭ�=�^�����o����p=�[��Ɵ�k��
/x��_��x}e����${� �%���FZ؎�i#.�p��;Ċ�.�|�C63R���wa<V�3ĭ|�nL�8��s����)�8Vl������``"�����9�f�[���.���a�LIW���Qf�g.r uk���@�9�o���/�Z�^H��kf���W2Hy)
{�-meQ�7��O��'c*��_͹_��58訢 �R����
q��S0$�[Z�b����{~�2s7ҵ��g��.V���V�t�5���	.R�mP��?�P:axEn�g&���u0ewH�Z�%�`��;��[5]u����i6n�9� sâl�&+L �e��s������ݼR۝s��܀<����������(�8k^��u��$���̾�b���%�i��?��lڜ{�enj�]0��`(^�/�J;W��T���8F��A�jQ�ʹ��t~y����>�c�����ʬM��-O���j�z�����_�������8A�׿V$f����)lӿ��\�����h�|N�^�݀�)VP`O`y���C ێ0c�[9i���x���	��<o�CPU���VS�i���wR3	Zw����R���H*.Fdg�u���PӒ��c�x��a�~)@Ɍ
r�KMH�v��8���,�V�s��n�������r��(Na��մi����������&I�>��(W��l�u�ы �K+�Y��$�1�'��0N✾��w�ҳLs`�T���]��d�kNO��i���1e#ؕ,iJ����o����j����d9X�3�}��_!��It��+�S=w��#�������+#ߨ�D�%;5JD�Ac@�´�����Zv��?�(H����<�b�Y��mծ�:�N�y�*,��^?��P����v>&�`3k|�:B�D1͑R����6j}��j��G]jp��tax1�a�j<����e���e�O�q�]ҘU��K����ťWIz����_�����I�B+�[j�x��x>4�s?��͎�)���.�H%穨f���JD��}pK�{�F�����G����;V�ާ�*��B�Vq3��oǄ��/4Ѷ�W`O��`[��Nn�ZG�E��x7���xf���g3�l~b���D�>�m#�uJ���m;U���i�������\�u5�?N&2�/���M���Oθ�Q�2"[P���T���Ш�m�ZҺF kLL��h(�z�V
�$Z�¤z<�R
A���m=SG�/:]��"�ÿRUѰΖ�$����=�a|'/� +��do�zk�j�=
te����{�.gpu"�b��g�`���lb���^�NH��Mj ��qv����w�pÌ������ܳKkL�:��d���#�9&��|�:����,�1�$�[,U�o���F�,�Or|�M�(ܱ-���v}� ��1�i�^���▶#�Sa��@�=`3jȲ'��7瑚C.]���M�笀pܯ����f�_�?Q����`��9r���f �+��ӵ�Zi/p�ˤ���\�53�OL
q��0�ｋ��?<@�|P��j��åi�2/T �1vȧ:���Y*F���t;��k%��rc�)#v 	�y�t����]+�e�]&z�V��%���yh0�2eh��0�Y�.֨ڗ��4���\�)N7�ܱ�JT�p`Ίx\F�{�׵�g|�.K����X�������Yix)R,r%_�xF;�H�hUо�P�M�ᨺ>�����|�Q�-	�5[���k�r��.N雌H�v�9YfХ���~��L�K	�p}ԉk܃�&�F��r���f���Qw���Yob7��o�W�R�8�ͷ1�I-��|��F֑ ��	:RRS��ԲG���rKqsv�{+�� ��D���>n�1��;뼓G�C�O���"o���-4����Z��6�^7E�D�=L@{̙`3�s������SH��ID����K��sҽ-�B�t��i� z���j �7�R;�C�߁Sf�Zb!�4�?�N��w,����_�m�/�X�0�g�s}g�#v�On�2�Q��K߰u�:�� ,޾L��	r��`�58x�wȅń'�	/�u�Rл�
7�p��.�X?��=�ο�Y��߃�L�����ò��W
h=�jx������U�)�]���������2z�p�8u�u�	@ <�@V�?м ��o���wG�zR��н����r�]tq������M�ĉ�P���T�H,�X?9hi|/gK���_K"wX�BX����&�QfO�Tm�H'��e�����	x��2��Ht�;e)�:�҉�'��ۑ����.9B	\Y��Լ���a�pq���g��EՀ9�,��Ɵbݹ�"�[��8����_[u�1�5�?k��JT���*�(�T��H5~e���Z�t�3���!� �,�Wɪ<x�<���̭��4�vy�����AZ\D2z�L��&Ǳ#�"��@\��>��پ+���M�In��9�!��zKM�o+2�gj$u�^�c�u���j�s�+E$Ϥ0��'?�t҂�w�
�hC�������G�\(_@t��/	ݗ*lT�D�R�vG��������/�w<��UB�c.,y�,z�pR>X�m��kݩ݁k+$?@�:���0��u���յ+�N?'�39�G��N4z��j�	^D('�b�@�1��C��<�U�i=��7���|U�;�$1�����}�$j��d�g�A�����#j��P��?�����R��o�6��]OM%�6��h\T2	�.*H����	3�ϟ
��K��X��>w}�Og�d�4'��k����J	�E�˕?��o�V�]4_�)\�u�.�A~��o��$�?���E�S�$	���^��Ɠy���'�賾�F����;�""�����T��:�[�|�0��̹��I��p㲁��.����<�z�vV��!o�%6��"ho�����I�%� rka�8+��Ff,㍖7ξ�%O\K5���rƦ^�e���P$k�D�!42� T��2�`$ym���H����oA80���Q��g�?]��x����"`}M6 �#m��r(#�kO��'@n��5�ށ�&v����,��D�Rx�d-���t��Ju��(g���5�ʠM�d���瘧�&λQQ���tT�nב����+���1��rS�J ��eH*����o�مc��P�{����k������v�G��~@���ʰ ���k'@ťԍ���.��O��$OJ�XF��P�g����6Y�묭bnH�@��=&�i3y/��z�c�S�|s��0�v1�TY�ዣõ~D�/�iVl{�����CÆ���n\̎/&�mM��Ők�h2o	��K�J�
x�)	CVq�Ѱ�B�k�����Orݤ��)�׹���L���/ �Z�n:i~=�����I�X���Ң6ܙ��$\;'֤��'3�\�K�r���̸ճ��O=�r~�~�p��i��|�PaEŏA(��_��m���R�ߞ6ˋ�_���/��`Y���'�)OZ{zӴEݴ���������d%O����#���M�L �:�S��:��"���A�щp�,���!V�;�@'���o���si�q� U�b��K��O\�l�\vַ�tm�F8.	�'Ճ�ڙ�5��f��)�2��슝�oвސ�\V_��'3�m&;�&�9[(XF�T���vE�v�n�g���\�@��R8ie�G
{P��֡�<�r��Y�@��u8�uG>D�~���
9��.�c[����2�*���@��ޮ��{pU�O�y�*��� cC�u�O	�\�`���N9��ֻI�,��K�������Jz9�7�iU�P�$�ތ���	���i
�r����c�;p0�b�L����:3�5/���=����� �7�����b�đ�F3��!�?����b�sO7���f�۰	��O5�œi�)�"�A?�=T
�.S���s1�t^��^ޑY�5;m�[~	C�p�^�n�<RW�_��Qy�0�ÙV���ʇ���w�]�*�� �p�d�e�ۦ�;�*H�q�бY!��"��_g$A�#R3���I�j�+�@l�yD�����[
3\o_)7�t���r}�܋�B��{us���A�I��+���L�9��}Ƿ^�+�� ����xg�� <�B����>*�� �1*'���`���Q�~�L�+'�i� V{���6&��$�>n�f��hb�H4^kv��������_@ۀZ��l�zS���7Q�o����9��������=�z�}U��-KPM���拨C2K�%FT�	�.�aP����y2=f�)���[m܏�'���u�}c�`S�ᑡ)��;r1HÝ��RI��1fI-08Q.�2"���K#Ǵa����~h�@Ҫ^ߪf���8H�CqM裡$���}�/�������y��9Ir��H�=��^i8���ݔ8K�u���'��T�DuC�S�zw�5����y�}>� LbP�Q���/X�VcX�&p����A���|v��-9����'�持"؂�T�����O�=�pĐ����@S�'�,Uc�+!��-��#�>k9���0">�G(���֮�&n}�BT8�ص���+r���ov��!6:�vhM-ׂjN��:���E��	-���%���;\�˥��Ҿ�M�
�Q��]x�R�&���	H�6m:el�)�*Jy��[�pC�&t� ��H�X��(�81��(e�u9KYu��6*|gi)���mp�T�I�DN��mt�������x�~@��]�b��$������M�:P>���(�X�J9�U&ԚFE��NŽH7��,��B8<f�>a�wz�η�MyO}���H�[��������;�6G�v.NO�K
��B�S�cm�[��mIv�#ou|,��8����Ĉ���=� �>�^TS���#M_Ǣ��}�E��	9�!8���-ط�B�-9\ޞ��R�K�H]Ӝ��4�ڙ�^T�ɽ;��M�Pfk7��������H��B�<G�d��O�t�ɏɯa��qr��^�]�c��U�����6jS���E�j�Ed����[�,�V���r@NNu���W~t�7��:�Mf:`�Q�HꝂ���[�.��̹�Ѧ_�"��ˬ�m�ଷy�'$
���Qԫ�9���������5� K:R'čO��R��Q�N,1�DT��[qy'ʿ��G���O�ѹ�9^���Qqbbas�.H�S$_���d�i�|�f�@ŤŨ8wqg��׺]���L��/�e�;K��p���8�B������,G�ܤ�eC�������������P�gy~��-��	�C�Bl�*ׁx�/�rg���Q�.8Y��1��)��8o��e�'}�����j*rR�6��K�N�߀���W�g��b��P�Rئ�v���}^��3��a�\/$�Y.��qih-ґ�c)&�ƻ�?�7�[��k�̬7�j6y��Y�=��j����,�&4,��o⊟�kq9d�E=&q�pI��g�,ڴnH���y.�'�d�syS+�\��U�h�qm�r�g���>��8�i��A�����*���^7�G���^ ���E�ER��W��"s|�q?��K����֓	��o�k�����dd9%�2����\��Y0�5G���>>�]0��Wf� �e�Օ�f����U7`�z�*��)�;�|V���13�^"I����wR���D�]����6^�Q��`��~Yگ��Ar8]/[j�G|NGқ�H���ƵX���a��cV��x:���R�+�*� E���D�|��Sh�E��g�RLuܽ8���ьS>�����js��`�I�<>M�8����.j�B��m7�ӟ7Ԏ�]�ƞSݦ[E#�2��i����j=B���6��k�~XI���r�nA�y�Q�R���L<�;����2h�2L?'��n�dP0��}����v�x�e(M�	'���qP�)G��l�����0��8-3��f������
�K��F��O2xp=����+ߊB�rӿ#t{�Mrd�!d*P�����8_*�k�
���mlR�	�d���ޮ�g��)�w�������u����6��%*>U`l���U}��ܺ%��פ^��Y�%�c�"��+�(#�����X\����sne��)���F�;HCsX�<�rb̴*yW�]��"��F#ӁV����l�6�df��u[�	���=��ֹ�����bt�O׫r�V�r�|!7�'��\�<)$�o���ۉ���?���������hm�	~�~�Ǡ�i��3�?6v�6�vU,o�c����XVvȖ��K��NK����&�}�Ȟ��J��R��a�����g��_z�ޏڤ#s�4g|UԞ���R8p�ea�uTԨ6B�x	��QE.m���{�Gnb�W��6`���`�[��JI�	+E�2[*���|	�?�~K2_���:d�;s'�m4,9���J�/;䃋 �>p��4h�M�"�9���y��eJt]去�����H�i��S�e0�&A�,.��!AE�~l{Y���X��E�>�u=0@r�D��-�>�FL���J�Q�,��`;�#��o�b���0p�5��������Ԕ��ɶ ��oٮ�ڊ���>KˏO_�[�)4��N����^{r��Q��!��M��(l��[��$6� �D���k_ܴ���<]Lꟑ0���Y.�gI3���$2}o��n#`qK ��+q�8��/DC�OӍ�=�]F6���n�s��Q�ʪ1 �gh}��{/����0��1�E��o����3g��_��"2�����[�U�����J��P!a�<6�7�]T�tNA�"3�);l��]��]��N'�O��/�J۹Y��N[��<9���%�M9l~s���C��Hl��q6�^�z���qJ��a�Ioݗ�s��Ѹ�.Q�ª���p��G.j��CqQ aa��n���V�7�.)����4%ԀW;	��3~3U�5�j�J�Mgy���ϋ(9��2�E��6;� �nҭ���l��$�pN�㡂c0���Tl�:���/���{���� �3��C�X9�G��s�k�?��s���J朒S�������-(0���@�]� ��ڟd���%c+��
��G���)8l&v/0I9�d��!�E|�|�t�
��L��Y �xy]����榀"�@i���{&K:�f�q"ŝN9GLv����w��?��#QӚ�a�V�e�a���:s�n��={f��RG���RNWvEwħ@&���ig��֖Pu�\������K���c�OuN���ͦuSnf�:[_Y*��JJ��Ђ�y���0|�\aN-4��u�����I0��NEo�����r�f�I�!�9K.�g'��m�u�ߢB�%2v��bf�x�D�)�>���3����|��O�FT��z��iA��Y���uL��B4�O�1���&���T6�&՛L�4a"'�z�!������X��׀5j�^<([Ur�?��Ҭs��.:V� �(�a�5���,�[�]XSd�;xO���%욚;Q�n����S�3�ǫ��XX���MK��氺1����	~k?�P�΃������G�����S����к����x��FN;��icwe�U�Ό�l<�d~��"z�&�଍��#������t:���x�V�*q�)f���۰�jZ���D���q�-�d��C&H�M��q�(j3�7�R��ʒ�5DpWy=N�ճ������Q����Y���+��mA�(�/��59�yCz����8{����M
����9p
$��x�9�/*Ȅ�v��K�ElM7������f�=�P�c�&�M������F�����UZ/f"�A�ž�����r�[���gt�NJH0��#��&u4�^��໰�����\����`��Ŝ!�/"��ՌU��o��+k���Iy�;e)�nM$�9%�(|��av�]�Im�!�� ��a��88 ~�c[��V����_�}�QT;�i��� Og����2�crЗ�i�X�j�_C��rq4�ۀ�`� 3�/�[��}zVܳEm�G�5,�s�k$~��C�Ϸ�Fcj�LԈy�C{���Ti1�9�wZ�
��C+�
�2G� �#oC�=b�t	��ݼU���j*�.�8�	R�hϩ�t���^4?b�P"��1V��E�[=��`iZ��<�'�3H�%�+�Y�f
�#5m��\w��(�5=��^=�j87u��FIr�G�MH�x�$B5f	8y�׉���@�v���Ƭ#�1�><����q#��{U���6!���z����l�D����5;�)���䫪�ڛ����.	���Vk	�.J{��!�0�`��K:��12��%�s
���Ŝc2��O��)s�,�A3�Ψ�p��R�@��vn�IojO�����dM&ڙoD����$(|��K`o�#�m s����8�?͔������F�G9K\X'�?��{J6;�Ot�6�xw�V�(Ylj�!�������ɺ��m��fA	TG<�E*�2�%j1�p�#<G`� ��뼌;d�F�#RՎ�L�� ���R�pV�ub2r��gM8��z�mr�5c7L$�V9e}E���P�0��8.���E�$q�ךb�%��;�A�/��!�)L��uz_�n�_��̤�ʺ}���G�i��|�R���4.�K�'��L�Ȝ!k�U�}���~_%��E�s���Ϡ��aܭ�1�$�W��9?S V��N� Ȋ��{��B�!����B6[w?���]Qp~���=��Q��i�����ŏ��^ o��>[����87YO�c�G'�
�2��T)���f�t���ep�B��z �ޥ'm�9��d`Jë�la��j����:i!H�8*^c��-�ˊzl��V�Q$I��'�W�"�Aj���T�X�a����#����T`H`Ei�6监}�D. �������(��I�
��?��LF8��� �U"R��^C&����K�q�#����A���7��*��&-�K��A}��
��?��X;���f��_wbX��k4����q��@ʖ�����,G���n�|��������Ҡ�q��k",H��Gћ��+A��x2V.�!��_���Wϖ��}Z�U�p�y[yE!�G�0S_.�����r��wC�I��_��d��U���
�V.zỰI%�3,_�m��튗�{���Q�����\@������h-�e��,�~���T��%l5���7�nM�Ϩ���y!J!(��D�[��QG�&���&���9
m,ه�&���ܿ-}�_��M�2��W`�q-tU ����*8���H@79 t4㡂���2(�v��E�{�_����R�Inza������3g	�6����K��/r4�cVT������C�=p�Jw'M��i�F�w[�IW,�+��|�,��2��"��b����w$���φ�����g�D�+�Q�>������OA:ro��d���^����ŉ6-�K�SQ��|�7��l�"��Y�w+xd��0~T{�z�a\0q�,���Cْ�f�9q	�-���
JH��8n�""1*�yj�x��ϗm|:�J��O�k*�0�m�Y������K�MY�_��l���+/��f�Du�s�N#���?1N��ڭ2�ٗh S�M�7nK�H�\	e�	�c�s��%d���|�щĶ�t�w�`o�0
Y�K��M�ȣҥa���8V��M��
EԹX��9�JHrTYG�����ҙ������;��k��Wg�H����N-��p����� �x�aZ$���!!+l:���wY.O�BgP�I�<��U��]�<,i*Z�����S��w�z�����r�8"�JP<��I�K�Þw����ز��Q4�[�g�^��N��(m�w���eY0��O�vL3`<�qb!1��.<��9G!��:ӡD�������$��T2�6�`��K�I'���W�~���H�ͨ�^H��·�^��2���O'P�q�:��{�g
��n?��,��"�W�F/�����C�|D>阾qH���%�w��w��{�A�~ɿ�6��TU�ŉ�`����p:�)#c�R�o��:��wS(kE�Y�JT�,��������8����	�8||�M��;P)�x��wQT	��2mQ�H��t5a
�>2"˼���A�3|��]l��"�C.�i-���00rS��OfC/��O;�/B�aڜ�?}m�Vӌi߆���m�󃣨)�SAA��)}�:Q�V�6�^U�1Iʉ}[���i���*'g]�f%q�LdV�!c��H�G��4A�[�łP��U�@9l2)�K��T��+�]ӓ�@!��9��,�ܫ]\tB��&j���!��*ȵ�_q��u `x���N�[d�7��d���'S	H�����aK����]Y�u�8���p}�K���߈_$�2�9ÿb;K��,���>�� Al�C����J͞�ͺPĔ`��E�؍��6:��R�(��%w�dpDL��5���e����=��E��p4w7V��פD�fs��C���|���v�͞w���Qg�4:�b��i�&�V<��Ppl4x(�hT�)��bj����@�&�'`�!um	
��vI�ih���VwF�.9~�n�){@��M#��f��(�vE3�����M�%��Y[�V\��p�%��[G�6����~g({$�"kƇ�������D������J��l����] ln)X���Dj��t%{LKm��۸#���ϭe�������T9r�i�;Y��4b{i9��%��^��]�l��72'K��^�i���jE��{I��@�k1�d�>AeMlQd]�981��4]pߧل�,4�V+ ������aLD���Oֵ\����^.�{�o�N!N!�r�۟�0b���rΊ��L������"Ap�>SS-��q*�֊���Tų6��fH��L7�.��+A�E�[��[8���OOH;���PPr-틸��JV$�;��@t���Ɏ̈Ts)�Vi@(c��s�e���(����?�Z,#J������)�C%��ApO�����p_	�U�ˠ@1Fsޖ�A~!GO7Z��?e���� �Q��Kg��m��w#�"�9M9REKg.�ꉹ�"�z�/Ș�Wܚ�v�|�2ͮ�I�懡IFE�+e��%���K���
�Ҁ�����E�;��)5����["�:�w�l�����?��n[e`;-/.��e��f�/�1���n�N%���Q�\�p�wZ���
[<9�!�\���L� �	��?��v�_)Qg_3�9X��#��)�$�,���&^����ʂ^�X�����`/��j3]�����:ĉ�|�N"vX�RP���92g֨
��!U=�X����[/-��i���]�a�7��ˎ���z^G���GX#x/�Q�fn|S��|��ٿ�=�����m��$S��F§��z���+�jU/j�5�ћά�57��Yi#&�=h�a�D�iQ���80G�^�=�;�a�������<�ZJ�l���aǿ�����f���d{V;��+��?�7���wpw�p0f���u_��D�~�ɰQ�m$'C����N��䗌�T�N��?��ؙ�N@`�JB�*�<Ӵs��.�WOf�uEs'PS�O����tg2�wQ۽P��t/nlWU9m���:|4K�x��Di������N�ja��%e	E�U��qY@x[��2�n8���[D�6�d��dr�!�>f5QE�$J\�����T_�W��S?�l�?�QOh�z���G�K�r��Ѥ)}����?$�4.d����s�~Jl������Mh� �WR�Q�S�6�Âh��-���7�@щ����2��ziܬ��*�hCGڿP�q�5��yg���}�2�'�16�N,m ���g��ʨ�b�R4B��X��#Dd)�,��z̅L��_����G��ܹ?�&/��S$x}'���2�f�]��w}�΀���ۑP~�޴�UJi���Y�D-���oZ�="<�^0[+������""�1��}HF�񪿱B��R�7�-N��:� �Hbq֦����◟��33��y���f�	t�#�=5T#*#B�jDbS��֭��߶E�è_�SR�����v��nڪ�$�{��¡��o/bIP�xД���]��L�WRn2�rJ��>�L��i�����ۺ���/R푿G
Xa��%�� ���+�b��
S�w�x`7��F�`�~�jyG��WU��!D$�n��=�Z�]kk<�_1�VlV����ͭG��j��p�b���
�'����� ���F���"�62�Sl�{L��z���\m�o+E��\��:�b-��?e���MK5�h����aO�Eͫi�~���ߊ/�fC����i.	P
�����X���e�x�`"�巄:��k����KR��*�%�E���\[�q�D-y�����o~�i�7
��Dh/����x�q2D}���L�(��U�)\��0�9�7-�Bx��dvfn7:^�Ӳ@�vK˕�13��qh5����O[�]�!x#�L'��w���X�����'�O��Q��2Ό����f,��d���ޅ�x�n4��HEmkݶ	NX���J�j�E��@0e8.�cq�Q��()����+9%LN���?SM�b�<��ow�Іw�y�e���J=���a+�
JOk��k��\r��xo,�lq�>4(1�%�1���������J~�BB`F�|������=*V�W����_.a4�l��~_[�-X�*�XG���e���p���v�Pp��=�a�e
Ҥn߳9.�
z��2���-�g�?�����f�
#��bR�2�yu�����Q��	�d�1p��t`#���Gb���w��PE�4W����t%�:u����;o	+:>����!�-��gP�nVͦ�L��,�z��M?E���2!�"�;������bvT6�i��ݻ�p�3��a#l�[�<D�U�z�[��.���m�ͦPz�	�~e1.D���ͷ�z�$#m��mUR�W�[|F����>0�4�`#1�T��:���U�=V�ڴĦx܄:���.��ϳT}����X�kOǜ&�@׮0����֌��=���z�M?Ge��g
Vc0��5��x�)���5�usæc��l�d������D��謵�z��1��Xs@Y_�jh�`&^�IidiOb�d�n, 't�L�^^����h��ϓ�P|RP��7��'��=i&�-��k����y�E�]}�V��>��Ώbt��K��������G�qe�,yd�$�G�q����orQspr�S"4#�ho�]��Lu�✜C,|��{2���D"�E�o�������+4��+��,�}j/
�����o���~�%X�u �◛A
ʉ�|þ㜇M��h5�5�������N��@�Ó��L_��+h�cG�ը!�����J/��
��~��N*�J3}��h+F.ܫ\�����V���v�;���憐?C��/4�1'D��RuD7�a��z		�p���a?ۗ�a_ 
��j���q1��nE�;%�	a��P�qX9�_��-xP��}�N��{\$���8>w�N�o?v��~E�L���n���ƌCq�/��*k82r"�	�q�ͮ��S*C8���w�!�����"�����ko�P�����gP�j8d�9����5Ir�L"AF�b����=#t�2W�290K��0Ҫ��>��02�u^��ҋ�9��F���3GN���
�0����s���W�����0F�JٲT�=v@o�<q��&�O������$���I�fZ�`��z�eW�C�<����3Q��|�E]����;�����b�G`D�4����)�R~�:�������r�ϥ�Ƕ֮%E���W5�2� |Y��
mТ�*�&ʻe�(�Vr���G9�#�/���?m�Ԅ�$�E�����e����ި=nds2�i�<�}�QІ��|y?a�#�������9bBD����6-:�Q�l�J�ڣ����!��>��p6��R��	�l���bKN(r��"��pv���N�ɠ�ciM�o^/������L05Fd�:\C7�(�g�^L���\���EJx������+�v���.��,7'
F�mϱg�1��EtQ�C֠~`.zf`��2#�a%U�r�ӈG������}�����0z���X�QG@���#�L=s�}�H.���.w��8	�q<Y�e����sP	��"aZ�!���:~�D��ٽ/�Z]�1��`1��#X�g%��e ����τóL "�k��GV��n�hvc�l�X2��m�@�n��x����<�\!t���YZ��������J��'3����y��q��#�3�b/p��鿺����nFN1���m5M]�pY�v>ao�J�h�ߟ�S�y5b�(�:ǜؽr���z���/����fV:���4�v�_��%x�TN��a'T�9B�T���ȇ�X��M8�{G�V�{�&;p����>�w��5��ܷ�2�M9�3��C&�0��������j퐞��x=�q��q�\�&VF�~Ƣđ� �p`�H!�Y��3f��z��Ú%m����	%��=g����S5�I��[@͟_w�T��h����B(c���f&�8O�'?��K{���y_��1�
i��/���'� ���m�Ej7q���>+��A %����yOk�k(�-�T-8e�;���?.�]��8������z�L��|���?��߼+�ڌNs�BzIӭE��8��P�x�Hc�Iǔ:`��� 	�Z��`R���Z�K��q	G|ſ��Zf���ǁZ�"��F�.6)T�{ɒ庍��5m$J��T#���K-蓌���d~&P6�@Ɏ�q������a�&��D,�;��v�T����YY�֛qƂ�*����3*�~N^g��
���V��,-�ߏQg�$v2���
 w]ݎ�-��� ��"��4 k��Цܨ�`ٜ{7��I����UR�s]�1N��mt�^���7�'��;�SK����n�A�=�A^5c���K�:5\��Q�о k�`�l��x�z�ŋ��"j�׷�ˏ��U�q���#�?��H��m��¥Lf���T8���1F��V,�)���ERQY�(������6���+y ����^E[�'Y���9T㦵zHB @��X*�i��M$U� n������Uϛ�18�����g�͛��%�s�f-�(�\��䏁�P��e�s��3���?�.�bC�������t1B|�o ���ʈWnQBݏ��a<����Tx���4��=ą� ���d��~Պ㐧>l�ŝ��AB�2�c���活�V��O��|�|�� �������hָ]H��+Y������&w����W콸UG���=6n�2�Ա..EU�<�`�%dc��o�[MbF~sO@D)˜�vE��K�X�R�U�����y`T�N�t���3+�G�W]sB͔����P�SŎç^|����T��b�˰\O���	9�\\������?l=�
1�I�c��r�Х��Ƿ�vy�lBbRY4X�N��z��tW�"u���h|<�(fy���i�/�#��dW�1Eqd��G٥�jE�W�~0ae�3+E*�[�ݰ�l���c1v|�H��
�n��V�r1���H�oj�S��B�%z<��M�C}�87�E�x�i��Ⱥ�z���86jx�Ǹ�.J>�	�X4�wY*��x�l����n����Qě����c�.Q"Iv5C]�� .�����~.y��j�⧇+G�D��d���(&:O�̡&�oF1��|�4��w��q�w��~97����>��@{�Rbbe+$5�\��D1u?l��UT�6�Z�x�͆��N:ps�}���i�Ւ��_��Q�_�=�X���:�4���B�$��v���?G<ʽ��]$���!H���ٗ��> �3�a�][�l#�EՀh�O���(�	^O���td�o@���V�G0�cV���{>�=DGe*��gq3����9�}�I<^��rZ{#�߹u)���-B��g��C�۷����a���1w����7Jkz*�׸���,v�� 6��㏎ڎT4��ҽ:$���ҬΠ�,3Qe>�?���Mު��h�<���.�8P�PdC�p_S�(��ɗM���^g厜�,k4�҄R��E-q��*��;w��p�S�_	�C�1��0s�Vz�3����VP/�v��gqq�����Yz�ֻ����)�~��E��eD�k8*��? T��gLֱ�{��*申�s���0ط�� ez������S�d/��x]�1IGnTT>��p
1U܀���	a@Rh�ϑ����K��!�h�tG�[���:Tl��DdVSkW�]WS����A�A��V��E<����7���Ĉ-wG�mPݡ��<����5���~�}��[0l���	&�P�dQϿ[��-!Q�
�˝�f9�V!�$Z_��hm��������/fIՉ�T��н����0%��M�C^��A�'�};�oH�������Ǜ 4v*�!�H{&A�%����q��W�4��\�b�q��X�s|��$�Ӵ��P��{��؂��}����%1���`����5�R#*f"�����ݷd=J�M@��I��_�S>���&5�Gx��,�0��K��Q֌*�v۶����Ʀ�.�+Fa�?��#T����|�g%D6���r��6�_̇Z^x#�r庄���E�[���9ԇ�O��欍C�UZi�.T�g�����P�U;����>�+r K��{��֧� ���4���Μ��k�#��_/�A�JUqC*G.γ�����6�E�!�� ��������a����7
��b��ma�q�I���a���i�gޖ����dp �_*�L3:���y�7@6�9{�L	�L��Q#��k�bqχa �~M"��b�u�BD�A<=��}�1�4��� e��#8���SdZ�=0��Q:$z�/+�<�S�iz�5�^d ̭��m�	�V�W�Oj|EȎ²Z��AS�"��O{#�g˓������vL��;��Z��>s�Q/]�Κ����~(�⾉�@5�em��+���i���׳���PV��>��Gj�ۜ�}Y��kGi3�M#�3����.�����S�.(B@��b\^LAy�4��nz��폵7ē#�!�X�`���"�w�����ك��N&*:�8�s8��J��G�����|��#��e�U1��`�̔=k�(�$赗��qJ���{ A�\��Tl��rW�HΥ���a�L��t�ը�K�s�&�ik����zU@"���c�����w��zr"���m�K&]�@�2W��v���࢔
)����Ru�#1O�j�*v�����(����k>>L�Y�P֩�(�C���3�SC�:ً��qb�@����Qe� ���VP��w�æ	 ��5�H����L���(�jHB�r�3��p����֧���aMw�|�V��t�@D�vF�p�Q�q]��E�g�����?Pp�v��&Nt�CK� /k�Y?
�sM��0�@�N�	�'Y��,�8^���`P��#��v����d�o��(b��U7����|�J-Bk1=�Fy)z���*�%^("�R����RWe�k>��A8�)ަ�j�R���L5�T�0Jd�H��^��[��e����DʍZ{�9x�Z)���t�w�@�:�`Vۓ@ԈN����j��>�.r���
 J�=E���i.�:�Kj���HL���{��:�(���1}6&�����w���w{6VQ)�&��'��|Ƿ��a���|4ȦJ06�i��8?���Ff�^�0����>3�K�_~�}�E�}��IΒ|1gYΞ�ρ�ehգ�/�E�%"��Z}�Bމ3Vyh��|Ď[`�G`�3�����$���q��3ʩ�*�b�z����'�*6�7B��0��9R����UZ��^�#�l��hq<M��V��U��3��<"�
Sβ���؛`�:Ds{U1�y;��#/;�2<���9�8\+>������a!�C��33�$Ғq�5
Y�0e��$־eLF���y;��+����
��^���������'JQ��R2ʇ1E�K��ㅻ��e�o�t��{�L�^Yh�]�C����|��i�~Hn�ƺ��[�9��F��YVm1���Dp�1M���Ù���r�b�9��>Ʀ���s�|�k	�����L��m�'&�3�rb�cؘXظ�DN����}3�a�b�[h��������f�u#xD"qJ�I(/@�I�P�l���%���'��c��ͻ�vk���rW��!��ɏ���Ѕ�~!|�`�G^)�ߣ�^�������hR̩_��|�H�	{�����H
��)�fy�cTzp� �s:�Z��VNZ'��$�f�t=�N��P`h{��@󊝐��|N�.s�VdTR��FWt�Tu1ڕ�1de��y$k,-?�	ݲ��=]�Pv�w�Ĭ�R��bI6j��]h�x$��Q�RFi��ۍaNӪ���.�B��?��_0O�s\�!f�& E�SlWC���&�>�J|��-��n���s�'j�,��Pb��W��|�\���<h��=�^�,՜v?0ʔ$gST��o&n
_�l��f���f!ڣ�Fn�'��~#8���8�R��3���p�TXV�h��+��,�ͩֱ˅��5�\{t��%����[T�{��������_K����� Ug?ogK���ƨ
�=�(�'�|��N��J���7Ԍ~I���#v�10A��n�kH��=g��^_��'�ر�8Ws�n���������O-x��l��ynsf!�J{*�>�F"����!֚�����3~K[> ��Q;p�d���~*�2�%^՘�3�4�����ZKO���{��7�v�����\�7�|\�zX��.$�1��l�c/S������W��_R<lX�/-*j�a.�Dr�ѫI�~���~"�]_U�ɯr�<������/%2��ȕַi�(�uu���3����=/�(>�?�j�W�e��� +1��"����$Z��	����3�R����R�9X�� ���4pd8�0el@�᧗�L҂�Kma�A��n�g���b�8�������3|�
*R��K&7B�Ff��Î�:�$�s�o;�������d|�x�&׏n�8�����!UΪq�^	ݘ���}�6]��s�H,EY1�U�m��_ܶm���y��S�d���_aD���
�'��{V_Z���*��#Ց���Z_�M��-�rZju�24�x��V��D��+ф�1rT�*2RhAe�v��6?�>�����V����SF�����^�|���1^d-��M|TE��u؊��Ԉ\s�_Rt�2`����^`w��
�K�ភc�|�u	�����=i�q���+��$3�M�<����l4��;����5�q�B�Έ,���U�-QxZ(v(��m�߀�aw^>'�K��
Ta�$�έue��7(=M��<���j��'��X�޾�m	,�E�	�����@12�dE躔*�VU�O\auԄ���uZNCt/�Vm�&�g8!NGI zwˑJ'���I�;S���m��|l)�j.<K%Оvy�n�)��������/�0����B��9@�7^O������'��2�ʰز��ww�r���.]����D���M����\+#��Ŧ��P�a�\�:�[��0O4�����U�4W�'eyH�M�.x�W��<�Gv;��Z'��l<���ƿGY�;�b����"�������x4L��-�t��tR|%�#�b���+>7�Ϻ3�= �v /"Jt$: sU�J���Y#�
�f���h'�B��#�8�N�'׮��~��ɣ�%뚵�P C���؍n7��v�_�=LIG�5x�I�)�}G� 
L��g���	�6T�}�Z�,Vω��ZhQ�ךF������h_�c��A�Et�k�|��]�6 ��Z����X�����ȏ�F=����b��-�׿G�͖L��	���I3mfeK
ة�˅"vVO#3l��p�ob_}��WE�i��{fN��)+��ҡ���%�}�"�����K�#�;2�U��%����IMK��k��������|�ݒ~ͳH�Y�g���w�X�J�B�wL�ב0*F᠒"��b���j�튆#`Q���F�O߷ͨEc�
\�Me���B���������^]Gk������#�-ۡЎ|��+]�b�d��{��	�Op)�����W7i�[����^<����m�<��ڕ����ZEѡ��薕�{�Y|4�LkM����Z&R��ݝ����ƣZ�_h�)���U�6����JU7&�%:)�2�m�~t�r�/v_�l{kZ�B��%͚�`�(1{�~'pg�{�܅=C�_���8���.(e�u.�|q��ni�X��y0�3���i����q�ɕ�Ȕ��`�l֜ƿ<Cüg��������<�{b�	�E�ǉ���ʧ�9�FB9ӿ�!ɤ����,[M�L�
�Ag%���>��i�oZ�[�V�ik�`E7�4k*���,P�b.K]]m��`̺����c~�j��h#D���	tэN���K��6��<�V��/}K���&w}���^�VS^�ZOBX�r;���"�����l� ��:s��YȨ�lAHKd�wOc.X�2���p8��Ir�2Ӿ���`��5���5�&���9��|���<���=�!,�is ˺[�h�|x6�B�C�ZWV�c���W����^���J�I�G%�Y��E�,R�_�!2.�_������_�;�d �,GIX��Uՠ�#���wl�-�{�����x�e%YX2%�V�Uw�����R�n�$��om#2Q}+G����ڧ�Awm2��5�Y)��Őn��Ŝ����j�b���0�S�o͖��.�X�~.h6�5�	����:��c�-���X��I_��B�y�O��͌A2��t������j����8�B�wuBF��x�������Mܕ���h7b�5x)~��պY.�'�EP,s��?���f*=������#w�Q�b���F0j��S�[��T�V�]�Tg����,
S������;Ø�c�F���cF�	�Q��J�����x��2��|�Z2�O� ��r_-\�s�k���}X������������B�_	�6�k��!�a��I��.�X������k=g�ՎQ��#���?��g�.�O��~��v�
?`:���4B�K��-O�D��<
5E�iMH��h� ���ơ�J�t��Y����b1����,��U�xo�rc�}��H�yNO��Ƞ�g'�~��vLj�G��$��$�C��w/�$o��x��\��1�����J�JE�1�H�S0\0�f=uӋ�s�7��g@��H�͚eڐF�.�g_iM!ɪ������,Ypr�+���:pH+D�Oڊ����m&/�e�
`&]%G��Op.��d�-�6/�Ŕ
�n�2}Qv��ˤ�&��_�!+��Q�P1��|��J��9���jO���KI��z�LX�/§#���1Z��5р�s�@��v�B\c�h�C��F��3ȃ�JH�>�����R_����K�Tn�D[�duWЦn�ey��K�%5I7qw���(�#.b�q��רQd�0��Te���pt ���߃�l��S�2 #o�����<VWd�a|z�z�]5�o����og��I2���檀tõ������R䡼s���wf\,�XI,h��b%�u^�t�K���ҁ�uE���%ȑ@��d��O�B�P��"k�P+_l菋�w}bD&�m��)�fkK�5� f�}�:W,1���F5i�N����M��iٳ��<$~ wG��$*�cv��g"W���q�2O�a,���u.�'�@�4Jՙp����nbW^d6�ǈxk��Ah=
�|̣d�X���ٟ!Ā�ކmj����؊��b)��u٣ErD���W-���^��CL��@\�N0���X�<b���T�	C�[7]���q'�s��*������G�)k�ۤ���O*�cձ�\�d�j���սG%���ܭD}�67h��w[l�@��#O�t6{]"��,��Q�2~�NH+�x�N�e�:~��	�r��,%�蒡\�cn�ƹ��{~���/Mi#S�5v�G�#�x*l�r�B���a#��n�ؙ�r�7�cϹ�ҁZ��Q;q����)�`� 0�<���g-|���"�G�Ӵ�9��K_����;A����ٓRI=#R�.ӡg� ��C`_�w�'�(����	�z��D�.0���v�R�x�X�W�(AgU�5����(���d�=��s����O�\�a��hr}/��w T:8����ec�����.�YB� r&�G��J `�����0�g��A�˛���^R����j>����6˭	%�B�pY�Ni��O�E��ۖ���XwZ�c}�`��~�A��0E�a��D=�	lņ����V#pxU�L\����ȫkQk��>�y��<�¡o1'X��)�"�˗g"m!xL�r��RnPaݠ.�d�ޛ��62�g�9�5���cs�����{g�0��q���B�B�o����=�����c�w��b@&�w}V�ܸ�t��k!�ȔR2p�|v����
�����Rj��>9��Z�<|,O���<6����rhb?"xYq�~ǒ/�q<�b����虌uq7k�Mlv��@Ӌ���=`�3���|0d�׈��Ve�μ�"IX)�tT����#��m1�#KS@:ɭ�-����L=f��}� ��̥���Ts\t�ޞ�ܡ�1j�R~�r>��u���~�क़�y����O��R���!�(�T푿[D��`�G�٢�$'�MHTy�L��y���:�	��X�N�R�=�Z��>>�>]�=Ot#u�{_�#B6@�Z�-�k8m����DE�t�^��$��G��J<�I`���(Uh��Y�1�i��Q�ދ�=o�.��gaXc�$����9d�o�,�8�Yn�Г�p�C����g���Y'���e�# ���&�W�Wd�X_�����7���@5R8&3P�']M�FD����� ��N;W�h�����*)�0jP@���z��]�7K+�)}q���tC��m����=�T"��X<UE�N��Nɣ� ��-�;����(#���A��A���r r��W���Ouu�t���	�>�_v�)6����e�D,j�|`{@�Ҿ1�y�%���2�̰,B[^s\q6rj�w�d��Ǟq��ڮ�]�?�f��-�]�t�F��˄�c�������h[
���������%;�����	oD�sʚ4�"���O!/���D%]��8�}J�����g}}.���Aq��(�p����aF���W^��!�p��E-���'�`\�^o}*�o^�{%[���P�Q� \�1���Ԧ�[�[�4C�z��jR��<��DhЇ"������
kvݞb.9L���b�jWU��hG��-M�P�0�t�K�h
���5(ZnJ���s�4^S������*��Sj�uc|G���_=��^�)�ղ���ś���O̹OѦ���H}]���h�U��g,�pR���؃�/�J�4�����M-����`�Sr�:7�U��U��� �/zlRI6�B�#��Z�B�䴚���g���hx�d�Z�<u���v��í�,���l]�ݘ�wT��T��	@XdMA�=^����&:0=�LP�>x9����֭�[��=v͜GqϾ�a|���+�Cf꘡�K�R���}i�d�ۻ��i_\�Mi�_j\������F���ZVl�Ƃ���MS�A����K�S���O�R����G�n����g�<t��2��]�q�9 Yݜ*T���y�c��R�b�_mq�1C�>��yc��r��VWU�)8q��3�O̫\�Q}���h�8�k�F�h1�qN�X��c%�m黒���p�ť��	Ѻ�o�����k*�Cs�23h�-'�"��\�aR�_i�^j�2H��),�Ġ[qE�ik)��ь�E�u��r���D��oc{��D���AoY���]�&xp.�e��|��=_����\�Y��@S���Mˌ���r�H�Oe6���81p��V�Ѫr�Ɉ�l?bZO���4��}z�P��dً�]I.չ�萘+{#1����wP'k~&�|p�����|�
��o��Gh��H�d/�?�"Y�=�e(�I��Y&��o&���� Bϴ�g���d7���;�Λ� ����JT�G���@��΍���ןFv�r �3j?�`�e���Q�̜�����6!DL�USnR���ֵ[���;�Ǽx�Uo�U<�Iogڿl�-*���v�3���?�ѧ���$P�a�4֨T/u��%��|vT�נ�0\�1_h�ʲ�v;��(a���S6x��aq�k�سN��{H���'4���*52A1�҅A�в9��S�eR����r7��ɞ`.y��e�ii��"C"=eN�'�J�)k��h¼v�zz�A�W�NԦp�!�{���{� ���`�,�콇~�@W)�a��+���=v6�g����<�TLM+�_�ښ#b$ɎUC�D�ҝQ�94�y������VI�]`�μΛ�F� J?^���< ���M`-�GJ��
 ���!��i.T�w&X�s�X�y�sE��F��P(-X���j_'|)��/�#V_^�"G���7�҅`x�p�rx�EN��8wN����ub�a+�X":����s�ժ,#�4Rd�!��R~�$[Fq�xb���l)��a_���1���ѡ�D�2��^K��?4��f�wt�@+�
��q�7�#-R[ytK>O�ii�UV�}G��"8���D���n<��n��f���������;��0�I�n�3ծ��ino"蔚D���?�S,$�c�y����@B��jm$��\���� ��8�G��h�V]�i����(ISc��ç�
	\C�'��Q�|��<Y�z�,-P�1~Ya��
����o;v��n����aӆw~�������l1�ʷָ2�T{��4B���̴�7��|<����?�@�ѫ�J��S�hdK\��E2σN�x;c�Qb񠒧�ҵ�I2>��n�A}3צ�lؒr)�b�a�L3��F����oE���y�Wd����:��=�|�N�Û��.+d��,�_)m29
�jF� ��,�~Jzz�����3��25]5��|������r�rT$X�'W8�+���̼������.~�������i��M��kV,(�z���&�V�]���Qə��|>-����g�H��H�ٜr�^����iqz�����z[��N��۸޾�@�ȑ�+�1uQ]�@��lcM��1Ud�*�?U���0DۼO����\�.`�g.V���%Q������~� -���nBQg�MT�qp�*���
�7�<��-�dB���;�ٴn�3U��������s�4�	�!dV]?����T�׽��!j�Req���ȨE	?�O��Zu{�$^}=�`����6��TO���L��|�,r��2�X)e7n�n'OyοE�r��	��.w`��*\��Ox��e�� �_����J�O��5zG�7P���.�6���ٶR�K &BP�����n��G��"�&[n�#�*�����"���\��� ����{׏����[�9P�ÿ
�ySŁ�a��he�{����X�T�;/�����3"�kx���gv�q�ϲ�~@ �#8�b����3_�U&�l	���d����+���C}i4m�)�Ef���(d@6���-A7*�z!�1ދ~�.C�q�����S�w
��;9wW}��~��T��������zwͲ_3����"Q�}���!~�)dM�˯*��7Bj�����y=���@p����6��Iq}	����ƹ���}0 [���b��TJ�Q�'
�Ə�HM���\Ҥ{�C��sY,���la[�� �����h4���j���Ε���[`��V��uKS��(��A2��l*M ����Xin�:��y�#��3C| ^��cYM�/p�*�xFN�;�����	ym���VW����x�c�˙D h��<��Gx���~�J���_?�0C��Q�mhL/���HU�$
�64�X����_Yv��ѯ�^�,�?6��6ȶ�aS�*?�fYC|R.&���̿�b�� �X�l���]o/�$�Dc[uךW0�y/PT�[�ֲ�˂]T����4�l�+#1�����x��?bh�XcD=:�zY��g_������Y�� �NH�x�x�q���T�p�/���*!��j����5?��q4� �ң0�����#�#�t�ѽi�1��o\��G�N��]��4�^q����~yDR_�=a;��<��N��Bd�1 7��Z>�^�ܡcxᙖ�2�:XX�0�q��^gV���3�ڬz�d������&8�+��uG���b�Qǃ���
�����f?��1Z�q�/k�,���z �.�;�o�����v�ё�~���%p	R����C���+�����t[Uǿ@Uꗕ�#�3��jؽY�kG��݆"&��i � $�=�M�ݬ
�a�� �Z�0�&�0��7����OHʳ�X�2úb嫘y|�@��bzI�w�E,��~٭��w3z���F�P�k�)С�5M$SUa��.���!���\��xa�U�c.�|����^�|��*Q;���;��?��{49�l�>�x��]�'i�b༬�y�����p.dйT�YH=����di�����8�1��ks�(Hv��E�^���0�ɖ�#��6�ηv3��#�'���`Ŗ���L��n�"|j�U�,e�)s����T�j����`១H>d�6#N�Tu�?=
�Wr�=#
γܨ|�ե�����g�IE�}��ǁh�t������.�X�B���z^B"������tڎ��T���g���V���S��;�^L��1'��x֔"�:F��hW�㰪��ZH��|�aM�q��vsH����i쾕u����MYeC3
R���\��/�
"m�͝��n�\�.v�3Y>� �V��Ǥȁ�.F��Ԏen_��+w��QH:�Z�o�����i�YNaԎUz3��2�=܍�7ϬՐ�GagfA�u�ϒ�� �W�U>�	�T���qRe#���P���a��2�8�p~���q��"����c��A,6.�_�\,��n���js��.9�{B3����M.8�K0C�
�S�oF��������oc";/���L�N�&���,��!� }��J��`�_D���缚P��;�Q@<�"��/�4?����$�������>/[�������d\�%�M;B6������������y.А:���*e
���8By2L�禭4�k%>0꥓��'��>џ�!�'��2j��P�۷Ԉk�[˟g�\�/�X!��rN��0��&��qMsˆ^�Q��n�����}�y�&!��D
�t�K)D���V�� ���gў4����<��d`3߇�E.w� )*w/:�1P��5���������C���/Iޘ������p=k8�ý�d�B�i^�ED��}�5W��uw�CE8e�"�59����n��6�s��U��s�xaL	,~�o0�������{��o�
P���{�iۦ���������H�kF��k"��Ɉa����������q/'��.�"�S�Rp}�Fz�rs�c=��D��8�-�ƕEq�ꭋo�H��wu�ܸ��pE�Ҭ�H�����_Plr7돕(:�ߊ��Jz5�f3(rIq����0�_9oR��8I�eE2�M(� 	�v�"���DQ�nܡUX��s�Z8�H���k�۵~@��_V"�)�>���*�d�aǱ%@C�����R�9V2��Sf����g�}Y�*�q�2=
t���H�!��M�xۨ�EB&��l��������Z�Ru�I=�N��l���!��j�q�MEJ�'�[���a��X�m��?�a�e�=ӆ������f���;E��~�$�PN�gqT�1������^���T�w\3F����1eQ��/�A[�b5�X�)̯��ª�~�#ik�X&�]�"�F]�i�d4��P�=դ�!Y�DL��$݂��0Q�������NbX��_��o�<�4\�/��y,�S�e���-���?�q��zL+�+Zs�v:��ti�1�	�9?�����Pm{��ϻ4�XBO/7�d�.�-M2����1���y�JB�u	e��e2���%�
h��45K1$�&И˖��b��8=i���1Ih�0���2y �����B7Jkzj$���RV�I#����6Xҹr��]��C�v��sd��Į�����+�Hy��޷G�I��p�iQy��q�bU�7(8��;�GZ�F�Z�2@�t��}�|ܙ�:��v���9�(+�{��ObxM=2~��w2��zG>�D��װ)��e�����лL���M�|G��W%rI@�b��"?�1�"5'�������GI�v�X;Ձ��d�3�*<ٵ\�o#�c�P�j7:Y��}��jPJ�����t(jRR����`��L�sԨ�(�R1O:uf�iWv�
�͍o�����ql3��,+�M`:�~�H���~�Y5K�"�s��F/��L�#�a'�#'t�-�>Z���Џ��$�^X�~AV�����gPCMt����Z���,l�K���%�o1��0�1�a�V�B]աOdX�![�0�pt>�4�g�s{�]�n���R�GY�@�4> ������8�G7DηR{�ѽhd�g�&��J�n?�VfhZ�4����r�� ��ګcP�(ˆLi(�;~����3� �^QH�U��Dܓ'��e3	B���CQ����)d�K����������L��c�	l�6/���l-}#���I��1=[�VS@^�-u�ڱJ1�bB9������n�������H�sU_�/����S���� ����������6Z��%x�ƀ���\��OH����Q�{<3)GAe�	�"Փ�鰣�vQpwaޝ���3�)�4aޣ����t�����y�c�Y7���AO�n� T� ��Ⱦy�\ ���cPaJC�1�A���R��o�Hma��y�>�,(��R������>Zj]���Ҡ��;�+���(3d�Zt��-�+�?k;��TH���i3�Wf��z�@�_|�CS ����h� 
�i�k}��Eg����SA�cj!|��$+���8��^�b�h����2ǋL�eA��������"��@�H�����-�-�T�Hy�GV�,,�^���~����].eF�7Zc'�D߇�`����xb2�3m�	/�3����RNQD��}��d�z��]�s�"�_o���9�"&F����v>CY�ߣ��]*��OV���+�ey�r��ǳC!��RoD��¥1~?흟O=Թ�qW~9%D[�W����7(��U������z�O�J�9�u�S!��}W��D�w:�<��5F;��FE��y���<�?�� �^{R����\Y90�6���tBkn��o8-�2zVGx�h���4%ƅ-�gnx�=!��O����Z,t�;*ƹ�h'�D�69�K���E��3�Zo��+^�'R#�����6�Jr�H
�[^��z��"S�u�0<-�A���DX\�H����ޓK�t���T�	�4�*
�}�x���h����?s�j��p�E��
O�ē�GT�؋�ʈ@�3}�m��e�l眢 �ͪ��D��Oy��-˾�_��e��v�����M3�P�	HZ@��ӈ&*u�'OD1d��P���<��'�:��n��b���v�? �)M��Uyv�xP�F��Tz�.ǑL�S��M꬧jj��"�V|�G�!}݂����BXL&ϓ�Uxq���$̧R,~�ab:"�k�Ή���tHE��ݲ��@��Y����}��JzK�ֿ4�u4�B����8��";=��K�0Ϩ�u�i�.H���m�d�����V�R�ŕ�w�y|U�$��B�֥w�<\�y�CK�a�d�U�9����i-����1ހ���P*�<-����0J\��,���&'p�}����x��Y�.'�4����'*�r��( ;��k���`4��vz}e��Z�-��uA]�%0�^j �0��$�W:��Ci�^�
�Re�T(����WK}#9�vS�i>���Z�Ƅ������o#���cA��S)�'���c��y.q���v�$�=�Z�U蓜�8�A���@��&���ro�������a���S3'�60뜜Ť1��SʌB8stbSc�Iyu�h&�"�5A�/�T��lpq}�U`W�K��_O�v�8�F!s)j��7��$�����r�$�Tnm�!����^h%�Ay��|=��6��2`3�X���#~q�j
5㺸�q���T�'k�a�Z�n����a��&E��RDT�Y���|M/� Gf<f�?|�bȡ0�'3+�P�Z T���똟��m�g���v�*{�CbWT8f�MȐ�;]xIb�3O��6+׃���$�p�=	q���*���<Hx����&m���P��[�V'� �
h�����������蘒��e��`�p� ����ɖ&�C@w�`!B&���;Q������ڲ�Bm-J�4c꽓�x|�+v#���5m�%����;�"�"�m<8V����հ!_<���E��d~��]愳i�ٔs�$!1f�n��R��>���m�r�WJ�MH��V�����h�Y���g�֬Mq�G�n�@}�̟km	}7�.L&�P���0M2k�l<���}��k�n�nq��K&�8���}��s�C7'�o�c��ܯmը�[�D�O%ߎ	�6�_(�\�\�ek�������S�=���_f-��h�(x��T�2�"�[����d��{A!������+p���Ca�����Tͷ���:�1N$FԝtD�\�O�w��k��h�nh��A� ����E�Gy4Ζ���"W�h��S/��`֧��Vޒ&�����R�\�b￥+~.�Dr1PH�[�y^��c��{j?�{J͹I5�z};�/�d��4}iУ�?�y�*N���N��ry�yr��F���Ѫe��z���k�j�+"�yIb��IR�;<oe�˯��,g�K��ը���e��$�x�缑�gvFI��{i�.��z���	�v���I�"M����@,Y�ߴ�m4�h,�\�(�u#Hc?,6�p�%ڏ��[y[���^���#�9�b�8���$j��L�!["9Kл�j�j�`T�?ԍ��Oo�5 �]zC�-+���܃�g��oSa�]��P�� &��S�V^<@;������RED�k����b�;ppĻ�9l� vu����	� 2L��f@Ӄ���1]���bD�r�$�c�M\��D���_��Z_�883%/��}�ừ�o[�2�نUy�����	��)V��}��&�K�D9�mcd�O䡰+Ɗx#P�l�UW7좊G1q�ب;�U5RE;O|B�Xh7������A�
ڲ�r#cU+�OZX���*���C�ȥGY�D�X��{���d�+jak�l���4I�vz�YF�P	6���"wT0f����ہ�/_-(tj�����)����̆h4��sz?�
�;_L�ʂlTqq#�|"�v���S�ˏ	��t�iB�>t=m�-E5�2�5p�0��#q��w���ƻR�u���`-v��Kh��(�R�Ո����Ք+W�w���˶a��i����;w��0!� ���/>  *���?=�PC�6��-H�������v�`8���y�E�{o\��C�fJr�Q��M�Ꮑ�W[=;���H>_�cӶ��K|�kN�W��5��� Κ|�ޞ#*1Ծ>3���O+�A�e4*�!%�V0>s#�B��D�3`95j�/yz`�Ġ�'�S��U�
��G���ƾ�I��4
�d����#��Xch��G���u6Y�z�����,��es[�����vY.��ʐ>�EM��'_��{P����Je1�'�ՋAT�T�G~1��ʣ��DOJe)d��� �?h{�Q<��"��x�`����	�p��[�=�׳B{f[�z*�'��LQO(��ڼ�z��YJ{�����Ae@T���L��Qy�.�ܠ΀���xV��c�=�R���s �SZcVg'+ph�`ߌ�1��-(B�I��M� �Ϯ��tp�-
RF���n�r�q N=Y6#��qְ�r�d��Hp�2���zD���`�}Ƙ��2+�({W̱�g�k9 Ja�:ekQ�s���,[ăH�mu�B�VcL�=�r�`���MԦ��vI�}㼿��XZ��rR�vo��zk��B��@�5���O��=v?	��+O���n��9?�Y����JHk�7$�^�؁������BE�&l��=|��e|?�2�<|���+%�$�Қ�"$^�4-C���"�e#��Y9'����������Z$\��6TR�	wwõ���^�ȵ��?:o�V{(�F��lp���0:~��k�Dl�~��o�E���Bo0* 2�c�;Ξ���cx.]YD;�z� <^q�t�:Wap ���P$BGWME���ov^o�
jS~Cq�H[�}�<���n=�eqk�:{�����c��%V^���h!��'��7z�J�4QCL\P��K��`�EG<,�^n<v�`��wFuv8�,;$�^�t��ӟ� .�[���^J?3��m��)�o��= t��wAe�'?���A��+Y���2$���\D��QS�(�ߒV���_�ǅ�4q���AC��?��og��b Jp�o��>����h��-�hi���$�o^�xs���,N��������}?����^�C3u�>���_�F�vT�$�������e�QWƬ7<��c�Q	��?˃������>��m�l�6(W�Vs�s�_�Bo�� ��W�Z��q<�i�����r�!��T"W�����4�F���o�J�h�uxۇRa"J�9�����J�7�*��C��vm�n`5ɝ���Ϧ\mX?��趩������f1�w[�H?7�1�'��*��.'���b�G����F�?j�pEŉ��"�:@Rt.xy6p@��F���F����=��լ��r�?��OG�\�����=%�Y����� G��<�kar=�l�x��;�p��^��l�G1���
7PVPB�)ch���E�ة;7��ǯ�$�ξ!�ڛ��!Z�yd����Y�a���V��t��X��X��t��,�8��X\��-��ٌ��عv�x�c҃�v4 t�N����YX�]���A��4v�#�W����5�˲��b5ٍ�L}oͧ��`��0KC=ȑ��1�iIͣ�?<�נ��BK���"�8l��)�b-���/�A�%�:0'��+P������<L��%O�x�	�	�����A(*H�f���j��|��溶�}��=U[݆}Zmh�ev��������Y� ��}ۭ�LK���k���$;��K��g��2(3���A2ׯ>��VL�3��3�6�~�B��^x����h3�etvZ�5%����x�e��CJ�z5�{��	ͳ/�	�,�AdLhm����Z=�Ni_ے)^:ř��j(��UX��e���co�j�䱞T&��Bܥ�_m���b�(�v>����X�J��8��}��O���o�P>7���Mu.Y���F��JJم:_�4�;W�ߟ
HH���)K�� >E@cҀ��J��r�gȝu���ܞ�?}Ӫ�֑9K�qgɱ.i��>��Ǌ=��Mi� �w÷d <d�d7�T��3����yO���w�ME.P��]��}k(џ�D�r`a��4(�r��T�'v)q�zCYT����P���k��r>[e����G� E��q��U��7dȍ��e�up>j�e-\�"n9���g�y v�.��iw�,�2O���I�D:��ŵ�3�6\�/n�g���NBHn	Z��CVe�W	L��恣�{������� Y����1�]�{�������+�	G�<�Z��������E"����
c{�J��lbUW4N����~T��=B)ʰv0)�MX���P���$FqZ�l�<���ez���C���R������c��3�d^��+�)��z�Sr��"IxԚ����4���;�Z�*x�����v�2�C��r]�4���q?��,�p��$�BM�j|��7�(�?�H̝!3	 LP�6�����̃���o�=��M�m���6����Q��X(R��j|ݥI�ʩ�
��D3���T_�>�FӨ����D�^�K+\�5�b�b�91q�E��ƱǦ[�2?-=��.�nQ�-��0�ã\���;f�y�9�3��V��S3M���c��ƽmC�y 2�!��n,�$V�����{\;wL��R��*t��-R��	�Z虠��Wp��B�⡇?����I����_�9v,Ͳ��^�/��ր��C���a��$י��?�`�n�Tm5[:��T�@�Y�zm�`Q��qh.J'�v�޳���8�&qE�=q�:�P�* J����	��R���`����sp�l&����}G�°��y��P., i����݊݊�g~C�F[oK�S03�WCZ?�D{��S=�s�{(�<M@�;0<�n��3(�Qd&��R�7_�r��2��ד��dҚX:�<N�y�&�:�mrF�A���ۧ�����i�&�fy	;����>[�=~QZ�I�r�"S�׿Y��ɣDňpI>��('�?�V7��*�2�+kV��m��EǛ���[P@���9�w�#l˂D�:vFr��juɖ����wA��Tu�q��ij���-9���?�<������%LF��v�%�^E&oI�$��z.���ĽJ&�-M��q��eR��[��d��(�A��+өDH���s��(���sJ̟̕d�17��=�.���C�5#�v<A4 BSaa*h�����KE$4�V���O��*YhM��)o�a!�;�y*4�t6݌���8���3$U:�&:�%am���?.x`�c��a�I�	\=6l�	.O3�@�J.#K}1��"DL2:�"��W�	c`��O���0���1�(���ڋ�&ʍ�;�M�������3��]��k��O��<����0��$0O=h��!Р�^l0H�0&���ww�d���d���N`�}���"��뷵r	�Ly��Q9 �˚:#]�����k���N�8Op��-_� Gç��BaG�[�Or;q�
�Q��:֗�`��Ȉt�z'�Q�R�^h����\g�N+��1����P����4b�Cs�P�����M^�׸?{��=�S+�Qvp}}��%}�i�"ُ#���y��.3 .|�خ�S��<Ul�l?��FF���x�t��r�Xf��a5ǩ�X���&�@p�����xe�t�Hjν��9$���x	���FfR_�����'t�U?UW�B��M d+	�ܰ&�kL�-��9����k�=i�b+�A�@A�&�NϺ��(��lD���b��;ͯ�U��ѳ���ҁ�w��B-&!�a�WU@���Q�-ЭS
 #�s��~���ȟ4(Ij��4���D���+�^0y{���^dj����x�Vq��oOb&��z�|͋`H��J>h�;'de�- �*�&t��j@�ٵ��T0w��R{�dO{�o��o�>7�ѭhHZ�����r��-�<�U ��%tcm޹��k]�xpɹ��ʢu*KRxUc������Ϙ]����N}I\�4o�2;hP-*C+���GQ���d\���
Ө?�L�
�
�\qg�K�0cbe�۟�ξ�\!Z�e^d]�U_<5<TjxOٞ(;d�E�o���T�W���?�ث?�R�v+��̥/�C��S:�i�� �	&]hw��s���r!\]E�SV@Ϭ���Z�.S0�l�g� �Ym��&�G��	S�Z�~�^�
T/�5��#�#�<P��0��C��}����߉�>M]i$���{��s��2/�k*k��ѐ���ߦ�Ur�¯O+�pS
��4���i`�٪�Z�sY�k������l
�C~ͻ�)G!L��L����a�`��I�l�P���7b�yy[��6�Pe�g��C�G>̼j`�<J1gW��a��q�_�wpD��+��\l~-+���\[��m�@�+x�I������*��!��~��Rx;�
�R�w� �%8��`1��8Ra)���@G��\wc����jy2��#Q<��}��)��8߹q��5gGR|Ў�w��@����7*�J}g,M<�Ѱۦ���?%��u�r|���;��B�}e4�*�n�h�s��:���>�{C��É� ���J<�"���JPF}�M�)�������D3�����z��9N��y	ư8`j
<��	h������qJ���m������fY7�u�ׅL���k��h�t�sM
�~$��'�B�d̹n9cw#���	�*v�T��.�M5/Rc<�(��m5�n���*�Hb�fWQ`���?"�g���-�8O�����`�$�VA�O���6(�%ew��Y5��1�O��i��٠HP���>� 0X�Χƫ�Q���T�<���W���P�`�zuñ��%��&{���\n�b��a�ۯ�S�#��H�]d�<T�l���YԾ����cG�|�,h��_\�rZ��|�x�Ϥ�+�W�<����n�m!}��-oK��>�ܦ^N��y��]��#>�QdH�hz�JVa������cS��e��]�Қ����9T1�a�</v������[��׏��E����M_�Ja�h��X���7<<�F{+�R5�o���� �{z�]q
C}���Zi���_�S:�ݥ���Kn-��n�)��X���W~1�/dD?~*qݥ��ȃ��ߥ1���p�ɵ�+O�n�t@�:�Oc�C�<� =��Bv%P��a�_��N�z��]S?��?�)s4:&oz�\���epe~&(�R�dV��d��r ԝQV@k�Z�WN�>h�(�p�������6�*5�e�	Pg��dnn��R�F�q�H6�`9��Ns͉_ol� ]?��[k2]�ӧ�NR�+���X�2%i���j��g���`$���tS��;� [��	��f�0��n���b]?������òߔ�)���t��nd˥pF���C#D"���05!)�0��qv �N��;{8�n7��o�Q �a�n��fm�s0�b}�
Ϯ�}�Ċ�R�]k��um�>��!$��I{� ֈ�b��*Ή,��[hX>��YKm
�lv'�yH����R9�u��&��5�-E�����"�s��/tK׉b��oyKj6�m�9eд�ʖcbX��L)���rCG��D��P��c�zڶ�^�J���H�`�R��H@�ɦ�v��	~��˂4\����i�U�N��,�I\6Ǐ����@$d�>�����:I�FQ�ˍ\���� �hգ�=�T^SM.ON�G�K�AҳG,�JM����F��StW���I�wN �V,�T�N��T�Ps��^�u�ORM忰.<��}]�
�����;��$=�'Z��ْ��'Nw&���O춬�0�c5BNC���%�]�31��+�).�4�MRy+ϒ��E���4�mL�@����F��H�)�6�0���vlh_�Be���O$���d����c{$�����c0���-"KVK�B����j�_�?c�@�<Ao|6d0I�|�eXcz=[�F�	��m�lln:����~1*�c��Y�Mo��+ۛ𥩳�����GԺa�D��@��2m��#�7M��_*�Ȳ��f�%��+�{�<l�l��z~N�#�d<���.�����r珝_
�O�M��lG|6���Q
Xx�0-[�?�}����I��J#e��-Q�^�\"[�X�|��ׁ��K8DW'T�ѺW�,zX�mY�UZ���z&s�u��L�w(���mo2\�E�ˮ����W�ɔp���2ϴ���.��0İbf�HCK;}���x���d��0�G*�m�B�`����v�&�<��(VTTAL.����eS=k�1�>3�q��|h
�\�'����z���[h�u=�j1��M�%QN��,��IyJ�><v>~�Q��@�`��k�tז]W6�ç��/��̞�C��>�۷���� ��uc��"Dc��t� vB�uWݶ@*�%��17����R��o���rY�=5�?R:ʬ��O�"������h��8�ڤ���Yfή��C����o�'KY��	��E�LxҾ-ǝ�z.�t�g�بD㎐�<�{
��m�ܦa��F�	�x���c9��'S���u�;�R\,��2IhC���b��m�_ XUg�;��h�G*��YD[��ؙ�~�
Ǵ��˽�,[#��'�"��4W1'�L��҇jN�۳��+���Ⴢ����쩐2�۶�z�2FR�V�4�%G�p��	�:���ŴJY���B�`�1�#��G�HF=u��\E��kZ���y��u�N����יɟ?w�W�d*Sגw!���g�c��h����4�� �]t�<4�Fޏq3�=<3�y)�p�r����$�gn�97��X*FS[���} �T�P���1/���~k��*��W'���
��?x>�FTz��\�Q��l�=~3��1D���Pe�%�#�k�彻x�E�%�,�8�d�'��T&���h�)��Ұ�o�@��ߜ��P����~�^�_����";j�U.�@}~�[s��O�0�mQ��w����5:_�kW�y_�	 v��3�U/���|_�䗠�a`�P�-!��,z��I�1���f��@_:�Ko��!&8�.e�ˉ�%v{�oGC@�bEծ[����5�f:�#5+>�Ӓ.��Qd�@C*y�h�
�$ʋWث|�1�\�����j�WY<&�	^�!�� �;v�/$����u��ͭ��D�$�D�]!�zc�Q=���4o�����M���#��1���j��iV����N��1�����R	[4��ͤNiw��x��4�
L�n���tr��2WE��ŀe�'_M���>������u=�H��:��B�Fٗ������͛�Ղ��v��'���m�����˞��lcE/ՈatP��#�l2�eL�=fx�����/S��S1��Z��'�"�����4c}6'A4j���Tg�q8���_�.��s���\ƌ;�Ӭ���_�8�h�~�2�z�v�t��}D�:ma)���f�4�[3�K
'�����U��m������׫EA���Q�S)M�dx���Ǧ���;ٷ}�I;^�<2t�_�{�w%�� J�d{�$�n/�͐!������.���w�b(��O��Vţ�>��#�{����U�״�"LT�)S�;�_�6&���57	��X��C�.��bΣ��#���ѡ{����� � �rp��D�.]���ilqK1*��@���'e�1q�����|?l4B�C���xG��첀�Q77~j q��[��z.�z1��+@����y���D�~���p��nH�Y��SYÉ�b����x1������1m����N;�rb��ZJ�XpEkw+2�L;�!����DV����>�7 ��s��	ߵ��/���ɇ��Bl���gH���m�ޚ�Z��uu.G���|E�Ox%�����Wi�A�V�d
5-2	d4���HF��M'�C��)X��ծ����.��!��I�Ԥ1ƴ���D���f�i���Ʋtd���N"xcVA��t}h�lh�z�2�2�]|�P�T�Y���B���5z���$�ta��Õ��joGY=v�/²0��h��A/�>�s,Q�Ȋ���>5����Α�X�-���ie_��;a��Ԡs8��c��>�/Q�Q&�] 3��<�\��B��w�\L|��zC�دKD�Ϋ�}n�2�J�����Jdѽ$'gr.e����'���,�!O��|Wr�n�G&�W�)�"��b[�E�T�*�:�lw�6��a1��=��,��g���21�1�L�ن� Z���eo.Ў��7��G[��`p?u'e�s��di��'��4�Y��:ߡȖ^�/�=L	O���o�%��8w��yE��О�E�?g�J��z�4�$��"bk��vv֚��^��t&���O�
��}�X�qӽ{�;l]��[���LK�(a��=j��RS5~��ɥ�8�<@;�}؜�N����ý��Y�,	�mG\~�z-T��4�q�K���h/vA.2'� �W��Zod�q�m���B�}�F��b��V9�p�=�;��x�}-<�]Kޕ����r�u�L�$��e��#Ϊ��-�=���jC9��x��SIm�F��Ǫkе�t~���+��� ��=�pA;.�	�V,F_v:����V�h�.��{�	��`]ϕ�l82��� !
���z�2�JN`��ɣ�L-]<	�J�S����7|z�<g���?坥��Џʥ������)s`�>^�NXT4���M�Q���2�M��9�*�钦sA˭��H,��P��QD��ڝ����N�Ly��PO���>�N �xu�oDԥ��U��s����@�=b;M�R��ᱬ��	�k�f� Ū-��f�z;�z�I�e���<Ӻ,Aǖ���\7�<��{K��f���m�ͬr��\'Ӕ��g{�`j��E�9������
��D�*Y�pj:�m�͒��c�$+v�]�$��0ͭd�@:�I�f�[,t��|=��n6
{�9�q�9��_n7W�8��姏�}%O�j�<��c������$nc3��r(弐��,c�mHh���W� PS�Y�04�|��O�M�`��ၹ���C��Ω��i����n�%��$������|�N����3
?��uT�,ڮR���	�H��'}�?'6(-I�0��M۽2P����!x�7�PN.�8���u��i}���ѓs�DA-�:Z�B/��ʾ?g�i)�g�M�-LZ)w~|����8�65�m�cm�wu�h��S����v�A'�X��J�k3#K���h�;�����X�r����G0�HJ�1��.�{�n���Ņu��vqG�F�˖���饌Յv��*]��NwR?�X	QC��r�p!�T��D��j`uC<bmKy�
��nUL��?v-v	fcxǍhq\XǶ�������[;�_�
lū��8���zÛ���i60���U8yHf��A��S	%��NBdU��33U^1_��iش}����1
���(y��d"\'ɺt�����ao�E.<��k�ț�;��}�M9:��l�K=�b���{T�02����=�I�:�A���h�z)��\��'�j??��w�:��Bl��f!���|E&�	g7ĵ��3bZ8��	XC_L�u��*Dx!�֏浸��֤�A���>jvm����"r��jo)J���w0����f_��F���p���Kf�T(���O(J���nB2��V��g2H��lx)� � T�����@�7��#�����с�xq�oժ8�w�J���GՖ6`���y�回��K�.C� �s�i!�,#vM!:S��߹aH�����)��QU��[���4�ʎ��)��ė #}����nk�g������>H��l�/!��'�P1r�<��{󈿏'2�݄ͭi��	.��_�K~t����/2�T�%'�K��=���e����g)�j�lZN�yv��pF�ѹ;F�	��²\v�5�6�y.�@尵�S������f���	SWev�&��x�x ,���>��E������=��EB�sπ��R�C�$-?�BE�Ͻ�K���qd���ɺb!SZ��i}�z��Z�ƈ3��w�j@�8���o��;� ��yl�2�'������E�"��nlxn*��Wh��q�� �㩸��iN��)���d���n��G\!��cf��\�v�$�yû����<x^_��~�`�_A���I;�Cuۮc+Ts�l� �{�D�_�)	Y1B��[x�?aŚ�ԡ� �bX375��-�t�]��i�|9T���~9��{U�`!@�pĿ�~�`o��^?%(v;����i��$��k�iO�܆�J�^e0$�%��?.#�Ds	��0���` ��=��~�e�y������hK�0�Yk}$�f����o1i���taF��z��1՝����4t9^Mj��0՗��m�jNDk�������n���D�&͎��fYU�o�}�I?LG��YI����<��ޣZ"��-�"���.p�U��`Ǡ/��ɹ_38����g�s��C::�89j������p�)�9�K5K`%�0���'����f�?�1�<̺4������B�H08-�  ~�r�y9C��U�s>��p�K5�#D��J6�$�a}f��*W�LV&��ꎐ��E�?"���3���r�&���}�aEx\k_��/�5/�T���!�d��8H�~��Mi�=�Ufltq��g@Ӱ��}�27	6��s���۠�u�û�F��L��`�~��)�!��0&����M�� �2V�]��0����H�PQ��b��c;忓�T�ɯ�H�<���ŖWvb^�#�f���6!�W��[����c̑ �FE����bgSi��2_�s*n��Mu�JhI!�x����),t���"�\ �S-�<���L���jV�[o���KY�Dl��-ʗ�"l5�Ogq~ɼ��v�m[�(�إ�vm7^�sԭ��h����wcùy�rT�x�$�
�"�{�����#3�W��A����d����X_)h���Ix����4�LNsV�R�S%���K�M);��R�y���a�$�������V�g%�G�/X��T)�Qs	�W�% G�a6�H^
jg��&ؘ��w�W(����~+���>Ԍ�ip�Lލ^�ū9���4��&�3;�.�#m�=�jS�u;և�Œ3���H|���Z:�_&����x�K2\�t~ ?R���$jH5w��(�%H2I��EB���*tV��˵�T�-��_���q{����3U���ð��*����.�Zӱ>߾�i�8���)&\G��'��Is�Z2]�J�٤��c<)��ŧ}����wU-4I^x&q���AI���5m��aZ��Swa�����l��%kp��o�k>�&Kq���+}ks��yR��6��>&���B`y�����o�^ۆ̯��<5G|oPт���&Ǧ.Ǣ��5�$B9cu�5�w��о��t�>H-��Yg�/��IB	�͓/S��hs�e��>Ƶ�i�O�-
��v�����PH�MI.����:��4OMn��Z^$Z�D&g���%M����KW?񍎜w�	���(�
�a>����	�I@%���QX��#�a��I?" ���X�5R���H	��7��7la�%V��������Ը�����r���:/kv�sr����Y�Vԁ~&��/R�)��^y�2�)��_+�������fcW�"f?��ar��0k�Ni��
���y�>�$�_�1^�A�.U�������W���2*D�K׸�[� ��*{�@����,ሜ.��%�3|*`�2{��f��{�A�mG����ZJe*�$wZ��Q"� ��ww��_:N
1�I@'����?��z0�^v���&�ej�p-��x�s�Y6���X1�#���BD�u��l���������IBȣK5���$R.3NFS5P����bX��ٯ�*���CA�8^����3	E'?�O��#��[��>Q�*�h�E��؊̰����7��䃫~�gr�p>�ul�����t����*)�(�{�'>Ya��}��F�f�b��&'�	"]ٵ������?��aj�֒����ċ��c�[o3\��^�un��<��z�FQ�t:��+{y��i���#��=1��%�3u �n��$���%ӗ����C6�z��<YN4�{�{.����:j��ֲ�)��@��5{�<����;���EY���\.���c�@�"��ԟ.��͠����&[A�*ZX�m�b�js{�fYH�TO��k��
4C�"a2�P�V:[�~,L����K4fP3���uS��9���Lbh��޻��>�$��Q�����k��
�c�8-b
\�N���:֡�߈�H�)��̼��id��ʣ��ԑ���Bj/F^ｄ��CY�\+	�#FHm*�y������[�@�dh�V�**+��}����9�y��3�z"9�8zV�jZ��	?���i�Tjo=�t�-��AK����&9��6�� Nl�	�T�����>@��Ľ��K��D�����|�WJ�| �TVD��BXq�$Jb.�!RoeK���M�	����c=����� ŞW�{tSWؘb,��i@�V�a��a[��q٣\ �@Kp_�_�>���� >��ųɩ��ֆQ㹷3�����?�-�˂6��D:��j)���4���$x�U�� � a��j]��MC���<[#����R��" �}UU?���n��q))��&_�����7	���|�֬a?�ִ�Ȃ1))��V��O��i
�2�v�����:�B�'���\O��\@)�"��(���iC5�/k�f�z��_!��G�k�u���Ԧ�S?�C�Y &"~m2�O�ܶ����LX-c@S������ڙ*�/����Ȑc�y�)~���#��V�db�u:��>0#�������m!�N�kbW�ft������@�xl���4@UM�q�$�""�����;��V��H�b��7��R��E	R`}�bI�=;�CN�8Q-�����'�F�ց�d�RQ��F�)BDy���@[�V�rFOʫ���y���G38�I�_�ޝ����;���m�TE������b/.^nlB��<��ν>�ۃ
��0�?�?r��2�2��9?cư{����5_���_+��#��M���}�M;΂( ��AC�c}Bb��;t#����;�"����8��)z=�(����x���i�bo�W�QU�9���J\3s	5�T��/����4$E�3��̗y�TF#���t�/�˨5?�;����r��fy?��T�q֚hϽ%����TR���(|n?�훺\�"b��9#q�e7&���]����5�h�e�����_����vҝN����,,��?�,�WGOD<���i�.5:Ăj��1�o��H��߃�9��%Y�=y9���m*��)����6�vu�P�lໃ<�Q��N��Mk)Hh���ʨ���b4i�{��⟡�c�e���*�E�	4:O�hdS���{�8Iu��q��r'��	�O_���a��u�Wތٔ/����O�4I_��_+�T�F��UaR���ā�m��7u�L�Km<���^������'V���5�N;D%�h�iE�J9���9��đ|�Ԛ�1�Չ�I8�)�~Km��W�����7��J����f�쨨k�=U�x��Y��6*T�=�b���$���s}(ܯB�9�ؘO_!v�U4O�PH�ٲ�`�J�]��mm<s��v�y������<�Tq���o'E��"Q`�ҁ��\7>�H !�C@�蘨k@절1^<���ǿ��;b���ַf�y5�tt�n�u7΅-ۏV&��Y�F���׽�����=�ĶP�8�wD'���S������s�D��>|f�ck����:�$�+��5R4��_� �ѝ~5��|�d�6�On��]�~J�6M��	&�
�Ҷ*��iЄsfT&~)��	���j�MAl-Ŝ>ĳ $�F��8�{D���5�2ׇr��dZ�c�Q�_�V��
�C��{�f��5�����a^����@Rڹ�c��fБ6"��w=_ܠ��l+/�͵�t;l�'���w
4�|:1i�l;��"���I��d������H1����ni����^�6�	�����_i�gU���\�h�c��/�1�i(��p�Ϗ� �I�n@\��)�xt��`Qv5g�L1�0�y(���a��5!a�L.�J�K���U��kP�&��f��A�;
.�!��n�G]ei� �4>kC��>�˘���X�GJT3�ǝ�}؈�)�W"��MV�&������Z�U��䔠(���󠚿��I�r�nӃ�P�^\ja�+�Gx(���+)5��1�cse[�ɋ��%��Ğ����0� ُ=�v���c���s�ז��(R.c�d����T`�����7O���G�'��ҩ�&MxC#'9q��O��σ��r��l��e�t0h�(.jd�x�)@j"��kz�P���x�����ԡ5�H"v��u%<�ҋ�!�i�jrƆ����	��$�.Q��×�Qz�M��[VH�B���n ,W�]��2�ݲ���b��v<�GC�<9��i��YN��v4nO�#V���$�n��a�,�Uȫ��X��D8���}�W"�Ŋ��4��d�0ie�����HW ������b7����I}�/�ǚO� ,���Q��K��xt�����T��|*�[����ʥΉo�/;�M��1w`��x;�%ЧK ۏ�ū~����7��ft�e� �����m<Z"�h�}����r���я�2_��3	jG��n&��+]y1�U-DjC�Qhs��X�N�hI �x�[���v�<�t��Ԭ��zK��y�f$H�/�b�#����C���'d�1{#��T'rJ���4�Ո;f0���˧0:�ϋ��YS/��6e������D����Zf�`~��0�Q��a�PPp�3O�̉��5��sw�,�4ƍ�'�o�M�U��}���W'�[q
-����ѠE�8���9�n�d �C�R��(�� g
��z���ğ0]aR����_`�(�H��j�V��uE��=6	��^��] ;����!m��ڧ%�g��!A+������kH��q���v�&ȃ|P�ҰT)�gSP��X�� e0w�	ZC�p.|r]1�GƏbס�Cqb�V�{��̡����;a^E6�0+�q���D�|m���2Y�l|�X�ڴ��Mɇ�s��f�IYG͈(K��-�E~�r����$`UT���t#^�r������ U/� ��u���z�1m:�ug ���6�+��h��s.��A�����6%�È���G[)�}f�D1��[���	C�e����Dj, 0U��}�H���ˑ�-
�֋�x�1%L6D�/R�c�ׁ���N�[�cP��+0��q�Q������KU��rx�GdpC?�!�g����lF�iT���/r��G|C�XS��Ͽ�&wo�V7d,sǧ�B".6���<�
Q���R:0.oi�ɚ��Ƚv"��A��}��!?
���uو-d� ����\���O��C����}�p��j���P���U?o���ԞƇK#� ��[��F{�M��_V����b�����b♳�� ���n�/�:��~����W/�j���+��R��;����+�Z�院!��
�Oca7ņX��yf�S�q#y��:�B�p�\;��$g�}��}g�����T�Q�98�:0$R�NV_z`�(һ$3��&Z���S^؎i�X������L�"�rґ(�g��� �跠����wQt$d֎���l�ڔ'��t/Z���n���&&޵2�o�n��71�u�l�vtNb�W��OpY���g�S���p�N\5���e�E����R�}\l�)�8�k��`9oív'a?�4�Kԙ3��7�c�*�`	�W��l������] �u���W�TT7tG87��֭|�j��l��?���x���n,��bC�M�#���G����`��S��sA�(�G�E>Ni������̺��_`��dMv<�uVQ�ܧ���y뀕�����*��^C��v�C��豽�hP���/�֭�>�T��ge9��H��;���k~ڷ@�BJ�\��b��04�a9p�x�r�(@���_Ml4b,���vC��
L��-ñe�Dc�`舙��$
�[�HT���γ���Z9�Q�6V��������j^P�>,X�Y�$� H�%z�
����0�j�ͤol�'��Q	��H��h�c����R�5��^3[8U����$�9Q\��ց�H��@Z��p>����l�%ƿ��բaT}�s��&f�z�ѥ`�!<���L��RΕYnS�l�~�!J&����(_�Ƽ�i�_�����x}�1eTM��0�c�q����=㋓C��}	 jgr�4��juC�{��w�D�޸�^L7�0w9�����1h�b9x�9赟S��aB �E��*j��(ʧ�C�ʏ<� JȌ�2��[��M������C����_dKZ� ����,�mq�ɋ�yL��+"��9��cD$�:�I(�`!���;�j��w>���G�K>W�R2*ۙ������o}�9��~Ø��u����Y��`�w�27��`݃3Ƒ��XK�CI���f��G���_�57Ʒ���,:��U��d�D�T����v�r3�f?�F�%� �Nf�Ϋ 3��xi�a���`2��v���v����$�ƣubm���&��͆3�԰��A����`�L��o)��]\s]�KY����@"g�ul�X�ϞDl���ԣ��()���Q6V�˺^��d��(*���Tn��Y�'}ቹ����U@���F�2S@�YU+��u@�J��{�ҍ�A���g�&ӿ1T]{�E��
K�0{�%Œ�B�@A��U�]ۉ}��uY��� �)&�nG�s�z��E��A�1)m�0���m"
�zq�J��[�ok��{�<Mm�u=�})�]ˤ�(ɯ�,<��,��I��d=�����'���\h[�\�4��$�d��,����G���y���$ ���$��BȀ���Ze�@8o]��Dw���P��#f+c���7]��KT7�O]�_Nm��+G���"Zeu����������Sy����u>#�շ!\h������Az-�Ѽ��ro�� ��� ��qc��>#b.���s�%����tg���>i�]�r�I<}�
P.��M�%yi:|���E����Iנ�e�H���૎�Q`��9��-��n�%M��5��,&�?� ��X-4�g���y�߼[�0w�xi$���7$t��9��m.��l����I4��@JJ��U�V�S�1�O�{M�����$�mrI�.�	��z:x)x��F�(�v��'OI;�m�RL���M�t�r5믤�� k�'h�M����,X��	7�� 1���#�}D�HQc�a܇�9���O����R�����������(����U��wF�/�M��HL䰉����Oē���d��J���2�}�Z� >�����A�'��5�V���`;qC"h�}zT�}�+���>!q~���V�'�#�A ��Y[�^IX�*�z��z"*f��_b�c�҆k��cq& ���]l"X���<�)��g9%�(Ȣ8[�VZ��U9�.��R���{��-�l>���s���Bs9���?�D
��᥻vnQ���hIG\�����=�h��ޝ��
�N9IJ�-��Xo?��93ʼ��W�r���J�X�v�M��*�u���i��jh����ʍaz��dɬ�C��b�#����+�wɠ���G~\��AF��{��a؀T�KZ���E�y�q���<؟��1�2��i�vU^#Cdyc�C�L�K�vC�@����E�+�~�^0S�t��j�*.~w��[�3�;�m��s~��hͥM(,܌&0�x�?�l5��S
���O �T�������5,9����h�ޠExv�'br��q��T����l�p鱞���x�A*��&LԦ�Lߚ��+pz��l�������k~���B��ۏ+���
l�N��������lp(3��r���&{*@\cdS��5u#,x�<�k��\wBFb��?u�wal��9��QQ=p�q��}�"`��z�4JY?�>1h���B�����b#���:���!������Y�Ӿ��� ���}�+k�_4��)ř;2�����v�:�V��Y�e�JX�a[�[�:<�q�~��s���|!MՆx�X�

z���:ڕ��:����({�6V%��SC�F�G����TDUQ(i�Yo�A�5+�ׂV������͆Nť�X��Ҥ��Eן߈+k*�J!���h<�ĵ.���ܼ��^"���FT���A���мiN7L61���Ե�S�`�']�CeT�;��=ʬ6v�Y=fHQ����tf�z>��]��dk�<bm�����!�wh�,�=B��L_x~!�D82���;�(��VtiJ%��w��f��9�n�Q�� ��J��.�\p�K�~��˺��Ĉ�ZebZ�X%��s��!6k��DAJ�TA��^�G�z%��oִ�3���-�k�T�n���g�A͵[���{����x���dȼ�"u��o0�<_7č|D1��&�ʎ~�ձS�F���^�tjbN]��ӳ��j1�MWv 1}��j�!쫷\����<���y�M�]c�-è��;�����K�|
��Vߵm���Se0�TSd��ΛZ�K���C�̸\���j�T�p��jɞ�d1�0i��PO� �؉H����L�L����|d�qu�Es X��B����f��F�(P�"u�>��-�]��98��0�4F��㚗y��v�d�Q'r'��������?Ԓj���h(���P�06��G�oP��e���(�*��T��+P'@ ��oC��	�^f,�Ll��2�#�Q�k>4i?4g�q�Y��4^ݸQ
�t W���"�]��o�>`�X:{V[.��U�3�C3��Dp��kC�VYzS<�4��Eԅ�Y'��*���en<��2�F�m��#�Y>�׫�Q��_�]���#�N�{�N�T}�v1u�V�0�ԥe6�.Ry2�V5#��B�n�*�2�./H�A��=+�9����=>�iK��дo�r�u?`)�|���+�����s59�=��r�����WH� ��<[ׯY�v�ǟ�hv���,���B���J{����i���!I�L�:t�|��x��CV���Nle��,e+��.��8���9Y~<��du7ww$08{ՊgPl�����1'o�Қ��w%^V��z�<�8+�3�XT٘���/W�W�YWn$s�EL����c�e֕n��f�!��^_��5�u`⁾�QT�_7F����$+Y>p�<t7�_��'���A�҅���vn��ؠ�`�|���K�;0����j��,��#Uߩ����\�m����!Y�����UZE�����E����Ѳ�p�t�|0e]C���3P��4n���z晡2g�U;b�fF���rNA�~G�8|������2���^u�K�_m{��P��ar�xhx	�ˁ���*dT��#�rc�r��8�c˯�f�PD���,V~h7!!t�XyV�'>���u9Uhn�D��S%D!Z���!G{��;a�Le}p>g+����Oj�(�
D�R�MO\�|�Q�+�J�꫗�n���.NȖ)�,�w2MA�Pr�}�K��/b�8��J�s�5j7%7�5,�j��Ɔ���n�f����c;q�	���� O̐������pq����S���Y Қ��27L�95\؀���O��`,]'�8�1�4	3�@��� �\�8o�kQ�XL~7�6�V:<�q���.%=�p�pl5 ��FMG�r)�Je~ ���ǯ���(����h F��Ó��C1ly1���m�ݢ)
��z5���d��Vھ Rݎ�|�9��Ȏ��<��C�Ne��#]բ����(����Iĸ�^�@�=s�g�13�֍�����C��?��hY1+���x9P�B	�wl��� �%A�J곓1}c�y����Ǻ.�اz���.G*��/k�C��> � �w*2�l9�}�����Zy��	����l����� f��F�/ʈ��͂L#��L��.0�ݻU�pbZ|��9�;��1����t1K��S���T�U���k�r�^_�����:�����w�����
`M���:x[�B!�0����Xs�p���J3���s;Y��U�2�eRqi�K�����}�"���dQy�5�Va���Z��Ъ��F�ij� 	c����;ٲ�pIXZz��D�dgtO3׶�J� v�
<�]�iØ��"(7�/:LA=���iJ%C�gO�J?k����X4L��1��ũ�>Q��)�Aq^��b"'����b<����ZK��[�o>�#E#�S5���/|���݆���N+:��ᄞ�uY.��y%��`�����a{"�<�傾,��O;h{ku���y0����UXE�� ^
��:Y9 l?*�^I�T�q��7����T�,��<���s�O��eP%�l�bf��AYX3+�U���V`�
��:H-����0��eo V�����o��H�x�6�� ��P���;�̵ug���w��f\�Oĥ_�t>`O��,��E`d���:ǘ��-, VT�!�ټ[C�:&Lj �����սz���m��'Y�w/�3� �A@��+&a d%H����#D�UK����@���w_"Z��k�I̅�p��HwJ
J�}&���6䒍 t#��@���3�ߺnL�IKi�&�|J�0=��ۥN܃a$�q��ԻK�U��0�+nj'X0��` ���[���=DΊ��׻�x��ӊ8�f�h�ORX�Y�p��dsd�&�l�B������N���&��&���M�����	htW)ĥ� ��bT���!MI�����qr�q�Wg�Z���� -�1�C	�F�����ԅ�G�����}��Z�&�;�Ұ���`�����c��[���(X��F�3��Лz_�{��(}�>lE�Z�^,@����Bfr+��)Y�la�%S��R֙l�ٹ�=�O�xI*X�����uܢ��j��bh�u-�p���	^��я�d��SS}���t���uMA/�� ��DžA-!�h�p/+�9]���P��+z�;<�����
���y��,q�B��9} y�0�j$D����X�Go>_E��x�:�'��!R�2��S����%��p��hq��>B>��-�)��I�h|�+�����W��j'IE�}���I���`4�g��y���<=���]Ӄ:�Sv8��1P�������L�'�����$�7qS"�$Ö��e����WE�4mF5�k�Z��0��(�&�-Z+]�g�n#7Fc�y��2��ŷ��<,��M{�S��ߎp�x�5��m��0Z��899�c4��j|�pw=wufLI�! �;h�ZC���J7M4��*������V��L��}.�Z�VxO������)C�tބ	�t����5}�NW��2�ۅLKǡ.�r��t�I�jڶ���*Ţ��+?�Qݖ��G޻��~��l�}�Eh	��n�����{���&�XF!Q����I��+	�D@i(/k�8���=��q������U�͠���{��p�]�t�N4�n;��@J�;h�"�53����`���u�y�Ѓ�a�����m�-,B��r���PG��w�nY;q+�����_��6�ga��j��pigry�Y�:͕{��ugC�Z����{�����$��hÌ�9��?oux�IM[����h��Dn�EKj��z��Zb1>x�wM�YmM�ty��FJS�:�B���(��<�-�l[��^��d���'cW,I���l��ȉ[��Aﲛ�	꒼�#+W��8/hfF�*�Y9Yͣ��ᮇ\t[�|�q�[�Gn��$�0w����Q���gv���z4��T�M�)�ѽb4Z���3�ݫr����g0��p_��
�+t�7��i��<��{7)d�ji��7�=q8���~J�/sY�d��\��g%��I�]���5u�h�
3-E��vL��cc�h@O��(��}4�*��GU�g'J�T�£q��tH�<�h~@��u�,g�^^���jV[q^{��l�.��E�Qe1v~m����`�y�s�h«f�]5�P͒���1O���O����O�ԝת���@�e0���x�H0ܶJXh%E���Uv'��9%�����,�FW1�P���<ؖ�����1��B��~�D�� ����:�?��)L�y���	�n����q�;�6�L�.O�����
A{�����B����lb⨽�R���5���1.��c�8&�[Λ$(
���r8�aޘ�� ������~r����bJ�W���p�z�kz���nЎd����h67�5^��@!'�*�����^�'�$~_&�uAW���Җ'��aH9�H�h�H(A.�+�ʱ#@ׇ�g.>��j�C���&Mx�X���a�t�UEi�0��t~s����LM�J
E���l��ѿ��w����.��s���y<�)V,[j� �mi��T����L]:��`���]�~�����9,�h�e�=�st���r:84IЁF�� �ջɉ�2ԧ\ϟ�]DQ�����B�;V�x<W�w�kE���&Ø{���%{�s}�g��M���Ϸ:VBe����IGX�^l9* <��p䦨��9���g��Vxw�W�+o}|5!��9$%�v=�~�"��j�\#�<��t4_�H��1���B��f�����WM�] ���N���p���a�Xw�9.��	i(��`�do�_u�&b|��''>�Z|���(���
8a5��� �Z�����,���Hf՟�԰H8]�şw�(֗�a1h�;tm:��9�s�D��o����(��pw�rݽ�0���E���o�:�#�y��?��5b���s?IDrz�غ!�{����+�%��1{j�3O�>�Q.�Rg�&�$�QtG����u-Ҳ�+*X}��骝�7y�����V�"
{qa^�9"�; �d��l�f��o����6�n�D������EH&��q|A��a�К8�h���[w��iS����л1}��O�l���Y򂛭�;���,�0$#��.�w�>_��kh4��
�GC��ӦE�p�q�0�X�^�S���(��P�W;�a���jz��4R���X(>]n3kv��%��8T=.\���5w�B���lI��rU�VY��A9� c�%�\�2p��(W6����l�H����s�����=/�9�MKn�/T"��h+�|X%��@�����C�Ւ��8 ��p�u��v��j�K�6����;�҄׫7򽍯���-}{'ے��`�������\�~�x�q��x?�֗ǰ�l:��`�y����'V�o�Ur���s}�2����;f!����~-@�l��6/A%"}�6����h3�۩�M���I����=}�����>)�(��Bp��n����I�Ư������k�T�[���)�-
v�B��5]�寎׍�mE2_qp�]��l�5JЎ%���|M�UM #���ǲ���v�H���P��-��{�5����;/�-�La�f�:4���f�&dtB�������/�D��3����� L|e���a���.|6��%(o� $(vƉ�;�<D�2�%9�i��w������a�<k�@:��^T��n�!]��+ڕ��� �d�����2�'1:8f�J'��~$�$`6kĒn�.܁`�2� �%
*!��Ŏ)Do�����[I�a#zc���9�W�q���	9��k_��M9���H�o��4��d`W�^UCS
 N۳�����[��n��n�5�_�MJ�@�:&k����n�؜�>���_�U�b=��y�6��i�&N��]Lr?�G��ҬB�s(�Kc��b��n�^֢���4;��w�Dɓ��1��~���M ��#Z��\Wz�=`.-�< �ڹ�U���{�3��2�&.�[����y.]�"�6M���ʂeuߝ��+��F�W�`���+��z�8��
�W ]k��"������� ��j<lm� �a��~ mz>���&S��ʜ��_�hgpXIԹCe*nv�%��X	;L�	����8h�p|麊n����% Qa�x�~%b��� �r06ˠ����gA�j2E�0�b�o���>��Fx� �K6^�Kj}�g��  ����%pk������(t"3WrE��8"���w��v$��Î}�xE (��(F��F��.���Q+nm菑ss�\�r� �r�1�*�ڰSYC�?���I�uv)�������|�o8=O�[-���~��L1_��%M��{3j�Y�H䘦��ڋ�>g�o\!zk��s'��RB�2k;`�(VF�Iޓ�1��~BFGW���_�e����L����X�=";����IDk#^t ����;_��M��o�Y�	�:K]刑�D����gmm5_-ҟҾŧQNY�Qb�ޖۤ�G@0�_����SpiA�1���0h&��N�N@*�Y��-���������R��'���phӃ��L��0 ���%��������
7�y�M𤢸�+�VZ�l]&,8�٠6�Ԗ��֣&sg����围���k9.�;W�*^?����z�����[�trU�t,�36�l̏ߡ2�dGGÔ�*1B`]�^���P���e�]����jPu�F\8�G������3�b��l�5�w|�d�YO0MP�;��x���#ꖰB$��2��u;�"&�rZ�+�/:y�LA=���6��mYe��~�vj����ϓr��z%x��"�;�(�8��������x�g��<����DA\������\�[mX���G�"��,29�8�j@�:oC��ț�y���/Z^6S1
�©�礰o	�c�0��)��{E�ύ3c,8�'6��U<�,K=�O1��܃V�I%�}��yX�O��qj@�	��1�' I.�@{�G�J��S�0�s"st�L���WED�UM{F� Gh"�"��<�>�WϦ��(~m�ʑ�nR:�"k3�
�o��f���c�u��`ŵ�Y��e,{t,2���]Q���e�n����̏6���oJ���1G�n�%�uK���<ї4&�b��
�Ңl_CK��@�>�D /��E��v##�
�.'@���C�_x�d��lWfR�k][�����;!�\J��(3��x�ë�ƼHFX�3k�� �s%vK�TGQ���)��h��ŗ1 �ikNFq��8V���8����iT�%/==����߰(+����Lc��s��f7M/k�K�'9j<��>G��Q[b��P�}�;0X�m�EG�Vߘ�0��*|���ސ��$7��xǡA��F�{G����T>��j. �7��d�t
7Ӻ�@{�f���@�
��䴳q�u��}�k���|� � �wF�]�����\�#M?m<P�t�0Ꙥ��z8��380�}���_X��������2Z�t7��L8�ڧH��CG�z��0E�h��ԍ'4+�h�.�<��T�7˰[�g`��|����o�-�ź�]���f=�M��w1�a3R�d(�u1rK?Z�gU{�A8��p����!�4�9���p'�]J�b6
Ѣv�4T������N��A��):]d�q�q�3@+r	`8�s�Q}9��[9��^@�����f!)K�ʵ6���v�D�N`�0�v��s�3,sUå���2��A6�9K��L��ðL�"Ԍ��Ǳ%��@B��[�����Θui��to�*<v�4��?:��T�B.�08`�6+�sꨠ��'�`��E�:�`�6��i������H�+>a?�yaO���	���J���X@�$�c���� ��ힴhC�B V�㎣�������5�_�w'�V�������=�x�p9��x�A���J�&�yc�b�k�܏��'G�XqZ���-I*��E�%UVPsk�W�P��:{������@�̦�'�
nz����3R5���:�cAbB�F��[��h����6 ^۞r�#���90�,{QɃ?m�k�_ �a�Ȯh��rD���z�v�ս٤.-/�(�!1�˞D�-]\���mx�Hf� \���ݭ>�/�5lv�H 7r:�6���� ���@FY��MЊ�}Z��	�D�{��T�U����T��uhD
ű�! ���J�gmB�-qI5�I ]��-A�B�tY��l6���s���*@�fh:9��k��&(~�aO_��h�h��y{*�j�%s�͢#��qL	�y{\*G��D��@�
�ʜ�^ ,5���
a�	�")X�����Sy�����C�Yfh� |�[}A�����0�5+���Q��;�1��)����3\1�r�ǻ���5�XZi{���vQ���v���Sb��	a�m[��wh�&W���9�������=��D�݀+BC�c��%;����`�������9v$�3�r��;�
�UBu��:�=&�F������H[�lx������9� �E�I�*�Fh�W�X���oCωM����! ��9�?�:�lu];������r�emzd<5w��R˕�螇zA�C0�b$��lg���4��_�d<8�Ԍ"67���nۜ�y�xV/G��kǬH������t"��L�1��L2""����:�p&䃣7��l�9���EگfQˬZ2�#�osIP���"Yb��C58�)�*��K�2<
��bS���$����y�\S���02�Z>�Ѽqi��~l#(���I���f`���S��DԪ:�����	��TR�T0�^5�N�*q�-:R�ֺz�����,��3��y�S��t�UKy(ϛ$ �-�h�)���M���؞�M|�[�C�/l����b��S�r��0v6��e���x O�5|��#5h��U���uAj+RHa�&a�E��?w��g�P
)jqk�:@�V�a4�-��h���j��__���ޞA��b�o�YNJuR��p�&����&x�,���
?��!_p�)q[���Cg��}�B��kO= a�I�s�e>H�K;.Ӂ<��O�R@�ǳn��;���4u$��p
�d��)���@�gd$�`���f%9�%�k!9QL�5C�{Jφ�2)g�J�G�����ui�BZ�#�2�y�S��`�==!WA��O��p�Jv�Q���
�������qV%��p-^a�$(���p���D�(�L�&
�`ӖJ�?�10
H��ܠ��W%��	����=��=�����^�*����;���<t�cWyFP�ط��u�t>��Z�+m2>r�vO`���*��T�� `��&2���'5cǌ�>�n��~Y��G�h��y�؂�o�������A�E�-�,���H��9CȪ"8��6�W+��^-LI4�>���5�d7�i� �c@��*��aAhKWj$����.�ܕ��b�v}-@pss�%�;��	��f��yI�,^D�&�T�� �"��Fi���/�u�_�|��H�+)��k/$�A�?g0�7�+��Ճ��]YmE���Y��a�]���A2�)y���r��Fd�v�?���)q�zIW���=�h�7�i%����Rحd�_q�������p�D4�e�E|������
�HZ��`��� {v�>@!D��o>���m�$u'>�
��F�+`8�0?��v�8�$�h�����İ��,L�뾢 }2Xqzˎ^P�mC��f:�:hNS1ͅ1|��y��A�!����yҰ�S��0d����ym�@ 0�n����/��v�����j�	�T�'S`�'�u�.I�)f��]��d�L��pQ;�������W���TS�������9mVfOu6{n�a����@n�1��5���67N�t�+�X�)J�����ٕD,;���)	S6zJ􂥘a=]��a��*{����(m��n%o�n"��p�_;���	�_�ߖ�	���ɦ�����[��bGER�2�� �HJ� ~��F[+�xo&���|��xQ-w����_�m��C�?����i��} bV��7f����N�R�|�?DRܵX���#t�c.�X��l�Ԏ�p���me�pr�P��'����?�Ӑ������+�]����t��L�R��1ۅ�R<ITB>���͛�����J���W;q��\MS+�|oā����ʽ�r��*�;ɘ�	��.)0`���N�� i���5_�BScS�:E/�!�I\F"��
�!�� �vjpwj�<x�i�F�d��-ݓ:�oJ��ۛ�}���v&���tC'������bw���z��>���8�q�q�#�nEf�;�;�=[���$�TQ�Z�P�^(���u
�e�����=~�(���g�ܮ(����<T�}��&�L���z��M}��){�R.b}_q��I�0
B5}dt�٩�	�N�9����6T?��\K�4���3~��F�4[�
߉��\e8��H���
�[QK&R�đ��%�2��"9���@��
���^Ap�O���U�������zP�P�j���URhm��Z&(B�RZVK�g���-.n���i%���B�[b�*{Uv�Qō�X�̿;Qt�m~�.���|���zU��ɀ\��%�X0xa7�� �A2������JXM��T�ٓ�9fD`�D'7@�q����q�e���=���z��է�R ����k�(Á�I��������O**p�N�0�g����c͊}�Ե�P&������E%K�(w�V�c;)4{h~G�Z�8̊���ْE������bj����e��u���V��+ó�-/�5\�4�L�/|��W��#��=Y[��N�]^�Lv.����;|���R���j]7,!���9k���F�x#A�4�θg�5R���L[����%L�gA����݂M������b@�9�v�fa��)�N+�X��Zňƨ�|��8~@� VJ�爬KI�<|�K�J�p�|��LdzT谧b>��-b�_�\�h��-R��'��>�s��ƃa�f/fj���l�Xq.�<_��;k�Ʒk¦�6�"��>�Ԕ�W6:%��9����zs�eg��}���.1/�NؿL=^K#� �ͩ �=���k�D�-�B�K�'6B������0�������b䟕�&� h^�D�Ӆ�wt�%� 3����m�C�ՃMb�i?��0�m�{>{J�lV�L�RK�G�zU��_ˌֶ�j��\�	"*��胮�^׷Գo{��~Q��ٟ_��V!�N�u�zE@$?��q�>)¸�
3|��lMԢY=g2���*�X��`����^�۪���;���}�pģ���` D @�觸c$�͔d����y"�Ʋ���P�՞���@�Q-�)�IMq�����}6/m�5GN�ɫ�4he�FL��4$��E�y��}%�^ܫE
���'N�'1<:�G*&�AH��r/5q懭2e'{ΰ��%V������ﶳnm�|��\7��3��_�#=u�����+y�*��;�{�m`hAwd�+�͡,��������9�/ѹ�HŻ#F��4G�9��k#����."��ά ���'!i]V�U&���6#�T�΍5;Y���#���,$��E4��=����:�b�r#�ͯıD�7����@/�`EJ͡{�:�6���J�γ˵��P����I�QJ���i�N��ߒ��Ws��Wa���r0.�j�V���j'\�r�-g]!������$n�}fg���-��L�D�����c�lR�PX�Y�	?�t.�������ԡ2�!��2�����XDxl����/]n��{@��Ņ��m��6�忧V���w����2H�>B���(3�*����g��
�}b�0f�ѽ��KP�����j�˩�c!���Ȣ�B��Xc����n���:�� �5��9@�hؽ"X���-.�]C?~�f�R�U��~x����L�p�N�Ǎ�#�^�<G䭗A�o^pb)t��Kc��G��t��T�k�i�Mf����R&
Jm��u�0������L�AX��c��m�[�U��v�#�����azR���~eA-*��������CTwl���jQ� P��<`+��O���YV�9f �����'��yw'��d�
*'�ؔ4�Me wF5pxXr#؅��@&����G�j/�ލ����&�	�Z���!��*x������w�֨�E傎�~
ۯT�PO���+@�\���\�98Oj�e�������p�.�z�|
sO�<�{�$Fŗ~�ZmQND9�D�r���/S��g�a�� ���V.2�g2B�*�j�����u�w
��-�K�rp񙸫�|�$�����<�޽n����� 	�~Bk{mG ���RA�;$G��6i;{D4K� _��RU n�E��ĹnD��Ȝ#�ٿʁu�6�߸�܍���z�V,�R+&(;N���{��+f	����W+1Z��¨U����7+�7�y���it�]�3�1~Ŵ#K=�)`J%�[N��|�����@!�:�R�?�-~�N[�n����??�a�	MXn��A�}#����=��Be�X�I��H�5�-�͎�)P%w�zq�c�d����ڡT�{(Q��UL�W� �S���6��K�拋ZE��}��C@��海!]T��oD(�B�s +�&��"�Y%A��S?8C��>��~	b�;kͭ����	ŧ��A�{�ܿ���S��v�H���8Rz��!1��kεg�l��&^6��D#��ۇm�3��qP�	m'��l+d��.߷�R�-�?uy:΃�,��jV�ࣸ���U*K�I
���V󤴴��YM;^�#\�K;Y`�h/�D�ʵf���o7�(Z~���*~2n��G"�;J��r
R�Ĵ��4>F	��_��/���k�b�"�IH#cܢB��o�'�8��н��0C�c'S3�8H���n�(C89l�&�j��;�1�oTQC6�ȧlJ�����\,E	j4!���+%d�.��ʓ����k
4�8�on��II�8w�2E&�l���.�r<��C��D ���j�K���)��[$Z���+U��-,����B�5���B?Na�T���[��m�w���O4�ֹ���x����i&�
`�e���縁��-�&�nT�"��d�7��֮*�H��Cb����3�}Y��dD�,Qg �8��D�ć�i�X����0���\��bZ;����#p`�Ǿ�Z���)ZǓf����o�
����[�h�0A*�Y#x鿴�~Q��b�9e�E��x�q�3v;�,M��M�@W|��������P��i�Jլ�pto
?���,/Lp��#3�r��H�m��3�0�b�誅����er�A��\�j���HDE�,\O`����^Q)���U6ؗzh��+0���� l`U��\n>QꞜ��ؙ� f!	�wF�u\��se�O;)���Xe���
�O��f�rd^��J�~U��Y�O���?�X��
��mJ)h�E"3�)��$(Lw��"�S�O�"�B��A��`Bzl:��상�(��k�jp���zf}��@�G9C��f�߻�ͮ�iH0֝�=XܪY�+���gNGu9�[�w�O7+�hOb�!�m\���2 �6�&�%=�N�<����b
�`���
M�@���ĝ����A� �/ي�y��ӆ��;���TI05���J�1���*�3��gU��ͳ�O^c�n<g�1�@�c;�$q�r[�[id�$�[���R��|�AY�vpE5zւ�!�����e4�ܐ��YỊ��?�2�w�2��U�՗�ٹ#,�y�҃��A
��6�OX���gZ��/
X�����h���u�x�gQ�At�&���Ԑ+�#y�E�h1�޸��[��K7��ˎ{]�f8��Ǉl�I(]���eQ�������ĴW�I�IL����g��k�`b�	|엂�a�/����N �b{Ii����3N{��&�+�����%�5����IC���%!�:r�:���l��U"۵̫	�\�"dx�@�E�*��kƩ��1I�8Q�����o�6F ��r�� �/z��0ӧ?����O����l�s�\f��,�#1�M�s�"5χ�h8����LDj��'P�r�,J~�����TO�wZ�n�6��xM,�#$��Bq!�.�x:�惄�����9�f\N8$$�GK�Zqi@I,��������J��	-����KG����""q�������������.?8�;��M��Q'}�@Á6H
�#��H�����g"��X�(H	�G��#�à5��a��˭t���5
���
��1�0�������n��(l&�?f��o`Q, ��P��ԕY���{4`��z���)�M�e7
��^� ;qi}����z7�+�>\�V����)Eկ8n��`�&H���'�V{�0C�^�%���ҒZ}�2�"[x�3�Fgg�"�%�Zw&+�K Љ�m��a�Y����?�w��Z|�Ԡ�%�K�kN��nw�������&MoΫ�(/Ac�p�������zb�3X����
�?�\�Rj_ǲO[DKxA.�"���!�8�w���tx0P��/�@[�M&�$sϡ�k�7:���M|ݦu��x�xx��X�s$Q+�y��~8�p7�N��*I��H�Mc�!���%y2j���j�l<�:)�ȷ�AN�����'n9f0Wy��p��ѿ�v� sķ���{����"���L@@7S'���_v}�g��ɭ��Mϱ%߹�/�����^�m��Tj ΅օ�W �*���w ��%-�XeNI|�|;8Z\�F�A�uD�Q���zm@��~��������渡�v��vN^�ŝ�X��]����z�"��<�ty��G#?�L�W	i�[��2D�nB�U��V�h�~��_�ѡ�������Gȸf!���#��,���A�"��.���R�8@��w6�D�O�֏I��i�L���Zz'��S@�H�� ʂ犰a���QYێ�k���ص���'&xP�3J"���09���	+	>zČ���{kϙ���r~���P>�����8]�g��3G�#E���b���z��k�<J��?��F�NEe/���GN��T�Qtc]��~`G���w�V'���@���*��je��]9p�=+_R�N �Y��>@~j��Z̾dF1O�gቬjW�2$!��l	�6z�/�ӕjQ�_�JS�-,e��sqe�*�AcaS�кf��-%p�3���������$w�_[?Pg	�,����s�퓸0�A�ѷ����bQb� ����6Z�v7Q4Z�!��_a��J'�5��
�N_W�r�.�W�{��&4�wgG��"�s2Wp���Դ��.�:Dl�� �����Z�垵�_�-k��H��? ���_��b6�jc��~��:$w\9��>���nT�N�>}�$u������i/s�0V�� D���2J���i,�(���E����(9�)s�I��@��eP�F�@�����ƙč^5�bH��ҏ:�2�â����x��j�<��I��i��w�k�sfS�������D�V0;@�!��;�;)�Ց�r��oh�~�ah:�Y������R�P1����^7���9���W]M�S��d5 0�F���@	q`���>�w�q{��K�܂aW�JPG��ҍ�,|&��Y�/�Yj��eT��2���M�(�7;Kقߒm����c�t��i ���U<�xe�y����p'�����<���� �R��'�RC�*]�~�Pso��l��F*�c�33���l�K��}�8!%d�>3�2�Cg}.�v٭�!U��I�z����JlRMsR�M+� O���|�bc�:�iQ��7Uչ�՚�{ #��9����;�T]��/\W�+�>!�����(���&)�m>�mulF;*2�'��2ή�%?�%+��VTr��_[.�}�`1E�;`^PHU�<�h�x���i!�.w�Y�o[7خ_�ޭ`�{/�#T�,h���2rí�J��]�=�CS�������R�%V��q,m<�yf���F@�yQ�tEGJy�8cv ���8�J������:,l�О�#��ֿ�1Ua����s0�m�ZL�y�-m��1���6N�*���u�"N3���ᢑ�,]q-�>�xL�� r�R��$81_3��zޟb#D�5����f۱����B;�c���L���Oi��/��e 6��q8�jk����#)hN����I+:�?�9�u�I��x�=f�TԦ�)��m�#��ޘ��E�ٖU<���I��q�ç���`����P`�k$
2�B��X�na<1�����X�[3����j�����(�l�^ht����l_
_О�@��-�Q�HZ8��� ^��]�gʅ���:e�:�Zmm�6�gbl])>���f��n��S/X�)��m2rb�5�秝.)m����&���䶞ahA4]S3	/p��%�0'��n\M�T�p']�����\�u��X�V�]fw=�����Pb*E�^����؉���h��	���DfVz+���]�Y����������>�-Z��U���ZP+�P@\E��bޯQ6<�?��7�I���k����LDJ�|�@�`N; �Tp}tJ�L��P}j�_�bd#8:
�1�)fͣ~��ζ�9��{B-�`m��<��۽�K��7!�1�4��Ц1��O�+���3���ae�I��M�셽[hM/�P��KM}��ˋȎ�jA����<v��L� �&ژ�8����C���ᒓ���XVĝd���]	E?�_��N?�Q*��Yu�����;1��I��<`m�������+Z�
b��L- �9��D��țçL�D�yc���(u�O�U3�^{���}��R����^̫�*VA��0�0S�J��W�L���vMJ@%�b^�%�W4Q�7���d���ͨ���<���j����	\�(��NK�%�������[�?#:{�V��5���gdW�Lx��6��4p%���N��2�92�gȴi�͐͵����C��#�,��9a��tF�|�I�^<j������y.�fz��f��?���r�Z�zj���{�Cd�Cj)\j��fנ��'�0}�����"qC���M���a�����tXW�O���E�l%�=#��mʷ�qbi�z����$b�Y���m=tO�2H�--e/��A碠w�ߤr���� ZǞ���7�(��(�×c--�U>zˠkÛ:��ZR�E�|R�c���J��������M>���u\Z��׾��/�v��v�j�����Ee��FQ�Պ��<��O/��(�ڽ�mD�>m� k2b+L�T�Ѱߧ*эU*5�pc�������s0��W��^�[[Ol���q7�@ߒMg2��$��M"�Mq<5+�:A�:��Y$NR�e�_^n����V�Ll�Y�3�:�b��,ś���#�5��F&��\�I�~��s����Pq�����
�}&>����)�'�	��yaL,X(���ey#��0��J�ؖ$5풮���- ��Ԃ� ���G��Z����&��c��16j�؂���WG%;Xi���oMi���x�lMO�#�V[����Z@:��_���ldv�.#o�d��I��^y���y�u�}I�f�����<&/\�~T��n��Y�y���T}��G7�u���V�q7��+l��\� �,�H�-�L�8�/@�Y�*uu�k�E��j(IwH5���X�#
zX��]A�TF�l% ;ײ�h�
;qꖇ�8!�-��9�]�D��=�\f���~6�� 
8�|�C�P�qX��qMOd��#����$c��7~&�kw����S�!]c >��d�z�ZD��+���B��y��V��=���;�_8=��>�c
Ǡ�?;"2Z|�=�k)����$R>i�f�nW�V�t���o
6��8�I�Y6�_���?�DY����J��y.I�B�Jw��H{���QC�Cfw��j���+G����R�L��$�8����HXK\�?��BH������jPe�6Gc�
gC"� W_��3v����?�AD| ���y�e��&I헠�ORP���#���0��GyG�8������V�Pt1�[�l��eA��R�����e�I�k�W3�q_{��/U�bE��Ȧt�)�� ۛ����6:7��[�V�C�/�����K��;D����#0B|��&�"�N7�dmp5���yR
��������b��uG����ȋ���m��*�ܺ�P��S���}EvS��o���X�7�l?� c4$y�p�����3��$K�����(�Y]�3��נ�&�؆���p�S�ӁGq}i{q��6�weV��ړ�V6Q��!W7c�	��bP���2f̙����+�W�:�t��O-�w�v^�:%���V&�Et���±�9�g�trɛ���@�:]�u�8[Sz����n�ظj��T�#����aU��̕�M7j��Ǘ�M K �.�[�I�ѵ�k>s7�H������K�~J�����m�W&�˴!#"��7-�w�e��q��z�f^O]�/��p�5�� h�w in�̛au�L�t� ��.Y��E�?���d�U��y���4�A$����+���a�3�6�<m�"b��������B�aL_/�=.��/�7��	u�%̥�\�i�n�]qL�T�6�pP��%�5���P1?�:�	�T�@�]U���cGzف�6����{�|{�k�P��߿�j>���|jy-�}&<�: �քs\+�a�.���\���Bmd��^���q*|����mV��'��̿[�9݊�����R��de�40��t���=2�Ud����RIM����A���)a�.�A%_��_�i�>|�q����ێ����%��9�7����אʦ����o�T����ž�D�t���ySi����EҐi�����##j�]��2C�]ݞS<��e=�F�C]�Q��B���X�B_0���l]�����:�ڳ�t+�'냽�h5�4��sHY�)��'��3�����Y�3p��r��\Rg�Y��l����Xr���ڑ��"��
m׹Xe�Hu�4 �z�x'�!��$��6u�z�<x�5�eE ��a��kϡ�a� �ʩ_��"�94���]O_��4�,rU�bPݵv�e<�L�]�*�^�����!�q��uU�.(��pbH�3�)~S͝ҥ��x�IP	�����A�!��V2!��$��q��U(+����G������￼M���r9�LEU=}P�D�b��v$�������|)��s�y֛��VN�T�,4���{R�0�h�xr���,�k��&���<�ݔ�#�@��տ\$Y�>�S��Qv����P9US���c4�n�Փ#���k:��/�CS��=���`agj!$�/P?��C���1Teʰ�q��;G3�U������T��)�����~��I���P���5��?��D����oU��{�����h����Ƀtz���R��>���㰅fs�
��+����W�L�bJ�23��Z��Em�Kk�F�rA+,+A�4�����*P9k$��qF��C�(!vm�|�Z��-W����h��uC�HȒ��]�(Sڿ��L��ޭ�M
�4xHC3�m᭑ٸ)z�S9�`rS�/
_��FEm�{�v�k�#;�F������u����(ZŭXOv��[,.�wրA�1 re�4F��\h�!f'h������G?f>&�P7ΝX� 0��a �r⢼�����i�xI�,�:[i)�,!���pf!��9���9e����E[y�,���=OY����󂈩nO�����'0�X��`��S?���E���Z��y�׳n�U,.��5I�Qj9A�'sEuT+OZ�-��r���F�M��WW�և�t-8���)�l�v�1��*c��(�w2=H�����x? �%{';�ů���-j\N�YM~�J�	�f���NB�;�U	&����7��F����R���1D(Ce֏�=�[�=��1�������oTf�jiz\$by�[@��]:\U��~_W���*�aPאK�S���MGOTbY��Ԡ� ���J�jgt�������Iʔ�������F��ю�P�sI���� �
�����/ߙ��k�cX����F#Az�C���L��*�]b���M�)�ۛ-���˨{B>s6!����_\Mʟ���]q�a��u\�� 5����3��d��c�_M���^Fo���֫�O	mM�!�B'=o�%6�Eҭ�������v�K��z|�	���@hK�J�5�G���qMQa��+�e<'�dO&Ͻ��X��ݳ/��S�?R��\#�7�pi�[H.�)�׼�G��!�c7{:v{�"�oг�6��t��WԘ��m��RKt��4oʯU�f����������K��}�,�p�����n�_��d��cEE���9�(ED� �-V오m�	���-tg���C��r;���F�k���=��&�xT���=X���,�O�����ʮ]�V�
��`�X|���6D���H�hV�$�a���.+c�3�!��(g	y����Z��]qbN�x�}¹=�4�e%"}Ee㩔+��=�e�#�� ���G_����{�B(�V5�U��W���#��	��Y���Nf94nhr	�g1���k7����Z�;^��|��9�������ՌL%Ǽ��x���i&P؇��b1�|b� �=�L$�X@Y?\��b��@���{q��c���L�w��,aU�DDL2z��:��6C2�kN��e:��tϡ��G�r�́ȊLj�����10ص2���ꇫ#��Z�C,3U�Mi����kN���,�%�k�d'𬗺������B�aT~�߈U�iJ{Ϡ��<X�M?��[)�� I��V&�.B18e���һe���)�h��=w�a��+\��s�}�QɌ�!q/򣉊�Ů�#Z��a
D�Қ?�jڱ�14�r��(fuI����R��Ȃh�4���pMD9��@RѹR��<LI�M���h����IͰi�a?
o�ސE�!��&�Ϸ�?I��ɦ	�1��d��������ە��V���;W����|t���o�d��e���V{���^��f��&�'�w���U��7h�A�j=)y~>�T��t��)N=�P�XG�6H��f��y�S&�V��H�6���Ã61��G���H�F��h�21�n�Ā��Xr
D��U�3MK�wJvo�S��{� ������S=ڈA���ʢ�z��H=Z-�:��ձ�KU7e3�O���{�TuB�4uyܚ������D�I��&��v�t&����2�b������a�4G�qD5ȶCWRX�3ޚ<�����#���d��� �r�pO�K(��K�:�:�����^�qIf?��L�TQ3����qU���AS�n��e��Tg�I��t��*�Mo��[Zig΃�$�p�V{�X���*��q7�!��Y�	s"ײ5䅪L<�EB!R�}K#��s~����b6>
�g%?R	�h������b'Y�p`B�4�!��M|Ҟ�����39�E�p8��.;�X;�_���Ȯ�^�������7nIf�r��<�8���G�G�</�dGP�t�i���5�B^|L�	���
��Z��������-��=aj���qW�� 5�[�i�i��C�R]�{��q썐b���������;�z�iC�����+�V3%��j ���)��U϶��O�a7�7�b��.޲���,�5sR�i\��E����wޯV��o�/��?�I+0���7j3/�pS:މBv�H6��ގum�
ƌ��8��>�z�Sq�P�f,�b�5ZF|�8�{98s�̕���6GN�X1Q]ގB�§�����M�+g�ƧQ�Q��[�>��-�9/G��<����g'�A'���o�|��w��C�/���J6� iץ��V��x���ܬ��B&�X�� Lbv����Mɞ'�E�>d��}���Ői ��ޓHB5$Vvs�&+�����%[q�	�ɂ�?�4o.���:���+<R{�I�hA������=��}�!J� ��@���/<o��ʄ�đ�vw|'��)��o
�ٖ ��/��v]H�d� ���H�!��ВF�]Z�Q��9�gv-YzʊÈ븣���9�/Ȗr?z���6�"���bc;7��)(��W���W�����a�W��籷��c�H� ug��ֈ0�"�g��~kV��^O+��BPR2FO��,��{9=�U�&�Z���-Y5Q�.'y��yj�]���*H�1>���v�����_�S�� ��H~�f�AV>&T�gE<l�F�zb,�s�����
S���d�X�Z�h�v��ٷ�B����#	�Abi>��n���ǐ�xA߸���{qz=Ł���3�����S"U��K#l��	M�B��b�k�����e��}v����f)���}!]pL}˛bcv���Y�H������Ҏ�bNsЖ��vzÌƭk��G���c��$�M���+�s]�n��p�@Ä��>�W�I�`����Y%��#d{�Fx�
)q��=�X��ͭ�h}f�|�bn�X��gY��
�ԛ�o�uݰ�v�)�.�H�ݗ�P��zI�im�{�Y�������Iu�,��"l��?�Q'��<yడVr�����;��o�'�����Yw/`f���"�M�Ȉ����=Uv휛��,�+WHt��Lx�� �G|�'�똁���M��0vdy�M�)���K�N��8|8��hJjG�إ�M�S(���t��fBD���b�3x��L3PY���9U=����}H��l's`�߈4.$��~&��03���A/͞�������}���E@�vC�I�4�awS�Ң|⬖?�R@8C秮��|�^�/��3��<�_s%/�ͪ��B�.�����LW{��$֦J()�{(���s`�F��!��%�Xh4{aa��d(������(|�a�_�H������T��Ѥ��� ֖������^^�4��L�)X���J0�B��6Kc�9�+���;s�-��F'�4ײ?�eo2���r��Br0;=6�E�ܦOَn�[#���г��3��*�M�����7���&B��RZ]��m},SҋiL�IO˚�V~�\�%���
&���8e,���1R��́Aj������S'T�	��+В 
}�x�2��CD��(U�����fr�kF��0��+����SX��A�4�w�V�;�CV_�ĐG��O�W
�Կ��UV�e�0t`Ʊ�j�r��γ����_�f��3�Џ�AF��8��I�����Y��n�C�u���F\��\��u҉��қ'ΐ!U�ͱ�Rl��\�$0v�f��uF�����D*7�|ſ��q`�T��<�� 6�nQTĕ�V�	ޕ���4��q�Qo*��k�^Ċc��K)�d�~����$���CaX�NS�9���jy*�sD�b˜�ں�����������6�>6O��5I��nd�l)y��NdG��׵�%��|eD3Q�=�t�E�����N�m:ޛ�|�� ����w��̬�2���}�I����`�0ydJ��4R����Lm�Te�_/M���6��c!���(�h��ݤ�|�{?��Y���z���&�`~lF2ߨ��~eT-�F�[�����;n��Ȯ�B��Sq���?��U��_��Hs)G�Qu������<e%�b�׿��
P���B�1��22���y#�f��W��^�k� �r *{�h�]�e\���m�����Ԣۙ��!R���My�'���c]sK��_�<98>(�s~]s�;�ʘg��tZ���жi�C �"�kV�>��i�(E�ho��Cw��Ϸe��Np��n�Jl�^��bd������% �r�w_��#�Ѡs`�4ڜ�Y 7�fWYُ��Z��m�`�i�d���H�������9�F��f\�O=�@`Jd�sb����KT�4m��d&���ՆE���=(.��Ӎ����՝j�D������Y���C�!Y�
�]-�"�0���]����h��а����Ƈhpqp�;qݎ{�\�����J�3��pڤ�l��;��lކ��a��D@�)m@<.�1�ZĒ�ً
�J9 �:x���L
����V�Ջ�!mȁ�4 ��'��c���˶F��?R|��/�3u17*[H�]q�C��۬v�-I�4R�qU^����e��;�WDa\�vh&�2M:�t�a�h�4�ϑo0�s���w7 �unue�Z�ʲ����k�h\B,>Su�����̞d�?Ǜ1M5l�Dr�9w��5��k�C�9�$�� 1��JC.�z� �w
 �BĎ``:��0��O&��8����C�������t��$<�V�hs`��n�}���6��gp'��a,b��JgD���a��"Z,��SM��n��ネ.	�}4�ʤ��U������
SF|������h�ۭgA�s�^��ħI�[u&��z��M=7U�xX�U�+�t�؏T��1ۿC��� ���$ܻu�~��ey���d^���i꿘is�W�0�Y�)m�U�n%E�2�El�X�>J�E}�Bݱ`�96"��^�Sʈ)�{�ע���V�y,��~�0y¢�RDJ�4ұ�C�	����k����4�_԰�*���g7��x��S!��r����S�t�`�`�t��W��Ad�0!X���B���<-��q��輳'�+�X�6<��37X$YëSl�F�0W��J�ȳ��{q��L-�1����q.���#���bܟ���護�"$F�\F3���va�Z�7��[Zh�l[{4�����N�%3�rh�FL7�h���3�����>��� �o+M� �����LfA�j_�1�P�#���2f��8%6���1�#�Y�_jh���N��/[�:X*�� =��/�i�Sjj8�Ir!�q�� n+�;Ҝ����v.7B*�Z�_ߟ����!�IU`���B�"���Eڙ;�؎���U�T2WHc
Fo�+x,z��^b��Z�<�����������E{����6����:�i��%;�0 �էĺF���3YLF`D��g$#F.wj�_re%0�ڞJMuIj
Xy��xn���`����}��:)�<����ZC���2l�-;:܉!������j� w~M�Iy��9������I@c����%��\�t�=�8��@B}`���V)|�t�C�H���j���%֐�b-mt?@!u�h��4��$# ���:w���{���;����k�붌��Ѭ/j��c��-�hE'�K�.�Ň�|�11���<�"sjQ�	LA|%I�$&� !9l��z�ru!���k5�?�@�{��k�5!|w�5�<{3�_�����ǳ!y�}��	�}��t��O0��PF���[Mg����i��}1���
.�E�h�\ �4��LW3ʹj�58��PmPAŃ��Ҋ�s���D~�I�4G�[Z�J�
�J	�mM�qSns	7>�Q�e@ h���ܑ|O�t}�̡�WW`V���=�T[ �ځ	.��X"���.�u�⊳�X�h[_���YE:�
��4�"l�;��%^g���vݫ�Ā��0���h("���uL"o7������O��Hϸ�Ö�� ���M�Bzk�
��vkb�eVp���Y7�Eqb��nQ\b��W���˷b�2�#��i�O��
��lP�������M�*��w]�B��`�Ɵ?�c���5�	)�Aɰ��s6��'U_�}��0�~�����kf��o�S�G�6��`���Ƽ����:�/�V�WJ��D���i�Pj��*�#eJ�8ƙX��+�50 9��v��僬gY^tFi���ߔY75�������|��w��z���y]��U�g��Ni�g[Qdk��i�L��,�C
�u��[�F��lW���Y��ӌ�ݔ�s?^�e� ��׫�'N��9���ěId�{�ݍ\�K��l}p�;�
��[�^{ʮ��m�,�uA��5y�Z�h�����a�HV:ð�}��@�s&���y!��~�!|�z��a=ʜ_�x�d!���!x?�[T.6��i8>S�T	�5x�������qbB� �i	|��
�)��mY�~��l�������tQ��p�*3d	��jqä1�*#���I�t����W[�؏��ކ]]zz����	D�:$�cA������T�����U��7y�*�}��TJu���{�35�Ϸ��%v*������J)�N��ĺ�]�όں��0��g��G�$b��mkS��,h�Q4[; ��،�������{!��/�OR� �/-��$��pFA�Zeƌ����&%���M���"l���]������x�����l#�p�>�����h��N#
���u��B*�G�q��4���ת�M��j�Z�
v���FU�W!���VHtJMm��	�E�ՔRa+U��tҁ�ьyg4��p
�{J����7v�5��y�S"��oxH|8���Lq��pЫ��K������$%'E�GS1��EA����%�J�1��M=X�+�I�,�(wބ�8�'Hǂ6!�/|.O����y�o^A|ARm֠�v�O��ܮEa�YH��V����[)!�����[��Xa�x�dO�p1P>�ߦ��qq��c�/��n�W:֩s9�?���~s�
��ڏ�����ҋ�-N���Ϻ'��yd1�A�+pR�Я%k��m9U�X�ǖڰ�,��T<�d�&�6&!h!&;;+K7)��2<,'�z��)m����M�S�K�ӣ}��{���B7�g��U�[�[?�c���G����Ge�j.7}0� }MфXB ��{�}q�?Qg!��x$�S�޷��Y�b������"b�j��ɽ���%�%�$�G5u��y8�r��#Y��:b���_@B�)��o>tGn�}=@�|��/Y���d�oO��jf�du�bO�s�H��[�g;V����J���r�� �꟯����^�)p�ӂW�5ݎ�i,��%$�3Xx�9a%�@&���Iek\%�[t��4{��G�FY�����ә�F/A�}r"+����h�a�/��i^�p�r��Nѩ���x{]��+Y��p���45�F���
���\����b�թ�f���?�܏��S�����[�����O*
zr\�e3g5��h"���z?v��PP)~��4�ۑ�(&�}�Z��	�	X��Ύ��w>7�I�g�a\ۯ�!U�'�ǖ��Ҙ"�S1se�����Ξ���1R�HM�O^�����a�q��Bz�ڜ�k	x���Pr	
J;|C�"a� _�a��Ă�'y�B�gy����QsFȇ{����Z��2#�[P���p05F�\������EU�U�����UGl㶖1���Υ��[�<�BV�Ny�H����8���� ǂ/n���3A��8�s������7�:}Э�$�F��������b����zݙ�i�3�NNK�Z�#�I��Ν����1Ո�ӈ<�``fuN!_P)'O�s)P\Ϩ�`̓�D,������եK�c�\5d��>�6���\`V�fR��d���e�`u�F���6�p_��_.��锢��&��h�b*�NJ�2������s�G�{�V��h�T���Y�d�^��Ux���+�G��`x��wSsmVl����Zg.k��Ɗ3a���'�ՁЖ��j��Ƌ�x�7� �4��Ɍ�lǍ���x��~�%7è�8D\dZۀP}��U���������?]��x&�j۽���<b�]��<��E˺��f�3�r��:�0��A�U�|��*�7OU�/�M�j�t������9����^���b."b�MP�W2�#��7���?_3zT�[���3��M(�������\��+�З9o���O�۱�џ	��M���Ö\���\m_�g`����zK�b��D_�}�dr�w<%�f�6��ڻ�cv����%&��1�ÆBY�ڭ����R���X�'u�;�8Ĕ\5�cѨ��������R�*&9�4���u�����>E����2/
���3�9��4��ԓ��Qnro�a����?3k\ݴ�7C����~m�LqQ�)	����A���&�J�^��''qg��&"�rc1R�x9���ۼ��Y�&ϢT8kQ,�?��GJ��X0���&ol,�[O�1���v'm����M�ڵ���r��&`�0������Vd8����@��9VZ�r����iOB�P����R��!`� ^��g�$���(�;"ov�(c!�I�lE�֚�/��Ji���^��n���90�/`�F �E��x" �����M�ٹ���W�N�r,���o��ZI��l�A���G�8�WA?"� �j���Q�uBd����ՁJ:�����V��?��|��HU�������@hi���#U����?͚��v���|�����"Q:��QڤάvB�;7�3��"�7.�����T�=����:�[���Ň��W[�;؜����FF�G7RO�J�l���<�����Tz4�Q^t�np������bq���\d g���������D��#+���Ҫ��8�!/:%�}'�x���[�:��ɤ�&���9�(�IV;䫊�x+�m�z��a�����A����]��+��G(���������[�
l �Ua{؅^�Тe�|�U����Ę ����]�Aib�ѨJ�����3���d�.�T��o��kT�\��!�	^4���z�J2��W��Eq����Q�������\�B��;i?%�HD��K͵Ca��b��9�+8&�!BQVO�s��|�=�|�&m����㹷�J���d��:-3����]�7
��D���h���<�`�I�^��X��u���ɔ}�������x)2"^`�Ϲ���a��4Y{IE�%^��'�!\F��m�G�!rwG���i��s-A�	b<+[�I�v��2��%�Yk���LҌSE�	�ٜxe�h��#�7ރX����@��@-����A� ��;E�=*�'*��k��.]��Hߍ�ɴp<lx Q1@^T
�� ([M�ǌ���ܴ,��V�0�#�9  ��f2��p��ҽ�1�R@7��y+�vF��g=����_��Y{�B���x�[::��f�I�`馮yR��+���,��!�>p�����ϙ��U�9q<�Fr)cR�*��]$�w�@�����qL�b��1G��f�;���YZ�'瀏�^}:[�ҩ�\��v >?��m�'v������S��|Xt�3��ܩ:aW��v����;�,��qlhEo��B}�%����o�o��7�%L��J3*2�G\�������G\����_$81�������Q/x����fVq�md�;����dBO7���=�
	S���i�U4Ўq��^{�:�`[��t����Y��in�EbK2?]�$�&��� oR?�O��]Ua���rg��3������O��Z��ߩ��l�}�uB'2�̔m��\p���j6FF�3�Mu�����G�.�ƩP���B�G#��lu�+�Fc怊0a(�%�לH����*�AxNߑ[2-YA ���>E$=��t�ʵV)6d���� �t�Qv�qz��C�4�/SF�/������xڒ�͞09���*4�K�<��9�^�y��4"��0A�1Z4�Q�B���<������G[�x;��
]�S�]��t�R�����U�o�"�=�]ݴ����`�o�J6<sKu?��i�$�Sm��a�d*$jt����\�D��M��Xt<�Tį1L��N��ǒkB~��km�bK �a��&Hڲ�߫�v.�;+������?mY[Y��b�Q5
2�i^A��cw�X������eeﺯ��Rp�\�&������*��<��U���	���{Q�C�Ȅ�t"�l��@"���Mda�~xbI)��=)�c	uB�Rq�"���rs�d����椥��x"���TC�"�u��0�U��u���tmWt_�,(��]�6tB�:M�i��1^�aa�j6&^�*˕B��%�2˵B��N��Kd�n�IhuY{�@�8�NN���(����{�Q���<i@�2�8�
��0Ǆn(��~N��WiO��t�n�|�"gck-�qvF|[X#Ȫצ~��{'�;��K��G�.�R;���KG�����i�w���zY�`_��]�4P�ך��'1�7˄<���B0���}�N1J���X�˕�ߎ_<���b��^�Q�-����6����h�2/�iL�����BS<�*�I�(!�K��9.�e�4"lq��*�N&BLPT~��_�����T�=�\�9����%AvnL��z��#Yle��[���=N���Gk��F�Eq�S��ɂ�g>1�1:K�=�?����� D�)r���͛��4�!�$ɶ6�����_2�/�n,M�/�g>�]�Y|T�F�\
����,pD
����#9�B-�'��kny����[�WD��&k�r1^]o��O_��XȎ%�@�C6�����x�Cb�t�f����e�s�GbB�GQ��pk^RY���!@JC'�LB|�|�"�8N��S��ryj[粠,�7)z+`��SػvZ�˰��%)���|��a�a�H4�>/���ĺ�"x�-��/2Ȕ�H��:XZ�j�M�Y������Z@�y,��s�?v� �z"F(��u����-�!M_p�z �U7#+�Ѥ�|��X����9	�����H�Ӛ��'oCD��@�됹��6<��U���e���e��ZbJ��e~���:'K�w��V{�~!��S��SBB1ez���R�̾���[?n3ڒy7��Sa����4�~�@�v����Vk�c�_�_�!q��#e�)K`�W���hܰe;L�p��}�ڂ�E2�rh�.[2�\I���)`�s̫��N`CJ�n��$���z�0^��)����Hh��;�,*�"-#���5++c3bE6�*��滏v��%ӑu6DUgw���C��	���w���v��o��$���-��_	!}�>d!�q6UQNő�4"�i']�k���ͼ�n�<b�r�x� kH�z.<����N����.�-��o�B�i~�^=B2h����u�~̍��)��=?���#��Ćj���[�&t��g����oU>�;h>"~�k{E���/�W�J����r�o�رf�\H�!�g\@�$#�4���Q"#���D��Z@@ܦ&��:�H�j��'��r\	lw�
/��VX�p�?��㳫>k.�>_��b�B��S�O����y��+2x\U�����X�7��|��o�8Dk0����pmkP���p�Q{������q���:�^���V�}p����_�����)'���v~��TLkP�{���J<�T!X�F�.��Ԁ�N�ҳ=uY��s�u���� ���r5˝J��\����[�
>��z_v��[�OҬ��J^Q�m^Ot��`�� ��,�W��V��7��V7�ʚ�z�*����
T����/
����(��=�ɤ�x��THh��˨ER8���d��۾�0#��X�Z�3�8	�'��%��#�=��'b*=!U9�P��v����%��u*�W�|�k�;����ؿ��娞[@���{�I4Z>����˻ɵ�n�l'Pj��`0�C�6�I(��O���$���8F���s�9�36��;:!?�I�K���0��kw���!����]٤����7dl�
�Fz>�%b M���Y��*��ϨITkI���<����j�e��.�]��na��z{f�;˧m�z�8-�F�ڄ��4�ӏ�y��Ws ����K�;���Γ����>���(�)�2FAל��:<�Ϧe���<!-��s�����"t�{����|8�D�I�fo!�f���@�7���.�+��\hrqz���w�\iO4Q��{HP�t��b��<I$��f�Ȳao!>:�qR��o�P ��p�W�Ï�Y�/0����v�����]`�V�=�@��k����}�\f�hrx
3�%ح@?�H�:�����d�SD6I���OGж�Tu^З)Dk��c�)B�4<Fțm�F~z�l���f���n����<O���ޚ�IY�7bW�C�Xo���E�ʝ�Rch�����wB��q`�p7�A�����S�UA1ʥ`�x��1�i`yL_�Y!JB�at��t��B[��ze�[�\JԴ8�\����V�99���w�, ~Y���Q��%v�F)<�T���p�19��~lwD�h`c�5�M;�zh�v��n�.���d�`x�yh��s �+*q�Y4��sT!�����/���_<�IO�ae��P���o����Ǟ�ٮZZ�7{����O.,��ң��J�\�Xd?�zQaj�q���~��g>��È�ѣ����f��UFK�j�,~7��lt�w��"Ѳ�X��o�-)����凔���B�E�%Gw�e�_j����M�Qx�o�J�d@�+$���}�}�TjI�k�"�� -D�;8&G愝���]2j5V���!�d��m��~��ʐ	a+k��kv�-�%6�1j��1. ���0e�@�
^ܥ,���~c;t�4��hm[��P%b�C���,t@Vqj�'�h36P���$���lA��*��O�@4eyퟘ��׼�0o��Xa��4u	E|B�0G�7��B�Er<�j𾽿l֯E7�ڡߩ��ǅ���b#���:_u�vc$�>�t��}�g��-�{�U���(�_Mt�^j���b%%<�S��> ��z�I�DZe��F|���2Թ�Xgnf���in
d�C��Ba6��>PHVM�����r�*�Hr����
Ɯ��`5799ޣrQ��#g�kF���-�c;Q;�^,��J��«M�`�u���q:���]ފL�T�& Zm֠S>��Mbe�ޕ��z���MHr�)E-�{�<��^)� ����}�gV.��ewFB5=�)k�H��?�Cw�n�sj��|/2�Y��
Jf'�JI�کG��/ ���o�����v5���N���m����O�2ad�5~ճo�b���ul@9"?i�Ib� a�Ru�Sn���n�.�F�w1&�+��\d����7�D���t�X�%}48�\�"w�2֤��Buv�f;��>����w�A~�$Y��+3I�o ΅;/��t���iuzi^�&y��G}?���;Q��á��"��FG7�hD}�u��D������"n�؃yPb��+��N.b@.�WZ������?V�rZ#�s05�&�����F���J���B=xX1&gѩJQf�T�G6ENV:�,75��UyڇE83���	��u�$�"�{ D���k@�ΕsC}��C���ί��;�g|*�*�w�bC�>��ב���ײӵ�4�g�n�q�rj��X�0����o�
�V1.1��~���WD���{[@��,������@����4����gT;��N��tj,?��j&Y����9�?y���;�FH��/�Q��z���ҷ�Y �� ��Q�玩�m��Dk�S�x1��'�*wy�#�k�BNO�U>�	b�ОE�&�Y !���_��xo�It��}��PsT5P�5��i�o̠vYj��t�-�Q��HB��q�tϕd�:���s�R��V:y�bͯ�2��a��V�~a������S�E��]pM�.��3��S��W�wg���-g�Z�ܚ��^/~�I9}?)p4���w�`��PT.r�q����B���#]�զ�gNk�Dau/��K���ےwL�蒍��
3؊���>��<����1��u�|DE��}��h����yיR�'YYB-<1�Z�Zf�\�GE�U&0<!Y�Q�E��j�X��Ҧ{����dj����7�f�L�܏��-��o5rޘ(��� �s�J�8�l0�����P�b�g}@?���v�Q�wi����C6�3O�+-l x�) ��0}�i��B��-31���%���_i�6���@R��o�V���FQ����c� D�l�G�n �z%yUN�����s����8@�&��D��]�Az.`�3��ec�w����E�����ଠ���2���dRe�1���D�^:�K�K�i�u���Q�<(�'���I{6����mN�~s��ƄC�F�0��	Q
��F]���h���n4���T��e�4�>>���w�r�"��9��ɥ�6)ڽ~)@#y� ��l��*v�{�L�~t�bܙ�`�>�~�w�̱�u���vp�M�^"�|���	Ī�5'��UOL���է�����l4x�b�@ԡC�\�0rC���<i������o;���,��'�E'����M�"��Br����BlR��`*�PIz�Iʋ�ӳ*�x|˃`���n���k����rs�M�.ѿ��F�#XF��M�:�wgn�VS�����`��7���oC���w3Y��J��]���-����l¯�;�!7*zG��������_L0�JMV�PIie�Ț$�s!��0ۆ䥷���Y.��,~t�mɧ$�D�7���*Coڈ?�}Ŋ����j��N.?)�X!��Bd�6&�C�������"�%�f�/��˭�"��C���	��z���W9�*��{�����Z����F��VUFF�Q͠��L��;/^�����^y�6�T*)����.�^@��X֡NI)�R���(6ɵ�b[n͎�V��E2S�u��U]��ڍ(�����33ng|ePi�V��F����p����<��>���!}�t�h�}+����z�j����:��ps�~�	X~)��K��@:�<$T����uFk�������Lq��u��o�Jy����	'��S������-*��~��n�B���Xz k�,#�%:Ac���]E����S��)j]~���0���ωA˶Ccu3%�K��f��f�a!�o�Ѩ���T��!h��O<[��S���h^
M�Ql�R:@�00=�L� }9ȓ�
"I�`�sWMNزDϞ����%��u'|Uղ��lŲ�6߯b���C�Foȳ=�r�7���f|��=Mb5����#��q�f�g�8 ��Zf���yjO	�c����F���R�a831���oVTғ_)❯�qp��m��KR��l)U��L$\��8���L��9	��(��nvK�Mܮ�N�]3��$�{o�R.�z�G�a�1�Nr7��O?������Y�<|蠩~J�P{�m}'Ey�15�f��E"=z��-��P�
�8򛚃I�����/�!�o/�Mr3���)KK IJ붳|-�;<ꌼ��"ti�L��������l�$�H�� ȑIĎ�=h?e`�}X�5���x�ݩPR�̦��!�yY�1����t�>�ԡq��o4��6���L_0��r��`x;�X��>���~�k@"EQOїݾ�W��Q"�� �SvT��)�.���v�[��_��E�u��o՜�o,�e
����%�ׄ�D���M��_^��N.�B9��`1���W�S�{s�'d�<��S[PW�iPT]����h+wR;�ۿ�N����Z���cfF; 
8-A� �C�I)�Pi��h|��ݳ�_E�/��zz�i��|�����^8��izO��=�72Z]u�&HNT)�i?���)E���7�Ŭ)N�w�]��%�y�;�:�\�z�?�����e�e�A�j��M�B��Q�莤f��s^˅&bW�H[t�2��|{8@9��o��}�e��aVHNs����}��vI��t!)����}�t/����~�4o�{���҆�t4������4A�E�y��m}Q���hR8B��DS�sYz1�y���U��ݤ��� �uQ6��h8�+a�Kz�'�i6��i�Yv��Yt0t�cQ�P�����n�_���3�&Y틴�07p�Зrǟ���XR�ҖQ�'Հ��R�N*c��V������P��<� �!�j�k�!�R=�0A�	��Cm痼��� ���
��(�m��Y��h^�@f�Dy
~,����5חxKG<���������eڹ�X*	R�B�����4b7�z��+
��f�TC�ֽH��t9���s�����cwS�@�t'����h�YјK~2�Yg "��Y�Ui@�[�G���Y��:���b�~A�r�s1VO�xF�(i��`�����.ىs���  aU�����y�� b���L�W7�L��m6�������!m6�Ô<�j�����Ì�Ã�[s'!���E^��?�V��&��N_���� ��j�#T��F���NH��R:jR
�*����~�  '�����@}�Mm��5����xa��p��ɰ��{�
l"�M���z�ߔ��S�~���Ss��M��".�L��f؉��On�#^b���(����Uw �W�at����3t�V/o�-���2n�^�޴��_���#��w��	���2��k�fN�y���R��ax����Y��`�vH�ur�Ke��.3�(aA�]A��4hXjdA-Ӗ�`��6�;�:	>�$	������� ��݃)�{h���3A�D)> ��#A�����?K�O���")El�)V��l��tw4_���s9�������͌�$|�� �H1�)9η^�/�.+)g�q�b�Fy���y��s��L����cl|i�ҷj�ܙ��*Z`��פ�^U�k��6Ў�ZY:+���DW��VY"��j�'i����")���x6'����,l���ڗʭ,ro+�Sʂ=����54k�c��G����[Ehq��鶜����ca�-7���(�T�K�L!���v���pP�t�R��m�OQY
 d2JLȤ�`�ǧ!���γ�9�L`�K����(4�>c��=�i��K*����mv�=���p�6�V�C<ar��_�1�چ��z2��*�gɁR:��n4V�^5�%4��X�B7N�����	+,"˝�5�!�:u�Q^�����퐡J$���!̀w����vD�G�ܯo�u��М.��dǦ�R��#�̎6������|zB!�'<�)�����J��(�?R��+��0)��y����z��ɥ#�NL�L��)r��:b�D&�9��s�hC��C?��ӵ,&��'�;IϧA>�NĨd!���!W*�EgO�"ҩC&�|������[X�oo�)1u�(���"g[63��3�"��sJ~9!Q}k�φ^9��j��%uQx�b���/��7A�����C/YUպ��_�x���|��\2��G�����p{�PK3~s����&d��v��i��L�K��%�O�L���[���y�b,Ѧm�So:w( %Tژ,m[S���	�3�+�fyבz��	��c+A�6n���L��Y
2�̽Ui_�.b\	��D:�m�L��Y���p�ESo��j2	w��:�ke����� �GW�g�m�`�!Y��i�f�G�%��ݳ���tDFΗ�즏�Wmfs�M.��x��j�>����>n�|�Q�g`#9s��M�O^�b�R$�>�\5��5�������hR}-M��S`z�w֝��{"��jj�����%g��.�������������g���_�_?�Y�=�Y9��9��pZ���0ȁk��s����VRs���2��&�K�v'h] ��҂ر�����0���e� �0��M�I��:�̼����4��{�Z�{���4�O��l��Eh`��6����M,��`�!�t����(�M_A���C�ܝ���-���%��p�sЉ;��N�h5�MU���c�D!��|5��!�c�Cn#�T�]�)�-0W �H7��]F|��}�%($JtD��P�.�ld�.Ħ_��IK����5ӵ=���c�k+���W�c�X�K�?����l��,Ký��4|0k�B>�\�y�1������M��7j����Q] ��Z�aԌA�?{J�4�����(�4=�+xu�y��m[��[׀��v��l3R���vq�X��*�'���$����� &b}V�A<j�U��
�9�� ����tM��N٢���M�f�o|	� o�!��Nw��rh6����z�䀃}���ݍ�๛+��^%�ﭶOj�be��B4�����P�^�|��n�S�����/�� yf��k:<���Qz��^�M���?�B�cD�b�����e�`�T�(����9d>z�x����0c��sU�}T�pλj���Y[m��D6����o8����D%��`��?�{@��~�䋽Ù���c&��o��LU�}%謧��}�����Hv��Q"��~�y�gxT��>�V2".�
f�P=q��%S�|�"�©V�2���o
��Q�64��A	�q�<@qkd�9QM� ]Feզ/�-��)���,�_�D�7��jU�⍐�K��  ���N����z�_���E'�Ob4p"2ɚ� �Z4���P"(���@\G�
І��JHW�&@�HыG��,(�b�@�&��l�}A��WZ�2�����1��^����ȡx9�����-��y�?q�1�7�`͐y^)(�y��fg��&K@��k`@���8�=:_�B�f�ާ���!�!��n0�^�*������&�t�v� b��w�8�m��:�7���PB]����:��e�\y�D���MnQ#n��u�˔8Ƨ���\[�*���ڗ�[�ҁ�H1[t;�@\�4�w���ܥ!�0}��W�kk�I<_��ȾU9E�n)L�;�h�����c�3�ޡ�X������&Kc�?�dx�D9=�0�*Ϳ{iFJ8�|�����;�?e�B ̒�Q�h���LW��
�:��Fk����z-0x���svV�e��AQ���V�J�����@>�B�L��]a��Y��B�k�q"�o� ���F\S|g���ER���e�]
�ܚ�v���Y0N9/zS�i\���.���Vt��Vf83qy ŝ���Q��I/#���eLzz�[�����p�ʸ�)5p*��%��f�}��R7��F�˫e20�M�ʈX�+v��fXގ�m��Ȗ���}E�դs�$M��̙P?U�:����o=��fn�-_�I�-V0�����E�5��ՂuZ:�2!��1�O��JB��d�F�I�ZHޅ�H���K�NB�x�����U'N3�B5�ݖ���O�n'g_(�����x����^�#�S�>��i�j@J��+�c9�}N^��'�͂�W!�爀�1N�(%���&��D�4���"��"�����.��w��.3�0�����g�%�ll�z��zDm�����5������I�cv����ߒ������I��$��i��`w�	J���]�� ��;�xc�xg�At5b�P;󿃑�R�I����:���u"Gؓ{��$R�51�#�?`�S(�t#��$n��?|�������Y�-EEz��d�*�nR,J#YiC 9�ɡ&���CyC�� ]�1��g�JNg�7����^��^D( �~@�Ƶ;����xن;t��a4E��Z��
*u>�**��?l�����6���T�m���Gy�jI=q�{����iۥۣqf��\ʭ3�]����ղ1���}]iKhi=W�	���d��7�`�2�FY>�����:?!:���F����>��p����t/�Iul�%�����6y{�\h0~��p7vɒ~icNM4���/��TM�p6=d:I����w�`x�0�L)|QA����!�%\������p���sv�L�_�|�z�+�ϋ�p7�R
V��WhU�> ���0Ӛk!Қ�w&0�in ��V�#�Z��Z�&Њ߁N{US6So/f�s��r��v��EU�&\G��%�.��~�J�����ТV�Ā}sʤ���N-w!�i�NRKz_d�`��I��Z�%�D�&G��V�&4�QP���=U�ޏ�z+<'yA���a^-�#��Sr8Rc�_�e��45�fl=d{�7��q�Txݶ�5ٯ����~����Xf`gx��y��С�0کE���6�S���]8=u��k��� ���o�u�CC���E��o{�qr�"=�L���rwA� �XbT���p��f�fj2Sq��]ԥ6~�6ְ���i��&���/	Z��u*²�Qam	Y{35{�����9���a���jya���l��$�)�
��q��*�lwbŲ�$qbԊ��qb����v��ZqH���mmѓ����;�cv�������i�"a�H �w-�/A9�ÂI����	b`U�CuF�"��}1�O��{��d��Yq~HM���g�E���Wk��\de˯�|�tS�5#!��p��,uC���k���8=~��p)�FPO��(lc/���lfZ��Pd�V$���m��"9�{D/�K�]i�x�
�rv�������=i�K!��xo&�HR{ki�,�,�u�\�Յ5+��x��t��hM]��g�z�~���o�EQ�r�n#��m���'�yb�NN���i�2�c�mQ����e�R�|����?c�f�m��[�!w��M�Y��xe�6.�{[�y��zQ��6H�|�3�I����~� �N��<,CL>qv��m�Q�+�*h-�7fH�C�����La�[J���wE�F�t���VJW��Z,��s�|��)ˆ��ש�IS�m�9@`�����!�Tw�U.0�c����.��uw�zO�CΫ���^�@�X} f���s�����ƣ��`��}	:
8�g����.(�5M:�����e���<��+ʟ3�ϋ�7s�������C���`��e�n��ѵ��	��*�a.A���}��~`�1�U:8���)���}�y���|lh�Twd{+"�a�����	D���㯫��մ��&��L����0�#ĸg|��m��3@�WӨ��@�B��s�"N��	�Z1Ū������ �å�U�dIi;�y���^:B��]��1�-V?��Y�%�D s�^��E��wv�՚�fAx�`>x	��8QΗl��y$),�l�ªH>�ԡ[���5Soċ�4�r��R�r�G$:yv��RLڛNt������wvҎ>�-�qYdv����G;>"��$%BB,d�{imt<@���Ü6m�ݱ	�Kn�	B��ى�ܙʓ������	�������|E��9��(�Yй|�WP���D6��֩Zk	�����s+�`�� Zղ��OM7K���F���ʉ{�$�_�R�"�Ԁ2�>�D��y;�Ϸ(~�G�	�h
Ӟ�݁����
�m��/F��A7끓vk?8<���/��0u����GD�|���"m��g�A+8�%�v�́@�遺�����vH�߫�����}<���=J�����a_�Y^�`3�툽;�WA�ey�t
�LA{���y����=V<R�B���0�l>VID���aP�~*��TZ\[R��ذ�D�i�$��uY߫��υ�����q�+��h�PwJ�9�����p�1M�����nه�Oщ��Z~yu�踘��=G��� �4r�՚)����j��;`1���G�)Y?r��W+H�W�)����G�O\iPcZ\�9�#���3�GK\l�}Ɵ͕�A5�{s��e��v@?��ru���C�O`���P �*���x�����]���Q�g��Z�K(�t�s�[@0n�~��h_��g,O\˼��zR�>|��A��E�s'���a ��9D`H�ܷ���/�\n�'��r��S�,L�wl4��t�\�3«���[Z�ߵ�an��a:�b�Yo�G���*���?%='�,�<q��������ږ�v��V�K�o`]r�;Dͷṕ��"�L�%�+��}=F(�;���쬀�6y������|��6x��$tP�!o�������o��!�Ǧbb�G�5�*��u��{���ۚ���&;9)��6�r��s���ʦ�`?Q���oa�nF��/
��a���="o�F�B�ϦB]��}
�4|3"��	�l.����,c�µ��Y�+A\,��Glg�H6"�����jM�V�_WO��c ���_��(�1mJa�+���,��0b���l�L�g���Ȓ��/a[S/�cn�z�C��$>�V��ym���,FнvAiL�C@� /!��4 8� ���M����
g{��؜\A�J�E4�����@��)����B!����Yə�:�a,�3��X�D)nC�.n�G�΅�`�@Z�!|H�f �V��V�#�<`m��AX[Vv;�W�]�H|���V\J)�~ב��%m�zR�8֭fb{I9�&m�ק�X�3��]>���o3�r�2�%@I9�� ����?4��x�Z������+|�,��a�4��5��+�Z����Y:���3�]��9=��)��!�Z�7V�[,�B��'6�6�p�t+ǝ'�������T>��	Ϭg2�di%��?�=�=>t�����
	Mx�0��@Υ#�{�O��	'�T$y��c�� �νĝ��M'��R�5���t����4I��ViT�[�ȁV���y�cٲ�m<�u�p��K���
~&v�SFGh�T�T-Q�+��֑����0F��x�Za���d^kFy������� ��M�mހK��_�,�
�]����a�/�7���KN/e�(x9E�W��i{����Dz�A����!0.W�>����V����ֈ�H�2+�e̏<�,�ffO�k'hp;�
)[]g��C�*h����J�&Ji�9����D�o++b˚r|ъH��P�Cu�������WR"��
#�j�z�ʐe�����\�e�&�uD����'E2z���O��j�x%�	܆�皎)�,�)r����G�~�?$��� ����t�����t+ɵ6u��hw�>U���le`@0"�4`�g���Uc-���d����!7�v�Q�ZU*�:��Č���A󏈫�����]W*�~��.cl�R�L*����(MK]d?FY̌o4Տ�l�°����`����tP]'�+����R�"�sUi-5��IӦ�o�,�B+���h�y�ۉ��HI��7*Zxx<���C��"�vU�DwMӿ,XW$-��+=�ć�*�#���1$-�\���g���:&��7!��cgE�-�b���Ŋ�ű�/�%Y�8�#�󙧮E 7�~q9��yFֲ�gʖ�<;�ѣ���:c�����W���פirS�MvA!j_���t "W����`�/�p˩�n@KRSF��|��mO�|=q4���!�_��yE�Q��y�HJ#��P�=����V���@�D2 ��"�����6[J���-)��yy�����u�z��[�~C^Ä.y�5�����x�E�S��lǂ�4���o����[2���=����xe�<����h���0����}���(�0~�ឞj!��p1�	r��6��i!2����l5�ҫ7�H�������q���^gn
����`"�@��X��65L����+��3���=]*%�*�"������*46���w��Q�ٝ�Scj�y���kxj��f&�_Hk�l"��m�hόТd��g�[s~I?���$��\�#"�㺶���}��6;�.%���Η"�6c2"�凴�A�EUӀ���FR������z0�XUuH�&*��,����fo�f���IΟ�2Ķ����f���G3����X<��c�����n-Nݜ����������-��1#�3��Gھ��*�E�
������	�����#ȓ����.�i8�7����	n-q�c��M��ar�Х,�_�*}z��Q퓣J�i����խ+Y.C(���؈�_�����i[���$�!�d����}%a�A_(�8�dW��4�TPƌ���#�r�}��Q�Ys&��7��`_s��x}C{i�NN�l��ݠѭ�Uv��[%\�5x���nb�������N���d�t�*Tr�_�i�ǥ�㤙�}(���9a��ڝ;�L+&��ʕ�b/w�H����XR���� �ȋ^!��\��L/o�as�~6.DC���llC6]� #��'�D,�^6��)��-�X�}�5�)�Щ1��O�q"�l~�`?��*�A�R+I��_C��qn Ɣ��ͬ�9	I�%+���gH5m����K�0 �W+D�EHQ�q������l�+j�}6����s��2{��`��k}���E-��R���=�H#I����a��s�XMg�����)6�&.1.H����c������LLVh���/"��F�p�L�\�����E��L�E�$1vޜl;�'�Ug�gя2�N��L�ß\����^B�~z�	���P	�	����m�����z[U�%��K��]�e�9(��&_��1�o&�M��r2��ԅ5r��BI����T�°>M9�k<�e�F�H���)�ZA�B�_,n�n����f7_ա'���k�M�Y�1WH�Ω(�S�_��ڐu��#�����^����q�RL�y�a��fOD��5F�\i�5+B���a+P|A�Y�5���n��mݰ>[)G��?1@������F�m�t�W@�|�]H�� �9WT�c!;��s��XZT�	�f�r5�
�u�;��S~�~b�MZ��B�*���������s�-g��^H=�)�|Ն�eP�1V�n9��Є�as��{A�\��E@�~��k��MS6�8�|-+n2�>t4�E�Xw�+\3����S�v�y�鷢����Ɓ�q:��P�����k�:l����ՙ^��E��wJ�p��Sj=�g@��"�Q����&�Oq�ʮ���=8$���&2���~��:���cun�P��0ƫ� +�]Dˮh�5յk�d�= ��KF���|������B	G��e���ksp ��&��o�ډ��?�Lpk'B%�S�B��� ��~���?3���v��h*�b�
 |M�9����p7v1-�w��i��@�(D�2��|��)7�tΤ��uG�K']Ri�瑶�9��74"([�9��W�K#�)ڡ�
z�<6If�0�"�ތk�(.,��m()@@ˈg����&=`=���1����C��ՀT���߆��/{�#��0,hP��12����
���,a�e�Y�rO,�	��.����/�:�i����>l��e��͇Kc�a|�i#����QλO ��]���մ��)\�K��)J_�V��5��|��ي�5ԍqjX���Ƿ'd���G�_G$d@^<��q޸spW~��"G�AԤ{���6�$5�R�m��և����dO�M"	/�!6(��o}�H�"z�z��6][�!�1���rSr�\�PnoCc.]��)b�?	I�n~�?��8��DA�[s|�3ص���n�:�L���6�@|+e>�r�	+�����Z(�~Oؤ�F�t�6�2�$�%4�7�mb ��jZd�̥��\��~_�Fh��������s�*ub��y/�n�x\��OtaY@�IM�J���m��F�Xz�\��s�q+�/�ɐЧ�9�U�QFѨ�}"�\�D���\g��
b�'��!sH��[�M�����9�yU8�G;����3$�d�
ƌ��\��ҷ�z	-�\��;�2t��{2�N���<�HT�eL���_n�8����Xp��z�\�{]��tj�_�9؞'�|��O�'I��C�ϩ�V�ܻ�g��猂-j�[�{����?a�W��31VX��ҁ�/g�!�� ��3�5���K���x�=��!���Bf[�q�f���H\F�լ���&�:���#q�΃��Ҋ��.&�)�}&�;���]����`z����T�c��KL}��-�I*ecQ;�ع��"6�I�{��z�-����}�@�.�&��Y�03D�"G��4oT[�0p�}�ؓѥ&���&u�(*�{��.Dn��H��F�2�Є���"����^$�y.���H �S��)"�3���g�1�$��TXV�	�43�n���k$�����ic�,����%|��jHN	v,|}$��qx�{Kr�|����O�d��[�6��V���A.�#y�x�m���$;�<	�M���v� �|�t^�@D.�D"Z��b�iɖ,V2XM8�#F��V�Xn� K�P[�h�� ��NiH[8��+Gʯ���h��g[�����e��c���b��
������&>�9r	�Cc3�t`�C{�ZրׯS�+�뭥um�k��.*Y gً���eo�:3q���4!�`k4u'��������M�<2ܛ�Tz�a�x�E.��qB��kX�yQ�0��R#��Gq�UmD�,�f�j�$��.?B�rN��
�~-ܣA@'qz��Kr�="Q����K�]䲖����i=�g��g6b'��Bv����X��of��C�m�͑D3��T��:i*�(�HS6��m��k�㊊�e�͂�| �ˠy����~6t%Yn=/΍)+��C��F��H��gY
�8�c�8zǰ�8������TO9�`I�) `��
(�tv wi����x㼌 ?�Tߌ�a%���{N8��̰o��H��x?5���ȃ�
�XE��Q��<6���"Z�ߢ��9\FYn8q9���席q w�ëaDC��8�۝�qn��۸p�rp��^�T����s�+�L����l�D|�Y�N�V��D�E�����=�;��Pb�P�OXE�UF�F��é�����(�c~�ł���*�|�݋��H�ܕ�;;��~�a�|�O���GH�R��I|�T=��<�#2;Щ�A�M2�@\���pm��̩؅ƿ*�])S|�����R�Zպ �e2�;g�؝�2�,W��� Z9�"*�c;�A�G�`�:��8G�b�]��S�M}�5�pc6x2���-�E�=J,\��#�P�8�z� F�
m���˚Mr����Y=xt8����� ��
�r�d2�@�<�������ڀ� TP�i�n��K�Ήɜ�h������[N�qW���n;x�2ͣa,������q�@+��!���������oBA�,���_���C�:B�r�Sr�<�2T���k	���vM� �aѐ%��j�1�j׭[�c\�A�ܟ��<���0B�v��9�"_,�-����	G�l��q� c�[�'��3$�=.�����Lm~�o({���B�z�!V�,t�wZ��M�c�`>=9�G{�XЛ�,���9��l�-�v��*���X��xgjqj��;d�I3�m�/NX^ó�9�@������!Ba -��Nj3T�\�ω���(����n��~�����ubu��o�E&^��G!^Ə�=
_����`qn�O�y���6�����i7u��\�����o�<uA�@)7U̸3(�SnGF�h؜T煾a�o��f�^��%H�^a�&�uV~��� :��4v��n^8W��56Z���U$���e����`���b<�[�D%�yk��[���8��!7�
Xx��x���%\�;4�Idr-[�g:p��$��҅�r�A�Ae� ���#+\�p���s�>�&���rF��ar��7���W�'\�U���M��t�2K�}��t ,���au?
��Ӯ�7����6yɱcX�0��y�WG�X�m|Bv���bP�N�@��y��F�F�㸪�I:���߫����[w�ho��'밣�q�"�����`P	g@k�'a�@ݱ�ǦX��9htƈ��)�4o��WĳA6݆�]��/5N#�h/-�W@�O���cx���A��n���G�� OC ��z3����О��}m�k��TJ�f���1�+н�q�"(d��z�d�/���([2�@T�e���{���1�)��mkf��!��Y�a�-2�����63%�m�D8���u�9D�R]�h��c��Ю ���^�@��i��O���$3�5`I�o�)��7.M��F|BX�y�u� 4	�L��.S,��b�Mv���^X$���f�"~�Z�aZ���O9+0[�jN`��6�y}aQ1��e�8��i]��(������c����N�H��"�m��wB���J3u�����b����Rl��{է�j�3�&�,��Ň��VV�Vׅ{͑�,~I����d]��V�ւɢP��ŋ��ps����
��� Jd>�R��B*�qu<U`����V�Z��H�c]p�=��V{�Т�m�y���n6�>�Q�#
_+]�M�]O<W���\D"�rPSwwp��C0�&`}��?�+�l���b��׮C�Qx;&|���h��.�2�3���	Y;HEv�w�n|xR�j�S�j����c�[i��L��6@����?w�gg���F�wޑ/�}#����k��"����&��!���d�X���sb]�|�|y��6�8�5�a��#���?�W�1����qݐ��1F��>v��8���S�_�����Ɣʨ[��d�;{��Y�GsO���E��!#���b�R��ݦ.1�j�����������W��lP��2��t?H:�1�^T��� ���,�/7C'��x�5���W�
�.4+Y�'��$�n"� �Z&W@ �@m����O!��{�\2DQ�v@t�1�u�@c�͖��{�y̱��Wn���?�U��R��䬅t�%��6�{�&�?3�.��Y�~V�(�XQ� ���2��Ɖ;�@��7W���x��/�Lw����]��P�NᲵ>
����o�?D����F��(���F��t�w	(q+�U`�����.���/��q�J/� �bFЬ!�ޮ�t�V^�d��sb!�50W�	-�
�jb�>wi(�ͭ���\-���E��ڜǌ�6=?)+@uJM0p?��G����U�A���Ի�U����T�`-������Bl�$ک��U�ӌoݺ�KW����K��������b��¯>c(�R�H�Hzͤ^���;w��,Ӷ�&aU_��'|($'4o��9���x?^/=�bJ���%nք��?]39 ~[HVe���4վ��>�o>lցn�s�BzT���,�2�����c4�!.gkt�vX>YPٚ�Y�>{�\��0��֝(IZ�S�;,���gp����M���=���F{�>i�
I��u����3o�0}���LB� ����6i�+id�;� L��W��*N�1LG}�1h��'�����?/	��:궸�*�M��h��K�ͪqB�4�������?+����b@��mٕ�r�h��Oxd=ɇ�j��{%��jq߭��Yt@x%WR���]�2���L�A���vu���hp/�g�ߙ~P���10�3��@X���;�[�EHE��JbK���X҄��ӯ��t9!?���5qi�U�z��X���
`,��J����.�������a
u-M�3��]�.@��2�r�59���Od�Wbϗ�4�b6�	U"M�WVNQ�����:�������"L����~DΡ�H��ˠ��G�i2�~�ٓ}�Wm��r롌�:�M�#R��g�8�$"u�g��N�>`��7U q���a�y!�sB�6o9:�D0��(i�h�c�pp�KP�䋑d�y?aAc���4����r�Ҝ���}���v�l�y�C���QX�#߄��=u�K1k����%����uZ(��C���o��n�zuIb,���PN=ֈ7һ�G �o0\!��ڀ�k��K�V�
3lf���@/:�+b�qgقz���#�ԖgÆ���<�M�2������q>�T�?ʜ���$TG��v�Y�Â��b.��T��ϖ�K^z���Lۧ7�{v�ݽ�X껳�];��e���~�*���(I�GY�7���>h�eD���~f���g��z����-M<g���v�Z�lD ��L����G�P�,��N��Ħ�)1Y������������V0UCh�xPɰ	HD�Pu�vrZ��q��i-�gdD��}}G���r���_l�$İ�6�6�l�[A{�B����:�&D�@���m��+�7�G���2@�.f��&��(�i�EO�Y
>]�i~�Bg����&�x<��2��#��u#�X*�t}��5���ª֢¯MӄBrzyG|\>j�ٷuh@�	`���U޻���<�1��9�P-�����(괚������(�����ؕ�v�B�E�9��Z�>M�}������uf���3BX��Db帩��1��ّzs��)���ba�	ē����nJ�XU!t��Ѡg:iG���FwޣE+�iP��nT��r��YSڲW��gkCY^�0��-wD	�X�L������/��L+dn�t�����tKzSΖ��O��F�������FBV�x���	����[�����$6a$��si��p�T� �x����S�,�˕���6��K6ȕ�f��w���.3���f���_�9������gln�q
���o��$��x�="V�<���1(�x�$���4�Di������;^:˦6��lvH�������~�P�Gz0���������0�,RM��$f�
�%�+�$�ite�mM��!���?*Qf�-x��KM(�,�Z��s3��M��RǞzB0/O0I� �=`'�����.n#&	y�������;,ȯ��_~o+p���$8e��9t���&�}0��g���D�w�,������	yV܄��Aб����Y���P`׶&,�C�}��@\��#\lt���EF�#3su��]0nW�xp�����&1
"�6 �)�ǳ%@J�-��X�P,(N�1#�k���2R�8�P^�J8m�5�c�ٝ:0�B�d�(�x� ��V���k*z���X��\>���aD}��%+�U�no�+x��%��W���\�Y���C�����Fȁ3��a�-��M�?{s,����LT�;��В�:u]2<��e�U��B��&�2PO&�J�l�|G8(+#���^��&��>D4ﱵD�H�������ɐe3�� �Ҝ��F�K���"��l��A`��#ٍ��ѿ�����D������ ����𶶕x���Z�Uj|��>غk��!���T�- ի�Mo�1j�f�o�P
�T�+�ґ(��8��Byℷw%��X��)��6�Wr�E�nn��I�o�(���KE~b�� ��v��mA��ʼNK�}G���h���;UBj24�4�-:�V�H̤z�~ش�'���zYpjb�P�~Z:�AMÕ �V9�C1|��%�vѼqM�����Z�kd{	�tb�P�%�����Z�5⸍o{L�l�I�����,��J'l_�)�<���06v�B��9��t_�����b;��q�+�𖝠�a�82<TY�$Ȝ�j�$���4-~2��؇�h�>=�/�kgvWR�D�r��Qf�)߶�}���KJ�D&�Q�gM��5%k/%��M���7���j��Y�U��r�eQ����0�k"l��"��uHR˘�v�B�c$��)�aW��ϫ�=�_9S���r����l�6I4l5���`��шNA�[G�^�yn�5���y�$Wlؕ������/�7LL~g����*�9d��Xp��۴	�r�n��%��	j�Ǚ`Ke�I�%aB�씸�'�g�>R���Q��g�������Րe~���}.r`Ъ��$�h������˝I��Z��Df	���r���d3J��ի���;��P�>:b�����ȫrCey�%�>��<P��x�S��E~�$���T�E�t�Al�MBf?=�=���۝~�A�`G��������b�����_A ��Ŵw���'�dٲ�?V��d���x��#�R��1�NG��]��a6��orG��|�:ކxYe����7���Ϸ�+u��- ���� N�ZC�I��qr�����S�I:�+H:�%��,^I��|_δ>����.�3�p�h�iY����;���Ҽ����L
z��_���m~��e��ዴ����XV���%7^��Z7͡F9���B�c�fj���uqK:y:z���G�`�g8U�Y^��	MI�:��	�W��G6/t�H�%�vO���@�u[友?��	U����[҅X�H2���J�I��v��ڱ��͐Cʳs�3��xS=}o)?H�w�4��Ƃ� �t�з�}֞	3�7��:�A�M-��!��1���3���q]?��+�X����5ir������k�% ��^��h���&Po�6��W�zi��I5~�>��R�T������(�="�����D�r�P&S6�I�;���#�j�s9��`�L6b6oD���p�T<�ke��nW;�����lN�{P�i1�ڍ���7�O�l�x:�%n�,Ab�Rοu�K'gŎ�O{^ �t^_������Q!��>Pr�)��T@~�*�y[�0�g0.�7VOhx������/����ڸv�|)�k�(D�*^�m�
�3��GIT6U �oPV(�͎�|�7�uJ�7�X)9�`4�f��-J=}�����FH�� Gÿ�{M��׫钣��y3�ďYA{�X�^P 3�!�������;&b�K�L`5���	��[Ӆ���k�_�4l��CZPS�R�p]�פ��y�S���^w��2
���g��N��:K��r�����f�N��J���@;�t_����P� fd�^��i�/����K����-�	�����Ķ��Nի�6��HZ��eD����ڬ�]*8�	���>�X�x��@m�:�����6��#�qeJAGDJ�-�����i�&����O�,l��y�2�|ܣGރ��a��~���Fz�hII�ر ĹV��FxB"�&���޵����A�@kG��دd���w�`��?�kiҵU)O0�fi��X�����B!$$��2@��A�O�2�j%�F]�廐B{,X~,HH¯�
{� �{ y�P��?���_.8���*	~����b�T����%':���afS����r�������z�[�\�̧d'����|r�;YG�j�h�H�kpؼ�KC&<~g�F"�1��g~�'bb�� u	��p�iS��Ф�Ы���֝y俊l%#Q|J�x�
��,##�&@Yu/�Y,���<��Ts��X6�/�t���Y�X1޴Q�V'xP��^��U��!2Lo}|k�r!o݀��<��s|��"	:�q�2��8IbB����mj ^��������M-�Oŝ����Q�
�b�ь]�,���~ȷ��q��o0	� ��%��$o�������2u�f"����&�{Ll]o	��M�� �l��z%t��@վ����I������j��g��k����!n%�F��c���+$H��}����N����v�/P_%�7(��~A��li&j@�4�9у�?�4;]���¡#�ڂ���]��#���I�d�I�6�'���nLͰŲkĸ߂ϫ�i��Q���6���/�o �P(��	��ᜲ�8���K��>�nH^����Q��*�q�i�R�Y��w�-�ۯ!j����-�JW��,;�W�uϠ��P.P�,����DU\�E�cL���v�)衼�9���+������`xbg=&LOi���*�V�fl���sv�3SP�M�nl��g�Y����D��'	�Ed��*�s��rn+M�%,�����d��W+>�l�ջS��%Of�.ҏ�;OBA}SK|+�hS��X�Gb���U0i����YfY�����G�5���Ly�@Uw#h'dߡ̊#�3ka�Ng�r����q|QG����5q���s�Fճ@2�D�$N<{��\*�h{v.��\�V
jA�ȗ�C�&RҚ�R��T�ݪ��:�`���<%�x��Kl,��Pf( �����ZO#8��������l�� ����፤atN�@�`)����b�d�F	���P�+Ҍ��.�&P�Cld�`H�pMKAO�&�����Kus:��4~� ���ڢ��^fJ#������������#veE�������=�F�>-�n�6����P5��4#eE��U�͵sR�m>SQ��Z�w$��*C�Ć��	ɱQ˴O�K�f�@a�t��]���>b��Y��X��fQ�d��GM����}��"�	��Ǌ���Y�7�G��B�ܤ�d=�ZK�D�G��+���`����`��'N��:d��/1�5�T�o�w���B�� ��%P\��Ш�'�.C���߽�exh��XE�[-�((i~c=�Wy����%}qx6���o�}���(��c9�z��8.�٪4㤻If�_�#o�!�ί':�Y�`��cl��%��R�� 	��I�,d���t�GX�u
�,6��j�Hkdg�1� ���M="� 	)��Ys��U���_���^�#���F�W�_s�%��t
B�8.ROd���b���~�k����{�q�͋[���Pvc�������7kRB�or[F�!AQ�4�Jut����V9@@J��xY���X�d�ܰCǺ��m�C�9A�.c�	��^}t��XՅ�Q��S���o���qt�*�e��*;��^�1��t%i�)B�h�(��SPʭX�-��M�@w�P&pD��}Wp8<h�y��k��ʄ��'E�f�Bʆ���t�ϒ����1���/�rE0�|Vm7���Nv�_�s.�z��~ܥw������ɦ�^��}�*��fl@�I7�bb��c|Ǿ�Ot�4���{��KG�Sf���!�MD!���>��R�V���i`>z�#D�>rP?1��@/ƨZU[}>���������l�����w��r�6
��]e«Zi ��4���N�87qi'𬁀Jq#:�v6�c�c���Qo��G�8���u�WD��˒�Q�
��T96Xl����'4�^_N���B't��[i�p��w	,�(���]�9�GXe�e!��M��w�LL'Q^��:'dE��`��- 'f�Xͩ��Їn:r�y̥�T7���?Ē�U!ŭ�o,|x$���_��L���K���N}ML���봻*�F��x��P�0��e4��WI�T�~N�g�7��+w��Me�WA`p����-{�Ӵ6�^����MZ�"l4ot ����|p*�X#�GC�;�����_��=l5�Pg�Q�UN����#� �mD53K���!������G�ލ�k�O����e��v�L^�&^�% �7� E�z����A�b2�M�:i�V��Fl���oO-���V*(K���:}��Z�Zt���"Ͻ��x��P�!��f�aW��!������O���l��o{ܞ}��/2g�����^m���Ҏr:�e�氾���:�Wx���m霫�\ ��ᱰ��ܧmᢅ����^C�/�J>;3�` ���u�+����x�/l05���e�M'�5�`���:�:���K�8��N;,�s�e��cD�Z��$����e���B���|���eF����`.�3Ss����J��I/�_�Xs}��!+��B�QEۭ�;���y>\��Q�	19��/�u���������ի0V��ys�?���7C�%�=5���i[�j̽�lh��#�$�%����f<j�����ͪ��ι��%�S��R7ޚ���鐬���[���"�죉RF����T�U�+��Z'T�+Dx��>d;�a��C���Oُ���7jB��2K@&$�9�++:8?IT�#n� }U�=�۸ �ĵZ��2�Q��춪[q��b�Z��@o�(s]�%6�0@Z��&Q���I<}Eq�����k� 
��V8w�s������
��*����Ȉ�rJ �:É1�_��YYt%�k�Lﻧ�,C��*�u��h޳�;a^[��I!��cU��p� \�)�hA�%
(� p/ ��h��f;�`ֺ¾ea#i��a�[�:��5y-��y���*"���غ7���K�T^r����C��|�E���@aZ��iB��Aj��6)6����v�X�`y�B"��
���M��t��Z[{oTȥc	BA�!!�<��,�t�jo���;ʮ+��2%4��W����&87C�h����!&m���,��Vr9e�r��K���:��h/�Caz���i�H�|9����&��Z����m���G��'J'�#�x���(�
_�y�-��+��NH��j�-�$���d����}���Y�b����WIS�1�2�Z��5~�.�?�l:g���7P]x^ά�T���8�Y����S�{�����0�����wp���˻~������+X���H�E�(�WX����#f� ��Z��N������Y�I���ӎ!������ܵQ�?�R����a����^�V�[�K61kJC�����1X�	�=�Z��c��[Y����Ƈ�a+�g�e��6߂;�}�^�&J���:�wHH�a���1�Sj,�b�ЈU��w��,1;?�88<��I$N��~��E�]u)�į]�u*�����<��e���vJ+%C�a�{��c�Ry���w�X��	�����/Q�#K���������MV��^1)�p)MA"���c�z�����a"'���34H�ݥ�ȼz���&V�R��&a�a"u(G)C���o�C]|�A�t ��~��8�.�c>�-�;�|b�[��8b*L��[O�bd�/DJƦ����_q��M&{t[�/d�Y2b�
���)���.���O�MiD���2�$nJ�`Gћ�$�����#S~(o��x;������u���3���}�;2W�C^f����<��[�v� !��ٷ����4V�vx+=�Ȃ��rp�[������U�`x<�a�a�zg[���G���
��6{��Da��XR���;f��;]�86���M(	"�7$ йul�#$@�7a쳩���ר��O2c���tI]t(�dJ�����;�_%AA�G���V����T���ua������I���7��������HVG�e�1yd%A~�W�\;�TeZ��-5w����[���|�L�e���ާ	�:g���,�_�� �C�5�<�����J������c�&��a/�J_h��ь}�N��Mi�&s�{F&XӪT�{�&�y��w����AT�f�FߓN
U|��t4�қ��lKA�k�1�0/����(i�h<��g�r�,с:�0�?�]E��q��"?�we�	^Є�"2�ύ,:p{��&-;��ĜH�!=z�G��W��#���X-����wI�)���j �m�0���<�)4��/n�8HA�����m�/$b�33>E�$�U�&Cq�Z�ωc�C!�lKai�>�ƣ�`��~�ώ��)Um��6��g��]�RbU�R\��mK��H�׆(�rU����:	Ќ�Rڦ�+���ׁE���8\��Q9�$��F�·l�@�-sĹ�+���C��&�n�ߋ���p4�&��OaY�6�л�����Q�S�X7>o�?��|Ɲ�087D��NhX>*�\̟4:w$vx`a����)<�
����c�+�D F����-�Q�< �� �mS
��Q��	� 3d<(�����[X�:�+�R��plL@�I��H���߁��ф��<cu�
�������|��Ϭ숎ߔ����
�����N\]��Aj����2u1J��yE�q��_�9v�^���4�E|�"x�*5�3]Q�3Kz�(�W4��=.l^�#�o�� ��ѹ�-�U��=�m0��<W��="���� |Z��a�S��e�)�C�oV�Z&�}���T��+w���W�^��8�@v�K¾�%Z.�䚂�0�'�EG���܉Wk��0�S5������n�	;�<�s�Tc
�Cn���Z�3?e�ǭ鏸�w56Ϻ�y���2_ͭG�5�9���Ⱦs�����E�� �al����v��c�����L���.�s����|��y6GV���cl������VĘ_��%��!fAE����j1���Y�=R�{�qT}>-�E&�D��?j=����&2������!�cW����̖	3B����7q&^ۋ�)J94�>�c�������ŉ�K��W<�H�p@3�H@e@֎��_�3�ތo��p����^�hL*P=�n�o��˚כ7���=k/m-��+�[�@&M����h΅���_K
�,>��"^�Q�4q
�K��.���J�+�
2u�'{��Ǹp�*�En_�<��V�xt{�(;O%��u�s�h�,���y^#P�O�{�p�]������+�
o���c,���V�;�c��Sp�F��3C��X�?���N�l��A������A��zv���M�,y��K��Z[���$�l��^�/X(~i!D��T�$2R��Hq~�:��]��Z��&u�Rڻ�-%��7��c��Gkצ5�]���P��Մ�c�HI� �hIj�F{6�v����2��z�c�����Zߋ�Lp	���g@��U���__�f֘I�Rݙ]XC[�l=�'�
d�7������gÌ��;�gk�g�W�jc��Mغ��u���JHJ]YH����3(L,
.��so�&)���|�]I��-IІ�U?��:(��]���XCO���I�Z��7�| �I�1��7�?���%��D�HL���iQ�˜p�8�^H��&�Hs{����E7	$�tQX�6nϯu�X ��O.K��ܷS�BD�t��ʝ>s���(&�m��t}F!��G�_�%�m|0 ���I7��Y���-ŋ�}cʧ�.Hj������_�Ͻ��}l��%�f��M�_O�ᑂ���XL��U��L,'ۍ z���yM
t�qޫX�^g��+N3�Ǧ���L�7-���xI]��Ǿֿe��e6��PE�	��z�9���K��X��u��#j/�'����P#��
7M��{`��_� �<����Ŭ���-Z�"7`�0w�&R�"��n�FQ������;�P#u��:�,M�9w^�����1���G�Z�6���]9�OqnuDa�A�9�ک_�	������h�v`���'��J��UWY���7q"��0.�6�c%r�C_%Cl�$�H7dr���ҴТΛW���{*^���;���Q�g�ሽ�໛)��sz�A�A�rP\ѡ��%y�����%pZ���"�h+̈z*��Lk�_TfV��4雫b}B��U�?*F#���S��&�H��EP��0��^�E��JN�������H��	c��/&Z�A-,(��9+�&Ϋ�}�����q�y�e)�X[_&�`nd~#�@;���h���g��/uM9����6����n��	{{	]Z�,>��v��I/z6���b4�i�+Lۤ��[u�uk�z�g����6�rʀ=-|i (��bZ���D�[�����7�Jlm$�IJCr����4��y�3�UT0 ���9����/m �P�ZčL��"��Ϳyn^�$H��ٝ@O���{� -:�^��?�M� �ܒ�� ����^@[�[�&X'Uai�%��c"9눰���~�/G8,OU�@bP�G�����T��o񫨏��=�.�ҿ���2�� �8L� � �.��o�ƕ��Z�����D~
���`�L���a,�T���}r`�~�3��+��и�E9`b_�IK��k �SN��%	Ǉ�KhUnȍ������)��Op ^
���q��G@9R���N�,Зn�2A��u����B���^O�'��i�t?Iվ��:Zr�h��%�"�]C���"-1ߚ�1U�����g}nFl��X�%Ϭe��?�t�CZَ��3)=+[��vuݘ(�6�RZca�4MnJ�W�G+Ib
o�顨U�|��Hriً2M$��+�K�z({i�yu�S1|�'M�'T���L9�"2w7t�VctHQ�u�cί�����e��}��qiϛ����2��H��"�Ƕ7�x*r�˷a�K��WnG�g�cYcd�z�O�&��{+^�"��!�dܔ�L�N4[�,�e"E�gU�˜|B����	oH,JTJ�������Gl?x7�v�,V5�͸����Xho��_�B�優��kƚ�tl˙"џ�M:��'�\,����Q.��DQN�탚1t
:�e�]��#y'���Ƥn�֊�bB1�b 7��pnFm��E�hg�����%�<�°�g�t��N�iK�J��q��W���~��J}�-��8f-����®���Z׮K02�^�BN�?O�.7�(�0��j�9��Rͳ��9
pH��I�ݔ���`ޭ�#!�r�N�{�8���=��E�[֣B_���5uq!{�T���C>,ߏ�}\_y�6�'Pl*�C<�kL��^rjk ��Y ��eczvJ����K�z\Ad*��]�,#����m�+gc��[mu���0��4��Kx(V���j��q*�t��6ݪ�(k%�m��y�?��ǰk���
�����X����}z�[���[�řF�U)�ٓ/,�=�%�$���Uŗ�ӱ�|�T���r�9�h�f���9�3�P��f'q��������c1����[��b�Q����Ϸ�� r��v����˅�a�QK�F�`�1���BB�k҆r�i�o�Y���j#Κ9&��e�˿�k�s�K���f	���	�	 ��a�n�/�7��祤3�R�H}�|мQͮ'K�t�k�>�[�4�����p�+{�JA�J`�8f����c\�f�3��i��KX�pq�5���d���Z-���bb��,�P�h����g��0O��A�Y��qRՊ�CR��Ä+"C����ț��6g-ܜ�L�N��:X�8�ՃLԨ�<ȉ�.�1lUojpW6x�~k��g��w0��n�u�����m��Cכݫ�?=S�?Z�;Fe��W�U���dR�ڬtM�k��,���L�t✜�|�ē�4�@CA��G��Gڠe�@�B�E��5µ꼒�8�
��wl��zX���`|��ݛ��q�9۪D�խ�~=kwb�K�)��/�u>(��n��N���i�V�-�r_���T^��[��o ���V����Co@������Iѣ���<S�����>�4yR��vI�
x��Zd���y(?Y�F2�!L�y����~�h9�EEu�������B�^�Om��b�E�loq{�^4���A�u8԰�Ǽj��2�R7�|����-S�	>���;�l�n��RI`f_��X��h,��g��{FviN��?<OK��M�]�Fh�01���78��_qxY������B��B0c����eZ_g���K�͌�5�J�~b�Zpc7�-���e���|p85K�Kï.<a�`��*-/�}�r�:M�ɶ,�f%�fA��<^X��8�1m�V�t�Ժ݄RaG>x����^�O� �֊�`�����26i2X�"A:t�v�Vڗs¾�.ݐ�&�V��ԥ��:�����"�&'����{>WMP1ַpp%m��䟉O,dxg�f�G�L�iF��-�t0L����C��|��2:u�c)���tp�\�36����2dd!7@A�3�t>9~��9!5�˝m1G�
�TrDF��9�@X٣�%���j����c�1͍JN�e|���L���dhH��9�%�$m�9!at��li�H�n�v��aRJ�R؎Hm9ns�+#csJ/r̽o��Y��������G�Dd*���Gi6�cН�9;��i�;Akz-B,�xxV��p���k��#��N��I�.I��7OI�d��؎��(Q�����Ӵ��m�#�f�D����/�h�!�m�5��Itr����.	��z`a%v��.�2���\Q4�0ĉUF����vE���j(����V<B��U�Y��c�Y��x��зq�z�?kO�l�x�Vt�e�ڢE`^Fh�2 ��oD�d%���lJ�B
�9	���r�^/r��l��^F���6)P��`/��0^���FON_ �));iF�S�bBL��=X�Mߋ�����XI|������CQ�0��4�Z���N�}������j����w�o�;L��1��42�n�qI]�Nn?\�����;����X��CE�|�ot�G��ʐ�2�	=@V4\����Z;Xu5Te:�*�|�~Y��e-�u�gȷ'�Ķ���Y��O����=���{!�.��b����)
B}�oeӓP�7���I��!��a��߂OSC/��e'�p~�$�j�f	���cͰb^��=�%���W�{�Y�!!�$�':%��q��� ���.#0z->��b���#Uu�4rU|[7��M������V��VC�U�mI-�����%�|aP�O$�3�����FI璕��}�.�v�j����Ecn�O�����ӟ�~��OqQi��uY�^Q�E2�����jCFq��Q�؎r�;�C"Dm�}��t}����fT�`M=�6Ɏyŀ�Ց��Y���O�'��W,#�:]K8�|o}� zs��&���e�L����D�(�%�+惠~np;���U:��(6eA3������� �k���:Z'���	�@�2����o��l���^�/3Á)�����ݦ�GRY���Z6��?ؒ����&�Eآ	�M�?0G�ܰ�]R�]s]!�:Ҝ��z��Ё�:����#�0yS�@i�N��V��:f�~@}��%{ܺ3w�.B`ugv��{����$D ��ۨ�����0�,F��I���A<��5K)��[�m�m%U�f�V��8Dv�->���^d�a���q�c	->�vs���p=��OK�Ʊ���3#������)7��Z!�:���fY��>��"gHA����� ۿ��D,
%G��b�÷6�H$�i_�B�3lR�|^���@��I�:aR�;h�����#����=Y)���Y��`p������A;D,�;y��T�3�x>����>1������K["�VSֈ|YnO�S�(�U�0����_��ڡsp��$`��#�Y�=��C�hf�)�a�s~���t}U�ڽ|EV�E��+C��=j<�L�Pϝq����6W����J��f�O�ϣ�m��ٶD��VG�~�D����3@�4�$*����܆�e6�m���d�ᕪ�f1��۾�z�p'�ՒݏF/�[��e�F�a��O�T�Y�9��Z�b�l_{�#��Z�B�{J��Y�6�^e����9H��}���	+�2��E��� �:B�%\�F:�*|��Q��g��J��\��e���3�r����B1��:��čˏ��e�6[��R��=��^�M���rz������"m��̶��^��.|��Ϊ`{���	���r���h@�M�5/�I4r��Ǒ\�8S̉i���?���֚�Q��hQ=�����4�m�3AF:����!�hal$/D��f�/��P��P=��6���U�^o���l��R����K�p�KD#�	����`l��`����<�������% �U�-��{��-�84�������=��3�r�>���)��#��N�v��D+��	(��_<�C����������d���J��6I'U3�S8c����9*��O�h�v�˛�$�_�nAN=$�`��|��Ğ��*J�:1Ѧ(�Ÿb�!�7|�`=lԄ�ic��_���ZD��d�<�����aZ���U�c�-,��`S��98���z~
�M��D�^�IY��^!�1�G:�<�a����C,֭ދH��!���в�bd�A������	-��k@��7W��vk�_�!'����r�q��Ɋ�����:d�SQ����fS�$XD=+���N#�aj.�u���RY��)8$ah�R�@�ʥ�k;�H	����&ظ�⺐SW�e'5��/R�L/�25<���宫J[�<_��w~��s:�x��C�����@[集��W�}n�@#�hƴB�B!��U�'O8���z�9r7�r`��؉�RJC�\
=��
��P�;�s�A������_�h�1?������cq�ς�l�^���u𷋗;.2������6A�h��o��N=�/˾���*%ڋ�������t^����W�,�b�y��#�;E���4��h�+Q�S��f���pY�eq(va�Ķ�:����S�� �~i6���i�2u��	@������p >�VHQ���ߍ�[ji�M��]�0.8�^cm�����~�9�)���\ZP0sl��J��yer�J��l��.h��)���%���l��7��B:�@Ϻ���f�/ޖ<�����(�R�R9��d`L����7(R�!� �yY�A�2w�BE|�"��#G����������o�S�ơ/X�N7�O�ӫ��zƥg��-��p��ky^��ؙݺ8'�P�\��LW+��T`���(��Q�9G���xu2��6��Ǉyq�e:��x �]����K�|IFt�Q�V�CQA�h�$�����=��b�d�w�a�c���j�,��Y�C9�e��GvV`{n;�� ��?�D�'�M���|�����*�H�P4h~b���$-�02�| �ƥ�l��oi�e2�I���&�Ԍ
!����=�pƊ&���k��.i�3e!A�5����Y5mkCI�
�z f�>����aq��l"D�I��0�����ڳ^␲�JC%��-O�I�@�)!��5�6M����ae����T5�R��0����W�Z��Fђ�ʂ�L���+L �cd����uݣR@��n�|3'_iѴ����W�Ɖv�����#�h�X�pHr�v&��2!ʄ�Ӌ�a��"iC�'�ӿ���͍.�V�u럨��t��b#l�lW`����5�8Tvr�7hĂS���	�Ԑ�v5|�P 4
i3X��~O2�����;n�-2�؂��_]��P#������e�%v93M�����4]��6�98qG�ķ�+���Iɋᡖ�ї�؈��ɲ�c�-�h9�2�����6��܎�0��Ɛ[3�qg.��_�����`ށS�m[�^ <�OSИE�j� c��?d,c���(�7.�Y'af!#U��HV��&�j�e=�1E�fHöa�R�O��chɮ=�L	FԸ�����P��	-�H���YV%k��.���j!�,w��H��y]Z����ߓOxg�iԒ�EcQ�����ˬ�<JGA�6�V���76�[|��v���Ʃ�Of��zΰ:*z{��k��}��B����4t	�|��j�ʜ��"����������1Q�����ݐ��d?��Ĝ^���!-sD�^K\��d�W4����
Sq���h�@%~:8�$�:��BaE�ʐ<��X7	�W�������U8�+�šʿ������T]f�.5�)����239��[��a�6�5�j�rNk�4�co�&Q��Z+���XB�����ݨ��<#g�]>c-D-L�r{�M�T���c5�� �]�r"�0���I��W%)���T�2k���^N�C/�x�y)0
��)YLA�m��9#[��*�K㶋����v}�qfuL������ݬev����0�h�r\<f�E̘��E��qB�m�U�J��s1T�30u��0K�@�G�	�='�Vj$�"��[���#E�`�,`4݆��$zBn�h�sN�_
���Ͽ�s�!���Ge�,�O��J,��g�Uߡ��dyV�Rv��{�1�����۟��흮�u��yE��M��>Wf:"��OK1�"��@hZ)e��e��)z�N����Alt��ZH"�+�1N8~�ޠZu��S�Ș&�|c�(B}��}��`H�)Z�)�NO��(6G�*�%a��mͧ�R��59S^��Ǹ,���b[­�q8��gzT���qE+eJ����o ���-���@�̈́h�M+7�$�W�' �vn���8�P���0UM�y+�K�VTG�sydWIT�@���]{8�(f�~Gf�sG��&��ct��φk��Y��ٶ&B����ϗ��)�J�}�V�P��A�L�*��$\^�B󦢾���g+��]6_ ��>ڻ�<�4F����6�[(�����V�����w�����<�O��a�&�+^�6��-�Ǵ习�I\9�ۍ �{b�B�� 1)����O���y7�Ҿ�����`�mX�U���n�Ln��֒�N�B$�~ܑ��qN-rV�#��{�B[N^ lB�2�*��;��K��.9)V���uS@�c7 *d<K;F�`���BP�ٛ���pG^�T��@Ƌ���;L2�oI*(lT;+kfeRT^A	GSk-�����ƁWً�)V�C8.;�5X+�`J���`B�������~�{�Kr��'2�l�w������NI弳J2�9̲�*���e�� �8��L»���a��5��v���Fρp�yL�Z����~|���r����D��(!'�,?&se���;
�]43��Y2���id���k�"�ykŦ�3�^l�Y��E�1�G���W���3�r�<�|��x�=m9�������K&dϸ���V���jem+y�)J��Xb����DAfN�m��8�WEq������~��
te�@k�Z�v�PEpy�� ������h�L�;��R5D��Rx���2�U�ٙBc�Z�C �x�_��O!,��:�/Oɢ#�Ǥ\���2	e�$�!]��Xe"�����n34�ʄ�6x�.��w��y�����ר�-�!{��ؒ��o�L����V���(����ދ\���Om | }N�z%]N��ǻ綧U���`��C͘L��u5�n&H���+��#g���)H
r�B��2�*�oe�l�K��XSl�n0I.r�gu�'$1��u��4��}Į7�É�^-��."P	F�9�m���MM#&���jk�m�6�jb2Na j�aZ�M��w�0���u����Te��+O}{��[^SU��xB��R��?Zod#�l�0B�{���˛���@��G��gn�w��	��a����0�l�ʦ0>c\���{<�X]�y�K�u⎬��������Uԩ�3�(�Vc��l2�]���r�\\�j��B7$Hf�oI��O�����VpV�	I)�W�����5ЌQW��{`�o���흑��Js��?8��w�r�{�Z��۞�ő5��l/����U9��t��g�1�T�u��2�߬��oi��%�A�6R��f~�?B�%�m;'t��-��*�)�������[����=�Xb4.�4�]狀Q���\�Z�n��Қ���n�O�m1S�LY�j�D�6;�=s������C�/C+��
��ox�s%(2&�R��"-ՙ/�U�kYD��-�~��c�杌��p�*�5,*xr���JeV=�d�u�C-�f��!Gf���V�0g�ݛ�SEG�#Fjg��+���'�\���5���uO�_˝m�<�?		2�-c�t����"� 3T��� �ղ����
-f�9��ºi�{�0#l��v ?mӐ�H��j,Eә���g^Մg�V�u�>yc�7����m`R�%�!���[����@M���|E��@�͚h����Ex��خR��3��[a�CĬ}֮�6�k�M�uCsSTRQ(�H�Ηz䦜+)����lO��>���+W�-�R���'�e�dXy�m�𫉤���ז>�L���4� ��C� ������gqv�y�dm���F��/w��B�I�q�;E,k���`��3�^(#���0|�]i9&ds�F��9�[��,q�Z�\* q
AE+f���b�|l�=�;�Tt��4�vЮM轠!���{}S�
�X)����ʻ:L��)j�"Ԭuǎ��`xwҡ��O��e��=����[����,����=Y�e~ u�e�X�����r!�=�}w�~�0�"�-)�ZLKp��Ԧ�80�.���/>��N�|.WA�%��"vxb��J���������hs���
�2�M�su�E��ѯc8�&�/�}�[��n|�dZ-E2>F /劗m�_K��.�},ꢂ��K�!y�_1�/���5=5�J������h�������u�	|*Z����hԃi<���\�&a�ۭ�/@I���EN�{�+&i�C�1�]�H�G�^j�NS=��H�����"vmA��T0�Ě����@���,H�4Z?S�<!g�6����*RF�n�I�8^
�/i:�l�"�@VBeb�#��#�H�'ɖ?�ge�������:>�>���_p%�� �$f�b\F-Q�6Ϟ�3;��-V�n�;������9
�|�N8����໨�.��ǜ^�e��U���>�w�V�m�y�Y�v����T�C7��Í"Y�*���N�,�6=�%���=aÁ��5���	@,_����M����,@���������ٽ�-�CF>�ed�o����~���gy��';��	��D>�Z����{���P��}�@\Ď�����O��@�V�d�4)�䏾�+JX)���A�[]#ok��� O�AD����4V-�Z[A�г=����(9.�q� ����:�L�O�1Sx��;��2l
��*����I�V�+�=B�ћVǹ�K��5�����ad�n`ٟ	yý�Fm��^��gf@WO�)�ɷiy�u���[p<3B�=PE3$�x�c`Op�mEJ{��$fb��s��k8>�P#O٭r�b/��t��i~�NaY ��o�~�U�N�*�5�R0y8f��5� ��>-�B�p��CN�� �rj���0�W��l�������e��['x�V�W�Ć���O���$A�D��[�+�!�%���)+ܧ�'hq1��jN0;U��������7�!��o��ەE2$.�R�⇷���z���N&K�)�T�Q
'��s9�w'�gt�s¸��Ӯe��^�H^F!�rE*���V��xw*fT�<M�	��Ƅ�-��'��q�k�cQ���9�6yF��;����s�����)�o�������<��ì�K/U�D/�8,������yF����}��n*�-�i~!��x���̅���no��Ϻ�;�D��(r���s�l1����7r�N�XPKꝇ���t��Y����4�<곂R�r�K�}Roq]���lˏ�+4M&<��_�s;���PR)�����oB-e�8B��pѫ��׹�(��W-�N�m5u�� �`��I�.��� O}/M\		i��F86��o���<9������>	�U�3�ⲻb/�u/��M}D;���o�qbI[��ԌJ8*����ʱ��}�
� ��)�f�ʍ�,9Z[e#�6��)�	�V7���}O�ٯ���.)u��j_:���G@P��H׻5r׬�CF��ǚ E3�ok�����Yo-�!!@�R���|��vw.�<L1G�����2,b������~�<�Ǚv#����"⧾<�u-㬝�1T��R11�2Vg��l�J��S`;�h�XpS�a	���(�2卥ӭ��x��)e�Q,��0�B�����
1|��[�쮙V- 0���j2~Cy�>/����zP5Ã6�w���	(*!����5���x͓�Y�����,��{�� }:���3�)��:��l�RZ=��B�5OX
��7���U���^�aG)�&j��sz �I��@��� ��ፒ{��O���'+L#?��*�&�]�M�ER08[�꒿ %��|���SZ�H��D❬±�_����@��fv����"�f��Z�/PϹA�v7�u?y_yղ���X��M�h��#�W?��Ɇ Ұ���qp���Q�4�P�TN&� �@"%|�����+�R�0�R�N��dS��.3����0;�'LHn�!�	����NI�J3���r�K�鷕6���z�on �����~~�wR�
x�b�z���e� ���)K���"��pS��,���~��K����fZ���֜EAh�l�N0x����ޓB${��q�]ܚ�<Dmhg��fĕHtb�-Y�������HY�:��8��.ttԢ�_N+� E��قN�d��@S�o'M�y��E�������,��kU��}�0��k"`#w����$�|�S7+�_�C�'S���C�mh�^��Н �c���6;��_1�����R�p�۳��D�h�9[Sx�X���j��NB<Wc��V�(�6�呹<�'S�����п�Krx��%y^Y�0��N���P}(�s�ڈ���ܕV�D3*p��ьg�p&�U�x5*Y��`��M�<�,�4f�ә����;�,���9D�r�qI٪u�E����3�~�2h�0U8���Ւ�q[U�R���h&y��
,�!�t�FU���sYw���X�u`_�Ʊ	0����H7��9*�7�7I'V�X?$��Ή��Y}�ǊM�_��v��(.B��ς@��W� Ă���ةO�&�&̔
u`U��]`*��Q�2po]�x�[������q��J���X�"�<܄��b6�w�����J���]׍��vwݹ%|�sҗq�1���dC� ���Qv}�����WȔ�G���5�4��_
��0�b������ &�yBt�h�
ʷ�B�3�g�њx,���#�v���I�z��sՐG��ښ���-�b��*�����S�T� I*}��,�xfO
.9�m�7,/y)HT8h�a�{=#�
�֫�"�u�H�Y��P"��?�F�?�Nͩ����*�qˤ��P"'�s~��Ѐe{�W�ke�5ĳY�J�t�s;or97��u�	E4���?ڞZLNׁOt�ι�5�^X�j�k8�*$o����n�2y  Z�e>�*
����l����f�p�+w9?�&{y� o��l��<N�<�l����ӳThLG�Э^(��e�x��q����Pj�i%&�{ڸ�ZS�U��+^�D)ɑN��!�e�w��Yh΂�Go�"��J�������DS�frqY��h�p8��Ƈ+�؀ٰ4���	=.5	^���������=i�*�J�������)Zu8�[8QZ�n,���t^����w!ͩ�-6[K�f�Az<�Sިq)�1�����A������|�v~�tO8h�/�xt���-��~�$�x����%l%O��eU�p2���V} ��3�%S�|M�e��W��傡8�+�f����S�&TYOI�oe�؎^Z����Z��P��&l�y��͇�5��RB�)^�8�<&�l��%�&A���^��?���\���;�i"Z�͐&�lvS,�cE�m���頤��4zA���;��_�BD��X�B��(k#-��&-��QWu�#Ϸ�B� <��5v��U�D�nm�6��w�x��� �������v�e��(�dr����"s���JT��b�_�!ɀ�� ��PGF{Q�
ӗ_x�I��!+S�'φo�����V����I��uZ�h�3Ӟ�rH�,ϕ7�n7�~��?�� %�+�?�p�=�**�?�爛֌���{M�DY}�D��ɇ�jM9�8�{Zu��nrF
j�J9�]
�������X�Q�1�.��k�B��.6?A�@�����D�qn~C�>DZx��8�^�jo�^�@m�_y=��F��e'�Y��"���)��|��|В2`�����e��maY�k~}��6����|�G��m�'�[o]a���^�~��ٹ��W�S�b�� �TQ��/��*m���/6��6���j�Cm�	��F���mJ['�!���_)��c���eN�l6���H��[0�l�K\��6����?�g�t4�}��V��Ǻ�S����>���YJ9�uPP7����+j��Hׇ/�/�-���-��kK���;3��q��J�B"Ǧ���3��}agm����H�$HM\,T܎B�~ �;*�)�j:DU�����>�E�_U�������)��~�e���Y��N�+�k�@tD�f	\����ܣr��y��<Y8�k��#�`~���K�K�F(�`�?L�K%�-�T-p|���f�O1��AVO�io�M�s��~��R-�(�������ک��c�W�Dcy�ŔCTPAΣ^!�$V YM7d?aL-��K�� 9�x��_}F��/�ji��k���W����(��]e�W�:��DC��#+�"��n \����
�-
���.+?R���to�i9��j@Y��d��C��_�,�����9��>U��z⣨Ϡ6��چ�K�TS��p)m��U_���>,|����ޢg���)=���k�0e���J�vm����" �"<����gxx���~6��kx����x@�+b����4�0�����Ύ��9�dR�c�:�E���>!]�����uj'��g�Ly߿��{Zv��<�r�-�d4�?D�rҤ���S����Fݠ��<�~�Leyx7�^�"Q7���`-���.</�汽F�$����M�F�.�m ɘ�O-�4K��$�h��g��w������ƚ��e+�c�~��&u���@�h%�Ю�i�vM9-~e>;���2b¡��b쭜ЈE�<��[V��ô<�3Ã�)�D[��G�=eX�L�ۼ�d���o�h"����)�K@VS�j�jŬ����h?=��5�M]H�/Y�!S>Tv��PW�;����AwC�Q���NJl�u���N��f\+"� ����q¥���}���P��h���v��oΙ$�ƆF��@�_�@l����E)��=��JAfymK-z�6��}L��"f�~��z2��2�������K����1
�Y�p�#���<YV«U6���	��8����"��B������,�o
��T�R���x�x�5�S&�|���.*�t*~�2�x#,�r>_dz�7��k;�����SթƠ���b��V�'�h]'-ž2�oX�7�nF�b@=�ן�>�?Ƴ���?��-���{��&�˶�_e6ـ�ϣ��1
	���S�/,h,����m��~E��o����S�nH���/��TJ��|�}Z�+i��f����a���� �v�+����@i���3�7�����5��fo����~N���(Z��+s���qO�~�~#�"�3<`���ud�>̟d�jsy)nF�����<���=|���~р�u��b;����K�&x�}����E'E�,� :KԲ,[��h���<�;�h=�IB=�%���n�\�e�P��s�^`��y`|�����r6���0�\3��� /'�y�o?*� &Czlm����k됲"������w��]ߗ�sjXh6��l����%�Ĳse?r�W�L��`�^�'�v�Hg�i�	���y��C�O�!�t)�}$�k"�rAT�ݓ�68�!����۠1hPӇ�.�{PW�T��T��t�3T��F:SԐgEXo��"m�Q���)#�p��ʛ�,�0ZS��'~�]�E���૖�$w��X�/1�c�^��y+Oz��$�6��f^L��W��q�{j��I��'T�a���vEL��+�O�k���*@���,�U�g�V6�r�����s4y�B�}��TL������?�Q�-7ׁG��]޻LH��ۢ��6|�J�O4��r-S�3�ȣ*(���B6�v����˩�~�,�cJ�����˲��>Q�J�Hw�g��~G�j��ߨ�(|:(1�-v�P� �q&i�S(F*����?tA�P�7*@k�Q��u�햩�j�N�9������dk�y��s����ZX3
-=V$��щ���ɇY�)VX�Q��3Jح���
�P򒢈ݰ/��b8�j��������Em�9 )Մb�V�C�+^ܮ�4�
�-!s!�s?~Q���ǈ�.�Xh�{ ���;�GNw�\c��a��eU/z�f|�����\ZC?R���l�����g�?sg.h�N:���x�+�����Z"$@*�>��}7��z��U`/�l�t�)���^&�݅ױ �g��PR���͕��k/�A�����hj�V�V!�K��F���6)�ܴ.��ŕ��z�#�(lc}c�=ѭ{�Y�75QdFe�҇K���V?���k��g'J��߆�9�%�S�4�jgᬓ�>�Q/��_Ǥ��د2b�X���?���˂��O,#e�ʪ�ή��V58O��ԓ��p��7�F�:���
6��I�g,KMwr�3�@�f��A,y�K�IO*���^}��ix�C�M��֑%���ky�XÑ�t�$|�|q��� �&ꦛ���d�9�:dC�@8��N	���ǯ�0y�,E�B"25���$> �i��D�>�tJ\��/kS����:��?��f�+�w�5�{^ W��$H��Q��(��o�d���㦋�ć�W�=����)h�OL�3��HU�`�(%2F��gw@�(\^�'E����yY� ���^0Y,me���$��I�O��9�Zi��'.���E�{0�qɢ�N^`DJ�ovNI &�Wv�]�猠�.y<�u!�ݎ�E&�r��N���]���M���ћ$+��V�B��L�F�9�ű8}�ѦS�@�8�4H}r�p`�k��n��?>u���������KG��5z[�K�9ǔx���P���TJ��@˟T��?-z����9���d�۠�Ae�0喁�]1P�&�e���u�*��r��I'N���j��$T�AZ�/��r�^!�p�e�]qh¦Ӽ#Y0����]}��/�l�1�HӰd
�@U��Mt��B�z���L5룓*jm(���������{�R D���jr���(+l�]/� j���t�p��jTHiw����P C�^|c���˲�JÏ묠��0����9gC�UTF��]�g�1m>���c��@�n�oR�s��?�~&�6ÆVں��Q~�	E���a�鸳��b��t�A���,�#q=-�0�d���Q���^�������D�
����c�3"X�P ����)嬝����U|`p�I[t�����\��ؘe�u�B�i9ȡ[��+�\�z��e��X�=�>��HSY�.xV�>}^Y����L`S8��x�(�n��@ef9�ޣ`����3]��<��DY�Q	5�� �I
�'�9B[�'Q BjEʡ�ff,�T"|(V�5���CZ����t������;7�y���O�&P�?GC}��%�#�^�!&�U"Z?M�p��%�.~R �m��[-<BӬ���/g�֮\|L���tf�e/!�jr��a,�ʓ�h�Y��eX�M$�S f�i�
Z��(I^�sY_�C}�i������i{f$�Y��ζ��=�ց�T ���
�m�o�dF1�r�=O��YP�=��	�y�9��w0ބ�5�g�@5�[��.�W���k�I�|�_��dkZ�.��kӋ7nE�,+1z���������a�j���'��'�{AHPjEwK�:����҆Լ������--Q��:f,6N��)�&@rD_ �P#�acT�E���)��«�������ڏw�' /�'��Z/1K�j��������u�L��
��"���d?�Qk�� ��A��"�j�:��Cw�h�ቧK�n��L���{Gѡ�e�2_m�~2z1���@aVH����T9j�+�����y�Jf"���9�xo�*'~�X��M����-�C�ו ��#g����r���P�.�E��]�0���cl�b]E ���"������>��X5�9B��,R��օ�b��ηuvzՕ4��S����Zu�.�j�P�6"'���.��)��K���wMbWg#a�Y&�+���m�n�D;�_y��p��Bn/q�紃�{�?ν����pH-�&^b(a"y�K�,ܢ�"�C���[^a�5�آu��x��N_nV�>>����h���K�b��Y�F[a?C�{h"��x*���!�(��d:�4	��^��O�L�,:>�_,qF^E��,��������AmW��sx&�����g��_z�pg���[}��f��O<4X�֮O3�Q�i�K}[��%���K�q3,P)��f��/��t��U����'��m�צZ[�7�c���qjuO�I|=�`�rȨ��Gx̉ZL�v�6ϥ����<�&xWB���#��\���M���r���/�o�S�q��8d�����D��{�Egl�lO'�k]Ж �����nvםTb�!K��D�X�F�F�1i}��Kw'���c����M���wЃ�k�Q�~�d��Y^'��Qk0y��Eæ�!��h(]'�;ﰎ2����ۍ�l�^��?a���W%�]y��"�p�����M�nx����ה�*'}��GEd�ۯ�v�3 v���h/�Ȋ�h�⚢y��q�K��?�<h=��΁��X	~��yQ"H
@��%�R?ư��8}�v���w�^9������XmǷ�mQ�RF��9rgupb�q�L�Q���d/��ձf^d���73�[�`Y���}ࡴ-q��ޤ���Nw)ua\w�T��A��4��55/O�5�@�J��~�w�,���F �oONk7L&[de��\;��o�� ����sM�v��)�3q��� �Gz���ࢹ9���3�m��h����rǁE�i�ǆ꿊��j��E�4� }�X�P�8�"OŜ�Vi���&�I���2X/��u��W@��Y=��%�����H�^e�ǝ����(�\�����ht�T�c L�C�e�}���^��sf�K������D�<e��˿��{h"�hZ�n۝f-#��LI�8P��+9��xGGb���}���<��|��K�ɵŗ�Ƞ5��t�K���R��(�A��Yy>��r{�����>!��BkX�*&��l@޲`�*P��|�7�8t#���q�7���z~��l�T)��}%7s��:�ɌT�z1ϓ���Zp�����;kd)�;�bBk�Ȝ��YQ	�("�.���QR�-�W����~���n�,pRDW8�>�2H�\	����>ac�A���F�HDd��4�tR���B��ލ��ŭ��")�����M[��!�^2�m��������9E�����V�2�T�F�C+��Ýd�Z�D�:���w�=3�� zUh؞�]�50Ʒj/"y�K*��7����0��HK9w>� _�ȎH?��7P��'�f��$�sr�1RG�`�,����w���AH����D����{wώ����6=�9���ܪg���nAg�*QH���?�u�����f��
+�9���}̳���&4K>U_Z�.ߺ�_/eP�T������L�
���E�w�\�����r�%I0� �J��Щ@vg	��������1����z�����p粋H�u���,����1dމӿj���k1��}�D2@I[��S��������Գ���\���1_2�z����F5A�􁙎�M�F�����AuK)`��:���h��)���)}��z;�s�w�"�"�un��z��|����o����>��ދ |Yݔ�_�_�r18-����gP�� [� ��b��mH�e��B�	���}���0{T�#�L&�ګw0��-�BI
Ү*9�6{����{T�Ů}%OB��!/�����"	Q�B6bD�c�jj^�Q�ǆhͰ@@X�g��["�����g��֫�֣��^�*�5����߶�� "\4j�B~�r�K]bk4y�!�|��E`��s]��;0�竃2?������F�����͐�:SD^Sz��@��Bȵ��!kɼ֢��c8�+�y���'��.UˠrrU�T�*�MX�ޣ�R��u�i
	����$ޖG��l	olʴ\�V�L���n=�4���H�|%]�;1���L�_7��G�g��*#A0��0��Ǧ�2�1��Ѐ���߄]����H�t����;�xZ <W�6�ª3r!]�`e�!�"S����.k�-�/g$5�u4�N@�5�u�H�1��[؈ʸf�x�stp+�}�A64�Z�TA� ���;ePo|
gc���l�>�`J d!MsR�cߪ�[��ҕ�T��t�Ő[�|��GB�7��hքDjȂx�N�v�����h^��.wQ�x��S��?��2�������>KVm�n!<;�g"�(f�ȺN��HTK��?���Y��d9vnl�0��m ��s���)�W�Ů��D(?�Ԉ��c�x��-�Yx#��/�eY/�k���B=�͕w JOd���4�|�j���W�?�ù�}YWJ�&hF�04���EHXr�j�]UMܐw��$Lt���y=Ro�s�o�ũ�����%^A����F��Y��dP��J#��JE��w��/oؚ�zD���0;�$�����X��t��������gŉ��F툯����Vr�~�IY �Ώ촦K;��ޏ�$�4S�=(��n���3J�"����W���z�I�J��1�������%��.\5H|>�mzG�7>��至E �� N
K��(U8�&�#0��|B���6�$8��!w�yb���T%�K�PN�f?z�c
��(��/�'�Y4�dh�Fg����� ���jfu����N�y�,3/ ���OVx�� ��>���i�i�hv�Pl+E�}#}��Л s�HO�"�q}��)�0��O艖Ŋ?��1�܊t?���>��˼c|椂�n��,��ho��j�æ�/G9
���}�idG5O�I�D���_����`8k��] ��,�s?�P�>Z����!^sk��A�F}ڷ �|[1���4F���E�U�-d���V�-�K"�3F�ϸy��%@Sl��294�J�=d��Ű͒
�,��k������Qժt6Rl�`ts�B����Q���������Ji�Q����G�g�͏��;?x?��.� �">��#>k�)��4�ӷ=���	��mdP\��"��E!�+)\U�HS�	�_Q[���Ʋ�y-�uq�8�L�#���6W��(��ՏB� �΍$�]�9@�%֘݇tUJ�������	<f��^t���j{ gC��.�=�p�\.3�5��vq��M�k;��-����m&��9�`)s���/�ITP�(�SN�������]k�h�tG�<�D�_^��SnTJ���@T�ʚ	�b!e�uM�J�l�dl�X���p�A���{���qn��#�R�fܝ΅���R��OT�	�q�u~��Hq�������-oI�5��J�g?��sI�zJ��.�b!��2YS	��T�Z�<�4;�83n>'$�|5~ז�Pݹ*
�H��Rf����l��%��U��u�κ�s~�}\aFo�~2��[;+���W�5ѭ��)͹@�A�!惡��׽|���5�k<�UM��-�����˜�g�nE&��^J^�w�G|��Wr�Ws�����*@+��D x�G�m�^l�T��UQb�T=�nu
�i1�H�����P"��Ga�"!^|�:�N�! N�=c�p~Mϊkf}X�e�u�,��:#r��P�N�Vb�O �볫��t�X�t��4 w/����<�]�#��vO����޲��.� l3�p��H���|v�#y�Ct/� PnȒ�Y&�T{3��F���:� 2��]3��Z�������-���.�̴g"�}�n�a~|��$�:�
c/2���E���| H&.�E���t��P4��9�`�84Ʌ�I��n�*��K�D ��-q|q���j�Ȇ�����Np#Dfx�Za ���h�."]�׏
?X�5eJ�-؈��x�0�a��yc����_�M;�d�������ґ��P�h�x?e�� #`�lk�P�o�Oe�FLk(���7)!��:�$�4���-lA- JI�Q_�{|0����!�V;�w����S��sb����]��U�a�V#���/5��I��3s��%�~������b?�_�ҢMm��!r�ǖ���\��,�ɒ��s���u|��a,�c���q�3E�Q�n�PAM�,X��;�6p�2�`���[�bk����q~`P���V��}N#ꌯ���q�-ǏXu��r�V��3�}��y������GJ&H�>ن�X�9���P
�nÖD�:*-΋���3�z�heK�"���n�{��Ѫ��Y2N>�Ys�̉���<�������DL��ގ�����,�tl��$萐 `�����)�����>�K�'�G�uH��t��iXY��39���%�u����#!b�Y!a㲹���ƒ�8��޷�I��<ɪ����-����u��q�_;:���4�A����k1^b3E6/�(�������������Cݍ���I���G݁Q�wC��M���(��^���0�c\=��"@	x#�5�_�9�q��]J�/�����'Ra�
}��)<a��eI}�
T,�3޼Τ�� oN#�fqa�ғ�hj����AKb,".VC��eԈ!n�I��=��3J�,Uw��-��:�=�-����l���] �)���^�
��.�#΍����W�|i��~�.�g���ϡ��:	��mG�cUW�;���[���^t{������X�8p���f]�_H_8�K�Ȓ�<�9Sq�^�)oh�-��/HG�IcE���!�y@���{$w�,�1
�^>pU~�	uPn(�V��Bd(�*�	�B��Cp���Y������ܖW���>�h��K�)�0�mrl�ޅ˯a�M�_��M.sݮ���{�> �� �C>�dUHN��>0q�tGtֱ���L�و ����^�B� O�9a�?���?{C�F��?�M'���9��T�=�b����1�'<�.�S��eT�Y�o�#6�a�2�ձν��5Ffn�˴�*.���Ta3�{v+�k�]�Ʀ	��L(�"\�ӄT�TRB򜦈�m������n�����~�?k:��9|;��Q�׋4Tχt���*��	��xy��	 �Y�9z��!�Mۂ�|�ȝ��/��.m�N�m�$�pxw@��\��;��%y�٪�֋�@�+�qrG���-$�5�γ�|ɥ�7|��3T�������^���1����#.)o^~V�T�{���^�F����
`/�0���C!�I#��d(�3�^.%�s��#r`+uo�k��4(�u��9¬g'RE7�^���d��ݭ��A�4��f�?-u��Yp�F-���O!f/Qm�N(�˦��"�������/�.�!�VE-|���mXcF�5����&��}3,U7��\!$��	��n�5H��E)u�
��Mrf��ڋ��˅Ι�3��0�@�}���JcM=�-��M?�ʂg��RY9��D���BZ!�;����ye��@��_�v����*�2�7U O�E	�!��o��Ϯ���n)@�f��wc�߳��->)��*	�q߉F�h�����^�`��`z�@�GB�F>��H�/GJzK�93g�X�
4*&�2%!+����俈u�Ի޾׵��t^�j/,K�^6��%�W���'�ϋ����'�$�ˊ{�T@{K-��ޯ�z�@{���ܥb ��cc����O��8�V���GI���rχ���c;��.��<�F���6Z{JFgb%��Z��ќ�����v���D�dM���kq����ԧ-F��d8Ҋ��cc�b�������h
��G�� ��*�.�5ḡ9U'w��4�K�9b���AL·�S�8�������w30X��Na��\��%����^R�R�e{����t��#��������kH��h�f��%�ZJ�8�'��H��BJ-�O`*�)o�ٍ��,���T���n?�/;Wq��0c��Z��3���/JS [�_g2������h**,W~̌���*�	Mׯ1O�e�W]��e�^��w���,jO{�K�&���Ktu�Ra%Y�����G�mh���t�hdﵣ��e'c��X�k��߇�'��n >���{�D��L$���pp���"�Gxٵ�G��O+�/d��	����.T긷��[/�o���Vn�Br�jl!���/���[�H�,~2���_�����$z]A��� ���1;T�*F���J;���"�Yb;,�#7�]���C�~�+�KZ��`k�L� ¥�ܨ C��A��x���1-?�8�*�p]�KbЗ�~k��LͿK�6:�x�N�LU�!a8%�G�I�jd�i���acE���P�0>Ѵ^�馐[�2Z�a�F7�ȗY�Z��]vxS�E��$M4[�8%<��A����g���dP�¾��vN��g�7�M��M��y�nѴkW��T�z8���r�P@�)D���93p�6jwZ]����H�t��& �P�d��0�{@��x;�i��x����b���u\9Q�m���9l���f�B�}$S�̀�nM�^^9ZgP���� (��X�`�i=�#s�@�q(
b �4h�n�v.��Tt��������\�ZK��������\{ҍip��|w�~�+�B'8���e�(r����_��X��h+���R�m���$OL	Y�7�m���ʟ�( ��q��ۥ6�d&sKǕ�4e.6��5m/0..#v��'"��'��P��=�L&6:��b�L�2$1aGXY<�H6�f��H�oƆ"��`��~�d>�V�YC��ZQK� �J�f7�xF�A��#|�@}
���%��T1G_�}e?u�k8�ҝ�5R���<}[<t��������Ā�a	����-;���?�N^П����~�w!U�����]._�����i@�	��ߐ����n��!�	*7Ua��8��W>O������VzB����:�2#j��3�\�@L~�>��o�I-��%��4��Q<]�2틇�T���h�D�˰_���_���È@��Vy�|[n�zQ�rX�JEY�u�A��! V��9>&|)��2��z<��gq��4�����#qe&-c��5���tH�=��NN;�f$NYK���;c- �~��������	Alji�ki�(F����G5��i�6�`1�U��[�ĕJ_�T#��}�m=��w"8an�S�E2��ڕ|��H5e��	�;+X�MM������Sp�\2	@�ѳ;��t��%=���A�S 5+���
�
�>R}�G�C�{v�TbLҾ(����!�d����o_�F�L�b#0�a��^�\M�\[-b	�3IK��k��@R� T�R�p�*�d&X�
@�Dl0��^�u�2�V!?)t����J�;��%�l�����^�,��j:�S���/W��;V�IΧ�����L}8��KWDZ�jCZ��j��;7(��I��ד�?��+�cO���� �m��~���а9T�UrӃ+�k�46�юiE0�b_A���;�+$!�h�o��L��H<(��o�3$9�S���sJqޤz�>z����Ǹ�B�8F��AmZ�[̿D:�a}>�Q���
�pe�&����AB|"���B�����4��˜����n-� ����+0=�ҁ��\k[z .�b��Iwh���o� �@j���čmH_�^��ф����ND���(������\��3&~`N��A�x4HؐgPp����ؕ��㳺�)_�ƥEY�LW>G�C���ł�65���+k��_�8їJc(�ұ�NÒ,R�\��m��+���=Mfm�\N�T�IEu��iZ s����K��矬YE��>#��2����#��)�����!b��U���/�Fk*�$'^;�g��R2���P�����Bޠ"{����	�śkN��ow�Dr�2��h��@$o	�\ɡa_��A�ֻ��T_��̯}gM�R<�u��ٔ�4�<�_����!gJ�K������P+ ����h�}�fZ�_���$5ts�����r�}�:Z�+�z�=<lJ�F�Zy[uV�?5���e;5(߃�3��{-<��̏��]I����p��]c�0"�h7߳�k����)���>�*�"���=s�IM5"�5���W.�C˃؀�#������gK:��y�ۂ|!8jUx�j����8�Ysb����ʭL>.(����zG4��0�l_`���e�!lۨo}N��	Bi�����o�6���-��Ċߒ���հې���S���C�yҔQ�\3|�f$�
_��ץ"�e�y�3��D�z��f'�/H&���o�Q�%KU���󹝸�=��'!OL]}��,
�Y�6� �F�	%�h�ZWЭj�KyC����ڔ���ґ�����f�����l%��8M��YIr$3�0Tk��3��@���K�}<(�������2�C��<A/���+_��"�0���I������%s���nM��R3�%�KI�u&�9���^mz\�9dk#g�ק+{q�b��-������������#��K��r���9�U̴�p#EY}+�^L'}��do�7����iZ�?���ajg�ɇͲ���W����$�'�dmr���R���A��u��'!�uw��	�k8���|���-ߒ��)�/�Հ�o.��DA�K������_�' !�j
Z{I���P�1@9�:9�{҈[���P��xF�������<�c�����4&��x���ܕ��ft�i����_�.�:#,��Dc#I�4�����p�<�H�w�oLg�M��f�� �~Ȏ�P�֡n +�Դ
��;�����&sX�{
�])��r���p�#�����Vy�5�F��i�fb��V��R��
v'�p��y�~xY�s��͒��^�743�{&�&��>�����g�2;�%�2�|�U�_��l�uU�����TƳ�|3��XV�.U}F��.ǁSLb��3ߍ���z,շ7�Ռ'S�zxG�;#:)"(�#wb>��G���c�J5�����6��/'��y�fקj��5�$"��w��Jee�(�d�^�U��CF�4ރ4ʫ���@���:��R���+5����D&�I�-8��OC�ޫ'-�!B�/yV��\�<�[?K:y��sRV7F7��*/;���1��J_Un\	�>Mz��^�am���)*x��
�x`��ٳ����N���7#�Q)R�wo���D��*)�����%�� ��3��Ť�Џ;��O��e�~o�q@r�%{LDwB+S�dMQ)9�<���"[U�*!�PQY�����7f�\E��y)� �NbCE�
G�vM
u�h�%0f<.�݃h��RZ��[��L��m�A�7V�$6r�V^c 2��ֱ�������Mq�y������;�Q����8����j�ݚ�G�}-��~��;�&�.JP`�$����닔/> ���p�Cm� �H�	��E����OiJ�j����L�ޥC�EC������d�'���ys����Z+14��j-�����>Ǎ�<���%�B�q\�2U}R�Wf|;��g�o�x��V	��gZ�T�Y��ZB������2��x Wq��0���m�qU�:������&?�$7Nk��C�p�*�씛f.���JE���:�>�e� e��t�8�%�T��D��=��`��ŧ~�٢�����~`[��oeD�6�\��n�]�vW]vT�M�]�-������{1��|�K��`��7�H^	6�|Vjj!�����R�*���W$�4����Q��|&E)�b�L�*�Ql}hH�Ըv�rZ�F�ϙ��1>��AJ�1����V7,P"I6uRL����ki��:c�d�v�z�a<�Z_dהvOqJj�h����K��:@�#��/6^j�.g�Pr�ӍԬ��}[C�Z�n�m�w-�\�7��Wl��۹X{�)E*�3� ������:�@Ѫ��ȝy{^k�R�U��M�A����K�3uj�N����x1T��_A�X9a���⣘��b~5���`3&^�Dh4�Xu��]T�t[���j�@�Ͽo�du/ g�����䂙q{n7y���<$�,��&�����H W����"���ܼ4�B�nӾb,�9�=C�1LR��Re���S���E .e
r�ɋ���ȷaL�7̦��I��g��o5)	�4�$_.�L����:�9��,+x��M�D�ens�Z�/R��w.��1{��YE�JY���|���,h�|9
g�`��vGa'+;�v^��RX�p�BmO��+|"
�*^��{"�~ӣh¢!�9����&A��W��fp�}=��k�5O�~^Ne�'Sh+�M����j��Q�X(�kAa��{����K����?�w��cAe��!�#���sc㲾��7��h<��I�j7(���%\�Y-��a@D���T���*�-�(���P��z�K�:�-F5��;���\�-�`|���pߌ�p>���BX���������Zae��(Zb!�*\Jl9�	S�� �P�f�'��#<��^|C�S��pݷȑ	�"/��8������-��q,�(DlIΕ�n�R#�w��(й�����~�/�k
��ҽ�V�s��s��Y��z�v�v���P��w%�F��^��<���&U3�D�l»�^���xo�=x�ڴ2�d���(�a>I�Ct���-;j���C�\ �[8�|�+�t� tP�A��U�}�8�-�/��u��>�C��y���jˎ�^:�>�aE5�,hj=��ϞM����ӏQ��=���,���N��'w�9Mԫ,��5��'�/0"8�?4�V��-�Ћ$�*����8m��0G_hk�/V�������z3p����c鷻��g�C���)��A3@9��,�8<�o���6��	|�g�b�>��w�6�X��uJ��D|���U��D[��S��G+c%d6�Tg5���pl.*���5_��@���c�����G�u��g/�	?Gr-�=��6�Q23�Ш��� ������Y7c���/x��a�v���g3�f�%NxSBC���u��9h�W��\�1ꏳ����g�j���#��� �A��7:�L
����G�_�N�W�TW�!�2ͺ��z9'�'��k�H��!��*�=�qA��HQ.[��'Z��#3�*����\x�%�]�J���Ѩ���@��?,53S �3-�Y�0�n���>�-�K,_,m�y�����{�+ERo��Tꔔ�����{,$cs��؄^ΊB<c�!������37�Z����
+�/�&�B{.Z �9M]�J�:�L�_ ��fO��5���
|mճq8��10q�Aܥ���XT8o(��&Ҫ;Τ j~�Z:[5D�#�B����`�6u�&�G49򇭠�������tL���8���Jg�PQl6BK�=���ĦY k#$��X$ܯ�e���F��=���Huai�8#puV(��	�5Н�<P��������B�'������1j#I$Nm"[���c�w0�d��&s	@V�l�V/d!��S�{U0�\�˳U�t'����D]����qL��%���WΨ˼=�ƪ�>�N ����Fc��Fu7���������0����d�av�FX��o�^Q��R����|�����������|�ږ�k�w]�x�Ҽ�� �P�kqF}���
�N��� �C���<SS�94>Ws�1��(�K�����DjB���YH ے����!' �#�����ݎ�鷰>�vH�S�tp����C��h.ku�o���&��ΰ��CnF;�7U����D��N�9x9��;�1�M��c:GZ5���i���9"W�����y�f{n����qb�D)��~T[��/q�y��]�Տ��V�+̞�\���w|5/�)���A��!���Z1Y7��\ĮT3����W~e5��	|�Ue�Gm��1�j!Ghw�lv�%2��׾ML�o���/#TD"��3���
�8��(��3��=�큘##ō3����¶���$So>N�!h��5����1��4�B>�hV�&�h�ˍ[�It�Ǜ����	�;]�.�d}�]�2�M_��.R�Hh��� �>�Iqy�xEݡ�|I_�Ț�26�������@SqM��71Z}�iR�9S�Ńv
��6�=�!�J݉nJ;_w�M7��r�*a�*��~r})�-H�hsg A5*�d�G���ۺ��z�텇ٞY�����Y,ZH��=�?�3]��Ɩ��7)�4qiE㙺	����K��4_F�˸Tl�0v��h#�n�a9�%�_�`5�������3j*�G�\Vä����g��맳��9{5�4T�c(��Zq�bz[� ���S�'X&�҂m�u�?'\H{>C��~�g3F m�<�(!X�(�J�%dW�R-�����(t���WΈf�}�x2I�w���R��(XNb9�I�;W�0�BX��%[%0--"�Vx@U�?���_�������{~a�aVX�[�`�pZ`K�c�������lC�����m �?���xUB���H�GV^����tgw9��|�<c$7����]8�*�	�2�W��-�Xg39�ID�7��I��xcy�N�W
qL�r���R#��p~�����x�����Hm%\tL�d�9�5m����^��y�=�g��SKc���o�N|ӑ���"����ran
!#����r"����1�QS�,?b�6�0��H[�����c�CI���r�5iY�b�.؞E�}�B|b%����]Fc�tu f��Q���(�Id�Ov3�����=�`�a��:�Ւ�e}�+pq�	%/nL|�ɛ��XeU%�	�Rur���w�E��x����e����"��d�Ap�W��rų�x��h���[�,�Iʄ@���9J���K �YRn�a\r�G�v,�L�䛱QX4�Iʑ�aK�ѱ}9��u�>����F��W¦�T����t3���ROڽ��q_�wW���"���gl�����ˎ	D5T=MjY��|��5r�ſ�z�.�#�#�B49A�����Ӟ�V_�s����8���jM,
	d5����Lk���wj�宐�t�ofs�oF",1�\1a�,�
j������������9e-z�TI�6(MF`.���J�\���.7� �
 JH,�0�:	PK5ŭ_X��W%l����g�˲e)�n�.,RE,2�c��FC���'N��9��|�����9�'��[Ng�L�Y��ZuUb���W"ݫ��"+��\�"���=��B�~]���B�w����u���`W����`��
p]:-��F,���'��g*-��a��"e �G����w.R:�l)3kABE���]rҤإt���P
JZi�!4����1�g��I�����5ʆ2'4Xz�+�|d��L+ɢ���dX���k TBH�ENE*錱���H5��!��&iR�n� Wڰn��у���i.vUt-�� l��~Ʃ�Z�Z��L�s�-��Ƙ|��cF�A?��V���#5���QXr����6^\Ey��⽱�@����M�W�����=��7���>�/��������6m|d���ֳT����[R��	�ύ�Щuaۘ��?� � �l�6\[.�~!u�m�@�E	�ra��\���Gr�3�Ȣ�~�!o#�1���>��V�C��NY]���]Z��9���Pg��<L5���T�_��F�Ʒ����ܫ��;T;�e�zB�BA����f���a[��JI�H�"����P��� ��(�a�Y���H�/��CY;��`
�_}0�B;Y�lZu���_�Gjٱ�0g�����}T��`��A�)�F<o��ec�bNR�ctr���3�o��u�z�t�]<c�0���}����
!)�II�3��rՌiKyB�6A��dD�-#o�t�&I>t8rF�`��7���4�-��nb�@ ��E���CZg.Z���f��?��wr���
��z*��"w��u4|>�󣸫�ofF�¿Ǉ�iCȤ��t����K�n#�ne�4��kc��6I:E.�}o���cL㬋�P�:'}IX��"��x��|�h]������MŅ����W�Ɇ�'�F�:,�p�h���,�p��!��cNM���ލ/"[б�A�1��q"+�R�<����Q�ם��Pz4���^�Ğ�/B0���;��%j�}K1U����+�;p�'�t��me��X���d��|{�Q����Z�����rk������4W�J�γ�%� ��=�����ܣ��@���`#���v��LD<�An�1����ub��MױB������a���6�� �ΧS�4LU�JѸv���\�L5jŁ;��bo�;Ŗ��	Vy���l����aerH�x��S�E��h�� �a�D�eg���k�c���2�7�d��\�������^H�Y��y<#�#�}N�C�����������k07�3ȱqA<��ʏn8H����wȏ��eݪ����8���ɵi�6���^Pu���m��X2|����y
���6���_�da³����]��3g���4�"���A_%������Z!+�v�]��!����vND��˪�PH�*�׎�lH�(���H�$���d�2�ȭ�g_!U�n���<i��;�Ig���OY,�ջ"h���;(�	�1#[�|#��@�D}����yUȗ8<��l0����;��FU/$հ��=č9l������5f]:����޾H�!�aE�) ��������lt�k+���'�L����!ˆ�<@P���.���3����BB�w��J��ee�a����ʴW����2yj�uo�[lX<�B��]j���;a]ޥ�u��$|�̉�fXa��!{C�RB�q����m��J�;���-Bq�r�K�� ��"����>O슂*�:�j�f�ᗟ�]ͱ��"/��)��Z~*x΢��(R~b賳T�RK���Xϖn]��lR�N�4��Yk��%��z�&,x��8�
s�����EG�L�{D���by��-}��> ��VN�yy~O���-�8�L;�����񉈩����A�T����Q���k���$tW�-J�3Q�k�N�V���t�eږ�10�4���I��n$�����O,�C��w����v�;%�ۚX��ẕ����*#�Αʇ����=�M���Q��|
m���wE�#`��e4Hz(���Y5�I�� �&bIuhtN��e4�����,�榏�S3<����`�}�g�]<V}4���$� ٵv�2���������a�A�����6�7�1t�]��Bk�*��JQ��)���a�|��2�������#r�MY�J_	d�ݬ7Ȝ9���]�`�V�͔��;�W�圥�G���"�A����oTA����4������� ?`���xD�?�x6�	F��Ɯ�Q�Oص/Z�*c�r�Z��/�\?Z��s�n�'3E�GG�KOށ���-��8ԦpqI޹�
���K>��5e�uzC�ŒH�L�`�P��iS��L1�����=֣�e��}d���_K�%w�5'Ps�\2g�׾L����lRֲ\��>h�,ZG�F�Y����/����؝�:_I@Z�E�?x�uSLeQ��-��댌��!k����9O��!��<�����|��Jr�t���H��M&��Wn&rgaBs�@v����@�e��QR��s|��}�㧋��8l�U2�l��/Q=]i����{���1�t�6�������)<3����"�V>U`���	Y�;Y4h��ެ	R��,�P��F�Lm�4M�0�3IA��Z��ע4���U?8���M@4��/��������(��2�HdD�3u)Ȏ���k�#0qŒ����rM?�:���
���%���b������?_�'�o��)�4���}�%�+�k�;��el��`��3��x@��ӫ�P�l�T� wV���j_lJ�v��Y;����?�Q3g�qOջ�/r�w���./=Ǿ��E�m��RZ@�c-���`yF��Z�o��|x����}՛
�]U%���![&�7JbN�6j%��!���BJoI�ʀc��\���Y��5a�>H3�<���Q\�49����=fV�7et>�جNV��<&�í�C vM
$��������x9q����\��]��4ݭpO��/i�|���2ó��Xe�-D��m+}���l|�ho�X��]d⬂,��hӓ����/8x�&�^K_�׽�<�A���F@�b�?����<I��l`�_"Mg�J&���It��'�1�������K%��2�4ӖR���,���k�x�{k�>��xbYBE���<�l]=��[sI�������	�]QkG.Ziإ�V��o�My9㕤�����~&��T_(��]�6���9����G'� ����
_��[K�Ѝ��d��t������P*�V�K	=�8w�,I�{�4�&Z�},$�����T�����H�~AHΦ�Wa�y��T�nI��W�m�K(v�� j��������f3__PЧ!;L�@|��4q�2ːP�����!�d;[w8��à��I�1��O*�?ÕEio�D��aKp��?��k��E��W8�1��[3k6��b�����H��)��Y�|����
#��owp>��Tm!@�h�����U�U�:TE� CL��a�`.X�V�a��o��݇�f)��b W�(F*�����t�y���3ӫN���}�F� ��"��<m�k.�{�{�c���
�����82"Qڕ�+ٝ౉
m����j!���z�O8t�z.��Q�k��=E~f�D��X�e��؞Gj`B�7H`Q8������v8j;����f�a�@s�I�b�#��*�7m�zL�5���އO,n�� c�Rw3F�%�v�2m!.�}���j�d�z"��b�j/������mX�o�؁Ή$��_	W�)=��sn�.$Lpe�"O�F�t7Ha+|dI�j��0U�0�d< Q�%}D-C$#��}�ه�=Ǔe�+$	K: �p�͋<x��-T����F񎍌3��]t
���~�*����/���UB�p��������i�dʿ�� jz�K�H�[�|�k��XXC\�-�>�� A%��7}��҂{��̺��RI��2�Ŏc7ީ���nvYP��@���x�ӿ$��-�u�,~��|��3,��
xV��\п�tSmQ4�z�V��!E�n�w����+3@��v�n�tZ�2�Y��;[~#]m��J�7�\��m��
P�����%5�����U����0=��1�����E��2�1	�&�Lm�%[.4�%uhu�z2��f%��x�0ν=Qpt������_>��d� ���|R������e�����@����3+��H�(C!��\Y�d�m--,��Q�ۭ˖q%�*3���<��"+��m1�tN�Ç�ji�7��c�J+"K��`f�݃.U� ˏMCq��4d��aȽ� -	Em}�e�����F��p@�޴�%���`/T���ʡЏ3���F��=�_�(�;ع&�p���=�ʂ3�~A�-s��0�yOӆ`�&�rI���r\W���D~���A�GwB��L�a���e4E��)I��55"���GH?�1��:�����Pױ�)R��hdko)�_ns�m�z�+��T9��
Q�G�a_�G�]굁��ĮmD������)_��vI�R��_�Ia�d���:�.h{S�2�e�1��4�\v��E�P~�\�M
@O(g���F��J�(}|�4g�j�@���~fBT`�E�(�i[�.(V�gt�?S�h�,���?`�C�����<?p%�3u�1�ҧg���8�	��7�2s8��	p{�p�-'�ߞূj�/aZ��r���[Ol���gc6�����k
��rծ���vyن�=�U�!�q@�=x�и^���m[�&�W)�`��m���O���J�FН���%�{�C���Y��"�)��D#�Fq�yD		E��is��젇�������L��\I�%���m,/���=��q�J���-Ӡ4��( �?��$ :�����o��<dis��Fn��z�δ���Q��f�"<Tv-w��J��΃���dع���>F?_���� \c"��2Jm-���pz���*�
�r�+6�d�H�G��0/�j�	��Z=#��3w �#���jw�ԯ���������ܓg�.Kj�VS>��$��E��U��iJ�&�	�?l���+���$���Qx�(V��:%PH�@�0P��Ŧ����^R_fy;Ku)@F�b�+c��)��.}��&T}n=�`QA+Q�!w�_�gSp���	�����+>Y	�G���1�v�8d��|�@����%�%�f�ra%]�=��ȏHۅ���� ���!<���U�,���M�M���8F��
'�gm��1�<ӽ@wR/]�T�Bǜ�\5�r0��@�C7�W�� �x��ھ.��ǽ�d�ؐZ1���k9^�{b�ۃ�E*����"k�K��#��uzЀ�81lo�ug�B���#�W���^H���AQZ��B�W��ڻ������i�ӡ���+����(T	>�Q�8��D}����p�NL�|� �Ţ�5�gwvhMF��5�ݪ6������O
���C] '������ �����?5^&(S���'Jƻ�������í��T�&��48����!ٹ�UA��|�'=k?����+�x���+��"7E_=7wCT���hLա�j���6�K�M��K<�Ӫ:3S5�C���Yq.d������Rk��!�����X{�`�	7H��j�h{��+�vUe�I`v�Zi>�,RM(��d���� ����OԜn}D�S�uL*�)9n~P�VC�~GHh�ͦ9�n@�F��c4Z��V�ռܸ�/C(n��!`u'7��-���$8,G��]�VKq��կ�EZ�	��|-�l�R��
��#O.�ILZ8�~�]��zQ��V�4��W�/_����(-�J8�G�
��I.!�2���chrm��E�[��F�����;v��M/�AU±3Z�y�/���� �c�=�*�p�ˉT6H��j��E�Z�w����#j���Mn(�+���1bp��;XiZ�Qd~Z�Th�gi��&���c�TX�/��zR�sƮ��)��������+;Xŵ;�r5M�*��?¶�}H�[ס����R	v�o(��"�_���.�;ј�C�>��ӁO�P�4����+�ܚ8G��pA׍�W�3�U�R�����)`;Rux?���u�98*-v�����/'���U��� ��:�|�R �����#�h�iD��cVj��7�U��x"��}I�<hF,�����;��Ί~3 k=a�/>�g�G��q�3��4����\ ����BB��
�"}V�q�Z��x7�����O>�y�SA�1�b��5G��!4뵢j���	lv@o�0��ίκ	�Y(e-{��o��K̓4�zWc�7��'] B��h�]6��+�QQ:E��d�5���1��wŨ #��������3��/0*9t��j���|_[�P�d%�^��qA���'�^�N2���+�{xc�):������2�s�О���g���s�g��$�1n����m�
�'��-F���N��ފ`�-���Xп�Q����N��;P�.��8�5T&���s�ޓ�����X�������z���2	�x�Y�T�ǔ��CBr~B";��*5���x�h���4�ʲy���{�Al�NzVi�rnQ�'�Z��~a�0���)�S���[�)b��M+�͓A$��B�0�G�mA|�%�����(�j�=.?�j��Sq9��{��W�ܓw���ϟq ��!��u��a�A���v��a��H�+bn�=蕣�	B����]�F�w������T����ث2��90$��W"��J�bo�a�(�{�'����Q�Q�%Ya�K��a���\d�ؘ�Vj?��y�G	a�Q}��S��1i����=T��X
/Ժ	�4�{]�S�1��Y/5�7U)+���ZǺ+�bn��@Mb��?��G���:���h̎L�Lo�f
���.�{Н���e͇F��Qj-B���gN�Ӛ4"֕`����;1�͉@77�-0SUت(�� 	OIܿ��ӠJ��츣{Z*)vu%n���>N2�
jb�
����?/��9\D������8kj�1��U���ZJ?�hN=�XT�Z.�,�Pש,�0�-U��R��?O��G�v"d�0��i��:���!X��ø�FοQ�~Z��� �r+�,!�z��m�S٬�}��ʼ?�ۅľ�*�W���N�a�ƃ�����Ȓ�Q��'_^s��'�UŎ��P\�M�6�Kb�l�:Y����	c2J�m*������7KKK��&-�s9�{����hJWj��G�5'���q_pL����� ��
]�m֛<��y������[,ߞp�r��|G �zOSTV	L��bz��(�hq=��;�
^"(��Z�?8�A؛��'�a>�Z8MP���T
T�]���F�����t�Υ�p�X	W�G��G`��9fy�&�b�����W�f�u��k-���[�ͅt��˦��R��m&��?�<���FdEYU�l�����1�F��r�@��־�%PGɋ�Ox���D���/T�kҊ���s���}!xq?���3�ߪ������qD�w�jsxPf��m��A�k��N��$� ���^6Ti#�۞��:i����D���	���9��苢���}0�l���3�����%g&�jO!�ubgW
�A��;�eݕc��);e\�n�����[� ���������0��=����D��?&�S�n���I.X8��~M�YL3��������l�� ��;i�4V$�0�T��~�Q�6��Z5 �r�1W��Aэ^�|Vq���u1ڀlr�^�����p�f��EP���'�B�ѩH�i�//��E(�ߑa�μ�Mv�J�������)z3�\{yYӫ�����,R�䙞t��0C��uмQ]��,��1ˬ_��/:��F�
x &�W�ڌEt	P#)]:wRA�Dq����A3��u�%/���z1�U�֙���ȇ��v!t���rz���ԯ���_8�Sfq�F��0�h��_R�z���*�6"x��nP��R�rD�}c�����A|�AHn�͋a>)��NOϻ��P^J�tLhLY��P῱������� cV^jW�3U�=;��C���r��/L��f/[�D^cխG�߇P��w3�C�<��?���w�n�5�[�˗�B�짗�3�8�R�{��s��|l�L0`M�*5~���J��q�*��՞ͼVL?k 3&�G��q+^AJA#T�������I3���~��PN �ɢ[�Z�%zO�(,�#�CŹ�(�l]�֍��Xb+�'�kOK�9���8���_s輋-G_�,,=L[	�)��\ d����R��G��q�����N�^2L�ǔ�q�@_L���d����rTwyG5��}��r�����R^�;a�e_���l�Xg�-�N>�N =J��������\x:SH�q4��03��
�#�v��u�^��b��M%�(��oQ���`��7תv�x��� �Q��A,��0�b�5�*�i��4��aHH�@ڐ�.l(<��3��~J��˻a�` �J��'�"���0ԽsG<W����+ܡ��W=8ѕV^i7$� ��`�芆��rW�����$oڤ��D7�*a�A�*A����_/�\��rJ&���"���ݲ�τ���VQF�*��<b�KOfz���O��!��d)�V�LX�R	����P 0���<��� x�ٛ�/YDi&����/�J�V��/��,�X��%j�x=�pR������/\����UOJT����{^і�#/]����MqAR�j�PI�4���$���.��X���TDy2���#���RTb��0 �����Ll����w�8���sR=�3$�g�2�x�'�"k���m�_z�"��̘���Ƿ��U��bfb���`f-g�V�s�SW]��u��@<!s���W�_'���Z��r|�tQ.9af���k{*�w#}3��$Ci��
�{p{0d~� ��.���0?�Ֆk��
b�u�hG	oo�=���1sA!2�d��,���P&���u���tE���ۊ��H��N?ڋ����B��	�c-�[c�n�~�k�}?�B��D�N:"JJL!��3�e����2���=Eg;*�����`臸9�&�9��}���4�:L�	$��D�x�X���X�>X���q�;vMԔ�u��W�V��`d�'SxO�c/�;&�W(ly�.�>J17�g��T]�"4��ʠ7�rb�R������yɪL�;��	�#j�-Nc[�\�3�I�1>Û�t��dO9��i���de��:W3-��c*D��.n�!M�>��7Yn6`��犆@#��ʔ�5��Ծj�D�����*���ܤs0�T�(�}8�]7{�V����3x�4�%G��3��K���VdJڣ� d�눤ld���!�_�Y!��
�d$"J�i�uSC6�{]N'T.���?�˷0t��Ny3�����A��67��<	_��Z�� ig�|���2W�G�_��6�=Q����5���R�9n�B��VJ���������@��;��/J��\FuA��+C�o.�Bf��R�������S���i�NJ%����Ա:M�g\�e�B��K.(����>l��&�&e���F{�M��s�7^��׌Xb5m�����QiV.��`X�vő���Y) ���R(Ϟ(6~�pvm4�E�
?!�ڭ|�_��>#[���P&���N��d��I
X+i�I�bۃ�d�_�*�y	��:}�~\]��X	�9� g1�4^�cM哢s�ĩ�A"x�l�����1淂dp�_TWG㏾?�t�ܹ��*��.e�*eҝP��,�kUY�o� 6H�E�j<�S�B�6�	r��Z���J�"�Q�	�ް��8�u��ok�J��ꊐ��yII<��jeT���^�^-4zc��Z��3crw�G���">h���RvB� ����Z���+�?�atTsH������+0��\��=(�s��,J���Y.�\�.Gzμ��D�?���=Km,�N{��	Thye�Έ;�Ǖl *{�>˳NU��O��4�l��עjs���x\'���E����yV���;�O~a�o����ި�ʍ�>V*h� Q�h]��&�Δz=#�-��~��i>����1 ��2;�f�K��c��W~�RU��tI>��6i�����L������u$D��N����@��t���d$A��[*L-ڀ0�u�u�e dt���c���ta��Q���cJ��Q��J��0\q�����ZT�dƝ����B�Ł-B�u�����r�C|�j�g��"2��g�͇���!��@�q���h�9+Ws�	����˓޼�*1+�~r���!�}�/���*��f3zd}y���� �v���@��M⪯���d\���Fv�9'F�����$�	�|���c�]���r�Yt�_��)���f�2�8��{!�l���S��"Z2E���)*?z<ڄ�X@j`n[,�=#���V�z����}����vhac!���k{�+���h��)y�D^���r+(`�^~�N�A1~?p�_�L�����Ϗ�3��+�(�z�'&�ȵ��]��g�߲�������Hr��i�\�Wĉ��}(p\轉#5e��l�m�5�t�D"C��?�����}q�Z�V�K�\����9��ؖ��;y��kJ-?և^ÔK����1(ȸ��'��_yb<3��|�̾!ޤ �Ggd�U� sE��e,��SVz�=d����>�v���,�C��(ʛi���[�b�_�w���_��m�䵼�����.�����J�U�?Z�c+
N:�_F�E��fIj�%ub�������t)QG����k#�r�o���*��e��
�� M[�(OKz���)���T'Ad�V5X
ϣ��愁��Y�t���z8��9%�u�����L��z4�+o	�v4�S�(;tWl����X kV�(aX;���/P�p�1, ![�5�	_�6]�XN颮��Z[|�Џ����U�89}�X�*���ә*�E�0Tl~�E#,>�+!�NW���jx��W��&�b�t4�9fd�W��9�tE3@�9y�]��h"gFU��� P���v<�����nn�̈́�[C.Y)˞�E��1�_�1��Q�����b��5���{�} |0��պ���B�ѻ�|l:ܳ���ל&�M�d��l!p����0�6��kra��:f{����[N���{g�BeHњ��, �ԯ��Ѳ�)�z���m���ݼ�KR�L� �"��I�!s�EWC��\OB���H;��]..Ur��M֪�݅ę�kOϛ�p���l�V��{�� ��ʩ��lY\q��b�{��zM�u$*} ���q�֒лb/��Ȫ:��'�@d�1ާ��Gu���I[��h=_BP|�%�?f�*4�(��(�N����|D(z9�;gN~ *�~O��=�j���՝K�d��˿����Cݔ=��OE���U!��LCC��ӃQ@�f{��FU������vK� Z%���b<�˺��8�;�~9�	;�x�'���3�/��V m[��B�I���B�U�Nhs�&�n���YA%#�(��`"{3�Ay/�����a��H���)�Y�Q�h-���☑��V��� g�1��r=c�/S�Ԥ����8�b�X(��m��M͡cO�hRZ5�]U*�#�P�<�I�$@	ˇzgp�6A���AK8��i���$�_,A3�|�h�fB�_���'�f�KK�B���=�A"R2�F�elb ԩ�	݂�d��/qL3�!��NR�d�O�c!6I/1-NP^}���r��&�Clnp��)��1A�'W�� u�m���)��s��j�|���x�d�D6�p��VPh�b�yf⋂��N^�ƭ=Y-�?
�n/f�[:+��Jѫ�TWq�����Q�iM��QW�|Ŀ�x��ɑ�#��B��T�k	d1;��D�珮��'�`:=����^��VQ���E�g%���h�Ɇ5�F�KcP�Q�~��37I��/-q�.���>"{��28��+�S���i�N�H>��Pj��Je�JOQ?�_Q��Ztoob=��$?�1�o*�}�;+<c��Г��l��ԁJ�����FD(�+[,���^�`N���J�I���S�sDel��E!�΋ȟI��'�E��y`��܂LTB�4�d*kVq4Ad�[Ɯ�up:�_�3�{�ٟ)��ZY�Y&��wg@1t��CEe�� ��b�^�@ ���#!{ew^��w��ዖk��I�!&7Z��OE��;����b@>���"|�$ηu)�?�H!q����>�PYI&��e7��9�����lY�/���Q -�C�d��j����v̉$�v�e��7��R����+�L������u	��[S�p+����M��v�y�k�
	ЃGE�:X�G���Î[g<��= n��-�l�	�:�@@!��),�SPQ��h�ܠ�~����U����HM�.��x�bW�Ra���H�7��;!3F����7��<�;����v�ֳ�n		_�:�'�.���b����ZYB��)��PK*A��G�9��*ǰ+W�v�f[�C���6gx�w��i������zV�p&AC�[W��f�d������
�-�TDV$3c�Г�N�8�o���f��!&� )�������7/"��!V�~y�(�O�oSZ��i��=��C�O�Q�Pt�l����L��m�LC�X,z�r� �1	Խ�b0�и�T-Ío��=�]����&�T�*&�������M���O������]��_#�%Fc�����P����w���9�I��UZV��x��>t��OO|�j���п�l V���&[�1x�q3��<J`-��}lсX�����圉��^���mtQd�S��
C�� $+����8c�bR��VpmS��OQ(��g#խ�6�����E���n��r
З�e{���sW��4v�1hp���"�`a�cn�����<�y���� ��?������=`k3�*�&wy��K�����W��İ�x�^=�"���p
��tJ�c(��_����0�E�,u�#����
�S�Xmr�Z���Oz^����ăzM)�R&b!1W@,���c��s��J�I*C�*�� ��@�+�J
z�y7Q�$W7��R��Z�6�]��4U���]��p(�X육].���4Is}tTC�_ޕP_r����;�����!Z���0�x����(	̔*��������"�^� ��^���-ve��t���L�`"�8�X/�̤s+�I�W��J����/ZJ$�;��@�Gi�*X��]h��=����T������t�PZk����Y �SO�4�ܞ������Z��3�f�	���ّ�ԡh�ŜBő��,��,T��5��
��gY�q�j�|n��}����Y�����h���Od�TsΈɯ+�.�(���"�=԰z���܄@t
볥>���+$�ny�k�^��~�m��b��"`�*yV�d��?B[e{$�2b�H:h|B��C+��p�Aj�%�F�9C���a��1Dt<�-+:�ݣn����M�h��+��c�ץ؜�|Hּ7�l��3m;޼�>2�y��LK�Q�h)걝�d� �f��������'���R~c�Ox�,�����1���Y�.�����8����c]�Xa�ǆz�����aNVb�u�`̷WD���8khu�`S�����, ��_n׸@�W})�����A̯�7s�ڂ묣�O���i���_�xX��G�K�@�g�d�~���WhN�K�VEC c��I'Q�i�����x~�z'��=�
�߭X����N(h�[����ˬ ��J��H��~hs�h�W�"�j3�i�| ���?���,���T�l ws���|Ab�4���g�'B� j)��ƫ��=L0듮dd*�n��'7� ��5|e���g��k�sPL�6o��H�v F�*fF÷�A=@Z7� ��Rw�R�LDˀ�A���e��0�C�46Tx�f��B-!/B�?x��v�����N��n 7MT?�q��1�+�&Qh���7k��p�A����A�P������ӊ>46��R\믦��,����-�UdJW'b��C��+���bW�E��̟���Ř�{��e� �<��[����:#��2f|˂f(��`�R��4��L@n����<n�f ��	�������r����C�����p/����+���~�[kX�@]N>�qk��%7J�ז�{46�c���睥'KQ�G��4���@�苁�I���~?���nZ�Y�?˩^[�/}�ڽ���z���������I��`JzyH�@��|\�_����^uQ�l]�����z�/� A�;<ƕ����a{Fg-���ǯ+k�qL��>��U��I�1���:g^��wbA���Ur�ۢs
��;��-&�:�u� ��+l�f7W�L��@�bش�p�-o1���O�p�� LLJ��&���]jǻUϦs���
#���1���ss��)6�HD�Lp���a"m���q��R,.�Y�1�Z�k��!��������nL�V�j���,�$(���-@U=�5�8�9���_Yg�{+��r?��p��)��w����:�ֵ�����4�n�A�a��JN��,3�'$v��{\8�{&�?	�ū����Z��`�2 �a��Эz�j�.�	jGѶ3��;��i��{�¤$#�{ȱ�������q���9,�(��'+�8����,�D��c��0�j��։�Q�E�.&����G.�Lo�x���ܤA��;��(�������=����;?b�i@o���%@DPO�&�'�|�z�C��͔o�wM���,��#�s��G1y�1ʆ���{5i��X�&�v�C�>og��:�5Ja��x�ͣV�$��	rU Խ`�K(>���ڍ�8X�<���ZH����Y)�4-2����inw��������'?�������1���Z�_Oƀ��t��P1������`x�ꞿ���5�Is��b�6�vI�E��	�Ȭ�<��Sz��\[~�f�mP�����L�p�:�>���,/��К�;!({��'08ݧ'�k*�g�0���}{��t�#�!Z��i`�֚$;��E1W _���D��O�\���l'�iR�G�z~=z�H�|�wZ#�o��~7-��Jﺗb̎�ya�u��$	��XG,�q����,�QL�?\<Q��u�6p�z������y`���ɿ�O��7aK���jRt?s7]��F��ȹ��]���u�k<�#��%R��i)���ϔ��ʯS�_ޜ��-��i�Y�3�Z���O���o4�|9E�r�u^�l ��p�ԉ�GR���S��?�f��ݮ������._{�K��7ss5M[Y>���GN�IK�'�q~�N�	Q�bq.v3��z�SW�I`S�Z	yG�T~'ګ��&K7���SR�v�Ծ��rP�3��sH"c:*�ݒ������ܺ�u�hy3h���#�䵁�&a9A�_<��T��@y��S�<$���gZ{��=F�E"����9h3���C|����@�69��$�9�i!��9��YdOW���"�@46��VNXR����kC������${�NW�q{� U{0�����z�j��:<����/��c����7��ӵ/������+E������ɭt	���!E1B6TE
A`2l�46��>�.4@}{И��6ղ�J��{NP��Z���R'Q6mآ>�����9x�k��J64�����~��㖛�w�G�i4?�f���ڃEe�ߎ,4w��f
$D��@i��	��!ӂM	`#Y���3��nZ�HX���`�M{�`�2&�#德�j��=��bY*&l�����Wc[x���B���w�L!1�P܈�!���DB�,EU��Kx��.�a���v�U��ܠ���Uf����1���Q;�P��*?p4�_ ���V������j��wf��M�`�pG�R)�	�P�gM"@�r��L���H.�`B�hE���G@��e���6 U�P��ZR���rE���(||9�+���Z�,18&%U:���SN4����z����)8b�S[g�U�Q�N�&��5� �L�[q; w[��L�Ũ�����h4�X�x�
��k>�4�������a4E�����Z�H[b|����{H;�	kjaS\h����۝"�^s�F�=wz���W@��p'L��(����E��
*�sF�Ծ�c�ղ���&�'�RL2�*��J��J^�F��I9�A�X���M��'KG+-�{�<Sd� ����:������R+����K N%�^���������e.��Ҋ7��A^ʑހ,�H~�ot*n�]�8���'m���U~p"�0��&;�h�K�2L�t��ص>V��1M���=�0���JR��=����g�EO���Ť*N�6?k�B�1JAzZ�+��l|������=9Yɀ�]vㆠ��@B�e�:�p�8A_�9nr�>�+�����-e*RhB@9�c��W�~��^J'$���*�E%�fp@Ǔ�t}�b�����@�ZKt�� 7�R�\�|���������Mﭜ���<򼑲�,�a� �jLuʟ�-5�o,n��f�K?�Li/Y���2Ch��h�]�4׈���,��� /VZ��x�b%b�y�c�S�(�:�yc���L�{���s��-У=:�^ym��nQYdT�;<���j}�9��J+\ �/�-Ģ���t����9@��>�/�5e�3'�~=�y���X��"� �b,Z{�&D�	�%-0�(��OvR�i��cq;�K��c�MY����cq��.�Aַ��H�\�碶�\U#��w��'�H��Ui���w��jf�mb���EUj hfH+�*��@_�(ԉ�(��W�fE��`��z#Rp�No
���gyK�UǺ�PAw� `�q�v@7����/�<��bj�B+�c � �4��e �Wpf��L�Οv_���[UA��� �R���6�<���5��x2':��C���c��a�c����x��ףx�p}y��f~��4�����G���1�>Γ���1�d���T]�E;#�b�p�[w�i�b}�)�9Ak�4ݐ�u����k�?�ӑxt�k�b9Z��s�F<���j��s�X����x�bQi���ƫ����V��qJӍ��c�Xo�j�K�h:-B ��J�i���`�H컹�'ھ�MY�ue�zC�A���N���&�;���8H\@��5V	���h�=�S
�Vѓ H�ƍq�=�NȜK"�%���;K����+ho$vn��պ3k~؜u��L���xɉ�-2J+\�`~ը�T���#�f`[�`�)�.���TyE[f+��؂��]5��Fnai�x�<���/t�`�Cw�5A���'��7K��z&��w�`6�}p�[��3�7��1	�-�"�ʵ��;������N�ǎ�.��h"¬v�28�V����N�"� .B'��x�l�1�����r�p�5���Ϙc/�<~:����\Hg�}fCO�E'�;怕�b�Y��������Ɔ����Y�Pw�\���<��� W� �n������~��x��V�����%���T#B	�}�PHfR$�fVt��)��~�-�˸_��7���LT��o]f�̱ж�����`#Gx1K�\�?� ����v�[8"c��+�������_������+�E����K��e�i_FT���lF��.ɮ�?���g1Rf�dt�����SSY�a��o?��1nH,٨�&�Hz�˶�*3*��on�(���w����QyW��ߤO�-hp�sƱūo��%$#�b����"�TG�@m��P5X��,�J2{��I��kk��������J�����c�>J(�����hN�5�vO��xT��쒍��!���u��E�Q��μ �!��U���Mӊ�(t�?Aof���VA�z2��-�W?�H+�,��.�w��o��k)��E~X��#�{z唖��	�^��B����ohR6Oʮ���m\�A�	$t0r5k|�.�|�}t���f��mya���Y�Nv�:%P�J��@�d�j����L�>e���)�`��6m�8�?�#�H`]ɬ��(��~&���2��(H� g.�E�il�3��-��$E�n�gW}46��v����`5�):U)�#.LA�_ѫ�CU��9��$uv���3k����7��:��{r���&����|]T����G�v����PZ��6��A����v�s7�P8�G��{�L $���;�\��e@wL�����MLm�\�,��G�Wm��y����|� ���O�â���b@�5�@��~��RE�k�ʜ'�)�B�ɤ��?}M}��f�7�k�l-L ՚O����|��?~�7U��񙒻"���6�����\��FO?ǀ��\�&��AR1��I��5"�ڏ���ȍ̥���8�r���M �mp�|A7���t�E�z���r�FRjF���	�1��S�ɮ+�5l����hT�Z�sv��0W�J YZ��~ٿxP�UqR @��|��(�j��l���9�)�L�&{G8כ��'��K���rLE��]EaD9\�h{���5^8�����}��1� �V-ݲя��Jf�oٶ�I/0èչ�4�&Hw��Y3M�*
P˴<��p�0�gu!Op��Q|�7�g��]C�!UI�f��~v'�g��>�%}�Z�#�g2����'���~�^�Hp��H�Y��ꈄ_�2p�h_�H�Z�K^�"�p|�H�1V���M~�4x���y�Y}#d�'�77��B��C?W@��"��k�4_�_s쌺���Q�mj�9J��Ϝ�U#.'��w�â!#I��pw��2����=`�v�R?��p:��@��0��78��C��K'ã}]Jl2 �L��%�GՅ�³��N*1B�ʟ����J�tƏ�ߗ�p����qT�0"n���Cjf�r�8�`du�.��H,��=첎+�'�������KP>#쾺m ͞@�����{��V� 늅6��FV#E�楠��N}�������F�`Qo�?�+�u�N���%��p�����љ7����D����6G��l��e*e��4 ���ن��3i�ɵ���� Vq����"G@ �S`SV���m�w��b�3��������W�'�Y�n�5�� k!��nY�E���{�8�]k3�+���t8қ[^ Ėm�bD#d��0�<D��zt�qj�_���m�	G��;�\�����
��ͳ���#O���g�y/ ��~8�I�90b���ִU�W��r���/�u�h�b��÷ѿ"�nj����S��wF`-(bsO}�hq�*~]�WC�W��[,nX��K�'�E����(���݉��S�F�.��>���"�kқ��
|�[�_^i��2��63\9�8Y=l��'=@�eO�O�y�e��6�H�3���֧�Ŭ%���R��6��^���m4��V�xs$l1�s�G�T����1$&���6���p��5�^g��|!?�Y���������`���a��ϑ�o���)�]����Π꥗g��b?# @6��y�,�i���#29J��x���f��ׇ\� ܭд�w����>����3��X������u��ی�pr�Q�X��9���[��b��r�@8}�eN�EK����<fVkj�Kmv�g�� }��_����"�d�M���Љ?gG��nрcl �H'Y:���:�D���E%���f5�}�XB�������OCW.S�VM��vP���aZ�|bN "��{�5���"PO�@Si~�6��(�S�z<j!�,�OH����/{��/�p��-f�@˧�(�E����X����5P��,�N�Y����qõ����c���c��S�x+���Y��
H��߫Rgjr��%�@�±{�.N�c��e�j{4f䱺����Z>
�L��̛��!�}>+`�/��m�@V��V��(�掩&b�zcǖ�ޚ�ѵ9i�ҰF$�g�u�a��8,߂�@���0"V9�!��R�� ��S�楄���򮒼c�S�00��J�~0��N���#�������/^���`��#�={t�Ư����/0k�<���_�ѥ(Q�-�\B��7l��37T���S!��#وqE�K���ن���h�NT7(��5���j��4�c�3�#�6���aa����c ��$C��l�y1��]ϱ#��]�0��ό�G��^I)��;)g�L�R�х(3�0[u��H�Ԁ�E*D'�rj���*&Ѳz*1���b7v	.��Ru�d�$P]xYb$9�x��Ӂ���	�ɰzD��F'd�Y;K(�I?,;Bʽ���>Q������U�۱B����I�s�)Y{1_��j3.��&�����B+��YT�����O�W���R���P���<۬�BQ6g���tf�# 3��/�{	�=�'}�y��=���v�*����,��Vזd ����a ��f��]�W�����88qz��i[�ї;!ŋ��E���Q����Y7*ZI�ђ�A�c]:�>�LۃDj.T��7�'��h�=�
�A�D?��4#O^�:��>�Q�e<��G��"8�9A���0S��?P���I9tE#�>
�h��%8@o��M墕�36� � �  4�ܕ��>=�(�Vg���;$�ٞ8��d������=��^��D�ɾ;�(O \����!!v+hȜ��$��[�����I�:�f`��ÆA^����L���!"��$�︂7k$n<)D�}�k�����_�=��2�9�l��|Hƾ���R)Bn`�~IE���~��_�hxW����}P���9��m9���z�ƨ1�)�d(�Zڙ[�C��K]���N��ұ�r2�P���Š~8�\M��!�����>���ڡ���>��p�g�D�)m|r��
6I�"L��PG1�3��i���Ԥ0=*���Z�N��a�6�K]`�+-1�ڇ���Z�v�+�A�]+E����/�ĥG&^ԁ�Y ��1~��c�i���D����n�pќب�87���K��x��-�w�U�&�n��	p�`�ʺ2H��qT̾��m/`�HQ�a��HE���Y4:N#9� �.Y�_Z/��'�5���Y}��r ���jގ��O���3�l��������0�Y���,�ޫ�2�#��^�,�v��̀����
	c	���`S�}�K3M��_32'�/mR� �9N����(C��/5���+�X�el�ݖ?n�C�YvE������@�Q2%N��"�g�v�e�?D�x03!���%Bt�P���79�a�R��ǚ�6(r��7HY���@r!�}{����xoR����m���h��cv�7��X�}.X�7,y�L�7ظr�@�5�#G��-w�M�q�����ױ�J{!�o#J��f�,��*�Mp������xy�se)4�_���ݰ�N)��,7�w��S�8o�|��kj�6,�3l�G���d'RIq�Ǜ�.]����X�|��I��h���ub���u��HO�vNK�!�Ů*�Ɗ�S�ߔ�]ZamKr��G�_Vt�r>ǣ��p��L��Lv}{~��|���ӛ<�\P��x�e��]g�Z��W��^d���~���� ����(��S�j��f���m~8��|t%ȴ�x��/#�A:o*����&B��U���7�s���5��ۼ�q<�8.*��`��5Ʒ���Cb�6qLt�k�d�'�Q�"mV����'��n xR�a���'	ҷ��9*}s���_{��qF�B��mNktj����I����ص��}��O�z������u;D�8PJ��:������ve���)��9��H5�FJ��������0��v�2��=e�=Q�8e��"3�f����"���sxD|cK��Y���J�&T��f��q���k��.�=�!���f�!�n���(����(��L��|��GKw�?�U2G@'a]ǐn��s�9��;�}�Xy�$�%Վ�,7u��ߦ��R�Z���(�[���~zj����R^�[���Ō�Rc�s�݌�#9Z���EzQ�&������N1Q騔�t�^ev�����aw��$�����P����ts=D0e�]� N�*Hӳ�/�\�"΢R����������� ���1�)\(��R���G�z��Ì�g
������7�L��[�l��.8���֣�Ծ~���F��W����#��"$Ќ�0�y��i�f��G���9�%�.�O�K.�EiS�`�-�=~�rrA�X6��V��b��} S��3�����Q/�������|�g�ȗ_�.tWmj��ex�Rl" s��F�3�����`Ú�;"�vh>�j�l��I���a�	cyF�OU_�$����<� �.?��%븆�iA3��n�u�>au���A;|ɮ[U'�A��c;���D�D�����t�vf�2J+9^�1�̌u�������Bǧ�YL�w��Z�=�� �xr��J��%yJ��~"�E�mc�o��9)�����B��8���\5��ڑ������v�Lz��^Rt	D�֤��&5��[Ry,��J�PͿ�C];{��Zp�1��-x�����ȓ=N;Xu�#Z��a��=ø�jj�<�<�S��w:�T��iS�Y������o�]�4z���E!<YSI�jc:��b;�O�ر��7 U� 1�<��s�I�x���BW�W>H���.����22����6���t�rē��xmw�X���8.�e�5F�.��O�8���P��I���F.z�å��`54`	�8([#ɽ���hYL�h9��ر4_��<q��b�⧂�- Iz�v�Z�	ٗZH�>{��⥧0O͝bP�Ar��}]K�V�؃l�i�	d�z�'�L��ĩ�(��4�IgL����Z��V���虒K�mے���d�fȷ�<�ai3���S������=~��P��E�0 d��`��b�T��
��i��tԺ��x�%����*��@�3&���E�`�O0���F�{!IB䓣�_��}�$�Y<�V�.�����7�\:wrj�;brYL�X&n�����)o?�d+W��,�8����)p�8�xU��)cۊl'�ݣ��D�+�D��Z�c�&�Y�'�oEM�V���o�	>h����˅�B���Jߗ���%D^���"A�8W�|���Ῑ���:&�Y�������Om�H�0c���a|a�q��OeJC)I�l���~қ�~]�t��k��+�$a�����y�L�8Ksn��Ja��ܹfeZ��~�j5q֙p�����Q�Em�H����!13n��s6��(G��I�r�t�8cڨ��VYz�z5������W���o�����%�xo���T����~�K�7���je�L�:�����8�P����^{�it^���5���$'�:7:�(�H�a�b���h:bƴ�)0� y%pI;����ߗp�ֱ�+8k�sﾎ�r���{�9<�c�~�'������O�����Qf���{�V���~-���Zx���Blsyf���ҩi=j�8��?�.˦�&#uX��o�d%i�f�v�q5K������N�R��x�Ms����g�1�Ӌ��}��{.���?FC\W��eĭ%8F� ]ȆV�ե�����t�u���,1M���nR|k�a����9u��Q�!���ny�^��y���!�xH˷ZKP�Ü����D4�d�|��5�{��}/�P��� ��ASmk�X[�IS�>�b���A?�J�ι�/U�Gnd/zMS&�>1�:�ߦ�j͔m5�4�UjIѺ��e�w�#�La~���=�����e����n�qb9|��.�D�� Gᔬ
-p�&�"��A7Ϯ�t������+J�|��9���OC�1w^nK�i ��B��m^2C�b��x�Ŵ-��,>-�DT4�lR���9���\�孡]�� Sk����cW�e=��0�#N@� �|��c�.^֑���"���P�&���%�iȵ�ң�Sx��X�]|'�hD�̖�;��������rL�����@�.uDuUjN55�<�ո�������o������i��ʿ��Zc�?����6F�_Z��%�P_c�I��1����GǙ9�T+GiZ'�4�/7�d|<�}�`!�os�hڧ|� �9gtP
��)u��k�+#m.�6$]z�7�B�4#8TMҽ-Z�Z�F�v5\����lIY�����/O-�4ǳ��:�um�o�z�"uH��jCLبtl����c���/�[j����Q�6��\�/idO@��A�Rs�˙�
� q�-5�* ��@��{����^@��/^q� ��|d���4|��v��~Z#׽d�J����������8j4Aa*�h]4�H)[/).;Fђ�}=�G��!{tp��5&�)V(��f]u*����d��ɑ��K.l7�4�?�|�*U�Sr�PB�N�@@��L�m:%���#q�O�m�O��A��j"\S)E���o>����<�N�_apeə+�>��)����\AG_s74��8�=�W��V筛���bņ�l�ǉq�r`>����XC"��L���ώ����n���O�����Q�A��*T�H�D�7�ӂ{�C�}�����S����Yhʗ�b˩|�;3S C>��� 3):���c�{��u�C��]����h	W���P˜5ݼo��!ֻQ+"�>�k�)y�$�\IM��d����_j��PyA̫��L	�=�ZQeB�7���q��5oS�l�u����& <o���A��;�·����E�b=�kD�x�1q�Q"�1���9݅��3���&n�%��!��:���Y������n��[[�����ӄ@V�ʢPBps�&�U�}H��뵞������
���݄�e_�V����ȑ�juqT��wrF���W~�K����>Ƃ�`��&��?M�����39�ౢ���5|#nF�K�$Ur�)��E
I2�b%f����X֮	�� ��.1�@�2�L�~��e��3b2{ͻoC� �|�J���������}-�>�7�	����E%�<������]��Hf�G�y�k�aW����t����V�Λ�����nd&_p����Ƈ�������\$6uvyb��Z�g�����K��u����T���Qf�_�`�FYG�n/�T�C�����I�~�x����sU
�����_Z �C��OJpv���P2&�R�m�FFy�}�0�Df�ZƠH.����@@)M4 s�s��]Y�#Z��9���u\��c 얻ghs�zXɖ�<�����`:I�Y|Ӓ�~���v�sfY��ėAkxk�+l_�=���z!RW��ہ*8���JKT
��Vt�JK[T�
��`�ߢ�74�˻%K�AR2��x�;c��?F��F�1<���c y]���"
8�D&ާ$XFl���ݧ� ����J��6h�k��������	�o9��i��3CI�	|�|9(ڣ��G�ٚ4Q~I��	�Wh��_��<�boSJ.]b�*���*,;����ɼ\8D����Zx;,b��"�f��W����y�RQ/�O�p�m��ѲSɇx���
����v�c��5�U�A��2>�2� ����ԸsR������Xp�q9�6Q�ՇZ`���l����-�e�Q�9׮�����3�r�2EE����c-.������F��f����(��K6��<�;0HZ[���8�Nq���П~�����L�N�Qu��@H�P�Eo`�r�ӝ��"��A�y�X.ԟ�5�ҷ�
��e9q��D!HE��o���d����ആ��^��p�`�����X,�-W��$*%�阈�Q(�c�BO������~��:�����d��꧅+��w'`��7������́i�&�k�uƇl�N��,���������R���=�mJ
�&h��p|�AY$�Ʒ{1���z�<��kd,��'�L���U����L8�]�q �_��2�;씋�7�Ì�dJ���ZG���G0-���q�s2���g.ӕ_��3���CGɆ�=�82�.K����ߋ�H����L#8����@��vc2b5Wڪ�`�k��u/�S�]��=��首5�FRV|�Xp�{��)�F���/U��}r�w	k<oi7m�5���O��s)Ww]��l603J
�����+x��4�����pt�'*�K�d �C����(9gr'+X�E��+`�̗��\�yzb)�gF|�k�n�9 �{`��Io��O�~w>��:�d �Z��'S|�w�=���%5���X�1�����ʳ
{�T2�$w�h��]��ey��t>Q���ńFV����-���?���׳���)�wwf{U�~T�2���������L���.��$8���9����m�������).8/L���W����_"7c�YS��P0�FO�������3>��K�r�����!N�^�_+�9�cܧ�ߖ�/O
��,�@��|ֶ�h@	aɜd����<Ҭ��#峿Q�W�r$�?�VP}E/�^�����p^��Z��D���U.���Ӥ�{ZI��aׯ �$"�y�)JGXD������ve��xl�!���_t�ާ�a�d#$5Q,�$v�U�E�pyr��_�)^�ޝ&y�9V��Yd�wy�8w*��U�'��'l��H��<gC��@�~�?T:����lm<�]����L�/a�V�㍷_B�/3���1��W���Ȧ%݆���^�;.�Ÿ[[��� �ִA;�1�8�8O~���@]v7�2���ۑZ(��K~��Dp�S�;�]Tܹ����~X�a.��|��P`�dTt66=�Bpڄ��d��:C]�<��ed�.?#��}�tU������;v�n�(h��������J"ur%��;��譴[.n'y.*�iC��!3�I�t�%nX�{�����T�ߚqJɅ���@uy��U�eW�����-!��;mr�@M��Ql����4<Ydz��W�G4�f������^ ��࠶�C�Nt�Zj�xVgB��m]�X�q�~�� �PN��~��_ao�X�O��.=����2����v�h����|��^�<��{R@�!�#�#��6��{	���:ֽ~�����z{E�0D�v�l@�����y(G��6܂�G��XU����cR�x={[	S`��Ts�rό��� ��z~�OР)$ 	�~�T����۝�c]朝��(:��5�����CE�q�O���20�`	�s�y����)
��s�'t!g0�G��1R�UM[��l�g���ٮؔig�F����[+Ew��v~x�ĦWN���.���I]F�>�z*��
�6x�Fx3�4��8�@QQҦ�s�|��@��� �ep����殎�)��v��[��βO:_ѰH�nV�N��]K#��q'��X
��x�<e.�4:��0�
jY���(*\��������'y+�� �b�?��;����e� ����r��?�c�B"&���z�����Xݡ���Q��.I��e�9�,i=,�(�۝ޫ��IG�A?��׭�$��{��E;�J�'�ח��g{o�j��i1����.��j�ihg��%d�gp��|"tch�![S�}P͎��N��.�/�g�M&<2]�J&�,�.��;��țl�5u�]J�0�����ͪ� �^�3~�@>�p�H���Zm���J9�����lT��p�^�ܱ98���>W�b;��ڍ��1S�o2lSn�ax��%�:�@���qM�4���
_@�YO�`C���B\�d����t�2�)�A���N�r��6�s�d��8�˾���PS��䦄��%*ZM�f1�YqOH��������v�a� �6u<�X�vM�m�����턤�a�1�xc��q��lN��6G�4�B���b ���
}��l�+���#"6��������M�b��#�zkmւ���i�y�xOٗ��w�/�8ЯI�|\�`U�ѭn�e�I��(���>~�U¹��v�#=n`�fs�"L�k|H��'e�-�J�Ç�N=.�M��c#MZ�v�S� Nk@��hz�dPƊ�����<����O�\��ҊIZR�9�W0�ʽ�SsQ���]<�،g��k�kf��U=e�,��st�E���ڸ{@ ǋZ��]ܞ.C�C�>�tV����Y�)\E���� �n�W&\�B����6�|�:���V�	��m+��0�[^��Sʡ�+�Gq؍������d�tUr�Qj{�o��x�a_�S�1���M���&���d^��}~�GH�v^���(W
�&둣t�'ݯ�y)�+[i�L��Gb�D�L{����x2��/�r0���=:��n���_֐29�(��>e�F�mQgӀ@�$clȴ�D%����E��ƹ6N�ur4�]�Y�%W$Ϳ���+"�����-pw��w��"o��THk�5���H_ߖm����������ƞs ����.!�)�*��%W&�Ցe��T�6��N1���QgO�������:���Y{�+`�ɱ���!��ި�>S���m@�{�>{t��v?z�d�QV�|�Ԡ�e+�\��Vc�Ӹ��v�jx�-d��;�]sZ�Xь�M�6�ig��Ƅ���+>֜R|i�b�o�m�]u=ަ�c�������2d�y�^�0,Vx�Ga4�M��D�3��b2'��S��g_j�� ���~��U�ƾ��h�b`��H4{Y���k~.*i��t:�C^�+�Ӱ��U�Ił�c����$2�\Ӕ	wrR=FE	9,�9�L0���V��m	m� \��`szU<É�q{t�w!���LT�Uz��x
�c��U�g)$��
��/�3\V(Ņ���Po�q���(��#�UP�e��\�T���]?'�
!7#+�L�n��9({���J��Cݏ#)2�cY�
�o1ZmxB�!@���߻���ޖ9�wP�F��ƴ���H�9A�O�����?e�-���14>��dfA���������p`u�$�CH�}�'<�_�̘-����}�~i�ԡQ��9{5��d���ɍM���9=��3O6���oc�d*aL�E0�t+�����\Ҹ�+����,g��gO'71h�k��!Ү�k0_�����'7��Z��4�]-�k3��9��9'���w�~�3����t��Ȱ	�3��N|����V�	n�*�e�o��ɷ�}�+q�H�c�Z���,�d�,̆\߾=�ے�u��TC��s)��Yn�|������fͺ�v�'7�Z���7��~9��f�_&�#��o������&�B�<���t�%{�W-�.�k��f��+X� I���H�x&#�����k:��@Q����8��鈇��yOm���* ���}�uo�w7��Sӯ]H��TXR.�P�JLZ�S���pc���o1�3\����v�H�LQ@:���P��L����wa2ѻW6��,rQZ��-�ב�,D�}�J�=�_�A�̀6(I�(�a�{h�A��
+V|�$j��b;�aS6C/����
I���Ȣ���2�]��'��C�����q��С��2��ܶ��7���R9T[�R�2n/#|�KNl�';²g����\q#ڍ��svS�&��+JE�)���9@V���v�'��=^Z���|�ϦX��P�1��,��j��ԟ+�C�V�},�
T��JB�icO`��4��M0)��̒�G�6Ю~c��v��݈p>�������NS�B����!�Ԏöǟe�TF��,��j���* �C�Rg�Ȭ��jƲ4Ɉ?����d��{ך�fko��gE�z�B�S�L��������}�
�gJ�9PR�॔��<t Ƽ�.���Y��;a���(	��ԵB��B��/8&��I�y�
޶�I��(�I�1jc|:��޵u����Z�K��](��i�{1Z%t9��2	�F��v9 Os���#���S8e���6�O�ӭ�4���T��$�wL�}a�!�E4��?� �w<���3��я��\B����x��`�Ӆ-o㺮����)hX����mb��+�&o],�qĐ�ݱW�W�^�%Cg���pPVCUp2�Fl�S�L��9�ZhJ o�� "v�k	�����8_��h�ʣ=���5��[�U����&{��6v��c��f VY�q�b;�X˪����QO�
������ ��h�N�h�oo����F<�t��]��BR��q�?��,�O�f��KB{ƽߨ:l��X��z���Z9����I�����6�a �*4:�w�������|�,�.2*I�ҍK�ʠ�����W&���z��sn^��'-��f��4�rŴ=ʾ�<5���XP�YՅ�%���'�4�g	��p�3�Pak?����*����Ǐ����_並w
��К��H�	t���u���uD��~� c�&��G���w�`ӓi:����AV`���5���������=�9�<��7�]g1�Ρ=͊���t���f�6$�W��ib!N����N ;]�*La��
)u�+�Ī�I4�))�RM�!^���ґ�u��>�����!S�֏�JԪӅB�ܳ�S'��G(��P#�Mܕm��Kw���D��B1�X���G����0y)��fV�{��C.p�:s8�-���4�yx,�g\��>�ORX�M[5�͋.�sC*�8�Jk�x���R��4!V!DZX��{y��o���q�q��|��%Z�0|y7ueCD�|�5
7�f�4�.�J���lũl��(
�7Z����͑��������U�V�,�ӛ�3��B#���?�<���$��>�㮉�D�m�j�f���"Eŝ�#Mrw(�W��e��
Fgn��S�w�y8��Kh�)7����d���x��Dh�����g��8�;$M�9'��,��ȕZ¸���`R��;����"Ǳ���:7�p��t���I��T��h�vcTS��[���:'���0r�K�וٚ3/��LmTik����T�j����;h���l0�u� ��f��N�B�8��QO�R�Cv&���}���h�P�م�e����hU��ߤ@ϊjʙ$�s�e	���R��
U�ML�9�]�M��*>�Q����-�k��0�j��?�>�2˷�N|����E�cl�Xc��Z՟�&;�8�m�­���8��/92�M/�`m�GJy�;6��s���h:0���N>��<����zf����ӳ�@u�Ǌ!�.�Xn��A��n1�e��W]�QB��A��`��nA��<|��:!d���f��eJw����B�P˴��/���"i(�m�1�2j#2�6gi郥qe�i"��a�w��i� 6[���V�r�������
l͝��Z�G�]p63q�|n0q�r� �if��ogj�Ke4�V6ln7V��q��#�F=�/M�����B���|�����T���x��łd2�[�T��0�Ӱ��=]����cF�� �dF��l�^ti���b[jɐv���ת�]�A!u	�#Hۓ�����������m��oTO3O�����6�}h���ף�'�F��sͥ�4�9'x��.D�Fg�?�28���=�Qvъ@��c���^��ʯ��6���k�L3D
U���&n����+��n���'�r=$�>�3�b�	+o���hܡ�;/��*�oD*�����47X�=�}�����G�~ؠE���6Z������_���M�����w���m<p�ͩ?���Juf:���w�G��dG�%�N<#u�D���2�Ұ�E�I��[�{.�fm��UV����$bE��{�K�XѺ}Q�T۴��,��/,�H���,r��l��<^3,S���Ō5g_^洠C~p�F�Ki��@3�RWi�[�xJ\0����� <*��3P1\F�y����i�a���?wKɗ܃��"f�}�b��#>GD�]nxq�m�}���8���+��b���s޲�PB�*6�*��L�?de�������O
����G]����ī}�iV�_g2�+���>\,is^��G0�U�Bbe�w5��{���.<l�6.곾��/�%�]�tQ^���E��B�+If-�\�)4?��0�E��>K5g:��L�^��W�`۱���eo�"������^b�[>��E���*��c�c����x/<�"�cw�����Y�$@��Y�!ٶ�T��� #�7�@	�E�v����d��9d�}_f<�si�Q����ьNT�z����1�m�IJ_
K� ����������|G��L��ޭy)����Y���K��D��$R]7X�t�K|�V�!;t�;��E�x	�u�劜����;�>o|vG���ėC�[����,��U�YB�	)�)X�9��)��d[����$q��F�0�Uī�M~�qR���m�2m.X.q���q\����~�������k� �l9��ϔ��Mq[���Ĩׅ*�±�@Y����#9�
�� ]�y�3H����E�M?t
�@ITS`�-�%׬�|��-��po�"���MpPm�
���FV���!�Ӕ	1���aTc�v��Q��H�ydZ��c�xꥬ��66����rG�5j��N����d��{����_��\��l?+�Q'���;>_%s̳�Vt�b[�Z�X�".f^�X5\�[*v@(�@�������l*f�%2��W5�������(I��)��hQ�K�5:5�	�_�z�U�[��������vru�N�$�D���/�[p������?H<VA�@���/jL�E�
~��ݩ��)�dZ��V�]�jS�vr��%n�>�Ex�o�0�P[%x	�7�� 8�/����Lo���H(�y��\��w^zt��Q���5�ʰ�q� ��HM�`�r���O���a_����Iw��Qr����v�M�"���;�d���0��ps;�Us�?��NE��"8����HҔ��⛱���o����bx��/S�R�T�����a�� ����H�"�M�
��]-��J�n�Z�TϦ�����!�T����UR�(1�����npꡝѮ�E��X�G�=���D��BLG�˟�m��p�B�����۳�f���I��늛���sYq�`�P3+���� �|}+���f�iOualN��"-ZCOi�Θ8j�0��qE�����#��@E�9�-(1щ0�lM�a�@E�3�"Sء	2��5*�o-t�H�����A��j��
�A0�{dOAƜ���#w�ls�?񆯁�K���ܡD��x2�{j��(����qlHBU��)�j�P%�J�ͤ'���H�h~��3�����\,2�Ի$;�([�t�4��~	g*��t9�����Ȁ�G���F{�Gj�$��qF�Mߛ0�i$���H�9{=��7�� C������C���P�q��.�5��&�>�?��Se�l���y���>��(a�|�77��	�8�]F�9/��"��V�h��W�N�r������M��g�j'���c��ҟp<��b��Ё8-u:�Y x�7J�%��
�%L\��-mߞw־3�'�Wvzě)}^��3�4�����$�m�ucO���%3A7�U[oë,x\lά�#iP/P%�/��@��k����ץ� հ�=���(��p,�}#�I��i��Tj����@S�-���{���ՠ
�;�{D+P,�BYg��ĸ�"���;cu�N/�������B��`��tr�T{iUx���JrY�ا��SW�?>L�
LkP�G|l͊;I:wY�o�`��s}��� �jVD@�dЌ4�2�P��90��`ǜ�e�x����[>]%w.䧑���젝�݀B�p�14��>�Ռ�)4~�n��5�C�(1WsU;6��	�1����_�ԧ��o��&3'���4��A���tel��Bp)v�C��m_�_��,�q�(��^,Z��E��r����fQY����%[�L��AZ3!���.@2
-ɏ���R�DŎ<�"��ߎ1ˇ�
�habv@?�F���ty8y�� �`t��H�v��/�4T�]��hbz�ʖ��8RnDq�K8�A�`,�l�6�IY$2�SB���F��)=���?VE�O�����|�cm��[�5o�������&L�8�=�|c�P��~��ñ�u��]9`�S&ď����W9J�3��D�/��N5��x�$����\�ޘ��G�dS�v�"	����^���(�g#|��i���tP���w{�X�X#�������3v"Tw��ZO��0���׭�G��j�4hCP=�������P�^��7[*(��� r~$�ro}}�бp ��Z:�wr�8��%(��T�`�ZH}F�AK�;oyV�ȋ��:�i!�@*��R�j��>`����y�R���R3��2�i1P[�_�|�xѦQ
���ǯ�c�a�o�Z`0��Bp�����%����cq�~�u�Aaܜө�Ӻ@p������Uظ'��w(���-N�l4v;{�ɴ��	ل�~�T�1+�
�F_tc��X�WT�S/Fv�m�"Z�`ұ�� 1�Z�Ip����7f��I�^��mg�j)�5�F�����TwwlS6��:�p�g��eVX�W�P�R�9#������� �Fq� �x��a�swJ��Upvf,R�q�*�*��KX��#�����H�0'A��%�@�j�v�e�����.9����As̸ " _vļj���$�b�pq���x~Ҧ���85l�10��vHΈ�N�H�68�_jo��(Qf(�yt�/�����U?�=�#~��=&��ŕ�#lt�Y][�E��ف�G��i��Q�<��A�v?^�Ղ�ᅹ�?�h9���4���AEp�J�2�=�%M*J�\/���ʂ��Kbq��k�����-�L����Yѐ $�I�&�y� o:�=�V���k��JjH�阩JM$�g�5�ʺ9Ɣ���;6����Q��Q�t9������F=jr@�%YOx���rR�M�QP���]���L��u<�4�wf����$�.~�� %��;T�<^[Ɩ�-i�K���h��_�g��x�4}���7Z�~u	��|]s]-�S��u���.9�z�F��ьiCL}N��ˊkoz�c���]e]X5�뉴�R����b~���`9�ҡ��R��e�cq�mrc@�ZP�-L���B����c�2�zc���sZ��(�0at%�k�R���@��k��E��x�%��>:�60]"1#Hg�ǃuY�%CS��f�,�����N�HM�Ƣ�_T1۷���s�y|yy.!Mu6�n��x��N�%17TP#�;gƻ_�w���26WE��N�ԍ�j�rȄ�,����]����j�&MBҡ1��xD&���mZS�]`���2��Z9��${^�J���&��#���A���)^��Vf}p����1�og��s�N����Ҩ�.o�-�b[8�����Z�S��ʤi`�=������ޮE ؂HUt�)���x�k@߈�Oh��s�l�w���^���C\��z�硺aE�����G�뎋SC�U7���'�tA'P�@q+���Sj�k0�o'��1�xx�kR?~��g���Y	��(5�I��5�G���$z�tѬC���@�]���jK�������Й�:�M��ph�N`"���l#�K��F§2�&��?ss:Þՠ���P�E��?
iBm�卒�Z}n���)v3a �+y&�EjY�d��U�6?�b.R��by(�v�Q2Lo���ٺ7�R������r��}W�����qX����i�>o "��/+���+R��z>8�Cte��X��Ʀ~�ê��ȷ�TL�X��H��n��y��3Bo<���x����.�S��h���r�'�D�Of�8I���K0�,1�cz�
��5���3ԅq�7��?PM~<�Pw�B�IA�3�Ճ���a�Ӟ�)�.q�LI% vu��3�7��:��Ru����b�o:r��&J4��k5ʋf�ߖ��w˵���!�e�#�S3���M\yf�<����f E6��	���}n(�fo��`}95��-bg�BX�Q6㶦R����LF��Ϝ���iY���qFos�63�>�7P�z�	u�������:�ȵc:�q�y~��qê+1O$��w�f��KPBJ�O��b7����`���p�!���nj�3L��$��ko��g h <�RK���8�灝�X3�����Ƅ���U��l��Uo�5��:S�Ѷ"��ձ�xkD�n"?�Pa3d�b�j`���;P�%�2�1(���<@��t��m3���5,'�p��ug�F^�q� �>
x?X<��*y4��/W�~/q�1��H��Ⱥ�1@;��l�ߩk�=8i�aԹ��;�sHf;"�J���Fo��>Dg��)Ҝ�F��"�����6�Ҵ��q�I�QA���.��7{ƿ�84h޳a�y��(9w�7�WO����BNe�p��vU/j�A��i��nj4�pF��H��ac�˷�T�N&�k�'8\荍��=}����9��)M��3wEh(.f��i{`��hDz-i��35�`s�f�=~b~f0��#��AL�36��a�w�s�Gih�.@�W ת��� U��B��U=�X���)�B�F85mD4�}F�7�w[": ?��ylѦNRhd2�W�r;*5�j[,�6�R��7+8�{uǡu;v~���� BA�Kv���d�G91)�Xk�D�(�e�ru_�ǩ����0��>!���;�oQ��H��M:'`P�;֪߶��W�u�'4|
j�ȑ<6��Z�ǝ|B����=��͙�ɇ�ŧT�|DdY�q�A��CR��W�H��X!�Su�M-ȗ�)S��ԘK�Pd}�V�Ҿ�t��v�)o;I.�)J�j�D(���O�&�Y�E���I��ޓ*�K���w{syq�ۛ�>puI�/���C�5�'����z�nw�#6J	?�$BD��~�����^��M(	!�0t�/a}b�ޣZ=�r[��J�(�Kb�����V%KU-����8nUuRx{��7p���?n/8�rm�)#�,�C�s����s����12R/���U/'���^�P����)}��ݚ|�ᡤf7� ��2k���6
(-�e�m��D�O�rdB]�#촐�@���56Fq�	�ݹ}��/�T^��9���$��(�e	)`�.{c�Q�7�2yi��`^��A���)��)>���:��¼Zq���~*F&MlҨ���&�~��������#�P<?4rL{����u�)��3�$��\k]ع�	����������^�6`�xA��3��-�@"K�q�zȨ�59�����G���l	�ue�ͤ=c�%�םg��)P"x&Fa��>+VG��1	r0�3�[F��]=8�Ե��x�g�d�fp��zw��<|z'Y��~�K�~�gE�2F�XG���h����kgP!3��6��V4 �[`#s�ᮅ߯|E��U�Z<�Ȯ2�D	k�ӥ�ֲS�ʫj�uU�%2�<���t���p��[+ܳ{��8_�F��O��t⏽��un�P�,�R'2���0b�b�� ��|�������f%�ԩa�������ཐُ#O՟�����
)��
�A��;�֔.4�o~��[MׄvB<���*6��2�ѢOT\E�O��X��ڕ��\7�|�wE������z���K?��w�Ws��(*Sx2{�s��f,��9[��nʾ�՝�%7!��<���h��� 
��-�JX=d���,� ���ѐ �D��f��X�dM�m�䊻@�@C�b�u]����F�>,"��.�~OV�^Q#��b�C7�8�΋���G(KR�K��b	��(\��惈Q�I[�H�4�;֩�v^lO:�,�Ώr9UE�k���Z��H6H��p?�A@ ��ڔ?��ܩX�ӊ1!�f�-jX{��*�:�js�_�qn!�՗z�3��"٬p���1�O����StS��p?n>��/���u��o)rg����������k[ oDC�d���"���*��ŷ6�,h���#l��.꽚�;`8��<���D&ӞNaF��� PB�-��&�t��U;��i]5{�5C�1�3�����V�A靗�����=6m���Xki�~mV{�`�d�^��/�vTo��(��u5^�_>��o��0��QGki�괍�^�+�X4>��7�(^͎�_~l
�X��L_�f�ΰ�]@~�>�
2��Z���>yg��1g��+����v�����gOʞNIR�U�:(��9�bs���^�Bw	�X�A2qY=l�N|�~��=(l���RL�0/I�XK-vA��h\ݞB�R��&Y3�G�<�̯�D3P7X⒞�/�� �{XM��`��qgs�F��۲��p��X����'��$ݥhI�T4*�����& J�WGMX>�O�Z��p��������O���Sld�m㯞_�{m�.����BQ�,l�9���	���}nZ��K��]/$p�G�\h`���KM�?fd�I��d�Ð���|�b���#�"ȡ���T�<۲8n�F>���`P����~��&��W��<�z*Ӱ4���Z �[ꠂ+��8��������v��_u�<y�W���@&��>�I�s�p���LA�Ҏ��/ے��
pEL�T��Ҫ�$�vģ�G����bA�z�vZ��M@�(����m�;�����#&�ZT
���r2�Tq���M�/�&Np2`����b]���]����p�L� �e����{F*A�W�')�zt�2`a�7�����%N�ё��m�mHI*K~7�x� YD��[��+f�S����|4-L���̼&3�����J���Ǫ�	v	S(�G,�凊������pLڃJq%��
=9�^�aw��P|ܷR�/�T�`	sг�y�K+�@PHe>���w�^��X�$9&d<k��]͘�O��ϲ������R����u�Z���s��u��Y��C�7�< �C�r��Ӗ��L�"?-x�����+x.e�ԘK�x���^��B�~v)�#���2�͕J�R�Qo�oqy��{�����N�w�
U\��+�[_�Kp
,~�N�-�T�L�l7���f���L9m?Rh��
�|��<�"m������b�()��9Є��v�r[��aӭ૗;9x,.rv{���b�i�5
N��s�@7�S�i���ϼ�:�մ�I�ٶ�o��o��Pj_:��=2�(yTa����m0�ؕ���R0��&=���mM�Y�[�-�p�7�!ٟ��fٙ
� |�,"�Ƃ��Zv�/�i�yh�t��W]���;0��L�����p| ǈI�	�	H�|���A�B�c��L��P������"Lu�~�:���87'��t��Vg[��xM��6`�������o��|U��ݱ3t�j8WI��=�+��|Gԕ�=�=O�t�V��������as�x_q����b ���ə��*�$�q?+�M�����F��.��S3e2�v��[�����A'�HHo�*�Vo���\W�>
�z�V��������%~N��:ۣ�5�[�p����ֳ�R����I�;��}Z�	��7�Ye=R�����Le�?���[i�vHt����'�bR�d=��$~O��2����;�5�+�j�H���wܷ��_���~-֦��,;L��"@����2��;S4B=.O�D�������SC%bބRЏ���� s�ԕ���ҕ�7B@h�8vx7���/(�f�R1�li�R���m4deZ�7��<��/�V�X8U�G�H�U𳍨 �V�c�7+~s9���u�jh��LE��OV�ܰ⏗)VJ��յ��}A9�=]�º:aR�����w#}�i�ە/�.kR�ʥ�>k�[���0��G~аD��ߋڃ������T
�����!��Q�GO��J>�~�3C Լ$�^Cg8�03����
�0g�;vzN������z�u�ؖ�m�c!�����PSr�[�0`��[�}�o�_y�_�c+�z&\L��ޞe�H�;S���K��0z���g�p�2��/�REIfpх�*��w2��K���|�G&bЫVaR^4G�B�c5��ڈ�8��uIGv2	L(m�<6��	8h��J�uJK�jF�F��6n�_<��D��Gai�^�'#l=č-���gN���a.Q�1L��3in)����L��u-o+%2]�Lw�s�S����[b�>F��������b�1%�~j���Q =�`m�ݓ��љV�дMcj�[\i
��{Gj�����Ɲ���|>[���n��DI/xo��9����fm�nU,��1o�f��ffqJ07����é�$�Qb8Oal 	DM�H`���*�1s��3���΀����
��b!�����ŋ|RVL[��d;0��ĝgs�}��%�0)�Q�����L�3Z�5��wdk�c�+ݍ�B�5�g��(��hP7��%g6Gٖ��ԣ���Y{����[,"l_�*7lܓEr>T�lx�i�������4�w ���������%�R�Z�9Q.�]%qړL�a�df�L!+: ZJ\�
DԜC�@F9�ǧ�:���`�=E���Q]Ԗ�X�v�S(/ ���E�D=�I%�d���K�Gﵠ�����9hz�����HT&��V�%���h# _���� ����Z]rUo���)��שUc[��CT�.���A���Dp�z��5"�?#IO�}F���	�B�d���60�F��_�"�����bդ�|�v�7��U���YH^����6���ě��"�JRk�3�7�9�8�k o��2b�c��IEyVN�7��q�ؐ����?QZ���@k�4�K�+���{�B�nn��Hw��l��Q���)����8�vQ�G�x��S�\���-�(��&'��3����G���(����P������&�:sRP���x�p��]�V��享��di�9eį�Z�I� �����/�R&�ͱ��RF"i�S����"l�u��]?,k|���)����/ߠj\��:>y%��MW��?�%D'Y�I ������
�Ih�ґ��L�@ȹ(aU���W,��'���I���'I��L���� a���1�j�+7��&J*���N�� ��x��/J�û��軹�-�2%��<��?���WS�A��s������S鵫�����2��1����-��hnߕ	Z�=a�?����I���6{6C�*��_�ȉ�:	\�Yy_�Op<�T��e���Z`b�ml��w�(���)�]l�����qyi�4_܇���Q�����:A���W�Pk�.|9�Uɔ�;Hɪ-�K9E"f6ײBP����.$>�ZA�LL�`�L��ܮeu�G�o��M��>�%FT�5O]b:`S:?X��3����a�lB�%�i 
)�pja-x���KӤq�����cer�(�?�v��#��F(ܭ�"�����k�a6��kc:d���.а�*��Ĵ���=���S���z���l
z�/�&l	�G��Q�?�XƁ�Ͱ��|Ԅ,����A�P���b�y>��E����M��c7�\yC[O$K�Kg�����V��xu���K�IE��O�څ���W��X��u��A�qP�r��ZY9�|��X
#��L�8){�\��$5J�����g���T�2�g�ca4����6ep� �����S��@�_�1���+q�������q	o�.2�2@=����֧)ȵ]�.X��~�K�SȌ��c]��f$ O	D�i~��K��3�dI�ɽM�%��6��X�T"��&˴ww��:8ܷ�O	M��/i��s�0�����=	Ȇ:+1RJ�}��2(k��֠y���'�>���h������5duh<���NE��e�r��Áx� '��±��o��I�$���I���-���կ�0x�h��a�)����_WM��
�>f�E��B��1���N�G��|&�����&V�L�PM<R0 �>����Pz��w���JkMvP�>:���J�[�����-����A��z��4�u�hV�򞬱	r��7���ļrƫ��~���ґN�(��2�3��v>@O�r�h^
�I�V��<�ֹ�Z����!��c!wnB���n�v�rw��#g�p�#<��W���Kt�)Cq�Q�(KC>bq^9;�Q�E�ء���&��|�R�q}��2L�m���hl����OxT5لL�����GoT�E��_1^���CFX��|d"�G�.O�)�=9a��W?�'�zW)�z(��N�m��z_�=^���GpL����<��F�M~�뫯�����G��4^6f
v�:tT�����	H��:�S!��Z�]"�:,Թ�;�!����p��a��33�t��xZ<�v+���^Jhr9k�:<�0���ɓN�t8�|�.d?;����Og��b�&��=;�����4��ӖP�:�����%$����I���@�mW��!6���c6�;��]����xn�7��CO������6���{����H�iK�qG??O��~q��!YD��O�ܪ��k~��7�xf����N��$��ÚG�q1f�*���\1	��ݨ8׳�̞�/���쭚���Ĵ8.�$�9P�32�?1�Q Y�K�� ʲ���C���\B��G���&�ꕥ-�� �{8�bV�t��Ȗ�F`+I
 Z�+~2�,�;=��cP��q��~���g��͙!����@�qRC���%Ɗ$��@��{�u��ь$��Z:�%�o�3oAYjp=���h_f"��\%ӄ(qN+���i�Y�!!��r��s��F��T�ȵ��Q�Y�U=�K�r:�|مa�{�<n8���2�.vϕ��&�j�>ʦAn1���xإ���E���W���*ȪU�4�	���,O��N�)��l��P�R�81>�gG�����qgZc��B$Ҵa�����Y�,����PD��Cv�������&�JMj���n� q�9�"�R�O֘�G�n���_�_"Ҭ�_x�~��X�]�$��ǲ�A�3Ր:�%�RТKܴ������4;����Hrt�b��f��r�/�g5�!��nwD�PM�7g��{���_a���s�O�����ꪗEBr�Xn�붣��LeSxZ�_�t���%�v4��������3�.�|������;��+�
�	@��ee��bl��5��wr�S��6�H��00�X����?N/Ř�����78�j�)�SZ��EZ"!��'N�5 �|Ď-�7�X�Fd�⯟���	a�3��=E����kcTO<@���?I�ʹ�I����d�5�gwu�.����n뮜==�j���QK�-i�ضA�C�����h@�+�ʞD.�&��P�*)\�F��rǛ���Q��o���|_7���x���ٴq��MT8�Tr |Ӥ�>�p�w	/%�S�b(ųޠ�3���E����>��X���%{p�4^e�QSM��S��=��������C�s�u�}��F��VA��2�
 G ��w)����p,;jv�r��\�,��ү�~�jӅ��?G��\(K�p�H���z��7�6���f3~�x�/)"X����N����ȫ}�ί��`����`�����?�`u�~�G�Θ��#�X}��J~dq�O��U��2;�`yQG��c�U]��;�6��A�P��o�$�ϾJ�fVԚ}���U�NN���|�*���o�s�C	[&�Q�$��6�y$���q�x3�5r%��x��}�;�����s�o'ڜ=�.��(݁�H�*�;v��?�m�ᖀ�\����� �.���X%#(��/hyk�w��T����&{E-F��=�K��HF�8��ׄ����r{���\ �Q�OW���I#���Py(%�ZȊJjtc6s%�OJ��
yT���4L�I�|\���O8��Q_j8�>�?�����"�ͻ�\�b�Ѐ�<����K�HF�h("-�2\�����/i��G.'�����yKM�GUi�,H�^��I�BY��mE%�d��5����r#�Y���I��Q8�˂Ԭ�J��dJ��_C��0�	(�0Z��,�bڻ� �WHb~`�H7����Y.<?' \���!���5�wj�ahxUyc7|����sifE���� ��.~9�p����2qT���k�J=�9�മ����4��n�R+����0K6�����$/1��4"�P
	�����B�J_g�~¢���Ĥc
S�;7<Zlh����7)��,o����g�B�	���rC_\��ĳ�ԠR/�3�nH�{=q��u�f�V������͚��]q�4G�S�)��XϪ#�8�XS��,B��m��%Ӓ�g��;b�4���8��o��t�`1��e�Ȅ�m3��~M��}^9ǘ���@t(�e��.z�d�LRI ꏈUW�Y�}r�����h�}����p(�X�*��t�x���m����7�)���'S	l�(�ޗZ4�6)�ȹ�׍}E�U`�$s���V���������T�_*�#UG�2�A�M/a�jl����ȅ������&�_e��u.t�&P�#Lĳ!GP��˳=����x����O幏ե#�v,��L}��
�����H�)*�؅U�����b	��)'��K�~�0�U�0���_ 2A�p,Phpy���`�U�×m�呃��D�,}��)�ɶ�ʀ�Eu������M8U<\ഽ�W�O�]\�����g�2�8Ʋ��
�Fv�f��F�Nt��i��J8;>��Gd@��a�L���p��|{�h� �&Jfú�>k��R�
��O�� ���gj���Q�+��;��n�b��D��C����J�lQ�fT�*t� ���C�</�U���	��u{�x�RF��b�A�q�����KĞ<���#���l���5�E���{�>�j�����'�C�ۥ�{w�총+�G����~4�����ѥkΰx�ဌ)&Ҟ�]`g"v�)�pyP�>Ez��vA��O�����OÁ���������ZPJ�a���x!*���� ��*�ɧ�b�^�Z������b^T�k�T�@Č�<*	!�ue6͵E?�/FTF�+�C<p���<:��3_���J�X�4}|>��%���W �R<f{��=�3q4�'߄?Yz�Sqq̥Q:�g@�M���j�>�M��Ť,�!��H�������[�WlCRyP�z�(��>C��A0�`���cc��K�mO��,c#��X�:+�C���U̦�"%��K\ ~*�t��nũ��C��ǽ��}��]H�'�{�D�ɪ����+��^�w?�t�|�������ng�7���ɐۜ���OQ�28W@� �w-;KAzƱ����;O���^b:8�G��:uFH�Ӏ9<m���Pz�uW2�f��K*���e�.(LUA�l�f��S+(����#�,W�h2��\W؏�1�;m�e���e��4���.�� �a��r��ZoL���؋��^*�s��U�	�����oS�P�"{mޤ�X$�첫�z��Ej�] *}uGd酗%6Ͻ ^��u���2�h�NfI���av�N�Θ��hw8��־��jL�ݬ����8��	u�*�J�A<���AY�-��a��)Y�K��i���G]_�o���-�A�%��<,dR}�(��ؗ-���S����U�\����iA�&+�'�k��8�O�C}/��W�#)�������A�'�������{�Ϥ����4Q��ҕ8��"��G���dZ9\�Z����/O�_u~Gs%�C�[�'��?�΃��ة�=�eO���(=.��F�~2)�I��,�`b͗w^#Я}@D(A�xL�bw�i_�t��u�&�0�B)�Ŝ���"��x�y4!�)M�X���i���5�ή0�[�L�8?
6~�J�.�c��&Я����̖�7<�*�>B�(~6��KZxIu�X�(�oK��m����˧S��UP
�L>�RO)z���M��[��6���dj�]�sK�6y/[C�c�d?����Lt�Fs0G�32V[�����W	�][al�9t����އ�� J��r"R�gnD١�8[�&��� 0E��-K��y�S�
�袭��ώ�e|����^�;c��짿�P����rp����\�v��i�	�niݾ	˪S� ��[jc��1N��*p<���	������cjNԮ�i�*�&�+��Ϗφ%�wκ&��`�%����PP�_c�A2��J�
|�hq���G@�As#�oj��}1afѺJ�g���q�	~�9@��T*���82a�,LD�'/p�2� �0s�����9Wkj�D���y�n��ACi�f��8�!ۮ ��R��["��U�ȫ�#��X��40���E�X���p�P�^iE:�z�6})O��ƃ�A5�Ӥ��4s��ʮ兠��n;X�\N���&����ޯ����Y�Ts:sI�t��f��~�U�h�&~�*�0T���Bٻ��D؀�|�n��`�Ϣ�ϐ�kB����"�B���7�԰�-8P�*�f��	dml\&x�I.t�@%GLZ+�=~����u.RxZ��ЊG�O�&���*�I���2�֒q3��+
EW �!)�=)�z]>|Yڽ��wCK�/7����E����)ΌWcT��L�E-�ڢ���S�k�%I�
���jy��`Pf5ߟίy�Y�ħ����P'^�h�^�ݟ����X3���%�J<\_v�k�бĵ�!-8�F]�c9I"��{�.ac��&\ =�T�(ې�a�C��&*~j5jv�u(
a:�#��ed:�F&?N#=ra�-R��q��:�5�!m>��x�[G�؍4��Yk>�ߔ�_d��+Nb�8j�K�n�3+�i�h�)r=`��k}�E���3�����Y��	�E�`Y�pЯP�����3�{�BI��b��mׁ0��U�߮��bz&b2ܝ���9%���&ؿ3��1|�0����jɛ�\��=��[E�q0�ˇ+���`��,C��{���&�<S#CCc><��˵W��R�wI�H'��'�C�+�2���e.r�b�Y��Ub�\�sŧ��	J��"Joi(�W+?�Ţ؟�yniK�3G�1��/.��7�偤c����"#H��$���N�`U^d�6�<�B��Q�!��
�g��}eW��p��	6�Dɔj�c���HԄ���Ο D��t��X�%�vX��¤gL��~E5�ܬqj#߷-�r��mi��f�HBa�\k	2zXc���c6����#��o��>)���N�!��ֿM*ɢ��ZC��e�a�,҃�
�-�1G	Db|��GО"O_����zՋ"Y��T%��K��.��D������:��ó��� _[=Cm�?�+��%eӻwK����!��iH�|8$[-�m|c|;N���M�ڝ+�h���l5?�{OG��|cD���Ϭ5�!�˷�ӻ���]���$���%����D���/}be��	#<!Ԇ��[�髍 ?�e���ۨ>�!�'��R���49������v��L��\�d}�0���LP����䶥��IP�(���C�L;6x6��}���퇢yUSj��6jE�7�tC��m���04̺-��ޥ2x@L.� �.os ��#�jP�y��۴k�I�}����#��Q�Kؑ��n��G��ġW��^��k��	�KwAa=�(�����`J��V�΅�����V3�&���ϒ�z�/U��cB�X�_hn�@z>x0]y�f��Q�x\ 5 !KЛ�~�3+h���l*��0]d ���i�5���y��x���`h&2����j�:���.��0�-? �9wEp?`yJ�Ӷ�9���Ub���'�8T���,>�;����\�u�bL�=�^��
0��u����?XN�#{�8
2����xo:ؓ���.�����&�Dx�����l��
�e�j�ێ`��A2�|.���6��(m�.�~�*�$��5q�]UJ�1U�j3�1���U���d�N<���h�z������������������e�S��7��qe�7_��>��o�mX�nzk�"�� Y����W�u�(b���0�Rĸ�S4k���qx�p9��	�c�6�N��t!V��p���2�4��Ѵ�d�QcPR�b�V�j����<���iƺ�9�{�@\���7?a�\v�+��D��7Z�}9ؾ#�U�	3y]�->?x�XC&;���TC�j~H�Dߖ�h��𨕹����w��=-�y���S���*����e޶k�d��v �9B�O�����t��8�F���7�ra.���"{�SO�}�9hg`��^$Z���V�W����1��m�)}l	�)���v��LU�b���F�$�0iS-�w�3aWɟ��}��a�]�q���u�����Y��Y�<r��Ows�yş���/r�x��|]�fb{�N��n�5���wD_ǖGW�\*�:b3#�>����� <��ˉ�׻̂#�?��Sd�Ӡގ7g2Ë��� xOG
����T��1����{O��:���O�]�Mb#��u?�Ů�$��صvu��S�U���8�?R�k�)�ȸ�S�U�~�C
.�<%����|ua?�s�6k*�Rq�&�<�ČY��UX5�jY��v�w���P�>�T�S���û�'ĊO�K��R%����� ��W�:��\��v�s��d���|�}3s.��y�f��z�K��܆X��{�p�Q�z,�^�ܝP��Y��=�ϒ��
�����7��"��F��.� T7�7gv�W<䮕��� %2f�s����>f��U��~c�>��y/S��S79��吇�h]vןEEh���^iaCE��r`��Cp���W�F@�`%�Y'�g�.ic)��T��+�{��8F]�����]=�,?�:�Q�u�л@�o>�",��L�2u��I��tm�T�ω���Yv�p��*"��m�/VHY�[��c�;t
_[��!6�j�^��K��߾�,�#�^ ��K
gظ`�/���D`G�$�{��,���]tRa�YoE@���Bp���r�M��'���|��7�A�>��������0��Zp
��zۣ'g���N5䠸���E��c�G+���oN�6�3 �n��S����119� 1�~�|�ť���<T��Z'2�V됐�@��D�,����No�I��ܦ�YQ�UN}@{�N�T�_��5���>�0�G^�7uIEeb���mH��%S�D��V��#o6w�O���"e@A��4�׺\�c��pw���@=�ɘ
����J��vO;� x����dRR�t��Q+3�"�>�R�
��C��sq<��Uf��;��2RDT�����R��".+@C���/Wx��.��!a1�C�P%~w�/�[lIr1<=����/1q���K��A���D;"k��k6Z��t��U#\�:�[N� ��,n�3e��t�)�9u�l�G����������BQR�Ђ�*�ﮀi��q��ǘ2��c%��ZG��V��I�!�e�Giq��F���`B�T�:�#�`��T}�&����p���I�q�[�[�YKzB��[Uh���R{]��6y�3̇yK����'�!J�Y�n�;9,�xb���^�٤�H�f�ջ)���$B�!H����n\#���&�2��&a�����z�!T��Z�Vp�<<slN��R\y�GsQ0>�.W���(����YZ��D������
rt��!�I��e3�IR}LS{ɅE��\S�{��k-aK`�^i;��1�w�����旫]6�6��\Pm}g2���:�� rF��\+���\W����х�����l�2~��ǎB�Cд��x���`CHNw�l!A��j+�,�i���(8H��"�e�B������`�=�IR.·�0�H�"?d}%���hbDh�l���Xւ(.�L�d*̆AI��f�����;%	�ٴ��g�㛜E+Մ�6��E�8?+���J�m�P�����!�G��>��$ņ����X^��FV��H$���=n���`���d�(fV��p'Z$�`��8������8�h��]yG	C�K!<1I� ��%�ݖ��9���]�L�� �MƖ�㢪�=� ��=ly��8R�N)lնߠp�
	���,\�m��+���b��x����4%Z��P�70�Yz��Z��i�rj����:5s�X9V`�_�� �j`&��:����T��̑Y�L�e�'<x��Xe�������2U"�n��j�e՞Dn֞�<AD��� _�t��Vm1xkK� pk�2ci� /`����LQ8�T��P܅���c�v0ѷZ?��]6	�ǳ�
��A	0ˡ=X�[[	�4�V�^�"�ւVu5n(
ٖ��t/�u��vW.s��yv����|4�B�h{H,[�r��@G[>�,�BC�M"&fz�����_d^�cu������f�	�>�i��"��-��^�JLg�L��q���,�qL���{�xCugV�A	'�S�oX��z*�wT�-����)L����y�}�G�]0qі�ۼ'�>�Y������*j7�B1˟I��1B��˓�3���橢#Ж�/��h�ʽ�|�c�3���Y�%�m�l)�b��~D���jA�A�n2���R~��`���v9$�=��	��'�#N�������}
�./���9��O
K�{Պ�O9�psKټ԰�������vM&"�
���i7�4���t�z*W2Y���Ng\�:1 F"0[������������So%	�#R��i$��%��A3C*�G��C�Vs���Bp	�Mg^���������XY�p�k��0n�>�z��E!������Y���Kc��Ԗ9b�O-s��a���s��}��\����,jw�豻���y�\�d˃��T&��ɹ̋YWUzTK[�sX��Zl��^�9hb$(g�ÿ!m->����9�ԕ�m�C��!�:�@����:m&t+�?+K7�*�C£�AP:��힡a���M��!?΋�����U�;�����-^�5r?���(��)4�`W�}�-�.�(���6d���o�C5�+*�&ǵ�}p�������{�ӑ`�?����a����	�KG��r[���GPb�W@����O<	zx>��I�g*1,�4�R�U�:"3K��b"%�M%������I��Ȝ9Yh�0�����N��݉�� g���a�K�r�e�7z9�H�U��� ��kƑ�~N������Znp����ęڭ"J��'���nn��hf���܉-��Fg�k��a<*�?��C�ë��v����5�`qŞL�Ϡۗ�kt(� L]�[z?��y��D���#/
� !�1ɭ5�1QGN�7�{�P��F-�Y@]�UUk� ���.�?�����08��nPoy-��$OOQ�EG�{v�qbV�!��T*�� I���,��(L���(�&����
�����s��=v�%Cڲ�}���z$g��c識BN�qYǰY�����1��ٕH�?��Z9N��i�%����K��uޣP*DMK�	�j=m�qs���e��@hc�-Nr�i��=��VFz� �,����O�#�.e4�������,Ĝ1@/�ZD)J�d�wZ��e�^QN[�F���� 9���%�3I��4w
m����T�j�/�d1U���3����0cuZBp���!���-^ �	�v��1ۚ���=6e�'�P�5�öq_~�������u�m�!fs�]�lӏ>�}�x'�Q0�S8�>��]P؈؇��S�:�aV���JCY?��xm���AD��掕����[7��̧ �aR9۵ m	��b �Rѳ#f첝s.j�S&�^�b�1���4R�~|R%�E\]�0�[�/9�u/�u� B*q�n����ͅG�p��ۄ�*��8j�@%̇�_CW��yw^�foE����)Q����>�f�ie6!�h��3^�٘M�Nr˷s�!�0(�S����6tt�is���`��;��\06<-<=��xh���I4��r���镢�,��:���������H2�*Č[O�Ma�r)�|�SI�[6�IB�c�AޑSK�b��Pȶ����+�_}�д�Ga8��R��t�qܛ��ƣз�5��|���O�F|�їv��֐8[�S��G?�������&��s���Q1 ���`W�{��N��F0���#DB�N%�ZJo���.(��p��;V��m"E�Ŋč�g�,9eFzc�i���A�x���]LKQdk��g��8Dt8�`O�f����vB�K��'�'+'R0C"-�cC$a��c���m�&Ukc��+n��%n�1�	5�JY�W-i�F�<�p	�k�SMgH�>x����)�am)x?O���݃D�'����= �wF<[��hgW@s��A"�	�QvƤ��e%�Z@H4����m��l��\c<N�%ekPZ�4�5�U{@c����R�0%K4��{:o��83�?Max�ؗ����p#�&�t	��D6�]�Y8��2�=��'6b.Z7�r��V�JG�v��L��w>ҦO�/z|�^P�V�$����R1AIM!A����k"���^qwQ4��w�7%bO�Έ`�t>�mv��eL�7�;���RSO��B3n�@�G�=[�����4�%tx�~9���p��p��\H�P�Pޠ��-���;ݮ�#@,4��7tA��R9Oo�c�TE,rJ��;dk�\���o��K������)ƠV��g��G>��:�����Gt�N|��K~��'i�2��H�x��y�x������/qN$�96�Qگ��fN��1�Z����Af9�J58����/�[������Q�FP�`��y$����ʳ��6{(�pqP��a��o!�/�ȘuNF�4o���d�@:cR�d2;6�(g�h;�]���r�Ё�,��8��Ɖw�����&r��ʫym��3�joR��x���H4�Ĳ$>/�u�<]�p�WAj�8�
a���]�A�&��FR��OZŝ(�D���b쪑��A�-�y`=��ƚ�s0f�F��Y�ՓqFw��d�<�~��3�����]��k�3���O(8��t4��JV�FdJC��x�`���DFl��+󁤑v�$e�߀ۊ�o��ǼBM�����U��8��A�#q�û����xu`�&H(g�f�J�%nJ����Y[�V̽��Y�@��r��aƾ3boNd�i�\�W8-����(D�PJ���?������[���G��Hr"�hi�%R��ˮ��Dy@kD��_��g��U޳�`�k�q��9�ݠ<�r�h�V��dYr�^���M���!�z�2���V��Z�]RR��m��z�������0��Ǫ(_e%I �g��f,�(���:���a�����<ႱL��\�uw���~T%�g=�f�D{��N����ۃ�$ֈ�k��z�ZC��~��P9�Isf�1��3klt�q�^YK��M2/C�e<~.�&��n�c	OoG����f�}L���T��I�����X����l��h)䚑	\�x�5)�{I�!��Q1o5:9�B���H�-@7Y�B�%pS����C}7�A=��e���KNAW-%��t͂���� �i
."���!:�Ȫ�?- D��u�Q�4��1���6U�$m�A$7P�*�=ڬ���i������q���̶7��[A4�y�=6��5�vu�<�@2u�Us^r[�
�7��"��A=��L7\�-t��jX�I�v0�>�6�%R�ۼ��̃>��R,��u��ãH;��6��n5ˣĘ�������z����=t�>V�W��FZ�/���2�Z�x�N,�o+�ҵX�,ѷhH�N��㆐gRTv�(�X� �f�����<�v�pL�>7�c��P���t×�7G�o,�H@*'�*M�-�~��{���اsɪv��mmjej��bS5p�U��m�b���u�8_�Wu�^�C���'wD-0o��i_�z~�&�f��}��N����V��g%B�QM�g��?��������XsD0=��]o���R��܇~�S0]��`�sz#%���#��^מJf��{R���,q"��돣t1���fi��Q�y⒩�C-�(����p*�&.��p XA$kV���;Mt��g�&��m<�19�4_^�'����f���rΚ���}��E�	6����܉�+~NX-�Mj{gӝd6�l�Ķ��عOWi������s2[�L#���h	���C�T���a�3�-���;���}�b��_��ӷ
̠B�n��Z ����ؗ���.%`b�|q�d1Kkj��4*d�lX�[~��z�б�; �02}�i�����zDȷ� N�
�	i^|*�[�/�;�2�P</�6���nr�F��A8��Uד���A$�����Pp2������v��J��fʄ(Q��KM���z�B3nJ&��X��2Ҳ���l䤣�'Vn�lm!�3
�.)^R�:��
�^]��f�y����o��d��O#hR���_�X�����`��D:�3�t�j���\�������Zg�B��$i	�F���ҟ���*�~��1U�����U�T� �����E!3*�xQ��qf�t[��x`�t����}�zHU�iL5Wu�[��5	�'᥂aOs9��SY�����]������4��cl��7-�qh�q�lA�����Ä�85���C03S��	��0�s�h��4H���u�sz�����D��N�$�o�l?��Ґ8�hGH�j��yZ��}Ɂ)[J}�/��kȯ 	�O�eG�j���mX&^cne��.��`����3�#ZƩ��Y*5�:1+�K^(�ʒ��R�dc���%���?��:[|W��ҙ"�F+�dL�5`N]��t��5y~%��y��.͹3��l���ı��\=@R��:�;��P�q��ZE&�T���胅�-�����,����`�v�j�-Mi�SM��\h����'�oEC��$Rz���%-&+݄�ˌ|�V����z/Q���Fs<�s�a���� (�)�0���n|�w��#��7V��7����ؔ�v�0U�b�D�5	���aib7�,�=wsi��F�"l�����玑���uq�J 4�5#��
풔3��A~�T��Şb��V�淵�3��<���S+ �b����� �Xc�U���o����p�	�1s��/N�]���vĘI�Qn�������Nd5��yF����K��iStD���9(λFW�3���.ɩ�t~Ӻ֑����Z�����&��n$=x���o�}�H¢T_-��J4������$bE�>�`�)m9M#D5�wGT��md&	з�����(�
=�l���~��������V�>=��8R�����D*7�H�-Z" ��dcY�'��ʔ�6��n�a�Z�!wU��frY�2����'���.���o�Sx�R���!ݙ�'�c��B���dt�G��pBA��5�|2�� ��]�Qb3蚲���Qqȟ�{���s�	0�ۋ%�:�ޖ�1[��&���r���/� 	�s?,��}�2P��+s��k*R3���s;�3U+��χf�lT�E�o��ʔ��H��3�[�����E�G_	�4��I�}\ 쏤>�v��:����6X#5���;�����	a�����=�)�z]��o�vg��x���"��2-��^���c����\r�I��i}�EɅX�擺\�3GZ��0v:��X�Rv�f.��?�jfV����ׄ��O��6�-p��7B:��13?^�
I�
�A�*S
h�"�no��7���G�M��h!r��H�U�/���ӟ��tQ������Ũ,��`06.�vD��TI�:2��?[��S'^W7�c��B��:A_�	�[�a@�|4	S9ڿ�$!"Kg�KOCo\tZ���s�����T\0�5>-
��2%遷�³��������N���*��Z��X�,H��F���Zo���,��<|�ln������b2��߱�c���\��n�0����5is�� �6@
7������Z$�w������Mm@��8aɳr�1Z���up����Zս�j�Y)$'?e��6ղ	���^�q��G�0z�7�.��|3L��и����/�o���Z�d��ጢ1˂ȈY �Oߙ�݇�m�Pp*�Dʮ!�փ�������}������d��U�����Bx�|6�jL������sg4�.|h�E��[E��!5��g�sf!y��ω�2S�m�sl���2]�e��æ�+�"Zpl�ֿ��R�C�i�Ռ2�)��,�����{[��A�������B^���
h�6�fwF���k�u�/���Z�������^�+y]��%����䃄�{k�����+����RKQ!�� ��{�GW$�W��\g�,n�gZs:K��7c٫C�wX8��4�5ǩ�pD��|fg�.�|�e*C�*�қ��'4�	�g����ՠ��e��l�+1>�(�g!`���Ǵo�c�"��"N��i�}#X�7F�����*XnD�2��D��EN1��w��浿����ifs��ɉ�Ò��G��mgW�i�%�?�eʕ>���A�k���|����L)���o]�KgB'/X�l�S�S-�w���ZŃ��r>���Ê����{���+(#ts�@��G|�Vq��r�|�2v���o��d�c��-�.�����]�A��7^��پЦ����9&��Qޘ�	Z�?�,�v:GGt���7�ta)���N�-����ƄN���Z;8���)I�G�Iq��;a�	�}2p�?Wւ6�#2]m{9y�$P>����2
~0v�XX��p��I\*clb�d�	�ڷ\�ڤ�j��ZXBG��uxFQ�0�4U]:%`��o.~�V��P�ez�E~��e�����Ӣ����tW{�ޝ���t�ӂ�|<Ա�,0r0�o�ɪz�����W�
M."���*��m��o�:�M���Ч��v�\�-���˵T��lt�ܥC.����|I��<���!f^�2ob��ܔ��d��~��;ZW����K'�r��{8q&�b��9��E�ďő��9&�M�b�=[�K����L��� �РPU�	�C���:��[��?���R"9�fZ�yY9XPEo����y �Sz-;��9��)\uZ�;iX��H"_I{zK�y��-Jꚰ')����*VZ�C�@5�����	K�� �ht�CT�n���:��cކ@�{�g_��ޡv-��~�.9���G���
:�O��b=B�vx	}�<�H��N���Rb�7�n�G�n9���<�� �<4�=r� �UZ�������kc����×�n)�� ��"/��p_�h��,dے9�rP/�#`K�	l�N�ؔ5�?D����["j @�"U����y��z�'Wb<���W͆:;`���,F�)�9���2Z�7�R��ʦ?�l���}8�Ε�)&)(��������>7�3�OU��`WB�ǀ������L�%h�ʀ�~	�ֵ�q�pp>_6h��ku~ -�� �a6�
�h���nV��lb��󲋲��x�z����w�b|!f@])�"�x�� �Ͷ�����wsD\�h��%QS��apA|
��+�$h�n���mUW�C.[���u�$D�5�Y{D�Eb��K��GA�n/�7O��,��f|>��	�� �ݫ1�[)��o��tЌ��?W�R������;�ۖ����������W(-�`kQ�m���۸(��_��/o=nj�3�' _�[>��I�'�c��=`"����02J���ė>�)�iH�L�2�A�>P�h��8�ԗAR=�U �!m�a�"c�����b�
�pjNy3Eemt�������ȥ��\�\C��?�Ѽ��4a���c!(y�����n�+:�
b`B8������I-.��Կ�������;���l��u�H��_��Y�����v��z�젆�F7j��IW	g��v�G�*������Cp�F/������B�6A�Rdc�˿�KK�y��s�a�
ɨ��]܇@!�1j ��&�1A��\�w�½�s쎍���%<Zp�:��޺�,�0 �g���F=&v��1�\�Y��1���v���J@�J�n)����ny��A�\��\7o�q��%S �9�������,C�h���YVI��\̓�@xo,��)�ƔX���q��J���N�*�!v�����������?ѝ��46�b��؏�nY�pλe��5��=���7�,P���Ƌ�}������������l��3_H2nz&�.hb��a`Qoou�y�,����H��4#�Ӏ�07�WE���i�7L�p�������	�6u(t3N��E����I�f��-�=�e<y��<y�Ǉ\�5�����]`�n$��s��l,c�\Jc(gJ�.o2��'O����h²�(�������C�_(2_�Y�Ǔ�`Y���S�>���Q0f�]�S$�&�V�s@)�z$p�gsj*�ub�=����9{��o��X��j��\C	G�A[GB�'z?0�1̩j����,Wʢ
���Ҵϟ<��C�
��{���O0�M|������u"+WT��+����e��e��=��u9)�V���g5��]{���U��1���5����C��L�krq$Ғ�и�=U}׳,{V��}`č-c��p8Q>#u}����r��i_aB4n_X�=��)!�u�=\��F%���cc�'��#:���0�$!?���eA�U���1Nt���`�x&t]56֟����_St����CW�$_zB�^�!���m�PϤMŕ�}[8W,\��e����kN{6F���OB��3򬱀�)�����bY~#"�����[��R`���S
��P^s�S�κYʎ܃;~פ�|�b��9�q���6�|x�֛1����Go�Z�F��*8��<��jgd"mR����o���#B�N�j�M$r
GH�� 	Q�y����|�����z����j�"46�@%	G��-?�4�O�P����a�"
#�2��%p|���a���~�`�$�HqL�}��Xԗ]����#+�@��'Őu{.,�i���ob<��v� �3��R�t2�w�w3hy0'�3��ǉ�f^�}�vߦ/�eX����w�T�{1P�T�xJ w?�Y��.�G*!�%��:N����MB{I�:�Ƕ���R!�}��S�t��s	ƶ�o����0�x�h�g�U�ы��J��-��c���_f-�J�X��Gx�8
u�U�'b��ք��n���[3�@������J%? ՞�J���cޘ5��/Ԙd	�L���5��M�k�tY±�{�!�!
CA��O^k�:�n9��n˘���I-)'��,�'�GvvΙ�i�5X�_�!��^���e�|��Q}��=!���Y�ӗl���gϮC�h.�6Q� ǖB�T-&>�,�,v������m���Mt)�:^�g`��-鼩m
t\뉊6@�'��w�D��5�T�I@�����y�{0�y�H�!b���g��b��]��(�UU\�b����&P�`-�� �l�7]�3{Y��1�3�bs���T�w��\�@_U
��#�� ��͜�3#��+����J��q�x���Ǹ�ԝ��`���~ҩ�A���G2D	�̭F��O@	��օ�n�Ͽ�*���ˠ�/xjiY�\�k��]i�x�W�<��-xԹ�Ak&f�g�$� MCN�"��ÏL�$n�eMŧC�$FI.
ν�.ז�n"<��*t�]oeP0I����#�-��ԋ��^��|��r��x)�>�JsмS����5B��#8�T�������{
\fihiߚ_�>Y��b/������|���ܘz~x���^��yU/�u�c�Q7�&���!SU��>T2`��ȗ�C.�ܘ`H�%�ev�5Q��*b�9"�2L����U.n�X�����s��m�K�]��zYŁ�!< �Qm֡�A&�� ���a�Ӏr��2�(��S�"����o`�4:J��� �Cݕ�b��⿰�0"��URF��.�(����
5�ѳlO>�.�q���7�M��\z�N�S�1�+g�J��O�b�xzg��MF=��.�������}�B�׍����TI�0�r���]�@~�
�8�&u8��:c�io3p�����b�"�贵ph
�H��}���Ih:<vZ�2�BZk�R��u��iSD-*����l���f��"��q��)2���?���c�4��c��Aq�3ٞwu��8� �jC��8Ȅ���?N���kk�#�#c��˺�,����6H�ܺ���N�]Ue�H�0J�#��`�lށ4|�X��F�j���m�-��Iȑ��'��N�tXxp�:��6j���o��5H��}�l�Y�SU�������:�>q稰�V��eX��Gˋ������h��c�Q\�D>R����L'8�0��{��*����r]�ZEj�hu)c����S)sy���n�ׅ�M�cq���~X��-� c,��ˉ� �8Ǫ)�x.и�Q���4�w����+�%�"lh$Dx�ai�w�c�NiV����{��ZC�祤*�愅����Ř�9���,z[7/��,&Vr{�m���_a:�����غ�	m��O�ʖ�#�:�<ԉ�:]�\��S�������5�\ݴQC���{('E	�'�w"ބ�o��5?�r��Dw����s�s�z��>n���}p(��Jv�j�G�mw�<W;�7��������.m�X��w�CP'�o�[C��헲�ʜ�#EQV���<��B�ì�r!�^UW�VX�(!�����Nb(�ԋ?I>�#�{��yMɢ�w+쀾�ټ�k���B
����) �H�?��.a�Ч��ʟҵ;�QE�V�N�Kp'�i��U�i���m��ɐ�g�*|W�	�	X8��N����"��[�E;]���-I��P�;(�|�*�� "��Q�[�5���__�f=�����DJ�$Ѫ�K�ӿ�A�1�=�k	-�I�^�l����އd9��⑻�w/'"��[E�:<o�9�+v�^J��L� [�q=�|�O%Kġ���gX9>ty�V�%�c+���HYF�[#UՍ������,�9N������������,o��dN�m#꼺'#��Cp�]}��N��5I�4��:/���$��%����bE�E�N"o�4�Y���P��P�|(%��ζ(ͪ�v��\��T���X�vH/�aŪba���5����<�eٛ����l��쀬`�7�#��V�A�i�'�g�@��uh����n .Pc(
��
��r�!� ��|�}l�R.�o�(���P��|���y�w��ގn	��8]٘��U�^v���$3C���TM�7��.N%0D��BD9�t��.��aٲ����H�:�8�s�p���Tk9�l�
����]P3������ό�%���]T5D6O�E2e��.;p&Z���ꍄ�7	�ht��z�������9�/B�
����I����lR�	���^�@���t�BJuO0�i�S%�r���)|��v�*��KhLRG�(�ܒbu���-������C*�����'Ah��AyJ��	q�q���a��j�>��d�@^��|���uT��@��3凌q�E1W
ޜ���w'�ʲ%����Wky�#՜�|�\�W��{�)���*�&H�%c''�ZA���bM^
��� ���W7G�%N|)�(?h��ؖ5oڮbfv���Ux�]V��� }Is�颕A}⟚Vť7�s�m;d�Au=��X���7����D�쐶��6�u��1��75��^��������`�1K��� i�\���R�%rx3+���-s�ҷ�{3�3����Z]8�+�8�3�"ka� Vj�΢j{����l7;��_r���6�/	q�Y��?NB�񏽪���LL��C����	*y�W��iE"��$C�}���.J������:�w���A�Oӭ���s��`��0j':tt�m�~�~"1��X!����/�i�{N��d�$��豌b'QR>�;����o����OA�P�.�x򦀗}��W�K���"�mi�&�f���T��Q�iū�e��&#�t8?$���%�䰁�"�ZXi�=��+���c�e7P�@8@�����-x��R7�ϯo�+�v�[ӆq�%N�\OMʰ���ކ�l�1p�ec7�l��@�	�|��p]�)D;��K�������}Y:�f�����S�%�t���z��l�� .dckqv�60�xR���S�x����'a(	OO�4���xW����
��X~�Jg�CfCە�>!�J?���g���3q.Ξ�����2oo�����~�,ᙐYXn���1A8c������~�׸�&B�l�Β�+dz2xP){�cE�2��T����k��O�ТXI�UT�^�Si�~ �ӐH�9�c�Z���m �G�n.k�I}�"&�3���/�����}?��w3�2#ylʰ�F�M�����r����0\r&�&��7ʉl5D���{6�<�&_�qx`��z�����E�{�"�~xyV��K)y�ik�G����0ڜ4H���u��Qm4��_��L�R{@%�@�}��ňI��#z�_�;�uo��'K��T���X���n�J��)�-N�G{ �U��'��I�^R3�癜���6N���s��a2�_��r/M|p_'2s�jc��Ϝ��ٜ*��
{K>_7�\򄋁�c����l�����Q��¥�°qH|�z��SI=R#I�#=Z1R���*���{U�j���z�G�����p����]�;x�)�e8a%�X�Ze� _Y���.�(��8$�!��ᳮŏ����n���opf*���a���)��I\n��,.���)�z�A����l��ܯgSF	_ː1@��s�YO:�S2����6N�r�m�sC���v����$��#����X�g�z�_�N� q\�՚1re���L��x�u�\�*�&�����X�Ys^�#r*��#͎���$��ps���?tv�M�	����>_4����4oL�n��˅�Ƒ���?g!�1��1�i�=�U)L��� ��aS�<r�OHZE��zH�[�r�i�r����Ց�9��3��Ϧ^�E8�5���LHZ�\�y�dɂ�������"$���+��e�Xm�Q㺷oi�C�b��>��j?u�C�5�{:��1���x&X9�V�y�2{3�`�c���ψ+R������<ɸSGy˄�.��r3r���Ā��=�0�d�9�83)�b����Ufu|�j��O�����%�Ž����<?���0^w].7G��x���)?�����!�������W5�;c$(�6_B�,��;��̓h��g3��מ���Y��}sQ��2��r�z�8�kQ&0�=��g�3]��vS�%�)5���h����5�O|�c�+�".�E�lYx��v�F�I�L�&>o�G�{�å8����&2��H��Uq��cI�DC}���i���]�]���+����]�y4?r+fw�՟
�y��ն�kDt�WZ�q$I�vßX��b��p�9�0@��H�o��M�"I)�ߺ��z����X�F[�OZ�Ӕ�+�W��/�l7���)� � c��Q��M67���(��D}��W�1���>K��ҕj�B����d���^# ��.QEJ���9 �ʞf�fmPi:3�E�������Z�f�֠�<B�7�+�B�hU�u^ƼøW�i2��޹������F��X~��u<!�
-N<��`�Ș��6�?-�O`�����F���R�F	���>F0Dv �{9���+$nD�GoP����#��FS��MU�o B�=������p��W�i����JI)�Ow����Ai����K�H����2.ӟ��i��i�M<���������g����H��B�lf����f&^u�`��0v� ��kP'7���|ڬV���f�!Oʭ(�-_r*�k� �3��gz@���c]X�P<�@ �5v�<�Cm�{p��?�<��b!�l���Q�A>Z�f�7/��S�Т����c0��-� ]9d�x��#Cʳ\<�7"� ��_o]�.O5#��/�Pj-�����*��h{��bI��GujZK�W@���F,;z3�)q�.m�"�4�������)�l,�h��^���c|�1_�8�Ϸ(���N���'7q�t��1�%��y��=d�͢jS�w�<�n��oʷ���E�~�Y�`(Y�[����8�(C^U��w|���h��E�d�ׇ[��  ���>yvs������%`=sX:b�31Z���)Lꡑ���6�cS����y��E4 ]ţR�N�Ŵ���r�=��m_@���W��Z�Jk���(�u*ڈ��T��4�b��ag��Mgؖ�u����t"�n��x�;SC�W�s(�W���.j�ibP�֜�����|z��L[z�ӝ���y�� �0bF�悋͝Y�HT����ԮLxI�Nxӗ�H�PD��5e����`/��!؆���A��5=��మ$GC�c
������刜���@K�ē��&jl��]q�����)6 o"r� ߮�j���H3�N�NU��q��GMΝ���.�}�ȽKh�c����{#�h����"������a�Hʍ?�v�ɪެ�:Ш
"�����C�K�Dh1珳����N��+��H�p�N�	�O�e�gB��|��hH���(w1=,F�`�(���9���Õ�	�s5�"���g
���r�Cd`��ϮvY�L�^�����_'	�#� B�I+W'��� �+�r&ӪL%;!��в��ڶmx����b��c�vx�-3��Z�d�v���z�d�L�S�	#�� ݚ�{�w�8s�&�#g�m�'�l��x��8q�OXW�9J�����2�H\}5Ј�d�ͩ����D���>=ﾐ	��9��}� �1U�'l�{:��W�~�/صIP^Ԯ��+i�`��C�X���"b��_6r��o	�"���
ᵂMb�m`��FgƆf�|7��أq䭆`��]Su�Wo�C�h삵�Ef��ø�N�ESmܘ&{��˪�CD7(�=�[�O+�h%���2`k'Hm>�@�bܧ�nJgQ��zɡ�z]u�M��3k�A�B!��qr���Я*3��
�R�[nñ�����8>��J}f���Z�J�jVD�m��o�:�E�to~�P$�G� ��n"�:��	���r�:)U=5�-�g4�:9���6	,�����f8 �]��.��#���o�w�a�UL(9��
DJu���[���=,�+y^��l�$�-"}-"d��4�JJ|&*��'��~��m=JS}H4y�vg���+EZd�\W�>� ���8RO�֠wL�0�s[T����R�0��B
�9f��C����.ߌ(s��2?t� �<8yaT)Y?��D��n���#��q�:	G�F6�IpAsV�Z2�3��:�BPY����5r�()���0Au))C�f��LvE��EeȐf�����e�:a9��`�;�<P��K��ļ2�
4����I�jS���S~� <��f$X�=�:��6�]�G�T���0$i#m�tE�M~�Kϟ��ްL���(�J	�Y�~�,_`Ynθ�}D���%�g[�k�ҕ��۪��;ÁoJ�
8	��7	�]���+T��A	��9��K�!���E�V_���D!9���7�%?/Ǵ�8�W$"�aZO9$��#_{ �C޿Ξ�����EPy+����B��%h��08�?L�Ep�uO���KH���qx	�Rv=Fҷ�_E���A���*Vl��v��1y�N�?��������y��)X��or��h$�I�Z������e��Q�&n�q�YJ=�g8ʂ\'Ga�n�&{�7����gaS��zn0�����^I����G.��ӓA�����$y����e��}Op��5�V,J��&6�7�����Q�c�yF��ZhaPco�5TY�Bt�E)��02��.Xu�4w�e�j��Q/`�:Y�2��9�����{�����8��}�EL�Pv�� b���:B��bՀ<u����h����	���#����L�����)ݿ����8 �A�A�au���ѧV���[�f�gw��A��L�?K������Z���{S���L�R}�0/-V�I4	��r�������1��n~���K���%_���r�L�kİC��ȞH^�Sp�Ǔ����)���A͉�1ޭ��k*��Ӟ
�����-��g����P��WՑ�U�/�C�T����)��n�z�*BO����"��"���
H�l�~�1�[����Jv_[nk���b�93[X����Q+pU�
�a��n��
����5�d�����lv�+i|I���e^�����>2��Pa9��j�_�?� ��ǒ�bp�/�����E���Ui����]�bo���f�h�[)�:S_Wm���3tE)�l!25_��k͈�}�W6ޒT"F�ÉI�]B؅^6���`�6P�����N����E&y��E�IIgO�ua�P�
�l ���y��t�:��L
�~�#g-�h����H�(ۿ�pp�����9��0)iG�\1v$.����T������֥F܉�~�D��x��5э����j&��ݤ��)�z)Ty��Ng�/�?
q~�ჺ	B!f�!��+j���Z*�l�cU6\$5ȓ8�C����ؠ=s���_(���i�.Ǳ���2y��-wS\v:c�v����m��A�	��Kk��^�������̝�^���#�e�h^u<7�x�|Y�)�G!b4�ov�Q���8��&�CnS�����qQ5X�/�4{��t�����# �q�NF~æ�";@c��b�7c}����	2�&�����T��{�f[���9�ɡ� ���:[�	g���{�w�JI�$6F��fv&)~�|ر=���2Z���mb	X�t��$�QP��`��A��}�;'e����n�@Ό���N��[i>y�����-���:���_⹄��˘O3�!}E��X_R���k�ֶ�&[l6�|����&��5�'��l*�*��^7!�B�����0�G��/!k�{�-Gy������ZƓ��U�O��dR�Y=���V��F��+G3 ʁ��!�g��b�����g�TFO����&�xk���r�iSfv�9�ц��=�Z�n�f�p��>!�A?��/�Q��S�0�>K��U!2�5���̓z�:Ӿ��cj���R��x�G�(���50�^N�p?F72S�5/OAf斮ϺnJ�K1O:@k����d��J��9)��&�כb�[�I��Ά��u��6��_R��,$ڳ!� r7shS�����X�C5����ң�P��O �AYn Y��ǅ4U�7ݑ��l�5e�q�Ծ�c��8��Zى��.��K���z�Ԋp\�Qg�>j|� w�IAXnh�|���Z"��i��ժ��+-�M'��hJ=��K��{~�$;�fE�D-�+�F�]*V�b��q_]�)Ո���Q�ϳ�ߗ)�Gĉ�v���;P Lf�W��7����1+y�<��b�_L-�Z�[��#+�<�Y�(�J7�պC��I���L⍅K�1�@�o]ڵ��hΧL�M�`3��ʘWDY�%���|>�z4�>��AO�NM\Ur,���a�']�P.fٮj�`���Lps]�"�zп�휑׈������/Q��	@ �?��l)��PO*����:W� i����b1+�=��F�>_���F�,U����"Qa&2#��sԕ�%�ʗ�.��>����N���ZХ����q��-U��i�`��o	kMb{,���vz��`Š�\����x�9� vR>o��t=�ߥ�>�<���7��1�|j�X��������N����@`�%͛)n�>䠧��3��)\9
.�:|�s'q�[tg�(����<Q��^��Q=i���٪��ԉ��7�����{���]�Z~Oh=Ĥ	U9j���⇐�M�z@S�����_K���=6��o�Ϩ��ؽ�'�^�g�s^0	n�C�EE�r�m�i)��t%�������b�#��m��]2u���nM����Hb �h�1�)��R��xn�(,�r]����D�?����{��]�ҋh�fxV\�Y�{Rg����Ќ}\�B�:D��{0+i���,�F�+Q�\��� (�K���Z٢�Y�H	��V�����t�v������_iБ󿭘��t{�ܚ�oT싑J��>�*�؟�9���l{:.-��{ ��,Z
���k��p3�Pd�0J�����ʻ����o��CD�}�ls�@Uq��an�_ \Q��(�����E��<QL��@#V�B�X*��z"��C<�+��fm���μ�b$�6��$弻w�7ڭ �m�A64~n�Sgj��D>P������D��I6��Q *=����z�c)Jن̹�؊��ڒ�dj��X��_]�uVZR�;�g�<ݙ1�b�*���]l˄�r<��w����F���j�n{��h�Rߵ����z���壔��">���ov��p���f��hDz��k��%���V�d[�L�
�m�$��Yܮ�w�.�7��^�fJʭ�a�5�z�Gx�*n�e�@��4k���1���F�6���3=��[���=��W�6O��KHMܵ���okv>��Y����lAzW��e�ǜ�>|�b�H�Ո���.��Q�7B�ӂ�>*��59/����4ʝ|Ϣ�;�˪���I@�������m>K��Q�����ܵ|�3������\/k�M��dJ�d�]�n�z��L�5������f�fZ7��vG����-�
��e���h~G�!�sf���2^@��������ڡ�:�œ.������|�I���pO'�!F��-�)q�{�0G.NH� Wַ�~��8���n�PdR�G�GF��Q����B>^�>��h��*}����U�_�.!��s}��ϳ�}��V���{+�~<vU�w���2��b��ٲ*ͥT�T]?JQRc��g_�E��[3%������o�:�1��3E_�3q�v��j�^�T��eh�b5dM����u�0����squ�u��g~{�i��v#��,Y��	4Ŧ��8�i��4v�FEl-�����>�L� ���.1>�q��� O7��9I�<3J���k& LC�U�^���I��h��S �zI�e�S_I��-L+˘��!7Iր�����U������b��'�D�rO���x��M��,#} ������w��ꡒ��Yb{qR�ݟ��}�����7���2�Kl2ef��T���b�hI �H�ѝ���<L�oz%>�X̗^�ԫ�����P�m=Dwg! ����wN��>sӐ��)ߌ��C�������ځ�HHJ����++� ��C�6Q�fmꯦ���M�Iz!�mh~Β��Fo��Sz�i^|Y��>�� i��p�*Z.>�g�(�F����Ja!�����h��/�:������[)s�R��!K��)�O���_��#���D�^䯦����f�5�*�t���2�A/]�,�Մ�����o8y��gh#�p�u��ۜ��:td <?,��4���50k�B"0`[W��n2��_�y*�
\$c�Xl�-&��ITpMd�G���R�>r�Z:�Cz�I����o7�~���̠���K��	~\"rf�� �!��!u���>pjk��l&_��c�c��m	�1.�z�m��^pT��	AjD4�!*քWq���aw�V/y�YSi�L\|���7�Ƌ�Hw��p�����㳞m�(e*�.}e�,iqx����"���p�7�J��q<�������phKĈ ��r��qԕ��~�xB�G��l��#�7�V��'pCн;��io�ȓv��$�:�-Yi)G���#,;���h��$�o�b^<2�#��7�E�7��N��+_���qJI1~^�K��ɬs'w�����<�/;-
�T��FG�48%f]T�)0�ٞ�h�-���L6�V���D�V���%��cI<�:֐�����!�ԣ���:g��@���İ��`�d4���=�BQ5��_s���u�B�}�/���v ��{N��Z#(�VU�2ޔ�u��hv<&3"n�_G���W�&a������}:\{�3�7�~�\��p	}���L`uxʽt�u�!���\����>����UK��|�Vq��.1���I�c-��8pA��˪�)G�$�r�˒�wI���7��hc�����/��q>�A��s�Bzu���e$mN
!�m���h���)���6�t�Tǵ�fe���;�?"{��Ә��R�eȫЛ& �sr��|�Z�:�N��=��mF�Yu X��|=U���^�
����'�2oU�֠}4�5��pG��9Ja#J��ru��vaW%H%jy8j$��_
40�@yc����wo�؏xu��|z�o��\�1���Y�{Ż��,��m����p��3Р/�W**��j_�0�_lEߨ��[��O<JB�6l>2�����"|>����1�-�[��A�����l���7 �P-���Wp�jN����N��hq=��e4(pq�8��g� \��)c+�5;G{������*�F�.�)Qƿ�D�Kf�Y=�<���ʰA0ݜ�YTf4�+�~|�-V��)�l����� ������G�R`�:�nȏ弾��9�r���U��J6U��K�e��k#_VC�9���?ק�eH������>���m��c�`k�Ġ<x/�I���f~8�u���#a�e�",�K��6��/AO>~�h���X��G�h����g�*4/8Q�Jghy�W�C[Q�x�������nv��%Y��l4&{ڧ�Z���I(D�����,o{޻o?{����NەCt���0�Df���EڱiD���yy@~��ĉ*��<I�o��*��LI����OMko<CV�sэ�d����y ��Ab9���ҏaKt34Fݫ�8Z�Z�6�b�k-A�虝�{	�8Qܹ_ᨀ�l�#�B����߶-8)�:Dj���t{��&Jt��m�Q��bBc(�͢t申��#X�FHoa��Z�`+l�A�o:�X-,E��%��ل:倮�������h%\���X�ew��O-��u�dF�.����ݕ����-DiNxP�:�ھe�?�S����D
�X��>1n�A�!�=�~@T�q�RS�1�by���%�F�N�0�.7�����%"㤬=�H��Zv��!Պڽo���j(�d9�����}�d�5����B�6��)�tgO���Cd��Mg�������V�E�di��I.�/�]}z�ȝ"��f�~H��=u�
9�R�^"f[F��:Ä�}��koU�[JpHJw�Y|�&�p逕���kTO1@��j�t@b/��.�I^��k�9L�%�M��jn����k���u��+_nt��Ɂ�0�8�1[
�@���ڳ��Fg�sj�gU?�E)�^d|>�И@��*gς�G5���/�o�~�������0F�q�j=QG�;�������x�ޅ5�W�i	>�� 1%��/��7��
e$�@��_���ȼ)T����P��B0D�>�2̓0si�����aʃ6�U����nI�F���t�b=�*�!�R���-�g	E]u�\�����3�_���J��0��EsJ�^h���e-�>�z�A�9��g�/ou�_	ES|�Њ&�˿%�@���kV���
��ý��ڗ,q�e�Zd�I@���g<�2�����dm!��h�?]ǵE9N�t'��!�3I��w��ɋ��S{Ֆ�V���'b�<N�Y�d�2hfÐ�����wչ{.�y�oC2#����uw 7�4�L2F� =C�dĆ�|Y�`ć#*�?�mV)� 2�$�_�Ôc
H/�ꢕI��������+b�-�=��7��[`D$�7�~7��y��ʐ˴��NI`,��̰�u�l�˜�4����/ɶ&���:����bG�'6l�/:��E���R1�Ԑr� ��u	FX��ל.��2�\2�}��{�pj��-|ƻ0j7=so	�r��&U�!�T7n8W�j�l,��W�98������f��J�g�ߜ���5Z��@V�&G�=����˛s�*lM�Lz8$Ҧ��(�w%Xu$�<Z{T&�4��b�_��I���8�y��N`�2�o7�J��+l����]��5oiX���Ě�n9���[\����g3T�<Ay�w �X@���Nz��>�
�_��;�.���u��an�A]�f<�~�_�C;�^I�{���qe�z�S�٨N�$�����,bw�Ze�}���&Z�o�u��{DU�`u�6���(�Ď�t4���_�vv	+
��M��N����{�ƀ���_��(ƛL���l=�w��Þ�4�!2�}*_�h=e�� ��/wm�Z��mD�����/!a3�-���/�#�zh��:l|"�_�{"���#�����~0���4ܟ�jڣ���쫑,�ᕉ<��Y�|�҃�Ɔ��]lY��T*����2�F[.�1�TD���y�z�"��V�����&W�<��e��-_\t 0F�;����2�G�Csk�P«m#RB2<ɤ���E�2Ձ�Xj�]��T�H�}q���dm���h�Z%"	�5'��d��_wL�/�P�}G;E�UP��Ք�K��7|�[�=�&���e��tH:K��>ј���|R5[���Z���w����I��X�D�S2V����/��yɝ����{�m�!�br�aS<u��r#S![�&�n���]�����=����ex�q�m.K��d����JKN��|bW��� �"4y���x�-����:�_�@ևZR�1pB�ػ�QrK �dD�Ҟ�c(`�Qb2E�O���ڃ� +���j��
�=���ٲ��L\�|D�h��R���Y���νUv�Ҳz�=O���f�{���
ʋKN^�H��s<sr�Z6�^��C㓰=���+x�K!	S�펟�F�<B������j����=��Wa�� �j��zC)�I�jlt�
 b�����p�����j�qB��]��
��y&;�ٕ|P8���C�j�h�N�-)�q�p����	��ލ����1��3.ׄ��S�5S�Mbp�D���_D���b�0ȭ���")@ �uX_ʭ�=TA��{�PWJ7�������N����ΎF�9�h24KmK'�������
*�zS�X�N��Mc�jWo�C|�)������̣����"J��ƽ��u%}���f����FE��R�d����P����C�ɟO�&�$fŋ��6C ��N�r��Ǜ�(��f�T�|$!V���1�a��o�LR"��{�^��!"1NV9����;ս���~��P<�"��*ڼ~9�^Y��o>)`6�D�G���i�W�M:;o�2����%������0\l�,��5Ȫ7�Qy׎x<���)ȵItN����2���ݽsdJ�r (k�"q�H�+zfcx{�Fr���**�jF4BՈ���ci�J1S�X��_ç�� q�D!G�3�|I�k����k�VwQ�G~C���>>^;s�3�����4�.p�W��0
�4}��"����)���w܍����k؝u���	k�f�$l��}`��e���@��w����h���)Ʒٌ�$\J�b�	����bƀ���(�Z�Z��ٴ[��H���KȀ�D�$�\�g��>���W���,Xf���8鎼0�0�e�RﻴB�z�4��ogB�������l�d�J͏����8RLE�$e�65ψ�A�'[�n��9�F-�'�?Q����9��RM��4K��;�@�y��D�'���(L0�G�o�>gY�)w�-$.�ZB	݌k}�oZ�rOtt���!��"�u�Mz�أE��<����%*����)�*�f嬴g l������v;߈������{1O���&�q{���1f߮$�طt;N��rBj'�*S�y�e5I���X��zn�p��J�X��� ��,�%k��m0'ݍ(������6��&�/��������'����S�&�=�|+�:��*�&��N��4(�|D��
n�a��,��d��s�>�FH_�ݙo`:�jhl��3O�hj��R�]��j� �� ���W7x�[H��}Q��8�Oj����uJö5j x3v7�?�.����I
����F�� l�P��ǹ}8$%D�9�\T� �gQ�Rh�Mt���x��������iWl!�[�5Y�Fr�#a�w��a���5i���r<����(��0�"�ˊ1�+��|�#V ��v���z��JV߈v(EȦf��D^����a@g}R�N�vz���Ɖ�o�CA��zj���� �%g�u؈8����������[�h����b��{�JzQ���KfҩI��Z���h�9��ib�$Z�ƹ���&o�m�0~3��ç����?�$$N'�e��V�]�w��3Y�\$����\����ZF�Vq6����)�4]�~��d�E������K�"�F�O�<"0�/|CΊ��/��M8}�m�Ɨ�,Xb�H���1��՘ښh�\��KO���T�\ׄ�1���;��W	 ��g�F���:.��ڱ��u��B�C@�������)01��'��[�J�q�/hk=��CX�yg�w�4�|�*؈��z�q�Y�9'W�$~�ة"�TS;��[�s�^,M;�������x��p]���J��g�/�p�)%O��~w��J[��_B|�!�-��4�E��[`�hR=.�\Ŏ�-XI2���B�aj��#}���&��"��k�	��4�Ϊ����!��Ǿ୎XYd�,�9���@��W�Zv��a���u���))�k�P�����.����:��`l�yЏh/�$�o��n�Ϊ��!�3�z���+�����H�-����ɃՇ
�>���$�62<DF�w�֑�P���ƷD�X��-��U^�`Cy7��3}��&,~��M�l;�k��*�Mi9�%r���ҿ[t[`�C��К�ҧF3@'�Y���!P[����K'��� R@E0���/��!����qv�X��N�H�.�w��O
��:ҿO�(�ɷW�UC�b��٬$S��1ȧ	��r}�D��U�`h��e���z{��[_1����ؔ�����`I
Hp��*�	�C4��A���E�0w-l|KY�����AQ�r�X��2�O��s�}�:�/[�5Άmhz~rX�*)\��S�)0+.���X9sT8��*�����	�mk�ZJ���lH�sE��٣�8��R��h��6��I�5'b��.���.�f��;�	��F�7���pfw����`�I#��w�|t�r�%6j,���,�y�C?u��AX�b��2��=�Vum�tN��T.C��]*�Qx1��(�Ԛ򲅰�0�U�	�3�������E��OV���a�`�&��q�~,P��Ⱦ��]V9�gP��g?{���׷O����!��HiV�YC&��_�+��m��P���$A�<2�%���%��!'���ݧ�Co7���e9ޓ�^�T��ŢbG������|�pb�Hl��������K��1N� �zBL��G�vnF�$!�g����)Ȏ&:IH�3U�%�8ҙ��u8���`�P/J��q:�Fܶ��R���*��7��������4OW偼q�AF@]��^~x��;tH�� 筓�H���x)�9d�t)Bw~K�g��(S+�q�~I����`�J�)�OB����[7��kq.���$����!-�I[��(�.R�a=�{4|���ǇZG��U�5��7\��+�z���D����˸�AX�9�5�8������C�pBi��r����7�( ��q�Cj~]�O���C��%����'�ֶ7� |&�b�k�r��(���u����~�_=`I����(���r�j�[J���:�m
��-vD"�QZ֦$9�Da��b����0��JԊ��/!�"���:��W|��y�<�s�����X��-�':b|G��4�N��i��"�Y㢉���Fd@BJ���L�C�ζ��%�?���R;�gڞ���aq���/uvk�7XM���o����4ch�i��C�젔�U4Ҍ��͟G%���fq�4T�X̊3fA|ƞ{�te�g�0]k6ΒzmkE�@��OB��ܒ�F�%ޣ�P�k�#c梤��g�=����D���}ךTR�&���&�LD����x���1M3?K]��E� �3Lh_i��FF��6�w�^��ü�֑����Z�q�7,�`*J�du��X�E�!�%%��\>3�ᱷ ��\r�̹�� ��W�v��
c�C�@T���
�2[W3&m��(Ց�N�{���a�����x"��u�d4�5`ngv�v��Ev�D��x��\FE� jk�29N�b��̵fe��?�3�jBlG��]�Y�j?Fy��5*��Тo��ˎ���ᬞ�č�z�3�{�ĉ���3?�C���rҮp�u�W�Il�]Y3���t�Y�v&���\�1�Oî�[��E�%.��wAK��,,��b����R�ΎO4$�$�?w�q̤�(fb��q����
;���{P�iG�A�yDx��y:��ەB���uX���#��G+L�^�*z�m�:~em��lR�FÓ�n���Ws^j&���x��h6��X4>z�r��F�Al�]�#�]�N����*n��R�_t��/�&;�|Z�G��.����q$o.�
4q�jW;�v�Tң�_wwj=*��s���O�a&PE^\�in֣b:o����/}�����B�?��m��)� ��V���S����$�o�,��>MI*�1�坥�8���P4��J�F�>���ho�<�����yn/6c%�@�,_� ��܃Y��r�?����f~�{�(p��嚔K�]�s���ŉ������鎚�z���k��GG?��g�$�c+��u[��I*���<����	A(�x��m�����'Bml����~')���i���V�	���4��f������PεZ=ΧN��I:Y8�ǎ�MUgK 7��+ ��t�+�K$���6&�*�sh�~I�����A�ڲ)D���c�\UH��l�����m:wiMJ�Em�?�� ���Dk2SU�� {8P�t2�+�`�E�(ҫ(�h�Y���V ^4������Ǻ7C�X��u�C�ÿF�3i��Лk8����ޥYC*�����%�0�
�gd#ιӚ�qrCx8����MW�����ݦZ�|��CӐ$ �p���,
���0�"�I*T��(� �.��s���(�=����&h�a�g�k���F 5��ϑ��	ޫ5��da�?�9�����S`(z���s�����vͮd��a3�D.L���:��d�t�ߑ�{�p��\^�x�G��'����׃Nf0}�b�G�8��]au��|�	#
o�N�0<<p������(�{W[���F%u���^c
�����D��i?ҭ�C���Rڼ�tG��>��>F<@��u�Fg&ҋ��텱����Ջ�c��ſ�ҍ*3 �$�1�H��̃Ɉw�L�@e�{�j�zu�\��G~����u"��L}A�ca�
���k��/:(���U<{aaշ7��O����C������9�Z�����{"$����[i|�z�ؗ/��
}=�����-�V�gr�|�z/�����t$��4\�1D���xc��!(N��9e���,���_���?��=OM3�_�zE�<���[D�s��,#��o$�4ϭ�p��Fl|�b&=E���2"�bw�7���fO=��7| g\�Q�+Ȱס��������]�*���mN@/�����!�DqXz^�����W'�+]��$�mO�+?�z��*0#���ՙE^%�<�����$]_3��\�H�G[u�,}(L,���3L&[�ak���Z���p�P�q��ά1$X�ޑ����u�8A<={fv�&O�8v���swŅ�N[���\�#~�P�M؅��RZ?�{آF�b���nkXX�������������tV��
�W�K���1��񆡃T�[����W�B�ݧ4-�����0��Đ�f��d��B��ueV,9�/A���s0)���E��#̢Z��3�3�)��a|.���E}��� �����i�K��~rdd<Ҡ�	b VhU����D������l�Q����h�p��7*�Ş�O؅i��1eλ3Y�c4�Y��N�~ ��� �Mz����D����n��J��<�>ɷ0���6�TR�8LF}��P�Խ�>o	c�ޔQ�S��
��f�r�6!#恧��n���;�x���p]
4��Trkۡ��o��?�HD̬�����2�J���8�],�z!��o.�TI��� �؆W62#t
:
�j
_72�F����~���mgd�D8�d���Nˁ�t��������*���7�ȺU9O|İ���"��\^��7�x>f�`!��SH>��jc�Z���U�Js�������������G�
�H��� ��7پ|-���7c����t'�P�!�b{�ѻG%,�vh�0��SJb�f��w��};�o-�S��z�m�)aJBr���浲��mq'�
n�]�Ąs��T��Y����P��ou��%_X�_/2e��-6�-e����zj`Q
9��0'�.tqњ�=���:4�pc�M^���~���U�̥����CG������j�����Λ�����b6��ܢ�1a�]!�7���!2.v��:�@�ǗIN��ՌV�7i�xջ�[����U߈C����z+���%%-.�%|,�;[Y�y�k��{�r[@,a����i�D�9�Ԫg��q�R���%����8E{ھGm?wT��ߴ���c���:�%CJ*���զ��϶�[=�aA�\���A^�X�ZC�.P)e�z��Q�Ϸ_���b;6b"�cމ��2�Ǿ�𒢦A-=���#	9��y[K!g��a 9"�P�d��O:2�}w��^x�(Ƭ����<�90��fӰJ�p�`a��&�+q>s�OB��:'��(]�	�C(��A0D\�����`'^�r�,� f��o�L��ℑT�	�s�qᆁ�{�n�Sݚ���g)A����),ZF�8�j�#���|�f���Y����d���7����g�P��\&}`��R,+SL�Mi�����䑉�A�k���t9ֈ��
�_^��\d$����l�Q�6�VE��[�H k�4��ШII�5����Y�v�ZH��t��"i bH�OwE}vIr<�[rĈ��Z	c(�.~�E�(����.v_���#&Ӆ�3 xKR�Vn;\
#�C��ā�ٱ��F$D������Jq3� �F��}X����͇�n��s����� ������	�ץf�y��[�b~g@,��yV��	D������!���s��5Q��rs,��ۭa�#M�:ཷ�(�aӤр�{�8�+-�zW�P]���^̩�{��
���#���]LƬ���U��ɔ�g3k6��{���*�nw������3����]�!:/'\k.N�CN{H�c�&�;�mn���
_� �L�!���?�UrH�II�*��4&��ZݶTh��� �='�'ʼ����G9FN��Y`t�<��B�%|Y��w�BT�?�Ț%����V6tU׍3M|!J�29�]g	e��*��y�� +q'y�����\��p͡(��mT���k��Q%�*�*X^����v�&�ߠ�)��8���t����ʸ��V-�H�@o�-A�Q��Q���b/+��������!C��y�A\�.�S��h�����HWys���|�<fQz�X�7��,�pN�e�Ni�/����pU��`�ls���r2`{ǒ��������Dv&��R��1�uTr+���څ�e���X`�i����_�^d�t�RPz��Ѯy5�O[�s�����Q�&����88a������c$�I�����f�;�W��]h"��?�W���x�d�0��IX��f���P.9h�pU,�1����ߣ�i���bs$�]�?�{����-��/͍���͖��|/	(���G�H��̝+��_c�FR�<������k�+�aő�Mg��E�����~]=֮d\-p����@�Qee2A|�k�9szqksy��XY�V"[��(����Τ��_'�E��F��x��R�[m�2w�_��-�k��m�..d�a�p^P����b6���=�V�kò�ZdQd`��z^V�}����:I��y?������^㟳��R�<?p\�'jq��H)&vV3������|�1�A���U�Z4�Y�y�<�k�B��&Mg����8nqS��'/���p�2�1|/��*�N)ǹ��<����W��/�v�P���\+1%բ]S6�����A���eo��z�3��)]J����'�m��� ؜��?U�)�8�:mһ�lȥRUC��/�Ӽ�
��v����B"3�Ne���x-�N�]�o.u�ܚQ����q[��K�8�����m"wC�~ѻ���8/2ג��b�#҃��� c���
�W�%7;�*|7�WS�A��޿ZL�]�D��T[��Obef3��ɯC������DQހ���\p�vH��<�O�?��W�P������
�'x#�����"A#�=v�:Y���t鳀���Z������K�%����dO�
�����H{�zhf�.�nX���㑇v��K�z���}l�n�ƿ���An#E$(�dM���73�����qP�5�q-�Y�'���n�d^HGO?�FzQ����O$��F�~��.e�B�u�7�����>�4�c�k(!�*�w��H����R�("� �����r+�J��C)�G�7��y��O��=���Q�v���6-0GQ�2~l�����������l�wAD"�e��7P�Y�������PhJ}�ѱ����m["���ާ*h/R+����Hv����8�c�eJ�4W�R�T�8γ����B�+�1���+�>���3��4����d���_,�V����ZW2��[rL\�g��`h q �$ɝHe���%��'^ ����\�wq .��W��'X���W+� #1��o]��?��iQ�Tj@IE��R������?���8�Sk��8|�:�_������Z���$�p-G�b� ��I�F�0P��@I���Ld�G<���e�J�5x	)���7&�=�q�ѽ����q�!��V�?]��K,�e�EV<x]?7�s��3բGU�� �~'�r��\�EvT�,#m�o�w�о��8�L���E��&���?2��'˝��[���	{?/�=�'h�}��ҷ�b����sI���X/@�Δ!�������^vh&O�?�6?�3aq��T�@�ɳ��w�Q�K�FOyG�Ly:�Qg#fO%>n��Ȥ5����+x�'��J��=P	@�aW�SĐ%x����������DB$ʝ`�x��|���G6=a�#h%Įe��A���V��r����`ep�.�I�|�h$���)�hbvUc���t�;�="�k���\�:?��S�|��B���8�������@��{�]����݃����z�溇1�{�m���OFPwu5B��{����PE
:��h�B�võ}A���?l�jﮚ_��6䥬�~^.�M@���TrQZ=��/���4w���/4�C<�%<W]��EW��*�ս,R����2o�)!�);t�t&DZǤpu�ٔ�%|����]�|��jh��̘8���3��l'��tf^<�������'G$h�]�qĠ��^��7����s�3Me&]	��#і�n�~1[�f�:��aG|b�� A��`���A��bU� y�~s#�P��!l��bj�xF�,x]}��+���z(��g�k5o����;�SW��	�|F����w Al)�B2�������9*�mz�g�\������#{��G��9l�^n�wG��T�,i�K�֔�/���b]��z5!9z,��8�x�_��=oہi t�S }�ݘ>����/(q�����-ߺ�����X�^ҙ��']�����d%8F�o�z�<g��U�l�b*�Wd+pSu�ަG��f
��t�a�VF�&�R��YK�y::��8X��X�e�x�J�2��z��jOR�����P�L^��8�_�K��������S�⺇�=.�?������^ߺRQm�ߵ�Bs~������b�1.�iN����z[xDR ˌo2Țq�R,9nڠ�� ��;���	����g�_R�x'Aw$j���r��r+���J�?�u($��Q�|{] 6��#��@JI��[z��DP�D�QD{�o��7�� ��/�.���7b����ø㌭��/I;C��n@�ߵ3U{sh����A�Aͷ#D�;�f��I�������SEt˧����K��Íg�q��LgXu:kH�]J������k�A6� ��$0s�_���8^NQ�����Br���(�Z6��|%՟�D�啥�'���{�>��x*��f����r��DĚr��D�>�T%���I��ص�2���'G�}��t��@?:<��Y9�H�I����4��2rH�'���B���8����fG�i\6���~i�$C�jQ�-�S���;(�³�mZ��lsF﮴x(�<#�����ܓ]l{��*��Zц��sg�	����j�5��]Ŭ�ɉL{�>�lj=I��Җ�P��syq�0��2��m��b����1��"R0v1UH~��3LeŽ�T���쐰?���^Դ�xg̔�7v���]��|m�p�Ω���g}r��x?o�n� ����v���,c� ������g���2�zgv���ޡ��5���ͣ�_d���0Y�;$3�8��o�G�n����zJ*i��)D�iMaHN���{7o{T������l�d��$��ѧ�21����REI+ܟr��M�PP�#pʜ[��DB�r�=ȸl��)G%f���Kb���l� E���W�Qio/�!Yp�qS���S�#�5���$��������WyuT�}P�D$��N�OV�U,�1:�r�>ΛޘI�I{����z^]����&��0�o6�r�r���f��ADO̎]��?��;�`ꌫM�%Wi�J���c� �|Xd���;����ZYW��=�����=B���+K��#o*�������i�������¸�� �!�sNWv�.���,�
\Ez�=f��N���f�Y�'%~��n,Y�gQ6��1���.Eg;ʆ=;��"��)��.Օ/�Ս�'�cD� �����IC�E�2ѡ=���o�K��R�����U�1K�>���UO!%�94�ٓ�����m	�=X6�BATe�7�G��f�ѝi�FIf�_e�.�ag����ͤ�#���'���V�����F�v2�h�k$e{ɕoYk.�R�AN[|������s�[ongML�+���T�9�|�b��N�Y#	�r�3��Z�{z�� c8Ď��w7l����t9��ŗ����'����N�i]�p
�o�;��-�z'���!ZV�E��z��Sk�"�tb��G�Sr�+r6���GΞ���N�l��y��D<C�9I�����J��������6��[�oH��zv!<(K�g:H�#9�b��y���>G!��ֵ�X�I�m�f�E_��a7#T�/�� *�s�n��X����c��/h�=�Kt������vPߺ�R)`���G!L�Y\� r�{Y�-^����r�H���":DGϖp�Z��	�$�<�R�$����}��!ǧn��-��o?6�|�es!~�X�-ΥYL��N|eٕ
#(�g>-�	�X���
�f��ȑ���}{+�3@��$6���%�%
�s <m�Yjz(u�wn�;@m�a)Ը���$�B͠��~�z7b�����(��3�ԯ�i?E^��SQ:��"�V&��0&0�W��T�q"8*�6�1��}��π|8�^��@�4�3�*1�o�o�,�f
ܕC>��:�p'i��KeQmni*��&� nVx[u�q���q�����W��.��v��H�8\S�Ot�"���'~wm~L;"����\�WUP�����T&/>��UQpX'Q������
N�fH�Z`��dD|��<B�y�c{+�aAF��?C�����Ȏc�-A�����ensO�G�;�Y?�]٠͐�6�"p�i�9��|���n~���$�ƪ���]j�m3ܹ�-�-�c�6��7����x	�W���M��b��9�Д泶�_HK%�3ă��&Pl�)iO��wC�C��Y��q^FT�z�vU�-�uf<��P�Z��Au׎(X`h!v �z��4*£K����=F���Q�s�Z.4�m�x���� �bVb����tyPw��4��m6�-�pZ�3D^�1���o�k٨ Ͷ0�_Y�R�7M���;�2$�ͰD�4Ӳ�i!J����tܞS�&Zu�N@υ�\�F#�N}��jE��Fz7[��?��_��I�h�~��GkT���T��F��M�8��0(�6/-0`�L���d�R3n�S���=����K��$��<����z.6�������^�X��N�8�i�y�b ��f�M]Ԗ�@�5�T�kǹ��J�ڶ�����s���.q+���ON_}���:0@�ݲ�;M��"�bN�Ǵl�Q"�|��Ј���qA�C�8ʋ�5@�j�a�i�9N�DqᎣ�i���e(�nQ���e^+�����#�U���v���y��3S�&)���W&$[
޾S;��.J>�9/�rYx�M���E�`�L7ӈޭ�j���>�**�4_G���^��^���`Mi�״�5ҟ"Z��͋M�y`��|��k!ɇ��EA��*C���gׯ�.z/Efh�YWRh=�r4���
v �L���O��ْ���;�֮^�K��������N-��r���0�=/Ϊ�E�e9��X]ҧ��^�F�vv� >�H�SV��U������b��4������kL��n��XD�� 
IW�2GD�NpV�Y������e��MaXw��4Ϧ���(`����Ɠ2���Å9��X~>$���z6��=a^���i9-�"� �[V�nǁ�������_�����
sR7���-{��V��hCZ>�Ha��[H���ӾV�:UT� �#t�))xʘP#��u؋-d�|�R�i��j��0��}]+X�t�6��N��k���B���Ij�c�D�C�7��q��A�"p��=4�o!o�M3���)T��x^A���mR/A<k�� aܡ@e��lJ�M鼦���aL��6�.�~w��9���E�I��ͶA�C
����t }Ht��>�\���K�:_�u}Z�6+@��4U��0�ߕ9��4n�����U�O�̖�mw���b�.؃cgn�|�W��
*�����'s������5[��tY:��p�'P�@Tr8�ȭ^��H�'��N+F�b�)��8!I�
��%s��(�I�4I�%fc�O�<	�l�)���ۭӝ` ���X��߀Đ�-#���sV�����U��F_����C���X���LX�.�&%W��#G���1V�r��P���3�����@2�\\ۍ�xq��F�����-�z�ej��Wc��Շ>�[`�����]+>=K�N�W7��og�}$��̾7����ӛ�p~3��a��ܝ��)Mr�� �s�0(���m<�3�����&�YT0&�\ ��UA{3�F*��(��F7�n��Y_]�{��x/;����:y�%4�V�8�A�=iL�:{k��hx#��7sr�g�����7+b<�\Y�4#���CQ����n�}I�����(��E�wڄ�(�l�gϘ#؆��}Ji1mWyI1�φC?xj��A�6V�n�Eә%n��
=>m�8��9��0�����������������x�cr���]���h[$(�b�"�*,ܢm$x=�Ф��<��bT%��>';��6���-�xv�}W�[U�`\5�ؗN�2��x�����+��-:V�1a[�򺟏	JG��X݆&�@Sx$FǱ�ף�r5b+q�DA�ʕ��|vI@0v�4"7����;?�#>�rl��lhCضu(ws�#�"v����knt2gaӏ�k8!�U=���$E��s|�ޫ+��qU)�2g���G֍¿eI�v�H�KG�v~7��m(���?yo'}�����Є�ye��e�cA��.KD�J6ΊТ[����|p��ő1��w,n'�˪t!j��ĚƇӺ��"������7�r�AO��AQ0�����i�"���U[�i�
�v�@ayZf�?q�4U���ߑoC�i�Y���]�l����o��V)��2%ȵ��iM���8� �s[Ҫ������+��c��-�6(�~+��A��ŃY��-��fXB C��h�2#�qB-F�b�lǿ�n#���F���S�]�~�}9�%mYc��~u]=2�E�2_&�JӗU���ی���~x�Ok����5�sV�ǢdD02���"� FJ��Y��jF@��tC�F������`&|W�F=n�W�tJR����J=kzR��m.��V�}+V.� �riNޛ�b�>��}F�˰w'ɠ�S��X�\}Z������0s!����������i��ɚAW"x���������i� �MQ�t�7tZ����A8l���p�S~�R;Ea߰V
䙅���s�N��T10^O!��Vc����y�t����1ɋ��2ڥ�1V��5gu��1W�	�_	�CX`=-On޽����.�|�9�Jk;P�j�{G��!ǣG]�$y��ӵ*p#r�wޤ��ƺ��5���EAZ�	��k7�ɬ!ۯ$�F\�؟b��}Fy��Kd�+���Èl���O�"	�:1��ݵڰ�H��Cnz⻒����8���$��B���ڊ#
��DX�,����+~\�H�:��J�OF���z_��qu��:4�J�b�ɀ�C�������5��p�2��?K��5��B�bzN��b�0�ا�o��)�0�4l$p��M�&��y��:��U:��b�ed�%ߓk��:��z����qYk���޽��܉!�N+�ȸ���,�0[))��(�����0��~1��r$��s�tu��t͍#{\�����|�ޟg��j"\��T�B�t���ҙ�V��h����2�E�f�W�Q������f�G���X*�������>I��݃�mw9�a:n�=��` ���~nl�/H��0�Y#�)tQ=��n��*�b��S��ZE��̵y'\	��m�:1G̏����*��6HI���֐�x����`�C.+�� ��u�h��{�ɡM�`����B�(��w����O�?�����4�~<���.���7h�!3?��_?2�U[���G�= �@���&l|$��v����f�t&�M�4���Z��d�����$�)^cg�%��)�g
N)�OTu�����C3��w�
i,�3�����7z���N��"�.)��퓖�8)��~C�rn��%��m��i��$X�'�dO�KѿDv�sA0%�2��S�2�\����K�M�_�Ri�����]��A3+g��̿�����I8���$K���糍��ُo=�}T�)�Bz�[)d�1�����K�Vt�F���!���}��#��ehf���mF�s�gԡ5��,N���;HX�������$�:ǆ�x:0��UO����xCް����6_V�؂>�7@��T4Í�wL�wXF��1��Y��&�����|o�R�J����MW ��Fᑛ)Г#`��&���*$�����r�휲�CKX���M�+��`���OB�AYc��%�/t�h�+^�������l]��Ɗ/?Y��!6�3y��KL�g��rTі���7	]�Y�"��3����Φm����gѪQ�b��,��Z��������o됺DԘ� H�1��6�5�P�~$T$���(�{�?ƅ���%KCsͳG�#�:�u@�չ����M[�^����%[�1&��R�#Չ��^�P������@�gi >��Ԑ�Y5��]֊��?�˴��7.��i�H@�o#�8R�(w	/y�.�#���X�n��X\�[�%W+	Ԍ��@g���d8L�fJ�q׸�Qzk��[��Bǣ��yS���%YcCM��q�#���_���:������3s�Mk0:����ԉu&�p�]E��<��(��Vm���6>ab�{�gM��հF���p<��@ÙJ�GĪ��b ���4<�ɀk�ñ?� �8g��A7+��K9��m<�iw�U:��z=�5�CQ8Fo�������|捙n@�D�DJ'�YPQf��9Q���r�������͚\�n~�A�}�zf/Ƀ?JpBF�����:��@jt4�Ԃ�x���"���CM�;S4k�[�/݃��WX�S��k�k�\�O�����?��2�t#E��X4դ�v������]�0H}t��o�D��� �x�-���`�]�h��q�7S�-��Ϯ����S�@R�!��H>�&r��5	r>�=O�W�b����OA���|�[Q@6���S=�>A�(�j�8�}��L��.��VΒ���̔��C�]���1p!���8y��K��W��#���2hI7~Vk�����Zv�?�D���%Y��Vh�p����ȝ�����Rr��S���/1󺺣��Ċ����/�]�����=5V�;��io���	e
���B�P��6ftsd�#�"��h��V+�6�}�V�6���4��9i6�eɷ�}�[�qv���G�NC��B�6���l�077s���C��hsw�{(�9�d۬�E�jN|f��$����]�C4�{��e�TV�ί�<t&�������银��L��l��>1���ŉ�����xlY���(k���O��<�P=ɚ���s��e����C.\rl?��Yc����X�0֓nF���x������|���!Ge�M��x�<:��D�Q�T��B�	�`�P�5q�CLa�Zm3�x4�)��Z]�r�(E g�xރ���њ	Q���d}`_Y���L�Za��p>?�Q}~\]�P/��"H�i8O*�
�b
Z3.��� l*I���_���ĸ�8�C9��Y]ëe�׌}�ټ?K�VL����\f���F�?�4�,|������5$h�Q)��셄:�%�#�����B`��3]��p��M���b����pJ��VJe�+%�_D���R��8���0����!��DL+��d0mz"7|/�D��h��<lzBq���͵�ev�{���XNꄼ[�mi���_%�/�4�Rj/N�c�}�i0����:	VM	e����~x�)�D�� ��cm��:��NxS�P��.X�tx�L��A��=�q�F�i��G����s("iTךOƴ.��ْ�|C�4��t7���
�"�Ƚy�꬛�t&��/͏�y:�o�f�C�x'���c;���f�){�����n1T��n�5]�󌝹g��"��h�`Q���BG�6E3���:u��I���<ИF��l̰<�ã9R��%�D�W���h�d��I�gd��wpV=Q�6��rׄ��q,K[�V>J\o�$�z\�A�R3>��q�t���or7�]����-�(;6��B O�ZrLʱ�HR�Z�w��=Չh�2f,����8p�IZ����z���0�Y�3�,l� [�2P�����?��gQ?2���W=C��n9�z	AƊ��U����a�X6 b���B����x�
]�W��1��Ǵ�m��ý�+��r�O�Y#>�rkO �C婹����%5�X.��O}����kU%V�����g1J���[���r����3�{�J#���O�`	���������Ƭ��
nh�|j�y��V��X8"Mr��!G=�!�\'!����R�xe����P<��x�Q�F�@IUX��ΔB=�������U�e�J���E�B������7.~e*7���������AT���_�,S�󉭼�/�������8ј~%?�O? ��0#�Qgd�W C��k�C�f�҈W�}��O �*�E����H���`,H嫁:C��3��
З��t�huѰ��'�|�]�pV��5tȁ���J)tM���phAٱ��$캆F��� �O�TO�޼�85{uoU	��!���vA��{!���O�pR�T��*бe�@�\5��d%�����MM�<�{�6���ESA�-��8�츂R��W�5�� �*(�vt��g�=��ͩ�ĳ'�pࠑ~�יP��sܣ�d�����L��!DY�2�,�nT��MU�.��p�vF� �;ن�p|R�a
{t6s������u�h�O"��Xw�R9�`[�HA�uN���h\�H��ʼ�e�B�d��Y��$��ֱ����OR�w����.��4$��ӖLn���|­o�t�8��o�9u�ɦH���S.X�F�����V�b�a����p��������F|�}�$g0�8�ϓE�
��^|,�.qļ�u����k��F���l=��U9����+�@`�:��Y4Ja}v�-�����p��+n�
�������.Z���j�A�N���i�JE�2�b�ru��W8]6��_|Y�RD�|��ɤ,���b@)�2�n���u��6�`j�}	�z�2��[*����>���z�Λ��s���F�Xׇ���"̔e��yEI�Ub�������Wo��&Si�������2Ĕ0�XG!�qy��A�Kp����(���iB.���[b��q�׹�8lck��o@ds����L��3��4��槤�}�^l�Z�����кq��w�wtUŸ��%�ΊX��mB��;��J���U��z�����U�2�e����-l�l-�7KD�o>(�{�������nR�I��)�4}Aήn�J/���ʖc�4D0��7�:T�/kN7���Sx�Ĩ��i�Sw�`W��q�|�}�gf<�VU�=�7[E^���S]}�.)E\����R5� �{��TQ���D�o�27n�ԨK�Q�JVa�$I�E�P������3�s�k�J!T���s >ㅈ�ڄ����E��Y�[��a<���R�Ric�;�Y+�#N�6�\{��C����)g<�>d�Sz�8H���ً���$)����(�]4h�ږ�*���f�!�EZ�f��<���l�voE�k���������1�����p$��L[�1Ս��d��q%��R�\gg��'eǽ�=t$�Z!+$�.��-���nU�P���3w�ɒ?`���\7��],6���ewٰ��b�pv����*���հ|�H�F2v���NW�R�9��|EA�\d��D~h%I4|��([�e���a�^�lH�jޤ�p�����Q�! ���ZS�X�ur_�Lm��\��b����I���j*���0����@��U�'��x
��	Z{ŷZ���K'��1RZ�\��e��gX�?ȋpA����IX�*V��t�*E�}Y9�ϷՋ,`�4�7�@�P����lg��^� I;�g-�K���^�����Wݸ�ƈxb^ꌲ�� n+�jH�ɍ{�p���\yMz��R2(Ɏ�8E$�l��\�_��2*ܫ�1�t��6�L�#L<n�ݴ�`�$�٨����;g�-�В�/����S{�"����Y!�BW&�Y��6v&��o�4_��QQdnƉk��<��Խ�%��wY]N�M8b�E{�ai�KQ�r�������"�lFܩ]�y�xJS�A:[�LZr�1}�\*tlЁ����0P呯�D����ɻ	�vk�rk�P>�R�Y�l��QG
�6G��}�p{�~�M��}�M�%�������I��w�}�lܤ����B���A�&W7*���{�*�������w�D6�dU�	�Lp%�<����Θm��H�9�����U߮��OK
�	
ੜ�I���\("��DUs�E��c��FÑ�E�3�ݑ+���):�3�u_S(��]kmö���V�x"�d9vRkr2S�f��Ϛ�͈L����N�vpM3��Ay�&"��˝�~�C��u&��op�&G�_2t1���˙g)'Q�l�b����$Ó0�P3�zf���9I� �pO:�y�PҨ��i˦�6�&+��c��2�"�ض5b�}����w`İj :��=���"ҊC�G�T|��EܷP@����K�y���-��"�I?���y�Ԩ������&/��KWg�R�E;YB�:��K��~_�X�)�\5b�P:�i(��.}�;C���:� qJDT{�x��r�>7?x��$+U]��g�Z'��ġ:��b�*&��l��y��m��.���`���'��̱�2]���#c�pu�އl�|r�
���e�������.���<U����9+(Y�� (2v���@& �eq��#i�A����a�R�
����$�Z�R���B�*��ג��B��hq��5U�_qa7���2��'�w�9���a$�HK'��"w�tlςwV��L�x�������/����p(���s���d�:R3�#��c0�W뢍���JP��'�d�]fp.:O?�c�վۧ7�kޭ��J�|����'Cߒ� �T�hx&��φ�݁g���nT^P��Bԁ�_�w�)5B@8�W[���	aN���bGK�nY�D���e�\��<��,��"Sh��
�n�	gy)�Q�5�_�`��?V�C,{���	�.5I/媃�ٮ��*ܑ�&���Cl�0������N�cL-�Fb���n��O�KF8I.�}
�Bfh0�� w����u�{�[7�����G��q����W#N̕{B�z���7�����‟�g�g���0nWa���Ok5c��n�>x��VA�Ό�UEJ ��������+�?b�VDVʴ�Y�ݐ�eww��+���Hr3d ���9/;��)ę�T�u+3;�t������Ko���T�fz^t{��N��s(�f퐿=҆���n|z�!瞯6�y"o�@I����������g�/)��bdj�@�Ϊ,t�)�E��)&�kf�S�B�Ѭ�t0u��ik����2ӆB-z_��
�L���O�GR��͌���p\X=�8�����>�Vw^�N���Y+o{�*ĒX��uX�rA�v�|��y`�TH���YeO���C�!�;�ԘvI��w��m/�A5x~��m�' ^f��n�;,Sr�5Х9 쥄��������k�c��%�RIs�sG!%�D���@��Z���$�;�$�jeT�cxD���Lx|ٔ=�ǲ&�]2O��G���7յU�^�Uyh�����\���:��sW��=nv>��F	!����Δ�%%�x��c�G�y�Jt��J��f��7�s\�^��Av�Y*�$�O.q���5'eK|(Ǖp�1��6Mxi�Å{/K}�(�Qjٺ�A��L~qFx��q�ǩ&/�W9�@>�n��`��Ŕ��Ā����R�;$��V��q/��m�2�B�>�@���P��K�>��/c�O�G���*�l�!Jk�5@�^lw���5��a7���E�� ���Hc�F7Az�L�=H+]8���$���ݖ�8�3�I�s�Ar��P��M7�q����^HJbO����v��;G�&���k͜ocf�[RӢ���l%VNt�w�:�F�X�� r��&���%�|3���m ���f�8T��h~Z�(W�������j��~���"��7��~�܊skp}����B��D����1Y��ŤY�[?j�7;}h�xt�w����j�(��y�� ?��f�$��;�X1�i8J
ʌ|Q�"u�:�'�G7�Q������,*�t��0��q���6tE�H�J@̠�p�a�cr�8��:�e��F�*�ͬ�2�u� X�
01����q�n�,تH=->�S�S`]�;��F��a�^�Y��WSr�f�^�3�T���$@p�����}��AǄ�n�798:T,Ѫӫ���ɹل)1��KjV�K���D��C|uD���C<���^���5t��(o=5�l�IM���Φ������}�.�D8[��q�T��J�|#�ޒ9V����Y�бO��Ns����v��a '��ۆIr��QmXM��0{[�<sWvh���ހJLaYj �����;���9�/3AZ;7_�����byf>_0��ÄN��V�3�3�ltmI	���)\�n��J�,JԴ�[clp�����/M��ށ�B�4��`���ëb��tR=w�#���,w�m��!>������|���UA휐p5K�&7��`xG�~X�����r����lJ�VG���J�΋6[�A�>n���ש��I&��$N������Q\�\(���ד��-�N��NH"y)I]�$,l�6FoWj�pKr`�X7�4Q��1�G�#��?]�t��Q[�1�����4M�ү|i�8�2���}y)�aD+j�ۧw<�&�n��Pj;̉u�DxZo
Y�g��awp�h)*J>����N�k���>ŧo蝦��><%�_d# :Q2��Z�@����ʓay<��$�]����f'О�ed�j�;����@���<!�ө2+Z7�5�G����2xr��]߰��q�?�I)�u2:7��*$�1_�yE����i�� $�7��z��٨H��x������ |6�X�`�.E�\`�.����j��Q�;�.��������v�җ�t�Ȁ�����@�&|�٤{�-�����}nV���"_�?����ʱL>1�H_�h�b=��V�T�y�x�[���n�{��+�W������=W����ȕ:«����I�h�7�)�)���W�R=��c���$"�$�����8�vkA���Ȼռͷ�����%6Z�n�,�Q�}���˪��=~͠���}c�m�:E���n���6��C��1p�H�@m���؋v*� ѯ<��;�p�T��LF��	@[s_��C�5�4L�O ���>�x�`�Pvo�����DOO�1w�҉�Wjίk��$@����4�.�1s�B�%��.����`�Urhm�D�ʄ��*Vr��+�P�:��Q�Č�� ���ӹ���()��F?�Q)�����`Ej���� @8�~H�����Rg �l;����\��\$%�`N(H|[�~�����a�wS�h?܂H�u�������`�\�9�φt�|;0����
�b���]�"<�)��L����s��M�O&����H��rC~��n���5�������S������;������>y�rȲ�����9-K M�����9���I���������6D�����+C�Kz��9�j">� �43Kc�R�)V������:q3K��+Q�@z��HRx0p�O'ˉ���;@܉�Y�
p�]l��� q��_[^�(��m�'��H�L�ą����6R_�7�g�;"m�$@��Kվ��o�!���[�ތ>.�ƭI]>-��}�Yn� e��Մ��æ��&Ja2y��9'��B:�й�σ,</��B�7WA��|�w�Y�Ճ�0��Tt,/��@�h�`�ƙ��8E��
�@�w.��M�m�o��I�
˔Ǭ�m�ޓ��<_�(L�v[��I����UK+	U��os��Lw�-q��d��X�z��|EA,ӺRy�BH �X��@Ϡ��6Jk�N��Zc7z;�*>Q�����=M?<�q$�!����S)��b�i�{H[W�:�+��j���B��J�'j���y>�D�A!������"��]P
��\�.Z���ļ�W�h3��/ҌQ���&�3Ā������`LA� $+c&@mAԨ�N��N����eR"v�U��H�Ώe5O��8�V]�R�%�U1FӢ�Y��Q�P"p�YkL[J�Zԏ�6�v�o�����q�/#tW'@{�l��)��\ĳ~��c]��6��B�B�
�!a�ܥ(���*{���P=��;����p���nh�C?�km*�W��I	vM`S�)Q^�4�3C7 ~h���1'D�-��#�Q�M�ܷ/a��������)4�����^.���l8��'*�K�1p=�T2�ux�(S��A&*�^ 2I�2T҈����
Ê��GZ�f��ߓ|.�|�`�MRNta �m�ڈƗ�)G?Tj����B\]Kw��a���J��w�0uH�_LO��&� �!�����*J�"��OX�C����Pw �U$�i���uu�S$G����!�[���P��eZ���XZ�������Dw��uf\p���=��IUɾ��<����Jak�$aU����H.}'��q�´��EJ�Q��"�[�5�`��_����M:�	��}�>��k�%��\�Gn��*�!B2'�b"ڇ}�C*ϰ
���5(Z{����/c��j�t�U;-1�9W}�r�j�u.L�Dt�8K�{�L�eY�鳣ӬDKUn�g��%՝�r�Ff��Z�$q�p>O�骗�6[SL}}�� ���Br����H��`�h�9�D���Wp���q��)d�Q�lnj���%�L�t�j�Qy�i�3�(�ZtB�XE�;�=�є�gpͣ��N�q���#�b�*��?�t��]t��Ԍ�S�=�E�������Q</t��Y!Ë"�C�����p� Y�Kܧ�������H�w���5�{_���3-5�J���t�\���4���F���NO�E#�VK�r��w�W
JO9*bT2�#{T_�K�����-v�Ң@x6e�S��qU��@��8>6	s�a����!S.�+��n��YZ����+�F\h���9&[&�|S��T�n�����1�NZ@��a��;���fu�Ci,u�>/�XE�����O���V:;<���6̷}��s����O��O�SE��.K�8�?��r��)f�C�Z!�ދ����:�?���j֗v{fN�]`��PbX��$�ښX��~��LP��n5��PUM3!W}��%$�n����Au��@�^�&�	�%T'��K�+�&�Ìن���/����H>|	���L(k�/��e�q!*V~$����J�¡��-
eW��RT�8C��v�7��m�a��V���XC�yKU0����t��Z@n���F	;�<Nkml�*���������aQ^Y�|���e��kųC�q���:XM����^�S5|�F��,�5;����{B~�<�gɯU�L��\�-����AV�{i�;.�Wy�N9�E�OH/���4={������ŵ?�. 높&
��-#f��&��?Q�.d�j�&��
/���!ł����%A^8p�[�]����5X�� �Lr3DR�<$t�ƽ�	3�����LW|�DV�9`�=D�s��ǽ'Ű�����2#�S��fxt���l�-Bu���~.��L�~ײ9�͗�|����`�oV���UV�$��^��Ev=d�M�Z�(����?��\�������c.&��6��m�W�)�ϕw̹�e�-Lv��G+n�
���V���6w�.�r���A���?�C\�/p�-%��B����E^Ȟ9�Pm���o���G��D�ነ_�Ub6�%���� B�J7	�ֿ����ې��v#ȇ!��j��5���'�w�^bf�.�+��ՕI��*��o2�$>+�����?_�x��e��x�Vg �g�}��]��jvx�E��7�d�/��YG�WZwيG�V�.1��o����3�����0	����l[��r�	�d^���Z)�-*o�c8r����I������I���=q9�C?KS�X�E�9L�gj��K'=��ؐ��j�+��c�����`m�@�+d����%�P�z�kPGmJ��!�T���؈�D�iM�:a/J��f���4|��｛Q��T^鐗	���%�M�U�7B��2w��tV*_µ�_�I�ɧ�/�ZD"�V\N����$�Z��C�mĕKЏ��=���xo��Cܯ�Ǡ�Xlq�H�@.����l�ޙ��yX��"��ڃ�r���(��e[�1%���)&�[��×k�k���xX<z���ѐtyE�*�m�o���oL�T�|�+s��&�̳?0��T_O�D�>�, �Vq�V�&�s��	68���,�z1�u@�i8���1G���X�L
�5��.��	V`��I| ���8��<�5����\PI�TֵYrjr�_̷K(�oTx�;��#�"���2V��B���Nq_*�Ed-7�k�(=�0�ٗB2���;�9Z�en���;���X_����J5�-��@AQP��Ő�
d[��tZ/H6R5��n�2HF��h�rA
���`�!�����v������NUY/�U>35�M�����'�;T[f��i�^n��<�0y=?��\�P{�1A�FbG��ϕ�׿�2��j�D%k���h	ۘ�R���,��h&U�^�~���j�1�m���?�q���cV 8a�h1�5����Ǡrm��M�i�M�ʎ��^�6 NB8���d|��P��S�T^�v}�9�R�����-#p":~3]��8�=Ę�	s��i�7�	 �N�xsX='"7I���4��0t���J�:��V�b������]���Cr�kČIv�& �~�����TU�۪%��� �ڬׂi��
[����_"�E"�m��1���o�J��(WZ��$��~��*gV(�^�|ݲ�?�,G��E�)��l���7dKh�˸��*�S�Z�	�^=K��j��m
��]��*d��=a��S�E�� G�$=NӤzs���#�����S��W�w�an~�NP�ੱ������l�d��.�L-��2�R��Z���<��0���o���,j��ĸ�!�Q�T�����vͻU)��)#�A�]J�6�7�1U��Ĝ����D<��&H*�[Y*�`W@.�.���k+tJ�ɓK�~��	�ݧ�������6��L��2e�Y��^����-6�mB|e���K�gh�B�l5�1�@��J���5g�X��&t�,b�d����gv
�D�ĭ�<jK�ıf?6���M�:q���W;����aO��a�?��L0u��<�9V#.�΅�a�*b}f�V#NHHT�4�>I�{)�A�ͺ�M�52bY�S�����1|����\ש��gYJ>c�q3�w	���;	}��o%1[�Ix�u��g�:(��/^�D��8(�6��r:6���%1�E��x'���y��u�l�s4ڿ9(��5�x87$��&̗�^�Ѵ�����C�.����*�w���;��_;��yv�j>���\DK� �c9W���Xy���kz�wuY�R�'��.Hh�Y�O�ڭ�Qx�y��t�×��$�_o��'���8�T�r�jsZ�\gh]�lɮ1��Q���8�
 '���ڦ�f%�����P\=�&����6���Y�mx��p����*�P7pJȽR��(�w`��ԏ��(�@���!͕�R.�v�Po�h��!������bEp�q+��0�ӡ-���L�,�e���I�X*�`����w6lP��\��3�)4`�� j���l���
�(TlQ{��������5�Kcݬ��g���j����wu�d�آ�D�������R[#�6~Ơ�%�h�Z$����n ��=�]��Nf�%�aH	��qy���F����}��fXz̓"�� �a�w��{�� ���	�ĺN�E݄�m^��%���"�N�{+>ʐ��/�yk���,���/��EJ�:,��e�V���5�Ϧ��
�����=Ę߅��S�[�l����^�>�/Q���Vn�c��`)�]���7� ��G�"�]�>hX�
!$7/	�m�⧝_�b�%@)���J=m/�q,�u �Q�����?)a@���$���J��6�b���f g�u��lǡ�6>�?�ҧ�q�
�f�q�r�V�7�F�o�XM8�����!	^����p�d���$�g�囂8"k�f���Υ�����%E78�36"��m�'^!���C��G��S������F&���aC5a3�l��@��p�G�՜N��-��r����:D�H�J��n�"���D�Qߋ��L'Q`����p}�t7ծF���x��˨m7��d1�\e�qd�!�]*�����>�����Ё�G��
5x�i���F1?\���9iB�uͻ�h?�AX�����QaZ(�R=5�)U������e�K�eu�?\������u���(D�P��GE̾y��{�YTh{�\<�0l��"���o2
B���hms�(��7�g�+Q�Q�4~_��
��	�n{�]D�E��.-P����l�k�Y8�f�F���n����a�]wQ�bc����~�����G߻�:q�/������xQ�F�?��0�渪S�ҳ[�����a��?��}�:�s{��o�����*��g�7@���8x!Q���_x�6����Dɪ�a��`
lF��ن�R�p��W�`�.�7�m��"�c|A���-S>$#��j�}��>���Ns�	��� s���.��-M�
�=�۽ӥ�-OBd�t#ӟR�Ȣ�㚉�o2��k"{�(UQ�h*,�l����SK�L�j���@�U�<[f�~ұ΁��p�`V��%�v^��TB��s�� ;��I�X��/w��be� ����nNs�z�7��W�0&����W��J��6!
F?�0�y*�;������> d% C j�ˊ;4{STE��MP�����,�Y��6a{�%}V�(F�!��3�SJ_����@ �� nI)=� 2彞�p_����~5�dyt!� �}.�<�y���:��������_�ڈ*�X�S�B�?�F�����H�� ��dr�����JD�Vo�Bu�ӌ���4m�B3�����qwm4N��j���@�Pf�ei��2]^��h? 97l䗠���@�.�Ie�"�����t<��6v��ҭu0KW�R�oJ?r��2�E۵�.���۩�g>@���|�DI��o��C.��St&�?���=�+$9C]��r�m3I%s��3��s�%)��@
J�(}���GrIt�B�A���S�?ݢ�L����y���k	 ��07O� �@5�%m�a����O�:��Ba� )��ݬ젘�&�ٌO�|�@����⨙	Ͽ��@�/K���.;s�3�H_���E�]-�.[oYi��O��$!�0M����2�������o;�t[�_'����NBgߎ�O����Φr�����^PA��Bt�a�5q4yϿ'��s�z(�'5��[�SZ�T�E���j:��Pt]��zd_�T�	u'!+��e�
�����߀/�1��
X��,�˰ب=��Bg�De�	V�R~�AV�ó�Dr,��#�I_}�Z���Ƚ��$�ێ߇Y�u
&��i��Y^73vi4���┞dx,6���\v.��n��\�x�ʭgy}u�&K�t3�A��+����'�K-�~�4�3[B;����i(�Ə\a��.�ey���7>R�i���O���r�r�T�D��A���h�Ò/��$���	��ß	��>]�����6p�B�톘������%-X�[o]˕������Qo��畫x��v�"�ce�a��#�,�j��s��0	с�؋��ESX[7W�=�yم,0��lM��W��齤Q��kǻ�tx�>�9�`r�I��T�w͇^.��~��l���$؆CJ���&= ��O§�����j�6�p}��i�gן�*�-b9	��שA����Gù,���8ߪk�����F�ƘܴŮ�5m��h%����/�z��b���ܷ��)=�o ��6YNW3��7�j�1's����7�����:�.���(Z�3�w�7�ia#2+&؁�ٴ`�����|�V}J���_��
��*{�d�����ӿa�p�I&4zjAR�s�
�y�Ϡ�q��l��L�;��)T>t������j�n[P�*B�,�Oa�^�'�k,��v�M9�m`;��e@`1Y����� fZ<"g��&���	��SqU#��2>�R�=�W���2![�I����������j�a˖��X6�6�[���-]�q�?��RAQ���?Z��q��s��`.����/�Z|�{Q��eqb�|~��	��`�X�8F����M���]\h:��G�29��1�Lpc0���4M�'�eA���"�9Xї�a�5�@�I�v�p�Wp<�Ef>�+0�!l�7��]�.��冘���P`���Rcң�Ʌ_{c�=�Oop$6'm�ەйiWW(�	v�K"K�s}U�Jg��t�Ie���\M���Z'_�B~H\�:t�6�kF�6SB�ߒzx����\�����Q����E�ָO?�V�Rn�����G�ά����e�~�g=�ڏc��\�>J6͔��x̮� cPWRI�X̑Uq��b�4�u��Q��t�//M���:+)`-��s�No�vg�o������\!� #��te��*k/)���@[����St
�2$jO'���������ĭh��
zS��N����G8��QԜX���<'�p�Ǖ/�쒴�g1U�����?S���0��ZGOM�p�z�wB1�A�,vK ��d���tUd s����xO���s��y�[Ar����a>�7��ڈ����Z��[�U�ҒS�[wO�\�\{�.���;�T��l,�$�Z)V�2息㈲����0 ��+>�LYs����m�L�w{y��s4��t`9��Cy�j�m��5����r
�'�����+Ys!��F0tSXJ���+h�����}�BT$��@��k�=U<�[5SJFy�)�����\E��*�8-�� k�p�v��o~����!�u��p�>p���~<�����]������I@���TŔo��
.�O��ܿ��]��%c%#ۢ���ʏ�}����fKq�A��UT��w-�IEvO��Š'�M���:+�Y�"�~�^��0W����nA(�_b�(�.3c\w��ʘ���X��u�y��K�S�by��)�d��{�ٲ7��ķ4�AN.����������$�24��r�_�rpY��a5g�sbC����x#��,WVK�Z�]�겿�{�уy��u�˃���:��$n[��n����Lu+��r��d���C�IV��{�:���Q߬��6$L��Ӽ���kO��<�j{����:OH��a�����&�Gp^��('�D^@9
"v��[7_�����PY=�|���&2���a�/��L����b.�P���u@BՒ���<�.���t�A�®P�����90�.i]'ⷕ'�P`uX<ϸ�^�H+X!<�8�KtD ��]{���"���<����W�JU�A{S�u��^TF8m^H��Oװ�+�0�N���s�K׈����S޲�vu�7�/��[1� o�x�~f �x���6>�-χ�Z���-D.�>�g�dN��ZID�?H����͖v�vU_Qr�i_J�`���VB=?.~ğm��*��]c�) Xw��q���^|��z��OH��3*u</����	��(�|p�ڷ�������P��xO<+Tx��@^O��M�rŖ����c��� �P�"�ԛ�+�?_��x�N9���ov[8��}�H�>�f~u±B���	�m�ɵ�`�X*�0PS�i7�%s��:/$��z�~�����<]"�t^䇱Q)È�A�Pk��!VL���<��ǋ��>���m[��s�����Z����r�<P�t	�h)E��kйC[g�}���`��z�����&5�t��8�s�©�&-�bODi�[q��}Imd�n��xD�4܇"�Xe&M�<���v�b&{G�6\!cXY�WNZ�4�+��ԭ��(�+����;.�ӻ8���3��z�u�q��n�a�CG��m��_��ۏ���_~0���>31�,����F�T�Q}�n%1B������O��!���+�-�8��O^�2?��.dy����Q���b�P�L�]���g�W'�N�����D�T����5!�٢
Է�$[ ���eOqᠸ��e�}�r=��O�½��;����`���n���\\=�1u��<�G��C�Hg,!����B��Ղ4DH��z���)Y��S4i	e�E��P[M�폚��W���C�:�<�0zo"�V�*:5Kks�7�#��ܣ�|O��8�LbJV-��4����֡���RF�S�Ш���W��1]�Ỳ�u97
QK�d"�g�,�)Qʞ1L� ����}�jK���J@=���~E��}JU�G�D��k8�"��g(�R��ܕ4�H�:��p���\ѯ�6�vb�� f�+c[�AxEM�l�U�ë�e��F��Q֌_��.5�'8MML~��;3K�� Y T��Q'1ap��]�^�jf��{��/�:W��b��Xsr�R������Kb?�~���C�ʀ��WN-�������^�!`5�ۓ�kC@�ƺ�%����&d���˩l;�����W>����SA���w|2ȧj��^l~7�-�����~Sx�r��,h�/m"!��8#d�-K�f��<B�ۏM+=�:�5�ޅr��/hG�aS���:g iN��<�R���(D�����)�(���Z-!�+̈́6�}�E�G�����#��	kA/���1u ��*��m!�\M�,��-�ǚв���?8�ὓf���+ ���YX�EV�Gg��9��0���Wc�&�;�t�.A��p��jS*F�������h���o�h��}i�H�S���>+�f�0��;;���������p[Bf1�
"3	��uo�r��fM\�K��+�|�@It;')˴B�e��1[G80�`��+���`�9OD<QS�_B1&cZ>���m�r���a$CS�	"�Q<�X�y+l�C0���X#z�ܪ�L�Xa-b����/;�v������k���2�!<o_�� ��,8��cY�Iʲ��[$����VJȘ��u��i�[?�:�ԗ��$�R�M�+t�F���Z��|���(���UԐ��g �e'�U�k`�HV���+BV�6(�E?�e	U�^E�jr�R}$�l�4��/�� c����7�Φ�qzK-m���O���69o�0����*#�S��D "1T�!����A�<��G�Hv��^�a8��9��z5��v��$��S@���y����S:2uQW-3>��*S�vG���긮ָًa��6U��
���k��t0nͬ�pMΕ�j��p�Z���>��+��Xe_���i�0�I'L=�1�~; m�^$|�wN��h���kp��^���m�ѯ!ERN'�Ǳ��'����A�s�OM�C�h�|<�@i�d�����ќw��˄Ւ����I��g�Q�u�lDX-�_������?��04������Wm���u,����Ky8��6��h�)�X��3��F��;"@�WP�Ӛ����X�Y�+j.·�B�����:��؂�5����ی�Z�t�ʚ?i�av�7U=�1w�v��*x��WG��(�y%yygȳ��#�Ĵ���J\j�<��(f�G��� ��J�g�"����T�[E~���=^T�-إ�qu(��D[Q���e�8�m����S��b�z3��s����ң@ R�*�醸	���� ��@�B�i"[QKd��`��mQ}�j�cEK�t>BSCkI9;��q�3g��.�f�~]��W�nW�f#v��%bj9�`gD4��_/DϤ'BJb�|.�^�Ȗ>������	�y�%SA��g[�̢E�ɿ��:tS	Y���R���,<L�X����NX;Z���O�����D��rrK�t_A�,=e�m	�����g����׀ee�\��"M��F�n��F�fbI�ʺQ�%͜��\/k��w�ںk��1ύd�&�[p"q��(]f6K�4��2s=�6>&�i���6<ω��Ri��E&��|�����_�>u�6FxA_�
��y�.z��3O���(x�7Ѐ���내\�wG"�����=?t0�L�-��x%�(�C��a:�Y+¸�GY��$qn)�K�1b�Ϳ�f�ν�˂�j��cJ)n�X_<�2��-]�t+�N��ҝI�����)�S��a�3����f'z�&���DE����rE7�6����]c�Qj
���jv`���1��t�m;����Y��f!�f$��3�_lq��L�a���S��6&�d ���Ad�D?�)��꼩��������EOx��Q�9I?f�K�xZ׎~��{Z��q���4u�5����<̑�>΃G�=E~/h��>����O��� �����D����3x�&�k�f3o�2u��:ݴ��E;ӫ�cj���Ps�( y�(Юb��x9q��؉KODo�#��4�_��	?~��L���>����W-��[����)�Ak��l��c�pL�� ��+m�6}{��)꣞��B�	B}�N�l
��ޓ�κZ�+5ݴ/#}�^_�;Cށ"A|'R�d����s���)U�Ɩo���|�TC�O���+���ꆆ	�7?�5=�
�,���@��[2�Qw��Z�4� �騸�6!0WL�w:�|K �A+�5�͌sm���;C�c(�+����]3�b��{g�X����0(UԵ�^6NҺb�9�p�ќ#+�_�x�Ǧ��7|R#�D%�e�ȥ?A��SYG�бfn��~�p̪���+����!��ɷi6���<yg<#�*N՟9�R(^��"�!�Vc����9�����N����`z
:�I�>���2��FY\�����;�&������=bzJ&����܄�Ѐ0�"���X�Y���%(O��d���[23�2�a���5�@8 p�Ћ)-���_`\�L�Q,2>��3#p���5�������: .����)�<�o�/Ñ�{�����;�m�Ƒ�$�l|��S�)�h�$I Tf5����lEbλ���#����U�٭W������S�r��=�H���Dn���=.O@@�\P��➖<�'ué?��s!S��c2�kD���\���ah�N� ����������;�]T&�$��[����l����FI�Pa`�\����ςI��f.��b�hR�I,�+���,�B�Y�z��܉�4���N�x/����
[�n����n,h�`=�h�L���!��%p���a�z7��1�w$O���c�_ �U�h��p؏�:�1�52�2J�Q$�������3��|6.�9�&�3K�;�Ѕ����kB��:��,�ד6���%�H��7Nyp��4!/��7W�.¾1IZ&�q���	%�Q*aѹ�F˄�Y���!w#(^�x�^���`a�ś��q�&����>�h�>�C��N�s˄����a�O_������p�R���'��_���C٥���
)ݶ��w���U�{p�2���D�����z+tx
��/�4�N�l�(98}O��w���c�
��Q�nH�z��,�
�0��8!�_�Q$�����>l��/V������UhP�w�(x��p�����j, �:[����F���������p.ĕ+��i��}�R�}nRus��0y켱����i���"ATGs�H�Wjݟ�q�W����A����J�[#R�6ƦX�]6�8z%�h�'̗^��"׈�	��l|x��q{�&#���Z[�7��D,[�<uw?��������T�VMc���[o�|x�̈&
\��TX�H�	TX"B�Yj���['uW���G�Տ�>���w��H������R)đ�o�����˨XXP੽��c���� ��io�I��� �a�)��zZy�5���%�\�`�|�'ؤ�]J��y���[i���'=��a�P�R�͞��u	ӫ����\�U���q�Df3+�lɦۑ|�o2�������0дߙ�{/a�
�]kWӪ�Yμ,>i�R��hG��Š`=��*;�����""� �����#a|F��{v\5�Kk+�j�Tr���S�O�$��0N
�	3�N��*dv�ㄝ2����G͝Ĩ�6�wVz�i�v�n0 Z�w	��nAJv~�g���kܣ�b����)Ke�ûL~�M�>�b��W���D�ؗ���/���[�g
�R%����-�c6KROVs݋�i��EP���eW�S��2C�,�a� RhG�[����n�G�p�M�����"ym?C�=�IEK�`�j"]�y&����]�.ˆz0�@d��#QyiL��LZe �����u�7k����p����L���S�xjE�/����gݞ��#YQ=�>l[�XA�&��%{ǎI�#��L�:CgP�
V$�P�P�v�v��R�"�jY�5��X�jJ�|$֕ ��+�c�nK��6p2���+k-2��k &�l�Nf0�&ԍ6��8R� 6uS���GTE�b��'_�?y�T��������a��5�*�wp*.��t�Ҩ)�di�0k�w�U͙b �u? {v�����T����*�e-_����`�nqf��d����YM@ĐO	�{��&�Q��x�d=���a#m�|<b�>[�C�ڻ"���ؗ�|x�V�p���!�R�t�]��Ġ,�u�嵖�G4u-ϕkjC�3y�Z��ǟ��'Kh�d����Ђ�p����F�1�@3��_ƨ\F*��M�k�P�`|Gc��U�*��a4 ���������6LP����W����ex�ʂ����}7�����a%6�d �Q��wZzt��S��at�i�Xg.���k���RWn8�o$�TRk�J�f�
`�sz�by�4�b�|��J$0i�+ecWJj�{.YM�����$:���P��-�gq
/�7�x�wë�{�zR޺X��|�uW`�����Y�mȞ���ra��>�/c�x�|>2T��e����j�w���6��}�{W�����b��?ry�����Y�w���j��"xKm`Q��ת/�F	�c����03�H����"�^߉Y�dɶ�ć(���\�L1�wG�>&Q����``4�p�ʷ\PJ5�0x�d�+�l$}�
k��W���d������	B��8WW]�t��+���4��T�� �vi	��C�^xj%�Ny��'�]d�� �7����c��6����G.3���T?�1 �d>5R��J�F���6�=�E�������ۋ�N��XQ��>�������q{xA"�w��l8�b�^�p��\������"��ŧ�T�Q���u�ET9��=�Â�,9W���Qb �c�)���b�}m3�����m���SA�@ �n�з�n�l�C���/x���.1c�k��Z�p'�
C�2��2攛��Yf$��mI�B	_��_�uB�S��a0}x�g�˥�wCsTa�,�s;�%Ga��������j\��(� ���/��˄�q2a��~�±�V����w7�<�{�Q�![��Z�Ց
���ݚ��څ/�L�!n�WW�ӱ}���#�bΔ��|���8��0�YC���eA�)m�L�g:<sm2lB(�l�\��R8V��Z�%h�[��C���*��������z5�.��mp��;���,�_��Ȯ~�N���w6�|�+;7{�R�����-�>P��̶���U{q��,�0Tl-��t'���~l�s���tQe�}�T���iB�;\տ\��������_���2vD���z:a��V��c���v9�<2t��k
4ԩ{Q��-;�g��~`� �^�vYxߊ��,����U���C��@K��&�"9�إ���5n6�)�*i���V$�� en_���I�����0*2p��~�"q�����>�3O	�&�(�+�z�u����8x����x�X���d���3%�M�	=l��]3�>�s2�V�@*������26I^���tT����7��	�z��o�g��:������YܑQ/���~��n %1v�u���:-	�%7�X°��
e��-�����q)�C��3� �,� j�&"�;7^K"�EhF�r+�?ˤ�)���S���r�:�d_2�#�BFLv3��x7ө{;:mi�{8�j9�a��x��ٰ��t&��"��,��9���t/e��:y�/E7���y��ѧ��Q�p��|-&{��G�g�B���C����Kes[�S�n{W����n�S�=b,��#�|�c�Ef��:�hk��p�s��O��I��Kd޷�f�@C��h�.M�ܵ�C�=g+�"�=�^H���G���h͐�њ{�A!#ԍA����w>91�����mw�鏌'����'v	�@\�A)�,$V$���[���JS����T��4%�~Y���As�$ϟ�@T{~� JQ0�#C(����_6�OF��]�t��)N�W��VL��o����^c�W��S!m�t��H���+��繶P=p��¸���p��/�ҁ̅�����캽���B�K��ݠ���)��� ��=!��q,>�}�<D��L���{Sw�xkc��Tx ��� sa���ٖf'�X}�?�ߧ��^��#�<8����T�8�@�h:���B`D��-s�r:�g��ى>�UT�C�u�g6��	��N��7�$=�[�&)%��2�3B�
^a�h��f�շ�&��qu�_tƼa�����º����ҋ���0\�I�]����T#]x�����;-����ә���:�b-���^����3���$≌�ٔ�%���<'�����}m,�띳6��2��	��6Ηfce����s����WI��!��+�Q�u�V_ۅ0�o]��e�v��'r�ׯ�z����2w�N���F���JѡK�J�)O��G��F6H�K�q_�*��LH�ES�_M����g�1m�r�[1��T�U���j�Pcۢ�������m�3[��ؔ����ͣ�bKe�x�@&��8�=l����|:6GV�\O���^�.UqAJS,	c:��!��T"��-Κ���9���QB�ZD{�hby.�z�Q9L��o��#OB���ef��d�qgIt��M�CQ�aՇ�'�~�5�
���;���s�E��r(�d�9�%ͪ���@�\��b7���2�x���.��#D\#�B�[ej�P8�fY\�EM��:��{%9}GcY�K`�g��n5�l`��R�Y0��2��9��"드测%���7�E�����t���~>�ċ=����3{�50����m#
�+�����Ivv�E����ϡ�w�&'�����Xmlu�8��2��h���?c~T�����K8�@We֯rG�w|@
a�"�8���v�cD����Ni�۱bj⟷6�2Ծ��d�>X&���?17�̮d��O��rf�l��G(�6H��:"�B���\�u5��6����{��g�+4| ������y��R|bR�*1�Tp�|�5�juzXɘ���DFrY�>Q��l���O��s]� L��Q�Es�r�!�ڇ�o(��~���U~�y�v���(�kG�0�o-��|��h�*.C��^%��`㩥ru�\��.$c���)��pa}��rj7������*j/m[��*����t���HC�A/��yQV[+i��\����[:g뒛6ٚVv��G�������;��U�%���ڏ�Q�l��4��yw۫���>2�͛�n֭����N�2^�,�|.��Y��:y�>(8}�D}*I16�=�B��i�O���S����Avm�C�cGh%|��Y"q9���V�4׺9k�����UMx.>��y:sT�޳�8��dS3��z�r�!
�-Q�қ���Ϊ!�k����4� m	�X�2
����H��)}gIe繄��ʩK�^�wC?=CD�k��d!Fv��C���(���_�P����ퟧE^�[�o/��d�v�$\��O*y�r�nG�T^7�M}��:���9/�2A�,⮷=֧�[1�X�/V����yo-��৊���G����F��Ѡ�=-�ᢏ&�/ha��̅����;�ͩ$��Ki��N�xxR�6�O6g)C��"~G�b
9U�Ƽ!:�9�OZ0m��F�z�"�åe�főH�)����������i�^"����b���᜺�v��Ly�A����w�����Hx���Ч�#����E$�ܩbx�h�(�s$:���l�3�1V	C��y�e"A�1�;9�P��G�����3'�	��
믘��a��|�jM�έh�9ب� �7���7z�O!#{Go��=i�ad��U�i��|�o>b.w�sJ�3c�:�xpvT@�)���k��rABO"�OyN�:�M�Z 4�������9I��g�"�� pe:z�$'�P����se�l�,:����P���0oK(�bL[�w��4@b�P��:��iOQ^�=h�=d3r~���wfII�q\O�w�� Y!=�OȽ���=����]=�TF�4<?*y:�.������x*I+އ�D Ff*��I�4���Y��|gG2��c�P�KR��亚kc2db�����էӥ>G�����]m_<�T�R�lR_^�4�K���zC��d�^�2YI�����p~�XS�u�*��]Ɯ�=��\D�� �C7�{�GV.��e5�?>�<f���@«�E��!�����dMFF���u4�w�ۇ���\�6T\$ƴ0�1Z:�7�MtO3��4"3W_�n����`�3�]eN�B�l�،�JG�������6`�,,o95uZ�:*��}n ��R{��Q�w0�g�Lٵ�<��4CW��SyRr i����%\��B3ԋRQ({��B� 6��N#���P��rLw��o��G�	�Rsz�LB%��9���$W��2t�DZ>�ǁ����yڑ�7��8*=��o>|�9��n�b�_��I��.�pi�u�ڂ��D��bԹ�G�Ҕ��$z�d�u���:R�{���������XWA��g�� ����{Օ5��E:Ι)[��w��?9A�L���c�W��2����[�_��eR�|�\���ub�w��HG6�|ĥ&n���@��w�oa%���".�*	��+euf�.76���Yq?ÕvΆ�j��)$���r$�&1�L��}�5d�\�8��f�.蟅���ט%j��kݱE1�0���3	?G笪��e�E�U��|î��*�U㊤�WOB�A�F�I��i	�2����~�a����$#Z$cS��.ºHc=�׻!";؂���=�?���?�--9�juDV�N�����3�g��$�/w\&�#���R8�6}����tI�)��
L��}��܈�Аs�P���2�((��oٞ��^�#(	m��ƀ�߯�9��Ǌ@�=.y���o^�-��\���}Y$�9�c�}|�WYe������+8�;��(-����#
��:�S���3^/ʰ>�¯����p�W����Dr?��'��s����SBLU��A�fP�ؚ!~���7?�cE�|R�Gy=A���y k0y-���W��x����W��ٍQP�*��RlD�q�[�94K�"T��q�����5���W:�n��hߎ1����_���~>�H��ˎ�R?
aV`p ��_�ѯ���G�nx�P\����Տ7�w�D�w���Jf�<�P]"������u��O�Ÿ=��fI{%�sb8���@���6BV�e�H�t�#ߩ�(�����Q��� ���ܧFXX���9mZ�&u��[!�t.ݪ�uccW��#��Գ���%�4c摞Q�R�L�qL\�T,/��JCw-�O�!C�xK�M �1@ tMq[5�9P_����O��3a>�&J;(BJ)���s�-�l�H��v՞�+`������t7��q�j�����c���1��F�XK@���3�A�[P�/G"���E �1�,���ۮ$TC_L��Q
S�������\Xŕ;����MS'Hl��{�l�]>�MOP��N�����`�0�%�Y��b{����<�q��S=|2���˦������yh>O�H�X��p�� B�Dj@1N�;�S�����*W >�4&,�i� ��r,��m,<_#��N	�k�<H�K� ��2r�p�볊�Ig�=���"������ ���汈�V�� ��D��Mh����u��u������MLCnk�M�.�4��6�)�'E��;�J|���K�BF�E��e�`S(�� 9[��z�����2h� V��R�I�@D���v>q�CZڎVY�SWV���詋�^}=�m�_�M���#�J|C�V���a�(�(�Z5�s�
׉�� ���U�^G��K��;�!�d������<AGe���\�<�$s�g���vV��6�d�=]�dT:�
��mrV���B�Qj0A��(N����T����G��k7�|��
o����(hR��2o�m�V�X~�.@�J��l֘�^6Df�Yr���v�cb|���c^f�.*�.��d�8U_fcnk���'U��F��{�gHѥ����S���]��	gU����o+�?1K˫)aأB�� }%P���$Ee�H�����{#�A�ٓ���Տ�f����2xf�-}�a�ٖ1�G���ڰ~U�	��A��f��uT�_u�q	��ø���ܓ>��bci��`m,@/iQ�z��Zplm"p���E��)�*֏�^f�XO=V����A�q����nӳO��ӂ�pd�"�b�_�jt癮�T�#/hd�ʶޭ4mQqF��]� H��=���������nFjX~\�:Y8K-i����v�kM��Ɍ���)z���*8{Yl,J9Ho0���D���/���t,xf�L��\$s��r��3�H>�m�)��?1��qO��FO	D�5݀A��^�e�P������3č;���(&�P�x+�\"�V[�\�7&�n��=��K�����0����N�\X��$r�S}f�S�����P0��4^5�>�,�b��v�9ncy4T���w�j�Sщ{�m��B�3e��<m
JjX� �������F�yq�������o�����u�5�d��uv�?-�N<��,WB�H��4�'��>ٟ9$~�ďqsSj�}�'Mp'7�@=Θc����U	Mw�(�m�$�)"����!�-�F�EG��SR���>>���&1*�����z���y�wsۮ��8��8����l�r͋�t�%��d}e�[0v�!gL?� w�/��.�>w��������⸌��ZlR5g�l��ˠh����z�M�/͈���{��њp_��U8_x�� ,Wϓ���r�EFJ@�������q���o�Z-[�	���g�`�돓����U?�P�.�V+��(�"o�Q������]�~�)�=W�:0+������-�4��Afhn����F��Esle�M5���H_���5�6�oڕr�@�p�[�sE���:`�m����
)!
eV����D�}��=~'n�;����xȢ�����x)�"t�dyL�_"��t��`Dp��n���f�}��!�i+!g���989�������ۨЂ��}Λh�7KI��wO���K�-�\;��ւ�U2�r~�3�)���׹�d���	1�R~w��̨tC�h�m[l}R?�L�����L� ٬�\G��ր�@e<���-���%�	ɑ�����e�����of-r-�mFT`<"�i���=��g�T�k���Fz/����h��¼�v��ԅ��RC�&�fq�ZB�|�&2����l�>�C�lc����/╤���k�]�4���L�.�{Ij��6�Vv��ݸv��uL�y{G�0�W� �.�4����5��1��Sn�f4?��
�#6���7�A�!�yI.��o�J+g���z��B�%����u��|�p��\c���چ�!Ԭ�e��	Q D!&#5�$�����d/<�ƙ< �psz��!aE灶��k8;�I�݁���M�,,��8n
���F�k���;o*��q��5"�	=p��!1�!�+�1|�S�x�놽!�84I���ĵ@��`-��.��X�l�#�����N��}؏5���t�FW��,�+5��jP$�{.I�&_g{��eh@�Ym1�پ�Q-)��n/%��*b2F:ĊG�ކ�˳��EO��T������`�MjQ�6 !�
���;����Ci��̡7ի�r�ģ \W"9fA}�t!�2r�t��lK�:xWc����/̡��ʲĖt�N$���� TR0݃Cɞ>Mމ�<k��׈�Ń�L��e1cD6�q2��O��)WN@o�Fsj����՜�<8��ܸ����,��d��5��d׳ׯ��L)R�19& ���+�:\`����D����\QaB6��<��g�@���`U��7WN7�ϟ�	M��AI�w\TN��f�v�PC�/:"�
(� �䄓�U���,�5e�"1v�v�Z�[fM�����3��j�~��o��c��O^�m5H�f1RӒ���4�u��@��݀2�:��k`��� ��G��,ƽL�6�۵��>�sFa��j��f��$����c�9?��9a�D����P�n�!�J�q�3l�����R�h?�T���S�s�Il�mGr��ή*l0�#�|6	�a/��}���R�<�� �u���b�+��i,���c�L��A~��ٺ�߶������J~�p��
9���Fx�t�1a�{r�MK���558����H9~�u����N&ߴ6K�8trAtci�lM_.~�Dd�p�o
�!�#FD{�6-��!��Q�g����(�s����XL�}ϯ�RVKY��2�����g�ր��w����x4�غ4I��
Ox��&Gʗ�A��������"�����e߽�}w�4
ɸ���Y4 \x�\L,���x�{�w���S�D�D�_�4n6�'�`�я�3=28��֧�Kb���Ұt�fZv�)\������Z{:c S���,[$H������V���l� m�.\]\ �%�0�=+���&�70����u:�y�ë-��Q����A]ķ����&i#fqZ7u�0:�h`֢��k�BE	��k����I�jgK��C\��a���������5�e���Wq�ą��M��X�?��pyZxᖒޢtK�l���:.r�W�Ն��L��m���Y�(���C,�R�ٿ^|�j�#��W���ט���U�m�2���U���2� >��x�j��U�=ޓu:���6��Ro���ȑ�3^�������]̺������#/cja��iT<�� �}B��G����w�Mj�����E��X��u��0Z��S;�A�7ns��%�b��5�^V;�U���t�׫^�r X9&0����=+��_b�3	�H#����gl�%	�@t��Ψ��e�3G�B`~x�!$6s�S�7Ξj~Bܙ��д�-�`�/o�=�CX`���L	�6����F�!��ƍ��e�mГ�>B��$�י\�[b�jk�L�ՈM��-�e)��k���>��򼑐�����Ɔ�����U#� -�/�o��v��am�Ť-_��v$��3*y��u�y��q@�.��&���q�+�i�+�����BJM�d�wSw��;?�[��[�^)����7v���@�c��|�؇ԣ�6Sj�������y�0�ب9	cq��r&^.kk����?VbВ���,���p�w®}��\ʓ��O��K�ā���'���~�e}+G�2�焺��,f���~��j]�N�t����/��������u�����EHz�n�凸�?���݇1�S����'�f�8��s8Ɂ�{���hb�REb�ۙ���m�����ރXp��e� z���NM8S.<�9Pd����j�SC�j��yY�}rx�������mO`�z,Ę�����P�.)2���S���{t�D��-����:e�D�.WkA�Q�ھ�pCn;G�-v�	�>��j4�uoĤ��M��d�1��L��1��b���z�l��R=%��L�~�0�$u�P��u@�����~�CuLWBNHg��J�Ct���9bb-�=s|biVqC�]�e��*x�Șr濍����.�=�0�%Q8W����8Aή}����PXa��cT�r&��Vw�.EB��KK�GTJ:�7��+17e�@^s�(�����>a�a�?`U3|0a
�G׆�QR�ڎ>��ɬ�{�ۮ�C�/�3�l����f_e�w�Sij�7;8Dd qTDW��@���\Xʎd:ɬs�z>6;Wo]o T]w�{�X�Ӽ��"X�l�|��бk��-30��4wwd�'�r�Dc�����d�BK*�%N�Gn��g�}��yYl�($��צK"����6�٠���:ĉWg�����Q�Q�HV3$�Pϣ����̎0�T3lY+OݸZ�vd�U��u��.2	P�?*<>�ʑ�Ʊ���;x�M��ᕚ�_��BJ3�k8��'LG�.��>{xz���?L���6�p����Y������#rGR�� ʖ(\�[W���ry�(�:3��)_.�!F㞡�p&m��S���%�#%�М�ٳ�m�|�$�Ш��k�;�_�ds�~���n$8�b�W ú~I���g��l=�Xx{�6���/�7��E�~���
;]@�/Y�>�Ė\D�hry�y|���o�>+�Z���/ɷ'Ж�����8
o����Ҝ�(�8���g�x9���z^ʹP�E��}����2�c�|�nB������ >��ڰ�K��iO�p��	_��y��/���z�d�Oyp�a<�c��9޲X�h'�n�rT�<C"�*a���_܇H��z�U�܂vb� J�B��$!	m����ny�1�8+E�'��!y����C��XY�Kn��a���.f���LX�ӛ	���X�=O������U1&X�;��ܱ,K��Lղ;��p_�F��d�5�ZH�������/���d��L�kh�	:�c>���ղ��VK�\Rԃ�m�IB�=�E�U�b��oy�eb�����SHO�y&�a[t��!|��� رw�Tfb�4���aC����	 �������ll"=fD<�C|��V��i%�� ǻ�_~����n�v'I�D���v�� 粀�|��j�\鱬�%�	E �`�}��!�r(P�/�#���5��,3w�,5]�Q���,� �C�\���HJE��ߖ�^�Z᝼�A��h��,�4bR��I��Ǵ.�-�~�r\9VO�?�-%_��y��E��Z7��G�;������;�v&�2g�ۼ6WxBSw����͔��6���$OE����Z�����B�L�W��)�j���#Ӗ�F��<ms���G�?�����%Y�2��(� �{^3Q�t�d̀��PI�؎�
`�Y�����Ifa�?��Nx��6�,���t�@�w�+���И�̩Tȯ�m��C�Ĺ0=5�rY0ipk�&��K����Ӗ����g�(�RZ�̫����+��v�O���9�vZ��͝�Ɣ��ߧ��i����kE�]}�"�Kmft.	FeA4/{{�H���Oަ�>��V�`���]0�w�"���q>@��H�vu�
�*ĿΎ�Bߏ�_�������ֵ��sR�����]~`<�I��V)G�7D�*:X1�L��57o���0�ɰL���ɻ��ၐ1V�i7�d�d�?l/'GUo��lF#1-x������8�aI���l���z|_��tQ���W�`��J�&z��+��( �I�ɮ!񉖨)�B���|�cK�"��YG�y��m��e�7�{H�'�8��v/U����[�M���њ��h	�X�N^ү~�?�i>��d�����7�nX*Ez��Gb�/C�����I�C0T�P��_���	�Q����k�7���H��,@�B�}@a��֮[Dp��3j�%>�>:��s�G1�H��͉���F�-6Qt�;�bG��EZ��ܭ�;C�~>7l>��`�L����(���h���u��N$dJT��`�����t<�ys�Rbe�}/[���������?�F����h���쌄:1����?���	$�HZ6?:�mx̦edg��A�L�!i��w/�����֒��b������߱�=���1�t��>j�`)Y�R���{/����5�V�K�Ե����Z1�{�YROA�gׁ���S]����<�md��"~���= ������$%�ϼ���$z���JT[4��[jn�p45t����(���*�B:�Me�{�5�y��=^}~Vj��Y�<MNjv��v�ȝ>��� ��^��m���~�Upo��Z���r�1-��k;ɺ��e	e���r�Fa�;�V�!hBJS���d2-��컗�]�7��v�1��ȩ��˸�\IL�e���vk�����z
�!�e��?��̛9���P�W�����**k�n^"�O�p�~�z�Ln�VY�8m���������US6�^���:���>�1�Ĺ��|Kq�l�t3D�z��ѻ��)S�V%h�KH��h�H�Y3�tU�W��M�Y�FY$��9�����x˰������>#,��Fu�ۦ4p&ҕX�����o$�{�xS����^��Ho�uGz��<|+B��U��ۧe���6E+��9]/F�P�O�+�F�^Nɐ2l�����؞����ڌ'�!����}c �SLc�W��}p��M�
�_����(a�*�V�K��̰�A��о�L���2t��d޺E�1�*df��}<�点�B��%�"�~:�Y���)�Q����S\'_���$/rg+�YrC��c���?B���d�&G�2�pj(Ш�ꍥ܄x/6��B`U�0�����>\!�73cy��9�+��m����m�v�Ҥc��&2�ܗ�X�힯+����떗s/K,v�(���h�٨bމ�������
�4ڽ��5g�k�m8Q�`R��B ;��M��Q�-�H��~���Xk��f�|�o����*;�w�p/�B��0x���b�I��F�sQ�f���B�/vy�֒*1�������J�s��v&/+�޼h;�H�Z����.�!p����Ye+�Yo�A��x����)4;@��Z�2C��S���\��n|C�HT��%WcT��r�1�.g��O@ܹ*(�pt7�X�uo�cz�u�-�7���#��?�^�E��=ԫ1���]{u�`@�&�it�yH+���G���@\_���(	��]a�Y�lxF��:P�uG�A5z��ލaK�.�NCf5�U��}�6޾>ٽ�t�-��u0s��'��ZN8-���)^@��I��H\�����]n���li�kФ1@	6��Z����"����rKu�5L�=b����������s'����S�"K�J��>�D�SꘅE�Ɨ��K�S�Fi�T��c��:�"�7�ا!�#��$<������|@8٥&�N辤�4_��w�CR&�l�Z�J�B�<��w���T]yϾ���ylܛ���o��o�������[�jq-�7�"���~ADp�G.�}Ea.E+�y�M9e���ޱ�s9�֡@�OAb��aZ�0e��k�]���_$�Q�-�O���$��[�>�G";��Ҟ�D�����"�R.��nʶ+@���L/k��P��sX�,�F���%�d��;x͂����_Lǣ	���u��zچ����w�a��῭_���������oУ�1O�&��S�W��,�H��g��~������5i�n�c3�d8^��mG����J7�}�8	�,RO'��!��P���M�:�F�t݈�5��^mîj(�6BCo�?g�[|�#�<��a���N�����x��9��Ou��Ii�f֝~�ۄ���q$���u�V�T��ǩG��\�ǈ�(�3�tq'�"ѻ��e�I�~�捳�!K�N������O�.lO�?��mE�Ir|\����G���<#OuL�n��r�:>	��WZdPǝ ��²�*���2���J��Y�z���nP߰��O�]G#ǰ+f~�A!�f�s4�M��/i���   N�J�I�F��[V�J���8l��~����(,8&z�o���`�5'��>�\�|��E�6�e�*;(�L!b6�:����U#Vk�z�e�N�/]	�w�<�F�jOe�xa�0F.����ʢ�½��UI-*ry����c�dP)c7v�B��i�'��El���z�A\7>&q�Yڔ��Vp9)���r�M���Y)�"]�!~/���e9� �h=C�����f�  d0�I�o{���I��v�ۅ���|� ��V��yAE��T�A(�2�E1�T�@��!3";ua!D�����"]�Y��a� �f����\i0Ez"ozv}�3�ɲ����_���Za�+хy��G���X��I��% 0})���?����	צN��l�[���Z��b&�h��;�Ű����J[WϢnf��/-��L�U���N �~�~Pވ�XY��ˡ1�vw^���B��Z1��Tke���b����}l������gwМ����bj���C�M�Nú~�1��6v�/]l;h�\�	���{��=ܙ��7d���
e��|�5P6n>r�R�T%��EXae5�ސ>@1{9��H���Y�8�O�)Ib8!ts�+����L%�ڳvB�j�_ ==��6��ȑӰ��Q,b/ڼ3�t���<�w�[�����##���K0�|�N��[\X�Z�]�y��͹�|�)���\��nD<���ٲ���LK�'ީ�܄eV��ʯW(�lZ�G��n��x��\��1��YF�����|�1�A�c�J�H ��d��<��Ț"ф�Z��(x�RŦ[0�%$�ܡY��D����[��� �-B�G���oMuPB��0~%�HW�σjk�q-�-�ރ{�C�����9]�1=��B�J|�p�gp�)�+�@�V /���ǲvJ6�1���t:�Q"��|�����UĦf�����5,����"FRL��zX�A�KP��Q7m�b��[��U�TV����f�����Y�&o���/�p��C��
��]�d��Q������ɫ�:�ؠX���Z�k䜰�X_yJ��r&�n_?�*�8�%F�l�2��)ԵZ))��dPnɩ���ޖ�@�_�2y�[��G�Ol[rL���A6��n��uX�rՐ3�'���6
���R��\��z-R�Σ��->|HhR#�a�~��=pS\0ڬ��M�dU�u��zS0{��,�Z�}F�)��̟=x�)�59-$���4f$.2&��_ln���Xu���N8r串�&q��&��;�>O{�v[&\�U酱���>���k��@��(�2HV�-�"�����DH�#Q!&[�C��[\�<hҶp�܏o��tȴ��>�5����j<�S�>�<�"i�]޻CϬ�q��mE!ق#��Y��ֽT�J��ՙ��)N��]v9 �_�&���
"e�b�������h���j�g���4q@�=�:2��pXf�����m/DQG���@�1��7?1iϥ�.�N�_
$;s�_6,t��L�Kc���=~ ?Y���~��Y��STi����v+�	z	8~[Pb����
��t��gn~BOp2�~�u CU�Wr�Z������91���{�<n܂e�軱0&��`�f�?P�����$+�/��<�d1Y}g���g,�Pa+Q��V1S&;UMS<�
����++R�j#/�`�G�lxǠ5�A��ﺘ��3A��l+1�)]��kBmO㽛6`�����>�J����X	]L�<�JﰪZ�|��}i5�����Γ�����FyT��:��l�#�wp8�l��}
��N�[��dB���l�i�i�~D1@g�*x�2[1�M�W��~:��A���j2�r��W�T��,s�+;��O`[�v�~S�x�+�R��fod�A�]jx`��Fk�P-�I�Ja�y�\��G'Y,%�D�Kx]��/��/��Lfj��18�Gc�� k�RnpYW�8��p� P�'	�ׅ��l{��d��.�FX���<�j�PT��j%]��$�M�|��p�_j����"k�=]%��yõ0�������"��!@�������#�%��ӓ� k������~6MQ%��Dd��\��M��Le�O��H��#��J�T4��!�y��NMس9�`�m.��@jcH���BH��[�2�N�D{6SM-Nu��8�k�f"�^���Q��m��:�v���~'���`������c�,$	3�<���_�]\5|��� 89�S=NS/�)D
�Dՙ����� i,*P�;3�p`�Uy"D��~���}F �v�M��¥[P	Gu�l��ڲ�q-]5
Z'��C2~o�l�e�}�Cs�⣺U�9d�iJ�������j�4��/!N-ʢ���������!%sz�`1�!��Ŏ��ˢ��Ԥ�=�S*(
��uo�~�#@�1^dGl�Q@���m)�{϶bJ3���T�'6>LmH�-ڴ���DS�4���}��R�^���.�85�sa꬗6wd�ˌ�?�8Q*�@�z�b�kmb�I�sjc�x5'X���m��k?���VE���B�K0<F�|tʹc�u�3���g��.�<��UY9���f׼�c�(��1�8a�BTZ���¿ǋ��O���C�N��Yא#-��)����[��{xX32�;�I��#X�λ�F]I�T
%�����'=E�e����&T!n�Lw�XEJ��f��K/}��ڵ:w����B��Vx%�_+00��!O76$-���T	��Dv%
q�u�sʱ%e�я[�T����_�g���ű0�8.7rB��rBS�j���ǉ�CN.g����~��xh8zg��<!��~n���.��>f>�l#
�N܃��?˘��0^#��'��ap��#a�떖�H.FG����d���-d�'eB`�X��G��|�j,��{�!nCnŸ<fde3L��v�L�F��׃�'�٩�B�9�Q9�@\��f��cW�6W�b�,j������D�Nc��vCa�%|���2��'A�QX�;�c�-m�>fm�Þi6W�.��Օ���eQz��,��4w�9�mu�k�����Y'��]|j����EL���kej.7�IY���#;K�����~UP�g�)c5�ߎ^5��ݖ����$t��%6X�� �O�[W��o��L�d(�`�}��l�j�z5Y�bB-=j�ݕ��	�մ�����a1&:j�>��j�������^ IFs��!��r%f��,V�֫`��B��;/�K��v�Y�n>��� � �jB����J��.&���1Pa������1;q�vT=��<My-�b�D��������-���: �LB�����c��=�5(ؚ�d+0� 6���5B�３|r�f
��+�!��KW��RU�&(�y��~�w ��Q��8
�o��Ƒ�����	�jRdO{��>>-��}�Tgir�#/5ˢP�#����1�����u���eէ�y��y.��X��;Xs�a��������by�O�\��&wn�b��fK^ U���S�ਉc�䢣FyvT��E�H��8Fgޥo��Լ�c]	������WS�C��2��#l�����iFS�@��O!�����
S���B1
�趩#*_.e�}u�m���z͹�g�Z>���φ���C�ጜ��H
�r��f	kd�֚s�YDpPU�iD��Q.S��!+9*���&�=w�R_#9�����kX�R(^z���8�2�<ʶ��Z8oҒR�`񋉒�Ԍ���;|��0�_���{�"$H�YwX��	�$����ܧm�o�եLy�L��&=zzK�f��j��^c�7^�^V�v���.��qD���9�w_��y4>1s9u���]���c6�vL�� ��[#��O*�!�l�����(�M�ĠŬy�?�^�<dxj�o�q'��O�-���
}��AC�<$�� ��jݖZ4=+���]��G}5�����N}�`�ψ�.*�Nٰgi��Œo�
R����Mx̰v"�%�ٟ�����2���$�� 1tӞ�@���g�����A�e-�/�:�!���J�п���u؀�Y^�'���ۑc��?����&z��"�f�����*k鱭��ù!M^��ꛝG�� `y�r���v��ޓ�w\�9aIiyX���jl��܄d�T���FT�m�sL;����s���������CW�5c��Y�����8ÿky�wّw��8c�4�q>A"���n�W[���v)M�$��㌜�=N�� kP��@f9�!��� �Nq�L����=Nu�Y�qb-�b�',R��5{㳊��`MTu�GQ�z⟀��9��=���H!]�����X�緅�"�О(�1����^�����y
s�#�������ɜo�p���䇲���;�R�[����T��,�-����A�?�i�E�����h��9�$���� �r|E���*�R�Z.kdJ&�R�UD�6�m�zP����c���(p�G�� Y�.qk�@$�N�T&X��gg�n�,4���Z��=.~� �7�s	5N+�X�����.���l�� TxG	NNuCըG���?����_uF.��lY3?E�{ʅم��8��f�
�W���@e��ޅ�e�[�V��'� %���\����K��v%&z�U��2}�PI|p��H?1@B��~6�G��7�Wqb˟�M*#SX��}�!��3�(��ko(H��y[ڣt�mԠ-(x�V��Om��j`�<m� fy��U*�w[�i�2�'\����=�J���/{0�� ���Io�h�©����ŀ$��$ �����~�iR.��.<&����)���j�c�.[x���D�����e4��<���,����Q��T�o��h���ϣR��"{�v�8OV
�L��k�#�/g|��ӑ+政gK��ђ��`"��ä:��ʢKF����roJY�#0MNs%����2=u���vEe��EL�.ϸ�/���n`�ڧE�?���H�a��>���t�%��(	�,���%���w��N]���S��)|,ѵp��[O�G�u�u����y1o�+͝V������Δ<��<�g��6���
>��l�=:<-���3�Trw&�&wSl�
�&�Yɭ@��r`ȓ�X `�%�=�n��m�v;�PZ���<�&ݎ~��I� s\5J��X�i��� ��nX7�Ϟ#%��l��&	����~r�yW�}�=���|h�)�rSS�扉��er7
���� ��S�x����CBd9��d����z�W����K���s�zd�9-ء[��]�k��ݐ�eO��2B%ƈ�!~�Mo'��P�Rƫ��H~a3�8��on�9$q��w���^0-�z� �Uo��?���3���o������]�R:�t��L,�z��aZ(8���Z[�n�/���M�}��MG,�A��z0�~�:�ޟA��|V�>�d`�e�L�M���E��a��s\#|�u��N��Y�j-�|N��ݖ|�'e�@�?r�Y��My�/!�.����n@H�L��M����;���n��/��Uk�ःweI���
�� ���q�Ss���E����e�Όy.�x��+�"[���׫	��}�X:�����$�l�<�q���V�C7G��T	��y����aqͦ5ᄪێ���H��/\�S�Ѳ�Y�ʦ���OܠP�������[B\���2Y���۬z��| �AyK��]��R�0U~y�ߩb�V��)�N���fھC|M�?%��&��y��Qh������~q��� ���W���@� lySH���w��G�l�t������yU�xX����}����	E���A�G�E�W��Г�+�@�1ߎ��:aճ�����=B%)c8�CtO�w#�|�4�*k�G�W�,�,��%�0��C���P�/��!%�U(�y�	����������90ڔ�ɶ�~���83�jϑ�>�z:��"���3'�G_�c�!	ܗ�RN|��p���uD���O�'� �}o��2i�a ���o:J���Ѐ49aQ�H�9[��5��OzO�]�������k�Ī�D�b��<<v�����@5:����=DD��JI����+���Q��TFȖ�� �����(o�ZOc��"�֧�d�&����oT?n*�468��8�ɕ+x��.Xw��>��������[��?e���j2�(`T�6�n��PP! ��J�(zn[���L��)8rp���_h��rc%��3P�Xy(9�S)v/�����+�\��P{L˧�!Q�_?�N*��&�͒��T�s����H��蜹1�`�v1-��r��P�V
I����ZDͶ"��>��1��UP���Rb��JC��������i���<��j�K�����`�M�m$�[�R��ϑ��jKԦ���"�r@Sv�ڨ2<�
�F>��k�e�*M�����zC��4����,��睘�D����#�U(qu�t����,��m�G���%o�zJ9�e�~y+��]�j8k��h?1�H�g+���HO�E1������o�Rw��GHC��\�j�W�z�xR���/_�W![v!�3�AI�>c��ڬ[�K� ���)w���Z�G%5�K�@��l���=1�!,�6�_�'��
��'��t�>�z;?L/�U�Z�	Ң>�d���=K��S"�fTZ2�HA'W�JY�*�/_���B|rN�̼��b�gAb���/��j2�[�;�H^a��ObF�mv̼�v��{��j��5�?�O�a.x*T��X��9�{���4��[�W�~���n���)5Sn<���f���8����>(wc��^��3)�c���)G{���秗)�VA��@�6|��d�=���ƣ2�y�A5@�w�5�R����ةǗ)zڙ��;�T`�!v����pp�9z�#�S����e��a�yUgy�@�Sdf���T�XBbS�goaGb��P�r�GT�5H/ɳ�v������]���y���L�T��p����)���{J���(Z��Ң-A�)�o^�vʤ���1�すMȾ���j�d����,]l�"u��(�É�B{�#fP�iC&�=���m��V�þ�3��t/Q|��[$���U�5m��j��%��W�18z�z� ��U}�8o$%_�=1Qgg���94�C|<�&���?4���Em0w���k��x~d�B�o..�gR�F�aJ;d�Kd&�࿘��������:֒߬�ײI�X��γ��il��^И��8�s*A�b�_��k���@�)%�2���*J�iu�)���J�kLQ�] ��L�G���+����ԮB� K�l�LX�$��f�����!7���t��8hD�h�լ�7-��p�B�k�$|_x���NTǎ��S#]�|�A�ᐼ�!j�_��A.�ѡ_���ʻ�Q�S��
Z��R{��:�������^�?�\�~��Is�}I��V� N6!����'�涠��5s���_Ҳ�׾{ǉ�����L���n��� ϲ�a&�Ɨ��E����o���\F������:Mc�yn��^մ- 
�b��jV���(��Ɋ�;*��,��"]��4�u#��lS���"kT�#,���S�����h(lI��B��V9g�̘�F� ^2q�!X,���c�O���u.��ʘ1�_
}��S<�m�^�a�PxYﾭ��l�=V����2��	���o~S A�_���LΖ��*䀳�
- {�8В*����߷��nXV~i&F>�8��U�;O��&�(��q�g2B�*"�I�Ò`J^��*�A!�_1_�?�c�2�$�\�8�����T��g�
��+�˼�jDɮ��m���y���wÚ��C���P�f���@���	�c�:��O��t7�e�|z)�o�엒��P"��q	ﵓp.W�Z�)$�r���Ͼ�B9H�o�%7� �#����✕�n���A9��B�;Co�A9�}t���D�;��ؒ:��۝��"���C�H?9A�4 �L��jG���52�HJ_��X=�|x|�#Y��Y�.��V��Xk>��2�M��V�G����D����&k�.k��$g_���}gZ/�G����7��0X�YovXM�[�Y1�\���J^���na�CzQ�73_�/��wB��]?��k�]h�Z]Ã?�G��3��|�$���Ag� ���1�$�/ V̠��YS�c�Ct����R>����e�-�0�4Y�����9@s���=�_�B2a���� �4Qs:aL�3�r�5)�6�6�����c�h�[Ҟ�"��\a]�ݒ��+'<���\�x�y�0@�Z��cLQ4�j ��2*�J��f��*<�>�&*Ը������[I�2�fP��Hv���~����"N2�wsش��D�b#��zk��hԻ�F�ʩn�f�ׂ�����>�ܠ��L��'Un���;h�T[�8��]W�'p��fψR�7�k5��JwN}y��f�Y�!�Ir1Kq�m�,���.�墍�%9>{�)��>��L��Q8K;��{�%W%�v���|��^q�̭.dH#�{-��}lrߴ����P��Ӓ��{i�t�O:��r��)�4rE>���s�44�sw-�\mA&��R���9���[0����t�ێYn׼$��s{���/q�'Y8y�F��~1.]��ϰ�&*r�޵|��V��=�%�gR� �n�Eb��%y'˦<��we�3UL28,h@��d���b�<%�*ء�����	��4s�W����ί�V��%�Ů�1`p�־�(�>ݓ�����F%�� �_�����v�ru7���4���V���H1wj�i�N�W�e_R�l��Ǡ-[�����6�\�p⇖6��Q��` ʔ쳭�* ��J0�W��,�gIR�HB�kQ��/Ҹ�w��x��[a���~�=��cfpg%�i��E���L4�#���}��Έ���(w�kժ���F&}K�����4��+0̧;�N��1 ����Y����OJ�Ҹ���/������)p}Q�
����'I���U?�q�vs��uH�l�'�IF���2�䟚��{Pd!��U�Ю
=t��t�2�U墋{����X":� ��U�,w�h���-�Fc{�����<Z�9�F .q}j
��D�gD����jHe_��S�=��*;�i������{p��,�::>3�^�S=��}���H�^hd�Ċ��ha�{cHk<$��}��[8l���6���Iw*�� Nطw�z��P��@{��-B�&�CӶ�Ix�]o	��om5����+���[y!�X1�Do/� S���p�+�(��h�]u�����]�t�������)�ބH}�\�y��&�i��Is�#;�R0��WR,��	���ޙR�������=�r;��\:à�U�����(j�	�m��8�*\��p6d57p��RK�<��đ��1�<���o�l��>L��"�ʡ�u��ڀ��}1�g�5P=�G��ԡ�@�j�leV�Dn�Bلu�x^�vzrǩ�>��wQ���P»˰�T�����I�B��UX��Q3�R��d��q\:��\�O��Q�m�(�N�G(���l��n��g<|������1����i�_�c=v�4iY�ꀅ�'��̡עmfԮ�sTX��sM��?��4����=��}qU�R��8wc/)�7�K�~`�)6�C��b��ι�v�5��"�!!����cc��O�how��-%�	������Z�T�9AC�Aoښ^R:�����O�Bt��D[snr^�c���C�,��2�2N��>��*� {R� �Ô��]�uM`�y��Am</+Z�Ѯ�������d��	Itȣ"{u��� t�iv%0{��P>D�ٖh��:�{b���g��9Y/�P�Q@	�l�AG˅���%|�Ѕ!-lץ�<I��@�Q<���p&�cp�2������UGm�2�T9],����l��Hp�I]v�$z��i� �O��/�&�xgu;���0�J&���I�i��k�>Wף&�/"3��Z��lq�4�k�R�">�Rv�[�MjKS�0�N)P��8�n�нP	fSeƆ{B�wRArz;9����t��U������o�s�Ϻ�Dn;s� �႗�����b�B�m�B)*4QOoAj�{�\�o�^�Y00�n�5C���:'mo&D�ϲb��=�Ӛ����s��B[_4e]e��Ï4�m���ȯ�e���y�uq�: �)�*R~��������b)9��K�}��j���������\No�9[O��!ۋ-�M�Rr�.f2�-�/�����㙣5u
dE�L��e
V x���'¿�x�!>�*���=.s�u�9���x�^��q���ck$]&����ټԖa�U1���o��rj�HcT殻L��<�d������ͻ��#�>GF��֤�IUk������~뒣c�"���%�%����%�����G}�A����`Z(�xɒ8��,�l)LQG��m��\AȤa_�׎���p�[��D���,F��)�3���8�HZ��uKm$Zb3�xS�0մ�,�䭲�&�_�P<�w�����9�(c�|IT��K0")������p���$"�I&R����¦ �N�q6T5����mn��ZT�0�sw�AO�4�v�df�J:^;���]N���D�ce��֊���i0 ������aST��=�S���e��&'_�٪�Xj�d��uˍ��.�qȴ�P��,�xO/���LV�)��Э_�z9�5�����c# %9�{��8�v���O�E�i�a�z@[]>WTC����3T�ྠt���729B8Wg�oW�O�`N��	(RO�S!i6?y;�g��Z��dĆzT��� Nn��޹paj.L3h��+�������&���N3l�q܏��X��h	��N �����=��#s�յc*U0���R���i�v��ek�+��<�x����Ծ���D�;�b1jF֝4�dȰb�RB�G������<��сc�R�V����lM�&@uA�K��f;tԉ6�G�� ��Z��˒��P<=q��d��,=���X��)u�a�Dѡ��ޢ��(� s+4���vS�X�bY���o���c�uŨ�L~q����48�0���*��G����$?��!d�X��*h�/�J�,��2�l�ؖ�+�C��*EJBfR`/U1��^�鏛;��#C���c���EQYW�J���-d{�w��h�(=g��b�mu�s;��'���w�Vp�Ǣ�*���d����c ��Q0���8T� �����㧯g8畩��C�^yD*������ŷ��m�fivؔ�<G���켗�p�Z2sc�^�\|�
�c�?.M�˹̣x��N�%�ﭞ���@܄��u��G�B 
�{��(P��:/a���Bϙ���,�QR���ZfJdY�P�s��+��^���Ly~�|᭗'@��s��,ة���G�F�AZ\Nl��=�6(����\M��V
�A|��L��:
�C-{uyĕ��.o����Jyq��i��7@�Ⱦ���l� {�����e�Z}h��MDxkM�W��-�Op�xc�eЯ��}r�-=�c�o:#�p�_���^�
�����9B�Ify�-�}�M�����4�Ft�?����e���=]����CHd�U����J 瞸-C��/�D��3T���Ë!%�y��5 ����z����½����m&1�E���f��v�s��<�޴Ks��G��E
�d\ƾEeU���
����Q���2��B2z�����K�KǫPߞ�	���#	����q�{��!���>Da���k��(�[�\�j0Dn_)�٭�a�
G��*���\t�7-\����Ǒ��ARu;tX��Ue.M��\<�W�ˑj����[��%iñ����i�z0U�w.ϺE7C{�E�[�S��r�Y�0Σ*o��&�G�IC�4��	7e����P�L#�Х�E!މޘ&�.܉ĥ:�I�����n<5`�#�[�^�P,q�I�Ik�|�&�eBY���Ys.�����i�=�>������2n��)?Sc��{�Tl�A�D���.�a��*R���c��nՌ� 74߶��Aֺb�;��Z)�Np���$���;���a��w���kТn�?��,
Zf��W(����I�����~J�S]m'T�V[?_<.����a�vA+�1����n=u��7�8���8c�����I�G\����@���H2����GI+/���ٗz=�ZƘ���J��6�w��?�{�h��4�Ƨm*�մf5�� ��?�*[j֫��o�t��	Q�D;��NH3y-�`�k���CS�N��O;ֻ~�b{W���T!r뫽�D�Aam��E��`DI�vDP�r�$t,gWAz*"�����m��͡u3hutn"i7[��Jg�!��(̱jU���}�?m�s��3T�OM���|�qatd��0]w��f@9!j�#��k*���aX2˴�X \8�
�hp]^�s#�s`�*T���/�k��*��������������R�͵���S��<�gú".]���i"�騉ғs:��C^�J�������eo&��jT99�E:M00���{�9�R	e��%9}���1C�R��¨�+������t�]��-�i�;'2����2a~2y��߀]��K5W6��Z����VA�I!��YŐ8Ac����w߻�2�ҥ�40�r�Ko3(��y�M&)����.� i�>�8�9C�� �=uE�������a:�8��� J}�T2�s?'jڂ�{>J~ǌ�2mS���!q�����n�Q_�B�y�ն"nj
�w���5s�κ�n��5NT�����C�GB��I�N噏^���t�M����rדG{z �!��)�I��f�K_�0�&�]�mK���?|��4�CN�l�L��-Ĺa+� aY�p%ХY�l5��r�0<6�`yVԤG�X=|Ux��}>H?U
��[.j���P3�zT�=@ۤNB���*�_�\�8�V�d�erWT=�/�:���c��mὙ.��۪G���4��MrN�к�&nX\���� ��bƓ�b��V��Ӗw���A��b1�N�,)CLY9��숰 m�#-����<�qX�$��U��� �>Ix�|n��_O]+Bs��#�;��i�QgE>O������P��B+0�»��9	<0|b��p�;D�̱�nY�S�`$l~��|&❙{�S4�Pd��y�z�wmO�!�zr����ʦ!|�кw�U���y
��r��+_֤��I�J[�4�78|O�N���~	��+7�g�~��.ty�q��ąӀw_�K�Ӓ
�_��HrJ����� �2Sf�J+���׎�!���S���G�D����3����t����I�����'ļN�GP����{T���p�*hNh�G��4��+"���"�J�_s�����[x\�-�g�K��<��_�ͤ"}�Ӝ̋o�&{���=�OE�M�"cn1�¯�d�jyx��v8ȴtL�PܹP$�0R�k��%js�e\�j������О]�dn`�8�
C�+#k�2qSU�?�SX��˹�6L%�QQ���0��Q|�m���ysb_�bJ���_�n� ��DѾ1�������֠�f��$m���5���㺏�x5�s�r�/�O��v�����`?EHI�6�z�INBv�=�����4�K��ʖ�j�AV��(\@Yw>[͌=��,"I���n�v �	����:��Q2�	A ����w��,?=qnJG� F�F���l]�7���j	(��њz�G\#,�?�[�J��iG����6T-��g�,�qF`	�%vb{b����;v!I�<[��lz���&NB��^ca�T�',F��7���e���
)��ھ�K#�������JO���gF)�H��]�1�Gr� J��]f��\\�/t������7��Ӱ�������ڄ�js ��F�Fi��G;wٳb���Շ`7���$ԡ|e@6�N�k�\�&���]�wH��f�?��=VS��@�r.d�ZG����fQFRXB5᪐3�J���DT(���Ve�l	A�iͧ,g'LA� V�>�at�f�N�-����૤RƲ>wJ���*�5"*����	�~�t������wa���5����^�fL��٧l���Z�����(#���;����=D�}P��[e8:@��L�EvҬ�mV8�ji���� �z��/#,�⠥pZ��;1��]<�6,v�Q���ǥ�e$������]���D����Mw&��'k��3��e�������d���i�<��k#%>2���wjL�g��Q���H�j����8(�K>�St4�9�V]Y����E��oD0�3��@�=���VZZ����^���!��-��Ű=�k�y��"�T�%+�\H���$Mr`��*�]��0������F&���e�"ъ�*&ئ'V���q���$}>��z�5 �On �����a��1Ф��'3 Ge*�HE�KW�Ђ/T
B��؝�l4�̏���j���4��'X�:vY�54U7��e���ʦ�%buDg���T��r��'2�1�m:~ұ87P����Η=e<GSeǮ�}ߨ�G��ͼ[������\��}M=偂�"Ì!���O���)�ǵj�:EOٸ�Qݪg-@7k4��@��g�2D蝳��(�a�H+·�?�VTUi,���4O�oe�^N��`� ������O��S�4~H�=f�^��Nr���jx��.U*�e( ��j��H�XA�cg[�뻞A9��2�����$�%����[.б��L�"6>�:B ����r~۩�_������-X�LER;�r%o-��B'����u J���S��.j�'2 ��$�<R��D*ݪWS`x����""5�J�=e�j�/Å�aD㒱l	^*��v0_�p�@��S!�.jq}"詤�����_3-G\%}��Q��������h8$��M6(�j˗옅���3`�%����:�=��Z��i'!�}�pf6��p�����Q,<�N[3��)�A.!B��d���װe�|ה���?.�>��9���t�/����
x�v�� #���^��"~L2�ӵ?1�f��X�&��ͲPT/���8[�h�♴[߶��c<h��vl=Ba��(9 ^z�X 򍣫���%z!�ҷEX"�+���YG㐃�Ů(�2x%t����J�w�*�U�a�c%.ƶ����[�1	���M8� e{^מJ��q�pu�����WV�
]O����d�TV��t�d/p�mN��G.7[�\\3.��+�dt.���[�����j�pǦ3	���HYP�Mkn���sC�{��N��� ���+ҩ9'v�4VYZ⹔ �r!��g�9�h�H��%���c������T����L�GS�.F�_P`�-��*�7�=3�_#�ҝ�jĽ1w;�q�`+c�Z'�b7A��[�i�e�C�H�^_ �(f����0�������s��8�^s�$}��@4�J_.{�{He5��F�`Y�ۅ�� 1�6�zbb �'�^Lxo*�hg��}+	lχ�K�%+�:�������u}b|핾�'������3�]RX\���9���Ⴘ�x�</]V�嘾J6X�H�N	q�|���) �v�/ޣ/Q�^WȦ��]hfQw��%��S�+��m�����:o�v���+=���x��xm�v�j��{�c��͂;��G���]#��L]�\Z����(�����Tz_:8�B�%��	x���!(�M�La�M�ы5r�"(b��������+�˵i� � �|s�7��a��f��P��;Zz�BbY �)���7D$��m���NR���F�w#Of�5*܇��fEͽ���?t�
����P2��P�����q��h�vP�^�]і��_���	������T�+̚Q�֚��!��_�M{F�2%�ʠT-@�y,Ĩ+���R~�Utny~^�Ǌ��-�rz���<��d4Zm_�	b��Z7�F%����p���J��a��� ʛT����;-��"l��{��C�q��*�/2M����CUG&�O�E_��1+;L�ow�*���l����_@o����ٚ%R�_�w�x�)j���Fq7�S��e���h����z�R§��MC�G� ��g�f��F"+c%��0�C���L��Uvg�|L86��ri�Ρ���A{�\����l����LYAd����ɰj���],a�mx6%�G<���2���+����W��c9}F�PWp�_�G}��s�]z��b����r�8�phc�b��/��(n2����̪>�;�������x�t�5�.��O�t�D�p��zy׬S������5KqM��^e ��sI�	"Z�2���&�'C� \�&�%󔘛8���{B����,R]^Qܤ�ԙH'����������dHg�z�(��P�?l4��o�O�I��<'�� 4�F��Ӟ�������^�_iµ��ֶ�Qp6��c�9������#�mRn��b�kG�~B�\�7����eǎw�֧�$�J�:C�L
���	�N9�~4;`���w�P9�b�q�n/GU�� �0�9�"����u|���-��ΰ���4}vҌ�W��N1�{�#[X��H7���Z@6�4$O�+jQ����Z|�A�g �Y*�\�Fŵ$�/r���f��d)�X��zucd?�չ���5����fZC� Y꣨���gj�Y�K���{�} &N��
m���ϪF�Km�~-+<cZj̧�����Z�`�1���7Y���
�m��_Sxڦ|������2�#��~�eX]�����+�ٟ�{�O������a���e���;��͘ @��\����J#+���*��peWD>��������S�Y'	 �R5r�rڀ�����p ���t�zJk�z�o:�,W )J�ޏ�U��Kl���7�ܛT����@�:P�w�������n8|���ž�Үc[��3Zm[17ֹh���A���%�O�3f�C�s)������C�h�	/E�9�r��?��QsT��6�eIk�õ�#a3>��R6T6tX8�9|TT^��V@|Ur2C.M�+
Ý%]� m8z�n��������ڟB|@̗u;�\[w����k'?�"�����C>S�>�ZTmc��3�FK�6�VPO$�C�d>�yHs�-7t-���,�����F��h0x������T7-y�5 ���|��A���ﻪ�ﴴy��5��kf&��]j8���r)�#����=?�յ4 ��/���+��C��M$M�F)�㾎^�o� �`/�&J'#�F�M���Bs�6�ڞ����ta�x�V��v�.��4:K��`�7(�}8wWW>��l�f�Bf��`��w��;�-�'��Ŕ�T�n���8�sXѪ���?A���f�ۜcx��E����?3�E�պ�ԑ�.5��	~5���qFJ�Ѫ�<��˛��hC-��RPL�$)ʇu�ӘG��i}�SRD~Om��G��	�e�l���s��Ս���>U�V:dx���#N��ӫ>K�8���v�5��d�2v9~� U$�8��b���((�k�K{�[X�n���\cI���d*p7+s M���_/G�^��PϜ���!� s�4õcD���r��k�c~�Vw]�R�����b+!c%,|�ʢ��gy�X�`\\+�fd0w9�}P<��IhHb�JM��������dF��yL��No~�i��Pn{|�A�rh�*��֒.��}qO[��w�hwC�x�8i��(�B������H5�:�V�?!� km�φ-�e�{ɐ�N���
�U�z�n��$�h����q!wb^�����ڋE�}z��zW�����0d,8�<0ce�N�f��m�H��!+�;�V�q�Bn�SO5�j�A�k�=�u�/���A#���@Ni�ݓ��� w��)��\�����������9-w�6�Z��]�S-������~a��#Z-*�q�q��g�
�@!8��@���w��]0mfCQr��J
I���qS�ӟ�9`�b�_�#������v�i�4W|1���B;�V�s'��ٚ��{N��i�[�y?�3�@RA�Ey�k[��$]�z�E�WA���x��	O�B��8�ه���\��>zh|�b|����ac�.���f�����5,��F�Svlũ�1B2ÒEM'��pGvCaE=cAb8œꉶU"��vftk!�k���n,�&�g{�7.DM0t���}�ϭU�MC0>�潛�Qr�Ϸ]v�!���=�I7��W�\
�d�J��M�	�7�`ˋW��YS��14�y��I�iU�����f��s����Mi��j��ǥ�Qg!�O�X��d�/�;��Y��_�R��LQv �kĦ�`�J��*��A.2��d(	y�}�7�����[�$v��첲�dBuKxvx`=�}ۏ�D��a#�;º��Y���S�kDV����+Y�(���v�:<�cԿ�J�����1�3)�����<��,L�׼Ik�Ļv�B���hE�J.�wj:$�5H�%T���(��'�Г�I���	���U���Ϳ�m'h-/��e8�u�s����F]ܴ.��~&����[�׷KH9,�C8�G�`��f���|'9��6�0�>��ذ\�MT��ċjz��D����c��_O푲��_���[�@����k��ײ;与���;Jjd������w�0Xкp��͟�4�0����JVjk�;��#)L7bK�e�G2Iլڤ� �n��*�6�8�Y�@�_��������T0+L���ǻ��q���v|{�*q��E�US��=i)�­a���^d�n%� ��K��O/�_�]��}! �`"�S�S<��Fj����R��t�Ĝ�1�#�?�S��DBS�&������^�kW9Xg���2��tǗl��M</���I�D����@�KdXc��tD��ѣ-�
;odH�زl�{��\�asY/�:P���q�9|���f&e����A�
������\zJvq��E[�rt7�f%�e�zm��N0u@�98e%u)M�bq��_lV7,�s�����c��VX�,�X����b� }qslz�֒�EA��8��i�tҝ�����&#��^�VuR�ín�F�0)��?B\���	AUt;\k�ω��G����%{����<#�[��0�<��]n-��a��->Ob��<ń��jx�]ל����x���SmgG��Y�e���^S�nS���u�S��c��OJ��~��	&뚼�L�e�U�V�ń.R�@A*� ���~;R��*�EB�q����it7��.=7m�0	��i�X���(EO�� �4��`�%��e$R�W���<2��Ɋ���7h�V����-θO����Q gº�yzC���K�]��"a��?����@�r����o�Á^����k�9X�e{\��ST��p�t/MB�ڳ�l�c�uo�˔T����y���<O��.*6 �e��4C:?V=2Z���~�e+��\��=����e��3ꆊ^]���?%4꧿����е�/*���a1B5:Y�� ׈�@�b#�O?_:s��<�>��1��q'����0�Ff��}�/X(�5����;�FL� �p
D�÷����g��0+�(,U���B}�c�N���}d���=s=o�*��!A�V:iēvdHi�Q�J��|<o��#�s�犙{j=�>��..���k�-�g�#�7���s�t�?*Ի@O�lh+��5X�;s@~�l_t<�'J<3 :��;o��C+�L�Hv���}��p��n�GA�fT�7�肋1)��:�<��j�>>/;���.�ԤJT$3!��-B� ݕ�W��ç���9���� N��6��r_�>0���Yޟ��ZxP%g\�[h͜�?��������%���zh��: �����a)?E���A�]m��,z�7jH����2Ih%�<�)&�ӁR�<z�Pn��Wޜ���N>�ٌܔ�$�b�؝��ƟG��ˮ^&��ˈ�3��yEhE{�@?�4�e�ZX�XA�f��������}�4�l;b�T'!E?�k�1s�Ƨ����B�t*�ࠆچ���T��{`�z�R�Ls�Y�Bz���KHm�exѨ)��_����j�t�`�y���&��.z���M���^{�М�YR�?�y�Fu4?�Yf�#Q�
��ӌ�@Ў���X{�!�
> e�}�"u#6��EY����on����I/��DCY���nH�����p��}��j1�=Z�w��)��B^2��J����������AH���-�';������%&T"��|Z�j�JZ\�a}-����כ�'%�P��U�؄�V,�b̦c���`c�Iob��LpL�1�pM�q!o{ Y�������qO}� �K�k�7+��ol[\����Ĥ�]�'�U�,&G�Y	h�AXc��&2^I�5��"�Cܜ"s�iܚ�Kg������N$G>�K��[k��;x��j7��DF���oZ"������*��m�'p�߮G#E���=���sQ�^P�㸃���+OTym�:��x� 7䆞^�RH�]k��v�
���BB��C�I����+Wd$(�����`�0��(�����e�r]u�i�ݓKT��@Ϩ�%� �L<ـ� ��|�H<oӌjK��1��`e�[���MB�u�-�z8�_ٞb+�#�C�{�v���̓l��b���+�&d��둅mO��a���o*pw�G�m����̘�m�"�������0��c��?���@*�r���JԜR�1����c��f����xvL��_�m���(~�u�i8F���j'h�ER������xz���O#��o�|�5��U&�o#9#�"l8�D�\HD�}�E�@�%���R��Uԟ��T`C0��(��>ɚ
�L�F�=P[I`���CWk�p���WE���H�#����)�Ҵ��1�j��0�4�#�:}}9`lQu�5�~r函f�ԣY�A�6}LvR�ǟ�q������5�$�o͡b��FsQP"�=��㎳e�9�"]���ĥ��k����/��Zs�����H2"ݕ>o�����vf�,!D����L!@�dBū�	�=����a%�3X� ك�o�/6ܚ�ц����K� �Pk�)O{�ȵ̓��<��P��k1�i0�.��:|����	�^��Y��0�G�����?�[�.����^�=�2(�|��XEwJ��n9�{d,��,�r01�B���DQq�L��hW���z�%M� �BϦhĎ�1s=ٗ}��d]l�WJi�8�����#L��J��I���ξ�L����� �^�׀��c�"���^0ԁ?Pk(����������d���\���?|p!}���aS������q��w�C����#�{��bA���'=������m���M(<�q���l��+�l{Zg}]"��B�:�ƪi㵔"���tN
�I��)$gZ¿����;P�Z����ބ(1��e�/N�z����Q�z6���~XpsH�$u��@�b&"��cI��d(���:m4	�[c�
ʐ1�T������?2���f(Cb��������B�K>�q�)��˚�����o��d�Kr���%��&��(?�O��%	���c_���|�3A��a���(VC�������V�_��u=7߳����w���̀�9�7�ՈjJ'�
hRV��)@�pG|��SFu�d�~B��H���}xa�o(���8\s��_��3@�e����}�)�3���W�g��ѱ���D@
��O`{�v��џw_��]iS�ДYr�$��J\�L�o�=��Y�8q]���K��%��~qī�XA?��#{��P^r��}>��7�˃�QfUJ�p��Q.ָ�B�|�`�c����~F ��I��,3iȴ�L��qT�Z��$�zPw	�&����8߬��M�_~�=A�r��/u��m#�^!��ǼJ4NFB��p�JcDE��p�՟9>l����ks�_�J��_�1o��!Z��PXhn��y�����g��0M�m7yW��8��n���0JȞ�5��4�ui��$sy���M�I�<j�,�krw	}��\��8��q����M�+d�"�
�p�C>�9�«<�6=a�]����M�u!`��t�,���΁����'����-Ӂ�������$�	]��9D�+*��oru�S�����m!ۨ�YƄj�]:+�G�A�3��q����ǘ�c�1����AR	C�h�߫[Ψi��v�+'&p�nr��գ?l�#@�^
����d��W^7��1������疹�g�W4@֘ӑEHt��?5���b�!� v�g�ɗe.0:�@5"J�D:U=|�|D<}@7&�^�*k��A�ϓ3%R[��C`���-��^�u"<�#�����U[���V�3��QD�mk�a�'�+0U��O���p��v�"�@t(i�x���VZ2�[g��l$��|�6iM�#٘�S��3 �����+��5|~>}����|��nl�l�zM=�����
(U�{pgE`����;���f0�u6P��m�@�#�g?�YV��)n��"C�W����W�\����&��`u0D��a#�Wp��81K���,�љ�����ABa�G�;���+鍍0�սd=l�h�C$�#ʬ�;�� $}�(w���?A��MĽ�$�itV,`∛���Y��e�E?��W��z��%��i�d�FU�b=+��^��{*�wPD�O�r�Um��0�����wbP3f 	Y��"gn���k�T6C7^L��u�R�5��a��?�s���C�K��F`)����	�Gg1B1)3;y���fEh}kN��B\YıAq����ԳK}��	��Q�9���[��oL��x$]Q�sD��ыT�ކL�����|1�*[���JiY�K����)����w�G��P��g��8�(���>�d� n�c�B����F���:J}Ľ2��!-dPp0������]k�%��޴���D�G��=�`��<�#����w����U�¿�=Y�D��d���:�Uu��m���'��u�*����r&�K���Pw8Cv�q�I���q:g0ٓ�u��O���d ƀ�:�K�ӕ���Q�,�jV4~iߤs�j_wGk:�S�)��@u�k���͢�}C%^t�%1�A�I����fe�^ϬU늳�y�}�������XW\?�4�@������l�>A��b��*|��-vpˈ�m��Q���E�ݱC{I"�bn�E����h�rMg��`ĩ�O�� }�­�C\���c�/��h�� 2�	 ~��:^����:6��m�[e�J�|?w�#�8��+�r�]'�{^���v�(E���w}�ƊI��~X����pЪ����&��?���<^`.�(�{8��/���Ы��x~�1�?�6�VG��6�.�%� ����V����(��	�m#�r]ày�ڝz����T�[8hL��������qk&���粟��Vm�GP�a_�J5�[��X��]�����FM�(��m��nPMf�J^��I$4,N��Ě�c�o��D�G��M<��f?��p��Z�ӥ�W�E޵��m��jzc{��������ߏ#LN�5v�XG]��mOӭ��j�z��̣X�ŁQ�Ζ6"QjO�1Ѯ��Z�$�
�j:L�^�礂�$����Gc�'N�뢧���8z�r_��%�@0�d���`��2Z`��<;L
�Ս4��wW7	A/�����&Mp0e��$�-%mv�"ɶP�x5[qsϸ�]T�ッ�{���t!��i�v�D�K	u�:}*}ǭ��^�L�*�b���W�@��l.N���`��Z�v-k�U✤�cZI5�o��yc��>�̙0N�CbLK쌰���_�_]yϔ%h��L��Nw�8S���Y�c9��I^�%/`WdX����>|���c/K|! H��&j�/8��͙�����I",d/N%�G��wc�}VM\҃ŠqhP/����-&���־���;A4[ϋ�XAN�d�B%���zm#SkΩ�- �k*��Q��Y��媰5r���߭w�:�NV2h�΍�L`T�S��I�7��m��χ��uE�	�i�(�������@وVZ:�Sʃ)��o�2����I"&)l��/#ߍ��e hW-a�=F���͆��q���rA�o��=!�j���P%�A�Sv���Q8S�|b��'�4�%�G'��*��,-���M�:�V�<����O�J��?D�(�S�k�3��@�Z�d8�l�'���~/�K,"X���=>��9[p-6ۖ��CH�F��������T\$��K� %.����;��f]&5���~-�C~O��1=��c�9|�)�� ��\v�@��}�@�Wlnu��4)`eץ�*�_�+4�����+�8|[G�z+=WU�k���8�xi��ۯ��}�a��v��-ܟӅ�E����1�s6`E��s�.5a�
C�y���<�U��>�O�]��_���%ǧ��y�>�)����k�%T��.0�ó��ސ_@���w�a���^AX%�!��߈����-&Q����=�lJϷ>v(#�f!a��2��2&�Ⱥ���ͻEP�FK�:��&��h|���P�ly��T׾�^��4r\���a����
}�,��]�$m�"��r��@v���_3Ǝ�L������^gN�����2����#��%�bh=k������qa� Ȭ��<�aA=%�K)h�gb�6�Z:�f�P�Fs��Lu�����3��=�ki�j�a���ߦ�^<�h'A}e4w�T�|R�\��Q�1Cـ�|d�8Xڛ�XXe�Զ��-/�~d����`e��O0"ND�j7If}No>���19DP�E'];��&l��ɭU�ͼ�a��Гrc�}]��#�e)?��İ��0[��We�z�P�w[O<z5�����N�D*�ڠ�p��tH\dٮ�	�o��ϤV0?n�m�rέ���/!:����{�tpQ�[��,�M
� ����+hԚܦP��j+L��w<����[�)�_��2ӯߝ��q��$\���+NH&���s|>h1w���	��MoёdX�u�N���	�� ]К�I��ѹ�y�D��	~�nyo���4?�@�T�Q�T�ه]�_jfk��U�~�]y��C��U�o�A ����&#G)�β��ON(߯�W�d��z;�p�S� � ��N"vv,n5���	X���)Ҳ
�v��A���"�40\��2���[!|?�KԻ(�ѹXF����;i!w����Or7�\{���V���?��x,��f�'cf�~Oi߄`��5��yP.Ki��['pO��Jd��`/L�����%Q{&)�.5P����"�,#�E���q�GHJCK�ߓ�qj�׋NP�)���RA���l�1���7gJW�y"8܂S3�����e-a�90>���&A�pr��ۦ!"I}9�y8���{o҃aKϒ�'�%t�?�>��(��3�q�o����p��?��]�POP:�l��c~������_��C��B�o0����!�[.̈́�)���N!�7膌ðĺ�4�n�Y8�F�,q�f����W��,1�LVs�8D9"h���O�ݐ�|@���� ���[�Dh�Ǉ��c�RRпv
��r��I�<�����C�R��׌�
'N����頧��z����缝�"}EElᙀ��ɏ��c;R���}M�6�O �Dr"=l6m(�"EJVB3�Q,�?���=��x\E��a�%Gsٱsś�c2_s��M����+^�a�����7��7R�@�B��`Eĉ���mIt��A�ca����}�b����d��D�+0�^'+�j	���z_{[����QYUÒ��c�����jS7&���D>��R(��7�|K��؟�H_��k[��Ȼ���Q��k�����D� #S�T�V�f����x�)j�΀��l�U��!A�d5n}���Z Ik����9ۏ_ II��7����q]��w��ȶ0F����q���Z*��oUi�X4=��v�nm��:G<Q`G���� ��?H*gT����ٕ���>���{��͈ y F2������Z[E�V{O���I1�s�*��>�C�6cz<��v+lN��F�z$�bU�U'֥��� ��:ɯ�$̚9�����Ν��fy���@����l
�g��A�r�\;;U�_�Ɲs(!�@�m����8�$$��%���oV��J����Y۫����Y�|e��Ϳ�q���4X�Ս�?e��c*>��s�AV:�~L���uX����rD,�Q���TOo��F��jrW4Y��Q?"�ahG�5(�,{T�A��	��RO˝�AV~���?�5�1�l������ �kT�y� ��wea���W�.����)4����'��'?J�0�p�{��n�N>�m)�Ӧ��$�b�w��
����%�u��F��:O0��B�7��_��葸bn�:Z ]:����02����L��o��L��1Qn&���hgi����4ƤM�E��Dm�i�
�-��}���~tt $s������T԰�C�<��|n�kբ��iu��^`�Uʚ��o��l��ʵ�O��$�&���6Ih��_�UO ���N��C.l�I@Hk`��V~���4�r*`�ֆ��X�2��S~� i�E't;��.#��0˽�xC���xp7�L�Q&z�o�t��	Z8D��n�#H�W��3rm)�o��J"D$ؖ�|���Ì7Ǒ�����^vU��k�������g	�\�~vm'��)"$\�/�G]���?t�"X"8~1b���L��45�)�Ӆ[�c�o!@�������[���/]/
�/0bZ���O��G.|�5+�v�v����̘�b��U�� ? �w�vYoC%��9z_ҫ �dL�� )�h[��)�잛���T�
Q�8hW��鮛
VH�����3�+�2y�-��Ri��g|,����T��;Z�^>vg7�p�������\���fp��W��;.Rcم�z�%����:0���8���h��]Q�Y��A�Tt����6Ԋ<�D0$���'\23DfȲ���ps�g�D�g��D�El *��h7��<�sp(3��P�<D&C_ɠL%�6��Z}�U:��d������/�p�r����v��T��>��B�����Z$�x�І}Tرu*���E4�����L+�����YI� ~k%{��#h�} 'a2�5S	�D v'�;���x�X�@7���ۄK��Ƙ&_]:��g�톶��~b���wq�M@��T0�����G�ezͪ ����������2RU�uY��v��� �������?��P0��|��� 
��^��s�T̮m�g�*����j���'�3��73��J�K�s���ߪ?3���]�2���C���y�9$��a���Fu��r�\������W#iHa�nle�Ѥ����/���^�7"�Y��_����&��M��:���2���L�&Ȼ��}Z	�þw�W�ai�4��y)�!�dJT��@2dX�ˏ�rzI׽F����=&�M��n2|Fh�dfAPi������W�2C^Ih>�j�;�(`��
�I�����Y"�,�F�f)x�vc��o�!��lo\F�μ1�@ٟ��]���K�ʲ�'L�-ۆ1A�e󼏉���#��۟.Y;9��e.�ŀ��͏�	P��덂r!D[�����H�� �|��,Į�M����~�����l�4�%#?��{5d�/f$+�/�S�ll8Q��P�5T�H��v�p���
�^c�7�0�Tʠ�8n�������/�=��M��<i"&������������{ݣ}su<��R}|ź�K����r��MYG[~ւ?yj"{4��g�ޛ߀���px�Ϡ��ܤ��mV�#O�C��s���`!\��éj��ت�g:�yY%q}�����VE�t��:�+P������1dI����q�����3���.�ɩ1?`1WՄ�N�C�\q�u'���ϖ&wK�F���5���(�/fY��ؼ;�޺N�؇&H�,�m��{�w���[Xvxx��7�{#e��E8��d��'����i��"�4{��T��dd���}��k�lҰ�����K*F�L+���9u��hm�dS�[���^h�,]��m,+ܳ�b���[��
CM���t���H�qGh��~�:靵�w�iBFFVi�@�؉%��jj�A�U|l�Ѕ�=f,aɞ��1ٕ��/�OO��<��==|0"�J�;�,	�e�nO�qTֿ�r��	v�{ۛ�A��ʭ.8-�"��Ŝ"��snޝ�+�?�?���B���#�z+�ZӅ�ٝW�\g5&W��9n������w�غ�	�m�P�O�������E���
�+4��Q�:��L��P7�C1W��-�y�Oھ���z9��Ċ������2��'I�RΗV�GN��[������f3�C�H�̛���ى̋��_dӑ]�%��D��"4�<촦�)F��Dk��|E�����]��<Z�EHe�q@��X�����,��K2��`5��5�P�l֛���:ܾ��I��!�����ד�zb�߭��)`*���K�0��:=mv����ҩ��!�Jʯ!��岋!�u�Ġ���VY�N�`�۬z<���Q���]���q�rҾ#�*Ӏ��fwv����lz]|��U"��|�� QkI��h,YV��[�����s��B�K��?Gl�>td��=��۷K�	�	��ge0>,�s�z��iS�?�Wm�[Q�uaM!�% X��_EI�\����yDO���W���%����@c�*'f�x��d�lJ!�3�4�A��$L���ń�N鑬d].��\;m����W����d�sީ}�HW�2r�o���1 ���SW�U:�,tɆ������HLbx��(�Kv�^ޠ����P_�FeL!տG��k�G8�E��LS�~���-��1�5�;gmX+�8�lD�C4��0p�koa�yX�mD`��=��CbD)/���?�y
�\���L�-�o�"p�	y����:]�JF�B�`b d�Ԕ�*F12N����26��%��4Km$��K��O̱��V�����K� ���*g�y]�Ym����B�! ��I���B��,VG	��v6Qś������(�Dlw�I���a  �~ �Jx�Xh�������Oŀ+�y��.Ve�"��c��zl��O������yI�a37���c��}Oj�kU�R�$��ƹ wqH����hwO��r�,C̄�얖���<!}8��Y�:�ݑΖ@wx�)�C�m���rJ��*[:nR���33��7�ţ�U#�u���Tq]=�����S�4�e�p�or��K���Cg�Q~�ĉPn��Yo �LF��v���q�� R�
U=N�*B�i~�`�;�eg�_���-��b�R��&��>�]�*M�ό^5��To���\��"}��hp.}��@ �%�ݭ�SZ��H"+a\פ0|#�����'Ǝ�nP�E�t��:��<�	ڸ ��֬�8պp��XFi���e���Ǫ�~h'�X���wyᲀ_B35G��p�]=KOS�h��D
�e,|��k�
�Q�(�!FB�^�>*?S$b��֫�n�#�RO��5�8�pʱ�e�G�1]	�#lq�@S�Bw�r9�AJ�P�틬	uDh"D�"�+����D
7��v�E��uM�@r�t�lG�iӦ�-��D����T)��<t4�a�p�8K��k����UqU<r��2���Gܑ�������6�W���Z��z����j�Ąq�ݢ�����0\I��=ʂ볔�5��=�+{E7�،�5ND���29A���\9᰾�%������疇�gM�&0�S��5��lV�,sy��n�vwDwKd0��K{����[�M��g�k�~ .����ʡ=^�*�fhD��Aѵw
X痆o%��4��P˖�k-K�m��D@�o�_�p��3�[���x#h��v	1������{�������Gbٯ5�fkΚ��wL�%L���/x�	M~n��X�M��8Cr[�*�:[д7{4��E&��s��M~�YK��?rϒ뒼�ϑ"��&���PKXS�"�M��OO��I����>�#f&���'4�T�����S.����s�C���Z9kkj?/t�I��I����O�$sX'��J4��V+s�4��9a�����)~� ��u?�j�v�C�湖{�@��]W9C� ���/|��Q���
�W��~g����<��(Yރ�1mpT����X:cK���$���s+�z)Rh���|K\L���"��_�+���]|좂<�[�V��yk���$���K��M�����d�0}TP�i5A��e�,�BkqH<>]4�K�i���m���j/�׬>3��z�u��s:1������[�����V��~����=s�-��zF+��g�xVR�io�t��)؝e�o��6�}Ƒ�j")Q�R0�ɢe������.g+-v�T���)gؔ�����y�[p�훁l��`!I�'Q2�٪`AB\Ι�8��ߞ�{�=��k�Gn�f�R��G!Xg��y��@��ɭ�f�}��=0ä-Qw_�jȵ�0�썼�#{��&Pj�"�\�,'�DWD�W��I��#=\��� "�����E�#��l�p��~o�3�a�r?<��-�;�2s�dwF��V#����x��Q}w(�2{o�a���m�VIx����(������U��X�Z���3v�CAif(g�k~�ʌ��L"`/���֛���@6�� }���2V�	�nMs)�%�����Ji�=Cj�e܎x�_u	b$M��T���1�����X��&�F�FӍ+�*m����qW�M딵��{��p���T�Jbr����a2/$��dwZU��:%2V�Å�Mf�%����� 6Y1(�-�'d A�x�R�L�oMTf�+B�����+(��Π'a��lʱ��O���:GV�Ν��p�S�|�9���Gf-����JУ=��+9G�ހ�'}rMD���c�.pn���H��A4�Eq��W�)��䭼[y��a�@��~�J�H��Vf��~��W���Ù��!�#���N@,q;zsY|z\&KqI�rkzyŚ�:԰j�'}��9+ �w�#dc�BnBh�^�ͲK��}�%�e)\lY銷�Zi<�h^Lf���)RO(v�q-���8�R&UU���,�'0V���F�5Z9��Ү�&�fk﮵���-�]���6�>���
{[�F�_��&�s��F���r� �1Dn��$��~� �����&�}�����:狥w�N/G��|T�^�T�'��P��V&�r�9A��W]S��
���]6�5%)x�e1r{ۮ��O��L�(0tW	��ꔷ��ݻ�?�Pw�J	��|���t�^pc��gxx����##��&P��[dO@-����m�|}_��5��m͖�� ��~Wx�p��z��3��x����n�/�)��g1�ŨЭ�{�y6�y=-�s`�Ǆ��>�8kU�YqŇ35�7j��@G�=��\]�^�d� t �,���q&#�IX�ɿp��R�{�Ri�p�Qcd�����z�D��I�����
����xYt����+`�v�H�I�'5s��bp��$s,6K�A[(������`�^����i��sK��������`%eO�(��Z�6m>�
�� ��C�P���tj	�}�n��N@�U�=��)�1�W�'�@ykU7cnkU�5���Ȇu,G&�[Q��}1L�"����LLlf"X�w�+�R��<1�2�w#���vǏoR/���N�
�
z���.�f]b��ͭĹ,W�m�Cb�4-F:���%�^U�l^G$�]���O�2 8�|�f�kB`��BA���೭������X�t_�?Uu�/e{$	b+�v��RE7c�#׺vz�qs��>6GG���rNzu��%�f|I��ç�Q�K�T}u��٦\�kӰco�M�tZʙ��U���������h����������]�^2�Ȫ1��k��' Մ��{gv=/z#R��kՍ�t~���΢��c�Ӥ�x�V�K'PZM����?�8{*V���5-ȃL��1�؎���Z�𤽭TW�R8�l[и��2��[�.�z�,� ;v�3�1�m����S�2Y�ޡ�����)]ɞ'�y[��78NUj'���␼ב�Ļ�gڥ�^,ϐč��
-����;��+��`b��_i'ι��D��X��3�%e׆�m�<ѠAp*T�H�{�ft2&s�������=? ze���ز� 3�4�Y�7�>Wj(�;]�DH|��Cղ�R�iv~�(�����E1 ��g�ޒO]��l����7� :ܝ�O�-�Bj�iܐ�Y��>��Zm豫�.q�QW"V;���/����Ѿ0�4���厢�BwTU�H��񦗩�Aն.*�,��"	�ڻ��]��QBo��6��1�a9�_��:fFPw�5N�	�SF���&n�:Eo��سͅb�/���w������	b�Ùqb�r�rw��Y���i�@_D�8��̎U��;a���X�#�_�G�lF!^��y�����~���x�GxyD]��͌!B��	әǠY�^�A���J}E�������(Ӑgo�{�&vY�S
��"J����_/m]
�%��$$����WF揖-��^a� } 1�8|=� ��C�oLEx��a��}{�s���ct��m/��X�%���)!��| �����k��_���ؘ���~�*<��n:M�mǃh��^��ʻ	k�|K���otߩ�OGc��;�%�?���%`������92g��ϱ��9ߴ�U9ZJ(ˠA�A�ۓU�q��]ɢ�(ȇ;�^s5Z!�h�`c�C�r���	?�k�'��2u��,}���h�����������`����ы���F+y1O�ߩ������h7;�U{E�b6J+t�ө�l�D�3�*��K���U QF�>��+��Og���m"�:���e�	H�f�����]Zi���;����8>#����_c�<Z�_�L2A��'�����mQ*�Dʊ��T��|_a��^ZE�0:��P�m�we+r���z nm�G�J:	4�E8� c�px�'a�I�d���4����B����8���0�j��3�"DJ0�c����so�n ��{c �$M\�Ah{'�[�ıT�7��LCJZ3!?���e�(7�(��@��w��f��Zz�t�
��p%[`_V��;��<���U���͊Q�6�u*,����?f~M&,�"X~�Pm�E�p;� �f�t��$t��R�NM�,�q>�fJ�;x}��Z�C��ۆ컳A�����
 ����Ʊ�� ���y����P��젒�%ZV8�^�<�˄�>�^�mE����1��3�����Ae�1dL�h��*<�3U5(����] ��� ���H����/��v�������o�T��aHp�
*��t��
ŉ^������qZ����E����ѭ#�: �dDTjy�:�����L���n	L%�����O둮������b���t�%�2�1j�Z����?ȫ�ʻ�o���YcТ���o(�{��U��'H� ��^Ou�<7a�w�mS�K�zL蝺Û}�؅�Z�'(��>(���3++t�oXY�K���>����
��j��&.s 0�ڞ���@@�:��$����_g}z�ʞq��gɲdN,��#y�I��\HI��$gD�Z�NB:�M�cSc�6s���w�p��i߳]_���X)���8�+a�8�&�]������8GDዯ��y�bn�����]0Q�b�(dM�� 4�c�k �\�tHL��@̸� `��D+���	b�C	\c�C����,�C|	�D��M�ф
D�R�!��*M��W\j	�)F� ���e�R�,7��v��*��w׸��;΋?��<1�Kf�C0�-h
����2���|��l�z�բ��Ϙ�(����M��d!<׺H��7}� \��.6�#0�y�ͳ5��Ė���_�f�'�KI�%�7D���};y���9T�e�b�kSx�֭����*�$EWHG���tl��f�e-��������Q��aJ�1ޗ�8��3�ǀfg5�+�� ���w��NP6N������'1:����*�s;R5!fO�Α;ĝ�<��雲��~=�A9��a^��T��ks�Rb�m�������Ԓ�gN/�~�%a�S<���������s��3���&!Mn�wNb�>m��vw>;��Ӆ�Z��X6M9�/=_Ujt���4h_�����Ļ��"O�ڇ�l.@�����R��V*C�?(�7^|��K[�ҍX�bW�5�>�P3uǺ+�_<(H�>�v�{��b���o��H�f]���AU&��#��?��E�g��@m������:���6�����&�TF��깩��I�RS)��*�1{b���NK ��:��wX4��m!/HkX�*L8��^�� 45�����,���!�L���4_��.Ku�L����Ξ�#�AcI�W�H�1�r��9aA�x�D;�/��c}��c����S���Nƒ?��*���b<!�:f�(#\�/��#�N��-�16^���+Wy{c�d�����#�j���O	�W���զ�hR�1LNaYd,�ɝ(�) k��B�v�x�xI�UU<�5	��ćYҬm	�'	��B_�u�E�u�j���9^�ܭ@al?tFE�Ӗ1���S�q�G���O��;���@�J,�H���Q�?@H�7�h�1�6����Ś	�K�6gi)|�/�K�5�7(�^??� ��O�@핎e0���O8��W���uBc��f�V��ߨ��H�v��7��[��3����Hk�K���h��?��᛼c�	�����U���[���
V���:E��2�X���c"Q�y,g9�v��I{�U��[eEM����	ڄ�[A�_��o�7u� �|Z�����q��I����a�Cǿ1�Ǔ�?�d<`y>���~ =E�0����Q�AW�����(��R��3��zk@*��"t����Ƴ�Ɍ�(��T��c�¹q�7>�Q85�s��{x�ǲ{�֌Z?�`n��1��f��PW�î�`�l ����D�X�-Ax�7{Pjjp��tmL��h�eY������7-�0�'���]&(�#h�k�~�FDp1����a�&�QҲފ�i�x�=,m7���&@"�g��}ni�K�W*o�&n��E��i������o�@��N���U^O�Z���e]�BC»[o����`R���/�oR�k���i�% ?��[ ЫG`Z�>C[G�1�.��5�ț��*�I��CS���C0��?TQ����@��$&@:p'�h���v��@`���gmA*b�M	��R��g!�J(n`�l��;�%�$iw�`�o�cľ-�I�:�O!�z�Ss�c����X�@���A�H�P)և�gj�tֈ]� Р^4���bw5D��0$6T�<'��zs��^F"Q/e�@,M��'�k�c�܉�JD�]��Y㫫�	�{��®'��z&܂U��_���q��j����W��0-�Ƚ��o�9h�"9�9�,RĂ�۳LGU��iT��j�"����C�\�F�3:2@C��B���<�ʙm����x6��R���Z���UgX�e:�F�Xy���r��y�i`�S�y�-�ӳQ�u�w�Gb�KȔ�L ���	ZD6���Y���Kܵ�uAl#�_)ǚ.�Y����:z�0���Mx=F_lf��
���w����K}:ˑ�o�LRA����m���$.`ob{���j�w�	�6u��؆�O��6�7^�c���-��̳��[�}Yb��1��*��+�u�I7�Q]WT8)��7)��z�ɶ�o�F�����N���^�6̢���&9���y���/;�<U��wkʢf��r��^�w�C
[�a{���6��[nx�j!}S&�����u�T�E��xwF�yP[�Q�Z��y��qϠj�A�I�$&�Y�nь�C��C����c�\��#�+3cf�(|�&e�Cs:��G���I:8��pp���ʛ�����JHL�/�,��!��a�F�"����&����ũ�/vt(�ߣW����#4	��׎ƭ �f:yϓ����H;o�K�ƕʧ�^�	��M9�G>��Lܽ͢��������Y�0ި��\���]=!��ܥ����fF#dg��5A4�<�Dg�i�[~��ec��I9�q�6
`���Ol�A�Cؓ�� y��s�L����N�&�E� <�[Z�V<�~����5Y�����jA58m`���f؏����&���eG�I�Kf��G����Xg�n,�?-��&H8����S`B��0P�t����q} ��!3p1�)��uS�<ȵW��y�k��1 �:�P3�y��Nֿ�<������9�ޠO�\���K4|?K8��*{ܩ
}�LfL����E�A��&��P�[^ �=�XU�g^+��������A�HeT�-���^��X�I>�Xr<֥��$� �rf�N����ֲg?�`p�;OphsT2�VQy���߉a�B�y�*_C6����
"�t��λo�ͦnG!���YPgLrnq*6%Y�a��~�㣄G�(�ׁ��@�G��XA����B�\Uy>m|��GC�t/��`�p�pu}������������e7��ƭ�+0c]�j4�G����Q\*�2��M|tܨo��tJ���Gw���OZ���w���n*�?/<x:*�A+����+g"h����.�$* z͏9nBmr"iL_��G����-R߇f��0!��R��`e0S6���$�,��� ���α�.�A!�/�
�����Y��`�]R}?�fM���?���Ʀ��c^W�����;��sU��8w����o/�yf��H����I��U��uj3�GL�u3�.�:���T�*�㋮%]t���"eF�݅@�}��5���!��۰2�K���"����'�
<t�\L�ՔP�N��8�J}�N�`X�c����oE���7w̴'��9q��\`�_�������k�FRBU��i	l1��{�0���p{��"}&^J�..-��0?h���漥6KY����0��wWI�����/�h,=��NLpQ�ȅ��@ �[%j�-5��d���A'^�88yk4v9_���n�Y@�T�N��|�+�5[	��O�:Vh�fN��%l������R�9ލ5\-���'Į3����"�y݌GX����J;֚ܐ*����J�ori�_�0�ڽ-�.ο�JRIh��nWZ�\��$0��6f��9˹%i��v���{����D�Z�?P��y�����V���A����Fם#�T�x�Yk�tJ!���]i9�
�S,�&���]���m4"��8����rgm#z�"���M2዆�{�0IR-d	�=N�޸�W(2~{�� ���X�t�s���s��O!@���o�&�������c�+�b��O=�JƗ�6š�:��%��]ůP*;BQs�+�R�Μ��m/!�3-g�:q���.�N?E:�A%�sq#x (���
�t;�#��	�����Q!�TC�_�lZ��J�Rࠜ.��V�5O���t-���B��Kq9�y�ŋ��^�G<�Ӝr�_�֎
ҏk�4\�'�m�����F�;!)�T�'���G@�v�)_9�ҽNo��J�+�/ޘ����+���U���F��4�2�X���bS��e<�㯡�Z����P���e��s9��[�.���xW��]r��_r��½����g�}��ťR�8��-�F�����?�ȷ TC7�h <������汫�lb�7A�r��0L�����lʳ��-������_�=�cr�XƐ�p�e�ꚃ��D�/eR̖����ެ���S�l�~�1����QP��Q�r��p*"i���f��D��'�`R����Aʱ�OY���,��&��=�^
ǁ�q0�]<�ȥQO�i(�:���C��[��������V�����)�i��n]�t���@,&�(%P���<߁x���1�K�}����ѩ(b#Ԥ������댵ς��
����y,q0���9����a���(_�,E]"��Z��|��-3Ʀ�g��k3�����0�z'ZQ�P13a�y��3W���(-DB���|�����Y�YKճ��q��y5��J�U>|�J�ަ�BT�P��	@n����=m=Eic]�o�=.y�.��C���W��vrb�4T� (�q��� ���.�6:v� �5�4ؘ��6 ¢mD�0��T/Ca�(�*�����`���A)o?ϝ;�����2I��?/%�m��B;*���Z�3����`�ʲIN@��m����.²�9�w�ߦnq�[˱�)�o-���w�AƔ�f4����][� �b��c�Kq��|��)`8��~3��e��`�����۾`#�6��a9�\f8I1�����^�3���N�tF�T;Z�hƱ�!�.�_��1蓊�O8>��/U�����ӣ�<��2DD8Nm���F1(������h�r����z�:���^p:�������S�f���d�=�7G�HJ�[�Q��ٙ��T{O��ޯsW���A8ӡ�"	4�͟
E�g��d���&�EvC��lI����Y�6'I���u�?��!����=:�r���]
*[�Gپ(���\/�2T�����j���m.�l릧��q�����/Y��7)U�`��~b��|��Wp��dp+�K�<M��<����i�����ώvM�f���V�f�����h,�P��s౲ڒ�c��H�:I�a��Y�UEԥ}-(א�#�.�-��)����>ZlW�N�6����ӳ�d��/��E�4���u���h0�����E�K�t��^���E���$�I��dvl�H�CW�M7���R��-�h�?V'�]�{w>�@<�=7n���շ&�{	������Z��--�h��t�p��{��S�N�7�@��~��;���A9!������ �4�#�D���Y2o���ٚ�![i���G;����B���4P��l>���!Zw��WA&N�*���{@�,��A�0��o��gW��f��X������u��;6�Z������O@g%��b;����Gu��|��%���P(�E���ƭ��܎a�5�n���Zp��}������F�:���_n��� ��=��>Jr󨮎�#;p~����k�)�C,�&2 ���5ZP�q0�٨Q�;L�!Y�=+��]JX���$���laL���kBۆ�y\�:$�N��Q$�[�p�������$�	���曛��0��ї��#��Jc�3��׍w�]��U�k����iC^�e.�X��<�{���V�P��6OF�p-�N��gNVa��Ut�$}ѱ�B�/��X�eY�d��Xa��	E��&��m@{�����)���b�13��'�ũ�E��m��ە�������%���]����{��Ss}a�B`���R�)����^;2���H�#Al�1V]D��W&� ���z1alP�
�Ki��C���������kk�m Q-��8Xv��~-��7.7��qE�&��%VoO��e��ϕiE+f�g*ë�m ����$o`p#�	��l���;T�u�U�1��c4Fm��#R���Б�u<�V
@�mIe��"�e���a���\�[V#Y����� ��t�����C����fl�Y�$K���H�9(z.ё=�������{ke�wǹg$�yN�S���P��G�m�&@��=wE�ԹF�l�{�,��9�/��S�T@��؊�f�]��_Ѷ,�tbUF�abRf�(<	�g7��f�8��Ƴn�h�Bk�Z$~ۊP)�G�*Ȓ���t�W;��]����D�{L�eaQ}KH�rR���HL��+��Z�5F��M\+81]̲P4��ީYBiX����DS��{��c)��>��r%ū�$�í��j*O8�����2X��t(u#*��{�S���{�͔x�نd�Y�!�[�*�������Y����)M~�eQ:�\���eG�-a�,�É�h;qI�|稢*�T�{gOU����۔�5 k(b�������5j[9�oG�E3��S��R��8���D�pՐ�hs��~��<	I�h��m��I�2/aoc�MM��Et״I��$#��&���K�(gKT�B;�T�N�A[Z\œ���e3T�?h�}�"7����Ɯ���lp�r�������-�jt����b8����Iy%�&����f��-�.�J���%8�O�Q���\L�8M�����]7X<aݛ��vk�����]�N�ՙ�Lِu蓠�T2�9 Ǫb0�����9��	�*�^�����?%����]5�:.$�1�SR]�OaewhH��hHz�o��#�(�.�EaT�LLt��s��O��~��(��5�G40a��|b�{�.4�I[�`d^��,qnZ5+�a�>�eY��`������еD��F�؉�l�u.�)�ٵ�9��Q06F�JvYq���]��'0��6$I�x�� ~2T7M*U_#�Bx�x�?���͕4_���\ʕ��,��H�L�i��#�9�X�`�%�&�8�X@�D��|L��l&�`��a|�z�Z��I�����ѲC����Ÿ�٬��K���H���#�e�RH���6\�;�%)�,�5O5�`�H��J%���`,%�X7?b���5�Z��\��H8��wZu���\�3�)��oGy �;�3� r@�,��%��l�= ۾v����`b��I���E�&�^;�T�c���W�Di�U�|���T�C�މ`�k���?a�f�
m�E?��all�����mD� �(�W�cO�L��dЧ�.�t�d�Zt�DM�N(݅:�n��qa9ox�5��\*/K����ؤ�Fp6�o���V׳�R���_������<�]%��9cW#�p�-�Y���w}���Z�qvʘ���m���GP[qQl�1��t��@�PA��mD���#�'k�����<&�Γ�;/�le���`+�W�#��rᩯX�s��N�:.��˚��@U���#�W���m�}��ЬF���N�ͤ��3�C�	If���!����>�G��=t�7<�k�m���(�i�1E�-��n%\Q�[w=t��B{ǀ�OS����2sr[7Z)��Vi7
3�,��'�}�9c��~��1o���7��)!-l]�2�X��WJ7Px$h���PΡ1�L/Sʄ��Mˣ�3�L�7�|ďz�m���8���3[���g��TW~A�IzsH��#�z_�>�D�&襉�z������tD.�*���xW[1��Sy��p��+�	�m����)�r!
2��B�ř��+��:p��x>��EͰY��������A�&���[�Cui*�8^��[�o��Uq:�W<C�����ll����XAeB{Db�~.��h�XR�w�A�[Pa��ҽ��Y�&hM��NZ{z��ߟ\�p��Hl��(+~"! j|��X��l��P��8���Au'jr����ʈ:���6���lP$<g�H(z'$.���
����z�Z�t_�mg{��븪Ipq>�ͼ���v'L�������+au"}H.P�3Ԋ���)����w)Δ�u�?o�ۡ��k�J&�;Q
[����xx��x�'��zH\�F.@���s�#a� eW��P�t6��CU���.�����nU�r�jh�_'!y�Ý,-DC9P�Ȟ���Z===����B�,�d`Gv�<������7)���������.�N�`��ȃ�{�(���z� J��u��+0���f�����g`i�.p��[�V;3ª�*��u<�0��x�|ϱ7'	��%���/e��ǨLac}�\�ɮ��L%���ϭ�&���&�3WV#�T-��zz=jR�8Nح`'�X�h,yjl���SnGRh��[>]�>�`�g�-t�0 |d����af�┗�[3�7;^��;��K��iJ���g$��1�e������Py���=a(7���,������!kt�/�=�1Yaq��L�`H�@G�tO�2�0������Vx�`�c��75�^`��Q�(����Cq�9u��~	���:>�tn�7�J���HT�7Q�����Qxd����?MC������]t�:�UYS�o4&+�n��C��������̖���� ���ߵT��hUڠɲ#=̞��r�n�5��Wf�����!yb�2F������C�0T�kY��%F�g��!�d�۟����01��K��~v��?��38x/NbטP�ϩ��)	XB�C��Bw��ڶ%-�yuo���#il@Y��g�O�[���{�[@R��xؠQG�ψwX�ݤƕV6M��x���|<�h���m�<�9.,)��#i���p���Ʃog��]B?��-��(LOa�_��޵�����eأf�y���6�EZ��x�h��
H�������VL�- ��G#�lα�:�ĤR�t��X�RIK& ��V�����	�s�$A�B@�55�JZ�t^��i+6�A56T�Y��������P�r�[�'��*�zgk�Vup��!�b�,���1ց��9�qD5���Ӈ.lCi5�9����1M@vYõ���Q�G��iˁIy��/?�׶ �c���-�uֶKF�@$ �0�Q�9�L�/̟f�F+��;�`.;!��7��=�(�-	q4�+@O�7[�s��Bx��Z�鱚��x�H�8����N�eDz���~t�����
�K�P�Xaۆ-�.�/�C��Σ@Z���2��(�T|^g��Het���?�d��)#�E�08;����,_GPz!*ʹ��/�.^���z�8����Bs�l�� M��c.:,F8���(է�/�/Ȁ�x
M�AL�۪x���gW�^T��0��2}C#tF���S?|��f?x�4�Cvҫ�ό^+O�yڊ�l�F�\����U?�?�\���ۧAʜ�!��g	��
��!z6]``%%[@ݶ�;͗��j:����*nfg��ß3������/(�������
n���%��p#ZR��ľ�x��I�)��N "1��vl�8G�'' ���J �������˚����ZN�ؘ��R�O�孄]'̛��[�R���֩�e�L��F"���w�&�^d�78�_W������;,���'�P�֘�A��Ⱥ013��W�(�쏬Ҿ*7ݩ���ca�V�� ����Iz6��1Y_7"�6Ġ�(�{f��*����e�{���(p����ͫ����G2�B*Y@�nU�(1WoqR�#�?��t�p��y�N������~~���=ta�������{����iŉ����u�jÕh��/CBd���h������?��]򇉥����r	��n7vn��Y�pQ�Y%��"��醈'턍v�/�l����~��cؠ�2��R��9�7]����}���T�_�`U�]�"K��l�5k+LT>�#b�g�4C͍A�@ϖ���\њ��u������J����N{���C�`�yX�J3GRT6ɍu��F�KU�i��l���=�9n`37�[��ДB�{�0LfC�f��R<2]���R����Fp�v�0>�����;G՛a�.ȓ�a�g��ֳ2@��ڞR)E��ߞ���9��j���F��1�rc^�T�GC��,��/�t;a���L�C��^���I�#������8Q�ʬ�����Ji��[����������K��FF޹}�#1������ �dFh#��"'Dܞ���hVmIT����C�>bKL�{%��\�vN�1�<���\�	T;�<z�}�/�ʮ1} Gy�%3}D���|�X��C��6-�!i!��3��Z�9���kB�Q�.��1�j n�Ѵ�=^xD���/�X�$&_fM7w����"t����{�*mo�l�q\�;�z�P��*�qSz��Y'���l8	^ʍ��*&�����r%4�c9�|�h)گ�4�����e|6}T<�^<lj�T�d6�"�7b���-�p����N�aﳳp_��k��2hU����N)�
�_�i�ɜ�*�ɳ0
5Gڑ]��r���H�1��i�3�s�~ý�bOR��!��	OT��e`[kN�����ASx"t`
I��ET�w}�ˌ[{#�"�BXt�֑�VΏ@&�'m�3OB�P�3���?�r�7��W���g�,�Ʉn@xLWc�G\]@7jڝ��]58G�W�βQ�"��(c�A:��	��̷��5oUҏ��	.N�N	֪�����׿vA�Y"���	��L�R��Ȑ����3.�;hfjtǠt����k��6CzY�̆#�꩜>-�)�~M"�J掻���c�玙��Q=XI (�;
ArtCj҉�|���c�pd�w
�����n6�aβUe�h�D�f�)"�ct�GU���Y�p�l�25lP�(ِ�p܃�c+��i�|~�;#�_Z�JB:V:����S+Jm��ݦ}�R����F�`���b�ղH�Eu�_C� E0W���x���}<�YٌA�Kߏ�%�k�B����2��\)u�L�)ڟ�F�@�
��;���v���ўN��T�Ԛ�w������O��oE�Q\%f�2T�T�?0����טi�.�՚�K3�'R�̡��q�n�շ،��?|Jf�4'y�潫$�X+�+?􃐺�/`y��7
��;g��������@؄U��9����/e_�)<0���-.�cJ<LP1����K�#BN����r?{[f'�̴�o�0E~��^������&0f?ҩ6RCm��a���6��j�{@��*+�BiIe�j-���8��j�Ă)͂��DE'؄�CL�[W�a��6�?%p��6���]�������e>��tN�6�FrA��<�={���4Yϓ��A�`����!F���+���AE��.h��;�]�a������h��XA�R��}BC�'B¡�72�Mb����z��@Ct��W���}�u��u��Ga�:e6󛞠9s+�n*IӇ�0�qT�R.�b�����8r��Ȱ��6���X�1P�H�e-L��|�<����u�t��v+_
={2i�C�ׇ��a5z�܇?m�|���8^Pr,�lW?��5+A���㟬yu�c�nY��䥂�ÿ�^��L[@e�jy�n�� )n�rU�ء�z�6��lר8(>�߲��Q~�Mj����ĳH���Jq�����{�}���a�8h�l�y�{�Tt� _*�Pf���A���#�' �l�DFF��[���Zɭm̅��P2P���@�K�)Rr�<���1�y���L�{�w�&���?2'�c��B�v͌��Q�^�V^�����Ȝ��� Q�3C��W���d��pp�}64�]�Ґ���P/�]�=���J�g=��q׾�ci��nl"���Mj�j��H���NLJ�SY�s���Ơ��iP�U:���nkx���ΒB�6���2�x��� �ɀjT_��-�<�RF����k��+F�X��7�Z-%�Z�6��[r8?Ƒ�>��[���[��ӯ���mJ��y\�z��;�brT}��awg����ߛJ��ڶ؈#��副q	��#ebW��[�^9��u�#�v��w.I�@d�����,�J�iP��g��jm(�m���/�����?l#]�UÔ�#S�:�]%p��"�v�OZ����7^IaId�^d�ђ���9,����N��cx�y��g�F<H1kG������N��sF�p����/@�����w��N��#����Z���W������� O.O[�l�����w�����1��,f�^Kx���)]u1����_����r�d���x��R��I���Bu�m"��J��`6m��9�8G.W\ղ!�g�}��vY�1;��'���=�,iN�7a)N��A.{'V�c%����9�Qߥ!�m�#C�C���r'.$�2kj�׋%�po�m�rP��,��Oڜ��n"~��9��^���w�S�U5<n�?�T�Ǧ]C�0�9;i��E�(	�!2��G2��lU\�C�_Դ}'����h	xj4�;H{N6k�7�"n�u����qꂼ�Z�m��#�b�0�?lb�8[��i�l3y�m��W�U�D�O�H��/�� �d�u@o]l�W@q~�!��ħ��f�qVu.:�_�E5�15���,V�B&d��%+K斶?����%�~UR	��{���s޲���G^����K�`1��|������ ����'�@H���Ʊ!8���vu�琨 �)Ր�3C�+�61t�+3�]�c3�;c���5�N69@�U��佼��F�6����LOi�=UQF�{m6�-��E��eh�O0�SY"f�aܯO��%k�O�;�8ӡʯl��q��,7p.�[�C��Ƀ���MH��������<h�����/�cñ��i�`Gf�j�u�hhIT�xv�Nj��F���	�`Z>G�OxxX ��J:,�Eҍ�!P����o�%����;A�� N3���/6w������&@�U5��HtO�dl�iN�P�g���u��N#��1�#Xx���;`S���L5�K�C�ۂ��ý\q�h<��B,tW�Ĉ���*���֭�.L��*����
p��k__����8�����7Mu��l����_��u|s��cN�>\��c����ҋ�nG$�{�zMj��x���p�D��s�r,5�	����}"z�U��j�\�y�Vg`�����fM��	0�cXt1PҔf�)�}��(C7c�We��n\�;v��{gדƝ*�F�Gf��tH����� B� <�m�7���W^`Q�A��n�"����wx"	�@�`s��)��,������t�dzS�ߊ{7?S�:2�U~&pv���txh&�2��UoPݬ���x6�^S)-�^Ԥ��=&�+�	@�G���f�Tn)/�4�dDQ����<��$/��}eNU<D�q�b�-���>c�V��o,�~�t��~h��MP��^�'����|8�Pea��9��|,����	x��ԏsw �U����CCsR�X�+�	 �9��+5P�����g�SS!	�ُ�M\.l�w�����L�*8{�Q ���r��*f��;q�.i4����O�p������_�qR�lin�ϼЌT{Ti�&��Z-��-M���j_D�I�N�`�d�y��9��L1��rޮ&����$�Ǡ��8�L�Ll�>�V���,���0�yVOI�B9���@!w&�W���{^��<g}�L")XiE
�J�T�pϏy0e�/���V���d�o\�XU�L��ӧ2�fvYi�#k%�y�y��gռE�f�̱�@=xx��1g����߄���I����� *Ph���=�~�R���J�)��ǿ�䵗k��[xo4)0�EфAz�=�]ޏ.Fm��M���^ޗ�����ݭ�.��^��2r�hֳT����|m�a�G����Y�L�ƽ���B̩�hs"��Ac�n|�>�M!)�_I�� v �_�$�6��"���b	/`���}(T\���j�E�H-�bB�PJ�_jP�<��نO�d�G���c揹�k�b[�2�I�.r�#ğ�i·�̈́�]7� �^'�Z������~z�n=��H����V�߈� ���6�D�-[���R�1Yr��Ui��@���Y�H>�/{������b��e:��g=��˹���`���.����*0c�s��%p ��H:fI�������m���ܽ��psc{z�1iyX��lߚM���Ȥ^c���~C�*m{r<@B��zo�*3y5/���7`+��#�ӄG�xf*ժr9��U�����\��Gk@��4f�@g;�2���nʟB��!�F���-r�(��2�q�6S�����&�ua8ǰ�,L� WIR=F��,߀�.��+�	D�}IM��&�Յx()٫��r���g0�)(;
�J)�V��C��;��΅ �W���(��V8Tu��z(�M���
BzQsR<�X�_�\�A�9��M[n�:!��`��4�d;��'���ׅe� ��ݶ�L�P-�  ��r�Y�x� ˗���DzG�vIN�d��p`��n�o��E�[�лD2Q�Vx���.�W:׃��@�3��3�wn�<7���s wF4�<��LbLT��L���OZ#�Z<[Z�h�=Б���|�B���^ȩO�Y� � ���B]Pk��w
_��� ==��d�Z_B����I��p̖��~�{O���r3�X�~��q�N9�z����H&6/�g?�|�ɉ��TOV�Ks����8#'�v0���_���m_���GO�b�J�
JRg)�xzV�+���kQ��V�3�-߶̽z����c{K/�f~��N����΢�[�Q���J��Պ=����0q�kr�y�>�d�����~��Y�<B�!9��ل�.�Y�'�ޔJӴ����~.�}g��3"��[Pic�Я�Q/.x/ƫ2�Q���	޸�C�����s�����2=�K�0�"�^��[:������o�ֽh"T��rY����ނ��x�gH���)���W8����`Z�\��*��U�� �dE�9�S�>���gPO�>N�$�] P���fju%��qb������N��^]�q"=P��LU�C�K�ҧM`��s�PW-���k����������p�G^e����rT�b���:��f�ћuD z�T��A��͞��BK�.+��&�K��]���3����n ����>�.z�o�l��?����3����k/*�1�ꡒ���~������[a%���ฺ)c�Vo��7K@m���A|���+?US5�@�����ǐܚ��mF��yV���:�8��0�j��j S����*��l��s�@�Q���H�b�p��{H�|&r�Xw�b
�f_�f�K�]�lC)�0�x}p��0�I���2���@3�jxo�t�C%��{2���[G;|�)�'b��4�.����
�4P^/K&�������K���s8�6^��/�d6�%�b?�y�� �GD�cy@!�S�U~+bC�k��v�b����g���}/�vI�y��v�o����%@g/���������7��v�Qm����?��c�˔�0��~v�5��H��	i?�/�ն�}�BF�$F��k��t¥�t%5u9�逡�٭����#3��V��%!M��p*���!ɬ�_y�Pi�������Gz9@I,���11b�XOQB;OM�jKPۦ��kٯ�RG�r��F��Z~To��Q{.gΝI�:cQ����.J�#n���p'-��'�Т���>�?��T�9T<��%͹J�%�wt���F�}mٻ����XESA@P����4c귙Q^"6�A�oV��ԕ��6-u 6��6<9�7��E�U˳�a�=��K&!˿a?�^6qi�1\3�s�Sӫҗ��?:;LP�����/Xq\��ۼ�K��p���ݹ����m�u7N83�bmD�O��oB�K�GWƜ����p�U3�g�Ҥ~_�.Z*О�P����t� O�'��k�©F���S|M�����Y�A0ʬ_B)��03iie�� حyߒ񗘸���گ��F�	Y�rb�x��0��TH$�"}k��z]���P�R��	%"���b�� ��B�+�.A�%'��Rp��ȟ%s`S"�
�[��& x�d���KA�l�г�@JR�̥�R����׌p���	�W���K�H�][`�y�dϮ��X_�:�w�l�`��?hD�@  ��X�~�]���ӌ�xh�w*����5d���D��u�V�;���/,!���gh�4������x<���>�U��2䶆�q 6�C��W���Z�5q�
R�z�2q���R�%�aO���h�Eu��%��z:���*���=m��u�#�=��LA�%	��Z.%��a}G�U���
��퉃�?��x�<�d��n;��jj!��Bw%(cn��C�����\�@jX�b�=Aa������*$��7M��y��3&ԍTa�y~|�o��E�v�t(P������#��W��'��DDm��X�阡�V<�����9HyQ��@I�n��-�e{zZ�-h��[�WÅ݀�-$���n\3����Lk�fl�X���?��}ٞF$w�<X�O_J�?�a6+�GTC3��|Jb^��ObMq6W�qC��~q�i�����G�_�<fM蕨��)"_�����<Oy�Ε��_N������ħ_ɾT	�d�J؃���2ITDE�/��?�yN����OKw�� �is�,�F��D�MN�0cy�(^iX�@*wRu�)���k��?���MI��,� ��Ķ�����AN�7�  �B�opz��Λ�89C�^�D?�xA;4n�Z�00op�g�y��0���++Ͳ煝,��7w*��RV�W�E `�P��Jdbz%���^S2��L�2
Q��H��O�ם��P�ټ�NE���ٌ;ř1,����H���ŷ��/�l�P��z?=<&�9����9��8�^��ե#����ėW��DC���QUV�Շ��l�=랐���̕9}4жB��}������M�#��{bn�au�X�Ԓ������`������(�D��U��ן��Ӭ�bfB�D�W�f`��ȳ�E�Wr&8� �(�B��:\iՇ:��~��Co:�d0��0ǘ�]h9;�4FQ\�
����ɸP�u�G�O��}
�?w��c<�15��$�xc�]௫���ֺ�}�����[��}�!ڌ1�~��L8��%l��]�į����y��BF�	>����&T�$gQq{ʥ8�ʾ|�	`�������7p�Ky�?̉�v��_�+y��%�"��u��� ;��X17a�������RePߖ�i�e�l��}C�Cb��9��be長Ŋ]B�T��ޑ��Ţ\p-�0�#�Ʈ�g��4k�a��
,p0s���-]E�z�U+�v袍���R�a�C?�n��D�q�^s�)�G���8�9��<�����
j&kw?�_]Hby�b�=O��Â1��������̈́v���{[�c	�xނ��r���F<Ǵ�k����0L��1!��..(C?e�~�!|)�U�#�M�	�a:\ �Nxsܤ}l`�)���$%��ӄ^����-��@��؊P���;���RR�{7ry�@x1R�ig������K8?�M���f�!�g��B�ڍ���}[^�~�+�D��D�]�{!;���c���J�C�oMW]��!L_��lZF��y�l���m� ݺ�Rջ>�a�����Z��Z,����k���b?Q4Yj�E�jp@>�43��hk�$��%��ap���p��0s]���M	rXuC���r����
3~�����:����zm���ވ��wo���3E�G��Q�6&�b=�^ ��T~d�)�d��G�
�LX�[���o>�ѐ�a�Xv�7T�����&X�����~�q���������0(��7t�`�tӥ�6ĺ4 "{ݰ�Ş��>  ]���M��#L�1�:!��uEg�̤5�zM�	�v�=�Yh��n�h+�H�FRs�2��p[�6&.���P�(���L\CZR�h�;l�9���-�t��8���T����&I�L�݊$ �U��ж'�_X@^V;�c����BWqk�NO�&�1�ꃦj���5V9��V=�Ǉe�i�m�}�J���k�ȭiA�����}P��g�4�� \e�y�KR�0�E�!f����:�ykI���PcrN*��JT��pl��7�	H��|�(���Y�Jw��qBJރ�9��
�4���/U�2�"k|:��S<�e4_G��wyȗ�7'wԊo�xpA<Y\�����݃�[��{�c��.5h^���n�^�0rTM��Q.�����0�R�����	>�J���a�l�� �+χ�y���hr �WH� ��%S1>��E�p�Nnh�*�y3�Kbɺ�ԧ�5]e��M�!�~1)>en�<m�lY�؏/�~d8=����������;y��Ϸ���<�Y��U�!==l1��CN� Ū�c�4��#"�qDWʃ��z7zP��H�6tI	(68��!{U�G,gx�
_5�-�h����T���C��!�E���BZ:G��Z_�}���!q'�T��@�_PH�aK䇖��Z�8ʼ�v5�W<!r�rE@��B���׿���!e�rΗ|�ȍçV���t˽No��2�	�mLx�M����1��h�eˁd 4os����M�&���$��r��i�ɳ��\P"z�<��1nU�wf��dX�:���r^�j��L8A�ʛ������9�XhS�b8j|��&R�.���c�v��̷H�j��遂5:�@�6�S�s���w�Q�z�O$N�� ��-t���*��"Z��G�h�?�����}��u��0��s��]+!�Fi���݋�uER)5(`}2�O�Xo��䋛�������T���@]/�˲�@��(�!î��v�"�QI�4őz��b����r�T<
��ĳ�-n>��Y�Oc�W�ɠ!��	�`���Bh�~����/Wҵ�a(,��Nk&�kJ�ߎ�"u ��ȣr��T�KV�2�:~�8-�7l�����cOQ���C�A�Lr�l9�cT��mC�s������Z6���yF���cUƅKl�#Řw�	�Q��(v�|O��U=�Ňcx�~olU��͹.��^�;챬���}�>�+4F�-�m�{U��g]'~�ֿ9}lX�E?c�k�?�~<_�C������������YǓ�4��/ǒ��ۥ�'�+�D	�ɤ ���A�!y�` #!��7CI�M�~4f$�{��������2M���έ^);.J�����P��DR���ɷ�F}s�Q����Ee���W��}3�����N��C��������m�e����^���I�֏T�' �ͮjc�$b���K�^>y�Q[|�����ӣ�ܲ�"g&g��V��Ѡa|>�� ���2H��S���"�Q�U�'!~	8�QyB&n]k��Sf��_�A�{��@����5��s�,-���Zn�������'�D;�
�R��L& �;.���G�1�ӊL��k�խ쇘�D�aq��V<S����.<��6�^�)U��Cݩ3*Ǌ�X7cV�".�ؐ�@L����z�^�.�N '���l��F��wuTg���9F��x��rc��4�~��ܰ�<�DG�_@�U�@�"��- B��ǉ~�e���f	,}h>z&�>~�%��]��6�e�	d�l�?��@�}�D��ܮ��\��R��ϴ�Ωp����HM��R�"/�L��"|޳#)~����^e�e6���r"z�
�Iѫ{����$�:��n�{j��'5�C�ߵ�����}ې��}Ng����s��Y�Ti��sKu�B��y�D>��Q���(�2���N����Q��&~P��b#���-����=
Wװ�d�(<ZW��TZ�˸�C�&c�)�9��o�Q/4Wy)-�C�n����	�+z�����'��!\��CWJY	S(��}<�9#��R|�^#�L)l��Գ�_����8�N�hf�5��7o`�QO�|1f��<M�h��>���"�y�d���
;��)�����Kl���ie����!�`�L�t��5��_��\M�c&���Z��� ��{V
|�}~(����t��9����.�qݔ�x��w�8��2:�ذ6� 9w��ܱ�:�%ʭS�yW�a�ր�H{��H�8]к�c)���f�����������k�-E�#�D������<Sy��)�n��k�~�|A!KF�WR�+q��q�5?͝x׉P�b͝1z����_�w���[w�&��"�WO�y�,r^	(nް������Z�^5�1�c��.��l,��m�,x�] ����6�tH�
Cː���!l���qZ>���Ӈcc$���u�סPv�B5�ˌ���;�Y<�a��E&���t�X���L��`u]�� ��	,zj%�ItJ������<�hb���4�J��q�J����B�G/2��/^�切����	ũ0�`�ʵ�!����l��L]K��0�\���E�Iو�,`������6^^����t˺HO��U��D�XB1K�LIh7�bg��S�<�R��zx�hD�a��&:x�̋��sKr(�o�`�A$}�(&��,́o��Ӡ��(�v��A'k��4f_�?\�a��+���,�S����bBն�ų��湢o���J����+��_�V_�_�؅����������g����萰SC��A� ��-_���,@#�U�P{����Qm�+_d�w����	�Q���VߞN���V�� p���$�o�%������Q�׏�1].���*ەR���H��<�hb��SL���@�g���m��S0�X?L�n��oJ�(��c(^��B��m��j�Ӈ���`BZ{���B�����>v��Χ۴�qw�W)��t`$YQ�!7���\�7��
�p������@D#W�,�7�Mt�X6��a>Ob(bJ0��	��Սn�# JS�y����]��L�~�Y���*l�����h��Ä��8�趃_ݖbu���ل���{}ƚU �ϸ��?5�uY��=�C�s	�T[A���W��_:���Q�wԈƝ�,�Z7�U������m�,��.�B��C5R�{GSN��L}�&�S		��b�?����E�R�{ӻ����vϩ�|p�PN�p����2=����<�c!� �61Ki�I]�G��1�(Р[��3ۅI�'MXD��Q�̭�lD��3������w�R���Wx�t�{�B*�&=���(.���(ݝ��;��w��V<�3i��� KT��e�r���FE	��X5D�ٿ:e�O���w�w�|^(����zRX#9�OK"������S~d�*(�q�s�K�x]J�����<D�Һ�A�^��ks����	��z@���Y��w*��Ç�Q��9�/�ΊS9!^`�}�0l��uL���#Ї��
)�k,Wˏ��� ��R�O��Mͷ�K"z26G��w,o���ńpF+pZl0l�(�Ry���
p��W��/���u�Y���P�ꃀ��ie�_�sv�.�9��u�SҪ閊��׼  j��ܠ�2)���琚�G�UӸ}����Tj�?�3`�
/�W �	�*�X�{m����{wH�%(X�<l+�b���fƝ|�ɗ(��iBU;��ȷ�[&�X?D��bX��u���̺��]���F�x�Vϰ���]ظ0N�-�qR��Y���&?�C�p"?���+�F�s�gu�w�Rj� ��q�����R�B�sa�^�E'����p2����*������%����u�LG�g��1oZ}��2<0�"r/��G���t�ih�.O3-C�L0�+o!5�d|�5!��"��c0��&bR/���u�l�I2�4a�n��D�[�X0,͜��$�����3��~uBEye��c��6��D�{�c�^��^�Kw�ϻ�U���	��%s�!���H�\v@�\$����q�|�!iߨxd�oj��Z�(-)w����F0y�~�Irvi��!�m8/ᓾ3����T'1��<����A�c8����R��hې�O/	A���$�݄|x��{�3Ԕ GѤ�E���;p�X+�6��i!��?
 l�P?�;PO�{	�4�a���#Rr���G���qF�b��
���J���9��׺`���}YcS��������#�Ӊ!1�61�]\-IdE1"�[�(��hX�v�^3��j�l75T�gc�"���������0
��+C���6�>]���u�E���n#��;|���Ar"q��C�z~����3�ya�h��\1�������jW8��/9HgL�;�)#H��v��ue�B�׼�u���ȗ�&�@�X�7aA���T��7�JĻ3"7�B�?i��	i\6�[@��Ȃ[Q!��9�ރ��_�$: H{��� y��C|v�S��)�R�$`b�������k�d2�C�9��P��Y{p���&�y��Hf>bAn�C2��M��7P�����p�3ߒ~�|^��)�΁б��ݥ�]G�nf�f��އ�V��R�n:��őv���׀[r�c�%�[#�Z1�����[Rp�)�Hb8�����������
 ����qg�SYk��Ѯ�Q���R*J�~�z���6���vI�A�N
HIf�}Ɔ�1�bʹ��㳹f���r�Hn9q�f�&c`� ��S��Rp#�4wQ�w���s춧ǽ�(���M�\��׻J`XQ�<�(��s2g_����f;�Z��π�~h�Qa~�b������
�<N]ĥ�FXe�K�Z6Bñ)u��pϿ,��ǌ��Z���7S���l3�������c&,��4���4�|	�����t���.�C� �yU���e؂�e	;gx�F�v�6��0#��-���}�)n�'�tt�X�Wa�<��
�c7�`��l��puֵ�D��\���}�$�3�8u-�Z|3���|�YQ๣Mtf��{�M����iTS��;��)t鋤7�?�^������(86*t�p+�����1��)�h��k�^ԕj�EoW�-��l"s�	��gc��,�ݻ�srHzD~ui���t~}�%^W�C�t*�i��1؀>1M�B��O��ms��ٮ��\ �8�	]ȗ�3�����U�~�d
��V�.�Z=�y{��6M"��z��K��x���E����?�0�n%]�22���hVr�_�|3�;*�7"�q�7ih�I?ӆȮ#hvz�v���r������v�w�?�Y1�m�#��!i1�/��<=x�s���s��6ǹ�n��}ܬx����TuG�b�?�9��{s������?y���/SGK���5��g��aC*駘~O	*�R���黧��n�Q�g`	lmR�{:��zi9�����ǉhNjfӥbO)�#���H�
�~�΋�͘�A���t(�x2�ɴ�ue�8�bYiK�	�X
�� �����
�'��+�����K)=u�ӏe7�}�cc.gA~��`_hN,.��cw<�:N��'J�Íԯ��OL��ї��d�5�o����)��Ջ��<8��5힤6����~Ot}�S�"{M+��V�YaE���^MZ C8�vKF�	�A�e�^�� X?06K7b�|��G ι��!iY��C�cRO�<z�z%�Z9����T�Ɇg��f[{l+��X�2^d�ӫ4J�[g�{i��C����}�Eb���k�R�'v�!���B?f���DN�����Q�،�S�<��7R(����3�'�q�M5tk�TQ"Z-xUq����V/��K�n���tA��_���p�`�][�2/�Ԭ&Rz~)O�tK�ψ%|��#�ѵ�k�:��
y��e��C�t�_��`������x�PA�hA?�\���g|;d�r�\�7����,�aT�OB�ʷE�aKN�����:M�q��V�o�āf���a6����VD�զ2�YT�C� ��� 
�kl.Ņ!��F�~�$\7[�����*��~����A������{���q�7s��%͒פm��-�EN������Y��x #��e4YOc���Ί��X��']�F�"�	���QL��V����(�\3��Pº�����b���۞�v8�W{r��&S*v-'֘Z��7F�ZR�w�=ZBqH�}ʒ|'0��b \���7���B*)^�u��%
��X�I�8�;Hί�5gb�۪h{��ݝX�a'I��C��s�S�*�!s7G�!�ȿ�)��	��`�򚬥i�s3�J*]D�z�6_���M�dڨ)�`�� �7��u!��x��y�j��tݖR��s�C@��`#��xd�Y)ŀg��z~bU�"��}K "���8�_��o�-�1�O½֎5H��} [c�} y.k�f5�V�v/�A%���r�T#;gF�n|?UIx�>���]H��X3�v5�a��4��x�2_�2��fe/�t�IZ_�M�)I��Y!�w!*��%Uz�_9��W�j��1��������	�!-5~��Q_I�"�oM��ģ�N����Uܦi:m?���ѯ���Atܧ:�t�k(�K�V�dIn��9�*Zn.冒)����ޡo��D��r?MHV 4������&;�N��
>W??E���'v����7�j����▪�E"��P2�t$�����"����ݾ��RQ�~f���m zN� ����������V=F�f]n.�w�I��R�h0ģ�>2 ��� �nV��8�F�i�1/�G�ۿҿ�_�y~��s�(�׀��d]���C�_I2�/�Es�-BLyc�}7`��25�ˮ��xFeN��V-��B��Ì��P�>��H��Ww�9{/&&(H^v���d�'0֗�1Ie7G�bF�����p���4󇶅��P}��T�n���a㯒��]Np�@�2��FJ�O=U���T؛)Pp��勋n���|6�U���2ߌ���L+�֏x���rX�x5����$UՓ�ڮM�uU.�X+��4�Sֱ�'�,D���4�k��c���O��m<*8��?۹��d��#sx��(9��$@fFJC}�t3yݾ�<�Q��/�ny�S}��\�?�2 Jm���i�"��k�J�E���N�_<�ct�%���=U2r������.�ے�3�~y$K��� g�8�lN4nw���R��)z꽏�!��G�u���q��3����0bt�K�C�|/�B�_M��fD,I��}O����pÌ��)���x��7��w��Ȑ�*��n�{D�"�,�7�M��P�d#u:��ag��׀r��&s�[�2;gws���`/���
��WI��c2�t\��'B�h�B&���.Og�"��{J��v�'J�0F�T����MbR:�qd�����x�W�2A��/s^=�ڼ��P����<�6�X�2��I�w�ɀ�S'C<����o&�R�:��wsh^b�Gz��~Z��}�x�}�}(�g���I��y�G����\XӪ�(���8����o��<y����'�bI7��L��0��N ���,�>��M,�w���[A���)lmη2K�<!p�.���'ҘT@y�*#Du�64�n��92��{�:=�)ץ��eq�����?���71�3~O�M��|s��[�Ch7�_�2.���)j�I!wF��@@ppK�w V����i������c"� -�\2#�1�;a�������b+��Mz�lzyx�R�0�l�D����sb�[e�c��bּ��g���Z�d�'#'�.N�|w�3	��JJK���Ii�ƛ뼡���7�e����|�'��O�� ��q�W�*�~fmtg��$��Z�2/�����ҁ��IcN���jϖ$j��>�V*�?�'rNs6�X������Ć�-��Wc]=9�Zܢ�@5*���R7�ÖY���/���.�J��*5$�'�h��+�;�2
_I�C�r`�l�Rl���`D�G�_5��d*�b̮�ql��5�#�S�WW^�JD��m���s��#� ��u�+�*��_��F�!����N�����T�
wwX�ϡ��y5GC-yv���/L�k���Κt��Be�~(��y�!�°��|ܐ�% �]�6��TG��}\ȑ. ү�ڄuptŮXQ�SK���s A<K��eu��a�T+�.�@��-w[���ǃ\O���g�ʪ谓��>Cp�Ql�����y�2t�5���*Ki&�-�ot%��n����	("�@+P/�騛zȒk�e�/�d
4�&?[i %'��hO��4�JG7����g�e��6J� N�0�2���d_E�$|��8�2���=�O
�f7�e؁�g�T�����Y�1D�L$w*�
rP撜"��P49V�gAkB�u8��FU",{6��:�g���y�K����d=y�څ4�X�MzD<g���6jp�|����W�%��~��H�d��U���/{� z����I�ǼE���'��Q�	`pG�H0LX�,�5H�}NPi�Wj�pԄ�[�qoX��-�Qa�tYT0��]�Zu��b����#j�K7�z|};_�טf<�,R[v�����1��!w60~�z=(j�=�d@bA�84�����MI�kأ=ȏw�������ׂ����a5D#�rٻN����W�Y���Ĭu���@C�5Yӑ�H�u�yt���AHY:�K�?�}C�Np
_N]��s�	|��Blֻ�&�L[e�ƐI�|�j2�	�Y��c-R|]��oFGX���t������&���h�bnvp1��5Ğ�hRc��v�+��a�^�h�!�|�pz��ƪR5���+�YGȘ`���5��H���6V�,��+���'��Va䘣]�<�b04�`vZ����!q��U������Yo0�+��&;DRU��0hG�n��I$?���S*18����Z�M�(m�ɑ�I�������U�soz�qVHU;�q,t��X�H�9C�D�G
?
vQ�T����V���X�[xs	ϗ!I�e�FrK�X;Rp!U���Oߟ��,��-pB����������t��ɣ��.�o��Xi�I�Hrf{M�y潦.{����1pd�+��J�4#_)��3x���H�p�fE F�鮾vZix&H���g1YPBU�u0q�#��ʌ V �-P]9(� 
�j�x�^��nOM0]^"W|u⇀O���G�9��N��s�Օ�OΨv�.������Έ7�*O���zZ3D\+ F�Sc�F�,���_���9o�j��CqK�{jб&����Ǜ�KΌw|d[��|��%[|�h��s���J�0u��8�FV⹳�uw��S�q�:7i��²��P�EHU��i���)b����	_U0��f�H��#K�`� !�d�<C�3#�Ni���$�ְ`�t5�-a�Y
�.� �[j_G�a�)��qS�Oy�v{������
��/%�	-$��` ��� ��e�1��6v��J�%l�߇,���L%۬s=X��b�O��h��������gvXT����_�0�p6�a�(G�]���={_�T����S� �9͜-n!@xE.#����X;@<ET>�Z����Љ�F��6����	g���[!�-��
�;r� 'F�=�`%���?3;��I�s�G�&3�;h��	��8����7{ԕ(���Q�K�!���g5���:6�D�Q�Ɩ�Zb,JX��i�����_^�R��3@\g
/��Oj�y1�!q�% �d���O�z|������$��/-oMƇ�u�s��ۅ���o�z��5�S\�1�x2ϣ�с���oa-�]_.�e��d9V��GK
�k4-�@	��Ŕ�	�#<����b:%S,zMk摬���L<Pl(fr��p�~j�v#Q=��v�=�l�@�f ��,�\���G|Zxevai���kgq��'N?"��8��Zx�w�/�ו6�e���f�����������ו��`��&�lA*>Q�c@�9�#"D�I�e�&��_�cZ�F���3��E�u��:��ʌ��3�l����x�w.T��@U�z
���``�^�XȺ!pPH��8�fW[,~�l��!t�%m�g���S,o�����t��ŘP�ػv��F�2�Ņ%��a�\��x�o�3j��U�-��Zr�w�
��p�ϯ�a3��/k���A��	�^�u쇮���� 8�n������qf��g���#KS��G9�A �ε����4����[u���e�]ce�ͨ�����p���	,�:%߀YZ"d�W2���'/���+TI
y��P�g�1�jv�)ƌ�14�����w��uD&'�h�p��1S8G����c�Fls��c���~i�-�v��'ԭ���q۸��sD����B�"��ńcH���O��s���d���O���6��(ݍ�$ge%��D�!G��=������w�c��1��	�ĕၟ1+�7
W=N����;�ʲ�� ��:c�Ќ�p~�7��h�Ȫ����!l�F������׈�_jB�-z2�� �{�oXm�2@7p٠�*-��{��ͷ濮�������լ(Hϲ8�E�	GA����CYE7y�����������b�'�BҰ����m�������L��$zc�c���/(6�	ں��c��w}���Z1����Vڱ\��iO�c�S���$ӻ����Otԥ&-2���D����w���3�MBa_�Ң+���%j&�JL_��L8�ηP`��)�|�"�}�t6)�V}Z�92g$�{���U���_�[M��+��Ԯ/�;��	�P]��Izc�֍:�M:k%������a�r�;4���ך�z��[Ч�6d-��VT�\��XO5�C�b�G+5%�Ĉ���}��x�K�?�BB�s	�hVg䭲�SB@��`�4),��):�};f�3d�N�n�<E�?�-w���i�p�y��=��O�R|��ISGr.���r���G�u&6 ����s?]��f�����Ut*�xuU�M�
n�TA
|d��7j�������0��@��Ȯ�#snn��q�-�k����Q٘�SLV�]Z�&�\}�Ǒ0�Ŵ�H\���&:��'\��'��	ZR���O7e���g|@�5a+���,4%�2Y�	x9�}V?���ur�������3�zm��d�E1�E{��?�������g�s~��(^I��_���vГ��΅�la�0ǟ���D��pa��R��H�\�G�)~V"�2���|�=��\��[�s�i�dat�>XB�c6���t�a��.\�@�_./�f!�9�cK��T��gϕ�&�$��Zm,��N3̇]�+e;F�%[Dd��M�sq�����z$�=����R=U�_8Ҟl��!ˬ��)	�r��e_�vh1�x�Z���֌�?�D5�4�AŤ�9�P&�9������F��\8h�4�.^A���5���X=$@nU�����6��Ҷ�u��/:T������]%|���Yf�m�J�H,�H�Tt��B}���Q^%y�"�g:��;��C�($�U��n.��a���=k^^V�HC�6��1�5� �.�����(�^�H�u�1�ǰ�o!������v�τ��=�>t���� ���X�s�*�f�	���e�L���f{��o_?
�d��8O>:f�Ï�0�ňO?���$'�������gM+�Y0�4)�#PL|��9g,V
�t�hz�t1�Q�RO5}hN�����4��H�p$NB[Z��>����y� $�Q[��Dǣ�9�ʪZ�C�D���	\;�������|,b��a0��Xɣ4���:�e�{Ĩ�Qӹğ+թ��M��^d�v-�6���5@S�/eሧ�@W�o<&��nc�_��de.��Ns���I��8ac�A|�z�����{���S��X��I���̬�ռZ�����ZW��Ps3/�
^0����oq�I͢�#��/�W²w]'�BG��hs.�a	�	�����'�m��_�i�B��i.o�h���j�
A���u��jڝ��͡�p�Uz�g�LW�Z�<|��m'��@��r�E�Ž5���"(i��n=��g�1����j���5w�����G�O�]dd�-�kg�s0T1��B��]��B^*�m����k�L�W��8����
Ss#�l{kX;��
�n!��^�D���!9ӆZ`VO�*�tީ��uy>���S(�H�&���R�F�7�ӄ�|g�{L1OK���0��o��nb��fc��bC��N]k�BV(DO<=��lAS�^�+!j����GI#\�ѫZ�z���>x�%[��ߥ���K,��W�$#��@��:_���,�%c�+i�0hu[O��jΑ�_��=�t�'���r�>�m��T��I�M&�K����*���-�:~��cØ�D��i�����	��i�K{<�f�υ���ǥ�3A�W�<�Ԍ?�wD�����,��-������(�M�3V�-��F��Bs�>�u����z%^���?�����t��b�c��+2W�y�r�1�?����L��gE��_����T�l(Z�[��]��S����*`�rf=�
O�q�FL�_M��DU��� �q;F�8b����t��bq����^���cvZ���.4�x$0w�4�0ߓ�A��Q�e�G��Kx�KcΎ}|��a�0����n�MEYdx������tTΚ�"�}��j��s�R�ԍ�n���&;x�-�?+��Zf�8��ϳ��mQ�l���t}��-+�1��J;��3#�V�)o<��N[�(ɖp�/�����_��9�aI4]S`^"O�1 ��rq8�)?��$��S�V@5�j5�����ȉ�:�!jfI'�� G��)B����^����l�o"0f��|H���d�L�Q���/���w4��9����hMh?3�8��p��TP�..4��X���9[֘�j@�!5��U�#�T�L��O���~�wL	�? ;��#�\��as��	�XE�T�C)�10��4'�����W���f��|Nڴϣ�=�dK�zQaq1i_�2�P��B��8��s�����Z�AF8뙯>p�y�t��O,�؜c�*����C(qx�D�Y����~��*Y� ��ՅX�{p9�r7���p��,~ `4����0��v5���w4dZ�Q��1���iU�1"��WŎ&)�+�iF�1���x�"�5��v��<#�m;;j�5���3�+����0���XG�y��w���u��q~�㟫�:ǃ�c�������K���W�^� z	u�.�u"4Q��@G��Z&r[�6�l����l��x^�������^qH-��t't`k �pA�җ�R�*��:q�R����a�%
P�$I^���Ų;=�ifd<����C?ܵ�Ţ;&6��2���J�KOn#���j�b�ߞ�+��iཊ�P���F빀}����ڜ���=��M����#xw��l;8��8�Z�#zRw�AEZ�1��7m��=��X��=�1=� ���N�U��)��TA����Lk��<���U��ܶxv�f:e�ޤ�g�mx ��m����ۈ1����I�ֹ�0O�$�'��}��wɓ��� ��̡J<ɥ�?��zT���Y���Y��o]v6�
|��۱�.ت H޼A[X}^kz��t�\N6�L��o����A�&T��*E�!���W�#9'E����68�D�����1�s����8oW(� I�7`����ɶLP���F�ޜ���ڷ�'N���l}0>
��(R4��H�H������b��X��-s��I��	�>��#�a��[��%�s)����$�k@[p4�����K��0
�E-��֚���/�m��-�d�.�����7�<j[�1��خ���|ZQ�jK�k<�	ܣ��!�p�Fd�i�������F'Fe(�1W�N�����|�tgÖ2Ym�rB�z���4�F�n6�A���1��x/׾r��DG ] �	J�p7肓�N]E�J���.+po��3��Fg�1��B,�4ɓl�B1/l�������4�����.W�;�� �*:8���||���r}(�:�p�U�\�3+54�:��������D���?�r.<)��T5�GzvR�Mc.�����!U��*;���d�H4�r�� �h�L�@�E#<)Ke���º-�}���<�&u��ر/<�,�l1�e�/�f�X�O�=���M����G����ϔ�������w�$��7��q�݈���S�ת_˛n�4�_n<_)�>������Q9������
K��!ޟk=�U�aC�ɨ��.�`B��^'�Z�]�l�AHB]O��|? �ү���t����������v��\���ҢԶF�'�l�F����"ؔ.di��/l��4K�%��7J~�Ǹ1�l�w4�f� 5���`u���?#`�=�;1n�u��q0_(Q_���(�{w��cW��.6?�����4B��&�������{�3�lyEM���u��?�{ ���t=�2��CC�*E�'X����X%L����X^J�[�˱��0<�e�����1���-י���\� �P�`>}}����i�X!�������!�Ƴ틫��ىR�(wOC�@��M~"���`��Ɠ�I/&l	&E �!� J��y�wS�ޖ�8��ZY�]�=GlKb6k���'���i"֗Ņg�[~����K�(c'JQ��Z��9Hk^c��	���~�;Q"w����4C�B�Abo������b���U�\�v�+�p�z^�66���hݞD��V��e �m5B��d�nQ����o3� �`'���n5�Ԙ;�^FQ9.�"L%p�c�»K��0�6i"1k2��,O�<�1
fIw.-�_�cs�KN^}���g�j���bч����bU��7~�49��51���� !\l`���He��M`Ď�\k����+uD�?�7�e�/��(�&���P�9I����a��6�nT�C�"xJ����=q������a�����E����s������1��m;�,~� �����n&�k9�$T��`ꨮe�آ*����;��i����l���0��5�2��n�}�O�3 w)`V�L�L ��=�Z/�+��o|�n��LL��Dpa1�0uS�J�qD19 �����vx�-�|b�\ʧ��3�v�O��c��R�{��m'-/�7,?���n�ԛ�c 2ｋY���)�B�� I�E�$W�;�.HI{��7C�r�`>���W��������-�yF�䆺i���4}�?Lڅ��?�B)̚�Ojm�=��b���(C}�8{�gq���������������˹��B�����Q��y��]�J�#�A��%�H,��8�ȡ���R>�Z�o��(&3a���s�=���9#������Ϳ�E�> 
�hmK��#bxV������8� ��?�y��Ε���ERut�&�(˓�n��F�����a���^��i-@s�97���P?ayk�^ Z	[�.����w�	��:�p� <0VK�=�no� ;x�M]�"��jxZ��n��;KAr��PT���M��i��].��wI�v��ph���Xr40y�_˦'N�H�z*d8���E�m�C�>~�G��@�	�c����@�
@2WQ�����-n���r��;�;��]R�i[��'d#�J쨲7��.�c;c���ֶt�0��#Sl����4��7 	k,!������L4D��i1Z��٘:I����4v����gÓu�@p ��M����x�㘡C�Ѓܠ2��q �p�L2�3K���U�3<"`������%�*��،ђ[����3�c������5����!������V�~P���?*�~�ù��M��8Zz�N�u8R.ރ�k�u~k�Aǭ�R6�����[<�9j	�����^��=����*�fe��Wq����NM�r��L�s��=\8��T�j��A�K}w�1,Kq��ّ������R��wy�t�f�Kv�(#z�h$�����D�	�@g_����z�q�2e�L�:�o�
��N#`i9[/T������[�s(��j�Z�F�Z]9��g��l�oۀ�q��̏��٦�S�2�#a��ζ2ʲ(�W�/��ϫדlg�K���od�%P���'�&Ӎԛ�n�oH���J�TmjYG��~:Cq�|8�FⅤ��ܯE��.���� ��I��B�Wk*��E���mp���|�E/q�j�҄�oE�W��'�~~� �P�K�um���|��iZ�K��P1��S3�s��BE���U����7���3BǬdS�D��'��u��cGN�f���x�j��FY"�ů�Ց���Y���7"��Ka5����bJ�'�&�J��\���YF ��"q�0`#t��X�u�#�S��w��ٱ��w�Qhb����;[�n/�̯Y� ���7�%��1nD`�� �Y������Z��Kϋu��!
�:�e�+�wsMs��#����Ad�	�D�4��J�Îwz���6\�d�[YJ�Һk̮����ߓ.�vf�y4�_�i��_�!ХI��K0�6V����T+��UĿ�<G�� \*�{JF=�t�L��;�SX0�I��Ž9���2�3f�d�}����Nv�Ր#��t:/��OK��O�7fڙgg�0��x1�i��(�C�n������Ĝ�x��S3�x���f�|�Ϧ��<-M�b{Cy,�+Dp��U�\�z�O�t� -���D��0�\�
s"~��!��E�B:+ۂ`���-GF阅gK��ݦY��TQ3�0��5W�o�D�[��V�I�������a��
}�r�\�ÐfOw�ߝ�>t�_�p�=ݠ�H�jI9
,'S�h�R��0~��`���ޢ�[�b`�&lۉ�~c�W�r�-֮��f�Z��d���+�����D���D"��\�ċ��#�I.����2���	�+ŏ�b���(��3��Z��PL@�e\�H��+�6�PH�qJE���A��a����ð���$^�*E���y��X�϶id�
j2����0Q��	o/�tT����]��Օ-Nh���a~K_�i���CC4�4eU�b,u�i�@RCAۣ�z���{�4C�"�!��ȧ{��u�������$��)cAlGU���P��A�$�"��2�Ƅ�l��c��ŷ�h���q�Va�T���KF����>�i��g9��`y����.�66'^]e!��*�y���f�����A�W��.�F��+���|�]5Cq0{��+ �[]`��%���6��^p�1��49�a���$���'�ݳc���T,�'��#w�˾0�ӥ�ﭘ�顕F�����(�a�|��B�N6�����WV�jRE.�PvM�!S�G�a��|���h�m��'�E����O|���	���0�h��D\o���Tj�e��5�CJO�ݣ�o'�-A��1$$��_�H�������u���L ��y�4��V��L��wdW{	!�(�"-��0S��$p��F9q���	�
?���f���I?��XY�A�1z����-U�s~�<7w-q$�Z�KΖ׫'��\�0�C��O|��4���ܭ��w!��-iW�+2	�Y�z��8;B�#��<� qpF��?ڃ�g�������C����&��Ё�"
p)��^Y+����,�:6]:�N�qj/k�o�A�t���%�C��S;�R��6V����_��Kbdo�:`C:�u��aS��dt��4n�/6'��a%�4ЦE^�007�\'8h�9���ٲf�7.t)7�c�v��˧k�̮&WgFJ��c{���\�J�������w�CU��M���:[*|�e�ნ)C��|cf��P=� ��EWSi?t���E�@fF��
C�X5�$+ W8,.}bN��F>n����i=d���jW��P�PCL>h\��~\P4�D�dx�IT�Tx: EyсW3n�l�� ��[�N���T	܅OQ�������2�͈�>������ˡ'C����H$���L?Y����(S��8(��+ 9�!�)�|�k�S�����)U0u�r����x�Z�����L&⟡��i����ОmU��Sl�~�9�sZ����?��8�]��?��Y�h�̣���Xk�2���U���ђ��Z�bJ(���r��	j�'!8�K�����o&��9���L�%��` ��KHD��	F9���V>�p� ����`l���c|���A����g���Qü6>&��&6�F5�.Z��B�(���٧O��{�}.Z|�5�pK��C���6���y0�\��k�6�U�8,���?����c~��Ak�� !�~���w���;H�<�ˡ~i'%+eq��E�$Rt;��y&�\�[H�7f��0M��S�$3<��?��e?'�yT�Z�k�%��}{jh�#~�dU�;�^U��	V�w�g=��m�@�z����!�\oGD݇/1�NB�i���xh_�M&~z0]���(q���|C�cU�ڴ6�/�!�K��޸�Z8�`V��{�#0�C�	��sX��;8���ŷ���f���N�
��f��@��ύ@�呗�"6m���2��+d���vv�=A�<q J"�u�7@��G�O��Q"bU)A�<�ٰ�F���g��n2C�{\���6jlcMy:k�C�_��J�Ϙ��2*^��وN��Tt:�3{�.hs�VȯF)��=?Eϋ^���L>3Ļr������uT��g���'������ �n(�ӟH�̏"$�P2]�Lb]0�b'dLߨ���b�]�K���U��7��x�h4TTi�"^���C�aܝ��`(�ĝM�	b�\~�be?�ruu�c�֣��0�<w=�A'�yƛ7\�vT� �jƶ7�aڤ�n� ��,�����.��]�u�
z�X敖����̍"ݸ�рz ��*V�(	��q���c�9c8�V�~mh��^iN��Rm?E����DB��&�H�%bRQ��{��.	~�KZ�ۅ�+!ĸ?����֠��7�-��6�>k�w�x�,GX�t�G�mN��)�P\�(��~S%ɗ��	o*�nܜt�㏬�ϝwA	|+Z'|$�����P�-��L$��X�j��+ܕp+����@w��t ������������7��& ��酬W��#�*�S4&�l�m�h����7-O�	�&@/m,]BM�F�Z�osRӞ�hP���q�O!}�f8P����=�����Ͽn�����F�n�1���>h)�d�-���_�"ZO�C
Ib�
���f�J�������h�l| ���P��[�f�zF�S�H���{��`��Ce���Q��W��^�����̑�
S�[����ĎC�k�+��"�I�>�(���RD�YX�|Bi+�y�ƥ�դFn�;�p�������X����9���;Ō R�t�$��?`i�D�S~]�C�Ω3��s�}��&[��������v������C������3�,���;u_Ў�x�7ͣA6��F.H�V:R`RVɔ�r1�Oȩ�2<�wm�?���A�m��*����᷊>r`�G�?`8Il�l�.Dʓ��Q�	f�t�F��붿���ݚ(�W���ݬE��zx�0����OiO���%~��s�^R�5�s�..�T\�N�!y@��t����e�+>Y�%ڇ���c���MP	��nj$�1��v}�$�����k;�6Td[sM�
��������vz|��g>f�u&�ؖoq���6�B}�9�k>�Ѭ�v��E��2(�V�m݇��2���*��Vyz��1y�Q�[l7ѫV�����1��+ө�P�d̘�*μae�h�r����H�9{m+�a�9���S���e��I?�L��E�آ�	R��٦�.Oۯ>�d� �l�i>�[��\�tE3��ǽ�o��z/*���*`��\U��I7?���Y����mH3bq�o�Y�b\g��#�8�,㌑��q�ϫv��_�3Pt����l���a�흽�Ƹ/�hޠ;93�QW�J�KB��v��y��l�������$I3茙�u�Z�o@�Wt��&Jn~����Q	����І��� $b��")� ��tn�K��;�TYI�~�Q�lZ�z!t�����h|���:���F���d�'�A�� �(˛�J��@Xv�xZT�z�W��%��о�-��)��nB�uY����gWэ�)��2G�l>6����ۼ��t�������Q�_s�+��iY.�#��cW����w��g��%wĠ�n���-�;Z7�~�>�@���Y��J����׶�����Һ��� ݆������I>�����E�X�i!]���O�yU��Iy�����9ȩ��0F^��
<�*zr��*��ݿ,a!������ڦ�	g5���̗O�/X�-���*��zT2
�ye���_�T��~�eZ�����9pZ��X�Ú�^�f�hhak�7I'g�D��: bGn��	#h�w'L/-���0UF����*��A�m��uf8y��uȈ��YL
�9D���W*�a\%�g��RI� I;	?�cW�.����`�(�2��=�F`P\��@�} F���=_�-(jT�,؏�DO�;0qI�IM���N�Ň\���h�?��������x�\?`g>]�>���]�g�D{�d��̆��(� ���$��Z�D�jx���0hD�$-k�wL��-)A�Ԅ�mDDݱ�wK�ّR%��r[��I��uq:�5l#�!=���	5�~kIK�TU���{\6�\B�j֏qg"�sa\�/$'�U�����a�@(�d�j���4��>��{�q��%O�_��w��gL�ς�Mt����dA���sF�9��5��G5��O�<��9���O��zR�v�^1e(��{<��+�z�f����~�#X���B���#���i�K��<�]=�P�S��!:�P��<��ګ0 �F�)��T�x�:��S���?휊E����I?ˌ_���_��j�����Q��Y�nr�>.A�Q79�K7-�+��	X����hnD�f�*O�l�gp�P��Y��ĩ[z߮�ߺ����i���:;	C$�$Wl��]��"Mhь�6��-�	�\;x��������<���%v��2��ߴ��nf�X�e�1�:�FpЌ��W��βV�)e�]#2ܷ�5����ƴ-�D.��?]��D�{UXK�?������b������|o�u<U�zM�#��U�S���	S��*�&F���B��uO�@��Z�Ux���ܺ��yY���Ǜ#�"�^��>U�]�)�\+0ަ�O����,�ơ��Φ�l��7��ؚ�k����z4�����WZ�@�Nh�M���1
굆7ѵo�+Ӳ>>�WV.OQ���0L쨛�"vq:xS���9"�?��b ��������@ڃ�c0Vk�jZ��^�C�^3�����������ɞYuP���z�D��nD2N�:��	!�B"G�����J�W�:/����B�h?z���(�D��DoL7�5�|	4�rK��Qk�(���2�Y�?��ΊbxvB��Ε]2�i�8]$�(�8ERJ^�r���K�D��*�5.�4`�Z�zQ��%�Z�n� 9�ab����W���j����#��np�[MfxV�����R����N��X��XuN�ѝ���*g,r[�ɬ�>�^r �p�#9�cP����Q�AE�dt��;��/ڀ�:O�I?��Z�|��C��Mr��H�~YS��
�^�Ѝ�9����o�~'�X�yy�\�k��Y�Ɏ<sq�!o��īZ�P�C7�%d*d� r|	}L��X��O�>CvS�-AqQ~��s_h�($4���u�*ʺ����ݶP�䠁�o��-�.]ЭOH? |���.�e�J`B��$)�b(�e4��7O.7\A~��sF�n\��A����r?�;�?c[Fӹ	=��ʲPz��q��Ԍ�T�/q��wQ��$�]}�U���WP��K�[q�k��+�	�<�� �`�%��E�&�5͆����7����ę��J��m3��k �rhf&�K]�"�D�n��Q��?�2��������{�蘚^�fT^�	��4V<b�y����CW�
�#����V^��E�C��w?�2&33!�Z��I��f kl��K �jg���z�	-�C�M�=����?�Gf� 9�{e��C�$8�[�m�~�I�4�O�x�# ,E�Z�b��4���
��UO��\8����"���6�Xxcl��)ǄU+K�
��o5��a,6���҄v���^��%��(ރ�	E��7*-����?�\��L��K=j��,��De[�>l��!��R���|����.w��^�!D�a�v܈6�:R��2mN�ʤ�fO����r���d.YF{���؉6� $_�+����π���fg/�5�s�����1����M큱B�?�A%>c�ȣ6�WS�g;�J�4���y�	���H�EHK��X�}��w#ҺV~%�r��|���]���PJ<$-��4�j�9>�w`b�����������A_���G]�^�/{�a��s�f~@�u$�P�S���+�񋭓9�ItU�F��*��lz--�Y�V��U���Yv<�}�bVȋ�a��'$��G)�zך�l> �]����YL�t��V��1�Ez�0G#�t��>Y�N�pͱ<�}��>�o]���r��WR��v���`��r�6���LS�_�^('L��,2���ш��$��/s<�C1)P��O�%�BZ�~z	�����������M��sn<�Ǣx��'X��X��r�/3�*Pg�����
繡�?�(�Ut 	���k�HsATܘ���3�r6FQ���؂Ǯ��v1�mA�[f�qA�Y�"d쏂�*j��6����)
�W���i���ڞ����в�N�&ZJ�a���=_�͔*F�j!�!j)'��T�|;lpl�B�C����A^����I���Z_��-2|#ͷ�G�A��3���e*��}��Y
��P��N���">�a2�z%m���͐��F؆LAs6%"b����|`�S���c�/�Z�J���z�������#��w=�; �6 wk7��_�>��RAgq��,qq����`�Qа'��0,Y�9��睮7���l�>~&,��&9��xz�N�����6�3�l�;(u@w�� 1��3��4W�d/|7, �a���E�S7�@RO���X��uw����v�g��ݭ(�����TT}θ.Ր����<�u��^Nr�F��ò�������:`Y��zaB\c'齣[k���P=��SK�^"�!��d��a�	�fޞ�z��0fx%CR��	#-m�a�B�Á][d�XVXr�{�Q��uj>j����:ɴ�ɩ�+Sro�F���&jf���t*Qjh�� 4F��`�����ӏ�˘�/C@��B
C%�!:���2s@���9��]��{��էoq1�Ca1+�����f�N�g��Tê������O�D<�������ǃ��_�n۸���5	;�fp8�(�/��1��A�&��4�Bl�
m�nM���o�g�ԟ��h�-T-T��oZGT�Ҿ�~K1	�
��j@�V�,���qׁ�q��d��uNP�_�M�Y������0	u3F�:��:���!���x��k�A����A8�����e�͒=��E��JX�M��ސ�
�8�.����QB��"����{g,�#�̘�>��.a����Y�/|��r[�_���(C�R��ƛ�V���F�PQ��-M��.�����U��:|c��òp�Ϥx�K�P[zC7�4AD�����MW9��6~hh�q".Me���j�C-�{s(K��|�������J�Ol ��`�8}��6k�D5����(����L
ܕR9���>���}5��.ky EDX�90>����k�ߙ%\�9Q���u�+�UCYq���-���q>���|�n7L8����\^�h��)}oQx�9_i<Z��G�̞&9��]�N�Gg��������=k�jJ�x��U0dO[�3AAňl{I�f{���x�B��k>-+7�gk�<������2��t&Ӈ
	�^y�U@?E/�q��/e�����fK���="A�v�6#��N3���>�� �+�wW�P�&��ν�m찷���J��z���
2�٦�����=};��Y.���N3y꧌)D+!�i숞�]�G�N5�m�շ���L?oe�w��B�r��S����f=z�F���뜡�I���z��-�<�H`�S������)CI#/ :�Y^�[�iO�(Tbk̛�E:�SZ �ȬΈy�:�7�9Y8����Q�>��ڔ91�n�Ø-);\�p�P���Jq?T�����ƈ��R���Q�s؜C�&�7p� ��zKE�Ӊz0�ǇOrX!�{_kC���]�;b���9Lܠ�d,�^~�vG�8��.ح����3c$N.� ��;�'��h��|˳t�me�k��,���O��I1�KJ�<z<���E?�hK�䃈��W?׿v4Vק2�s$�Z�(G/���\/��ΤF����۵4�luJ���_����'θ��ߚa�e�g�p���Ok�//+T���8'���C&��n���~;��=n�:=�Um�5"�fm� ��G�A�&�p�E�"�
X1�-`�?�KP���d��l�":1@K��	I-}�`�E���g2�,VF{����p۫h��PTi��#��Ǒ��G���}z�9�rO�5o]�ʌ�ϛ�Q .����ˤ3fD��
�9��ʢM�$��'��J�k#��
J��+>@`b�zr�Q�dӋ�
��IW��*�`���YB�Y��_Cˊ)"��kI�`O=�>;3��无v֓�3P���u]�A��V���uBe�Z'w���C��h���E&qK�%u!<0ڬS5�A����t�慭���m���!EUjD#O��UTϪ����aؚn���g\�"�O'��z���r"�s;,�^y���l�����~�~����'O���F`��v�)�י�����_��Ǥ��Ӂ#�/�$�-�+<m6�0��Qym7��;�J���2/�'�N�vU+5�  ����b�۱9z ��N��9zSޏg-
#�i��j�?�OE�1�eW�{�����F��p��S�h)�t�J4�7�,V���&E�=bp�JT��+
䨒@��;�xW���XP���OQ�"�TPY�����W(1�g�dnܯbXzB?�o�ڿPSq���m��o-?���`����ٛ��#�ֵ��g�%�������'8�^� ��3��y���,�n� �<�X-z�t�y�O��e��ژ� t�����C��hߴ y0*��*q ��6�)�[��u
��S]����:���h&M�����㊋1:���o�x)�o0�562�8�[x� ��v�"�A�%����c�3�F�n�.�2s�����ي�ľ�G��)��>9��� rm$�F����>�I�M��h���dఎC��ǆa�0�{����V��G�A�?㑵�Yj-*"r� KF���AyV3^%K�h�W#�ˉi4��t�R����C��W�<�!�Di%����W�Ut\J������o��l�d~����&	���d��Mq:��7�]��[d
�ԛ�{���C�H�<ST\�͆7��)�O&�06+�~�=�������-J65Ωa�g��Qpp�;B�2��t!0R�BdPV��x���x�`�n���e��{�pK='�T������o�pbo���^HM�i��ԴD�j��'N��v%��2��m�p(���G�?��UOY�S�TW97%�E�Ļz�H�31*��e�����2p-�M���Ί���E�#%o�Ŷ����W����5Q4�9ԛ� ߞ6s)q�����H�:�c�����@s�}�4Ś����r?{~�T��n�99��$��d5��!;�[�JFɧ��"������ж�SG�#��X����n��v�����k��lL�i����M��}3U�M�«V��
{U�H)<��:_�[��;�qo��KԷ�֛nT�,ml�I��M�G��?�oAl_�l��س�ؾ�;'��Ek��a���	��Ы�/�\�&'�����������@r��cڻ�r��]�RzNeF{�k���Wy�&����.+�(�`)�H��2.PU��D������F=ZM����⒞�f�IF#J�d��E�hY�[)�c� ����������ȵ�x��;�:�0|�n���,ؤ_ꭈ8�w���?QX �ʄk���M�	��n�6W��`�	�ͣ�8�Z�����
�$xw��Yp_�!�E���ߤ��]K�؂���8���.�x!����¡������VKy��U�"���UF0}5��#�}�!�
l���~�	`u��h�\V��M�j���_�]��n��Aa {�w<Rd)��r{ � ��o=v9��$��H|�rV�SD�[�h|����ԃc��"w[��
��H��'@��|��Um�C.@8sym�7G��w��`aFY<�1E;Zj�R|�3�^V�ڽ���`I�]�أ�e��PJ�L܌<}N���bs�
$���m8�FA�ʑ���@����r�U�rcz,�t�$�Ľ"@cX>��I���"Z��ƴ���h����j���6y��H�j��;{��I�����r�`:�6�5�3%.@�^���#H%\�"�)��G�8���Q�m,3ڜ�˘d 9�~%X߻<k[�4�g.e�xǓTojS~~]��:H�H<���˟V��C�2�a�d��B��� �����흢�Iڥ&K�i��rz�o8L��Ϳ�>,=܉ґsKD�XV ����-����S��%�������P�lՠ�5'�`�B�ȇ�D��i��ݝ��s�-�@�c�<���V��q��#& �rٞ�䌹��8�'=���x%a�2� �3�Nq�҃��}��!��@.��Q8B��w�q�v�K�GeM�i�|\o�D�ߛu��h�-�D����R��)<N�;�}堝�o�m�p^t���C�}~5��h�4�s� ��"CK�]�w`,.�}���A<I��Ǚ�>����P�P���y�����^ϼ徊D{��s����H�{E"�D5���Ïy��x�.ӌ�_R���K&q8I�T�F�9I8&�{��� hą.V�ɬG^I2VƎ����8�@@�`�(�t��~���W:a�nQ���p{<����lrP2���l��E}\���\}ՙuvԭ�1ڪ�2z ���8:��C�or���M�h�6v�|�#���]�a�b�Z7�t�띅�����܋����/_�Z���E�KKJ�kl�ۜ�ڈ��av�m�撢��C�ٝ��;����+��ѥ &Q I��=�*��G��_z�;���r<�#خ�c��`Uzʙ������z����'�_,�y5ʛǬ�Ԁ�0�V�h�7R4�Hr������ʫL�= �?�q�݅�g����=�/�+�*
���(�C��BIE*u���_�]/>�i�A9��2�qq��IDf*�o������#���e�+e\��bJ��D�p�$�����C�@�����|֋�8Q������ɪ���Q���K�.��|�
�\H@�ݑWҜ;X�-Xt���^�j/�^Nȥ��R^s|�PN}@��k��>��ʎߏ�$��l�3�F�/�9�K��`4>����,�<�S���a��]D̲�.�[tk�;��ay�e�b�5���#�����P8��3��қ+�1f�H���Q]�ķ �+x��+�R ��5���V�*�M�P�W:ӡ�68>��-��Ɍ�	�%'���ێ�WV������qD?'��3&���*>�с�^���Q*:���H�ve퇅E~�w�&i�ڹh�ܟ�Xf�����q����(F��>�6��kw��.�p=9���-_~���f@o�1��Y��-@/��'�~����9�Ǜ�/l�=,��BEW.x p�X>����U�ï��Wȋ�9���P6z��'@N2aJӚ <�W[�x ��i����oi1龲�8��H���{7W��hw�4Km�2�H�1/"C<[��"�c�Ec�����g���d*%8�;�M��1g����B֕�?8�]�@�)�}kC�k���W��x}@�[;�~&�b���γ�;>�=Y���_r:�c�$����3������d�I�s���x��f��2Jj9��à��;%�F��ӝ��ݓys�����B�}�],��7�{�;���Q  8ss%���zr�)'0�9��A`mҤ�&�����p���l��ޘ9t"�0v�
�ܺ������8�o6���{�DPq%��ׇ��*�a Ss�;*[�����n	��Y��v�L���6U	1`�J �L��;!������ܛ�x�y�a�U���$X��'R�uhos�R8��2^77��q����E���uJ�Y��ԓ4�a}E B��_���V����P�tȣ�9t�R(�1A�!�s���썸�A,yU8#Њ�S���B���QX`gґ� g���AR��HT����L=���8`�-�_��*�LR�ǅ�{y8ɓg�>�������AJ8�����AAn�~�ؐ�OP>.�S�Ci:*����J:�~�'��Cv�ۅk�H��3��e�Q�q�������2��^����cBTF>PVXXbk��"�h����CS�8��]���;��/��$)�������	���E�������38��������R�x��e	D�gYG"�>��A������!�2q�
אmx�8
2QAu!{y �Cg��.�?XQ�W�����zsLT��i���(C00�a�[[�8}��v���J ��Ӣ^���WY������,���5d/饳�ɻW(���h��%F��`E�#>�
�	���l�9SX�m����`� ��qY�xB�`��e�|x�6����R���5�ߐ�˘���!��[ͪFN�p�utqh��"�����=(��
��u�g�KIFO�L�Y�UD+7�1���0�Q�ǫ��g)�枫!xX�w�n\2���-|�^Ê"��_�8�yq��a���APh��&��+�j&]��K��l�2;ɦ����)��O�/��3/x:��S�Q�P�?Y����/i�kG.ܦ.�a��S'V�����d�s$
�O	&��i�����b�}Q��L��!��GɃ�tD.%,�=n!C���к��N����8���SBV�[U���z�#W��<-+N��vo�R9C
�C4sk���N�Z�|�OP����x�����^y8��+���ȳb��1��}8��=�HUh,ݒ��D�ųr��O���ꉵ5�]�b-������ 3OJ/2��!��]�Oв86aw�*Us�&�j6��b�!����Ƅr�B�����Zc���,�<!���+��a�'�=��v�ƈЌ��R�[z_�\b������'F]�kjS���Ҍ��zOY������~-eF��y�����B���m��dM�Ю�g�h�l��ۃJ-��pF�}DgK~��;0�[2�c� ���yڧ�h�7�g���ȷ4;p֞�ct
�P�e�C7�����g�BK)�#E����V�9]]ۿ����|����&a�8�?K0���(�
3RK��
B�Y �x�p`�ىQ��=�U��7J�X����
WSu���+��'�g��-�~��$2����H�R�=n��z$�)Fyu*+S�����G�	��c"Џ�[I	\j+J��D��ʦ��~�]5]�X�
���1]��Y�{֠���҈�sq=��X	�'���\!�hW*iI�s��e�ӻ�P��z^������!�*Ƭ#e���
=�P��I�L��d&W�!�!d�Fj�|���M�&2�E�ɻ�WD�o� ���Mmjo ���t����T��%c������'Y�ʢO>� CJ�ؚ�uUC�F��7�d�\�G��u�2��M�+�C �I���NPE�_�!��U��y3-,�r܉�k@��o�N�t��?bR�
�^�ݠ��|<�s��+�
�jk�Φ<�~&\����ã�g@�9?#�|}�&��wU\�lh��9�nW�R�n:���yV1l�q�%�[��������0O�+�)\�7,	��{�S��L=���6�C�j��Ӣp�۶��Uri�o��7��	��L��iw��WP|��~�ѷ���q�^��)�{Ѩ)K�pe=k{��(# :}n#=%�G"@wZ#P�&r���b���A�ok7�g|�n<��*���-�pb��F.Q��]=�s�-����q�J�	�#�v�O�VpB~� �ͯ�h�i� E������^[��HD>����YB��8���~[�ҫ�1�1muk��@j2����m��8��g��,�4��d��s�g��+j��. r����Y�A~�wo����-f�3SY�M��;�
�/�2�>k���k:7{�q{���[���z_9|�TLK�D0���R�}��Ҥ��i��
�����>�a�f��m���� ���U#�}����j"z�%���0��9��:�V����T�y�\`�ɳ�%���N^�����iXu�x�z��0A�p:��C��j�$�š�@�#_����Sk�Z�5�u�q�tܲj7s%#TaQ`�(Ǟqz�<�'���q�����Nz����Ex���FZJ����۰���i4s�ö���ԫ��-
!��Ym��,��A�R8��V��{��i����t�X�>w>�����~-�������>��s(\�6d�%QABE���Z���.K�`~��3��l嬲f�Wo�@{�<�q�_�Ϫe�H��4������4�}*k�(.1ӿ���'��'5y�����~���u���
y��S<�g�; "QU���͋.����/�E�8O�*b�"?$�WMD\�=�}Ǭc�Ē�5�O ~<��51��+"�`��q&Z/�v��?���l��|��D���N�oǣݍ˖Q��P�-��j-c��X%T}��T{��}��P|oy�>Rs�[Qq�$�D!Ⱦ�tٕ�	X�y��Jb�ۏm��\�f�2��q����wr��Ţ+���D����QuT�rJ	�h�m��q\�
z�p��l��͍�*o%�p���mr���pr��C�	us%.j-f��R��K�,<�/.�B�d!t��A��̛�WnBg&�V�8UIM)��=#L2��5tĝ��;�۠8���o��Bd_��[�o�(UvhFq�:,�]G����
�i�SWc[r	m�*��`�pzSښ��}�£���[�Ĭ�YW}�hSx�I�7�QW1g��Zy#�5�z����(�g]&�ڦ�8�Cbz산�����VZ��g��.hrQ�WNR�+dhb�Q��M�zy���ç�'�82�I3J�st�ÊmJ%��j2!�S�l3���Χ��c��w���Rؔ&����#w�R�ͫLG	�W���L�M%�cu��J<M�!�%%�oF(�� ��FmtV��]��:;IߚD���n��y)����}�h����$Di�n�v�P0�2�t�N��Ҙ��|�	/q_|����q�K������TZ�>A׭$"��vl�����YM�ۇ�����a�r�դ'��w?���ɺC���B��m��\EU���^�܂�0�WLe��Б�>l���"��B㚁��_@�ڸ������a����J��@7��N�����d�P�2���(1�/�k���tM4T�ݔ�^���z����[��W���L!β8F���s�q�cr`���/u[9c��
h��`}8��G*�F�?vA]�dA/�Ay:3O<��/c�4����;=E
;<��Q9}�*l/E�1h�e#l��`&U��G��[�=�E�/���y��y(��G�-�|Q*�����N ��8�����i�8.UU���S����Ӏ[2��
kd��*ʹN.<f�!ѭGv,�8�OeԃqR1��^�_ECjQ����4J��Y�#k��K�:GXXZ�{�pD~�.+:+�[5�s��"�%�������o���b��]��Kͅ������-oQKb������}_+�BH^``�Ċ�'w�K;*c����:�������K?�=����.כw��{�Y�Fo�3�I����WZ/J����|s}?��F�<�g���9�[� ��\I�C�"�I	��=�H�+$Ϙ�z[���������0���}c����:��nvV�c[-*�A�a��dN�����^����L�,~,�3o̜!)�J��'nԷ��4t/���;B1#��4��3�:�4zV�>�)�-�UN������nyJ%o��|~g�uQճ]���9�qQ�WLo�0Y�L�c�b���x8dm�)�`�a�:����Q%H�� Å*K�Κ$WS(פ��@���8!�s���y�%%�q%T��A5�4l��(���>�A����:��R"-Jg	tF�nW�e�7̦�C�a&o����է����';�W%�o�	q�g�2pl��zn�o��O�.u��nk�Ͼ�7u�9�4M�y|������p��b�b����q����_���i>����U�a�kN���9� u���ܲ}��{��unnMO{ sP
��1��]�M;(�"i�89|v�A!6qؐ�b��K{�p�_S���|OW�ugkL&>��2+i��a`|(�,��D�<�����9��:��1���4�6R}WFYR��D�4���H)=C��.�������Hi��xe�4~=I�]�8����dj?�P�yxu��$x3�
�����BU�>�h�EU^�Ax%��%�B�
������B+b9텠a�@�LX��H3�?^l�D	�-{����E��xeĜ�vND1��ݰ��T�X��Bn<�GD�5j͸�a�#�����7�Ԝ�a���v�	E:�����%X~��
Rz���s��@(��4~�Ӥ�{�VV��M�{�4d*j�� 9�k�:z0��<r����=6��#�Q
6l�O�o�$��$,9����l�p]����E:	�;1�Wt�b�a朲�k6�7��[��� ���Ls3�� E+��ѭ<�/6��P<_�0E~�	�ѣ����6�lm��N>�/@q�HV~�&S��}���'1���� ,�(_�������NN���4WE��L�fN�����$��H)���[)W����?j]���I�9�}Z�i�1;��NA'ps2ѽ �+�~(;��ӛ�H�W��?�-�(yL瀊Я_-�c��[�����S=��q��C��_��#G�tAI�V�N�=OR��yT@����`r�|�O�̭���* ��U3_���+��,�٨
U�ό|�������α�+������%�y)۵���p1XG�U�WR��4bE܃�'Jc�%7��Vk���`�4$_R!a�������/��YF��^�eC=���'�`@�I�D�CŬ���0��5��Ɨ�J�n�,,�N+�lo+��m�`1�E�����9s���$�H�P8<�Rѿ����d���>�f�8�?¾
ɢ {& k5��P�@��^	�B��M�(pq�D!͌�^�ɮCu��y,8�G {��k�}0~�u�7�Tu8�,&����yFd������`к���h %����L�3d�G�<��x�B�]��_x�}�u���_��5��U��v
���l@��o��M%h����v���O�<f���X����Y/}1� \���Y}����ee���n� v�������	M391�.��a��I�\Q�A�(DB6� g��4������l.[�o�cse'��,�PU����
�;�|� )��ʠ^�~���'<���$���:f\�$YWX�0�*�8 w˴�0�7d�T"N���$���� ���C�GK���l����E�o4-3���Ց���D���J���t�+`%&L �-��l�<+u����v,�=:��x� �d�%�h��v��m�V=x���yU�ZH��0Ui06	K)�������g����qل5�@.O4������|��+������x+T� ���Vv���턾����'�hd�RWH(0&�`��+o�o �%��%)0��=x����7^��ff�ˉ�9_#3d?$�@4q�������j=+1l�K%$�#��!�c��qc�H��:�[�@�ݭ{�.���%'��D���Rv�l�S��;e��� 맒�u�Z��]��ա��W�0:�o�R��M���Y�!I�`�TҬ����i��5�z]��h/���m���l&)�-Z"���UDj�$ԯ3����~&�E��Zb�hװäo&f�}�=��bl���*�ȡ�[�\K��|sJ�� Ds��d��\`L.�a�P���z����_}��(��.j�p-!my��- �w	"x���?)��+M�G��>���u�gZ��� �T�CS��d��t=�0�77r� �׺ָ@�Of�~`9y����3�隐�n�H��ݢ�g�>��v�l}���d�>������?B�РkH|�9xFj�b	ٽ�e�k��.�M!�)��Oť;�gwh���
��ޤ�hC.U$�|4�t?MP����VM�B�"��\���xv��9���F-�)�>vn�M�� �.��<i݅� �����l��"o��~��Z8�����2���$�R�u�; ľ�zټ��Bh�Dl��<��Ĕ@�y"�ʡ�?msw��,<�Z��c��*Bm��/�Wrj�wԐ�#�o4�׍��u^k��d9#i�,un}�Ӱغ�s��D�=���� �y�-�ʇ�鶠Hՠ4������_�Q�{��H��P3O5y�������%B�Mx4�a�ϏWG�{�l�z"|b�S��T�KriA۰�tΛ�VVC(gG%�͞pT$f�E�*Ļ�/d�cD_�15���*����H�w��C�<G�TR��*��GLC^�����ow��ѳ;(�i��Xz}��^3#�9 .���,���&�Kv��@�vG��Z�p��P���c@�ǟ'B�vY�25�? �%�f~�Z��M���=�xT�� ��}�ٱ��o��-�i y@��r\��~�2��6��	�H���,a��~��kD��;�|J=D��LPS���N~2�E���3Bf��NQ�ʸE���)�x�A#��3$W�AE�Ȑ������@��+�G�m�"��f�vlk��)��)�n	q\jP&�Չ�����{��-�����0V	6^�H_/�U��W��ъ8���O^�%�~��A�u���a��f�J��m��4dpЎ�4���� �ٙ���8m������ߪ$�(L����l�+�cdG��_�%z�(�2����s�bE��KlE��0���4w!�)估"AT���<������&5*!U|"�1-�>$��n��4�j7��%E�QZ�$�co;�tIK�N�Y^�jA��?�����T@�$�r�K�Q���쒶{��x�1ߟ��2���"��(v����.��LNv�MA���E[�� 0`��T�g\�_��dl��n�i��:��=p����f�B��K)%C��I
�z&6������h��I�tf�$@ҳ�$j5�g=N+@������q8!g��%"E��.�Y�r�:E���8Bk`Oѐn�OU<y��*[p����M�b'�cK^Zw2�uD�-@���y�����$,��8:x�(���R>Ï̐2sEU�����A�Y�,��k�"0��M��/B��>1uk��Oat1��#�B�>L��x��k M��c����� ]J�D��59R�j��J����!R���E|�1�n�����I}��R<ݶ�$I�hl�4!�b���k<�U6��<�t�oDK��+�����v>N��yT�OS�$%��$��)�����O�I��i��m�К�5.����,�6�)o;����.ꀺ�n}�ӥ ���{ b�*FB}���6�U���۞;�?_��	e��w�@gyf>e@��9q�c�-ɘ��QP��t�gp��B��B�1)�l-�VƇ:,�'����&�"ٚ�o��6�i��w��y��~����M�!'m$����)���:�-B��HП��ǕGԲ]
](��W��o�Kj3|{%�'��48�	[�y_����O+|��z�f�y�i�d&��}�nՙ" �C���#�����g��`c�tՍ��*��>�ijX�gZ;���)_�+�܉)�߿Y���5�^�j��'�۱�r���Q�A�/:�_�J�dL͗
|��
�gY��P5$���V��4>\�|ʰ�i��a8���(ֳ�z{�e�&6s�	{z�hmv4v��v���T�W���|]8��|E�p/v��A˪r�8�=#��~.l�S�A�6��M��-�P�F�X:d�]q�MP�[5���{E�u]�����)܏�N)�
k�����o�>�TC���}�(��3�@�D��(2���̰³q�G�.h��*�ʑ�n,���n��F6���
hت�C7ؙq�� �f��q�A�<���74�z���z����,*���h]U.�q�k<�7���d:DV�������R_T�c[b8ɔYq����yt8���!��ջ���$�����	�l��05lZ<�]�%�g@��
\����ۉ�d��8%��H4Fnh)dxo���4��a	��B�A�#'yK���e�TNK~��f�w��o�����C��<���ǗǓ֋O]�dGՃ��f��n\��*��O�X��f�3��{ҕ��Z���~ycA���:�y��0�q�p�v����5h;�߇E"�e��[�����Rn$C݆@%��E4��$��c0,d7y'r ��P��yr�zx��uKt�G��g�>�y�P]�����u)��x�j`"��rՋyq��vYW�T��d/t<5���s���������ۄ�an�&W�ڠx�`L»��ଶ���� ��3xX�B��I���߫�k��wf���A�_�媘	ɏ;Q*G���+�b�����8Fm�5� �`9UQX[��TM����}�,����ݝ^�+y~�D��O�� �u��KKJ��W�w�=g �z1�O�i���{?�F�+�<�&)[�Y�J�~��3�ӄd9`�"Ȧ�F!M��s���+�Mc���̶�pip%�7��!�]\p��Ö����Hh���v���*�T�3Z�������{��d�-����~�,������������r�z��\�6�V�J���������\�J�{��ҚZ�u��J$Xo	���s��H�����PW�P��y_#����Ee�ȳ�נ��
�2������:��>���A	z�_��M�(PbIŖ0��f0޺����e�Zd2G��K%����BB՟����7�[@<܈Bф}�\��"�m5��A��c��-J��{�i�F7J|d\�tv��BM���z$gA�F0%���eY�HX�@�{�IEam��k���mTi���/P�;��Ł�l=��t�g�R�[
	�<�Ί3+��;�+"�T�_6pc���M��X!�O���7�����l�zfȭ� ���y�O�W�
�j�Y|�)ĺ�S�8���;���T�\!-�|0��E��m�,�=U2�^Y�N;�tKi�^�Т	�lA�y\|o��qM���|ubJJ��
�	�"(t-�7�zI���LpkYVj�asj�b�bg�T�N��kP!!���>_Zf�Q���Yo޸�2��͇��!��fǤVM�������x�������(J]��$UK57�d��	�mG�<1V�iF�/��O_Al؛�G��/ 0�m"�Z��+5�9�[��xuU&�0DHB,�?��Y�i���.Ϛ|t%�h.@Օ�(��o=�SjVM���af
��pI�;�B���BA��,=�菧�v��hO�"if
˜���>�(���S�(���K��Q�+z�������,S�K0�wi���׉�gx�y��l��,�"P*�%0�l����ܟ��؎`	)w�n�p��C��C,ؽ�dJ��>��9�P�X�m�ER��E#�Q�!����Xx�u~B�m����m3���h[�b�~�E\u���@0:Ŕx�-�6�z��Ȯ�k�J�w6:��&nG
�d��w�<Vg��8�o��o ��#B���ׁh�c�G�L>�@�H6��(,X�Usuގ���p��z%Rl�|:V~���t���]���GP�Z
�U�.R�F �N�/d��tv�XAC����є�}���7��}��RT�T�ˈ�*�4qA�َ�Q��nay�Dh��k�O���p��ńF���6�E�&`�3=�$�V�`>�\�E{lσ~�<�T鹍DĢ6F6��e�MOW�}-��W�!<}����@n|�]��hAq���}1���4��(�4�R&D�۽k	ޠ'���?e��9���V���h�HQg�pxT�R?rcއ���0N{��S�iF��|�c���$��;M�Q���T�p����̵�����XEl�\t� [wxv<��n;�N+Ni�Л^*�����\��/1��˵�>�i%���@-[+v|@�J���2w)�<Y4xarN�