��/  ��Q(���]G%�B�C��G�1�*�$�^�Z��%�������[�Wq�~`�	v�.@s�Yꥱ��+[q�~�����h\x�W�f��O�盁G{b�]���i {����~.q}<�	���`�� �)���(�c�,��e�طɍq�޳n���6�����������HZڠ�I��Ƃ�b�_��c�hd��N��q�f�M����t9���཮�l�rF�$E���`sQ��<#��:��嶺&$��pwe��������0�%�)�u�2wű2�"x_GC$u^��#�X�f����X�r�{@�����.:�iC���^1�2pi���l[�}cZϰ'I�8�Q*��9'�G��,�os��T%��>�H��M7Iqf�x�� ���ǵ�X�L��I��SF}�΢��Lz�
����c���3���b7E��������~aiiۙ�]i��ʎ�ay�8e�*�T���δ,�J�0#i�ԯ/t�5_}����؀�ŀ�LEi���0���C�Q�3T\���ӊ�`������*���hXf��BU�I��Y?̡sW�§�w�d���1��<�Ж�QM�:=d�l��'f��(�"�'��[іm������k��q~�l^K�;����qW8L.���$Q<̛j�|����=�gjUOԫ�����{���ɞ��sǓ���_/��Ԩ��|�������Gx7������(�`ݵ"o�t~��2)�D5E���ZW�H�/m��ks���-�����2��,g6�/�gl��9��wn�tF{�$LU�;� KC��+X�yE��8 �F��Q���0�y���oW	��B��y�"i��c	k�Q�����˒�vx�E��i�)>|h;U6�~ԝ87z�)�s8s�ȁ�zn�z4�+�<K�x�>¸F�F|i�OhOӈv�
(.F��l�B��n{)Y6�B�y��v*���N<]8��6�S��ƻY�����U8[��'�ط����&�[?�Àu�;Gj�j<���5��H��mj2���Z�����W�AE ��֘�{�9��Yd�!,��T3ް#��h;��vS�agt�^'���t�x�:7c?ƞ�P���&`aH�����)z��M����g4!Mۇ�tw���cp��._q�?�N�G����-7o&�A��dH�T�h/WL�	S'���Az������v�Yc��Q8nQ��>ӿ�::h��9Q�(����y��ϳ5J�JQ����$�XQ�{:�S]����ol�Ĝ�{�׆��i�f!�0�/̂Bt���z{~n%H�������t.��i�rb�C�`�$��9�=k҄bFCۍb+���YC+9/���v��%���9{j���~�� ��H/�;�&z�ùZ�r�Q��=��~��am�{1֥��_$�@�D`?Y|�d��NY�r ́��W��<$1n�%��'�]0���6�V��Z�8�4��-B��9�k?R� ���1W�y��@��9�,vv�T:����x�Oa���6�/%]Q�Ew�C�8�K���E��0�C���&��`�"���&��Y�5g��ۤ��p�w���Σ�'���rE�&~���a�Bhl�$�wL(�,����6g�w��vm��~t����bqQd����kR�!����Z.��̦5�N�[�ÕL=��eZL�F��փ9�V�eB� !6�5y��8��1qdHZ�y>��1d�h#�'�m��3��A��^�W��	(P�٭�?(���� ~��Z-�:���VFFq�����~�ol����q�7�RNU���m���ewb�?��F��ך@�;�D�i;�;�f�L	a�q">
��8B.���$�C�#��m%IhuQ7��-�B���T�йy�*6��
k��|���;DnR2ƒ���3#�т:k�M�xC��"[�ou5��Ƨ���ˁ�w(��C�<M�_�1��p� R�� >g`�>X��ua0B]�,6����&�/�pG04{)G��������G<Frn+��gK���Q?����5s�:��h
��T�>�b��{q ���zu��zr��o�E�gs���p�-�+wG�i9���)n$�ּ��<5a��"��kx���h�U�E�q�N��ae��]8u/���6�K��G�����_��n>7~ns9e'}�Z�Uȁ�6|چ�[��Ú~;BP���zNFύ�c�y�����z���#H��z�.����$��8$�W���Z�d���tr� ZN*y$N����Y	�v���~�yqA3��Bs�����)�\�2����~N�Tf�U4���^�q�i��U��o�'E�^��u�[(j�5ޓ����Q�Z�ECUl��@c?ȧ8����碍��IU�F h"�cG�N)��K��#a�8*�\��dbp�(���<�����;v`�"�K�	ya+�>�!���7��4�q��1��Z���Q���P����s�\l�TCuq�M����p:g�a
�Zi��7��O1��?@>k}Ը�yU.Ġ���H�����Ys�=��V��KCY+�6
Ǚ6��.`h��� nch,��x�'�7�Je7�܃�uY�%�c��n�"8&���;���R�屢s��N�"��i�ǐc�V�Fg5z-W�)��F����Yy���ax���/rh��]sL�bl5
Ժ�슥�?[EL �݆�6�հ���߳U����
���:�GT�C���8%p���G�GysM�O���Y,~q��$�Ȝ	�w�EA�iGc��+��F������Mg?o}�/�G����3�)��2���L_�h
{�a�=dM�_�yu{}�i��<��\��7��~��q������֠�`��7�Oۢ= ����SM7|_�.�Y��_�BTu�h �O�(@IdꐁzTTx���и�8Jp�\�lR-PqF&x( ��u�H��->����yEG@�,r�\*y�Y���q�P���x.�J��bJ9b\+�#F� ��+�/��0e��Ю��9'�V_���M7���T���Em�l�j�c����bí�ս�c9]9����0s����A��I�)}�E}A]�7W�ض`J�R ���
��Pob�T�N��}��z�:�F�i�I�6)<)���5��g�˄F�H?Cw���1�O��[�p�x����0*�0VL�4�y�C�V�w������Ԥs9�Y����ğ?!�]���E��
Z�&Ο����1��KB���M5�@�����-�����38k��p���0�Q�� |��c�N}�^�ߛ~"�Ű�N=�_:�#pU�1�;���k6�m0�	N�[]s3����cت��-px���Z��ߏ��&���U��R]ʀ��I�F��l(�S �s��!�ʬ�"�R->@t�U�ʔ��*�T��
kp��ƛ� dc_P6h�՘�t�3�|9��-��R~����;�@;���b"Ey|��)T���q�rm�~��n&2���.�ur��H��٨��c�]��<��4��	g��a+)�M��I/�&q�`X$+� �i!��:�瘅��.m9��C	�6/�u���_�`To��1��f�B��n��Q�%�Uւ634irSU�\�!/�A���)<�O��D0b�ڬnH�����N+5AK��o(O�j��~uEc�ϯ�@LsL_�>*F�����9'��6��'���jAi3m'��C	b��1�{8��q�)_�2���$���>F���s�SI���.��BG���*t�>���xqyN\�<�<lq��uIq>�ݾ�W���Q$y��&LQ1,4���J��/U��ޛ�*�6*ጤD/�^��H'<c�Ǒ�f�'w	D_���wQE�D"~�O¢�@��h����?�Kp٤�;ù��H3-p��v�U���J�coS��j7Px��`�`�N~Cx8HP����b	<Fy�u ����G���^��zO�`�����<H,	�����8n+��H)���9=]<p�Z/�פ�"ٖ�{V$��8A+�������N����'%�~�r���i���n�����ڕ42_\b������7�P�00�5�9(��ډ�d���֬�h��X>Yl�Z��j���;6��;x���ǵ,>��>Vw��W$Y��NC \�Z�B��]Do�^p�����P�~�/ʼ� ~ܥ����O�ߡ� J
������"�R%O�f�� ��Ӊdk�D��4�މ�����?=0����q��E���0X�ju�v�5�%�%<ޞ�;Е�$�ܐ �1���n�eŘp��NkFĚ��Y���7E9�pD���j47�����.�_�J
N�f�fG���*J[�MK�,��������I�{�1~B�WH���1��՞�N���	.k��YB���[,�4��F�����p�ǈ~vꇔ��'�w:�h�C��>�{��G�_*ѠvZ�7ͅ�E�R]\J?GF�M�oc��N��W<��v�9�n��8�4\-p�y���Y���Y��W^ޢ��yd�n�� A�פ�ԑɃm����K�
�s�O������[K�3@u�p�cFi7O�9��E� &��Od=�n���N=�I�Oް���,����;.��#zR�0�٩�)֏�vSi". ��z��*��Ԓ�Lڊ�= O���TK/^u`�oCj���p�sm"9���Z�ɂ�Q�DN��8��0�Mw�#�̅����/���)�Y���N�G5�Cc��O�/XB0iU�	��g�x-*�VJZX����.-U���P��wV�ωz؃$�>T�7q9
����~ܓO����u��K)h�
��lU�`}@�_h��㲋��x�>��a'�� N�K�䱭y��WsV�t�3�ώ��+�y�;�}���B����Rl!@�B(S�r����VF����y�F��zz����ĹE{�%���3�5�'ښO��y�bX�����ŝ�Z�=���~!q����m���3��1Lp�7[g��P��l��eG>����穼�UU;�xUAI���t�#�Ϟ^��H#FǂN�Y��Iw��<���g?��GC��&tzNY[�ظSq�����}�����E�r��[o���#�֢M��1���S���u�&�pu��Nq�s݌�
��$�1#����͡��Ǽ��$|;/�\K����{�#s�.�۠v�N$�wESQ�^�rNv-.I��W��XF��T&�����X�I���n�Ѧ�wp0��$3�g�L)��=�<tWOc(ΐ's��8��'���
���L����Ln]�(4��A`�Sٶ�7R��sT���-�G�%���Wd��U�E����Rw�n�b�j|7i1^������*����<:�α�h��S8\'�tF�<���R�,�H�L�~�1�H>�آvSxң�l5����^���巚���N���|dJv?=+�c�ߡ_a�IR��(E��( ہ�DI��&PU6��D*�
� p��DB��<�[}��k㠆gx��P�A�c��7z\ۉEǬ�uv!+�O���_K+7�t�é�Ok�f�(�0m+i��4��R�A4���ƬL����PS\ ��W�cW���O���z�i�lXCq��NϵY���H��7<ɼ���l��,�<���z���I�P��2|�Y\E?l��w<�=�a�����,�+��Ɇ�dP�Y���ҙ��G��޲�B7R�^��`�����!�wX\A' lƃ�能���9��}��b�!�C��dN	.9�ϸf;��/ T��3��D Y\@WO�W̣�\�=�4���9�b��b�x.�s�"kR���;ܲ���]�.UqU���.������1B���&�S+Ү�M�Ֆ]�j�'�]�����S3�)5b��ZY-��}�&FJ�p�(ދ� �#x��L���7�K<hլ��6nK��Қ�~���1��{�'��)��p!���f��VK�<{��#��91 sI8���\�6��~h�si[���i�4���������j[��TN9���S����h8� �K!"TkX<b)u���"K|���)�����T k8U1O������̋Ĕ���O�<��u�!E	����U�(ޡY��o�l7��
��|�����8S���7*���IN��������5���#%q$g6Pa`0 �:n���K�W��k�)�T�#GQ*��T �>� ��.���
@��Z@���ڀz?x�
�x�� yutQ���A�hT��&�-��!�;��Lm����J%̐�D�����S�>5J��+m,�3-��nm��I}o!&�=��l-�V9v0K� {�L����O��:I8�4p��-�;Y�����_��(C'1Ii�A���L�À<v.�d&:ii4E���J5�u�����P�I�6:�N�����2
��#�f�~hW�ɽ��쥢x��w_����łH�J�ܧy�c������'}�ГU�N�?��$�����@����;A�ع�ï8*_�rq�#A�X^�G'�q^�zJ����Yi|xIӳ��xڐ�*�2���o��h$�]×���)	�∜�B��5lH�\�$%�8|%��W���r���h��JN\,u��悸��z��ђ10��\��{]䤄(�%Ҵ����Ɛ)�j���G0E4-~h��88��
< 4������>JU��X�vFf��,T�ш�?�<��᧙�d���r�K������������E��֎.��g�1uq��̥��L��J����j���2��&>i҂���M]V��]�(������ץ�N�=�I&�~��>��<�rP$�|Z�-�<ڜ-�;�y(V�y��L�e�oڿ_:��8JxJpb��U��K��$���b�q����,^��B�c�|}a�5wO���\�����#�y�A��`f���J����F���T�3��bM��6�p�!n$����hS���!�,}���;2T���W�tI����WÞ�kR��l�c�9Q��.�-�~>�v6��m,�q�w��z�� i�@LMtHҎxP���=����$�Ω���v0�#Sslb9�EƄ�ض���&G{#�Lp�^��=n��j!F��\�p���w����\�T)����u��ES��ZK�� �(v��[>���0D%�ϼMG0��fxu,�
���9+��7��Բ$����Ì�1�`Ѱ?�q�T��0�D��������)�ߦ��K<:��dd;R@���+ �����g�y 
X��:����=W�^� �;�ut�	�<^C[���LN���q~��9��&�[�O��1t[���
}s�܃��#���h�`u���ͫ7�WI�l�o8l��g�׈/]ҝ	����M�nd�f�8Ju�'-��((� ٫Ya���Ю�@Hψ�Q�`��F���L_���rp�t�Ε��f��;��r���MQ�7��f��^�U)�a���t�A�h洂�;��V���vR����);�^T�@>V����P_�%$��o=t+]�4b��H^	W��H�5�]Z�ݚArI��H�2��tY��}�>U�u��'/��M�R�G(�kO{'	�`,�d��9}$�L_!�a�p>���Y�fDk�Yf�ڃ�
���8�Rݎ?�Y��Z)i�Q|ڰ�HѪ�~ܽGPx�*���K�����r�J������؂[;N��YE��/�#�m>��&���dTz�ُ�߇=�qIE��7r���˲��^d����h<�_7�{�p �ɡR�� ~��&C����P�?	|Ï|�븻�(@�U[�!40�T�������r�T5q��{�J���h�{����d.z]R�u���;M|��х��aի��&�Q�d���Q-M�p��]�d����q�y�=K4<�e��Y�
�_�!��F;�OuJzM1��|�LW3u	0�*�Ld6�_9U`dXV�`�⃭�sz񌦙��i!	�=�m�������z�	s�/�%w��K�4�c�|Q�n���h
ruI�'��K��+���*iMՕ݌�U�i������^�"�u).���S��ӎ@Q��dA�7#ʐ��!z|����_Ê���K.?�q�foL�nh8���CNA����R��>
~-�J�������*e�œN,�K�-BNu�E�2��i��f:4�ƳG1�Ww7�ǨV9G)4"|Z�?��庿P����x���i�
��ᨽƖ���KS:'�g�[�R'��֋��WU�]��Y���)X�<�Z[QS�ו+��Fk�2Y�Fo��M��ϼ���y�6��IE�)�e�`k��x���~&`�ǔ�'!^�����9��jdU���_�V���(���]�sP�]n��Z��.㎨X�b+��<'� ���,��{�d��'��ƕ�%��0:1��9��������͸���pǐH�����@G�zj��=n~�Mu����-���7ĉ!���͵o�/6�l�H����_EJ��x�Ml>��YQY�:���k�ZdY{���،��(;�8�ǜ�D
�M�T �#f@h����bZ�i��P�U)�8��7s����I}��������ۖ��co�p
n��Syk�Ѕ���U�מ@�gl��ӡ�������� c5F�yz�D^p0�+�F��}��8��>_��4!��'dr�Ԑ7��5����}�|t�y���(D�U� ?��S�K�Z�{Oh�΂A�
r�Y��+$F���Sxid������Z���j�Fl P�5w����T��y$g�"��)�Jt}�9Wk��mY�k�+�R�Z���cg#����NSP��n]�ǣr.���2���_8�i�Ϛ�O�_���h+�yE�m�l�ȫT�5��=�kX`�ݽ"��D�ϫ^S��z��m9��܂"�|��t��:{{��/Pxμ��D=	H
p��fV�:��
����_%��i�6������=T|��%	� �Ѫ�2|	ht3W6]2l���ͅ����7�1)'�i1N��ߢY����@�''h�
i�uTfB@�K�+���Xp��Ҹ�Z���/��S^��
��o&P�f:T)�[J�&�.��oR�=�T$>�DIU!����N���+��$H��r��-H�Ku�J���@�x�eZ�G0ݚ�>��.0�0k_�cPDZ�>�,��խ��Y@�>S"��U=(��ˆГ|N�������a\�6W_KSN�fEL�F,�������^au�/��J� X�]S^��x����0�lVu�����F�(N�4Ǻ\I�=��e[�u\�D۵z[Ϳ�i��a��H�&�Y�c{�&���h�i�	~��u.�&�����x/��X�SH����Y ���~���Ց�)��������^Lق6�%�t-����7�^m@ɉ*nz)r�Ee��s ���p�d>z�ϫ�A�O�z�~ELΑ\�Ӱ�emYe(�!��}LX�d~�Ƕ�/k�)�����Cj��9����4��I��7���b*a�r-Az��匩�gzB�G��\ό�����j}Y���p�r����]ڬf�)��0H`� �p�Λ�sc���O~9f���.^2�?��`� {��c�,��zgf���g�N�+�Y��6�u��S�Օ?�(�=6^!�l�0�*�4�]�F>[�O�m.
U��B�)5�o-��;���h ��
2��n����g	Wf7j�R�m2<#=_y$1�[l���&��7u�铕	i�)@��AvՉ9���Ғ��z7�g��RΤ���'q�8�2�v7qP�9�bc2��&�M%�|�mO�[���W(������r݉�Z�#��a�(��O��~X@��%7oq���#)祺�I��j����]7B�=�kM��j@��]L�)�Kc���� �t#���1!���$|�Ðe#�Y��G�;}
�y�I�J�v���$7��z�֤���n��j�
�tݴ�Ym����L����a2��a2:l5f��;�'M���� �&xT)��P�%�#�T�[W�����we]x�e\F�4\�����3O�#"�,Aj���P̰E���Xi$R)���e=/뫪'�����W�	"��7
9�lq�4�Օ;��ەn��Y�*|�Z9�MY'-"#�[f*@ڵ�л��͈�"��x9��9+L�?��¾�q�L�qj�"m�=�R�+v�N�&�`q[�������?q���?h����W��*�����b���-M�#�7kBγ���� �8~���u[ǋf�����d�p�т_7䪣��'G�H�K���*!����yо�Q�$1���ػ�8JU�m�%��^�Oe���~���L�})%jz�,,z��j��y��8����3�Ե��O|�abǔ�A�M�S�K~��i'���=�b�T<!E*ԁ��_(�:�>_;o�m��sgH�f+�'8�	upy"���f&̹0G������>]��*Ƹ�����v��dm:��A߿8���N���B�X%ڤ�zV�\�����U�$ (j��g85�h����s���U��T��
h�d�aD�UY l��q	����xt]���Dߨ�[�h�ό��`|�i6���@�Ũ"�(��	���@�;��<�E�����vgvUI�Ke���r�>*IaJ��������l�ꟲ���W墙v$(<�=���C�>�3@&�����٢��A�#�}�ňGo�p�`�A �(�����ޒ1 �i~%h� I}Ƶ(�6�)6e�9^�#���?��`��6q��b�!�k����#�v����+ÿ�4v�`WL�RP�&W	Ϭk _f�Z<�Ķ��Þ�z�
H���n��Q��.%��'(�å&1�#���AAE�-��l Ch>���w~�H^��)t[�а`�ߚ.IqPMw��쨋�[�W�̏�{e{󫣶[�<f�  �)Z��f��fj����z � �f��|��TQe��M2�����6��Q�U������obJ'X}���K�p�h����"Ү�͑%���mE�Cup��%Oڹ\d^e&�鈺}�|��B��+�����k�7ν���s�x�٠s��|[g�R�n�6�Z�s�z�t��6�q�g�q�o��U��A��x<M��f�i�J$�˵�	>]?z
�E�ԫꡞm��k�g����3�F��/�����7��N�f��=��G��x�1��Z�˧}�&l����5�g�7Z�&V�Hak�=�RdѨ�9�?����
	!��¤�hM&+����R�����j�a�$g�hEV�er��c����N��'�g,N�M�#�edޘB>G��4S3�d\fS�v�.e}TŞۏR�j��}u��q�7Md\y�)JI��`
�ڮ$�U��E"_�T��m�ŗg�D~�R�޴��N�YMA�z	�&��
�{�,��4�  ��eF�s��Lro�@T�����ܖ��\�'fO���8b��T�]��kjW	����H���@���������W��U;%jr�&��͝�⬘��U�t�!u� ����2���,���t��`(h���n�hm�8�%`���i?�w��]y��B��T.��R�M��R�Ƣ*᭸#ã����׳�TK�w|D�-�?�HAB�vd�T@��?r�*z��T�r�U�������%�2O���h����}��/�Y��#�\�0�"se?��1��{����L��+?V*��Q��=C�{��@�� ]k��p�����Q����H%�(/7�E�5�њ��J�q���G����#���Z�6�Q��$[
0n;��jLq-��"��FP��	3�r���	��]�3v��9�^�_���l�E�D,J��ܐ�5�E�G�.��iL�y@�u��!�"d�	fw��"��̣O`!w��������5�~���V���(��n �y�Nk:ԴL�[;wϭ	n�!v=���[:����!&w�$:W�_9�g�VjS���O�R�\���lI;�֞&�i��]�s�O��~ ���m[��i7rٸ���I����(�`�e��ڧ���n^��b���yV�H����9���mtûL�f�Q�>}N����C\��_=��x����.Vz1����f(w���9��ȴ.���[e�-��&�ƔK��!*���~���`ҫ���o���{}?�l^�=��r:��3��vےT�q�vF1�&���2�z����HQt[�Ym���E�GJx�X�W�(�\ ^�N�;�r�0�-j����<nu7����oʋ>����O.��^���ʊM�`E<#�F�~c�L��
 ������KA-���@��L�p�+����X�x44�?t����6󖡒h�o�Vy#���c�@@��o$�Ƨ,�cwD�	kQxϧᇼ/�D/����A�e�}�s/�rS+�ħ#����b�ҶDCW�d*w���%���f�(�So@Ĺw��b#�zZ�	���<�#�����RL��C��3b�/��$̠�R<��,z�D ��M�)�0��1b����Ya��+F�r�>nX7��u�kZ���#�8Wt{k9�V�r$]�s�O[�a
sK(�/��v؋��ƍ:)F7W��	R��b6΀�\�.�_gz�]�=K>��fN���>�p՝n+����V^�򩇴��"=�ߓ�@��f09`C]��T6F`��C{�<:J��E�}B'��?
Q�
v/�4)::���� ��;��Y��9�C���B�k�k��7Y�QH���x�#��lo�H�x���;8J�&�o�W*�&��m���/f h8�������g��4�$É&Ԩez�#�j�j���hQ%����g���Y��ę�����0�>ý�='�_���:�+?���B�h:��A���Me~J9*����Z�a&��S�H�}�C���`�I_�`�����7b��+mŁGFPިFlyE�?	XUQ�[���'���>�W�Sjgl���u\�tR�d	L�dz��5���ʘB^�"�Okp�\Y(H�RT�3����Ɂ�Z�s/�I+˴
�=:��%p�Ɋ��q�0;ŧp���ռ�J-�2v�.tX���~߯��`
�0u�;Stj������mŋP9�+�U�Nڊ&s˒��-G���iHc�}�� sV�ů�>�c�x�v�Ȥ�W�L��l���R��{���A�V�zլV�S�R��dR�Bc��@wd��&�B#J�S�_v��\��kFҎ�7ß'\W�8��L�y3؛&�ɬK`�6|�	j7z�*�LE���YB`th����2�Z�J��=���,�D�E���ʥ����i\��'�{"��t�
w�;�U�.�@!6��b�Z��X��V˙{�5�{��W�飛SN��AF_���3�'ˑG&�;��.�-�ݐ;��	y���1=�f�9��ގ4�Y�j gH0�Jo�Dt�x�n��t���#:Z��s�W`Rb܍�5}��O�������ru��"X�O|X-1��a�!Գ-����J�%}=�l��b��
#؇w6���>���&�Ymǲ�TERa�r��N1�[�pK�z�E[;]9�a�?�2��?��N�`�������1F�!�mx��2iA��ai�pG��{��l��$"���յ܅y'��H��������i2_�mi��晣���R�]X�}�ծ����8��,7�VBSS��OT��>Z����@1�� n����T0>��-����h�E��+_'|�Y�[���5?��&A�F���3GhZ"�����Jۭ����o$MG��K������;�?�3
>߫���eq��G�·�VJHܦ�S�S���;���\����?,��$O�y��[��^�0=�C���ॎűF�������ٱ�<�FF��q���s'�]�}��qU}���Ir�����~kI
凷�4D.c	�1���ݢ-�[�|��^N]-�M�J�ǔ����L@��֜�iTC�ac�w�<T�7�3��3<��R���U��ͥ�?��tgE���;��|�����k	E�&�.K
bnÕ��$�����5�đV�8�]����LS[e��H�����U
�p3gvF��A��c����q�3��.ט�y�ש�܃����7������֛���R�7�ƴߜ�Q��C@2�ʳ>�fZ�V�9p��e%�����2O$q !?"�)��irE��GY��7�H6@�n��I���F���z�#h���)�*E�E�O�.Bh���	�\�����AqlI�~�MZ�=(�<?�b�7�;�MuS�̽�-i�+�9���=�t�uh��]-�j�?�5chM���L��F}�{�%T�K�������xK1<�0�������Ʋ]����o#��p�q�:��A$�G�j̍z�kQ�\���	�C�'����:��w������W����V[��ʀNt~�&<�7gĪ]��>� ��簳��L�r�ZA^6�F#z]����97�A܂���ǝi�p8�;pG���'��(����'a�m��1k���"���m�����g�ì78ajq;QT�X�+�� ©�g|�}~��Ly�2(��o{��4!��EA���|~L�כ�8��U��h��#�R���E��9��z~3s���z%_� �[Z+Z�[}�����cX>�����wZ�LhΙPȘ�)&AI3�u\�.��S�/5a�/I='�R�{��u�6�}A~G����	���2�J�y�� �l�����mW4:�(y8��v����̘�v�2��jeX1|X)7"]�vW���3����;#;��m��f�?A�l��A�M�+��j'���LZ_N�J6��v��c��G�-/���$M�	��y�_>�U�#�*ފi9,Z&K�@U��\j�0��b���d�{?�N���[=v�Y����q^~E��z%�-25����wP�(ͦ�	uG)�m�.dlQߙ
��(�z������|m�h'H*�|�>��β������:}��_��?��vW�eiϖ�/� kۖ��-�~]�
E�]d��^��r[�I�f���	�8	L�iꇯO�K%�G�U�ȍ 6G�e1���S��1����H���c�hB�:(��|��B�֛��&8,���%�;��l�c�&Y��uL)K���&ͼ��F찜�-��K$�&٫�� ���&��zq�I��F�.#����R����]'
oUt��rk��)�g�#�]*Żp��1	Z|R�b�UbĮ '��@�y�h1����6
`�u��M)K(U���Y+a�j�ىBW_D؉��S����Y��#d��<����0E�����`B�K�~u.�7?^�9�ջ�|�Ǘb��~���[ ��I��8MD�Z8F����]ƶ�2Rإr�l��FQ�����҉��t-���l�
;;x��e�R�L?޻��w|2G9����ntM(�&�����To�e��AK�I���[\��c1��"���p��h�59��k�R4�-�V�${��K}>��1��75`��]���.`XHP����s�V�w�*�c�!��\�t�CD��T~���Iz�d�"�	�L8�p� �`�|n�`r1��@E�1��n�잎�B(y2�\�a��9��S��5��}9��~ɼ;k\.�{�#�$Z��J?�B��z�����-�i��,||�G�f4WmGefߩ�:�`~�I�S��64a[Prj��v��&��Fd�{��PF�OX7�gVɤůn�Y&�^���ºc�����܆ĭ5���o48�8���\��B�_���s����������v�X�m=��
��8���Ho_��T�w4��.RQ��kkӲ��r$���&�!yð@�x^`u�jz̰b�t�T��x� Ԯ�r�8�l���)�!?]"���I翾�7J)򭕓eqyL���XY��"�#�&v���Ϯ���7-�P6��3H�k\�5<[���ku�fg;�.K��y�}O^T��ǣ�����R<Y���/�С,>�f9�vo7a/�����ݜ+�p��BR)yë��x����'%\���SN.���֋4�[�����r���h�@�CX�Vt����s�Z�5�\��/�B"�9z��U8N��J�����χ3��0�AQ�y�������GV�~�r�e�mނ�Y���KŒSxH���[���V)��dr�u%�Z斬h4B&�c��]�d�%�z�K���R}mOr��Zb��PO�w���p�*���"����҂��tS1_^����}��%!<�뼰׬G"��Z�b&�N)���9�P��[:��.��3�!����m��c���ԫp��!>.TINl��2��u�l�槗�Ǎ�IF�G`������w$��
ܸ�� W6<��R�'l����#_?�����VS���>+���	]�xaI����Ժ��N�UH��	�������,�$߉��4Fa$ڽ�'���b�/����E�����8�ۜڟ�a���ľ/��0��������[,�L̀�լ�Ϛ���[r��������v���L8�O��'�3e�VF��<�{�NL�lg��x�5������î��=.��D�|4�0V^�-_��{i=��
��6<7�Zcl������� !C�{�����iE�Wp��)a��,|ꍾ���p4F��1�Q�L���L
!m{MM��D9s!�l�gW~���oȏ���:(-Bc��H�������c
�S)��Xں� ��^\Q�ow>HE?�½��}���!���U�cP[9 	KG���Jr(�X��n��s�@%Oj㰸�����&��$�.T���ec�x�UҴ����� �ޤ���jL���7�W�4��a���4��f�3'@�л�E��^��c1�@�/��od��ؒs��"+]|�h��{@Y���Ot}��
7my��;�BQ�)e��mH�g��s>��i�fҹҵ= ��te��d�Xt�^<H�v=�6m�K'�_�&ϴB}����42B?0@s1�Ϊg��I���;V�[�LP����5��t�-�qz\�?!��U�Xۻ��*���8�c��F���(a����P� �^fi�B�9����Ф����V�O֜�AW�]zn�T\����Z���5诌#Y+���Z�zA���i�G��q�Q�R����U<7j����֘�X�(�x4�!:\�A޲�)����ao'ū�D�A���,��}J�h8�%K��m(�F��+��[4�����]4��]�inQ��7�Uc�������̨��MW�ŀr�����ө 
[��"/�c��v۟N/Ql�e)�UD�y���[Wq��\[h���<��=��py\�{ d}G��6W_+[Ƌ���HÍ��ޡ�%��5ϯ%������
R��b�0���'"B��I<�=wa"�*I�%}�A�7fa�����y+)�f턤�/ (U�ck��,Ϳ��rtϡ˗�S�1�e1 ����Dm���W�g��k�.�W�yz���gPV����9Fi0:`�JS���$a��M�X�vm~�M ��i�ԁ�g����b#�jw����1��G9���@�_�ڶ����&�V�<z'�Q]�VE����hk�T^��*A�Bn��4�>B���7�-_��m�{ �ȟ�Yl���b�wӔ �ɠ瞀���\�}Ώ��7}7������Q�BO��bP��3��dբ9��[��?f���w�p��� ϾX-_o���yI $��<�(�ة�F���v:H��
HեN�8�-�D���%ݾiiY�;w���C�w?��|,AeӉ�����\��8���^��(����Ғ�@�Ϭ=��m;B��X,;S�F��ʂD|�N�4i�6�m�����l�E�\ ^B��"���ĐGR����ץ�������h[a��՚��2�L����G|�m���޻r��Y�1������XVg)��@��kl��g��7�}5�Y�1��:z�������r�i&����ҟ��e����_��~|TXF��FA�\���4�+�I���!�4����u��� jʗ��j�O�)c}��mlz��?�g�Q���;f�uj\��Hu��s0$��t��^����8��_:���Y��l�ۗ�0�ݟm���Z���n�c�]�P}#���L�d[��1[k AF�B���OY����k���jk��C棃U�Ev�>L����Zv3H�Z��� �m�IP'q�jw�����+�e9�#.rE68������Ã��n����K�*�C�jC�̑\u�s�tó���G��֮�V Uo-�U*	���vm�p�f��;��P����K��Z�����n��7=��CG�I��	-Z9+CF����z�g���(@�)�l"���D��ڔ|A�����!'�܍�3פ��
?ڵPE
��Ͳ:��[d��X���r� e���^X!8�(�y�?&$c�#���1�	.��e�Bt�j2!*J����ƵA��?�r��	(H���(�M��ͯ�'E� �}[��g�W���O�$~;1��^�6!�?y���e���3�������)[�դ�Ez�B�:=v�K�����`��5F���pg2�~z����^�@��d��C��l�yA.���7�Q�	�Wn�ާ@�ƄƉZ��&�ݢk��x�����?b3��;�DH�M�"��'��ǰ'�V�i�M т�ߠ�#�N�1P+ə7�n���na|p�LS �x?Yv���ϰ�]�,}��s)��c��l��$����r��8V0�j��<���z/�K�Pٸ �q�]�T�E��]��a,�K���^Ei?��,�Q	�U��3�S3���4���]]E��SsGR�;V�_�9~A��~�ôr5��N�H!,p�[��F��π̰bGg���%*J�h �ufX)�Z�$7,Q�VS�I��uO� ��EO_P�Fan@q~�c_����Mx���D�Y�Q/�g�0?r�W�@B��e2��l��y�@��9N-�K\棁M䤭Ki��c��v�5L2���.��Rk��qSٳ��N9���|�!��{ُ�8�Y�O�2T���r/���,�{�W0�8=�VF� &�N�h���2�����BqZ��Y\��#O�5$�������g�i�w3���n����P�D��kS2�G,j�1+�l����ݞ3ny)]�_���֝��@���i�_��y-b��P���,��~fz�
s'��PG����^x��9�9$3�sO1K��n�;�Ӧ����5�'�� ���5]<���}���/|dR\��4Ϧŀ��x�i9�*�{$#'�Om��gG��k���Ak���{1�4m��˄ČLs�7Ӿ=��eT��N���*���<������\��b3˓,�.��ߛ��?Y^�����������v��SW��ۙ���#��[ ���v/��"pa�� �r��P$,���1�ƙv]8Rt[ֲ��߼u����!����͝q����9𑱊�L�]L�`���+�+�~<�!��u��>�׾UY���Q���p��������ε���T?b�Ckh���vE�j�[ ]0�=�)��.+����'�"?	U6�+7�D��n�+'*�lp�	�}ŬD����ݵ��'��d��i����-=�N,�>a�(Y9�*���ufx9�L����!al�? �c����Cd{�	�
Y���!=��-}�~����0���ɧ-_He��-�s���7��s}�\���P"_a#�M��cR?�f�G��r�uVeBT�hg%K!l�����e�`QE;���2�s�y�!ʤx?R��*':Ƈj��ک����F�S\g����C�d���jD�_�l�B�΃5=\����+�c�O`�І�`l��t$+І��cX'��!*'���~�?��t"�Zd�pC`���Mm[�а�_���~W6y= ������yj�)杧cB�N?W8J���T�,���(o�O }�%�݈E��d.�2����H��p�e�a��0�O����Y?�l�aW��䑕��x#���]�C���`�o�gJW��&�K�:lA�����n�t�;�o�d��p��Գ��s�����h�}�{�"�ӗ��}���� B����RK�q[�%Jo���W䊞��UD|��i7-�K��lQG�,�EZ�-?ip�ɶo�aі?����z�g���~�5�J�|���*���$��%/��k�"Mc�w�,�.�P��fq�c�L�A���FkY�p0����k-7u��F3�ryi�ڜY� ���[��� E����Y�B���@���.�rY���<\q�����vcЏ�������]�qoh��s��j[������~��-�=T��ŧ�L�:���~ǷGn!)�!��r����/��U__���l|�7����N
tQg/��V���c¯�x�m:8�t{!f�CA�ÃK㙆~Z0�t_�:dC��>����	?���ʶ�V��O����jC��
�גpJ�!��'u�&D��Q:/!������%/]0�	���9R�OL�:X�9�m�2���9ǭ����ؼCtwa�
�򢔱� ��aO�xVj�*�6��F����G���x=O�5��)z�}�/��[mk��q�����:z�n�k�;�d��ޤ]�s�zz���Tx�V�5��#~�����S����$Ir)pb����M���j��)A/����G�aE^�A�$���%��y�;��j�"�(5� 2{��������6>�|0���Yf��?_]�V��q�Nl�B,]+N��#u-�kTw����_aek���0k�1�o&��	 �x�g%�J^	�0�Waa�6v�8����~h$������Q�m�⯰
��&�q��<?��t���GÐ�>]��`A@�Ġ���}���mN�ޟ���%2h��2��Y�wL�zpvM�~���V��M�F�V�� ?��2|JwAԹ㕙sXs��M��2@Ѽ6��q`���~�M��%^�x�&���6o�7�����{�8�M�g���$��0��~�P���tF���J�l�JT̫�U�:���x���]�Z����/�u�c)�~���N�j�?�x���~ V�~��̄C�Y�+	f��9��N�C
- L�!o�5���M��J����[讄"������;�O�W��a��������J��]Sx�7 �	�h����!�"� �zK�pWk@�+���E�4㘡N$g,��'�}���M�u�U��{w��^�{�%&>�!�RI4���{��+������*�b��Q�ЪYPEUXA|�v�:{��@���ܹl�P�:��5��݆��b�Zc�$�LؿV�躴o�Af�m}�D��;$w�ڙ *q��V�0˛�)��CM���h!�o��/�vC��PsL0SB���zP��`�-WH���
�߲�K ����T{�m3M�����{�M�����R�y��C,H]�δ�97�̦���J�)P�
�턒��M٠�+ϴ��b/�sHϛZ�O���j��K\�]��BL�5C?���9��
t`.4BuvD_QCP�˺<-���]��x믾;��$�ϵ�n�g�d�쟈��af��Ma�]���u�<o4F�z	���sX�yˣ^���O\���Oy>C2D��>�g��_�]��^�4�Ȃ�~h9xT������j��9��nc���]�/m�2=���ߍ�-���*��T��
��I�'@=5� ����x��;��)�	#j&9X!������e1J�x�̗��7�kJI(��v�u�K�~��PM ��Вs���$wǙL�l�Jj�>	]8_ڇj��B�d�A��D�T���'�w�[&��Τ.;S���R;.�E1;�Pq�i�R�	E�ME�v.���Ϝ�l�7��ڤntE�U�AQ%�[����:��m���A�ޡ�l<�i�����E5���笶����;���2C��h������*ȕ�����	�����ƙ��9�&~^o%
����#NX��),�X�����Q�b�N=,
m��W͕��-�ܼl(7�sI���4����<4K�w�6}��	B�/W�J��4��'刢����`^�j^,@Z�!P -�E	���ת�Sy��L۴�M��K$;���1^Z�RC��%+N\��\{q��-ud@JOv���
<w3YM��6+d۰��.A=OqrP%�<'��r����*ޢ��y%ԯB�u���������-���~$����g?my�QX��֊6P���R���KT�8xG �#���X�����	�ֺ���##����'�8�M�^����E���o\ܹq6�y�+,t���/F|c�0�Z���Y�`և�r�i���4�E��.�ژ\Y�*ʬ1�l��|�ܭ� Ƞ���-/�Uy]u
�F��l�4k멜M +z��^�&ƂD�K�̛	�����ʧ���=�d�ʠ��U(�T���V�x/�P�B������cV����M��3�x�-��{�p�c51��4�j/���*��(�Xr��e�<��4NmK��9��9�qv�~l.�&֫6��Z�9ӹ�᡺/�yf��C�i����F��;�2��3J�W�a� ��A��d�7l��$��;⪙L���8����y��r�p�1��\E��[7�o����3 ����>2J�2��+���<@p|B�dҧ�2tԂi8�CΣ���Er���M,����^��L6l�~N�O!rz?l����$�kG@.<��G�՘ױc�';k�Ó�2l
^"qD���o~��!�K/TӉ�cTs�I8�	�)*[��ƟNFa�*�zT���u�UG���"W��(d��ed�0�+�)����d}�?��d��&b,$���3�V��F��́`w�P6�����죂PU>G}/H����P�`��j+w1"7L�����1q�!&��\�vf�Z��_��0x�(��1���4���՝�Iar��B^���4�}����,5j�;���3ڮ�(����I#�)t�[6��$r����w�a��A���n����x=�� ^ޛ��U�E�y�K���<��]�<���*g�]{5�qt��QC��2.�KT�H�ͧ�^�|�������~(��RBR�̙_�6�)J6s�r@o�)�ήm���
ڸ�Ά�~���u6��w�0)Ɵ��#�E:�������������Xi)��?ܚZ�e�b��uT\��fy�$�e!�
V�����:3P�8����.�J_���(�g1�i����!N�0y5�Ǉ�s��9> .�ao������Bd�g2����E��OG�����jC������=�E�%��^��l#t�w�O7��<縞͑�3��SΛ��R_ܤ�β����w��$~1w�������<��y�R[���=n��M�$=��Ѐ�.��.�	�m�au��tԇ�.��~�s��z��Z��+R$�롽�@P�1N�k�'��	�u:�i٪��ӌ�L=o�O=��OH�?l�
�������|�����Ldx�S��)jA�с`�ص�'��Vk�v�v�PI��=駏�g0_�_���?;\C����\Rm�]�>��i����~�]�!`p�,P�E��!��XC���(��c ���@J�P�._��J0�1�%��C�݁����c-��}Q@s��J�#�e�a��`%[i�;�i���P��!���ek*�`R�$��~@mx����;>�;�z����њ��:H���&�����Z�2'�j`Fg��M>d {��zNP2bW���d��L@$�R��x,̻+_J�� P%��nՑ�܇�lЖO��nebV;���;���ര$�ˈ	g��c��O��H���?y~�](�(vҮ�И�7�$���|頁��}㣋��ѪU]���������}����T���C��B�%~�<�g�Y�ml8V�XѲN厪^N���{/��{^kU�WGb0"H��\fHpD�m8k�Y��~����)�59�#=�&2��^MF2�:#��~Ģ<0��UEǔ�uoj�@Wv� ���ߕ,��.9����׭����g[�bѻڱ�*5f?�e�
F��)���)w��;�����LUԩ�s�i�J^���iOÚͲs�[�g��/i��
��u5��O��1��UK���](�#�pn��r2ss�FVm�j�o<���_��W@�@������<G8�@@�[�Z(�CR��H��CE�z�,�P����!��^�o�8:rycn�@s.����<�m_�/}�H)l�4�|k��U��.:V�2?/�7	�Y���,���,:��VO�{�bm�ȕ�Fa6����Z�J�0��J���nS%�s�-X^̜9�B����`��,D@�����Z�]�����C�~K��|��	b_|[�b�#�����Z�)ܘ������)���'��up�5Y��g�;%q�>�Nx�[ E|5�!�&�@5�a0���%���^l@L�ˤɒ���k��h�S/�_<$�H������rc:�]I\�l%��Ep��|}`xa����Wc+���6��tʷ"��Q��!��J�+P�����1ɩz����w�;
_IK���ҔI|k��nQA�/������+���x�>1���R~��NFx���Da=w���ϼ�D{��o,2�')vH��I�cn�������}�f���*E�2�V��]Y��-�;��l��b��7W���S�z*��/V���w]�f=t�Q��S�W���M껎�4O0ȼ��!R�v�x7���M�>�xX�`�[��|�_K�T7��ۑ8��~(,_����N?V�K{#Ͼ4�J+&A-��bD4��%E�v�����I���
��N!�9�՜l?�b�m/#H�����-���e�y&�QsE,���9���7�'�b���J�6(6���5κ�,��e����x�ɫ�x�5����q}�d/�>v�/�I���("�G�#/�dY�/�m9P�=�r(�w�G#��h�#D֟����Z����ۂ�����SC�V�<I��U�*�����?�or�ь�����	c�F�����yX��^Z���"~��4)��vȶ�Y�.�&�֯	��Vk加r�B��)`ہO�o����ClH�:؈�4D�L��RXV�#���2������s+{�G��\]߀(�k��e��'�*<�y�1:O��*����ʕڒ(4.S�.��������A�\WQ�⇜oTM(,�wn���-U%M�������l	;O(���,Y�G�lpN_J惶'�߹�(Np���E_��#�0�#}|��s�٦s(&�^�SW3��?����k�jh��7����T�+�5G��$���`��)uMz�gn�f��:��g�Ld��IX�+�1`	�#3���b�&�C�KCw��v���W�����eǪ���3�F��FO��s
��"E)���QV�[A,�h/ʋ�V�%�nk�V"!��}�a��B�4����dc M��շr��m�ߡ���Ⱦ��#F)����L�B}L��i�껾?h�,���S93_P�v�4�0��~dȧ8�����)�X0 opYU��w�{�c��:�����$AǊ��Fɰ�{��٦�ݳ�3��9	�V��A�.�q5�N{���oJ��f����H�~[>�zJjnJ�@�L��a��O6Eaz'�Y�o��aFڰ�`$��6�TO�{�&%9�Zn�/5rP�l�}VL\z ��7���ti7	A��}�j��@)V@�9��'. �l6T٧2�r��H�ʱ�)j��y� D����=���j�6��W�?��?�<�.��v���{��"ϓ٪�p�.EGa�1��;`�d�0��v'ζM�`�����[�-��;��)���C��O�/D�o%sJF�ǟ�/�~�m��ag��s�'���r��3�]K8��\q��p���F<���J�B��T�[��W|Bb$���)�����,Ӝ�49D"�ۚ��y���r=�b�����r��/�t� �Ύ0s��c�� O��*�E#���ꍩG���n)�m\0�uI���Г���ޫ��=����Fv��t<k~��:[7��=N)3G=��f�įy�<x�}��톁����9<����'Ԅ'�i��'�t;��p�����=��=Q�U���1��u᧹����Gsk׽'��1<Q~�&y:.���S-�f����ywY��x�I>�VĂm�G�yy��b_�4}#^�d���c��
8�G�)���eZ���I�N���<FSE(��8Ĉ�8����eo��Gj��23guu8�cz�ݮ�#������u˳H�v�#�e�*�|�p(m��ɺ�OC��ԙ�������堩~ '1T^��m]��ak�ގf�]>�F�Z,cѡ�F���$�5Y,�V��Cr�(ju"��[�������d��*E���)<W4|�%a��x�je�m�!6U;h�/�V����M���Ԉ������R�t��k�j氆���e��p�eWZ&*�X�6tҶ�f@N\����x^�L�3r�=���;���0���[(B�v�e��}��Ǫt0�7���
� H� g9V���x\ݥx��_��,w���2�8Gr��uکf|n~� v��%<��ʀ,�P�8��eB��g+$�}�8���0hw�t�LzkW�"��u}�.N�ޭ �E�=r�a���v��λ1�~N�
܋�ʀ��vǶ�����R���x�ۢ�/"�,x$���lf�b`�F��`&w?~8�Ґ~;�i\���Z��3M��E���Y��dV3_�>w�u%02/�kHQ�s�J�?5��Kmjoьh�jr\Y�&�e�]�8d�1`�-R�'"�`�h,p�y�#w�����:̞�����q��9�R�\������uE��N�.L�_�\
�_.�o���V'�
���D�=�1YތbO]��r#[�'+.=(��˙bG�`�ک�&J3�%����wÂ�2^��A�	M&)O�*�w4I�F�}�V���*4A-�6�d�(*2&G��EA�f�6^Auu�I�
9�c�U�v�+��&\J���,�>��W�a��t�QA���G�����<-���0�ȅ���V��m�Wr]���}C�K9�ȡ�K��(�(9��K�)�q����܎�7Ǡnzב�7X���w���!+Ĵ<M�;'8��v�t�œB��ڡ��'��Go��``;�����ޡ��P�� (Mx��+,|lӛ�*��O�	r-��=3�R�F�T0g��#�AN������E��j�q���ˋӢ��.'�W�!Ϸ�T~ު�>z��M�al���U4vjm�V���q��:!h��(�/ �'�%�N��!%HU�r��$��Gy��Μ���n1h�&������n�u��Vf�m�B�ۯ�r�<�k��1��YS=�S��6-e��W��V�HYܹj2pu=�#�PT�"��h�����Hx�'��쮙Z"W�B���]��K��b��iib�t�m�$�����5�W"c�k/�����dÃYP��UA�F��I�Q'�(P������&����nȖ���~fh�<�->�4i�-���_{���9�y΁x�Sqo�-.aJ�A1��H{��r.���dڅ���H�G���i�f���ĠPn�D��g�;]�on�^ �cX��mn�9*��%�{}�"��C�`��ǛZ�3��
�I����K�<dM� ׊�.����c�C�}�����
�)&ȑ���Um
(d
��xH{D��ovh"P=m_�f%���Y)T\� ���3<����x��wr,�����*�� ���4	�3t�K��`9gH�����L�������n�1��c^yT~�{��1B-я_��6��������Z���q b��=H۞.�}@�ʶ�X�3�g�.�͘Ҿ�1��jvyF�/�@�b���&�J���=}�����84~��IuvA23�2��d���d�n��7�l�ADVK�%3���������E<9��#FzD�xeH��|�-7=�����~p��Rķ�z��TT�P��������d�6Py��n���B��TZ�Ag5�!zR^w/4��Yƞ���ޟ��6<�G�����e�2��֣Ǘ�&z|HeK��Yl�l�o29}��g�bO�΋�j)�J ���ѐ�,��Ϸ�[{[㏹�L�Mv�:����꨻\V7��O��x�{H(y�U͊)�myᏵ< ��N��M��F�|DfB�x��tX M��o$��Qu���HX!Ԫېz(�Y��/*G��J5���?��[�Ǳ�x���H)t��.2�Sb�6g�5�LC�Vx�޺��u���/,T26�'��w�R]$��k>DH�CN��R;A���kV_J�c����A�5�֡��}�D�izx�����b��`O�d�l�aI��׵W'|��N\C7x�xi�;6ȞAZhi��ڤ
N�3˔gÁ��nΔk�k�/d�8�(�dJ6�;��	5w�հ&��5��,�k�=�̤5���ɑzH�~4`C<?����X����W����@��ڻ�,��/�a�L��3��:���rM�;��ÞR�)T����4�s�?�7�l�˧�����k�]n�L�րlH��p�8�����Yc	�_Y�&$�a'87��/Q@�gD	�թ�;���\����a�Gu��Y��= �Ӽ��8F7�Qy���6�}�Xu׼�~&/+cGA4$�M�S�ڔޛ�D+�}eKܣM�S������  �����N�Y@����Y�JS� ��J����l�'u�2���^9kM���L��ߔS�G�/Tδd��G��8�վm�#pHgMͲ6���!��C��&�#*�٫�*�_�I��C�l{��������	vP!S.%9j�U��0�d�@+����hUǀ9�7�د��^�Tl*�[�-'2�����h����(՞C�m��:%N�|��H��h�!y���ŖP�1Cr���5~��+�`Z�C�7>23�{�Y|C�ѕ��d���ܵ�Չ�������v���M3�Ey�x��wG������F��ifO���F��a�8�Ё��L�ɛ��k��a[��-c+PR���gm"8��(��Z�E�\x���_!�oœ��
?�Z��$�Ѷ���8pO6r)"�4�J�-*$Ө{��m��D��oz�c�mk��Gl"�[�\�t&�e9M	�v��"[㒆�?���k^�=�10�W#`9�6}�Cf
�z-i�7�T�/'#���n��`N��o-`O�߇���� TM��b��E�X@��]��;�Ra)�\�6'Z�`"k����~a�v=����(��B�t��!p}7W�}���&���:{9��s�]���xF�\�KE�pOF嗴7?g&����I��,��A��G�}���D�+N�K����H�����UZ�B��e,e�wX��3̮|O�eS�j1�� �tkU*����y=T�.&o�)d3
�n�;�8�U�!�Z2]�T���ʉ�}3]��+\��wD�^`�c�VE%����y[�a]��a�a��'$�KFYP���L԰�z>�t��b;+����u�UEt&(������<�aP�z�H���]�����i�s �7�ܫ���6��_�ȧ�؊Е#���K}>�	� Y��C�?�ZyOg8�x�8PƢJ��XtŪ�sB-ODC[�����'�w�Є� ;��o(|u�{�s}E��e#�=
ℝ{���c!Y�8ǟ�}�:�M�2i���[@�`P��b�H�L\/�W��v�ux0g��hk����`���G��S�+���@e�w �Oe��}(�s�SJLB>�]凑�d�U�/	��J�U\��$M��t�4%�-,�g�ۙĩYk�hʅ������u�^��ʏ��d8=�rSՍ���抑�Z�"@��%����@6��,����qRRx�:	2�R�����tm�I?������ٖC����@�Dt�7�nb!�:�А;T �v):+T�9��ϣ������[�$�=���R�|y�+�"�����R�oع��	�#�>����Ӫ����y��N\̭����Gi��UtC��F5�f�QX��!��J=/c��(A7m���ZcZ�U�G�����8�����9b�Ԑ�؅�/dWj�b�(�S7����e(��E�UńG�(t�:m��1�*&q埣EC��9��TT�y��<E�%X��L���y������A��]�B�����$��?R"��O�&��PU4�����AX��X��]'�B�G��y�l������ji݃`�[���0�lh�}�5{;;I*�9��F'��*�.Y�p�۷���yx��j��ܮѓPd�����[����3�z%u(4�?��wm�`��8~�=%��_� ��
��(Y#�Z���Z��?9S�� ��7����ry�PA����"��FD���G#�{Y�����1��w��>�]�/Hs䄝1<���d\x�i����<�瀞��-��(쿟4(���)�!{1!ͬ��k�y�O��UC{"�$�[纙�ջ$�/1���c�s�i�[D���XU$égd��ZՋ� 4�#7H 5���0�@�;A�$z}]�@l�T��i8D�*l��0cQ���[���E��s���w������F�[c~`;6�ѷ���������x��ˡ�8�7O���Ġ)�u�[��aI|-^��gPr�]H����	b�|Rr�� "�DrQ�6���~��/<1l�s�+�b�$����"��}v���n?|�����;��K��ox�FbN���8[?{�-Q�*����w��d[����a+�\�4x֐�x��6��A�:@d�;e�Ƀ7R��X d�p:�+ϒ�w����p� �M�S�'��A�P�q��5e���!�k�����CkN��F�m�\�K6��;���r$�&���ȫ�}��ʙ�֝� �;7�T�Yk�x5����
(tT]m�0F���(��W��yq�f+�Ak,dȌQ��5�{fRB�*�'�-\껨�.i��0vYk�+c��y�,�u���a�c'|����������Vb�j��;U'W7:յ��.������O��.|P+�oH ��Y�vÙT���~;�	x]��1S��Kj�������B��mG���/�w�I�I⊆s4)��k��@i�6�|sl1��;O�r��no���%ns��7ۍ�>Tp#���<5�)+�n�/��˸���!,*ݽ�ᲃe���%�ᔙ�>��iX�U��+�g�E�m��28(��qNDO��0m�M8:y��@+ �Q�d9�κ�5����9K"�Ӡ�̃��듏g���[�פ��+%�f���E�i����#�d�x�o���R��fu�Pjz��xC�[�P�㬙CVἂѧ�Q�,�zt0�#���d��&	��(��b[>���}���W:N��QV��*�ho��
�XC����b
nPb�t�j�E�B2��mజ!���^7
^\��^#�%|5�$S�R���mc�7>�0h���:�K��;aZPl�Ծ�J ������7-��E��1_��y��:��g��H���;�L�f�^�(Z��C�+~��
Z6"$VTn���S��g�
9���λ��e/��V���K Lh<,A���~ӄ��e����g�R���ʛ~���Q�9P�S@'iZ�����M�`��ʗD�#�����QDt�m�kR8G{��g�ȩ��-�$����"z����e5�ݠO�����x̨����t����b��X�ˣ5����@���\��m��_�T��nlIwR|m6�Ǡ`�j�JZ�-��w�E��u�lIU�~���d�C:�9"�������^PUT|N-{���q���X�,���*6g�o9:�tV.\�0�F��c���cK���w/>2��h"�p.Y���X�W�1���s1ϰ�ld�$p�`����Aߠ���*zH��$�ɕs�W�0�s��+ּUV�z�1������_�	e���{�ږ���*���@�yߨ|ժ�2���V~DN����FPH!��*K�����02�&�z�-�F=�sW>��j�GOzn��~>��e�X��M	�b2p/}�ͦ�%x������G��K�3~��'@�$���c�V��B܇��\5Eu��]�����^��ˁ��<�?犭m���p*�n�F�LsN~�Q)ݝo=Fp�_ZV`a_�5���ŏ��m����*(�k�ײ��lP3���<�!�t
�=��$�z&�5R�iy�p�14�]>��4s�|������7^� 		O+Fr���������vį�AX�,9�m�U�~J<̀�}��lrV��I�M�����f���*�r�0�I�fE�$9�-VH�.cܵf� x���)L�|����c�9�ng�E�J��~��`�K����5�ƪ��Q�h:v^w"�9��qB�[�H��?&]%�ְ߸J_� y�G��*��Y�o�#�D��EϬ��'1a�`T_�C�++eR��˓������Z�}	I�&&�W�j�6	��w8�>�:q�=r+^1U�c�a������!{����!n:��b����foah�����M �ʗk�dL>D�C��J�q8�eY3ןvֹ#��(ۊ�ME����Y���֣��#}���j�n�7�ͺ*C�*Y̨&T�7FZ���A�2�i�֊��<�0�\���Z;��͜J]R�t.lb��ڄf��e�:l|�����tK������^��䴋|� ��K�s�ܶ�m2$������J�5�@k��|�@:F:?��KF@o�8�)R�Tm!�c���¢�ז�*��I�ڸ:�(vq����Xv/L`�-��@�݇+�}�ߕ6� 6���r	�LL/`�C9.	�����E���9-��W7�U�I���&�#���[�I����M�r�Xh�ƨ�s���A��r���y$�,;���A�~�PE�;Nu�� ?L�u���`؅~� ��[�.�O��c�?h\�Ȓ���/76�#�Ji�e}�"qH�p��wn��=��R�����'�	*�rq�"�3�T����Յ��1�=E]C!=_�p�K
����)ޣ+,�r���g�~ suMG~�U�'��M��s?�Ih�ϐ��62�u�n�f� �&��Pa}*��S��J�$�'�j!���̌J����W�U���`�tY�@d &;	O�0X��*����xa�G�`*Wg�����.X�>��6��f�Y�β�D2��tM,Ј���e�����5�4x�q6х|��k?���/|O��s���rc���TZp�(�\�J�z�D(Pڶ-�W��v���"���0�_k���w~|
�Z�f�2%������0Dj?����������e�����`kA��͹����z�|E����U��K��7]cl���0ȟksm̷��?@�ZR�e3�?;�{[W�`���TC앃q
{	�����K08�L?�ښ7�wT�'�g�T���T�E����qʠ&6:���2�8"Z�k@}Dg�a��b�G�𙍂]D��T�Ԍ7[�� �t(�\��r���h���ᙲM�\�$Z8����=�!bƙ�t�F%�ツ;¶~�Q�*m5{��w�@ ��) $:KN���{�������!?[CNG{A�/�Se�`Z�Cv���S�JԦp
b���Տ��C9`1Tl�+w��:lěː��t��PYr�%P�#�
��}��t/� =�*���˰;�} !`���\Ӫ�?+ҕ�`������Y�_����O�B&|�z\>{O��xN�����v�T�9t4���"c,N�����)؂-�aBљ0����+��@ד���M���U�Jj�|x:1^�P��Re�� ��r�Q��1��/Tc�-�j~N	��f�W��(1y:�ۓ�uޥU����׆&������|.9�R����\FB��"uU��Կ�H3#��*�L�E�j�8�f� ��k��R�vU�$(C���)��G��:ȕ-���-�e��㐎�i�Ę���J��k�b��[&@��U�\�K�קw�R�}{�͵$\�4r�S��iH5b���:b���@z�w�%Iv<��v	����g����B����a�&죇��s��%��"�������H���sc�~��1;Fi�T��GϹW_K�(�1�A�8_���t�2� m:�m��m?Ҵ@dԷ�mv�
����(���Q-�|�ܫ6��+�l]�O��\�ɘ����⋧1��_���k9�=��7�)�W£ �_>w��j(;b.D�,7�Nźq9К�\�;P׺��C)Ɯ, ^9E&��]��Wm	B�j�S�F��#�M���X�|c�˃<��1�]-�B����;z��s�Z&J��t�JvS羹��M8���V)�io�Nm�b�Q2��$)��6�����(*l���:���9V5���8��oh}�3߱hw��qX���{Ǉ-G�HAW>����^M7oo�A����ZBZ.l�<��P��wW�=�GV�<ok	���iπ�M�{;7�?���I�����B-E��z;�z-^�F���20�N�j^r��R�G�j��3UO"R`�G�>^Y}4�%���I5꽁2���U�dV|������p{�w"pg_iM�1� r�K"�vttS�3p[Ư��Dc	'Q��ѷ�V"&�3`����1<��N�5&��\	�q��9����TLqLn��cR�E�O;�D�y��*��E��B�=�F�w�@��e��^�-�嬒x��q��ڟ�&���_���l�u��-C ��ս��� ��У8'����4�r���J� b���hہ���tN���&K2cF��["�.bx�'�����xE}�uRn���d�|SY=����,���*���e�ٸq���gh�{�ɒ�}��^�Ɯu��2&Ņ���%�Q�i���${-�i�^����,�ǔ��>���T.�&��� Tr�IÕNj}?��o����{���"����R)c����E�߀T��qj�}0���p����z�Z�N+Ϥ�N��n� XZ�x2�)^��/�1�)*��Q]��h�9i���-6�5�׋-��E>!�-۰�;�,�N�5 ��԰�)��6����lGQ_+��������{k}�gё~ #Bh��\�\|�f.ǭ������8!��o�W��?&�V�CuO��~ڡsc(�v��@��P�nU��Ƭ�*$,�Bצ1����Hz�B>��8��H���|D�#�)�j9�u���A���/-�tC�
�,��BBD�h�]����uұRVR"���D�-��L\oo6��|�=Ln��"��J�M)o^$5���*]�X�X��9y�%߮�%��%�'?(�q~��vl??_p�Ko��:���p =@�k��+�Ǭ���)���Œg��g�Ũ�	qW�\����(���u�4*s���ზ yw�=�A2�/)�pXN4sU��7�":��т�)m��_��xѓW�������0'���,��~�(7��X+�� n��Ͽ�W/����S<�rh a YQ�n4���� p�ȫ������`��^Hnc�Cvc�{�@^&��aI��<��{!{�t�6�H�d��́!a�C�<�Ug�b�FY����f`��ub�����i��rA�N]��tl=�_3�JvxWX�������e�YO��U!���5��l����"�X�������#4{"	k��8l��Ե)�)�e���B��S������F��A����.�����謑IP�UY@�����dZB��"��Vͦd��g�+fh�B=�5(�(6�������b�f��ӿ��.��FH�)5�Z�g]�Z�=~EXU��l�$tM��}�_�+4@��4	���1P���~)�o*Ң>^���9oU 8'�n��B1����q���������)�0���̤X/+���&��:Ў�K������
�V�&}-˙�4��`�"��3��=2�J}a�@�Gy:e����.v�Dq�/����A�	�'��J�b�<��w*L�]:� ���!y���;V����X&���A��\�q�׃���p3�����fQQDu��Ը��K���i��u�=*W�$�b�x�͢-x��$?�~N�D��j���5(�P��,�?��r(�������EW�P��}h��D������.L������I��}}���(��.%�4aSU'ȉ��k3'������^��
x��f���b�w�bˌaҰ���2�Γv�����|��\������j��9T�(ay$���� `^]u��2�=\w�C�LkK�i�{��`�����*����.L�����3�R��jO�
=������r��&H��*��>��%�"��6�Y��C�\��q������Ӥ:�8!�2E;�N��0���
��R=�q�Sr��O��K�E�2���S�O�ZV^s��#I|���~��x�M���) EO�@8��wq�lk
��@�'@`5�}�
�����۲w� K�9���m��zBF��#H]�8��Y~$��xx�z��̃��2�6�k3��'��Җ�UjB2=1�H�J��;Xv1�Y�]��Ӑ��OO���4��i��ӆWe��|�٫K�2��˂������Cy9*v���N��D���Xs���GQsJ3��ڵ=�C�����Ŝ�i����������t����ڻ���$� ��vH���a��,U�y�v���M�}�4�"���j�)g�����>��e�AK����J�gy����OR{0�Up�ZDEN�g`+��P-���ǖS�h$&����W��>��0�.(ɡ�}r�*��Gi�Na���saIޛ���Q�}X�LZ�=�6�wD��}Ԧ�F@g�xޘ%��z�
I;�f?�N�U��LH����k��6�`����=u�EZ����Ȓ�Q�����!c�ׄ87�9��-|�>G�Φ2ٸfT_4�x\~T.����]�Ų�;�|z��_9��܇i��X�9�-��6Eb1�v�$& m<�_Y����s��S⁣��*&1��O lRm���`(��r��R;d :A��[����ӣ��FOWNU� �AzN),]�j�4� ~ �o �|tĀ���l�}��J���CE�*�T!`����<କ�Dyﰷ����m� w*{1;�/�,T���	C��f��P����P�:y쐿�ٚ�X,�2*�{`��`٥��
�������.d&���ن�!��s�w	����w\���/]&��<�ִr��zF˪�3綱)����V3�"���7�P�{/�A�6����^��/q��"�Et���� 
U�Ӂ�%p��ԡ���˫�(P�����m��1�4m�} �G�S���c�QǻJOٍf'pk8z�0.,e4\�"Z�0�Q';��G��;�2����������-j����j��h�qQ��5�~�Oқ���r�IS#�{x�F���	!͡�@��v�W�x�K
�pU`�-Z���"������I$�� �W�Q����3AӅ���~ʠ�D�jς���(6��\�nߞ9���C�ˤ��IM�'N(.�܁�T��!�ů{S����٫�OF�3¬�s��C�k���P9����Ok �nf�[�&u����,�>N��Y��C\���
��{!z���M�L=�{ ,[?�CN��wm��yy��w_5A}�UN:z;�[FNgrˇx��6�j�����]�#�ٮ�X�e��Zj�Ւ����<-��K~�(g������rB݈��}�"Ꝑ�z�0���1��~9�Ij���R�%4
QZs~�eҞn�� ΅�f��j��\�)���]4�ΈX�N�D!�zY�䍈��qS۪���Q8�����C�&^�����A�-�qڦ ���}7�~:0����_�������=�e�$�p����!�X~gL];dg.���,O&��?��;'��+��9{����aw�����a���%�I���Eo��s;\� \�T�O���q��wq\���֦�#�3Ԑ<��&(�QX{��x�M�k,CKح��d*VI���9��r�a�� ���#�b�%����9�h����u�{f���ښ�m}��bS\qkUh��D��$�VY��۴qä6��Y a*�g� ����,}���s@�+n�X.���%����a��:ru�7�i� e]���J���wD���)�����Ϸ�zIIQ�󣤮f�W[��D����ML���(��|���|2�i�*>�皻M�T�m���<8�dN ҍ�Z�0y�NX�������ks����|˫-����G�=9���n1���RH��s��w�l�C���m��}ow@jZD�{�#A��u��{B#&()l�������ٿ���2�(�K<]i������`vl�ҸVV�� SPm����&�L���ʹ�f��"e�Y$4)������3�/<�����9�[l`�.������š�澪�)�&o_�>�k����0�F���W������tT�b,ٵ�Pc��M��[�	暤-D�4�;f�'�Ȗ���1�	�[���$]�1w�-vsϨ����[c��oo|�ډ�e&%�T\ڠ�?�\ù�*Ic��m�y*��X�<˼����^��żы�]Q�!����O	�ó�s�9�QR�o:����Cul��,uvb��Ϊ��S���A�革����W�p=��]cf��V���F�|��q��A���)�� ?R�-�����D�h�u�E�'K'
$DU�6J�����]������~8���u
g�^
����������$7_������1�i�g%�fy�s<�n�UH�G>���A��o]�|�m�D=��u>gj�4)#�����P���_l$v�:�}�d��$�����J�qG�����R��uj�����K�LS7�i�kGN����s�!�tH�����Y�^�Ԟ�ٛ�h�����;%�V�m�X��R:Xey���i�ӽ�0T9�T��|�^}���2G�z�V��<�]O>`��D��GO_����(6�f��+���Ao�t��M�~���¡Y�)mz���y�v������6뎛:��/ecTZ��/�=6ye׺ѼR�@���O\�W�gαR�߉R��DS��8����;�v��f5�Z���Z`⥒��m��A����� ��S�ʹ���T)�����,ױˮe��nĈbK�b�N�/ ���y�>��0��ڪ���#ֱ hJ���G끰���\1�<D(��Ԅ'g�v;���|�3]&������ߕe�l��C�א	U��^���0��$\4B0hcN1Y�f�z-R�����o�^x��+���n�W�..�wg�2f7��w��q=��x�B9OߞW7xx/��;l����������FJ�Nn�pH�kN0未%$�ș�и��!h����Ϭ]0Y�����_�2S�SR?m��/	/�̽M��E�"�5�������h r25����oXȲi�c��d~�!����0|��=�ns�.��0�_� �<�wJ��uѸ��-������~�3��q}�X/Ȍ��b�ʹ�.V�h����V٩D��VF	�!��e�_�`��>gK {�?��Ğq�����.>��������3��At�@>E�t�:�$X�<Y��5k��oO��O�
�+���|�_��B��nrf*��p��^dG���Uy���+��e1䋢���~�w��Q���0��m��JC��n̹ׅด�H�@>?�h��]�>�e.��K�������V�c%���O9��x+'��u�w^���!Vk�5Ѻț5��\�6gP���(���0���Y�g�sv2���!q.�Dh��u�P�?�D��S�����a�q�ɻ銻�����T �Yo�;��]�l�)Pq
���-��	T��L)/�&e�������9poc��)���(�C!�ߞq/J#%�Q<o%?
�Y�+}wSN
���-�D����!t��\-�uaU���&��(�vVF��@��~ҁKW��~A�`,tb�*?���:����4F�彩�0yU:�
�ت\�n��e��Q� ��G�e/������)���E|�()�@>���H
2�ٰ��)�����Q�>�%_�]��}�M���>��.t�ڲ�R�62���
H�k�2O3�An�������z��؇d8���t����U�"��9{�x�*��_5r(��K���ֵ�r�S4�9��5�vC��}�[�����A���!7�����iOڎ.���g��K��ѐݣՙ�3����v��m��ڹ��'$��&��=�Ov|Q3W�^Ԉ��qrۚm)�|^�m����'�o��g4K���I��<J�h)�0��dp&��Ѐ�9���e��i���/"h�=��Y���,��y���T�1 ��69m9�oZ�S}d��tKLb���9��J�H��m���dߎb��هr��>D3��|�z�]v��y��S`C�"���s����Ӂ�U�;E+sP��S)�����0��8L�}ϴ�,��ݲe��N�WcY���=Ⱥ���֪��)�\�j�1�%k�� �A�y�4�Vo�_�����41J��'_,�W-F���x3�{�B0u�f�Hճ|��梛H�<G�yfB"��i�Rd�ꊅb	�6��9!݇��N�Θ�eM��*�G�JDo(`R���h�zv��� &�U���84+�~ߴ���Bj�>R��yD�I)�uf`d1&J����=5Z���@"���^)bPT{��Y������+���Y]9�\��B�pj=޷M���M�4�[�6�;�L�+E1 1l��Ɓ�2h�c�Ph�t瘁ãu㐔�·���Dr�?Q����	P5��;{���{�p6�kuB�������N`�F&; �Yܲqݒ|t=a\mw.[��">���[&�������qAr9����Ҹ�y�K6�_�T�`@(1�F���	�#��sl����yY��˽���Ȝ��l�&��}��L�-��;T�_�7=٨�B�!��7���� �a�d��2H��<N��c?�9S�(+'V�^NdUL�2���ɚ[�)�Ya���&�Nh Y�PA|?8����CY�lh��I¬S����{L��
j(�B�b�o���ߺ�<��\��v��?o~��o
١���G{�N%�����W�WA��������7��f��h?�4-vխC�$����h������B�y�R����R1�'�-Ԧ�J��g��Ζ�yl��x�����\��yj�����Y�5�>5�!G�IW����-y&N�ZK^��4��ɇp��N�1�vo�n�P�_\�cFS%�9�p�S<��!t�k�@Do����h.�pFx�i��7���k��O�nP��?�!�B9�����7>��{�l���:Q�v�H��c�B���k@QY�ɑ������9��;���P��/I�NC�8�P@�a!N�Yݿ:���oiF4��5���({�V�P��?l�Coy�2rm%<���鍄��jjo�a�p������_E�5��j�;dy�[?���7��n�m�%��D�
���D'�p5�ȍ ,��x�7҂"Y8���$�R�$�D�o�,5�H �+nN���t�$�~�x0�G:�uR�~)���<��4��
���hP�ʅV���3�&��$�a�r��e-���z���;2�w���`��*��4�uv4D�b�Ŭ�VS��)����4L��e�J�x,�Xcآm�"__��r#�����(�b�$��:�W�o�wȖW��)b{�؞���ޡ��k����X�9WJ-M
J��C�}�u���5�^\;F�rP79a�,��M��g��9���r1�~��|>��P���z��)9��B�4�g�良羕���_���8�\������"�-k:dY�������_H\�����M��J~l��Uf�����L���x7�B9[[0
�.���B��y���l<1���(�cYF�4���c�`��^�/��w�mJ��[:64^b*\>����+b��=��u��dn��%�쐑�g����>��m�C�8Y�1��88ws�O/���O��p�nxg2�ύ�x,2�$c/�:����hܗ�T���!g��M�:��
�}��Ɓi�=���Y96B� `�s�۷�[&�s��`�!��<)3/Z�λ�^oE��ġBb=Cz���*pp�k[]�Q����.̵c�}_\%φK�%F��/QxLDD9�$��-X6�n��U�K�5ݗD��o��^��?nъ�D�pN">�\���%U\bDğ�%������1d�p��-��u�𿔐h��{v��z�;��Qi�k�c��m�8G{=�7wQr.ж}�Tgj}N��Q��9OM�=%S�n�
�\]�$� �mպPYUoV#)1﹖ޛg��
�l_@{��9�_{��i�u��9��;Oͻ���p�9�$ʾu;�o�/��5{| �ؙ�r(���o�sg�a���G%��K�@�̏���Y@?���������Yr	D��'9��Ųo�E�
7�!��4$Z�թE�N�K�B�i5jXΎ�)q*C?�� �����2�\_w�4���b����q�.j0�&�QxF>!���j���U�$���Џ@d&�;�IEA�~M#M��Ȭ�H�zK�y��	����s�-BHy�!e7��k�RT���ۯ[M���4exOH�>x���P��%[38�����7p�H��&}s��= ����v�R��Ib�f�?���*����a��V�}����u*������R��Z�T �Z�۽�����gHM��}"�<���w�H������}ƍ�%6�V�s�4�}����Jd=)u1Lf@�̖E�Y�=QPak�jX�K��ug��i�{�ǘ�shK�\�FĠ�d)q0��t�`۽��<Ǜ'-�\kύ�{�!��^̻Q9!*fو�M�dt��5��`t�-�9:$� �|:��?D���C�@�
����!�\Ax����O7ԅ�������Y�!W*��]��/F�K��j�%�e��N�����m�i1IKu�<a�v.c�kL����h�mK���R����Pt>@5.}H��gdӪE��0�p/:8!���n�9H�	=�]� �a����R�TO����#<vkqQd�A�)���ϩ�xz�յ��f���򘑞��j��Ƨ�j�DS9j%~���k�w�D]Yr�S�ml��jںFO��N'�U=Zy�O;�����\$��sr͖2���}����+����)6̿��9;��;�]vF��˚� �BUl)|_箷���(,��a�y�c���<'m�1}Z����T����;0��7T��#�I(W*�����Ms	:�z4��Z�^1]x��ʪ$�p6z�y�W<N��'��>!:��7����r�`
.wL+�9I0��qj f�EP�-Z��PZ�$n��z]�!UwF��-����Ĵ��	!�ާ���a�bv�]c�u<��x4�k}��=w�h��	@���6��@b"�*�,����+��W��En/1~�
��
h�,u�誯�Xqr�6�L8zpd��;�"AH^m�,����,�6�Z��Q��j�ᒞ�89�B�`bi�0�
���C�,�0��R��������������{��;$�IX�w|�c�KiG���{y=w�=��ᝁ���pٲ��<�e [��twbߞ-�h��0�{�йr�a3��b][�BiS�2kL����р�LwK�����x��ǖ��髐k�������0)`m��(�m7�����+�,,_a,�3` �.�4[��/����3�oo���]qą�����s�n������Լ <���:@�ߒenB;P.�=Z�)�{�`��Hm�X�X���f�F?r��B�0
��m�u�4
-�=�?;Ϟ\l��=�L�-�Z��}�C;�B��b=�;n��v��a M��RX�����w�:��v�Thi��}���1��[y$E��LP97rDk��X*hի��M��8�x�k��s��J�&l���t��@��f���a&���X�Y�ȴP
+��Y�8�*�CX��3]x�߽�LA��mۼl�x�T�������퇪����.oe�pҪ�r��-��U�G:&Ê~�2����:�9�_Z2C��ZW�M{�d�����#���9�<��\��AFL+e��i<~�<�����2rHaY�h�/�^�u���kP��Y�i����S��)3�&7�!٫k���oA���M"�)2�6�6���41��f��!3�f�~�YG8�;
����6�BI����-�D�|�LG�E�i��"]��|64;S�I���+�+�;&�o�oO�� ±D�i�^b^xaU�9m$ISq�z.�^��j�W��H�K�(�N�O�%eoŘ��3�NJ��pp6ȫ�f��7�]@��𻊓l*�^;�X4l[�Kugal�z��^�IǷt������omqHO�U�н?���
ht�fl���gtcy��K�4���z�?@\�g�cl�!3h0�Jq�Y���A��(1F�q�m�Ԓ_Sl�V������)H��x;	�~��_ֿ#&��7�^Ąsn�Jv��v?3E�w�l�˜�k�H!��ꮳ�»d`�B�o�~���r��i`:d�\���Y�Ʉ> �f�Hq�[-W|�@:���t�M�M��}��EΑC��Pg Ti8���m�zѤ�g�X�n\��V�`
�uq����U�}� [IM�5���F.�?Xϓi�2��K)n!f�[4�@�N����y��!��n�X��.�&��)PP�D壘��<���|[����{T���{cy��,�j��.�������m��G`<ˀ�G�֠u�'U��0Pդ�a����u(ngFo�T$���6x�
C�-d<r�O}͠����E�Mз�N����=�c*��]Iy�!��\�`��]����L���5�L��W°e�[�y�iQn��uFdR����	�p���z��`=!����[����q��}��ک�>��EQ*o=�"���'*Vő|�p�O��R��^��P�����9�Cɭf9���?RP�GP5��N���Y�	�:V���i�7ԡ�����L�5yV��R�aq�����(^QI�u��'"��qρE�%�� ��A�iX�v��a,�:���o���v�(_���#�w����+'���EReh�ހ����.Ӂ?>êħ��9fQ��dSe�p���T���kxޟ�; ���fz��WD9k�GXj<���uo�
�b�l�]*G���y�6��S~"��פ����|�i0�p�1�A[f��ٖ�|�6��ԸoA7��c^fj,�h��2�d(�7&���J�d���6�c�!]��{���[�Fs��U���1��H?�M�=�nRF��1�P4�-n0h�Q�~lĎz�1�S��fG�N����*��h�..2�����Ɓ�Ir�9�A�e��B�1����4�b�ߵ�G�0�h<܀K���P�*�jG�D�`�b�[l�`{L��1�v�1��u�4�;� =��m�2F�u����\�j�s�D���\��0��W����m��!��4�-'�3]���<*�ҙ��AL��:`�|sY� +!VF��;Hxe�A�}`3����]H� ��P���m�g2��Irb�M�WFse'TL��e��+ܜQ�a=��P:�PϐJsչ*��еmIY"�	l�1��J�ղ��D��815�r�����a>oG�|�Y���G1�HMҧ�|�)�ӳ`�@20��۾��-�<ͽ�Ӫ�b��,�@@�?��Ӝ���$<!�yc&o�)/^�7�gʋ�[�L�m���W�����M��h
V�@�)%t��w����QS�!�$EK~���Y�O@��Ŀ�!��7�
412�Rф����9-�(�VU ��˺��tՖ>�
�&���qkUM���w<�QU:AhyϯW�k��hx��Vgp�ܷ��~)A�B����u��)�� s互�?��W�-���C6���MoY��P�\���	[`�E8���,8�~�ں��x��}��.r��~;�[Y���J�rmX��U1���:~r'��FSϬ����� �H��/�;}|;��5�8�KS~���!Pސ� �f����T%�ęDߊ�y7&�ו'���:0$��
u������t��Ϛ�HuA͖��N���~�B��8�R�w��̈́�ɫ'���EX��N�ɤ:�,u{��nH�����ef�����E7T���;Tb��=HwM%t�z�>�U�.P��cF�iA�t惚#qUX��PVy�"����]��I�/� �b0R�:��S����(�z������j��<v�.�|��9��U38I��]����?���y��
���?��o�c���P�\D�ǔJ��h�O�@�N�.-����1@��z���s�/�<�~)_}�Y蓋����C%m	����@�4��~i�o����i�����h*rN���{��+7Mg��<����ƛ�F-�d�+��Jc�9z-���5b+��P��"����b\�=n|$��B��e`䜊��4�X
�r���D����U�#���L��Hn(�D~��?/4�SR�w
�	���X�Y"����)c���;G'<��	�������q�l�eeq�wJQ��ȳ���6�?�y�ǩjZ���N���E�b=�)gb�0�21ÃUuy_a���&�~}���Ul����$�Dr��}���|��<�O\�]9�ͻa�Mh'��x�K�>Eff�����X��?�P�9�:�l�1�2��U�I)`_�,�%�dZ�	�d:0�&���1E��hx�|�~�u��������n�g�H-�������?��Q�z���6�`5-,��s ���$��1�{J����sPn[=�l�`��[`��9�HB�et-�L9�ʷ�vzV���/�����~����ٗ��*TY�������~���i�h_\-PGC�F%U���
T�5����v��t��Lԣ{<5�D��#�?�Nn��3K�X��3�[Q#<���!�+���~W�Ŧ�0��WKV��!������Y�'�rK�U4���q�gfm<	`�ij�jl"[t��v��OZ-P�؁�����H�xO����3��dq��-RQ�f�2��Gp&������ToQ{�d�T��;����D;cn���;޹�-EOZL�����7��ȗ=�ޟ�r4���\��EB^;ti_�o���h.9`��,����6���Y��骛��	VV�HZUD&-��{��� ć�>=��B����e�T	�O��ӆԙf܇6�#�W+��vٌ��O_f���e�>*sl]z�ѡ U�m$X���cP$��-�����x0�^d�L����ل��Xk2|����gX#]�G_BkB����U���p��	�_Ć�sZ���c�V�w�s�-�Qw�����Q�������Ռ��!ox���
<DҥVf�3h�]a���2�Ϳ�(�#ͺ����i��tjE-��%��Է��Gr�_�99d�<4��2>;E|�d�G��=;�HϪ�oQes���v��D�:���6���g���3%x���p	�؊������-y���qa��{�_"�������~�'�bC���,29~MYε�DA��o��ag9�.�X(f� 4/��v&P��%��{��zD���^U�bk��_�M��Љ]�"M�Cυ���.|�F���������ꙍT�B�o}�p�Λ�~��d��ʹv߇������� Q�(�H�;QD���U���W�T�Z��F�-�up����R���J8o	�?y�!�T�|G��D;���u����,ѓ<���xA� �t�*j�O�F1R/�"��5�#pٹH0�˿�#vē�͑m�ܕ#����!g�D��#w�oxKb�WV�G*���-�I{F�6�~	+�b���oʖ�k�7���>J���d ���q���i�?=�!����Wp����i"bA������S�6����� m�Q��CĬ�cp��&7�E�����ƅ�c�����	s��;���h�E
��@6�Tp8�ٻT �
O�J�,���M��_�
��Q��/xIN	;��})�S��`H1���3�3���h�8��K7��F���xqk�j�򌦇���1F��?�����ñiӖ��U"�����_"I���N@T�Y��E�R�,��c5�m��b��h9�%���Vŭ돧�;!�5���}�s�������O�#F��?A���SR)�k���Kߌ� ��46>\������h,���:?�O#沈��p'�g�F���*v�cm�<�!8�9;��bj�>5������Nڒ:��"��E	��K�A���D���yd��R2Uy͕|��t������R�qB�G�V<;9ZO����p�7@y	 ����>5n�R?Ƒ��$r(��	G
֧��k 4����\Ohy�#�ѭ�_��M[$���RW�2_�Ð(f�O����zT#,��[��{��?���h��$��*��|gn�<��A/s\3�(=�K&�J�C�X�}��-�I�8�b��Ѿ&<���[����O�*��S�.�]�Ţz��gXޛ�Zoo�����r�b�;1f8�+��\�|�M����]�D�˜߷��$j����s�!&��i�7iKZ���fwW�9R	�"f��I�x+�����ɡ��+SXF�vzZ��@_�b�;&cE�B����quŔ���w��̗�M?�Yo����c� ���zU2���(��p̀���2��h"��5���:�)Tsh�	�.��zOg�3>�/(��@K��T�
QT���@PG]i��~��aP:,c�`_|�q��lf=+2C�͖U�:��W�\��9��n���<��_"7
Be��ݛy5l7 ��!��)�����Y���wD�*>�D�D�Vr4i���\8w�}r��Z�;j ��aE<�:
��L�nM:���I��y���٦���w�F��ۚ���=��N��Gƌ;=Q�`�������#��;��A"Kas9�XPf�u�:#gL.���2�p��WL�4���k#i�u�\����=K��.J ��zOk@�p�i�]���aXY�e�fb�����K�C�{Ẕ9Wf5L�Sp�K��$���U���ŉ�}�8%������tSCa�V�T����,Qn%s"s�R�ȡ���/"˴W�{73$�b���.*�Kn�h�=�?�<�����L���dYK��
���R��~;�\, �����71��F���H�bK����^�\b ���0����I��r�f��Dݺ@��@���8|�YW�y���^������،���C�jZ��=�3�j>�{=S�t[fs=c]�
���[��z$!`~şg�),��A�H������%V����m@����RP���f�W��$���[��5C6�ƦRA���_zF!�c$��J2�q��V2��D��S]�%���oh^E./��ja�(co���k��	ܷ�@��J}~l���.b������Ü�Ry�5b�A�\?��\�/���@XbS� 3�^0Ի�.���Ȉ�d�s��V>�.��ʜZl}�J3������p(�W>#�O��i�t�\��v�q�n#��5_\���
<ErJ�$J���}Q]�[�5{L�:K/Ȱ���S���~��{Lّ��ނ�m�YO�=��`-: \\�y����LBNՑfm�v��� �;&�`���Ji���q��|E�BY�' �Jzu&?,��;.2��w������RH��N�;�4��� �`��(�����c~3��fq&�{�B�MX]3��N{S�����w��Y尚�(*�|T�R:$4��Ư靶,躌%�ۤ-n���θK&4E'τ�n.$i�M��&��+�D_�4��uG5�l��f���c���'g��ě��lVBњyX����Mj��9�
� ���g��A������=3Pu�mu��v�DE��i�PN�p���W��g6�K_7�f�/e͵x�:�~�=��,xjG|K�[u`�=&\O�K�����	�����]T�g&�������0��/5_�n���K�EB���/������qi�����W}FLo��6�}�ClL��U�ϩ��e���:U�:(�)�Z5i����-.���imHz�X��r�����.Y��hk�t�#�R�^~shV��ҹ�TR[���7�x?@�Y���=�U}���^�$��?��[ `ֆJ��E�?4��`b�t+D�yC 8�_$60���r����n;,�|�����t<Ќw�Y%���?������33��
F+��&�6�7uB5*�y&o�J��a>a��l��d�� ���VrE�$�,���;� �|�.ڇT4��P~�5����.ӹ�)i"�g�q̠@�;�%�5#����`��/�������9Ė�z�� �K*�-s�jⶻq/��k �2����c%`<�U�ืK��1!t�?3�]�-��<M3:�)Z�q�F�UK͖~z9�;ي ;Y8m�P��bD[�����Pd"+�5�12�.�3���/0Y²S=��bƎ�x�u�k8���)A[:A��}��	��*���i��NQqm>"�?h��z7,��'J
��;
��E��$�\W,��-2�d]����\= �j�[,(�E���&�M�WI]="DDn8�AMC��p�V�J���9��q�A#�v�r��M��=�����sQ�{d�����<&�Jt�YF}�"lcs�n:�:9Y;A���L����8MaeoS��s����W�B)��M��~���������p#�p�TY��v�(R$��7�@.~�������>�'g^�% LD8�"8��ny3��x�(ZÊ��W�a�iˢ��4(pK�ȼʿ	0�W���9�Ҥ�6�L7������	�I%a����p_B�X>Hjk�ҧ}���f����9beK��t�t�+�W�R�sؖ���=gT��5+Y5(ݵL�51BN��A��3jGI����?G��d[ڝV�@Y~�S�/i����I7,FF���i��]���l������fSz><75���4>C{%�;%�6�=�\*l�A�(n<��ȃ~�N��a�]���@�|�R��tj�\�ڲ&���@�ί���7���(�t����W�C�3����=ϼε��1�2Ut&0�GЮ?Y����x��܊����Y�;��[z[��[�#ߎ�������/��
w<� UA'��N�2��m���U5��l�_��ӏuO�����Z�fu�'����PA���������������Y�w9���>�k��T޻�����#>>��R#w�V�@��v��C�����.Nl����V�x��1�_��𑏐�4�g��2O$+�q��5x�Q���8B� ��!7M�|���y�*�MXܡ�������Մ%f�ڗT�	�I,��ee����`̽x�ǦC~h��WV�C%ð3��@�e3���)�p��G��mY�P#���I��*��N?�������M�����W�oz��h�ncE�S&/|C��T��� 5TW��)
%�:��o&Wѣ�3q�Pq�n#����Q� g�g~�=��BK)��fc�*0���2k/���0��%`J-Ƹ��6~�����?�&�������>=���8{{c���O"�_��V�.���I�T?ܰ.꾊A�OHB��/�c�n ����{��G���%�'zݎ�r��F]��T;Xv�%*ԏKB��rAH�n�fsY���@
@¨�����_�e�0�%���G4�!������i3�Ψ�ʖ�8��B�Ֆ@�\=Qf
g��C�`dė�巅���J ��Q�D����+��+a����\2�1�_��ӂA���:��nQ�0�L�X�&�p����s������fb��-2�L19([���d�q���L|=Z1(�_5�RŌ�����<;��׍��UhNv��Y����%�}��u��T�$�z*|�z��!�K�u���s�,�W��OGJ�3��;��;�o|O�rFUNN�M�>2h�K.�"��lE�PM��#�\��o�&�����ľ���{��	�	z�۬��w��B4K1��Т���zh�>�K֌h}��3v_��� U�)A{W��� ]�2 tR�>0�6��h؀�ٔg���J0<A:�D����(��,n�9�v I&:֜���%GY(=����ϢD~�����>ũd�o�}4�
SY�][��m�HTW|���ɀ2���ɵ�ov\�E�{���}l�����y���5�[�K���>>�δ�0*$Rϻ��FX>�*��hF�G�wXmx��&��P`={�0��o8:�ma���ϸ6N�YD�����f�p��q������:���`��خ�v�������#0B' I�ui0PL�Ǆt� T�7�ki�Jm�ˁ�&sER&z��?\4W����רhu�X
i嵖|�N} ^M�G݊�^OP�&�׎(ixY�욙�9"j��!���t�u)6�Ln�����?-'5fD}D^�p�������νSҲ^�4��v�o�%��VH�M�E���B4�8��a�W� ��Zu�ų�-��3uB%ɡR�_�@�&nG�mQU�G\=�ErZAc{�lE�<��aL�MB;W;-<�$�?!pP%T[�����90|4$��wۣ�Z�$�~xzO�>�n}��{��79(��ǆ�rL-|���B�G����M��DfH�'[�2�H����4V���|7��E��g��$Q_&��lʄp^���h�.0���KFxfp聏��|�	.o�t��	l��p}F��v�mD��X";��5O�):�vR�8{�imſٌS .�m�s|0b�(� f�ߓ��8�W�~���<`J����I��_�����ﵨ����B�����1��@�r`hLr�0�Ą���T�&�
�PkiY޷ț���eP)&KY͵M��mFrA�&�|��heM�-	@��OG	h�%3�0̔m
7����0Υ6Y���fb��K�����_��p�z@`�ǰ������]	M&Y�O"��=�e��)p������<F��^��?־]$D�P}��@�E�/�b�J	Z���� �<�'��ґ�i��`"U�9�8��P�!�v�H0q��J@��p�ȕ�� }��C�i�3r�8_[
-1��8%�E�N�`�����!b��糭Ba�`rB��*�#�^���q����,pI'�'└�'ӳc�ض�<��.��I��~G�l�a����v���ܼ��c��j�!���yvй²�?ZL� ���EJț�H�7Hܬ@nͧ*��1 �(�>���^Κ)|�'l��T�Ȑ��Cu�����k�\�i��ށ��5<9�^n��0Ͷ�;� �\�Q��U!d.��K�������?�KK	0��h��/�ރ �m?f��K�Q���~6�=j�7�K���$M}��뵰�E��q$����U�D"v�����dԩ"���&�wIhns�sA�3�qЗ�b��4��3�\v�f��e	��JP���O4�L���K�Mc-Y 7� �|F�vAxeM6x���4��r���-f]C_[U�"�)��*�$���G�F�|�֥�$��m�'>\3 I��T+���9�t
L0%����;���S.̓�:;R�խT�h:��j�A�'l�j��JV`:�$oCJ�_��� *� p�`�͊q��Dr��h�C�vۢT����Z��#�I9��y"����	�N�ᓁ��w8M�k�Np��l�8��l��~�b��qM����B��]f��V�Q{A��f��6o�2���_�5g�sE����$[l��#������諍�&���6�\��e��Ʉԟ��7ʩ��*B ���G)�:���d�ff�Q/^�i��cdZ��S�� ��  ��c�JK�2E�7ը��3�4_[���B,Avn���n�J�JU��=I\a�=g��rjǑ?Q^��z�1��Ĳ��{Z���|�R�᜖Z�_�4ԡ�d�bN{@�����m+rx��#yp��� KD��u.'��^S?"��X���p����&��Sc
bg�X�q���m��r��e0���c,���;'.ʷ�^�u���Gp
�D���j3�|��|^�E�e�Y�}|	�=tX�oY��V<�3 $�Cw�Y���@������5
�i���*&��)�_�̦��v���M�_SW�%��Q��� }M�*�����r�J��[�W~�/UO\du��bԔ������Ӡ���P�n�Џ4��Q���0R_�$ =F�"U�1*c��s0VA7�I�Z�]q��t�1e���l��LJ�3�!�~~4S톐�J�Sbp�bTPLdx��<mzn:���h��<�����@_^=�ӂ;>_�T�:��Q���m�,���Ze�\XӤRiO0�.����k��w���p�kcK�o�W�6W��붶,�?Y螂0�@���;/�ng�ɵ��e��{W5އ;�k��Щ�ۛ�?��>�Q��X|�Aa�ͧ���4ь�������ɍѪ"��?�h%��t8�8�Β ��qi��\�K���Y)�����%
u1D=�%�ލ|΢S�I�8S��%I��|��lҒ� ��+��S�;��%|�� �O,�C�	�׻�}��&��M+�6��!+~�k���!	b=�=��B�dbT�H���Կb�����(��g7����J�H6@��0��x�"W�Dz����~�e�-�gS>��Iq��[��3�ubts?�[)m��t)�L���/�,w[��s�=��3>�,�Ӑ��&� �a�E��7J�Ջ���-�p�cMF0������T���?���p۱��鷳i��r2�^�M�߻ݻ��@aCw�s�#˱
e��8p1���B8V�a)�/�I��e|� ��O�C?�a�`�d_(N7`P�O[2 rT�&�m�K��'���m^!�h7�o��F ��C\��E�>��M3��o���C�[���� :���;R���ڪ�<�Ŵ}�D���d.��an����^���"�3�!��܍IH��n�.����Z�ga8?f���h�u���_h@8��u�.~�-�X�LfX�`�!�S�R?�ё��m���!�����J�
T��	��K�o��T��(3�|�I�N��
�5�"P4i�i�{Ğ/' � ܨxհ��ZJE�o��0��F���1�����H]��9��b�b��Hzr�����C�
c;~��)r�Ա>����7��,��S�(rRP�Ak�P�L+�}R�^T��~�e!����t,8E\oH��x���}Pb$n�U�.Pկl��D�R���#�'����b9:��&=���_��
�DZA�JS.O�`�F��N�?���'��X�����4+�p�h��3�����l����1Ow"� ����h���I���`���7����3%E�k�\��U�]�q�~i�c�㸕�|�B���?������t�W������/X)���OЈ�l���'�3�Yk5��u'CN���J��@ ���L[�{�%#\
���{X��ϞR���z_V-��3��}([j��i��	����Y�'!��PT�7�(����;)�^�r��0�D��A���m�!V�U�9�/t�_� �ș�ϖ����Xd ����b.�gm�,v��/�k�"Q�ѡ�L .��c���L��p	ь�\=���	�'aF]ģ$ �S:,W������6��vv5����B�0��æa_�bh����O$z��W�њw o���������o��:kX��������5x���w�b������n�� v-�f����;1�|d�XyGdL~�ʱ��ˋ��0��^a�xO6��w9j7C�x�y��P�=(�#S���oW�U������~ Z��r�����x��ictO `9<�)���'9�/:���.6��d�Xyp�G�i¼�,�r�n�TF_�g��Ǣ�;x�Q,��mzSH���`X�Sծ����?�x*�&\`D��ajf��n ��r�e�������7T�ݢN.^~�Vطj�SK0��h|{�����
?�cY%-2��d�<�/=�K]G_�%��Q�,���x��l��j�=�c��?��g�2>&rx!x���)�Z6�9�X���H5y"���q}����Ϭ�Z+�����o?���U/�ӾE�'wϛs��N��B�tX
�êE!5E5V�� �;���7�X",�& ������Q��|"� �э�'ml̫C�
&��e~�&�rU#�s�Y��M�e��(1��Q��C���?4�r�[� ��/�ш��Վ�?�it������*�5�*D�;~-�p�\
`jK? ��Zg79���Eg��Fa�	��b��}LIW��k���j0��(Š����5��~w�7n$���ķ֜	�!%g�Գ�&�.�C�1v[6�"؄�C���R�9��b-�Ex6�y1���0r���A�
��N���b��k�x��8کSa�'y�d���'�ě�>%�*Z��Hݏ����)@ns�UM���|�S����Y�,�j����0k+h��燦��D��(@��hb�E�x˲�W�"��+Gz�2�.��Jh�8�w�^���u:�o�W�
+q�{���y���ec�,�����S- o��21K�9B<B�0�@���<S�֒�pv7�<�p��Ғ�vm��x���?td���ϴ.+��A�A�����7P�� ��D==�T�䠉כ��N�6H���u,��＝ı����Ce�� C�Z�{?�-we��R��#/��r"�4ZS��E�~5 �w<�w )L�#X&����'40��`��oa���5U�Z���`���@�?�e��e x0��� �K[p/���{�k�23�p^�G]kճ=��TJYH�sQ��!0�U^���
:}���:7��Tا��}Z��W�-'���b�q��i��{��6��a��<�q�K))�x�ǚ�uZd��ؑ�u,,ք��`���v��J�,��� �I�P�8S	��$��I�h��$@L-���#�5����`���J��?�L�
rPmY�u��]aKSS�Ҽ�Ƃ���4S��[3�?��|������2GS�{����hD
c��'��=�
����`�F�S
Gќ ��;E�k��2�HGX��XO23Xc���\F]y��GB
W���4�镌+�8L����Rj����Z;NJ��tLV��'W��ȇ)i?[c����%4�oM	�́���L�58��C��'X/Z����&�0�$)�|H�-Ǝ���~Xz���ܕ�τӲ^׆;4��v��'��%�-�y!=��5����_���9m�����h>�e�Pv�;	µ^���{��M�����á���{��o"e���|=��U�(Z��uGB,RJMַ�S��	Vg�"�5�,�g�0[G@'m�g	�"��J+���,��ŨE�k4_��}ٔ3�ޔ���2Ɔ�@N<W���p��w'qh��fޏ9z�� �������{
�a3��g�u*�79���s��̂�;
s�
 ��v�����~��m�&��%z�1��q����EP.�1ߌ����C���"�ɨ��!=(��tO�p=��-��[�T�a&v�x�����Xg?v�/���%ҹQ������>*Fx�������-'����:�kܹ�?�۷�~�-k���ߠh5&��;�ZpQ�b!-\���q_��[$aW�\EHS~�Ef����j{���9c��6������'-ׇ"�~U-�������q+��K����m��W9��^A�x�,$+�m�F�<+6����|�{�\�:��RQڂ,	G��&q��a=��xܬN[���aw����xL��
�ɱ�X�=֤v������H����(���������w�� �|����%�w�?r�_�l92^2����bF8�B�&�(+)қE��#E@7e�O*q��$[���}���5�@
+���1Ku�{� o���.D�|
I
l,���t��k3��k����(B��Bpgm/I�s�|ld�\ݙ�,8��ME�&�h�H-F���HVN&>�-	���:�E6���D-�{���-X�����Ym��#��j��iΒ��)�zH�ⱉ���;ͷ�,i�(j��B�mI�!�J��T���	U.'�U]�g�wGZl�	���>�ɇ�^j��$��(]n;���nڒT�D�86�4O9�3�~z
p�z������+n�/Z&�	~�+���� D�� Ղ?]���vG-O�҈E���i2�}��+���Y4#�
Wz��w'�Z��C�G%�a8��>�}w��7O ���f�/:s$��@���V���*6���֣۸װ��*z��Z���\���R�ߤL�#�So»E�T>�!��T̎	���x��g�9����lsӉ}��,��<} �!��ۿ�����Jf���u����;k��Z����F�T\��l���bJ��%6D[������s*g�Y�y�Æ��-��\@�y�?ܗD��SRz�Q=��F��
�P	pt��\|�k����$��`��i�����[�����F&�W�,���Ƌ�J��ߕg�m����7��"FV+�v�{A��ئ�8^v�㬃�J��IND��L�s��i��c�n����D�t�,-���sY�Q}�M��\�d�c�ݑ����J,�@�Rmk�r��N��j���\B��h"~$<�����5�z��z�oA;'s2:�:�֬���tL;�G�]�p��=��K�-�z>�5d|��ʣ�=F ?<h;0�a?J��fϿ[��8? ��e��L�"��nb�.���$�;��y�}D}̆����>gX�g0}<NmR�ޮQR��c��^����'�в<�SY�� ���@}�|G�	%?��ir/��0�]2���F���(4a�0��G��Z0i�|���& d��8O���ݮ��g���L�J�-lQ�kb�B�$�G��r@uOMp��N>eP�~d�����*E��H��!.T{�� ��"&�Ȏ6bQ���4������)vtuBش�ɑ����E�C:�5��<�+Qm�r�(�}�xԜ�*��U���F�o�*���z̧�4[��MD�p�T��m�\j��={�,�1�" �@��`#�Eo��R�4�5��Z]��P��.�~M�MֆITRܮh�\���)���w��H��M0�py���%,�'�.bn�-ZX��.,l
K���lg�)��O�9aĈ�C@-Ia���S�(�&D���h|)Ю�a;�ڲ�/�ų2.�m�mQ�:��"YDmҢ7EAs5���� ��N2Q���!�Kd�_h����;��3E�f�!�h3Çq���B�e����,��0�K[!�3��������,��+�c������k~=����X�HQ��z��Z&L�i�_x�7%��Ίݑ��P�"??��`��p�N�!���%�.nA���T�8�]�9��yχ���8|`J
b�R�7V�Cs�j��|y6_�:�]�|��/J۱')t��?�� 0+�kzJER�̸�:�.j�ؗ!�z�	��0s�:'i�$���|=�TDx�(�D��9�����&Tk!3�lʷ�}?E�cL��d��7���%�R,h�c��%c6E1�|"�xO^�X��S�|����F���-Z�H;0�u��)�z�e��� ���E�f�T�)R`��!O`��QO$�^u�2�p$���l�C,lf�]8q�<|d 4g���g1���}+��D�{et�9o2�����6�dS,����i�7��wq�[���Vr�6WO)�s�à�0\��qe��\�]��W��Rɉ���Oq��w>y�=�W6��e't�	��ʈ^�Hph��@滽��]
���VC����)�)�FZ;����|y�)H����c�܋�Ty{ d�N̯p����ize��)�h�c= I�v��u�'�u��^W�v��Trd�Kk:��ș1%��Ms��E:��$�o�"dTYo�G�2�dB鐪�ݻ�B���� � 2շt�
��P,���~��V���~����lf��9�)�!�O���;�z�0o�k��{Ð�+g@�:�������[�{wM�H��K����ٺ�k��Yͮ*46^jI��w�
��F��3��X���_덆��1��]^�TqN8tT�^j�r����^q*�S.���g�V��{p��"YkT$�f���5`����Nvcjӌ� :��]�]��<��	����(u�u�m�;���o�$�4ۊ�0������r�{�ت�����@����6E������x[Ѥ��Z�%E�B�w�Ō56��Θ��O����Ry���"�w��r�;��5��:��\��>�jK�bwu��f9�f��1���'�w��j�i��8�t���e�;	���H(�u�ތ�M���P�5]ܧI���i]e6��t�9@(C==�e0����wkt�Ga���V�ܐR����Pw+�a�[�� t��Ȳ�Ъ�Av*��� ��_2�~�ٕB.���q��gLC�9N�[L0H��ڻHI��$��0kp�lIf���O^��bs�����<é�_�W)S�Io(V�T}��²Iʽx��|��jCQ��\���*j��$+�tg�������Z7�A�
d��� �
H�@��
�򮹐���o����.ˡNǊ�v������a���v	���&�a�M�n�u<Z��������{���&������2@�z4�:��&���khwՌ�K0Ӟ��j��l��l�_Y����*�hw˚'A�]�v�C3�9�[��� ����|�w��'��,��ϕ��B[����p�0TG~������w�tF�R��Bpm��O󚋣��Gݛ$���L�`q��	�ߴ�b~~��˿�'g�^j$Z�����sF��+��gc�Lj�!��
�OC��t�a��Z5�0��\%T�Bdu��#"��)��%OĖ�z(dS�jW|�X�ȩ�®y�½��}8����o�n��q3�����ik�?q���Zu��P�bI���B�#���ͱ�Z"=I�cJ�O�oHot�����p�R��{�Z�s+z�r'F�8� ���t�#?��#���V9R2r��J�DGB)
��k}r6����,ꫭ,_�uU����י�ٗ�����Ê݇`�]#D�'I�a>GW����6-G�v�L�a^&�fP��S�ƨ��0�c�~�����x�
�����X�r�P9t7����ؕ�9�ۻi�� ���r���P���Bc��GM�c�rK� Q�3��J����n�G
Z�����F�\�\�3����)b�#�b�d@�WRT�:u�7�� �\����}�i��ε��(~ 0�����������I�w��%�-��I�z�\�71n�W)���++�Q��FcB�A�)�0�W����6w恛�S����l��b�<��x���s/��3�
�'+~�%�[H�΢%��=,Wm�Ӂ�wE�+"�`�9E`WS��y��M|ut�~���m]�Ĺ}f����:�A��̣�����_;Ңk�� ����Y�Hd�'��h��SM(�H轚0$J����D`��[��;_~+[\�W5�B-�eBB����F� ����/��U���0J,�avYSq��oP������5���f�i��W�����9�C/�}#�����S+E_�����,��'��B?V�˿B�Y�)	Hd֙;_
����s$���ut�GH
�k�<e�2���O��۽g���+R�X~���=cl<QL+"Q:���7g](��/�^,�y�0S��,QQ���Ӥ�!�����Z��U⸝E�?§�V���⋕
8�׾S..vU�hC�J[�І�^�~-����JLH���9ۙ �	3�-����9��� |�+Zv�*H"٭R!��	�d/�f�aM��Z�=Ja�a���T����졞�Ҙl!t1�<�_�=����8x6ʣ�Y�j�/^�g,�"��wDv������%�47+e�*}Q����7��Gv
��u�[`��������RM��[���)��0F��Ps���4(J���NUmK}�Q�1�XD"0:�GS�/�:.��y�)-��0�D���2��.{*�1s�{P��v茠��(2�����&,#��δ�
�4F�K���� �mK3���3�M,ɉi/c*�R�`
H՝���� |6x�y�r��I�v..�\�3�9�>�����X�%���wn�O�ڛ�hn��ʄۗB�����xhN��>T�Gv��/>�h�z��*�J��f!U��n3�eҭ�	\>?��!��DD�ԡ�����y�F5BM�ُ�R�Uj�*MA`��P�����TS�$�Y��T@
Yp���+��Ĕ�R�2��P����z�(�U���l�V�P������B~;^i�����k�B��4��h����|��9�~œ50�pF��H��j��c@hU�`Oo�mT���mx3�<�g����p~��.��T��l�C��I�ϊC��
�Έj{e�:���𗇃�؇�:�{>&�T�R��D?R
sE��Tc�^��%A���ӣ�d��y��r�f���RO�N]��S�J�i�e��P��j�,ㆎ(���2���BM'�f�m�{昨L�h+�1��՟�y��/�����{��]�.�'UT8x��]Ny|1�zW:q�~�7�67I��I�Y��Ҵ
/:Ɋ�ˌ9ٻM�AR*��-.DQ�S���p��Ehʢ��aw�".�c!"�߂�uE8����_6�9�'}�Cs��o��yi���'�0z����Zm,v����u��)�SW��C�q_�Z�`˄\�0؅��zKH�2�� ;����f�$�SR�F����? ��lۥY#�Dg;� .�e�PDE!cM��ښc��bR��kx��"O�^_�EG�(^�l�).5?Dw���WWJ�o���o�N:R[;	n��5��+�%��x���)�E%�:�ˢ]cN��y(����P��,���_s}'mr�>�������"���~��%�G����cf�rl��ǽ�{���5P�3
��r=���s���ڛ�����8B���f��V|Zg���$�yUO��V��{��G�R���p}Cc'=r��`�b�B�r�Mҋ����K<����%�jIiJ��d&�2tj$U<��,m��]��]�>�h���k�:"J�V���.�r��D��Xېk�(�{N��ƕ�F�]A/n�&"� �l���jS��=�rau�#���*�°���# ��\,�>{f��k\���j���}�v��,�)��_���ز¶�2��_�JJC�f�m&���aɄ
�{U��{ʮ�D�E��{�瘘�J�&�r���T��0�"l:.��$q[ʁ�^���/�k�Y�$[��������.�!zvam��><��0�����J3��e�����U$�Ks�	]�9���x�@ �����R>�o��Jx˻_!^p&��e^���U�����dj�ȡar����TW����0�ǒ��\%s�����8
Q���i�$�Ea�ѤXJ�m���n�֙�ű?�\��e3��Ǌ�R�������GD�����{�i@��vw�%�F���d��F��������GQA�YO;>@�5u񃷆�e `���p(�����z��;�� h�d�c�&�k��$��)g����1v
D���d�r����	���Dm�!5�Y ���j�سb��6K#������?��� w����Iϸٍ_HX�0�]��~� ���j�o��kG5۰V"'u�Z���OcV+0A�����Ź\�)@2 eEFhm��C�h���_��?+��_�tW�+��A�p.M���Rl��f�5^�u�gR��QE�٥pg��w/7��R*��Z�K|b�-[3섥<zE^��ƞe�z�K��R�r���p�/~��}�qS����_��OJJ��~q��A:L*�1�8�n������3uTHk5:�7V����{%�P3�j���;j�9�x���R���6&!Y��� IHY��D�.�����G.큐��F�?i{��=aC�����"e*�}Ԭx��&�� ǀR��q�'m��䴖uJ=K��\���n�\0���`#���8~��2���4�񦧁�ψ��Z������|N[���T��#�Vحt�-�
t�ax_T�>Qw�#��>�sD�. �l��e
��n3?y��_�O��W��mhj�\<��R�m}},����CU���0S���L�m}��!r��0m��.�D�����4���$�h��Pm~��)�x���p���K���\_`.�_9���֜"�翙4pNB�l�,H"
3�塬���:̈my60!����c.NKJ��Yܺ��PL%�#��E���6��L�s���>����NRS���ݪ>+x�ucB��/Ыg9��y��y:�Y����^���X��E�K[�\�A0�ꚫT�ׯ�9Ȋ�#D�h�lK�z{�����w2fAcQw
���ꡦU�9[��s�8�*]��l�x3�N�
D�x���(x$���,X���P��d}���ә��T	H^{w>Y�l���~�f����-���D�T��hӏ����m0����&�0�,G�s3+�B�����k����l*��}�	Mw�EAi���o�2�=d}�Y�F�,ѫ@3S@��*���F2�~umT>��mo���JR����$Βؤ��m%�C����ǁ�$܆��it����1ϛ�1�hn���g�jy��u��4㺅8�Y�(x��s�N@{3�Z5C�O~�ig����`�(G�0�SA,��:ERx2>s��.�#Br����d�4�/<�>�G�JR.@��Ҏc��K�8A���w��Ci��*�ي��g`�H�>�{6]S4����>��X�6�V�	(�4.'��P'u����ך����o�\��)��8Vi��s���`�*���ʉ\ݷ�Ϗ2�8�Tx���1�9��3S�_ro�����hv��l��4�6�%�#xI��O[p�/C@]"��B��a�����T�	���ߞ�v��5m�Q|�Df��]��$��F}ܜ	R�����g�%q	��9���3���{-e�2l�V��Q ����ޫ�n�O�� �B�$8t�G�r4�b{6 ��*J.��>_/}U�rb��l��i��U>W}ॠ�5�XQ����C$��;�~ta��[3�̞x���tU�c�%BV�ãEfv�:��p�J�,Wv�fWE�C�L]o�E���/]��������zX����q�MO���T.�1|[����1��ƹ������|`�xG�t��_,>�1���N$Е*u�=T4]���%a�kî�v�.��!+EM�I�32�I�����Um�Z�*
�5��[���Q�|y(([V!�Qc2�6wX�P�Y��C#4n�޿T�DF��o�A�7�'؄�������_@���w�UË�\��#���xZ��6��h�̪\Q�;����|!�B�w����{�Q�u�E>M�g��
�R��
zV�'������\/�*�I��nyJ��\�.;�5��M�qȪŊ�?��lW,�祢��"�c�y��\�+F|Y�&A\��Eވ��n����#�c�~|*|1/�:������<Dyg��߻�,V Kڝ��">h3�g��q�������Y��M��������>o�%Bġ�<���B~�5�rn8��B�{����k�r�SZ����1�K �L�2�Ɏ��h7���ρmG�H��E[�V�N��'�ʘ%��c	����\��X��������-N�Ӫ�d]hK�CH�d�eJ�uo�`��ꃷS���Y�8�i�KY�(=����t]-��qz��۶fl,�U��+��S��ȶd�*�!R�UD�B��M~�]��s{��4--p�;�4�eq
��ʲ�Pf-�n�k9|=�IG��Q!\R��!��/�MR=��_'ʕ_Gqcb�q�b U�LS���$a��(l�U�br����G0�輈���*
�Gm�l��Z!���PQZ$b��{����h̭*A���k�P��e�0����6$X� ����D[� ao�S���\6)T�<F��~�QD�-�6�!�oǑ(&�~	�r�G���h'j�L�b��"�{Lm�\6	��ɱ =��!V����Bِ��+FD�w��z��!e�K2i���W��3(�ܰ.�$)��$�5��׿S%H��%�B/���S;��X��(j�()F�? �}+c{F>��4ԡ�ǝj`y>C�/N�s,<*K�]/+�"V�m���N@(�O�䪍�.K�&�˯�3��ٓ�/p]����;y�:���N%��7+x�WU+oI_!HI'0ګD�:T�T�������$&��}�J�L~Un+d���� Ŭۗ+)RW�0&k՟�F?�\�C0�jYJ�H���14� �Ϡ3����mB ��s���r�U3s�|rGPa�IO�w�ſe�����l���l�
�0a���5Uä�
*�1���5�Ns�K��CraK"��|L��-��/�fGl���tcßR�ݲ���bH�-���wiȰ���+���?a��4d��*���r$yv*o!�_{���1�f�9��{
���U�����LJ4����>< �0�[Դv��k�Z�{�9�����v*�tT���#܃q�� ޱ#���,�U���t5V`��.�D���xz/��H�d˚��?��K'}_f�Ȕљ���WM��(XˇV�y�X����$W�3��	\iG�.��)�=�.���� K�3�z. �$��ϹV��I۪��oaHT�Y��tBQ�O� �	"t��l�}ޒ�n��Kk�;���g��4�pr��d�🡥���o#�P�:�0ګO��
��i&$�4"�h�GB-FҠ��u��ZA���.کY�5�!Qb����������;۩_�;�{�q�lj�Oa ��W�'��}k���g�� ~�b�����L%�cjJ����X���}F$��U�� bwa6�ډ��F��az!�B=bD�n�L�%19DƟ�������x���K$Xj��k#{�r3�Ulbܱ�hD�AG��o\���0�Č��#�)�Ƅ!���Vၔ���N��b�:6ñ�4kf�Ά�}�.,�)�Hm�[��^��,��Yj.�)Њ�G���'@������2��-�b�cmh�sA����-����]�1lGƒE�^�ɋ�f��6����\K�d����G2؈�Iό�G���K��-��H�����KXkl9���Y�*�ށajҐ��{C��Rm�u0�V7b~%�2<��K-76U�}4d�y
��d֫�G	׎����/!z�����CT G9o� XE6|��{�˪p�%(�Pf$��c���%�^��=�8(�~r�1���g�$�Bt�N����Y4(h�r�=x_FD�󲮨����ZjXoEFJ�J�ʴ��g�-B3��]��c`�|ؔe���
	�\	
�P����W����w�YB8�?����dq �H1�v�/f�lX��$%[���{YW3<�MM��4�%|
�xû�g�K��*k�������֬dǋ]IS&Ta΅*t.�\뚨t�t)J俸c%���QS !��}��P�����)�b2~�p!�(�*y���h���U�,�ve�>��Eɴ�>�Fa�6D�א����߹�?;�1��)l���ğ�&t��P��b.DI�a��[wZ�޲�Q�GRw�Ep&�"ax��:d����z�PUk0:EU���C���]�����k�"]{ܮC�P�FBy��84���
�mF����?�@l鳴�Ԉ�_�t�o�˝�JI$W���[�v�relc�f(Z}p�����2ے�� ����WǬV7W����'����n�c���Z����J���ׂ����!H��-�ִ��UP��r��y����ۙ�Y^|)}��1��p����Dܛ�*�y�3Ϩ ��4�_�y��f�}tG�ŵ��7��V�f�+�&�7�>�.3 �0{S�����nqu���f	�՗粬���}�v�C�Ėq�������$���(��H1K"�MȰ ��]:b8�$�&�����.jr�GiFe4�G����x�*��������5��]��ü�)�p�5��?���׺<�m�k��������e�g��`��pp�C����$�3�����;׷V
8����=8��U�"��۩��Q��L,����m ��%s-`9Y�R��� �<�닑�b�Z�w$�������,�¨���w��>���0z��%�b�{���o��,xQV&�$t<�r�[��tX_��:��Q�k����I���&�KAD�]�-�8��)���7�j�A�xD�9�G.e6��JS�����m:m��,f��q��L�+X�@�0��v��S�`��K�`��8��O�t~4����K�	?˛�OC8F~�	;c��C��}Ė�.�3��b�t�]#͆��a�q��q�Ę���@�M�9u��WM���m5T�2��<�|�J|[G�	�� �0���U�i��	�s{��(��r���#~!��r�BI�˴��O~+c�'�n:CJ��r�o�ztъ��v���,9�c�I�%�{�$��n3�G��=��~���&����p��nKO��5����,�פՉbm�QMX�TB��O.�=�X�B��JJ��\Kͨ�޵g�@�o/���8*U�Ƥɤ?���aF�������G�{KG���ym���jז:׮D���h�c��������Q��i��fa�%R��;�m��}�"�58�Ջ~'�c����R�i�RZS�z�8�")i0�ۂ��!�%S�*��8����#�ŤQ�_ʦ�P��ԇ�Ȍc-Н�3�#n~0�$~�-;z�ץ�Y{������Wm<Vo(��Ws&b�C=W*f��zLb檊I�ڢL���^�����N2"���FS��� u,�X̠ӄ�4�����s)F�;��I�N�k�:Q�
���?�{���T1g��H�P4y~��Q��2�i�� "�&��]_�*z�����zy�H���rDa��1?^��K#��ڥ���0KB9��)��?��\�M�!!?��;@�Qp�{��o$Dk�0%�2K_b~{���v��� E=��i�Z�"9�8R�!�sȯ��j��5#�7�1��p7b#!k�'R�36�[���k��b���g�|�������r&Ƈ$�d�ChS�K��6_��X��`6m��!�/Y-��{�Z�����&�|���Ű8��/�7�tV,|3���l�����������Kî�����q8D'|��C6��ơ�YL���5u�[kv�b��u���~g������x�I�`��_E���c~�;p��fpg�1��� .遒�����ȎY��R�~
���I%�B���,���z�c���)F+��[��� a-�{��{C�?;�~ty�n���50�U�H�.��ǇR�� IC@��Xk5���^��-p��C��W����0���wp��t�Mp�61/���!P�6���VN���P$Sޥ��!��BgX�?݈��Ψ^^"%������n4}����`�3̓�~Ǌ1�1�ս��W��^�����)7����*�OL�Q����% ���"+A�P�s{ɂ�P���n�j�Ÿk^�����E��bL�Y��o�������f��0d�	���\KP�?5;��Q��w�=(h��L
��4Hh����T�ӝI�WS(�[ⴈf}�e0�ڥ��zp^
�E�������=SM!'�)�&�l�|�.�,�S��F@qƝZI�6mxɎP`�[�$`�t�H�ȟ� ����c�=�[�c�)�3`(�m~҇R�L[pS�Ъ��lZ�#YErD��I�<���r�]C`�Ic����,`�".��2�x��H�:�=���;���G-�Rv8�u�Ud?}��Фe�u�k�-V�dA�*��Қ�6ӳŘ���I0���/��j���a]v�]&X3��Q�t{�Zq�j�Y�k�	�����̈�&���y�0|4���<\vO�!2D��=Đf���q�r��3�N�.N@%nRKs�vf!��N�p���D�[.I������9Ր�of��?��)�ӵ�7LZ90��_����	+���Y`5���U�Ll>�%�~ۮ�(�zKe�6)w�'ϟ��dL���C�b�Px����<��0�G�]��z��)}R���ɐ��cA:F���Z��.�"����%�B���54�j8�a�=�n�-5إlo�F`c>��x �{QF+Y\A]+P%A_K��~�"F�AG�F]Z%�[�D�Ê#MB�%�8�ʀ����0��xi�c~�JX�V�da�udu�m&J�5A�E�����H�ϴF%��}�6���i��� ����@��i�2u|���,��Z�L����1�O���/�Q�ϲ'�G��RR��2#>�-%�M�n�� :~ުTŎӥ��������~��Y��_���ّKe-�Ck��> ����\RviÚ4���,���w�A)&��W�o*%;~�`̶r��3��4��Jm��Qu��v�̍l��t���
�Lz��0޶�.��562rO��2��N��ˁ�B��Y{s1�%�A6)o�'���.� �	���X�ۦO�k�!�O�?�o#!��hj�MF���m�a�¬,�"	s+?��$��p���~z��U�����������<��W�
P.߉�l��Ű?B���&��M>m�&-ل0ES��3Ǜ������U������Bf6bW��y��ψ5�ѥ].�ѥ;�j�E�'O��P+�cio�NBKV���:�7��$�3$��Ͼ`܏+�L=h,>O�,�8h���>h��3yeq�|�c�Շj�e5i prQD^e���㕮ӿ��7jy����I{�i�����[��]�ּ�M�������|B��B#�6��*[>��GC�e�&؏�l��7z��+^�1��/K���!�}���m�.���%��������`魱�g��"�����\)�\�TZ<���\�=�����6�R�~2k�����"UN\�A՚�GeH���?��y7A�N��-Ϩ��=I��G���{�O[�����u%��I�"�}�7w�XͷR�]����׻�� ��b�3v��A� ��F*�ٴ�g�_���:��j:�� ʀ������d1�[�fp�En=}������Ej턱�2AT��MZ+]e�QK�c�$A�W!�R�y �*�ֶ����)���ˬ�G�rms96	[�=ʇ���+:1�~���BI��`OM��S@�jV���n��)���B�(*u�0��9UlF-hx ���j��Qa65����a���u��DXe�'��8'9�8)�2�,ߗ���P�ö燦}л���[$}+�yF�6| �M����Ո��LU�j?��Y�+��7��=���˥[:�8�2�Y)��uU$�d�ѢS@J�R:���l�i��Us^���(׍iq�cf�L~��O�+F!ݱ�#ۢ�ğ�E�޵����={�(K�j ��f�/���.x��J�U�#lVOվ�E���?	�UQ&�+yF�&<���*L�D���I����f���B�%�$��	`>݌U���`aj�*3��o��-R�`e!���>�2~v�Yw+�W�d���O� 9�+;/�ۢDQ@|@�ę�2^i�ҽ&4�� :n]=�a��[|� ��w���m�h�`��Z���| -�ѿ�)ZBIzH�b�_Yb�}��HF.�Wg��;���o�9����2	Qhp� ����e�U�d��4��qnG�_�������#ܩ�1�p��u���e�yi����z��f�v�g��������#q:��_�hM.��3(�>�͌��ѹ T�B#�:�ջ��m�)T�o��ϫ�=U��aL���u~����a����'
�z�Vxu�r���4�f7�H5���>dxQ��_S5��X]�26�z]mA��dj$�4Eyh�'P?:9��j����F��=��#imz�Bk����7�Do��8� Ym��h�_�4���W���'g� �#'��^�,�f!����c$_���wï�r�Q�U��Ԗ/�+���:cN�&t~0?2�W(�)�,_Oޤ�+�l��D+�B+�veW�T�<�ܻ�|�q�T�߾�����y9k�:��l"s/?�FV�dec�
ny>j-��pȸ��,d��<W���A�<1��cXq�5��B,�h�8r5~|���i��4�Z�?���EAo�~ã�
����R��f�ω��Ӫȯ(Jݛ��XC���ܳ��P--�����S�,��g��e/�v�[�Gt ��V��$أ�DЧ��iI�&�_�'���Y�!�m�<���W%v�Zުe��Q<99 )+Bd�F���L�HhFxW�2�g}� ��H���ϯ���XLrt,�{�P`� ��+F�џƮ��R��C�Z����|O�<�W������f��_�
2�0���G����
��}������|����z.��8:���h>xzN�R(���~dF2�|}��h�zD{C���s)r�ĵ3\M'mpCR"��5�_���\غ��V!Ɯ���&x�~�0Q��W���5�߲��S:u/W�wܛ�W1[a����h���,{#.���r:�ۜ��9��B��j��Q��(+z�Ə�G�t��?,\[�F�sy���1V���(Yn�PX�y��CX���dA�xj��k
-��+�eP=��3��=l��T�K��u���&�������!,P[�w)ۡ(�p"��{�w�R�_ŷ�ui�R�F�Ay4�u�j-�f��<�ğ�ʡ��㰊��On��}C�{�H���&��G�k���Ԣ����@���y�C3N�pP�F�h��A�!�L=H���Z���~��&-0�����S�M����ڇ��X��=��=�T���VX}��p�B���0uӴFʕ���Ζ T:�c_�x�[J	 |Q�f����0��b�-�ʦ:��%��*z<��Q���	kr�8>5�%��u��My��&��
��oy�r�H�Ǥ�uP��n�g�����re.<$Gs�Cd���u�j�h�����A�H�3,n��E�%���|����U� S K�aX�Rm��C�� �)6����|iW~��[+��tȹ�j	�u��%yka��]�+���ӎ@�|�4FuY�-��|AV����&a�L���
�N\�2��������j��q���N#e?���9�/����;��<��jjh��To��\1vh8�p�A>�:��R3/�F��@�?������ �1�j��ڑ�fp�+ N��OW�q���/�̊(�o�0�ʎvS�>?B!��a�ƫ�8�S�5�m�a:�!C�1�6?R��J��y���Ev1���(��G�.�L̜녷�H��a���e�a�aT]��"��mD�F�;�Qz��&-��OAgW��c�O��WQ���1߀�+������ؒ��S�y�zMOxB�vY��qF����!nT+@M�i���`��#I$��E�)�+p��R�a�o0�~�٠�K���l+6G9[����yoYC1R̕����y���� i�#S����F��qu���p��#i���A�3�����n��TK���	3(��P�
�0X3M~��^<���t��U��M2%Pj�+7}��륦��\z|\[Z�I�������/�+N�� ���m�(k�##�v��e��-΄���37���,�����)G�qY������%%f��l$x�?)��(�Ĥw":�
0��K���Yٝ^/2���"����e7��bh������B�#мo�D~����pw�����=��ӗRf��'-?��RI8��+��uR��6�13����o�]����;��zQ�,��%&�, ���Ȃa�Ç�YcB�+����ieV3>BV��/?�K'cҏ;���&�v!7@5ɔ�}?B8�lW�����Ql�R.�>�u��i7yxO��u>�M�#������7��%�\r�z�ǹ�*��ډt6����8��D�G�m##ˊS.���ȞO���c1�3V��ɫ��%{1�b�����	η��ﳯ��;�]\�J�,�_))g8g<�t��p�_Y�A-V'+*>��}����7�CjU�t6��WU$���CG]�yz��`���3F
7�!7�`@����Ftgk�Y}ۄ��O�^���2h��&@�!���Q�"S9&cq���"���Vs���`Y[�w�C�S0{��k�ڔ��6Z�8
�tv�`G�r�%e�J%F�����D��ƻ�H<'�:�6��4V��5��3�5Ѐ�!|a*������P����
�1wf@����,4�8���C�dz�1GOlEs�7E��Ǌ��Ɉ�e&9c�B��_*Cvg��Nx��l�J�m��<�{)�fŵ�H�ԪD&�6�_^@���R��I=�/�	8�V�D	_ sz=*��[����Y^W��H��!mߊa��%�?�tOe3�qc�ٕ��	�:�/Oꂓ/�7���u�}�TG�0޼���>���iJ�|��O�B���z����avl�>�a�v��l�!�����9�o$p)��mOڤ��T^���2���k�Ru�Α��Z r|,���o=����J��!���Ɛ&�d�rR���[]�1�2�c��h-�+�d��U����/A��xZb8��Y�'�%��K�;�Р�CF��a8�:A|�z���W����Č����y��c��sT�c�h�&v��}o�]4�܃�����c�
\�q��?�I{e����$�;(�T��x���Y�vbT9,-��J��fдL@\u�mj�i۰����6�J�,a�tS���s����A��F�,�Q9�ѵ^�,��"X
),��~J�����>֪�����ջ��l;u"�����ۚ��*0�АS���:ny&�ǐ.:���$P���1���{�$��T������q8���ǆ�з�W�Wi2�J��tE1" JH������t�A��3u[f��^jpNW�h���\����%����J\��u
��#���aۥ<�w­��V� �oB�@����fT��s	���yFh~��6���J���g[��`���k]�VS��҂����a$5��D/��ǌy��K��p4��'�(�.b;4��3�G��P(���H���T���x��]E$���f�L=ҷ��[���l���O�*��f�QX���N�"$U0�p�RG�R�D�T�FˋHsd߈�������|���?�/�&׳}��#T�X��3�
��[��ltl��[�����+��wυ�A o���:Ї��"�F>(��|�R��A-_�qol@�(�>�tQd�B��'dRRҋ��l!f��	K��+	~{�M7��{�IP3�<Y���8�@K�J�B��T��^��WS!�}��2� u�ߌS��t���ey���Gʮf�/u�! _���65�5��o��և~(~�?wC�Ё@;~��V$q�b���mW8��$�ƣj�9�Qt�ٸ�l���ӳ+}�I
���{x��D�H{,����Y�)G�a�ї����y;�19�����3��Z2�p�.���7��`qg��VS���,�Y ����������{���Jݿ����B�#�Ճ�\m!ļғ���|�����$;,@�k{�,;�������q����/�:B�҅81s��PDo�?�8+��ς1��y���Q�;��&��b�sHOP�o#鋉�5�12�hg�lxDf�AK�"H���d�\s�e��)�5,m��j�?$�-�(�E*V��Yz���<e���`d�o����E�I�$i{Vc�D��t��X�J�T�ܳy�tr+����v��ض��3{�E�+�D(��M�w�`\����b�{����v�0�L;��̃zs|H`'��kN12oK��Iy��=�&?��p�}U�~D"��2���p��#,E��n=<����ſ�*���]����L�+��'�Q�Hy�b1�¾uу�Av�vj�Ȩm��K�>���T�+`坣.g�iF�+��-�#����Q��CNأ��NX����W3����8���f����=��g�t�["�݌r�.��_.��'�m6��NV����=w4Y�����>�]��.Tz#Q�?�}���Z�uf��mb�lP\
h%~��u�s%������u�I��*_ER�"���%+[A�].�kɁ��~�m��"�둣*� �8�W�u�� ��M���a�V+:�kTP���0S�;�L�P,#�:x���k����@K��TF�o�O��l^d*C�1��(I���k�Ϣ#�B]�&5FzX/Ⱦ�r}}f]�s��v.+1�ϴ}~=�4��!%��^�p�B�^{܂���5��J�Cϴ[�����ӀPm�T�D�fZ�Y6j5N�����*u%�ʶ���"*�lRm��ۛ���g��E8p��~M�(@4U���1K;��˅w6��p��%�HOa�C��=��ͪ���ɤ���Kjb����v�6O�8����/�+])�^��h��#W4ʚ�<j�4+oPe׵x(��N������hQ3��� �i��x�Kn�<RY�q6H�ֳ��w�m�*}�j�Y�G����w���#_�h�ڕӨ�Y�<η��zf�_\qr�Đ��A��hÏ�'M���Ԥ!�V�-#������TK(9��A�L�T����u~���b�'�Eі��4F���:N;�o=���ae��>U������ 	�a�B�ѐ,�A��\�_�^��y�=��ڞ��!�o�{df�1��J�����S�����Rj�n̎S��p�0��sN�޲����>Y9���k4GtӍh5^�nX�Ћ�\�����<�s�EX"�>����9�B0��@���@e�!!D$tYt��HuI�S��p�9jb�k���4GG�i��z�P�|����iY���=�6�`p1�/�ܿ�J��IY䄒���� ���d����K�>�s��?F�ykQ~el�6��b�d����'h���*�AH�W�^�y���?\6C���팤��-����ۣ ��lo��۪�Bj ���b"%e�\�\����$��m��Wx��*�jANl
B�.j�H�H���m��<���{/�w�{%Ll�6Fp�0�U�.�%]v?S��臄n�h�ݸ$\��]Z2�a����rM��@D�ceh*�ܬ[�n�����($R��=t�3H(��@d��{��:���F�W��.�a�P�g6�
2�?��G�V��;t{����a�OV����_=���-�>t�C�+�6�޶�kV��iC��x�N��a^x�����j�M�}�ʎ�[{����28�G�x׉�%^y��H޶�4׮�)tQ�W=�x�#[W� �ļҝ��#�!Ӕaw#KU5���O���x�u{z��"+Lg�~�-�����)�I���m�>�m��;���Y�Ѕ�`���[>��"�}��?`��x{�XP�~(��"��d���fQm�Of�Q���)V�l��$W����ip��3L��%n�����O��7Mae��\�jJ��Y)�DX bf�����y�A9��I�X�G�v��l	�Cy����Tq�(R�8���J��σis"�$�N�^���T�����8�p�e2E+z���2��L����=Yy!��e�x�$X��$�ee�y����Գ��@�����ݯ9��tVJ�mZ�_�?�1�Ld��}��/�:/.�3���c�3d7gt�l<
��H�
f�ܼG_�>��WС�5����:� ��.`1]*�<�>���)���t�2�6���A>�%zTc%�DW�!�rD��*�{���C��	�OJ�3h�C���C�_��#�ybH��;�ebkӼ��,!`ܓ:Ч��[�
cS?���,=y���6�R���B�S�`��T�6�d���Ń���x���|������=��W����G�a�H�-W���0�|�/*�H>���k��SK�ȹ��ܕt�uvS"FYP� �e�3���4?��u�cu\��rW�a����`�b �A'��'R͈�2���`�A� /�	��v����)��x��F6��~^��zi�S�z��K� d@]�_�ѵٛ�(��&l��>/:s�������4n:��	]J�f�H�g9��i���l]C���׶~!';C-��Ϲ��,Y >4ih��3�7Y��_d41� ��c��p��6-�PP�S�&e���1��qh�Ո�39�3�gFP"X4]�U��"��.q,�n?�],�x�W��a����Y�#����F��h��8~��#�^G�(���>��t�\ۇU�@��n�LNf�`)ך�����)�'��Xcn�E�-[��۝|�>\�����OC�eހ;=o���M@n�{5�?�L��-�1Sۨ楬�s��-�HG]��-� �n�x�j��:�������S�h+��Bў�4W9e��l�����[�O��`�wN���:6���;���%�jL��;-pnP�iK�ЊX�*s��sȯ�^�kV[����1����Կ�]�V@���aV=�#�0�,\%�߶��r��1>��;�a���{{��X�2�7q�
��i���|0�^"w�e��]Msˠ+��h�릉E _I�9��W��")��X��'n/F���\�yk#��;��1܄eK���|��ߚQӝ��?���S�
Un��P/Jz�zDti�T�Y!Ɠ���މ�KW�M��[�.�����cAQ�ı�`}$�9>/���[��&�.C����t��d��E�h��Jvzi�o5Ú�@�+]5�@��9�sQ&�RxON�"�^��<|�Q��NH���[b��Ц�O�iA����i�Ŝ�"N0|�cR�os����Թ9�af�zZ܆��J�Q0T]�}��\s��o\�v(_ϖfЇ�<]��?l?5�Q���;�ndK�R�w�;?Uq�ۧ���qQ�� <����R,5��oE�^�b�a�LB4Q��Ɍl+�v�7r4�\t���y�s��f9�Ȯ�|?��4�s}qP��A+�F��������L�������K�&����S�+����.���^�9[$e�;�N�8S�����(�
�E�㈼6�:Q�U�A	�HKx�?,J��X�Z�¼g�Pm}+G+��v3�=�F�sO�	�(2KW����1ejhX5��&$F�I/s7�6Ð�|���9P�N������mik8�{�N����a⨐���_�M�㖠4�K��{��]�a��H���Ks8�ς�d�M���.�9~�\v�r�I��@8".U�U��=�?Q��Xb	R��G�zծ�[��cy�$�0�fD�ܙ[���[O �Ӊ�Z��*ʨ�6���d����q�Ϭ>w�lː���!�JUlH�i���ǵJ��t�d�iy�[G�E�=�6���F��H��ձ��|m��ꗿ�:	o��)���|]�V�O��U��Tu�c�B�}*�>�}��_*X�֥�yI��l� Dc�,�����t`���0�V\��u���#���.��w��F����g��S��<t\�.�#��~G,�܊:�o^,eY"��`m�p��8lҡ&�"���(�)�v�$����q��,x����8���>��	2!���9�2zoI�icV�B�i�HQ�oہ�>�|����<.���O��������\�-�4c!4��sW � �o����"
��8��o�y�t�j6!��B!��t�fI:)���L��ة�[i���n�����\bdeh�z��!g�GI�|;֗���O�~�*(8����i+/_;m�9���>�O$�2N���s�G2�Q2f�|.C�i����y/W2X3w�.�����ѡp��u�D�óG_��`O�Kw�&S��BMa�6&"���T`z������:���jruM��]��:a ,,�ГhX���I�B1]&��	쁆�GӃjfz[X���&ju]� ��T�Q���]8��"@v_Q��fQ� �9��R�ة�pR�/e<�
������ɸ��>�AT����`Dٜ"ys��ܴAJ�Ϩ�ź���Y��X!u�0Ye�	o�R���u"j��׿%��$�kFA��oӅc���iC�*\�|�i�VV�9�	����A���y*LR����-��X$�&���7̆|p��Db*�|���IлKy>������]J�ŀ�������^0�<�]�99b�$^:�;T�5??�:C�C�*�ۈs��;:�g&���)&D�zH���mG�)V���R����E��ė}ϻn�g�}	��y�I�Q�6$��u!������LZ��1�n�p� ��b%E��]�,�q(�ٚ4j��v�����uZz��e��8�{�d=����2��r���8�-ڻ�2���В�hK�i�� ���zSu��K�v=!�������Uu˗��= �&gCY�Zy?��jw�0RMz�ȸ�n�/���N�.���3��UՓ3��g.<
Lť�o�e4��G��0n�.2���E�+>k�!��V��G�'���c]�[�A] ����)�7)���?�d��`Vl�Ց�;�y��Z��v�ݞ�o4��Z�E_��o�cܥ�:���*n���utYe�G�E����/��Z1R���X	��y�]bH�K�m���p��2<E�����Q��>t���؏LA5E ��Q�;i*�5-���)Iǆhl�:�by����H�<Q�y�WW�mxa�.����n�wyMI~�o*�S��{j11�����t�?�l�5#[r�`[�Q�f�mw��Q�I?�~|��{�\c��B�aW`�x���>1�	=Y)��Nؿ���0��0�����M���I����q����{L�x7*��O?�3�czn�^��s׿��3{a�D�rh�0�!���z<��`i�t?/@5Y(ʁ�u�ݵ_E�A���1������X���a`E0:orW=j/ @r�������G��"`y)ԙQ4:�T��`�~��	WPV��	��턦���
Kw�D��c�A��s�{���!z"@����6�}��A���N���\�q+k#�i��߹��E��.�j�&����2o�����j��.[���/�FK�I>T����ڵԬ�i�􄢥����S�O{Ď����NhA(����_-�@.T�z�e��P﹃�v��Ƽ��xߥa����<q���2����U�=n�I� �˛�M���t�gc�Ek��g�G���n5� m����itE�젱�C��"%;��+�p��ש�8�͞Ѧ)@ϴ��I�OS�(��mDZl�ĩv�M�`l�\��H�fG����s�&R�gs�P����߰���-�<v��t��#t�My�|=nv�SϨ�xF�8p�5��!�M�)/;����St<<.�K*><����/8�
8�D(�-գ�+�w"cMԒ
\����h�6���6u�Qj6�����%}�ۢ0f����j!�a��­ڃt7.��ȃ�p��SܷN%����;il��>�&7`��`���C��ؽ�2����Nϼ�2�>��'/��i��S�&�#p��E����U��+�q.�U�����n ׀��d���IQrB�ӂ�TrR�|�YXJ�Ŕ��zVũ)���q�@VL��k�hRC��By*��o�(亂��J(V�-�-��Y(
���{[��ήE�y�
B����#c�1p�P@|%�[� �&u�9$�g+w�ūx���D�G��������7��.F�M�t�%�����շ�1ݫ*����� Z��/�n�U7K����.ъ�z���wj�����7=S�	��1P��e����zU�x,�=�1{q����Z�C�2�=���-=�iiʃ���X��]ҙ㺂�'�����W�����	6Y�o�w���ܲ��^�6fշ?=d\8g97�P_hn��2��ك��9�ȃ%�n�J�U�,*�Ajlr�03Y�m��R)���k*#�O(��-ڃ9�҃�A���TJ��\�����.(�y�->�#��E���.���rڐ�����/H#	���-Q���:�8!�	��nXw��A��rF��co�a�Хs�C�x�u�N�����
T��9���<�!�!��xbk%Hb���X5t1�/�`L�K���� �� PV� �����D��ޙe3}�F������9ǻf���\<e�^,�m��bj(�h��@zt8�d�RzwЋ�f�G"����/#h�T��cRq|:��yùJ��i�e�O���n)^���$�\|f �W p� )z��y2�#���Ǩ���
l����Ol1�Z���/�������Iꅮ������f�瓫}­�NI�=�ȋ_l�8��
;��
Z�/�������P��������_ߣy8]#;pz�OR��E�(��'4�~DO�+���������\� b��7߉H��X9!G�Z�O|V�%T�;��9�uB��Ih�^o���m�5#�P�<zݸ�� d���Eo|�V�p7uW���SY"�2�A�N�H<���x��89�'n�І�F�Z�����_��3�B����iV$�L��`�'�x�ܮH;'�яBNp�??�+b��u�����utV���T<�i�B�l�]�3F��2a-�f���C��>{�I��*����T3������{7�L�un��xV��/����������D5��~*V�g	�E�	V�Z����T�c����1���ѣ8�ɜ�=��Ƹcl�֣���9�9W���#u�� �n����F��V�ȚK�K9��Cdk?��C��1���⨓�5q��O���À0K�Ki[#����<�!V&5CT��r)�RQ�K�̚���deW�����,�����ka�6�R�_��J�P�7 �loX_JW�y��l�(�0��K ��-H��6�HuR�A`��N��z}	b7�8�QQO;F{"�Y���t����?���=`|��0.h�����S������j��F�OՅY����t��D �8����&��tY�B��wf����H��3?u�griњ��h"�s����u�j�ZջN5�(U�N�	7`�eu�]�R����<�����|��-��ڍ���y0�]�Jf�T���»��4�+�m�0\R`T&IN��T`>Ղ�
�HX1r���&�?�J����l�8��������d�L�����(�˯*���_:Os(��R�%Plg�6��W����]b��o�����'�4�U�o�O���qL	��c�T�xh�E@;V6�^w��~�ΰ���w��Z\7B�N����=�p���%,���l�La=�"���  )�*Ia�̲��֮���g�P�\���Q��ls��&7���3E��PQ�$%eHW _���˯�ix���W�W����ȩ��H2M�g ��� �o0�bnT�2r��p��v����#2�@��B�#-+Yu��b�࿈�����+�`g
�U/��_X�t�*K{�w�÷r��L����Z@
2�C����48�f:�Rldۖ�d��� K�kʳ�n�"��W��3��_f���1>b���G�]dWs_�*�'<_9���j�q�OI���[��r�rTl�WƯ0a��M�%�!��+ !"��U۳�:�G�y�s�O�伔 $v)sEg�0K*�����y���Y���W=;��`�{�׮�q��\�n�W��ɾ�lMQM��(�_�\���v0���$Q-U�Fd^����U�CRu�O<N�ϵ$�����'��_��ٿhG����z�q����s8��p BYx.W�H�<@���s�
4�f�uh3� �<]���odч��Eď)A�wgɗ
"��)yp@�!~+s9��WG�U� ���5er/C�q�T���B�-���uq���0~�m/{�6�@B���z�x}>c��T�v�1Ec�'ܔ�R�����܊��C�7��#�S�~��S6�ؚ�u����)�Ȏ͞�0�����/��r�Mth4F��4K�Ƴ� ^���~4�����ou�Ip�ܐ����&WωOG%
�{@O�!	���z>���a��!��l�tHZmdT�΋Ȅ��$�I�q��5k���eb	����8�`+����[��پ�4°%���`�W�y~��A�k�=�=��\�	|0K��=��]��5A��F��ۍ��̖������V�z]��W�������K�n��߄"�Җ3w�J�v�?����E�"�Q�'cqwV9J{�S���W8{����x��+��C�,��Z�DA�~ܞ�H��?4x��x/�j'.&M��!jj����ֱ͞��`;a�Xt�ҦD��:�K^�N�i=[����������B ��d\l����_�M��% �Mj�PGWv���9��ͪ;cQv�Ѽ{[��j1�^����|9�F��m�1�,k�q��%^%���7K���S�}��{НJ`5����^�:ܯ��n�E�zA(=�-	�?�yLU:�'��P
O�p/Ʊ$t� �-etkw{mDGx�g)�B���!r�<�� �(���*j�?��[���{�_n͡G���);�m��W�H�n������2O
͚ˡ��1�m���
���s����?�Kr<x���<K�kՇ��񠹨��DJ#���p)�ʼ�������� ���ʮ6��EA�?j�l�5ĖX�I_��d.���{�v��'#�Z���uM���eM)\���*.F�|��7��_�&�4I���DAГv@޾�\Yn�ѷT>���-�C$~y͚������q���q���!F?	2P�Oõ��R��[����B֙�����lA9��rHZW�nW��b'��L�Z��'�1Jw�z��C��颤��ll��+B���՛�(J4)b���qܡ��ˤ#{�i�m�6��y�)K�ʰ�w�ʋ�<
fa]ؿt�B��$θ�[��Z�BJ�!��S����3��FE|�f��H*�]I8��>+�'3J�c�� �gDv��>cǋ>^/�Y���إ�S��#Z�s��g&��Î���;
��쎮�(��ʄ-�r�4 �?�Dgu�����! �弪�J�`��ͬS6�\'��0?��Xd���4�:-�r�O�u��
�OZ[���81c�g�k��!(Tr^�TN*B $xȨ5���m��b���[Ɵ2��L(���wGh6'�G|���*k|!(k0���A\�j�����>�}s��q�݂���^��>��v��'DҸ��] $3i�Ƌ`qPa3��䈣.1�L�K�2��}8d����Ge騇�XZĚ ͬ3��x���|���%T� ��QLN�#�!QO6F����l�1�3�Q� �k�.�`t*뢯s��V<j��-��lV%4����^Ǐ:<���2����`F��b&�����g6�3�A��{�����EVa[�}��k�'��E�
��Se��*-��{
�V�Q���mH�-LR��? ڨ���6�|��?jĂ�-&�&��R3��TT�^+������$�	�҂�S��H |;�E�o�Z	g.dI��N\����
p�z1.������K�G�u����������2���4��1�UtI<�C�F�k8h�1<��{��U>K� �y
�ϻ
���*zK2�H�yt�_~��h�~꒟�+N�,�G����G^b%���~/�n�at́�)�����tWMxб�ߴf���˵ �r5`$V���`jG!��޲R���Z��q�i�7Žu���n���%úax ��wp�W4�X4�iu���[��ϣR�eqA��W���-�@����dzƆseob@�Q=���`Fc2hVPU�Zg�-�=�C=3EL�ޏt��O}%��ta�~5�j�l4��My��9���&�a����e˾��_r��.����j	�NՊ#����V��5���k���9�-sv P��Jŋ�p��'�9�VV��>��A>Ik���盃���W�-+�i�E�(yJHu���v�~�[���D{�f�c�@�Fv��4W�~�����)	�怹	~�oG1&�i���ø�OO�Y�?r�7�h�cW�p|A߳f\����Y����t6�=�J�'�E�j9�^���t�:��\xQ�0\��5� �~�KʕA��M=�4�"\lk\xVk7!�;��Ӡ*,_��^�`�@�$�t&�L��L%��'�s��]4 �=p-��M4����"p7��i�FF��E��ަ~XI�8&H�6��|���W��5Ԛbb�x�vv�C`���+��z�02T���er�6�D4\~�D�@���v��̜��V٨�H��� ���$,۹�k��lf�w̏s���r
�MI�����.��~���&��`�ʹD�
甕�����f�~=���ۻ7<TCg���Zk��\�:�����e�U:S����&�d�8 +��t��+j��+a�Q�������U�i4�M�0q�A{zp�A\��#��teC��j�>���.�Ǖ]^��E?�/x�U��^��*LoL��a���S��]�������mo0L�F�,� ����2,�m(��Ksi�?�U�/�������)���He�0�g6L�)��I�}~lp��q���"U�sK�%=��<���3�V^�L6>w�*��7d��/����X��L~DӪ��01���
k�q�S�b� ��ذgÛ�EJ��>�Մ.b�/w�wPSBػg5;���	fR)�#j�1�l�ש�/�"���-��~���Ո�p�&��v�?���ۯ�W�>������C��E�zd��Vv<|
�����}������sWX�Bp�Gp�O�t���6�y��O�உs������@�E�����j+䕉��T��W�5iߓ�QXn���^jw
F 2`�r��c\��Tkj���u�X���`g��Y@=��<-�<�&����N���Y�.�N�Ζ�M����(I��'1a�MB�4!l����I���3t,҆��!B�r�c���uq�Ƙ9(��.���9e�&A����t~�nJ�c�ȏ������iD
���R߆ejT��al�㟙�ZS�nB�c�5�0�g�>pf[��n�	��ꏹ�z��beޜ��$0|@�{�J�!��n���1`r}(�d�!9	�T�<qU����b@.��J�������.��#�Þ�B|~��#s�KD%�����]�h�Nl�o�寍�HJ�7��n�Փ
+���mY��W�J�Rzz�X��u2�U���Z�b��gkM)�=�@�n���ؓ&R��'�~	�T��
�Ӱ����){��l���Bvm=ak);z�({���C�Z�6`a�v(<�(p���zHut*�zNH27�M4��b�0��D�����b$�e��x�>�vJ�I��V�Z���P@����i��7"���駻{��`Z�Gn8j?�C�:��Ѻ�����
T�N ,�@��RDy��l*�="y��Џ�R��S:�tt�'c�WP�@o�2Ȍk�Ѧ����P�0����V��ޱ��7oUd��Tǳ��yH�9u@`u�]gaNfc�Cl��7=;�M�k0^	Q��9��� �R��in�u
����P���*T"�����jr�m��,�
zc�0?*bj�޷O�KP�4j���X]3�T�,o�#gŮ�y��7���&�牦��[����4��p}
�%��Y�yd���݅�*�a��	�Ef`6$K����N� �i�����3���z�\Z�Q}W��<�!�l<M��M�{���i�JW��Ň���Z����
� "��&�����ǎ�˛Bۜ2�a$��hS�@����	*�&��Ȇ��I�KM�k5��h�G"���/��ڮC�vз�1�Z��	�s�m��n�#P��e�\D����i�����܄d��h/1� M�:�\�Z:��0�X�-�`�/ؐ��*H�i�̀����޶ qM����?�@�@{_B���8I��U��M�ʳ8�~T��C�\!hCϏc3zU����;�jIM��E��m��М������R��-�%�C�t��)�@4���an�as�w�+�\�n;�i�f�����
����6�V[M�m-A�VJ�Ǎ�6�n��NF�ئ0�5yzNq���_��7��Som��mUq�k� ������ܘ����z�#KK!�]� ̤\1|N��]+�럅���:��]ޣl,�O��)m�:u7n$���(3#���Mڹ4(
��Ve�H��5���"�9���v�	=H��
�ժ�	P��3��6p�@i,>@R�	?��|D�]ၑߍ�mQ��P��H����e�d���q/7[��v�O�����y��W�:�e�{Z�"�ez�؅��M*_��.�]�GW M	�+|_�x�Uv�+Q�������71�l4儞0���<2�,Ѳ����D���j/��f�y�_�!=��L~��jhTq~E�*?#W[�	*	�)V��]��W(�ɸ�Հ����L��,֭A_�V�sK���|%5�i���Z���'�6v�A=�:��<ZV@��7hL}�[�����_&���@�/xhwv{�/�<����JH iZ� ���Јt٧�ϳ�ʘ:�������BF<����;�V=��[�qd�h�}R�!�oE{eJ�1�=�j���K���NI�9D<z2w�.H��0���~��z2�p4�D�98�J�>�� �kο��YikM�����˯0Œ���Y����сӘ�Z���PlW�cR	d܌�=5@�ޤ��jy�����w���|��C�8o��)a�ڎ�jk������]�K�����#3i�awv|�3*#o��SO��v,����ɔ��P.J�O�� 0 ����!j��Q���t�}%Vp8�?~��L��m��P
1=[�<%`%ٔ�Xf��;����MP��<����>�8Qs[h�mp� �t���K|ƛ���,�E9���Ζ`�	?����2 �R��a����ٞ' �8ۛ�H��6������&��Z�% �G���A�;�����7_�ð�[�*aHG��8���&�ݞ,��7��Jks��b�LmX��+X�E@�aӢ��x�EQ-���X�Ij2a��"�"��^{)���[�M4�>���3o2���1�p&V?��������xE�m4�vMCQ���\���H�fU�m]�4�v(��'3 u���V�.F���2ޔ�q��n޳u;B����nM����e������;0#�-;}jbL�wʹZ�q�����pQ:�q�S�)���2#'��H��F"��d�$}���N�?{�,�}|4��k�V���F�u���
z��Զ�I�G1���&�|=�-d�e���XBQ�s��'>��ܪ��i2�<h�df�"��O�<��n|�@�W�2]�������߾��g��B%ҡ^�k�t�TW����P�L�6D��'A�$�����@JC��3��[CH�	����l��'~��y�r��_,�j)!����1b~C���1cRBR����7L���t,s����˯�����H�f gW��{�_�h�x+}����Io��
��8@#��s����yX�0^�h�|q��[�Yso�����ʠ�΄=`��l����>''� i��`v�Z@��k5�������'t_8���Z�g�)=���n~ZF��\�U�4�Q��4��w�T1�7�A]�,���1��fP������/�e��H6�	��k�_��dU�q���j�t��|�~a���=�I�k/����8+n�y����\ ��0��ڬ
�mԘL~�T�7�m:,�4 ��?�˵+&j|d�R�Yu��J��ͫŹK��*Ջȏi�vn�M[��o�(��4����|H���,�i�ŕ��I�/�(w5΢�8�E�k������WBy�n��|�i�a�f9��vGZɶ�h	=�. Ŧ����7����Qyd�?�UsB��rw�O)'��&c8<�{�r�4@l$��Qm�1�Ɠ�>�v���� D?U��͊�&����/Xv����]	��)�ܵڅ����$���+7S=�Tn�,�0v0�-V��K�Ը`B��Ys6_�y+*��sr%]7�{��� TMU���n#��U�]c�o�~2��s<����ЌK���6��~����'Q	�Җ��|l�te�ǢU�0Ű3������9���r�r��g�\�¦ �л�Ky��`�˻2!+L�2��a?xR��nV;U꒞�7"� ����=�$�2��P�M'ZE��Y��yx"�"��k�g�ሜ�<K�n�q�R��$k��)�)m]����S�㝡?�6�����s��xa2B�a��لs�e���}�. 7�G�8���"���<�Ǒ����_��OW	�(�p� �5"Wۺ������8Szhq� R��9�?�X�����V�m�И�<��(-�Ԓ$�A}���G�+�#:��wՙ4�֋v��u�{(��&ʀ�������&�ו(� 

�	ե��CH2�j��k��(���gQ��^i��J�����i��3JV��
	���h��	ݩ=�ud�+<�Y(�I�P�tn�M���ǐ)+���Ά:�d��*@	G��w��?��T�8|Be3��q[�ϱ�.@s4��3�xٟ�i
��_M�"��%4碞"H�o,5f��Z8An:�r&6��sg��ؿ0��`��g�].=�T�v��)Ak�W��?,�6�����5'\����('�W��I �E	�5DZ�s��i ���	WrQ�n�����3�O�ￍeٰyg]�D㰏+n��>�Sp�r�����I�󼩫��f�ֆ⧊Y��A�Ƽ6w�خ�e��s���^h��f+��v��S1�'��9��Ⰿ6�a�gY�%6(� ��HS����1���DN9\]�? ��cW��?���	��d�.s��%���80�֥�1�߇����ʹ��k5�.~S�MېB�]�BͶ;�&ILw�ė�\tƖ��N*��P-�a�)B�f����?ˌlμ<���9b9
w�E�U�L5ojm9X�Rz��@G���ⷻ��[N�-,?a�<���RE>���u�q
Y8GjBC��MII��(��G����%������ĸ48x8���������W��v��º�}j�8���F�_Ȼ}'�h�������DSlx�2�R4+�1���)�0��(I�v>vł5�5��|���b��O�9�8Ro��BT<�ږP��ޢH�U��h�O�L&1z�3��7�.�a7a;u���IkW(A�uI���#3��<ϐu��TE^Y��0���H�����nƳ�t�g���A�}[Մ�;��I��g��z�]ӠU��0ڄM�-U?�F&��Ʀ}c4#��pD9����|����9ѧ�9
��2���;ƶ�g�Q���M���ǒPN��
"�f��r�w�(�n��C�N�{ʹ9x����؈_AdM�p�}�����?7у�Uā�|���	= ᛶ�!� r������,�A�w���o�K�G5��-+��Q��ȟ�N|��ւY�k�g�Ts3��d�3��~�j��/���ݒ[�6i|����Wk���1.Ri8�+���u7��L ���U�o�_��!��;�gaߴ;ھ]aG�
��{IY�A�#R�i�Z:>�G������yw����=��P~^���0������yԛ��O6�%݈�Jöo��=���.�'`�؇�N��j�����{@ܤb��w�M�{���2ۂw<T��f���5	03�]�xѪH�r���_��K���Ht�S�%?F��D�n����n}:�s_��pvI�'7�������F���՗?��ng�,3��1b��.8q�Մ_j,]Ϝ�����d�4�L�a���M��Ҙ�_��!�}@����R�h���GD8�YY�0�@��f���p�c�G��ё�zT����+`a�"��aGD��8�A!L���f�ޗ�a]+�J��l`H?3y�2�y�Z.+�܊��Љ��������Ӎ��z�H��Ψ�����p�z���
��F1\ϛX���w�A���Ѯ&�>��F�RN�E�B[١5�`Q�-�8�������箜���[3ɿ���t� ߖXѸ-[�x�f.�.�;ÂW1�!����7x9UN,K�660\r}��ʕ�е:��
�I�=p'��Cf��Ã�<~D�� �w��s��No�QZ�&}d���	lw�����j=f��(��cȌ>�(�c���FUj��%	ֳ���>j�0Z1��ĸ�4�H�N]���� �.�1}��_}B�@fJ罽���}�NȐ�|�0!�Vj-Ð�����o�G�B��&�|	��倁�Z|Č�ziG�3nO�8KS���v�=��!��!eD^�m�
�3�>�����Zu�c�J��-�_x�*��f˿�OԄ���DYi�����cYT~��R4��Ų�T�ߚU���͘7a�I�+��BNX�Q�8O�{#jRnnW��m;���y>�"��(	a�,бg~�ɏs+)&�SW�Ҹ���`�O�%P(�u/�۬O	�ZW;�dG�B�f�6��n�F [��K�t?-ϭQ4$�75��G�'����q3���u=��p�r�7Md�=������0�ummֿ$J�fnS˓�kH�qJ���џ+x�K3h1�0��1n��fס�Ǟ�C{��_|�"����آD8І����L�-����S��_%#��s�+�*cWS#oW(�ͳ���7:gЊ��vs���^:]<l�-P6xJil��]��ܷ���������	�h_f/?��Bv4��Q�.�_� l=�ۈ$���UbՁ
��9�kl�pJ�c�
�#$�/]�	ɗ}CӶ��tH��������4<E���p���j�J��V��A��iB���C������ұ���h�@f�78�N�� ���q����Y�[5�I��n��W�e�j�[���}�t��}��" �ux:"UC�aA����
�߲~oP�����Rߗ4��������k-ÿ'��ŝFK3�u��܎��mKX�Be�
��������7�O���K�&��=6��z}$�8<oA�n����,��*��BbX,%3�Ӝ`�Eڱh�F�23�GJV�.�E��6�f�E����u�f����3T�񻴎Ö/��ௐ}�w�0���
��7�k��Y�7&mIx�F�������ԩ1�W��Ɯ�QV�aҷS��[�ya)�#^�T�.Q�q����Rp������d��
'�0��^�=w�f���'�\��xX�%��L�0���15ݚ�� e��5Pvi�f5h���N_�Pk�O�(���T)X{gE�=�?��]<]�'L��Ŧd�f���7��o4QܽL�uiʇh�`���e#�C�ʧT'��L 湋XL+G�P*�`�����M~��zdܵ=�Ę�W��y� ٥+��8��}����R��%��6YZ��}#��0�tlΈ�����)J�%8�sڀ��B��ο�Y���IX�U�~��{��h:	�X���<����ָAI��2T;4�+ò>]�Q�SJ���H̤�kY�X�n�j-�5��g�@N�Ȍt���Z,�n�zć���/:a�H��X%�'eݶ4wϝ�`ub�5�˼Qy]�;��Q�/i*H�Y��#�>Q3�E�qFi�)�h�R�ê���yBbJ�'X��M�"J}��Q���ã��r�[_�/�\0�3�~m"��hSb��}_�\E���B�(�����:>Z�U��U��/5U͗�k�X˧썐8I��?@��o:nZ�-|�ì��1QA�m��ہ2�,\ؙq>����_i��K0�Q&^U��~���-khezu,��ٗ���%�]�w4��.�.S��z/�Y�S)P��_4YfǼ���4z{�ZX]7W��Kx��~T_uC�	mR��.�dw&S��y8��1b�nx��P��r��¾�{FV��{��ݥu���J�x��s�E��[�Z�ESyS-�ݘ���3D��)��?d��T���K(��\��!�MG𯄕�H̬#��F�Ddi& ��(��q���n�lt�M�!�0Y�iĴy��'bMt3(֪"�Cs)U4>Z�(�}bM��T��q��M���C�X�x-���0$��;U)F�׸&�n1����� ��#��������G�ۗ�P�\�Y�YZ�ٜ00"Mt�=h�sWH��[HQ/�F���>D�*��Ժ/`�s�#�^?k9���԰t�?J����&�OB���L�i[z�R�W��_��
�&���~^�oqpy���CL�%|�#H ��P&_��{���E�T` `N9��T~d��s���J�ܤ�Q��E>)�Q�K�[�	Ac]��Ҵ/K|�o�M/�������f-������(R\��ӻJ�lY�b��M�w�?�O������6��i�`xZ=/�X)��Hn�H��(x��\ķ��he]>f��}���A��U���:TyY�����h� ^�Y����Ї f��p*���st���0�2�}
b����,rSts���օ�U���I����jq�í���㣟go�lN�(� J�z:����c��s�r`���|-�����\DC����4����	�p
h��'hX�8��ٛ��G�t0�G\���|8r[��.xz/xI�_	b�H�
mru�c\xt��RC��gq�R{i�FDS�t��f��6(��Z�#��q�� ��j�x�RW�#$�g��OqԼ�����(�:4�+�*�ܾ�V����z����ߌ�����;��㮡 ��� �?|n�A���2�?��h}ή�wK��v����+#cd�{�1�*���l�����1}wy��[�~�〪:o�Eh�`yc�v����H,���ہ%i�
)j������z�|��R<y����%��wW,����We��?i�0����ZW�L}�cZ��.��6:	��"m��@��ZL��{����hq� ��ľ�t��4 .Y-VPb�E'�3��
��نb:N�	�a���h�fW�-p/r�[D��r$ɶ�Nm�@����,��S��A��4ns��Yx,c����t��<6Qo%��0���ewЖEm$c�	���N��B��RƪIszH�<�E�Y�B�ی][V��g���Ѵ)lꟘ	Lx?�O���aW������Tk���椸X�T�`���A�k����z�J�d&��|?���ܘ,���8D��4z�e:Ne��BJ�N�q-�������-��wZ��Ƣ/�u>�
��ר����w�,�rV6�jOLFՙ.�&�>Z�뷯�jʄ1+%C�[L(�T��Y%��«�6z��H#�b���TJ6�� �����7ƨ�JU{z����]��[�$�[K���TY��}\�<��^6i+�EF� �K�EGA��T�"b΁O[B*l�)�@C=P������',�a�X���\t�a������g���x7�e$(-�4�h:D�_5���c_SΌ ���RKJ��b��@�Y<��C�%:H-dߌ�I��iɸ1�_ՙ_4��)�Uv��K�[N�է����4o�M�@��IK�)�Ņ�2�O!�_�$���Ms��C�~QK�9s�⨾5e�<��!�ɲ�˄v&�{���Q��?������0&�y�* �I�ƾ�LuV6�Cg�K	r�lKĨ�Q��Q�}��N.�	T�?���Y)=,���
�*�F���h���X���{��⁕͒f�/���
N�I�A�u�1q3��ߵa�q�ԓ�Q�4�ے���+�I�m {ޥ�(�wg9xq�Cb�˹|>�)�8�8M��.�� �X2�a�,�~yU�P]����$���4����-���DQ{菾h�J�rtO˝~f�������hy��]�i����m�	����V�9�z�{�R�� 2=x����V[���j�C�p�D�|���� ��=��Ƴ�#ٓewѐ$ྲྀ���.P?;Ô�]z��9�w�l����\���n�EQ������"Dw���&4J��Y^Q�;��d�xݰ���Y?+?�̾���,�T{-�R}x���(��%N'J�=�Q���T�r~�U�5�2 e@R�l@�o��[A����Q��2��)���E�q�O�r�h�_�Y8�r�q*�NE�N!V�Qߊ	���+�	�v�tJ�]*�IN/�UC6����}M��<��uxB��:t��b�]�o����Z�dȱO�B��8 ��@?��-�i����5��|m먯��8�$K[�`�̸�D��i���ü2[U�Y?�T>B�/�\����ӝ��N�n2�Dq!�b�?�2��6Y¸%�����G�d��:���~�ǽ#R�wq�i�P8��_�0}4����P@?�G7GqW����;U����+���ȋ
K_�]^A[C;N����B��co&�| z����{Ǿ�$����'�_(��f�s<W�\kL�t"c�:�.S�l���]Ymь��?0r@�`S?R�^�Ѷ�L5��D*8���Ҕ���i���P4&���=��;�p��F�����)���!�s�@��q��\"y��_	,��U�:X (��CIq�����)������-���<�� �DM}'~
�u���.Zq�;��/G���o~vKE��^�5|�0YI�\>�A�� P��WȢ�,#٭R�S��=�++��q𱌘6zk9�|ի�`�C�+�" g2�w��-�h��|B�;�U�R8��ƈ�u��_���kwz��>��zo)��o��c�D�{��(�
ߺte ��N&*�U4�kn@���.�����VTE}�E�������KT�J9����H|1�����j'�J�g�/�Ͳq��W(��!+R�R�R���'&:L^�X��:��0EE��7U�CU����4�H�B�K�o��4���+��%���e��D���ߍ��|�Q��A��QV?Ne������eX�Ȑ]�=�;/��I�3ky+c��AY�v-����NLޯ��h�4XA����k�b�p�iZD|+p�\_6خ�*I��YZ�֙�4�-pfm��������1���֔>%	ܨ5�k>�)�e�(ŕ��+$��v=�ޏ����C�ͨ�QG�}�M��v�&�.6#V�BC6����ɖ-9�( �#�+��s�˅(�a�M�\Ӟ���S�xM�٫,~�T�3��	�t�7ز��"�>�4Ԋ�`� 7j8���y�əh3�mDdֳ�|.���(���5P(>,���յ�[������ج��/:w\n�8͛rg�Yw���Apqz7�CE���9�M�Z�-�k����`�E��w��M�R�(�!��t�[�'��J:�b�]�[=���>�Z�=�����5qJB��Ua��#k�e�*��,��>��S[oO�گϽ_�L���,+�B?k`�4�[���̣4�����ւ�4V�#�&���|����O�(�Ƃ����O��S�n�˓?���,ږwa�L[}-Y<�=���Հ$�|��3�޲x��~ �?"Jɲ?K�@��6P�E�j���^��
�7X q+�4�iL �Oi�kz�1_�
|����k��He��+9�����*��f.���L�c�#-4e�͌�zG�Ȑ��vh�	�����|���&�W�މ��<%6�ÌG`���he;:�6�u!���
�zaZ;��a�,��]qQF�������ԭ��tn �l]
PMڎA\�بi�TjG�U��eu͞ �jJ0�W9������{�(_�9y����z#�r�U�s�JU`l����/!6]j�h�SUR��&(;�=PZ�"�݊Gȱw�SPg�5j�w�J� m���aE�&�������J����zK/v��?��ڈ�ˀ2�̈U��H�0�a�k�b���d�՞�Ck�4����?:�5p�*E�	��nl)�ų��X������h�@�9�j��biՋ��3͔r�����1%�wȕO'�1�� ���y�|�0���5���XܡyU����,��gO�D1�����Puׅ��Μ�z1ףƊ���<j��*�e��4��\�<�Ȧ�lFxw�O�c��������������X�ݮ�dk<r}�b[~��a�S-R�x��/��Y��P�:%ʢ�3���P&�/�8eخ?�ik���0��$�D������l/O�4& Qg�j0˴�YH*��r�7�)x���S^����Q��y<-���z��@)�}}1��g� �)Wm��;Wlr��w�Zh��&USZ6^������fC��I:>" `j�y>خ���y���rNs�I��G��_MEZ���Qǝ����B��� m���+{�4>*o:1��A�57~*X�� Q�E[�Z]{�X_�urO�Μ2�G@��Q���e��)s8 Ӛ�N��u �γA �l.�g��x����=�0[g4��O���� 4 hO:��&5�N�h@��l"����������A+�u�����;+�G�����d��Jg�اom�)ܥ*��[w�����0��ߓ���Q_�=K�����̴S0�i�U�a$#�yO2{�G�TB�,��I+�=NN�U�.�#������7���nUFv�Y���Q�qz�������;�+�ۚ:��Z|b"{�Vױ�LV�	��-r�_@st��=S~D�Ғ�9�Ň��d�泥rE>�)7P��^S��KHW�x`:@3�@�n��g*�|�ߙ���˳(��>DK�eN_4�^/OB�=�c�.���n�4��_���!]
�ؒ�,��Ƅ�Q��2���U���F� �`�D�Bۈ����+��]�l,2���&� ��!��AϲJf��JԵ�
�M��AC���Ț5���;�C3 Ke]�6���E�V\ߩ�~�?�\�:d�a}����&��W ���
���ˡ���U�k��NM������L�ԂΚ2�I-`:�����>l	U�}s����#�2t3E�	G�6�����A H��1����7s`7�=>��A�jwy����b���n��Kg�dr��D��sig��-6�<��$ޢ�k��Z\���D�h%a����H@��%�lƙ��j�+���YF�4���"3Gu���Iܶ��	i!����෮~��aى��� .��S(b�[))��
��� `�&,;�R?�+ˑ���ݼm���:B��YL���7�#���S�VhV{�T�Q��Uu��'s��=C�H�l<��8�g~K.)��U���1x/�Wt���P������J�Sy/��К�k~�@PB
�d�բ�a"pq��@��ӛG�Y ��#+�X�Z��������z� r���)�%��~:��S��ԯ�bih�]H��^
�.��W������	�ff��D�p���G�K��@������9ߏ�9��?�Q'����8�ֺ��Dj!�q�3F�B�`ьzY�=\&���Z|1S�L����z����_e�G����g�<f��M�����I��i��qa	�of�� ��W�.�k��`^�Ђ��H�b�sl�gǏ�K�{p蒅t,̓����X���eà��b���}s^*��g��z��Ki;��J����Al��	���ѼF�R�f�]D86w�E��x�L�l�ݫ����4NBuï�$^|p=ӆ�L�u�TYz����-��!�0�.b����{�s��ݧP�<3�p�?���]+6������O��Q-��v��r����Y�ʨ��]��D[�ѡe�>��t��(_h��چ��cQqI��I�k0;�Zp"B��"�F� �#�1�r'��؇�/KQnzlm�=�
���5,��;8���B�)��}�c�LpUp�;��c�d����I�������O���F�����~ZZ�!�f,��x�㐵��KX��+�s������:{����-����x�Ir�Q�M����kܒ����59ѽtBh�'��IXP�=��Hb��g�*O�����!����7;%�=���)Ć�<B*#����+\�l�3���~3��3݆�G] �ӬO@�WJ0`.Z��l5Y���G�l{����4n��.0���؉�Jx<�Q>e7��GlK��O�R�`�ǌ�f�U����	���+����p�!*W���Tim�^��B��1Ӑ~^O᠕Mj!l [G��U�����`�-?NPo�b$s!V��؍rHp��a\(�����(��	NN�Zƃ�AG �/�iYhA�L���K�S+�`6Q�çfz8��7��6��ZA��Ɋ-�)�}#uQ�i_��y�~[�+�������-|��1���W�@tʏ>X�������A@�w�ˤ���4�G���=���?B*C��
w=�U�c���{l�h�=\��K�U�A�t�F:����H2x�E��.���c߆�[ Š��49�ݶ,@��y�Tu���Y��B��:�	�،�gӒ�G�/�>�^w#]�:�ʇ�#K;��E�f�یy���1�Ⱦⴋ�)!B�ǚf�샠��WTڒ��Ӎ�6�١����m�!�-_,W��Y��h�KN�%���׻�Bm �Tӯ����/2;H�S͡"�`e����j�ԃ}zE��n��6�W�٦�&�ľ�"�;�d1Jq�םJQ�?���1���H�(9׾vŒ��"������{�X$̽�FN��t�H�S<*�$�T}�*�T��Y-�r�=u��(�U�E	������&���K���G�j8B��- �tH�"�i{l�����Bp�aG�K</����'�)��ﮅG�3:�,��&�D�il�0��������(��-�:5����A��N���0�5yQ����e��9�)��a���Ձ��ʷ�ގ��b��1�O��;����/�AlK|X1��A4�A�<��Ik�GWkT���
��,�@��)��n$�7�Q�x�7gYE`p]˚��rWv�Z�Z�" ?�"����qyS��H4�j�^v�F�<�W�N�˙�������	����>)�7zKX[�	4i�lUB�L�̇��v�5;=(��VJs_a>)Y[��/�/稫�)����|g�9KA�e�M(��$�>����a璉ʅåp��ST�xX[R�r��z�0߰sR��k����	�3���|/�U���'���I]W
�+p[^e��>�[_��Bc�JuN%��O���)3�⃜W��pO���#g��v��p;w��0O�@�}�c��c��3��V�u�ό'R,�HT�'��ٔ�F�;��?�������B4wܗ���gqZ�Y��Rw� [ܖc��QHwo�(�4F��O�S���W[��m�=���]�-f���½$.�t�;��8��~@�\m�h3���c"a��������H���~�l	��WDF��2�E�q+�
o/�\ZSm���}>�*�k�ڹ�_g��kQ�G�ل,�?؇w~�œ5x�]��{)��	��Y�&t���i�X��!� �$���b��� �k(Z�;�X�!�F��>c������0���o��#�(�3��[�G|� ������p��@���9447]�e��pγ���;��)vs��W�ͼ|���������n'�\PQF-��F�"��Cg����ӟ���)y8��?6-�hW)U��3@�@x!Ǭ��2n�%�g~谎P'&P�6���v���k/��xXhP4��
j�?ET�a���r5�4�e�4n�O�IoH>��oX��Mj�|Z��<����^R.��7ꯀ�����-]=]��VhE0���
X��JԤ
xA�����0��A�րT��h���xE���ZC����Σ&p-����3�X��:�̓�I���V�UO���g�R�/f�&�s���ˈ�iJ���@@rǒ�ĉ�ڬ�H���:XV�0�B��+���$~N-/,�@P��k���B�]�cO'���A��v��Ե���T梫kJԠ���ZS��n�'�������+x"I�� �b�d��=���9G�=J�����P,��\q-�֒yg��4ϡ&�ZMK"�׺�=�=�H]UJ���=���
��w�K��9�
��n�Ҷ.JP�����yGU+�u�ާ��a ��I\W2W�%��dT!OYbEa�^��;�yK� =V5���Fgi��l���K8a�cH28Ѐ�R%Y[��!�,ښ�h��&)���gX��Tw�>��4(��A ��g Z�n&�:h�XY��&vD;������W1��':��Y%֕������k9�LAǉ��/�k_%���!�WM��`^��3��*��k=+U��^y�u��AI�k`�P�쏣���A��'���S�D*�([�,�j s���h�3Il�u�B��:��~�,_��ћ��rӄ%������B�*2�$�G�G[�`��8|���2�	4�j�&8n�B�6I8��� 	EѼM9`�_�Vf�t3�.1�p�kP��rل_+�
8y��=�VX��L�����{Hp�a�y���0x�Ա���L`�sP�jsj��?r��p���*"L��M��@G�+�	-5�:���lAz#H����)Ӟ$��.���0�
�� f���W�h�c��@'�@ӓb<�)a.��Tո=�X���F��q�X�<r�倳�\�uAg�O��S��M��� qJ�S�u����n*f�[iN{��� �P�oP���g\�]�@U��w5�2�AN�tD�*�6��=�>nl�Ll!�ɦ=d��7�k#7����|Pw�v�Ҁc�S3���$�Fj�XO��Z�{�|�'��(y�hȁ��5r�_8�.��)�E�
��s����}S���Y�-Q�B��>�!y!|�S�Ā��b3�����|��.��˓)��*��\��P!�oE"G�	��wN���3�m��7�Л��<�X��Φ�u滛�*ə����SC��:�6�R����^)�c��} �F?�+�#�â!6���LR+��4É9�-��Nʛ��Y�>%�f̞��-1�J\r�p�A|%�[-JT�W�ϧ7�Ԃl�Ak����%zk�*F������b���-���w]�!�[%�6w�]��H*���7�
�B��X�L��lj��`�T�E���~�F���a�;Q��V��־Ea��}Q5u��A��k~��e���K��b$88d��l?�S~��%t��Xn�0�	���&7�Y<��&aA��h�.HMC�D}
k��fXfL=�k�I��ց�;����"0���B?��Ju1��ۡ���(7��8�����D�,���/c���7KӆT��bo�C���fR?D!��g@���cؚ���!]5ð[��*��^˃�ԉ�4���5(�������'�!�B�ibʎ�"J��8���(�c�K�����(�S��s��+�]�ӃL������Ĕ�v���Ԏ��U��0��)�q&����kҖ�0 �9��	��굶��)���� �𔀰i�?wp��j2P�,��S��wN!�
���W���]�&��~�I}O��Z����G8���H�Z5g������gk�o��!�vL~�u"��I�Q�5ҙ�8m4kY((�	���d�hV�L�A�l�J������r@/����N�V��H{J�+��ѷW��K7f��X� t������wW��6e�gnv��ܾ B�&�|�RԒ�"2K!g�P�?]JD��H�C��o��Ir��`��i�!���K*�ne��������9ð�ek��8C��E��0fGu�p;�@����Lb�?�|e|J�.��7��#%�F.E�V���)��q�!ME�1c��q�Hߒ��.���,b��"�=�`-=�Q�"M�r����`��rb�ݱ8�e�qbx�*u�V����C =���=p�T����i��X��&[��[��MM�}H�������
3 JDdrt�٥�/�h;��
r��b�}L�iZ���f(�����.#�ᆴ���z�v�G՟~.��[�g눩SUx@�l�
�m���U��Ó��AA�Z���h��ڔ";ڿ�:� �lb�&�M����_H{�r=B����C�rPܟ��ΰ���*�r���~����7����u)y�l�f)�\�ϕ��^��S�YsG���(/Hw3(w^�o߭OD�q��lۉ��-��ɸ|�	B-c"W|R��Pi1�\S�v$~��/������%�����:Q�כ�7�
w��@��p��������?O��(+ jK��ϓ1R=�\%ђ���+jf�_�v�	��,������^ʖ��ms���fU�ë�ɢo\��x��H�!�۱M�����?���ΟSu��YYW�k][�T����m�Ϙ�e�����V��0�4��,[�mK|qgV4S:��ƠN�y�*x�Ѹ$���O"WlO�QB!@H�0��7��,W������Y��`ѡ�A�þ(�4�76�>��9x�����=�U�<��{ux�A�x��Jwz:�6�E7��}(gzi���
�1$/c��žHǟ-@��~��������Z��~��uA,lV��͈)�y5>і|r�̒�3 ��m�A�l���n�@:J���3+��-�����������d}V6%���x�/"�þ�1��߹x�΀%��Am�l��ڰ�"�y�M �ݹ�։�3������mp�5gw��hWM�(�r?�������m1��*�Gt��������4��a�p�����Z�t�Mn��g`���Y���]|Zq|�e')i�\W��VGC���x�Is���2Rf��A(r��W��erv��p�X�h�-4�j��Oi��M�hVY �Ճ ����Bd]�Nt�A���e��
��~V���H�͡;9��ɾ��,�_l�+Swb� 8�K����x�q��4$�ϒl�`w�=X��� erp��!OI�Yc>^�Ȓ����*���*V?�Fmϟ�B��8�4�@&���}�T��Con��������e!�,�����L�K6x�*K���V�R��������cM���;��T�5 +*b�naD����Ѱg��c��!�a|5��c�����A�mX��ܣ5�1+���{Sں�9�=9�~d ��#	�*�<E�,X�pԳ���
�o���̓HƗ���![RN����N�]���'�	�������,hV���6�
q�=� ��L���L�� ������)�!�/�g�<AhX���8�!��<]ĝ�������-¨�U��g��h��Mk��#&�P`����w��a����[�j�`���<�Y��G�c~�өY�Sq�^ϸR%���kU���_��Sl'i)W^g>�/�o�[�Xr������ġ<�&}ڰN��t�@�pX���#�.R��&����9	y�b��#F}�$�eΈ��{�L,���w��dø\w�
Qѧ)�`
�n���G�ޥ���3GJ�r_:\�<��x��s}n�	��8[��c=a��H��6��#��lk�1���¢���o.�M%�z��١إ>rjW���t"�V��w٪���BNT�l���c�٩�6�>�2��Ck��9;�A�a�\o+���^>�>���ׄ�7e!���Q_���|���1WzΑ�Y)�@��?����l�9}U�R�\�?� K
P��/�T��=J=��2I���C��S��됇QO�^�ˣR���b��/�j�b�����u�Bn�)(���T�p5�I�	��M'�x�k6[* Rq;�;���kgyӪ�)�RB������&ѯ+� �Q��oe��u5<A����Y?�����H'YM�I�g�!���< �:8�̱��+6�I�ܐ�i�D/E�'/>�w-3E.�R'WH&��G8{w�k1�3:F/&y*�|����S��{W��:��%ݓ���F�\"h�$=��H���/r�ft�hA��8_}�$��h X*��cI�dgo���5���5{�$��L��wj��[~�4���3��� ��)�q�8X��䱬�*(������D�W՟�P󔚒F1� ���7����@���C�+�-��;
�����s�7�K�d��B�c�)/���@U,1�<�&���E��ؼ�JeCh��l0+����C��ÿf�������o��M�U���1��\+?ݩ��c��+7�n���%�i����kj ��^���Q�h^0�7�&��;�@���C��}2s��b�*�=�ȓ�jErQ��x�̃]^���s=�w\��_�j���EeCID���K�Em����-��,ӆe0c%BӠNE����i�m��s4�g�B�ڃ��^��EM(���r��(7�� u�>��]E1ZQe{W�"������Њz�:�n;j���bn�>�@5�a��P!Њ�&r)��DB#��h���E#��."�s =�W%�L"��~Q�3��GAq7�������ZNU�qƨj'r���u{C�uGJ�`	���o�a�z
^�Fu^�n�$2V�b�(���cԿ��:�I/#M�
Y!~D�Չ'z��(��v�:^��k�`���$�9�a
���~r���;��~�`B���}pA����#���ﺆ�]T�{���@�'oB�?���5���
X�7i�}�����%�AҐ��CM�+@�.V��_Uee�?�"y�d|@;"H[C�19q�tkê�t�Vl�[u�63k��jM%��8+U-�5�y��0Ck��F-b�`�����z.Z�|v�YEtE�
Y�+xq���_��&G�%�15I�Ėʻ�/I�^����6�ED����ل���0���K-�66�缘�}h�!A�J0O%6)p�����@\'��#�[�h��g� �%��V���Ncq%�&~B�� ß�閾�ũ�cy��
~7�]c�=a�y�!a&	�$�N���ZR�Ǔ��$~��quA-|O�Tn�ࡣG�	�Y�w�Ŝ�.J2�-Z^��"P:��ch	�+��u��Lu�hL�E?/�O�9qZZkn�9��X�Ɉъ�ە6��\����P�p�-Q�v5�X'�=�d`��g���We�P���ڱ8*qZ�|]S��c�~\酿3�@͗!m<�FyI4��
'�Ѽ�U=m�/fч�,PغL@D3�������'@� +�z��!�ۚ���DǈS�l�}x��vn�7t��"����c��d�K6` ��k[�%��X�ϧY��B�����惛ߑ��(m�O�ã��":��s�f�X:���#�$5�����S�8����´)�ى���!�.�N&�d˒��Kd����I�n���Y���ԑ��:&F$�%�P��G��Px�q�Rr�]+�5��t�(8�-ڦdK�{�b"!)��!�c�.#���6P�����ʩ��gS<�͎+�옠2�����u|H�����d����Z����/ܟ�<�k)��#��t���"pX�]'(;4�� |VZ��]xgI�h���0{���㧆W�'uͥu�~o�����eJ]ڃ9���{��Z�vk���V�̵*�_�h>��z�,�BQ��h�$AG�x"�ú�@;�C�Y �@ɠ&W)�uH�d�����׳�}�Ċ��Q%m1e��tWj�گ� $H&J�ԫ��~�c(��߉�3���@ck�B,&fj�
/z�1�髧_I3��Aٸ ��x�ʴ��i�EE]����G�,��ܣ�s.]����KP��U�w������)6�K�v���P��S��B�ꐙt�YXb7��̝b���+sHz�@:�!���.j��Pؙ���m��1�O��s�=�o֏P�%S�������b%�Ze߱Ҡ�����[�@���i{<U�(��['����s��3���ho��4$��(��a��1ٞ� äĖ�0�{�����oX�j�w{A�%M[|JÝ��g� ���Ql"`96�H�z*6~ ���[��cY����%Yc_���,4�3���c"�3 �O�
�p֭���#ٓ����Pz6��}訮�����W�u�+�X�v�Bۑs`^���e�
*��O�dT8��w�[}���<=j�uK��P��@�;�ܶ�}���𾋚��H�kq /�e^E�UqwG����䤥`�|�7�y'��7��ZZ�8aISZA'�ص߿n=�ݩ�pK��P�P�<�ɥ �&x+.4Nޔ�G��eM�K�]@��A�|�i����]�_uhS��+	�Z�uዝ#OP�����6�p�I�O&3ɳ�m��6����ua��+�{�J��X�Q��2�"e���*�G��WFtGJ):Rs:�G�H�0�Л��V�}��c#��h��sPVa2ab��r��=i�ٔ�P�G-~����Q9��֦�i����3D	�9�Þt1L�r�^��*�s�E�]��Ҏ1���G1��m~�G1���!���4����FQ��v����9�U��B�@��`���.>�Q�i�~~�<�q½J�z2^���b�8<#u�|�T@>vӄ�,a��=L��� ���M�F�� �H��u2xw����μ�k��_c�~�Tk~K�����ȏ��Bodo�u���M.�Z�U����7yY����6�y�f�=D�^l�G�Sӫ��*���E%ãx��\b���0V�q\�uUu?�a���J��%X�7!�FM����s�w��h��CQ�ym9��i�0�q��$���Hvd?�	�Q��O>�/�D.��$V��������k_UQ�'�h�6M4S�Һϻ=�ʚq����w!F�Y -��\���b�g�6�"�tHoC�"	fg�0��L��Q����A����t!Fn=����ӫc-�9.V�}K{@̇��ʻ��Q��K�8� S�UO\�`b/��`��۵��j^ZU��������o����ܘ��!�+��m�N+	�"����%zUAc�$�I�0S��Z�W�p�Ae"��9Ed��A#�8wxG��&,��`����zJ-�+ѱǁGݓYmLY�t{�+�A�:�[آM�;�Zjpk�G�g��CET-��RP�$wc���z��W�-��"~Zv1��b[�h!H{�4��xZ��v�s�����6G��]^�&$�Q��-�*P^#�E٘��D����T��S�2q�o�	
�w�3�E��<�k��.Q��d�a)z�%�� �mS�h [��W�}�\,�A����\����7���~�~0�-e�	Q��� �<�H�	t��b���G,�0�G91�h��H!B����$˂��$=�R`U�0L2�8�)9FȆ
]F$�s�_Dj�^���ex� ���R���2����wU�xa��"Uh¹5ɭ	}�J�*�x=`�.f�ޥ�H���K;qᇝ�m�M/�v��H�Y|�p�;�}�M	�� 
���.��w�W��l/C
q�D�hpR��T-�O��
�Y�j%^S��␩�.On�	���R��)�EX�@[ �$�� �,x�Յ��G������1SŁ� x[�^�g�eu�����!��{�G�1�0���}b0�X�n�'><���N���w����]��#�)v��u!K��Ce�O��A��齱�0�2�G��~	ރS�g�y�F��)�M��!���/�βOxR��N��4����<��ͫڸB��̎��Χv(X�Z��z�U~��%؁��r.�
N�E>u���i��ab�$��H
��ָ��^δy_��eB����J:G;l�<9�	օ-��!��_@и�����#�e��T��~���z�Y���Fp�\NE~��'�s�Z��F����|�0�c��g����.iI���(lŴ�����J5�N
V��N�ë>�rj��Yn�!� 6�8W�j-��ƥ&��0�{�츹i#�����yq��#Qmy�Fڅ�U����IQ�Z?��F�6��q�Q0�7tc}^��v\[d��QW��b�'�[�z^	g�E�Q�Ɇ��K,��-}������ �*�\}�1�{��2X��'Œc�����9�^6���u<_	Qb���R��G�t,,�/�l?�/�T%�v%�D"��i�#�ʟ�B��U��4MY�1Q�wTA�^Oq�Y����9�'� �<[�^JV84��`ti�|�NsGA�U���= _Ɨ���@x��e�"���Rq�|D���ɇ�ZҌ}���X�p�7'�K>���%�Uڇ� �ED��ġ�jd���SX�%M2�0������2��k�՛�GC����K�Mұ`��}7x�.&+��oڊ��U�Vf�q����q��0:�tޏ�ub�9I&]��_�fDFB����q�g�I_5I�h���r=J��YX c5������T~���=iB 5�UO).��y��f�ԋ
�캠��%��hݕ�����J���_����`%q� ��֔8��
c�f)�ֱ1�L�yC��������1����>�7z�Īt��%g������ߠ�h�f_�ǄO�sF�Nۛ��G�_�ei�ӻ?7��-�[��o������6�Ι�K�\�۬?����53���jB�R4��2E�~���c�� P4��t�@K7�Z��>��<*���h����H�}UEv�]v�{�{�;�O�����N�<�[��c� ����;B�d[�fȜ7~��7r����Y#'$*���w%w��:u�'�&�9��9�eՇ@.�KVD%�1пӔ<l 0l�Z"l�|j9Wǈ�ɗkE�V�[4�ȥ��(��֗2A����X��d���lm��:{}����ʖ鎕���	��&�ϥD���0b)쨶���Zw�{w�Nu&�5d�09��9M�%�\ej�I8��:r���UR�|��t���a��)�G#���?ݡn̖<Ͻ�p���H��4�����n�6�o<F˖��)r�q�^6:� ���{��l��+TL;��	��L���m�=����hL%4݁���N�Fu�圂��Dh�T��E\��lF��]/��M�B^�ᖚ�o�������`���ae[���s����$����S�t�������1Z^��L��:���,��H���f��ؗ�#\�`��&0���2�a�0ؚ��4�I�UG��L���uu�K�MO��d�Nz�2�e�6�zw��ݚj`�;�A�y���(��.wV��7*��n3#�I?�1�&e^C���)ܓ���]�FL3�d�r۴Ԍ)V���&�Y���m�rΤ���.���c)k1��׉O	�m�������{�8�&��*8s����Z��ʸl���6xJ >\���P"�y�f���?������#��Xl|>V��	�*����O��&qAC,�7���RB�]0��"�$D��w;z��tJ�HIU�t�-�&F授����ERB��ez�7��E|�@�2�2.v_tV�,U����C�������������9*�G��� ��ev0�<%�N%�Ht<@+�;������[5&��<���(mLGGcR� �/���D:�����\�h����I��<H&3�zU�)]Cp�u^V�	3�k�»�VW���J�i\�sz�a��D�=���ՠ���j%<��J�p��IHBi_��}G�����|�u��.C�SÝ͎��fW3��(?���H�U]*�+�<˳�
���n{�!�)��U��a����0����V$�̨ ��-��K�N,|#|�b��`�,%>0ۑ�4՗*ޞ�rL�������P&��� Lhtt���=�l	���Ɵ"��$pu�I.;����(���3M���͹*�+�qWj�%�z��>�K^�$�'D�o4]'��=�¼PhBn\��)k����^�����rQ~=�;����|ht��t���"Q#޻����y\xh�h�j4	*�n�ﮥ:i��dHYd>��Z��8&�d�LZъ�]�ǻ�z�F��6h��I	��ѷg���vK<�Kt賒��#|r�@�Tv�WH�F�	D�M�����2gNT� �;��O��r��S�Q#��j;��{@:�,�=f���i=e��q��r8	��x��hvhPh}�F����<���?}�t� q�<�+�2ˎ�;�ѫ���`��9��e�9Ȃ���z�V�v �6��fV�P��&���T��+`Pn9s	���&B@�MS������i��fW#t<#���XX�����pQ>��%5� �Py3�깨�Ƈ���3��9�ÏO��߄����
"��^������q����\�jj�Nv1�����yPDڇ'��uY�p�]�[)/Y�y��&K�8-8kBW��$A�#�P/�ra�u\��un�F3�sE��o�s9վ"���`Y��υq@nu�|~"�no7�Թ�����	0O�L��3��\Q������� ]�3�U�PfC�ذ��yu��X��_Iv�rfiI�&r�^����;��Ln�^ [�/thݣM"o&�)R%h��)(fq<�GĴ{s`E�5Vr�݄@��YO�s?Z�߾a�	o�6@�� �-�\�QҠDL^�<3<t���=�$�FKg���cN)'2Y5W�̆	�0T ��1h1�qJ�)���6`�]���x ̓7�X/-屌Mg�A����I�-���/��c6�R5��(Ȅ��<�uKga>j6��J�S/�5X�vF\��ך�|�6��X>%�^�W^F���y>���Y������ک�"�/,�Ohk2ɝq̝g�陨fj�L��u��0���d�$F	Qͬ��r��u��+a,c'M:�yØj䓯�Дާ�c��lh���G��B[�J�O��oN�K(��N�;&��dI ��阡>��� ���ݽ�A�:��®@�t�KyF'�k�OU�Ӫ1��p���+�% dp�C�}����մ��$-<QSZ���Z�Ĵj�ƪ�6���o\!��u�b��흥��u���緆¹/�����b�-�N޼�Y��\�K��+/�����)�>$�j���|���D��Й	�L����Xs�N�V�Ԧ}�fD� ӌ�_p�A�_35\�9�ؘl<ߪ���?��a
"�F+�%}�0U �)c��D�3�F�,�מ���X�M��uaeRo���<�|4?7��1�S����˻�T�/\��l����֤����ЂY�5�E}W�����6L�խ�&���A�Yɢm�p��as�2"��3.��a@z
�w�I�K:��K�=��f=�w��3��Dmo%��QV��S6��ce/�lay�uY���-�!GF¡�3<���Et?��]�(�=Q�/Utw1bbs�l1���'rSzH߱}����c�9��r���uj�x�d������'���?sԈ�,���˘X7iy�_5E�J��|Z�C�旘�SM��*��Ab\\C���@�͜_�႒��y����iF��
���$�CrZ��Em���wdK/�8Q��
*�d�	���E!+6��Dj���e���l�\4��G=�g�`W��Q��Rax
�C>-���V9���,T������ >���r4dY�F��� �m��A��֧k�0kp�[B2tV��|�z4`�~�"�Sp�'Nm���^g�~��1���6�rHo��Z�q��ь��<u�'���������,u�����G�「�n��̥�L/9F�v@�S�C��l� )q�H�������E����O�`.2��62a@n����1�����33�I�f��S�DB��ZζėI,|B�2��1�b��Y3��s���&�վ��S�t�bϷ��l{���0/�92Mq?�V|y�Z�{�'�݇����;Ddi���j�j毋�'%����N3�l�7�����T�g҄fpW�B[���8ٳe6*:���$5�J���%��׵פ��I{�Ѐi�i�����5��@��ܕ����Q���܅�VCb;K����6km7ל�Z.�"�dX�C�l�hv[Zam+�H�)�@O3Ձr �Ĉ�l����!�+
�&��
�ԝ�![��ҟ<����H���OUgx;�3��t���{���2�J�qӭo�m���F�r���9�.�q:�=����l>"y��6��D�j�5_�Ⱥg��v;�'�"�T���r'm)k���B���kq������v �]WD�˜��%�-�N��5*ܙf�j�Mq���<e�����je��q�������' x�p1}�����#�c�-�{��ܧ����J'�����',{)�����g6��{#c@?@?%���52*�V�  3���y��ή��4����Ń��1���\R�$�]֩?�ͳ��
u}���y3�<W�2�)aS(���Jb~�m�$��:�C��7������jY'R��s"�K2��<E&�NӍ��l0��ڎ�	��
r��xO��Ԯ��%�Q}n�Er��W�]#��H���B���6�PQcs�mo)�#�Ç����T@�M��2��6�B�T�&m=���Q�(�s��� �萙��5����1�̎�|{,�נ	��+�:#��]xߢ��E��S����-�YH?�t��ynd� �$I÷at��]����|���/[O�sg�)ȴ�$��-��H�_�5�6�Cy�=�ṉ�ݯUI!5�9~���w��G�Jn(��c�_y���D��+���J`�ԺRJ����)|$�O�ʹ��V�G�;4�����/�^_���%����X?h���|�\9��BӲ�8b�-�DŚ7�=6���Wm�)���-]g>���i�ͷS)��5x�s!M ��k�q��Gs�9��y��Y��CZ��4��x�G�����������m���{�{�&�(z�p,�!���:{���>���Z��HQ
6kԦ�~�-.�������|�C�R���os��\z)oq� X+����L�P;b����4�F�`�_F�6c�z�ט��~����=%�RL�R�i���.w�W���ϝ^%�ܣ"Ә�(�̔��l7XT*�>|𢥌�=Y��-��c9� :�P1x��%�� &���6�^�M�;��B������LS<�}��;���FX`�3e�o�vtf�O9)=�����=�"W[�Z�6��p#�0�Cݕ���\��Z�qhw ��Tt2�Ih��;������X���pv��ׅ�O$5�}���S�Т$��X��U��/�0��5�����2?m]���9�P94晕Z������َ�W��I�m���z�|pG�W�Բ�D�Qt�b��4��j`��Fx�Q�g�o���憐gT��	͛���d�og�U���gN�Y��$�d'Nng�>aۊWoT��Ӷ!ZV1����F��3Z*d��k=�����8~�4�AC����]�38�r#�a\����{�JDB�� 7QDf���cQ�S0zF���ex��2�r����|E��衻�^�/d���YZ:>��zr�VF��ρ�(�4��M.^�˗�, ��MM"�r����GY�n2���q�8���a�C��x��~3$�||���!��w�v��
�/P(��ME�{Jq�Fp��FE����R7���͛~^��W	���/�Z�R�&���'+1�#�5q_�ku����h/���<���E q�ߛ�{-b��AH �:u^�hUU���2_L�Ju��k����[�N`Y������Ue������^��#O�4X���X.��6x�4W0Apg�%�a��U:���.�s�aBT��;%�:.'�ġ��
��0���ôLZ_�j]r�C����øU���6=a����H����q]��:��@�B'�?5�%^W@0?7��gE�71U�䊒��'4�J�^�}�$�fq���״,��V�����C'�A\�ZZ<�R},��_�>�hi�|�0*�C�lm��"�����]�i�����"/��f]Z��4A�=XЈ�d��W�;U��P�9�D��:!����?[#->;?���o�[�$�1̐��Ţ��Oh��Q��3��JX�m_��.� K����F�"j3��p���O����5�r�2��I��:�}��/�� յi�#/P&�,�]�βn�g����oC_�Q�.&��)	��"��AD ��ΰ���k��恋�X3|s�"�+8uU��l���9m�/#w��e?��,k��s��d���Y8�e�l@v�<ZR�q�vC�vQ���}����6�]��.@�D�/��g��-&W�22���2/wB
߆?���xL��˅=��16�V<M��3�)��`�H���u�r�[�'��tT� �2q����<?3´�ߜ�;j�d�u���;�q�=3�;��n�n�Aq9~��:7p^WM[��K�aА��^��t|qf��M��)3��Vˀ���=s�"Ȅ�+�/pϐ�z,�T��fh���?2��Z7�g���7�2���b/.1�G��6<_�:�^sZ9�	~!�@�c�5rnK�m:��{�+��`�W�d�4�����q��N��o~56E��!��Z��#rJ�
������{�"2أ����UVS�a�뀣<��Cߌ,�๫.�~�ɰsY����0��Pl�ͼ �r���(<�$R��.�?�4���#1�E�(J����%F�m��/WL�E�ۄb�&�3�T�s�s�n��t��Ak7��q^2�0^U�Ԉ��Dq�>�%��p�RS-H��!A��8k.�c�>�p�[��4t���&�K��Y���ܬ�K2Е�l��$����K-1>�j٣��� t�� �d��-���e���G��#��|dQ����W��2MԋxAכ�]YMas1���2r����ᴉ�Xכ1q�&)NW�h�����B���ŵ�fц�lM���>,ؑD5%>�8
�#c���\���ȃ灪�pd�'\*��/M�"��1��*k��>w���ܿo���猂 X� �R�Ƃ���;�Z���;��f�� ��t��a)��- H/�l�)���Xx6�E���4~�ޜ��_�D�	~�GY}ju�.J����z}]�'����g���g��u���2Gm;gZC�K��2k%z7�w����1	<뷝�pJZ�@�r{�~�AX� �1c�3�����{��a��ῥe>S�h.�z�X���
�ދ��z���ï�	u>j�	i����8���N�Fj�P���`��E�<��e���S"Tj��+����Ӗ�C�G�{P��G7Ǔ(�� q�G?��J+T��h!sr��8���¬�V�ND��0��f��{���ܾЉ���L��0�E c�N5��chA����,p�/_%��Ɩ���ϰ)��9$9�@����������y�(_��	k���7�gd��+}h��u��.V xl������׵b�]�Bz�>A�-*m�X{��G�[���_5�*t��h��zm��7��`����Ǻ%�;HyIR:�"l�{�� ���ݧD���r�}Hr��tڃC���G�$w"�d+��5�$S]�Q@_��,X�D���z�mB5�|��o3P�o�/, <(�b��"�*�.���
%�($M$0��mOL�o��Ŕ]�2�%�Y:��=LM�3�2���A?hsV��-e\�t�u�Xj&uo8�k9S��_P���S6Ⳟ��qyr�7�h��<��)c�܍��"���~�j��z��}�� {j��_4�[�0A	WEV }ce'����2��kYa@����ƀ��&���5���U��3�@�,0	T%̣�Fw�|����g�-�2�b|B&�Y�-[}��MZ��Wh��놦�0DSѯ��Z_Ϊ�x����J�̍Zi��b]�]O/�o�tTz�DpZڞz�����)���(� 2�� ��،d��q`��s��Z7ՉU�NQP�<ӟ��}���ǜJ>/�8�/�����Γ^!��m�֍��Y�Y�	X&%�+����-n�J���n�in�QzgɖƝ�֒���2���G�D��������C:N�g��\����<�;p)����m���#7߶<�N^rȺ&�v���\�f���I�R����&f��:�l�!�1�[���R0�Q���e�@����b���[E}����R~���g�����0*�{�hJ��V�U���4(��1���/���;2"�ĺ�6`B�h�TW��GZ�����E��4Zm���óI�R/5z�-�a��kl���V����sOHzՋ~Mx�1@Z�"��j�g��e���F��*c�U�U�x�߀gb�]��&�����0}``�M�	��l5�N.e,�%�s��4t��<��#�M��.;{4�x&{0�0�6̪[I�r%�5�"�p -d#�Jt�����T����dK2&�:��\_�lEN���/g��m��_��N��|6�!���-F�"m�،"�
�H��B�xH�9Lv0��m�������
̞�u���5��{�,/;�V��l.��2ۏ���9`�./����ݯX��1v�,���[�JE�cW&�i�ս�����d�ߴ�eɭܠ�H��̉�n0{����I9t��7	<�7I`p_��w0	�
��]��г����9���x9gM��Pv9�*�2)��~|����~���\�z�@����
��N<��ER�6�5|��Ϧ�yR���*,���N�'���Y�#�7�W(U�N>\ �m�f�+V@���#��D��c}eȰ�|���d����fg�JI�y��2e�C������B��i�2�+~0��dq��[	s`&��������gbD��g����l$�ӽ����*�FB����8a!�
_7�K�8_��3�V\�i�8�]`Ӈ`�5�@�y�8�'
�@u�J��F$t9F�b|!�25�^ ?���3�q�����4�prf�����t�*���#��fq�?��ܔ�x!��/�"��B�EvJ�%"�Ekv1ڛ��}o����������r&5o��&N�������>������;��%o�&Tj����:�8��+�9"�НA�&�Jf�0��5��J"+[Y/�v`�'�ۑz�큪�x�Ԑ�	�a��S���R��>BT�}�V䨮�d-����l�r'��b�q�w؊�0G蟻�!ɁÊ���?͉j�ji]R�x����ᝁ�Gs�����,ތ�Zi��z��R��_�)�뮿x	_w[�ڰ+�O.�H��������A���ö1�&�o,�ה?/�B;l�)�>i
˅�� �9��8v>+��SO�y�$u1��m�8l�N0��)����e�}Ƅ�<�8.��!Ѿsuћ����l\���%zgt��"��Xt��F����I^L�6��˳O����Y����`Y'��^�Ѿ�xL4�`:�6;C�;�|�u�˔�}����.�������ɶ�b�p��?���ބXh���!��� ���Y���j�ͭ{EzU�+��Hw'������"�^0`΢ b�iOտ�_� �F�z�Q+6�wԳ�ך��w���{Α������� ^������}6*ܪ]R��p�J�� 1��y���5�a���u���$́jUB����#�c)g?�hF�G��i�Yj����Rُ������M���Ò�gO;�!�%�.z�` ԙq�������R
;�c�"������r���A�K�G�n�P���ա!0���2�JX�}��X�q/n����jkmXM���/9��(|�B�����"�Y�CX3k'9>��a'�#>W���;�>]�ā�` �\�t�A=�4<(&a�� �,�f��P�1R����㒘|���M+� -*������1��j������X2�а�)�N۴W5<�@���B%��$�;��������o���J�u��6˒�ߖ��Ma�of�5VR��)p�u�.p�P��z؎�d�3��! }c�C֣<�9"���%��_�+�c�d~r�w  �j�l`J���ޜcV~q����D��G?�㚉6{M��1r���V}�2��	k���|+� �w�at��8����&����y��[(�s�rx����Q�"ZX6�R�W���d��L�'i��1 �U;�ax��CF��>�v����ϑG�q�pS��7�P�-�^W�ck�HO0�G���q��-���d��X�N��5�;M㥉u�3�����Q��=�h���O&�sd�!�K#�c��|u��0w�p���V�k)W�Ǌ�ZX�<�¤���55����;�-�N� u��Rp#���8�␋Ea�|ʞJ�׌��J��vQ����P���'��)��B�)�B|9�A�n�9r�~�BYfF3V��2v츶�fu�+���������%�A�!��C��q�ýo(չV6�)�+ȗ�Wȗ��f!�۹jp^˨�V��w����81�e:������2��a�ި�\�u�0A�)��dIs8�`�K�[�{mcL+m�� �<fG�^��O�M4ǲ�#͌v���])��bs��K��e��[���o�%��ht����k^Yݕ� r�ϙo�;oQp���)EV2y���a�E��5�/k:>bge��k�`��ݑ�r����YD�T�Q\��mu�_\��r���}eO�^��v��R������g���%�v2O�dí���D�xZ��[7ڰ�EF�:�@f�쌱����*ĎO�zy���o��Y����n^�ص%����	�W�gj��~O1d�0ܶB��`n�ȫd��s�X)Wd�2�&���50��9��-$��b�LG��^��R����I�%z��������T��u�+f�W��&�`���{>�@^�_�`���G�#4�֠=��v�QXh���&wqj���88�/�EhT�=�C���?���HlK>XA�j����pM3����Q��u����n���.<:���,�(�������
�y	b��Ѥ~	���^��٥��Tv����7}�xwLp]{���^�'RQ-_�LT�LV��')&������.��8?�d��.ע촞b�����������;t���h�f9��q���ah8 k"��Nw���!�2���g�o����he����ޅ5yư��)�;������Dz�q+�ς��y*�:�^f�9�1����\� ΚGѫ���P�!��4�8ۻ�������A������}	�i��3й&�S��ү���o�W4:�&
ң��Q�pҬ��L5�&;��G�DԒt�ٯ[����Q|Ƞ֩�� `�UI�/7���h����Vx��6t���vN>.j.�X/�X~���Xi�����K��S�����}�/jf�Ɔ�n�=��SA@<�TLLgP4����*Ǡ�?�'��v1�>��WmbW�!�����S�ڑ����/�M_�ԅ�FTI'!��wP7�jť9�^�5��4�C�G�4�ˢ��N��)��k���-3Ç޺�L����|�6~�#o�"l1�9�8mӐVG{��߬Z<�}���c���ԉ���e:�$��-U�E!&��eD�Ɋ:ì�C�dB��`���lu��88(�`�# {����w�\?�R��$w�\����{}��C(���d�$�����oO�R	�%2�7�x��������/��p�ۍ',����^Ӳ�sra�Vј��jS�癌t������Щj�R�!n�9aO����'�i����:�� �5<���˅ %��Y �&���R���f#Bd^=H&������&��;tA�8p�Z�@�vŘ�uK�A��4�	I�A@Ma��![�S��'o<Nkjc�0��eä�ӚD�|��I���X��Pġ.^�J�X��H��`�<P&�ŎS[��3��{�a/C�uX���F��EgMϝ�bW9�#tu�mlkKB�,Y$#��L�V�X��F BߕF�[_	pY�}IP�T�ˏ6��n��&S�ZlgB�I�@�}��~=���]^��;R�_��G�m�����/�ȳ��T�Iٛ yy6����1!-#9`�@Ҵz�?�%t��	0ׯ]P��Ѻ������!G����5�������}s$�v�Vf¼!.���_Ċz������Q��I@�DN(�sj��m���4JL���>�fV�,|vt����4nM��q;.P�����J�
���;��2	�C�8Ɉ��
'��.��z��3��ڡa�1�D����' `�T��srQ��L�X,�;:3X�^E���Ņ�ʶ��[�,�X����b,�op^rÇ�R�]t\F�W�M�����aw�X��kiF��ܗ�*�k���r}���˔+��0�ѽ?.���E\|*1f�������m	�N���7�м�h�ZZ�x���ދOEб�NG�=E�� �Ü�Y$�Bs�=�SOCt��C�˩`�1�e����V.��g�X��3w��?�yJ�g���/��on�Jv�������D k�w��	�}�,��vI�ÕE�.b=���9|���L	�Q۴�����¿��~\�����*�N���+�O{|���!W,�.�_�%�/�\�_���I���z�\�����;;�����-�c{���AF�M|Q��8��yN�2��rf�X�{�>} �z5m�R'RLœ�&�/򐙋AՓ5I��Vd�@#}�(3��j�-
��������߆�_	�m�� 2­�iY�J��o�jpm�z��;]tO���%f68��$p�&���?�l/����͎U��Фݓl�q{Մ�J'� �cH�����}w;g����k�\��ڢx�����o���i���Ѧ�O{��h�8H7�_I<���E)RWTY�B&���j�J�g^�o���Q�{����_�BR~E� `�9xkǌ�5'b8�A�/Sn+(����9���9��Ȼ�Qw�#�O= /T��,,�]���Q��X�:��2[�ߠ� ���
��H���tCK�+��	��o�R� ��-��WM�/��&N�TkjtMS�c#�Fc��-|Sꦤm��� �P�:�#��^Y�����ۋ�E��FP�.�]E���iPN�M�On�����ǉV��][U��o m[�����x������zЇ�;M+���Ω�+�wv�t�!������,En��D�7��%;k���0�����e?�OE|���Kx�ܭ�-��tŻ�Ħ����mRx���˭�^ܩ���2EN�y|�H���x����A18�o�����|�dVQ����(iHƆB�62���e���k}��8
�����3i[Є��::��h7���I���7�T���N�-c�{��i��R2EWt�(��K��g�"1�b�h�;���kƮ�a,��3��]�+����ydOI�{r�\?�ɂ-Fn{7r�H��5��&_�9{���J;t+��卧�z��"-F0�e��z���f]O��x��{�w;�l�ј�X��&-��G��h`�j�/G��̺�\BK<zhMSζ'_(��q�L'���&� a"[�K�]� �~O^u�Y�7�O.�A[�j���c�]���:af�4�/�e�H����q���v9k��zBA^B����X��|=�v_
*�0B���-��u�g\�LF�$s
捘��4�eh�[v��U��C�&�xL��/��iK���w�؟�WQ�A0G��-jXZM��'}�d�K��cj4��_bBŏ�����L���Q8԰KF��\�yqca\�@ C��#�A�SC+���I��� l�$�@��D1Y`��9�KF ���8�t��@s
���.���ڧ�EWޛ	2�k���<_Ə��Nr��|i������Q�����Q4��.��l�E.2́,pIc"0��z�?7�	�@�Υ�Q�Ǘ3�q��.�G��Q��D!��s1�P�qun*ǦB��V#4�o �F8�5�2��wgv_$`���^���	{E��B���
�6T���6#_��R�\�Ӑ�=�t�o,`E)����`ty�G��߄ˁH����n�y�倌��o��(B	��ox����t���D���&RH�8��	턄Y�U���QA�`��^��Yme${�KU���"��1��㊶2,�~�vɐ���,6鎙u]�a ���u�dL�r֛��Wg��������1퀲GP��~+��v� 4�;�6�\�����8����'��,ؠV!�n�s��j+���Śe=�6���Z��YMT�m8��e��"^h��	�Ǻx?2�g#�f�G��\��;�e�>�A�^���wR����B�[/��U���#X��B��:,�X�=D�sϫ,�&2#T����ޱ\�s�I�}�_��s���<��!���Hv^�9�ހqR�l�Ƴ�D^8I�эN8~E:�w��J�b��9Ȓ�v)�˟�l����$jo��������d��RXuQq�f:ϥ͇�7{ܖ��Ɨ��Ϲ@]Z�h�����C�l�eq��hu���$�4���C��.��vC���+�Ҹ=YK�h��h���M�RҢB����M�gL�NuyE�������R�^ Y�
�e���)��]���v����9���)��ܧZ�h��?X
��ض�FC�A{��F�������D�5o��m�]��jB�=m$�G!��Q-������r#`~J�~6�B�Aƒ�m.OOV��\� 3���#OY�i�>%i� AC b�(����h<>sw2c�����>��Һy�3��;W�*�ޚ���?c������~�bz]I1p«6ΰ�=7v����K�=���k�?�LQ�Ү��g�)x��"�{$\/Ƀ9��������}�+Ԃ.�A�8^U˸����X9�B�&䆧�g#K�a�[�
��5Or'U�E�Q�*�48:VJ�H�9�z9wU�E�q�Yʘq�H2D���=6���J�7#��7�{(�i�MnY��;�.1;t�DweG��H�:��9����u��6�w�)����͕�\��Fĵ?����1�6���]�M/�/%dLA�N���5v�C�!�7�D���3QM���+��	�Z�������)`H�?���6�~� ����y�����������c+~��PX"�i&� �L��'CE�HC�Тc㚞J�ɯ�,��1~�4`�v(���"G��Uwtº��0�P�����p���p���zg�d�1����I�
��_01lScA&n)��tM<�
�4s��֯?'��ͨ*.�F�߹/N��v����,��{�;�'��A�~;��h_ �~3F�B�l�	%�UC�<]�)������I=*Vgyd�k�y.'�Q?����5��h�5�« X��s�X�E1U)���#�?˦�|{b��nuǊ�a�z��$+&� ��Ն�c��{��k�":c$�Q�V�� Tk%���\��=R٭ n%��}[���[Տv
[{R	�Hh�F~���H=�QI���RV��S ��Ђ�%���
O�˦k�k�X��HôH�J�>�G�gv�֐�:F�qj��X�T>7P�;�	A��mx�vnр_Aɑ"�_��b� ?8�#�M�m���]�f-/O��8:'�fO�m�[���L�����{��e?���;�т�'l������%~�6�-@� �L�O?��WC�"�&Q:�m�'&)�	���+��:9��
��ݴJ���B��a�bfq������� Yg�.�^�N��j�*!�fML�1�Ҥ�0q��=__�R��8U�Z�	�>��� �OQ�S�9r�ѩ�H��F��	��C+�X[��SP�*3v�=Q���wѷ�Q������8�=g�P��N�/w�����8�CQ�Y�~r4A%�.�����ׯ�4:2�L��7��i[���i����
4���[��&ɘT����W^n�*�S?W6[a��B�UM6Ǽ4ǖN���}����ܵ�u����N�~g�������gT��2��X��t&�ʜ9�h	G��/5�*HO��N=�Fz�^1�x8y^�5��'Vצqߜ~��R��0s��"��a��:��UC?h�o�9K�����_��2"3�7)}6²���#k���u�?r9���l*`�/���~7yvD�I���JL:a�`��Ռ��pI��S�51ioú�%�~�{l*���Emn�_d."Bq�UE�uB��Rb8��\?Pݍz)U���	��N���FFJGH Y�O�v`���������PX�:`ӆ��Ȏy�~8v� ��}�#��"e������,�e�na5ͼic8��E/�_���yE�����m7̏������[%y��T�ޚ��ݔJ�rF�\~��e8�сV�E�E�>�Vo1?���j�5U��!��$�g�Fg{fc'�!C+W+3t�i��W�)g�¹�n�(U�˛
4�$�':k��^k�Q2Ud��g�CX:�>������󭲌��I���S#���xOPoN�A(y�u=�8�>Q�@QD+���Z�-�;0���M	z;w��2�d�Ŗ�l|�&2}�D0'�C��΍�1�`�҉���y �8�� 7.:O<D���M	��K�P�O(���?M����ȯ�P���!R��y|���֞���#����p�K�)�Wr� ����Z௱מ�J҄Fh��\ӽ�)�]�H�(���h���u�
�
k��5�����T��H���UȽ6XM�96��y�{��p����BsV2����µ�2^�>
�C�	0�#�Z[~�_xd��ں���E��HZ�xn�R�3�u�����Q>�XH�ǀ���z��΃��V{�vYc�ߚao� �U�q��Y��J���3���w����n�AVֽ)V�ȭo�����_h�y�-EԦ.QX�����7;}�h��~A�G�˖Zg��E�T����%	��}�v�l�W}M�*#�;DE�4�GD��=a�硜-u=���w�����7���h 
����#���l0�O��#i��(��^�t�_�<�Aͦ��1������؞lG%T���
��K9�d|㟈��Db0�! ��U�a��ء���ƿ���q@���MҰ��Ϛ����
m�@��_���f�T�\|��wk�fX_>��0�G��c�>�	G-�ѠbWm��A�*Җ�V&�@azn�gA��W.�{rX�Y;ΐ�v�Y�g�=�]Ϫsg�<'�=;���}6���N��<L~<dxTRR��������t7$=MB�Y+u�=ұ�s�K����_���Xdwv�Fаz�k��U����U�5�rla>��P��$��A�
��Y��<��v<��;9�g�Qo��ވ�m�RB�U�S������}�-�6Ͳ�}��x�R�ۙ� �X	�"̪�&/�w�	�����X
"JK�����蟸W�}�KGO߃3Y=���34�-��;�.f\F��>Y^e�'�)/|��d�ym�!�:��N�A�	&d�	Ⱦ8I֬�퀹qJϫ�i�I��PMjuf�w}hM�5����#7�����_���=$��!��<��A��p�z��<0ۃڵ��%�5Ny����\9C���Et}�z��� W\�b+;؜�O�sNt�o$��%�Z��}��d�����o���(�QW7�m���*ٻ�+:������3Kb�#/�b�����!�L��y�\�ׅ/$�Y��<ͽ@��]���T�$	�ds��ί�$�o=�ׇYM�mp%��
�ѕ9ȯp��H�;X(C�4 @�Ģ�جD��u}��$��p��=P������b՟��34�a4��_��Z��.��r�f*��]����)g�?�����Г����j���ir�Xh!ٸ��J�n��Y����'n�j�����	I)��M��$n���5��X��Vu�@����2��m��]�����P�XR�m��ӈ�����r��)�R��J� �k]k���~z��"�y=DG퐐�:ȴ;.�`�-�:��O��:�_�2x�G�$?�F�E���|��]���k0{�DK4��F����f�k`��Gu>�(_y:o_bY�G�'8�Ts�SS �����s�]%H��^+d��v#�=���92��&�v��o]�"v\O����4d���N��M)G`�1
�A�����4�J����s�������w"�rg�����A4�b���=�S�M<���&��ZB�'���U�3+���!sB���}:���z��W��O���&���t�A%�`U���dTUK2��?�l>?���bP��+�IM3�3[cI�zt
��ۭ�8m�]�6�H�F��_ l�^ה#ӱ>�'�wO%x�Xx�q���*��k+���O�$7�uǘC�(�F/ ]Vz�����cU�T��3���q����(�O��d����Hy-}�2}���ϙO�cʘh��>���Ҽ7~s��D����[�A���場B�,�8{G��k�
�����~��ߩ�qUM��biM0�k"<�0E)�KH�B��U�&$�X�v7SnC�n�%rE��J��g.0��N�F��U)�AB {�[|jN�J1H���m�!��)�Ez:-�$�4�1/���F�t���aL	u.���_s8��R�E��$W�M	�&�����J+� �s��,tަJ-��tK׭�)��8x��)S-�ֱ��+!�T�ή!�΋�OҖ��f��r�Ǎ4ue�jSǬ����"І ���-fi�Z;����r�2���+��z��8�(�*�Wc	ʽ�H��)X� 5!�&%��t�L0�	����7�5|/q�� ��  >��d��ߊ04/!�ոI�y��+� S����&P?Y�+�`P=�i3b�tu-C�$�l�8�����
q��c�]�}`x�-�X�{�˯�CX{j���U��z��?�������v�! �L��h'犞OPM#�Y,8��*��D	$+Z<���HUHzM���\zr�_Z�� Wa�E�(~q�9�G�-�wS�M m��0��,�������%��~"q	0� x�{g�bÃ���� ��_��^�,���F�3{:Dq{�%
�2���<4�ڠA���	����uZ(��.��,v}�R�I'6��5�����DQm%��t��J�O� ��Db����1���wf���x>��7�1�Ĳ`�Bb*G5��G���RZ�{�,?�6�2�%�}�Tnw�o��:�/bub;;���j�/li{�jaH4wd�~�`���[y����P3!��8:?���������;��a2����G�?������ǒg��B� �kC4���]~�;⑅26l�-��O��i�/o3��'۟��P�W�����
ǈq�E~�x���5��Jq}#f-�sy�8�z���l��T���G��WӔrgW��F��6v��,�W��S[��ﾊ
�h5'��jL��Uފ\�C,��M��P2�5�P΃ߠ(��K� $_L[���P5��'z>�rn#�CM `t
�ܣ��K��#Ò�˸����jl��l �3E#�C,�ԇ3A��g7����Vx���ڠ��r7��劊kЀ�W>�9*"�Ҭb|t���a�q��yz�#$n�����2CX�]���9]ݚ87�5��+)�o�q�_�!{X��ǎ?ZXò�AR�з��u�]_g�8�lӅ�܄�%l9��@͑����KC{�"[vc���
�|�ܦ��s4�G��j� խu>#�T�tq�����;xК��8NM��� >L�,,K$`"�5����ϋ�T6;��g� d{ѭ�r��]�|�]Fm���6�����^y�=@�G�a�'Z� n��^p�I4�BW��=�ŔN����Q��j����4���2�}ќ��v��ֱ�yn���E�:����쐇U'���n��>�.D�,[���̾ژ�_�.�c�E�S� �I�B���r�t��B�z屦��S:���R�����VK֩��x6�����Ty��Q�����إ=3b_# fI��Y\F�~ٗԞ�v��w�o┵�[����E�z�X�!��?��!� �Mm��T7��������%:�����N�<RY��^?W:Y�l��hȺ^'�,�ƷM�C?�ٔF�VB�^�oJ��R}�z��b��ߟN��Cٕ0J4%0t	L��}�/�(/$Fx+��.�#� ]�c�U:b�\rw.^5���Ϯ�+
�]��`���b��'n�Iᮼ��/1�_��h�s�&��PlJ[+5��8��x�Y�wQ�;?��G��&������g(�`[^�O����]��a;����P���ڙG�O}�����sΜ�2/V�+d���~��%#8�p��N�/��~��\E�MY_��	巫ʔ�3�0B�#,�P�|O�0O�E����j� �[�`��ۛ;G=�o'Tྎ����6�1g�E�7�V�5� �O��2�M�h;\w��O�L���Pih�J�&zn�+q�B�^sOW`t�-t j�
�W%��߀+��\?��'d0�����y�7��!�/�c�!�yT�L�[yt)@8�3���2�%YoS��z�T^1J��B���0̶�"T��	9�_�;�5Sj�����z�oR���m&��5l�ae���Z��B�I�
�%�z[�w�����\�������R6��8h��Fkͱ�W,��lE�����L�p#ė:ݷ�wB��20/�����I�z������_|��D��ڨJ������[�* ��9��6$�?�/��->���g�I�FՌy������h����{+�WS�h��?k��cd�;��d��h�{�<�O��E,���;N��a�ʟr#P�V���]K����޾s��#n� ~�H:Q�5)�z�N	��L���D2��{��o���_�#$��6��@����<ּ̼sqK�1�Oa���i)�D���h��z��g6��Q�����
 A�|:]N� >u6Ҫ�G��G�s#���'2��1�p��j�6Lu+|�I��F�xF̖S<��%c̻)7d�+�  ����W֐�_�c�CD*�i��x�Վ�?����5��/�Ϙ1�iaSf����� �<	t�IUU�ü�`��ӏ2����O�4�PޚO����S�0m�[��z���I���*!�5f:��rc������3~E7@%�c�<�m�7,�Q����=kp�	+�m~����/P�&��1 
n�ǃ�Moa��=%�e��&�x�&�爲P�Zi�@��3PG��=�;��.���t7����W�,\��nd��|0��^��1<�&��
����B�B���≹�D��㺖>�;�����
��F�|��y��u=�����8��W�*�=���0�]B��|�=5�Y#�/m�)�C
�����I����tv1_���,*�! ����q�M!��	���E ����.:�Gz�E�0xĶ��u�jmG���an�r|KV��k�3��U^K*��<=�X���X�mɸ�4´�W��20H�0�m뜋�B�&�*N�_t��:�S��p<6���f����ȩ} ����U��{��(c{c���Ʋq蘜�P[����Na��Y�K)�o�b^��i|�\ޥ� ��F�~/��\�u�!���6�u�u��V.l�ձ$�s���6� ��_<@(6�M�����ӂ��LI�+�&Ӵ�K��;���&�Ē~$��-���&�G[���<+��_�=]�{i�[�"��D�bT9�4ņ�촲�va���(�BV�o�dm�f��!��X�և8����B4�p��j�(ћR�[ۭ��U+Q��솭_N95�o'� #+��6��D��d8�w@/�M�r3F��s21}�;���;�O��������O٦��� <����s^�p� ���"bﵘ�8��_�n���C��i$b�m�e�ü}� ͯMP���W�����o=Ξ�زW�?�����|D�_^������NJM���~���i*��4�q������⢙d0�NH^a���Ϋ�Y;P�tTG>�~��n���N�4c|H�m��E(��'	
<�}��1����\�~�K��$Q���1w�T����!��Vs6���Q�y�l��O-����bP�)j��o��`L� eN��Q7O^��_��s��Ӹ��<��%b�C�&g����v����o��!��o�8��v�`DpMT9
�7f�҈T�
e����Rj��0*����\�Z��X�.�/3�x��ɟ�F�2�% ��j��O��N�7�M�.��zd+t^�KM�����y'H�Pʄ��^����ܒje�f�-��i���ӨR���yLB.͸�UC25�?��ǭx�2Q�� VQ��:����jW~��/]4jTΝ6t��	�u|VB�uC6�9bm�����+��yN�D�pC�qE�aT߯��z�5�K�����)�yW�Z~Gw���D?��SC�m�e�M$Pt��t-����7x6׃�H\�I�<W�ݪ�v��k$4X$����R���D�ݸ^%*S�Kᓲ�£o��H��- 4����d�JB��S�W��L�2��3kCEΐ"!�����4��垀
�}�F�p#>����&դ��1�g�hw�Hj�����\df0�>���Uwc9V�,)	LPeH�ϡ$�7@@��R���V ��C�t�k$��QAm��+.EG�➤��-��(��A��d����1�_����'�S��}~.flR��Q�[���i�Rt����=|,����YX�3�$О��1E	�D�r��@�N�d���zW�5�ǛPy9��'`$+�3���=I��5�b�h����bl?Aw���)i��7<!�<��@�fX�G_����T��Vɏ�Q�0x~���l��R���q�
[�������*b�}
���~�z���T�Z�AH=��A��%I�:���#��r��k~C�j���O�NϺŀQc�� fb���Gf����'��cP_\��'RB��G��}��:�j�d`����_��Q���bj��T6�Z�Q�q�꣘`�=n�H�����r7V���~>Ł����i�ê=#��L��З�����
�C�d��E出>��K+\TIs��4�;d�j��`pV��(�g��[8s�s"����/EK:!x�ZO�{��Ug��{f<����e���s�+hb��+���v�~�BF�/�㟚c%dԘM�E�B�D �B�o�4�ø�c����{[���~<$��(5�a9z>�b�ލH�Y/衣�wK�N�!��A�^X'�䩺���s˶e��`�����= kJ�u�P�G����1S�ѓ)fF�w�ߢ�S�6Ɖ�W����$���c���t���mU�DyC�GP�5Kf���z?�lAM��mn��
�����OZ�����$��V� �O&>!�sXy<X+r�g7Ѽ���.Sh3����������@��|.��R�6��3[9�FFQ'��T������%�qYν��|x�+`�(0�Z�((�0d$��-���se�ʵ"� ��ZW�@5c%aM[�)b�J�y�h����|1M�K��c*>p�u����hdD����Օ즋.t�w�����PN�YU������Sr��G�^��f5�ҹ�.�<�降�[�%ĜC�3v};��p�&4ܞΪ[���%zC��بf	'��Ŀ��cg�l���v�5/�\lٞz��o�q�iHL�����Z��m(
���B��9>O����7N*�%�l�Q:&�E����f�pZqYp�g�i�uٝ��?�EF��$v܈��҉��^�.��j.C����vD&m��������(U��o\բ��P��[&�q�Uަp�r3Og笫�p��FP�z�&mte@a��[�������³iW0��G�υ�P�e.�[m ݾi� h}�d��37V=�Q$9%������_	<%���Y�+&ݩ�N�t;m�(a�~����7;��{-�����۔e{�Yÿ��.ff$��2��!�^�.6d�Os�p=���t�[�������Zo�'RG���%�(��4�����j��]�Q$&%��b�����/]�د�߸tSc�~�D1����#�B�`�n�����ƍ��Ia�t��`sn��VM����L"U5A}�nf��1�#<�o�/B�uȔ/x���q�]��7*�H�����_WN�-!/y��w�K���n%������3��z�Z �XOX�@7#X�(�oP�N�÷/��j�2UD�X�90��z��3&��)U��`��[K�����2�d&��*�Ѐ*`��3�/�r�Eƞ��[���k`�$z58�������q._�3���5�����gY����Cv1�C�_Șz%3�h��~��X��b\ T~&�#\�-�� ��?
��ɪ���hɏC��({	"����)!(d�$5߫�3��k�*��7�.�����Z�h/���tkM�����cz$�K�Z��i^4���:��q���M�*�����9+�t
�[�m%�S5�`TZ�Yx�G�|Wm������C�X����Quԓ���A�x0(��pcռ�x	H�������I�%ӯ�I�DIߝC:j&��c���bI��$\(Q�5̽����%�#/d�P��+G�&+&<=xC�S��[�Lv�s(���Λ��p|��'"�U&�A��sV�$���:L�����H�������9�b�a��@�[��r+��ހdq.'�K�{����5�K\�޻w�S�6�;���a@��P��!���0���HP���@fL�]�`�_u\6�ə{����5
����lD��=��	����iAa�o W�ŕ�+���FA��d������A��O�pؠR���Yh�F���Dg��f� 	��)�n`��A�4��y�L �%����-�F!��i�����O7��R1����$��CU�W@���i�?c���.�߸�6<��e���1Ţ��.I�L녉�A�z��)��%(V;��m1^1:S�[G��j��Չ͟��9��S����;�3����t�8�`q��^���>n�9��o~�[W+'���G������}
π4�Y��-i�n�OփQ�����Kϋ0[	Q����@-[�4��`�ia�ғ��&ʌ�fjP��̎�����fd[h�s&"M�Yq���]I;{�ܽ	�����l����_!�w��bt�#FS�p��B�c��ŵ�2~�Nާ崬�n$93��'���/?i�X�e�ܥ�f���o�����|
LG����FQ(��C^��m,���0:��kkv&�,V��½�9x�]Q7���i,E����7���mr�� �W�m�?��x:�={�n�[2����#�z7���& y��qM�S�f��	C,Cr��8��)���i�Y��/�>C�uwt�?7Z'�t���F���&���U�w����括��f�d��&^����ڞ⎿;�_+v�4I�VO���S�� ��ߟ�qi�h�:!ӥ𙣖�<��X�d]�{���P.���~z�^9G[K�aTh���'�Ja�����6	�~h�����\;nN#Fă�Q$�2	�J����5YX'R�O`3�,�բ�XJ ���(���v�kK�"R��]�y]Zq���Fh5�o.6":�ޛ��
o�`w[ɫ�h�����Bu���ן����(�^����K�߱��>R%)���W<�~6�j�P�3�������F8F���a ���(h�&~c� ,\t�;:�z�,�I�2��гPms��Y����~7vO�Rs�B�T�/n	�7��n�����Q�Xf��Tp��sP�%��d��#)����p�"�j �D���W�ٛӱ[����=����a�-�:
�x�S���=Ʌ�*�P���]A�j*���h����칙w���}8[�h���OT�Ee�u���V���ǁ^ �t�G�L�������*�0�xb
���c����ec�r�}xzBt'�U����>
��(l�*�7R΂���{�݇��b��ϫ+�s�[M]ʷy�<�������e���)B��kbt?3�d�1��Q@���okYPi�:l�]��y��<��k�e��2��<�s�ކ}ZYŻյR�+f�XA�����iK����[<Q�nKȵ�V��-u
��޽̔Κ�,`i�k���T���c�DR�����QrR$�D9����oje��4�n\��a������Y��|>q� ����y8�kyt0�M�20�X���^7�+M��N���P��e`tpH�m<������߮�e�S���$���9���r��>��+���o��f�U���i7��ߏd����U�*�U"�\�e���$�`liT0z>�W�?���V��a�C,�vRSy������\�e�;�Љ��p�GM����a�s)����t�Z�jM~X�����`��x�$P��.s�'N6�%iJ��^��w�p�������9xT��S�s[s�����j�E#��?���n���lPv ����I�N��v*���T�ĀN�r~]�(sx@S9n�l,�᣿N���p���u�}��8�.w�k�8[a�x��q�� ��bUQ4�8�z�����pڎ�D�/�.T?,X>�rMu�y��k�~T�V:;
"��/�[�g�I�R��E�y��ē�Z�!^�5��_��:o�f��$p߱χ��B(��m��RV�9�O$��J��x �1
�zA+� ��B�60���<����^ٽ��ߊ6]ڴW?���&f+y�hme3�/��b�Rq�pH�ܮm,�u�Tۄz�u�����T�\ƛ5(F!H�%^�0�,�\���`l~�܉��ϔ�,������/Jӗ"��|1�s]��1����o�^������tW1#�[�e$ʢ7�F�=�d�ӡ�2���Io�2� Wt��-;��l�^��/s��¾Kԓ.��LyOXϸ�!h �:���gt�<��V[��ȍ�={��6�C²S������>�R�/��=�T?C��\�mk� �V���<�ש��1�V���Jqmm	�)J�}> �iaH��{pM���"aQ�ؤ	��r�A]��>����V�n{EK��D'@�����5����B�O��mԤ��7;P����*ک���-�-i�H\ҡЦ��U�^ܤ׸ �F�.�u4���!%,bF ��"�:$²�!9m2!7�Ր�g~��ם��(��O�MM�e��Ύ5���S�6�Ñ�
<��b����Y�a�;F�����Ϣ�Q�l���/�.�=sƻgZ$1Mh"����.�������Нo4i�������H:6a���I�47/�Y�U��J�]L�ӎ��U)�7����OMd�Y�\]�A�>@9N5hS�ӟ��0s�L�x�w����u��9�6���-�~�R��l��T�p��a�{#i�7�����>F�+]�]�"}O0<�q<k	�%/پY,�������Ov0�G��T&����+J0H"�����r�ݤ�`� Q��8�b��i����P!;�����8�ͱ`���n���ҶO/��V��B}���Tv�4�۩4p���;N��S��q��}oƘD�'�yO��n�Jl���8��S�}��nt�ө���S"�+m�D��aZo_
�>S�{�bm��O�A�fguZټË ��f
�$� �-ʴ`
s,:�Ŷ���٫3�?1L�Q���2dS�qX�M��NN�sn
N����Brȗ��(�{����&�h|f�Yh�5;��y?tF"�gD�Ľ��3D��*O��u��3�F�N:�B������~��U
?ڕ�����6� L�_�r}��N�[4��`'��Y~�d?�!����_4�Lh��)Œq����-�S�g���Fv��{��T�؉�������ś�iϊ��@0�|�9��PM�R�������4��F|�-."�h��'ߒ�d�Z��D�"͇&w3������JSV;�F��L������������*C \�#P)H����xG�y���ߪ�u2F���kP���}�~ͭ��J�`����4�GĞ��y� "�.�g����J;��6�G��4���<>�lp�Wy�2k�WJc�U0����R��'��=#Q��uOJ3|W�G.G"㙍��2��0�",P�1�4h��jyn�0�2�	�p8 �����b�i��"Ldq����Z���hFQ=�Ę��cd�M��{��l}U1�v`��5AO�B}O5WD�֡Moۑ�� ���lj`do��D��H�wlF���d6*���k'�ww�I�W�Y� U����n�t];�[9b��"�G`l��˾���t��Ӳ,�ss]�&n�0�0`Vtb��yk.�=��$ jZ5�N,X����"�Y�&������H٬.>�BZ��pc����^�H��6��S��:�\>��G�O4*��.�S�ǥ�2�q�Y�eY��;���mk8��1��ƱA�	�Z!�M:F��w��W ��$�bK�	(9� ���G�FkE�>���z��R���'��Y���N��a��n\�������=�7W�����C^�"�6�|*L�/_��	��͛�i[P�U��K�l��M8���_�t���*�4'��,+/��ƴ�cO�@X����Q�����S�)�7��si��^�5�|�c��_���M��Y��[�g�(�H��'y�{<��o�X]Y�HM��\��H��(��D�A��B��f�.���㈌U�b[I�J�j��.��̖qE�u�I5X�{��<��e	6E��WM�=Ѧt6��h|]�EqJK�������y;,`ޏ|�;�d���K�k�w(��M�� �砎P���"�l	6����܀&���ku�m]� -�kK8������vU��HE��L��(fT<u
�����6�0li�)�����/��O� e�����5p�J1�zډ}l*:�}�(�箱!O��w��Y�����C(5��Fn��	
I[F%d�ʊ�<�An؈�N����!_�#�S!��Ҁ�Z�q�Ѝ�-�����o"�"��+��]/�d*(Ir��~F��%���gg 2��1�v	�i�"�z׷��_�+?��><��+`ќ�DDP:��Z  U��$y6�Ʌ�
���z��9�,E-��U�9rĬE"숋��K�ko��G�=�yʼ�g�� 6U����(L���O�:!@x�Of���q8��;Rs4�Mq�cR�.��-�8��������}��F�j'�f�O�SP�N���vU	���1:���m�D#�(���w�~4i���;gF������f��ON���9�h���
�n��s+x��K�y�AVo������.��w!,{MH QZ4��� ���-�^^�_��$I�����v���2,fz�K���i�LEq]������HZ4I:�}�7bZ���6WV�-��PQs���4��}��Zڄy��9Ma�P ��崊�52���}�A:B��t:Q��7�{��}��X����)'��Z���])P+��W�9e� ��F�ӡ;�n�}Y���t��?\���!��� De�yK�S�5%<�-7���S%b��]�����{\lu��d��@�`��׽K��Lש�uo�FaL�}�L��O"��f���ة�2B�a��ŠX�`g��x���lX�m0�7�2�,�ǻ�\�>�j�*oO�BG �m�N��SE�ŞM�\-������#��5_T�J��6��a{�0º��U��RVPTW���\Ӿ<����]K�yx@�K���TF\�ToV${A� d�ʟ���n����S:�d�������@z�=DE��o�j��y�]G���d�tP1�sđY������Njp�X?}�����3| �I�Y~�k��ӈB&�h�HG�pCٸ�3g�K���ϥe�*޽:6�`90�ԕ▸�}�D�a���N�%��r}�C1)L�%�Ѓ�- �j{���QcOv�P+��Q��ɛ�@������Iׂ*��\��'Qjiǜ�<��$�X�,��|lہ`�+;]�����p�=�K��JB^/���h�^d���U��!BORӾ��a#+V�,3�rRqu�b5G.�� ��ܻn�L?�lFv`ΎU����v ��zS����$rk}OA��]�z�\��<�BMRv9d�2ͱ�f�4�7�v^��"\��g8Ma�U�g=d�;�/�ذ�1�Cq��;S<��C;B"oKvRp����zd5M����'`F�md�>1������n�Ct�����'R(������7EY���?�2=�y��9Θ��	�y*��d�^���S��!r.�(	�B*�+@k�F�-�V�j�oIhTj�4��p�/%�lq$���傳�S���7և�J�~aE��R�4^m�A��֦��I��[��/�8�)�w��D�>���sR��b�|���e��H"�m����B!�d����s�<�m�Ϯ�`$����?X2��d��7 ����/s?�6���b&�c����í�N"�f��!������UN[��rj��O�����9T-�
��+-
=)č�L௣����{��<�)q��IS W-)��.ڻ(�J�LҀ��+k��(S���H�;�S+��3��-R��C}����733��8���$��dD5���}�hn���H��m�����."���5�.�ܶ��XǴ�'�_8�2fp��M�b>��(�d�.�����]#<6�ȡ$k�Vk�Y�C���fˈ`YT����ǂ�o/]�r�����+6��g�����zV�6]�t�x�w��\"���0W�<;,�X�ei[B9�5��"k�S�>�z��1���E�����(�+,y���#[HVԲÄ������OY�@Q�����l�q����o��嚨i�J��~�|�V�I�/�	���3#�h����!�Tg�zP�Uz��ٵ�t1x� �u�a��t3���cĠ�i�]�p��ݗP.�a��'Ȭ�JmO��֍��h�0�Z�to� ���rT1S`ѵ�ƕ����L��c�Oʢ=�9p�id�2�_S=��!�d�ʜ��Wl���mf/O�jYT(�k K�O��7H����-aV-ۥ ��$#�yjg�x�W~�a�Y&G`� Sm(�������}
�ˀP��V
�H�n3�]�rN;?�m���,T�bZ��]��}��b�܂Y�P8�U�E@��d��؀�/��怏B�4�el?ly���+�Y[\wM%ʄ��a�@� bɅ���C��>E�؀4�)d0�h��������n��*�<���l�?�8f�@���$�Z??�	� ��,�Κ��kd�
%���΄�M�u+RR�lv�V]B���Nb�����P=���qm���si��L:���H}��A�_�3s��r9?܈,����k�T��ն����jp1�n��*��h�{y��A� �\��:�,��)ܫP��0�n�k��`-h.���dXI�hPq�5��z`�#[�	v �� n'q�z����-����J�aY`�SN��Ѷ7���3�>g���������5�"OZ[0Y�ӫ�,��4y��rgd�P�������,�:��y/�a|�1������'�u����hU���EumT��S	�ܽ�H�2�`2�xksE@�s��o��D9���h+�x��8>��0n1t�X�E
�����I�5��Ge����_8o���Ɵ*�̹�O'e�2e�`x��6|���lЛoE��fO�%�$gJ�ֻ�_��d\��#��#���S�ml��� Ζ�>q_wU��9����Fq��<:�P�J��:����.�����X����S� T�s�-����GiM<D��ʚ�Pk�2��E�0a'Z�)c�/�p�
)�֗��`Pn���ƽ�\P�󻯿��z�?O���g;˪_Xď��7��l�D�i��b fr�d�G���|�aZ7�7^��$��P�l˰�9�`���r�/���/�M(�]����dݴ�d'�9*�&C��y��9*]�}(��+1�������N7$֔��i�!ԺIމ��cL0�jTG��g��|��i��l=~8��Nj����E�:� �3�ΘDM'OZA hs�#T�+Ў�5�E�Y��t4aǹS̱r͚��b(ԓwDv�fS��[��V�>��5'����Mr�����JjZ;�?�l�'�,u7�9t�1k:�F=��~H�~ľie��a��X����:|�0T�M��U��lo�M�����+g���]K2��O�DB�+����fk���q��ZIB�9����)� �?p��ƙ31i:ۯA�����s����/%�O!f��|N딁$�w["��vn�H�G��᢫2�]e�C�H/�̃~��~�?�v$C�����t�7sJ9k�_:Gv�/=�(j�UJ�^�v$ěF��] C}� @K�� ����KɌOs�z'�2����	�E̘[dS2A�n�0�ƶn���T����e��XE�
��q�mBn����,O� x�,�v?�<�FN���̲c�����:y�p�o�Zd�1���UZ6�ԿO�Z���k�#R =(���w����[���"�C�,�\z%���ć�@�>����r�@7$���a2x�A�B盖�� `�C��= ju��C,�}�f
��l���}���*y�a��\�|g���I*�
�����-A)�O)��-.�}�r�Y��~�B�|E}��R3���z�x��>��1�G`�]�1�4c��@-N���"�F�|ļ	6�$*��=��6�a�,sy:I��q;=��Z�60�te�)��Q=����Om=�����Es�F��VAa5=��L-g�_�]+R�l��6r����l(�a&+0W�����,K贪�H���he����(Z1O�Sz��W���6�#�n0-�%��;��x,f���������X�q%�d��MѾ�����-����a�k�߼�~����#o	�1�%x���d���e�lJ��ZU ~��2���AB��1R���Ajpaw����M>�Ϣ�]^��˺;�i9��	�����4�l������:�8�T�8��¼��S#���u�W9�R���A�(�f���4K��0 ����9�?	�$�- �����5��_+���$�#��F�u��Ԃ^��1��̼ȖH6�ݑ�m�NA{�����F�	ؙ��G�z��)+m S���׾-v.�,5�������I
	�H��^sK�,Q�����^ɢ!#��h�PgR1QE�7�����pl�O���M��&�F5^7��?9<����J����,�؄nZ�ҟ�C�2�*?��,�����u�jV�)-�������t��f,_O�X4��[8v�� ռ���:F���$��zMp�IאJQD?U?4?1�b����`��(��M}z�B��X&�P��	�p�ʹ�\%�m��O�`�r��sŋ,�V�Y��m��QweX��^�k�)���|�}���`�O�/[���@���+��h����wQ�2o���-��Z��eսP��0�y5B�;i����h�57��� �O2l�|�r��o��Wd��#��85���I�Z�	R2L5~��P�I��2.Aē���AȈ�����V��H��4x�˒<�hj�4D��kHdQV�������{�g�I�9k�m~�dEͩE�[Y�V3jGj��Ģ��b��q8I�~�YȀ9�?�N��X� �i��˄��*k#�G��+$��EQ3��*s���$��gϊ�9'�^й�5?����E�$p	 �Sy��ف4�Q����tr����Mh�}�wޠ�s�@5`zצ��ֈ����`~x�`���ݦe����N69��m�5	��[��ej��~�;�����P��b�}Ѡ�e�p�!es!�mjr2�V���ֺ	�/�]�Z�2Vy�g�p����W����9��x$e�/X�k�^p�9�KI>����~�:���ڹz�7U�q�0t�3�ص�\4��r�ǛR�%�4��|й� /�8~��2i�`3X��;9�D-�y�b�gq#����/�"Q��8>52�m��� �yGP�d�8I �~��ixD5䪑��ǔ�K&f��`H�K\/c��M�G�2�8����:�xc�B��kPCf��dg�q488���gu��_�?:ص�
1�C�*G��.;��/v�1���MosG�<��/6`��1
��9���Q�=�n=KNx���y:�$�����z���| Q����5t�����ATA�J�h�L�}$�^��U�k�l��iU�F7��A71�x �� ��U���%D�Ra�^4�y�,0���G#�L�BH�����z~֎6�z|^v(���z�tu��zR[W�Ŗ$����߬^� v9��d���'3D�Y��O�NHֵ�yD�j½�x�bNv�`�Csg�o+��c���BݥPȦ��������60�b�#�Q�r=�T;��ʮ-���痢&���������(H72�s�ܰ`����W�0�.���x�ܿ��g�mS�7��Bq��S*��&��)@z%�Qܩ�vt�]3�kE`��^�p�d�,�����5T����I�+$���?e)Ǡ�������jLt �΂�0�6�xu�}�>��j:%���k!�
}��{�掠�^��?�w�+���C�x��o�ڳ�v�3/K}�� B`��b��h>`ڣNr(����A7�*Y���w&��"y���S�^�s1���PX%Rb����Kl@�R]��}d݉ �iM��o�m�|r��ϩJ��j/5�K�����j�(����Ҝ����$�]L�)��������aٺ�$�a��/�s�bRu0w����_��@Uw��ĭYC ���
���Y�Q`yh�״��'-�_D%(F�cN�R~[�7M ��f�~T �Hu�0qP� FW,Op�"r30|CT�$�ih�:���!�^U vAr����v9͑:zre u��?�ﶯהc ܡv���������4;�X>���K.�,�fC�m3�9�e��L��ӴF�Yr/�9@�Ԫ����~'�X�5��l��ߧ/�}C��ۺ
��Ȅ"(xy�uV��~��5�І�sVr*�} #$L�>���Ǖ�S ᙀxX�E{h��c^"C�����m���)����jT*�}��H��׀��qe�{qw��`vK�<�����] �Uo6�޲Q��|�!`�n�.g��}�PQu�F�ȿ\9F>�ʺ95�U@���B:�� �
�����([�p�d�j�_�k�^[���@�YPXK�wv�A�8j���8�s�k�'�� �����d�6��D��K��h��uÝB���HI�(_�:��'/s����IF��:1-�-%!��N!_���K��u�Þ���Xr`�8=�$v���l�S�tӤl�"�S�
�b'��A��"�3�<��?ށ S���d��v��K<^�ۀ+T���I�u�fd�����	����i	f7��+�S���Q>�b/���ȳ�19��]<����3g�E���Z$��d��VY����D��-&��[2�m�,^���r�_��B�w���ޚv���F�+�+C��42�#]�G�d�%�<�G��28�5W��ox�T*��K�tBVO��+�_�}�7�%���3������%h���rT5sDL�d���Z[H��  ��]��\�Y>{�(�^Σl��a$"?mU��`�e��]<�Do�F c;�c��qG���r�2#��y���{��i�#�����՘!�ߎ�O��ڒ��<æ���5����z�0W4��{�5�7w�7�@<
�ĝ>MUl󤖈�	޾���=x�&�J!�N5�Q5!�|���3M�BE�e�ӵjpbw����P���a	�<,V��WΦ�s�������B�=Wh9��U���%���l؊`R��l��!"����2k�^; �RQ*AIS���xV���ul��h�hL��G�q΍�B���k��s��ǹ�gcA���|[**�2=��2���n����Mׇ���n��9I�UT��8/hG&xE�`k��y�.�����mJ$��w�ѭ��������,�e*@�.\��C%m�3:���p�W��f_́W}|�@�	0�}��������`Ძ�ͧlJ���:�8���Y����e�̨��1_���l������St�f�ވ�W������:�E��J"M��u߇����*
����&��ͺi���ȅQ��s��q��1����������-���32h�4�%>��z�^�vL��^��' ��\0k���Ԋ,���N� �L��4��ԆMav#Z����\�`%r(z��
��!l\#�<��+���¯���r��������j���k��ʬK��ќ��Wy�jk=��P��z<0l�9��	d
�J��_�E�1�v��1���Y�_��w���w(�.���1 ���9�;�7�j�u�6@��B���j���'nڶ�q�o�jr2�1Y���+d���;ӟL�8��W3C$���)�]}���5h�����@!�m�\۶%��8�rq8!�Vj!��j1�t�j��\�����%VE<x�޺��B���.�K�]��`r5xFL��Dv��=��&&.H�M�a��1��n�>^Yt��Z����,�pFU�Sp'H�K�������^?��23��i�=T�O�zVC1c��Դ�cA?c�����f�Y�i]�������i%�!�4�_}''U��0�c�HTZMkU�S8�ʓ���=L:K�BŊ�Q�������|�ŝ��ݗ�M��R�e��"Y*����u���5�,��Q,��{\�W��H��T����2��1A:𶶌��!�UF�о���e�?L��E�0�cjqU!w)F兕�q��'��29��u)��t2�l�i����c�b�֛b�R�B:�{�O��潭,�O������D�#oB�:x0�q{� x )��PE�҇�#�0��G�y��|>�Hǈ��{qT�<�*"��&��>��HH�pˊo!���~��2��;ϊ�nԲ��� �]�\�c!b l4+r�e4�@��~TAp[�����)�-��>��̗�u��(nqxg~WC�KXbb��	�
a������A�o�&�ݏT�бP^P>�����(`��:D�����6��=��ڗ,x�$���ړ���QK0e���t��I1?]A� �iSx�h�Yx9`=�pL�"�+"�	)<�H�6�����WDa�bq��Z'g`����ږ&�kA��3B�L�U~Țs����PN���sO��`���Q��S&e�5���wߌ���t��ܲ�T��<� �b6[s���lˣT`M�����e����o:zt��]�!�E�8���&�E}gE�n�g����859� �ނ�����WնS��
725.�e�l$Js��B�㡪v<��w��u�id�i��L�?�Z�QS1��G���1rq ����S��&�dD��\���&<כ.����8�5�l�P5�3�U������
𯺓��I�7U��X�@��bz��l��<�D��͛֩�y�� ��Z��C�KO�~�*jb��;�oPo�|���8���)��#�}m�k���3k�ǌ1�+��+Mְ������6�$�]�i�@ci�_im3O�ckzl�%�Y����Ԣ~�For
��>��ڈ��
���Z�+ �	ww���W���: &�/���Z��"h?���F����H�^J�����v0�Wk?�JwO���m����������(�n�;!��+����SxZ��
����1��{dq�U��5�-=��N�d��M	`�����]���b�r�=�L��@�4�,��ot'�h�C�sC$��\u\�tl?��ud�!:�.��$��>�&3��#%���!ufg�
�L(.)��n�s���.��zࢽ]�// �-���!X� ê�Ī��Y���3+��T��W��],ɩ�t���i?U��`�aZ؉�_��顭��3&����00xC@b��r0	@h���~�^xn��;&�ӝR7���5�|�=u���h`P4�P��}�(����޽M�����[|��X�qg��Y����/��b�[�Na�"[���$�M�8��"M�4��Q�������� �3�(P�
"�Op�N�%�մ؊��Aƞ�����H�W�o(p�E%�s8����"]��s�!�Rb�A���>oV��4e�`��Y�0$
��l*J��+�1��:�}���g�侣n�]�������KV�t�KF�!2�c+� K�F᳿�f��m%�����;Mw��ל����uqbF�7�v����s�t�ֲ
��č��ka���#k9�J�qӷ�J��Þ�kI9P�*~y%�6؟0��c�t�(O�S�`��*�\�0_��/͟�M�R�"`�JGl�_����ʴ��K_�!$7(��&ChG�K�N���̚�L��IR�]
k�5[@[:I���Z�Z������4��Zwy] �VFy��ٱ�HP�!6�W�������k	��i��AI�B����󉺀<�l��^5W�<����u�3`}2���>���s�ˑl#���bFiц�0p��$7'Cڤe�Pˎ�?�k<��'�p�?%n��@{�f�O-fp���u��j/�D�o��������
_{����M!�4�`	�2,�4�|b5���~���y�.�O���;���[
v�I(�N���{Y�K��I�� �+rH���\Z�K�x�h\=9���W���d�:����>�H��w�7�5���<KfX戉�Jlz�>��-�`a��Wš�{��~E�S=��K{���1>��c
:Jʰr���s�p��?N#vm?dF���"�Q���vUw�TE�9+~�.ݨ��>��/����s�:4r�e)���aO��/6�N�֯��L{5I�>�>6����
�mjR-�73�P�:Ugľ�af[m������3X�>�B��0��@�~��v�
~� ;<��yT�8�@l��۩K�Íz/����a��&��)\H�$�k��]f0f�{Kcn��ee�aQ�:~�~�:z܄���:o]ǐ�~O��w]�KQ��};zk�@�g�W��*y4��bW�R?	_�E>X�&/g����襧�U�MG�ޒ���[�_�6kh���b�{��E9��������l�α��ɿ��#' � z��1,x�Ed�ý����W4:
;��s���,AN�U���5�ք�y��v��� �Q�c�u@0$���j=h��b�;��h���Ar���c�C��> ��P�[�iɶ���4;�ǁmSx �����*3��;�F�*�,O�;M�dm��ޑ���U���IY >A21M��r��s?4q͟lĵ�9���x���b w���h|>�B�����E������.�-oN�U�l"u�gZ��@o=�:�ŹdS��~\��l����V)�;?� ��qL���
��AG����S�Ӯ˜Y$A1��aԹʳ��'�L�w��Ge�"�_�66	@���'��#3�<�`ex��7f�m��M2�*X ��ef��0df.ƛd*�_���g�9��Wu��C�xF��6��M���YȾꭍ��P�����?RcM�q���M��I��'`��B���[�z[�q�����������	�3:�>r��V�8�G
i8<�3��i),��tc�`����P<�@ԸQ���j�m��c�B�G~��� l5���v
PEW!:��Ĭ�}�J�1���D趜��a{'n(��.�&�lh��Y��ղ���d�y�}ǃ��@��Ro��=�S4t��o����j��'�_:6شO4~��x/)��-_��$�K�ה= V� �S��#R#��sE�|&]��X��((��M�R%�T�(��a;��!�7Rㆺ���KTX1E��[�MlF\7 �a6�����8;�3�c����bܢ�5:������ F1[ն)��z�n�eMy�[��k��	���
Sn���'��IfO��U$���5��p?��-��Ӓ�H�3��~S���.�~I8b�������;Nfc��1�@E��+T �����C��g^h:��	���]t�v��|eI��G�%��"�:q���X��Re��)�Vpo�@|t:>�H=�r6V����Y��Au�@2�&ڿ;�_'f�)�?x)�4 �W$pE-흨���h�[:��9�����}�[֫,�Me�W�$3*�*��>�z!��Y��Vjy�H֘�Pf�.��c�<�V�m��L(=8�A4��;A�%��XV�m���8Eb9c(;�n?cB9��_)8���Z@8~���;��CXB��2ZG���*�$���Wֲ�{J-m�8�iކ��IT��qиޢ�������EAlUr��I4},������8��>�|�%���ѯ�|ۥ~��o�����R��P[M�d�:�����f���8�*�z豴߾��pW\�N�O8���BL�RO�П��'7N���H`�#{�j���}���%���B=��y��Gg�,����t*�k?3;�&g��R^�O�N�6ջnw3]<�L𒥧I����KX<������D��1����K4�a�(�]��(��)Q���� u -}��N�O���,@��T�5�����X2��Xu[�d���B�1ms<>����
�^WR*5�67F�%$��E�+�x�3J�HTK����ťH��f��Ə�-�*�^�G�[�<m��	���F�c|��,V~k�҆41�H�0��I�y��,<e�T��٪�-FK}����i�95�3!3UW���;��ٯ!�ͦ\^�.��x���\P���t1�+��#��!��d���J�vF3�=����Z���mӿc�����G�q�S�C'�Z*�p��1�5\��2�����A7���eoL�����#�*E�|�9`.2�'9_	>�\h��S~:&�D$K3���X�?.��mO���6�9\��#�����?����ᛟ�5W��|�2�1�+:j�y����hu���r	�����;" qih����_h�CV��	���V tK���Y�,�%^�^BpKsp�C`YҒo�����6��qH֊�=�JI�S�MA˜�h��G,w�7 yn/���ry��L�a�k��-�Ku)ZL��q��[u� ���}�L�h�mڼ�Tm�`$	��)ǜ�K_�S����sR�iW�T���lक़g~RA�TGvs����<�Ȓ�Ո[Ѯr�<ͣ��SIh�����w��U,m���������Z6���7�"E?�yɫ���Ӊ��>�v���;�"��N�L���>�冋.S�H>x�[qF���k��p�o0S<�������gr����M���(��9���K}�3�I�ej�6*/�toT�-76^�h���֨tJ���_�o���)ƏʆI�:��kO�m2_��x5���FdMp���P_��Y�����|V�Y~)�^Y��U�N�d�U���Q±Z���\o8�k�xV��_T�9�$�C��x�m��o�]u
��vЪ��b����U	ॲӎ�	~��Q	��)��sJ�T�P��N�b�����&� �n֠�}UX�� 4�
_3�	�Na�(=�����[����T�6�v�l��M�~S�Ʒ��nr�]�˹�N����O,kc��f8]{L�ے9��5���;����u��Qjݹ.�
�)Y@�	��~�Pz�Pg���T} w�@�H���F���7�ki���D�^�Z�\�2�]�/k���j��XwN��`7���-�<y.���9�-!7)ȏ
��*m�gMJ\�Z_����i��Z`Lb�-��Ǻ��v�X<�˚8��r��X/�#�$���u���{�o��ZqB�8X�yC�.X���~%�3Z�+���X����X:�ߍX��t��P+ x���p�N}�ǉ���'e�m�<����wm�jC�g%�����}Q�S���E�ŏ�����:�J&A�,&}�|XF�~(ўNr�=�a��Y�,TE�$tV�Y��Oe��'�4������h�-�:ٿ�Ne�HX�rz��Ⳬ���J{YQ�[����cX��J�MC����1;�&�?�[ݍ���sl��{��(67�]��feڃ=X�gُ�F�S�SU���kk��0��/ �2�E�iC��'�����nj���r�#̗Z�����~�.A�S=��������&*�
�?�6+��.Tҩ V5��w��R�.H�댙}o���ȅ�E�H�(��Me_���}\���c�H��G�!�/�,�e���!즺\���0
P?/��ߓ���T���9�ъ�Ώ7Q���g�9����1�<4��o�d걲�d���&9���sI(P	�7o��	�ܪ����&������f��)3�+�e�B��J���7tz&?]j9�&���Xԭf�}h�P.\�:g��>���*�X�`G�V�p>� >l�0����A.Ѹ��F�|����lK��cl���A}YsM�o�C�� Ǯ��S��ޚ&�Y6D_J��	���~LE�k���*(ǅ��؁�<��"��F��ӌ(��Bps�q4�c�&�])m�-ūh�xY^l��Aq�>'(sFlpՙ�~m3T'j}sxImU8���+4�i6�og=�ל.��ׇ��}U���9C��F�����̳�6�ŀ|qXM8�K��­���o���ͬ�_oN޲Yʬ
Q��cz O
o$h�ѹ}(�9��K�ї�ZA�3q�<�Ձ�`@ Oo�a儯K����S놰4V
��ا�K�F�۴A5�%�l��ј����C��˻���L	�ؓA��$5>������}�{c�SOz�T= �Jy��ݸ�� !g�O�BϦN=~Һ��n��Vա��P��>`=c��Gz\e�]��ݍ�[w
t:����+bYp��FX4��q@Q@�5Lcv��;�)H������KJ�1��6(��@�"��X%�*�~@�T���!�p�t"s��]\�0$԰�%:�T� �۹��$j5�-Y �*�z��6���5*��;���> ~h �u��M$�m^f-���Ї�Ń��{�W�#Ot�Q�(q�`��P AMylc�®Y�1<��L��L�&'-S)��Cs��D
��ϴ�(K��<]FrE�����+���{�u���1�x��rLr��RՙS��I4s'\�1��������/0!����EϮ�-%�"I�<��#X��u{��-���������^;׌}ě�w��z�?�Bf�����|OM�#FiHJ�Rٰޔ��Ʊ&� �b)!��*�2/�Z��-�����H�QNN5	��H6���}��� | x��B��2�����K�v|������_��jT<�i-��_{�;�J^ܰ �5j;�0�i���;�

�O�d+0���HKM�!�iㅒ�;�=_�iR�D4[�!���_�d�/��6�f0�1�uk[WdE����ݞ1C2���2���2Z�Eh'�ID�}o����&��˯���b���T���ZL+�l���3���^�V.���nm[ ��bl�\(y#�$�G�5�{�SE]���Pg��Y����Hj��ΏK��l��t9��K�K=��p�+�6-n���1jz\�o��ťv�,�F� >��X3i�d�`�hf�ԫ�O���" ��I�$}e�UHGغ�?"rO=��jY����	ض� �������jmÖ*wNݢo�~�"��H�Zj�Дa��3s���C���N\]4�f�1�ח.�-��(A�M��z�K��m��'��ׁ|H�a��6'^2`���U�	>�pC�\�g����ʫvi8�E6��H%/&��h���q���k
R�����P�V�u�9j�I��;j8D���g�0��Т�˳d8��<H�����G���W�|ځ�ѡ��,H��v�j���#�m`Rv�)g#|�k��di�[R�lCC�g�׿�T:�?���\��+g66Art�ʙ��CbA�F6�.�#��� �ܳ���~��!�I>��Ew,��U�st�� `i~ݥ c}#�2�`k�*H�'� R4�?�9��ؾ�Zҋ`0$�K����,����ɝNoZMJ���˛�
���6^��'c%/d�.sk����z��{7i�w]����c���9Mv��FF���m�:t���Z��J������!�k�&�ͺhV�w��GWB��2���a��pm�I�s��V�g�)��B^[�w� ��<�c����P�\���"��ݯ�^$�ы����To c���h{���QMc1'*��9N�r�L����s9p��۬���Ф/4���zFE7�ܯ���ػ<�w�F�3:+����[g�i:��9ٶ#)�cKX@��m4_ґ 9?��Fݹ�(���5	��k�)������v��e�3����ЇB���QTꬆ��e[���?��B����\y���T���G�$�:D՜aA��/I��)�p�9`��Z<*�X�L�=I
��8�$f���G|�Zg�7*k����l�s�v�`���i�Z��Zb�Z�[�A�^2!� �yj�-��f!����@��bCܫSg���H����{�8u���R��H�I,���
Z��`��p�@��86Q;�1�P��\e���V9���k�e���Z��h�Jܟ�L�[%`�6�CM�:�?��1?F�,hE�(,�e�l���;�{�L�d��J�n� ѬJ�;��+Kzk�%g�u˟(�u2֐�;mK�R��r�+�ly�p4OOb�^������7xY��c?z�
"_��ż/R��~�:ڣ3nBx��'m�f-�_Z�Z�;�	����}81�� v��B���ߤ;>�[�j(� (�eG$}_=��-�lŐ�ϳ����M>�Qr��o�����Y3��ZBi�{ߑ2�Fnh㪰/��|�X�̞��F�YXն8�L&�w�����t���py����k��_��;�,��G�j#*:=�;�tތ"�@�D}��A�1@��Y�$����=C�$�ad\���j��\��o�+�g�P�O��gz�9%�^c.H��`�_���?ݱr1O�<M�`E�;��~Kb{a�[��!,�q"��լæk�i!�'���3]�%bG�"<�&�C:��A��_�����lr��Z��	"��o�����sV3�v��*S��T�E�{M[�>a��T��6�{�4ƹU_d�1T���V��U�)݁8�:&��Rtn� 7���ߓ�p�W7�J]��D�'��oh���n����ɛ��Bpu?ˇ]#�Sp�:��fד�ĹY|��׽K�L��M!�Ś��F�E�+�b��"hEW�օ��Rd��עh\�nH�����7j�^w&�Y��m�K�%�L�Im��_탱��BBe
��wyZ�4~֩?.�Eu�Oa�0�J�U�����D�+ya��	@ ���(y�t���L���lF�5��N��J��� Xm=���DTK�O1���]��;�9���=h����( �4��M���L�4sJn�y���0���c�B�4`nSa� �T�uȦ0����$��(�U[؜ >4g�ނ�A�Ԏ�0%�Qj�A�i��u8wi��n���Ȃ��+��"�����e ��h���,���P�� cX��s�o�<Q[Z	�į煚�#���IF�Ќ�g��"�`s+J[�/���w�l�U��"��̍�u5;g�.^��ή��ykue<� bu5]�ܱj���U��=�K���NЋ�Ă�ގ�BO��d�(9;��(�Ze u9ʕke��s���Q�\u���h@p��vA-s)�;4�w#�* !�P֘��Ij��1�"�*!����?������4fP#�2��.M���ǅ��l�����t��f�d#�w���U/a�a����>[_�mAjCxXP��,+�A�"r�VN1�3�d��nN�����t��Y�^�"E�҂+P�1d�X�W�`�
M��<�(�>Dnӏ* X�����{<�Zċ�K�ĉ1�0W;+(��J	��C�>}ckڥ�$ք=���+��J�8��u1!=�ǜY���PH�V?nژ�@
��#�� �A��� �I���~��W AhB`ƙTs����jEW�0��l�eu;�;�@��q��f�>6����!�#��]�t��b(BΜu�I���o�� Cۧ7D}�,N��٘��N�TJ1�ۇF7(�TTLg�:P.J�ޟ��|�&(/��.�ץ�C#ģ��8��4@�ר��#��Z4�1�X̸�nlu�Zn{H܀&tl��Ɲ��q�D��~�"�H��S��HQ�ί���Ǹ=�0R�#�TO蒴̎��z�Ńޔ4?p��@j{���S�7��Lon�r%�ûOT��N �	ee�X��Ma��7����x_��i������YOyh�K�z���Hɤj��팶���"��h��Vhn�G��r������J�˒i�Xq���I�|!o��S�|�,�*vS�E�|���i5�7xA|���19n�{(bkWs˘�3��P��wy�7��h5��z%#m����)@D�0������]�T����[����FEk�y�8����X�n���Ds��C�����	� �T����ia�Of�)�{�S؀�L��p��� $�K�C	e��h>����o�c��kŭ"�����*iM�ͻ\�1��U�r�ėl].4��]񍔋(���l������B�#D�t�9�o�!J�M<�j.���]j���)6��T�q�vw\JI�DdՄfaj5}o^ eW��k�Y׊��8kˬ��\F����gP�~���`K�Er�N0P�EYMFF�٫@���C�Ɣ��%ZsA�Jx{&Y��yS��N8.��
��מGJ䩍T��{���qI����S�ԧ\����\qW��dأ�v�$���Bo[#�YP{n����rb��v��G�[�߶Z�_1}��%��U��@Y��0�q�c�gb��X*�׸�g=W��zw �X�>{��%�cǕ~F���t��|d.Xhy������m��Z���vS�{��1��
'%��!8W����,������}�����e h�����^���Y�rV�m���VJ8��:�-�q]��.��c]�h7�g9lJ�z�̔zfO���l����̱ʃ�s�TZ(/�f=׋x�b����E��bӵA���?ʃD	��̙�w5���D��8�����J˂�&+A����+�:b��ɲ�}�c��ǃ& �ʨ6���]z��-;%�<T����U��x��`l_���8r�[<Ƨ-vT�������޳]zù*Rlv����3��@���&|ϱX�/x:�}�Y������<�4��xy%���@�O�v/R��w0��������+�
�9�F�F�M@��+|@Ʈ1���T8���X�_����[\�A���N㔵�V�JC�Q���5g�bWd�ly=�4&A���sp*5�"q,5��00iΤ���}��g��P�CbM,��5�տ�3�~�O��>6��U6�3��jw��)�IZ9��sM��8��;!+�W�X&��l�@�Om�a�<����:S��ݵ��V���m��i��&���CO����g�����,H��/�*-Y�����WC��b�JL�2��3މ�����������#�+�|�Q+��T<E��L�eQ�7���p˓%�M�{j6Kp���s�#o�H�~o�V�hl��#��M�WI[L�GX��g�Z�l�� ����q�9�'��cՓ�aO�.�dC�"�7�P�Ab�m���fo���ɴ����͘��aV#�y.�$w�mp���䒪���A���SV�D]�qG|Yξu1��ʊ�.IТf{ ��E��;~�G,��>fG�����9Ꞗ���01��ޫ��&)���+t��XN��n��q$��C8z�D����Cp��/NC���,�y�Q?�Iֺ��'���� ����jQGz�M�"s��vMmI-������(���������:��}$g�����k��8�e��p�lh���,o��nC�c ��u�#��� $;D��p��]#�zO�/�0T���'%�q�RbX���:�
y�Ɉ���}�M
��㥌��w�y�%v8��h�n{���[��܀s�#yv����g��̎FS:i���j�n���P���u��<l)q� i�@:�\�:�s�k'�wMM&-��Ni��=%�Ja� X�O+��S��@��v�łD.m���J��� j������DX]_@j����T��ƽ5D�1�&b�|�D��b��\���F�j�
�0�ܦ��ږ@{{���_����uP�XE�	w�4a�@��I:�I�����O:������ױ'�r�|���W��w��F$��.�#�0Q��:F�Y�����F��?���]��_q<SV&#\�08���6�v6/m{#��Vȭ�	{?�I�*᫝��j;Q����=��6�0y�c ޓ��v�x33�2�B���ќoK����׷�dDsoJ3��}�� ��k!��z|8����Of�T�TliuRC�������>��6aŭ4�e�>����������[�fjs� �'h��m�UO¦�ݪ�v�(�sڗ�٧�x�I�8��g`�����]�ے�F^sb7)�iϺue��j���R�
q�0��5P��G��"m�Dc�h��}Ps����z�[ɾh4
�9��S���:x^��T,�2�d����?�!5����,i�3ӓ(B��x!�IU�m�s5F�jS��V����]d�Z�Y�҅l�t���.n�Y:{������P��z��ZD#W`����aS65�G�݁�:��Q����(o�}žw�����7�G3�D�;z�cyv�k�u��ÑF`id�yq�L��_m i��S�d/ܛ.�*=Kb۽V:������<6�� ��Hqc���^�x�����K�}u�u.����+��D#�+��W��8��Cܕ��l��sZt^f��cF^Ф�.� �N�RB�,v���th|�������� ��t��j�J �L�I��lY|(�P{a��}G��N���@e�恁��r�S���ntۅ�H�{+���%:r����
'��Ee+��
=g�P.�z�����T�p�S�@	x[���z��X���}o����ya,6�@*~��i�^��F1b���d�M�ࢥ%�ĦJ�Y��0NAX���	�ә��瀡+Λ�Ḓw�+��G���M�Z���1Ӧ�k��R]�k��H�Խ_+��_2�s�q�|a�_�oU�_�分y���:���?����
m/s,�>}�װ�@`9���
�D��E����8εE�b����޲Ld��h�h�>�Dm�ؓ�c%^x�n���j8������[l��s���!O�;���U>�)�K�
qKf�����dxS"ʟ�f�GF�L��2�'���|���Y9���n}{
�gy?`�窫������Kw4:@x~���
�#��R��cBo&���"�������������5�����+B�7X�_�%	�{��94$��v���D���ɛ�?���&��6��Q/�b� ��U�!@�� B��e��0C"80����l>�������&����-����uO�����y�e=��˪�J?�*�,Up�fb�AZ�ԬVsΌV��Q+�g�6�Z�i(���/Y.�T��o:��!}鎾�h�u�����q+��� �j��	��1���YI��S�s���k}l!���v��;���j�_ظ�}��׵=�������cn�G�e9kW�װ���M�I,^��fS���Y�HM@	�\�����͊������{���R�W��P���:���p�������N!X����P,����^�PK���ljhb�dK��CAr�-�ǿ�P�(�qs��E�����ȯ<���N�m��-�?] Q��k�|��#�z|� 8�����F�n�t/���4�$i����+��R�&���(7��Y�ym�Ky0���!CQ��KS����ք]���˞�2��|�eb��ҫz��q�*"�CO��?����T��,Wh��Y�X�N�4r�
��s�JH�L�o�9p<.;kɨ�jYe~��5Q;w��؍��}�����?!�|��Ί��ؖ/��KX�ǽޯ~w���N�Z�ӏ:M�W����V�)�H�ʯ�_�� 5��x=���φ��"i�}��VRc���?S0.)�N�)���~I����Խ�O�P�se?��=����$�\Q�b���U1O9H8���azhQhM����.]�F�ǧ���--|[j>�0�����<�*��@w²w?�D�U����(�ofq�E��&�mS�4��) ��Xx(u4VL�*�q��#��M6��wb��(����|�#��Y�L5-m�3h^�,�0^�t�c�^��^ ݻ�����E5wǨw�(�(bRcn^V3��;�4��J�X����Yq��g�NR�5 &��Пl��{ӗZZ�,�1U^Ҵ*j.R:��6Ia�4 ��C���ì%�*}��J+��}��Zz�pѫS8�f����C����z�M��Z�"7F)R�T@��\5É?>�ܲ�B�D��K��ǓJǠ��7�$q�&u��/��xB��U��̒f�Es}t��r�ː]R�rl��P����*�S��|b�0��JwW�?p~E���fqp��x�G$����)+ CL"���&�5�����e�+�䋥?#��"�D�����ud #��N�2�PqǐO�� s����2w�`_�g���w�����2����.��ǯUH�� F��g�d��ӡ�� ��Ƥ�L��<F�A�R��=Xq:D_#��W�F.�I�d?�7�ww���S��Be�&��F|��)�W�ϫw��ڴ��L�hW��A+o��6]nWD�!"��p]�x׫]W H�F����	�L����C���U'G@$��('?]��&�z��`֌��'�=���pk���v�)�\�۬s&��q\�մ|�k�D��Ə�����0����ei{��_۰1˶�:�E�����#�J���Qhff}���C/`f� /��L�؏�n�>�6WN�;���Q��m��p�-�{}!s�6�����d��n�U�Ɍ���.v�͋����d���}-pa>?�2dQТ/��#xM2�������Ү�z>�U��*�/4?��o��/	���.�Yn�1������7wd�1�C6J���"�.IZ7F������JȦ��..�7��n@P�t���RG�E�:q~�=dT�m3���t������{����m!b����T��Pqk���+-���y?��y��nK����Yg�,��T����rb�y�e}ƊU�l4�W�����G�f´�E��t�V�0�8e2�2u���� �;�m o ��'cQ�ȥm�d�ɫ���=��1\��#W���\�U��t�Gǡ��2N}�w1f�Fk�i���r3z�I��m^���d���p�=���As�^@`l��}���A����9������P
1�����.���'AQ� !(�'eCЦ_F�^��ͅ�D���D��^Li�g�B�ڔD�Ѽl݌E���5;�1�tر}�=������/��<��� )����8m�=��ȍ�}��o�;!w�^�]s���3��Mq�o9E�u��aFۨ��	I�'��hn�[v�%�<T�^�h�\�6��������K&��c�M(����*��|����ih�Y03�$?2�	NG����8WuJd����������E�}A7��f�Z K����u�h��F7AfDq�F��*�;�C5�T(.��!7�x���ʋ㜔�=y�ղtg�A����=D��I�C�ӷIEu������~�sx��yld�}��%lst�F�JW)x�+#qsw�A��4��Hl��o]~����@/�$�z�S�}��kG����
����I��\�7�ic4�؆�ޭ5�6��qM��m�\D
@�8����ϑк4�Q����K5#T`��r�����
	���1�U5��|���^bl��g�-��KQ�Rfߖ���%�@����	^)�6}a0�uJnTvA2*}��r��dE��H�J�
�r�\D1l���Cg	*��o�7�'����k8o�"d���q��nكC(�DAc��&����z�-�θ6_�pN��ah���e���m�	B\FhY���W{�[q��Ѷy'=h�	������/\cR�|窻�4�o��f�yb�#!�k�qq�N�D���,�Z���Q��𒎓x��Ҿ�QqB2������˺]D-!�;��O��C�*� Ly����S�1��z��~��
[o�G�����X�o��y�C�5����Q�@FCh��c�zæ�1�č�追�K��bP�HjL�e�=�������k����g�}�k�u����;�	7�δ5Ȍ�a\S�0(i�3A�m��}��Eg�0�j��I�O��������E �>@"m;�����C|S��~�4WS��������kIF>�b��w�J�*�o����ܟIz���L��.	�LW"������E0+�i��k2˭u�E��^��F���z�]��<��Y�.E����?�,�GH^U�
�ha��P}��6wF���V� 񆭈���t��J��c��*�Pnܮŷ�a\�-�+�g`�x$2��<�nXF��+�ӏ����gbm$��X8�ț�?���҉Fg�Zc�ũ��ݒ��U;�����V��8���M7����]R��əL��t*�y � C�&���)�}����'�.�F�?L�`�>�j�?c��Γ�}?��*���m:V�7��Ǜ}�2/�BˌM3����((�&y�2)2C/B��sΛ.σ�.r:��Kٓ�C����ieH��W�X�ƶ*�T�D7����+ 
���%gп7f9�tZ�X�B>_l�b��QQL4�T���2c--xR��1��nѳ��8�-��-�Ճ욁���/q'��B�n��|9F��bG$.S�{�X'�ѕ	�o�p$�Iq���E2~������)���0�*�\���X�i㟱N7�J�El���v<�8r�=��'��&���2Kq����B�;����[%B��!QGz�w%8f���$��)�J�z>� �;��RJyβ�$KA��W�lRwi�*���*��A���G��6�`q�0����^`�	9���^�O>��t�su �'k*2��"��%�ϭc.���g�p�!Y��Ƕ1��w�?���X;^+��f
�eo�t���[<�X �-�I{̏Fr�h5/��]e��m+��<L�yQ��OP���{a���-��Y�'j��CQ�����l]�E[��3����/a�v�Yp��[q�����������.[^�QP�D���}+�u��w^�Ϙ�2�IC�H�`�Zħ�ݑ�B���P/�[��^ޗ��7��zı�'2�5kc�.�l�������tDO���E*�A3�k
&��#�;T��X������V��WUx��/4R#p�^�d���]�-�L��
�phݣ+��#���V#so���	��?�� �>
Q�藝>(�n�Κ��Ov-ϝbN+2���|WZ81���q]�pV���:JBu������Hә�#}Y��|U�T��/à�b�]���E*�hg0�?�2W�_����X����&�0xú-�����4MJ��9(��OvӮ/�c��*�í�/��
�J����4cK=q-����:�d���rO�T��G��Q��|���o_[�!o"3@$=h���ɯ�.Q!u��#�Qn0	���TR��<
���J�w��~�H�ai~����A�k�·6��a��%�`�xG���a<%�4@?�J�`��Dj���ز�����趾XY�+7�L��-Ap� �@�p���Bq�6d�2l��9`z���� Յ���v�lo�'�u0���	�+:�/2{I�$V���ԫjW1��խ�
���
���F�e��H���g��s;莝���(�	�&󯙋��c[$�\�6�>a�M�^���^o���
]���B�QP�e�X���a̸\>���C� ��4&�2Gw�4��Ƽ���D�s������0ڵvY~[�
��;��>�S�_�*�Z9�n�Z���[u�����0!Y:N�m�ޙC671Cy��U)��BhJ5�3�"���cx�2��"���5����$3�tv	l�/�w��T�R�.jb�A�k�������5gm0`��V����{w��8a<��mġ�NB��Zw)yo-�t���t�Ja�����p7ГS�H����8͘�o�_-���D�_h	 ]G���2&�#�Ut�,���0�_+|�"�������>w�KL5H��}��#p��0M��Ob�[Y��^���I�8����+'��o�{P�Q���,�4�Z���`k�2���	n��c��{_ʢ
Y3�A���-�xӾ��W�Z���K{{�Kv�.#���V�t-^��f��J�KY&�����TFԋB�@^��.�!���*R���I��V�����ᄋ;_0��UA�o���;l���ٞ���$��������D6I��	��Z5(�x�|ٹ|y�G4#^KwP�!�Լfӽ�
�:8���к���fW�@��]ʆh*�)M'�e�v��祱Fx�^ɲqq!_R=I���av X��[��~{�Ɍmr���x��$U�;����i� ں�����&o�Y��W���谕K_/h�bA�u�HBA��Y֒۞W�����,H�ǔc>c��?���$������wb{�-r&��]Qf������+sEU�eʘ��e6��Ԩwn�Y4�pI�T�8�<��� ��]0U���Ns�qO�?���x7�JZ��3�q??�:f�%�r���E�|����¬�+h[��NQ9�	���Aw2�6�������w?��0�Q}�.�iz���y�����+���i�PPR�9�`���3�˩w��P|m0���`���#�Ɂ��]g�^���-Bt���������D�����Zſ�iU�=��0���i��=�:�BP���Af�8�=Ĺ}��8E�CC�.A�K
���W��|r���\]�¯�6je��Mٹ·�C��u������R}�tQ���ȡ�s��#�cןmD�O��i����&����e�șt���٩���v�h�n�;�� �L3q@#�xĽ���:�����o�N%��&�H
�CQ^?���?�4�ū��(dڎ���n��L�d�O���ve1���Vh��q�O�C��H�HD��m���_؏����Y�I��0����+�Am�ɧ"���5V�ѽ��]��V⺢��g��ჩ� ��^�L�Ro#u|./�YX�j��D_B�_��3h�� $oi�R��m����t���y��$9p�6F���G�0(�B�d�˙��.�[��v��/�őg�9h��+�&z^rQrh����GB�/�]�AhлfH[׎�A
^���~ZG�^�Yu ������Z��Ⱥ�)�f�@��<a�p��Y��.�(�n;/w��2�,%��v��Re��/��a>"���p�b�%��L��#a�=��Cؽ5v�J�TЊ��ŦtN�[/A,��g�*��@0�6�����.�p�$���r`A6�d��R��'���������5H��s�[/+��P��|`p1�7At��3I�Q� ՞B��W�.�B˳���̈́�?S��N�$��-���v���-�����O�wK2�V�/+~�}�&8��<Ys��3ag���N9I3�1V��QG�C�0]���ոn��̗�K��b�6Z;06@.��$?s�i���:ݺHH��� i�|L�j��n*�HA^/��*�����_d��+�R���aH�A/`�ť����@�����0��yB���NBx�s�ķa��D�Ö�f^�آѣ|U��Q֚1);|y7�tb*rT�X����ݮ��H2A$Z��/��+*
�iL:���x_�Z�/�+H^t�_� �͈�����������Γq.Л˗�𖎣��
��Ow$�K|�XQ�툼���T(]j{ ��fW�Va�Z�ǉw	�rp�٠)}9I$Y�B[���y	P,!�P%׺�`��+�?�Ec[u{^��ѿ���X��U�{���������0�p-���UI#�..@K�%��K�L��Tv�� �E`��)�;mT[Gt��?�N*n����nĽ%����+F�9���oDktҰ�#Pc��	Im�-���wT��~]��tZYxk�����>���P|�.�r�i�ǄU�0 ��}��d
��q�9y�Nl���� �w		p��KB� ��y��{�)���$��I�݃�o�*�2�:�U�>�������`�K��ge�Qs�쏞gD�:�q�M�<��iË�u/.W�CU�SVP�eK.�s	�`m1����R�.m0 W.�$�X�w��?�(/���x}א#��8dW��O�9ND��{_r���/�o	׸{�>5[��_ڱ1�$�
���*�<���.""����0@t���M8�e�;Ǚ%&Z�M��[w�\#��u��۾Ng6�-7��_k#�k�])��x۳��ޠ-8l��1�U-0�un��@2X����dE%�jS����ă�+}�8�?ޗg�٤/7�M��S��L�
�x~�6�J�v0Hy!V6t5��9pW���DzWM��7u��A��x��'���� 	�q���I8?��r'�$?V��k�dxY��ZQ�Z�<|I�� @][\����jBZ�t�m5�#��*&Q���38�zh�*�0�������';�;�b7^����ٵ���]͸�>/��3���w�z��R�}'�$��S��������D�i*��[_�;p�4z�P$�kL��8�읝�ʇ|�f�� ?��Jy��Y��U�)25��"����H�zKjOv+��'4�b�}6 ��{���af��@Fs�Sš��7Y�ȫ;�@ld|��dB!E�_ˬZ�c:4[(�UW�)�l�5�~����B�8�lI!��N�Q�&�Ƚ�4ݒ>�I@�y�g�)�`�+�����c��� ����BA\���қ�Tʈ�7A�1%�8�\�����:��{d-Q��w�l*��V��~�B�;�!|<�j�l>4m6ڤO�|?�j�Źݚ�*<�h���2ޝIU�O�Ѽ�8�o����L)�F��x��3�fB�&�H9! ��J0��Ӓ�����fo��?3ԧ [I␼y�I�g���
I_y�����FP�n�L��cS����O����F�D
�l�ܼOSI5��%�$lu��0���	�)sdtR��L��J��K�u7W�>V�+�-/V�0���8z�Q<y�YR�>Q=yd��dܔ����n;�&�����\��J�O*U�����'����{�굏�a�ȴ�x�,��V�Zs�J��u��F4	�;N��v9"�ڠ���=J5�5ny:��ĮK��H�K$���0$�ݸy�2�����	�P<�'4!���5Xb%c� �3����>�`�qBdtc6tM���_gB*'�w�YU���,�&��QW-S��-29
Y��rL�.����V�h�q5f��o� e���x�ծx��*�L������ҕ�	������﷮���P@�/�rq�a*zj��e�D���R��;Q/�� .7���M�E��y"�g� �Cn��6C��>5��i�us�h2�����Rl�}݌gT��q�鴝%�D�-4c�ֺ.'U+��lJ���U�*�Tc�Z���U-��cZE�{�X ��C��AO07^�_�&�1�� y�{7�G8�����j�v�$X��d����B߷�WB���ݗ�v�WK��=��������*]���&���lw
H^%�C����Vk��3udD��<�LSd��� �V��S�� D�X�G`���^7�P��2gr
Z���xwA� �P�T3�������If@�t�� ֯*��/�޳�6��Kk4!-.�s�M�z�j,�����΃�g�j�"�-���p:���5u��+b塆�H�rc��i_�n�=��/1P ���n�)75����7���&|K� ү9���}�t��
m!�zFZ�$�4R��t�ÐT��[I��������Y~,6a�Ui��� SrK��v5�$�
�z�@\�	��͘�Z��r�IfWo�┮�U�d�����о�U�M�+�Vu${�� �2
)ņ!�,��輸Y�K�?aL̞3y�`�������3�������@���ޭz�>�.�\/
DI
��赴#4 �U��׽ ޜ7�wd�lʀ�!��o(/9��NΏ������m����1Hi�!�e��������(ı2xt5�r)8�_����亶��#a�H	sDm��3y�	U%�FM�+X�H���4ZX	s�v���4�����A�&+�XgY&f���Ӓc�.��I�|7�?�Jg����^?4�T�ڽC0����{�w�d}F��if��08b�B��\]W�c�M� ��A����,�˙�n���\#h�U[$��/V\�rVHNY��ǰ@A0Ȕ�;�/�f��b<+J��d~�kb�����#�J52Ug�F!��
���|)e������LP�7l�*U:�ƠP���AVJF��Iq�@���A��v�wb��.�y�˃
�6�vVUĨ��UC�7��ŵ�l)3%`?+�vS�4�@�������L�Kݮ�M��7�����Ł*7��&�\J���)�ׄ/v8��9�9+¹��)P�l�}*�o���(�6�e~'��#�u3 {�����zi�`F	��5U��-ꄯ�E���`~ΉQ�'^�3�{��AS.H���*�e�/��8	���8B�I�R ��:q|����甹��JK����rxn��d�}�;�k$�3{-��V���� n��Izaή!��^��Gժ�J�#!y��â���;��I>'��@��e��êR|���Wb9�e0��f�^�4��/�v�I�����=5wCo�l��[��T���f��of�6r�4��(�M�v_U���B�W�X��6nHi���Ն��EZ������C��%����b%��E����?ǵ�w���sk���>� )�ё	|Q���|�*a`	����· �X��[y���L��3z��rK��Cp�jVx���{QuV�l`�_��<��ؙ+�SO'��+�~{�: �/"��1��-�1[YbF8	vøigxM���t��G4+��E��o�����_G�5w���ܲ��w��)C�T.�g��{V��P:�Q�]u�tՒC{W�B�;�S�l+�)8�g�1��ip��3E�ʡ-�<���2���N�#|���tѫe������0�>L>�X�|5�D������
�r�����+�; ^m�P]UF/��Z
���.#�}&��q�ޱ��<�U;d`�
���Zb�7d��O$���&r����b��46�Q����\l4��χ���A����v܅���J�%;f"��	�wģ-�ƌ���6���S-a�EZ/�/zfꎼ�Ώ2i�����!�#+ߋ��v�v�Y�9O��O� ���J�uj�ל��-.@���iw*`�7_��'A��Į�����z��W 9��".T�}�-4Ő U#��Y��>v�X� )��g��%[k��O���w��hj�~�}�>�	�t��<h���[\�#%��� �����N��c�<!\�`sh��X{�q-���֟A����`�Li������]N:ܢD�S>���{5W��u���C��Q��s�%����{"�Q�z3�|˵j-B��h-�}8;	��ohpm�k�Y�l��`F��-]���\-��=�SB<��;�Òz|;M��;?��W��V_�>��]o���v�%�x��W-夣�y���b!<� ݓ1D$�����1ߝ��~Ot^�ڈ:|T� �X�7K���%���uR0;�]��
�K=&���!�.�@�9PS��4�)�;t
	d"��$ŀ"ؗt��R� �^�xV���7'�V���0E�+�N�H�ً�����T԰�f�s�Aŕu�}���O���,	:������P����q�;-H�6S�B&�%Q���kB�� �$�h�1̧3?u8]&�C{*z�v�ĳ�An��j��Mdw��M�6:\�ìꎾ�{��e�e��ǔG#�4�}),n[�.���)m��m�]k�����������{�H��6M�����;Ǟ��+ ��$�
����2��y���X��8�wQ�&��Vx��E��yT���
p�eF�ራ�����Ƈų���X,U0���q4Ae8�ú�&7	�1�(�3Ƥ�VR>N~P����� ����V�z>Y0r��V��O�3PD�5M#�P�� �R�EkBr���Q>�/�b�R��w��ҹ�ܡ�ȑ�>�?�u�$�v>"��]�Y���R�L�rȺ�	�塏�w������H
�Zw��]1��tMӵ -��)��_��-��{��`ۼ�,ji���&Z�%��Љ�a�Z��y:n6K7��)C=ɑR�$�@��Wp���3
a<~��n��ųѠ�9C����������
H,f��A�< fU�T�r��t�6w4��O�+�:k��҈p"xA�7�+��5�do:����:8��6wr
oi0�:$�d}9Z|���X ;B�иxf��v7�586]f��l�o6�wJϣ�%ָߒ+�H/�Mf��C���_j��:|	&�gh1�S��� ������|�����cc��q'�T��:9�[5���l��m��L�UE�U��X���̓*3�`c4�l��D2r�����]���� ��彫|�h?�n��]�/��s�+vi?^`f���F�g��0�kq+Ml;�ǣI}��L�8�����mE���4��'�b���/N+=���	�[���{H��Q�^���&]��$Wr�I0Z���egU��GrW�O��I�b��۳�a9�%�7�kob�'f�=�_;���(�2�=t �u�(�ia^�:�'#&="\��Q�"���j&Xp{��؍;M���6	5_��F�����eL*�g���a�FAji�+r/��}��}B��7j��O���i�J�A�>!�����	����S�/LV	�J��Mi��S�!��Q����U������.�;��XK����1]j�S,���8@�wT�/~�;P8�>��w��W
���}�f鶡|Q�� ���@/P0i0h�2��D��k�l�EA��D��w����È�>&�WR��!���R��dǹD�T�e|�cӔ���e���o'eL��,�k��W^)�{7`RV�O�TFB��U���x�j�E<K�f�hLV��;~j��B�$�rz�B�pߍLn ����⼭�gJ�A0��b���|Kd��*�f,�]�����E�d���旰i��	�*u�e ��.���G���U{�B{�f�*�N[}DwN��.21������to/��c&����.Po���Ri�b���"��Q"ɟ���tNGV?j�5c*h�Ah���BN�b'4�>�sLM�M�#*���������C�@���
�,��/���P:IB��M��ǧ#w��` ��6��:�B`*GT&�#�H��]���9+sԓFd�q��"�p�3��@-c�3�����$�oOFǻ �Q��9���]���ۤ��p"� Y_��������)�M�m�eN�6�fQ�C?�A/��f�����`!ޙ̞l�����PZlܬt��
ơ:#?��O��0�0Y�v/�I��y\�N$J��Wg��]\{<!��5�r����ʫ��0�:G��%�+�P<��=�%'�����W��@��%�z�I��a�;�sGu���q��)]�;��'y#>m����^I����>� $��3���w��ӊ�؉O�;�ÑC�����Î\A����ٓ=y'f��K��[=k[	�N�x�S�wuE*�yz9��-�hD����� qi*U0�c�v��G1	���4Áц��F�sK��D5�ߌ}6t�+��u���n���#F�w�=* ��9��:}v�����;H��Rs����c�l�a�<���Q�}vh�>��ѐ	�^�+݌�" �����X�,��qd��5{�| �j�jv6���wN�7.��z�،F��&���Ƨ�2*�v2�es,rI�H���E����r�.�؛��)�+��Gc'cJ�⫋�7�!�%jx:9�7O�0mZB<��1;g�bp/��	R�\�=768�7���D�� ��[aB���V����ǟ��q�[���"]��phi���4�m��cl��~�кt4}3I)8KL� ]H���I�E������i�L��?D�$��BU<I�v,b����'��эj�����~�������x��#IB�I�;kJ����$yW3�mh6�1�]��Ljq�9'���p�A.���quC �"�:��Y��g��.�~x@�j�-�����P��!*6�*[l�e�f�𺱞�1�� 8[5�_�&��f�A��лV�a�D3��m�L�'HN��nUG�O9[�:�bf4��"� �t��=���JYzǒ].m�� Yas'�wP��+K��7��a�;���w�T$˿���ߓ��-�g�}��V�OSF�r�?�h���6/�&�#�����.-q��S֭�����1+��T�߆�tWR���8�˶���x�q�t�Z��u'�v���2Ųۧ�2������Sv�e(1���,*s��e�tWx�Y��a̓���3�i����ǻv�	0~�Kn��)��
�uT����nY�nu��G�wk�!�$�np�Z�G-�ǥB�����'��7] �7�KjS���'��~*�z/�,T�H��3_jj�E>f�z����N�x��2�wX�&�B�/�j�>~�510������}�}H�,��� x:L���~�*C�\}J_���/hK}n��a�|���!�;$��꩔��ò�=[�����T�x�#*�z�}�0����H�qK6�s͇�K�s~���HW:�J��&�����],���g"�u�J:w����R߫�X<u�<�]fBp�)��&�$%N���;� �3ۘ�:�@���Ȉo+�t5���:g$4
Gīx��h��q%���|7<Q/c�|�]G<\���ā��"�H�����Z��V�츿��L�bUអ�{�4%[wZ�����%^E�`�<fp�Hu;���
z�_*!Q��G=�{�1A��5nR����wgӑr��L����~���.InB�]���U��K�.p�n��Z��6?-��ڽmy��K�A�ɜd�a��t2ɲ
=E��E��'��M�.I���9���bn��\?&N��5���,�@����Gb����̙���-n2�P�	y�s[���AUOT�/ �<����t�hux������n�}ZA��y!�����+*޲i=��Nw1r!�1�b�/�m���>B�4���C��M]�=���\�r�5SR�ZUAz����Cm�����8�_�vT!A�^� ����nAV.��M!�I��|���5\u�]+��2�>��_��O��ذk�J��l݈�z�pϵ�=Fu�z/���s�c�Z�i#uY�~I�_���?!O)U	t�ð��������O:��Ŋ�u��Wa�8�h/�<-h '�x��N�]��.�4�x4�L���״������\D8�|yxĚAfs˙' -� �Ek��{�ݕ�o7Q?��%o7?A���w��g�
R=�"0����ߌE�x
)�&ߤR֖��R"�3=m�o:֓����d?��5])��"w��͓t��^1o���q�u�q�����vP\��].3�iFrv
K�~?v �+�V젠����cV��M���	��\���:i��_L;���j&�*�@��rA���Wك ��i���ݡdX�>8�ų=HC�!�;]+�Nl����Qȫ�{�O����u:dS�t"}�J}R���i��U�{5M�쀦F���d5�&��η����\K�`�yY�it ��~?�>�%0r���v�.]��%v/���������[$��r�4�j���LF��0h���q⭏����/d�A���#{������sU\�1��v�O�a:��xwJ�=�� �w�d8p���	!�*�~�%��:��vV���V��C����IR�K�&�6iJJX �d�p� 6�fa�"6�(̽6Y��*D�'i�1��d�Q(,�����R����%*��Uil�fk��UP����E�X����е�&e��<d���D�ֹ��q��}�rC/��g�;����U�b)��W7%"njD�pvy��F�(���F��h������}i�Vk=����Y���d%�&+d(y}F�+��a��L�.ß��l��g CG(*P������-��~V�be��;�K�	��2Tp֬����QA���Q~�V�bj��WT���`-�!7A��&�G|��$�&6�<��>-G����. m�o��i:���5H|<��H|(��;�T̪�����7��D��qz1��z�E	���~p���Is����54���OJ~��B/e���������HȁBÜ��_v�,
tԁ��m�3}���Cݘ�Y�iA��U����}�k����e��ؑ�@�=9�>.��S�������'<��fM��7�'��C�� g���xO@�����腒V�A鰪�J��0���S��� u�b��躔��@��j�
�L���T] ���KdHă�3?���1�di�2߽o��Sy��X�2���������o����?rD���*�� ��˷�v~'<!��5�e�
��P[�5����\�z�cw����}�ę�?O���Y�++6ӆXiۻ�R�D�I+$ӹ��_�f�=pF�Ư����ɒLC�m�RbsB�rD�u�pA䨽�)x�k��q���$'������`�jo�0\��̚��&��t�D�y����?]$ƞ�ʷɋ�ҕ�,�6��pһ��tI�?X�roP .4`������Z���mF�*�~Fj����m��U���J���ȓ�N|�	��f�n�74�Gq����|n��N?p���q���j�s+a�AMYVY��
��%�-��yy"9�S���j2S��?�j��[�?�T��+X�9��3M����!9V�wH.x����(q~mm�¶Y0�[k��c�+�f�9��Ǵ�8��Nq�%�}8��W*ZU	�0K�:���M��C����)�v6��x�߉��0����0���Xs��(5��F��Y%Gql��wH�8]G\.C�:�|+�M�=��'%�����7%O����W��@��5���d¿�+_:�'�v"bA*Q`��,�"'i ;��H�gU�^�$i�[<36u�4d��،�i�����;�h���ތXB�ek�?-��J�u+��h�����S��ݶ�a#M@�I�>��N�#%D��A��	��cc��z�UF ���>.���o���p7�-f�'��J* $s3��i���jbO�3/�9������C؝f�\N��j��Wk�6anͭ��}�QX%!{S�H�s�mK�%����g+�o����Yp��n4�4�kF�-W(�q[�����z����t����!^���8wX��.��tS�7��}���M���|1_	���#u�*�Qp�x���7�C������ء��#R'�W�'�9q,阮���xMN�� ���yS�K��m�.z�D�gl��æ��TQV/��})�W��Г�rWT�y��,��$��t�pkq^����%7 M��'�	��]͋��O�/"�,��u�){QX֞Ax��+��Ϻ�}�_�	����^�z𥡐���id}6,�Z#���_�V?����Ɉ>zJD�s�W��M��^G{� ��IS�=� t1�,t�j��l[΢-�,qj���}�:E�������)��]Z���m���~���@D}k�t�1B�g�m1���u
Y��C���9�b��q9�j�r�����'��~(�m�z��F�
� f΂T��L��jA���8�rݾ­�zO������ۮW˵����n*}��ƃ!q� \byJ�Y�N䫯�8~n#f� ��S�O�:�Qo���q;�������s�ޔ�8	�4�d��`2j�\d?Ց�E�U�>����|�{Gfgݲw���TC���
��;��F�tC�Ī���b"���%�e����r^.#59Ф����p`q��阗j�E����(}g��^��5:���Nʑ� ��?�*��AL �N��K�F9\���[�ڻE��%\l���_N~�.賏�5�F�>>ZW�)Bor�{ʻip4����:���W�M�x�ڲ-�"R7�n�20�.#�L�]ɭȀ��" ��Y���X��h��q����7~s�����`9c[��X��Em/KcPGt�ý��>�=�2O^o��]OT* a@�����S�A�t�V�1�����g��3��hWs_qmK�Wc�r�T���[L�HZ���;�<l�L�]�ϼ�,r���1���+q�%�x����t�#��"\TmƏ7
|w򄷲��l'K[W�纚���������?qV�(R >���2��l3$�X�PR�ّr��|W�vi�m,���mQ��ԭ'.I]�E�?G�&O�W�ES7�(w��}KN2���>��"�1%����t��A� �d�����H�avgmf��p���|�r?�(6^�M��Am2"�Fp������4|�qf��q�Y)u3�V�_l]������%��*�f�B,'�RY��7� ��rF�P��pH���77�����ؙQ춴��+g��Dnݨ�Fd����>����:V/��3��}�N��k�<R@��%�oq�g�)�f=��L��d�Q��ڮ]�V�prr*�|$o~�Y+v�� B,ZA������&i��^�������,^�Yq��-Ҭ~w��7�����JYJ�?T��b�t�Ւv��>�R���#( NS��Q=��5�N��B���q���44�ߺŪ*3�ݺ��{v?���D�o e�y�w,1�n�oi ٣#	}�X�O�lk�+iB6�$���M���ITCV�f�#��0���[) ~|��T̪�2�ζOvVڃ�(�f��^*�Nu�Q_����J��r�BA�*�=o���	��f��O�_%�^���#���=#�.����ho�eC����0 4�T#�%�''#{u ���Rߎ�
?�G�����Ѕ3X�A���dI�	B����{2^��V�$�<�L4�Y4�l�{���E}��egk�}'�Ғ52d� ʭ2+6��r��"���?&� &-VG����ւ@�%8~2���Dɿ�r8ﲗ���5�mf�u6A��W���5>
@;� ;u�_���ж�g� |����H5,d��U���/�� ޾�(Z�k,�\�����!
4l��� �괮۟��sI+et������tvC��|В���.;p�b����[e0_Fϸ��%����S�iO1���H���#VS�*�"v;k>�F��B:S��@CXJ��WbȔ�J��3i�	�K�Y��q�)U�\K���_�������>���f�1j�:��#ex�T6
�	�������O�έ1�p��^;AK��`�a+9;S%�䇘ľ�v����u��
�����\�O
�7��-_�qJ==/,�"�~�H�����cz5�6�鴊�۱l���]���8�j�w���x4�^|��B�A�K�����s�:�j��7Rׯ�K��9σGTϙ��t�O���CM|�C~�~_��w��dmNN1�*�ZSN���R�g��.�.b�JNw:TO����آt"�b�u�DH9�� ���Z�[sT�W�t~�+���n�,�I��h
��*���V�o:p�K����W������^)/�����=�|y�}>
�F��Hu�v^�<B��o��7�F�+�\ݕ�M  z�)����h�߭�s�#.����!4��%����Y�1b�}�v̝��=���n���ӝ�C��l�y�+�w28���Q.E5:)U��_t�ѱ��P �up�`�[��P2F���i۳�C�������3��[�������O�7)��zt�P�'�	[%��E�&X�����u���_�������+��`�WN�?�a����yxt�{�p�� lڦ���C�7�ea1���a����xK�sIZ ��h! �N�0�^�i��� ��#���� ��dS���d�¯�`�ASo�\Y0?�-��&}�7YV�px�T�S��䝎�P�	��9�t�#�w����Z�Y��ȯ��Ɓ��`I���jں�7�p%���nx�V
o�����w7f��p�d'p ��4W{-�вYNru�/m�]���a�hݭW�qѝ�My��<�����(����ITf_uy�t��]k��W�%bc��.�!��p^��7�Lo�������&?-D���{�/g���B�o^oAr�S/��X��B��^�8~ph�P���J����d�Q�R}���L�J��[��(�'vB]�1(;0t�UM[iI(TF#zlᡍ�:w.ea{6�-�����K��* �o(�J�`�ihU��x�y�獴�t�C6⢺�O|+v{J����h|E���־�����J�����{�]���l]��B�-��밅RbՐ����?۷1�N��1׊J���銢E����<���ʛG�;yB��C�`�boN�	�`g���� _O��� ��0�z@���'�@`{�e�M�!��I�����˂�>�C[���y�N�-���A�iU@�m`�J L�O�,>� ���s�A�D&�ݶàe;lgb$a����������a0�A�a:n����Bܗ�q��wx���a�a��M�`w������L��0 U�{�KXN*E
�jL带5p� t�3}�q��F����ݰ���K�4��zu�P�%��s�!�#��i���0�*��}~�+3T��Q�-z��K���������3����2��w	�A��E�{_{R�H�����GuɎ�!��F�?ߧ ��}��U^	~x��I�_Q���QFÖ���T��n0X��FǕ{B֓��u���*f���Fde�7{Kd ��kh 'k˰/r�v�My��i�����@�*l��C����c��=$D�LC��]���K��̪S�]��p��4�I)h6�-�q�Y��&{�b����N�-�%���;U�P�jrO�U�p3��Մ������/Z*0Eʧ�Lx� �〄By�� B�tF�{�Ùѵ�(.q���S�5A���p��X:���PCUl,C��.�h�X LT��Ew��6�ai#�>�Yp���#��&~�/�+I ���\�d�	<Z��7��}?e�ܬTe��M�Rl�z`��^N�J��.ުz�����O��vH�kb��w �=��zq�.	�TYW"?�8\�I^HU����Gv/&k5��Ad��lk�(SgHn��G���l�\�I�>���@�,�����E�"$_��d��Pc&�y����X�fGy/����,_�z�5�X@+g��S�vC��ʮW��tc�fNb�^�I��T�ol���+�����f5�puV!t�"#C������?�W�o�pY��w �O��I*P�ǃA�H�����4�����:b�ɹTl�N<;G
���d=�Bp��#�{�W-�jz���N��_9���A��{Aά��ʐ
�8�Hy�ן�^�J`��5��\a˓\[���$���Q�V�kIs��2k�P� >��&��@�l�.F�����S��u�S��.p�i�mf�\D FwD���l9�~`�}|
���%�|�ۃ�`�f `��{���A�)�Fv�HM8|ჲ҈mw�8�t ��?lPo��#�n�׀��`R�y�:�=�ã��.�_$�5�jNf%�Ӓ���]u�MH��
|#�d���.pJĳ���<9����b��S:�Xu�5;���Z���N�z�g��SZa�#K2w���Im�&A����C;��j���yUB6�4<��L�߉�l�<_�:1mB��+*�#�.���`b�O&$��v���R�~���'�Q�*Nˍb���-�ok���hf����9 �� ��<Tƥ���W��t�����Ň�y�>T=֘�� �E���] l�����G��c�|�o���{�<)�հI7�(0�3���%����y�g�h�h��`(E45Q��ic�ڪU6/�.F	]�43vA�B^����g��e#��!;�d/'^j	��ɾ�������%�<�wЬ�IfF��C����_+���$�$�@��s�,��<ģ���a���&��l� 6� ���h��=~1Q�8�vcHk#���
%�-�w_�ڑR�Me�p�ä2��jw�0�g(�)��-�G�O��n���#�H/q嬯t�~�z����U
!��He��40k�Z��'�9g���cq�����/��ZZ����Q��KT[;���s��!Ct����5"�^T���G�����W��u�/:��%����a��A����
��[�c�;g�2�Tc�9�5E:
"�g���T�-�z�G5 �����*P0YK��1u	G%BT�hEk��"��-ʶ��]U�;����vݲO�wZJ[�iA�(������4j���n�u�Z�Q�"�����������m�n�>^)���s1�u��6���/yj/3�a�����_��~�5�� ��jB��״�B�$��{p�<1���F�O��������ۻ��a[K?y�m"2Z�%�;�жZ�Z
K5?<S���\Ai��u<���#�2��1��9xp��x����gN�߾Y8�mtBm�0Qh{rN���=���<��&A|�)
��%�k�1���]��������-�N��J-��2�P��N͋
��HI�HF�H����X�|���}Hi�V�#�rV�54�2o�n�['��~s�)ꄸɢ��>��7���k7*�1e'��@�Atl�F.8!�e��'��Z�]g�}���y���i�8]��Ne�����óΪ�.���v���*�U����8� G�*�~U_k�XO�4�9�Cȟ��pt�okTI��ۯ/�P��X�������V�vw	KGҟ�u�S�Ȏ?L(s�>T�[�B��gQ��g]2B�Նdf:��{	��٨���N�ݹ�]��Q=�o�c&Ït8���fM!Wr�]Zcs��6�~�o�Z}���0m��9�B5�ko���%S|x��2r0�HH!��;�)�f����yh���gI��c�&׃�������Q�νnS߁��y�o�"v�M��{��1"'���	��p��x��x�i��i��\�!�h�Z�T[������5i@u��w�㢁���f�Y1�+C:ֿ��]gU�ߊ̍<؇��t��F��A�rh�z�Şd�nKt�B�Ȗ�ipK��!��C���2�v��[�YG�/:��{.zR����9��[;ڈr�N� 2L�͇���[�4:5.�pG:S��_������жK�N����cw�w���w� t�`�@O�VC�+R ;�4�ޞ�H�U���%��	R[Ԩ1n۬��]��w�f�#s9�W�ݴ2� �,�RZK;�� �
v��0�6ЖV;:vG�|��y���o���D�3��
xъ*��5�e��j_�㸼��[�p@y�ܦ����7R�Yݧl9�'�WI+]��?�B�2���O��:���}R$0,DD�g'>�<]3�� X��rܕ��&��M�d�-B�ފ.3{u�MJ�����m�/g��*�u��w�1�$����j{�����c��@����)t*���f��2Z�qmޗ�ڠ����Θ)��T���2�-t�h�z�/Z+�1E)�}Cz�-���/��o"_���-1�p� )�*��^g`�̬z�c�(��G���l�e����R��dX��-�vI�Ck���(ы���R+Gº��|
c��7!�K��bt����*���#�'�N�-�W��h�~�zjc����1&��>����{�8������FW�Y3G�_�q��(|*#�����|�Iص�����,�I�F������p�y��+g?C'�TBn\m�e�P�c�Kڅ�XN�9IHw>�65� M���t��]H��-�'������Y�x86�]*X^J0\	��҄_�2~�g;@�*@,h*�jRJ�B'(�����-K��y�:�,3aH�:'�ٱ"�$�h(��{)Q���6k�f~�<�-�
�&`X�I#d�&2ϕ=�(+wls��ɠ�k#r���|��e���^�j|D>|	"34�R\}�V?�b���	s��ܮ�& .{M���)S��c>DemL�
�\Nѵ�d
����N�pv��o�;o< �Z�L\�����e�B����M|����J��#@_(��l�ˤ����`ǳ���Ò͘$!#�T�鰣�n��,a��=�	���#h��^� :n��jٶ��Ef���Y�������y�%fqך��U��9?��" }'k��h����|�-kBa"��x���|3.]4�~$lI����볿�c�qm˒,9'�iέ崀�xGࠁa=����r�,��Am��7©ٶ�����r��,���!U�����7>���ب�t��_(P���f(�{�Q����M;��+��O9D36����UH/�7����G���fR���*�M��59|��? |�����U��Z����֥�(�0="�;!B�4t��yO�ˉ�ޖ�����V�����K��s�������b�]6�ffR�hHF�u�Hꅰ?���zA�ٚb���SA� ����Fw�$���?��[5��y
PoEq�T GI��K��t4*a�]����8x�[��]��*���Ֆc-��YQxecE02SAArQ�Q~��~Ζe��{*�G�b6%�t�
*���R���x�2I�9(��nzK��b�C�/6?%��l��Xt�U�i��AP��?��;y���,�nn�P��:.�&3�w���9Dɢs�k��Q�Wd�~�	��<~������IX}XL2�/�S��!��"�4!l�=J�"o�r�Ϯ|8���q�;C�$gp��#�4ƿ9�����[)A+��hg�>�x	��^NJs�����܃m�ŕ]CZ���}���nu�|��0����?Z�������]�k��Wi뱔d� ���4B1�L)�O�z�t1�1�����Rl)H{;���l��ܹҰ+�dRGC�Zx���#|�}�¢P�O^�:�n����B,��tr���k�7�ޓ��26vUz�'Aa�dz{Ɋ 
�����{v�ֳ�S>�ȅ��C$�Os�t��wYw�!�����1q<��Wd*s�YD!j�ѭÖЬ^>-�ี�F6�ӥs$��@�,F��a��Y;N��ޠ�̙�ոp}Ӧj�aS�7�"��4�~`�KNT��8��v.�#|G��+�k�Q�
(gO&��b� 6۳<K��?G��`r B����s	�;��?�ǡ\�0H�Q*ue?���������s�<�������J�5���㩃�D��~XNo�r{���Q>V���r�\�`�mk������P�$�B�(��&�ř��5����ڐ��ݯ�bio�C&"^�V��7�����S��y���+,�����r��R�[v�-��4�N��J��fGN{5#y�%j�d�8!6ͨ�e��̞�8�)��, �P���1 �S|�
y����O�bI����U*����E`���2��ωS����sB���J�jt'�D�魼��@| ��qQ&e�E-���+��*\����6��m�0������� �����M�M�l�gPa�uj��=�pU��1�V���7�� �$f;fq�<���,�4Z�А�J�?�lQ��J�Y�S�8���|Z]tSV����!>�]��h���Q;[�"Ȼyͼ�nc�=��8��.t^���a]	l~�"�-M��Ŀr)*o&'�n 9rJ����<!ЊWd�k�.�6�mxFG��p>��A�����)�R��/�+@ě|�jb�r~�EZBef:w��zi ������>�K�z%K��bc�:�n���/�J��xe>pDj��S$A�=]�'��EĊ,.Dl��#���u;z�~��
��P��N74��[I��сM�����ϴ,il�(�Ֆa[��,�$S��<��PpNs�M�Vh��ŏ��$Y��&s��K�S4��p�1dO��S�����Q;�����C��v�*�I޹����Y4�R���t�_޲��<��q���c�B��(��S�s� �k*X7C;3|V��V��x��
)}�U��WQ�p�EkF��к�#��t�H{�}�����O�0�����h��3Wq�2ޜ�SCv԰����l��Ǿ���,��p��ރpR`��+Hq����r����!�۰�=�0ɰ8�&РQ�Kr� �GMG<�$H��d>u����*Bg��Dh$�|�b�:{3�;K�|�]�E���p �֚��¸���S��.btP�n-*E�H���\ӧ^_��1�#������&��Y2���!_�]\qx��fи��x����^��vD�e���l��kP��'����Z$��I*�����)4!ȸ/�������wM���t�!����WG��>�|3�[L�:I{������K>Yf���0�S�@ӭ�������<��1�>��01�O/�n��l��b6s�=N���x�P�x]�+�K��l0TA9F�Z������-�Q'��fKlMq/��Ӣ�@ r�E�QU�3�a0�b]!B���(%��,��b�ON��.�}���>� �P�ԭv�Z����K#1���<b������7
&[N¢������VT;�����m���:���E��4�I���y�	�_fF�Zڇ�f�R�Mh	4qAr����y�~�\*#�4Pq_j���e$[��[e����؅�e
��Ի�>)�K'42���r!2�)$;J��*Զ?�P��r@�OMw��xJ~=�,Q���?c�8G��-�����v�*Ѕ��.�X����L��mKU��S[�5���F�ճ4��+Aj��0s.48W��*����)��p�_ͯ�8��Kx��4�$���4I�T�0(��:�G��s�S��b��O�qN��*�;�#��6*Ṉs�ٕo��F���?|!ƫ� �T]Ʀ����.{�@�@��O0��M�ʞK����c.@�Y�sc��Mvq�,�^wthg�;����@}�m��*�I�������68E��Ae%�֒J��;����&���,�&�r��b$�ADj1%���Վ;�+��<��	c�O��A��Aq#R�I�.��.��ip�?I�3��	Q�\��&?�Z���"M�6S�uQ=p.`����C��_�䶦ƛ�Xj�4�p>���`�4��N0|A8b����&�`U��edi�3QKa"*���щ�]'Z�sﲷ���.�w
�O�N�I�Z�
f�L�)֨+��֏b���ݺ׃X����'��f�ds�޶�W����2MI�!`�	cA��z�}�ָ0�Н�컥���:�۵y;��>D��*�o�flӔ�=���-�KT���p.= n�H� �Ȇ��7=��O���y��Ī:��t���<ds�Mg�E�}v��L"�`V���@i'2u���1,�2��D�Є�r+CN��'�hpX]U p�\fȜ�(V��UN/��s�����f3|�Y���s,pb|yJ<d�O˭Rj��#��N�v��֌��ݢ:AX��Ҙ����Xx�d>��ώ���>�,��b�?���"���δw��
�>;]�kM�o��28�D|s����T!*hn��W+�:��;��ťQȓ�l>B��g�P*O�ɐ!a)O2�_��g�e���f�% ��y��/��*�C���������$'x�?j������s�?��̹�a����XGzX��mHo?vͩf	!"
p,�Z���r�QL��{%��.�R�O0��L�7�K�O;��^G�7�ٚ����"�9X���F>ԁo��X��f8�U������3'���a��N�����-W���q�=�ZU X�$�C~�DY���B�ק�R,�@;�I�y�Z�Nv	Z�v����ԓ��қ0�2L�#�@�� $�`{�BRYuۆ8�f	�L�WBh�XM5ʰ�RܨB\@�˷�����3���ԯWE\R#A�=mDy
"��/փ����-�n�x�闗�\�~��}��p��5�� +`�N�����lY��B�f�x����7�c��5�Jj��=�!�	��/T:�qE4���G��*��l���T��	�U�$�u�~7�%����0��<E��^�g\�a��8���O�/��cp�!�wI���q��(�?�egǐ>�0��D��!�k����<`v;��������ν|����BMw�!:d��ϓ+�޿�X���Uc�|�Afp���w��|jbS`�/ZQ]��Ia�Gm�j��5[��Kn����^Cj��5ݛ�X��d�_�>��PF�^���kO-AZGCVS�w��+�e�R���h4�r���9�Ft�W �۹L�/�ss��:7'Sȫ��1������%0PF�;s�+�ç�ә�jQ���P;��k�p`��E�������-����/>V�W�/���W��甜��[_���[h�˩����T�a&v*���[��z8*P�s�Ȧ��ϩ�d�4�Fr�L�%����8UJ�CMѭq���e�+���5B��ꮳw���ߊ+U����x.00�ZCf�d,7�"K��2��Kn���|���
"�D��.�tʿ��v�*��n"��S��-S P+m��IZ)qz���6(-��������e�k&8�yV��ǋ��q��V��	�[���E�ck�λ�)��=4]��R�u����hk�t������M�s'^}0\H����:��	'T��s�F�sA��E���0���>��gr��@b<��+�OP%�qu�D��
����s5�W�� ���k�c�W�F'qz2`��/���O*@~�ՠ+V*�iFi�Z��M79	�*�$�z,��tQ:���!ّ)C3^���kmzITa�Y��ۥ��8$�q�@��
i�)��X~�;֌U�tT9O����Ws���)a ~X�*�ݘӣy��粇���?a=xKvֲ#��~��{��Cfr�~Ze@�8᥶E�~xJ�b׿$J����5�y� 5��&�����z�zbg=!�����KF��q:f�s���S�4�yw�r��U�x����M�ܠ����Vˇ�3����ћ"�a���/�~w�.m��"�7}��|�"����Pb)#��5��rjX��ԋ�+�D1�
�%X�r ��!���\H�����n�����o ��R',���b�'����~����;���#mH#���O;\�c��ڻ��_�y9�7����X�M���Q�3ο&yC%���!sz�����?����	�ۘ�/Z
����@i!�@��'��ap)��4���U���R4����,rN�%��[�^�3�d�`�%(�ei�%������n�ָ�J��ɲb�#�3���]�_�ĆJ�쭼�W�7�t�g'O�9��D�f��"q�G4�|���G�
���YZ��G��I�{F2aL�=M�o��3ӷ�،�|O�(�C��p<T܅J\����TO|f�w��6�O��a�FU�'�:<���cQ�A�-��k�s � ĉܘ���߻R����Z��mxRd�Y��9�K��d�^7#P��`��W��{�v��6��*�FF�e<U��cM�C8"������CWD'㷿R����,�Ŝ����� 6�!�%I�$RP���8��d�҃�q�P��	�\E�˚
����rW�ц�L�YL��Y�=	U�����m����"�^G	��s4��~���~��+�D�.6�{]�{������<�M�'�o�=Q[��@�H)
h���g��7���+(&}K���c��-)�+������$���K�(G&�t|Tf[�m۞bcB��ݰ^���g�	�B-A:�?�'X�7(��)|���H�@�����.W�M�c������jq2c��s�>�@���SO�h~��K�=}v%P$uY���]�"���s�2c���&t��f*��z��n3�d�n�>Cm��n�;��u����Go����T�s��si�����'�	[��Y�穦�( �L�e<�Q��P2M��2#,W�?=�Y��)����k�@
�yW���a{�Gw((Dzᢄ��y�-��٧ӫ���N&�Ϗ�����I\6kW)J;��!?���J���ې��#3���0��â?�4g<U�t{,���B v�/�!nbphFϱ���aN�y��O�-v��S��}�?d[�����H�"��W*��H���E1{��|�S.����	��-�,#o��6� 5#���Q��aJ�AtQ0���fV�|VҪ`
v��|�&_Os+w��\��,Q�� 7sqm�d�/]\���(��?��+L�#�SM;��H�o�W���x�W��b,;����7mڼ:��[��=�S�'%��YBz�BKg�볃�ЙBr^�/�d0��.��=��縔+h���oj�y�:d(����NTO�d%��P���G�
���V3b0�z O�Wl8��Cw<�jg��Ȩ|/���r��'ǯ�F��WW���T�3�R6��Y��#*����8�5��{dHP�t���]���ǜ� l۵A����DS��g��gs���%L4#�~v+�{��W?�q/"�ʬN�SM>�c��Y�R�eƇo�2��Osz��rp��P�&�]�� k&��@CZ}�%�Z�-�!�KK�%�!Y���:�=:i��n��Zm`���`l:v�ۑ2��)�sѺ͹���A�D�e���wh�&�:�����
.1�?[�E��j;�9�O9�\�[�����3�0BY=��?K��]wV@T�9�z� t��B��ŕ�vwW40��j=-�@��)�Ȗ����SLl��$�0~�'��hY��z���V��:@��� #�"$CFZ�[��E���@�
S�j��rS�.�\�	�� o�'%DR'���l�^��5�$�7ǽ�H�ɒ�-ԕfPAW���AZ@�$Tq�j�<S�6Ɩ Fr�j�j�G�L�~V�[:'2]Kq��*|b �����J�7���F��Qhޗ�f��i�R��x{ǑuH6��d�t�GNWQ/!�v��జ9%x��/'���(�{o�B��q��n��*�v��@UK����rx�����@�/�<�$)S�P�
eW.>��c�Ċ��v�(X���]���[�ڌ�7�=^�C�h7)Y�����Yz*y9�ܚ�8g���X�#�(TxE�ļ�����؆~��ȗ�%�|��I%��HJaX كo´)!�(S
>� ��Γ;��(���[���u�ն�KvS*��3Q(���(3$�0C{�0�������Wc|&��
��GZ��O�ґ��6$*#���#��1�-�MS���:���u'C0kt�34",�6GB��u:"�<Cu(b�Ft	�����������n�:� ��AQ����M'#�&'���w��(�p/�2�]�bJ�~a�I}��R�Fp����{��_���yӳ�/��d����r��o�i\�A�A�ss��8�]��eY(W�f����������\=�ff�r	���Igit��Wp�����%��]���X��DOA�#Y~^'LE�R"�Y`�(�7�����V�_O��wa�����K72MJm#�@r���'������b������/�<���Fhf���YT KZ^c�`c�(v�/Φ�U��}�ؖ0{W8��Rr�Y�:��	9��?�)��ym��tzՔ�7���H9���F�݇1�NQ��✰`э�.x��jz%]N�0�E����:�CV��i�*^sC�^�T�f[���d��n-܊Yw��/�Q�H)���}
�<�34�đEu`��l���$��\�/%���^+hTvi	V�ʯ|*r~��5�RtE�j=[��h� ��[�����t�\���k����\5`w��kJ�=�X���Rl-�p����sz�
Z�G͑�y���+}���'���K(1D>�۞VTQ������.��!�Ӂ��$�j,�
Sw:y8��2տ�#�	q��r�HS�8ϗ��#N�������;���Y���
Z��	���Y��K>#'Pp��>���F��W*��T�*Z|�����d��7��:�d��R�b��,`
�9��<�J�Ǟ;���pq�ԡ���,�C������n���bQM�����X{�5�ˉbt �vkɀ��%�$���<��3�����l�������\D��_��&k�,�K -Ð�	�Ru��ο ]�.9�|nr�z�KtXn�\@ﱟn�(��u�� �τ3I����m�8-�V���'��%C����	���`RM?�$[b��d��@��־y��3[A�rMT�+Nh#\����Ƭc��Ӌ�[.mʿ�;I.��Z�L��E���cֳ%J�ϙ�Ž�����xM�ͫ����:6��ojw��9��P^�@�i�x�ҧ�C�v5��4�5�1�|lA��
$_Qzh*�rk�(��\�]�/��.�#tG����_��UV�YR꾅���2�甶H"瞧�����XZ�����젒�h�m9�j���l��DH�� �o��V�r������e�sVZ�vޱ�oGfAܾ��.�����(�x�3��jC(c\��呑#����KA��Tc2���:�W�$^^UjǾl������Nt<�)�3��2l���/Hg��~g�EB�z�VIc�dku�H3�Xd0 h�H�ǸHe�V$�r�ԟ�>�� �E?_�Xv�����[r�Q�z��c��H��3�H~�ݽ�t����Ҳ�ǌ�o���P|�2���֔O.+���ީ'n��^����KXП��@>�D�#&sҰ#����4+�Yb%m�6@O:�*���'��P^D�d��*d�6`�4������e
�|� �E �$_W�~�z�n��m��$-l��x��~�/�&i�Gb�"��âH��ڬS_���J��RU �Q G��N[ߧ���'��u�y�[�r��S��4��>�K%�g-�mb��0!��%TFI����$q����7 &o�-��D�/����}l�F�d{E�W��K����,��X���2����u�'�B���Z�pbMa�����'����L�%�\ר���&B����x��^�7�h۔�p�����!'^(j;35����j+N$ܬU&!��|���dn�Џ[��I��F�m���'��j���Gy���s�S��3��8%����kET���@���Ii�����Af�����w�7��f��m��M�\�r��՗'ѵt(���4�dN:J��ɜ��*wn������:�S/l��g���h��������b��m���{p���K8�p��C�̹tUnܥ�պl��ü� tT量��r��/��@���p�ډ ��l�B
:�ާ����e�
�u����t�h�埦�"M�w�r�fܝV��{��[���n�ӓ�峍�2�x�G�fw�X؄t|)�>�x���V[$���Ŵ��[�����[�rsA5���~���@b��q0��W�R�J��ͦ�Y��~i8A��`�c�P��1N��Jҙ�Ѧ��^#9j5d�T�����b��L�A���ؚa2-|1sH�^�cW ��b �e��(bV;ԍ�����ǍCH�j@��DpDV�l߯�Ќj��X|=���L^NMz�����,d�q�*����K��60�u:�$r-r�P[����<�FV��~�n�q�V}��}�?�������0$F�k#Ǳ�r�#��Z遶x�-z5�Qs�pɽZCp7�O�PD�>�]�o�hȝ{�����Un�]c��#y��zJ�m��$=W���tZn��q˾��籮=Mk��VV`߲?.8&!	
��e���̨3�)�9����o��,���!ӥ���	�]�6g �u�8��t��X�4�qZ�����nQ�ฦ��vi�7)/�6�S�-Z�A
#������|�[>nEk��w;h6*�юcCaZрRX�
�2��.J,�3�*�"Y�Dq2�Y����������89x�d�)��Bᶺ<�B���(}����H]�����,G��ᬑʹˡV��&��U�wT�c�[c+l�drۀn�b���J4W��z�x��Eff@�d����H-r�Yi$�8����D�*�>�c���s���@����6�������V� �s�fX����2��Ǿq�:��S�wZ�;贱��e�mb���Q���!���^0��&��Aq�X�b(�]����о��24y�mz���J�F�o�I8g9�����!wC_G�]����e ���HK"[��=� �HN�4A���z<U{6":+P��d�^z��a/��f4�z��Cָ�ǘ{S��Ht���F('�[W����Qtݨ;��Nԑz��b����%���P.����-+��WW�u�)��m(�D��J�L�����z�A�kr�'�ɁX#M�*w�)93�[��^$A������<hI�a���~�D:�䙛��Gv�����>��nԵ��\��o��\�pU{��褆��d����!we�ʽ�S�&���譭x{��l�)-�Ʀ�A�nN��d�p�Z�w� މ��/��:vdB�(����ތ���|K�������j��G�K���*�������i��/ {Ѿ �}. �8�>��k"�S����"dhy?Z��;�K��#L�؀G�7E[�ĳŰ�8�$C���,Q2`4���B�`�J�C�މ��IS$lS2�X�1rP���&k1T�h��7�)S~Q����*��.=2� &	�I�2am�¡�-r[r���ph�6��J��}S�'���#Z��7��ǹ'K�럳_�0�埜���6#�F��-�ŖA�-���`[��ֿ
�-![`ԍ���"�0�).�n/��^ŝ!l�"腁S��J����0��F�v.�]���k�iN���jQ�^޳b�FyY�I��B ��EG9�\ہ�hus�R�q�ȩ����kۗ?P?�vZI���<K|���ח�Uڰ��k�k7ўa�ns�<�ƬM��L��[R��ZR5+��/FP�X�j�*�NA<���i�䌀V��9�3�{��-C�iW����Ml<wX���n���#��
C���'����G���$Ys�#�53���CIQ���ئvR��,���;�t�kTI:r)�� m,�r_�]c��K|�ݣH��$�L51-�5؏�0 i� 4q��U����r0�l񝮲�xk��,t�[�D�G����pM#���G �A4Q��Lz�	��y�����S`U'��2.h�g����>�f����o����X�n�&�B��C�0[Z?����o�l-�,p+Ə6���1�aN�a������ =B^�	sǌ�����mS
��#m�����3M�J��\��x�(�ut��D���`�q
��]�5ߌ���uH�Kէ�^�t�|�1
杻Y�3���}�~.�6T_e%���lK��N`�dH��������q���[�T��3�Cb?c����e��J!q�9��6 ����X�%��&7�{-�"���W<� �/A��a�9�Vań[��g'�z��p�V�LJ���o�q�C��]{�d�3�w�r1 =��`��ݝ��rcQ.7��L4�6��*�Y���B#����<��~ځ"J�)�$GL|�7 
�����K�@�͊?%���|�K%�R�����>���kV�x����:�IC��ɧ��$b�s� {� xv)��;m��k��h� v�����aG��R��As���cZ�� ��k�Zi�I���#�o�g����5CUM��k���3'8ӻ\���$K��F�Y��.xz�q�i|(W�?�e�H-.zaF�5[e��<[X�-�ނY�9Zj���@�V;��@���W\U�V�a�J�Y�S�*Y�.a~�}xF�@��^5�"9�r��\h�Ǻ9��ҭ܁
,U)a��W�[��Wb���.���҂m��XnP�������=zl��i�dݏ�RWW�A��F
��2UH��!>�~���֔����þ����.��'���6Y�����`��s��M���]6�N�kh��a�<��bрx-p��ָ}���/o�����wh���]�ߴ tj�K�F��Ҕ���gzٶ�+B�2�݁��7��Nר�@�^�]�E��f�`�1M;%�x,��:�\`���x=�^@��x�Р�Y�x|8��Ӧ�C���Tym�sqC�E�zL��4E�����ٝ,�V>�؏}|Aa�g��NK«�0�2�so��2׻�=��,�֟�Yٯ�C�" �
�U���>�`y��.d6�Qs��2$�NFrV��N���Is"
�RoX�#q�
���
C\ݏm.���D���N��9����.�:fxo�����d��zR���+��,)���Q��)����f`+��<���6�*�?"�!x0#��k�Z�<�~d s6m�ÇUc���|Џ�5IG�w難��Wd�4�@��/A8nA�L��M��x�-B��SF[%"�oO�9[i�4��g�	?̷�]�y(*~Z��JnL���z�jK�:�0Qnk�ҵ��.��q���㉸�; �C�2پLV8sho�+��9gI��K&����zNY�䊪�JoH�nƉ#��ih1?�����~i{N�_PM��`c.�hɏ{��COȮ��?%�^�5��G_΢ݑR�K��/V,aM��K�2�i�/��c�?�qqc�lE��|r�%�>�_
R���e�����i�|�3m������U��O0�gk/Jגg��t�{�m;|��Pb��䤤�R@��D� Ʋ�iw��-�*a��,�8c ȑ_h�Ў�̶j&��@~�M���|�	Ͳ�T�{K�4��:����X9G��*���Ծ,j�S��Z#�g��3�?Z�dh�_wO��l���Ö�֗^�m�uv���Vg��р��Q��y����h��B�)�E7]��Ĝ��c�OfSe1� U���<�㽸�Y4X�fys�P2�e%���m��o7¼��8�<��9��
�8����ME$#�d��_@�����%^�3{��cڿڊ]y�~>ì���Lw�-T��U;�.����$�bkXB�"4�N&>����P�ݥ���ut�C5�*�]ϴFp8���?1��d9-����,�s����o4x�'7��7s���ł�!˻g��#nV¤��oj�>q�8�b��@�)xݏ�q��gNG�������|���AIn�~� .��.p��is^h+�?,���L�_V�u��,�Av9���ӫlA���1��;�W��X�*`�h��Nu�0���3�H���p��j)Ω
W��ܻ֊�n�T*Ce�d�J3ہ_������]g�
0�fK\���n��0 r����D�X�u߉mԵ+l�I���UK���/�'@59�</`�����V��%:��	J������N���wGU 0�5�ɇ�l����1/��_��U,k�{�Qv�D�2����ztM���p�L�t���z�dC_��K���1�v�/.��K���Arz��B�����}�׫��.gބn��j�����p{�*�F�=��q&��Q�~����
��%~>���U�~��Bi#Q�Rl�l&�0��{j6�c����Pv"�y�V���Eq�ߺ�h��=�i �)��F+"˞J�����|���:?{�afUs�
������	P��P�Y�9��V������b7^#�~C������3���4����~g�b�Ao�����-�r�1	�Ux�c��KA���4�A	����U�cחֱ�g��N��G7��@=�w���9��[�AM;��2;��嵅��\@��x�	����,����o���~f'm�j�ᚓ�����a���N�~����ǵp��g0��/ZFľ5x���p
�������t�^N^�"�I���FeR�l�y\�>�>���:�\uav\���VEO���_���x�.�K2����D�"Y��з^*	o�-
Ҷ��Hu��où�H�W%��N(xbG2��U�-N�/v����	���~/	$Ѷ<�����~�
l��3씙Vj�w����4��Z��A�@��)�7��Mt�j0Ƌۓ�@��o�\Pn?T:���Ж��+���x�����uĪy��ӡb'�<('��y��=�ef)�5��� �@���b<�w����9����+���H���!��
|�*����9M��0<�;�!b��x�e�f�D�,Q[ƚ�Q
����+;�&1_P$��3)�DXP��?<-��I=z`��P_�ns��|�X6`�%�:��  ����Q�/��P� �7�Xk��^Al��g-��d�tピX�0��ԑ�4�y �Y�����]�CU5�'B2*֦�j��1�D�)��P�� ���V,�h�C,�3�i�����\h@O�1�@�V!��_���"��I�#��4�M-��Uj�T%�O��WK�hO����%r0��f�%�0�R�h�>�l(=,��@?3?Tq��]jb�ʋ\��36���V�R
��?�^��ވ~(��p�a�U���SܩA�k����/��}UK
����'�ݘk�G��w���4�n�ߑc��X����B���ղ�*�z0���X��u_l��2F����h�B�����?t�uf��AR`��{;�*cDMB�,��V��R�lR[H�P0P���P�\0�c�=H��Äߨ�(H�10*>��њ�����)A���A�4n�<0	�>&��x�0��P�
;�!�:�}ba��4.��
6T�y�UT���"�&t}��ˤ�1)��̋	p���)3��YĀ��$��bP����okb�HA�Do�����r�HktG/1�֖e������%nq�.�fhN�]E`�8�5-���ܠkX�O����x�,fD��h�0��~��wx?�ԃo�Y�����x�o$�'"���O������c��yN��z��Iw�(�#��͈wq�qwD�E�z�\�s��o���(�r=� U���/MV�Y#Q����ϻ���a�؈�	�(��{W�d��^��V��!Q5�C���^�gY-���J�������G�=��'�2Qw�C",5$s�,/;���tHY�ɲ\:/�$�Q	����c�ߛ<a��F-`Ve��-O:hn�	��@��,�R���jH�! ��er���� ��m��-��aa���:s�����K���z	2�7����7����B��v��-wx���L�![��UY�Q��AHE<�;
a��`������1^�/$��`��ZXp3�9�Q�`f�A�k��x��h;�������=�n%|�L��m�k2���R4ld4�{@KL}1=+�\Hdq8&յez�Fߕ��$�����1d3>��os��o��1�4+�)[=f��r�����e�l\`�z=XᎱ�ܻȤۥ�-��u1y��9�b ���}������V�:�>���6]���@��P����`&'��vꝣ���5�Q��8��٥e����͛��U�3!�0�3O�:�M�0������E�<u�;��R�v��X��+m��#U�`�u�.ǏJ�	�	��OJɳ����g���+0� y����׃uՕ���=c���	d�&�.���BG�f�_pewh�U�X�!e���\�lO����w�)g�8�E���ܖ�2P~��tz̫o9EAh�SlX��Y@��ڴ�}��|"h�BoY� N����N)fq��[K	��w%�j��u*���FO�F�0�:�M:��7��5h�m;+ͣ�20sE�D�Kf�:�	��������J
�j�e�D�1-�C��w���ф���n`�=F����>��.���NVk�$�m�4n�Im�1�w2��t�T踫������O�ɟLm��K�E�d�m��N��B��[�ir/i�u�WRjb�dX��x~et����"B�0bѱ�[���A����^�D��_�`W��#W�j�'�_(��f�@��ڒ�W�C� 	���k3g%��X���P�
h�����d㐞�D�A!��	׶YM�*�ɯ���ڸN{Jm&��M��J��Qf�މ��\i��������`n�JY�j���z��"��g��L*�$�?��Y��;�|&&q�b����O�	���nQԇ���z8��eBɪ�s��)E��%#�Ze�l-��H�a�#ſ�I�ݘ��Y黷(
h�@�|�:��Iʖ'VSH��ty��d��8�Q��d���N�d6l^�2��K�;�E��8�����mǆ`�Ɏ0���?����*�X=�rZ������ΖU�s'�}�L��]�+�Z|˒k@��ƽF� B�7��{H���$�]C��ot�a/?f77����5�t׊˭p��"�½�ʯɩ�m^ݶ9a��9X����O[�]�MV��	�C����/�z��z��N˽�ː1�y�ܡ�'m��J��U`t�:L���!��1���J��Q����`6vENO���d�:�����!��� �b�":a��c�zpL�u��"�V���7#�/��oxτ¼]����O�d��*72�WA�E�� �r��Uo�]�{��j�š��d��\�3�G��#*]a�z�+_��)p�&���_�\���A�V<�3~�9���vM�,��ks+#a[0�+u����K�:N�V۬P]��?�i�
h�"���c6T�.�:u�#�A4G����.���$0��@+�w��W&"��d��K$��U�
�G�����	<����,��v�(�~{x�[�*օ����b� ������wXL@J]k��E?�@	y�-����do�eL�+.<V�Ls�_P�r��v V�e	ٷL��r����Q��I7Z�RI���S?0����b:c���H2��]ZO!B�s��u<oL���l�9\��2��ݠO� �<ԉ�"ٽ�)ilG�r0M�^�!�d�C��j�^ڱNV8�~֐a�"/X�r��0���m���IrN�6)VU�a.�y��=��cᶣ��L\J=�	�D��]p��Q����"�*���0��I^C��'�5����M5��.e��V���;���)8X�k*�):������sG:p������a�o����HvWI
X�A��!�+�ߤc�\��*��0��Raf`#u��<�A5�E���{k0k��9Z���ߝ&Z�l�OU����~a��	��t����=������A���۰��z����}mnf �܉�2�o��vgR�UxP-�z6��@��j���@������l.��O��O���b��H����C�!A'9�����vOڟ��c��?h|7'Md�v&`2�
�C��8�E�1"���o�,X:nGA�PX�e1�l�gY���PO�ʏ���>�e;���×�:�%0\�д3��|N�\��X�?��������Yc��wu�D���H<f�$��-�K#�WU)���~�WB�ts�EE��}����0�ġn�&W��X",�t�93�}g���!�񶟌��]ʳ�vx���Ð#�i��B�c�mG��ֹ��p��z)3]t�;?��wm���+SZ:�h�@�>���؏Q=�}�i�e�u!�(����c/:u�hry7����3{�2:�MQ��zl�.��__��8A����S�M�t#�<�ڋ	��4(����#填�k�e��\C�m�)�$����h+�V�+ =^yǯL5���i����LVy/�st�;�l�p�KVA���\��CB��]f������3�Ȣnɜ��b�o��g���M��iv `��q�f>�3�PƴlG���U�.�m��Xv�fkȣ:�����).���@<��7X�%0�w�yF����"p�&�e!�T��D��{�q6vjT��hY����1�4�&�In�#���@�E,��tf99M.(!O�vn�K?6����NuqH1D2)�/F/BM�A�(�ql��!��@8�5�1ܱg��K�[���&��Xf���9a0]�i����Nf_䆬&(k�#Z}��� ��q��s�����A�tK�e�;6w��6�"'5Q�e��Q��� w�k �0�	1���5~ ��vꯜ�}YG:>�$�=�Vl�8�����:�V8���/tけR�`��|?�E^��bOt��7=��ȉ9��i�pʁ���>!�����2�}���.0�
�5��JxMCBx����������ӵɭ��OC����^�K���|��Rx���|��ٻ����-�hê�t�%�M�kψ��9Ck{�y�.����r�P4��e�����)ԛH��Ѫ��!�#	��S:���t����p�&�RO\����'��D$���K�t�eST��%��L*��`	�'V7��g��m�F���
q�Ե���=e�Bu{�C?�>,���v宪�H����$�8<p�.|�'TjX<S�%cal�}#ka��(����1Yo�q5WNҵ���0�.�{����i�fЎ�޸pBٜ
�t��?D��HOo\���f tC����'A����{Q�Yo]�<o���7�q����P��Q+�yh�ጱk�/�i�����ja���?.�a=4��(��u:(r�+�4
���V��2�%C�A�pu�=Ų�?,P�Q��fte�I®�BQ�&��&�B;��܃A_�~�8�t�1AD�h�I�\������N�q)�
d󣓦�F�"{�	R��s��p
m�ҰmQ�]�K&��»��w�Kk[��&W�q�;�V��l�j��4��< �<4e�|�U~��B��嚪+yY���s���4s�ȳ_�}�ٻP��m����x�`G�TZ�Г��h�N����!�qY�J� ch�-�����G���j�����Yg3]����ʼ�)�Y�W?P�P�3?+@7϶�9��Dt�"�Ѕ��G�����Yoh�o>ܦ�0�'�,N�����Ĝ�^�pt�C��F�Q�� <����-�������T��uT(�2CЅ�H�p�%�hn�x4�49D�����e�[0��C	dUu�m������'l
6�Mܑ�� .��^���萜���?ڲ��N���:��W�&cTz���E3�U�e9��-b&Xg�k�$���~��Ёo:`�����⳱���O�B�3�G�"59">�V�C���u%�ǀ����(�nfe��!�*j�5�>7s��L��>�a��7Hj׹��<���H��J���y���YЧ�v�7i�Z :��5���M�3ٌ=�C)�	�UM�3Ob����v��5Z3��\��;'Ņ��Td� �ۣq;���M�u]W�n.W���\��>X'�9��μ�Qʘ~�һ��~��`������jQ�^͍Z�an��2b映�y�28�C��@������;�)���{P�I�"��u���fv�Θ�t��y�m����ğZR�&Ue`��<ҝ���D$����� 	
ʼE�j�S�O���/��a����l-����_�u�'׹�x��a��I��/
ͫaS�ɸ��A�V%g!͆����k�~Ċ��<҈��KO�}���.q7�-�%��$ŉ�5~���+o���'����(jahF�UB�o�:e�,}_�ɬ<S?~/���So֌)��5]�)ۆ e�hX����-)�Ij�iT�c���D��p�Ď=�H� cm$�qʦ9;�
ٕ��¢�C�EEe�R�pjŴ��aG�gks��ɏ��߷y��-��mc�-G�X�e����̸��ޡy��=[\U̷�����WK��f@�]�谛/���V�b��D�p����EnN���FTtKA�(�~�\}ص�Y[� �q��H�;ԟ��Dn^����a��֒@�֑���n�x]k#:Kv-]%���yT�8{��������\WUwE� t8cf@�ln�(^�Ѯ�%0)��N�&�d��}��T���*�ǚs_.����@������n<k4[�� x�bB���:�Udl$�~Ax�� �l��8�%f�B����ή�-+��L+��/��Dm��� �הYJ��h��3���4�{�����S_�76�8g�G��IQ�d��*JC
7X���l�Rd�s��Ti�M9Rj̟m#z�e��GL?�ڦ�-}$(�˷?��ƂòF�H��ӊ�f���Iن��9�؉�x��:3�|����
|x�_�U7=�hs[�A��a����ej_�L�[�\�B�o̎S��g��h~�v崟~W|�;�咬݋��dΥ����bs2�+׺<u�e�7����W���d�?����2))����~0)�
�#O��Dƕv�2sпZ���>XTgйfvܲ~���O��X�8�_��S���p/�$�젻����<�6�U����D�4�r?�B0��<�8���ɫcE�\wP,��"�qҠF�Ĵw���,~0�)�r�{����c��|�`F"�3�y*��b�_�ԉ\6�-h��}N�z�����2�����#o|�Z����`���B#����6��mȯR�̻]"ʨ�v���Xм�c�8ǭ���}n��6B^m��Ƌ�=����4��O�A~���)������F|���²���fkH�Bh{��y�ki�K�d�K ��єe8{Oo�-�u���B�btZ��-x|[9{�Y#9�X�L�		C�=����1�{$K���<X`��Uq���[���vR�0�`��=k!Ua���r�.�4�$T�^Q@T6�z����_l�u��N۟0��}���G��*��g��#��|�*߾o�R(���82I z��~%�B�o����9.�v1���G9^��:z픘3�2��ϖT&�:-��4{�����5���9X��v}��:�6g���v��!��ډCߐ����� �ل��}���Qy���YNM)�FX�iX��f�$I�*���/�XA/s�ޕ��w>�Am��.�m����%*>1ݐ.�{`Pv�k����S!��#ˋ�m���j�m'�n[>i���H8%F�C�/2�쥰D��we�$��X���"	0ٍ��a��wu��t�]m27M��'��̠T����ց��*�O.��g-+>ښ@)e*)�|u�4cF�l\�g��]C�\pf�8�>�	���NY��`$�i�9�H+z�����$C��`n<��*W�A����o{ɭ�(�L��OB�1�r^w
�!�"�1{��Ԙ4�X���SD��#��|ŭ�����!E�u���K�����&�C�j�*�i���Ϗ��!ܗ`�wZe�j�9Y#9H��ם{WQ��#u��y��6<�.��0{^�9:�E4��pb���<렠{?�~�70�ثe7G��dÜ4�k����!��/�y8�m@���J���{R����Q״I�y��5�*l��ړ'�"Â�*�sW���Z�_���0��y% f�0�2��KJ���M��'�uC��눕h[?���~��i��|wI��r- ���2�ZN�3)絑d1�t/A6"(�GD�I���!M�X��>c"�A`l0'g����j~D�� S�����̩���b��*>�z���no�c0_ �������Ȩ�ԊcQ�ܣ{�E��߇�8�Ɉ�D��M'Oh��6��֙�0�R3�{�D�z'Y;W��F�O�x�� ��J��{�2s�7���Ņ裡jR)�2M����Ů���wA/�<�y��į�y迍��&���`����pHI���f��R��l�)�4!�f�T[�{�0!Di[	cj@@c�� ,�9�7�\,���r4���H�����mL�wV����;0Xۣ����P��k��e�#�n{dy.>O����\,b�UC���f"^��#iT��3��E�:� 8��}���< ��>�m�Q/�_H��Ǘ�y/M�S� ���
�ٚ��9��m� �Z��2�h4��B+��x�[/����F���N�����s��m���]u�6��&!�BY���5��8a��
)�(_EO�q�g��yKa�?���kׄ�����>�o�?��]�;7��&������dE���ůf�&Ht�j�ĺ� _u�c��u���O!��x�ل��,[Z6�=���3�r/bA��d3���t��]����̊��w�5~dxt�ro�z�"N�� 0�nքC�ܛL�<=ot��I�y�1cи!�:L�a�#u�\? ��[�b���-��5(�!���t��l�$� ;����Ҧ������N��k6/O�q���Ý��}M/��� ��@�LH���t0n'�U�����Ph�G��
cҞ��N?������%�3�4I��Օ��Tmq5�F�Wo�{�P3��96OV���ՉgH^�7�ߧ2@��Gz�z���^��-ۥ�WMB� >넦cg,G~H�Qi
}�X%Qh�ǋ���THY@����a�a�iw'�;�������X¥�x*Z���W�p�!�,��E�>���L�Sĸ�q�Y鎱�L#�$�F6♈vB��gb��;��B-��$���ئ|�z�_��`�l�RaJkx�#�!X+�%&��ڿ\���nW �A��o�X>�^݈cnI���&��Ќ�xJ��U0w�ۦ��n+;�w�3��:���3-A��=���T�84%K��˷����u�!Y�r>Ox>r�Jj%(x�������b2�l�i�?��[�t������t�%�� Ø{e|w�һ�E쀧�"�� AU+����[�On���ԝ�G5@T��ubxl�A�e!�,�P��5�w��ʿ-��<���ڝ�V�����D��s�_L)�٭���ZבΛ�س��Ky���LI���1�s�me��珑"�e�R�
>�Ye�<�0W1?�}�b�5Zġ�[�Q����w���qAx!D���s���Hԓ,�S�t�/�bT(o�=e;e�](��Nq6�h�=��Xޮ���;�9��T�.;�u���zf����� �P��<��v��9W��[T�~᠈�$\�.�Q�:"�gy���ɢ6Z��2���z�+I�ߒP�轀: ��.�ߎ��j�����_�P�&���`N/.r_�kh��L�q[~u{�. V-�|oh�����@Mh�צU{xP�w������Q��B��%n C��Vj�_1nz�Y<ɅH�������ֻ#�d\BO��e۵������^]�{H4��(���C�>b��qWz�����7r����F��	�y>X/��@n�Gqy���*���>�F4@i�b�
�Ai��s�v!�C�HL+����5�{�{���Ǖ��`F�?�T|j�c�ʙ�1��u =�c�̛I�3T��a�x��wW|5Ԁ8���}s�(F@t�7���W#�ba���RLC?^�/��0�	���B�sFʽ�-�r$l��J����L���Jܴ�Z��K�x]�3�G�˿���i����aVE$"���'l?e$
��;�.�ěQ,�gG�q���|~ݢг��>���ߢQ��-��+o&�IcsZS��ڑ�
80�:F/P㕇;3B��Z �}t��'Gv{y��npd���lg1<eGS""�ܔ?hp�żf�6��h�ĒRPi��f�Z\�_ܕs�:��[�X",V���ӭ=ht�8E:</g2����I� *Xn*�D�YNu�/`��p.��}r��\m�#��-�&B�2�k��%�#�\����D���cVu��o��Y�翮�eb;�������n�����������vSR���})�w���˅fgP��/���0�̫0H��(E��F*�vd]Y�����)Z�n���3-���H3O}�Q�ܰ�ǀZX�BlS݂���=�8�o2]�qv㸭ra#�*���mN�-u��5F	_���zhom�.�o�l�f��{�Jg�}<!m�[5RYa~�=)\l RW��z����6�-��E�Lƣ����X�9�*Z�B�1�u�r���lS<�iu �7A%�5H�m�k�)�	,j�y-8��yԃ�ݭHheٳ�Q|K�N�%���(i#�C��`�DS�{Ev�Ӱ��O�#��֋SAU��u�
��Bw�e���(]�5�0v��-*�;)\?�K#�˷"��k��(�I$�����"
����o�����(ѳZ	����?�F[�X�{���K�/A㚲�؃�u��X
�L	hj��M�@3H�!�mg�
�	�JI�����V�	��rz29�i��r�o>s�qm:�dy�����*�&�k#���ŉ�_]��?k��p��8�j�:Iڨ���/K�IUOC�B�{	��2�b���{kXK�{Ch��@�	z.��3��(E%�G(Vj��H2��Z,ڐ&��� �f�Uw�1�bG7���f$iX�۶i\py�s�e }%+�B8��
�I-\5�eX	�B�����_�.co+ �jF�x]���S3C�_F8�è���%N��x����(����=N���|���OĞ�A[Z�q~�:b$�?�"3��K�^����݁�`i�̔O�z���
�_����k/u������(tXޙ~�7FQ��B�޳;(���AFI��Y�D���uzo�C�=�?{�C����M�d���ĺov2Z�ڍ��l���Ot�ݎ��B�IM͕d㿲�i��p!D��T��Q���7iE4��r�.��i��4�x+�	8���Q~lp�o�׋3���Y(wǘ�Ћ�C�l��JU��IE.�IzAD���t��{{62-�B6�r����#�{ }���X��|9T�L��/����;zT��fuwDpMg�W���Sė���n,��]!�#��D%���/�3	�F����ʴ�z�a�5
�f l���i�0�=Ұ)�� �"`l":c��G�]tS�9���w�Xu|�y��E�h�U�39����W�K��F�Y��(�"�Kb��q�]����݊�L< �^��*N!��~��/�KN��r3�+&���&R��D��;v(HU89(q� R#�f�)�Á�4B�v�f/m{�ˤWv	�6����]�ڂ�4�<dX�&5����L�v��ẁ�Ѧ���)V}
�!��=�� ; ��@����Ѹy�1��(u/Dݵ3݂�Ñ��"������P��ϕ�vS�;5a�]0�1)=<p����r
�#�ԭ�F�`����/�M|���g���9m5�<�˯eQ�a�3ᅪ��,R�iP��f� ����WE58�_}�������ժ>4�������ahA6��S�?v���l�,����̈�0��o2�W��N�_X��,��.%�t�q-���e~|]�
1ґ��lv��B9PVI�R�;t���R�_��ɇM�Ry���)�.�hM����K���%#,���^��������t�o���0+�P#_�8S�9�-	}E��9�����%L�4�뢨�_^p:�~�Mgx�o�/H��W�/�0r|%����s�Q�?�V�7"�Fh�X���P�!@�U��m�2w�i	�U�^<�z��]c�\��}ګ*�������m� �"�Yh���z��x��o \��ٳ��k�Y])1���	k������%����9ô��T;J�:E������+-/����KY-$��C��Q:���I�K�����U���3k����[M�_(�/cl5���OhL��M��s-G�!�q��Jtdb;���h��4�d�/j#Y��)��\)�L}�����[u3�=�Mr܆�� �	[ªP41��h�zi��+�ù���wN /s%��S�t:�b�>Ʃ��'q�>6���غX?=��(Qձ�M��
���9�&��5��j�S!����}�Hp����������`�S�|$&���a!�i��L���c.?���h��'Y����#�`Op`�0nM�ր�Ux�X�!�{���JY[
�ٓ��Ѩ�oÍ���c��>��m�t	�	�~�����w�[��.���#�h4`��<������V����dV���ᧂ�A�x���q�(�n�S((��$7���*�Z�=����`_ߺ�Q��]�m�c:�3Q�d���8N��Z���{� 	��� �ɧ�����	e~����2Ѯ��j��w=?�ɟ����7{��$\�c�Y���K�]_M^���������>�¹h7�n�� ߍ���,["q8e�쉢�=�[+�DH{A�v��f���>����Ƴޚ V_�
�DGJ����A��)��'ĳ����V�)��~�Cg��"�0���Hs �5�~)��hR}&xx���^x�*���������v�r$����F��{JN��Q�}�P�iG�Ќ$'���p�R�Q��}�%J
��ʭ��UUh(\�X�^��W&�d��
�ҋ�9zj�;�0������p)���	Eް��%��"x9����>KB�Hc��U&�3ň_�$��[����Y��;�_D)g2���{��@�u�n���z�QBd��798z�"�~�3q���J3��
�����^ث��UL���5���IP�6,?��K�v�koS�h�)=�P��g�c`�o7�ǙNy�����-�a�~	2k�?Z��}q>j3�N�{PF0,O�f��`)*��R�k��8��׈$Aly�en��x�B��,�.��l(��-ym,8�$$vw	�O)� ��\s�g�_��)�&��u��q�)q��)�n��7�`�����gO��	�4���Arـc� -%ͳ�%�4h������8|_��GkRΆ4��i�Q,�Qұ{�Mo�l��C\�\�\�F���y��IW��N���b?�P���h:&'�u(��+Z'm���T7�a�_°v�M��ZI����N|�����Z�����ige�Xa=~�'gB1��/�1��̗�R�6�U��iX�"�`k�Dp3�V��H=���W�;�<\b���~ht��3ih�pS$Q���9p��������[	��˴w5f��i�I��8cƼ��M�pp��G��ϕ�l�(Vk�/�dVo���k�N|���g=4s�{P���?v��C��V�P�-��?	|:1^��O9S<�M�.yr0_s����愻���$V3���C�6d�,����E�������n�00���0R5�̪Ua�牢qbx�w�b��G�2m��c# "�
��iԍ���l�"������a�L�X#��c����,Ӄ��U�k�2�zwL�w1��y���)D�\mq�3
��)�n?�O���"<!w���\.��Х�U�8bJ!0�|���׋�e\�>��l���{�Y�!�5�z�1�mKB��x�	t�E���"��Z�������� L�4�ㄏ�q?��!�1�BX4e�J��&V�v��j9z�t���W��1�?�D���Õc���U��p����#8DJv
:�;z���_%���.R�,�TbA�;%Јp?!�a�B�^�q%9�ʻ��7����F���U%A�k��S<e ),ј:�\^H�i�Yó�(uh��5���$Z���d�Y�.�(������׼������ǌ%m�w$Qv���qAz����9��40���92ĥ�P���R*�%�][I�C���/t��J0��)���Vq)�n��'#}ˡJT�"3gsd1��ն��XlK1�bTa#�}P�R��A�C	"4.�Q�^� qH6NJ��H+ŞJ%�3������=�c�%zS�|�4�����z,Ꙕsr��l��7�&��W׋��.�V�?�-��|���"���"��}����n����@@=�]_5�t�VS
�*o��J��lM���,��m�辖	���ϯ$�Z2� �?^�q6xG�{T�Z�1�nFMc�N[�����s�]�0�������j���ؕ2�s�h7Lf�.�.$��D�䢨i^tGz^��v/�n<ԅ�4j�c̘A>�~��Y�z�,�u�Ql�w�k(�%��6V"x+!�cɻ���.�Ǵ��\��	�f�������ߟ��Y4�<���7�$��x��]�s���+P���Xi��;�J��.kp��MP�q-Fx=u8�C�?�G0�2yM[��JK&^{#}���k{�OT)ٷ�p��$�(����"�!	���'���n�YЂ촹��|�C*��PRq�2�5^ћ]�/$ªt�:S�_�����8�� �5��5k�3��	Y�j��+"F�[e�#�7h$8�n��"�Kt��5P��-oj�԰�ֲ`�r,�-$�J���~"��Q�wO�v!�rR�h7f֏"���.��Z:%�O��ŷ%��]�����l.�[�'�Q��
�5_�C澴�>$�w�Z���4[_v:�����I�Ν�[�
0Ͻ`�ld�
��$��|�I:���uݯ���L���:P�8��@����,��ݚ~�2x����VG��X��tA�����S�t��%5��3"�>�}�^�&P�-�Oh����kr,J�n(�����C勠�n>c����DΆ[�^�]b�o_�0L}�?] ��Qpl�!��W�Į�{�Bi亘0t�U��}NX�{d���� �I�\]*1�&8�]PT�܅z(+	��z1VA�e?{3��������h|誩y�F��Դ�jNL�kE�$�up@��[O9w?c���F8� GD~ '�i.�E�bn)QRk�e�^���kw(�M1qG,�l|�x�C�!��:׌�M�f"t?	�ڭv� ˗^�r��HT�N��D�5ab�J<� �I����)~q�Ξ���k`�[�`>h�����t��>>ıF� �J�f�H��?����<���񩧲c)�EJ�M5��g}�5m�ӝ�Ϥ�[}���������]�۠�����3wy qܛa\>*�i�S��}��&�%�k�B�Ӕ�$ij��!��aa����h�l��@V��S�2M�y�	ַ7���
�b�U.�$�9DJ1q=0����-i�����4�V����J��7���L8ȼ˗��Xڿ�G1�
*��z�N@[�~y$�w��0�Z���Z&(��v�4*�R#�x}?
�u�j�A�A�g�g�%.�䕌���J+��!����I5h^��J��G���{�=/�%MJS����i��}܆'��6I;�XY��V��qv�=,���_0P,��
�Tl@������w0��&��q�X��0�@^n����Y!b!����'��"E���K5���P�^vc��0Q:EДW���p�nS��>q��:_rӆ�4���<��.T#�!�G��Dhn���d6\����-x��y���I�i��P$�O�!/}�TY���L�O�{��e�pa{��fM�|,��;&*��D�m���G��#��\muBM�p��u؉��/ ��nCƯ��.o�B��@�yu�χ���ē�'F'S��6	WԓC��^�nhJwQqI�&ix���&��Xz�d�p��`�+r>i؅��?2��Mc%��;��a�P��3JC%�i��N0�� R}t}��X��'�s�Hr��	
�N)ߚ�!�τ�cu�$�µ��	P�s% z�[B0Hq�0PNn�%,"iJ���z����N	��:�Mɼ���	�N��Q$��r�R�x�,��((�Xo4v�I�Eg�`��Iz��֚�.�4?j呀��ſ$M����&����#|�^:�k0l��Q��b����@3EW��fNdOjkZq�ֺ867��Q�G?�&I	�K��e�fCr#]�k��������[A�΋!���&�����^5p:�?�J׻T:X��x���4�Gw��<��B=T���I�9n֚@w�pz�tKs\n2U�V�yM'�$��g�,�!ڿ'�w��,��偣WΧb?�$�兌�%iOk�}�+�7�p<U6ٹ��}"��.��5Q�	ө���L����,��ą�r?�F�[�-�br�,��NV�<�: �;�9b�s�gv�о%?
M��)u����Y9�V7R�+��;_�%7i0����N.�,1$~�(�{��jM�wx���^��fS�=���c$�Λ�ߗ�r��9�,�7 ���?�Wٯ�#����I3|��JЮ�S�K�r�[TM;6 g��#���5:)8���_�bڕ,W�-�����>5��;�*I��GPS�U"s1ZAm2g�ەtǛ}�v+)��9�KU�8�F$��]�;��M	�Q+g��] D�v�u��7��G�p	�f��`j%.u@Ś���#�������(]��J�΂��b�g�o��
5�-�M��B!w�=s���^;�G_n��)hBWo\Bd*�q����	�G#�ݫ��&�>?m�vz��.�t�orqIZe�� ���F�KI	�E��sT�uV�[5FA$;0�$�y@�wX�c. �jʑpP�u=���c�$�����쨐d�
j2��Bލ�����e�e2�gN��X8Ճ�����5DN"�9�N7�I��!��2?3���x�dd�E���b�ƽJ� !�8'�z�eDP��{m��o<i0D�BT]�#���o�|�U��~kP�<H�,g��h"WPP�ݨ�����@�T�J��f'�i��b���H���VK",��x\��ƇU�g��f���;���b��������-+�g 0A��q"vݣ�Z�Q�SqN����)6kZ�T\eVw����c�P�n�hp��� 5&
���NE����ppZ��P���
�&��j�[7��(��r#�F8O�$I��3������*�O ��^j�+�����^,�g.� g��z�jmQ�-�1�oV�fh�A�V���]�sRW�'�IB���o������O15zJc�]MDH�%���B��>����:��ďZՄ�;�c�k��=Q�{���D[�a�WfDY��A���O@��!ԫ2�).R����tIʵ��q��ۺQ��\K�q�w=�:�*�>�K�R� z�R�u���Se�H$�k�8���ZU/����L�;�C4��(*�M^��@K?}��<by@>ae�Y�hT4��խUd��[�5^+�SF���2�f�Y���St�LX�{���		.��|����-��Z��uQ�@<3C��g�^��u�I���R%�/Q �,L�$#�ǝ�+�d�x{'���^� ��M�:)���|"͑���9#'�*>��'k�REۉ����r	���3�kT'���*����;O�q�.��C�h �9�j�fV�.�R�oF��X�}��By�؇��w�����!9�#���Q�d6�r�5��R�H_�6�2M�����tX���8�c4�Uj�Fer2�i@�Ti@>���J58��rFx�������Y��]�ϮT~Ǟ;�,��[P���k+
t2��Ѯ�C�a�;��Wb�o%l��5�TU<5}��=�
�шwJ�'r����yC��+�k�|�̕�1�E.��[Gʜ��b�f _�~x^��t�c�9��jZK��.~q����^I�ʾId���"xC�׽�&��T�J�}�������ﰘe��p��!@�D-��G�5/�;@�"v� "o���b�&���(tr�z�.ܳp�*��0zUP1t�x�W�E��Pk)�p��P���7T�MCHm�ء�h>��I��6YΩ;�I������=�}jD�6�VI�cF1���ܶ��a<�l\	s�;��/��f�ӻNqO٥�7�1�2~k�-�f�������S�tIҹ����j!��!;���\�g��9�X���X�+�d_A�IC7����c�p2.Qѩσ���ޠj=[��e=��h&��مc��`�y����ſ�KU����%0) �t�ʀ�ޥ"�=��h9������J��4��#�°�D<o�ե�S$>��ns���#O 3+!@���=Ł���l&H�7V]I��W�*E	2!�SHt�
s���ڷ�*�~�NP�X�1�T��N���d��\K��?o�q�����,hD���&ٕF�E:ݨ��EY�`=�X�>	UčlDɍ���t�n���������u6�w�e�ځ�Cw�`4�ot�����abX�ܢ��m����]��?&��:�o*ň�%��+��e܈>��]�ƣt�=��T�?�3o�U�wu��+l�ʹT�j�
�ૃ��a��QB��(2��V���s�Ī%����c`B@�����g*��I(Ɂ����P5~c�S���I����������P!;�G��c^�l���`�!���[N
2}D�:�8C�(?\�����S7apÍ�>�Ws��Sa�݁�ܨ<w�����4U�� (
Y�˄B�P4犽�T��U���X`����j
@:�m��W��o��=9d��l/%if������羳���lT�^� {�9�<�+��<W'�Yj鵔��by�bG��(w����D�D�*��6 ���$��aIt�˞z�|ض\p�f92��󄡈$��x{�J܊%&j�?���G4�D�4R�}UHёG��`��s�x]� ���;��Mj���>�}��@꫎V����'h�:��R)��X�m������<"�� ��%�s�;˧]�:ɚ?��O�*Q�$6b"ohyM���y*�v6�+�s|�i���a�7"�阨��GLM��{�a������V�jO�:�rs�Z5��|��m�0f�T��CIo�9���t?t��Xơ*��`�#�@��R�j�c��~Ώ�*C:�?ڙ�{X��Lܠ��yo��@T����fn&!'���[�l�?�}6��.0׬l��f�� [�؋Wj��v�����CA
����N����ܓ�sB5�2�؊��d �۳�#w9&����M�n�J�;�W"��$7tW��Bj��ڱȴЖ�����Ȉ�5�b�f��q*�ˬ��u$��"�5J*�qteKTAO�N��%����1N�O����K�L̡�:��	�4���a�3_����C?�
?j�_bz��2�v�8����n*����ɧ19m�t:ͲfU]E5�/�D���k��8*�"����h� �*���+����Io�h��[f1c��̉^P�6��	 r�&y����d	u��Й�ț�mmz���#��?�N|J��U"\"�ː!<T�7.��!)���A��!�YN�+��yakx`�Ζ/��T\P2�E�#�mP��)�@��%��)��6����ŗ�����͘� �jEz^��}/V�N$����Wx/�3-Kup�}��C��/a	�����|L��v�IL�D�~��i�>�p����)5�(���mm�����C�W���[�m����� k�D� ��}9DE���=p�����s'�������	$�Y�d��L?�o���u��y:�E3jD�f�{��|�vp?�Ɋ�K�R�B�.י%z����@�ߛ��wK�Bx������4��1Z�͑k�#�ӆ^�����0PH���J�Ȥm�u5���l]k��a���e$On,'5�,�O�Nդ��g2�V�%~�q���Uj�]��1�@E�޼����!%��<`H2+b���5�Y�1S!yu�xm��i��8�/ ��$�ʭ3��v�J�0�y=��P�z�]j!� �:����פm�bn�Ӛ��rЫթQ��.���b�Kb�$d�?`�ƞL0��^��'�No�4<�Ơ��D��B���C�Z�/�9�I��̿PԀ��Q?���;k,A@�@:D9���๒H�w�	�wǡ�J����n�~¨)���/<�0�w�N �&Q���r��h/7O�v���zQ���Ah<�UTTKƙ����Yj�9��_���+�(D����`dz�u���:�{�Ʌfxe�u��5`�B�%$�Q�����I���󔲪ɞa�YgRF�<ө���Pp� �s5BN�.9K�@�<׶���j*RM�����M�0ԓ:���>v�R����A	�mn�0�V��js���M��w�1�i�_J}0^�$��)X?���fT����+V9�s��N���t�g�{l~uG|�?���3�|Ҥ�o����sF��Z�����1$^:��μ��|�t|��N����g�eڤg�Tj;����0{P8	�[���E,	i>�ԑ�a=tA�w����K����-o��n�>�v���0=��y�ZA�F�c���*�V��5���n?ԝo�¾�k�^�+s����5�z*?Ҙ��N���8G�&?�g��f�\��Ҩ��2����Xp�?1�#nΤ�����h�x�"idࠣK��mn�;Es�d
'=���|"������׬� <'-H��7,�b�tw.WB�b' }҇S�LUR�K3�:�-]���6�\��H<i��X�@�����i�nZM���&`�f���E��5d8�3��D�7��H$����W�z�_3���u�	tX �f��_?\�Ke�st�Z�]H�'��I�*i�-���;��9e[��ջ�@�D,C7�߾�He1_^���ڭ�����	#u�&ڰױ���y>�9�?{��L ���J=H�#/#/V�r/�(�3�e��2���퇡���Dia�L����~WGqQ�Y��֪�I�|G��;_	g��B�JX�/�s	?�;��G+�4��4��^����?��C��'K����H����H�&I��M�v�� �F�Ca�h@3�t��h�4/b��8������O��� ���6�er�$.�+*F��Hy����[x:4z_+*)T� ZY�F��tx�N��V}���g��Ӽ~�br���v��t+�S2T�Ϩ�ܥ��Ԩ[�x8�ux!�Ue>[>M�K�� 6���jֿ*��r"�(�p�.k:�� ����*X�۵u� �٘]�}5G��:=<Ș�ν�]���.�����n�F�jrk^�i�������柃W c8��W��]�^.�4���� �F*�j�����Ѵ�Ca� �b���ģ*�u����� \laffЭI��h ���O4��=7�f[�J���پs��{'k�3�E�E�Ks���΢���2�e�,�3~'�ٮo{�.8i���4�����K� �.-��֋>>��~`gW�eqv�� TM�B������^�M�g��H�L���p@Y��Sk<UE���qք�8������I��S� ��1��X�W����u��EC��R�7����nA�d�d��J�2�t�VU���YπDӇ�]"F8���i:�]Q��v��s���������d�:L�4m��5rB�m��ٓ/����'����H���xz@�i�u'�ƣnw�gO�� 8]묬�冿Gۉ���,s��O�
���9>l��ˣ���,J�s���8\�����܈?���B�۶�����)�r
*�r��,��=|*ۿ�r��&��H�嶌�3 z�c}�j��4QM���f�C�l[��g��<Z����d���+��>A�F�%ݼ'�0�^ƕ����\��nau+jk}K��mx�Kn¯�5���1��,bYc�v{CnXL2�sk5�Ű���7�r�A�j��9~�9u��ВTM��o���èn�i^->��gI&���-�=�!$�7���;F
!��KCD�X����$X��j-����7�q:�$�5�$u���x�G��ۛ���-�,y	D����F���Is���@���(̄���V�
��OUF]h�'�.H�Pe+����Ɲ��,���;S��>xi� o����y�Z���"�|��S� ��7~F�����i:G>з��X�W�	}nߋ]�9�Z�~�4�����@P�79�����r<UWcd��c*b�Rb�<aU]������p�Pj��T���م��[ê�n�/��Q�RR�����¢.(��c=��v@(���7���R��LZ�β�3�Y"!�R����3! ��pq\���3�zSTN��&Bh��ɳAj�\���k�vC�9���3�Pd>^g��k��7GQ��[���R�o����+;�3|��Ĵ�b�tw[{=,���WX�����^h�Cp�ey/k�ם��&�8�A�ks�BZsO�55U&�f�/���� 0F�[k�'�j(�<��A�K̡oވw|���yJi��,��-�6w�qN:�����ٴ<r��U=�] eۯ@e'��Pn�� bhqx"���.�&�.���7���=�Ͳ��e]c��b��\M(�Ħpry�ga�ZL+i#F}�"O2Y��{�t%ɓ��OK[�oN��ٯ���
�����JJi�uOICvCv�2����G�F7�
�ժ�3���;�TBb�����~94��q��(�_���
�Eg�@���<~4|�?�FD݀��&J�Sk�ʁ7�T�b�fm��N������� _/X-!6���pwm %��KA�Q3�f�+|�������#W��*g.�6��X��CP3��*��G�d4�R�{#��<}f�C��a�3FO\�R��m@�sPL�hO���Վ�}�z�i�=R���2\�{�̎`��Y�����
��í�(y�}C�!P� £H=j-.ش��O�}dW!��t!�{]2��-`O���a�fv6+W޾���U���آ]��M)�ŻdzI�d�r�.��r�����v�W�)գ������+' +M:����Pk���Ӵ%�ķ�ޟ�o�>_�f������HF`�>�F�=Y�TKؿD��?���(��P�O⪧+!N6_�d�&����a�S�
Vͯ<���3]��x�0��$0o�Z@�������p��&{�+��7�$Ƌ����d2ڳ'�xQN�{�����"�x��(�o�~�~I
�����E����;�������u&��ZE���Et�	�%��B,�c���HW8�:ƣ��K��s�H����N[H�S��ʦ!���J�w�l��!����PS�5����� ���P7 ����s�k!B�@귂W���� �s7�J$��6C�n���"}����>���������ok��M�?�SU�1+	��j�ʻ�Υ6t�A���uy��F�5I'�e9;����*A�`d��ǻԔ�>��>	��^yY[o�&��#ӝ�
���]�0B}�v��M�X����X��-(D�����Ny�|x�ԁ�����-XZP��-�Ԛ��~��tI��h���46�n�f7�@W`�M��	�j��gx�a:��U!��<��KT���
���GG���� +Y)u֘*�W[��3�h/�P3��~p�;by�΅��67v�T$��n��z)�aHA�y�d��ʥ��{�,&��^g���rw�Ɨ��~�ys��H~��FΨst��ti<��pl	>�~Kz���dcu����$޷��~j�(�����L>�8	E���u�UǉI��ɰ'c���p�9�>��=���6�񴴴�T�f#�V���j�!��fъ�P��j�e��Ţ����*�&�lU�	̅���ȳ��b�@'�	O�׾�����WlS��.p�b^�>�,ز���t�����	�y'F �����=���wװ�1�D �*'r��$��4�@��"��s���,�֘Dv�	���8|cV%���O��&�$�~�9�hP>ސ�J���v���ۤ+�UNc!e�� YwU�����zOs_Uѣt`�W�-E;�ٴ��o��y�;�J�j�9�z���B/��b�s�P�;ƙ��(��8����$6��}0��h�d���U`����uL3�N�Ii�-F#�\���;�8 ����XGtZ�B�P�`���48ИUV	n�埴<�L(:�-��.�b��I����e@���*��&��d�=/V$�g&����� ���JB1=�;t0"�afHG�=bԀ���A�f~�l�5��K��������K9eg8Q*��|�Ǆ#��	��������GB��t�F�P��AOS�++ɻ�Dc����M
�U��{������R���'[��j�#Q�\�*���Ћ2�X�Ga[9,��&��I��D]��Ѳ)mW��f�K�9��*b�%�M����]���x���<kNB�â��Ӛ�����=J���}(L�J�2�=4�K� !3�����"�ڞ4�����hxb�3�F�^.��#O֗����5/]�}�_ז͞�P�?�L8�[�K��4זA<O�**|���WGp&@L�G�A}%�]�U-[�R�ԧ�ÿ#1-�eǶw;��%�AB�L3�N0ɉ"	���#�_�K�*`��+3W$߀�O@(�t�d��O�N��8��`[��C����J���C��1����B'�?�ŷ�x�{�_[ƤUUnBS�Up�R҆��VEڷ�+h�YkE�2�6�̷�&�`���YFH;�KQ���`�Gr��R����c��:na�עYc�?�6X��Ĺ��p���=��R�I,��^*��Sٚ��:��/�B�ި<��v*�bE�&G�"�o�D6����	8��Ȋ��絣�q9��|���r�?�=������mķ�5�&Z&p�6���{��5�^�������3����^]�D��qz�$��P������ȩ�b�|?�lJc!p=cF]�R�D"�WSV����M������?1�A�K��S�����y~K��\��E,�Gڵ��ʑr�G�^m��]�%�g9����� �S�\���ϥAhk`�#�牴�e�L�z��=�,s���G�_ ��L���'_���wMa@��D��������|>4��'[�_Ԭ��h�#ؿ(j���ZΩ{�!���Cؿ*��ji�9J�{�q����ć���MR!���y��BU�!j�)���R���S�3��*���:��j�
�+ps��1���Ɦ��= a�/��_Z`J��1c�-s���(4�O���K���jAw0ɢ��ё[�Ś�W.�_{��KC�.oZg��	�R�f��'��Q�$ަeVX����e>ֽ�u=�N�Hq!��'���߁T|VOc[�B����
��[��m�����o���d!}��|?AH?�1h-�B`�D�BK{聱"�HTh0K����v�_b�Y��KIޔ4�y|���w�;����[��6 �2�W���=tA:�s���0���f~FIP�!r�f�����=T	ڐ�t�{�1�
�5,���
�1��7 ��+AF;���l�<X�73���R؉Mꌯ�E"�U�%��&��v'^37:������n����@�NZ��~�܎���վ?x�����t���Є���3����;"���r�,P�{��\�%�u�~*��&��6䆗��h.��י0���x.���(_�8Zl�s�,��,*�j�%h͓˘�"�`t�3�Qcѱ�Muʍzf��0���ВyTo�ʾ[�H��Ny�#+���4�;����ld1��7)����A� ��Ք�Ob(|�<�����r6ƑWt$�Sf�����Ti+�[|<��G�p�0맵�W���2K�<��+yW�ĵi�ళ(�[=KR�Ka�ԗ��Gzv�½3®]2u�\@�n!S�Jzn����>R5���Rh6�s]��m�|G8�Z&���M�<"f~���6�Y�E"F�JT�߀2�*漤��>��8>n��w���_��~/��;m��G�#ޒs�2����$�'搨�.�����Q�#�pc
�!��`�M�#π,��LVܙ/�Q�m�t����(�q�=�ѫ�-*��Λ�~��oH5�cs��0�~���B�i�+�*���SX��d��*б�^�;)V�5�| ��ς�V*?�����j)����9%�������j���-B4����̨�lh6?G''���Ws+2TKj��RX�a���j�M��!�bI��߾�Jo@(vlE[����ŏ�8]A(c���r_�\��w�_ʊ�f���|���_���-*�ڭk��`o՝wtZ�ś�[�3}��q~�V ���9�����Y�Eô��R����GCXI�G���΋^��-ڦ���k�eF�0}�w_,�pew�G�����2�(�#��������9?_Nي��g�y�K�M�I���R��ԝ��_�Aj��'��-���zM��
��	���#����2�uj.�+�>Q{o�zU�uٽ;zx�OT@����rs�b,7���2���X�>�M�ϑ��7�0.��"_>Sg�w9�Hi�RJ߱�GIe�9>�pqd��T����v�_�!�̾�)o*-��C����>��mc� Ua�L��o��ۖ�V0N�쁐�
�'��pc_��ߴ%w?ReU�D4߂�vq�Ed�}��Y�_�M�|B����|eAe�Ai8Jp�R��~&��)6#��1��������3��$0�ꏳN�1>h�N���>N�h&�<�����!t����׃˭=��_�],q?3f���j���Z#ur�����O^w���J��9bu� �������{�����B+�L��ǵ��%u�#\9���B3����$�)�"2��(^��4��m�P$(�MȊP��!>���j�OJ�}�Wp�E��^w4�*����|��Nz�M?p�ϴ:��u-�R��b��<|gЖ���+�ʽ�a.48�(q�`�����I=�}�P]j=k,��*��Do-ô�g��]���k�H慪�l�Qk�h�\��1� ց��+ijø��Dk�|-�b�ZOa�B���$�G
��%��n�~�-��ȉ��V�*��� �/�8/�I�"�.��ɘ�i�/�2�p�0��S�̑�����A�,�R�����~�����=fOn�������������Q�iYL��2��Vё�P�_�z�{Ud�;z�'�0�"`�c�Q.�&,� ��:�:����ȗ잘�Q�P���E/���Pmj�T����	��\�t̰�&3����")�5	FH������.\P@�N�&ÐYؓ�O�ƄPe� �bo:���6 `�(emֺ�j��U��?ɀ�=���P�0�x~���U��`\�®(�^��th^W7��	�0��,�<_�������|����^cؓ�&�Y����<T��
V��n�tU�V��8=4Q�·o1	�u��,I��S+�yjSU+���Yq�=0��P�a����A�|�]�ϭ��ĵjd�Ӈ�����`�tIץ�A��k�����6���9��]-mԷm��%��-�@��S�nXZ��]�ﮯ�^�B�e�10�8�'ݸ`��8�*Wg�X�� mn�5���Ƀ����T)�����P3e�^:kJ3�ʹ���>��^��p��S�5h��6�����F3��ؾd�z �:��ԉ =wne�����gMK ��H��L/���6�?����
�2��R��׬�-��ȹ�#4(k��sM�5@��� $=�&r�<�Ѷ�]�\�m���~��e=i�H�B�C5)�s��zB�a�=VH��%�B"v,���AM��95[�@�_
98�lXT����F�J�*�}�f	���$*�a�IKKH!�+u<�ɹL�կ�IK�Y�7� �����e/��_E�^�
a�!��)?dAHIp��k����� �v��7�6[�*h2�#!�W]������؞���C��b�^p����]��Z�!.��()MgFu�k��.'�u޿P��{ֹ�q/�C��_�u�~�Q^�ur:->��aj?+K��=�,_����T1`xzK��䧈2���Y.�Ϝ��Wp*aQ��	Ǆ����M�d��3Lͫ*o$����F�W�D�ٮ�`gW�,��&f�;�9�I���v�jB_E�D+k�8����"4��G�bTNٽ����1����� ���f�`;����v�U_E!�23��2��:�}�!�A��<�@�1���}�pՇs���*?�z�^�/VD��J���dLW�(�W��m.��Q�L��������ʩɭ��K6�,NAQ�`�����Qn��v���p܅W�v����NjB��:��T�c!�y�fI����|μ�H���D�^��~l�$K�ۚޢ�v�l�T:'�
FB������,1$��Ɓ}����b_�V1�;+������S*�TL����m�0��CM��o5�[6j�ˎ�Dp,�	֖�z&��ۂ�y�7�P�p~G��������h�����Z�u�Ǫ�l�B=Vhi���ᬖI)�Zhi��hkm�\�.2�� бF��oj�Z���۶��o�-:�h<X\���Qi<8=�br�0s�e���a��I����pȿ�F&1���B [��_dD�1��N.�,zM�(��%.��;ǒ���	�8�	y]�l�G~OAH3�\E�<�H�_�yFb���Ro���l@�N�:�j��r�]U�j�څ��M�i��&���	����V�h�%+(���$��������!���5�(S��E@Z+
>]��H�XP�yd��	
�0	!��ZI|'V΄��I&~y��Ɣ��^Ą<Gmoz:�
��
���3R�n������pI-�j:��׃7�#�>)���Z�%�@P��T�� 4Z~2�p��_Kf׍x3����D��o�����O��m�ǣ���e���l���E�[G�Vβ������m{%�<o$=(KF���؁o;���^�����W�᧟۫��ʭ�GuL�{�u;}��S��M��b~��:�\�Bl���-����Y,"�1̠pd�����?�p"�0FF�S7��* �C(�:�#�@n���D�J�-޷��["�ޫ`��|�y>2�l�AŌ�ڌ�Q|����e����\��;���XJ���-�AV'O�u��q�_ @S�T�5��y@Av�Q6�%���s� ~�m5�P��ٜ$��[�5�9ʏ�,���%����Ӫ7U`�a��s_|�8�'oC�>�ő���C'������2��Ł�3[�=%2���H�C��M>[�XH�A,ކ�9 J��
g}xwod���|��-��s�\Vrw���촳k��/�8�ZJ�C�mR݁G��z6�'���r��� 9l`��q��0SP��i��%p]iPr�ئ��[��ܮ��T �h�H��wI9����\�y�����6��s����	9���261�Uc�� �D����w���A�N{<���:�IC�/-á��N^A�|���㉾l�#"�������h
�Y�#��D����x1�����7�x�_���᳟���6��������WAik���a���2�b9��l�ww6԰��a����u �x�4�Zg�T�.�k ����O5�+	�D�푘�1]=���}�r��`8s8�I���:�\@����JU��s /��ҍB�U+��^ԁ*f@X�?���]�G~uS
���������V������?w�:��Y���F\$Vs��T��	C�Ab��iN����>�6�:9�%#oʭ�wџɁy��j�U����BEU3�e�\��4@�J���Ūc<� �X)�1�"��������7RH�m�����F�i:BB���u	D�>�c�S=`�
�a�*�6��.����i�|�1��W���E<�y��/�D$�#
�F�.tO�̸٘8�0V��}3��.!�v�a�������,�j$�7ex����쪌�^��H�����P��A�*g�8����Y���[$p���1zgc��rat|�'ہ�s��t���'��#��?�/(g�7_��
�������c�;��� ����Q�$	Ҝt]f	G��,y�!8��.�C��'��V�1��g���	{�~Ɉ�i+�t!v	����ԡ�,��#�ѐQ!��i�-��q�J5�P��j���_gߌ��� -ݼ�_�JӛW�5`)VFbh��B������E�WC�~f�f�5��7���4�������K�ۨ�	�Ond^�����O�#}��"�����c��>�۔�B}j��=�|7zm:�vE�^O�L�*3K�9�<'t�t��-]��<��<�a]�Ҭ"�e>�O���iH���x��lU��o�L�J;�'W�'�7�g�V�Քt��NE)�b�-���U��SG���~�c6�l�ĴV��w	����hm�87=aQg�g�g�uæ)��!խ�p�Ͷ�v��R������V��y�`W:�X�x/��M� �1��q2�@ǜ��~���7����'�uE��k�xN"���������C���MT1Z���$�G�BKP��������Ē�q$�ޅ��g�zN����U��6lz�?5������3��u0���(KrF�i('�
\�rt���*����>QڇMO��x��!�Y��/0��b���a��?��Pi��|@?j=���Z��֥VJ>}�����w�LӅ 6q���ED�x��:sJ1��������葧�C�x���^������O�������~X&.�����eB"�4(	;llr��Kf��ԅJެ*�n��%�:��h�I_X�0}��4Q�B�	��&2���ug��=y�5VMP�"d:�6�1H 8SC���;51��,��~�)/U[��1K#>	����8[W+�)͂u���x�¶viQ�;<.�Ӏq��RJ~�vEḨ���[�>y&EǢ��ǿsX���g��!*g� ѐ^^魥�Ͼ@7��g�2C_���rvU��S#<��Po'�S�D�N"z�n�-�dr���AdJ$Ư�B?���%Y-44Ͽ1���J���s�9��]n cs��2U��М�z��v���ث�*��]�� �kL�q�t?42W���|hWN�HKns/�o��I�g�����L�:�*�X�cH�}��}�Tt��	-d������#�6�n������E��V�ˎkU*o@��Ko^�zQ�L�m|I}d��C��_j򗦏Q��q]���������#3��p����3qeA��%('h_������k�Y�`>��\�sҍ�@���_�Ti\j���Z�k�Y�O���= L/ǆ鍫s��P`��p��4�Ub�봇������>��U|����(�$X�0y!���ˣ���{��� �f#���v!�LJ��ź�Ϛ���I���WC@Ժ���=���ݛTB6nӤ˂����Q甠"�{A+ܕ��"�|�D^�P0��o�U�ܳ�Ѽ�S�=��#���(:Cl,8V��%-��=�]��&�)��呂���ƴlڏ�pa�¶m��c�I��ҹ����2q9�r��(y�N�|T�C�*�c���X�-FܒM@.?P�%���]�C����"��
��N�V_���1�0���n�R'��sQF���X����.�L���u<_{c�����rrg�ڈ��:��0���l�܄�	B���!{�Ѻ�Q��8[@L�y�%!�!�z���C�VB��Pzp���u^a8��O>��_U���n��C�d9'��T!�<��L���&��0`S��Bhv��\��:�>ҕ��ٶ.�P;���X��(�_e�
�o�c졆�%��꼫x�y�Zj�U���0-k�&b3: ���	�+�� 	 kZ���+�CX �S0�M�;���QA��F@��4�@T�ޞ����|�����Pe\��� ���(���sx[\}>�ΦCt�;d��lZ/y�o���	6�r-u,�g/�$�}S�u7����^�|m�.�[��u��Ж�!er[uù�����Ĳ2�$'�f�#��mz}L�����ľ�Þ4��p�_�-�Y�
V�8uV��������p>�]�!���ឱ���H���6���Q	DWb��[�|�l�X��O�\ў$i�X<�l_ܲ��	�D����D�u�H͞�a���n\��kMځ����	x�Xhk!�E.��ӻ�c��4��צ<�_�D�EN�Ļ�.�q)�d��i�Y�A�+��l7���A�尭�x����l���fЀ�P������Ȥ�- �H��0�;tj�8�	���i�-k)ՆG��|zWc�t$�k-W'1����׾��*R息�c�Q���f�!�|�L
��I�֦�C󶘒�r�p<�N���s�!�EQFUߟ��t|�kTŐG�J!0Hn�r򴘸��>�-�v���� ��a0���d\�pI<���|-�#��i�^��p�EP��FHB���3k�Og�K�gTG���/�X�p�\�g���T�l�O��"5�j�Zf�J�Q���)`����Qp]��jr�Z�l.൙ FXT6��1��o�������Ϫ����������G�r�o�rzMn��Ks��Zْ���4:X�����Z��F��TU&I����3�Ow#�*<�`dT{IE�$*|���A��xN'��[��%�=#oR��^�ZCu�4�B��VG_��� �9.��7������d��J�$����Щ�����w�F�g#�6��3R4�`���=/;a[������Z9	ReYX��^��^��1����������N��H�h�R|��lvvK?4��0�20���*����"�D��%���[:�`�|s5��:|5�F�O��Sq5[����x#3]� ��G��Ol���y�~�`�[�s��#]�(��z�`��@:�i�ey����=���z�"��\�kh��� ��y�aݸ��*w��q��3��|��s�%'��nr�8�wK�p[뿨���D�Ӧ�l/g����Wf�*P���%�<�D�Ia�ds|UC!ԫ�}��`߽�\�łEe�d�P�^��4�	>�G�&��+>�N�1��}Ҷ�ʵ��7�e�9��Z)�ќ�e�c�-� ��O?��3��S N�r�����'��H�.'�����%�i?(Q�a��?��:���\B�|6��;o�����pL���b��tJo�4Ls�g��f��bW�ɶ�g�A�0<��>;"-	NH<Ll{�I]毽��S1���5���������	��L�ҭ[3�tO�賳����cP��@Ю����5�2w4لt�0�����O�z�*w���奚��|m[��/P!ˑ�����H�e_��3a`dː
�R0���k�u&�@��4n���I!,�&Tl2V8R
�Q/���j�_��	i+����Q9��I@a8&�&�hй�~|VtS�[�*���Le�O�º=� �p�8F5��
Tֳ�>�n��ۢ�s�_��֔�<sXQ�~CԞ?]��u_9��"m7��i�3Ly�Tڊ��T7r>n5�a��,Ai*J0x!�:F�S�t�\�Pc����M`:$������QX]�G�)s��;l(ѕ�O����N�j��ߓP~�G=B��j����>#��d�����B���}���K�J@~���F�H:v�!����;�wXtV۰0.��vQ >��Ëj��sV6�q��86	�lf���C�P7���?�%�3�/(�r�is��B���^N��'������)�2�,l���+GyU���͇�8\{V�<��,@V+�?4D��~��=�)�����N�QtȻ8����O5�hZS���ݏ��MV5���&T���E���W
㙐�r ߼m|��P4�cr����C;�F4�eY�h*�Đ�+�&P
&Jx���_J�-Lam�oB�wwv�M�R^I�iM�?,ժ���� �*x�X@!p�kC,T]��HnC9�����2��*�.%P�K�4~�?���x�Tt�+X��/*�.9�6��U�K���+G1��>�i֜��uj �@ٿ��֥�.��ݟ
����]aWN�X���ry�AO|4V�6vk�����܏l�O�⩾ω�ͩ������e�Yw�@��n|>�=��UEa�;��bK�C�e�	:y�&���Hw1tC�>�n2Ѱx��D!cw���V\-#����η�������h��93��p����߉�x��s�����Ud�੩p?fNǛ�n"�?҈��#��ה߫�������O���s����8���\ғO�6���lr��B2�A��kL�[��#����<��4�Ĺ����懟���8��"�e�����-��	�����XD629:H���4)L�b�I����]o�8k�M�O��M%��/ўr4e�:=��Jwla+����{��N9�*i�Ʀ*�
Nْ�[�A�!Y��h�[pq���P��ޥ�i�n�\��	��e�Z6K]��)B�V�^F@�� ����z��4�UFr?�&��2i�u��~�~%���w���Ŝ\*N��z�o`��@�����D"[.�si^ m\�x�=GG�x���E1�מ��x�;饍�4�� ��]u�SӝaX���}D`"��S���Wj�$�.�m�"�Kt���=����l���m�?�.%寤b?���w\�h���n:M�$ÑI�w���ܪ|^:���m!aeP�d����T-���5��!��q(��n�m�])����ز���bC���iǇ�ŷ�EZ�`�v��M'M}<FB�;^��dAsෘ�+������y簨�ʡxg��>C�J1�����Г8�yg�o�Z�?�*?������u'l�o3$'^�12�H�ةs<o�,��ҍ_-�=�W���#��$4�.�'b��ѭtc��4X�!A��e��5��H�$�������
���0,<��nf470�A4�t�L?MYC�0��'~���o��Q?������JZ^���=���k���$�"`�6�1H9�6�e����1M"ͼ�ܰv��v��C�5����ל]<�����آ׺��ε�8V��s��?u'�E��F ƃ�9�"��F?��{	4r��2��|d��O���j��_���"*6k�s<ź���wr�!���MB��]�S�oL�]3PĲD*PAݗqB��&�f�B��n�[bE�D��Q��-�؂q'caѶK���6�"�v_���x�ǅ5�m�*J�7z\�hA��N	���Ɲ�b�`p�xa�w�F;U�x�����L>ݐv�[���<��X�S*�~s~|ވ������E������<���^6GԚ���>5��� f�6ؼEBx��w�!Y�qyd����f&z�e�\,W�pֹ�;�p}��*��A�Md�� �9Qp�"���DO�W.)�u�!�G�B�H
�X˞�`�;�,��v 9���U���#3��~���	=����H��z��ۅ��dQ�@&�렙u��Ҧ13��<x�T|UN4�M��KT�SBLŁU+�p�p5���b����T߃��+9�u@�B�lc�e"�\Q��L�X�Ӿ�7O^][3�;����<�7��YS?�*y>�@�s���$�Z��"^�j���j�$z��ڂ׵���>��a���ZS�.�-F&�����Al#}"��A����X}C��:��U���ɶ��;����JI�Q�#�J�v��E����rw8��T>��aC�΋�:`�X�uN�Q  xׂ�~����ڊ	��x 
%,P|�}܏7�VI�$�?=0���H��9I��{��e��޷�^�#$4�J��)��&��7��,�w���%�SK�>��{�'�z_�ק7��n�y��Grysߣ�:H��Ń#/��t���3hm�M�bt;P7gVVD>~ژ�r|�a�Ƌ������R�T�,��~�0p�W��fRn��8���M�aV�{jV�q��H\0�Zt�/l5�S��a��,��=��ھ<�
�ui�,�g�b �W3j�`c�+� �`7��FH��q��Ұb�
�u�G��]#N}�	F怷z�"P�,8O�,��$�av3逩�f�$7S4�5��(z�J��Y�J�� ��1�i�����刯��)��\��H�IEN9���@R�V!ih�{�E��a!z����^�����"��Bn�ͳ|wP�.\��4���'e��ۏ՗@q��%n�)m�O��,�txV�J����*�u�"a��=���ӏ����/��_,.��i��k��<�io�dS��Dw׷��$�0��/���E� f��[����U��B��0�ƨ^��� =������[���O��-9叡N�'���K�����,�����-�Fҳ������������,�!����y��4�n��@�=�r��n�x���\�d��c���"=^���.�ڲB��X��T-0��w�%[JNәc�"��0k�aG�[%�����)�Y����7�Ç�%� �K�����q�e�bd&�iR���[_���t�d4��LJ��s���Пt|QCG�����6Z�T�r��D<�[���h�ʕ�8u�h2�d�!$rq,3QZM��J64�P(����t~8G����&�)5�Ws�r�׸:�:N���TNM
��{@�����95�!Li}tVb,��1����L� f��_�?�j�e+G�D4xv��]�:Rk18����<���nd�I4y5:�˱��q݄"��_'^���+m�7h=FĀ@X�;z�$�@�6�n���M�M�dmʕk"�;�����	�Y���I�'�t7�+ܣ�B���l�+Hّ��+���,���ZC+�;,����/�Z�������v:d���q'�M�s�J��-9??�E�i89W�e��G�qN���������Zx�!O��E�K-)�80�n�7!U����[݂e{��E��A�˲-���O���A�3Y�H^�(�T�S���LK�D�hR+
�"��kg^.��9�Vo���pX\�P)�o�-e��z�x.b���|KJO4�6�p�Ͽ�#�p�\[D��B��$��P`do����V�J��5!���������r�,�z :�C��eH�,��e�,��{w��ȟ���xms1����8��͋����v��o�RUw���$qFJF�yٽ"g����z(�ߨ]�A��9����<���i{C�����+�H-��`�Nѳ�i�}D{�qa�ʄ����v��q&���-ě6�aB3c���n��G)(�XܸӘ��)>���<����u�×�V����	����V8@�4�BC�样e��-R(�.��A������Sh�jj�ʠ�L��B��4���B��|T��W���X8ZY^�!�B����}�mJ���Zdaވ�1�����޴��8��0�p���l(P�1�da�Iu� �\������SB@����	��ـ�}m|&�(���@%�S���h��Zh�7-���@�-Bu��S�2]l5I�d>ާz[$y���+�N����m��B]��z@,"����\��)��lJ3U�(�TP��3ܦU����Q�M�TZ��=B�TzH9i<��PǪ��:FtJ!2�+A��һ_8�"P4��x���T��oq�~XWmi/Z���:V��*@�6�h�J}a]p��G�(�Л�f����F;��ܠ�W<�ۉr-khMh��Fc5ƹE��9��|o��r�'��1�f�k��[�u�^� �j�6� ��5�˾����|���]*�{y�/T�\����26���e��g�~�q*�l!ZO��*��n�%��%$�LW���&H�f����)kNTD�%|mTߊp�}��;o� �<��]/���}�[p��������pp��V�M꾲�3D��w�i�:�&��+�&���ߏi�{�ȗ�R���a�R�=�ic�Bz�PC�����z�'޵^c�%гy~2�~�h ]Z�B���8���u2�b�=���*��;��2����r�ʖ�2媨��þ����Â��jR<S���*Gc	��F8�!����8�@�θ��p�����������O�j�5��[Q⭌��)r�E�=���b�}�_-` ��
��(h�p@9��u7^@��ʪxd�ǩ[Xt#ջ+�E��<�r�Ep�ɠ/���d�¨����~�C�CI��k|��!C(`�:HK�=V�L�\
����#����ds?Y��
*�i��$��s�d6	���nfG8rO<ņ�k.	��dzF�@��b�cn�%�n��Ԡi�muI4y�l�Y��JJ���F�#�Is�A�JC����/�o	1�C�q�9�c{���J���[E��g���_4+z�6����;��)NK��T)j��}���ō5@ !�25/N�yu&2{>Y�-m{���� b�$�4����*��(k������\r��X��Z��N�:̡�l�l����|��!�o0d༯(�ӿ��	+�G}�E)a�!��|����>���Dy�`mo��D�xT���܏�98`,+����YU�7����� ��Ee��������� ~u���S<rc%�IBL4Jb[������oGT�ms.���~v���\@0{̻1��X�'��c؅�b��P�פ��f��b-�>a���E��75�����+���We<z(ت���ņ��}틔��N{c3�Ʈ&W���I�b�8l��G�`4 z$��8��.��2{�,�4;«D�t����_���C%p���?��3�LҏF"^}Nb������k#�J��n@�� d��g��YI�4����z�y@���~���)�B{��5v�ۀ+y��Ƴ,�ܠ�����|*I�{Y�>�Z��fz��/���2�'?�r�lQD{�n�"�y �YQz?�V���!�Dj���W�����	��Hm���M�6�gD|97�{��m�s�2vI ���1)���:��I��m���b��B�_�a����r�HJ�TrQ	�(���y3M��s���?�6��K>�3�ٝ�{'�i,*���?vF���W�T�w���&�D�A*�買/�F^_d���X�:�	9u״Z�])��%kӟ�.��.u���/��{=��Z������g��sbz �g���s�Ե�?+�ih�Y�'�m�b���}�D1��u���T�y��cX���4eT��o�5Դ�/"c����)ظ�n@�j�������XQI8ܹD�6��7��ʜ	�m����G#S��Yl!%L���?�E{�c�5<iP�����6��k����y�S*�1Q�$py��M��)hsԟ!w%�BJ�� ���=�mv�R�ra2�.7���t��6%���Wu��}=�Ь���/���쁵���f;,i������c��`B�`�?�%vF5:�!]V����&�'�	m���iA�+��*?p��!����$_��?�i����U� ������/�L�T�^l���(Ea4<*Z�����V���.w(�_������p:��4�V=��%��鉄��p�Z��ʋ�S ����/�T�e��ض�J�j��ȓ��̑���gR����̭nd��Hd'#z<Ό�>LǨYp�J֜�9éu�3;���fT�Q�11HC�C�O$:"�}��:[��ZRz��W��(P��vz���j=����1�x�.�7O#|���}B�w�[X���	o�4�
�[c�Yv)*�/�3��FJA��ӏ�)����*:�%���ԔB��u�\�4xA7�&�Ae١S�a�L���hQ�m�4TS�N�/�%�G<����bbJ6.:S�=,��|<6�7Na+�^�_���)�;-��v�)$!c�5���&˽Y��׏�?���D6Vt�]��ϙ���p���c��t��`!�A��� [vU��Tk[9������o�"d����Xԭ.T(kՎڂ�J7��QN���җ�eh�G���s��Y#_˨�s�`gǤ	6�{+2/ib�{�B�J�?} f��m��j�^��~����W�''����}���S�����Zɰt��y+$������S�{��%7�������=��Rq�J�0�]/�{��\��g4��Ȕ�in(O<O�y[H���>�N>j����� �|2��tArkӶ�,7������x�Y�o��C�r�_�n)�oٗ���}���m���u��FE�j���k+�e~��QF� hO�e����+���OkR*�7���J���'�܃�ͳ8��X�dz~3��oF�Mqf�����:�a]A2ufm�;�^��]MF��A!�Gm� R���T�%y�%�5��9��]HGB���Hz���c'���}:�P����}l�`G��������NT��Ug���Z|����U�ݵ}F�84�����:f��^۩ ��r������s�:N_��<�b��/v���9>���'�ϊ�NR	g:�?�Fz�lF}�l1�p�R(��H�,�'%�*fyZ�<���N���ǝ��4G�j�=��rp@y2A��i �N�'���W������i�>�z��f�ƒ�&���\������8��\�>� �:�������;%Z�@��A�d�P�I�5�x�h62���J�+:z��G����MU�B�$� ���7��� "��M?�VE�K^`J�����*�hv?o����������-�<N�0�E�����wk��_�6�A��±<����W:�%��ؙ��bȂ�]kj��k-���5�8x%z��N��$f]�F���8GG���� Q]Bx��e�m%���:��1�NyOY ٘�f��#�L��S�R2,(�m�W�1m�5�`}G�s#���@Z�ڎtF�=pX ����}��ǟ4��C��!a�Pʋv��ÂOI�|�1��H�&?�Z˘!��̓j��M������h9�g��z�O�J[G��K���
�⏦:]y;L�y��V㨜�dP��]&���U��N@���c�z�#���!V��,�N�V,C�DL��ȑ��\jY�Z+��5n�.r�� �)������Uv��Wڰ��� dAcv�H�i��)�S�{#섟���w�-�v�~�fp'T�U�I���D$i��ŉ)���#�7���n����zN;=��<b�0�X1�-�o���|gu$�u2"�^�玬�a�����,������2�r09X�������AM-��g����I*/�(E�%l�vZ� k�����Pߖ5��8i��A,�n;81��6⟎�,~���������#��Nal[KS��� J�Z팡�ʑ�r��������տ����w�t�g�G-\��YKFjz.w&���4,|-�`(��f���>���zv��O8���}>�-�S�"͝��x�I�{�@��S�
{��s�s4zR�c�2�s��B�����O;:�%�>�G���r�QJ�G�<�sV�,�����M�"Ҡk{��]U�@R3-Ӌ.=����q=�
� w:[��D������f'7�����*�w:���_�� ^�D�i��rcb����B���ʦ��%�m}�xP!��������b��6*�X�Ѥ�u��&M�5����=��9��If���#L�:����e�b�@͙~%T���d��`3�К����»04o�h�[��u�2��e6Ü"2���,>%���=���U�YU[�(�6ܱ��K)�>�٭ئT��E�Q� ��{P�䜡`!@���f�[G���:}7�U� Hg"x�@���/�Qw)/�U��F/r��n|3�Ա�ܮ� ����p����-�����L6P+�[u`z����[qu9T!
����C�]Zlp��&Sח�7�/��U�ubH�����ˑ8�1,u���n� �����䫈��Zk�O�%��r��S���g��=?2����J��8\v8�F[��f�6l��J֒Sz��0_�v�B�������O$�!(��W�1��5���}��ý�¢������d�b��XΘb ��jj��繚l�h48h{� ��Otf�Ǯ�Ep��� ��L�J:��Έu @�CA#_���N-*����k�x�KҤ��v�6{0GW�\�v��4�A�N<w#���>�N��7��Q��+�r���]S�9L^�_���3�t�uD�C�K���;o�+S5b@�mĔ*$XQ��0U�����b_��㑤��9nu�1� ���f��M53@O*�
ٓEg�Ķ�QƢl* Z.4?4ht�~X������ r
���w�U<_C�Ҫ��kJ�cǅ��1�	H{��kV�
4���Q�8��.z��� *��i��r=����/0u��{ޗdj�ņAh�H�o�U���P����9��A-RE�;�A�������m��mu�*g=P��w�<�,R�����T����l]R-��쩅�*��"��qw��	@P�ֿ"Tl{�ͦ64X�C����1�;6=�I��ͅãg�đm��`@��=Im�R����].�a噯Y�"����uU�=���.<f&��n3a��<h�H	$!�����r�%�ʅ�4@o�(w�T|�w ~s�NO��P��M5L��XL�(�#|�s�|�Q[�`9���[v{����R�R���7�dm��� �_;�f0C���O��?�?;�5x��Z��;���'������(	?k��0@��,�o����Y��:�>P>T�������g���};�M�:eW�h�B�T;bD��`C-M걩"�&����,���=L�ɏ\��ɷ5+5,I	��c�#LАz��)�&���C ��M�t��{�?��;�W]d�����U^1����R�YG������´[~�N
`���%֯�T˛����-��BQۚ��6�|w���e0ԁ������L^^�r�z?��xՖ��d=En«��R��xMZ/����o5����#֣oI���>��u��2P�+�Q�����i��u���
qK��(=�ӈ#�g��p@�*���URl2�pLrnX��^8Q���|��R��2�jK۝��	j�isu�.:Ҽ�=N�d}��U��b�K���v����lo)�� ��M2�W[��u�B��Ϗ����i��m�1O��
*�5 ��K6�����? tro���O�
�[_(=�t��N�s��B���V��̓X� Y�}T:�5��:=�LR���wBܪ��d�dơ�w�\k`�����z��*	��[��Qc��v���G	�m��A^����z��4�t��I�������(H�'pk��s�uhBR�+8�
�y@J��J�|)��<�8�������sj����L��@ܗ��N���Cx��;�u�ۣr�y�y�>˩K�{x!�c���1!v�a}~ߗ�B��Ɠ�����C=���@Y������آ�;g8~�����5F����n���+�FzoX8_��>���"�(�@�z6x*
�]<>.v���Tmw��6��B���)G� ��S}���?EPf�� >Q1ׯoX)L6qpf��tI�!uzW0��Z�����z(�j��-���Vv�+�^]�W��!J�t�K���eh�i׶�KV�3ũwǖ�G~�9��ję^�0�p�
c�cq�W=�":�V���"UH<��]2U���B�W�r{�^?����O�M�`0!���z�R��'+u�"��c'���ϡa#4�	}]��F��f3�\���כ�x�9Y� ���5&9��!�6��E��y���k��$<���U�>�n��+����b'3�{����~�܉,A���엁rm�o��5۬Z �,2�����/VI���1B:\�3�"��D]�:��d�n����S\/M2����P�"|(A��ּS��nt&I�d��D��!��}%�1��bfu���G��g�H�# �%�nOg�\�6Gc�9���Gr��FRm'İe�u�A�F� w���FPG�VVt�<�[�f���{d��k�;���l���Ӓ�
����A|B�IkcdSH=���h����=��g\}� �'�C�$<������4
�,u���oY=	oA��ʖ�4M�g	��g��QcX�	�8BМ�[��)D0��)>�����6� L:?#Q������)Bg?��81	ٜ�G�(����TKOU9Ett���4��#�7�X�@��h�I
�|4���^4�#�҃g�Un��	
������,��ʛ�_�:X Ĵg�X]�:1tv�:� �D��	�0iA^�o�sB����� � T���;�C�o�۸-�(W�<��E�L2̘�?��lrS��r��I��)~�� �{���ףV�������8Z�D��(��!��ai2��|z���;:��0°bs�����z��:�y�Ӊ!iȤ��7�i�Z��Q���@�nG�b�t��Ѫ��C��IK���r��Ųe�|se�l��2��9�@��4|�&�{'����s�}���E�Hǝ)�t��陕;�q%�e�4���z���Y��j���:�F��K���lGO�)ݡ4I��+��$�I2d�&�(�'g�ѳ%��"�YY��2��b��F��[i����/ł���Lě��ɞ��Q�!�mxũ�[�$[Rb��0�t�XBҝǖ	�� ��� Q2����^#���O��ۃp�g
�t�F�N��d*�@���,Y�UY�^M_�5�p��U��Wq�zcE��u�� Ve/�^�����gp���O���-r��W,�;ӖϬ�O.'3���G�����E�9*�b���r����2��i���{P�e�F'X����Z��~���3� q�R-�s(���TO'�sڷ�'� |��w�+�È<%7��b~f
+=[c�ﻰ(�ߌ�3RYVm�qи�V ��xɘ��u>���d:��a���
���fG����{UV� W��|u�����Xd �Z=��1�S�]C<A'����߻��)�J�e\u67]`[f.�@	��N�b/�/-V�ʽ�ha��(�ix�D�#-{Q����-�lTa����ec ���ZeA���̟:B
����qΦ�Cʆ����γc}�9Z��r�������'�!2�&qv?�},lQ���>�	�uJ���X�Y-e�2Ee���jx]͎��M���K4�� '����O?�'��L~�G�`?�C�$`][e2��ZCᅬ�u����2�QZ��_�W]���/���]�N���R�)�+�RgOE��s�Ҷ|�^$�9���UC�z�E�|��4�K���e85��4���q?l���!���qV׵Bn@�d$'���4{���4��Ğ�u�}a#Փh�St2�p?N����@�/���)e.]o�#�iBeÉu����YV���c�h�c���`�J�O��Ub�ǿFb�8dJ��&����f�t���*�؏��ؚq���u-&��]�@�����`�f��̉F}��4n]ħ3��o���6��8ߍKF�=�8 o��Df^
sF1]��GM�e�o!Q
Эw��G9Q N�6�Q�T�;�|��ŘƄ����yu�;�3����r�J&�;�xM���f��b��^6kr��W��ᙿ�r��53kx�uA*k��<င��'���Q��%M��<������z���)%�q�꟪��)��� �t��GF=up��s��y��4�p`�y���C�:Wz1�"0��<B�p�Nݥ��4j�k�)z�����xq��Yױ�y�z�'�� ��Y����'���3���X!~�'�p��0�:��lc�&�X6���·�:D.��r[]	��Un"g��m�rV+�}2�|��Jih���aI����*�)���wf���a����g,� �o�����V����)%�-�Ɩ�����sa�,�=�u�N�c�y��:�*�%��;6_z��(������or$�I�q�\.\�Z,I���22<y��]�姽G�zU�����=lj[|��J�ڿ�Ci�_���%�ʒ��k:�r��ʹ�W��� E�D�,$���=�~��}8���Rٵ��g�!j81>-�I|p�]%iY�ˏ'��3�i>�r�}N3��R�}P�?�����^�\j���5):��)A.�ֳ����a-���18O�#�e0;Z^�X���vh�_�W��䯽��YFf�Y�Pw���<�H�]�,Z+۟P\Q؃���b�V��,SG��̔�73\��h�C�Z7Q�sb���Y�?�jW�u* �d�9�3}%E2"���}�<nR	n�%��e]���VM�1��̄��a�L|������FV��K%5[˩�
W�e���AV��X��q5�U���p�T�1�3t�nO�Z�>G�FMZJӲ�&X����I	wj1�L����\>h����hkAdǛ}�
=oWgu/�>D��Z@$���X�gq�^���W��I4��|S?�ɂzO	)O�y���^g�y4�����`՝�"�X�d��!y�i2XD�a�s�Y�p6��"��\��+�+�}W6(	⮮)-�<>?yo�$����%���˧�5���vy�-���Ul9w,����aq&'J�\��˸��V��y�<[ ű���P4��K�U�p7�A�j�7R��6���Dn�EF�KH����ne�H��¶�c�`�q�B�5@�r!TQ�d�DR� 6Vϒ�ۀ�uZ9��ܑK Ӛ���B�b)�y����v�MhŎuO��S�Sa�'���HωB2��sV�	��S�aPO����w-���"��1�aZ��E�/�q�첄���ӗ>[�+Bt<�-�/ߺ`�������<T/�$H���}xh��L��'�1��@/��8� ֿu����Ȓ�m* Lދ�(Ӹ��-��Ý(�%=P���q.k-yW�{N�~{�)>�q��ѱ�v.�琢\+���e�����Э�T�ެ�,���Ѱ���j�(e���lf+�n���`x��#���e�D"���j�0���]�i;�Q�Z�:��M��9u��z]��M�57z>�v�|]�_��'Z�����'���ޤMM�!�=�a�vV<N�,�wG�-/��G�R�V��"Ś`\�Ȓ�U(���������8c�\�\�'��v�_�'�����Rz6�B���WI(�|D�n!:����t�ξc���a�oz9�/�_�h������-j,W{`���������h|'�O��E�"f��*�p`�b������M�4���ihf��$�U�mX�2B�7��=@8|���8��\�%�L�_�]�.���3�s��Tܡ�q�*�z���� c>�;If(�8��B�]$�t�߯-ha�bLͥ	��cJ�W4\.]�����g�߆4-?�Д���hO���YfխS��B�
I�Ύ�t:4�Hk��;l��t��N���&@����C��޺q��Bm�Q��_/��6[���ć���zE���ݿ�1!h�D���(4w6~m�v���w�ʳW�;�Ġ�]�޾5����.��>�ҽ7�XL6��,}�t��F���e�dL��˨%co�����=`A��������!���8�)����yzߧ�zj�L�I�M��=�1A�* �� KY����S�X�]����q%��Z�3�ZDl�WV����hr(�*\����4j�L�?2�o`	�i�4�`	:u*\�KKVxhm��#����x�y-<�������m�?��Q�c��Z�8r1��N���%x�����{B�+�`>ٜl tSuA}�>����K��=��W8ف�?��Q����>��wy���L��#��QԴJ8��П�����7v�f����5�a���PX����F�U��.#�'��5��yd�3���`B+�j:pO��nR�Ofܰ/�z��f�+ab������\���HB13X��.:�`�����ޞǧ�$ߘ�O�"Q^��e��w &2�HK���$����[��f\@��;�p!9p{�O����	i����2	l�|t�6�^�ƭ_ͱ��?��]`��撃���53�܌��#R�J��J��z�V��O$'}����ǋ���f��\��$�c�߃ň�� ���*?8�@֥-�C�ج�2�d� .]	��n�L�Uvňx\�v��\���K�S��0v�_�O���G,��g������l�ҩ��~�nk�S��ܗ��H_\�(��Q.�Qo��S����������������Ƽӹ��*��a4+�B�F�u~���-FQ��2U�]=�K��TA�%Thz;K
�Y�8����K�tL�l;:����z�~��e�L�z6 Rx��5�:Z_��;V�$�I�����Ǹ*: ?�/����ȳ��"��g�U�G�j�\����&��1M�9vnD���=� C�q�.�Q��i���i�v���U*��F5��^Q?��=�{g><��Z��7��_�����-��t���O��6�ƵS��8U�%$ȡŉY-p��HVj����<��%���B���x���.j�E�iD
�e��ZQ���l��'(�Δ
$���*�uW��b����,��o��m���u��1�J�x�XiB#�2tg8�O��;WfR�)�a;bԋt	�Ȑ|�5�Ӫ:��������Īq	8\t�����{�!	�Xնɮ�y��l+�[��3
nL��<���>�H�=���ɹA�4];U������0��e^�|�_豈c����~n���v�v�>Y�҇�]ҋ/;Mٛ��ʹ~����|��9����1����~VqUG��ȭ�/���zyubz���b�0G�Z��؄Q�O�ؙ�D@���=uՠ��H�ZJ����v�PJ4��Y��N9ա���$lM���`����;j�k���/���|u�$ƹ-��~U����&�n�6�(#PW�"���g�w���7��mi�z`R���!U�C��ݥ������k����҃��K�/"7�_��7&�aCǒ�/cBJ('�䢖��5��F�~���F��p'z��&�:h������M���V۬^z�6-������?}z��g��	��XK��z]#���ﬄ���R`��<^�.o�-�H����!F:��n�_�^	�!�>��V-&Fb�$~����-&��|����W��P_[BX���e::2/���ߤn����=��2v`{+>bh*Fy�����V����1�f��P�`y-�b9V5���o���i��1�	���k�SDqr�B V���A�!4b!�_�a�R�=�}�'|w��í*�oK�j;�	�w �'�= !���������=�|z�=�g�zMç�@	�(��xM7�7��$�>�)����E	�PU
��^Bc��j�5<1�`�������!bI�)���VC�D�l!���������O����^$qU��g��2(	�C��X7K)~d)�`G3=O����7b�Q��㔡���7�1�f��
	�Oڨ��Ұs���s`�܌H�z������<".�4S�٥|B8�R$�<�q͋��i�Ў�r��87mӝ5P^�
�~�n��#?��V���*��]�:�_fc���F��I�b)!{��8�>e����(Z��"�QM�����̛�}-�:n�5�LKW8�e&U�2*�i%�v8�y�WWm_㡘�;u�Bg>�{�;ӌ��l�1�J�F ёh�;-����h� &H����%����v-D��9�G�v��D�`Xa q�v���U�	/��F�i=��JE�=	u�"e�����}x_�xq�yk(
x�����7}��7|�2�{B�i=�|D�Y��9�;G�����)e�Kz�]xӻ�?�x�=�)4�`T�ՖD>�q\3�W���"����u	�0��Z*��m��X)�f��|�A):6+���!�b��h��D�T�g��f��3\C5B��=�Z��ؔi�x�I�@� .j�xUh��ђ�5'@���!�����æ�<"���e7��lP���$�1x��{Y��( �#��귤�*�M�}��œ5���%u6��#�g�g��<7\T���8x>�ѥ�>��r��� ��j��:{����"�9�SH�&z������6$�/�D p\)�dH�(B��j��)�A����YA\4-k{1`~!��P~y�Fh�>��վ���o-���E=,
� �IZ�N2enj.�!�;J�6�V�&������A�� �U���A.#���1r��"�10��dR@��.
͌��|�>�F�^�V]1
P.eM	<�p�|�]�<�B�?:X�zs�{xlU��o�r��hX�u�M\e6~�F�̶!o��,�� �5l��˖#�3X������(.:�6Vc-*J;q��o���"A*����"$P7���l���|8�=�у�=����i=I�$a�����?ȧD�^ΞB4�:e���9OD/ߝaR� �>gZ��!l�0�,'~ ����v�k�.V��LKߴ����1���8�D��� XZ����0��R<�I��B�\�?�p��ǅ�G�T�U���`*���-��	���4�)
/_ �ft��U�j���H{�/�"�ܡ�Yڃ!��Bx�c�aF*#;�M�`��'�p��$ǽo]�*^N�Z�w��*����y��09�z/��T��1�(UCPfW�x�z���ʘ$z:Z�*r͹��������L�>Q0?h�u��{�����Cx���5_���n����V���c�� J��� ;o�`#*����j���T�B�9�}��b���6)|k�_�W�"���4۳ԯ�z�~y�0�0):��e+`�RǴ��n��N�pd��	}�R��)H����@����SP���'�~��mX�C�,����|Jđ�pq�&��T�F�D��^}�Z�)�*�Sf�\� ����f@̍s2U����=�S��`x0��?oJ����M@�/�U����l(c6�u���~7?C�������&ڀ��^��.�Z��V�o5�ى��-���;����}X\HӮ�$�]n��f��ƈ�x�� 6OKc�'���G�9L]�:��/Oꦰ}S�u%tnT!����6���3��;��t�f��r�ψ8�q�A�n[�8i��׻���#$�L�O�.US>/˩QW����{ ��pЌ���'� �9� };+�{ �7�߿�<o����w���wq#T�
�^!�P��qx6�8>3��I�S���FؾeE����NF���3'�x��;B�@$W r$�|Q�����5�C���;�D���Ü�fPn���Q��?͢10 zcy$N����o�u�����=+�B�߷u�Aw��� zll�=���|��Cp�P�~��n"ɲŤ4g�sC��X8r��T���-1�U_��$zNT߹��m�<O�L��O'	�.Xd�Rp|axr"S�c�wi���b��(�s��F��Å�����{�R<�6Q��yc8�?ז�
x�o��F����Rr���d����R�M�X�h��C<�G�5���ơ2�u�~`���õ��S�{o\Փ�cr�`7���{�-���t�?C��{U�^ŷLo'�*�٤`ߎ[�`��n���VZ��sgf�g�^�7%=���K�S~�H_�4�W)�Ȟq��𪍆��*֋�|��!�/<]����Z9�)�ry���-�L��~)���NSZ��"���`�����Z�M�zq��,�S�a���`��ŽuZ�*�F����Z���o-}}?����؀��!�
E�n<�9����R�)P,�b����פ�>-2��٨|_֔1��jt�fj����y��N�YG�4�>�)��l%܅�C�A����5NV�ٳ��MN{��|�R��7ӊ|�%���TЧf�73�Fr7o�*b�}
ʑ:���rf�5 4T����
���ggQ߅&��J�s��чH�r��Wj�0୊/&'�ޕr�v~`���Å!5����إWêB��:�QǾ^�
TNЬ6�H3��"I��f���{���� |��[A���9C=���I����&ʁs�MĞ"�r��P,�ΐ�Ѯ%���nv�Ť�|a��I�S:��E*�sS*:��ӈ$�B��⛯q�Ƹ������ʶZ��ˏj2l�7%g��qT���7Hr��W�M��BO-<�c?B���������)�tJ����m;I_{��4�`5��_`ZNu��r�����X�#��2���0H��W~�;u��R�����-�P;�iB<E�&27�Z�V9.�xH�H���a���Cnʡ���ʘe=t���6¯!�*s��=��(R�G��x#oTw�x���LGJ���4$���bR� �[?�#���?ː�GE{&F��A����k�YqJ�
sI'�T"f�|t(x�M!b�ζ��*�����B���\L�u����� PU�iA�M�����%4Qd�S�ː5�������ӊRw�L�Z�^�e�aq%�=��*N���R�4���s������~��P���Ƹj�:��t8F5j^a��͗��% S�~o�T�u���dŅ�;[Z�F4�gˊ�+���2��a�"��N;]y�?����;�� ��4k�G�#ϳKtun#G���2��٫�#)�2po�f"y�xz��$�Һ����@��^���(&7X�n�v&�	����a���S��x��g竾�JѪ>?��>��<�X�6":F����(�+iM���%��K��0�p�6 4�����|�}���h}^�*&S�����D"Z�q��K�A���$6eQ��b�oc�*6g�	�/q�}|Dag��Qq�}���E�`�
���O�x`���	� [��X[��۰(B^��S8��Gx�]���*���%�.�N"�#A���rvI~�.���Y�3��9Fהr�qoLFRj歂��'
�@����[y���&<���B7X8N9Ĭ�/��3�T�yr):l�H]���d��0�n?��yi=��Ż�-��YATnb���U�u,�+u�YO����G-�=���J�W=���fa�p1DN#W����d�䔏zm4�����qCL>'_V2Yp�4���Ӊ��1��~�ZX˫��>L�*E� b�����Հ�vt��v�
z{v�-�	�����|LoT>FJ����Zk��r�}u���>;4�3�m9)�C�	IΎ��<�e����h�Z�2�N5i �Z~�cUx�&�s�U��؟�un�3�&�X�5^��p	>��@c���������`z�0����Y^���(:�y���_#�5�J�w�F���7���9Z��f�3�o����%�`j��쯤k5w�� ƽM��4�Wv�@)E!?��O��Y۽����`��v�lT�q�G�fa���m����9QNa��ކ���HE�4}|tW&U| �j -��<.aܼ-?�LW�r�Hǚx4Ϸ�JW�P����5�d���**�U8۷4^=/�0��x�!\������dILK�*�9��Ӌa`?�o={�珻�X($g�� ?�8wǐ�F��I*����H�C���\	�.;#^1��T�dO3�ODpR�FVqu�h����N�uW��Nb��b�z�R���
�h�M�����)e
����7�4>W�Z�i�d���x�\B�f�衊�d1S�%�N@4P]�-C<��'
$���{G�>�օ�Hp�8�,u�r�R��K���o(e;� ��2� bI�BG�hZ��AYn�OC̯�j���Zm[���YZخG�论cjci�'�]��AD��X>��>�7C�8D�A��˷� �B�->tj��7�[�Ⴠ���o�1�i��܅�$�බĮ���۠ME��sw=�w����}>��!y��b�o�/���gc.6R3���~%'��H2E���o�<6�i��'U����9�~W�.�j���+�!D���VPDI-^'��VT�L�`X�0Y�`��fX6�ևu�x�ӱ��_��B�QA��=�1���6PzOH#͢��o�&�?�H=l��!G�z���	f,��,j��{o���mR��zdr��
|Ot3���)E����z!&�l$��d�0>f�@�;Ma*��I!��f��[es���s��R�P��Cw5�=kS�aoѤ����������j��5�.|�Ʈ�~oտ��6 ĥ�@_��+�~@�~�l���6����' z�4�dB��"*����n�!�i��Km�ܽPd�ŷ����hț�4Bc�_�BW��es8A4/m�_d/_��Ы���%���>k��fABʿ�z��#�%c���q�!�:.�J-�����L���a���Pw���+��n�:��l��"��C<�����$6�AmYG�X�r�5,$���l&Q�&T��襡������*]�ԝ���{l��tcNѳ}��3���>W��R���,d,��|ʎ���s�і��i4��P����f��e_0�@	�duW��D��1��=4��������3�,e�����:xΘ,���ao^���s�!x�΍���i|k���\�2�>���,����UͬH|��N����;�8��w?>Y-�2�O�  �=��&��{�؛��o/%\8�-Y|�?,�տ�/BĄz�I�<^(��ij�>N	��^R<�uM��-��?�54ŀ�I FՈ�(C��W���e����_H9��Xȭ�K0��.6���.9Ls�e��/�̀I���U9j~��R׹yķc��ﭡ{��#�!|y�(�"�/A�3Gxl�m>R�v������v�#�x�l/�k�r�N!z���E
�� L(��Z�J�*7o-� ;�`����� �:�\�K�LE�fŸ������~��}���_�d��#��z�
MX�>Z��`9�8���I�A�`⦥*'&�{WoHpp��?21UN!b"o��XZ�_��4�2J��!���-MA�+�k����x�$l�d���l�����_�1~������*�|Awv���x��&���2�xKQ9�m��m��4m�2���k)����r�$3K$�C�Ӏ�>��gۋX��.�@��.C՘��C�@�T�
��j*���V� ���M9�za9�'��d �>D�I
x��3�e�&�`�\!�1����v�+�����#��7����W��c�>}�U~sax�����2(��cwmf}l|��G{8$vE^���_��!�qE��I��U'~B�	$������ �n��FX}�O�q�E,�\�ruX
{�´Q�h�hMխ��$'wM��\��+/U�9��:kө�\AB���U��5���4^㍪����峈 ��7_���a�Ը&�d2e���9�;~.�ر���Sln��"4�i� ����.ڞiS�Z��lU�7>�Q&�4U,�X��	�H��̐M>q1���@4����a@�I�!��i�dce�E���l<�x�$���=�o�r�i�	�_ih�FQI4��Eu�V;#���U��P��P���U�ڙ�������+���5&K6Z�`��uG@f���j�i*,�����XFJ�e�*N��k�B
�����B�Me�?�Tޭ$y����X����Z�8=I]A�V�p��W�v��H��~��B�'���<�ds������H�̙�m��s}_�4�t�]W�Z��H�t=�D��߂��YA������m������)k6�A��Ǆ�[���6�j�����w��'k#��e�:B_"�r�;��PF��U=<�ı=T��h�52��_m�EQސ�=N��`�Nz�V,<���$����ʧO�$JL�k�,�}Y�P��Q��aE�]���u���Z�H秐�[ށt�D.)^$�9��2��LI��);kJQ�t�4��;g�È�[!q 7���u]�Y�45�_���`�@jy����^&�Ga��iUZ�*D�*�e�Rp�W!���ͪe�$3z���C�����n��8��wS4�h�E.h�7"�Y2M�sgE�R�D��{*�܎�z�W�*@�jٗl �;�I�h.O����&�)i!)���t�fЉ� �x �UD�Ԁ�$^֛Kz��$�d�@9��/�.d���n��s>���Ѕ)��f#r!;�C���prv��dR��̃�8Wr�6X�\���H����w�Ŗ�"��p^}���&>��Ζ���K*�c89���[��n]v�%p�p�=C<d��w��P1���8��h)��q'��gW���lB��_qo���d���%�D�ȥ�� "f�3 ( �\��r&)�N���5ඤ�5G_�z���65`���d�:?{�|�����`��	��W����v���D�i�r�]�&��	���_(wm'�3އ��U%�`x�u�W�,uU����փ�I�?��DFߔy��p���{j:4�j܏Z|f��B��P76��}�q"�<$ܫ(���ބ��~�ۼP�|���)�Ũ�I-��4��LU�J)4��-Xع?`.�d�ua`	��O��W�9^7�d-�`��-x�e�����#b�~a�z^�^��"��H/�6�m`�\��3�R���t\�X[�$H��>(6�Tԫr���Ȁ:�_�h�I��[`%
�n�����`�䟏7�V;<Lg�����P��P��k_P��)�ہ\�،�i�5ԹuU��ģ#<���W��l�o�(�VQ���!���8�fа�4�|6�Exu$9&��	�{4��VD=LҘ���m��{$�����)�
��C�@���.;��4�|�C,jU�K��	D�ͳ��]���ux3��1���`��������0����� <���N���iK�-Bˮ�sɂ�B�Q��5�B����{�kb4!���p��6j������!3�.^��6���8�����>�����
v@+�c��a1�S;xbV�g�?5k
s�`bx����EO��Q0����AD�W��|,�Z�uoZ.�_�Qwh���� e�}+���!߳]9=�e�6�q�L��qs��Y�B�f �-j� ��lh��9`DɣԾa��N�z= J�Z�Z������a|#j�^EX�� �@N3}�@�� ���?�� �d�qv4O7P��:_2�X-R���A��}���?�j�D�z��� j��}�y�X�M����b85$e#^5y���D9Y_xU������!.&�E��LiJ�m2�//S��:z�~�#���N�UB'�Gb�Ȑ�^ ЈH�����yH�d�*0n�V�0��3����Vэ��IS���E�	��ߌ��X�r��~	ܴ�Ev���3/"N���{�9ǳ��>ĝ˻�v���%�J�����.)����J����x�t�,$MgV�̞ԍ�j��]9÷�?�|M���~h�"�z��Ur5��éCƃ�AHɵ�,�z]t�z0�@�!ϐ;����m?�2�km�����.S��
������s=��K��'Rv�~��Rs��'j���+�9���Z �Ǩ{A4�P�lY.����r4�6Ӳl b����s�����I�����*��������*{X�C��JS�k&�yg��+3w�#ɤ����/�l�n2�M�of�ϋ!Yx�@h�ܼ���"$qp�(�r�U�^w�L��Ƚ ��d4bZ�1
��=�Q�ڥ�bl/Y#I�*�F�J��r�����c��7Z
HDz��3JĖ����[���Ƃ�3^WinI�1���}�_-ra�K�T�ڢ�q�g��Jf�Gbzk����;%�|o�H��q�����h	���E-^����� ^ٷ�]
�<TXD�� �5a>���V�~��ɾ��k�U�?ZG�1Vuv}�l08R�l�<�|~��4��O���'�~��q
�� �[�a�rV�O^e�֎�!�1@��e�H�%��zS^��-%PsLDJ�����Ĝ'ӻ�MLA�m���1����C&�Y�yS�|?�x����L�g��$WC��ߵ�x%_�Z�)���~�E�h�6�r#�+Z=zjw#���y�fW��ր]_ӱ/C츅�s_��\�6��d�91�;����&�i��NV��m -a+w���*�iM�O]O��2��k�Е1MJ䆧p�qvw�x$�8w-��M�Ӽۦ��<�g�V�5_�>���P��VT��T9��JK�RQ�/�2��{4����gh�n�s�8I���v���^�@C��o�j�@W���`,�U����7"��$ɖ��竅%�?���Ց}�R
�7��\� [C-��ލD$(�gk�2�:� ��'�y�UW~-��l��ƚ�4�N� � �av!�����:]��	U%��)A(��]��z�
��i�.t��<sǁ�ѳ^d+C,�pݐ7E�#�������kh"���k����#�q�ҷ�^߲]���+�t9>�ˍD{��b����~9��4o��j-K��~Qr'�C�vV�y��ü[���G`Θ�.��/�r��/W���u���Lo �I�jv���SIvPG�(6�4�=M��B��양��}v�1k/ˉK�1�*v8<�d��]�<�����<gO�9{��"�ñ�q蔻`�Y��֪x%j`��ذ`�.U�j!D��yt�S;����1 ��z۾-cP}����[�ڎ��[�y�A�B;�fISh�͌b�$��C�b)Z<7m�Ʀ�����xwc�ۇ<Ç*޿�u�Ø��&&������F��S�WL	`�8�����#�H�k���#�|5�3IgZB̅�JJ�b��8�Ekt����s\`oRaʲ�s[�Rx�~��;,m��NwW�a�c�����3-
qpT^C���;�i��l�QH�z���ٰ=�����@�hEM��� cbɈ,�o,����E3�טZ~��vf�V�C�����/��	��n��M�N`M�DLG7�d�u�9�-�>Q��T��qP����U�{|>ps�.Tm�1m��F�}�&�e+�)�I��,�_�/��k�����,3��5xS�%�$�_V�I#�F�dj���\h���C�[��$�b=̕�1{�����ݍ*�VTH���J�d['�*I6�a�����w�#�H��I謋@��aS�}K�i��v�`.���r�+>���;�Π# ߾H�my�sF��<>��2&��'��!�.�ĕId1�Ynҏb�Ck��0{���3�ghIW����6��M+2�{�}�Q%Ybn��h�[3��E3�E��j_s�b�_��ݭ=+I��y\h:�Db�TU��t���[���s�Z���K�Ae�;�vR��Z>��$�V�� ��d���م�.�����U`^1�Z�*�ʗ��"���������eq�?�H�h����*�5�C�{�Ja?��f��%�^���G(<߻�p-�O�E�r;�*|f�:�����0����=�]�.x����O� �+�rg�����8���l<t���?G�x�i�у;�S�1rɧ�o������
a�p6�H��#�ҀV���{��6ayU�[%�s��nVM���x0�:�l��r
m����&��5���O�ӎ1K͓�Ty��J�w1A�U�(*Ъ�^t�nU�n�v��������M}��øl���¹t���E�"�D&�j�p���U�i�f-��|�w�D�`��o8���<��5'�"	B�ŵ��M�%�OѴS!��^/h"Y>�+X�]e���M��'��5W)4���Dn�6�4ף(�KJٶs�(��V�fU�>����2��./�ij��u,3<�mM!v��Wj!>���#8�
������r4bD�ƹ���4тDL��`���/�6 �Ky^G�1΋���Eh@�e.�,��1�A�Y����N�d�m����d_�z�a���ę�P��vy&W�[R���?���~g��^O9n)�K[o>�7Á��m��*�y���ˣ�@�;�_���??�y��������Ϗ���aK�fԨ�P��f��͛���f8:��Ν��KVLHE
��c��Qq��H!j=|��=�s�6$�����R�(�:Eפ�N��*Qǩ�lqn/:Y�Lsg2���x�$���X���x��(

7媓 �I�_�T��4�׵9�������~��u"�/����F��/z�Ri"Z?>���[�W���[�#�����ĥI�ˠk��7�����_����5��"\�\{���BY0XN�Z���3{��NV9�=�N��z�{�ݬe![`�W��r<��69�o�(�Q�����5��`vX8D�Im��y?E=wfd� q�l8P�����r[�����W��E��y�ޏccSu1�Ə�=������盧��^�&ҥ���܅9h�!����'B�6 ��X̮M��[�D�ٲ�x8!}{�x��`sS-R̎�vق��>��h�o�g)a��n\{3c�g- �qO�{$�+�cz���#
��ͅ��{q��[0��ّ�Z��>�|"��M�o���YNGYvU����g$7�,U����&h:K;���+��B5�?�ӊ�aDn4�:��TJ��U|h:�EG�Y�ː|<l)��Ҥa�R����D4E��B+���Դ6�ApB{�I�HP�ߩU7��?/5�c�~�a���LJ %��Tj=�zMA�)��?!�S����ou�ֳ'��6���~��Jr�u��K����!#$��`�yd0(m/$)D��Q���R��h��D2M6�NP>���mV�Zh�&6�sh�R����X�v%�(WOy�29��&�F+A�/n��w���F�i����9���;�Ud�#�Y�i�I������a9��.�u~�
1'�3��}Ui.� �7�m�WpWks��-ȡ�ځ���'^�ռ��?�`�{�R��̚m�x	�� �I�B@���oo���[�rS��y6'0���pض�PS~y)�@�9oB^������9�}^�o�`ᦿ|B&�ĶJA��:q�:??�m����'��@mb�(��D *����B�@Rb�/N��F@��E�>/��4���#��y�L\ �K��V���j��#=�NBj��K�2mdp��Gor��b���~����F.)Ko���k!���U_'���ڸ	�k�PN�6�a^�)�$�V�w�� �I�=
�6��B��u�(�'R�<vS��e\~&,�3=���6Zu��Ә+T��\���כh="RG�	�(+,"ɩ����?�t����WH�,{�w�Lu��^fW�](����i#���	ůH�|d��>|?	|����(+�u������gpoKrYʚ����V@A�WE)�ٿs�
9h��)8&$h�1ALD1.���^�`������`� �����:�IX�R��ר�0�������&P��TOO�5��DN%��ҵpj�7ԕ�\�q�*QCz?����ut�
�l�}����@����e�ϨZQ���S��U��+bq�|�o�{L0���H͑F�=r����g~Gh��\~XQ�w������������{���F��6�v�Թ�^$�xjd�+_f���xp��F`A��Q�'���s��w�(\��S�Et�Y�rѿn+��zn*@�d)�/ w��8skO�H�l���HM��4��S�m쓵ܻ�>�)��?�Q���� r�.�{>Ɏ9h�$dI!��������J��t���57��mFB�ھaӫc.x"�n��}1ŀ\�<0��bq�	bV��S#j�5�`�Х�8bx����%����pAc.B]m�pa�Wu��Y��p����̔v^� V�6�r�L<�(�m��Ib�>8dے �[�Ɍ�q�p���6��hb��Y�k��t'���X񷴂*By)+GC�vˏXVİa��m����lc,�s�TvQ��i�cj���O���b��߫�R�G-�?঴A�l�����<��k����4N[�����,�6fvX/��e}Hf�t����(�
����h�+:|�j�;_ۣ���6xDL�lt��J�`$pU=�
�9A(�wR�~�\)OJA�\RR���7��ˏm3�/��n��u�4�Qn�)��)���� .G�BB�_E�g�RƠ,�V� �nK��U���Iwvy`�� )ݱ� ԍ�x/ce<����� D!-=��C����A༕���sV���;Eһ�
�m�TJ�E�;� �� �[K�'�����V`�֓�w
�[�r��"���)'�,�)�N����d��aG�,vi��딱�93�V}_��V"v;���<�x��� ��g�&|*�O�w�}܋�b��|c��G�>�O�େа����{1���E�UH{��J[�����������k�a� �O�����B`��O��6�5V���.����3/BDB�)�_�k�-��8���vR���[���в.x� �た��!��g�澖�$7��Y?Yx4uId�;�v%`n[F]l�uz��u^Ѷ�ۜ9�=LrZߣ8�����Z>!��]�LX��Xފ�@>lK��Ir=�ʛ�9�!Z����������ww�!.~��H�J�7z�Os���>̘EBG$�=���a�eq#�۶�7���O a����l���8L+Z��Z8�_��DB\�k	��mSkO�o�ݡ��~�e��2��-hX��1����F�RZ��t`�Z����_� 5�m�s�|����(��?��;�\u+r��c��p�:�x��g}['vn��B,Gvc�4_u=BA�"�@��6����?M�/�V`�����eU�C ��fJu� ~��N��"�� c��Wy���$~������Bz�6�-r�˦�@����&���~H��
���ۋƋ&"~����V�XJ޲U�>��W�p�֠���-7�b-㏾mcS^,��u�U4���)AG?b<�F�	�iP$�ܩ�>�qm�M��*c��wkS+~�N������1g2��݇�ܯs��^d�h[�\ ʎ-O��+���N sɐ�>}=F%��+��v�0$g�k���/�nu�D���nJŨ�|�e�����Y�<���x8�V���S��)	@����@0��q�k�PҔ�R6�ԋ�/�ʽvl�ؒ	I�i X-��n��қ2�
���RD��e!݉��N�[���
I(l0wm1f$V�7z~r(�:�.��ip.��v]*��\We��}��ݨQɠ=��ح#FE0���[(��Pb�8�ޣ�/v���(~s �$�b�^6ӊ��Yg:�yɒ�,��J~���z��� B>�#�#��ԸЎ"l��)�i`�b͔5����x��=�i�
9Wb���|���֤ p���|x�RnaU����p�\�[�P�R�C��W.�s���V�
��37���i~&a�,��Q}7�0��'_�Pc	#"��D�*'�p���\-u��Kd� w~�w^�c*h{�y���n_j'\�0��+)![�a]h#��N.S�}OH�4�v����]굼�u�t�x50�[Y�\8�P����!�7�a�7�N,���)U�,A{�0��Ψ+>+ �JX�݀���5H��c��bf�[��Ī��T'{2��c5 ���s��X��-P/��Ӵ���$�b,�?��C�dLG���ƕe��,�s����N�s�I�{O�ɝ�Q��a���A	� �����fٔ!�R��{en_��@q����͟c�|�j�c�{���\#L�D}�[r�k�r�����r�6����˿Z;��>3�e/��i���K<�:�ѭhW�r�a���,��K�$���6��sܑ�p�;��o��xquƙ�<4��<�ˑ���k��M�m����?��ڟ=�v]N}��� �l���l���:�S'2�p��`Y

��}�|RX�crE��x)#t��	P��5&�
���Oז`���a8�P>��Zu�c���s�w���L�gEL̿�������3o3����.�j �HC��g:�kp^�W�(���g���K��K�u}
_-ؐX��g����ivD
E.���DJ8�W0�Q1����;��d����x���b�w����}�����]c�x��ﻝJݬ���TCd�+���)P�rB����\n�O"/Xw\8�#�:�s���쟈�&yaf�NZ�}����ψrt�K��c9�U�9��V$���("�o������)B�8c?ؖ'.V��+|ߕ�ԣ����� +1^Q��b���{M9c���=�1��
�Br��uY�*/o1�I7�d5r�L&Z6�U���H�~�~��'���	�Q�O'Ҙ����c@���b`n���ʗ��l�H����[�_�FZ�,����9��^l�}�"�ƣ憋3#����X�%�Յ��}��Ib�g��)נ`�gƔOH�B���p��CW=׊����xa���sW�5�+��&'�dUDaXː9n)��慲�r���%��K��U�t�� ��j2v��؞T�{�T ���L�ۉN_�����Uv3��=������E���6���!�'��Ԭ%�on�� >�X{x��_@������̙�Q(�a�?�v33��ӭ��RJ�ɺ���r�j�%�(o��;���uD���9�x�V%�%j�2#���h���3|���f`�q��c샳�=�ۓt1vS�ݍWi�@�i�Ë;b#�U�B���>��N����E�[���\�y�����>��u��K��R*�L��0'�]�K{�L���8{��R}��g���	cC�@�n��&@%*TO�k�"��"?}�tjg1=�t�c[W�t��Ow:s�7c\(����g鑦)��S8����~.�@H�'F�щ�p�O�hp1�D!���'6�_�r�@�
F�S��D��: $TvS��Ǩ�`����F{e�~f�-����� ���`-��f�
w@��2� H8"rF�k$��H����g��q�<�F�J����"������o����|�GI^p�8���oo�(ݲ�w��f�e�^r�����T�;3����Ҋ�e��4��X�d8��A�&cJ����	e7��6�. e�����2�Յ�r���� �=��P>Uv���"�a1�+C��I�E{��?j���I��$���╝x#��a����c�̣
H, �㰄�j'��:`�	���n��]��\qo�n���F����
���d:���HI�Ǯ�u�[�B�������`�+��ج#)��P��E�ԟv��&K���U�
Er#S�S{a62�]���%��2I	�w͋�9�9�$#0#�͗���y��aj�l4�ɳ�֖Au(m!%�j�O��2m�`�UnO 90�k$d7�xJύ�Ix:(`��QC*�����7  ������hI�]@V#8Oj��ɒe��&\��5��;��#�R ��[Eř���"�eG���(K��d!�	U����bx�\���������-zG�9����܍>/�0Q�)}A1�WX�AN���~�n��6����
��;<K��k%���f����?U��1(�t!� �Y ��a�=b��l�@��)�mt�NCLwB��Aw�]0�a���4�EZ���%�w�B�AC�62OpC�A,�V��7��$|��m�j����|��3E�&^��m�ў�B+�n2�VgP?���;Ԯ!�z�.ݨ��˚��v:���7�ׅmy�)̳.C�����+�Z�H��݅��$aE(���/��a��{���Z�W�[�)ư��7qm���}��z������B�H�(��LP�� b�Ȃ�������yW��8���b�fE/��1���:@)�@��^hh�:��:m�&�n���Il}�x�`�z�4���]r�e��T��s��?���M�:��p)�V��iY�]��H1F"(�%Mҋ4[��Y��R�LWW��|c�8YRڱ�����z�6�C�~A�Ζ`n�(�l��tp����!�l�w��bd\�� ��zhi��I���G(��iW���쟤!��P�0寵-�hh�v�X�L5�c�����?À0a�����<c��T��`p��b��md��KASEy����H�D������7��j-�6�N5���c>'@p�����*��C�?gU�Z��G�f3�A7�F��� �ƅk�`�!�� �Q���]t�+��l�$�͹]�+]J�J$�g#�3�d|�~��ѕ����w�P�vЌ���
'�;��������t>�5���j��ò#�LVkWl�g�>�*x����P0�K0ޙq�@���	�a}s7�I��/J���xшp�O��3�n�~7_7���fMp>����n�/�Y�ܜC.�"�s���}x#�I5�xvc�}׶�
:��l&�����e= #o����H?uM��et�t�k�xi�v�2��!WJ۝L��P�B��5��������?h6ZSH��<$�L���6��,ck�R��]N&�Vx|�2�&�l��"�g_���zx��W�sm��Q�a���G�j��6\�gOS䠑)�f֩�\�I���#�W�ȑ�*�Ĺ�V!���MW.���
��Ċ~���hZw��dĳ3������F%�3pp)JpW/�nV�V6��H�����Bpp?@�����'b=��P�&hJg 1ͩc}�����+�}SΕ<!�oi#�P�˳��TV}�ץ��&'0T���4]��L��0Z�Vmx���+f������^��Ea���w��D�>�-0dHU��T��~@���͛�]?�)��`�ny�S
�e��[ji�l��%P`�]��^GN���̺�}dw5uVN �ȴ["�f"Ukb�O�ÈD7�����|pC�|���J.�?h8ː��H�V�PG�~I�����{K�`��_mt���4��!�}�}�A�n�e�f O�j����)]8�=��Ʒ7�	V��Ӧ-,PG͸D�+ˡpVM*N��Ֆ��y�I��8^������i�`�c�u�z��J�CXl#�㟂~cB2�z҂ ����v,�YK����Y���2������T���_��e�(1x٠�Ky>Ƣf�����3���F�)�,��s9����cY�ǆ�UH;��`J&7��nƮ)�U.O��o&`�=�yA���pR	�-q�U��YCQ>����$7(#�9�N�ꎇ?uu�#@A<���v�@�6+]#끻��`hv��oFO~���������3��s�5�A���I\�!�V!g�	_7 )xdf�f�z7�(����c��5���h"���3p,7I����겱=�[d�����Bv���2nӢ�|���Pc�!q���Zh�u�}�|��̪����	hm��|�c��Z5`|��y��Ɨ^i%�\��d� .ڜ�܂JQ�`���a*����wE$�{yf������ߨ�b��W	�L��E}L
SS�[f���2P���@A�{l�%V~��&߯���{1�K�:�TڎH���9xzBKL��ٛ�S�U��AAX�3�$�s��3�U���� �p싀�C���C����Ep�	����b��⊥�P�G-���	
4r��K�ԛ�jR�=x2{���L��7[�,�A��{�v��oKR���7��N6�ü'��"�W�E��0e��W�?���E�#�e�E`rPq9��RD���b�V�'��xR�&c  �.as ��ҥ�(��)�k��7�A�@k��KgY��	���n��g'�����#5w��E�K��t,o�_��3#����ވ�#-�����T�n��Vؘ<WȰK�����{����̈��w���� �Q|U�������,����	p�����1�/'` ��5/�pf\��`�I��iUj�`�L��A����a�m�xӡ�`sU{��O�:�m���u��V�[Ud�2��G쨩�w��-�N�k�=�C�߉i�א�4O�� ��[G>����G(�riK	$.>4(���(�f�_�1^IΒU��[wR&�ٍQ��\'�^��̉"����B~�g����?�e�.(-���im'�X��5ֽ(Tz)��<��쉑e��ӹ���e�ࠟc����&��I������ɡ�� �]�L�Y�#�&_�=ˌ��]�v���w�%������D\�� ��z�\�r���W�i6���U��)����ͦt�K�h�� �Q?�J
ȗ&��m�ZA��k㚦q0��������dR�Y�|>D�/ی�H+�t��he:�����"ٽ8���NsЧ���
�EM��~��~�T��	Z,�����'�yW��nT'��ӈD�g�A������rќg�,!���@�0��7�12&ʈ�B)�cYdw٫�n��7���e�����K��'�M�(	�-e�ٵ����:_8��BҴ�,v�Zx"a8(��!7�'����x3(wK���r+�����A�+G����c2Ǖ��[��.�� p|���]�Y�8�lӡ��8�^h�#��/I����*}N�lt�#�����R�Is;�Ĳm���b��LgI��l2�)T��j���Z�LE��iCV�/��t��,�BBɉoEQ$K�_���}��D4m��L��_���?ٽ4�i!ֲ�ެy��P�3E�La��	�=nq�M����` u\}m,�4��xT���(=�.^ė�9���|�Ί���}�y�%-�~�0��HF;@Ǧ���dL0��rB���)!� �
�~f��9���w���F]M�e��o4��w�4'�}}N��K|P�Nf�U	 ���^��9d�����A�4}LQ�S���NG�5�RBg���`�p���y�"c�~�@ @D��%S��{�&(���`�)�O=O���tvm��)�H(�9���ʚ�� !��GI� �-Oo�۴��Ҍ�o*"��ΐ��_���v��q�|
Q���&�-~�ܳ.��� ��}����O��Y �¡fs�p-�gpج6u��=�$�4���Q%����W��#k&��K��>S��g� ���3k2��C��=,�}����-��;�$Mr�M�}���#Z�'F��-q�t�ǭ@���F~:�'�Lw�`���95'��R%JyqϾ�4O���z��Ȍ�<A� )�7+�4�e��?��,� =�Z���Hz�d]�F�Y�����5�Ṙ���A�=C��|-/&�Bg,��<J|���R���IZi�WC��1�-+�����/�C��*61��'u�����/���`��z�DP�sO+��wr)��|t�2]�&���Z�ps������K,͘�i3�|LF�8��T�wJx�k|ƈ�E����>/
�,&�g�Vy�E�F��)z�mH��h�#s3l��1����2���z*?�~�/*�����Z�z&_�6y�+'�#?��\�t�{s��7O�ϟs��{q�.'ﱦ�� �
�=H�����7ɹ!��VT	�e�t�B�}=����µC5��ޑ����KY�}��.Y�N��4����b���� �ngL��K����I��7����
&��ܴ�~,N��qlH`a'l�F��<3T�}��Y��̨���z��7�ڞ���.��|ȣӘ-���E,n/�UD�KV�ˑ�N'Y=����(8%ܮ[�S$M+�"���@ƚ�y�rC�N=��r2W
��(�J�,�{�1<�~�y�"����<@����P�o�w�>1��:k8��f���Ml�Ɂa%�"��)P��V�L*ꞑ"]WV3��bҵ��~�I�'��i ����D��rG����Ѩ���@+C�S$��i���oc"o8f��dW<�E� I��$����o�5�.�,��suHBl.�O������SR9e[Ƥ��T�?�A�����t@�߃*%���޷k���T���so��O�)W�5�xK�_R� ����!��Kf:}[ӓ����}�Z�{f{��!��+���٤�JTl��0���݇��̼9��%������g/�~���,���9\�y�"X$q�m��3��&*D��
���f��W��z͎2�R%���4t�Ї���=?���@H�&�����4�3U����o����������L�;�(s�W(�#�����|�SR߳���$�g�4�ǡ���W�}N�Glɣ���X<2���ؙ���΅Q�1�Ļ����I ��]�P��09��pnG����c�<�N�;?�w� cr�Y�ρ~����bbc���'z�����)���V,�E)���r[AQ{&7v�1G�*��sՓ�&����r��ϳ1uWE8�5�O�*������'�bPIe@L3�`o$���9��D��ma��ؙWy�x(����f��Ү�Ą�D�$��n��@#�B�u0�_�.�Ӕ�E��O�xU~�5u��v]��$��M�:�B�-z4�e�4k�۳/MM�T�V�i�,PB�� h��V�$W�zhpm���������SD)�("R��)	��V^��J�~�L*3�&�U��7���]k-�yz{4�#�h�\I��@��ݴ]��.=��A8��Ok=����s��[i�n�՞@<Ib�C���@�Mq6Ƀ�D�����s����2�J)�2��� !ȅ�vu���st[!Q�
v����^ם��
�C*��O��mb�1[>�%_�#q��=�kG*�D�&��"��� ��}���T>�/=��\�W�Nn(�Dw����	�I;L��w��@;�Q�F�r���bǽ��u_���L�]a:6��	�A����z�������YWd�����Anuh7�.��7�C�X���[]x|��5�����˫������x�\�PYc��l���9O�Z ��W�x1�+����C��QcX�HW��0�)���;��3��j/��6��q��3��JW�i���}��h�L�#�#L�n����j�vt�PK	λ�A켄��O��͢MB�?�;���a�Q�[j>$���68�:瑐eqy�["�}�,5˩O�Ag�qdd׆T�⛻t�r�
�	��ˡ"a�M/-s�}P�X���6[ة6���:g4�M�yb��)�·�Gݽ2�1<j�4��iP��{��� ^f�jȒ"��T��jg@oq�n��H싐Pr|L80�>a�c �!��>��P �qUO�[?����W;;a �14�x���U_��_L��TY��a�P>'%�Z�Ya�h|y�A�B�q�w��X�-J�+������Lj�Y�0�V&ɏthm@�-��6���'�$g��d<n9O��n���n#��c��Pb�Í[)�����u_�E����M��H�R8�#:H��߁��f����9C
G.������ �x�ZNB��Haa�><������t`�/m�N��#C��^��L��v�e�iw�$-�Ht��0l�=�����r���=t^�;�D	Q��ԲңfRbd|GTt>����<��z����W��ՆAW��y�".�I�!��2˓D���sZ[�>��d�h{���|�ER]����,x�e�Ш`&�b�9N���\̃	L"�N�~;���R����4�{�4Q���\������9�N&����XLݕR�A����Y|0H��n���Fl�
ǪB��U�Lk5�^���wk,���^\������}]�R��,��n>|.E���3��DҦ̘c}J�fk��B��U�9�p�M�����]r`ĄW��P'۞-}�[�c�Hu�s�@�&`�:rI�ODM5(�n�2��N�3m<ǏAz!�%w?�����	�f�Ѣ���O�ӣ�z� �ܙ�X�*��#�;~{i���k
s��y`'a7���09�W���tb=FV��J�@]�k�PU�*?e�)��������b#r ��7 ��mrb�7��T5/���(Z�]dd�oJ�T��7��-��������?�k��wG�7q��'�-�m�C2����#"`>�f]��ëD�c&M���{�� ��	5�*\z�o�5� od�L���|}��I���u#C�8]3T�0���@Z�G��ޝua��ٻؗb��6��x`�l�"��Q�����x���P�J%��*ƨܨ	a�������	�U�z�U4gz��V�l�������ީ��5��\��'�w��^�]�H@9�����&�qu���m&D��I(xǎ�/D��(���p��Ⱦ�J�BSS�%,��"}I��a@YOI�T���;{�[Zn0��F\B.�	)�QU�Eb��i���[�:��sg+_l�K�4�䥜��;}����}�ᦻk�]�0/
q?�0|:��w �}���ӂ=�[v�( �Ţ`�	���`ôy��pz㏆\3��싚>�Ww�/�:�Y���\�
�0⛭��ݩ�j)�T��)���o����E\PM�7G�3�LC�[�7L�k����,.)nx��N�+�h����3�b�V���CkU0�����R��L?¼���g���MqT�9>�������`(-7xo�!`�o}�o�P�� �K ��$Vsm�l���{�g��k�r�-0\�S����A��*oD$�ik횊�:��B���+(Q�nʟ��]9��a�ڔF'YD
o°���A����id�9�Ub���$=�rrA���	��m�$���B�cP���X��o�["�ˎq蜹_eq_�H�?�:��T�&]�@>ɲ^c�Y�c�D�o�vY�#����l������X�734��@
9^�).1�x��=o��t��6��0�?�,�TFR��_�dFd8<J�s�Ÿp!��r寝]��q;�"�[�~�A�e�M��^�.�B_�#u�:�m:����j�����Û�uP@�>���t}�% �R?^���Z)��l��_t��4��ڸc�ߓC�$��
L~�<j僻3����2����eB
�Rr	�A�nsW��8�oRM���,A`0'��=�#��+#>/f<��D��!>�F����K�3��{F�k�R;�љJ����BU�'�C"]��{�$���7���5��VO9�v��S�3��
,�O�w����sT����t3�����F9>�a���Fv�y<��f6����M]~Sx����Q���Q<q�-�,®Vl��w�E�)>��y�Y�/%s7Uj�(����C6ʠ�����vЂ���Q0(	z6II-OZ�z���	Y�FI�8.�I2���Pѣ7P��N������� x�讧�E���5;qBW��e�nMƖ�4�8��!n��^nƹ�ߨQ���A�8,��.�`?��|�mE��ʣHWt�X�CA���%�꙳��-&��§�[��k/L��;H}a���b�wC�'=�)c���n��`���$�"�l�O�;\�HzPc�.�W�fh�aHC��mK��]�>�m$h����G0����؜��g,K3-�^�}�rC��O;�U����U�`lgƞ���Ub\���_I#
�a4����6�\�ᅉ�æ&q.Xu3>������ދ����ls�ԅiU �E����Y<���8\�s���v��c|�U���l^��(}f���9��T�,��v�+�_�R�j�����ty��9�� �i���^���w�ǢOq�G
9z{S�D�|�J��DQ�C��֪v#�d�/p}�J1tW�n�YSե�v�o��\�]��g��>�Ů.�-���j�	�X�\��p��ũ�?E�)�𶻸ARk���)`�����9��������BZ��qӾ�k��D�����]�
ف�r6���y�˼��V*�٩4��jQa���.��=H�U!IW�D�Y�^ycO��֌!R�p�����w-�R�G[mJܕ*,���4�i�9��Y<�@F�+}�<�{��� �qA�a4������n8��8Ћ��
�l����kP�����s�/u�$_��G<�'���b�?"#1>�vճ���s��S�J����/b7J��rD�	����Β�oX����x�* �N`9��n3�;@bO/�&��2'����)%F�?��mn�\$)�5��3pm�S�k�N:�N�U��üʜаw>n�yU��/<��4��<zP���zKq���PMk$��)�Ͷy�Ne!�A��t-�4������kD�Q���"p�c�b��/�1��/43G���D��w�s�����ok�B{#���ew��&a��@�7G9K�(UD�������U�'�G ����D"���Q��%'�
�,܏bqCzW��#c>t	��2���3��Ր
qʜ&x�� g����sum�?Ф������c�4�ƿ.5�)~c�t|�߬V@g��sq���2S.��Z�/V#*�����%;D'�z��8�3a/�h�ЕU���l���G[�D)'Lڧk��[x�tΈ� b��Ŋ3�,<����z�
ˀc�An��7�2�W)���x��:�>`���Fj�Ԭ�����S�7�ќ�aIc���м�F��i�Q�����ny��Ĳ.pU��
`�`�<�`٪
�����~�]1�,����:"]ˀ&!+8�Z�`�=�)�@0'bO��p�%�����JB���au2�[��XH��F�wߊ�Ǔf]f��T���'w��G/�9��9}pD�����r�5S�s�J�Q��l���ވtv��h��+��y.����У�J6���+����&��1�߹�?�E��7�c���m��"���6Ih�0c�`�i��2��Q�V�~Syߦ���,
W���a�;��+�%��.wQ7>��{����Œ�?�u�慄|�7p���ǳ ������zQ���T;A�Ncg��\#��z^�1��:���/��iM� -]�d� ���k�"�T�ڏ��� �Փ�L���>"j���I�%P��%[̟C���
�t��'�w����z�ST�J��]P�=�M4�ڸ8�;5�]��"��yq����8-���oUV\!+/ff�Z�L[���'���>�7�{� ��γc�o�fҨ���U|1��4@�ǻ��^��.h�����	� )����כ1Q���:�wG�~���.	V�C�ҤY�^�T��,4¬��g��}\d�%T��d�.+��$�X<GE��r���>�Pjs�i��gP:ѣ��K�5>F��`�ׄ�Vg�S���/?�X�'��/=4�z�l�c�\;�ztT@��:��q�)�^�wB7��q,����=���,1=G�7G��Ps<E�����`~�	]��T�x?�A$�S���y�q�_r��0�?�7G��pE1Xg�49��Jcd �9��R�E+�ʴ
�ȈHY�p��F�^�����W,��ZY].b�ڸUDFy�Ƽ����ѵ�P�S-�*a_�q)"A`���&L�R�m[C���0_����ᶦX���Oy���)� �.�^�+�U-P�s��*I��r�����$��������+E�dܱ�����(ftj�V�TXvtbNܝ�����z��5����Ӽ�҂��� ܒ����U���=��\kw��7C�msL��u� ^u�����n�ڀ�����2W E�84l\�{Nm�Bm_�\}�^hg�G��3t�Ⱦҍ��hh#ӣ����AᛚA�z\� ��:��1���k@�6زm�Q3�fU�T����{���,��lEb��,�Qr�LA�k5�Ά�0�� LYs�2�zU)����h.�q�԰��"&zʚ���c���f���A$�;�!w[��nL+�x3��n�pg+�']�}�����+2��*�Ş��S1x�3�#1��uA�'�4"T����oI�g�����_gX�`Q�> Q�4�X�w'�~����ح��0����]�K_.�8>�n�kXR�����HU�N|�f-�K��DH��
03���NX�h�����X���!yI6��#�Uq�7��ǁ��F���<�v�K�4Oֱ�{4�5m��b�:�kk0PO��h�=��E�\��"j;a�z	�.��?\���<����s����X���r�����5:�����PA`�f���n�\pu��!��j���p����܉%c�̵�0Aj%���c;~[��̷k���^=��}|	fS|MZl/Q�H�YJi�Ǌ��;�:K�`�c�F�R�kF{�1%)�`�߇��$�O�e��$�����;.��a|�6z�.�.�C�Űws/n X�pw�W�9_�,AI�e�����H!�K(��"����7���T5�:��7Õ[$�3���(_uɸ:�H�`�Ƌz��L�f�s�������i�	X=s�0���f?["'C|�_M��.��_2�h0\j�¢�:��{�%!F*8VP���0rN|��T%��5e�����ڹ���6aW�&�'	�v�k��ﶠ�,����^�&���]7|��m�v���j�-�ⷺ%2rAq(4�{(?��xNn�~�L�����ѤVp�u�9��F?�l��^�8��z��!n;�݇@{�g���z� ?���^���o=6e�P�L�E��˱k����\��lµ�)�$$�;g���ɮh��6[lM߬�����̐��M��l�{���o<w�sG	@�M\�AT���<�H*6S����F�� ���7�qg�z�Uh�+�8W!��:+��v2��!����ۡ���̓KX�5�D �ZA:]U�O����t������(���J֙�2^$k�H�
����VU�L`�ɀ��QY�D;�d����d�)	�r�]�V�Vl"Dec�'qr�$�a9��(�{puC��꽸Z\K²�,sT�>H���>^�-� ��K�O�|���
da����M�Ew|�k�i|�#�@��bj[s� �"O
C��)�y��ƓJ}�8F9�&�2�<#����Y�%=4�;��An����F��Tr�W6��d�r����X
6��=eddH���yE>�Aa~zq"�K���%!�CP�kˑ�e��=�e}��-���Ē~��S��=����J��4"O0�o�)l5��>rg�?��Zʴ�z���!1��6�4�K�0�Jw�\��S�g�4ޜ'4�M���m%�4Ed����y��0��1�2��� wu��f��zf�LY��T���ơ�"�X�{/ 0�"K'%���
�a[��Ǳ� �I��AX��U`�HP]0_���L�f�m��� �]͋Rڟ����$t�ICE숄8��2&L��}+e ���F�R���\f?ͣ��Nh��+���r��K
�@:����<��T�Ng���,E�SC4��(�m�0�<`���-�,ړaz��.z٥�ᙼJJ�"�5M��`�X�/CSGM���{*�F�Q��V�i5H÷z#�!1�r���]~��s����[ހ��e����Z�
������5ye�@��\���M���v�|u}��ur@��B�A�Y����'�}5��ʘ�å�35w� �]D��؝g��>T\б[ucwFZ��ޝ��E���]N��0ݚS]����W���jY>�t�~�t$<�F�9��ԡ��|�_��7��S���I�+�X�@���4
��\.|0��>��ikm�J�;�C�8�T�̌���ճ�+CH�	P�t?���J�T@z�wcW[x!N��U��O>W��!�Q�3o�,����(�Ws���c"�Cʑ�N���k�66�hq7�׀?e##�8Z�:�<�!1��
h���Ə:�L��"=�vX����"��.����v�E}���'i	��^n�o�C�������l��ֳ�PB�KBI3Y���$:����S��P��[z����~1�w�T��4}9�+��<D�/�K`�����K���Sf<F�2�K��Nr�RQ�p�O��މB�:��-�a�o���N�G��8SB�V��6p��$�����f��$��=�wVnpm)~>����J+��9|�.]vA��R�?��{��,Io�M?��;;AӞ�Ǩ���˯��#݆B�}%�:b�x�Cr�Xc9����(6`2��O9�f��:�F��sj��5Q�<uLJp���B���mү=�͇�U('K���D�\�9��W�S(�V�5��UY�ߙe������t�$�������`�o�m|qb4�PP��&+��Ǥ�vtҍS�IM/S�#j�;v�Ŵ�� �N{a���t.����}�Vڋ�5\���)4aӡ��28��l:r���C��J+^�۝��:l��=�]���2%�羵�p�f-	|x��)Y��Q��ʈ�cE c��(@.N�,�f�AlF��U&3�;CTv���|��w*�#�w�������B���L�B@J#1R�OZc'n���t<˪��Z����W���P��B�&)e:<G�1�|=�E�@Ӱp'���my�@>.�>��Cъԝq��V|!P�9�������=u�x���L|�W��:5�S0"�Ձ���hf��T���P��������V��R	J :��H����>��}�(�����`O����� �G��'Պ�p��.&����s��lfe
�`b�nX��3�m��ߜ�L���%�t¡��n`/L�rQ������2��T�1�g!f9z�$)�	�4,ߡH]$�'�Cc��s=��W��̯���N۬w93�/=���(Z8�	=�=j?�N���H�!I���L�d�?�b\��^���u>��t�G�s��,4T��t'�@o������#"�'�1�q+�m�A�µo�N�#��̢� �cK�:�ΰ8$���%���Z�jy��������rLM������]@��L�u+���3�"�r�˂��� �T���r�Jሼ�[�%%J�t5Ŷ.(�m�w��ۋ
/��o��� ��!_^
�Z@�)iD��KA��D�/P
fS��N��#,ۉ:'ǆ��ϊ���D�	�s<���0���F�/�j������dy^_�X���DK��Z��ݢ,�s�"��8 ��˄��lفR�4��2��������30y+�RYkH��$��lY͹y�pk�OП'9M�

LI1!Q�ѓ��(�췲W䙎����ʧ���-��0�!"�MxCBU���NV�@�_eI�3<�}UZ�3a�4=i�и~o#<Jggِ݋��?m����y�,���"��!/�.�|�03@;��7�Y�$8W�/d�!'�b�#4u�ő �=�6� �J����q�.�59�T�V5� �̭ ����{:�0;�7M`=����A�P�]l�z0�y�t�T��;��n���l5�z>`f����#�rr����+̬��EB���c�!��� ��͡�cD\�2qp�^���VWz���ôV�j��#GO��t��C0 ����92Q0M��K��sN�(�h���j��F����̶�=�_1lL��o#*k��y(����Wm����*��:�<u���78 P�[ǹl[�U��Gʙ��S�**���g���HP�l���-]�N�H2>U�N�w!`��iP��^��<\�3!l�����1�P��4�3�IP��'��+�Z�.�m���������ĺ8�PW��}�p�ش���x�r�� �G�8-�,�@B�����&���1L�;�6��$y)��2.J8���I�"tظ��3�O끕�2�WRl� Te��c�m�F�v��KY�1�[�D�������f<�GA&7�?c`���#�;K)p>���f`��o�Pm��i^F��G��S	G�G��b�vӂsNw�j�P�'��t�d�1('��O����j�(�0~L��I�`�K��X�.J�=�� �L�U$��1bJ�d��l�el������ZrK,�cC��*oP)]�e���U��ݕ�Y���9��g��[*X�q����p�Jl@V�}�z�4{�>�yzʢ�2i��B���������N;�R����ux��x��hK�ʄU(	ћoݡ6��n�BR�~.���wIVm��:�<�e���lo-ؐ���(E-Y"5'���W��p)K^V]�E|-����9lY��~uf�߬3���Ci7�n�Wp��%}s�d�/����㷽�e��{��5]єL&s8e��^'#8�c~ �(i��0����;{���j��t_�Ei:w�
��j��4~��D����8��A�q�9L��tS����R��~�@?Y�-�[�0|�l��Q���o�~��"��]"��*���'GS�^VP����;�Eq�-
n
; �h�LW�����_��15Fi�
�K�W���E#KYp{�kK{Pn�E&]��d����4�-��x�����z���q�S���L�L|/*�]h�f�� m�ZF}���<��lrw8g�o��ʃ@<-���	��m=�p��+򇙘x`y����]Vh��J�����B�L£^֟��p{�Hf�^g�	���"�T��٘��Y5��^���z�U���>ى��^ӊrS�j�k$X�����&�laįʾ�<��փ/VF��3�c�*8��D�l�l1��uD��.t��e *?=�a��_.����g� �F�����,N���;J����i��J>��GU��3�F%�����O�s�!������Ho}��&,�:Q ���R�m䥣��LrdLIԜA�손н��ڿ�c��Y/��ܻ�T� �t����k�=�����������_��M�z�<y�����,����� �Y�&�ȗ�0";�*�/|!���鐩��Ҽ�V&�ʂW���t�� i�F鼦�5�lL���'�M��J���'���+M� l�.���"LI�o#d-����Oi�B�N/�	t9W�JB�����0��]/��J�����{���`2�9��N����ɪ��h��3��SG��������d��#��7�U�#�@�[8��٫2ȃ��6r�P�B��B+���`�&���g?-��Q#�\e�8	sZ,���u���S�U����q�Ԃ�����k�dR�g�%Р^�ʵ�p��&��)?�_��:��b��ێ�˲��)�q�������h.�oQ[��5���{K�����~[�俊��dHQ���0��"�lS7��0|$F|}4��w��tVS8�e����Е��>���������p ��:�\)2�d����*w$?�j�9Q	�����{� ��&�^w��Q�&���v����Si�VC��(���zܺpi�9p���%"�"U�Z��$��3[p�[d�n��8���M��fk%���A��/�!��|���.%���T�����(I��"���%�q�E� ��=e�su�M:V�KΣ3�ͧ�F1H��D'2s,�L�%��Y��׮�C�ngEѓ���v��QKC�n?�5؇������h�Q2�漿7ӌ�uX����?V�N�rU�Y�<��#,��6'.μ���FJ�o���W�܆d�<yVm�$��vz��4���{�c��3��� ���}��Ե���h��3�;�!��mr�L)�J��z�z���yO��(馷��ʬEM�)�~��y3e��m�8G���[��!��H rfA�R����nksv���\�l�"~���D�3���@����}:�B+���	���%'����WE�7n���G�V� �fT�o*E	� �jT��v^2��Q\�ف�E�O������y�tSw����e�C�	5og�Ӥ^v��ea�9ብ�:l �j>�M�ry�} CG�r������nTn.����s��ޞl�0/����1���)Đ�xp�ԯ�c�8JEG��k��IBZVPݼR0�M�����M?ҕ?��8�mW�E 9�t�Xm2j"�Ͷ.�.pt�L�*��-�/�B�;�}.!�,=�x�GMK������+���1G��� �E燇�} �X�����`UFP�6�>`�Q;��#�нI��]�C�3b\�4�Qւ�B��jXdx`8���Ƴ��Hm��z�o�gz\n*&Ef����/�Tz�Hr�F��Ȗ�����(��f��JF�.[�ܜ�b�����:뉑|1�y��,�SN	��Ht'��J�`�Z_�f���Fm� _�n_���t}���p@��11���F?�cX	hb Z#�bR�n�`��H�����g�{x���Գ�Ƙ�k�O5��a����ś}3-/��D� �`����=��M��|�U���:+�!���{�Mi�H/3s>Q.Lz;MEB�TW^��ؿ��J/��Y������8�+��t�{�}�=���%��7��q�w
���>����iK-n��@�׼�hi��2����_�6}�3%��E��y;��@!H��gM��<��#�!ʙ�����Yi��H-�bś6�p �����C�8r� ��6�n��:<����q�nR��*5���ϢF��et�F�
_ͪ�k��;���k����rnY�1�C��?ߜ0��O�7b��3T�Zf��n43�a�i}��.�Ҳ�8�Y�9!,��r��ڊ�K�i��h���U�p~g�M��A0�,C
9�ІU�owF���z���b�J��H���yclִ�����ω�fe7y�$��x��%�휻rn�W���4�r��B���t���\��ba�'�����N��|{��������(���\3�O�X�n-�c>`P�r=i�F���D���<�!{g�xP���z��އ�ٽx�� UqE|�{�����x�����6��o����f2Dx��O;�cOHǭˡt:q)r^������3#Ȋ���Z�ƕ���P	X����n)g'M�`���W�x%�~l>�5�a�FH��,\Xi���P'�낵]��|B����n�ڶA��9n��]ط��Eo��+�0֏m��5Tګ�cB�b����������u��(�g��H����HpJ�3[;ycu���5�8�F�u.��?��������~̐���4j�3���^�D'	*h���Nॎ�R|[��>�-,�W�ek��&�3p_��d�.��R+w3DP�
Q�:L]	;Kw�Y�>A��."(������X�z��NJR�5s49��~��e�$�}qB���2�(`
��q��^��k�:�G;�9vz���Gp��j�8%t]hܐ\��B������k�0�����66�cMQ�%V���E��pY�����B��FSn����{&e����Kl:~b��K�xa\
؊ۖ����R�hυ�J��H�b^��]3�L�`|SI�2LK�]�a`�T�ܭ3m�ڏ� ��˂�we����v�jK�=@VLKK������5���������t�8ex�5C��VQ��^8t��äx��Pg���]�����#e��}o�D�H�:����,�W?�#u�����ݦ�rޚv�^�_� sM�g�ˈ9�����E�C76������N��{��i� �-�-�w�2���S_����>�^}� 7�E��f�S:��w�Y(*��d���i�3��`���W2f���՛ ~G9��z;�D�*�Z
FI]/��N�n��K���QQ$��܁o,��;a?����E2�͒-��p��Y��3��fjZ�oFiݘ���k�0~6|M���?Ƥ	�J��9=�2鳹�|�Lq�Q�p��F�NCq�юQdK$�(�+3AFm&R�z<�/�1� ���L�14a|]�/��5�t&�X��kC��E��C��B���]�3��A<��j�yNs�̝��xE>�&�&~�ɫ�	�o�d4��=�KNc�P8�զ+������-�	��9V�1��+̦�Edqcr\�[�B�O���6b}0d��7=�Γ��}@��!���\L����G�Q�f|�K�
9M�4���ޕ�p�A%�x ��֙(�!�*��gV�Ꮺ[��f�	�R5�lt[�s�� �_~g�q�O�ꀋ�d�M;��S4bW��4�"5��Zb���1����&���jS��uj�c�>�p��>"G4\�ޗ1�����]e�?�A,tB\\�����F��<j���7�	)H���gR� ��L]h�Ư �q��4͇N��zki�u�݊�r��ƊF)���1�uy���S��QQ'CB�A�m �CM����a����&�����v� �`'>��H���Q�J��`�n��#9o �9�U�H�6�U�d��F�k�GJ�wDdET^�,�Ɍa���GC��S�//GQ�*x��^�}�8�.��$��Z1ٺ-���!���iЀ����P�&�[�r-Z�4�}%��2�"����'��Ǯ�È���M (���񹺖�z�(#/0;�[ٚ���V�$(4`R����N�p�ð���ԋ, ��Hd �]{]�[%_��.E���S�ӶQ���RU��ƺ�-�=����r��C�r.6�i�����3)*'�=����
0��h�d{ڦ�Ԟ:M���$�E�-%�}Ap�x�$/����-sk����(���^@��iC��dt[9`�p�*�ݟ��VMC�����/�#K@�+���^��0<��t|��޿���ސ'��ߑ���]ܹt���^��9�gUg���ؐ���R$ʎ��lq�7)�����_aưϕN�q/$`0�:��X�x��J�hQ6o����YX���V��cfW�V�����:����m���&�u���9��<H0�F�M�W�T�D�?d�2�)��N�A�7Ҽ�gn+D�|�aA��B^��j�0�������p��=j(�*k�Зv)��}�u���7�
�k������i��<��x��8��%�=Ϙj�N�B��f^kF�G�����YG��W��#���Y�c>l�
��Ź��yQ�b_ �.���_���f����WΦk�V@�9	���(��a_� ����\�n�'��=j����zx
��x�9.��J;G"�p�NA椒2mG^��!,'�e�6�͘N�Ɓ$T��.�YS�;DZy&^'f4�A�2�>,	ó���f5�C���"���������%�n�$΂N�q���$�
�-]ڇ�V
TI獤{V.,^��E��NF�u	��D?uu��,��산�����X���~	���^��
���1�/}P�߻��O�$��k2 5j�<vZBX�Yu�r��Ve�a��g��x���x�'��|���&kVm۝=�o38)X�E����ԉ�𺶠�x���*��tP�]O��m1����8�.�Jl����/�F�~�O�4�I���=�@|	B^$k�!����= ���v���`��״A��`멶�<��jfD�	K�,�ټ�.~�� ���L>#� ������z���NGc���c:�OEjֆu��'Z"���+�� �}c��\�h^4��:2�����A�+��6��yi�V ǣ���ĵ�4w�[�~2�&�ӊ6"4̊Ǉ�-����EddnF{�I  Q�(W
ظ�6!�)U3קm𩫖 �魉�Եv�0��9�Qk�za��p60�U�}����r:'DSŚ��G�]� �n��U��&n��"ue�T�~"N�JM�՟������e������5n�z�b� �N���ݐ�������5�h����L��f�[��q4��]�$��UꜨʶ1X�E^U�Z��Q��X�K��*�(�L����8�[�޴��ߦ߷1���L��$�Ƌk���M}+)jT����Q4��ɿ+���\�d���C�>��:Gj���@+t�rd�ǘР�S�Cm# ߈7Kw�/t�
�����|�Ve<T�H" e��W�#�gk��ӊ��]��tg���
���IbgP�Ț�82�e�@Y�P� Z1�k`,7a�:o��1j�F�I�o��eѣ|;h6(&߹%��oQ(8S�g�S*����2�Z�$cC���'�SȰ����|���N�}_��
+��+��RL+���	��6��P_�o��-��p��"�$|~��1ofv,"X7���DP�s���ݼ���K�H�̲υ /��mD�	CXp�KA��9�7L��iL��b�r�vn���c��[[7r�#ŉA�X�V\���I��;_bt�Ust�Qn[x	c�����
��% [Ǵ�R��؋{o�@������o�m���\�$v�3���J�*]��۲l ���5�]���k�@�H���e����GMI�i|s�h��
����S#������+.5&[ؐ���䶉�ӷu*����K�nS��	dd��ྟ�	.�n^��ct�����S,��2&�c�������0vh�֎��G��9����ղQ�-� L"��|Et������#�5? -'���T��;�ս��Iiz�>#����}:_W1�H�7��$_�׵Ј����s`"��n8B�U��sy	q�*��Х,�{�Qi�w��!Y������G�%�o�.�W(�M�Ȓ[��L��Θv"������[2�|0�Bc�i�͞�|P:[�aȀ��l���
�W��M!WS*F-���. w�3}C2���N]c-dv0�g����:̌�.ۇ�ВuRsy�{;�^����vyK�eD�n<�m�G֯x�6��w������;h�Ǿ�Ӣ�,;�A�un�O�ha����bA��9T𙫙X��`��Q�	�	-�H)X���w�,>����Qh�4��)N�J�[��V]`��$����Օ�<ͦ�*=`��+�%������$�^o����L2֨֕>»ɲ�ތ�x���ݿ�;_��2)������dQ��pl8`�4����ơ��֦����
)�W�J˼d��Q^n������&(g�(=�"r���܄w���e�>��ŧX�H�P�œ,Ek*�u'9�-m�+�xv�.Dt��.�a����S��2�on�7�5T�}�����k��¶po��K����P���o.��i(�d2�f�XH�d��ɖ�8�O�qN�*������rz��
�͛3�62g"�В���/4�y�y dSz��o8CO��p��o���(!��쁛�����<�~5H�`G�iqr�u����1�R8��۟�y�9T�dM�A#z�fN-1��w���=T�^����BQ%�1�|�g�ȋ�h�1ѶG��V�`�R�ī4:lKI��o�R�_|gzJ�����@�۶�bi�4٠I��#����<D�XHg���EF�T����8T#��V���Ҳ9��<nMOt0��*�L(rL(�Z�#�o�"~�:�(#��[�m�D�>1g>�� "����<��P��X�u5�q��hk:k���:pg?����.��B�ȿS9�7�r���nͳs�τ*],Lw��>���2�l|�����dxB�ǲx��ß�*a��|�p�E�p��PV��ӧ�m�?$g���}��o�X鈃��������<7�ʝ٤C9�����fZ։�����uPFF���orO�9^�\��lx4}_<�^ZZE�vo�����%Z�	
]m�+^���*Vڿ���S��]�)V���hî2֎~qij}��Nu��f����A�1khR�s&��8���p�U���G�����P�@je�8��m���Xe�wANg�#K �c���W�-�V��cݍ%�Qm_6���t�UH���QS�� A�Ggu�;���u�G?�c��>��緐}����߉l�!�8�[z����C�K�Jat���$xd�L���:'W�
U���'�a�My�H���yo�����4�ĉ���f��S�z���=e�^N�G������P��c��<��i���ʷ�u�$��>x�o�*l����'�T[\�~b2m�q�:
�Hcqz�l���$�8�����Y�&�!���v,�.��C[T|y("�#�]�u��ih�ȧ�씶/>#Ѫ�OJ�$Uo�r���H�p���_ώս�*3,?���y��aE�6N�Y�����Hk�2��&X?cnF�]	k<�a��o��M��si���	Je��XHꥎ���}(dE�xŬ�T˩�5[H��v*�v���ֶu�GM+@�����k�GQ�n���c;Y3����f:�{�A�16,��!����9���3������<�g4��v�B�3.W�"�Y�MQ�)�-�|X��!��:��V3T���E�^�����\��h�E3�d�J�s�X�/��8eTL/�W���/Ӫ��U|�Kd�� �
� ���aJb{��7�� lP����f�������L�Ȕm�5��yq^ץ�	��d����8a�k#�7�%K'K�^� ������ ��	�Lr�3:�E�Y���dB�
�˶Hhg-~2�qu�쾢�4��[X���,�����j�i|��F:$�$�ߠ��'�]�}��..�$����D�μ�ۺ�*]{���Mb�I��r9�U�jD��l�IcAp�'Y���\�W�5�ep�Z���uA�]�0<TgP�[Dܰ�s���IZ�^}T����qR���]�Z:c&�
{9&��"�;1�D����)7ɂt	%��w#�N;+�-��	~��s)����W;�fFo� )�����	���p�V�gw9H��fK�}�)�f]6�ˍ����!�f�鏡1�%Y��$̉�,ʺH�Q	3q��ەG+o��G?�'6g�M�{�H��u5�i�x�c���qiv�����Z}zf�f��a9��K���N�R��ՙ�������$�ǜ�J!n2�Ш1F	�]����W	j�!�n���r^qJP2�y5�@@�]�'3m]�)��3�(��g���C��u���l$f]�ŕ)Ų����a��̲�	3Ht�[}瓼rV�fo�x�+�s�sA�b��3�UԪS����\F����P��7jz(����p�_�Ø��g�hw#���i�����-˞3҂ه��&�<.�)���?��I04hu�`�3;_{�/P�M��nJ E�H��<[^�L)S�"n|<�M�2��BMd>�۔5_��)@������ؙd��گ��!�ٮ�ԩ !f��1AWU8L"�<ԙ;J��Q?��lP�~����C�
V�CL�H�&��xibfu��~��~����wO�k��=�V&O3Q#P���d�1��F��Vκ���Xt��nD b��Fk�%�]ԝU�٦�'���KB4C�j{�.��V�u�γp���,ÞHj*ޢ�?��C5�
��sV"(h1�����x	�9�ý�ZwA�����D�g�cp��4K�8|�%�x���%D�q�c+SB~�󢄴_���p5�TY���7�ɿ�n�WH�!�DI��v��
p��PIj|�������Һ�G��L���hL�mX5u�;����5�L�x�� �4Л=�J�fM	��0j X��SSѨ�~�������HW8��?`�-��\��fb�Q8�|�<{&�X�G;D3��w�Jڕ�|@���박��]كN�Az_k��pf�IQ���w:�6��Eo�#�(��U�7�l�M��^�NuT�y�_�G<�$�.�j X��oXw�;����Y6�J�f�;��]Qg[�^�v|*�Ǐԅ��PV_2ΞHv���:�Ӹ���z�B]Y���ݽ/-��sk��2�T��|	��j�����u����%�f��-+���93'`��!B��%}&O����������(6t�Î�@�Q:��ù9��w���oξ��qQ�`�/�m��|4���P
nv�,�lD�v���zF�+��aA��D'xͧqBs��G�t�"]	�W��(���X�?�tH�o4 )��5~��_i	x<�:��$��H	�Њ/�~���6x�����A��F���ϘU��G��Lv��Ϊ�u +��Ea�2����ۣ�y	��__��Ҩjz�ƿ��xV�����k���.Z`RN�-|PT�΁'�]Ɉ��S�ƋG;�K�i�H�/p
�2Ȍ�R�-'�^Q�.�L����$T`3����䏾~(~p�T�. �N�Ir�,%���_P�X�;�~��f~�N,��P V��f��/�)c@t����V��	\ŕ��~A�\c��/���1��Vpj� �$��d�G�T�Q(ݼ��Rę@��}F#�B
_&�d<��<�i��c��n�kT��f|cW��'G~�Kph�b	����K��a<.f �5��֦J�o���>���v��1q.(>�:�9�\A+�׾dp�7��f�}M��7ۼb��p�+,C�V�f	��֊�d���e������� 2"ʏ_�RZ ��͢^v�`��q͇��׶R�u���ՠ�� ���8��������NS3_h�k�	]u��A<q�M!{R�s0�1��E�`M��������{�I�@b�d�R/!�g뾑b��^�#���C��=�#�T��gE@ԛ�V�XXڒ�E��(z��=
NaJDCr&�.yr�ͭ�^$8:N�n|˰Y��qBS[�O�TI֚�Ό���d���?~�6h�(&�z��Y'�c8�/Z849G0��(GS5e��4}�\��$��<��,k������r��9��e�X侶P��e��8��D���´%��Ռ��W�Sv�����>rr/���`��Zn���U�'���7Dod���4�t~�W�N���h�Ϣ�aop�%�C�^ړ��>$)��e�h,�^w�%z'�CETb��4IE��p�����E�����Z�����62djمұ<&���V���h�'������vT�k8��T�����)gREXJ����T#�ʒ�8�#�̹�g,�Ld�.�3�ap�ki	>~�W� �oGgh��(��j?��,��r�)y[A��G��2�14LQ� Ұv���l�a-u�>���+q����%�;���PPBB_~y��f�)#xrf?g�'�vf^[O�~78����Mӧ`N2-^�vY,��S'(@dn]�?��[1�)~a;��B2y�&��Q�8vec|��X�j�MU�m')j�����(�Uq)\4�&z�,=z�e9Fp�H�|G����sH�f�u�����g�,�����	[]?EO���k�����ᄊ(l���G���"�U�w��w���u�%oB��,w+�6�q���}EOC�T 6�A٫e}�A|h�ۦ�v�]q�S�a�h���"�!���)~�4��������5��ث�&��(y��u_���kD�����Jl:���]�K@ݤv�����*î�K��T�M^Gj0�X�����:#�E��ŀ7�=�JN�4l¶��(�l���k�䰀���NE�=�C�wj��8~B{k��H�F�/����3�ļ�>˹y���`��QG�>#&�_W�r�&|���Q/.�1I}�����б�K��2><uh�M�w���1|��-{|Z�Kb�_�"��4���|d�{���1���\u{rԐ�J*)	�#�w|��F����,�'��Ļ�����uUc�jN��D�b���Jw���R���R�r���oGd�3ɡPB����]���[����Gݗ�!�]��`%x|�Y�G�X���M6�b�Lݿ!�"l��'h�ơ;��_}���K2�@*l�Xv�����5����iQ�/�a�6��D4t|�[�QF��۸ԭ4x����=���"�G+1�M3,'Z��H��#�{����_OY�5�nM`U���?��-U�G�\�֓�é�"��A�� ��Z�M+����J,�6�&�!K���s|m��XK8d�〗��#'e�����@�NL�$[�A���r�'ϢLBc�vQ��6o�j�T5�:cv����"hN xzpdoĵE�p��8�-�.�#�Y<Q|h��A3'ǧ��)�oH��]^b+����{���|�:�2C���y��c[z��d�t�x��7���$��B}�Ӑ�z��/���nP���k���/p|� ��Yc�ʧ�0�p��hi�_b�S�'U|[����&Kp�����F2޻����L�Q-�� ������v�z�'���Z7�H.X�k�������!u(l�>�1w'!/�&UF�U�n&Y��~�R�@����f�pw��mTlu������KS�Z�U|r��P�M�B�R�|����.���7��$��2�LIqJ.��Ѽ�T�}A���������/�}~�5.�!��rA���S�NTvQ�#�ଘ�TO���ZZ���ep2����'�m�v��=�!�� y=�w/U{�YA�>������Z3*��{�q�EK��@i>7X�B�m����yl&6x=���Y��y�"���K�鯦Q矬��X�j����	�>d$�r_SX	"1$
2�8ŉ>����s����Y觱-u�x��z�K���,��0�z��J��b�t�_��"�DYyq�mk�v����Ou9�� �lt�P�A�����%PGU:�&���$��j�\{��;��҈��QY��Q���vwI�"z�R���S�>k�U������T}�V�?��M~#�����T #��m\�3�"5����#1#���j�4��@��단P���Bd��c����<r�8a���t�!6��6����/�ym�	����e�R��h�ƥ*mjR���2yU�CO�`��|<O0��9P��g?H�aa>r3X���z�?8�w�{CP��(&&����+\D�A=Ǎn�a���<L��aY�3�5e���䢶�,:Vb�3)<܉]u@���A��b�{�y��T[��D����1U�;�VZ�͇���E���ՆP]�uV�2<�'�u�JΑMh��0Pվ���)���ˣ��ۅ�z��G{.�Ǭ���ք@xt�[U���M��������_��((ʑx�g�A��I�c����^4'��h��/Ҥ��TZ��$�1��`�t��e�����z�8-���7_�\ǝ?dLc`#���O���R�r����K��a�4����z!���rj&�\�G�$��p�������>I~ 4MJPN{����d�[Հ��ܬ�:��@wd˨yi&�ْ����Jw��u�E�E:/~�]�`?ßTg��%v|ߵ�W�XCΌ�k�e��F&.(��aur�r��^���	hw�vt���}�6(�����})�%��T���|s�'�\^�ڿ���ehul��i�u�+��	��)��pɉ#C~6M7��������ר��]�7��]GQߠ3/z��e!��.'%x�5��������3%�������m����sJ�40�0���q�OG�[?	����W�Zcl�ֹ����_Q�M���}\T�E+�hN�N�l0w4�A���f-
�0��L�Ԧ�n�~��җ��(C��2iW[�5�
WV�����(��SXž@�=�*����Z�2�<n3���|7�ܓ���# 1"$٣��	o�?����Ȱ�J�
~���b�V\�
��.�K�I�O��XL.�]L �_s��lK	����\̑��e���L���n������ZF)Ϣ�c�n֥�>,��{�D��M�*$��Έݡ�x�ċK���ߑW*��2�`>�hkr�(��F�������D�E�	�'eń�|_�ĵ���gi$���[���N�,�c4-�p�s��ݨϴF��K����8ϯ�I����뻿1lXxЄsW������5x?v>�O�����(i��6b�f-"���\�M_�Ao"ZD�8����ϊJ_�ʹ���Xk�$�K6�%S>T��1r]��c��LE_��U_������IG�������&�z���]��O�Gl�l�0���B}FM�ojb��sy%����4��"��<?vcɬ'��� ��Ц��w[���a�55C�D�m�b(sc%�X%G�W}�3�E�pHhP�T7d0�<��q���Hl,��I��P�ׄn�������!��r��-���8g�b���g��@�����TS�=]���J)�w�ˣ����^�-�^&mlZ������"������0�|q l�"B�����F9��Gn�x�~�R���c��#��f��=p �(-�8��{qv��e�l�=����8��l���<�	��/Ƅ��eר�*�_�Д�'u������FE
3k_&1���
�k�S���hT����(A�ѓ��w��G#���c'i����>�ֿ9��$��������7dh�㒅,䨽���;�ZͿeLO�'��6����<�1Çfat�iO, ��u<ƌ̆G��W9(29��-s��t��_�1���QV��M��^%6uj��ى���Iz���t��V�]�㳩~��F�ċ��.�#�k0��|�4����z(��6�S_�xb�ɿw՛ � 41�1���ۗ�'����$|?�%�hf���:�MإR�?���Z��6���1NHQ���m��(�}:�_;8��U.�#�2c�R��ލj�шӒ*�LڳG�ް1�q��/����R�oUsn�;_�DF��-\�Y���]�.�{g�^��qP� �)�86�G�k/�Ё"(I�9����M�k���y���H�{*6���׎�bT�3�H���8��	�bhO����g�m�^�{��=����:���[Sz.8��紊w�`6K�ES��ţ�O\|��J�Ϝ��l�����w�,�8>H�s4��=N=x;�P���/��E�k��;k�"��^���u�B�$����N��Bщ�N�������j�>��ZT`eí|$u|��G���V\}��?��=�����M3��n�V ����?��n�$�⤘�-�+��`�*�p���&��v��x��ȼ���D���5m����G@����q�̳&opX��~+ę|N��U�1,ۮ��������&<��B��E��DOr������.A�}׹B7j��/B��-+~e��@���u�Ǥ�b.1{$�����Q���S:��[�A��J�j�0*1(��]�#��RPj�����1k�U��K`��C~���WI��?�a�NY?�S5���} �N�Vܿ'D"�ut|��h�|�f��k���K���	9��1`��Ju�P��wΊ�=��~��_k��34�Lv���Ky|�F*p]��yM����A�zRNb� �07����S�9� &�.�q)�!O�Tq?ӪR/17h[)�L�U9���s[�Q��Qx�����N�@܌��b� W[��.l�P)� 8���~�Q����H�������.j6_��<��e�C�Ew�䥱�^��.o,W�����>V��
Js��l5��
mO�Y3H������qSc_^�n�(�%��mڇ����� �yV7o�7]��"���ç4r�I�B����[�K炋�~��w ��3��`Ӟ��)<�!���Hܾ��q���<Ǡ���
Ȼ|�ڴ�c�k�G@�i���=h%S������@e�J��)O�К="uHS�����Z�TE0���4��V��m�c�&c�&\�%��V��5�ov�*ɱsP�0�,<���P*+G������GT�/��H�q�ɇB�����S��K&�Ф�/���2ֵ*&(�}���3�G[��V���� G/��juc�7#�)C�c\� ���E�_��y$��*�\5�wL���
|�(}{�]�@ͥhw��c`H�P�;�H�P�_����hV�W���d" ��v�A2����a�0�錍7H��k_z��P̡���T��'}I�J����Mx^�C����ҫ~'Љ�R���Q��x�|�M��H��uv��9�_��>|���/�4��*�މ�N%�W�K�tfx��6�����6륺M����p�6`C\ͼ�A'_{b��"�p�Ù8R�!�+�}7ǲܴ��$�,�u�o�x�s`9�T�?H��	���d�w���E���ts*�i����Wm`C!�G$���Wʤ��Z���Ќ��G7 �4�\�X�Ft���[�_��/���B/�ڃ�r� M+�� [�b\���\̓�6��	��z�Eٵ��/�>��2�,����Z����#V3w�y�I"�� ���1�ï�������fjJ�����ʲ4uDk�>�9�U��!�݆_52�=X�Į�۔7�JU��ס���ڏ�!���Ŗ�곦�js5�6�@�	Ona_M��"�ew ����U�لcB]Rܥ��mZB�W!C�ps ��;�ޑ4�W�]UL6�����ŋ��s����9��6g�,3k����uq��Rڙa�.���<���Y�)ɼ�Wz����"Zvq(�8K�C��y�q6۟�Mu��#ߑ��$~&�t�����֒��	�ye(��xmc��7,��b�CV.g�����w�֫����̉��8}ܚ�x�%���;5��|!|}��%U�A_o�#C���&�{������?U�x� �p:Wb�$���H�.B��X�O���\rS�%-p� &RO+��Fхn����]|D��0�ݼ����S�ܬ�(+��|3��ƔcT���<p>��J茿[�_q/crKbaت������KJύ3����g���v�`h�fNU�+��XF��q,tm,q���v���2�%?���qj��n����P
#��(�.���.�[Y�u9I��JB�%����
�(x@W}��sB��`��}D��YY��.�W!6)��KXet�������QϷ97�.��������?�#\)hdC�=gwZ�l=lb�Q�u�ɤaC1����<�p3V��HA��&;g_�S0��}HC�),
U�V\����M7D�6�&���%���a/���k��Ro�4et|0����*�i��I���m���`֔j�E�#l2D�sfԏ\�{;�E��G�����K���!�C\2��`�K�G�D���X�������H��H���n���=�ڧ�Pȫ~��{��H��۟\nI����lC��=�Db��A��������?��q���2蹐rS�ud,���*��5�,`�Z�� Ањ8o���BM<��<#��T�����ThaȖ�4�L���'
 K	���l�Wj� �;�FI���z��U�Ph��Y�(�Pp�b�� r`��̷�K������u�C�7Vz�.�Kr`���0���O���9�{�-�F(�������齌ѫ���ҩ�s�ޥ�֡�&�"0�7 ��zB6V�>
��͓E3SV�:��ٓI��7B����ֺ̞�S^�b'�x�I��X���%�,���A��a?<�sn���,�v�@��������fR�i���>�a�-���Bp��f�X��)�w��0��)�ٴ��~�GC0u�""�(X��o����v% �u�������$D�7y{Q�}�$H_J�v]����Ne�l��6eiMT���"�h��,,�p�J�i/+�>l�UϚ� ���!H��Jj�i�]�W�we���r��٣��b
㭭5A?�zsJ��p���ܽ0nz�������m���?�Q\��j�xԯ�>�ﰍ5�
�m�hBT��	!L��}�Bh��3��q�K��C��/\��*'�=1��SۗXc7k�.�Ǭ;�]|�.��\3��?�є�$#�Wr�(+�(��)����g�w�a gچ�%*�bD���ԥ+� �{��λ)o�{�����!�����c����i�*Y��u3���=�<�*ԉc~сV㨵 d�q�Ͷ��ۙG�G{�Nq���Aw�u)����ڿ������~�ۯ��#u�S���!��..qjͷ���!��d���A���h�-a�?�.Qn�́+�쒬wHJ�ҿU�g��c9�XC��:T�w�ˍ0jT9)��A�KY	�j�����qg����J�e%jL �ѽ����t�Y���w�h��QkJ0��<33[��y��B�������K-��A� j���g�S�S8V��Z@������G������Ō*o_B�Fŕ���"��X}"`4�Uߖ1��M�0�H���&��6HfJs`�(_��Ug�O%R�acH�`�t�~2
�4��dr�_���O�v����(�[�N��?�e�ߩ�p��U��A���FMsK��s��qA����5tS8㹂��/�X������j���\**��Ml�f����w���Q���;��Zc9֘B��R�II/�_��Z8]O��%8����\m��O��)5{�g�Β��b�U��)�n�bR$��k�Ӗ`gqqR}���G���}5{G,�X��!g`��!��{R�M�EI�ӝH��A^�uCP�e�y������{N�5���O��uH�M9�/��q�Bj{��F*�c�oç4�ـ�-8?
�Q%e��`ݵ��ȋ-`u�eD�vpͦۉ��F���$�d&�=M.	����R�&�;�h���D/��@�2"��)��l~��WDw�"�m��fP*�:j���<H�88>��0��L� j꬇��q��A4�^A$��z���4�Of��ː^] 7�f�`{�9H�#���{|�DD:��_v�l�&�Tbr�)�9��Pa�b�z0=%�=tp��#������?���au.^�p���Y����� ��ă>������pj�����P���L�&�Ȟ�|@0�ի'4X��%i���a�=m��u����9��)S�q�PT㒠X�nx��gu0��{��"P"�����,���־���8vxtc��ݨK�����U'6Q'r����Ҷ�T�#��k�0�En�#M���';��+0�J�s��3�n\�՟����H��h{�{.�?����kb��Իc<�t��3�X�k(G
T���y�-��#�t@�Pᩨ��h���-pd�r_K�|�1eYصt�=��@��(t�;:�ŏ�&A�%o�q�*�~i��Rsh�>�Q��<B�+R>׎��8�`|T���b>4��{�l�uM�B��k�%���t��$�F��&o����@�)��
��P�]������ t���L%G2X��n��F����Utm�k��ӊ�F
wS�A��9��Uo��j,mB��J o�
���1���g^(72���ԟ	��HN�\Q�7J���-eKw {��i*O��A�Y����i��!:ʋ���z�:Ǖ�j�.�@C�M�l�����4�l�BT����r��>�W�Ŧ�߹Ԩt�t�n8>�h�WO��c�i�S�JJL��Q�t����Uµk��)<�$�f��{zI��G��(�d�z>����ln{�WX���+	XM�Gs~��H'B@+A'�zIo�%$�{�}^F�>rq���D�D(�,�@ 
0�m%ҨU�\N��a.Aa��ZB�w�TP�p*y�N_� l��n����F�IB] �Ӥ�*�%ǂԍ������U�N_�T�:��ٖ@
���(o#B��������s��u�-��-�� �A>�I��Qaed�yTp�WWI~�Ӈ�fIk`mP�ڐt�˻�9�/�b�Io��?��/�Y�^�(�hY7ppo>�J���D��L�!K5�y�D��f���ۀy��y҉`b�b,FIZ�+%�KM�6�ƤL
+z�T�̢��C�=�ڕ�.��7�7��o.ua;U����~uמ�*�\���>�z�������Ӱ�`�~a�Yt;p���9�*q��r�q��,�ޭ���B2m�МcP�>�a�q)��k,�cw���6m���5��T-9�拈wQπ�
�F�L�K���++�i�x	Fr�ςn�Io`��%
����3[4ɑ���.9"�i|��)qS�<�{�y���Db��܆0�K,���$���<0V97��4
=���HC��aD�N�b�9��Jק��-�k9b�.#��sM�pp�k��>�!:�4���s�`��Ȅl�p\���#T��'����|����̩/�o��ԙ�kb�����������^�L^c���jlg�i�g
�
ٶXOl6��~�E��&ڙ��w�ok��z̀<��4NA�O��bD����Z��cy��&�Ha�J��mYA<\@JW���ڠ���'Gf)��B������S/k�r�
�9�A��Dota����/�Z���
��{$^��~r����˹���m��X��~�M��z�¹��4�����}
�&�+�Ay�Y�c`����K�+���δ�6Y�$������u��
$ �X�"��{e&�A߮15�ߵ�k�;�u�Ь����M(�Κ4Ǒ�m�'Y@�
��>'*!Y�كE��]��eWDI���}f�ه�*�!��rE}d�0���h�Y�Q�h`���bRC>sU��#_.��3z)C�N��i,^<)_�I���e��ݿ�|�a�C��T� �j)!+��nkh�ג��s�^]X:���g�I��)�MU��G={NMȻ�y_;R�y��ꙮ%yq̤�˗2�G	���6I�({�ٕ3��.�$xU�J������h���"U�/|�K�z�f�/�M�ZA�P��g�ԵP�z�}Z\Z9<�1В��;`����\e ,�'=������#�.�"���/�|�s���)~>�R���E'�FJ�V��E��.�nbt;�_jrcḠ�;d�F�={iE�ٴ�¯�7ib���<��C��ح5�c�.4<�~p{yA����0��<ͷ��^nIc�ՙ��]�:�֪�h�"a�&���N�o���Y,Ƨ�Z�7.}�!4$=@#
-����[Tӽ�>�|u�����xQ����xi��G��CƩۏH_�� ����8#�����k&��j2]+�q䒰&���@��ן6�������x�^�w��a��U�,�m�!\�4����c�]�E�,eiP��P����Le����=��΍KB�����ZQ2Knu	�h}�f������K��d�{-�ϰ�T�T�BV���t��������#L��-��+�iC��U����j�bZ�O{>�-8�;$-�d�'����m�D �5�%QB���ғēD�<Π��0C����|�0�[�3��SW{�J["�"8��pαJ�O���	N��r	��tp�1_���ⱖ���,��g+*�Z�U���f	)��,��`� �Ù���������Rأ��Q�&-n]�����$�z�X��҆�6px�"	Ӑ�]J�N�6{*Hd�p�@ �;��)Ů'�4?��ynh��0�o'0��_��펛�Ȃʺ~>t.�ǲ.�z$�u�0R�R��t��$���*̗Q(CR��I�4AH.���+�=�㸗S�v��)�y��;!0\�8���(�j)F�l��e���g�![��8���k�I����WsE�L���P�SY�>ߤ�^h��H~���5\T>G�?�'�B'}+���D�W!�҄��[&�d�4����W��9��$=k�;��}�����лt��pV���Z�-�CQ�6N�eE�|X�H��1�O_¼#��2p�?��?vǹ�"Uo*�l;^���O,XO�t��S�c�JrI�*��gKX�"�@����%s>��K|EA�r`pᄉzc��M�/_�%kɷ���䝬3���UT��H�ˎ*+Ǥ�y���*�,�r����UNMz��N|�rY��RN&*����y��a�E�Mk�W�岤�F�~s���qmxGoj��0i;d�]^Ծ4�d.�������qB3��N.C�?I�X�?��GBxSH${���갳����!GcFA|���Qw�����H�A��� HPc8������Ȉ!���\�ignO�R2Ʋ6����&n�ayc`t�䦅9C6X���������.U��aK�cN-�xr�B�[ާ7���صp۸K�÷x�k�=�Olk��z���\r`�	V�v�~V��Q>�S��X�lLym��"�ί"N��5v�%:�����<1c�`P
���t�VQ���x`{�ޝ�j:��E���$��cċ�h@�F��]p���jK9�ˮXk���vu�w�-��ӳ'm*9s�B������]^��C� �0F��3���R�GR�F�;,^ ޣp4iB�C+��N�EL������|M����5(6�����ݵ�>��#hb�r����~�����o�JQ[ݭ
�dO�Q�[�K�-@3��*3r-6��Me}�P���y34oǷ��_�A]>�ۄgW�A�G��`^`��O�LA��b�b�񎼟
u��@0��I��:锆�.(bz4"{/��_�7��1��6+U߇3���K�R�{4$����Eb�a��O!���V�J�S�{8�i�S�.n���w����{X"��aiZle�w5;0�f봱�X�'*�	��������Y���oS�h��LځL:�����"SW*j���*�.�����{�֝���52[lQ��G��,�/w<�"-�P�m�֑4�����C^�6�D�O"��/��H�ڀ��.��ŏy��>f��{Q󝤲T���|QD����+l�˳�F3��㺞�_x��u\��ww	�ȥf���> ��	U�SC4�����sl��d��8>�e�gqPl�V����R]�i�����L�xH��q{0G���i��$CF;v�������ܫ��}�Dg���� �qJ�L����;�[=���|��}����\e7�ϖ2K�ۥ\
<	H�\*��q�F#@��t�{�{\V�Y��J�����v�n���&v0����qu���ZO���Q��� ����i򂥨�P:���%�E͒�4_qm2NY9n�����5n�[����kY��ػ�[���d:,�k���Me�����\_Ak"Uc�ܼ���.��N��v�:�U`��+�O,�7@�~4P�������AA��]��l��b���8"]�<��Ŏ�N�s��_#�Q.�tjTg6�@}�^߁�4�ۦ�鄏L�l?PE˗��j��������B��?�aXP}���<�(���"W�LU]$n�Fv���eAk��
sq�ƪ6��^��8*�)��T�ɜ��&���p��o����ay�Emj�/i���/�yaZ����LV3�Ev>�������F��ٺ���]PS�sFnR��C���tdk���Jd�+s��Q�?N�e�s<�3\���؂��c����!s7�Xˋ>�!K�/&?����-:��	4�q�ci��k��t�K	�Yzw�~J�K��0�0�R�Ğx�9Q�5�Զ���U8�&֤x�jD*0��P�ͧ)���U~������C0�C�-ߥ^�d��v<9�!�@_���
>�r믿y7ӭHٔ���C�"�#Ϯ�F�%���]��[ܐ�Vk7aQ�O3q�=�/Y?9%M�:k��_%��t:#;���Ϥ��e��J�g����>2J��U�U�H�߰�hݲ$�y�aM��+ۼ�f�z���rUVZ$�����4oőW����T����h��?���;��Ħ4,ty����V��r���N������&�?-}n%�;F����0F�i�#`A2h�m�{����B���03�?���(�9�'��l�+6��Ud'�Ƣj�яL�ٗ��I������^J,����� M�P��2�7���|�)�H
��I�8�U��*��T+B��ڥ�y�o�6\pi����|���'�ی��JU�K�/&�<����}*�a��w��OlNc�Z�$���f�J�@�-{����^�*��6a_���9 Yd��aZoynx��[WQxgI�����r�
���p�d�(�r�p���ƈ��K����t����Ƶ�$u���t�a��r{<6�0�;�Yzїo�SV�ۡ���(j�;�	��}�PL8�df����6���UY�7��H{J�K�g��Y�l���go�J��:r��
z��K�9q�٪������$#�'�MPRDP"�DU`*��"���`��+�_!��ǂ�>��� n�v�$$`��k,�hm�GH��f$ſ�	(�q��Mp�W�u٦S[o���Oq*B�����Q�/��׵��	�&��4�S�2ʃE�` �k���wH*�(1�/'V2�����w��i���P��=�E����RӶ��_�� wf^f?�f:V͟]���R��խ�=@3Y���W-���	˒�U�,a���	qd���j���#�~{�Ѳ���q��B�R��Lk����>���j<f9�����N4�;ʌQRX�ם�[I��׿ܸ�3���w/n�U_��X�K4�-�eN)�ZA�S�:�O��H���cD�ǳ(N�(�*&�S����GQk�V5I,(��sT�֧��Ȏ��L�r��k"��r��"!# V�=�o2b-Qx��H�"��,|�����ue��b��B8���"�h��.��A:}H
��LJ����xf�G0�@�å��bw��$7�ju;C�l$b�4"~^,��<-Ê�|[�^	�x�M�Vu�4җ��Ja8۷&[�.�L9Vb����Y�̤/��l�m&�7�4��Fg5���fvK���I�`��x��/����\���e�P9o|zb���>3����<��	<U.���ڭg���Q�:b�!��(����ܭ#�>�7K�-�	�c��O�"Z+Qܖ�؀y~�m"����C�^��!���=X����V�G��>z�����`�����Wz���j��}~�5��w/YXx�}��h���u}*��~�u�;�_�9S�EIf2:�I�;ْ����d�pȋ��I-��������	8אl�B�*���07�f��"�1��6��Ҹ�'���v=I/�����>�s»K'��tWHֲ�=�V7f�HL)��_�,��ʖ��z� ����c�^$1��L��p={�9��h�D�����K��=m���`��~���i*c}P��@�W�B�)������s�:-�?-'�5'p� oT�F���/�k:��	��l������:PD�!WC8��x�W>2���৾we�3��~�w�S�d���'�#�q����<�b9��\�u�gYA�`��~��x~�J�ܦrWR�m�����HTiH�g�u���D쬻4�T���.��1����-��Mp�Q��e�V�ֹ�u�t���6`\O�{�iN&��UX�i�'�̿%rgިhñ���$�L6��}���<�Mg��k��5��J"���^�@�*P�ř*�R��U�3�Y���~!��5��M�`渆Be?n�wBN|Ҙ�'����s�-�M�o�TΏ��P�̬�0��|o9X�{G�9_�#��bVA��&���n�	���#%ו��E6����JF��\E��<P,Eͨ������ ��%T��8����T�+z��+���׏-a>���zMU�f�?����H
�%d5��m�mHc��KSp��ټ��-��&5d���ɩبV�/��֨��ԁ�ӧ��*]K�as��۸9����JcAq�x~�roV�������kP@q{��U�����p��q2}�Tv��
���#����S�)�>!��D��f��.��)5�P|ܵ'
1�D�j�%��ܘ��LkD�H�l!�vP�.��9��	ܟ4�<)���7R�n�NH�P��VB���4�\�S �E��]J�
��-|L�]����
]�ݜk�Irol;0�v��=�y"`�~\����b�1�r����@fH�e�'�4����!־�Z:y���8t�/_����xUF%�G�Ou��T��
ZF�GsX�� �o���E�z�ؔ2ݹ��Sa�����P��e����m\��s7h��}M����j�'�ɦ��"VUI�6h�!<w	�ʳ�u���/Ez���<���\L�����X�n��XC~�g�N�(�_�|�$b�o9�∱���ՠpal�5���L�L�Ae��;�Q��{t�4��`�V8�
��7���#I��M�����J�۹��R��A�ȉy��Y1��R��^_��� �E�b�2A%� {�P�ߋMpB�����ai:��+d���l�o'=�܇����ip������'F,�y��;n^�
1�[�$���3�W��7�B&��A���o�n[z�W����Ȱ$�2	Vl�J��;�xo�ħTL�D6�W�珫AO�%�Î��V���U¯�����uQ��8�H	xT��ؕ�|)Z�ſ��["񤩓�c��������O���XF�)����<�j���
[�a�y;U�䱪3���|�:\S��B֊+q+�����tO^��!@�Ɏ[l�ׁ��'���G4����8#�)x�D���?C��I�Av������mR~�����ʹ�r�@�kD9�K�'P��RٿI�y-
�@����3�?�F��k~}�5-�)Y����]"k(�Ҟ:e��s�7���.S]�[�w�����(PM���`�<�w(;Q�^��K%����vx��Q���Usˇ����wA�i�Ĵ��,��a'7l�<O	��vQ&}#��Y�b��R_���˄U��y�1+3��� ݐ��k@��hA�KUyh:C͸C2��j$���j���S�=�)%%��5�ըH��=ʢ;<�1R����pC����Jz,����s����ٺ8 �{ȁ�YBV�@2o���۟`���y�&�Hc$��oh���X+Fr�,��̨V5�Ny~�K������PD�A\�t�U��{F�BDk�T��$����(��NL�R���>�����ҿ�����o������޻Y�=�4��~8U�9�K�1�>�gNa|k�d�X]}���ޓ���[�7(��cJ��Q��eG��Wӈ�>�2P��,U��Y��7T��j�g���,�jh%s�A���9[���sc#:��쪗�cN���c��M��Qf�[�4����"�+���*��f���S�S2$Hk2Fz�r��� *D��y�g�h�]�x��$**��Z�cF�p��g��:m�iRbi�Kjf	�����^�IH-�J�<��#$��%���A��`�	'������W�;����)��K���^����=
4��}�"M�Ӽ���j��rpq�ˣ�%�v�$�WZi)C�N���S*#<���q�忉Zm{X4��$*��D�G��ﾄٽ�'/�i7߿����<��@f��~�x�U�|E�5��G���S<T���ӛδG�,y۵J��1:t\f�����p����T�p��tCE��E��Eq^<$�|�h{H�(��fk�4Z�B�L���!ޤ�{���7s%f���~i�% )n�'�3���H8f5�J���������z��{;�%$AuIg*!Yx����D��7Y*=��P�;�ez���X��}��05�;:�V�;����x[F�UI�8Ɖ���.�]�׹ܮ�G��b�6�B��.�H~Y�*�
�p0S:��
V(��!���@ l�z�A,�������D��K��̆4�=����B�\��J�Sz!'�7JWr�M7�G+t�h%B��}�|ʚɀz爨�N�8q��?�-ǚ$�ܠg�f�^��_߈n1���'��^����h'�`���E��ǘL��	�y7w����[�ea"�z�R�%�'�k��-��l���t?�k�DS�=�Ȗn ����?�C��%�Ox�5��ˇ�>ټVPQ�G�U���-������� xU�$��=I5?#{�F<�b��Q�+ʒ�4�A7�];ʣr�~���8���z� ��|��-FV�'Aš��Uo��k�|f��1'O�a�it(!أ���}�h��LV�r;n`ڬBpC*v.I�-U��v�N$\�0c����\��k��h�)*\�M��|8'�	�G�M��"n�c�!�օ�e�Æ��?�l��9�����(EC�����X���4H�J������9�6��#:.���)�ԧ�mW��.|��YoY���}������C7�S��u.3����''NP[CD��i�_�ٚR��?��B�]�ƕ�_�r�\��ؽ@/��7^���X�Q�����u�Cr�5荏B�;(;A�d��Lv���� +9�^�Xn����E/�� P���wo���K�4=�KF���˔���@1�ϓu{�	��rq9�2:iar/���r��H�jO��&5np��]��w}�Qۉ�%��L�_F�$�����U��oʩq�f��'b���b(UI����A%��(��Ĉ�z�,L�ѩ��>��j��
�����Rd�Bu_S���Yyq��PBmf�Z�12v>����{����N����ӎ��K�qs�Q5'h _V��HՅg��
��(�de3Z��ƶ)\�D3�v?�rqPm>��fb� ���f3}�δT�bQ{U�G�|6�|����H��E�fh=�3�@s0����j�!�|!n�y�t���:{�v��jil�X��-[�m�7k�G[���޴�ݒ�S-l�1+���Ů�<�9�/�Y9J�'��Q�re��r=}�.yb���z��`�݊�j�	7~L{0'�c߆B�^�˼��g�@������\�	u[ֺ��%Ng,�pP���B��:8�;��X�#WN������$���G�d1~�U����4�]��M4������ �kӘ'J�Yq�9��X �ϲ���T��43J�5\S+x�[���	����*�MV�M4�DOkP����3*m{�v&vt \^���i���g�4�N�e�v���C$�vz��c��ю't)br�=K%p���`�t��y��>���Ǆx_�~v��O����[����,~"��}T%xlC���[���[y�9���-i,o����:�O�3OK���.q!z\ �S��K~�3�3Sc>z<V�7������Ml�7�|�D����u������+���E��h[�;�v�������j/y�<�BK
	��<M?m&B �0�n\>W�كc��O8bao%4@�;�OAn��3���3cҩ�.f��3o�b�Z� 5�N���g��K��fM��n��AP�yw��vE�I.&�p<��r�Ԡ����1������׬��x��8��ĹĻS�=���%���ĳ��8ޕ��T͉�2p5tf.
I�a�*�0�Z�2�yEҒ_7�5�6Hݚ��a���f�f�uH؈��.�����0���@�{S���æ��6�/R+������TDb�����N��1�(գ��7G�I�#�s8�H���(�;"�["rB~)'��.��b	>&{��x`��
 �_!5���"��;y�$���I�qg��P� ���d�,��H��͡�7]ηD�V����pĥoM@k֒�?���<	�h�2�H}f�hc�jδ_#љ�t:�{tQo���������$�p���_�`G{�����w���;���ٛ��g�� ��X,��?�?���*��*z�we�A����)��^�������՜i��2�z}��&�&�Kir|��t!?
*���Wr1�빸�A4�ָ��|���N��k!�XXd(N��v�k�N�޼x�*zyi�~�!YkCJO�çڿ�����L,/v�7�K=��� �4��IJ� �~����S7����E�e���a��e�Wo�����3��
 qrn��~&?�ͲiR;5C��{�(XS$,�W��T��EV%�m�h�w~���}@X�y\���Ƒc�_�|\9�����U�*������sKZ�~dc�|d�4��0�Y�� �����f�
d��r�F�w�}���1�<W����O����f��:��P<<�o=��G��Xxcӣ������"�R�,7����<Z���1Q��Y���"T����(��ά�(\Ir��Sʹ9�g�9��$�*0$<(sp,Q���F���B���O��l�XQc,l5@��H�vb���	N��Z: g	@��w�H���і���ᆲ�*ZoOj��+��
L�W�*B����](�� ��-[�ʷ���հ�w�I���gqq��~�<�3H��mg�H�����)X�*�!Dh(��v8	��{Ս��Ô�G��*�K�
7+�j����G9��XG9Sf�QM>����/��qG:�c=k�4��G=�J�F��F��K��fT��jH���wtsv�U��Am��_�a�6���}*��� ��A�,�5���L�]Y���9�2)�W��2��C�ք�%f��)��Ce��;�E���E�C�%�^'�����0�oփ'��~�F�J��V�s�8��:�p��o��n���M[�.N:�O�+��K~�ȧ(THʂH�w�sY�`�o�����,�뿠q,�(	d�.c���FsH�������yi��8���O� rK��(%5<q���e��gD���{��yD��,���2����;�6�9���B�����k�>6����|�|W#	˱�Bu�e�!��@�y@l�7A��䨻zp(� �0WH�'�0�<;�B��b6��`��_���"]5C���"�C�	;��jg��I�����O|�iK��/D��ur��E>�ED�{���������#'����Tz%�R�]�G<���c��]�(X��w�u����d-<9ɹ~T^d����D��@���P�x�
Ys���zz�+]a�9؍r�m'kJz����U�z�z�ֿ[_i�.W��&@��"�L�C����Є��O��	���%e#�Z���x/2���D'�p��o��mu*��gپ�'��`�+�	.�(�4�6c#�/Qϸ)�v���.f/�@�L]�l1X�4���W:2���.�7k�x?��6�=09�:�ϓ�3�dh�`$����M�������`&MLW��{깢3ʝ� �5Zj���%�,`\�kd��e�E��e2�"r!Կ�ɨ/�殱P��0���:�t�Lx+�p@�������$�V�6����h�@��^�g����)"�'�LR#������{��)�e�,������s�;fx�Q��V��Xa�ȻW�]��o6�g�0�����lA]�@W��H�.0D��C�@��|������=v(�E����>�=�ky�[��'$�C�x.��ґm[��|��v�����V3#1E+c�7++���B83d�<-
X�0��﹙��\W�KU����*5���@�^�OT�5�u����%㺸ߪY�m��	�p^�:�u��w�� ʍ�4p�JSY��j��[��.�� ��F�M����🆂Ȉ���C���j��}m?~�R�肜�l��r���¤T����	���>��g^�v��5�l�8��\�q��(�z�xr`	�r7Q �F���Dv_�n�=.��Ѣ:&��	%�X,�qz&��"$����u^���S+�,�qI;xU�LH:��<N،�a��?
ڛ�%�[XP�<���g�ia4�Z��6���$�#kw�N���v�Yɸ(�b1!�g��ǆ��'��F�����e^��4rY�m�L;��x����K(��Y+�!fTZ�6#�E�+Pf��T�yn�Sw6� �Bv0��9ab8����|,�%�$��A����u
��pBF�`��o�c{ݝ�ؚ������o���%���?��e�Þ��1kϺ���uλG6�|�c�]@�sa�Z0G��ķ����˭�ab�R�ێ'�5�;he^����xwZ%����B;)B?����&���T���8lE˚�g�3����^����j<ƸȢ�� �u��M�]�Ã�y_�yM��OQm�c��+2�S@{ی��E�4P�؁�r��\h���NE��n9;�u�Z���������Os��N�x2���u>Wq=�s
<-���w}G��s�]:D��O)[�@.r����y!�v�yZY������^)�F(8����s����1Eʉ�.`�n�� B���:�y�2�2�]�\~�1	�D��C���$�@z^s��J�z1;ɖ�ú���+�"���W&{W�.����U�E��!m�M���i�`<`�~�>FT@Hl��=��R���Z T������7^���DR`h�fe�(���|�I��@�*͘k�͔�0K�ʮU���߭G+�(w�׍Wl<gK��V���ܿ,��t�0<w[�n܎-�H[������N���%$Y�g����?���c� +�U�q�Lr���x�S4m�ΞcZ��\���X$�N�_�I�z�T� b�u4�/��0�~SТ��A��SJE�H\�%gS�'���'Y$�I�-z��5�[����w��$��u�-^	��Q[ƪ��I��� D����ҁ.:��QGr�w�B2�(0�G��楜	YPD�)G�w���le���E%>�I�U�I�r�o����5F��[�ˢ�,V�Å�Ji&� �]J�� �����z�� (�fcSD?j��r�]�*��y�|aq ���@unl��d��e��H��4x��7��ڻ.=��\����H	�v�@�׷�B>�G��q�M5�N�&iy� ga��#{�\a��G+�*�T8� Lj�q�A�M�[�~
�]�i*3پ����B�G��Y"��������,0=�Ł���7:�颪!Y�Q�F�>��R��7��?_Hj��{'�%@��ך����f���2��|?u�w��n��d�C���;��awif��{�y���8+P���ir`�R.�e ��o=xnB�$�p�d��왐�am@�'5z��U���g�6"���bc�g�H�p$��!�B����<�Z:���5h��Ȉ��Ɖ�(���)$� t)p�y�]�{��t� ��P�x��=��&���eGE9���09�=����aGG���0coS�|ˤ.����)�:I��J�7D��y1��j��_T�c�~�f���g�VLsU�&^��� Q�tqQL�a���Ng�8e���3�����Ux�1|� 
&̊�Ǒ�>�3�9fj4��Q����*�9&�<��l����	B��v�.���м]��+'�Ζ���z,��T��#����j��R�Y��P����Jo]!�خT(IF�a���7�HN(�ù07��
�6�,�����4E�'�UgHF�!���PN�ZqU7�Xo�Ŀ�b�+��r;�VS��[0���!c��׌Ӻ�	@����H�!���W�qR�D9��~�`�J.��^< "� ut��`z���bC����٤`�u֒�X��6;�,���
F3�:�Qy��Ss�QI�d��+���zZ��Mt��u��qG6���6%�G��-���?7c;K��adh)yE�[`��"�1�y��c�q�
��+25k]��*� � �5P�P�S �����jlMd�4gG]*D��^w���6���s��nMo��2�yJ�s!�XWPPM�<�s�7���/���I�k��}�F�$E�D�@�� z����)�s���$�#)h���^���g�	тA�'�4��[���!�{�q��~"��+!@ֽ���vE,�F�V���9�%�����8����:�#Y���� H��:����dCS~���y�?��vД�\��%�<���%*�0ug2hY�l	�M�ǜ�9�1���d�!k&���@���b�A�о��kSD��J��v�f	�����?���"�J��N���f4�E4ӯWj_!r-OK7�X�1B������4"�UĬ�|�Chқ5��UUثSka�̃�'ED�W{��8��}$Ӄ]S�t�_o:re������n=b?K��ԴxY�XZv���:Ӝ������l��_1�e���/�<a�4�H���N�U�L��Lu�}.+���R0:d�n&";��WY��,!���2��w�����T���8�#eE��)�� xD�׊^��M����<�����ˎ�ڿ�\��w���7/VŒi!@Ja�N�e�
.��q�g��{�0���s*cF	���cx&�B���j��y���snt�6�`�h8�U�p�=\
\ebR�O1B,�ȠkԺ��!
���Cw�¾2��4���)e�{��/��x����������ֿ�sL�j�$f9j�	��xf[��� ��0�;s�2��i�i#�m�8��i���s6 �nsy��*{�m��  D��'vs�Qܔ��^�d�8E%~T5�h������w ��$��PHa���V�1�o"��W; Tj���F������q3k7c�}�z�N�-�|Gj�D!7> �f� R/l�Ո�R��M���\���]�3�.-18��1?O��R�,ro��&�i�\�������) �IE��@0G��$3�܃������4 �ċ�;��6�=P�� �H'�1����m�)r�����J���	Pe��?�9(7��%d����?�;���n��cxx��m+Y���r&��kU� �>
0W�+���֊E��-��}z���������N�:Կ�(����~B�d�UǛ��4"�3��i�G��j��H���(?AN�!��Fu��<;�w�0@P�E%`��\Un���ɘ*	q�R�ض3 L�[8��#���
�����/fډ��G]]��a��	$���ϙXgr�:ӧ�Q��Wd�#�A��y18���PL�H6�"��y��r��У{�����Q{C����㴲�})��L��HX]���-Ζ�w_�T����I�9�3y�] �M�3Te:��7�P��8_��zb�T���"������v��F�:�ۧm�e���|���<O�fT�v�I�"Vԃ��/UڊF%N��j�(�T���9]�x�H��F�SM��O~;?�0~�6������d6(��,ȉw�)�/|qS�b��X����Τ��w?�<�o�:To$�:@Ɗ=:�%Lu�9� �"�Ѻfd���� ��m����~��2�6J=n�0�~��n�w�C��G##�
�4}NOrlI1�+�6��fWt�o���X*�	����/d�P��@˄�?�	zV��~�������Uj��9�pL�zD2<K'uh�9�n�����9�9��eR� @�"3��q�'cC�ߊQ�=����"����~�$�=��l��E�֟�O��u�S��~�L	��en#&��E���p�)Y/������C�7P���
��͜�\��XO���|v�=����e�nL�+ȭi���i;���S ���F�QEN�Q{�W���R5��dB`�g/�������( R�WU�9�:v��7.R�� �� ^�͹q��NDX�<��j��QJ�c�*�ޜ^hra����Jꍚ�����7��߱�Ώg�[\�&7��0�\�3X�`�>��w���q 2�ٔ�x0皞E-:�g���j!�e����
�)*��55i}�+�����/�@�/n�g���f|�; 	�ϰ�Y<�ם�@������$Gs�/_���8c|B~]z8��"n��w"ο�8V7lB��X�#.�$���8�tį;1+����i����Ε���XC����ʻe�6�,�艭P�r�6��m,�G���KO���]X��Y;_l������Q��A<�Ж���F��Y֝�/�!�@R�����M#j��	V������%�3Q��
�.�
6�-ߓ��d}ʐ�o^	,����h�Aj:�gD�����}G��#�2�H�z��NM�5�J:��Q0-o�ޙ`؎���1}GN��C�������^࿰��=,�W�6:����arj%��M2��#*L��髏5��ȅB�����Q�y��G��Q����n��-��l��72���1�64k���-�rK��_�K����LJ�pi5C��T(��Ѣ����̑�����p契:ˀ�ľT�|װ�e��^���Y[G !E�PF����PD_?>��k?Q^NZ A]~���"?��K���feX�{xw�Wp��(��"�7wtl�0жl)���bB��6���q@��!��1�6�Y ;_0h�J������T�ʭ@
��tP:/��t���P@�z"�{7� W\E�x�W-\���l�&�i�P��!�S%�L5w5�����U=?�^��D��e@>�)�!tc5�Q3>}���)^�+����R��亴�r\�:��k�����wH���@�x����JU!���g�6��b!CJe��lz���0X�W��Nbd�k�7��(>��<)��T�>�~EҐ���gQ�"5}6|=^�yk�K�y>Ќ	�N�{�L.�����t#�[���gW�׾�-h�Űǰ}�+�W�i��xo�m��	���=�G<b�5_�@hr�����@LCo[xG��^��L���^��6A4d�T�(AF�A8���a���Q1	M���ӾhRQ��"�]Y���&c�@LTf ��F��/����u3�$Sߩ����
͂nr�k}�Or.f��gIP+��n�5�[ �m~��?=��1��ݗ�1�pY�2�LC�����p��n�P�� ��kl��L�`,�C!<X�Wl�����NJ���h���pc��;�W���T�ˬMz�A;�y��ʴ�XR�ɻ�$���Z�ی�ed?���D�t�VS���>՟��9R��{sE�nGҫ0]/��:�|3�W+��-���~���{Ęwh[���|����?hP�<%��x~M�B\X��'V�5#��]�Aθ`Q�e�ha�Yaʆ]'�&\c�P��^�|V3��,@�V7������1C�te�җ�h�`����E��E���º3ԣdi���gE���b�
�BXߤ3�V:�r��Ļ{5x~�����Y\	R�� ��4��Sdt��,cN�fۊ����맋Mg2�^��IlC�J��8�(0 H3)��HLwWN�v�Մ1�a��K�+�6_:g�"e�#��k�`��i-��paў6��}�륤lؔ��{��S#��G���pvrP�Ÿ��P������SW״�f0P�겣��6����O�7$�{�9��aN�i6�AU2{G:1t �0`<���Em�N�Nb���5�f����]9usD���(�7U�)�`����Y8�DZj��^�b���~��dS�����$�yq����V(�'�OA�5��<RG�%p�q�<��-y��G��qXU�LF���;B��.��2�C�׀�G\�5�}�E�-�?�G�����B������uI�����4���Q.v�J2G�Z�~43G�ss�S��]闣��@�7����}��Z	�������}����~I&t�۽�Q�*.���PR� Dae�ɝaS��%����n1i,�f \��4�9z?�%!=0�@245�^$� �g�-1�ǅ]���M>�53�^�`3J��L�[��r��&@�v"��ΛP�!��ViFs�����FQs2��񳝦锸�i�15�+����kՁ8�� �Y�]Y��P��f���^$cX���c|����$*�����j)ߍ�"�U?�X��]L�=I�]�a�*����G{�0�o3�y>:bͦ��x��v����i�u�/�}���t��B
>������R�]��;B���؋������3L�x���&��b2v77��;ش�0E��n��4]&����2��
&2cԑ�
�@�Xc;��?,���X��s�r8C.��������P
�u�j�1��bθ�2ʺR ��¿��4�����C�1͖áM�-��b�sX�������hԧ��/�	����rm0�~Q����Q^PC�E�1r O�f �K.-�F��@?:���|"q��ţ��B�sl ��Q�� r1Thc9�2g1C~���,=l��[���kd�N]T�	�Ncv���c$z
sC�V�Е��8����-Z�����UrW>�s �2�>��	�4��ȫ�}���Q���!Wd�
_u�z����T�6��,�!Q�@w6��A/ߣ�>G��'2���?�[xV �:=e�~,�F�ϓ���$��	�k_��	��x�(E$RI������ RN�9#�Z �^'H�I,J��}KǡB�B��v��3)���~�y�},�DKWyLa�'&�1�A�c9�A���>�x�� w�C��;G�-��Ǳc�k��T����bJc~�œs<Fٗt�nI��E9Sچ��^��f+V0�-�����N�O��4�����-%�j+��N�$�g%[/z>���#�>��#H��p������o�����5���r���~U6�S�X6R �zv�_oj��4F���㔚B>���T݇��{I����uՒ�>o��f�/TW����v�j3h>p=�(�;4�~}4ꌍԾ�KZ��y�?�S:�H�nJ�_p�� ۺ\bKyߌP����Q>����v�9�:�B����38��K��DlP��WQ'��Uj�d�<�a�]w�Zd���f4B�#%7/Sl�ا���(�����������n���a��c("�W��SEYu>�<�+b�)����(uÎ�L#���g@�������ԡ��2�_.���s�J��k?��dJn�` �sCM���x:F�k�z��6��h��е!�0Yq��{��X�<�blw�u���!����>	g��	��곇^7c\.���'eC��(���j������5�����Fݴ�ª d߀vb��F��1�^ƅ�`�'B�9�*n�	S}|Dע�O��{@���k۪�)z[�3�K�!\h��C���%Je���ry�Ҿ�F� ����Z�:MF���ɛ�{���7e�����u��W���m�A�bK^���s��K0�l^�.�$���y��'lT5�i6���C?s�z��v�x� ��G��J��*ko�e2g%�
I�ֻJ �"�y!�Z����ٷO�F�fD�����Z���Y�)� �P��`H 3s��<!dKd��<��ɟ8����}j�՜gք��P�W1�tY>bѲ�=���r�뢡����Ӎ�u6Fm��~	I��������ŵ����'�_w���ɩ�:W�~9h�M����B���<E��DP�Rc�9H*���?�ӛ��Rx2qq�N�8��@�E�(��BW��
m��@�����q&V.ڛי����-;���=;�l�0K̼@������6�.B���D̕#{��N��>ZzWu�r1��T�;�{ت����M�5~��gѶ������+��B�����f?�SP_���a�y��M��'��Tԟ'��`6���連gq����_v�+��XbH�jA�>�[I��]��{��&�:~;�"6����)�mӌ�-�]��w�i6���>�P�Ӄ3�2��_�x*e��^I�c9P@"�!�`�Ϙ}�U�F�_���%�9`���	H����bbtvK���$�7�~�L��ռ%lt�4x��)�,R��M�)"�q���EƯ��͕㏺7q��ZS$INn
��$b�^^�M��;*�zA�X(��Ykm\��/��/w
�S�/��e�g�����H�hd-_t(ld8��`��;�+��FH���2$"�-��*=���97gA8 ������E�y��
�	l{S���Yq�S��uC}}�iu��æ���1�n�
��O.˻�I��	�/(�ܵ��)�QS��°��k�>u�l�P�����a�9�՝	�+O ��K��ĕY����aM�pUH���\�x�Nf�<���0��
�W
��������O����[H��:/��m�|�]�	����?%~4:��s����"�V���R�훆�y��{!�;��t�8�2�7@��'j4!�ǐ�*ʬ��
5m��+������'o2�~�R��ހk�C�q4ZJ_U��_��s]�"_�����U���Y��B�opR��3LNJ#��'ah
G�ѷ���&��^ǳ���iX���
���Ti�X�N���u*���.L���[��e4"!�Ớ5e|�U����۲���`����6�xz}as��K]KA��~��M�!J��7��'�&��O�9�(X�|P6f�.�\�Ȝ�g�vr t��$�f�Y�����/���V�}T+?�Q��+ɿ{�g�!�d�^�A3�+L�pH��g����L�'H��r���J�7�ȿɿT:T<�����@J��"�0�y�6��T}CR��ڏ�k�"W�I���Tf焧��v>ZI7l��	gtEݟG ���P����IF��� �%��˱UK��Ia�pT�1]��?� �L�e�]��%YCAg����rrFb���b�
�V.�"@������$5�Nt��ݍ���3����ϡ��߹�Ӿ{9�0S�E����5��_�7N�0l�7�#��].�c��?��:ȗ�R:����3.}(��|��}	Q�*�_CL���I�T�Hя�����2�)�ڒ~h+|xO�o	�(��u�$<�Q?�g�Q��ɖ�O����4���|ä ��7���āw��ס�$��V�҄�4RQT��0�`��L�k���=�z�U"`8���m�%J�ֶ�M����8/�i��J�%���e2�:��9��f���}��:Zv���g�&����Ar�<��ť���	 5�Q!�|�������ar"�=/'����bRMb�h�P߃z�g*�K/ 1�.Ь��sD��8ʰd��� �U����u
&�n���C��f6� ���y����q���]�af�z��?�C�2-���K����Mk�IbM\QZ����o/6|$gUu��XGR�|I��M�ۣ�;�k��3�a�O��|t���)�
S����La�u�.GI��[¾�=S��h}�hS��i�k���/��ΐ��t:���P�
{ҵ�4\���Ӗ��9�H��E�6�d|�A>�C�K����p����X]%��=��J��::�v���vK�l�5�Ѕ�%7�|I�ӄ��9�������7�=f+D�k�uDZ[̏!7͑%]��af�M��	�z��Z6U�9cۊ*����lQ�k@Ife#!�h����1r��]4��II&	7���Yh8�{���W�m��E7Fn���c�l�
� )���;x�4lR�XbD6�J�Ǉl�/Es#
`A;�u��Y�쯛�8�4I<`�����QI��1�a9Y�r|͓��9��Lr"
��+~�r�)���~]��3׌��u~,��u�k΁�R�D>�$�z���>s���r|���1��^�2Ͳ��z�;�>�	���Sϒ�/�0a��w/Ϋ֘����S��t���>��y�$<��6s���,���wB��_1��.�6Sv��՛�fҎ;9���K�cv~�-+�G��rg��v���9% �Kݾ.C�#/�W�벥p�O�᳨��$��HUS���bWxcg|Ʃ}q�>���4��w�_�ȵ4�D	f������)_�%,��ɜ�FV��:<�b�w����*�PHs}X������kɳ!����=}7n����Zֱ��2t�ge����da�YK�8�-�O��d�X�����Վ�=V����+�g���MON@��U�(�%��}��
A/$�4�*�s{�`!K���ޏ�x��7l>,�,NBfsJ�I	[�rZ&^��/�x0�����Q�Tk/&�6r�=ַ��lIl)���AJ�6`�^0C��P,�r�`8]�r �b\E�2t밤L4p`����3��pI�oj���k���joS��?g�N�Pν���h'�7�)/ϕ%.� �$�KU�����I��㭈;���t�����	�r���X^�?]s���L�y"[oi z.9�=VYU2x����3�/���z �\���/�P���:��pF�'K�|V�?�`��&x�k>�0�g��\��-r���g��\�W��"�p�؏qգ\ɺ���ӑ�@�b�"O_VY���`�X:����#��*�^F�fM�ϑ_$P�q�Pv�V�� S�^��꧳�|	��$��~���I��ǘS ��Lo�?	���i�鮉�Ӣ�H�D��\;�FĨ����%�-G���n�3Ij��1��L:���2�z|z����Y��Aa��_$I�A���P �r�KT������Ej����P��)Ca�-�g�G�~�?��G�I��=�6��hwz�
�|����xҗ�5�3~��L{v�08&�SG��
��p�3f1	<���r��l��N�|���@?���~��r<)�Ý���&�a�G��;�x��X-@��K ���I�/�2�8!��M#0T��rU/L+�կo��f�!��z��F�:7ͬy�vK���Tl#�Ō�i��A<�s#^�c��d�e�M��M	Vh�'Ym�~[��w�1zk�&���ȷ�b�f���̐.�2��+���!�1"�~(F7�%+T�y�! ]g�-�a8哣��Ï.��cꗪ����y�\X���������/K��#Z=R���P��O�$��W�3+�ӽ
�'珹��� g������q#���T��؍�#�z�p+�m�*4h���8 B2�*�CN��k�<Bg5a��P�ð�gc`�m3Y���
,��kNU��G�ѱ�	w��g���z�m�P�u&�%۶=bt��˧j��gvEd��x�8�͏�ʭ�sXY��vWδ�ʹw�[�0R�nb��^���]8���i&4��������u�0��������9�7}��]��b"A�lR�6�m/�ߠ��n��i�EM�s[����
m��s1��+�J�]fbϮ5����q*]�Ux��h��_���x^V%���4�pL�Dm�r���3�ҳR�"у��r���l$�U`�(����'���O�H0H*j7� "?b��9@�9924�0|m�.w��ԠU��MO�B!ݽ��#[B饽aԐb��޵���8���l  �t+|
Dt�n�s�V��{E�V�T�S��7U�1@���Z6��j�0����:R]8�<���������3,u�� W�T\3��K�u���2�(�jp`ZP�F��� �=����	�;��.�Q���ƃ�1���w�=�@S�q������
���m+#�����ř�����ݑ�rj�(�HӬ	��������X���2�M`�8��R�I��\����������n��%�s���V/�byK�j�����^y�fR�V���5�iP9kRඵ��l�����uK���C��E�#�=�d��#:�;T�jo>���/;��/���~�A~�P�1�hA���ozY��`��ք��[�����a���PH�£IexqtL��/"Q��_{P��fE-���SH�/L��5�mW{9T����1�ϱ��U�oKp,�?���t.5}�F{f}	�����?��G�>�U���r�W�3�Q�;\�pq9��w�O�Jx4$�W�/*Տ��h 4�ޠz�8)<���
�Q_h`��O%Iոݿ�g#r�R�9ׄJ8�S1๵Ǌ��5�e|g���|�vI	��L�������T%����ã��:�)I��O�E�V$�F,��0�ڊ�o"-N�!�z���~VJ<��K�h��۽����i����ػ�r֚����ʳ!��a������e,4��t4ɺ�R���Q�d�'�JG��iG�'�.`�1X7�>�c����9d)�� ��vB��Em�� �`S�]-�}&�����h;��?K��R����X�aq����%��TׇD���ؒf�q����f�����L!���N�7�5)���dT�	5���<����{$��~H��Hݲ��H�$+[��h7=�;���{����g}ƛ/ļp>?��O#of7���I�'�9"A[4Ru�n�J�����Tz�N�_��+#r�NMC~Z�g �,��	-p̦�7���u�ȩ�����z[v���6�)^�ެ�.������w9���E�ث�,0��^X�fQ�����8���I'��m��� ��4�ҟ�e��Wht0�K��ƚ�>-�}������%�6��';z���k��햀�i&�S���U}Owzp��q�2I`��o`�E�{>�S�U��mRF��6c؀�A�"Ǿ}/lj���x|z������S������$y8z�FK�ݻ�?rSJ��5[�5^�v�3����v�b�v��cg�SW����%��|%r��fȅ��ee���bk�km����rw��;���s�톓e@b7��d\C� f%Ԁ��y��8`���a���_~&q����J�@A���^īz���/\��'HJ�a�_���D� ������.��K=��s@p"Z޿f���� ��Z�v���<��Ǣo�:k����,�
�� {�I�k���؀���gE�CP�l�")	C:O���� J?�]@�8o�&ܨ�~E�'~t������B���G�J���@�_�&	�Ȓ|��8t�d��=�A3���DLo#�b�$��d�b$�Fr�� �f^��/&��h��o��!d��vϓR�NB0���o3P*h]�Vqش�f>��"%����!��/�v�NA�1����X�I�F�ӓw��i߆ �����~����g6f�ȝ�|t��>�h㜇�A��.�b�j����K�z�H��蘟�&݅O�ѓ��K6F,*���Xd&���o�:@,\�[W�N5�k�
�G��G
����9rs�.��V�lSuh�O�Xnyڊ)���%�H���������̪U�N�J:*�U��	�G���"�P�8��~&:ܴ�>�
�4���+y�Q��6;�݃��&�ea��R�5��|-�ku�����w�sn��'�=����r_�w�Fq��ھ��z�0�4����b� ���=��Ù�<�V =�������Z�Z0��|��l[�$���A�(WV��M��̘�\e^b'\�w7IaB�T�,ll�]B3�/�q��]�>/��-�NE����ŵv�:��KL��s��X\�:�!Id.��)T�(F��!'-�eT
��[�-#�|1�eq�fxr�?��칳����~8�U��?L>��8D�����ܵ
!]߈��ІR"�P�	�~��Ȉ7b�L�@�Zez��`�S�h���;��1O��Z���p¡xV�)��-����x���}�',�� ;wUo�҇k=�#���_3��Q�0�����'�rb^TO�? #,/*5���
�n�V�]O:�(�����m��1�-�;j�
�#��+a�2v�v��{T�V���}lm$bga}�OH@�d���N��{��aB���'��.aShh�D�f���ѹ-���\{
	(�3@��tQy��a��l��7xS�y��T�w<�j��շ�>k�ի�֜.��6͂.3�����=..�?�s�0�D��#���N�z�_��=2ICf��L:��ZC�d�j����z���&q��cdC�|�UyI��ǉD�y���*��N��m�zP�K���Q׊����j�9��B;����X�<@�:������z`��LQ%�0w��V�������+�{
|�&�Y%��kN����w1�N�p�0'����v#���u^9��w��I#���K4S�������Ғ-��I7�zI��I�T�&�Wn�1���F`�If��ln�A��a0�{��p�:8��O*1Z��~8w�g�-FX���4�wL/;e	���ȑg�ǔ�Sb��!�^�S�2��4A�@��A7��m��F��W�H��s}p�T����/Bo����$�w/,�����2��~Z��������ѿVt��dG� c�x� ���SV�b��������>	�LmBǼ��}�Y����^$�E�q� -��4�]�x���Ad����杏f�j�a�I�&Q�&2yK��x|���7��o1wu�b��~��߳+4��kﭦ�J�w��P}�M�&q�l>�<��>�W0�G�p�4�%��X��k���7ʳL�q�OV�x\�xv'U�� �=0OC�b;ahy�%^��9�*P��>�V�,��ݬu2�;)�=|����sO�9ਓMG�Ei�#��+�x�@ˇ�"���:�Uq�Y�"� T�*���&F���rw�0�i�QmK�}k��ОT%d邾ei��#���}i�c�ab��>R�������/�_���{�~�?@���[7v����Ei%�8Ա�h}&P�3[ ��˥��_���5nwH�Ghr<�.�|�(�	���.#NQ�>�<tu˟�M��P]ͥ����Hf;������Y*xq��@��`p��#�K�L����TR��WDM��B���\Ӡ��)�NL���d.�>��a�b��z�/�g�^�{�g�tl@?�(|/�Z�IM|�z�{�����Q��s�O����>̲k�}_���P�\����Q��0�j0�=3�Q���.�ū��;1P�dE���&jB����bW��Ǳ���9N��~�Z+a�h*���g�������(&���ܧ�!Ϗ�����bv��xbq#qY$&	-R���}�͟i����s�H*Q�A2�C��mq _��Ʀ�)ӳ����<�4L�nB��W�Ps�R�p��R)f����p/VNɦ���e�"&��#�'poAgxק�eb��$TD��j�hC�'�t�dQ�.���չ��6@EK��+�N�<���33�8�QR��*OF�r4#�Cl�(��eKʆ� F�,bb�����W"�f���&si��oP��=���VC��N��5���s�Z@.5;�ݤMsB���]��h#�=J^�Ois�ן�-ځ��I36�
e���!4R^эC�<:�W2sTN;=�l��R݊�ʍ�Oe�MI%��.�鯋���X=��>i��}U��^�m�d�5����e�^�D�5��t�)کZ|@��.���Ko'�X���e�O�>�a������ɸv��4���m9�8��3+���ɠe�y~��q<AW�U��/�HG�,>}��?+������mgV4;��&�������B���ֽ�Iw��k���j]m�����Y�:0#���_`w�Z� Ps{�E�lFbl#;����ҖE�[փ�o������[A�û��a Y�|�E��cE˄�;O�<�Z�����ׯ����i��IIM�yrߢ_�o����-r���,ӫo'�<.6�m����U�\8
3.����ε;�nsk��_���M|���6c�(6Sᒹe�NH!����T�f��ٝ��?���K�-��=e{�@�Q܁}��!�g.��_]dy����g��P����VO��t��}�A���X)���=>�E@w8���)�;�1^������̭7)(�� A��W�6Ú��T�E,[+�|B�*��Z{�H����K@%�|I�u!�����HQ�4�����	�ʵ;�B|��~;�	��+<�el�	��H΀�<΍����(x���P���W�5�1��PZ ��lZ����n�gS�,b�c�f:�w}�E0��5��<�sק�w�CU[F����+�����T:V4��NB��N_��@t��N�b�7�l"��̱�����~�r��M�f��T{��l�%�E|�ǎe�@����%��q�1�RF��Ua/�þ���#g"�|�x�\V�=�'y��X��XP⽚���YW;��5oa>��4�u����%u���퉰71! ��($�@�b�+��5�]D���*`g�Ѧvt�������$h!|���|��!���5km ���zqXKm$rM�VPbDt�<�]L�ҩq�3!�%b�A����>�Q\?)���qBQ/a#����P�x�>'$oތ}�1�Z6�<jbr�)V�k.���c����cR.���Q�k��Ō|g���A9>���m��_ɡ�hↆm��7�M��=��Y:|�=�� w��eA�綽4��[�u�>�2�\�'&��&��qEy��a�d��@��C�� ����x�9��{��VQF+�y?�B)��cWPgc�����%��O�����I�!M���(��D��W6w?����ZJ�,V�����HS&�G���UhPg�̏Z�~���d�#��̼���rA�jLǬ��]�[˭�����=U�;([1+�p���z�g	�����u�>��N?��z3`��b��0gU��]Y��)���vm���ly��Vj�C��@'	�a�Fy��}�
�z�^-�~`�T�mM�+���ޱ4(� F@�)�������m9�[��1�8p��<����6�o򣒱�'~��huˢ�gN����[�J8�,�����6�_�Ƿ��m�r���3S( �)�'�(KQĂ��
߻g,���քƳ��\nt
�m�_)�=�[�^X@Ʃz�����X�3y�����8�Y�^�6�����I����~�Ǡ� ��fGs�g߰x�M:W���D5r>B|�C�6�@\۽^׼?�k��b��f��-Y�A�dU�|�̼s�Q�Stu��}w��KsD%�?7(9G.�OӺH�)�����4Z����9�,����� �Ѱou�a���in��/�X���T��/�/8��՛w��Zw�3C�����RV֡�pd��o�������>�QT��>�o��d����_i���AU~�����"�Jh*/�����?]���[���j̴s��/3-�����R'2hw���$��Rj1�6����:O�J���g@�ٗ��c~!�ȿnG��0�
+<-��h3�D\pv��=y}A��|�c̪ߞ ��f��y��Q�nu����)�.��Ma��w��!���*:
���t���^�Ә��#*���	�:l|�d�I�����_�]��i	땨������J�!���T�$C���� 7� ��ЋZ�:���8��xp<��5SѰ��4T��h��ɟ3p[������?���%��h�H*,�
�Uh�*	��w��9�z#��g~�M�
��΂� V!�E��o��^2$��U�R*{�/1 6�
1� Q��ƥ3�/n�fS�/[�W;9:D�(�V��>���#�d!�F��h7��}��~�ܩ���U�^��E^�&��<��#�qg�G:�]���]M:������[%_.���>ш�y�%���+#{Z�D�4�z����D)��F2tD�Ox��E?Zj�=�e9$�&YO��\H���Q;�v�r�z�B���X���^��Hy �5Ē�R�,<��L	���.B�P��G�/��5��k��M�G)��K;� X��U
�9M�!�	%F�{��7:��5��PG[�����	�%��A��r4?��B�lw�14�+.��kO?�i����4h�ps��D��X���R���/=G�fJ0��($-t�,D��
���L��Qێ�k�/`����>�ʱM刹���%ݧ�0D�֜m�S��_��`Q�9cLg���`GN�r������tR��)��"�(�;�yH���g!�������O>���|�i׼��V������)�-S����;�8iS�ϖ�_��d��l_�J��PVߴ�Ӿ���[�E-F�/ �3鮜�A�z�q�L�(��	��FFt3�pۃ�N��E�������$�%<�i�_�R���M���Z�OP�.��u ��z�{q>g��j,���w��o�YP�ʃ��P�Ww��]f�Օ]��8���xI�M��c �6[�D�0~�|��6ã�J%H]��{3/���>^o���H���+�"��\�(_u���,
��P.��Gs(a�⃔������)��.�+l�Txm�#A�*�H���b���������D}��K�?cQ����,\:���c$T�o��aL?��d��A��p��r᳡ܶ{�O�'�Tm#�M���ZC���Ѿ����툿�o� 'm`kt,�s�1���S�N[X�B7������۷"Q��Ey�������t�)�]Ţ���Zݦ�D:[+�n鉨W���p�<�#�ۼ�;�F/؇pLpK	+�-��+A쎑����	>�p��^A%?N��y) U��f��m)fc�K`aR��=�֘x6�#��XHۣk������7l�Xƥw�T��c5�6��?R��Z��y!�l]ży`�[V��\�����u��z�Lj0,���><�ZvJ��-r��F�����u��:�AY;�A@Sa4%]���<e<ݎ��S.�� �:[᫹,َ���Ǧ�����V-�URaj����Z_�B=�)>8a��y�'<�ҁA����oZ��+�~�;�(G=���W&��@{��9n	�І"ZО�XW�E����{T�'R��_�w� S ?�|�%ɦ�v�S������Xn����TxY@�A�8 �b����ؚ6�A/�l|>3D�ժ�q��#2GE��9@==��I���(��ꊿ�6K�!Rv�ε)��廖���ʘ���EyB{R��數��`�!ڹ���U߿���|6Wrٳ��j�����zu�Oz�?K"���-�5N�o������oW��M��$�4��Q�� ��+��,�)���x�4S���yf��\����֥ pGT�"�Y��W¯Z�R��r#�M�kx�	O��aŐ��y��
���\y S���6w"�t��#W����]k۵a�mPK#��	aܼ��}|��Ǥ���?�D���/गZ��88"c/?aӻɱBum\�����vK�Zĸ�Cr�� >��D3��#0ms��%�Ä@U����?O�Є�{�ɫw�|
cʡ��_��:�	�6.���A�<D�=��FO�H?ː�R��+�x3��=�����fW��)y���M����[R[l��M{5S��Ȏ�aT��|<�!�W��I�mJ9	����U�M�q����wk��ydr~u�/�|�@��%BE���
�(����F��q�P2���A�J�B���u�X�p�)l��S7����0)ꫤ�q.���ו��\K�(&��ĩ��(q�C���H;���vKN�~��N��ߴ.��Ú����:r��Ǚ)R��}��G�������:�����/F��Z�;wH�4m�E!"��*\tH˻�����YJa�m��&�iy]�~�7	N�W�Y��%(�8W0ѧJ"�2G��ߑP(�([p����;nOjݸد ��\\�Y�;��:}��ϑѣ�J]Z߽�:=�K����=)�㳓J�<�$�I�.GnV�/�ɱR9 >����;O8,�{]�Ra�?朗��m��9�u�ύ_[�/���s
*�Ȋ���E�=ܣ����8�՜\�*hZ��<�\Lhn�Ǘ���- "�o���=�?�4�2ڐ}?���K�YD��F����%�G�r�
J1�B��76S�G쩠�t%$��vƜY�s3v7�/."�1P��DMfﻳu�6�������h'&�oi��=dF ؼќ�o�`Sm`�t-��F�o�~��B���#.x�	��@oL���li�6t���^�?�#r����Db��H�E��2�pޤ����.�pUu�Q�wۧL0���zۗݼm?9�$���kc�� H��&ʩ��z5?����o�J�w�gK��s����G[��j:��P)�����̱�w�L�Ȫ<�Vy�S�1H���.q�S��Q���Y&~ ���U%�)��P,Ux�ֆ��E2�~y����Os��7v�-y���ΕGL�H�AapQ*�]d�=��m�Pu�S�K'Q�Ld�x ��i��u��2�YO���H$����* .�'�� 	�j��H�4~�/kjr��XOR|k2����A����{�E����ݷ�>�}��`�+��ܖ�6����L֣������i�~���	í���kX���tF�e��t��I���L4�����G����l�cTM8��b�s\E�؄_��/vu����{��h����[��2sr;?8�Д�4���GA�a�s"��?�A��{��E��]��p�SI�2y��y:7��m�d���mDRݹ�����5[�.�� �>�0�~��k�D�|7�%������S]*|)�p��b�� #�>/YJҀ!q�b)�ʓ<2g%�G�.�7F_af�W׏��Z�O[�]޲� ?C�"6�d���x����:?���ˈ�Ǟ��3m0|���,'��M�]+�@�=!��Sy�aJ������]���5�'F I�8��Su�ֲٸs�	�	$c7��B��˳�^�97�����-�	-uy	<�`����s
��0�y�wB�M ��d���˥�p��ե_S3��6��"[E�t[
�ĭΛ�eKw�Y�J� \��I��W"Z��f;x̍b6BL+��cj�����2���zl�Ť��7���	BN��8lՂ����G��K/z�j"���$��9%���H�� ���"���0'Ee�m���4I�,;k�d�&M��^*�DY����ŋ=K٧J�}3���̞�o8�Ixm�߫�j����gO8:{���3Q�G	�Y~?���6è��*V�됤���W��7��a�3+���h��)�'�x�E檺y�xM�A5٩����T�m~H��l#���~|����c��E`).̈�\*u��Vg��q������?��Ն�M����iyGe�F�r���������^9�Lݦ�p�H�.�����v�D�S�̦��"�	WT�Ta�����2^��� ��E	 d��P�x�Q��43��� qF�m�'0}�ԅR��\��~4bG3R�Ƶ��ZS����AE^;�9��^�v{2�|6�iD2A�;`<�r��h^��;���#E�����K?-��q��@k*�4������L�r�1N��=f0ϐ
��e=
�X�v_hxh��T��>�.G�l`G��׉;��TT�|�
cS	9����X�� �m��C�	�Ʃ)�"i�t��.s�'�<T|(;6�� ��x�˱��1�ؔ�fs�Y�*�׭[kƥ�)�H6�&O5㭍�Ri�آl��v���-����h�J�rԲ�\[�cHhs�|��
	��x/;�(�������r Q}���v��ʩ���q�ġ���"(���[B&b@� ��L]���G�% i�Q�[����󕆧+��T?1�u�T
�F�7#M�d]]��T*m90�4�����{�>��y��{�gg��%!��oќλ����*�^P�>�cr���!s=�0:SXw�]��q�ۦ�jϥg:�v���&���=ý���c	S,;51 ��48��(9۫Xkg�=S'��i;2/�W>��l�*\+�tm`z{�l&x���M��bt�g�U�J��"C�xc��EI.�dv.\�2b���+M������IT9L}I��V~�h�,ι�-_������d����l�vk|Wm+��8��ǁ�*�g�>������	1!�_��2���$�`�|_�pX?���V�M@1�O�6N�%�_2Ý:_6�i�2����x��m���?���|�_�#Y���
 GN5���� �"��#;3D��d���f�\����۶�sN0;���\�U�����yo���Z3��w���if�h"!.5"�c�'�1�}6Y�U���:grBfl�}�p"*G�J���w���n����G,��j؋V�8#"�c�OeI��Qd�|x}��vW��q�=2#� W��Bt{�$w�������l��r�}KO�~�s�q1V�I��.��`��_�g(Z%�l����;�i�[�$=\���B}.6��e E�ҧ0w��{�D4�4��dG�G%�d��G;�GW*�7Uc��UK"ٔ��I
o����`�M];"Sv��	�\��xN7Ƣ*��+�YN�|8Co�щ��ۛ��Ru��F�ҽ"��.��]�`R$A����P��=S@I(����-�y>������u�(����W2n����_�����N���H�jv�wzD��.�	-����]�XU+6��['�2��Լ�[%:����F�;i�gg��i\�r�83��^�݌ƽbR��u�2̌��`iiN�t��<�8"F�M��a�2����)�Ѷ�I}��lr7��i��0ʴl<�ˮ&�R��x��H���&���yԔ9���W�Q��ۉ�fǎD%;�Kx颏��� A��~d��6���Q�L9��l����q�r�Cћ8�g�<]J�y'�[6I���T�o11�T�̒���PM��|k��G;>�N	����G��]��0TGE�"U�Li����v�)B�gܺg��A4d��Id�w�Xg뻹�M��ׅ�n1W��*��D�D���޿Y�h����[̂1fվ��Q��D�@�h0]���pQ&J�ZgĘG�ϐ�o�B�̗��SB��0-�Uc���=��s3�5�n��Z/��i��r@�M?!�% `�cUQ`��<����}����!�;��TO8�E/�kJB�'����������v���x��F����UϔH��r����"��Jv��h�7I�,7�s�t)�*BBn���\�e(!����M�w,�w#MH���M���\��~��(��?�l��(E]xI���@���?�bA�e$2��C�F�:ȑ`��V.=*�\�g(m��`��{�]t:w�!�F5�E�Z)uAJ�������]k�T�ך�n����&���!A*U��rNy\j�����ү�;J��2؁���8�ړ�e��|`2�5�s͡ҊJ��i��'a��^��o�KQR��x^_��}����3+��Km�+�M�+2�X�8�y����*�Ry�;my4٫-{�
��`��쐎�Pĥ�M$�����+�w̰a^�b�F7Yb�X�5�H��7r�d���֭���Z�kIv���m_g�Gk5�����%�/��2[͞�B��qQ��M�'�o����O�'e\�"���W���C%�_��:�%^0�ә����F�M�-;���K��95�9 �6\���DrϾQ�7��$���@��!�R��I{Nch,�����	X@�k��4��?uU}wV�������e�#�
]	
���Q1���E�]G���-r��aK��XÃi��i�����<�3��~mŸŹt�����֮}��\ӹ�!��/9w&v;�Ā�48�jx/�$���b"?#��MQ�1���ʖ��G�&=D5�Y/s���6�r�w:x�5���xadg EL#�P�X�g�|��Y~��Mĝ�J`x��<�O�p���W���[�>M?��o9B�'��;*P��NK7�����D��ի��͉��P69�s��}y�4gweJ�,��e��a��G�^j�DEʿ0I����}����3�Np>���f������_KM�w7�\�eu�*����=ɉ���L�KD�J4\�n���eb��Z)C��r[��d��>��p��ꫢz�Z��z2��Yj�M�����n���5R������[�"�^5h�6�+��ƙ@�|�o�"���nw����q�;�lb�MC6��C�~P:�c�'�ގ7,�N*q/@8�,2m�σT���K�ԑ�����\1�!@��q��e�Sw��B1C6�H��y�dmq�AsT�SO�J�l��9�7(ԬĊ����$����ddif�-��-���إ��J�r ,��/7HM�"��3xY.�1�*7�sR��"�
86�og��ܡԈ�M�����O�LȢe��~ُ����%�V��߃�C"{Un���x�GW�X*��}:r��g�á{�G�b�6�)Y�q��O���-��k'�t��J�ݫz����̃��C5Sm��k��y�a?'K����'��/��B���d/�-ܬl�u�a��iuފ���{$��I6q:���K㋾?��Z�ܳ~�J�"�%h|� �]�X!���y�K�
 ������xgX�>���j��+�4j#SE}����v�<�Y��J��f���b�Z:�w9 �|���/	��X��ʌ��z:�Ͽ��ƅVډi��s(��s��U����x�𴸅 -sK{�T�pCQ��L�〬v��+>Z�=��0>Ɂc���^;+��JP�<��jT��+�煷Q�!Yo�BR��͢���]���7��(��5�g��=��J	A'�[}m����EO�2��|=�(�g�_���e���$y[�v��v	w�ͅQ��rv������'�H��i�0���5��Ճ�q��Z�޷�jh�u��]�U!n	U%Q��KJ�<B!�pֿ0���"#������@�a�% �������T[�07g��V;��ڌ�`^�᢯b	�S6�J�ͽ$&F�%�,1vk ���/F�u��������;h���B=���p�s<��
�0�����D�?޽x�mu�Fm�	�n��4s�5��k�Գoa]цE�1�p��Zr�vh�y�t���^��)�ޜ� ��V�钳ْ5�&���ì� ��'�B��`��)�ٚ�4L�޼����<�͂\���F�[�zo;�Oe�Y����,�4%}�� ���6*����C-Q_N�\^>D_��!�e��ǝ�E���pԻzn��@a�Faw�h�<�2��f:��G�u�^v-���(Eg��=R�4���������P�.�-�
ٔ�<��(�U��k�Fo)&4<��b�#�KJ����h��=�(2�l�iQ�y1���x�ɴ\�r�Z��,[ (�v�p��<�쨧��K:w m��w���XƐ��p�#�$>G������+e�Ji	���|�
K/��w���ƹk��.�I#�nw}��+c����D;��B�hoK@WR鎴�鲋A�1�Il ���e�t_�<@Ѻ��R�p���-�	��d>ԏ��A)�)��a��'�@ت��2���H;Qw4or�<�f�K��>����4A{���P��Z~Ȍվ���ߑ�%�,%��������-0rľ�,��6.<~��֬���O��=�Q��	j��f�y�4_3�g�[����E������zjU��.'��I�E7@�Do.�l��-�XA(#��~�AbF���ㅫ�:n�u*���F0n[�T��R}�+5u���(�u�U�GL8�(�2�%�j����$�	yv���$�T)P^M�/���N<k���1�J�`�P�s�VM��6�p3w������#��G�'rs��e�"�^�!�����ZޓHdJ/�A��-�=p�)��]�����7J^� ��2g|�� �G$BN�儎v]�{�"�W!o3Ԡ�@75hR��iwN��T.8ҙ`��6�0٣���]j�g�q��QН7d�
Ջ�zG?��q��㝏�J��p�A�7�-IK���I_�*	���e�o^��v�t��(������P�j��MJF�����8Ɉ �$�.��f�@ۊ������9���ժ�[�b}��:!�e_È�6�C���E�J�X����`�zy������g(
Sc�tf�&�(-� (8�7�w��<0�[A�(K"F�����`/:�����5�B������p~�-����������#�Y�Ei n�T�{�&�{��M2$�����}ryd#�/3�)�q�l�o��I�P���8`{�6ѧlVkĂj/`[���5��6_�Ԁ���C����@+�[��.��j��)7ٗV2ԦB��JtWKXt���m�u"��/eR�I�	M�=ط��ܵ�*W\n=bk!���ϒ)� !���2�w���~_
�0!����{	�Z��l�6��E��M�+<
:�>`�9�.�Xg�I�W�_�K��J�B*����V��!S���s�W�d���I���lC�1�W8�h�MK���~�B�aYi��y��:��o��5Ń	����b��ۓ�u�T�ʼ�(�c�s�������ӣ���}��N0�p�};e~��?��3pIDg,y�v{���h����"�A�R�0Dy2��,Td�3뇮��t�]�g��Ͻk.4TM��
1�F��68Xo�AG���V�0	�7�����fd_��<Ҡ���Ԓ���jҧ��"K
�^L��~�58���u˚{��r��m�����dzy*��sV��v����稽ۢ�_�Z��a�=d�h0=�=,�
4�U�^ �@�*���$I�Ջ�����Y�6|�*~��r3;r�����D�v�m��0�5Y�)=�{��vhC����J6�#E�V�f̓��aqEԪ���3l��<5�$��3r��#LSC�2B%��J/�����R.{nE�Eh�V��y#�r�lV.��t#��RӦ��]�M'� \>W���zb������G�V|�0ý\�cئ��>��<hs0ƣ1N�m�䇅�,(SI��x���}6e@�>�q��u����==(�w�xA�O'��L7��__W����U���ь���~�l�4y�6��O5˾�u>�.���7N��0]����(��
�R�D���7������L���k�3���t���ߢ�(�'�	���S!$1$|5ᘮ��{#��J�Z+Ӄ�%��$��_ *
��!j�̦��͙���$#Qj��:ނ4��|����%����ub��j^��~���Yt��
0�s�9ϬG����kM�����/��`�.�%H��H 9:�W
GdV��.篰�Q���h�p�|�-�y/�;	(g	K9�}���|Q���N��৮����釩I{����Q�m;=��P��dI��1���T�o>�́�O�ávfR�Lz�D)��&b���a�-����������]&JW���fV4�~�:�;Lg��T� 2?[{nX�a�����J�j��Q��c�L�>�UskLcG����!��o$m:&N�8�coUƒ�4�V4	Op���/��Ϻ�t�ؖ
T6����G��t��S,A��i-/x�٭ΎW5]�O49�{R��m�=B�[���,}٫LNN��'����q�F��?$g�<�~���nu�� B�����eP}4A��ޡy�r���Nő�Z%��D�9����:��l�ppEm����Њ�C�n:�1!����B��R	-֪y@N	�֚xQ�z�m�#�C5-��������U��8��k��0�"W�IW�B�NF�0��� �D8E,���
Ixv��I�+k�P#u��@�S3��2;
{�E�{�H� F�CN�I��Y�N��Q��G8ܚb�NNC6��SaA��̂Ta/9G���bTC[������~��-� h�!�/\;�����s�Ġ᯷I�V�H����s���w�Q��m�G�<�y�z8���q�1pZ�dPڰ>�Obܲ4�ʂMN�~���-��U�6c(���9Ze���'^�t�Q�[���`����[�u,�(�Q׸�3v�aFs��%�uQ��NO�:֝p�;����RK� 4S�d��(�4���m.�4����)�?1$��y9�A4�I���\��F�d�Q���+����㏹��
�/���gX��D�3�]��LQZ�ޟ],��W9��"���ϊ����sU^�BS�l�yf��R�MU��)3�%�U���E���~���S�1KV� �"E$�50�'���|�4^uSd�e��l�Cۓ�D�CR�/Jk0t*4H�8�����<+(^�}c*�b�@r\����LiЏ1)��}Y�
D�w�m�]2�N��~XT�~�ƭ�r���V�5�)�eG�_/I���E��~�?�/`�RB���k9��*�J�3�#�1Bu�܂�/S�m���R�5Y (jKQ��Ueb&;�Q+C�.;K�f�T`���$&����}��'O�
�G�ń1T�5��0�u���?�ݲ�o�.��Hɇ�t����h��S-�8��%��'��>���A:)��sb	����]6��Ii�ٵN�ɢ~8�f��+�z��X&��_[�U��#8-32ݻ���n�s�S� V���jR��-3�u�W��QwnE����^1��]z�����#	�jj�Յ�f�y ���(�xL�?3�$� ��Z"6S`�J3!o����Q�N�G����߽�w�מ#�
"'���Ձ��F��==�<\��z�6o�(��}�(�\Ia���~��z�xm�G��N���9{nq	V����+�<o���Ο��@/(K}������MC����&��MomyM�U[��8X녏#s=aJ_5�h��2"�B�"KJЅb.K�	���T'R���!�f���v���oc��AS���fQ�U�;��
�����%-dmD�W�D"�X��ї�C���e{��K�a�-��*��u��ze�U��1�]/���s��d&�H�ڸ^n�*US�R2�J*o��9�'9�"F�%DJ��ѹ5r�9��P�+k�lI��Y���ї�ĺiM��Nf<�� i'S��m#4�b�-gh5f+��}�~:%�3s�C�~��`!��j^���6�a����\=�}D(oJ�1rͱ�7�ֳ"ڜ��q�d�p� *M3q'���.د�n���*W��a�$,�Dt#��m:1��qNZ���<j��m�24Q���=�Ҷ�~`<�����L� ʧ@��nCW&6*���,��k��N�q"B��2n��ryR/�N�Jm(=4�:RY@�Rdp;��]���8�|��2 .�r�Q�o����-�'u��;"7��t�G]w�$������7���5�%����1#�E@U�z<!\�^K�s1�U�hݢ�*��޾⛟��s�(�X(co�[�*�ro湞��:�a���&htD�&2���(���Ũ��-��T��
�ަ�!H�P�ϔAka�"�*|`�.��E�&~�|���l�T�Ǘȳ�w��ހ|�A�
,��~��,8�mb{�����aRGr25!:�X�dT�D��'_���ϛ��˪2܃�$�\قռ�U���c���.�8O0���*jb������=O�����Y��mOhj놫��a�����1;�L#I���u��Zv��O�"�\���xP4K���'+ی���� 6C�vQ��7�1���|~�=#!�*V�����A��w��Ύ_��f��1�/ʌa�+�����30��A�6�>,�IKj�F�yZ��&LG���g;G�&��I*ǽ��S�Z�FC^̱�n�b��^�jOm�+�w�j��
�чqB������(#0�|f�YԶz�<>kp�}�Ԋ������n��c�Y�VN�e�ms�*drP�V�۟z���6��IZ|��&��>���8:۩�������7���E�"؁&�`��I�7���/X�vEJo����%n5t�-_�m������e$u�5U�� ��q����Y��F;\�&�ᾈq�M4�����8\+��8,}}س`щj@����-#~���q�EF�/蓼w�OCR̛W�Ql������?R��]�L=q���đ�ϝ�yg<���j4���B-&�Ou%;5�ӬXp(\F��$���ݶI�|�ro�ֺ>JfV�́��W�>=0C�/E�L]��!e��͊=>V�Y�Q�2k�X��]�f7���$L���y�Z��������T}�Kh�7-|)Y�m�ik:_SB����u�!�DoN�'b��uFM@���?}X����U����QpTa�ڴO�k��)(P74����p[ΦЦ�mkI-��Z��=r]h�(��#B�Ƴ_�;p�
�?�N���i>��C�x��O�v�Ŗ�-P���~>s�~l�����`:X�� ��p1�K�l�����똫aG���>݈K�ʤ[�
7l���q�w��e��U�&�Ó�����x�U#2�W0hUW,�t0�f�5�EFM$��;�X����0(�1FuhP&�cd����Y��-���oK��j7��9�"IW�V���5߭�0�N�4����&���1��'�w�ʇ]��%c�;�Ej�~�t�1ݮ��A7>E�������8 V6�MT���w�Տ�,`E��l��,���M����[=I���=����,y� d�6��-�H������X���Â���[rZii����r[e�Ʊ8�M�(��:L7|!hlJ�fլD�����sὮ�/7��ܲ�h3h{��"X]�X�"�v)�k^�p�
Pk�Pp��A θ���$?X&�h�or�4��S�a�	P���Q��t�S3=7y�/��䴎&D<?/���_�?0���	ݕ.аJYMB	�n�[kX��{��K�{�QMw�!C�[۷O�E:�V�����[GH�f�dk�Xn�8�P�/�k��� �c=���h�N��,V��z6��R�A��e�7Ñsc<����� B���]�lM�T�e�n��݂	�Z���@����;+x���_�	K����	�祝���3%2Tv���Ct���$���G�^̉�cr5L�Q�Y�P�#�L��!1EZ�Bl�a��<���jR�K��x>�'C0p"�ʠr���3꿕��'w�5%x��ߊV5t7R|P����N�ʸHy��!����$��:	��Z� >z�gi�55 8��B��T�$�JM�_��d�����7-.��	a���D��2�(x��-!q��ֹ� �A��.�s���n~
B8+�T��\�DN��S��l4��gë�z]MB�i�'�g�Wj\��������O�
��Hn��3��x�Y���pR%H��<c'\3�ɇ�К����%�}�M��G����a�_D����E"�O��h_���#��r�S�;�w��a��� �*��S��g���,Ϭڋ�A��7��%���<�K޻�K��D�W|�~�7�>�a��a��v���ţS ��斧����[�4I2��njU���H�K�jk����4�����P\�t�;���S�5�x�b]�7ç3�t6�/f��v�փ���F#���iq��Wk�2�a�<]�w��3Y��]�� ���9����`sO��Ӹ
W�JЗzO�>��]�ZI�$�d��B���)ӭ�b[���T�H'�J�A+p��tߧ�w>P<\������B�k� �Y���ܓ��)�`U�wɄk���h���T�����f�Ģ��)3�5j�,��A� h�K���6�'yc�5ǎW=�C�[Ƨk�bl���r`c`|t���� �W{����_�������N���^�`�t��W ���%�^�2N.I����ѕ0��kn礊��P,|7���)�V� *	RI�(�����"xf�jmXX�,I��x�-�;�F�'}|�(�]����[�e�_���+��}����N�+Ѧ���
`CQ�,#$� Uu�w�m�h��M�~e�i�eN��64L�$���̕�J�^�@ÃᑜH��N��rt楩|�� �A��A���Ȝ���Ѽ�wbO��^\��BlDP?,��]�T ;��/_�ڸ��e��Fݰ$e�?�FށPQ���2*?��_J��*k�R�lZ�$���m��A͸�7^��EMϢ؉�dE��MjEO���=��*�V.,N���Ҡx�<������"�WE�HC>mT ����K~�J��QphX���%����f�j��k�S��z_q��b*P��� Ait�[SZ#5�:-z6�����1@�y�2`2cJ*9�9G��c������t�+�3Oz�
GQT3�v	De۪�d>QH���96Ƥ�y���7n������[H�)�^ WV_�ٕ��^���|~�?f"<;��z�w/�~�^�ɪA-Mڗ�G��\�F��ڹ�|�W�&T�L���V�ns?���L�
l53��W2(�ǇjI�G!@w	B�����Ð���ڑ]�4���%���a�N�MK���`��tӖN�R�=2O;�^�;HxZ>Km��Dl^
�1&���f���EBifcF�*ᒗ�=���P��Y���cq�	j󮦾	S�1b�b<���;8i#���bi�r��ӶSn�CI�93���Ĩ+�qF��gIDڣ�&�����5�#�� ��k-U�G�NA�f�|�R����Zl�G	�+�e��E� Sa_=O�r���o���FYs�`kC��	'P
S�
�S��ޣ�Ad���)uh�4��A@�Q�N�؎{�pÙ�}����	|w6����"?��S&�Y}l�&�䉹�#3I�ǈ\sS�;�kn��1(��qA��n3����A㛳8B�0��sx4�kRW�����:\;�DX?�f���V�>���K.���X!n�����*s�Ӌ��@�lmh♭2ĀAe����f�K?�+2 ��/&�[���Bɉ�jз�bq�m��{M$Rc��@�Z�b�[l��y}BV���S�]r��ۊ&wp��G�G��'v\7m�`ڰC�/��dӼ�
�S=���M�`hK�`-h��Un�=4�%O���(E�-���p@�x��2���?�A��΋�<0D�K3�|��Jۄ�4I�<A,IsŔ�V8M�Y#�p���`�P������5�W<��>����oc�.�~�#鉺��D�ߒS�����$�0����)@Fb���#$��X��1�z�M\����N
�ٚ�L��wJ�k���&��?�eU��t��Ʌ�j%�B�����7JP@��Ql_�Y���=��0�p��z`iDd�C�YI�u9�JqjJ��x����'r���� �-���|��Qomo
J�t*���Bv,�R�b�D�@/p~њ�\I�2�����s�(\�����$�Z����T��5�y俹�me����]Ԃy�$���:C����蚐_�[A���9��fGJ�`h�ұ,�4_��R��;���x/�EF�|�A6E�;Q� ŷ�pF���:�E��!p;����>�|T�F�~_j��j|%/��m4�X�a����Jc&2o��f׳TU�lAԯ?��3��ő�/p5�Ic�g�A���N*�����
����{��=����E�k�'1n���8�RR��{�!�%�Y��P�j��)���HzX�xb�SؤUƻ�|���WJ�]MB��2{
_����D�ů,���b�B&O��W�@��&�U%�5�sH� (�p�ڤ�\fs�!������A⨀�^C�GqΡ$C�VH8>�e*��P=�[�[<,�>�1���.�H D�)�*r*FY� �t���u�*�("ү��8^�7�\�
��j/y=0"�a����[�Jk���0��̱!c�K\���0ﴕzC�8.ꜽ歀�Kl9��N��Q�-�J��sZ���9��?��?iQ�A�;��]캀�~?����}�wM����Y�={~F|v٤.��q�� �R����y0<a��U]E �$)�'p҇�y�/��@�C�����=a�_\W�(���-<o���K�ڡV��3%~����0ή7vO��$.ajrwW��	�i�e()X�8Ψ=ᎸHZ�)tPKS4�R�
�=�D떗0�=����4Z�y��t�"ռQ�[�k�\�V?|�&��2Z��6Q�m�7_̐4��l��㵠��l֭�;^��`b�������:�r�;3c<�澉�25�
kZp�]7�g_Ej���s���Y��F���VᑤEo��KQ^�:�;�D�TSc�穨.mdrgˉ�j�ɶ����`d���ȁ��� �2f�/&��@ʾ�����i��	�$R�"���bӕ�veB!�v"�9�5TsQ
���cg�� f�7iR金��-�dxם������Z���G`���F_op	����_��g&�P�Z%����e�D�]���D���!�䟅����*���i���>��V�`5����-�[>�\m��HP�`s��Z{�%�di~6���i)�*X�#�_�ì��:w�h����~mm�T���y_r>tj��=�<<D��Ŭ�k����h�O��A�3����X�B�&*ͣ�ãƜ63����k�f��s���_����s�aǫ�B�?C��a���(�~�U��*�H\A%��������]�)�d@^p�H�@	��m�pn,R�L�񬁋�_�CuR����:�.2��>1�NJT�r�#t`�W`O�Ĝ������mK�h ?z�$Ab_�U�$���V�0��,�
�6z�99�ʫ[>N�v�ߗ���lL�άE6+
�&a�G�Bs�`Ʊ�D%q}qFX�TT{�"*t���x�Ē��z٤�@��<��G=5����ə��Y����R��%��'n�c����CW�x\|��s��p�Qge���Y%������dT��z��%�.٧�u�T����?����V���K�$�����׳/�@��M8xv�'ӵJ>�=S��Y��,���J�'��Ѳ [f������.��9���)�La��jU�����T����e6[|���H����M�����9B*��9훈Xu�8q�e-�J��T��*��ts37��;T�`ҟ¨	� ^���vcu)%�㎾0M:~��:A�#���T��<;MT:�K������y����>��w����Уi�+:SW�\���׽G�3���S
,tŁ��BJ8.��5����D`�Y�����|�	�`����mB�{Y�2�xh7�*��'�/$�3F�UL����@ 0aM�aa�84�q֕��;��s�Bz+�9 ��X�:^,P���Ō�*�RԵˠ�lD���Х�U�4*��9D�+�i9�ߥ�V�@s���n�(�{�L(��!�h��/=�p�Z��f����^/BڶՏi楴%;��l�b-{��7Y�>
Bg_�2l�� �5?_���Ja��T���a� "`��P��9B}�����C���e�xK����J�����h��	ˍ�Q��Q1�,��CE�Գ~�d��=b;<����o��� �W��RˠU �MPq�K�#��En���N{�X(N�u9��M�|6�oҿ��|�#<l�v0�t)��4����˨ت��5(5@�6�S87�+�>z�����o���Xf����,����R�lO*;�u#���ѩ�_9nr|�:^h�\B8,�VuG�IR��~���6����զ�]��{��J��l�����cq+�Xg����i�H4�ek�asg�/x��\��%����ⅺ�Aq
:D6�����*U���ڈ���ћJF1��L�A��n����OGO^x�j �����=v6��3���)�$e���
;�	���(Ҍ'o��!�)��O/�(	�1����7���j�b��6ұ�sPe1��\)^'��5�!R�-Yb����;������/W���sH�|쾩ր�U����h��RB������5dBJ*	��1��'xx���B�:HM�j��sN�oh��d�O-��+�U�]&�!�����}#�Ԭ�
E������_��d�Sr<I?Nr�X 2�O���p��t��\j��xM�3&�G�1�<�nG|Q��D#�_A���;p.�KJҩY��\���?�t���S?�Z6��J�7O��}�qFB� KՓ�u̴����i��ҍɂ_� u��ʔ�"7�<$�al	�WA\ˠ��(��?3j9���:�H�c��`�e���>��i�dӼCi&r��4V��&upKR�J=wa�C����X�O��#RA�≶z�W��<y@	</�D��%"!t�PL	V����Tǣ���X^�v����h"��)�[H�o8{tʙS�L���(g�[_Jv����5SQ�A�G�4X)�[Lr��=Ū���]<^�T���@^kxK\'(����ZQ8|.�����?���=;!�h^�T-7��i�K�RJ������'�U���_d{��񈩵�4`��WT�z]|.����l��Ɣ�AxU�лQ�/qj�a�3`ŝ�/�<�?�`o��x����)��>z�[%�i�d�q���D�\�h�+�@�r�k�>�.�2r�/��һ ;��	�Q��n���ۈ���V�n�u�fK~r������3���Ơ�[W�O]��Z�dd�4�>I�u�:^TZp�iN2�W�������g�iOٳ��n��ⶔ4M�3glL�3��b�o�yh���S۲�91r�'�q��u��<���v@X�g
���v'�k5�����g��m���:����>6_Q.��1�����I ��������Iy���-k򾚾�i����ɐ��1�[�uM�a
��9�",'-�7R/u� �C-��fͶ{"F1C0�HuFA���;�pƗ�#Y���!�Ԝnԉן����1@�Q�3^�x�A�8����H�����k�Q���$��㧞(�@S��p��l|f��ՇN4�-~��]_gRM	1�SQ�g�u4a�ĝ���<Z��GT'*&����F �F�/h� 9p������/ ��F�q�*!�W(��3��v\]�����t�jX׉�gX��C��[R���.�L��#1�gť�^�uԈN�
�7����փ����xP�O���(���Fu�w��f�P�r����muA�]�S���RV��D��U;�<�HW�dL5H��Bs+}V#��C;�f�6d����~�@�Ahl@%i?�^���Wog�e|
S���k���w׻/���-�1�2A�8��� @ 81�UEx�12V�Vvno�J/���l]���Չ�%{�A�2����&'������]vlW�������FZ%%�O1�-��Гa��K߈8����7�M-��j���GS;3�D��v)��ە��yږR��M��p"
��q� ������F��R�2�Ȥ�.�YhMtuXH��c�VF9���4Α��F�u��cel�X�����U���X����g��9B�b�H+�����nv�i��7�|�*�������~z$t�H֚�#�>��%�i��R�
�ߧ�������
�JN"t,ƽ%�Kn�v�N߀�vc�a���F�������]wG��.f,v��~7�q���H�F�~�z�-�w �Z��o��DS�	N���@��^A@K�[�Sk~�:cv�H��|�Z�b�T��������k�b��'��ߦv���4�1Epp�!� 4(�r*x���W`ӲIN~�{8�iq͊$�2\Z�Ӄ\lM�*5&!z�Rwɭ:AxC��)!%�(��v��vQUB�'"ʀ��/�U���s�e�eK�{?�Yj���Qq����g���D*�/E4w���ya��Q�i(���۠�#�q�G�|�E�:���Ěl3��K�@����oD�0��WZ�e(�Z�~�򊓴K}T�]�FZ�:yW�G$�+��H�k�8Pݱ��*;t�ổ�|��r�|�+Iy	��6ϓH�z�T:����9�/�(�Ϥ�<�e��'��b4��8���V/�Z�f���<�eU�N;<�ϡ������1?w'���[���ƈ!?�xi-��\ʧ�d^y�?�1�X�r���2SW<�C�\+b�`�����[4�X�4�痔m$>r͈U��{��z�����8�&^��34������ ��g[��n�bx�Y�H��.~]�x�@m�>sX���
T\����1\�ʇ#���P~&r�Bfb�ߧ�%YWzpL��C�p�j�z0��Δi����"A:gp0�krHӌ4��,>,�|T�C9$�&q߿�vB>E�K���M��𱤙<4BN����l:m`��)M�*����dWs�k7���ˁٖ@t1�����C<4�ͣacA�Y��N��:��>=���P!�9���}����S�1��`�	�h�w���+�GQ*,�#���W� W����DYl���?��g���fI�j��iB
��� j�Q�ն7�Pݚ� ��?.�-1�Ac�O�?�P�eb~[q׍
�^
^��絉 ��g��2��]�n�iOe�<ш�D(������>�ʳWY���B�99ֈF�1��N?y����z#У*.��8~ѧ��s1����DB�(� '��I`��(�?�s� s`bP�9��W)���N�����!��j��m��/�~�4��h��rI�TbD����[_�P����q�����O��s�b����d:A!gӄ(����З/LB~Q~7��p�D�:�hk�XC�В7��;�1��>�,p��"�O��&oo�����h���1���j�
8"h��͘�M�_�&�a�N>��B���=��O��v�q�~}��XgU}8#tL����چ�}"@]��;�o=�;���YB��N�\ȷ�lH���'�U<�$�Rw�������5��֮�o����Pr�N�1>�b������������"�31�҇�C�|/��ʀ�������*S&�!��=U���ӫ��sb��B���D!�Am�P-!�?�˾�E���5��jH'��f5����,C�K�b	�)z��n:�'O;<e)[��6?0�lj�@ŕ3��xD�B=�ܭLU�t?�:f�����
g���w����V H ���I���:S�vE�C�ퟸK�R�v��lUa��SyJ��ne����[H�<éV�5����+�=���f��gQ�x�d}W�E����n ^���-���r�L�Z"�ǧw
�&�U��O��j#�HW�u)����k'��nbD����F�B�9ы��a�&�B��-��ՠ����uz����\h3�)"���bgh��?��
F���a���xru7Z[!��yE�<J��Oв�NF�
���JtiN(�2�`��� �l�R1�O/�����Z��)�qj���zq&�o��ocQ�y�'!e��l��K�H��|.W�c�{�^�n$R��>$P8K���R�u�;*��wbx6�J���;���m�J��*3��5�
GB@Y�I�5(���3���a}9N2�xN%*rZ�����:��ŋ�U��E�H��]�зWV_{�/����2^20� �}JZn�~G1L�7z�����6|���|�[��H�4���.�r���֑��-1gc�T��
3\��!���S������biU�o�J�2r�jg�)���!�3�{��<��r?���"�������j��긁��,׺ ����`��Aü�oZ�o�ś�;D@�g��
 *\�l&`�Ol$H?M4v����2�,aݏ$Y*f���E��ϊ�:�Kξ� �ۚ�u�|�{�O=�^�j(���Vi70��% ��:P9�A��y�ZG-��>W��BV8�x^ 0�r��B #�~uA7�BI��3�X��)��YlWz��G�i_�Ox��:Ll�c�WP�c{��H����,�4�-��B-�^!"*z�|1��b�:Ҙ-���UP�PT��O3^b�̃m���urCl<�n�(��y�c�<Z.�0����.�͂�zS�=�X��C_���C���s�,���HU�˼�d�yb�/��O�VvƓ�1����$�*$�;[3j�$f��x��&j.`o�l�0�R0� ���ڮ�"���:�0v�
n���-���)��n$�BI������!�������!���ݙ�WD�|�����Xx3j��7oWB��<|5���;���{er�0���0��k��ӓ6K��H�;.K4|W1����M��!Z�%���nF\4K#x�F^>� ��~ڰ_�9}���"�{C��}~��"�-�w�ng��,�k���Nz�&���u~���a:�Ozّ���Jà����MJBB�m�Vg����m����@nB(�ֳ�#E�s0���B��9$�A+����C"�Jȁ��]���*�_�� <��i������̗?+D"�b�B�K^Ф��yxWǿJ���
Lj��	E��tNL%�C�<� �V����}U,i��jrpF���[���8	�Ni�3P"@���PHgrm�=�?�����<+B�n�6�ԧp�7�b�L\�΋�:|�S*��D�b����+��J�j]�E"Do2�'�_��Q<���lh`L}�^�q
D�Q�Ƿ���ju]�!��7^�n�(�1IP���=��z{�Hq!#uE"m���˧m�&*8��b����a��t�~�Kz`�_�So2��6��D3|���׸g���:0|,�Ү�����{�l���y@aZt����մ��x=�������d���<z�(q T��FԹ�SA�=U�Q��β�@b(CK{�`7lE^H����eHG��c���(5�b"����-�4��y�N���uT�TCn���O$Cշ���"���C�0p�w�Q�4�4�v�#@�G(�
y�en.�����V�Nשv��&\�VŰa�:�8�C ���>;����q2ᶑ>��.�O�mF��ex�/{�O��� g.�l̼��a�k

iͿY
�L���7Bu3��ģ�ٰ���׏'	kF�`�<�9~����yh�E��o=����5�ڲ��J�Q��PJn<	��p"���½�vT"��g���7��A��HR����w�lb@�k��J)l����k�֭�@��卦uX��,!jl"z���_�"����[s��F�X���ڻ��_��Чa#-}|���$EB�:��IYQ�f����jl.��7X��\<��|���q�c����U){,���ڸ��:Fv5 R"�-�3��+K�_�����U�c�f���r(���[�I:_7��q��I��ؾ�#�YU��	[.�{&F Z-�^
DL-�i�������͎�n�-��D;�b��/i����eLv8��%��6Î�����7�R������J��3d���\��:�e���'K���r�u #�E?�*�_�<5����ߦ��$S*E��MjO�(���i�c����hZ��Vѷc�wRa5��@Z���,K�rg�Dߴ3��=�h�����h݃Q���с��ֵ���N�#�3���ora�R��K,y�o�`��-ً�5���"\%@ ��Ӫ�;ǥȠ�2�-�8ߧ�Hʠ��E�.�B3W�"`˙�b���P�S]������L��B�q[���=gB�pq����ڛ�q�f��K��3-!/O1E�HLՌ��×�DБ@!���՝��{[�-C}��l�u�Bc��[f �h~��ʼ��k�C9M^S���5^y�+5��e��[EE��N4A2�u=��Mf�X��?$�k� �H���m�ϑ��՚��N@FB]Q�iOt��ٷƾ�O~p��Ǉ���Qo�V ���;t�L�6�ORP��N� [�����{a���<�?�� 0�� KA��w�c�^�%T�|�<�A���;��4��c����Z?c5$l?��ҩ\7妬��f�����P!��WΝ\�#�e�I�C;�����:�Ju#��tR=�?�i��o�z��=v^����߱)P���;���h���T��8�A�R��ҏ��A�;I�SS"�����:J�E!�w%�|�:Y�S;v�
���`
������
(X�_�e_h3m?=n��K6�Z��yI�6~^�L�碯�?Y�۽I�X����B�@��YA�@Y ��4i+c�5�|�+y������?��^��,������5��j�1;��J�*������ ��S�Dj&J<���̋�7+��s�l�k����Tl�[g�]:�)K��^jnk�S>��Ҝl����馂C��r��vf���c�2�Hc� r��3Pr�Y�/�#7��*kqzE���.^ ��ͭ��y���4�z�ˊIov;'�nQ���#�uߡ'������,�N��� ���q)c4M�ʚu��Q�xǸq2"�c��ՠ9E��߉��81�ƴγ������oJ[j��D*�
We�R_�����C��]��x �Bj�_�7a�^3Lq�u��AY���QgK�%i �`�w`qY&�V���~x`�������9��h��Xx���Qk/�J����H"�D�}0��x���3j�w���P�}���w����נ�����	�$ݎ!��Xo�nΤ0��aN����v�[!ÆA��:��_K��*W��j2W� �u�Q�ʸ��e�_��;W��x��?��`����/ �<�.x��l��o����g�:�w���Q7�I�0tܲ���peR M�C$[�Kq���;��t�l��;KI�j��������� �vp�0�� B|�a��A/�ڡ���O�l����*�\��4vZ��*��-��LbIנ2��w��6�C�H~=*��~F�&�'|�E�N7(}�T�F�fr��t��k6m�k?{)��Lo��1�0��e�>��~���l~e�@:A	 N������ҍ�bF�C&���)r1�Z��o��k��KP�_��F�����Z 3� ;6O��R�{}�vĒ�����J5����Lʈy�S�؁�l%,U�i�[ζ~WP�a+������l�a��=�L�=#���Q�B��Q��\D��ۦjnPG������%p�~����K���.b��t
	���SGҰ|H��d�eLQ�A�����)ψR\[PV���a�5��?��iώ��
t�T���5Թ>=H�<UtI�b�+��*Éژ�Z"�J��YGC�cUJZ�F���{�%�J�J��}��J�p>KPr�����(X����� �^=�����}v40ë�LH�[	(݃:V�T��7�\G�,_��:�ˍ }'��	[�ڟ�JGY�W �a	
�e1{}�O�i��h�G��<W }�Eٱ`C vږ�"|�N�Ͳ�4S�?R�o��G�N�~ ��\Xu�?����#z�o�8|R�m��EMU�&�ݎ�n�u$��8���k����f�MFvo���wiIV$D�_���&wP.��-�Ӿ�TjU9��F[��f\,�m8yH���B�� Bh��@jZt @��� ��NԜ�����9r/s���2�l�� �7�(��>}��O�,��eo`�_~yS�<}iJ�����`� �|J�S���|Α�-a���Wkf_��re��c��xHo�ۮK��V5�]-d��d��:�Y�r�\�{�:nI�6�s^����D�F���w��i���#e�,���s�i�+��׼C�wѐF
uU2�������0=�X���%D�Bx������xu���W�5(M_[e�
�_�)	̄C5��ys��u�vDb�d/��# ���d h�V%Mf�t�cg2Bn��XH���ZA���0H*�B�D��u&ZG��Xx3۷���dS���d�mϥYZ��"��
U�/D��#�oA����Ѕt�1Y����~�)ڍ	�#r֫Q4��SV���H�[��x	0�#<���B-�B�CT����F�g�N1�faJ���
N�r;%�v�U[�P.����6|�����я��h�.$����������������84H.����t��-k/���/c�|���ہ�y:EH�R%�rBa��l��E-�}�S7,p7�������+�槏�\JZS�� E��Ga���QC5����,��O
Xl�UҤ�O����妊��BL�^>��(-&�9��fHw\�SP:�J�oU�m%��<��<c����b)&н��qm�M̙����⹳����M૜e��'�
��Ԛ��XM�ђ<G�C����t�9�d���5Wya��s:kU-2���k;7 ������<N�ΰ�9 �u4�/��+�+�Sxb?f���>_דo��(�ۥP0��s<�8�P=��Su;�SE�qOL���"E�Q��ȱJ<h˾�ٛ��%�w���1G��&Y��]��`�|\ �g%9#��͎ ����kk��6���������f�sCF����Te�b��g��d֛�Y���0�S�8"��
d.���@��By����/j�U4e�¢#����Hn#]���`P�w[�z5_��,aW&JȌ>@A��wT���|ިҏ��P�~��S2ѡS���g.��`r�WC8�߮%��c���z�B�p��	6�y1Lt�N�$xew]R$?A�1��~�&�z8���i�L�.�[R�7r:"�)�i�Ӌq���̸�B^�J�)��1��h:�Q"Lы~�99�n��>  �]��G��K�5<��9����!�|�Zk�\Q���<�-*����N�q�%aR�����+�����������*z���k��U�ʌ�����y6#D`k�I�V�DCy� T� �v��Х��m W�+W����9;6r|j�Ca�ǎzg@Z@X����6&�+�2���)3֌	>o�|2!�<�*����!}u�<G���`)j���ů�7=�w1S4�]Fj~���6ֻ-�Sم�)?����$SK���/�ݙ6�@ͼ���ԡ;�t�"lj�`㋋���T��+Y����=ؔ�|b�z�p���qOp-&�j
2���d#,_��>��k�ߍQc<G���lW�j���kkL�ȽB��1�+�[�Y=�e{�O;�t�;���� 2�֙O
��-��'3�F�d�ܠ� �[%�Ca^a����4���j�*�~]2�8�:?��ӿ���Do2�4�&��2@� �:�n)�<���;l3������?��ץ(���oy0�u����=�����A>Wج�(�Jr	�$p��� ��g�Bc�OV�v��tU���	��
��\h��6��?��3A�(�k-Nۭf�~"�v��@�C�����)����Y
�ubC�ԋԩT�.�7z>���!��'w�qj	i�6�	�T�O�,�y�׫^GS>��m5�����~��C&��a�u�X�%�����[SO"���Q\7N|a5���g�,Cjn�近�j
����ٿ�\é"���n�O��7�w'7��J�@�}9���a�D�1-ҳ�o�m_� Ê�ZR��h�#��#�"�;�����9	�SB�\�,����L��Ր��e�
�j�o��$�6�{P.�\�F5� @���E*�s�` ����$e�����Y�	���iVwƮs}�s�RY��>	�)�c0���Di!�K�Z��e�溲�>����x�`��ޯ��n����8�S��G� *�XG�4�Fw��Lk�NC��]��swa9�W��!rt�:��̲w3P=b:B�KI�#��g��zCL���ץ،���C	�$ ��PNK��މ�aҲ�|f���Ȃ�"0p�0��;�ʬ#F��]kKҚU�[�|~^�e��8�z>�Y�z6X�[��+���|%����5��'m�	���nW���D�ǳ/	iO�?P��l��P1�\���K��2�z��yQ��5�K����iVm	��ݍ�0�j�j��FJ�H�O�^D���0 7L�sY ��1V N[S-��	G.FȊ���>V%���ơ�IC���Kb�5?곮}3���׭��9�b���񗂵b��fL�(	�4+����ɤe
n!�9�#v�6b?ݰ�0{�����r5��uQ�I<��u��q/�P�6853s�Z?��������G����ˀ8����Ha��䀊��.���B���`��\\��Az����=�֕32�#�Mv�W�x)����B�P��0���[�����e x(�������^I��&6�ʾ��[��ǝhN8q�/�����ё��w��F~τ��{�	iON�eΧW�+��-��Y�=J�o�{X��2yrL��
\u5���r5qItJ�yժ��|C��f0��-O�^���*�5
~��R�u����p�K��wg�JvD�>8����#ݳ��3��?��߲peN�S�fF��'�����b�s��VS�_���Aej����$IE8l^���c�٦?�e����t�J�D���Y�NV�1�<��_�;��;(���A�P��;.��m�QA�յ���Y�Jn,NW�-f_*�+�n\��OB�&��V��45���O�M_k�8Lq���Un:��)M/�]2�K��w�����dR���n����T7dM�e���+����UՑI�[~hyb�;Y�nט��Bc��ӪB�V�h����u���{�����Z�������� ���s�߂�x����@׵#C�5=]aa
��W��p�DV@�j�_n���W;�xz� �n^�~�:\�I�����Z�ॏ;JPˍ|X�R�`w0��<�\���5���eЎ�<�u�mp"�j�~��h���LDM(��B��0�>�������{p��/�j���a[G����0|�3�z���st�S�˴�b���hYRbU��F��7��$���\t�~�scn���mkzZ�l˘W⃇Z�@��:�o�Nq\=Rm��h'����AP �*\N%��B���4�yn�>6����(�C���਋����qD�R�yY����Z�u����szd䦘s������鶛��2m��Z����޲ �8S�-N�)��lml��޺%���
<�ɳ�Y|
�,[���߽���G��]ʑ? b���,B��.f��Z}�$}�1�X����Hv����x�e^���H���(���F���$��u�e���Ϲf9
כֿ��P�d��+h���̉�7�A�����2��[����C�4��q���EoM�)�~�y�E�MY��m���Re�H����3A���.򿅢�h-�����!�����Q �����Y��X�U #>�L�>�'/��:c��U\��o�o5&C�5�s�
�읊�2\-&��yB���T���5$�zgI`�y�H�Q��]z�$�P��HхF����=is��\R���x�DUEdJ��x�EWGVt_��7aw�ޤ��%Z�N�U�����'%#o9+4�m���L}cx9���:�~i�� 1<�r�3��e�|IΚ\s�෺��@���Ѐ���y�8�ZwW�XmV�YT���(��a �g&����k�ɼys���i� b��{�_�*�;��4.=�R��l�8.�0�3�~c�V�2�}�+��h�(%�X���M��X��.���ǜ `���A2����O�7��޿�ۊ�������>|A#+{�E-����Hq>�����',�P���q"��Tf�]�hN���<*�g��VܔhOG�����Z�7����Y�n
��`,�'E�u��:N��%�����I*1P�_��J�`���X8������FЗ��!rQS5�f$:������N��ӊ�n2%������e>RFU,�ʽ�P)p{�������&�6y%�����"��5n����k%��r=�0A9�|Füsa&�\J�j�Us���$y��eqJ�;6��~�Ɲ'����Q���2-��2Ԁ$GQ�r7R�B�4=D5�� �~ԫ����|�O�v���b�gde��{����f:������E�����Ri��	��I�^m�7�s������S��z��/?e(TjS] �v�0���?ᅲAw�s![��E���T��Aޝ�b��մ�D#������F���b�6V蒬<2����K�m����ɫN�Z�0C�4��܀�;�����2 u�b��C��\�1bٟD���ו4�A�
5��Ѯ���k�l�M�;�H�8q��̌�6{`��'}Z{�9��ӻ�eg�|��e�NH#�wDqd�6y��@��*a&�X�����z�ʮe�ط`݄�Õ����׭�Sb�{ǄC�b��U��7n`�����?�MrSƧO1"���9l�����KX��у��f�^��!ʌ�lMI/=)�rdrĪ���)����}/�Z�C5F���%5C�aoT��+�͜x� 6��q/g�.8SФ�=�F��n^Gr��q�����E#�wO��ѵ�4V�� �rCK��N6�x��i�*��i �H�8�YϹ��J�La)�+�i<��h~�[�-����rES
�r�V��lW|���^�^�^a�e��}pZ�剣<]���X�vwe�M,��x �ܣzy�r���TX��ʳ ���2��7�ɝ������aP��z<�f�m��O4�7�Wv=a����r<��-�3��͑�����.�˫a�f�v�����Z���W���V��`��zr1������܇�g�>�q���WE�*y#��h1���/�ܙ Э
���pa*+�X-��BaE�4�<��XG9�@�Q[�t���m_����=�ز>����y�Ԡn���rL�e�~��~��������CG���;�"�G�#*Tf��>
�>��=e!�y"A�R��$�6��W�1�ô�U�%����?�C�i��\JXʇ�o�!W빋���h���������9�sw@~�aB��jp=ǿ6���յ�whhG�?|��䗝��J�)������zMp���=j����T���qv�z��nV�q���B�1�F��`�3�6�0�(-͝g°aetyL"u��s��o2��>�:��̈7k+Fy�R�~����f�N�!1�f8D��s�t��1l��~�V/2�8�ڌ�vWQ~�A�d��Q�*�PQ
���IjQ�Ip�"ܿ�鷶_y�XC���(���Ge�JcV��D]�c%������4NI�m�PC�� �=��`u��g^'���D�b/��������w`�ۡ�4�����rAjf ��I��pD�S����{�ցY.��
vD��=��-G���N��3����=zm��E�y��X?����+i�?E��O7UE�Ny�7f&Ԝ_� /M�	�s�v�vmH:ϺV%�u��ѣ���^�N�d:�RG-�XG�!�	[��oٛ��c�s6�ź_����.l�]�g�CvȔ�,�R��d�))=�I��ꁧ`������`Q$��V5�z��.ܚ�">q��x�Z�6���v�P��s/���f��`�P�R�4'ߠ�T���;��/�8`��C���UM���;i�'O�����O���=�C�mӱ����h���݊PI�Ao������r@05�Kv�B � ����Ɋ+�t�b<Q3l�����#�hؓ&ݐ�c���Wkf�\���t+�������d�7�O�5�h���Ug�FQ��<����Թ�� � �J��%�,=^�HrQ� �D�J�6�m!��F�͏�s�_y�(>z[����D��h�C�K��L��Jk�w�1L��1k�Ln)��V˙<Z�Q,�K���$���j�he�A*���,���j0m�ڤw�~l�r�5:G�(<a�������Xb`NX�ViNء��r �j 
�(^#Z��o�'܃o�o�R^�=	��h�/o<S�K�:vg���YpR���>�M���/��-��χ%� �ĵ�=Ob)��NR�;�<�U�W~֯E��"c�׍�ӆ_�)�#��y�B�E\��_���w�M�N�y�[+��YE�� =��4%��L�r���ɦXIff���F�gy���^� l�C?$���1����{����Лr�"��e:#�IH7v��"F��k�qŘ+���
�d���(��mcG��w�j���~����,*��W)z���N����O;�k �ǥC1]A���X��~eps`P0�Vaߑ[�7�2ztK��~�4����[�o<+�F�{.�C�|:TF~�&f2
d��8��]yxFp�V�2�'m�fI8;Z*��w�'b*����Tu펍@�<�����ܸ��08Z�'K�n�K(���*[4j� 3hPPa���d��Ј53�W��ݑ�
��5�#M�ٵ�&ֵ���e��I�aO��Qa����g�9^NPg�8�槑�԰����&�/B���8��3���u��Pp�zd����̃$��\�"c|�]5�v-���<�Y�~�Q���!��@6���yҎޱՂ	rl�O��O#���L�ƣ�Ӏ�+���R.��3��ڲn�D�l��-F�!M������[���k�_�r��Wr��0~�IziYxpI�[����(�?���#���2��
�
▲H�����_�O��2��{��zƃ*N��M��D�?�ƺ6lc�M��Í�8�]�,h�	�;�I�펄�)�o6�7]� ��g*������J�&O�!��d\�P��ٞ-�+��ď�Y$� ���)Au,�7�Ԑ*ӫ�8�j���a �?���<�ƒ���hA�\�*TF�[�:�y���h����@����B2�5k��vL@s�$i�|y4σ��F�Pހ��S�x������ ��<)�r*]�#�E �­ۢ�òKAt8��~9��q�[�G�ŇM'%`���MP�&��5�l��,D�e��]B��J���3�K��(�8Uh��rB��@r�9ڐ���򚒕p��ǿ��xY>�Li�h�S�:��I�ю�e�P&����ٍG�7�~	�"��U^��z�X;��.�W����?�����*~��j�s�L��uQ�����p�u$+��nEIC�@\�� zUj��Q�\ ��8�ὃA�*���_�m��>�'X�	r�e�@���8�P�:����_8҉�J���G��u�6���Q&&vK�LB(����!��3� �����f��)4�N��wWkf-�Q�U���wtB�����QLt޻dU���cdP�M2H���z�RV���Ȼ��
OfAwW�t�j�g��Ew�A4�^I��
��î�F���!5�I'�.3BGK׺P�mw��ǲ����*�T"���D���dr��_'�p��@
hNP�!j��60p��V�e�ܿK��d^ ���������sDKH��8?��
�4,p��s7��P�M����>�c�y8�ms����h�θw�,F��tȮYFnno�'���,ek��n����=�(@g�� �b�siX{r91l]�ܜ )f�DpT���3@V�ZR[G'DG����SQ��)�7w�������J�����q�`��7��h�*Qe.���$Q�ܰ yX-�U9fG��O*��Ev��� R<֫*|�&��x�h&﯑�\" ��!=8]�y��Iie�ՅW�8&������l�,����i!V���
j��`�:td��9�h���Լ����@s� dqN���@�x͔^LH���9~Lĵou�,��A	|;	X�K�f�<�tT�0�/@~~6 ��ƮR��P���#�z��1z�j�RC�J�x�!���K�f�}6��~H ,b�8	���ر ]st�	�Y%hT�^`ǩ<�6�=F�"ac���
��>)PlM��OƑ��AR�`(����"Cy5��Hv�X��" %��[~��e����d
��
����_�\z��aj�\��꼉Jf!C3�m��_V]v�~�)�@�8��\Ϡ�/��Cz��������|�����V	����Ȳ�c�,�Qł5��[���:U�Ŵp�L�o�-3"WL�[��\�5]�`(9`�Ѯ?(�8�x�T�f���)��37�L��v][�~�U�l��.���`t��P�!3��έ_d����'X-�CՑ��j$L����1)y5F��{7�y�h��R*h:�'+�.c?���M���"�2{������sդ�h�F)I����V��Z�.�˙��~8 }�2y+��(D�ZP�Y����h%��m4;P�埅�Q�k$, �ͩ!ZC�"	Lb���W��F��+ww�p�iN�Yi�8E}4�tP�{UiS�]��J[2M��;�þ�yp�����͊�p&�,�����-��"@��y�����=r J�d�5��yq��=����,ʵ��k��w��,t4&��x���Ľ�:A�0�X��VÙG{3��s$Ér���R�ii����Mq��$��)�c�_Xx���o6_�.h@��w����PlT ��@y%-�U{�c�}ǈN㐒��L����k�^o��>t���-���*�������Df�*\ �c���E�'���{$M^�)���`�7O���
_¶;m�yh����a5�6l��[|I���8���.?x��7�Ы��4@"G*-�*�/�$�J��j��M9�:D����O2�(q����9�g�ׄ�QN8���[a A�t�$/����f:Wu.a
'<���w-��8���O�EfD�T�Tc�S$1���v�A^L�g�K0��*������:�/L>�/���W%=��$�xXHU���;˹Jh~���_w�~� X�� 66� �x�6�87��=�V����w���*`+[��6[�\"�3Bdqd pQ�}��n��}Z��Y�y�H��إx�d��T�uL�ŲEJq��d�AMo#8=�u��%�<�:��V᳁
ec���g�e�h��Ra4�n�1�Pv�K�D9�������lY���so�P����!����ф�`0����!�/��y0���7Oem=�[	!��qB.�(+���6y��iw��_�T:)�o�f��&�x�w��h䷳�欮�-�hʞ��zLxC �>� "�3�Nx~SBݹ\��臃�i$��W� ���	)�{L��ۑ~,:�`�֖�g2"Hz/�JG���KL�\P�&�4�
�{�'�H�E��X�TUk�S�	r�x
��}-ӘrX[�\Ј��6�L�k�v�˗Y�;z���a[gp�vO)���D�*�فĺ��Ԙ�0l�qu�)6����˷+���H�=c�2. �m�:��d�A�7�ǹ�W����Y$uj��f��x �r�.(�4f�?��x���@ɊwڻY�mcV�U�^يvŏ�SL#+߈CR`�AW�q߁�����$�\�-(wv��ȴ^�[�m��)�����mW1�Ĥ�r�����%M�><� �#9�+����U6��`�>9�嘊�;줺�xK�h��şYڡ^���Dv�	hsq�rA��cs>E���e��st���A��q����*�Տ������j�T�f�g:�-^�a;'<�h`8�	������p|,h�.(p�75P?WP7T7w�9 �����u	����6B<T�|M����	H��~J� �^1��-�fP���w�q;3�x�cT�*�y$���� Y�Џ�19K��W|��y-�ȱy�I&n���v����L��!�f��2���zj����-vy�t2���h������d�Z��0�,��Ս0��*ݠ-x u��)�1W����� �)Қ���
���� ���
`b�I�BcH@oխ�0��������7f"��{���g�"���p�B`��7{[�&�HD�zFd;�Yէ���H�wlQ	{����.ʇ�.���Z�ɘ�M���^��?��Ö�@��MI�H�������e��d��c]�	�9kd�=;�Վ�p,2�бG������ ���P��!K�y���Ѡ�v�z�fO�������{L� /��Ͼ&�;Q����F��Lť׆3��9Y��jzqB'��t��(R?Iuϲw@f���|�szl��TjW����۵�x�� ^a&s&4#h�C-�(NCa�os� ���;�]q>�Fˇq��)�#p{ʸzC��;e�����ف+��!󈊛��*�BT7�G 謚!	ܼ�w���LL�jO����!V	�A� &����$WMS�'�a��9���V�9
C����6>1jW�y*7�W+�k�d�Uv#�G�t:���R�n�e"�m���T�0�FR*�Y��e[��o��ґN*Lwb��	e.̟ea���_�Տ��綩�&1�J��b�P�|nm7	^����͵��ꯥ!���R�ع�ip�����\ErM=m��� ['��is�Ѷ`r3K� u}p�Q$�7!̒u/��$���컗���E�y,�N��L�-��%w�
�	���w�[��ޟ(o����TB����ܫ'CZə~��Sc�t��>Y����I}��;`�e��t����^��=*~�� ��T\�� B�5�)�Z�ߍ���.�Kz�<��m�MκԼ9���=��67<����jq�Z�#��p�P$"k2j�A��D�g>G?p�v�]7��^�R�c�8��  
�ɰtoCȗ\T����rG���!��%��zQ&5y�F�����84\"ע�gi[M����|�&��4nF��ƹs�lʣ+!BáGs�~I�)�b��[�J:��{[!��&��ek˻>
M�O�52�R/��4���6��дPt?�T�C�1+�X����=SZ��5GېW&P�R���t��g���~�A����rH�A(r1����p��v��E����X�/#'^r��a�4����#��eI�WPv���WZ1��t��DˆZ/����)3��uHp� �0<��5�dM�e�c<�Ut�s'*��N��.�ob�|ό&gq9�@�_gn������5�}�t H���>{LZ�l��H�z�9��[3Z�%�l8=�PX_`b��A0��D1�.���Kա����ణ�(�[t��=���P���x��,�F�~Ց����c�d�5n���i���X(+�t���?����#1)E����������b{zʯ�����ҶZٜ�Ae�$~� �i�_ك�O�d�M�(-�����*c.@��W� #�a���O(x?���G@v�Yx%[�^��v���71��c Oyǡ��1���R�����8,xmb�`.y�֪q��Dn�P\0 ���\�����ifd��{�[
8E�yE<�S]e����i��ţE��^'1]�kp6;qxE|�N>,U�Ws\�
�
�"a[��$�v��E����� :��� t(;/�� ����6�-q���R��2�O�ϼLw�!���7K�-!�x��+RCEh�Us�I���W�_�s���h�|Ry�rx�ݙ��`r�T�-�����s4N��G�ܮ^��P�������+���`E^V����n�D,�����Ⱦ�����^_����W�{�����r_v�0��lv'<�
l�9a
-v�('�.��ؗu}� $SS`���0�/��?���n!W�?�&�a�ۃ]�M��y%0�I��$���I1P�ntT!ӄ�5X7�6��}�Y�ω�eU7Q����/'��bep>O�s�YJ���]����舻(@��oKQ)_�qT��Ϗ���]O���MQ3��3L�x��UYyX[��!�[t��T���1��Y���+	�ܧ�Ý�R�����L�˲�	�s�E泏�����]zI-rf+����H9˔X���S�JuG�(�^�Z�f"��;+���ӂηb��?�Nt�q�A��y��|����/**�ı�#�j=�kb�����������@��S�R��ec���U����:vb�S�Dq-���t�b�h�������U&8yc]	��毾'M^6;�E���I������a\������2tR���U*Lm7Y�s7n�u*��?�3��ꓧrAŌA		HPh����A8��W��Xsh���}�*��.��'�3� �k�?l�Y���A�Qh�d�pL�V�ՕQh�!�����-W�)�B�������E��h4�p-�k���Q"޻X�CUm������ Ȅ\x�����QV��r18?Ғ�.[�&��.��z��Q�wQF0W���leU�e��6�h\i<NS���t6����A���YYwh�s\�o:3� �*c����P�K���u�N�ˢH�K���f�*D�$�ߣq����>�+����J	�%����M3r�~���㦓�|۶IDƯ�6��v���nZ3�=l2���Q{p&?�Y(��w�!G@@��<����Mn�Ui<��ۡv�r����9�A{(���J���Lku{$��)����!1���̺�Pv�3���z�c����,M�2�N��o���
3�U�n�8N��*��4K�)%ƬeD$H�f��!,�Z���}�5|$|��bdfHG)��LDMiG��
��q�6,� �2�j��6�\��*��5��c��ϸC��dO�z�4~��d)<��@��DI�6U��J<�x���^��T Ic�gN���`��V!
�,���|
@\����ǹ	��X�ܪ����k���O�M�C�Iv_�[!��\�	�r�?�����O�31>m�ڬ����{RK����s��OϙWԠ�M�I�5д�;ཐ����XN&(s�m�$i���k��f��}�
��u��)g�l]j��/> N��@��	=��
V�˲��f�'����X�W��g�������e]sh��� d���\-&#�e�������O+T���ƧL�~'������(��/j�aI)���U�n}��{َ6����y��H�]B�b?K(�����E��1?����W�Y).������@~rBvw����毰��o��M����q>�]S��\)�"H��}<\>2�Hh�>�����F�-Q�'Ǝ9���$��e�����;f�7V@9�%g�d8�"3K��Tu��kŉ�0��s,g��.���;i��D29��ըk��sh��A�ա��?_XHO#��F`N�A��|9�]���$u���FԨa�}*��M��U fBW¤u��U4�d�Q�(��+�� =@cJ��2��C3���NMyP�k��x�iufk}/E0�ێ��#��+DǢGŉ#@�*wE���0c���yG��]��6��2ʇ���Rx��X�`��I���Z��P0@LH�1�F*#g�O�~6'Q�n�cW�U�S��4��41s,��;3j&�tKє�v�#�ȃb�� �."'/H{��;��}8J�^�R��|����*���v<W�P����n��E>w^�w����DJ�l���T���ƗY��`��)g1d����|~��a�
DBu��dGW��z�����r�o��T�rn����/����eb:�z��wтyi2�<�f�!$��ձN7�%Ҟ��o��?k��84ƀ���CH� |�)7��(��_	�$�m�T�׎ٮȖ��j��N_�H�g���C�	��0�N=�~�ُ�>�]-�8R�`�I��4��P��5R�������4G���uyQ���[�����օP���`� �����-p�
�Q��'��>�/��������C�w�O�|�=�G��e^�rW�d�B�~�'ܽ��PhN����:�,%�Rvs��5y�@����$Rgj�jƲ�{��R�?�ۖ��,���p��E��>�(Q9�z���� �xc>�{�-�Ê�\�W:���]6=��lƆ�|��'l�#a�����K�+���[\AQ�^�`c@�Q�3�Bq:r<�ȟ� �&'/� �z�N��}˿R�Xsje�ج��tAX}Ƈn(�a���� ����lb��_�c(E���tk�R�Y�����U��{�H
Q��$���dT �d�].bc#A��~�ō�c��Ź��ƙ�A\P^7B�{�r�o���?��V�e���p���!>6<�]���$Y{��sD1��TLNH62���+�amP�2v*�A1�)R��f(o
�n6X���VA~cG�4��6"̻/.>��ـ�`:��f;	
��-�d�d��PY��'�x��3�#f5\U���[&>�4~�Ep� �G�,B�(��b_�ը���ң��NMHƉ�U���:t
����� ^n@�L�a���WY����4 	@/��9�*P�Ԟ�����=��h�J���͔t�X�����7�cﲫ����&��"���7�-�Q*WR�
K'��<x�B�o,.�vS"׈T��0@HS�d�8��[��؟��zl^���C�iDt�e��+��.,9ߜ���$�ge��{ }jAsp��V��INy�i��T���HO���,��x�6e��o������mwSqA8/sH��]��._V�2�B��B�9U��l\PY�l@���D�Y�g�}�� <`������vI�o=�+�΍��	|��+I� ���W_*��B�� �����maȫ\��:h\��a����/�J�M�V(#�u�U�^`����b�3�FW��ׂ��23\x
ѡ�8^I�/�ĘRT�^� Z.�VgGu&i���Z�x��"�l�����ѡ ����r��BV��R�j��s��'ymF�r}��[	_;={>nc��
����K����������fT�u}<��m`��h��5Xڰ)���fҊ{��Rdc���_* ���ط�d��7��4Va+�_`�ԕ�����U��hs�˃���[F���@���\�N��Z?>�)�Qg.�U	h8����
Z)R�D��z,aV���> ���m:D��<ݴ�m��c<�d��"F�S'��z�_�BY8�}�/�n]�IyJ� �^��{�H�Gp�!6,~!���{*M5Mu��T}F��s՜��5�P�3O�����:G��u��$1�E��k�.i�����/�"�j�Z�*J�>TWV�m��o�u��1�š���f�Á��52+@#{3u݉���_�8�h*�i�&۱����XhenIAo�����o�Dg-��c���|��?-�x��)Z�H�k�O\�N%ҜejL�����q�&�U.1���;Ll�˛��qVN��aت(�*E��g��sJ���ܡ����%�q�*V/M������X49��b�W�t�:���Ե���m�o��E�@�C*!��S�o�d�[d�r�;���̿lN�q�A�6��c�9��d�s��k�q�����[SSG���6��]�����L+�ق�P��F�`"\�J�>k9����my2�4s鵴�{�+/�4�G��{#�a1��	o��F;�y����Ԥr3u��dRD�(S�8���j��}ǎįtֻ��@�x�-��<'��b�2�v���4�TIE��mX�>�1�۷��UN��0Nh;zθ����8��6�}�ljf.�ep���q�{t&{�����m�d��pp��\�Y�c�4֘�*"���Se䱠�`��0��g�q5E4�Z��u�A`i�u~�He�R�u�$�>]������9���bSϵ�ݧ�K��ڋ�d����+�ql��{;�i��E��c楀j��Q�{.�e�HQ�t�h�q�vE�靱B)7ClP�>�Q ?Ͽ��!{�ݴ#"owZt�渄����Lo'��xx�,̉5�'��� �&�W�x1I�HH{���=��:��O+�^}�S~_�����&9���)�/m?� X��2����7��#�F>�n���iO� d&|�����S[c��a��c��3�-R���*�U|Ƀ?�W89��B����H)�����9O�\:�7~2i�	wΗU�H��7�����4�H�ay�]�Z�S���/W�86�f�Nvx��ۚ�-��w'�u���kC��4��|/��ϊ�e7{C�i��.�3��t	kg�ͻ}cUk9G"�����#Щx�yaa���}��g#�����rm��IK���v�jmu�e�z��rq)�{B����������ҹS�
Hq�(D��?^S|ފRR獞f��}*K��Q�4AJ��'�l���Z�+k�F���Hw&�3�s(��O�1�9C�Ⱥ@��NT#]M(2":a	~�<ɤﱾ������lnx'��Y���ݎ����1GA���^����o��"�ƾ�z�GX���|�� b���iy��b��ŧ�΋�r�`1�|.���T_�7� �cH�͚<��ҕ\!�@�['��:����T�����f�����>�[U!O���xK#s�O؟�g��Q\�^�0�z��o1B��V�׳� ϼh��2=�G�٩ɶ(dkM-98����q>��f^O�q��.{�\����2J��$��� _~��t���n��
�?��ͺB��؄��,���W���.�-uqn^�����m��;Q��;)��>���������A���t2��Vw�$�����:-���	�s�GvL������g�?�߶M"5�(q�jiU��6�*\zT]F��.���yQ~���汃F4�NVO�J�W;{L�7C�n�ϱT��]+o�/�X^G�2��Sm�I�mڑ�2v��� I��+dj�F?>p/M�k��)g�bY��s4ٌ(��EB�zS�� V�C�	fsKIK5��h�� ��]��Z�OH�\��ZGtuiD;�x_'���*TKLD��!��q{�4��Q��Jq�`ĿV�gv�LC�A]�w���=l)57:�E��t�wx�θif[�-��Ұ������rMb�1�&���p�����hY~~O�1�Y�#�u����(�;%[��Ni��~]I�bG�У6������K�g~�
����'�X@Fǯ~�����WG��C3"V�F� ������Z+`�v7к@AQ�e�gq����?�v���c'7�9�n�r�֎��^�9���/]G+U7�������O7�k, &k��fr>=f&���v<�j8$�Cqa�O��r����Av�rm&:���,�e�׭<�xn�xė�X4;V����<��#��B֑v�N[�Ћ�����a�C��`�K�����G	�a�ny��hs�4��C��U
�q �vk����^�}fx�����ܓZ�V��h3ݏ,}먏N�ELk[�#��a�Z���˥]wl�(�F��*Ef� ly�"0���781 ���s��l�i��s�Ń����Ԝ��T��3*��f[\a9r�6N�����#n��^мT��eJ�މ���T��_D�*a�"��]o*#��<���HIɋsO�|/Uw�v��/�|�LGi���F�'|��F�����0�4d`�9�����ח�3˅�<o�6�k�j
I�S�Ri{�oO�d�(c���}\�i<S�C�!��v���'�h�"\�c�k����LK�gh\H�������H���)O�KҬ|��F�EP��X���y��^ �T�k�9аJz���w��F�m�3�ԯ>���t�q�\�f����<��K�SF���0�D���Ȣ[.�T�AwXb�}�m��� +����,l���>�:���\���_���#�My�P�%�姴��Qhp�,Ƙm!.0��{��BI]A�3����8�ɝ�?j36��̔�A(�%_@��I߮a}�Z�LK�5A���)k���I�N�қ��NQ�u4*��뷄�!`D�p*}	�� B|���1Y�^: �tQj�qH�c�In�I��fu���D�|ei �.�N�%i���F�ȇ�/������_�x�a~[�e�#�\��[��Lt�^͔��:��'���93W���u?���<԰����|]1bˠ�j�g��@�U$@b�O`
�^�f�,3�=�g��eՋF������I뙇����QЈ���)�u����d+�.u/������
(@�UVk�x���Y���XWwRQ�y���M1�I�~<�?GS9,��Sw��b�?�{����Z�t�S�9�� �:%nf�v���>YQ�<񴐍c�0E5��d+e0_9������?/�_��`̙*�-�ߺ����m��v���HBm�V��uҚ]�We�"�&�l<Uc�S4�����^?���[m�Y��e�+�v�*�&��>	s��`��%����n�,�
��ua�?0#bw$I��B
e�z�*A��pw�\���]өV�?��?L�.��P��T3طt��H����X��e;5�x��'zX'Ug�⤶
n{��a����-�ƽKI�C/�����q� T6��A�.zm �߲����N��"�w=/!��?��Hz�I]����� ��<��a�͛��ߤ�&������N�idc=g<�M�If� 67#��~����X�Gh���,e&����N��lMQia���%��c�w-���p�g�
�O-L$�w����<�)Ɖ���3Z~�߄<ʕP�����^Ac�(;M��%8�oY`��ₑ����2��	ֲ�n-�tQ�e� Ԇ�B�֒۠�%�F��)<�����G56C;�8K���TFF���ʖ���!\���An�_��ʻ�_oR�˜a¤glń����t=�E�o�������1ow�굹׾��h�u��"�?M������P�ړ��x.��E�O�H������̏�*�� �d���[�P? �h�G�����@�ĖŞ��C����R/����xu����E.�Apo�c�REv'Y~�81�-�6��K#bW�d�Z�0}sO�NI�R>֎��)<�]%�!�{s�q����E�lW�K������4���ʎ�"��'�(���/�����mF,��~P�8;�M&0�g8p`�{D9��U�J�����T���D����Dxb�%n�`%1U���(Pd�#Yy�NV�������w`���jG�FEpFbؐ^z����@R�̿�'�p�g������� �s?f"�,!ˉR	0��&�c}&���X`�~�':J+�|��۠D� ������]]m;�/�	�9d��-�[fKbf'�4��e��$�4<w$̿��c�8��5�-�Dwݒ��uʕ��ā�8)Y���O��vlqTB�u��5��� �~��oA)W҈�#T��{Z���wȉ��J-�bص��3���PٸW<�DV��T�V�E����nF����o�v��QK�C#M�Ǩ�pa��P��5c04Z`�7�C|^�@Uw/�Bo�I@���5�K �uH}��#�}t�a�Ma����Κ�H��ڐ�9yB/���e��>��14���pPcʫ�C��&�_��ĸ��?���O��d0�5<�����w�=kO�)Ŵ2h����O�uU^y,�H��ن�BC��=��V�!�F@�� s�����)�f�Ўi���=�"\C���2��{���[3��X�P��B��O�����_���S�� O2�Q(޲�E��Q_�q|=M&���]��-�dp�'��Z���x��s���/��"�h$�+`�!v5�a��Bf��>�e)d^_=xľ(�?�pb��G_�)�t�����=	i]&�B�|�pR:G�,�tR��ޛ��6t��z��j���Aپ���2�5�'�Wy}�S;�[�YG���6~�b]�4v�nŧ;{�ҘN�������os���A ��i:���|!�D�:v�?@���+n��h�1S�Q�|-�m필����Gn/N2n�N��	�>]oyO�W�?�8L�����p����,2媁'"�3c� �*PD����VN4�1A���Q�V��l_r!��\�O���Ϡ�	�"sjiT:��Cn+?����Ǉ�ee-K�ƚ!Z��U�~'s#���u����3�>������2��p�i|��/w^�Z�y���y�<�Z�3H����S��c�8�z�"$"��ߍ�4�C.r��ߘ����f^��]Y	�4���i;g#�?���A��A��Aa3����u�O�j�db��c���d�$����h麀�w�S�r@���e�a^���^$BL����R��
���W�
6%:���N���R%����|o��$p��X:Iq���s�-1�����
��0=�}RM`%��1��Jc�%y��c�϶��t���b�D�oz!SYO�l$�_A�Lv`��I��QP�|��9r}(4tu�\�XEª�i*��	Q# �kig��;fn<��	gp1�  Y�oQ�b@�{q�+��m:���3z�
����ty��0��P1����>�u@�EҖ�L���l4#Z�.(����AL���>�)_��4u.�dSiZ�.��:�AIџ�8'h[��ò+�h����A�`�i5�
�5�?��}���C53!�;.8���8B�b@����\{]%,<�D����h��1���J#:3�6j��*�ͫ{Mq�a;��_v:C�c�\��x�XACفH�b`��\�ӂe����~�m��F�'�Dԅ�3������M߁��?i�Ŏ{��^ ���Q�q���g���?��[�</�M�&5��;�hJQ@�~l�+��2�"��|�i)4�C��Z�o�ߵO���W�/��ۄ�x�keD����[�p���*py���힙!�y5|�Y��1�0�Tͮa��ٲ3�v�)�FJ+ɔ�)�a!��>��ʤrN)�m�ٶ��"F`�O"�"ӍPF�s�nB���fT�C	>��^!�T��Fg.Uߦ��x'F�2�5ʖj�R*זMd��i����03T�йd#F�%7�j��Y�\��VM��ĪH�^�a�I����O0/GA5�MD1�3HH��JZ>�������,�SjH�4�m!QX���X�  ;@�ѣ"�e�i��l�J]�,`@3�m0�RH�*K4����Dp�q	�g@m��9������k�ha����B���U{/�l���[���|GA��U��Q��Wd�?����鐖ʲ$$(b����yPyby� ��RGya(�d�̊��$��UR�;�J���,	o�}r�S���� �=�;уI���0���B�W5,M#����gL��oQR�u�.�ֶ����n���M���z��i�7���rE��������xj�
ie��HJ��[#�$�q(S\"���Ͷ7I�lDW�K
������6�}��/�И���
�V`��,��n��_K���x�a��D҇sm%��+�����ă�3�2�'X�E��g9���H��d��ߤj��0q���#t�%j�b�����
���ίE�$s<�6�z��|�=��2.K)�XJ��K�;~�����R���"�j�+�¢Y�@H��)y!������o8Q��A��`K狥)j_��P1{�Wۇ���}'��ۍ�1���85���{��K�$k�c�b�0ӾQ7z����)�Z�RB�
���ϔ��T�Q���a�ip�ePL�5/�/v�Ƣ�[�j�8;X�E�}�3��P�	<�ʸ�P�y�m�Y�{}�'W(����=��5a���K�r�R>�W�����=����`��b����h,�]#�k�aS��A	�{�X=|\hŐ��f��Wj�h��6p
Q	q1+����D�Hp#K鯮ֿ���w/�~ܰi�tP�_�*Gi�qc�M�@4̐}�˪�/��/ S�yM.&�P�o�T`��r��o�B��X����X���͍	�n��w1ym����p@����-W}�?j�s^���̢Ae�7���u��<?G�?��r�ƇZၓ��ȕ�fD��<�E��7)�Z�������87�8,�%�a�H�$Ox'ڳ��kW�)2�X���tAUw󞟔ި�I�Dݦ�Ip�~�/�~ΑAGDk�<t�V�'�!k�r`��{Iz�4�5���x�M�6	��`�%��9"�*�s<n�������<��޹.��w�F�YT6"�ƹ4D
.���k��2�j�w�s���&J,��6[U�S��bb���;7���	=CkqRم����(/�Y���
����/>q�4YnTh��F`�C��ѫX���Єt��*$�9��+��;9?R_�ުE�UG\�CƔ��|[��a⨼3��7;�O��M���ȟ��~�٠�t��f4k�w�Z���_��%ߵ#�i����g�4b��Ÿ�r[�U��� �nk���c�X7�f^�jz\�a�)��}�����-A=�h��=G�ү�G�|�l��Y��l; �b�vUR�й���ʉ!i��r��q������^���S/@��0�h�Vһ�_(^6+��9���!|<�Qh+�o�̶��Ȩ��W[�[(�6����R��I0���G�"_�=�aZ��pf*�M�X�Y+�E���f��@B��W�}?��'>�=�lc����xkܹ3}g��}q���.�$�E��Ӷ���F�罎ޭ�^�V��?0c�JW��d���5�ҹ�f�uK*W��m_��ɟ\��s���)u��P5X�^���� �b0�-q��UM@eQ>�#���2�q�P����
Sp�J�'��?��	3�n0�� ��tD��B��1R�pW��+�U���Ev-���[~rlG�/�:L���!JJ���O��5E�x�~�_�4{q,7�ohS��p�a����E�L�Ӯ㳝ׁO5�t6��1�R[.e��������:#`�j�}AL!�W@�^��� �̕o���%{����g�$�sE6�c-w7kл�8U�̓Iw2 �F��AdQ�͝�&����9��~��ߢ/����$O��c�D>#H_�Bl!�GQ(�ک���-�w'i�u:�ó�"K%^�j-�'t��h9;���a����7䰋2`�����C��P�@ճgd�G]8���������y:�DMG�ځB�T-z��#���z���\ȶ�$���mu؝�&��朩;U���Wfm�1D�f�-��י�qEp�~�X�ū6�Ĥ:��e�t5�<�����$M�; ����8������0hxXP���^������ֆ!oM឴-��z6	�^�Ը3/�\��"���'�G�����8��
h�2��`�g8�ʿ�'�@Z��2�QkЗͿ���s����C���oR�p��c��Ds�a���?�U�Tk�� y�+%��O�Z���B��M�.�4Dpe�$Z�s��0�򞢂��7<boz�����l�6���������,�#k�9B�fsHAQ�Ѡq!�CU�go��x�߬mϥ�#��c�C�!��c�c_��9��k�Bs˃�A�Ivv��(
��圽�as�q��.R.�uBO��p��K�.�6�*��o�;1O���ߪjϓ G"�/����[Y��7�1���5���k�<��-��}���-�% �	��)e�1�J�WI6M��}G�V���x \�wT�j�d2ڵ�m+"�	��ï����Vr��{5j� :�!|Ww��d��t�w��b�-�'z#�	0!���U��ӵW�X_r� ���^��U�jx�oݫ��=^S�h2�����3{�Z�Dy&2_W�
�ll�ctL��F8�rz6��z�[���|V*�7��-��q�ܙT�j9��0�y�0-�0�������	���i��>r��^������T3�{�w3�6U�̰O�o]ri����7�!&V{)�UmZ��/�<����ؼDB������u��x����v
� $�`�#��v�#�5{h�3 A�q+0,����>i�I$	ٴjV��E���ߢ����,ǳ!O�·/���l���`����1|-\kE�hJ@f!�J,��a'��#�a���J�U�N~�\��O�eU;����7j�=�EЅ=��1ug��x!���ᛲҗ����<�k���3��~}yƠn���ʷ+���[J޹S��&�)����+����Qg�Dk4�>�r����!)YV���h� �F�=A��d��0�/�ů�ȟ������j���a���bc���*��;⼁�3y�
Q��Z���L�6M	r{h�UH�5�(8��B�`ܪ�p��:>�\m��U�bDY$�rq=�ɴ�I�f�b�pjƢ@��CXX8��^�̪�m��5]�gQF�o���������tA~�#Hp�t�r�%SG��AX#����G)+m�ǋX�Fe�;[£�v*�x=�ҍ����°�(�6�T,�&�E�����%jߏ�5^������,�;m�۫X�
V�n��n��]#p���鴧��uy��|�c/�r�,Zq� s4�;.��+��Ù�O��	^)���w[+����ub�h��LFp��p)����h�L��<��'�2�5�yF�Ŭ/!�D�v��x��X�y�v�*�~8��*D�"}�2j���g\j���蜱�H��Cu#b5�ū%���? �u�m��:�8��C��WL�����o!����`�jս�zba��+Si�`�]�~��Ko!��+�Ƙ�7�W\�Պu�J���
��@w�Zb��ݨ���m�1\����y=箝Gd�+��豞����6H��$�4��:�	HI��P�2�"�@zo�7�#F_��D+|��k���4Y��T;��A����\B�r�oY���(�<�*��ZVu �������U���ڃތ$��I[���N�ӹ�J�έx�F��<t�9��z�-�$ \��c<]*��e�p�-�r��S%n.����&<�¤���ȳ���#K�a*]�>C-h��թv�L*t���Gw'���>�gaO��O��X����{�蛜p�z�]V�dW��#��~��xD�	��w�ҷ���Z&��S�W��2�<�'�M �S�d�w��r��)�9����d�4V����@�"�Hȃ	
%���{ʖ���m�TP�n�S0�mH���w�[�:��+r�C��(����!���ڄ�����Z8��e�(h�e�1YG����-��"R�q�r�)�L���ω>�_�$a6=L}�"г��=ܗ^�L%�"L���;����1Y/�ꓔb!�����z��OX��~ �䮱�i�x/K-T��ʻ`~����P�U���g�*)���a�� <4�7zq��,�c�'��T�� ЁE�RȠ���\3n�\�c(o��@�7{C2�^Z��̒����lę�Ͷ8����r33�6���Wr�V��dar
��c�#&}m���[Zu�����c�D�%(�z5��j;Nעa4L�roR)�y�����'�Z,�aF���D+�o�"K���r^(`�CL�6T���~%���պ�x�
 L�F]?%�����\�E�����9��Uׂ������z0	"�e��W1=z��M��`��i�+��a�Pc��
�XQ��!��"��'й�Qw㑊o���%�VD1��!�,n�V�-��2�2fT��ո�^G�����v�%W��(�IA힡$6A�/��	�[��\���l���r��xa��ᙼ�n��ef�b�0��ZmZ�rg3�����K%S_����z�'��D^ �͙�3ϱ�hֵ�@��a��0�-ov�6��iA*�ug��0�UcV>�}��yx���[��p��|��SCܺS���u�iA��c�*0����'�F��sA/�&n�.q)�O ��-��s�&P��4I�POu�ah�j�u��t?#�b�㉿@/��D�e#��8�(��3`L�Lr��^����S��2Z��ᰶ?��'	c)��k/l�-�j�9Ό�U?����YIM
c��Q�dT�ĩ.B�v��,�lW�a��U�QD�<*��q�n�hb�^D�q��㳲&�,W����q��՝��O��A��&k�5V�~46˸B�	�k)�&�a������a�0arP%�O���b��6H�S�V���99f~�h�ø�lC��_��aH���0;��Ί{�ҸJ��6���}� �"����Ks����vg�_��b���u��d����@��J��a�`�=3���Z;3�� |�-�+||��8Ը�j�nF�9�� ����<��Κ���� [��]!"%�s]=����(bx<o�M�p�V�'�#�K�P2��h�y)�wͪۗ��e��M
��r��-�=5lD�<j�+�,�+�L �A����i E�CLXz�̽���f!,Z�O^ͻVO{ō�VS,���AE˗X�)3�
!���.-�kL�|�����!�n}�<_��w+�󽂦�Y˛z�0%+[}
���>�3�85��Y� ]fKp�2j!]T���ի��e��v��$��b�ɚ�X�3�CN\@F�V�2'�hr������� I/1�u�Q���3���c��8�7��˥�\n�́.�E2{������e�Ze�_���0�#&)���)~&�u+o�����$Z�ޕԩ���	�7�c��>�h���2¯5�WߛR?)�e��,L����~���sb��v�,��+߭\�m�j��.�ļ�����v�w"�'��d0��Al�|�Y�FE�u�>�3���2�9�E��U�s�wFe3�؊�?P��8���[����K�f�O��#F [?HY���tY�����b�+4�Q�M4<�c>,���"�w6q��
S4���~�Xy$��a�c����~��_��f���iWM`\^L�:(�Y��@+����}�KW�K� 9<���l���52c}M��Bj�!BFb+{�ghC9xf�.2�-��G:�@�Ի�}ɡ;bH������P��LռO�]����x��#�V�pߛ���f}İ�i��s�e���3Z�T��VPF��� b���hV�����x|ka�VVJ�R-�6�2LiT�;=�}�-ip,��ʋ)�Hh���&*�-���A�`���/��U���72�CD�;`�6���#��lt�!fMr� zr�Xט�D�����
��"	k��U<e�	�[���c|������o�������q:��������.p���z\���i�1�x���]Twˉ'��[���#FS�����sj�l�6���s�c.�w~� �U����Rg%ɧ%���@�x��ƽ��þ0�HT�*�Eb�败}�	��:��4�C�RFL����x�� �ea�<7`� o�ǻK5"�	Zr6?c�!����p�Z�� 	���&ck��W�|�
4�=݁@�2�l @'<�c�-�=�,	��s��`�ܮJ��D�:�x�1J���:Ap̽;��9+����iA��9P7qf-Lo���DKI�A�`����!�#��j��vL�����R$}�V�V�N*Dl���{v����t��t��6�.�EL>˶%���l�
��JL�$W"/��O�ҋ*�9�pk� ֻ�� �,�����$�i(l~�i��Y-$5;<��%�/��AA/Xk�{�e���7^�V�k��C
(Sl̓��%�hX*ZF�1p�� �Ǔ���~�Z.�i`��15�7&1j���H��\��!��fB���y�;�#�����~pzʔ������A�z�i��KSj���1�(�u5�4�^�9o�K�[��e�ET��/�e#�ϪLN�0� e>;��^��:[}�&N�]��j��Z�R�3��y�������9BZ���h�'���Ne$Ю��PΑ)@ {��_������N�V�e�18/���iM����T6l�F��d^��?��#�.i>=@�~'x����d�v�<�(�v?߿��h��e���|ǟ�K��u^�Ї{� >h��:%�]e��Z� �)-�6��u��vv���s%��vD��r[YC�4��'-O�!]RU>I���n��Zv-NO6J�V* ;�3�Y�ȁ̼L�!��}�k	)Yw�4-Y�؈�U�)���^��>�"�q�����s�Sy�A��p�9��>�p���.\��f�FOZw�#	�Z�rqk�����e��d^;U�sL�N�sF���[��5�����+�&�mJi��`����,!��Tky� �6�9�	q[4��@fl�M�$OˌQY���<!��A|��)�%;�0d���J�[N�hH�^}�ކv[:�$�ɐ��*���>!:$�h���3���r��"�D�m�9�tF)�z�A_{a�ެ���Ea	82iJf�^�ӝ�`Ҷ������ia�����bJ	�-M{i&|z�D�1)��K��(NU����la��>A���f[���^��y�~\�>�O	Nk�O�����t�'���ݶ��)L1t]��`iW��a��P�%�yc1�s�`�В/��n��b>lҺ�Ɇ�x��(��+Bsg
���/?ШL	kL~�p{�2��?�0�F��� ���;#,�vH/$hBTw���1~��LC��{����E�ړ��A�Xנ6P��2Xjnf�����P�'��� �։���'xk�y���4�f�OF��J�waޕOt�J�-`��3�,x�-Bѹ�UI	L��Vă���*I&���\V���\���3��!#�z���ߍzr�at�'�7������@�[JŗT	P��ѻM�f޴u����:��Z�pd'��*�8e�&�q�#pn�t7�BdW"��Xb��v�xw�G�A� ��+&o��{���"�NhghS�w���ף�v�_�;��m�B��z��n���uF�@ܾ}4��og�!�C�>�n���`��@0_M�g�z
��������k�	_� ��L��{�n����)�+����n�v5a���T�=��Pp��bΞ@E9���>��vr+)0��UUB�
3mp*p[N�uQ�#�)<S/P�����{�D}�U�/#\%j��8��	�X� ���!ėh2�k�eE!e{�+���6��r���'ϔ�t�:܄�d1������}O7��mN>GI�g�&�#�? ��Kv��k�<�����ܷ��A%g.r�G��<?X��od_��þHY�����"M;�觗�$�?���G�����(V��8���w��cF�<JYE�����(|ԸXZ�4Il�S.c��8����	�-�L�V�T~�"o#�L ��]_����w��ģϔ;�Q|���Y�FoU���xg̒u)`0��a��̔�??�0�|���YN�o^���J�ԩ����`��9s���Ď���?q�(���<�Un�2;cݢ�{_	��J�?+����#����-���Q�q '8I�Z����p԰�[\'�H!"��?���B?hs���c�}��D��:F���U�)Q)&��q74#Ё����ς�%���C�T(�ţ��+c>��շ���A�
��\�����ӷ���wF�@(����/Ӫ>ܩ�"1[;EC]w<JEF�/���s<:�O�!^&q�M�����.yN��j���'�"DA�
�[g�O���*�2�?O�^k�\�T*�G�rxk5�2K{F�N	b�[
�0��Ε���W�;bUm<��U��[(��n�7$ڝ��ċ �I�z�R����w��T	��سF�m�Ag'eV�_?O1� �U��o_�0 ��0Y�0KhNU�����p$UӅ��������pz]`�P��>���d�gX��̼�?S<�a�������Z���TY�4w8�l��ak
h'�k��m_MB����T��"�b!���{_��ru���ý(MT?r� ��7�
0��k�mP�	i�O�(���R�֏���+�D����\GfN�+���_`� n����Ao�~s��]N!7B��������lj�>��+�D�d����J��YƯ|΀�l)����u��.�<��<�Nl��6mֵ󚶸N�wjQ��<��(�1��a�<���SVԱ�=Q,K�j[�:�0�U�m��-�@L��wJ[��Յ��L1��:���>܆��]�����|,���ݩ�\H�=��!
�Z�	�WU^`">�f�1�ˆ\lЍ�	���]!���
)֗vU�x�5�@��ų��P<o�L=�ԵF���n�	��(ied�mʚ
=i�9Lz���h�O��4�iNb�P-Z���;{`�t_�(|������Ȍ��I���<��F��E�$�23M\�X�$��1q 	mpnz���ucU������N��Е#�e4����̑��K��� b�(�,�;J��v.!�//�D�ه\W���ȟz��E���>6Z�\����#��3yK�� ؊X�-_�����t�ڛ)�:���$���bv�H г_�/1���y�L��?/�s��>v����++����k|��3��E���Cѐ|۠L��#ŻDҋ�>�Q+�ZΚ�XE�ʍ�>ۘ|)���Bh5���_�c����{ו+��$�������PM�|���I��FQɯ�r�Y��tL]�y���B��*�y���`�M�)�R�Y�(�7(����}R�Vby|�p4�Iq���L>3`R�D%�*�0G6��(w���X�����65�є݊�_3�D#�
\T���,�W��)�ب�j�&�����$�R�4݁�r(��j�Pm�B92�M��&e���Ś= ��h�3[n
}�����^��"�5#Gãy��c�x��"��h��a���uD>ȡ���^����'"�S�937�� Fנ\�N칠�|�!;F�J!�j=���ڳ��O,�����u�}���NW~�ؼ�m�1���m팆�a����t��n�Z��+^�!E��2nցs�AިS�/��T�J|�e��t�6X5��W��*�K��R���%�4U����Y_Lc�!����t�>���Ȇd0�1�3�&�X�d3^4�L���N��Y-�%G>�k�ڦ��r.���Yԍ�
��u�z=e��,?Nȭq�^OQ�ṋ�ؐ`Bu�칡�)4dU|t�^�}5`�
=.�(�<8�Q/��}�jC�Q��	��_��6/{"���� �$�1J�J��g/��&�k��<��Xa|	�R"x�����?۶��Q���&�j��Ӹ�.�ɍ�A���J��?J�wd�cw�n:����P��/�]�i�ʳ�˃�'�$đ[%����SDsrV��aL�,��N���VO����b}���݄�0�\K�0;�j�3��yz.��A*�;a��.
�l��O����1�[�-�nة4ny���~;}Gd��O';�M���"Sg*ѰB��Ny��Я������5�c�������L�j�J1T�Op���iĠ�7�jo�)��19�6�p�q�G�L%���%�>���`'�Mٛ���(�swśr�KC���[mWAhn�ϬX(vw�&�=R�2�$8���:����}i�5�|Is~�N��qhS���{�@{���?y��{zB`�S҆����Y]��$Ғ�p��/J����<��Ց��7�o���5�A ܔ%�����h�L+t�������������nԧ���z>����9�8�ܮ��c�W ]�ؓ�<^|�B���o+T9�� J�dل؃����t��j���
c�1��DQ���lW���[3�?K��MQ�t�|Z����yD�;bB�؊r��NC�E�nGg+G��X��=�C1k�vR�r0u?�3d�e�\p��Ps�q��{�!\��ث��D'1^%��G T̺�u�����,WG�wy�P�BI8���$Xy�S�+@��~��y�#Ü�%\�y��B7�N�?�����qqSk��:�i�^N�.(T%�=+��M$Ú6��S�����O9~�P�6�eߕ�h��,֯Td�%�\�p��=�a�d�'�/�6���7��9�����3J��l4���,ʠ��r��Q��Yf����������;�"+�뉄�Nm�w��^>���ke�>��2f��L���`:��<*�޳��ӗ�_�79
u�b�f��5bu�����@W�~��՚Sҙx�����7L�<#JUC +��<����w�/�P���:2�`�a��[���Lg"������';�#cm��?�-�q�Rf�	�p'�W���;߬��tb�Z[C5�����Ӌ�N �"Vx�UR"�M��t�E��@�֩�`��C?eRy��g��ǧݞC���n���6mq*4#��?����DLw�2�K��M��b�$�*r�̭E%z-Q��O����vū�,��#:� �rh.�,�4�k{��pw�O�%8�d��zu��������d�1�p5���&ξ��;�T����PD��=��]���kFk�M26��:t�����A�s���z�M����8]�@�=S��w��/ݐ�gA�Z�y;�,15�U!��I"�@�GL}�W�h:�	������ǚ�
�5M�����B��c�Z/�ת>}�OE�'��rHK~��n4�~�+χ�{�����0�n5��]S�Yܦ�F;i�p؈�F�{W�tW��.EhG�z�
+���
A�^>;�Ż�f��ܧ�.�5�|���4b4�0�Q�W��	`�r��K@���P��1�+�6zE��Ə`��I'��9ln{1��������D!c�3��e���bc�I����48��$p��ph�}�U.��m��Wײ����pg���5�����\� {GŌ��������Y�k^�
:Q���W���P�v�j�o��4�AA!�,�TP���V��;~TQfNl�V#@�X����[2�Љpt�"R$�YK}�6'n����6��S.l�~��Nɥw-�_���kw���sˍ�&�,VU�l�SWO���� ^Z��|���Q��zm(.A�v�,ûRWY�`i�{�i�)4�t�r{`e��5�������o��I�R��R�!���$"����I)b���p�	e�7�N��������!-]33�hіF��\J�,������^H͐�?�����c���ZmY��5d����2������䜖dȊ�|�	��fr"t��xTV�4꼔�����O��V>f���Q 6)Z��(č��Q.��{�e�9��v��0�o���0��h77����K{�IrD�Z^U�4Ý�)QC���%h�p|5)��\��D�~����+��i�ȫ!��(ÖS^��(�Q�N,�e M���:9?5#�ˬ��z��=�YFO끌>�F����BKKI��v�\�ﾛ+�Q�������Wh�7F����5x;
��F��>�L�%˫�(��p���l��d�~�5�ٛ����;x.��$�ž������v�P��"�B{�����'��ʝ���p��t�h=�t\���I���QF���Dt����?`�Ξ������K��8��ݪ^��M*!�X��cۍ����%�V)�p�9;ڲ��k�+�y�!��H����:4�Iʼ M��>	�� "��{����sg㐝��y9ߗw8Z�E(#��C9&n�8Ga�t���k!Ie-�����#"�#�{!<獰r����L��Z��ݸ������a�V��;������q/����TbD��K��A��h.^�{�yp8�|�硑�Ln>8u���c��F&�B%T����'�9Ukc�s��ɏ���7�es���wѻ��F�x��|�#�0�Y��3x��p,k� ,HD�Ub��gT�|0�����B�(H�#�5�1&:�����&ޘ�_=�?hݞg��+E�],��$d�Р�y!T@����g&�X߭��@���� ��~��nj�^D{�. HWt���q�u �7d'�G��Kk
5��Җ����l4��H��ޠ5��3 ��nx���ʑP��L]e�����Z�&	���/�Tδ��/�	|�vR���.���`h�WP�d[g@՟�W���"����>͇��Y�� ���$���M�܏�Ф�Y|�lA{̛���cMl��!	���Q�2"=�������)�O8l�H��r��9gV��g���墺�@1� �Y��L��}�gy�$�:lݗ7�3�1��mֵ��ǶU6r�3=�C�~:߰�P�依���x��#�Tc�G�8NJgq�h�mN��g���+���Ե�Et 3bJ-.��lb����%����G��"��'M��y�������A�	c�z;���j����؝�h�4��@S�*�H�����&��7�}��;�.|����4M��&����怚�!og��~�A8~%�!�+�ᇩ��< Z ݵ�����qi�����[�$�N����
�H�B��"I�Q%R�cZ�cmiZMy��g;�s�������`"�ˋP��_�''���O�!7K昤�(��7��fB�|��_�Ս�j��B׋ }Q` �p7�fU�,?psb�q���O�Nq��m�+�+OǧA��O �P�����5��ou%�!+aF�G:<yuRuS��=���y����|��^�[!���xK����\\8���YO#1�[,w�� D���˓���9:G3P�g|U1N��K@��BUx���yf���u�F� �j.�	M�8�Z�8�C|v�V�.���`��I�g�/�E*�ّ>��e:�m���G��c�m�r/;+�t��{��_9)ftO�/�ǩ���邭i�S�[��)\�O�4	.�����(����7���5�~ُ��z��\)�L䆂j,緵6*�v�4����Z����f�W�Gt7O��9Lk��kI�MRk�;Fp�Xl@��)�� a�"��F���9�ָ�L���v�� �����l��sC7\�@)�"�k�oXu��F��v4t !��3EQ���m�v�[�����!"*�r�����x �Տ�kc���(ۯ���7_M�6ު�C�":.,]s���l�?(�X��s�]�� e�Y'>��Dnp>�X����'������6�b\�U����s��7��x�5�B喦޸�S{e^�CY�H^g��e�Γ5�-��F�dù���$��L$�T�>B�������FG%`����fTC�F�ɣ�� ���iip�eW�;ux�ଝ��@J�7�4�����4뜝[s�Q��\�y��X�34':�yqv��8�ڀ�3�JUu��3���&a&�e�Cߑ4?� �ے��,�A�3޲�f���Z�%�փ�cmX�)���,�H�H�W�A�ⅅ+mNrj:�������j��=�+Y�
��~)g}���H�3sWY��?��]N��o�t~���'zH�p��'xH���X����w��$���������r��p���*Z՚��]y��uc�2��?cԼ9�v�� `EXv������Y຿�q�����}�.5B����3���_yxu(�׭�+�'>��~X�O�5se����T��c��;-��F"iJ�����$H&�:��t3�54#��1��[�u���+P�Z<���!������1iw�*���Z-.�+�10qs�>�w����ONsK��9�3�0�Qn�j�)|1��J�NT�k�0����"PMa�����KA����C/��L��=������m���F�ml�ש2���N�J�Nc�"+�׆�b��g���e���� �^cB���{2ɳ��1�8��,�)`���:���_틗���FB�WKc�F�<�M�w�㚻���0r�PJgȼu��7D��ex��w8��:!�$���-,b<QB�����(�_�"�m/� }���<�s�eTR���F��iq�J�5�06N8G�PB�I��)k�P5�;�w�?Nh�e��X������w,�*]���S}:�:Wx*��۔�j�Z蜖���6�Rl�	u�g�'���|��7��_�����["э}��}C}�%-#;\X&V��T���z��<�~�Ђu���Sú�0�_����Z�s�ڏn �l��#u���
F\�7X,J %�M�Fa��fH���ySJIcE�]75�?L4�H2zb�,c��~��Cdq
�]4�
���P�<'�$)�T�t���Ӵ|�ŝ�B�@���� r&hd�Ec�"B�'��*5�'��_4Pf-�����pu�y�F��������L��ޯs{������DlCr4��L�@���~���/����±3$ۼ֧�0����y}�r���삦�ۗ@4�����[Jʵֵ� ��k"b6p���0��.e_��/D�0:��?��ty�Y&2tvM���Ak� ͅ-<as@z9Y��)���
��Q��f���v�a՘����6��f��I�Y�i5v��
��� LS�R�W���h���̔ꨜ���B��P\��Kg�p�
W�"jT�N����ry�K��Vl�X�35�W�?�]�l��d������߅ B)+�˸�5ڞ9�	E<f=�Oſ&ƛ�P�\n����ӭ$N�F��>o40��1��� �黌{������o��>��$ib�Y��c+W�G��&?��Y$j�(�$��(�-~λF >_t�_�x�)2��}{H�O���@3�����nݣ0�ǖ��mP�l+����Qr��Y�Z$S	^�be#�t.Ext��4�.�.�7g�By�×T 2dmFp;�ڲ�"C�������C����6<ۿ��	���j�/u�3�����H�f8�x�����賢:Kr=�S.B����b]3�|�}��k����
Ϟ��đ@%��}���G/g�lT�X9.�������B���h>�Y������������!�e�9�<H��E��)�SG������*s�I�c��V�Nh��9�ʦ`��R�|g�җ��<%Rq0�^]&Ɨ�G,Gt���U�ZRD�d�%Sݼ�r���8^�C����0���Dp'��[���xoE��G~����J�0C�R����J7�'��	Nw}��7B���It0���8A��=�{���q��dc�:_c@�8���R� KM~�2��kv�`��i�������L��pA*�`�`�X�������=E"��:h��oQid���Us�BAK��#J[�[���BAD��ކN���l�V��M�1G`��N���N2�[��~�Ę���6��4[0&��ofZ�9-g�&uG�ɕȄ����-ɳ��Qqռዏh8��a���Z��$w�b��Hn��RNKO[�n����rghp����Hv�|��2����?ǄK�>�/�DEꢣ�b?�;��+iTk=���d+�'�;������_�N���}�
��U���,݊.�r�I/���c ���ds%���b�W!�o�b=X�Y�W4��;@���5�ρM����$u�cMX���~(� �m��g ^����!q�N1q�p��l��x�Ϩf;�f�Jyv;��I *H����\�f�����cS"ӷ7���G,��,�6��!\@��7���ۋЀ��%�'̚)�t�:o�^W���5�C�o����G-��������fR�l9dڄܐ	%ۗ2��r'�O��V���ӊ��n�%�o�^���]�/++�����C�g0�s���[3_oм�����/V�WXףٖ��I*�J	J�T7��� o�խ���^�ԋ޴�Xt��C�W�H8�M�=�e>{�y �=�ЇHȾ�/����&.c/͒��Mf���� ML����X}�*���o����L�Y�c�O:���^do����)N۔%�B]h�}S��+��"���K���U�۳Xn����a��ݥq{>#���j�j�\�i��<,��q�8h�1,5rQ�y�SQ���Rǉ}�����*+ĉ��u��j�5`�ںRב@P{��k�
��8uw�-��,WL_,;q]j��G�>/��0����<���e�f]�X����\2̵�-�VP?Uל+T {�'pM�G���t�~����q�� {x���#�$&>א!�:y$<ޓ�����[�V��<�r�`�7/ %֐kkV���㍅lf��x�9ŝ��-�~Mv������2��LK�Ϡ+Փg��!���AFu�{�O+v6_/^4J{f���BX!3�|�pO)�F�ٌc[�pc� ֱ������g��x��i}��Шʲ�Q���Ar07눿�ghߒ1���A�2̣_U.-oD�
�D��O�U#	�fnf�:��9�L��&(��ɱ��l֒��g��&
��Eh�"7\��o��攑Bi��R;b�Nb���'�m��2��B�QZ.���L���0jf����@=o!��G��r��(f�S��i�D+d��)�����j�F��vdU�m��d@+P��v�A��BCD�ww����
d��	x\��qM�N��1)ĥt����u���پK�'^�򳐳u�7����y	g�Q��O(�xQx�ڰ�z��s|�(�v�����f�)�m�S�n��L�������,Q�_�������v3���0�^��-�+wR�e��5�,���彬O׋?.m�f�Z���Ppk��&z�����c����g`m�yJ�?���Q����-��au*��,Y^H1�=��/Vɳ8���%?�A=��[Ѿ��3��F�xN/snUAJ��^��Ĵ)�V~ewb�XR�T�r=��ݍ'v`v�#i4�W��h ~��F���g�u�F{F셟7L*8�Y�-}�W���ʴi�<��$h�N`�\fF-h��
$���C��{�j��cR>~��fA*���j?�}5ߏ����}S���_�[c�.�C��A�^�í�k�j�S�u���a�����>�B�.�S�"��U���� k��'j��Q<R	��K�e�t�!���,ϰŃ~?��X���=����?����/)&��_)��+s��	/|Wpn�z@p������6�9���y7�zfF��S� �m2�fE�R�`Ǭ�p��?�4:Nv�;۶Qc�VEX/�'��y2�����FtP�W%�-E���f	-�V��f9<�mZ(yK�P"1a#Qۂ�T��u����|���H���F(���� ^�]F�� G�fiYP׍	s���h\�[�!~�FL�G]b�
�7���w�_7F~ �ȶ�4vps��ڡɯ��d��hT�f�-�!���Lw��DP�~���F��Wme3�R�Z�{�n*Jߴ�R)~�����(DO��9(�t�b+�d��t���|#��q���|���4�q"�D�z�A������7���ha��Q��a���a� خ>�0ۓ�@�>��t��f��Mz��iRU�����ݢ���k8���(������p���AMle�b�ǡ7�ݫ�-�$� ��v�qOP��A����%�gEũ*�*���(��^1Pg�����t雁���i[����ʧNJ��������P��
t��
ǻ]eli�~H��w� ���Q��C|�Ҽ�V�����"r7]��̃5�"p��Xͷb��)Eb����C�:p�)��!���������"��&~ 
ɚ:�L����| �%�E\�Ƴ��\j��P�yV�/�/iD.ڼ�*��(hE�(���Ӓ�l��C����x��	�	���8ea�j͓��H������?��%���m�<�{������"�6E��Sg͓�
Z����8R�(ѩ�plJ�[��z�d�;��On+Q�	��W��w�'�C*/L_����6�B��>���������5�o��r�����m3�5z��H}K�c�#����q���_[�Zk�� Cl�����E[�U	� ch#���!���?��o��/f���/��%I� ��pgp	��=�!�N�����0��V�|S�����I��;9�uq���3�N����&�_���o�BD�y�[ޛ�\.��/�_ x�S���d󳹋��"�1��;Hg���*��]
A�^o�h��]���p/N��������\��kѧ��1|��ǾT���ĝ�Ö6� �ֽ�4-�e��MS,��7��]�WY��-iL\_��'*�;b?�/Z���18��󝂨��M;�;"�-.p[9��$ ��j�1�\}J��p)��Ʉ�Y��?�$P��n�)L�����s���,_4�/��8�V�cQھ(����$�1ɐ��̰'�O�ZhCU�8-&���`X3�K����v6�{/��T3z>C�B���=4ŉ�@Y³�Q��u `$ӭ=ފ��%�?Fp����녰YEO�)6]�=���G���z���"��PG�._bآ��U�:L�x��[l�^]��ҘϘL���5>3�M1�l�<��V�{2ӣ���J��'l+}�a���x�B��CQU% $������*�ppdЄ@�q��ʣ�-mV��%�b��!�q`��H�{[*Nn�]���n�u����8�� �ceӨ� ,�.jD_���K�$���l��,�L27������
�� Pkz�;;cɰ���l#!RcL�Q�`�һO���2j%���&@���T�#���5X���N$���h�ӌ�y\�Q�6,6��nò	P��K1�=��H+In#�
<FF���R�R�`�i�;�d[�m�x�P�������;x(|o�?�6��� ���r���Fw�4�fnm�Qsi��4V�ç�}����J��`ᓮr2������8��)�r�z6�2P�K�|��#����=u��ű����$��P�%)Ö��"������(��(��^ߛ����<�A�R� c���[:����0��L���S]�ă����原���s.��Jڰ��b�#����T@>ڄ��˫��Ϻ���q������}־ϫ:1�P�ݞ�w� ��~U�� �h��|�Y�CI(׻$k��������g�ڇLf�N⿀<G��.�o9MD�V{�[/�C��&;�Yu�WL	4J����P�f*v��l+(�fO#�w�詧����5�BslW��{YG����y��Ma�*o��wl��ޢ2���
�_����-!��FOl^;�!�Ý�����P�Ʊ��v�OD��\&�X~�m6�e��Ya�9F�*�|�o}�bW|h��m����ޑjl��@4>�'b�\������T�:��̻Fϑ%N&�'� ��̾��p���6�IY�u��n��X��y�ަ*�0�7��(�r�ܥ��I�R��@@���r1g��*1mp>���h������i,��P��@�%,����⟓܃+�O�h�߰)����Y��g�7������Y��J��K��%�v!���Q�cAX��.���������*#�dؿ+��/���B���[�;��T�q�g����K��F#�i���(�ttƈ��
��Q2���>�S?]c��_3���X��(3�S�q��������B���v�����@�h٧�{5UQ���f�E��K���m��ܖ� �YcoaG�B��h �t#�Y��ew�%�/�a xoBFj��`����'���n�p;����o�ǘ��o|��>2���A.��j����sč��zH�%^��7\.�9�d�3�j2D:�`_��]S���%����DmD���]w�g�#̺e�	�Un��ww���= �e~z�<��U)v�JϫJ#dw�Ew.i��cՐشA�Sl[���L)��y_W���]���
Д/�p�S�=� %&A�7	��f"*<�J�n��Hd�B2` h�|���;+����Q�r�vV*,6����q�m������Al݅���%�.Ny�n��6s~N=vefDmX����.m<�P����}�	���
��L��cGw�E,����-ǡ������Tl���BBe���
6P
J�m�BW�T@�d��K	�	�Ф���qN�e��ջ�����1��(�*L�w:v4���B�y��L&T�2��h�c�sGfT.5!���4�Lae{�|�7���RD�f<h=:�����r��� ^U���oB/�]xc�qsxCq�����0�$�F����F���Cg�!/��T��'/��U���i����cl�{�9"cm��ħ�2�.+��[�L��� ��������(�!�2a�;Z������Y��q�1|F�=،M^Z��mC��M���/&�M[����V�3�V��< 5��m�wl���G�	:`y�P)�O��)���ŝB�q�;9sa�oL7	��`��eQY�M��^���*&��<J�)���;�� H��G<�1�}BҐ�Nc��U��2pN��%�2R���1f���	Lu�V\͌��z�۪o�t��r��!`���4��'g�j��HYw:��D�Dp�f]e���9/]$��c-��Xc��͇ڟ�2��G��}G�D8���]6�B�!�����j-fh�<�-�lrml�z�0���P��"�W�6@堙�q��jtM+��)���	�l����mzr��lL�G��ǣ�&rmS�<)��.�w��c�>Rю����^����*-纆��!	�
<�Q�}���е��^�ײ�-kFN�m�x�T<�fI@-U��s,8�kp��Me�B:Cg:u? ��
t7�k�gج�5�ȏ9�>~�VC)���M��*�=�_)���ɮJ��7l�,�eZ1��8T��9��%X���Mܩ@ǣ������Nri��f���_F�����ֶQ������vX��m�ſ�
�U�M&Yau�߸]�O��y"i��oyGA?9b���)��D��%Y�����31�:����3�'=@�w��Or�vl�H��}�uf�u����lb��u�����d-��Ҡ���_��Z�j�\d�~Y� �+���IK��d�����f3u�w��Nk�K_��ӹ���^�Fʠ�h��T�ƕU��aX����5�؜+��'T��l�T�*��%MR_��1+D(�A/��Ro}cx\��_|���������8'���Mx&��'|N���C����w� �Ò�$�x^�+���;}-�bݛ=`���0;`D��c��yӤ�鱰
����u� Ka-��n���kt_?%�ݓ�;s֒٣ck���	_�V����pn�!ִt��c���T��H�w�N���0T�~�����L�'���D�ʈ��t��jzp�NF�[�Lle6���i ��Z���Ts V��H9�	G��C$�2wdm��Ka�m2����hZ����B��E���vv'�u�O����%���aoÓؾKz�"@�Έ��ǉr'J
�������-{/��a�蹿u�gц/�J�z�gi�%{>3\��w�A��,�&>S༞`��4Ql&I�̩~�b����c��*z.a>��)b1��u�p;�Xc����Q���h��\�r+�
��-���9�=L#���`d�*��)<��?HN���n�!Y����Sl7�wՂ��c��빔�?&�6�h��y����^UPÚ�Nץ�(K�5���L֍UL����|�����Y1��7<-鮜 �"Ӓ���/�����`���А��K�mR+��O�$�[�����{0����m>EI���|���F��Xc�*@)�>����Q�������!k��9#��1K-V���,��ພ���Q�3`���'�t���T���h[^��4�blݞժ�b�0@RTv��9�4�O#�AA`ԖB���3������i�b܉��C�]P�t ��/������6����K���Do�׏��:&$�_x�|�[�Ps���ve��ً���Wo��F����
�;e�gͶS�@�[٘g����߽��KC�w\�JeA,�:B]=MAS;g�s�2,gi��jߗ�_�Y�Ŝh���+F6bt�4�����cr�gJ��<�KB��;&Ԓbm/�����t�_U�*��Eĝ)�(���q�_"�4n�y��#�s	�_��
xv-�Q�5w@UϦ��K�1��%T,f;�߶l���["��e�O�|�\oL�������&̵����0��Qi��_7��3���� $s�I�i�7ܵ��oy�5�	A?K6ū}@{}9Uqe��z��!�a�N&^��^�ؓZz�������pZ�<��g"Yt�S��;v!@�fa����>W�'��b����hz��"�ܬ[��{��i�z�&X�z1��
ɵL���7:�v+��Цž����?R�;]�d� �,e[�@�U珯�e}��+�4��@�;\D��:�E�g�!��U�1���5?'6+?���
S�?�~g�4y ���S�ydZg��r��Cƚh�� M��ϸ'A�<o)P�I��|)�.V���W�A(nqu� ��8܀�PU�*��S:�����)����"�����v��Z�j�������βF��2��o�]h���ǂ��K��6��gp�f��b3����Ο
7��m�lĳW�`�1R��'%�(��1�w��$ ��9Ĳ���T�|mk)��@�@"D-a���R���B��A��Gy������=N�sX	���n5���9m�lJ��O��e�Z��x�Y�������1���`�2�;z/��D~�]�Uk��Px�f�U��nAi"��'N���hX�s��&��2���Y����TO�[��3{�_N�wd{
�a]��SH�+k���Q����4���iV�H_��XW �y�(B�U0�j���H��T-z?�$������']:�7��k�9<�n�q���C�� ���Yx	a��ey$� ��J�Y���{�[�-���wE�noO�����hi-.���B��=Xd���h�B���/�شLTEH��ו$r~|��E��I�BեE��Cp���N+J��/���^�RE�I�D�LĆ��|E��5��Ӌ1ުw�P�
��(Q7�fX�y=�X��32��͐b�,!֠}M5�.J`���c*�D"�a_6�ʫ0�[`�ր���<�_�PU �Q\`�j����t.H�)�S:�iNOū���Р	&�KB@O�DY�1�$��Ä�ؤ_�E<��r��	��gj;��.�G}]G ׁ
y�_,�SPf|,�Hj}����Z
�ϡ<��R=�Lr��0�-�H��а8
w<��wkr��s��.����Wf>^y4@���cF�]����"�i:�����Z[��)�h̏О�+��-6��.S��x�&�
�p.�BV����B�3mW�k�޷Z �Í�h�bۈH��S��Z'}?��$Z�9�|�,�竀{r��`�:�7ԥ�ѣeO���&d��������UC�����8;��?�dE_r�S���Fg��)������츻T)k���&�����25����E8֡IF+�
5��S�KYy��;ـ�Ǒ*�'��s��=��E�.�b��`��ҕLi!|����=�3\g�<�Gy�tƭS��g�MWH���0����k������:D~�gA�ӡ��J��~�o�o`}:�@ĝ͒�چ�n��n$(��I}&�q���9�ONR�|c��4�@��-w���)뚆bk"��9��UL��8�c�8��?���hm}�-�$�y�7b�b��Ã��+|�cWu�J�S:�D����m��8�a+s!��
�}�RK�Q3	l&��� �d5���g؂`�o�&���+@s2��i�Ej4Fk�/*i��������ԟ���0j{�_8�`�
\�D��
o㾩�>7�[G�/�\�`�5y�9� xM�U2�g^���m-Y�����F�U��a]�qmɱߞ��>PK�\���-��M�	3P4.��r<�����o'�z����2L�ۂ���uY>͢�夬&�}���Еl�HV�-cqx1kTf_U����l@L�	���k��p�Y��`��:ٽpDm4d�~�렯��>~F���r�7`�?�`�1 �U�����1�N��e�$���L���dB��<L�k���KH����O"`7(���Pp}l;y�H��4���/y-Uԃ�!e,ֶ��>�@@W8�q-$;{��"� ������b��򦎢)���,������W�txqǦU�t�9����N@���g�OD����UFl�rp-�	��Jr����X`�tU�Ⱥ�t3LUJ�k���CG��8x���ͮJ|��H�]�~f�+��4�Կ�>p�y�Q>O�YS�Bb��d{-���c��%�d�=T���"�.�N�2g��yi�PY��<Am�~�҈���R�<�%)��5zY��S(�������]z�n����T�� �Ȓ%����8}��vtL���Dzve}�.��CV%�P��El�4�p4c����qz�cv5�þ��22h��N1�K�%-A��Ζ���{l⏌�!"@氒��T8r�L4Uζ����`�6W�ӧ�HH��L=g*~���-J�$~�9 �e�6�pS�c�U����8tE�ڪ��MVq˲�f����@�ޘs"GЂ}�J��tu�ʏ2��̊��e��������ezfw��^���ɣtP�SF��������w��@�/���P"楑
u$[�����rٝ��!ʨ�<���؂Q坿�< ��{2Q�Ñ ����Ҟ�v�cW���HD]V��n8@կݎ� �V,�@�HLȫ:7�;F��R��aA��)�:�f�źQ�Y=Xt��F�z���������]�*sYyq=Z�=}u�L���E���Bܵ�O��!���`�?�F��F�1q>u@�$,&bMFO�O�`�S�hm2c�6�s-�']t��|����tH����g��W��[)��
0c4�-����?������t̡|�	����h����#m��9�X��y!�_�ߨY��5�����=�t�n���)����f*<��D�]0�(���(���������`}_���ۿ21+����=byt��?�I"�#�}�5xY��ǚ�2�9,���g �Fok�Cj�t��Y�����Ǚ7�|pq����.�5������d�!쿡\~@%$�<r%���iT���`Ռ�#�4���(�y��*����[���ͧ���U���j�/�b�5�8�T0�u�	�	ls Me'r�E����W�N.X��sT�"t�zS�k�s<rV+p�{Q;`I:sz�v�8���fP�v)��'`�DB�>R�T���Cv���	ƻ%'������J�PL�IBN�TlԴ.ZԬ\��1kv��:�( ������^]��S� �:����on��F0�2lcP]w���y�5KO��mË��ԫ��v���ͧ���U�j?E ?3	�XF�k�2���S��n���]"�	��~8�gua��¤��X��9�R��� \�M�d�.�}nr�tr�W����N
��g�<m�־i���-t��o��87o��~�y��;S_���C��u/2��,�t�GNv$ealA!(	���!}SY��O6�~/,�@Us��7��3ʟ�;H��C@M4���}�Ϡ��ê|5O��H��g!,�X��ݏiGͦx�R��2������-:qY��d��m<,���0����_)Y�.� �
����#�w�m��� �]F����k\�ÂK5c�_�0Đ�s��#��-�MHw�#t>܃4�a:�c�آjw>ZJ��ԣ�m�<���v )g2m�F��[l�_�?Z@FI�
�q��S�Jt��@@�L���=NAA��	^x{[o9��˘@#�nk�z���x*�r��e��?�dSlV4�he�A��s3��_�z��^�[�&�kŐ�bC2�����o5���������8�������r���Hվ�x�KX�#��u����J��Q`#%O��O��B'���,��2��N?ZO��Hf�� ��S��RAV?�a<�J3�倅KY�"ȝ���Gi�9V��UC����I���7�3k�l�M)�X���{৹ ]�����EYo��4�^+#ʴ�m�Ӳ��w�~=��n���jMF�u�$�ު�;���}P�9��4��6�n�?��Q�'N��qQ*l�s*���3=6oH�è��ڒ�'�}<��&������.�QO�7�-��Vw�^/�39� �+�mv��2o��0��hoJJ�T����R����нv�A��h�& �q^-���N4!�m�[�,�}gȔ	�`S=��~�B��t���<2���qe�[�la��+���P�t��u5eHV�H����Dp�w�ey>`��N��PH�I����� �E���4��������A��U��Q5���ݹN|�۾�����X���������c�~��%�ຖ������`�H7�[�	������6��c3"f���I��D���+w���~���8�27[��u�����P����E���m����n?�@'��%Bd�x�	����KO�{����Qe��B<�IzqY�
O�q�[��Ny;P��XD?TxV�\�/����ToaX��(yZ���+�(��bR�[�;��sS�%N���ҷN蝠mdN�qQ��`x��6�`pE�,MD��R��o��������:He�R~�G<��.f��#��0
����� G���8�؇�*65�栕�/��΄��,�!�(�Njdw���U�J ��H�~����1����}x�{���c���B*��`�pF�C>�8fE�I���=Ip���7��#@�V��0�y�
D���}�7' Aj%Wk�+(D�u�^�:�cO������s�Sc;�6o��1��':��$v�k�:�4
�Ey�����s�ўK�K�V����y� �B�q�*�N:�p4�S9�S�|�.�ݬ�PJ��?��9�u�|T���-@�өEO��}���v�Ko����oz�E�͹��wܜ�����L;���@�Al��j��s�� `���ʵ�ym3�a�
(dT�=���A^����r��a"֔���h�H�%zvJxW_��{��*V�u��k�L���Z��?��a4>������8�KkK�k�(+pb-ux���7�p�nk�Rgc���~�'YN8��0q��q��8�R�0�H�#�ؕ�!��V���c�=����yb����f�E�� v{A
���*����
��a�Õ���b�m'z�J�uW������/�\m?->,WO|e����ʍoD1�A��"����Ruд.4� �Z��6<0��&��DAi�Y|z��	�5�Z�i��˅G襩�0P�O��3�+LNpZ����QXfXl*��l&��n��c Tt�v�P�� 6��A3�hj�7_a!�/��ch$鶠*�pz;ʧ���7�'( I�FWG�v�LO�u�A;���m�F[�������@��<d,�ε{�XV�灱�d^��X�2
w(�1{sǦ�oVo
ݠ$n�W`4YG�i;檰"A��}!�A)�����j}���|-|�kC�}%��"h>$��-��1��\�}��q֙�ڥ����vn�psZ�9�R�y�q�:�}����9�!b�YIJ@���mϕP_*�?�����O�BK
I�Fnn���8�2�,����Lε1�Ȋ��gl,�V�h���e>��$k����'$�Vc�Z�X4b<�^3�ʢo��h��c@�k�aR���ɋ�������[R��!�'�ڇ��}��s˙9]�TŸ��L�����6�vC�( * C#?D]G|d�+��4Z9@�W�_���"��x�����4�V������o/5>��+w��:2�$Oy�(�W��7X��������'1��lDA�7�H���"��H�I�m�|�R�������X�������`�od	��=��0���2���aS�=�b=�Z����9�%Vx�J���;����N\Z0);�c^Z�z����M�V��:�|c��M�����Q�����`lL���4��2�V��(���Kdl�:l��~�6��2�m~!�h���v�Af7��Z�~��c���	M��"�<�e�)_O:��i���>S~���n	���¾!3�	���j��b����A.Ĥ�j��C��`����w�vxG�[�����tI�������U��Лq�'S��������o���9Ŗ�ɱ�8����x�J���}�!E�se�$xs<�@�T�� '�x���-��k)ͦ�D�t��1�%�#x��o���;d��4�5���?�飪H�o�a�U����n?nt΂�w�A���%4 p�p�}��?�̎_���]bݾ\��V�����h�:\���7}Ѷ����'��
P�:�V�_Z�77_Ϯ�D+���VӤ�ᅛ%K�9��_� �����V�([9g󊝸Y��V�����?�a�E���A�.]�=
�퐘]�z����u}�͖�S��s��h�Jp�ߨ��k��]�Y"�y��75���=�a���(]�2Iդd�e�Y���x�5���YCP����A�r��T��pT{AvAZ�Ի?����.3?I�w L�����C/��o+���;�S�RG|g_$���H�D�ޡ���ˉ �����ۆ��I��y����[�����N%�M̷�E��O(�jnO7?	<uf��]}r�;R��_k=�
~6m����G7�&�_�Y�
z�+k275�3�'>�h$U��/X��5����Fz�;�J�V�ẙ�)�>�dG8��E�%k��˱�S	��=+f�4gm���}�N�ӆ)i'szo2A�<�Ţ�$e❩�DF� K@j7�"�R��50&�ش�$'��S�;�yR��ӺIS�0���������W(
�Z{z����t������I�a��ŗB�cH:c�	�����<��n��s����޿�c?3.�N~^O/��%�&���8��`
W��-6A��͜�@1xu��_k��S ���u�c���+i���q�cʸ�c;����2|O������]��`��c`[D�jI�]��m��'V�N9�ؠ��~��6�M�A����ХOF��M3M���������L�]K6D:��o�339�����YP�ט�����ր�"��ir�j��b]
AgÁ�"F4gѝEü�h_r*G�����zPn!>J|D���v����6T�T�B[���"�!�%[��l
�͹k{<��|&ֿY`�MX�?�yJB����,�$��/S�_X����p���`�nM����c��S/	sʠh�������n��_��M�b�-D���d��%�EH_�
���F�C=�Mw#@}��|� �֤�[>�3�]�"�8����I�L����� �)D��W9�rm�K�).��'�=��٧/�L�� �pGIn�W�0tq?�0�RPez�(�&oم��4�?k���9��ꎃ��keW�'̱B��11I�T�� V��Zo���p\G].��R�r�R���*�����SO�p�iy�§	��e�5�T�镕nl�ڸ���n؟��0�+X�w7?�;����U�z�Y�\X=ͱi�J@�F�2B�8�뿛ŉPn�ё�b�����ڎ�jb-w7�u�#��C��I]4�&l��ŤP���	k��u�B�c�:�q��95�g��I��4��%i��In��(��2��^�{3`"���b3f#�'&� (k�-ļ����Yx�Y��e��EX9��31��Nio��r�%���O/� C;�#01>b�1f��#5�iK�lT��e�-�~IQ��Ng�X7�@a���M��_57�i��w��gl�u2X�����h��q]^VW���E�ՙ*K̟d���]�dalEb�8��G�-نs�L[)|��P�]m��T��0EF�P��)�! 8����i����V��C���K�f�q�)d)��˲�ج��]zۆ���Y����� y�+����7�����|0Z�P�Έ��F�"�D�O�?��;HH�=��=gc���t��TP�y�?p�댋�������hoGaO]ř������?:�����U�"֊(���H�-D;�C���T�,��n>z���� ��&E����&
%�c��k�;N��Jʊ�}������|�V�X�D�*c����� ����;�X�A1#�	ܶ��C�<�?��	��If��K�y+(�I��L�8`�������V����H���o����Z�a3�kyZ�r�v�2�l�n�����Bۑ�J�|�j\����F�l��)��P1��qǸ��E}��վi
�\f5�i�[ae#���7�IG^΄X�2��GEZ���5�{}Zʜ�ʝg��LW-Bm��J*E�r��*�n��`:/�Y!(�]Ѽd��-"��{��wR�]��8p����Q/j:�>w����$�𫌘�	Dk�;�"�xw �b|�#u�u��eݪ�� ��v�7h�#���pp2�&���ZN��s�u���s��N��R M*!U����W�g��i�(��e�ɹ�&�(6Ie�bė�┶��}��{r��B�}�V���ܑE�rSP�r}���y�v�E�Ѿ�Ų,�1�:d����)Ay`2��?�GaU���ɦ8��MUV��G��.>du�=��a�+_�w3icWuϞ��
ۜN�O#q�`5O(TCꢌWzS�,��徜nqn���;4p��]�:�w����".'����3��H.��!.n�pR�\ˇ�b��bJ�5�=�����f	��i�V��lHj��3.�<O��2�$�� ��4�İ�}<b���҃}�~e�t��ƉTa�/)D�]|*�+Y�0���~lCr�-����W����a��x��
�d�:;�]�[�M�z�V8Ҹ녷�i�j�̖��H񀺁���*�)i���Y7�]Q�	��\U�K�1�wWn�Q����O��Wa$FB��=٩}O�F�yʒ@*���uB�ɺ�'Koʴ���A�W��x�)�S�y��~+cUQ���'�>-�©\�!��Ww�]�.h�hv��;R��3���}>�V����]�Y�`��1k:����ɍ��%�b�SrH�
e�ɽ�Ҵ<� lh6�3�x<��	�(���轕萋��Y��`׏��ƿ��I%yiY��P%r�ݑY�`Pa���L��-�q4�A"o^�̩@��Y�a�w�����41���b�k ����;��HW9��6��&��3�&���?��!�ʽY�3K9�����6�r�Ǟ݄k6Z O�H >c�m:��&��Z/�NV�j+x�C�u=��Z��!�G�4����_��k�|Tʸ����|��ˠ��hP�4�rj"�����dJ`��l ���2�ַ2��2ZR ��|Q�w���#�[��m?t=.+"�Fz����{�Na*�Wva��F���,��e쩬p*�����3>-x�a;���d���9�hB���^�h���� � �Bx�+�����s��nr��fi��,�й��Htl������������{�:&�M	�v>���@>����xM ��"��o ��r�YF?n��k��S��HJ?����U���Lak@4���UYv������P9��!W p!Uq��@�a�y�s�p��ߖ�#0���H��Ug�#h8�Ʃ�m��i��6�=D�X`	әS'�.)Z�G��w�*��hD;���i|�:ԙ���5�:���N����<¨}<{s/=�1�x�{z����þ��Ir� ۾���2��ߠ���}�kŚ\�$ΎC&����|"��n5cd9��]#Ń���[���'�N�B �]�я{����]�B@�	����H�*�˛�х�=�)�Kt��4��zj�h�����jN�!��͟�e�H����7���V�R�ݩ��E��E6���P$�$F��:���o��P��������{G�l���f�x�o?�$�d�%�	O3���jm���	i�c�Q�0i���I�oI&����[�t	�{
;��LvS
�{
���[����)ahn�����Y�Y��W���1�j����D��6�hۆ�=��$�~��@mM�(��7�2��˴�#����᳾���w���|�91�s��|�gƒ����o5(�t�-���#N���Q1vT�VkL�DX$}
�(��A�����@��������0]@�H��@qx���E��m[��h�h���%��b��N$��A�1BPב� ^Y�
gwL��Yp²<�=�?��p�s*���b�G}�}ѿ	�xYwս�F]�N�I��B��/�|����dJ�������N��EBO#�=�@ u�;\�1�G�S���=8�f��n�eY�L��7��^3������
�F�h�=/�_5e�AX�+uOL��"9����QNѤú�`�y��O�H�a����Eڻ��d��Y����Q �(�qr,C�|�@,<zo�L��/M.55�%��щG*Ld��1t .���R(�FZ>��U�0�����r���
�s�#���3�>�	a�7%������9�ؕ�m��,/������5���x(�*��J�Q8;Q%V�YXƃ �������0�u� �rv��TQ��r|��um3��֯�&F]�����P�*����h��1Nyo�D_��l�xdn�z��=� �Ⱦ���5�����59�bA�G-�EA�;����x6�_���5�.:��"�b�,�j��XC!�Hg0y�J:�Ȯ�M�k7ͼ(XM@*����17��^�MҾ���UK�P�ok�2�/��u$f��{��b�N�,��Ⱥ�#si×�ڵ��8ث�{���ߙ领Ž�������	bl��s7���M���U.�	��O�e���_���j׭u���{��SbS�n�9�S���u�;J�	՜&<>��̋|��;�0(�����ao&�DG��Vj�	4?#�J��Ha2ѿf<��J캑�y�Zpp%V�눧�9�Y귃ې0x���E��Z0�2�|��'�}�J�(]�ћ�q�+��Ԃs ��d�C���Cۂ�� �SD���� ��;l�faB�1���:T�b�<�*�+ ��9�6���?iNḟ^����G(NT��'0y��2wZ�n|jѐ*u�� ��H�����ix��ky��(0RCV����l���v�%_�e*����z5����h��C�z��p9Q�'���Tb�. ���\R�#�{��mf�����e7j)0�N��P���_d����{�`#�*�9��#�<̆�/��5����#衟��_�P>W��)\����<{��ƿ#a����&9�#ET�ᑧ�o��k_~���j��J�&:������jIug봱�!��c����i��0��z�����1��n�9>H,��g�k.H�'��dZґ��ߞ@{h�h�����Y�7v�{�d���]���I�Q��o��*�j���U��Oፔ�+��O�CY#T��@�(��~�[0=�n�0;%hXjX��.M[`-��T�u�o$��D�}Y�#U��,NU�*&"���˻�����7�]��>h�V�ɼF��X[!�sy�t����Hp��MRk:;X��n?��7��Ƌ���G������񹦉��sdip�B¥쌎��l����sB�ޚX�x7	j4�����p�D�()���y�5������8*1.bu������%a�[�a��?����Y&6��:�C�q��#��ɫV�Q�ʦ%�S����r�I%AG5>�9�k��Y��f�@�I/v��:���^�6�,<�}Q�J��<��N{7-�n�tPT>����Ď
�����R�����D�A��z�C�[�q�=Ja��?��T�󰯢ө{�uS][�="����%Kxr"���9jR�j�u�M���9\�k�q�G����zA���׊��F�;)��7�D�:Li�>	��q|��702�A �W}1kѷam�-s�_����C�O�	� ����}v��N0T��!6vW�m&�7�<v��X!���m#h.��,�����y+��ZIX�>��;��%�Ŝ �Q�?�2A��$�W���B��P�5�ℸ����H�m8y~�%^���Y��,sYr�� �@����z�*�� ��3�cb��+����h�hM_
���XϿ�x��F�B�Ǽ�5WT�}~�e|����^`=�S9�T'�lJ��W���ژ��C\x���h�8�H���#�v�����߱�ckӼ�j��
eg]z����T���
L.�JP=s���FQ<�U
�?�F�-g�M�(cJ�U��j�ߡKG�g���>��q���s������uHW��<��xt��}?`qҴ�q͐w�/֗Vjղ��0�;.��,���E��� 5�w	�v�0|�eS���{j�YB��.�)�O�{ײ@�x#��L��ܕ��g�ЙfL�� �E��~������������C�T��r8�*z�F=^ps�#\����)�ͻ\�PQ�̹ڣ@�]n볾}��*�B��>��Ce��~(
KM��x�&ɑ�6��l,53Q+)Ę�72�_�!�1r*Y��t_���]��0V��Ѕx��+"	M� ��� n��� �P�Fq�j2�Q"D��+��|41E���h�;�T��/!��S�W�5o���!��{��[�<BImJ=) �u�C�	.l`���Y���V�����V��OLX�X�1�i����)���W�W��ow�.���zg�i�*J��R��(jn4<ȟ7���s��31����߻Ro#+���,������-n��]�t�Q5�?Z��?F��p��Jme��bǯ�|�
W�x��0y*]�Z�Sm�,��	D[��O'�k���9��O ���o��_qx����׆	�^����G(�*�*�$g+��oS��!���VWUf�F��б�S7� �Lr�"}hfrm������CY�Æ4�"?�G'ު^���y�~�iJNe�eb�5���f4�y��6e
�G��nn�TR����vѾv[��{i�I!fk���Mǲ����{�f�)�V�N�/:]��B���0|����bq$�s#���h+�U�o�xථI��-L�7��P�wO�N;���炽A�\����_�D��a�۵3��E��Nu	$E��Sh��
��D�Us%5�43Y��R��������^��⃐q�/�S�H�mMM�
�>suc�թՅu��i��Xq�����R|:\I�tUt[:��R��ˠ���8�p�c������&5f�30a��w�t�W��C���d��G�p\�a�A��7�Ve?�&C��Uㇻe�M8� V��^�]�;�EZN��.^�Ay��Q`�[�d�U�`ᤋ��s�'�	�r%*��o�w�Q��k��#ڃU���f�u�u��/e�%EW�~��EQ�dj	'�

��rǄ���[�?w��@j� �8О���`:�Q�����շH2}�w��I�@�$�sNnqژQ:A0�:�
C�߇;��TX�׹,bio�Ofޏ���� Wh��j���E��*�YW,��`�r�,U�˓��uSI*�>HA	,T!}��˳$���A�*��'��>":�y��?;L��?���]�{{��� ���	��}U��������[W�U�d���qQ�Y|�a�6�Q��_�
u���B�%b��!��[SP(����c�B.<�IjU�.��`�.S�{� 5��n)lEF;+Z+� ɫ3)�E�}��t�r�ɌZ�) <A�V ��[���I��*��s`�⎚��Y^>�n��f�t�<�����_q����m<�1�Y��}�w����Ƞoz�̐q$5�5�J��}�5�;��4��:�-�5�@�;ť�B�CS����ˉ���+�ބ<Җ�F�������O�A�������f��ɹ�7&�n��^	6^ �X�F-���������؈<�T ;GK����N��A��Ѫ;$���[���yAhq7��9:��-#���F~��m�p�}��KCl��S�k�$���⾪���,���(���8활�Mg������߶�K&�Bm���U��i{�����\��.��<VI� �v�z�`�~-�A�^Fמ����@A�t��P/%����	�Lw����uF#oj;�GVZm�-�&'������V�A�eF�d��' T������U�G���s�k�(-���������~��.���w��b�>e���U��aA�A�oFaj�%Go= N��\��ݪ�R�0&����Db��������G1ͨ��&�J�,=V����(����[��4�$����Py�X���w'�SQ�M��V�W�K�p�?OBm�-A0źZv)�\�2�3]�T�C���|HL��	g8�]���q�)�o��t�5A\�>v��u� y�X�������5��I�?ࠛ�\�q�x�x�v�]����o^^���w`,{_��ԛY��Nl�N��=�}=��hT������y`�ԭQ]���c���]����즁z���US3���vܩ;�D�k?�;N�;��{�:�^����K��q�[�G��dy���؝�u��ibi}]�����Nʭ#N��ag�ܪ���;�,�'�˔j�������J��c��	��sň����ʬ�`��+�� J�_% �A/[�'��Ҭt>w'���D�e�>e�h���vN�2���M���^\��?��*����^s�L�K���<.kL��Z<��U��ז��X:{d��YX��N(~�3�,**�f��@f��}��O����@yt]r�p�g~�~JÝVI����ce���y���Wμ�{i��Dz�X������-�.{�Nm�*_�]�:ϼץҐZ����.Y̱��:��} �*����!��o�)�4�0 a���`���4�QmפQ8#�"��P��dV�5r�ם����:�ҙj�y�;LmB��J�z+��=��zn���:i#ΜKD	�6��5S����5��7� ��I�%T0�ÚE��-*�ˎSu�9�&Z�7���������	�0�� ��b���62o�������|��o5՚�'cGO��s���J�g�<�ʒ�� ��.�ݳ�ԯ-��K��)]�: \��h�I��l��ch7ِ��I�x2,��𦲺��vH�����kj�������5䣵��}'���O����_r���ԯ���ڟ ��b��Xm��3��Ц�	�6>�v�<�ɧ&��N��\(5^�14�V�=r����|�N�y���� �qh�	,�rhl2S�7{|��ti������8�*�W{0��}h��Cb�0�`�j;�~0�0�b؋��9Լ*�$%���Yߖ94:_�p�h(����?�;�]�b\��8x����T��[�X-�Ʋ��w_|�ϑ�?D1L����d��Q
8�A%3��7�������XE3	�O�m5bNnۖ�ωLqL&���6h�uʜ� �'�]��j�8�&t���
���Sh/�+e�5Uی?��1_�j~O�I��uьyiq�]ܩ_��i�)�J�n%���lw�U;�j	� IGPJ�nօ�����3C���;�${�^D|�g�����챈�[��P��1��:'�'�	3�2���G�|�`��^Օ@�ml�P1ĸ�}���}��V嚼�C:�_��5���HO��q�I;Eyu�v*���;f�&g�%7�fq�nOE>���Ʉ�P䝜�j��އ�3�do&��3�ev-k�ّt����S����5�Y��cœ�˦zs�6߱��he-퐉��}��o�QѦ����?�]���X֧?2��Kú����"�WBf�/��>Q����2�4]�S^�L���9�4�ǐ3�k��?�ڹ_Zы��һǁ�52�Y�=�,UyM��9��Ze}M�\D:���Q�I��U��º��
��v������|��࿆9�1�i٧N��m$vX�}���MU"�ƶjc��֙l N���ұ<�W�m0��;�~3ʚ�	u&��f���~���w�g�w��l��ѓ$I�µI��V��Ia��j�s�@K���_NVW�J$`��^dr�2P�R���H��g�ǜT����'e\��
�3VC���=ՉQ�����2x�q��I!�i�S��B�Lu*/�L)+�I�X �D����ʴ�n:[���N�aN/�}��2�8k�J�Z�'�j��:�5��>h�)�/*|ԋ�HJo�.1�Ŏ~�=J=�k�9��|��������UY�J�Sڝ��V���4I�X�s�V'	��dX�[��{Nr%E�i>��D�}��09�t���9��A�����]X�1d�q[�9ʉ&r����!��{��97cW�rJ#Z�}��Wun٣�!1�vJ�bQ,��Kڭ���-<
��O���g�i#�O� (j6�Zs����%&��!Y��c专���>��1��/W�.Ϻ�C㷒z��0z��bcGr-nL�v�3@��/n?�j�����" ��D�GyV�;��]��F�/���R�gd��俲L��6[��I�pi������VO2����*?L@b�WdG��!��o���Ԟ"so,�LΥWI������<>���}�`��u�@f����h"p��O��-��H�ۺ9���-�(m��Faaߜ����?bꦓ�o%������;�%�W�W�CV���Za�f8X�s�/�ص�'�U��'%VXA%ҹ����EE���<[a�����u)��M�[p���'���[�JM������Rn��;�ٌKJ��{1���@���r"8˟}����N.P���Ž�Ɔ3s����ma��w�?�?
��s�-;TmX�O9e��5N�j<�]�1�������!�K��?��,H����x;e?���6�P���*:iw���^T�̀&>Cu^=��_����n)��K�Fok��;��H���8��b���r�fXw�����q�t���2�ob�K^ZE��z���&K��5�R��� E����[6˱Nq�6
���b(,_m�/� �������Pq�_���l��c�Xq�!�mY� O\�E!z�	~��^?���P��|2B�|�=��N1Ӝ}A$$��n�3�E�N��C�T�b[��R�,���c�~��=���z����ʣ|\Q�XO"dt�<���>�X�۰K��2���RZ�N]t��5��~Ei"�$�FZJ1��"�-�a�]�cع
iS��έ^��s�X���;u�Qy��j���V݀�dj��avD1���zG��1\/2�4*�"�=y�S�)�����'���|�������ڎ,�Ӯ���M�S�q}�1;��S�7M�#{5�{mv.�jbk�Q[�ښ�k�"MXp�~�{����(����@BfVZ��1��@�L�yq�a��V�k�nE�"�:�n����@�Z7����܈��=bw�=n��g�F^���*�Eo9��آ-b__ݱJr����:�ђ�4j� �-v���K�M���7\� u_��o�N�͉��Ex�j�eE��3\��KӠ�'��fU��Bݐ=ɢM�4D���xPC�OfL���
a��f~Hoɉ�i`�}?욾C>�GJs+��MޑD��;G�p�L~5j֡l$�����+�	4X�W�K^�h�����܊�#�y���2�>B:��K�x@v�"V�1akc����9�\mi>��4�S���Q�ճ�PS��Z������4 �Pr����#\�x�
�[K�=�4]qل�0�}�6������-ǐ����ǎ�S�l�es��.A&�&��ri�ѡe�5�0J��u�}@��y��$k��5��Ms�TAwb/ɻ4�|��� 1���uv �_t���Vf^<��������f��yC� ��O��˯��e��wx*6�h#C����
�>
��	Tf�%)j�wAʗ��e8ܮ_n5|��Q|wUF���]$⋫.ȑ���6���o�C�wi�����S.�xa���}p�'��_�_9y1�i	�+�sݝGN���Â�i�T��y�����h1�u�������2�t�����n��jk���YX��VByL}���n��������⷇�"6L,H����KF��6��sʚy�G�b+���Qn�uH"��������:��gՁ��#C�OZ`��a�9)�%3��S�
�a�}�S���<J��6"�>�����?j%^�b�����-���%��;j|�� ͹pS-=9��$�>���BޠO_�Xѯ�jY/'�nN�?Q��0�;��fΐJ���ra��8�w#a��J�ez�z�c>���d�����\�TjZR��l[(�5��D�FyР�9�&��k�a!�=LT/.�
�Qa%�fҽ�~"�7���]h���G�~v�r�+?��()�n � ��{{�se�/-����:/���ZpO�z����S�|$���~�'~��[��N�
�#TN�XY��CK��	�R³�q�0��n��оu$�����y�9�4>����O��]m�d������:�����[��r�F�5l�g�����2�o�V)<ǧ���6-{�$��2@u?�H���!���{8�d�i&8'�9����"����W~:�w�;����	)|��*��U��m�pc5�m��U��P�C�7.�ޅ9=H��ֈټ=&m��~8���p�d {<�y���������Bw�FP4+T����Y�7g��M$����?٥dȠ�Ak]��O���)�a���K+��Ý�K
Ҩ�鮤�J:|��:�a�AUv��'|�}��e,�iH��i�� ^���Zs���=u�vQ5��d��Q�Z��C�f+ ��ɀ�x\���B�y��H���l��d�;1��$�s���ut�5�7(����m�-�hٜkϒ��}%�r�Ȭ/?��D���P�����H�ϳ�����s,�b��mu&�X��#�� |��_ə�t��W��_n��}Gm���q/�$$�Hq�lLMu����'��$�CԒ�N�*�R[�K���ŉ��u���l �Z-���C�*��f����R��F�2j�"9��f�� 7�A9�� ��>(QМ�Z�B���J��O���g���i����Ʋ)�o�,[6�%�z��7����%���0���%����@�$8`6|��l4�Ql��t�����Yh��#߂SI��v/duf鏧���͸��w���/@��Bo��=�(ė\��
I��y�u�
�#�g��w]V�D�X-a�%��9���G�z}����Ė��� vV6�0�ψD�7����V�ʨ�n�^�h���b�ی�#�"��Q������y
T�Ϟ��׬՜�p�)@����Q�惱\[4Ǭ/�W�H\0�r��k훜��8����c!&n�o��u{�7�Gv?cù+�����߇�'h�!����A>�]ӵ�O�Xӗ�1h�z�]
��p�2�	�w�T}�,��~c�fp�gׁ�2?Yd�Hw5Vdi%u���6�
U�����l6U*�銥����:�њ\�;�������^rW@��V[��U�ڳ��U�5#d���y]�+���T1��Z�Q�~�K	�9O�� Cy����H�����Қ<������d�J��㈺t��X�IE��n�	6<�I������,6�����&/���-'ӗ�F��|�+�,;��;K-zF��;ºF,٤��AH��Y`�i��s�����$}Ȩ/Z��6q�?n��5\3Y�ٴo�����z�����/��y�����lp߹9,=�߾SN6I����;��Q]^��n=�:��D�������	���Gԝu~��03�rZv%%����{+32�IGnN*����G��W��)�*�,��W&3�������(B�zt���N,ױptNE��K�n��/�:^"��GO�S����$:��)��t^R����Y�I�(��m�&���C��E'�o_�-*�H�Z�H�/V��5E��;��Pn\iQQL�Pv�' ��Wn\�~N�7N�q���2���݉�]Ǌ.O���5���'<�|��E�>�Ky����Uc�&�����`���\����Y��$��s%�L:"ԋ����g�W8U�<��k��i�F��<�s9�����tl�b�lՔ���ڞ���lC�}�'FU3�k`�6����N�RffW�,ǻ7�C�G�C�^�Nn����6�G�2��;���'�LSd���m1RL���h�̨;ƃ� ]��"��&ó�ݙږ�cnl%� k���X�q��4�D�7c���	-�"�S���I��"����)�2����f��zu��7_��
g�.j��,���s��I>��+g�Bҋ�p�~�^��,e��뚆{{+�\�ؘs�{ux��Ӱ-�Z��eh���~^�k�w�Ң<3rD��Օ)�
��=���H|�Y&���ۭ���[J�{����u��0�\y%f���b���iRO��G��4 r���ݎ������yQ�+_����#�{N�ۊ����3�&0��>,�O��O�^��7�{�>��4k���I�n����{������qڔ�$�[��T� ��8݌����S��B\���,@7��&v6Nt?6�t�o�2��y��	�n�"�7="��HՋ��.��NR�W-�LCҕ�g,���9Ϝ����K�K>/�n�!����8��+�Y�-p��?�3{0�_e����q�d��Z�����-�|_����A��Kb�Y��8�<�yN��BeR����ֱ"����Yl�Yզ�i��'}\�&|����3�GrP�c���:�H�T�5_f��'�A�:n���j����#���I[ܲ�Zd�\i�:�yA�ᶯ-�	��4Ѭ)��1)s��fo�l3�Y-�J)�QѢb#쑑ɝ��3�l> X�A,>9j��Ok�^�!!�ZtuU�΢jof��Zc���_�o�ݡUf�� �^?]�Q̣~�P��T���3���!�ߝ�
���\�5�zȊ}1����<���s4���T[�ݬMҪ>x��cv!��1�!@��Ń�F�Vx��[Cc
[�X��ܳc �р@���wq��&@b[C�E��aE�W�����#3(2(��g?@Ya���j�Y�T��|��q.�Q�x���⍢,')�jA���v-]��\e �NZOɚ@�(����
(�,v�=��E!;.C�ܟ����ܢ��]S����P����˜��]*J�u���o{U���ټg~݌x�
�($�@�^�=9�<	����8���^1��'�k]�y�.xi�&U>m�K��\ZR���~�܅�����39�-.�߈�� N �'�G��^��!�av	E�@��7��s��iX�IĮ��N�\�����q6L���8�=x>�+�F��5��Խ�Ĕ¥�������؍����R>���v������@�Â������F4��#zH�^G�^�?�0���J�4h�9�D֕����)@����w����Y,X0MtW=x�S$N�_Is5�#�]�͙"h��Br���Xx͉�5E?Լ�rAJ��c�V��+����.�ɸN.��E����t�f�f��>.�,�'�&�t(%l5���z�՞Ƣ�����%���u<ސ��<�q��㺓�\r��"x�'��H���܂R�4��"�n��QX������)Ll�&���s�X,RIg�P��O�J��l� ����{��*��Tr���N]��l����Q\w��f������X�ی��YT��șQDo��C+�#s�f*��Wѐ�8�<,�y�'��a�)����<}�����ӆK���N���(Z��?,|�?�kL� u�^L�|I.���˰�ST�jՒb�����<	���f�1r�� r�XM�	�5#E�p�K�����k�Du���]
����A���F����;	��B��|��?k5�Z��EUwVw㽆n��WK>Fc��AR݂t��Y=�6�|�pg��4uL��`�*��, �EO�����Nhftp�*���Q�a��݆eoR���������]������;y�$�Q��H��ٝ�#�Y&�kS���ϓ(n,���=)��D�~�"TX�v��kG��%Y��� @�ڏڧ��r��#�Y�u| �ᨤ���`p?���t��d�l	��d��5�^��!�7{ȋ����=�\�}o�GuOvqs�:��Ƿ&=�k��h��;���m� +% ���pK�>��֔*��.�c�I(T(ȱ�7|��(�Z��b��3rB���kY���@E��JP�m���J���Q�4�N�d~�!��̜�۰QZ�<��ĝ���3�����<�{���ǵ���0 �$iH� /����PJy�BC������6f�:A�M� �_ui�F��@g����|($Z��7)�����Q����Χ�j7���ϕ�
h��5l��ۗA� � mK��6H�QǨx�׎:�Bp��� ����="ۗ3n*��V�:]�U�AIj�X�.Ic�8�-�Y.��#�8^�伧cz�֧��=TK%,O�%%���SF�&4����zڶ9[ҟ�h-�c�d��'߷�2#X��i��N��eZ�P�՝�������c��v��2&�ס.5��˔�)��M=a,���E���,��!=�+�CF�UЃCset�ujk��Y�>8a�xUǃV�+G]6�{Xv�����
n(�tpu��<���_�L��;�Q�ۼ��)�i��0J5�3	K��&xJ	�K��c.q�֙�T���jV��!w�2�����Cg�o�,�Ѹ�1q�� �/0�F�d�
z%M�27�N�{k������>�n��G��� B�?gҰ���{N��q���=�Ҙ�OnOj� ��_ZB�_�_���R�j��F����>�k
[�e��ud�ڧj�'8}�$5-��뿦�WNOO�YfBp�� Bh��s1�+�rt~4�6s���w���NQ�9�u���4<���L���m��U����z�Y"�E!A1u��Soh���}A���"5�������I>h��^����x�( ��.��w����n�������o�nV��4Aah�:��1<߹Y�T��R	H������O��}ۑ�ڀ�(�w��,�?�30Ƕm�MH'[Vyg��ףbQ��iVf)-\O^Q�ޗQ1\f��uߏ����G��Yy�6�y㛮%����
(�;ٲ��i�$.�&�	�t#�Ҍ~l�%���1��ަ$��=%�5�*�o��1� H��q��9WO�u^eum�3�,��FmY�+�%��t �9lV���"Dv�wJ;���+~�0wt��=՞C說#�@+[y~��u��R(�@Ą�5
snΆm]x��c��bt��`���vn���e B��%�5᫦��D|���X]j��V��[R�4z�\@x���؀S���~6�� �K�}�'[�����u�� �����������N7-X��;�B�ͷu���V���+"�K���|F�#�ȳ�%��cd�k}�ִMΌK���]bK�M%�Ғ81�k��S�S���|���F�' kx.�SӽU�����@�^PX�4]��Ot�P��LOWf��M��hҒ�EESk���;	K�bT�ހJ#r����d��!J��>���)��f��!�~��Bc@?�N弸|��`�y�����߷�(�~�Lmʀ�1'����e�95s�|T��6`�ut��'�W�48��!;����M� Iu�rҰ��kB��}�4�a�u ���)���ƶFí�e��j[�����~�Jqi����l�3�'��t��X�j��i�x��U5}���9Ǘ,rc�n�y\#��#�k�9���j��/p��@���l�P������ ��������̭	Zv���H!aIB��%�����Z�8XN�E��\�:1�߉]`��#f��ƽ���E|A�s�t�ގ<=�C�_���uu/BשHO�n��������$t�=��,�E|U_�$oX@��##���)�L{f�2x`y��7��[*K�m��/�28�AMg�%WA���p�I��Ѭ��=�������2]�W���N�4�;6Aj*�"�+.�����=v!��}Vh��x&�jd�*�v���4��$�u\0��k�ëh���Q�쵡C.���i�/=�M�NN��f~V�b':h�I���Q�E٘��?��] ���h�K/*ʞ�b�K�be����cES�{���Z��ps*��:��`�{ �(@H�&�7�@�9�}zm�NCN�Dy��X�M�-���|�.�z�d"mC-��d�m����̎#��ⅿu�'Xl���UC�r{1�ق5zܿ�����Dw��J�����@A�����Hݍ��iP'���P�}�p��D ^���x�x5�Ta?���S:~����Ѡ+� �f�f뮶u�'2� {��ǎ�K�H�R5��@1�0C)�5y��H;j���~xF�&R�W!X�H?�������*��k;�\OX*f�Ļ�ip�4xE� o�\����~���_x~���$��p�sp�Q�}�[�pLu�A��G.~� 賆�q-RTG=���{K�(�`�KnKם[�ɯ/8Ԁ��U�֒v#�l,��lM�3w�|��3�}s)�Ʃ�Н}G<#_̲O8|��`�r�!�> Aҁ9�����8��eo�!c�>��G��$��|��KY�*���JH>�K�T�_չ.m��~nL���4���;��'4M)S���",���c�^"a]��X����t�:
�O��M�8[��[�,n�E�W	 I���7�Xs����6��A��K��h�xܣ��6�iŕ���8}���̗E����
K�z�A��m�B��H1�!ؓ�-/x���ۉPջ�+�^Q�V�4���§C����G��h���ȾFf�Zy��Y�@!��d)Q"
^0C�P�b]�R�%uN0�<;�
v��Y��̾���j`쭪J��;\���*:����t���z�'��D�~�C3D�/�P�@7�6{�S`XP����������>�^R�>V��z��S�.0"k��͌0dZ��K����5}���4)�Ka��R�����ۃ �0�B8���ţ�.wb���x��ZFP�*=r�m~0�<��� ��%�4բ�ц�Tv/dw{;D�oKl���e��}3B�x#���z~}6�mo�g�����ά��U�GR	�
r]��GR����{c����}���Tip�� �$�1.he��կ}�n��EQ�J㨝��X�j:tl���\�`��n�d��۾�j���d�rQj���mݫ ��U���*�2�ڡcs�.��-��=��%��f�=�ƷNz��qQӧ��H�m\\7�BǓO�{f�	y[,���m*�:TE�[�x�5i��T� N�U�Ω�%��O~������-C� | ���yo�ޒ�n�eˆ�>ƨ���$e��<���m�����R5O�ŏ&��l���pf�3�,��"HR?=���~���� ާ� ��w:��$�����+���	����B33�L��^����s�(�Czp�}�Yˇr������T�R�:��u,�S�"�g&H�(�8��!�o �zD�;x��)��e�1�����6;mʌi��a~�Q aB��Wʞɓfes��VH�jC���Y*����N��J�H=Xg��g}����V���ۍ�ᡸ+���^ ��Sd�𸤻�� ¯<D[�Jf�{A�r�.ݛn���A�ͼa��
�W��̏��� j���{%B��6�� j����X�>�P��,4ٰ."��"�v�$ːoë{����	�v�+���	M����?��:mey
��?*��3i_W��E�3.��(�.nR�`�#�	k��mV)$��}V���F��Px�^8�GQ�ΙћC��[|�L �y���P5Ud���/]>��� 2�a~+6�E4�3�=tC��A��8ʱ��7ݎeǧ��z��+�s�2W�fMH4��(�"El`�,�恚2x|�����I.�|?���O:�.�W{˦|�-���x��[�ɗ�6K;�B�Ֆ4l�_N�;�<���-�t>�cճ��5V�����Y�|E�ͻh7�ʌ/,(j�y�,:�ℤ��zZH:^��������]HRH�r*���Dƕ�~�>̦6F�sN���T埔�u*��2������b��
:��3pݔɥ��G<�Po�؊ +8/��c$�#m��g�Ip���m��3Ye��?Be��y�66@]�V�z����,�����2�}<7,U��-g���t���HV.Om���I�V,8��1��,��g$� �~�8�cV??�)G�؂��+�=�R+Q���jFޥ.��G����0~֭h����+��A�Q}�_�Q���Kq/������J���(|�Yy�(r�7�6S�I �*K��:a7:O��	i�|C�����p\-D�2u��&�j�o����0I4kæ�c��ê"�+<�����#�@�/ =ȏ��vlM������u��1�������MȺzXuY1ET�[	|~����q�E�~r�,[����!�O�T�e�=�pf���]M�`����Fs�J���ˈ=�J�
}�{��1d�oC� ���-�q ��[��v�-����I�F�@��N�[��0�:i�ϧ/\�~3B}V}��X�$11+�ҜKC�p(N��٬@Ot�g#�_Ȼ��b���֡ż��6s���1v�P�k�l2/�0�QW��ZGUd�GvfswN�U�q�Ѣ�����������V`N6��L��
4��![�<����������ܱ�PQ8�Ӝ�ޜ$Ng����j����������*��}����%F�2sQ1��H\Be]Rn��$�|MJk]�ít����ag"ڣ���&L>K�pL�����ť��K<�2u
`.�@E�|ޅ,�ܥA�k�%W�1��5�!Ў6����W���g�y8�$�:.����8KHB���[xjݹ�7gګ*پ���@����3i����0���"�V�T�B��,H{�ZP�n�ٓН��o��٢�[�75�5����c0:�:-+�ݍ�͖Jb�6��V�+�;3)A-6��$V��"&-���p;pFe���� <ҏҬ)k�sHZ��A�H�v>)�|��X��bɩ7�; bʞ3,�l� {{�#�ޥf��%t�՟�id��$+冞�%I�_�S٧��o�X�s�:����9
�����������B�j���4���}^8��[ �΢>	&W�lՄ�����O��B@~�G�I��-k���6Y��T���N�(SÓׇ0Ɣ�+��i��+�	���٧�A�2�B���v�Y��ucS�tXP	J^ˣ?���ydqxo��Je�<��$ ��>����63����4���l�������:b��p�c��X�G��?.Vg�Ou�ޒ4.wh\�=0�I"�܈󕕙	op�Jtd$:w�x�H�=�%>can
4RmlDi[�����"?��\
�3�3g�6�9��ϟ�2T�M؆xD�!�'&��x*��
k�e���DH!�#���/d;�8
'���a�h�����O��ճ�!f2��^-w��׭�w��*T� B�����o��~[�Q����>᷁#��𬲎?đ�QI�&&��r3��&0�n���ʙ%|�Y���7RG^'XL���eH�sx'#2��i����q��8}e��w��?Q-��n��>xê����֯�n�/�R�B|w-�b�sT���Go�,.��4���&������'XGso��_Ll��I4R���)�����N�	{X�#���8A�ěz��=��A���1�TP�̄�iVq�(�b'm���#����;��Ľ��OsO{{.���Nt���H׿0��iW���חBk��5��a}�K��\x�����#t��P�+4��,7y��)g�VSAQ��$�@�OkT���1��#	�j[���N �R�b�_a���,`,[}���%��֪ԛnoj�Ŕ}H��X\��lj�GL�x�Խ|�?�@e\���"ۤD��3B҅�m��23�!d��Ŷ��M�f�"�����bLz���fNu�7��3�Tl���k�
a�,�Z>�&��t�./�Kl�V��p#:�<�}��.�v˒�;�!O}CKo�͐v0�
r����8t�:�5W�BH<�v@����,�U�c��4��#g˙b<#V ��?o�&"&�2:�,��<��r@k-�.������ ���`~eJ�%��*8}䁨�j6��U��j֛�Y����ǳ�aj��A�����&��kd;���!��=,�����}��7��'`��7q[�k��[Ha�����G>. |h�MVK��$��?��B^,L�\�Ƽz���� ?���|_��t>n�WΫ�K�^5���d� Bc	?�C���-gv6
1Tg(���|�jg��烛�`��P��yn�	��,�������{�m�}�Kd��b�q���R�L'�+]I�^�~�;�j�la�G��p�2%PX�:k^߫�߯q~J9��^��� ��&E��9�tM?R���޸6��1ͿK}�VW���R%�eV/�P��V��v��b1�e`�s��\����0;���Jޘ�����I���:o=�R�$7�ڎ=�c�9)[��IS�U�9đ�1sj�y���	��G�����������+/ZoK������[�&��݈�`�r�|L>o�t�蔄'e`i"��T����ܖҼ��VR<u#�Kdx'd��y$hxF!'�'C�Ժ��c$�9u �͸������g�dx0~�����A>3>ȃ@�� H��s�=��i3�[�q�����Ο�s+�~7�EB�*p��*��> {�ێ˦����X ![��8K9pk��	b��7t��L����N�x�.�_&�/Q�qܙm��	���h������ HK��o6����D-�I�i@�dS0Zރ���hS娚��¦�be��r^
d��И=!ʫ�� x�~���뀔et�.~�:�s��1/p��Ӓ��u��W�l�
T�U/��g�w��R8|n<�%�#4�(\}��p&k/�J�$�Zo�kI���:���A�ʭ���(rg�.���:&�@:��۱��_+K�-�	���;o�<e��>))煬1i��aӳsY��V��]W�?cWC�:���<�[v
�?��ۙ�O�zFc~PG(���B1�A��AK#�v�;MRia<������P#�q�e��m@�N]�yM�)���S`,n��g) �^���T��ZR}F>���-�`Pl���n?oё�5N��	��{���9�g&�T��I��O3��#�\�]
)�=���������q���A�����D�A ����ahϫ�=���u¨YܧK/��?I�����SH���\b��m��3p�aD	]��p��j���z���=ͻ��e�7�k�S+F�D�����T�����lq�(U�4���~�D]����bv�v)Gs��2�SI�8�A�Z�K(��\L�y�8��T���l�n�t'�$��]����!B*��[~z�˧�FɍA�'�x"Ƙ�pJ��*ȫ����G{�z�{��7-b����ݲOe3�u�����X�,���ķBb���v`�9�5�����f��R�	ܭ:]�{G�2�>4�7���_�	X��g;}��m�����U�����B���������8͎�Aŝ��BFt�<]P���YC��E&ޘ�����h̊'��UF�L���Cw�nO�t�^5g�����g2��>�?����{�?:��j�ͼ�>tc���, �)��Y����?��fX�NDk=W3��&�[�5GY�.0A��LR�<x�(���b�tvOt�8D7�'���M.-��D�-�� /j�3�AU�$���������g����ǥ�H�zA�j@4�b{��6}cw%u��_쟤Ua}2n�>&�%�L�5u��N����ٻЪhG��|��HE+m�ڔ�,7*y� �r)�7N�Nݵ筻�)xKKd�x�s�����/PV.�����=�3g�� i*�#��l�8|r'��d�h��iz�5b���S�g���Y��v=��5׏>��ߛ�W�/�횝�׆�U�;l�����k­C�����h���xC��ތD��^�q�T{�X�I7�sVZ\nmX�B+Z��ҩ��%�d���J��7��k� �b!��XQ|_/�����|�<#<�2F��EQŗj�|�j阐����w�g1�}s�M�Uhj,'��|5"�-�UO�¦���J6H�4R|�'�;e�o^�
@ܬ�,[�k�sh��ͭ������JH]u�=�ާ�l��ƙ�c���vw��$� W֍w�K�W�c՚��|&ږ��5Q����A�����J86�V�'	�-ziVR�b<rS��f|�ڐ�槓�	B��֯	���&�~����y��i�#�!>�t)y�r4PE�Ic�����p��?'ME��.�$ >_��!���}M�R�X�j�|��U敜n^�F���Ԑ�oh+_Fe�:N���=d��']4�T��1NNٻ剝���PS������n�������o��NSb�7��xf�&-�w�����)�/�1(ތb�H&8Q�I��=�ݴ��Xإ�pu�'��ˬ[�8�ט~��bz:��&��Փ+K�%hq{�
@E>ws��2��c�_3��̊�;,��H.���AP�̼��;:�&]ǃ�*�;La�yH&g&���p�,�.�� �Ͱ���?NFnfK�	3���y�[��u�?(��uLZ=�N<d���G�8o!��|ǀ�6��t��,��>]Y.��Z��C���7�
)<H��U�%d;��o�uC�_ɽio�3��PJp�h�VH}�����!��A5������Aw��y/<��r��}%���jM!��;]���fvg�x�,�q\w��z>��&ң��ԅx��Т�`-/w���	�t�7�8�>`0*[��	y��X&NS�rղ�p�7�T2}�B�l30\����d ��bָ��u�qK!����Pc���_��V�ɬ�6�Z*��OL�ZUS��~=���z�B$��
GR��I���ꛞ<
�~d��J�b��O6<fx=]�:||D�j�R`��v��2O<b
bPU�Ӄ�hC��u[�$�G\�T�FEh����(�9�x������ߒB��E�)�E�P%�^PLvث��t�@�
71Z/1�Z�.�ӛ��ɇ&�)��6ܞ�z�Ŷ���v$0o�th~uvvi�6(��p����]�MzL��+� Q���W����3����S�����u��/����Y�g?���\k�)Sy1%�G�g��lz1�D���$��de�9�nO��.y{���~�#'��(y��"NO��7$E��6�d�H0��y��������!�p�l-���#*yȀ��ԝѹc\_�;1܁�9�*�YF-��:��hoީ�;�ZD���L������~�kϱC����:�E/V���[r�+%�q{>���z���b����fK�P����4m��ijZ��s>���]A����{� �fg)I�@WHE���Cۂʆ�oa�O��ҤEM
Ğ�]��қ|z�@�]��p�R7p���Yoɴ��o�	�㲹һ��P���c�wM2��╨��s��#%�F�4�\H��.4��Z7�;����ޯ�3"8mF��0�ƔW�цI$'H����4�.��\���'k5�v�3|#��s5�}�l�SӜm�r��L�i�<�[�:��<�ߨ}����{����D�����3�{h�,V���H�6`Z:���0b*�ꧬ?�>��7bΎK��������)fdè�L�Nmǈ����[��O�x��b͇�l?d#T�W��|Yq�y��|n��7Ii�E�'vt9��¨W�̈#��)pӅ����VK^�%V��j�,\�Dh�|���5w��I#	��j� ��*��������!�c�eV{\����*;A�1��:���/�<9����a<T$�����.�E�n�E�IX���~K�@|p����u�}�Z�?�fy�S�:��0�ޓ���W7RZQ~�GA�Y2+���|�j��H�@�b���G�O}����Y߂�N��5���tѬ��{MA�������<�-��=������������1
�L��W?4�^��������̳'��H��!Z�àҒ���d�d%k>;����gF�����"8��s=6.�͛�$'��<��%����e�������eǞf�q�jue[e-�d
�?S4R���(�C��2"��a�j��d�R*E�����R3IǮ�;4]�8���� D .:2�Iqd�.���x��?�����0"e��6,e���bn��̊�Q����R>�ptY�Ȇϊ��g���O�e��xa�&vk�����M	��+�Zko�EGU	.[|U۳w,��n+�_ ��ٿn�nvZ��mMt�I�w�oC�z0��ɸ5�=bvŔ��Z^[ʖ���b��;���Kb��Xk�W��;�Y9> Y*x����)t�'�6�WwX�����Ջ��lp�J�V����b�/B�}�^�1����)��H>���~��"���xMH���)�~�
�;��m�{��ى�]���St����1�@ӏL�������nI��L̅�Yo�E��*���:�����z2š�N�*�*,�A��{#Tk��e� x�~�a慇��d��3UbL7�q��X����d �C^cQQ�L�4T{H�H��� έ
=�̩��RA��?x�LD��E��qχ�Gy�kk٭Η+{Ut`�q��>�B�\ͷDV���n����X�#29h�S�.nhu����x�ՙ�~Z�a��E�/5��J3�@�{�B��
zC��`r(�����Na�4�rMxE�UG��ݴV?�;��/QQ���ҋ��
����ڸ.Jk�����^�iá(�ɝSk�s��{���wԺ�Af通����_�T���J�t}����%��������E��w��)��4L!�?FON�aS�QeO��	g�.1�=�n���88lr"���ObK�1mXu�s��q�gC:��V��bo#������;S��8���n���M%�L�rPA[��&3�M�z�����B#�2�i@��rVܹ/W?�g�����]ܼ�bs��}oi��Y�lH�+�"���4@n]Zt-=W˓y�nw�n{$���WC"Ŕ��b�gh9h>"����nАH��t�����,ͳ����p6����Ҵ�%����{uirǶ:~���g��i����D���r�� ����Aj|#$�;x�<��,�K Ƃ��u*p��v���%)c5������y��o�0�7����B�q�p۳�	I�X��HEQ��ݕ�St�O߇c`�6ZJd�p�*ΔߪD锁��_Ӕ��`�8�i���ȶ�,��P��הpLU#�Oଉ>��y�Q6��ٮb���/���&֥�~�Q����G}�hP��A�v;3��>煯,��`�'c6]A�:Cی3�l��{b������`A{IX!z���ۮ'`�z���R{j!kC�0����9�	���ɍ�(�C��>/�p�����ܪ������z������ �E�=XNa�# ���q��u�hCe>FPX�s0��ͤ+�)^���'�����D�CYF���/k[\��>o<#z�Ol#�73�׀��G6
.����ڻ&�m�`���N��I�����+�� WM�8���Z��P��+�����[��8g�T��*�߃���3��z`���Y����7�rS�|=�ъ����0u�&�_�m+q1-t�����0��z+���W���T��(�R��m��1���~f���j\'8�r�V��4�e��Z��X�&@����"W@��t�$�-�X+��~��`�+�>���CtȖ��<���^��0����*;m��Lۜ ��H6j��(&�:.�����iᣖ������:54^�����ȗy�eb!�Iz׊^�Bh����{�X?�7�<i�L�h9uB�t}m����L�s?דU��M��H�ፘWj[t�e�Z�!M�z�*'�wy�bЎf�`Ta�dG<�S�>�&�gJJ�u~F�	��):;����'����7�kM)_N���'�@j$�bV^8�)�F�����:�\���dp�FX��8�/�J=�� �Y�im����oϘ�;�a�Du�e�Lt<�2�;�RONX6f��g�:�B�gv��^3h��d�%����]���@c��F�FC��]o-��H�[1�D=� }~g(�sF�����x)o��u��l:F����[�x��q��ę4��2��՗�o�NG�lۺ�	Z%���9_�/�W9uqa�.�'�Z����o/�Jx�#F��A�RtX������+P8G����,�%Z��w���IIw�e�g��q%��>�;��-9iV� E��b��a,}�;�K�#ϓZ.����v�z�#z��A�L������jh�Dӏ�y�l[[jqf�}��x]j���Et�N�����¹���f�MzҜn�S���8M'�(5�Yx�ӹ���@	����"�c[���t��!ƣ��zt訂�qe��)���D�O�����e���j��ùP�!��bFۯ�p
o��j�����I4�~`��񩩭�6qWƵ�-e,�6(�g��uk#�����d̛ɱa��5��3�Y)��U}ϓHʏ���r5��Z��(�0�\%8��!�Ѫ�xl[������IM��5r��A9�w����2�Ģ��r��8�����$>V""_�F"�O.��\$D���zk��F���0� 1��yW[��k��q:4u im����0X�_-���k�F�[��P<E~Pl�{������O(8��O��s�C�	<Ǖ�.�s�v�0mn�4�7���������i��S��K1�y���u ��~S�-�E�M�l:�E��,� h
�����4b0��E�	e��HW��QX�����b�>7w���Y��XSqaauWD05�_%�	]^.`^�XS.��_8�?-l��j�����V@$�����������8���hۅ��ܪ�#�Βsކ����c1~�~�F��Ŭ�E�K^Ň5G\3�u�[ ��
�:`�J��CnD�Þ�5	�ΛL�r$ 嶘�~Z�8�/ �]�,?�l�,4���2�A� ��^AFI���Į���j<qd' �]�:T�5�~��ۈV�f�W%�-������:fDV��w�5��mr��d�0C�8A�n!!���p	�Ԯs�S;_���F5�/q��IL5ӧ�h�B����B-G�Y�M��{9����˛�v	����ak��/��-W{��]L�������WF����xfN����:�,�D�Y�$�h8w��mv3�Q�6�A/���j|�i4J� �� ҏ5�����Eb��Rd1(�F�-mq���{6!�xHf�[l�(�����Z�6�f��}�.����u�E@���i�m��C�|Wtjv�o�0%9���Ϳ��9���N����~�K���35e����<���.�-ҡ��	���~4GIʟ�qD�p�es�@�	��t��Q�X���v@��O�ʞ�˕��oxqX��g7���� {'0�Q��0�d��1 ���r�D�5��W����I-f,�4�+�VR�/2�'xw�ە�01lo�Q�����5x�d!$x�u�a�3�c��e$m� �yP7��^%O�ܬ��O�f,=���cV��u:4i�|������x�R�]L��&B~��6��/V̈���`<ن��&4g������(e рNQ��IJDupF������'�v,n�n�O��֨�.���L�2;7 j�Q:��(V1SK�;����:#:��-0���4�vUeQ�Nv\*�n}␮�%�	�u��;˻ ���}��{�.��P͓����
N��M��;��%��QͭDn7�UVf�������3�8�<�V,EU���e����wH7�CI����x.����H�2x_@D�\������.�����D�h�0�c�w��^�2�	�y������~4�Y��� ����`���{������'=	�w#5�7*�@��MUQ9i�� Ǎ�X[+��o[��w���=�w~+����F�5YL�eiK�[ZR\V��rJ�4������?����3Tԏ��1k
�=x��]�Zy�O�b����Q~�G���K�k�&�lm
��-ׅ����>�ef�9�斾 ��	����"󴇧��݉s�)�ȗ{�����}Y�l���N�����������m�Ja����c��{T��`��6IŬ��\��� C�|�d����煮�a�K@Ӭ�{��F������޽fe�p��k(�m��Sm�V��9E�7 W��g �k�A~z��c���W[��]��bn��9t��ʢB	��J=�*jzj]௦�x�6JE��8��Si��^{�w
6~�'��נ�ǈ��sԬ@F�Ϋ�f�
}�U�`��4b7��CX��贋82�N�q�Yst'����t��sʁ��s8�/�a��asQi~��3����Ä��e���S�0����W�p
/��S{d"k��s(F%�����}4�Z�T������@���6�s��;���������
I��W�	K�[<6����q��(��lk?���av�!#`+���sw:ê�u+R�@�+H%����o�+�GΛ��š{����i٦��5�*숚e�%.�![��pcn��&TS|~ۼe�1�٥kU�p>�.X��q��'wH]��� @����|�ȉ��lm�������h���v^!1��![�����BF�2��8Dfzĕ��e�b���]��JY�ؖC֩a��J*��.��Z��B�{����f�~K-�����V�}Ҟ���$�G�=vZB,tsw�xgd$��#��^�(�3T�;���8����Ë���`�̶�N��`y.{���3{�2V=(��`͞2�H�c=g���fMB
�F���C2�~g���x��������b�gs��X�n�������h0`>P�I]y(T[W�{��Gd��Ԉ<���֕R�ΰ8�*�T;��=�d9�I�d��F\�<����߰o��ׁ���\ĳ�v��n��]Z��fz�]o\dp�����KOv�4���L-���Ia:mpO�H�5�K)�	�����@e˕��cQ�N@���������G㦑{�V��V�,:�ѓ���9�F���vs�{��M���y�<z@�t��K��+?��Q_�L\Xh��2<����N�5��@$!'��x��>v�0�[Pqxfl��E�
z� ��]@�/�U�mc�u�)����1�5��>�)��	��+�hiȘ��$�wI�7gmBRH�kM��\	�d�v��d��Qx���s���+�SPWI��O��5���Z�D�*ү��>�K����b��T�(g	��_3C������x�i8�Y�ꙇx����� �Pޮ�<��y�%1�|%�Em������j�j�jV�xZ[�څ������9gʇK#v<�Ϫ m�Rxd�ʽ�X�=�D�9�υ�?��yC�\�6�Doo6[h�ԕ	ȏ�H��t�#��cB�7���{��k@bO�b>�.�"�Thi�2�(�֥9�u�H�z%;�8�rGE�׭��1��ސ���tw��H�g�
��޼ŝ\����6��m+�Pa������GQ����=v�fS(�l�+����+�{"��Z%��'����O����x�}Bk	���D��WWTP�¡�偿��;&�Lb�Q�M|wS�b^�O���ƠB��55�G���rjO��<\���$}�º{� ���<�P!�]��VJ�LI��vd��R�/�����Q���'0w�) �oW��mJ�Va�Q.�.w���C�v���/�1�[��R,�(d�'�`�w�
8ǲ�ׅnsF�UI�Ú�B�xޔ�8��C�x��o��p%�R,5����x�P8��LF�}?�]'>Z:<��-/[k��� �u�6q�tB��7� F�P��tf3��z�$����
�� 6h.=����>�5�a(B9�ĭ�XNX�A{4�-��Fv|�K����Dbd���φ��u�g���a�w�&gM~�m�kz��t��g*'5�yH�?����gR�������ZF�V�&4RA�.���n���z��(�]\u]�]��*-��lV�*�$8ا�n�_1!Dw��3��ʞ�2ƥ�&4��F?�w�{&��v.��e�v1�!��S�� �P4��X����"����I��J�MC���K��ķ�����ֈ)�R�^���>�}v�������	�Ȼyj�F��A3������RJұ�����CH�K�� ��ηnm
�6�x���Zf�[$��F�q�m��a��~n�:K? ��n{)�5Ix0����8�/r���u�5��ӊ�t��m1���ޙ�؝�U�|�		��6�g�fQM�Ͻ6���*�0P�
1Kݽ{�6Μ� qN2+�˩:�9�/��O^�
B<_l���W�%���L<E�"�$�F
= (��q*y���tS�4.h�h�V䶻f��6����gE{�U�J����i	��73��@�7헶~�K�A0+�x]�o�V��
/� C�a_�������v�v�;�X�6ٙ\�<_����Z��.�?�]/\�{u,ϫ{��DIPe�
��g����Pa&�<�?�Vx#��	�&�"�7�?b�C}�ғm�Z+���O�*)Ϸ�N�䠡R�Y���1?$.��ʊYF	+n�D,�T�\��������Y��03��0�'��A�+r�$�2�<��G����
�P�~-��F�􉠲囲��es�`�r��r@������܈��y]_�Dh�*Bi�tu�����O�){l��� ��>#J��f�%tN4݉���z&w��3r�=�ѰjV�N���DM�8�!_a��y��� ���n}�:���W8S��=�xO�,�>�%I�,�Z�f��+�"�0����]� ���a�d�JA��j7���R@&��(�1L���d��*-²x������Q�C��X��;���_��oJ>��&��P�o��t(��e�.�������_�N��e=2���β0a�W����lG��&Z�1���7��д�D�p��Fr��@b��*�3:�f�	}���E��g6���,;7;�������.��~��+�Upsz��{.�����ç�jp-���v-�ۚq�W�FU|�-X��Br类I`-C$�wO'�oYj������[������L�R��㉰(&��"˾�[{�V�U��U	��D����j�|�փ��U���h���/�I�ľ���g�e�)�)�ʓ�==L)�%��i�:Á�u� <�#C��-;���=�U�Ѷn�UF��I��wÁT����~�@�c˵ޚ���(�5����?_k��*z���e��ء@�Cx���lF"m�L��G�_z�;�|��8aE]����`�.�6K�Y҉l��h�H0onk����,��NS�4�Q�^v��\R�f�h<���������ӧ�ͮz� ߰#�Y>
2����޼@����M.���j�?/���
|7x��j�p~~�T�ͧ�֍|:�m�	a�@�v�Ջt�ͦh߂`�Ș�7����:�#�U�Ց���i�f{ć��W�|�(Cǜ{U�b��c�^�Pߡk�+���g�)+�J��2W�Ƀ�3��C�U�~mo��Ƈ��a#d�n��w(d���;��%:�^hĐ�eq�i��Ur���������s�A���:a�ꈄ��!V!�Q쇉 &�-\c�y��c�F�2e����8R�w�u��;95�{*��o*���GYd�xT�\%b�ݡ���p�AS���ـ��J%�#t1�\ę�g���?"���,2��g0�i�ꞑ����B$fgL~A9��2G�8��|���<�w������ws)�<�Or,\y��سoԞ��q�_�����k>���
ήīg*�,�����X�3��7�x�}X���`�[Ӈ�jA��I>�)��� ���ܹ�iK����N�����0�eKcA�����/A����*"�P6�y�ü�]�}���(�������Zj�2m^��j����:��U�p�Ee��6��Э���qHo�k��LЕ�Fd��
r����֬/to�AUƻ+�����UT�����]c���+����&>����I13��+ų�<��=]t\Ε��y?RM`덉��������~�晦����=��PX>z�������\��O\_����|���T�.FM�*��B�O!�e�&uA���+q;{�0c�� �=�{�#��I�fְD��r�>c�k�ghX⩣��:Cۇ��'#,��Ć(�+r�j����u�:�N��f��q�y�^�Z,�G�$�� &�h�!A�'p������o�'�o'��~j쫈�ȗ�<U�����fQ>)�׮=[圲+q�A�l�}�r�́�e;a9(�r&؀2=�J��
����n��&%ⱎ��>���>Dl��@}�!��n�&����{��[�v�7t";smo�c�|#�1F�����u�*p��eMO��ۉK���t��MAY\<��(��S��8f4q����v�(J�CB�[??c2�< �wT>Ǝ�$!#������: ��q-1r ���0���䅐�4���7�n�n���jg��y��JO2�ۋ�{Y%<[��W�}�R�o/yOFd
�s����M��uo�,l�n���S�`9���a�0-~V{O2Ǣ��V�H�N���%�SSm=���N���E&�`�N��TΌ���U�ncb�@�+����ëy�œU?@k0����ʴl�6����97���ys�U�/�#WX�\C��_4��q�����x`A#�z?��������t�!�uy� �^���j��SԻ����mi&X���RA[��-����{�-�xU�!u%��ȼ�d��8�2k�P�UM��%xƊ�Hص̩'.�������|21(�L
����TG�
	��J�R]�=ǥ!��=,��]sM�蚃��< V�׋���*Q0R�z�{)$�������*��
�`���q+�����al�"~�tPi������P{@R4�,�R��������
��V$�U��Vqo����I~�V�u��@Y�����ܜ����9��ͱ�c؟�X�*����T�b�C:���6��#C@��U����<M��]��i�}y��;BU��.�!�S��4�RƟ��i�{q̟r]F���)8iu��<��"�Fއ�7�h���+!��lÀ�m�6Ʉ������7�;f��ї�yh�ǽ�����=.U�Z��p}sx��0忧4^�WC���'�s�7� �N��ZӚ�]�ʼ�Y� ^�7�M�
t�+�Cf���7P�Fzb>wJ���Hy�<thI[��'����|�d"+����8���,h�1ܞ�A�I��UQ���ي�z�W0z���i~c(D	P������{�\Ġ�g0�b���C&5���(�� ��$�~ȅ�]�NF�{ۑ���k��d��ϔ�5��l"RgQ����>�`of�̈́��'�16sX �#e�fr���LUZ�1�֗3z�ÏYG��L(���H��Q�ڀ���}�\�0�.���i��G:�*`���?�0�ZQ{�"���Ř0�l���R^�!JF��l���i�kM:I+!Y���w��Aֺ7Hd���S�1=^1��C�mr�J$u����E����v�75���1ؤ���@E�%�+�e�"��h�5o�hYg�奾7�?��m�G�0�مeJ�F��aF���e�e��<���2R �k_�[<�V8_:��{�֖6��!I�Q�=Y�dx�x}� �cѯ�nn���D`��$b�u���}	(�6<�Vwȿa�`�@��%n�S����]G����b�����=!>f�9*������v��j{��7���c�$_&Y��9#�5����.J���|7�g���Ud���/qB�A��l�Yv�Hɑ��H^Ŀ���#99���a�t�M��L.4�ð7��2����-	��<�+U��ר?ؕV�CM��E�8�va�Eo�r|���G�q����LT�:ܐ����r4(c��<�w͆bh�%�ma?/Wl��컜 �kI:�i>>��k
�٧4-��k���J앶O�>��bG�{�B(�̮_vBć��[�������ӎI��bVyG���9~x�;"�PƶpKl�短�D��i�&[�|К��X�x���P��X��m`�o�����8�����5Zkf���K��հş��L�,at�=�T�\g�HP����gХ�Y� ��-f���n�@�k���'d8Y�6�1\a]BOc�k���4E�*�ZҾD2R:X0�7O�����Ş.��su/LU�5rS�P'}B�"��B�P�ע\Z~�ep%����IWks1J~�
�,yxK(��F���<��ӳ܍@-d������hA�S���K(��e�2�}��!�����ۑ��%��������� C�����ǡi��\�5)����
�'����'g0���1nZЍ��k���������U��3]�`K%�߄_gs��Ƅ퇞P[z,�H��@�^�Oɣ}��ۙٶZ�`���0�t�%m;W�&/F-�
���b��'�	�\|����l���`�o���cY"=����~?��,*�d����T-�w�D�������%�̰�����p^-����I\=�t��Z��6cF�9�,=F>�t�/��O�m�y��p
�����%�]Д�˲`�i�'Y�=�'�hӏ�E��v�;��i�t�i���*C,&�'(�w;s�P�����qp������ǻ�u�l^X����۸��T�;��"���q�&T�U㋇l��
ncC��\����tFUsl��Q\ˣx���(,��p_ٔiU&�r�<$�D��\���~a���;�&���%�Fe��'�K<^�\�_��H�08ة��R�UiiiΪAr�p�C/I�1=�r�^��=<���oÚ�I��-r�K�qܣ{�:T�h��z�CMq�B� S��^E���x���T=��]m2�0$$����y�*��Y��e���E�z��3~��c4}o�y�H6A�.`GNW�$LG������Š� �< F%�����(V���<s���n{Ώrn;M�jq���sDy�?�uZπ���h��@�y��Zf PE���r�Sզm����{x��=V+r�O}��F�4�(vX��p�YN�{N����1$��v�ı�N�`7!���ѱ�������)��nՆOp�(�P��H��i����'>�4g����ҫ+�KG|�j-9Ud�H�ƴ����;�n8ةOC�x�r�	RZ� `�.V8б�W4|V�z�8r��﶑�F�8ʜp���N��ּuk�R�>U�Q�KtaŢ��*9�m�?a�0n��p�����[�Kٹ4XS?�N{��mZ?������v�h�GZ�����*9��&��Y)�'�+>��GO+��XA�x|��w��Ux�`s�c!Ʈ!j���"Ƃ���b����d��
��a���x��`��[��(hN��HqĤ"ks+�ay^����{�K��;���I��mH	����{�X�<Lδg"6����"'px�1)���/r�uw�Bo�"79��-ߠ�IL�y�%��&�0w�FNs6Y_C�ltB	H���}I��^/���jc-vBX�A{�k��`"�!J�'��@m6����e�߀0���^�~���L�ZCQ�����4]n�O�S�B��J��v>��֊���Vl���&���!w��%�����)��;{���}�[��{�nn��q�T���8���r_�p]XF����n�ڹ��°���D����FU��D�<Ԉɡb�s>Cʾ�ϵ} ͈��Д�����ݔ\�+�D�����xm�g(`qw`�q]y�o�������%S�s�+��𵑈����y�g�%D�e8�=� �ˉ���d����-om�_�UB ���	(��}��<��7��90rV�-��~��7���ǚQ�;��-ε
�q�W�2E*߸\���3�F�wt�.V��c���\�KL�����3�^���*x;�6H]���0����LB�@n6f������'H���Z���oTm�?�n%����f?��^)4���B'*C���� �r���IWC��1���=[���%� ��05����ǂ�Pc��!S�7:�Sb:�B1��v�s��]��ߗ`@���N���g�����Hs�<�r��4���/��0A���jW�A�=0H�LFR���k��"h� �q�mQ��65�&z��!g/�n��+#�J%��x�����@��#�/�8��k�.k�t
�0�M�"�}dQ�?���i�bI�)! �.l���t𙆸$�e.�6�X]�gV ���I����Z)��3��i�� L�	���Ǉ�]�ç ���N\&'5�+��ܴ_B��do��R����>u��W=�w�������[O�/���X]���핽D�����wɋ���#�MQ}*D/�d@E�>2�_*�
��>u�5�)��J4<�ƌA������b��A�6�.�m: 5��XEW1E^������_�e��k�"���� �d�.Tʪ�xQ���<ʌ�7c��l��Q�K������bl��.�vjL&�Q�W�Kd���$�47�2a{`y�G��+|�B�IMO��tBr�z��E���K�e��`N6��� ؒ��GM����?�[� ŭ<9F/�i�-@�)��Qk� ����q;d�Q�,�ʩ���ю*wi�2T��@� ���@��{���eQPG�q��[�OA?6b2�d7��"r��g _�a�O��%�#��wT�仦�ya0~/m��|J�Z�G��Ñ����RQs�Wz��-eD����/���s�U���N��3��f��Y����loz����A8��y��>�w����yЍ� ���U�c֧~����&{=rF'Y���Ԟ�
K�Ȩ��U�����1�1`���[FeR��M�z�0��
`(J���z����*���܅�Cf���`[#�Ԅ��A�*Rfk����r�t�,��n����;�e�d/������v��Ѷ-��[aA��wR?�V·#u�o�(�L��N�*����A��9�#�8�5�y��5镢�(ޢ�>�X���2xX,�B�����,5��Z�f0c3T��;@��\�|$��GI�V���P�D��=���OY���Gm����Na-���c�g����.=h��"_�h�,M�\��T�1���VW������~kL��;�4���/ep�qY���	����=�U=����.� `e��{�R<d��0��� }s^'0$$7�~MŲ}��k��[BH#V�=�"�xs8]�x8m�`���Co�l7�+�L��*�A������aE��>=�����ő�k+�)�̺�h�ؕ�1�t�ϲ���,�aOX}��6^�-�F��S�*�~[�t9��^pG��7��t$��d~����8�Qp��bP�E��I��������!�g�yT�LV����T����vp�A��V�kPk����7������}ȢC��%Z6�N[t��z�����z����)@��&�<�z|�|�Fr,(6"q���#om^_�者Ȅ4������?a�v��4]��*�p�˕�$�í�pd����v�<�Kh<n/T
��6��2AUc
�r}��\�P[��	�j�DQ6y������4�:!2#9���=�Q�54n�qQ�<'v>�fɯgB�B���	���I�^}�[,3R0J�U��]��~�5c�
"�6�V���q�)+�\����
�a�����83B}�����x�����P�L�Z��j __�^�kH�0���|6�y��6������k��lJ��٘��X��$]�h��nb2F8���'ܟM����e��;b�[[��ON�&���E���� C��D{�i�CZ�!#���c4
I�Ҟ��ϋ!R�I�^Y⡏X�',�pvMb꓌�bB)��fR�v�M�ũçf�ʞk�o��_��Bt���m�By�vB����6�Ϛ�/��t&'�j6c��*Ġ@�#ч�pEr�óg=r�`�p��|O��%���dk?,�A@alk�%�������o�̂־���llH�J�8�2و�|0�����sr�9:�@�uBA�wG�H-|�J�$�7n�:EEn�"y��x~����P����6���q�HAk��E� !%�;`���h]u0��$�໓� &�m��
�eg�R3�������Q����9�|R��/$X�Q�w3F_O�I�MK��͒/�v���iMgz��}� ����L���zc:- $S9��@�����Y�Ɵ�㝾Sa%��W�͔'�:g�GN�rc���N��H�p�����30��D.I�藳�C��0�m������3�\��e����v����a�0^bD�Je1䫍����Vi:�����ƚ��WV�bbJyR� ��-[�-r�S�]F1��k�9���4^�F���o������,ִc��^�����_eH�Y~G;>l��-��4h/��яU]��H�z3NU&(�|4�^X�h Y7~R��t�Ga{Ry��^*�;��?^U�[�)���Q��+����0OPBX=X� ��_�Z���ĩ�,�-�2�.���ǯ�����HIw�/�cJ=�,9����n�&��[~���4W=f�e�l�s�`:�'�&�I�AΘ����F
y�
�ˬ�w7k�8���63��2��?U�KQy��+�tί�ʢ�rr$p5�X+�¦�Aۅ��M,P+��a&�������� �*k� I[x-�S�F�\�}��y������z����<�\�����< δn��6>�#���k8�$VG�|}�g�(���%�G�~�6zfy��R�M�	[�D�Pk�^�⽏�o!�!k�{�433.)����ˈ�9Q���Ye]������sp��iѐ"��B�U�s���"d[��.s�s�tӠ����TP<�t������]�pw��|�������Z�T"ִ0BA�RK�pٶ�Ī6%�1�c���5B�D���&
K��"��� ��7y�c��K)���X(��3.%v찿��8�׫9G>��0$�)�r�aw�󰷙��:�1T�
c8��]���K�0;���k��.��u�n�<�A��2�q�N��]R �[���j׺�uѵ��C]���r�N��oep���م>I�[I�[w=��g_��Ec�9�w���f⃆��MwM>�ʖ>��x�,9���'ls�ڏ�z��xE<�/9����\!�ئ�֋�Z�^��fD=.]HI���vvZR)��J9@R�G=ٗ��=��"��-bB�����,��ј�?��ᯯ��C�U��_W�?�N���G�zT�7���6�:�T�zi 2|jD¢�<?Zh�@��ɪ�Lw&�h�n���{�����<�π��>�oI���_("o�{���r�C���Mr��Pz�@����o]�y�f��!���mr�y}7g�ZaQo[$ 僑�\���o}W��q>�7�v@�r�X��f�$���ж�&d�Ť��Q?��cφ⑿A�z�������W��@-onb7��Q,Rj������5|S��YV� ���~r�v�y�!��Oe�vn��2��5�T=�N�I��M"W�f�[�����q�v�G��Z��R�P���bY@����KcH@�^������ /�"���c�C}���H\���ҨQˎ12�y�T���^�A���q�?z�؎B�'�˴>n�R��k Rf�u}��m*=�F��#*h�dG��.6D(�a|Ҋ3���ü�P���X9�2���`��8e,�6�����`G--�U�2���S�(Ġ�*sh��{���ASH��9J(E�!2���&d����e��Xx}n�k-����n]�����e�#�z�c�r�#3� �^jd�{���{l՟���6w���&�䑺��� �'_1@����b�e��o�޷%FA!��������P�MՐo��~*�O-Tg���ьHt��$�n"�H��5�#�s�����H)��v<v��	���{��\ZhJ�[�y0�*kc&y�A�&�]a��:����]�	P�ex�xe�3�N���Q����J��$�5E���ځ����\ĵ\������B��n}��y_�o������ȞO��ǫ�̭R��_9���Uj����u᫝}�9Z^�8�昺+�k,�n/� �[x�E�m<�匰��j)Ҁ��N1�3�5�+]��
yI@��L�F�%^XM��~�^J��3z;��m����k�	��#�Ե��xmN�ɛ�*�s�d�@�A˹��~P���K�a$��% ���cs�񅏲�@���.�����k�O:o@H���\Z:�L��N���\�ϘA>��4"�}���$&��Ds�����;<�{@J�z
Q�$Ȓ;�����>q�<���t�G"(��������`d��.4_�/*�4>(��7"g��ȸ�2���RR�U	���&�@.�.1Y;��.A�?`.͂ьOO�{#�ʝ���L����(+��Z��G�\z����;��0{��!��ø��|�K���s��s��.N$Ы��G�C2SK������}�83!Q����8�-����4	Q�U:"���B�Q�����ά��c�'����'�vB��������i�B���^�/Ҕ�f��Ų�2m�V��}7�i�+�8�˦!�+J�<h�a���}��vN���Pj��=rM�1�k	���?F��J�{ZJ��}iܟ�u����:����/��Q�ȗ�oǺw�աaX�HE5���y(_hH�Ύ��bE�nE���8yP�w��h�JM����"ڒ�
�H��	����A�?�U�Xh��JdnICS��I�rÉp�z��y����fF��wg�C�S|d�oC:��l�yS���T5������^�� W^�eƫ봎����$�f��E,����c�oG�%5>\sƜ�����Āx���bOw_���A�V���='&K��!)eXN�
��<|V6sT��iVtaW\��ŧޓޫ�3���GXk"
�f�D���1�������K�J`T%T�M���~�6�Z�뱚>E����2{q4�D��B��x+֋�T�o��-��)��ƿ�|.}����3N��麿��!�Ś��G��fȰ�ǘ�]���U_�q��2�
7	q�[�9���D����H�6��cbZ|Kя��4�B�Y��@wXe��%�P���-�<o�3/�`$�����zNkЦ��~��6g�-j���Iη;u�u�#Al{,v4���@�P؉j���k#��?3xH@��Y�`$��7���E��� M3<r�>.�xggv���K4}��q�m�Oӗ�ݷ��
@O{����@7�/N����-~ȮU�y1��PVD-����4�̉Tp�I�5��T6D��q"�x��,�#Za!�S�����'�u�m����cڢy��ˮo��cx%l��3�z��a�i$���uNڏv̄j�\4�\�qg��vӈ�e�c3,!D��6�!������D�Z|��M+q�N��;���h'��v�S��B{A��	b��3�FmU�ҮL�ꆢ|y�W�W<4@ؘ�BQP6����n�ӑ�:�0�	�䑤�g���E��P��\��@@��;�Z2'kA�m�Iu�����C�� �	K��h��R�"����A�ȯ�n &��ӄ#u#���t��/c�ԣP�O��Z�	�у� C�ڲs�6Ձ^=�x����E'�\蘯$+i�e.�>Ё`����8�����l8à�Ҟ�u�!�'�o�)��{�����ك���8��D-�y栦�t�����۞̫��k�*v}�, ��]�N�S�J~��q]�F��vqUd�J���e�
��ud�jJ�k�Irv�e@!4m1ߺ��}��A�)�BBP����o�XY���*ɏ�l)��l�b�zj��^:�P��ٱ�<kƱNw*��o�R���Wt��$P>r0����2�u%�S��lE�k�'C�� �yap��a	��矀�k�?[y.���Y����]��['V���R�e"�C���c� c��%$���9���������őL	H��k�ê�a���޼����s�M�QsQZJ
�>����,�Y�C�{G��hg�\�W�/�1��[�#P�`��êP.�T�����.�N �̙y�	��ށ:�$}�,K�f�Tv���P72�F3�A�~��Ї�7��{�g�q?�g�_i�Rev��')���ª�w�x}��"�r���u��SQ��6����`����3x��FU�!��Iz���R��>E�YA)���J^|�D��p���Y~�7h$>N�6H|� �*/��eٲ�9V��d����X~ǵ˛�5554�����*>��C�K����V��yޯ���ڪC��YD�&<!*YyG�h|ԶY�?�щjݼ��R�xLJC�z�^�>�Jb�����ު=_uY�H m�~�.F���6�WK�H�Y��uwS#�c�{Ƶ^5_1_�0�`�dRߴV1��J�_�}�S�-λ;��,�T�i�ѿm����T���d�V��#�v��Ma<�	��?ax�3��[����>[�`��u��W���?�������#�
�����~��i���Q�je���I�(;p�d5H��ي����i�>8�I%w�K�z���M�������x��Q�U� �Q�u�+}4��p���I�՘�O�gf�~��k��e��v%i�������r�xƕ`G�Ȧ_����LH��"0P<�5�2�a��iR�����t�z3��Tx��ӡwؽ�Q���?�S7�%�<���k���n5F���Y�̚�:��U-��a)�����A��;rK3����M.����wNսP����i� Hۀ�w�A�E�����)"m�)v�>�p���Kg�k�#��.~t�2v��<fI)���A�V�v�)٨���*1l���
!t��[��E�vL-���B|�.���L.�
�/ro80.�k`�Nr$�JK�� �I��e��{���A/YV�u������s(�����ux
S�\M�6?u��f5��8i��&���NPLh�[�����k}.�/�w/8.8sZٻ�ZQ��|�s�vjǾ���2�+�q���5\��c����)B�z�1b�.����W�C�F�]t�[U���f��oA��R�{�ح�&�W�иӽe����=�(�.�͏���	�Xc"�‒������7W9��U��O�*�4��(����O���c�w}y@�J���	��U%�� �0��n �nm��9��I�9��yw"�V��4��2�i���V�e���������n�d�J�&F�pͩ�����DS��ezB|@��PK�9h�5\O5�{/Ӣ"��+�^8�>�dT�#�@ ۑ�����և�sT��4���0R3 {����ļ�[�kRQ?<y�-<k����0|�6W�"�Qy�?FCS��{j�5ð6wi��>S���܀`{�H�\U�y-��D����	Wt�NPp���(����
!'{�>�v��;��T
P���T�Kb/5/���$�O!<�V'  ��d�����˱zhq8�8�
Zqw��j]���N@��Е���8����ʈ���kK�_w�h��CjN�
���c�I:m�A^4����kMz�֙L���e{١>IR)A����.�l:ܓ�&�t�)4l�Q4��e����*a���%#LoVey�p �v-����K��Wpy4�ܦzs�i�X7��� ���V�\�j�T�OG���4Q�+xC���"]m��l���� 44��O\\�`I�Fq���G��g����3������h�+s@�O@t{A�+Y���~t��R9��A��)J�A4���EC��^u={��M����,)�
�Յ��8/#4f@��=��x	��#��!���݃�X�ٵ�)'p;�m�U���A��bZ���[����T�Yy�RL5���S )*\���x3�<yw$�k�>��Kt#jC�>�j�r�H��� ��VJR�WD`�B����im��u�:���r��{��xTV�8ԩl�(0���&�Vv��_��:3�x�$� '�㹙"d��#s���u�в�ܡx��8�3;�zk>�s���/fӅ�rW:���p�`�e)�a��/D��<�����ξ�x8�!�A�|��]��q5�b��r@U��ܤ��m\�i|������J���:ձL���bӗ�嫀�v1���k�dL���yQ|6S0��+o�4�{7�)���9bO)Ka�L���o�t�TkKN�!9��U�^CY��xP@�9f+�v�$�]{a��f\�I�[\<>@���R�}�H�I���#5G�B��.���3�<�Q�kA�"&2�Z��bvw�P:�I�=��@�j�6�����Қ~���cv�8��J�)Y�C�����A�ۏ�/q"��Y8q�.� G.K����q����x��
EH`�m���r�t�I=)j���j�P���{x;��XהȌrN�]�G��z q~�+��7S葇�$;\!*�N��.EB|�~�d>����Ҫ���O�Oa~�^�W'�S�B�̩�*��HH�}0#�YL�zt?"�(wA�L8j*�$���g�ߘgE'2��T��E�VewJ\�6E��AF�u4P����w^��x&���؈T+�łZt��C�%l���mR�m��'$�����%i(�j�a�C$�z<,��� uc��5y��eӂ!�w��� E��2�֜��M=Q�����'y�]w���kFSs�Iټd�A�_9���|f��3�i����Vlu�q�0qT�g��|�4�H:MtQ�E��ѡ�_����Z�T��<�8�7�}1�\�7m����0�F�cW��}�7� ����hC)64
��s	��J�A���kf*���(s}s�cӷ��H$�e��_oʦABɽ��e�r�p₤�X.}����#��l�3�W,ʺZ�HO�o��G���O=|@Nd�y��b>���}L)�I�f��j��7!~8
���k8[�Ɯ���,D��e*��B�m��{E��LXV�_�o�i��|	�#��8򗵎�Y�͛�L���㪮);_%
���e�9H��:E,#W�Ⓧ�� m�pM���w�*�l�W�;�>�"]����D.�J����G|~B��B�3��Nf�,؞���ȷ�"����鈑M�r_���������!u��q�LU�(��'Ƃ�cO�<P�,ґ��R��͍vkޞ�� ����(�]��m�ԥƻ�ypu���=I;�Py�ׅ���ʻ9*
v��c�����0��G������p���t��3Z�S��|Y
���&��V�1����5�'�_u�;W�����2�B���\# A�].�s�ߠ�s!�ӏ�#a�T�6ݤ���"r-��3b�8��w���x`I
���3R��66o�x��K��Ҍ�ה/�N�x���g� HJ1�@G��jp!'L�H?z�9� �������W.�3ةnf��냗K �d�t	�IS3so�<\�P%��n7(h��ۇӤ3bG�Zx�nC���R9��ϲtjhԚ"�[]eyDb�J�x�gx��N�o'J:�ö�qVg�����?��6��#}��NsN���"��r4�P�I	��JC�ex��X�w���3�����n�� ����X�||zK�Q,�(~|������(nڋy׬�~���!2�:p�5�1xA���L��`�Fo�1�#̳��+/ �v��C��ig0�UUF��$Q�����^�{���ݙ/�M4&��O�	�e&;d�Z�B4���z{L�T-�Α��Y0riV����3l>ퟍ&�2(��Xs�[��n��>��ua��h~�+�<��z��g��_���+�B�š��Ҥ��S�Y@����m�Z���A�$�z��1us�I����+���u���})�(�A��	f���)�Cl2�����$᝛J�dAx�5������hT?95��G�������j�.Am�Oc� 6`��s:��@��� qKǴ8�J��[�]�1����Pa�t�,K���s�ַ��DP\�k�yb�ng��7���;�/[Tb�����a�#C���5�'��,��V��VQة6W��x쨟�AV�0�v��Q*e��|%�����U�G]4�._��em�E�ň
<�F"��OA�)�d��5AcX�U�L?!��V'�Z��.�̟�ǜ�{E��"Ug�=�-v�D���d�б�ӥ�@�j]
>�郦M{=��#'��}iȴ ����8 Yw�B�jl�Wj�����E��v,Y�����/w!^.Wt��?�0ۂ���"?���0�5�a����w����7�B�5�������%՘록T&<a�P��CX��~�y��CX�Ы�7|������6](G�ٔQ�]d�!�-m���
��]�R��j#R��c2����fhNԪ^���% D�� �N�Ϯ�*�ù�$A����(���<r�ZJ���t��s�H�N�ɳSN��t��72��i�ھ��q��{�� �Jw�-X׺c����\@"����TG��fU s�I>�����Y]-F���EO�[�H	�Tt^J����b��q���ݚ
$���)%���A��� A�?O�T +\P l65�P}�P�iR/hN��s��9E�m�d�V�^+&�zZ`�;j@3�=�D�j��!f�^�^�G��'p�	�����y�'��La�'.Q�U$x�~lOE����T��Z�#��k;�֩�v�]��a�cN���cu�ܥ��^�4{���C����h�"���c�&F:_� �*^���S�w+{����f�H�~��ױ3��4E�!pl�
���7nld��p/�\���U9|w��`7�ok�@�ʾI]���U3R���9������M�f���Q�gӼ���\f������<��B�C��y3$���٢.�Hα��􍶟�JY�1�3C"�_.�U�ꃌ%�	�N��f3Ɲ���E�ϸ7�7GN��0��Q�,�TP�$���j�ԯ
"��L%�U5�۬��a�������2�*�tMFݒ���Zh�H{U�q�]�����I5�� ����}�]p�cRo�3��v�rRŐ3t�oF�գ��,�t��B�]3�F"s���ʣ1�Q[�5E�#u���&���$����4I��D}DY���a��r�W�����1��g?	_����n2��D6,xG;��ܕ�&E�J%Wj�ne��W�3����,��bI˽�M�:6�}o���7w=����O���_��Wi�!���g�u�aZjNVp���?�^O	��3,�W���Y���5�<�$Z�u�Cpy*>��<v޼B��M�.�kƉ%�}{h�H���ˀe�PϘ�A���cpK�vn^�����m�Wn뷉*�M�Ã+R��FXݳ'C7�7��,j�'!0��@�/>��BL3���ۆ	�x">|��F��~ѥ� ĥ#d�#��@Y7��5��pp��fP�g���^�8R�xQFc�"]J���ϪO�>�����=�����+S*M=*B�Nz��sT��k#�(����C�<���E+>�5�g;���O�g�%{437�,�$�?�*�Zu��{��ը�=����QdϹ#!�3o�dR0���YH|��Q[�J��Gf�T�񺩨���׭>*<�M�g�wA5����-A��$��̤��E|5Sx�P	qP���n�}�(�D��*��EhC@� �#	&b?��p���*��&��:"�*D���NJ�Yv~bF2+��Ď2�N�B��&)��x�:G��`�
4�5��"���N�ܔ���Ű�v��i������*��~����b��Ѩ(��(�19TO�OHS
.�瑢k��-^)��@���!Fí��eTO��@����<��?'�=F��2��~�!���W�.�ٓ��$��C)6�lcݼ*�ѭ��	�:������	�d�D������*���/o�M��zņ<��U	kT�W��QOG^Xob͎6R^� �~���3����Ō�\HcE���{�v{hp�.ɟRjB{C,½����<���34�� �Zq�|����̠iU@��\�]�NA��Z���=�]>F ̪��g����-�V�֯;��)wJ�(�E�N���3��&u�t���w|57��;�8�7����V���5Ƚho��5i*@Z.�Xi��=�}DD㮩`8u'M�Ăn�k�� 6�m��-��[/���]9>¢C��n��mM��v��KZC9�ЌM`�Ӛ��b���✽�`�}8
u!���.��8���OUdg���KkX�j����$�̛����ӃL��R2nv���.AF���;��v������M���d���?M���=)��T'�l@`�3I�6퉯]��f��uJ�9�F��M'��9>�^>hs`�AҼ�\���e������^��
�sXv��c�����E�>�A��H{��*�x�������K;:�~d[<κ�K�:��dQӉ���T+������y$֔Ny�4�u��!lw��P�lt���x��4ӝL���Q~ U�:
��HM���3n����ϩ|)Պc��"S�O+Sz"�sbó/�g��aD�<��W��a������]cV}yq!L�c:��FG�o�Y���W�*}��ɣZZ>#4%��5�����Y����t�w�c��z���G?U�&��Ǽ�8���x,%��b���q�R19����~<��Gk6)�{��{Hw��|�r.�I�=����Ü��LGu�=�v(�<�k�/'���kz����'�d�R�l�ZᆪKv����m����צ��mE1�zфr��$�ň��D��х��U�Q6��\(0?h��>Z��}PD�Vcov�'v_q�W}b"�X��H��C�U=ƶ���	2I�v�f{�&߇���*dNGf�Og���k�x'�C.��YN��t���P�6z��jo�Nd��HQ��%�b>�MS9�d�K���鋬&@�6s��q[�$�m^b����Aw��%��)u��u��!�H�p�s���d}���n��3�@�A)wbU���ǻH�H}kf�kܗI�v�r����p���
KbH�a������z�i)5�!5g�)]���m�҈N�o!<=��3�a�����w>>��,�i��B҇{�䉎�/� �E6�PD����uuV3S��N���E$f�H\McZ�=f�\��q��K�z�T��6��Yƨ4��_�`K�+Yc��3V�ǀ5���!]���懲�hYy^�ބ��א(T�^e�{a���ֿ�U(إ�az�?|�:��Z����j�Y����J4a挮�,i�)z�#�!!���r�޷��D4��G}"b�G�ߌ���}�{d��9�6G�B�4�s�c :H(�z5r��hdF!'� V�[��GN�w(��(����4]�K��<����B�ԛ3�An'a���.�±�&�}�3tS���p|[{O�,zv�1�3�\�.96�d��7)i'�6��6��şw��!��^-����\L�5���f]#��pѪ?����v����hk%_�%Ԇ�x��oD�����(W����s����+�ZV_Q���Ԑ96�	���>�W�,>�zU�,'y�D;�������+��3���\�F��=40� �և ǨS|�M��V��2����
 .&VƊm6�w��&Q!V ��w���L�ȋ���qST���{'Gdn�/�`�f/q�����)J!��	�t����P3�>���Oy�����e�j�:QK�� yO+ڛ�����@���JG\R�R�������!N�?G��P��ƽ�SNC^��ڕA#vd��;WY]
�B5�U7X�yE'���2ԃ�"�W�\20V1�!�~9X6&B����P����2���g�����
a�6r�E���֬e9�=�X�} r�0�6Gd�h��rT����ɮ�7Vɩ͜�26������C O+E���#خ��I^R��C�l�~U���O�$ؿ���o��i��T�����(mP�����n��%\|�f�����=V����F
\�膇�Ư)�V7��9�q/ӷ���_jJ���$s#^��ʏ���V���i���(�[4j�^X��@%���ڻ���td^�C˫�Ǎ$c6�ΚlX����_r\�#vg�;ZU�DH�t�e�u�@����oWdѱ�ʔ����ā�q��rm�m�	U��H�?0�cl��̅E������#1����GTi\�X���^�Y���M2-��
!Fj���Z&�<�3��!v��d��{ ~���oȔ?�m���5����`��f{�s�qr��B���/��K7���eQM����%fG�/=]���l{��G�����U�w��ɀ+�~�L����?c�2t!:\{�z��M%
�>:����@��f~���� ��C�oS,ű����TV]�7�������B��L´N�Bz���
�I��S	�
�f���+���т�2� y�(` �3z��o_�l�֚��Ai�3`0�(��x�B���L��8���W����@�������c�>|��;�:�^�=U�m�����|����	@莓7�EKW��+��Tk���K���g�2�b�Չ�~%�$�j ����������M��#l[#r&�h?�_,M��K� ��u�;8S#U����_��R�8�!K;p���S��cG./�xڟ�^�?�wX��d�#���X���Ifɛ�x����6���̉�y�q�}���$���r���q�-W���+lhT�:B#�)��`�13�w���7�S�PfI���_vd*��Q���C���x�T��'0E�FS�I�����w�M�ҿ����i��Ġ�H�,��h����R����u
�K�I�wl|�����"�j�WaVExa���gРq���^qN�"a���Ƙ�+x��˃�բ#�":���+r�r��]bc�E���f�h��O���TP��uL���	���X'���{K��k'4DѬ�bXV~D?�i� ��,�Nu�.m*O\������J�RA)V����g_1jR���qh4����6��k4�zN�U�D�6����w�Mܹ�O�[?�Lθԁ��������ї�M�-�0���p�ݶ��O�z����'le ��)�9��ӣ�r��Yt)j������S�f�e��,�G0�M@����Е��6�� �1`�Ȗ<�yZ���"�5�ؙ�Z���	_ۂ�[ʰQ4_����g2��rAd�F�б��K�a�u.���l�h�ifIB� �_��%t�oY�uhqߏc��mls�ȱ�k^sdM�� ��3k$��h��;-���耊|�^j�qp;<Y���l�� ^��w3�^�z�v������U���F[��r�i��
��gA�3���N�4�;��p��
�eDׂJ�e��?����(ɽ�:��n��L��UI̢fu�څ���Dc'��Ƕ5�T���� H��p&1
�$7�����`f�l��]���3�"̚�E��:$�� �������=Rs�� q���d�sG�Q�1?�����^�NG�( ]䧬�V��Tۉ����F:��w&��k�ѓ2��w,6�%�o|F��{g�M���Э��eҀq���Q��~�ʵw�;�V+5�i�%G���q����7�`��谔���-�|q�
B+�oT/�k��ql"�MQ�3;������`��Ι�$�\��<�a5��)>F�]��c�hR����K���j��?��f_���J��`v� ZZ3<�D���x���9��>j��d޲K�2���m�m�fCؽRp��p�"Ֆ$6�����6Bk�"��'<����0��}�L��*�\��b�P���N*>b��dpq��d�(Bϙ2}���z�`����xLYm6VԲR"��;!:���#���။c§��#bYDrf�F�`�Lg��(��Τ�}J��([8����qA��?80~�ؑm�-��G��6����4+�?Q��H%tL�3�0M�6�90�R��,�։�E�ֽK.��m!���j���A �$�j�a��u*9I�Dr�&�I�M�����c�q�َ��y�!F5�>��}��Px[��VrX� ���j�.��m8�e%�ؑPf�S�����yZ�Я<�٢��
)����6�V����/3��c���I�=Ҕ��m���6ją�!�Kd�DXjE�ֱ&�$:A˟�^Q7��:?��!�P/�?N�،��'���>{{���i�<)������GQ~��w�xqF/��9�r�-S2A�y�
�A)�=�cB
t��a�}�%����l��n)�9�<��\��絳�Q�}����(�\�M���s�w���br���o�RL�,-�7�-�S�YSd�e��9%��w^�[�{��	]��\�t��ҫ�:��Μa1e'9�t���iB�!�>�>)�-˝L<R��.b�1�Q��[r��D/�S����'�>\�N8�� �͡p��ø�ݝ�*������U'��v�2�IZ#��d!��"t�M��d�b��ZAK��fOb�l���c�{�����g���D]��i` R�P�{�l��{��������Տ���:B���A�H*#;Ø�3��������z%;�IZ�v���Ј+����d5���9��0�{4E��u�^T�-�ZsdPjg��]<���p�A{-��g}F�|,��"6��(�q�槑��x�g �NRAh�a� II�	��`��� XṠ_�����'~�ONwX�8T�wO*YƧC�k�#����0��E6�W�oZxY���e��N�"��ߐo硍�
h'���U�\��[S��:��	Zůğt[�X�J�Np�C�儰V0 >z�:³�}t�\ї���D"�#�D������<�=~H	�b���-O-By�.�N�8nf��id͘���9��^&�SH��[�	s�c;۪f�Ny���'7����4[ӎyPWҩh�c��a��T.Pp�\g=d[�����X�8F5<9���D����_X;dN��b�:��kÎ��%K�t*3u��~}�g/)���4]���z[a��1�4'_y.h0���?+��Q���.�+ʑf�O2Jԏ,��9ch��qS;�Rg�G����d��"W#�y�[����:��v����0s� 2WMPd.�6�I?������!��W�B��{�u��+��n:�MZ�~_�e72�[0^s��s Zk��'_�~�s���'#���?9*�T�z�M�T�C���GQX�[�̸�\^�4��]�9"V��$�\�'������ůL�50�Z�����ҡN�������
�"Ʒ��D� ��k�
��/u\4���R�)_m���o�~���q#H�W�`#�q��G�����AhWe�¬W��-M0�P[�(ڛvB�p���^� 上�Ǥ3���d�s%c�f��h�c�1�-_�B:.�s����ļ�����N��A���7\G��{��jQt��lb5�MU��2��x�Q59?�����U�ʯZ���'�/: 6Lv��E�:�y�dċ�j��F�}"��P�T�˺�
�S�mk/&��Fa��������(�?�h����~��t��kƨ����^�jx}���כ�t����P��W�7���̂��B�.�31���e	J����?s�ֈ�zH����Q���A6�{����8���!6a��z��'����^�(�c�{ِ��("�+kU�eG��X�Qv~���/m�Ϟ�-b|�mͥ�a8j5
w ��2���>��g�
���, xl�}�����J���!�-�H��8��
�$��:��ӹ��H��l�/15$��0����{f���XWi|h���α��FQ���`H�sW� 1�3���B1���fp@��n��Й�j}p�5�pIG��-/�f���F�v�6n5���U��Jڟ����M��KoC��&dO���%��Ł��K]�? M�B8̧<Xⶨ�'��Y�.���6�n������ѳ�u�E�a2*d#�w�����[n�$�@×�����n=EW�w7~��Ҙ�M�$�w�]5Ԝ
qJ?젰w�j��/�8E�rr�����
9]%�6S��V/T#��(J�M�BL�����%»��@�,7���`����j�r�mi���P�/?�\-\)�|��S�OQ�X@]fS7_�0�?+���R���=S�ܿ��������ET�|�7A0'4�oW�ܜ���FUo�UTd��'�u_@jtS�� pw�����v.��?�MR�wJ��M)�D]%D��THdc��{�Mw։�t1}�_E����`�����8�.��v���4W�@U�i�:j��~�U��U&�Y*��^E-�����7���h����ؚ��H�����ٝY���>ǫ����w>bx���u����z�/��ދ%����ϗ�ydQua��Y�������*����ٸ�os���1]����l�/����1kѩs��۰B�`�F֓+�d���ߪ�A'èJ{a���[�C�����$��:D3Y�������Y����A�Guīʷ�-8�|���/*q�@��VԽ�U�J���6H`���V�D��Q����l��LM� 1�dW֦O���	�7.Q�Ѝk�cx'_�h\#I'̆��Nc��)@�lۨ�|�����"�:}��0��h�vo`�\���=����'X_s�E,<�� �-=�1�DZ8d��]�B����o�q��a�&���Q1�x �?��L43�!z$�>xUX��z:^�n4�V��kh�<C� YDQu��*���}�Ƙ��m~�:��+a*��X4�U� ��|տE��l��*�54��]�� �:v�-V G�=!T0Iē���@���.@:�O
��(t\zo�E�[��(�ga��A����ї�>j���kKi�sl��l(щ����GI=!�pP�0�!�c��W��r���48F�P��^��ǚ'hPE�<�R��p{�Y��~�MD	�� O��B�����ĄC=��O0�7[|ܑmg_ Q0�F;Q���
z���a�H���<F����F�=�Ւ������^n��{��}����Ǉ�}��Y���~�8���?���ec�.�m�p�j3�3�9}_���Ԁ����;��;�����:,[3{:�ϐDp�Kw: #��QW�2�o�䠍<��}o�(~�_4P���\E��m�V�͞(�l0�	��x"��t�,��}�9m�+h8�7�JhX�':���=���C����� �LS�(r��V#,��xjC�>-Z}��f�,�>Dl6m����N>��+P��z�����|H��[��]�s)�Wy�Ptt~H{��X�H�"�{�h�O.Zt��uY�'0�ϲ��D�)���N�����ŊpJv�v�b�Q��2TX쎈`�pP����xhHsf��d��K9t4`%n�5����oo��� �������6tC��v��~�G�m$H䬜�|�<O���h㰔�JwpX��ɛ��L�wZ���_Ygl` `'̙�Ԓ���6D��>|̶���1k7��$�.���i_���9h1�Đ��r�B�H�OG�����U��-7�x �0�������~U������T���G�.���A�Q�O���/�=�,��Y��!]���XGp�M����*�3Ǐ�V}��s��Ȫ�Τ&ї	`��^h:69Ìz�t��4l��ō���&`��8uS8aE���U���X<L��su��n�Z��`�#,C薸,cH*�\u����c̞<Ɓ��E@�Hm���>� �'�t�6d��eQo�T�%�m�D�jM�N�\�H� i����!7h�τ�1�RM����9ǝp�;����^�Ө�����V�~����O��Y�/5�o���pߠ!2���>+�֔�������R�`m�
�gD�l��4B�/I\�������.�����EB�>�$�_J��3��k�(�Xl`�O�6���<��%�?���kb3gN�k�Lw&�s�2$���V�vF�*$�U�Ί�WO;�IWF�U���
6��$L�\/��R;T�nǥ0��l#^�͞k��=Q�e���|�r��+�#'\=p.K
�l �l� 2�R%A�����E�chtډ ���NE�[떐#WљV�������7H�M*�Ty��N;Er���؞Ԡ±8ϴ�X�2�]����G�Z��;��L�T3+��l�ƛB�9���^Ss_�#(�����9	��+1tI��8�P�'�^�����B��_-����*�ID����:a��k��(� t���.���5WB��w�:�rɐ� h��#0����I��ۨ�9���I��[@�^䑾����4��r�K7�\{��ë�c���q��e&�MauF趶����^&$��v�޿P�z����R��:��="lN�M<����U���t�)�FYT��tԻ�i��vUӖ�0��*ԥn�����>(		$�Ft�i�8!�I^#���1ډ7:0��ݮ�ŵ�a�~y�Ҝ`����t��,YĶZ���Fe-�䈛����<�r��u� �A�@���V���a��W�t����ϱ����W����t�+'Zu�D���^����U�!��P��	��5�130����ӧ��5_{�8����Om	���CS��A��&֑��V��YO ����� �5��QK���`}���� 5��RBz�p#1���:���������W�r��"V0��U���w�E�ߡ�,��v�����Iѻ���Vq�6�L���-ω:UqM��i��B�+UVs&@�J	��0�m���t&�sJȫ���H�ߓEk]�~~�7��K<H�
�x	Y̠�al�`�d���wAbx�C��x':�d:���nx���4E��~�=`W���<� �\eB#гv� $m ����.�.����d�`�?#���8�:��K�|�5�f������R���pxH�=]M�&�js�[��J�@���g���[O��t\�P�F&���a6��RS�b.:�'�4�w���r�.w���?#�㒢���f����
��ǰc]�~��ouh����Je2P��Z�������"���[	 Ę,�i����EP�m��yS� ��C(?wɂ�Ufж�%����&H�P#%z"Е��b'a�5��
k}2�c����Q��@B.�n�����ǆ�m�˞g]�gQ'�ܐvV?8���x��Hg
.�mL+���]�^�~��Mp`���QO�U��|��_��Bz*��IN?�o�vC���h������&��`� ��j���:�� A'�K�����|�{��P[>�!���~K�!���{��lN��6K���s�`�+mXvu�l���)�6�ӭZ��KΥz�y� ����
���jѯ�;�'�B�6�;�:~ә��@�����'2��Ʈd��:�hc��,g�Q*b���~�ae��o�H0����@'F�H��8R�`?��°yL �r|M��c�ޤ�)��9�y�T���/a1vE�W-$FR+�U;�����C�c�H��`����w�v�]�=���C$�fd#�o���=�O�\ze���ksgԒ�d��%H���ǣ(�veF�(c.*	�UA�h(sH����%�����AK�5���a���d.�j^e�mӔ �w<B�C��lw�Ը&��֪��J>��Y	�!�0�ܩ�8\������OAC��*�La�����lk$�A���r�C��Z�<���1"j�j
j���3�AN���^�
������UTU���o_]D,����ޑڤ�R( �+�;�6�B��i���lw}�� V�j�|�*�������C�؅�uU4�ɚ���]� k!�`�샥���8/���ն�nE����w����k�~���$�9�ZF��k��_,�@U���f����D�"#�����AW�Ɣ�b�L��q���C�xz���*�D��+l���'�5�Tnjm�k&��!�t��	�q�%<�}��Yp*Y��$E<� I�n����Ť��36�{Y��<�2-ݯbt��.9���e0�����֕lN�z+�kح�*<�0��fR�;�\W�2sݙ�Oo�N^�H��CXb-��OV "�>����1^I�$�IҠHb�8�Z�T&¯s��q��`l@��ѣU�R�,h�s�m���;p�t���o
����S�o�Jp.!�m�Q[�ϏI�� �+���8��cQ�U)m~�~xp�EB���#x��� �������F�J�6VYD�G�_�E�=��ٝ���c��8ds�3e{됙��˺0��,+C�㗙���rc��m��b%�I��ySG**[�Zi�Ɓ��%-��7M�h�Rg��K����^�{h�~^�Atണn(Jj �����$�������O5W$�A�iH���%��;P^�Úz�>Kv�c�@Uį�9��S��M�@K�帙�0��n�&8��Z���t<�����y��	�f�~�|?��4�$����$��*��਒k���w��*b��D�Y�����D�"E�2a��F�ǧ9��xN�333��r�=Z���l��O���<j���y�p�h��="{q����	1qM����	ȵߕ��0�H�?0a�5�����ΤC�9T���4����L|�Qu�٠>eĠ�,X��:?s��"�z`��gܤ���ԑK�,�<��bH�>O�b(v�cD��U-�3i�����Fz�a;G����iLD �ߥ{z(�����O���8|���Ň������od������ho*�R�yg���Л�M���ZzIo�\0V��v\t"r9�zȐr����l.����J4��j�Z	����$�R��kk���C[iw�s΋tҖ�9&���`KP�i��!k�s��� �$#�����n%-Z��! �J�4�*��;��44�$���mi�"��սF�Ge|��� &����@/�g?�W6�,���Wt&����>J\���sӉ����Cf�]�_�}ڶH�
/�>��#���Hc ��� ���м�t�r�n2��o�~����8��m��~�׬����w#���*'/8�$�.��)���gO�Wba�a{��M)+b|�(���*�
=Z
w��p}���}��@�$�ze��"�>�|b���O_e��
�<�p�$�M���mߚ�V8��o�N�9�2���ec_����L#j/�!D˗Qk\�b���?��TQ|�'�S����4[y"��U����^�1�|�+upv;@�yINғN�~�	q�⭡�{�)�m!u�JSTM/���KPկ.B&��� j�9>E1t\���z\o�i����p�X ��������]%d�Æ��yn��.S�F�6a�}ST$�;�)��O��W_�$��u�򴠬�ۦ��gg��m!X���m�	Lo�m�`����$�~��KmQX���c�j@7����G'C�L�\4���H���
��(?}�>���,Pv,��,��i��i5�l���0L(Avu[��O�x`9��T��yA=ۑ��*��9����r����UW�d@r��F�i��7;�on�4���f��������/�q(��Ȅ�i+��d��8�6�:��y[%}Rp�����$#_Ȇ��%�P(�iŉ,w��qt�o�v�|�oG(���Bհ_,��r��&^\�)�,A��:x1���C���;�s쁻�����[��sR�������Fr�"�I��e+��"z�\'�����]�w5��ݒ�?{�߷�ngC�'R�^�@[�7�����؆IW�c��UQ���	�a��}S4`s��?tk��v�T8���b��[\���V���Mԯ�� �	Lb�1��F�RloA����ʨgf:T�����2c������>J
Ac���f4�A�!#���V(�(	/*ӱ_{��y�&8(.4��/�N�Ĕ3�?^i�2��N��<g��{� 4�˲��#
�ֽQ_hoNX�D��9t�ˑ����ʓm=�V������6OXO��8�ή�	�V����k�^�T����0`��wҙ�X/�N6���(����|���bh驋�a�Ysw{0��8���t�w����]�����}��� �^ＸF}_ԡ��_&#�lK�߳ҟz����!b�Ga?@��T�3W��β�ϝt�m &rӢ&�*�σ�jZ/du�-9�h�O�qA��g<���A%�	�YJa[l�uZ=E��	�㩣��\��ժѸ��؋%B�Aw^���S���	����~ms6_�� �=�����O�Iga)J�����*�!q��M�R�\�zk1�w�T7^U�.�X�]i���,캂<�3�d���T�"�${�A�pc�+�k�����|H|;f>��3 �A�sd��^a����t���+��^�M���R$�/�\����ZG���н@횃�d7Y&0�u��*�G[&�
��P(��k����l�@���M���jq�lp\�k�y�2O��}����)��_��Hb��CO��V�<en���R�?/�P!V��v�S��@1Ӏx�iw����<��m���cpw��w��s��.�)@��f�!x؏���{�@��#��@s57[dHTv��Y[r��-c�Oi�#Y��'�sߠ��x��10$U��>��qe3>�
nWN��&��Aɑ�g�M��/���K!���xJ���RʗҽE���Y�S.�M74�Q��ֱ���Z��OA�kC���)��ٵp%��Ⅼ���Nm>⭹����mx��*v��v4�݉�K8�����(�~��k�]	f��7
���!�*��!D �����(~Ĝ2�t�C��3ϝ/�4ݶ�Kr诨�o0r�b�Zmb�$��iv�AA�K�ZQ���$��~o=�R��GM�� ��4Q����'��m?��n4��pz�ĿR�7T �FR��Ĭ�<�)��KqU'�	����@>E�t8�����7��=s�P�!ht��o��v(X+�'q���+���[�JylQ�G3�!�V��h��n�Nx���{XV�Qc���o(<�oh�,���X".�)�Û[fGp�C[^���$�e�:(νAj���4G����y�t��~���qC�c}%��S�� ��6
T���
�V+*�4<XcA�w����`�
Y�؋�*G�O�B���H�j[@X���x��yP��տ��;�@�;��W�f�Jɶ�%b�����a����eb��w*`�@p8/�Y�
t����O�_�����'o��׋�r�Ɨ<�Y��J��)�G*|m��?-������j�N�QA�מeM	��ՙ)�5�'���3g4a�7����\ ��[R����k8���̸��\��V�G��Y��S���Q_�Qj�3!  \����!!a�SA��v�]d���Ԓ�y�)~x�J(8���}bk�Tf�ɧ�K|hH��f�_Ψ$��d�
	D.$&(	�]~\p�ofٽ'tu����-�mz�v��]�*����+c��o���\��Ń��`�N�G��ݎ��t�;��r��JJ�/��#�_a��!�F�U�#Z��� �u�R�����o� :&���q�k�C��CRG���Z�c�������
����-��E6� �W��j2�[QH��p�o�S~�t��o�VE��=ӻ%�k�{���5�#�\ $��H����pG� �j����4O�g0��ޣ����<��& �-l.��������`oӻ*J�Εg�0\��_�5h�ՙ%��I]_�[ ���jGU�Tf�l��	�@���3]�O�C
��$4�Ӛ.q��v�f+���ՉT�	[X��1�7H��ӸO�S(�
ʋ��Ww�A�SbkQ�9�y��_yj��Q�����uש(��v�X|o=Ҋ��C�G磠zY2�x�ZưJ"�c��ë��1
�bj*�9� |ub�1� ,{2���&ڑ5�B��.��u����P����Q{�_ ��캌����9��94�k��8{���x�2�g?lLS��B�5��Kb�0�P8��Q��*Z�t��&�d)=���t�V$?�Lt��pn5���1^1O`]��:��+�_�Tt�͟�)}��FЇ��9���ɠ9I�#1�џ.����x.I�b2T��i?�����AY�@?M�V����C�������zx���&��Xڴ�����DX��QXS�#�/��Fm#���n~e��e�k���y}��?���k���E���1ꪣ��8�^��u{J[���,��{�&�JW�N� �&��,�\�تn��!0}4�\��|iWa)l�(����~6�7�g�FEĠ��,�Ц �혟��뉵S�~����B쏸��ԙ���:F2v�������뿒����=�����Qu1�Y�s}e�K7��]B{��>0�^�b��Q����Z�*c3H�%�PM��f�3Ff��~|��7�[Ns�>@K�DM���f=&E`��}���֛�����p�J`�?4ʙz*;hi�*�H�o�x{a��jU�p�.E�i�G*ma���|;*�^��O�YFa7s �	��܏w7Q����<��J7�:���}5���~�A�#+����*X"����o��`�`M�Ueļ�{���ĺ�}Qc;�I���4�	����<�ťզ㸤��>�$��,���->ؼK*��Q�o͑N���Q�R�Uꮷ������Α&�a�/�w���c��5����;�(p_m�������Ps�v�i���w���ҥL�o�!�Ⱥ�f�adl�I\Z)�(�WHkve�S��uMP_1� k�����SFC�="r�r�É��P�Ǿ����(n�����������[.��N�+�
���T����2t&I�[Y�W��9�D16w����Zü���B�b2)�����p݄��y�%i���A(���':Kzg:�0�9����aJ�{���zփ��m� ��I��N�~�*�zm����B��Σ>���,���h���a��^78�/��`�(қH�8���������u�D��R�߲�W�*5�����+����4eo���bo,���~�v�P�aΰ�'����g�݅B���pp%����3	� ���3
:�bŅ2�1	]�Ψ�!�vU{@��0w���O �])ܱY�Q����b�Tҫ��'m���xT@�!q��Ó&�j<5O�8�]����������˴�L�ݺ\���x*׎(w�+1�y9�?S�j�01����B�c�������!�3�&�p)�5��F�!ۑfH&�	��
fbV�:�bq�r�SS(�w�Tbx�J��+�rI��5Bg����NP�~��J����RAP�D�K��1`���h�F��E-�XX��T5=�Ȋz��۾�2����I�c�pTj���|^�)&k�DwKA�?����c�`�?�L��x�E����w���;���nh.qkٓ֑[9��P��e(4Y�~ͳ���( �z
G.�%��,f���[�uZu6�5��- .Z�Ȯ���}��h���Gk�9x���G�龍�i�;K�lڽ������#�@B��6F�\�w����<�j
�ACҠ��Oj+���n�C��X��q�(Q�G�b�Wl��&x����I��p��b6`©�}�H���X��g	lOx��bŋ���׮:P������hԭ�+�i ���\B���p�b������6hp��^2-)��sz�(L�X�ۢ�^rY������PI~�%�	X��&�R^���ܧ耢
Ң������Htd�.n-\�b.�Ġg)��}�c�93*)�(�@,<��7BNŋ��D��QD>�yx���aĎ&㪑�2.�	=��X�i�/����,�b���y��e�,�.�+s�"��P�hN3��}�g�{3/1�X�pL�Cg������-�M�!�Y�'��0�R�'\�ѳ���)b%Щq�}�7ĳ�K)��a*��+!�$n>��]��M��Ԓ�<O��w¢G������ۆ>!H�`��� _e���JSf�z����jDꈱg��7�$��kƂ���ͼ%�Yn5��rr����Pb����;���(ei�S�W��4�t��O#��׋��'o�Q�)I�9_/�P�E�5d2����Pt��<˲w
�S�NMqN&���	hA� d	% k%��Sp�ܐ)�S?:$1<���6�jjeɕ߰��R���|���g��ДUfl��	�_���x�R!��'����0��@� <�8Sh�=���Ǫ6�ml{�n�J�)�r�>�	���E�m�'@�^"�U Je�k�F�˾8�����l&�E���� �����!:�N@g�p��4W8�!K��-�A{�J�d�Q�d͓:�%�i@S���� ���״a�,c�6��4n&&��Q�EO���8|��`�Ж��ߩB��d��������/��;E%��I�9��	����N �k��`�~~0���6lU:D�l��@���O��<�Rub�£��e��g�6y?� ��A- T�T�Y��	-��/;��~�O�A>L�%9t?���ڂ��ю9��׍�T֌E�,�Nz�Z�A�s��]4�^T�9&Sh�}5�MySz-���@�|� e�ƭ2wT�2���fၶEJS�����ZP�	�^�i�6��ϬS�2Ȳ�5O�&��r
�.�N�����z�6j���^ئ�S��f2�RБ�[H�W0�(B|Y�B0H��V��	�=l�MaU�!A$�� ;~a\��F*������U���	��U #Q����1�����S6�п���ދ��dz������M��<��:��褢+*����H�v6�X(��|�}N�A�n}�Jg�M������s���G��P}���ߌL������R�>�.x�d;ь{ߴejH$�>&Ĉ����H�Ǹ���A¾oap/$��ɗl]`䜃i6�.�O�����]8�}`W5��|��(H�Ȉ�W�B2�������[2����}��!�_8�dѷɫ^pAK���ج���8��غR�+�!����p?"n���A��A�C��h1ԝ':�.��j��*Ϋ�F���f{&E�M,�>N9<]�	��a3Ě�nȎ�;��N�l�B#�����,��X̞u�j���X:Ln�I���`>�~�ͯpT���2�9)(�c�6,�,�F &�׀aQ�ˍ� �t�U�xh�Oy�z�����#o���,C�C~P���6v���\�d�r
=uȪT�CrknVq0w��w����mu�f�%��3��WA��m��A����Z�kS(}��I63]�-<t`*�67���� � Np%ϗ�D~� ^�V'j��� /u���8nS������\O��T�5�ܒ����h�,�7�k}��
�'�a�L�p�FK�b.jr5����似n�B�܅����j��J���|�^&�0Y�Ӣ3}�e�9�b{��c��?PX��d��8yX�&�s*t��x,ۋ��n�g"�7d��&�`X{/���MlA�|@�Z�	sX��� '�I��H*����!:�k�y������l��T}~�[{h3�m�U[��FbY˂��Xkuj,(J��
b,��͑��P���̏)R��pÍVy񻏹�`"L��ݜ������)��Ӌν���&��;9ik}�[�����r4�����V&<+�ڳ�&Y2�Ѵ!I��c�0�.�G��\���:��/إ�<6�(e�8�D�_=V�H9��T9���&DbL�ZjOe1�C�a��������Ϳ�4E9�y9��^40�Y[���ޞ$Z�y��!v#c�P�4"�#�~��V7�g���\yҍq��҄» �~8w ��t�߬�0��<�+/fբ�`��}	3|�4̍o�Jr�)wN�
�Z�y��bTh����|���9���c-,��|� Qq�l�w��w$���h��ʭw�N<�N�Tw�q����M�o����s/
��;@e�Oo�.��Fҏ8��EL��z�����;�=6c���rh��<6�R~�+�<,�!8B�ZuK�.����:lb��A��o�Z\#IUJdM�wQP�B��㓎�٥�[Ha*ڽLc��G���ൡ�@s�kئ�|˨�{���v��a�M�CD%��NsH���XU���5���8;��@�}���L?0Co� �#c�Hl�5藫ڳ��Q������f��8@�%�ɠ��3|�cB�\�q��ր"�=�<�J�A�.�M�7�D�>� !�8��4l�ԐV&'��z�i���9y��P��%{e)�Sc���CcW;�
�r&�*�?N�y��#�i��	��eF3���*7���9�
 �t��>հ�/�|5����8}nK����=�x�ڸ�u�wdY8u�u%��+��N#>��oMQhόS�PV����oS3��Bk3���嬎���~�#��W��y�X3�생����Qb0=�~��h�uw328��^Ȍ$���!Sqn(�+�ׄK: Z�}�P�}�+��tf<�c|?��,�$���K�M�\�Q���|0NUJre?lb(�:��fZn}�V;r�m�����;�r��:B��u��4h�XvO��@�G<�g�0>�E�rP�m�Q�l�.��7h�݋79�5�FFhcd�,����՞0�&Ǝ�� V����{��Ρ�$��E4|���(��?�)��;l���C�a���čQC����{��/�q>��*x�N=R.'��+[��	a��tӠܘ��
�Hv�u���w�:V:ߙ����1�r廎1�[㎆�N��m܀ʌ}��6���+�� a�Z�iz��to�躼�^iW�Ѡd�y�|��TF�+���b��^�����-]�@%M?C�ܩP������l1�j[w��m܂�����O���[�R�������88����s�;�8 �� �D}�� ��F���fĝ	�Y�ظc֠�4XLZ�:ǁ���[���SW=��CgC��
!�^W^��������ZM)Ё>����d�?������h��]8�T�+R@-P$�w+���F��,P&���z��t
�R��f�a&��xg@Էg���~o�Bua���b��WE��B Q��ݤh0�;N⅄�q
>7?�T�9��Q<�\h���輙�v�2�/|��=pt�iv�p��F���/B܇sa��oK��D���YjQ����f6M�JW�x����?�Q�m�٦oʱ�?Y��`�6��7+�{��\�C>E�(�/�P_#!���2���wیިmF���𧐯�1<|��=<7ea�� ʼ7n�P�X��ޯL�L���:��;*_t��	o�@W,��0&����J�c7܌�/<\�T�ͷv��*���罁�[��z@o��bGB�5�8�c��=Q��D'��a�:��Pe-���|�v�юU�S>�q�{�
��A�ȉ���VQc+Հ�(�]|7|ٟ����0�7{;�b�QH����!�D
�1a�E*�k	]������4�8�C��:�4�(څ�p�Ƅ������j)����<��J���5
oQ��P�M�\P9���/t�'XO�\O�]�/�����u0�h�����6Tx<4������?+"E��f�N�%���X.�qޥ����:��C��b�	Rc�	ܚ�{Q �C��B��`��&�zzZ�Px��{7�g(�r݆_�"�%�m�+��W�����t��,@]p�㵠'�O�R�kA��N�ŉ�4�@���h��8,�d�NC��Ʒk�� �.z%i�Ŀ�b�B_����<%ew��2�ڣ�o�vq��l$4��HB�R�l!������7���0r��dM�ӼS���Pș���a�E��Ȼ����x p#��ɗ�})L�������]V�=�ς��)⺓X(����J�]�K��G��t�ɇ�w�l�� �,��WH����p@T1��1����^���["Jv�	�
ĳ�����iQ��x5�[��Մ��&@�(�mh��%uNG1v�6���9�K��C�Xqs;�k�Wo+���f(Y�+����;��#�H�upʕm�sm�$�J�ᶭ�r!���I�_=���������b{8��#:��9ޱ�$���PkO�X�r����"i����ي�^Bv՟���o��WhK	L�)S�/KVD񤢴�&����ϬW��p�,���C�a�Ksh)M��/��	�S��y�D��x4.=�����ʰ����0��QGW;DD�VM�U�5���p�t�wz�`9��/X3qG���t��oK-�+�CKu�9�6|}����'E�$s���\١#)8���P؟]B��^�������}G␱ *�H�6�k�"�|� ���.J��R��\�1�ǀ��:]5�3�S3G�̆�[�R�`��'t��&��Z ⌼n�f<�3Pj���'���d|҇��<G.�Ρ՘Cf0K��v=f 6�<�EE�,� 4���2ڶE�7<�#��)���~�RQ�w��������x"�b��YP߃<>,"�1����m�Qȟ��\�yCc~k�)5?�EK ��(�y.�8�aw ה� n�9u{�_��gq�PT���v��u�o��Z"���"�g����c��S���7���/�c�7W"�=2�;e�Lf��D�|�ut�@����
�Y��p�׊T��k3 (�R�������o!!�	�@�R3����U�و����yp���q!���(�B�OY�6�80J'��vM��J�#�*�y���f��,�w��
?�
E�~��$��-����;�����#2	�Zư�ͼ�����H�O� JKˌM���x�J)��y���ppϿ��422���P qt�`x�ё���5��l�p���	�{�m@���2Y�Ju�R/R���A=��|X*� ��Gk�ǀ�7��V��묧����2ǹ�oBqfp�^����&z-�A+a��{�T�Z]%j0S���e�D�d����C5���ro�#����
)���$`�s�l�P�&+��Eٙ2����Zg#}������*.L�Wt�.Ǳ�n��v��h�V9���O��R�-p��rE��d}�
Oߵ��BAG���s:d�KV�00,Η���O[� ��Oj�Qr��rϟ����9�G6��"�$��V��W��n�ǃ��<or6n��ċB��ʟ[=]W�iB�$I2�h��@�����׋���i�������q����]G��W��j�uh(�?ͬ��$v���so0<�����$e^\��N$E�V�p����'�7�N�S��>��Ş08�Pe�8�4�F�ƴ��M�:Ao���<�Sw��_��Yc�^ye��WQ�U�rW;�x��&@�w�q�[��%���K�#g��Y���0��Z�r%kR}A�Ѣ�$֫�_m�`j!�%�sS��G$��'ܰتshqY�D�go�Wa?���Ѽ�Tۺx��-P��2ݺ#�A6��Y.=��H�������,�Ҭr��A�ޛ'�-�j�c������qMQ��~Q)?�_���,�>G�&?�e?��iEv_&"�ɂ+Q&���[_�p^����ǔ�l�`�	�빻�5$��lX�2D�n��н�lY�҇+s�J�� V(>B�
f$�@"��i�d���8ۺ��/e0�)�������_TKV�#rf���*����0��`���R����_n�1h��j5��Y��zs�t͗� �K�SΠ��C��y�(�ςR��v��(M�����5_�&�jz?����������	$&~1<@���śu���L�QkH�G��	����4�bB���|�;����'���Jʘ�K�K�!m�e�b��1�~ ;imo��M�y�S���+I�x�̗㸣�]zO�rշ�t�xT�p}�Dj��fx,"c��,��Ο}{ǶA���i��T��S�n<}!;#�q љub�+���*��熵���A�)�O��e�~��J#"�E5&��R���5�Nάr>P�"��ݬ����N��K�,�~G2����\Rzo�+�\�UT~u�^0�M��}��)���W�"�'�Tp��6�
�q7�G�������C!�����,DMl��SV�9�[=I��40>O���L�ÿƲy�R��^eyl��	�'����҄z"�%�l?��㏏��L�PRZRG��m�ǒ0��y�eG߹� ����Ք�����F�ˤc2�m�X+U�`�iV����q�1=P�b[T��f��rU�殁[�(��?x[ʣ�	G(i��s�\���OcYh�n�
Tұ�1�<����~�����lgV۩鮾����Go�]Y�8g�O>o�d��@��J1�4�_�:�a	�ZO�7�X2�yv�ʙ&+�Ʌ�5p�*���N��iY�L����[}�8����~�og��ƴf�x�e�@d�z����n,0~���G;}���A�C5���z��z"|�l�ut�08�F�)Up�lׁ���>4���,�Af>��i�<.j��(Q��h���EaL<�V���%t�C[�������A�g�w�C�~�~���#�(W2p����B���~?i̛�vO�YG����
謾|�-�����S}jaE]?����Y,U��3ʆJF��id�얃�6P#P�˖���f}/��*�t2�"����c��.�����"OR�n�BU�yŉu@���X��s��!���,�@_�P��
Μ
�f;�p�S�j�x6>1K��s_}�8S�O�A�>}�I>���I;^t=ɶ#n *�+}D���I=%�.���f�"y!�\b�3~hSg.^m���i=�H����k�E�%ez��
џC��V)8���������=����Sn�繚������y7Ke�o!4��.~f��g��ߺ�=��G��PМ�s�tq��£T������qώ��xFž¤{�9w�D�=���~Z�6y��݌���� <��\S1��*9>	5gkacS��� ��`�[�l��cX`���
+�̯H�����E��|-ʼV`҄nqm���>·\�E�+4�w�M���3�:!ݣ+dƩ�u'�V[�^w�N��h�{��3����BA���o$ɖA�6����ֽ/�X�0V�sg�N�`q��� wǃ;LՕS:'x��bx����ײ��<�B�>x������1�"O���ނLz�����n�M@id[��s�Hi��E����6�/.ģ|Ce"E���~S��9,[�x����K�����S�kEW���(U�ڗ�ug���a}a�Cͨ,����֪��:�9�S���J�@�l�0�/������V>���Qvl������|;�����DT�~;�2tJ��Y���!d�B��\�^��?�-$#%�O\m(J���-x��eo�RpxT�p���:�&�����~�b%k���%���z��!���v3R�����ԍ}%���aFi��WhmW�>�l�|~����yd�to�c:�`�����\�B`p��<�6�,,P��ÔL�k	0�����2!'��qo|P���9�b�a����P��ꔙ�=�C���n�l��>��9��F���K;�HT)d"�5ց������{�-eI�����_k:�p	�|�M���SM�ql�ƧF���eV2�?���z<̹���p���J~�ǱO�E䉣�VL9mZI=�:�l{��5��X�Ϙ�]W}������!ȉ�YD�m�鼢Ɩ�]�ǰ���5�dc����s&M�ٟ��#K��	JƏ��q>M9����/�����sLZ�Φ�w���L����;�̾oDf��l��4�6ҧ�[p�v���3�k]$���98'י�1������_yQ� BjY�� �v�
�P�q�=�M ��2��6����(M5��?�5k1��!z������T���԰%�D�Y�L�9�h�$�����.��r����4V�~��QCX���1���ڂY� G�IN"tU0M�ZĮ�����$�~�]k�'��_N1����hTqT�s|��e�Գ�����=�������  ���]J�4��#�k�s3�(�WY�V=n�>�~8�D4,}"%Gz2i��K/$P{�7��L^m삀d��t�6
��.T�`8L�[�u���u��3م��`�w�O;��AV������S��D��~mN�Ϗ&����_�ɔN��D��A��8�� k@�����g1))y��$ҵ��k�~��J92i:�ꛨ���=Cz�f�[�yk��n����}~���=�%���_�j悬~��B.�N�Ft~���1�	Y�&��*�4]{�b��}����>�4��CM2�&G��k����}O	K@���Ѝa1.�%��������]Y����{B��h�+��]�$�Zv4I:�e]k}l�]�W�oi4l��8�O�����E*�~*I�ȶkNѳ=,�`m�O� �N���AuBGc;?|��,�Xi7�a��
ˏ7t"jD�]MC���?}�JCX�*� �5��!�ʨލ�N�A_�J��A����I�(p�J�x��8A&���X�F �yWڷ�ѩ�+(p6Q�nt���)7�zJl�ص�nZ���:����P<33�b�c�p�C%y�6�gWb4�9p���r(`�M��Ƿdb�ۇ���#;�Ago��~B@M��K�.�8�װW*%s��F�����-�>�Ɨ��oq�����k�R��coo��%������|�_��Қ��Mw�응�Jj�b�&q/l3A�I��vIn�)J9$�ȲzΗmq�XV�x�<���<�u\���7\)EI��:7v��1[����̌&����&?�X<������d#y�.�jk�⹥�f��V�jԝ����I��b
�^bqW����Q�r@��N��}��ٺ�e���R���iw_�[,��d�gh��=�-�_X�.?��?���*�",��)��/{&XdG�;��1ˬ;Ѩj.���+�(B�d�OX���'C���O�jρykϢ0�NO2�/&sQ�8���Le�/��3j��w�pN�K^.W���\�r�.�������y��E��ȱy��#ok���X���B��~ܦ�2�?�0��n�th���"0�[MR��n�mR�ķ��!Hs4��&DAWm�+ͳ핤{�?�萬��}z��S��f*2�/�j-�W��]��$e��P
�]�q�q��̉q����?�
��2Ws�9��e�v����_���@����ɢ�?9�{����Lּ>�+�)ٲ���������E�������g�OK�su?s@!�������\|���E�l7Mz%u"���s���º�
%��S皩�(w�$�!/���
��IX���ȆwǛ(m:Ҧ2I­�.�%W�v�����̋�}Iրڛ���a�U���tҢ@��,ɛ�s�O8´b�Sh��j8lr���M#x�)p�\~�[�eS6�s��f�Y@�$��χ�S�$���$1nW��b�4w�D��6���EbC"�u0�0�/5[�%�i��\�}��[���.�m��o�ɱ�5����r�������V�3�I;�~nt�%��}�a��jAA�^�<�c�`�yhP
.*��EZMsl�U��{Ȩ{�)�E����zw��n�"����1�?�&�f��G���	� �ԟ��۸�s�=���� [����H��[ݸ=?LI7��Hf&�[ˁ�2԰S�k��r��(�s� s��޶W��19j����!�!�<��2ٕQR�J���2G��W��'S�`}[���n�tc�S��#Z�Y�f��1�p�ߍ�k��f� ގ �⥠!�O�A���Z׎�+O��v���q=��^��Dk�*,���2�iȌg�WT��D���ײ��d�aY6�ɲ!�r�-z҇㚸��qyA�Ap�~��K���i�P�H�Tߛ�mݐ�����eJܷ��;W�b4K�̖�⵪���ӝ�/������|Y�ʻ�Qa��+T\����1;I���D=���Dmm;��(�I݌�"��@X����^���Y��W4K �6��^��v������T�<�[$��^d��N��y�;mC�F��N�+20lz���!%"PW��/�ۆD�r�����j@����f��'��qжlu,c��4���zJ�g���Kp �W��ҡ�S����+�^��'�����f�����M:Z��S��̆z���WT����y$�Ap�un�#��w�N���d��%
ql�޿�b��>��f6�&�T�-�����_I8�'2�>uxt��j���?��w)�|:q4eQ�;7��R�@�YW-s&[wHL6`hKF@WU����W�N�v��cm�-E�F���:�m���dh=� mP#���$�|�T^�A��O]�ٛc�ӑE�}�A��%]�\���ְNh��k�e�����|`ƾ��ph�<�A��QJr(f
;OLR���f|�m*�O���oT0�:3��Z��iJ�M��i73�Mi2�� f���� �"<��m�'��YaY�ί�#o����;K"�|ȐZ��n� h�]�Vo�	SrW��t$�7շ@X#�@�s�J���Z`_�eĉa�Hieek�<�Y~j[�ݬ6(��9���y�`�ͦ>��n>��t�5kޜ�fE<	55����l�2;�]����*g�]ӆC�FR�Dթ������$�I���X�q��Ō*�Isz)��z�ML���4��?�3�_�+H~��;z�+�-d a Ë.����*���e/ΨJ�)E_�M��q_<�ե/Z����')0�E3r�j�y��t�d�Fb�<�@G�?�5Z({�:%��Ԟ�D�A�o
~�,�͒�9J�'��{|8�^O��O�>š/ y䷔��w��	.��W�c���܎-��ކ�n�ZEf�&CD�%{�X�#B]��9���Ew/�^!k0����<U��B����g�$��ڍ"�o�K��;�_ٵ��� 7)k�k \�7:��iȀi�`4Z7��6tY(*��^�����U��\����A4Q2�х`�Z�� �A'�\C��������,8v#V��f	�V��ss!�?O�Z�6q����Et@L��` ��u��da�k���!|�w�p/ߺ)�,p|�$�6E���(��A�gN5�N��O^,��k� l�lr@��'(]�	ۛ�zJ/R7�s�8�e����H��="9�CS1��qlk~��Ӏjg�*�n��'h$��/ғd��ݘ���>+G��J��8J;%��^�Ԓ���}x�Q%^2r��}%�R�(��A��8�^{�d5}vy��L�<p7��;w^x���~G��;�p���|�"Q<;hT���ib�����C3���e�U�Ӭ�� ���D��yIQ����ͻ>�D,���N'�1������B�F���M��߰O�0�5�K�d��,��w�$|�E�<�Q��/i�Dzӥ��;t�xiq���9��rd���} �w/���yy't~�㛋�<17�3�A�ֱ���)y}��Ny�'����o��� �q���S�%
�nW��j�hI�rG�9^	Ƴ�pb�� ��H~jvEѲm0:�h�zG����ʁ�-� E��G����R������F������!�aI�<��.�W�A�tLJ��{��
�HZA�۶�㸃�U������Q5y��;�����I�E�:A�؃���=%���v���R�n�tz����5�'����_,H%*��}�] wc�c}xL�n�`B���Pt/ƍ�Dt%7�ˎ����h�4چ���֮v@�6[J[W�[���h׌�$q
��S�k��ByeL����C�OJ
7P9X�n��� ڧ[���%�{E�z^����<�{~E^�0*>�b��Tkd�'ޠ��ZE!� �Iб�1�G���TY.'�&{!���V�P
Xq�Q��A��-��,��ߋ���_ndE�l�(���Lm�N��c���_0fz%�g!�,�G��.�a�ی���̟���C�%IbwP�|�m��@]Ur,�[�X���0ѽ�����*յsY���p�sh��Z�^�qYVvڴRa^K,�L�.�mf(��D_��t�k+�]��\�*@ƒs�~.�']����N<}HT��>�4�U��x����='j�� L�"�>;I>􆙃��C挙GL
˱+�Mn2���F��~�,ֵM�-+��d���B�]�J���o(q\�����qX�e$i���=���Ʃ�7R��SF�����j.80�&ZT�C��k>`m#�Ө'��y�դ�j���X�wL���>������AOuA`p����N� aF�1��N=��e`,̀��[P�R%���>Pq�q�դ��uK*��
[������@��'�����p��̉�S\�NN���4�8�}'��G5�SF����o�$k<~��
�qؐ��� R)6̋��8��A���8��~^1A""�}������/���_�
N�������FRs��6��~�+v�t�-�o�f�Y� ��D�n����+_L�>�9-���IEl���j'�#J��"is��=��Y��LEf5T��G��+�t�u��]���0(IQQ��P�k;�(�%q:/�L�eBW��iC-XD�a��Q�p��\z�d)��~f30GG\�F�����XTvF�h*���3E�Ьh��gj�����8N���e�� 6J�D"�Ec��-aJ��HH��no9?1jP�R�]4��|%fm;�{tn�h��X�lO���W��,܏A:z�^�m蹀W�+x��IP��d���eVd%�tjȞ��͌���)1�$�~!볮$�RF z&�������0�%�/J|<�+��ަ��W_Kкӿ�42�-/�Qs)�e�9�S��r8I� ���NS'����P6���Z=3�M�z��>�y��	������U ��#Ƕqa���?�h?�x���d@l�]h���!�1`(�(��W�#��3Q	�Ma(l*�
^��@��y`��OPs����,n�
�{������p���xDQ��D��(oݣBQc}Tk�����,�}7�Ŵ��5�4�Yoxd��Q�T^oO!�������x�+��"u.���Q��?�3{ ��O)����4��r���1�z��V~f��,*���2����7��cN�����&������#�	�����u5q����cb5��#?���}�2%B�M��1�O�(l��-��"�9t:�0"��:FE7�Fk�|���|����KЛYۇ���%
�6`�؂��slg�@����/�����g����I�oz��duxX�q$��j���K��"s1\
8h�x���b�_�w��z�Ro=�;Yfܖ$�|�r=��b���xPLx�Og�.���䯮���@b
1���eҤtP)�0�|�,��V���dY�K�ؘ�����X�cK_kC�sM9����v�K�P�Fs�
��P�9֛��sA?s!	�-����*��]��|qh>^qF)�#GO�pFm���2��*D�]��y�,AO=��x7pT&��P'nV��Sѣ>V⪴�ꓔ��ߐ*�,sB��fNS�6�ȧ��$�Y}�3V��HB����t��W~�I�6]L'$�*]��hUi��1~��1$O�em҉ ��b{'�5bI,Y�8��H]�Hd���W}��tE*˖v����QfF�*E�u�+��%Q$lxj���� �����k˕�D���6q�k��݊�.��r�μ�-4�t<6Ba�F�W(�D�1}��n@A3��hZN����s	ۘS�4o7�/��5bU6"�82��qN�,���K�V�����u��-�%g��������Q�I�y��ic�����g����G�h�c�����,���W�?���{'��E�q��u^�Y_[���hM4ؒ���a�δ��� '�I�<�?��߯ ���6RPЭ�,��I3��І��qm�`��hM�� ��?��܈�~8�u��ƫ������J��|��eSƎ�Q�熝'aG=m7ɶ[-!�5j*G���R[�����)3�|V�h�6��F�����̰n�(�ܦaB�2$�v��GU��C�ܼ�҂�=���A~^c�w�R9�پ�'�1&p�w,�b�Ax�k��sWu�����ʈM/���`ӟ��eX����4�ƟMx�Yn���+	�j�$*O��m��=��L��tk[�&���������yt �W#-g�Hb�W�Fv��dr٦	����ݨ����8������~?MoJ�%U_bݥO��	�L�ƎV1�"�$�����8�kņ�
�c��
�t9�J�1���;��:��'���n����Q�)˝��E�
��еGm�����j_7%6Sz���� ��I�*���t�f��>���*$9"��JP�����,$Y��ț QfI>�L�?��Ο���(�ĩG�2��>ŝ�"�D1U'o���T���z Y��F"��ۙ
|~uMi��hn�N�Y�rL2�\P���^���c�b��w��W(����^@e�����H�-oXL��X0�U�s�*��6�B�J
������=3�@s�4�=G�ΰ\0�]��Ԧپւ@��ux;9�7�t�~���O���Z�X�4���[��?s�tժQ�NN�HR��i�;���+$��"i����kփ���93��	-����v�6�JK������½���lHUylxl9M��W>�Z2N�o�e��o<�~�!ڌH&���P��)D�.�,�>�}Ř")k
</<A�u�Z������)t]�����<�oM*$8`�<�����an�{��g5���;z��~�Z��78g�%R��m=:�+l�ȭ)����4=�]㵬W>�	�k���Y�#�x����N�B�>.}4�$�d��<��8!儫��Ӹ����;�����o��!=߶B��4��yi?���u�V�&	���Ӣā�1��@��?m�l4+�V$"
�������Zm�"��X�C	;���'G�*�3�z��"�"�^ϝ5�)����&2�W��2����H�2U�hy�$T|�*���`��+>�������i)-A��ftslrQ���~�ol�L���~TL�������(�Q8Q�4޴�KцhyԚ↶�4�d��:!�H��C3:�rE^f�d>ա��c>@�7e�p����h�s7���-����'�V�>Pݞ���;�Y^��M�8%C�	�Q\#S�Q�s��R��D�#҉�k�����HL��[�8
%A�W梙��		8.��!T
���/er����Gw����y&G٪"9�:,�H�,�5#�DÑw�VFK^9�?FD�E6�z�^Ė�X]�Tt.�˔�J��7�v`q=٘�4�]���Qd�5�>o�<q������3`�+���F��Q�Ґs�Z7�:K���uM����`H ^&2Bİk>	(6���M���4�F�Um��M]�K#�:�ϋS|�K�e��Q�[-�cѧ��1�Q�&t�Q�qA�+��9����<�X9�-D�)�A��BW,�JB���1q�����PV�I�M�7;-0���߼%��Ow}�V���5D�`��t�ҐJej�-�d���{뵰��wٌ�˝7*[����.�(u�J�G(�Mm�-����.�RX��z��x��yw?�uq�5�|�Ȏ2O����i�rB�I����ݦr�;�Y���u��u�W��"�.���ڗ*nI����?@�'u<����7?�ւ�!�����1���6����2O��p��������]�Rә��7bň�����3�qq+��γ�K�Km��	���JSR�U�G[k\�w���in��q[�N��sm"M���
�e�-�� �t�r�P<�g"��oÈ�#�1���Vj�=?[ζ	�P�a�R�΁pLZDvS�wJ8(�a4R8���Յ�J& ��/���@�P����ာsC\

%>0�x6C]�q45�,e�L�7�\)�9-��O?]D�?��=N6�^wbmF\��K�9����3��9Ѡ!��&P���Tw�����Ԙ�U���r��.o?�����#�]�_=�Ԓ��:^'ͥ�8�:�a���JGEW�/|�x��F���S�ZlI�sVY�H��������Q1�{��DG 
/��%��t�Z�i��|{!N5��/O��J�24�끕F�_����~8�ܣ8��4m�/�J�Kl�ґ���&�V����.�?J����I6��[�6���e��
���"D[����Z���3J����/5Ck+�Ռ�U��և�V�,P;[���MC�cE�H~^�	&�ں�QJ��2e%�a����
\nӐ��E�w� �7?J�x�J���4�H�n�c��V�u݀T�W6��&�Ŕ�p������Э�<Xń\�����OYY V'�w�y[A�B����6�pT��^����;����ϝ�)/�[�F�A���Ip�����-���!:�!�^�,hFF�!���m،y>$�s�]1�'���_�J�V3�Ʉ�V:y����?su`螁�� �@Ig��z�Yd���Tt&3[?ؿ�xf�V>���@���.��� 1�M	b-�&1s�m�c��w�@(%�W���z�U��~��H�Yə��[W���WGiv�$� ��s+��TH��}�Oi�0����������򸫂�4UD>˸�oF���v;���UZKf4���EH�Ʃ,YIH�8�@P�i�i�D ���`�i�{�ڴ<�t�+uKV^�B[,"��NYr�hY����}�GR8�"��p��U��bt�⇳#�<܂�>�����c1b�M���Մw���� 媻^U^��)Բ����؍5���L�X�&d������(>Kd�?LX��n*�9�0#j�/$
�18^����l��Yy���8*kXܣ.�����fIL�?4��k�`���ɑl����z�ϐ
n5xP3�T�6i#���,���3�xnd�%XU�
���V��d� 0~�'�?T�v]��_؁�´y�u���������4jq~��({�l�o�%<����up I약����|q��/O��W�45��a�7
�R{��%!�RJ%me�	e}ʖB�`O`2��;�WH�6�i})]mx���� ���@��N��Z��������'ꫝ�5�>uߺ���,
�$ǜ�ݳ��/���4�s�x�n���9JQ��6�䘞,M̫!'B�_m���7���PS1�Dϫ:��	���6����S�V�6�`qkl���V�,8EO�O�&�HB�����y_��!�N�gd�w{���AQwӝAZ��0�����i(�ϛ�o �����"��!<�h�ݖ�莆�9����THBGsf��B�:�vΒm�|����^�&b����L�2<=���I�k� �ۋ�_��Hy��xU��ӑ6W�p����<\�՛;m.�I�� �r����s����恪P�Q��i��3�:I8����1�Ŕ��R�;��3A����?�^��')�9�z��_���5� ��L(�ÄX�?Y�6���G*�'; �k�� ���I	8��$�T5�G3v-�?�+ƻ��?꾘Dc��1�]}��n�|�D=��
�j�^+���9e�5'�6R��j���eo'� ��B?�Q9��������#���:����p�{H� t��ڳ�����/8�t���E��h\�ǲ��i�M�Z6������K<�T#N�\����_6C5T[�N�l9@<���M�`o�1�/�ý�?0%��$4�	R��Kz��Rd��G��*������ɊkVQ�9�y�Dĺ�*ґ�7��(7���$���c���tmH�N�@�L�O�ŭ'��� ��>�z6�Z��"��7�Q�E�b���L�F9WfdCvo U��6���	{�I���q�wP'-�u��}u���x�5:�D ��N��⅛)$��h4)���_��r����>�,8�p�a���^Sm~�/JL�$k�*:'@\�hx�B/ÕE룿Q�!ų�Ǎ�f���7��Q%Jv�zueb�������W���P�e-�'���#wXK���C�O;���W���)���跫�z�_�����H�Ιi)ݍ
�.�~˞��Le)�:������<RM�X���Zy�%<;�38�g�"(pB1�n\�#W;&�����t�L��r�ֹ�[~F��~C'qTJPM�̥�c���g�Ĩ��)ﻖhL�*�=)�����:�,�'e�w3�hFv��tQRRp&t�իc6gJ �׺��M�4�*#�&C�3,7ۑ&WT�0�e-�d-u�o�/KRt��Q5��py��*a�@��$(W'�W=�QS?�kR_�J��=�敪��ɧ���4��2�Q8�d�<����Z\���.��`�
��*B���q�
��:��&����g�Z�r�j�v�pT]X? ��(G��y�5�/�x���fʱ��5��<�d���H�XýT�AԲ��ڽ��N*����U�]O�Y<�'��RP}�B���kc��2�3Kls1� G�J�����p�A���Dl���)չ�a�:�,�*�7+��(-��/A�O�~v��Ci"8��I�`|q8�1{W��F��A��z�Ts�.zS�����{�$��٧O�P��ݧ����I~�/K�\D-5)�8@�㬈��mؑG}�jm��j򰀸̡$�q��# �*k�M�oK�����+�NU7��.�4Vo�5�ë����(���:/��!�	>j|A�6w
BT+���v�����Y�2F�|�uE���eTe��f��F_:$�Z�0���Dg/��J�;��Z�2'`���]�Sփ�����ܲ����a��^U���1	��f��:x���q\������I:7�A_u���@n�V�@��B�!b��0�.,0MW7����9 �J�pɇt'1 �|K��v��&
�W����)��O���O�"uyG\s�c!�YI��
l2�F	^��Tu�[!љʹ:L/�p9��v���:��2��c�(��`Ŋ2�x
���X���:�����W��̟���,�Jhkd���mG:O�9�L$��5��H�8I�\���)��x�M�Z�e7�6�\s��G����dݤ��pfF9�ƴ��t$4�P��#:*��C�s	��"5�
�@	v���5�C�3�̯h�v�y��D�^ t�|��%�ᇀ;;/�����9��$F�/#�'����k9����o ˞�n�/�)�X�
����8,b�"j)�^S�!�,��w�N��¢�	��W��v���E~�kAz������+�>�@) 9�
o痫�m:@�ԥ0���i��^�ez|������VU���"
�v��6?��O
PLz���:��B]�<^��gD	��3�lp��K��_�l6j������;�����P-�7�cw��P�g�izO0FA���n3Z�r���2Sς��$���,�WCH��E���\Pո[ �P�V�0dP"f�b��Վ���DaYF��3#���)�7�Lj�G�[sn��RVA���i��5��!C=���׌�Ur#,�׷7&��d�t-�%�8_F�e ���@ҧ�^Z_Q�H��7]���ic��f��x�1�E�@��w��k�#��xG()!K'��h��qf�k���?BUA�}�Y ���U �{Q���g��;������o�8F���Qݳ8���Θ��ˍäj�i��-�ۘ!�'��p�_�>�K�zH�#t�Y.�TTZO����.�2X��^�֠�����~8���V�j��
�=\iV�ט��վ �}7�p�����f�D�u����C�;+�����ySAOp>�P1K]��[O� S�ۚs b 	[O�E��w��i.k��K���r�&=$�*�_��)���v��!.�m�Z�85+�f��z�R��d�:g��]��]{�)7�Q���G<J�d�ȧD�t�
N�E8���e�oa���7b�D�C�~��b~j�%�����ލ[|�t�.Wݑ;��>O|�����r�%�û7W^���̃�13My�&}�X��<V�\�!��fCQZ�7˨'+�*��917����<V�p̿�/Ў��� =y[��k�I�J��Uh�8�AnIZ_i��.b)�lr���[j�g~�Bbm Ž*�!����M݆|�cɞ�������܃��ٶ�M������a� ʚ�ƛ�ӫ5�≠
j�ߍ��s�(�i���a�O3�Dՠ=/����D���{���7d��4�m�}��~me"�����9x���o�)��[�L���/{�� �.�^~��8�~���ߠ)Jw�j�[�	[���L�P�|�*�F��W�$��p�uE;#aE��pA6��ɵ�;plIHh�vb���-�w6K����Ѱ8,�^C�m��K�@���~�2y7��Er��Îa�,f��3����Wd^�wY~�#$����\�7�QԒ�7�.����^w�LP��x2�!h�ƴ\��`+s�͙�ʽ�����*`��{-�5���Ze���2���ݳ��5�89}$�'q���&%mB�|��?F��K���K�U���lu����a�af��شUCT�i�|p�ʁ��V��#ೕ���)U�Z\��U�S%ieՖ��h=q�,@�<��:��b��Ldͩ���\�Jlq%ߞ�ޙ.�M�N���
\�K��Z�k���N{\�h�+���i ��"b^:�����0B�L=��P�	a+G.<)�*�Y�f
=�0��B���,&�w�Fj�k��[�c��b���w0@�lC�K��Lق��»�\'�ϩ�Ϛ�2�kR�먴���@��R�s��qٕ���d,/�C9�	�1WW�6H9{/א6U��݋?�y�����^��O�4�����J<&�y5���RwCT|�F�5=�pk���9'�����M�.�
h�#fǹF�����5Ū�ʵ>�j�����vY���;�����ߤ��L�ؑ���L6u��Y��z.n0���}�Mp��j���5� /�9���3CL�:3�O�|��m��
GY��5�b��Fb2/j>w�s���S�9��E�v�)8:�@�Kn#�^���'ݚ�6�/�! ��m3�h'�'�ng�#��26iE����
�^��V��^�H��rlPY�c#V����AB�y�LL���zS�-�I���1C4:J7�er1M�(P<儱�?�
�d�)�\��bkFB���z�:��%��#����qz�����?]Xd��0�M�A��7Ro�=��Ca:ǁz�x�'�쾲Q���YV /�<�h<�s-���|�1�!?;:�o�-�_O��$��D�K"��'y�\?_%ee�ڗ�K�?�0���7��#�����f$�?Ж/��4�>������A zV7&~�ȟ�sA�@[�}Z�*�d�l��3%,e0+�e���Ṃ��N�CFUo[�i�[<������	!9�� s�Ѭ�cT�X(b/9�]�Yi�|?�x��-u���[�p��Y��L;}�E8�8	����,f~�'zpB���2��3A� �����ش��~<E����W�.�����I\0|a����SGl����Ԟ(�n��M]���dDiu!��g�,�7|seן)�8 ��c�pn�Z}5<Dśe|��o����j�dQQ��b�
20[����=���̌7B���/��-;vg_S�AW���؄�`5�X^J�������q��tMe�q EI�e�����R�T��]h�kS@���8$��nX����M�8Y���Z'SN?P��)�K$,�v�[u�^��Vb:���J������o_�:*<�Pg�3Wi�lKa �q����DK��#L�yL�eBlG��-.>hv��%Aw�D�Mk �ɏr��/��>g*���o� ��$�ݿm���u�s������)�_wʾ~�V�����v��)���>:����9}M�o�(�'A�&����X�apx���N���]bE�Λttݔ�����Ř��0,�4����b�0!h
�������ე�PP6�8�;�Q�W�>��31.9Drλ��.-dE�00�k��ExL3�u�lG��	��W�Bi@�"��{���X�f�(׼c�MI�W���S��wI���m��fLg.���z��%���i�]Su*�B������F� ��[�B�6KN̻���5ɸT�ڙ�J;��>��ښ��|X�l֭��g95S'�kY�7�a�@g�=No�s\�n�O���N�`���'����^s92��)���~d�+*�oV�b�je���s�k��%[5����k0��;��!��d��6�J��q�G�񪉥��g�/k�48�}0ZpM����S�+9qѢ��O��q9 j�����o���Q��w�=�59y�cŬ�ո�����ĵ��t�2pF3^e8,%���c�����'D߮m5(�V�Q�$S�N�m�dSڸ���!�M� �Z6���ڔZ=�W �ъ�Uʧm��hb����,
���J(}q�qak��Р'�D� #0��>�۬$IkR�k��^ǡK�wg6�*�~Of�'�M	����ƥ�1��=n���	֌��l���f��|U,<�pۤ�Ь�e\�G,m����#���4��B�IH���	B��Z�	C?�ތ� �+���pE>����a,�3� �{����n��T��D�u+��d,�����k�t.f��}�O�-]y,��<\�k�],�ږ�]pw�7u��`Xg^>2��U��*�F�*y��й�����9|L<�v�"�bM���&�7ܮ\��Yy��	#���)�|	�(�Cz�>��=uAo蹠�:�-���q�Li�����î��8�+{�2�@��8q���#<����g�,�>���O3�&i�g���\�)ъ�]��@A4�E�_=)U���s���D�gШ�IY�����m<2/�/��~!޾��K\Щ g����B�N�Z�V(�9�x��������<R��	�Ɂ~ɲ�!z�S���� ��Y�1%��y�kغ�$Xl ��*�0�w����Um^��4�� h�k�3�Jd�RD*.K����Lc�.���꺄��Ǽ! i�h���hN��?��."�gH�E<���;7�ῑ���M)���ɒ��\�q�N1�6�?����怷�LS��N��su�aH�5 �!�B�]���wWڹ��`OO"���I1'�b�9��ڍfMp�9[NuK��?Q���$~�b�f:�pG6~�����6E��j���� ���R(�S?a���7���?�����
�,�l~�_���H��gK��3����W���kդ'���1�����Q�v��b���3���*�>1�'��tz�%��sI}���0ln�#�P�袦�ey�[�U#V�����ը��� ����b����
���X@HM�o;l*èD�y�#�]�.�X�ӭ�3��#�.�t�E~�F@��T`�f���}V�Z����lz��b6��L�t쑹vw�}�6�E�uBF�'�6N������4.��ȁ��ɶxa��D!�D�-�
Tb1׆�&�&��:�1\)�B�����.���C(p���qjծ�$���/�j(3s�o{��u�F�Q�dx�Uġ�"��L�j�_�E0g<�dA���~鋇b~����4�H�6^|���uv(�gr�KG����b�{x�D��݌[���������>��0�յ�)�C"R=zOX�5e�D�����V�Y���DT�d�~ѷb�����W~CKuv���^Q1��;0~�����SUĮʳ��m�����v&Y�r�J&��qT��y ���,s��A�P�te�/�D�V�q<�!���tP�@Wn��0<8p��wHru�Ȏ���1Ϗ1G#h
l�KmZP`M����`���l��/BAp��IaX���uc�ͮh���%()␬�mϊ��|�sx$%F�"�W:�DR����IZ>);ؙ��$��1ؖ�V��HG�De�9�-�ﾏ�>�C$B��1�!,����OWm���K�M�.��-h�7t���V��ZO
����`먛�(k/�ĚZ0Z��A�?D��]���vQ� ��9Ce/x���7�Z����8Dr���|C�Hp����M�'��s��
��'~��z�=�Vɳ���i$D�i��yA��%C�D���P|�(^���P88/L�cd4��Xq��#>x?��-Ɂ\�"ͳAY��{{ç�v`y��N`0\�z�� ��9]a�˻�l�-1��n1�:�������jeI%��Q<�`�������Dl����}S���-d�П1�{S�j�I}�f��T��{������R��Γv�ϣ22� ;ٶ��N����<:�2�6�K>�ހ���Q�4�T&
ƪ�0r�?"�� �xW�|���q4�^�8�Z|O1u��{�zDʿ���<{�9�X�;�P���g������ۆ9�ao"����1$���^����{T �2��w�y��r�k:�+#����1�4�W��3�h���٪)<�f舯#�`LMô�cA����6�+2�¬,�Z�ˮ�zi׎�@a����ՋC��S��k���tZ��~D��~AΡ~��!�OM�x�?�ω9�[�&Ĕ�V *�{�Y�K$c�w��5N(p�`�O7��)����	���i�Ф�`%}{�8jjc��W�p��N�ʱ��(�pz��o��M���Z�5#�a��ʮrB����R1��ܶ�f�cr�HT���r��~�)�?_�Rt01�H���복Suz��/a8tfO�V����A��HP�����AvKR���I��ؙ_XcBms��^����M�ݮ��C(%|	�y~y U�YuBK�jf�>X*6�wܚ�;�{���rg ��	}�J��ԗ"��M�0e���:p�n_+-�M�h�����HbX���)�����8���|Q�e�F���$*�k6�eLYEZa���f�V�FY>(ce��_��@3[�25���5��C^�ŀ�����j����
.�7P����+��8x����k�d$娐��K��'Fn�LD!���}��q_�j�]�
��z���fv��w4nc���@m���66���»?jo\����5H�j�����9�Dz�"`_�p`�k�vpLX�;�wf׋����2j��D�|���/^'|E�t�m�e�a��
2N�t���aQ�Sfc��A-�5���Q����������k�wk!rtgW�����_� k�UȢ��y���7�]�0Z=�=h�Q��	Ӈ�0,rs��A�7�����EL�3��s�Iv#�2�� 0)�����C:�kZ�)./��	�h�_��Ls�B8���d=�-*���=�m`�XuT���U�{�D��~5�!�nB�d�`6"����n��!�+��4�H*X%X>g�Ԋ�6��A��n�'�Ԏ�Dꃘ��z3�Ü��-^0g�s�ݴj ����;%*�g�v��e�]���6�t5QKG������}p�y����!숵.��*f��-���v��}AȒN�Z���xw F�G��v����Fci�]q�sp�a�&N�T����וc�C��/��=�2���,�M꺈6l�\�3��Nn���d����Ƌ�,�f���8���7�SyBm<IU�վ%鈃��7Y(�o���(�����p�!FR���e�dSo�U�`{�w
L�xsA�� ���;8m��"���5�ѹ�~'6�a\;��l��~������C+���H�x�zL�o�c@	"V�F�Ib�A<д���9N� Sw����*���>��*�˾1F�&�U�6±���8:a��;������3�WCi�ye�3D�;{��?�|��@�+V�y��̗B�*"f�� w�\o�}�3r*��s� �hX�A*��(4-K3I��|���������"�K�������vVVc*3#�<���qǊ��Ts8��ТQo&;�ݮwH<�֩�L� �0\D �l��{���qhi�u�n�w��^��:��HΜ�a�u��C�8N��OX9�b̡���R��o���+חؚ��uK����{��Xo�����o$��ov�Y|:������^ L����D(C�!���N�A�%��G����/r��	��Ƌ��C.i�����߮k�4��@�)������O��T\��v�ՃVt_�]7�ǯ��k���,���.��+�J�O?�H_<Q���{L������� "e_[$Jcy�`�c���/MW�������Bo��c�1���ǃ��N�#�� �$%��<[b��J�D�!��%���ɘb@��C	���G@���l�&j�EE|�5�����Z�a�%������Ȭ�/yˍQ �kQ�4�j�z`����xo/�k��а�|آ����{
)��,a�xi��u\�5<�*�����[�%s�-G�JVY��$�|���Q,��z�����P��b����a.:�d.Ո��,�a3|%�����\}l�=�LQ�(z���S�~b�l#Uѵǥ� ���&ڢ4���$e0�i�r��2�H+��X�>�B��U>la��B�NF R˷{��(�/|bE0��Ѭ
��7�����4�m2Hƙv ���^��dRܞ�rT�OE#�;�D�{�f�=w�8��|h �x���n�<��Y������?`��V�+	1���k[� 8��	t@M˧�HB��z���rV�g5�������V��iZ��-M����h�h�p-/_�o�R���}_�^:�BSښ���o��� `D�ǘ�x"˪r���X�}hJ�å7�؇��Μ�Q�%�v� ����ӿ/Q�����ѲkuJ��B�V��Ir:I(`[�鈨�P�<���Y�����Qt��K��^3c���Шu�0)�@}�Y��S\rv�<��|,n!&�W�
�H�u'�^��s�>�L�@ʮ���e�E���z�I��'Ƀ��vu��Xa�.��L���1�R)�9X�9\�T�C �C-��@,�	�'z���y���j��]k�P��b�Z�*h����L��Uvi���`���/�<��6ۜ���Gto��&�dK��=�W��^9�(���f)b�C#���!�9/F��%��&]�w3�~�X��k�qPc�N]n�
�
E�$u�K������J��xA~�_7Y���0�����V�.�=3��JC�k,�'�6�\Pt�;��#C`�b?C	�Xܖ�2�+��&���Mz�X
=�����N�by�r��(����]����$i+���\梑J�+rW��\���<Sԩ��}`���D!����j��N��c+'��ta�g]�	YǏ��	_�l-[�~�2�n��Ѝ�v�a ���������ޞ�2كq̑�ek8fA��;�*�r��3���l6tX3g� ͢
�D�0�\*w]d7(�M����$p���¿��F�t�$� 
U�P�;:q��� ޕ}��W]��
��u��U�p�,�'
:����4�buy��;�o�	4j�ȵ->1�J����\��4n���w>l+���52HC\��*J֨�����i밝p�T����5�����郱J�z��<d�0��krF��롢p��r�l3��&s5��m��ayk��ҧ|���3o2- �Ҏ��SO�%���?��4:���Ds�sa\�B{⎷ �,�X%�m@W��ɵ3�	��~
��W�Pu���������'�r��j�1}^�̱j�`�ύ��Z�+�2�~��A�E����l&&�W��ʩ�U�pXx^�k�^ ��A������Ã�pY�㷡/"������{��e��/���s)��vZc�%��Tg�ғ��Ą�"��Tq���HPD�*�A �R��3�%��f���nZ�~fI��1o������>�>X�&��<��1wS�����Kl$gAkw�7O�h��x>��@�&�k�c�]��n��N�[ᆵ�:2�4r�l�#ټd0"���ޙ�I>�@
��ҹ����Qa�����םPh|7(�b�UI��B��r`6]�ᄄv*u)S����F|���-�������ks'e���$�N�*��iGxr1)�؛{E�������,��Vq�V#�x�AJA3"�=q��d�v���=��s�7]r_OQ�2���l���bN=�+IX_�G�6yn�<<����?�,P`�ֵV�<���X��O��͛�9>�(ݷc5�;OPמA΃��=J[�*VE B��~v�L ����Ecu��s=N'�Zg�!_��b�<6�.�"����I�.HI�f:��)�(��ع�	�T���c��b�]�B��a�b���ٺ��4�evz}	��g&r'��x�[��2��ܩ����9 40�8Ѕ=<��'���+έ����Ի	�1���۰��8I[o�腭eoHL�9����M�д/)~�S,CJrakj�Q����z-�(�҃u��I3U�J喡��\��9�;���/��?�ž��U ��UI5J%�	Hh��l7�7���ā��ި��yqVJ�'� ���f��ybf��(fǴ��q@!�Ξ�{� ��@�Qoj��Ʀ�ΉǃNh��C���2����Q��>��`�.'��v;X-�c%� �'(�p�G���z�[��,���0搝!�9ӶK�,]��hP+g��ٽsJ��ɜ|}�J d���Z)U�9ԪT�*e�6���Q�5VN�������[��GA���g�B�IQgև�i�y�*�߅ź��|be3�
���~�na�6�AnY�(���U�qwF8�P�k͑�^�ڦ�?�l2��f�S1�5n�"AI�\�e�����������'� ~�Ѩ|tî��Д����[���y���QΗ�X�'���A��6O�	쭔����4\��/m�z`���`˭oBr[��`~�?4��c���u��x�w|��&uM����}ֲL��Nݙ7�*lzk`�yˠ�E�X�E|�y��m�m,��<G���Eg�`��un�ҹ��>�j����������u�ˑ��B!�%Q���U#�;� �|ѹV�}��E{��a�#�V/�3Y�]�q����Dt��>'9�N2��9�u9[?�+��\�dW,YS���ʸ�&h��zz:s�Ц�׭��o*�.��ׇ�#\��H�*Q����I+"3��'l�P�]0��y�����dy/�%UC��&!EٳI�	�TN����p!����Wh���y܋W�ʧO�A����~��T�Q����z���F$���Ra��߄����M����7K��}j�<]��~��u�
L`�zR8o=6_ �Ht�'��c4���%K�Nnc����_�����=�,�H�MR5U<�Ph<i��#b�p���*��^�٣g�@�,�qm�M���{�5�󹾩Ӓ�<1ª��� O�z��c�X�>i�Bon��ů҆���I�O������lꦄn��;��3׎��c9r�F�`[0��:z�G��$,!I�=-�NM)9��^��8�N�G�7��t�{�6kL(�尤��)z�����:��y5ߒ����,[;�N?k��H���� D��
�I�c�Le9��b�S���P9�q<�޵K��x�]09��3�*�����Ї+�W�/��x^�DJ��K��SZd������4�O�S`�r����9����{�H����Ӽ��7!+l��E+IJ ˟$7��D0��%�}xy�7'���V�#> �Ƿ�t���RK���_�#(l&����Gj��n��Ƴ���~0�mcr�D� ����1Kl�C�Cz!]��*�s^� &v�Қ* $^�M����4mB�~LB:kluž5&o�!�^w�J"a���<�����\sd>x��ʴm:���5�(�kX��I(�00���a�o������#�
`��}a�<c�a��/~z��І ���K/�uG5V[{~��w�IP9�plz)�����V]�wž"g�O��y����y/�Ab���(�o�Y�ox�@�p����3�?zS���Q$�.���Z�1;���Q6Z�Ĥ��!��=���835����ZWz_���:8�q\׭D/�n��_���������ޕ)� Z���,TA̿/p�hoc��"��Y�ӟ���S�Բ��KKᱍ�S��Y/Bi���\��Uw����c�@7.�A�W򹘦�
MX)冑�z��1D��I�-v��'tr�Q��A~'��G�8� M�nHu`]���%��-��K�� 1��	�}� �I��tN�:o�0\{��<\�����?=Z��Q��P 0��gs�V25 �� �]��rP�;ݿ�� 
�mʈ���Z�R q��_���0�*O*G����9�B��n�ɕ���
��|�#b~9�N�kJ�Vv�V�h�t���Y��ȵ4�a����[Y�,�\��Z��9&渴S��O�s��O�د�m���ȏ�5�g�!���w|���_���-q�L)��c�3�e��d咄SK�I@G^�ա�G*'���ϣ�؏p��x?���cS��m�ʨ�������n�<��r��������Z!���-0��Z�-�R{)Rן�=yx)Fwy��c
�l�p���
�G�E��(�Fg��]�ͩ����!7��l�r��oc�X0	��/0�iߒ��&Dx޷�1��*��߸���,s�ġ���	:�k�Q�FQ�1�+�#)(X�D�F�R�s��).ҟlH<Z�佹�7��\{�7
�-i@�1�T�� 3��+�q<e������▣��)9����p����G�h�j�t�5_�0C��~d�?FQ��T�F��+��n�S�}��ܨ 6���Ҩ���t�:�=iљV�X����{'���I�rS��w�	��Ǣ�_n8�+�\�㥎S��SSH��*ڸ1Hfi ����R�#d������|�x�S`
ϘEӧ�o��<���x�+�EH�d���"��j��ɇl��4��>gz���#ߍ�<Ec��3#���Ƌ��ϣ�V�:�Ҫr�}��KP>��-�Z��7�C糅������뺋\�/��FPwlD���(��'~���|�89,�Ϙ��Z�Ճ����v�(��L��*c��^d���P��}��@�}�ī�;%� s-4�O9@b-^>'������M"����GB���O��pϒL�Ю��������$�9(�3�
!sw�J$-1-��#�~�Pݠ�שn�ȕ�D�wI����գ��(X%e�6�q�b���k�ݛ�s��[�{v����Wq��'�x@:�;�Sl��--�Ub���<j����费'�ܖ}w�F�QU��X��ޡ�v������K����[͎{� �����wQ�P�Q7���ރ�Cr<��.�����;Cm��
P�;]?�,�\󮃋���Cj�tM^�d��bC"�M3�@�w���nϨb���l�ƒ�F	r<	�����D�
h Gat�7}��/vT���*W5��WJ?r�v`��I��r�C�fdcl鯡6�I_*�>٢�S����������d�i2�O
U�J:�l��$hǂ�[:�}���__�0��К�+� ��;۠�+��5C�H�M��:I��;I����;��|'���ɗ�P=�D�@ڿ�B�u����Ȏ$�z�W���XUL�?�G��I�Z������-��'C�Xm	���3��@禀km��NG(n�!���}�����#��4	�q�T6<�]�9	$@��8�D���a���lu�v�)�E�֏����0/�E({�+%�����Fx��O�9\e,���z$���d��UYEn�h)9���	x��X�4��c����1D�%��Ή�-)Z	�w�m)�B��}(�0'�"Zh ��8�x�I����y�ơ�#��T���b�(�O�smd���G���� ��^�jxhԟ
ط���,��aMF?��[᜕����}���VK��0��,�!��:��;%Zc���&�DT�f��jh�L���\|�n�_w����ʖ�3:/?��y�����#���GW_a���*?%��@M����N�����&*��٬֍ ZӮ��5�m���.AriB��Oz���L�|��ƌl��f���΁�c\�֎h6��r�3z�N$tѭ�y�|����q�?���$�}eá_u��ͯN�)�O٫��z��1Sr@�h�R�r�y�ˋ捂Z <�/�ͫ����QX��:P ���K�w(r��g��x㊖�yA�Z2���"HL>�'}瘣��^RZ�V$��؉��/ʦ2�i��3�Kt`+'3�S�ד��$�� r��� �b�Sۏ�#Sv��b�ː��)4�C����~�49�)�# �H#�mmc����M\��#p�3^	q$�B�"OHYWiy��IugAs�;DO�FBpn��+Oі��Ak��xV�!����!Z �N�`��|oP>JR�e-��~ݡP�ú։��Pͦ�?��971#*�ZM>���z��/E~����]�+vo-�{ ��O�)d��x��F$h4LA���k�6��@6��/�z�H����-�5��c�U\**1��$ܒn&�r�4<�eK��bkm��%\��[���԰*D��u���m��/ӝ��N"���04h1�^�����LH��+��i���-L�%K����~�h}�J%$^�!Z{h��;=�������������|�Su?2��^j��;B��)�z�k��.��X�B�A������x��a��|]�U�be�`A���)��^D#�_w�1��M(*�O����o޺s&���l3�UU[�!/�Eȷ}1�W)�O)\�wć<��5���f��zw16���7�	_��!vrܰ�IÒbV�<��v���'y��&D�K-I�ې	���G�����:x	�ޕ_@ni8{������B:�(�0����Yz����Mi����=����:P,��^�����Y0��|r#�3��ָhg��G�#���U{{���ͯ�Z�X|H޻`��g��	"��\�I='�0]�4CA�� 2�����?3��|����)�E��\�s���.�74��G���{#Q��};o
����;�u��q��AVh� S54���ޏ����ٯ]�8C�N�9�U�)��x��n>95FU�i
j;��7�㌏�O��J�
��YZ����0�im���XbT�||��G�ڧ�.��v�}p�Y<N�d/��jljw�a��s��%�-��N)�ޭ�����4�8ux	�)c������C�}�9{�3�x;����i	�+�Ă���R*��[0P��7���_)c%Z��p �Z	��k�نCG�M�~kY��a�>-j�\�Տ[��N��p7�T�����(��m[Ǖ�^d�������܁�rkN��'#<��XmE��^1���:����Hl�-
��-ex+�̞ա0U4Hynmj������╉åi$,�1�B��R�i\䓑k�G_c�r2#�j�Oz�Ĩ�HZ�;lJDI�v�f�0�#U��2��ŝ�	��iڇ�'����\F�!;�BA�6�׎Ϝ>Q�'��ȻW���Y2��b��,�o ���w(e���~�C£��֠�����+.�k��}|6�&R���k�sQ݊*�0�mmFN�N����Z�j�1�|�i���14$�W�v��َ�77NR>ЧMz-�؞�b0Dԣe0
%�kp%��JK�zaW�?&�qMI�0�'��,�R])i����'9�������m����	��n�Av�Y��?����>=�f�1E�Dُ�ۡ���D���r]�D����g�R�^�������� ������QQZZ���͝�J�I��I�6��u����/��ө
c�ܟ�z��Ρ{R��+��,:	Dh�	�6�Q	"ޫ��T��c% b���O��U��Í��FHlR��3םJ����w��Y����e.�Fi +0~�m����]+�7�G�ۛ?]G�E�:��=vG�=k<߀�8�ivnU�v�r�=3�Nێ����¬����O�s��8d3���OjyP�7�Ianǒ-��u�d q�l��F ±U	��鬉��W��J����r�o�^9�Oy����Қ�$�Q�3wC�L�'�@��Q]�5u�[�����F'�� 4<0�W�'jr}:0#Z�P�))���������x��G1JG��̢��(6�_��)��9���$rj�:�~Mk�>����Jƪg���,A[޵�.^-�,���lKX��U�cْ�����YW{(�l����*��M�s���䲏kXk�{
Z��LǇ�&�fP�F�V+��lN�֕ �V�+�
m��3yw�T�V	V�m-m�B�d���W��t86�S=�+t�Z�4w�$Sk��OL��ٍ`�(ĉ�`ʠ&�G׏ލ̓9�'8��(��&�"���6s��~��>���G���m��w���E��b
fx����I0蜬�ŝ,�WxS���	���V�i��J��	i��V{�ob��k�~=P#�ƻ�V�5��{����64y,�ڏa����=�dE�[�_=|��<�#)��Y�)퍶�\7aQ��0�܂���Oǀ�B����t��ѩ�3zkz��f��z�v��N��W�^�4���½�#I� V�A��\p%�h'x[�{O�}����^*h��.A�I��p}Ò��8Dg��d��k���y�,>Z<]�3��;�oa%�2�&�Oᖢ#�[4��\���i�i�koE���2��:�J��E����Y(5����[Qy�a=�m��-��/0Pg�T���g���5Ȉw,�S��v���>������,�ō*{��FSuߗ�����q����S��iA5��M�阽��G }I\�E����A
��Q�9��$���n�[��.��=�y��6�s�_���XE�ᓉ{d�� Q  �E'��>�m�����2:`�"�ۉ!�G� �ot������M�J�X厥�f�Q3�)uZ�x��s��hW�m3w�L1".܇�5���
��Ճ|�8��ݻo�C���[u��T��$c�!k���
rЅ�t����4U��ȃ$��xd�Gȷ�@���/�< ?	F� ����D�+�<�ͺj#,�aѪYƗ��lTy��U�)���?��Y��	H�Z�ն�����^�qhA�4���N��\���~QO]sՍJ�,���e#�iD U��<m�3��Z%�� d7���mf^�g[�V�c��L��g�
�x�7>����:v���{�j��a��]�h.8�a�s�����wi�>R/�_P���G�`|M"$au��$Z.4}!�su�ڍe�C��]}3��IRIe8������U�3nѾ�H	;��q�<)��SܛW��׶��e��@-*jm�V�Qz� �*�� ���6@����둗PCD��9R���H�D��1�s���HvH��� x�D� �ZZB�ǂ�Z��.v�E���{�"�B�4��1�'��t!�)�^HNx[���j�8�l�]t[3��g1^�0�~�i��!>jg��S�� �Fz쑞N?�Lf=���2̅��_�>S���K�	��1��+�^k��j(����vH}��x�C�5K�Ȁ����(��5�!Pz�X��ͨ���gU^F�+m��&��5jC[L�Xc��&e C�+��#]����S�Z�p��>O4�5���U���^c�t��Ђ>�x.��� /�0�,�r[��l���T�U�������R���3��;�E'�[��A��c�
�����03P"7נdQa�%xV"�9ùhT��Ȣ�������t�1�ӫ8v���w06�y�21�S�$����7>,]��#�V�.���n��f���b$�T 핓����Xo�Fzr�|� �\�	u��_�Wb���oU-��D���~��B���$�?./�l�Gs�}t�H���_Y��v�ݴ�ݟ�91y�C��03\|R~�v�:�z��l%�_��~�g|��`c1׬7).��S��sĭ��0@@��e����6C4�C�j��G��[��T=w���١E�C���������t7�:TG~y~Z!��+��T�"M�]��R�wP�Ej��X����:�������1����*
#+w���&l�i	x���T���ݯ;���b�lH8����,gv���*g�+�ŭ�_~ܒû1֬�rxo�K�S\3���6b��xXE�xA!�%�{�Xl��=��ƒ7��!,F$+o��En����ی`'�����Ǧ܉K1I>_6���4�Y���FE[�4iX�"X������{.ı�7�dO�ҙW�/��~�^H'4���2G�?���,ĐV�!�y�,�0�;+E9�҂2'����d��+�����3��Ny!){��|(��4u܅���y�����c�`}�����G�]X���:V�xdW��ű�a�ԃ���>����$-�m~͐��ޏ��*������
%us�X��6�bZ�gW7�>�s��ə�@���v���3>��-}j��` �v�G�+�)�?����Vj,�C�?^8\��u��Vw��v��г�j���~��6Cb���"�z�iM���v��x�0���\+�L��݅�䉇�w�r ͩ��N��3��C��.�QF�E�Pس�8��?��c�,U����l�h��U\�{����Q��L݀vP��m�)� ��9�#�?�Ug��B{z �����P�ze��w��HG�{�v�ha�M�`D$�'���F������G��sb9�<dDE�u,A��+6��<7�
���c{3(B�1�ai�KpIҐ���,�����%%�|��i>���1�o�F�P`�2�F����5�Q��lbdƈ0J1�Yր@0b�]�=���M�q2�L`���6�;V�p�[�m��'ʕEI3��nr���H˦�%��J-��y��s�r�E$�ASȥ��i
c�t���U�wDi�r���$��j�x�O�Tڳ^�>nrL)C��q]=���dj[���������}�x��P'?��� �E��l�
{{B+�-%�b�$BN�--����a?������k�� `U��t3�/���EC�ڪPC@�C�{�$R�/@H���i/�b6��c��Ȧm�y�8�c�y�*�_W77������S��θ8~iG1I�ƺZ�&|��$����؈�͂�;�=#ϐ����=Um4���aʪA	ޘ�pT0�f9b�����x�Z��<���G�e$v�;#s˚���@���g
+V⦭���*���ܤ���Kc�FY�h!�9@��@u]N���di�U_m�Q+��Cfc`;���x�%{8�G/�l'���[���8�����7�?��6�8�K�w��ܚ�׸9s��+E	}s��#�f[n�R���HI��3g7��sy�ɧN���Lz��kr���.N ��
R����c��z�QWw�s������FI�v�ZSw��ع�\8���Y�b!�a��k���0)U\��� ϖ��!�S�pN-�֔uV����P�XJ�MFmc���������(�i�v������N)�h�bR\E��(e���Z�Fe��ף1����tj��=��l�U*ш��/�'z��ɻ��mC.�8����EQ�T7$K��.�p���Hs�tc��T%��+i�i�� I�C��Z��2ē��B�O�<��`[w_�
kQ9�Hfȼwګ��-�#hQ?ǹ�t��9�oU���բ����OZ�H���K�PNc{�/£q!����J�;/�������7�%�?����hz���\΂~��E`���~
�O��ӗ/70��j}�w�h)g���܏ɘ}�{��r�O�u ʥ�e�=6B�t8�(m��/ֽ4&ߚ[=QA�Syi4���y�V�+�_�^�2�dAoӛ�OՒkT���9}��Yo�\���*nW��ަ�<c3��[��N��Kq|�S!���#>"�Px�fW�+��-���(���]P��g��T�m!��Aj�s9|�>�IHe��8��!��:(��f��lU�M�TI�Q��������ٌ���	J�삱�E��Ei��6��A�Q��߅��ы��6�nJqd셤���k�qP�`�!�X&�ޱ?k;d2���
�&ʦ�V�FD-~Z����m�iSMq��d_���1l�W-Y^��ƘPy�en���;��ν���4�q�(�{�F��	�����v��@��^k��>l?�����"����0�D̙�:�гv��ls��Zĳz0�-��$}�e����T�c�� �g�_�XO_n틺���"R�;��\�>v�;�@9A;�#�xQ����ؕ����6ϑ���N���!r�+��W�qo��c��h9W�[V�:��Ki�E��;t�����RL���v�cC-5&S�:udt�L}�5�M¯b�A������؆X)  ����.��K]�\y�^�GCh�Ȧ�&x?��>�<@�5�B�M�$�X�zZ:e�m�Έ5�iT֗���
$��L�j��S�W�$�� �ww�b9:�*�"L#OA��`��,S�P��Y/l�	U6��#�/�r�H�5��\�_n �"�*�#wp�_�Z:���� XF�����2�+�Z���j�b9��B�X��\B�V�06#��.���ak,��),N��;?�/�7���R��W+"Q�N����·�V=�k�P�c�'�JJD�o��B�?MTBHq͢�w)n���w4P����s��X�oe�����s%É}�m,�\��^~͖�������V79����,'�1ahC��j����Eg��3�l�¯�$�pH���w�l���"��g�C�B2���m���j7���{�R>1�5��(��3��*E�-�2�*;k�hb.��.;^t���3�C�rؔ�q���0��A�ϴBb��r51kP��}ᵊ�������kƆ��Q�^�!^Bt�����lr_�1?O���i�!������j糵�p)�#1Ǧ������`�X�A�p��CߴB�aSI7����	��\U�ܗ�m7�#�2�D��˽��3{��d����ڇ��L�ؠ�NҪ�g!�����s$��E�6�d�@�
�O+5��+	��ȉ����H�\�ޕ������B���dz�����|��R���|%�~ϤX�a��m̃m�k��V~2�S�ղ����W��"�}$��ѨOѐ,@tf9�7�2�w@\E��o;V #ȼ��pY!�b����T�~����09d�t �څ���(qk��T�c\�N��:�;Joɴ�]H��i������g ��X�6�ړ��7bׅ���s~��C��X�<�0�
;S�B��ՁPǈ_�	Em�9�̅sk��f����K�Bb�C@N-��g��( ��I[�w!{�!��hnhg�*�^}K�9Ռ4F&�ߜ)�/�z��\�+�����%��HS�z��B�L���?�Nu��/*sD0��U��Nl>�ǳ��i������/�O�s]Ѩ�V�f��~,�&|2[kK�t�o��� �?�ȇ��=us�Z4k|],��hT!h]X'�LJ-�����.���/5z]N�R���^��]|�1[�y��W��
�_���W��*�Xz�:��b���g�]&�p���uQܷ�h1AB���R��v*�~0>�^�����7@'d�f��H	Ed�Q%�$>�Qa��U%�����Z��Ĝ�$B}���g�j]��,e�)�߳.�k���k��m<�Oh�3C���ǟ$P��k�hp�\����Ȝ6D&�;g]�Y��}�k����"�|Q_����{�/[?��b���	XHcX
�V����N��N�y7�Ռ"tv\wA�nX׍i � �<NKdR���Vj�������O�/��т��ʵ�9W� ��w�dr��箓W5%��F��[.XD��j�yU������z�3q��Z�c�\ݗb�������Zt�9������5$��jJS�_b˓������(Ԏ������iQKD*�R�߅�u�F�]/��s�[��
l��f;�� �7�f�]��	�<z��ITG�:����.��UQ2SC��_��]љ��Ɗ�ȉ�7E��S ��~���i݌e>��?�շ�&!�$T&}�� �pohV�Lkᝋ�C@Da����ՃE1_o���@��5&� �_w�07����o�;��;ly{w�l"�^��'�hx��j�ST�j-��$��ڈM �(��){���jMY�lB�A�� �
�Q
Ӛ��$R�`1��.t�_t>ޫ�ˍq*����Tg�mr�����c�>�1 )��6J)��b��E�۟��+�_g5����Ɲ�ـ���=���I�S�z���`%Q.j� ��)s: �t�b@O��݃�+�5�{	��P?K a)#ţ~:�;õ!��?WQ��4x��~��H8�5������1�)��\�`6�_�ߟ�3��kYL`��u\���u�=��*�N�y�|+�h#*��@�x�-W��Wj��lM�[���-7�>����o�%�.�&����_�'\֢��j*�{��W�g��
�D ��C��5�/6����z*67),}�ۣ7y�x��@�'e�^�@�TuY�z�Ӡs�i���DT��Å�+f<5�������A�L2���࿅cJߕ=Q�.��9�S�~M��R�?]WfY���w�u`n@�o�T�w7J����JVԅ�
��*�P�,a@�wb��X��}/��]t�a
8�@�+��@m�^b��	D̴���+<ڠ�Qh��5���4�[5A��i]x"
� �@`���4�f���Z�޾��?y�N�0�?���$xL:K;RKJ��c��Y�+a�� Ix���"O���SP���n��1���_�5w�ӲC޼��͖��Tj������K(ͻ�#��<��	
�T��Z��.W�<ܖ�=ɇ�9�R�tՙJ!5.ZU��4�
�.Z�5`��]e�W�ꊑ��#"7:��e.\���5�7Oh0]��ٰ�G���͍���%�+T+���s�����bp�ݜ������nJ
E콂VJ���I}�OJ ��#�ۃ�'��O�7�6ȩ�h
(�8S' �}��8@ގ�5�{m`7�zyi��'�����52�X��߿)y�d�)��1$Q�H��U� P�wz@�Z*RA�M	��)[fP�;M���Hn~ɕ��4"��%�L�V[86˨x ž;
:`T�9���˓��Cʛ.7Gv\sb�HH�3����><;4�+���i�"h���4^���jk�#ψ??1�!Q�V�����1��J��@��=���^vlː��!�'��Kc#�<�8昁�!����PԎ��|�!�@Ȥ1�b
������|\�#�ѹ��r�L�G"y�������������:���s�{o�jm?�kڮ)����f��^���T͢��J�B�db�{{���2�\`��� �굖/Mq\aI�m�%�=_�'ݿ�@��c���H��Q)\�m>�� xg��MmG��M�0~�rw���6�u��n���K9K\�;�S���s=�G��d9u;�àK��h-G)��#�׋�R%�˾z�G)o��<�"P8Ci�%��i����%C�B�&��o�A�^�ۄ]�Z���ecO�Ql��`v�G��m����b���V>�Eb�cog��=9,�:C�)�U�Ak�̢�n_E4�b�8Z�N��ܧ�唑��$�mV6�WE��e����Bs����{�c��l/2�F�g�݀��rm�g�ߜB�(���*�t���d�ٔ�3�*\�.�y;ۥu?���n�m'����i/�:�t���}�	�n�Y�6Fy���A����H�Ƽ{�Q��m5T4��gd,�:@V�3��?�2��<��ƺ�i�$����h�r�g�^D�+tKoq�t���B\�ߒ���P۾;?^B��[5h�xc1]���6��s�g�����(�*��\��?$��߬��M�T{W#:R��W1�/��4.,���a��C0%9Ә4�7v����e]��p-�|�lX�τ6e�̸������K{�=i:/�Cxʉ~Xn�
U� ��Cd -E��
��X�E�5D�� a��C )��o�_y��y��q�\p��GVL�c6�" �;9K��!��=�(��L�Vg5�v�M�E��� o�(5��w�TE�;dN� �;zxo��w%)���X
�?�	���^b�J�Z��s�:'�A�01�\�
$�H��U�
w6��0���'�0̮�(�1��0�����r
�m��̄��t0�|�������$�!��iR�Q�K��ԡ� (�kM�X�}� ��x����~{"Z�?Q���`��J͞��5�����|~�DZ�<�ɴ8�vi��k�S��9�ݴY� �RDd��������6B2�����!��$�Q�YP6��i����{��td�,�Ͽ�W^l�s��4>Sb�w�.�<��ݽƳ}����EX�!O#��������5���֌BѵĊݯΨ+�����k��������� #�fj�TuXٞ�9�g��F�ǻ�a>w�ߌ�0�0���D��>����k��	�2T  |��7n`%!
o_D���5Jl~W�W��«��
�F�̦��6Ke���5sV#ZO^G����,kByk�h�ރ�v����.�l��� ��/�ݺ|s�*�T���;;�m?-�4+F'��kzL,&JȒ'|mGB������<j���l=����{�y���lm�ժ�$�x��n��V8������i@Ÿ +5!��oc*��A�V���+��t~^�YзC���<���jr�ivX��,��b�y�&�I+���ޖ�����×n?h��d�F�o0}멏_vХl�0>#����?zZ#�O˄0e��a�B��  ��n�WVnd"^�<���)�ɭ�HfG��~`��ʽOJ�m���'WNi>;L`��#�Fh�2�kD`
QR1��_n�v�k?^�� ��v>J��3	\$�s*��Z`�<��f���Cu�t42!w��.ǌ��zP�W�J

�%!�����i�6�5��){e�=�4��!����q���ct��M�H;��T�4 vA�h���cq^z�]�:Ƕ���b(��n����KohK���-�E��Z����{�F����8�����ـW[t}W��9���gv���<���B�9�,��Ɔ�&p�`��iT�]����㑺_m!�쉴7ZibG6�&r���C�П�B�J(]�(��,�F�s��LDZ`�l���R	g��脝O��Y�^�uW1�u��a�Cf|_6y%Ѐ�EI�&d�&�&���1I1�@@6r�������z��9�-�2�I�8�h����� A���,	��=lh��J������3a�6��A���r&f_��Rj�d͝}C��M���-ߺ�k��=ok�����'�hcy��An��g
��� N��q�1�v��Nؠ6�+�co`wI���yІ�l�]����Rr<��G��S��?S���O�ݛ���5v�+B��^4�L�iE7��I�հ`@>�q�n�(���\�#�l���;H6��\���d������|�=�	>`���0�4|�?�V9P�ތ�J(���m4��S�M>C����m�	��\=��kve�xʧJ�cY��9�Fh�L�ӈ���A��ْ���?��X5dk��RW�	�����w�f���'�Y�uD�!�򙗰�oM��*��|1=+�{!��O�V�v��2*�*$w���|Odv��GТ���c�!@HhC`�0#hI��wf�d��K� �<�c����?��I�Y���n�۟��C]v��:_��.�T%]���wfj�~zXw�/ YI�_�)���������Q���S�߈3Ny��x!���|�����2iC�d�svh�>pL#rk�5��H���3�Y��#]b𳮏ʯ8	sk��;��9Φ��z��z�C#%U�[P�4�,,���+/)W�9��x�K�����2~J>u'N��w(���"̈�Wu��k&I*9��Ճ�Y���vf�e=&�Qy_�1�HO�Zԧ��i}X,ST'����އ�W�)�K>��n�Ř\Sb�QA�/��2�~+m��H��70��8�C��d�ا��A��x� 1�댇WO4O��(`ycF��X���_��|��D�P�
���K��������!� �*Q�9=��O�@�5mu�箪p퀄��D�P&����+!�F�հ+g!&,�;���B��T
�Fdu	�ds#ᅝ*}h��w�����ʄ!~�_��2�����]��<��{���t�-�D�؈�k��,�Y4��FeH@�t�����Da������L��'�C�� ��N��B2I�/����{��av���.�vɸ�#��rgwO��iHf��mڞš@�O�oڸ-�炌m;!Jza-�ř
Kf���ؚӤ� 1����� e9'����"V����"<;h���}�iFxI��ф��U�G�L�o���қa���Y�_�ȶ�³`f��rg=���S�"<�nZ˄�U�B�\�$G?A1;9�3I=��ن�{%=��b��9��&��1S�����E����xw�	�_�!ג��=�}�bo�k j8Ť2�Qg���� �\�FB�}v$7����d����֔�3S�N�}��R���� ��_[�F�6�D�^y�V���{$s�6Qw�J�n0�e�37���vX�S����.R-����f�B*��*��v�d�UR� !�H�w2Թ��Ĺ���n���Ѓ���Z�#B5"�9.�!o��?��Q��}B)?L�R��@FQ����w33 ��������7h��oqIc�n�]��/ų���d{���gE�j� .�*�S���	��5$���gOC~�"	��5��.ʪb5�	C���$�8QU@J�̒C%L�־T�TM9�p�Y���W/�:�mZ7	�p"c�������<L�p����L���P�P���m�//u�@���؀�y��3 d�V���ܘ�෭�tԠ�Q�2g��ơo0�1"^��;�;h�s�@̉��q���T>��a4Xk���8�F�^1/=����y�Pi���x#I��F�u?�K�4�Z�Wj3�'U2�A��B9)Xo{�j)��R�W�yE�����y�r�sW�q�@��_�E3�A��s��G.R3�3&��������z߃�J+�m!6�n]ڇ���[��
�Z��Ha �ڞb������Ư��{]�<	�ڬ�~]KY��t�kBE�kY��Α�SL����f�hkq�;�v��y Pq��OU׮�;�S﬇D@U&)�����N8N�	@��K�]+�Q�]�POx0���K1���j�S����������)4�>WH�{���;�b����h��Q��J��&g܀Q�_S4G͵�lD��C�[�������ݴ7`��j�:��	��8u��M|�ݢ��I��:sl��o�cuߦY���Sv�+}�j ��%����`+��Ȑ�[uC��B��e	`����1�ҫ�F[��%�UA�����$�"(9���Q���uuܧK�ު�J��#`,WP6�,MT�7zh*�s߸OV��'��m1ML`Kr{"0C�i���h5ͺ�H�cڛG��:�d�a~jf\�{��bM&�.��)���¹b�d0�[�QLi�Jd�x��S��?�j����]������~���d�n���&�D���E�cҭ���xό,-�=M�s�6�AHOJ�J#C�ڢ��cC/ B��LШ��ړ��"�5x
��Y����M��������w"`��B�e�1v2�^ސ�3�VER�<��T=�E̦�]�]��b�ߖrm2�&���C�Q������=j�(���<v}(,�o{�Ss�:�o)2����e5���Iw�a ���u�^/!(#G?U�a��sN��PT�� ��k����8�}��\^k�J*Ѷ�ԟ��Dv�����q`G�,�5�D/�ʵ]�t|�����ԯߋ"�,��:�j�7	����z?D�l��uF�y�{Q�f����iP�R|$��]�pj*�U��|5l�{�1��y����.L��n?1��r�)v�ܿ�kAc37����|��L�+�]6o޿",��q�r���� Q���b��b��F��o���Bl�/D��'pprK,�D���NF�5�3|��N|
��`��^3V@\a'�l�+�������n��\#����ތ	��/"2��Zt><�Ov�;K�/SՎRR���"��9�F#~3c"�]��a9��y�[{���W�	��f�CL~r邽8�ɹ��<I8�o�cC�e$·:-a���	Co���������
�<h6u���fkȃ�_���7L��v�\�J]�-���+�:[o'�+��(?�5�}D�cȂV>O
I���j�.5a����U�ț�<�D|S�≆3T�� �`�(���<���{���A)��:@@5��! W�+�{Y�G�N}���e�9W�W�y�-W� �X��1=����;�ͲD' q�d-���X��_�ƚ�Q2�e�H��5����| �ߟ�I}t�s�O~	�av�䰭�"�q��'^U�q*�:dc�hA|(GU��@�{7	����s|1<*���=X֑QPp����[$ q\��ѵ� ������O8�+�Hh����(�
�ޣ�>��NC|���ǥ͊gNy ��Y�:����λ�Q����.K�&��5o"��A�\%]����p�MK��{v���U�(������������ M2ңH8I��6C�/�G\Ja�Gm�x	iYV�ay��G�@$姉b������(ٍ�f`�+,���k�J�v@�ۥ��X�Ʉ`	��
5����&Xo�y�����P��'394���M�Re��́��XP��N����وv9MB��L�d�~��^�aѺ�`�o@Rm�����c��:�xnػ�$#�*���s��(ʠh�XN��׃���;�vq���eh���Hw(K~aW����^����X��fr�/��I3FQ<BH0�a�p+oF-{���r1P�U��P�K��(Fˮ���PkӎS��VP�KW��k�
�+dCJA]�$��U8;��M�[�����qwj_��u%��Ɖ�f��x'�R���^X��q�k������G�X�ܝ���67*��v51�i+���6Ey'�T�e�t75X�+� O���I���5'�$G�q�_wf��E�Vn>��]����x��jF�t}�'&\�]Sp��gw��t�&��f��!�?�y���vn�	���gB�%GꡝJ��N�e8��-) s�ɞ��PC�4��	�2���$N�E0 ���\�fx�a�����8����4�ݎA��n���Ԍ��S��� '�ʔn�xsC�3�E���[J!;+�G�;u�.ĵ��(B/K<�2��K�h��[�UM-<H���ۖ��'��"���ߒ����uT���V7��:��.�|*:�,U���	rNC�֏̕�>e�ogrbf�������~��Y��]�W�e�t��/#����8GVG�B:0��_>An޾�~����n�u�� }]d(I�����d��d}`�J��*^@͙4hkw�\��*dYU��&�mL ��Y�F�K�C�.���`���Iu�9h�Z�m3��H4���|�5K�Z:l�����unqI�
Ir��K����v������G1K��kP�vΡ�R���!5����L�����'�jn�!���v
��	*�;u����JT��#aU�i&�]U���_��T�N�=˸�s�D�R�$��ϔ�dw�#�0:7!��Rq �$]����nu6qo?���Z�ވ\�R�40ԅu�.�����a~��y���(c �ht�p���`��}S�U��#�D/)%�^�B�rmt{�&�vן*H,{OŢ�q13��N��["ϫ�h�a�r� ������,`����7F�����j�gw�>hINQq��a1�b�$�7����5Ϝ���օ�x7N5�����<0=�t頱,Ab.����4+���J�+���s��V�/־�n���&���mǾ� �gX |���Ȳ(�������m�m�tx�H5�?�ތL��^�5�1�����@�y�9oW$����Bf�+yOî��U˄�+V���F��[@u���f�R���v�'�P	��m!p�%�<1�O��j�=���!�1{��vJ �`��nm�<gn-�_ED̓<�_	�,wp��9 0S��*"��&�5�S�`_�7�B��DS��P�P����+�g�L3y���$�u����L[l���[K�|}���#�O�Wz�5rB{n9:���@>IU�3���u��y��{g��v&t�o��QEB��ݰ�+W�%%9b��Cnն�O���ۘ倨߿�!���	��%�����p�ACn�o�x�����c�&Xb02�8�&������k�����̿���KTS�&��ݤ�r{E�-��k��T�-��}pֻ��O��i�y��94l8�٘�c_���B����e ���T4^F|��Ѭ�q2�&�o�eIJ�l�dQg^� 4}v^�z���a�P��%�c��S����Bk���Pi�Z�����Np5荔���8�,�/�A%o2��^`���%�S`k�,
5������y# {n-�C������0X��K܈��MĮ�[zPu�+��
w��� 5ک&��+�W&cB>u^ -�`�!��bF9�lDku�/:�k�<�/���R��qs�P��<<�_�Ό١P=�
,�dn/�"���H�LU�|S2N�)3G��-Β�
��2_{��1�<)<p�$��rΛ+ןs���`���R�[VJ<�6��K�]�,u��d���f��s��	����­�;�"�)(����lۡlf�<��yYQ@�P��ܝ��VH��T�]J9i��b�ԇjxX��r�G:��$�P��A�]�`0b�U,���Σ'<�Q6��Fn)�Z;�/��4x�Z�-yd铐��ܐ�*������/��`��He�1�zvٵ������ �!U�7�M�4��ἡEX7�_7�Z\KK��bS�G���9G�Ӌ:�t4瘄�PEzu� E�y�Y�+�W� ��(`��z�Y�,($�Y��,쐝�c)��v�Mc4F{����O{	�I�uنmu;}�n"�NS�^Ъ�= �rsyTTgh���#�R�/�N\�����:�?2�(W>k_t�Y�I'��8��Ύq���J Y���y�ṂW���>�\�$K7�;9��X?ץ�ý*�Q��+�a�9��E�IJ3^yU��nk8ʗ���|$��_�����I*���tj�����s/S`ed[���~� 1�M��H��{�e.�][�=coz?$��l���&�]�!]�9���p��Ds���:�����n�9%�����و���&�~�Y��Yd�g�������k_-|̆cV�i���>�PӬ~Vv�U��o��<��7�	Ә������6J�R.���S���q���]B0D��`��هX��}
>+���篨��ƍ0zY�A5��B;�'o]آ���%�����K3���
EP
��1��JscW��N�+��l����h��y=c�_�����a��ز�1y~|�[d�N���h��Nl��>N����O�=q��.��0���&ĕO�Q��wy.Ek���PlZ��}�@�ƺ�A>)�ޏl�)��L'�Ҥ0�APiJ�p6��+�K�xUG))�l_��º��J97��(������8��y_/��N��P�(�:9=����
�ВɠcUu>{ݟ�/\J���Y���ٵ�F�o~bȃO�/�����v#���GHi�N�zg�8I#�) 6���ֲ�	�ׄE�k+Rot�kTc$~�����2�Θ�)��^ٜ��r�z%í��o��gI�Nd׭<4�|��5�7ٚ1J��S)�P�܋#�>���=�V<��v��?:�s���*�_rĩ}�<��5��*��P������Ċo{�ֶ޴��ߺ��ps}XUM���@�;�p+00@[P��q��ռ0��|T�"4@yP�Oܰ�!��k5|g��3�s��u��~�cO�$��{��&v:7���1���hd��('FZ�̪�. ����5����r�	q�mL�n � �`�4i�J6/F��h=#)�u!����[��;TҥP��(�?t$X${kǽa�K�o��,���Z4��W�T,����Q�p^�o�Ps�$�&tAxD�w>�~�k����gw����� ���=_�����vI$%�A�1D0�w*r��<_Р��-�]����T��Cj`�5)��(��FÏ�)�-\p"�}�]MDۯӘ���c�c��;�_ɝFg�C��f��ț�v�����O�w�7��1{+��n�O ������H18�m۹���	�jg5c��f/�|�
VN��I��3�����L!���W����%�U��H܈	'�����.JJ���Y����	zW��z�Ʊ�r��g�J8;�m''i�L��J0�]4F��j8�FI���x��Dfe 5z_���Z%qj���GL�?<�Q0&����1�����	m�rA1���{-�(�����ۄ��/:����+��)b�v�����s�4;����Ϛ��x�/�ssxvĺ��b��6f=�����)Dφ]b2�x�X�d����'�K��D;h�t1hA�}B[�^�=����ø�%���I��9����G0�s��
t���y%yO�v9�h���Y��FYQ7�馅1��� ��U%<
 Z�"4�)ǥ���Kׯ�4�]�7����cƐ�*ַ��������W��h3�Wr�\3\��2@�ZY���Sܓ.'۷���Aw�24�7cj����k���G��c���vCŶ��)]�[X�����\�
�9�:�s;��2�n�bT��.]�@���	��Ͱ�|�S���[%'|#�&c�t�dvlC�: "V�W}��6d��C
푪k�G��:�2��l�n���'���1�^Fw�_��3��{����C�Q��Kv��j���?bh��îs3x�Tb�Ra!�Ώ���;uЪ�k1��~A! ��h_d�)��+�|T{,�R�M"yY���E}��UP�8?�dZĈ���TZ���K��%r�L���S��YF��,$mTjJs��X�Z�N2�
���o��d6���s�b:}��c#e�n�hB�����X����&�D�"Ĳ�uB���)Ю�ʛ� �S�H,�	�)�&�Y�n�B��H�+�/|<h( �b�ⱜ��%w���8�'7|kt�j$�4��In����~��n=o��d��&O�I=;s"|Ҩ�6��h������a�<ag<�Ih�p���8��1��Ը<������8��O���Ӯ�P�v�����������נ���yB�F��]Ȭ��� �5�n���F����gh���k�r�yQ���J��@�cRL�Q��)�����Īt�u�F@uUYRnF��͸���x&i��$����		����e/�X"�]n�8��y| x�v�ǭ�e��Ց֯�̬��-Ă���],��)S�1�TB��˳��F��}eYK.PG�3|���a�`�%���e8� ž���_cz�-�d!�j�i~!�]�֤ow �i��;
�co|_���b��v�[;2�]SqJtӆ�sU����9�n&�"g�I�ԃ�zso>�1g�Z����m̯ŗL�l�Kq��K�-�#, ��P�f`Y�Ub�D��;�+:�tc���Ue�r���6>i��a_�
�a�P���{�%_� ��4�v,1���'��I	z0HJ'�DVe�}���U�ģ�;5�bx��q�Nؾ�FFJZ1�@��hŧ��^�����=�p��;!W�1��0B������g��d;B�N&��PT����H�1'��PDq��T���:ցe�'�¸����Ci���B�n�7����������' f���V��&� E�p�kj1eA-��{ޜ9M�1(zm>����-ɱ�@�s�+O���y��Y�|��]��e���w-r=��62�J�6���g������W��G&�aB��Eׅ��-2S͔5�k'��Ʃ���.�S��W���a}B����4zQ�'c��?�SKK%j2���k�`u�����.���jS0}ku�B�w�ljc�Fkt3�����%=Rx����oZt��%΃{�:�+�fYj�v�څ�8I%2��l �G� ����	Ax��D^���Qq �EnWE���0�&�IZ9]
e:l����~x����a�S��4�lWu��X08��!8��q�\@���"���ـ�GB��6����w=9ձ~���"�&�uK�<����#���r��C��q�1�V,#L�d�����������ݿ^����^��wm�Ȳ�G�h�l��Z�L6��f&�a��o��}���!�� ��i-Z;?c'�3�!�c���+PTx���������6����qL�%6W�e>�ԋ̆{��3����4�o�6�fb� aj���^Uq��>�E#'��ɢ�e��,��%-,7���I�RyZq��jp�C'��*oֶ�&�����kZj�)��)�T����Ӎe@3E9?h3��0�'>�_§�j�����E���,�V���Ftg ����� �6h�ɺ�ų@F)��5��c�sɒ�l�9��M׊�O%`���� ��CK�-�ݜ��Y��n��{�����\�Fw���E^�S�Ø+M��uX͗ܦU��P�D����:�bC����8�f��P	�'T�:Uiٯ�!p����.�6�⌃��7�K�N�sd�G�k���cIK*�.^�c����.~��x��s�A�1B�C�Ű�� ��eH�v��Gک�D|����!{��������$G-�/���d2-�%c?4-��
͸�9~�����$Y����1y>L�m8�`Q��~"�Rd�2U�0 �~��y�4)$9���	W�f2I�]L�&�<3X:&W���U5!�9��RUzN�;�{�H�6��en")s����Σ]�*�0��%}G�t��>R��͒F��L����ϙ�dv���eV;w�)z��EI���Ї�$I�aS���`�b�VA�&�	W$ݻ� dt7�+fcM*�!6�+�)�k���
����������X��0Fw�G�~r�1�4it��;�z�u�����HN��DI �6��Y�
WW��8p��,ڛ�ɮ�~����?z��V`��Ӿ���c�l)���](常�C5L�4�fE̔�����L˕��O�_�͎w��x�{o0����T\����S=�nG��n� 꼚 ��s��2�)\��Ӏ<�Sk8��Vj� "E4ķ3}��9���Y���c����E0Sᯕ���@[~`������"9O�ٟ���Ҕ��H��p�;����-��Q��b�O^�%�VO���to�zz�*m�������y�C[��%�B������X�ۿ[�[���7��l+	�����Y��y������٤B�r!���~@�#�҈��ʘ�w%ݱS��5V�?�`�@�v��j�����b�׀��W�����@�j[�����A����\�~�ŉJ�It�#b=��x��Vǣ�im9R5�Ʀ��e�B�v���SlD�0)�:���S�Yy��jb�\c��Vү��dP�^PPm[�[���l��,s`Z�A`@�A�\H�:�Y.9�t�O����#frV(We<=}�|�:�p��� m)kpJ��G֘s-�7�/��$	}��t"���\�i��d�>�1�?}����^��~t/��V/�&UHŠ��:���?>�)��hA/;�d��୲���¥$�1��-����\� �f3���h��(��ǒ#`��"�+t�L �;������̄'����rg�,i�fƖ-�����l�\�����+)K[�T�ڟ�_���y}�+!�"��<��,�Sh#ӱ9�3�{8Pj̡�������.�zP~,��)X��+���T�%Y$ր�4Eu��-��[3K���KՍ:qvF�J1e:��Y|m�����1�����=AX�o~M����ǎT�@��nDǊ	e+���I�9H�o]��
#q��0�[�����	��>��h�c>�-ۛ�N[��?6�ҙU��RTf�`�D.�[�0*/�.������**�4F��w��Vۼ���Z�I��g�"%�+�l�O���|S���t���L���A�^e�db�>$�-\4�E2ݎ��h�=y�f숙4���MJ��d8>C� @�`D��$���?t�Kzŕ��߼][�y�Ȥ��œ���ڡa��Ԗ���xI����D��_�׹w�]�5����w�`����z{��@/���e;��Hй�.�&臣�����W���i�(!oO�v.#������w&�%g@���F�Uo���L�nm{v�kN�pQy�n�Q�f4|�������/�>Mc[GI� w�9(uf�+9ۃm�b��]k �x�'��>�q�	��[mvլ��2�P8��i+�=U�m�LF�V2Dac;�8�H>oĠmy�@`,����Ǳ��`0���(wYzsŝZam�ɖ��~jceG�G_w%�d�$�R���n6�6��tΚ5�/
m���\���U9,�9��e��s�Rrd�yoI�*���u��b����+��m�*$�#O�fq�x�%k1\@Q�{��h�D�{�I���5�ڱ�9H�:��7
�*�	ܓS"z�?�㨄QhUD+�˝��[����S�w����m�^ Ѽ!�X���&k4�^�ƽE}����3�K胊��]Wۻ��'�b�;|JAtQD�-�(Ŵ%Ԏ���SY��D���͊���C&��?��떸�$�b�@�L�	d+�
Ԕ����VO����4��`�!^x�E�~$�9d��uǀ�
�+b'������3=H����<�ԑ@�$��RGak�X�֙L�K�8Y[,02c-�!��R��������bh�֏ZV�W
3����;�#���!��b�%\�2?�̿��|%�W���3u *�
CW��-�BBne��O�Z�_��tsq,�*թ:�X��Q�¤�
��1��nDU.	��4��T��3N
�a4�%iE��k��e0�9f��_��F���Ys���{���(^oQ��и�߭*=���h~m�(
E��B�;���?<=
��'�'Q��Gܣ_h�����Ǭ>��`�q�e�$\�� S\�,���~Fc�nH��(�hmv�p�"f��ܤ������⿗��=�	$��ר����ҙ|H�idȏ�%�P��ᶟ,a�p�@i��V|��D;�Hfg���1x�U`T��O�l<��ϱ��+���a4����+�ɾ��wę�s[�^ꩽr��Bh��\ҙ�����ê'M)N�"z��`��UR�~������3���.��u����5V���
*��+�&v�;Z{�(Vw�����}5vI
�n�כ�@��RN��V�eD�2�(!p�1���(���t
�wlT.2ۆ"��������(�έ7�{*�6$˂�{{�Z���+ �'bkC�����(M�����������L���J_�����-��$��x�+鱷�{��>�>;�ˇ˴��;~��������w��:��KF��_s��q"F�yK2"�2鞢T�����İw矟��������B}L6�����We_�"R��-k���$��Owe�͂�Y-�]?%�O����Ή��t<�5���2�39F)��;��ו�c�u���Q���y�����|_�6�1�̊��D�`�f���7n�-���h�����EyԈ����.�&;��YW��SB�fGR��JN���f!���W��g��Tʵ�U�1 �%�n�͔Z���Gi��p�e�[(���t��aDZ���=2�a��7�Z��*/�R��YyzZQ��.�Tեc�.�:�G�U�/d5R��o�g��a@�=vu�ڲ"j�}�\��GYu�^�-��O����ЎL(W���s\��R�wQ�v�qn����vA����2�%w�G��Ђ��"�#���,
]��-�_
gP��"Ɵ��'�!N4N,�(π|����u�����5/Bp�.w�<���$��ɨWA���v��~x7�{�]*-�fa������FЍ>cf�`�-`�'[����n��kX���GsU{ݛ��pFZ��o��� �̌�s�T�0��
�&I�w�t`��Jkv-9HP� APѹ���>�RFn��1Z������x���_�W��ɳ���-���j�^p��,��*��M����}{n��eƱ�bИY&��d�0
�Ʃ���&�.�,�֌Zn_�,�*�W�/Ƹ�Ѻ!m����J�@1"\k��e��nT�=��82��*�B�mU$�S��Y�q kJ��<ӌ�1)��Q�!lCm��N��)�o��jr���b����/}��ƴ����f�È�_d��7Ͱ��s
�'�V�H�Y�]r�:B-�
�׭^ʮ{P ��k��so���_jO�K����wYF�7e�K+K�(5���_������ʡ��?>���ס9
��%pS'@��͈�D#�U�/��V�(����ӄľ��ܥ.&%@�{�)�m���z#�a�/��Q| `�ȝ��1RN�(��(�kȕ4�v<����ez�=�܎�Bv�X �&j�����>���7�4�"��21���5!�ߥ��d0z5�] �A���CӁ�C�k����,Z/ ̻IfYf�7����wHn
F�`}�k�'p*m��B-*f��d=�m3D��/^�����V[�6��0Xs��@����Y�WP)�ʄ32�0�<P���B�;�6�����SH��B���3�Ȫ�7���Ֆ�E�d�2�R�t�76"ɫE�}
����H"�n7���e����
�D�˽wqbb��S�Jk}�!�N�\I�
�U5=M�|>1~b��y���\�k�Kp�p�\���q�V�}=2	g\5��چ�~�v�v#�C<���� *X~['Wh(��8dC�����{vP���$K+�W�����PQ�D^ä���g�+�?ww���
��M�@��T����?�0��4����r�4�-~���桉yBpa�8����d�젞��J5��+��yt��B�0�E�ȟ�o!`�P�h0�7L�&���q���d%o%����@�#*�3�L��MjP���J�Q�n��ߵV��=��bq� 7���V`l�����21�9���T�$��9hlW��A3ns�<���0��0�k�]�d8d2�5o@"'�71��z�k��p��|�w��꠯ی�7�Ʋ���"�MA�i�#��e`�u�|tA�!7�����#4�`wH�#�8������:Ao#�gߍ>Rꁖ��wR�w�"���{���T�nozZ�����v��7Mh�,5�dZ3Emizsy�C��]���.E���y��z����ԀO�����;���l�Q�M6�un�_=�{
g)��GPB����J�C����X��x���� <ټ�Xu��r�Y�[ݻ�	�X�}7/�N䕛�OK�eĒ RN��i
�f�"G�%����eQ�^L�W�3�͏Kt'���w)@��ě87@�&��ʲx���E��X�v��
3l�0�����Lo˞����V�O�tMS�XS�5�,� ���m��Мh�Q���2�qg��fY
E�qV??��79&�`���M�U��H�p.l��y����z����;���x3�}�= � ��+�g�D.�B���2��q;<� �V�,�&���)+1l���1�~�(��W��xV*@؅���".&O�9j��CO�:���g�v�țђ�"�����Z�:��w�+��̆���YL��!������mg�H$|�GAѼ�������1Wes
+�����t�'�a#d�ͦ�J�/H�K���r�E�(���)��N������;��Di�/��7�,�N?���w[��N��c���<2�Va԰\��W���hߖ�c��X�fa� ��F/\*(��1G��@I
 p�'%���w��0�f�Xy�ب��믉�@�,���?��DE�0��*f�B����)H�c/���L��C�z*���q2�G'�*�u�������zH�q���(4Z辍���fL����bME���'ܝH���ߓ��!�4A�5A����s��K@�����|۪S�� ��b���Qt����	R8��/l�v�JkՇ)�p�pɑ
��o �(IEC����`ԝ��g��V0�V!��w���K�=���3���� $�̿�BE��Bt���T��F�z?9��0Du��ջL؂�(�h�TK�n�M�#k|�Yå��I��U8b�|�l�AL&��d�L�+�S(z�s�P�C�kWҷ�NPD�]�UJv'&E�ԁ����Ŷd8j�yw�X��/��0p�T�cvr��@�遣ǫ����1}�IR+=�$M�(��.�t`�P�����i!o�>��rKt�����T�Vi�.�PDK!�$2��D*���P�z6a�΅�Q>R��;������/�r�\�]��QC�U�
vx
u݅�w�5�l �P�/���tiɜ;(�fY�&���'�%E���;<R�[45�A��R����C�=�V��)k��`��xЙ_�.���d=���E<)�ZI�$| ���9,xH �ϣw��2�7[��mn�p|������-^��!����2m*?{3q�pR�b`��K���u��ɑ3���<p�9@Y2���^+���5�b1�B�. ^��NW���
6�kSM�q�,�2h�
�j�IY�����ֵ�b�ŗ�5������~�������9j�NNU\��8HWRLK�ge����/T�qt!��UK��==J�7w����ȭ�Q;>2m.[�_k���9�  p�h����@GT��=�*�u�i"[�ލXP?����aYM!�wSUDo��Y����n��="��x��
HxJTiyv���{"�
��[CII�K�:���|��I�0��cn�z#�,���4���f�J����F,_	{{���IE�#5����v���i���r�v�
+z�{�7� �S�����)���>�'ݏ�:.a<�NZ�c[�DW�gW8�Ÿ�ll4��E�9�������.g�C5O{%�m>�bg�5�VB�����W�71NhKeF�5Nd�������ك�H�g��Y.�O�y��o��D�hZ�@�4ۯ�m��ġs�ߔ��KW_B�X��i��z�;|���hħt���N1�n=?t,�����{xb�"�{=fսlX�� 8��i8��v�^����i��F#L��^�(��T?
l�I]d��U�2x�|�b���0���YҸC�p"����g��� �S{�쑅NU� ���W��t"����8��{kmY�=�?��p?�f�ţ�|�Rt���qT_O�Aޛ�, i�� �%9K���o v�]���G57&5%�q�e�ߴ���QH�����2���"ӉQ&��3]P:Pz��e�7(��<����VؗV���II�"jU�=����}k��b뷺��&6��In椭|�u �<��3�E�֬Hy������9�k(�An��l�%�n)פc��U�K�p����ZZ��]B�X��@�JJb�l�S������:�֙�����gp?�I�p9��.�d)�I���
�m䰼y�S3�u��"nYZT�� �r�I��}J��:�;���z��<8QQ8<�E�/0�`��<�?Ǹɟ}����r{I{[	��؍���R�J���7F����$JLUx��,�^Tx���!<�9��R�x�l>��1o[gGz̢$^� 3.Q��v>D_�KN�{A���ۚ�?Uʑ%�i��Jf9��=qR���]��~c��4�8(���(�R�0iS(�(#�j�?�IX��\Ԛ҅�sbH���<�TP�7��j�5��ǳ�(R�8�$4���=+�dS�g����G��A#m�:�6Q�D�B���Y�IXB�m��r�D��	RTo����rޮ��{� <�1�"�:����Ԛ�O�8�M������V�$���=r#�%�lۡ�K�Ρ��)�TX���4���W}#Ք�w�-&�TK ��%��i|��Y�!��ܝ^Kɿ�f��S�����-�]&vi[��WzF�(`"�o 0���_�}�݂'���Ґ�F#��i%Z��F�3��2�}I�@2����_�zp�2:��4YU+P�߷������l���`ϼ�mFԥ��-+��]��o�l_���JҸIN�S`:@�x!8@��dۂsV]H޺�l��0Y�����1����F��mꚢ~���֊n G�&�*�!q�X9�DI���3�"&�Dk��>��Lµ���-�	��Ow&ZK6:����"��l����LB>s0R�S_g7��A��:^{��3��"l�sԺt�����A�N����}q+�)�&�{m�`�=��{�=�]�m�Cԏ���<����d<��H- G��*;F�v�Z�z.�Z"h �,��к�n��"�e7}��&��C�4Vi��������A;uTd�<�X�Q���_l�aho`L���?���az{���4�Ŧ�c��B��Dm�w@��*M�����>[j�@�;�� ��,��1�$�5�������9ke��(���G_�L��h ��|��)�2x��x�N�4� R�N*��w�1^�� �Nn�����Y0���V�5>b�Y�.3][F�&�v��v��d�%�qC��
��P�|��g���A0��T����ƥ�����%Z|�;u�ᷔ���>����@�}R9mn�/��Yd�1a,%�j[[���q^��D�N���Z>}}�ã�N!l���RR:���9sy�dn9�]��WJ�.H7�����+����f��9�O���ɫ�ܬ�#ϓ�����Ru� +�ޱiw����
laqhs;��2ǯ�#��!iEx����\��b߬���-H�c��~'����WiU�7���bdW��ܟ��5�jy}xt�D����O`�:��d�oe���� �'�!Wu��J
�>��Z:�^V�p�,�����˼�����ìW�3w�Tx�tߑŐ�ݝ����;d����V�����yKL� x
d���9�<SS�o���~�>�@܃��Xf{羍�����[�/Q����Jw�:D�Y���x�(��8�gf�ڋﵫ���qOY\3 )�~�D�+X$]q.�OCDr6Z�_����b$�7�C�6>���!ԩ��U~��ݧ[x�R�Ɩ���Q�(`p��u��PD"��%a	�(������K>�҂�`D�ӚX��P$�Rj��3�GsY'�D�!���[}�-��U��i��J�H \��u`������Úȷ��|a��f�@����-���偁�EYc����er����2�u�?����Y��SF�<��4���x!T��\�u�d��-{��]�_�B�ܕ�eXja%��X���)�)^kP��eP,�uWɌa��tU��|q4R��F1����K�^���wm�	�Ӳ;�RC{g��]��B{i��W�T����R(�M�j���>�5����A줲J�^�y�i&��u���bT��wy�AR���R%��-�Y��'�N��'�J�(�A)kW��A�(T��9�]@,������0�������_�w-`<%ygNJ��c؝�Z��aI��+nmR�^#����7!�j�Sq4�"���5��]���KpF��i`��V���iM!�Q�,��膈�,�7}o�5h�J׺zG�x5��P}TEd0��G��1�>��|�����3�g��N��qaBf���6�4����1\Gz;���I�.L�[H<��Gm-�s{y;��3��iT���,�+�h����.	�Aγ��gC�@��g+}ܘ��L��j���ζ$i����)M�+����kGbN)e�L�U"���EqY�۰Js��2ѷ�58�
r��U�a���T8�MI��C���l/�]o�⯷c�Y���KҶ�A��w�r u���ږ�����ö�D:�2�� T`�pI;^�\@}8�!3��?,����������y��[�O�r��X��ݘ������g.����%	�S}7�2�W?>�qh��79m�č���#��JY#�&,����w��Q�<٣q�[����+���q����zn_�0�մ�����y�����M��e�*��N���Bi��XA���\��T`;឵�D9��r9JBQ�T��Yє[�5�4��!N0-.��GąV:`4d?cl�o�,}��J������ڿ��O���@��Y1@R�ǒ��/5�.$>��z�}�:Q�0;�4�lJ "��g�,��
q?fH��U9U�{#G���2�>1Ը����e���FY�&�%D�J��\�n���Z4�S��=Gmڌ�e��`hS��ye:&���- �P~m�0���3��`|h�ٞY���,���x:��2s)4��u~e�r.���BS�wYz�,�w����j�^�9��Lú*Ȑf��0] �p{�"��[���Ι_�����Nۋ
��<ˌ�E��\n���C�DLO"��Q����+9NB����7+���V�:'.1֞��O��??Wʫ���k>/��26���43���w��`���EG���&%��'���DKN^\��,�<	͡ �o�%G������a���<������4@o��3�� �:΂��)v��뱈Һvi��ik�%5���N�m��9#
�t拳:@'�_��Տ�=�Ji)d�[�/���t�?�5�Ok�4b���tB,��bn:��`wh�TwVa�1�\���zТQ�`�l�ҿc˖=��#�4S��:#�ր�r����2���.�^E(��~���3a7��=\B�'�az�8����7_��-�zۨ��sd��&�D+s���Q�E�|��&���ue�q��"w	 {q�H7�j���TdЬ�/�����LZ���<W#-�����w�V��#��>���g�r�Ӣ��qʅ�]�����l#�Ia.[)dkh�i袇���'+Moeo
2��ǅ|�#PFk�	�A�R����H)�Z���G�A�����e^+Y"VȨ�-T/�m���s�����F&�/�U�������ո���y]�[�3BO)\�{e䋜^!g�Q���I��I��uLd�g��90qԬ�Tߝf��C�<wo��{Nd��0_d��B��;Hn�r��o�A�ƹr����a��s���c����u ڌ�S�[x�Mb��q�}IH��~?��e,n�Jc]�����7e��4YS�.C����cakk~��Ө�`�Y���M��ֆ�T%��ڻݐ�m�������1���\��EHӧ�E�!�(ا�@�iH�[d��$_�wj{/������%�XM� @�
�+�:0T+��T�����Zo�A�W��+]��{E�{�A��O��8�pYoC�?�����4P'���(A��Z��,k�����5���k�4�5���|�$�!�)P���X�(�]��n5M��"S�a1�\,t�`�&43��!B����y���}U�ʑ� �a����$t�q�7Y������`kO�CC����͂34��L=۰4=%Hr�/���#�{��XE�Gޙ�N]���������'��L�5��_T����8�^�mM��P�ԯ�9����[��ǧ�����y�?rd���>�y)��O2P >�
�x 
�)����O��ˏ��%)�F�;�(4f�/<�Xet��L;b�6��8Y��:΢"�L��5���{h,�Q6ޜ�G��Z,��-<g������či��Zf2�6�Z�
���h�,���E �#}{�V����CB�]Ӂ�<P], me�
�ԪQ���ϥ�"�D)U(��v@S����O�E��|��?�EbUA���J0a�7��E������:�X� ՋvA�a�]+DС����7�$~@��ٜ@;�q�BP�{�[`�hn�}̢��o�w�LɆ������� ��4C�Q�������1�Lu�8wB�*����j�+ү�'�E7Ϧv�)Gh�V�^�{r Ia?)�3�Ү�J�	3h���'���L
A�NV��������Ji���uz�R/ҭ �v~%K�p�t��t�O~�y�s�5��������>!�-��gu�ز�'E���t�u}B�MX���>QR���o���n�7�he�u=�j�8*�P�*��\�sԆ#�p�o�F|IR�5*!w�5mjt������1Ǟ"k�2���+�w�y8�W�4�S=��x��-E��طIu��g�5C�����̋r,�hD�tߞPڎ�H	tBX&m��C�+�-E^_`�*���|=���da�-prs��*qZS4@�׆�A�FEY�M
���G��7JwV�l�|B�$xR��(F,�X�7kC�:�#��غ;J{@�"��]8��e�UĦ��U�C|=Ǭ���{V��8y����*��"�5I����J[��7,���n%荼Ɔ�zReyH�,$x���>lY�<}�̶�o�KTe�r�Z�&-��N�h�"��!?�{�LJ�&5�I�� �mv��Ֆi������|��i�����ɽQ� C��Q��+�K8�T�#��T���1�g��kq'�H�������M����)�h�^TՁ-���y2/��:�<������hʏ��	��B{	j�e[]�R��q���.�I4Ҝ&�2J���i��,zi������T�cb��J��1��e��1����_	��p���Y�y�`�'^G"y�&bJ	g�O��\�~8�7Fsc��e��g\�*�:̢���t`�s�?�#�Z�L ��i��$�`r�k�N��kcT�ډ�@�,��3�̓���+�C��f*��`�!f0wvo,f��K��y�!�Mc��TNi� 2S%�v�ۡR"��u�{l�*#�� r �,������;D��*�!�-�W'�.�c8���'�ے�Q�����'c��������Z�����ß$�`���3z��E5�ŗ�jSޑ�Ŋ�B��ox	�
|��0��+H�D�\5���{a�#?X���E��W� 3K�d��w/�C-���܊�7�Ҿ��/� �l��þ�k�Z��a��A3�Ob���>�#񍘢 R�A8�x9�4�@q�pBv��h �����)N	#��fy̷7��Aʸ;�/���Mr��}�P�a������Ȣ{�	�aK�F4Ɓ���r���*AeL�1t��D�9j\����*&~u�<��(q���*�:"�z[�m��ݍcG��Nˇ���\�Q�\Y<�iȯ�EZ��t]��,P�زA6���J���M��?ݦ�1�Ď&�� . �f�S6�^~豧
��{O>��=�Q�P���|��x�˕�\ҷ��eSD�A1_�K�9�T��ޯ`�(l7;�W�"u����	�}��5� �'���c[�]n�H�>���^�v�!s�J�v�'�6�9�!?G@��˹V�_z��ĉ�n���!GyXh*R&��؏�˩Vbl�܈����.V�VAO?_�����WnMҼ~QH	Iẻ;t�5��ѓ�P\W�2��1Jl������:����Ǹ��.�IR�6#�	��y=,l��*��������oSO�b.FK��� [ YY&U�(�2߱*?��|��^J��:T)��Þ3'�ES%W�O	h����6�W��;>�,^a�t^ܿ� iA���a`�^�}��t'���R��!�`%X 5�Á<�Q�HD=���F&:�TY����2�L�!�S� bQ�۫�$�"���Fڑ%�=�
�(�BBQDɫ�3�� -�<;d)�ܦ�����f�Q5��k�`UYf�|�Wӭ(�w��VL��R0��~�db�X��آ��$��D{&@a�謟�����mZ?�|�% ��I4�_�����ޘ~?3�������(��#��T��*��̭� �L��Z�r�#�����Mw_�jGv��U��������1Y���&�9 ��1^�IE痿XD�g�ï��Z"�>����r�2���3���6���}���(��?�4*�	��:��4v] ��H�u�q�}�
�S�}���v[��㉪��o���C��d�w_C��L���n!�������n�K�>E��6��j֜C��z)��M?���qMf��7��a�a?fn���dm�$E7�۷pHć ��uɻ����*��#���~��qg��J��V�i�7l�ג(S�ex-�s
.P�w�U��X�$�v�]_��f����ì��R����c�2���}�d�n)����p�EpA8}�� o@p@D���'Eq�h8A��)���B��[F�5�E��pm;��ܿ�r>�<c{v����N��}k��*�E},s},���Peʌt�x����ǭ�EJ�Z*�먍r�"��.�_�w0�	��2�B���p�b���!�4�%�Bz��P@�sy2>�D0�=�)&�P?x��k�f�I��V�w&��2���O6��P���Q^ ���Kp���ۚ
��7N�5�ĵ�+��BKp��rw���:�����^��RK����*��>/ EMKX"�~>9#�1·�tv#����o.MD�̱��u��S���!���C�Xn��,乊bLD+HHF!7��%��x�jM��aF��&%2�H�e�1�y	>�C 2zQV˦�G?�b9B�8��<h�\E�z~��jٴe�=5�P��<7{�~��LA��aʖ���=ǔ3]6!�@OA��(b�U�.'��/U��n+K�~��W�#vߓ�"�y�D5d7��vY��c�����s�)~ ���e��LXG�ъ�uEkʶ4����ѿ���-dl����KLX��3�NH���Rv4_q2�,�rۀCFڝf}�i)Oi꜀��.���y��l����J3�,��5���<��ΫQ�#���9jx�6'	Cu �#9}�%j"B6|���ڎ�H��u�	��U%��~ǏU���f��m��nW�����r%��G��:�����PFh�뛑?��?��{W3���
E7&ek��	�2&���S��`Y��q�W��n�6'�XLm��T���f��/<��e��dY��s�95m4��V�5��I'Y��#vى�ҦG�.H��
F��a#e~�bY����1���\?�c
{&��2A�0�k��Wސoy� �Ċ��9�W��u���?����:a_��+R~�n̈́��B/��{8�W:�����;L�>!�7��v�
[I�/JM�Hk����dg+3����M�ॹc�3�$�ͳ�k�*�N��&�L����?)j�9v=L�D5,��$/Ǆ'?K/�+�&h�&���a�*���+���P��F�O� �%\��X��yr%8�N�Dx�7t?mhbSA<��?����iP,@oUJɇ�lOC�d���	Z��fR����G#@�a�mZ�?�#Kn(J�֕���x�0=��)[#��ic�a�����CM����꫍�!�Q�����p�������.�k�,��� I'���)g��7�ǝ~�7]X_���k�r�;�Y��f���9��i�M���f�[EVzRJ����V���v�i��?��W8G���3���kqH�����RG�Dҿ����% ��:�����g���ధp��0�zL�?��Шצ�F�l�D����A3�7�E��%��d�$s�)ٱ�N������ɳ	��OR��~N�vn�65'�
�W85��R|V�i����v9Th��܆`��W4�*k̿��5	q���(���-� �
 ��(����7�L�������N���o{��_���q�4މ�,�F����'���|g��G��)��B�A&�B��:Ș*yOj0JSP�<)uN���	}�V���-�C�,υ}G����tRO�ӭ��Kz��}��RXz�0�?��򁝙��mk_�wb����=����M�lڼ:�b�C���y��n��l��A,� �*�>�+��[bƴ-X�(n�L�(�S7��K�A�a����ʲ����{�,�pG �V%u|��i-��������T�J݅n�z�H�=C'
��<LE�_����ꖏq��r��BDp�r�yl�ꙕE���X�ڦ�s!�O�cotP��	&�c�M��I���	-��w���r����nW^tn �t�������
�T�o�ۖ�I�`y&�AC�D7�*�E���C����*�w/�>2��K?%?�O ��g4ܕ�{4��P ]/��l��P����If������߃c�֧��h�8K��|^�+��QG�&�Vy3��K�,���:��Ӎ�оo�����@P4ݓ�ĝ��C�r�
9�/�6)��43"�!3�����%s��-.}�c�����3͛��|R���yW��_�����)�ʫ� �=�_2�(��r[En�fXK���K��7^��'�t!a9ԍĪ���N��n,��E����c��e��&gl�QΒ�:%��� �x�"�~K����]FX�W1��>�J<.'�������i��P���A�H�)�H`��I�/��t@w�|1�]�2��İ�U)�b>2�I����i��}nT�0;1��/^���ܚ��j܌rA�y;�F';[X"��2�(6����C�:R�4�������7�;-����ovϊq��å�'68�e=�K���M�kn<�w�a o�(�
08����t[�����ɏ��n�g��M�;�C}�DC%Ə�0Z� �c�UſH����&�:h��n�������wc�7����;-�z�F��w�d����+�gj�[f0� ���&��>k9R�cL3ކ��}�$ˢ�qH
v��|��]b�M?I�b ��QҶ.�����9?Ctt������?�Ļ��!��.�����q1Hh�c=�[��H1���+����� )���X����t��2��>Q�HQ� �+ �����f��dlx�%)��U
�K�`����{�� 9'Å=�*n� �W�s��T��uA�����V��k �9ׇs�9�Y~觩�90y��k�f
�3��ߣ�,�����Q�����`AȄ��C���Gبs���40c���eX�qLi��'Z2��@��3\@��FƆ��7�`�͊L��Q�˓U|��v R �����C�o�>��p/+<!�4dz������w�b�V�́[��G�.�B �yn��J�-��B��K����}������+X՟VP�;^�s�4��2 �`'�ya4���aa	b��%c���b�]O�P�^�t���B��?~���,<��¼��\����2L��z�ǂ��B�e{�k�!��T*!A�^��t���,��Z��
���J����,l����IN���ş�J��19B��1�g����"_VOzx�m��[�Ӡj��=6M�K�C���5WS�K�4�6����h�q���,R�Dһ�M��l�a�;��v��Y�k��h3���{w�9����`2��6�{
�����驕�ȩ�F޽�dz�P�0J�6xv���$V��Fv�~i�X�I���Źބ>Ԅ��7k(��p��5 _h���X�ڣ��hb �S����?�-���{� /7d"K��"�6�s�%Gh�&���r�f1B�x���oN@23!���N�.w���N��L?�P���yOJm$&g�}�Ro�W�:��W�#3+5Z�+�¯��,������ѥ�J��?��S$^?(�q����qr��v�?�}�q6�����)��w�t	�[���Z�c{ 5������B~�ͣƈV��F8\�jB����5i�.]����V��|�(�S������H�{��\����rl.G�e�d��k�^;�J�S�����e����%,ھ����������e�F����8A*�f����!Ij���_iEtO���/s�hg��.^������2�.���>TՀ'��-����8m�P�<�MN�yb*H���lT��Tv2�%Y��	�8�5�	�#3��8>?J��1Pm��������%�F:W�\�������68�uv�ݡ}%�aK�
9�/ɗJ������L���/m ���6�
OL�=��S0���5����cmp�:�q�*���M8t��wx�R_������u�]�9��.9�W��5�0ߒ6Z�A�� ��z�|½7u,!-�<Uei2+Pӄ��؅6x�;{�r<�e�*��@{%1��_T�Oě�>ڟSl����˧���L��*��S�}�1H�.��D�����]����l��� <�����j�e=��(0�O�hȊVކ�*��͝NƗ��W�y�!�_.�g��J*�qq���;�L��ޫ^۰�%����s���n��ކ�C`͈j��zs&XP���튦��=�e]� ��D6�A>�hMk�=�ݣ�E���t�=�^~�B�΃w!0.6==M�R��(��86K�Q���
���1R�T$�bF�^,"�380�8*���qyY���\K<�$��1��Q��y�Hw�����~��8�v:�~�4�r�y	��v�K���H]'��K}�j�c0���c�qE轲A�D.�dB���	<Hp4�F.��]u��P5X[~�aA�1� :�����Hm�H[#R
�_E�a_�1�(i��x���H���=A��|��W�̿�@_���V>d[\!�d%^E��J��P�a�7���z���HT`��X�>ꆙ�[���Z�X���,����KHkF���B�a��ΘZ�z�O�sX�7�£���/~wK�2`�jˤ�m* 3�l��&�!ki<�/����g!��rm��0]��PzUj�Fy$�`�V����	}x�֓'f;���Z�kg@�*r�:�֌�����a�p�v�b�p^�Jy
kω���0PY�����1�T畩ЄMlo1��:pr?�6����!}�JoN )7���W\��E�,�Ivj�?�c;�%�|��*�3+e���\v�O���C}��<y�h�X=�.���?tW6�e�:G�_hZ<c��!�/��H
5m�e���X�Q.�x1����O���|���U͍8�.�����^2qQך�'x�Z��8d6S��fA�������(f�����"��"���N޹�w����4�\�I7��T��D?>��u<��M�]}�}��-E��e����e�����g�s�+�<mf�����ӚbA����o[�!4(d�#�յ�.,�ڡГ�Y��z��l�&N�iL��P�?�礝n`�;rsn`����-:qp�Ÿd���ͷ�� +d'G����ڍ�`5İ<�L�/t}�.��>��!  ���Fo7`��D�^�v�B�����!|P���u�
nN7�?D�kO�zz_j6��*���7�>�Ŧ@Uc�ʑ��m�~ʟ��X�A��!9ج&����0 �dq��������%�ਫ਼����T�!I��&�(DiX��� R.0b"��A���ob˵�9�T9��_���X{;1H�ZJt�R�O��y�o�2}ƺ��B�㷶=�~Η��\�k�6.�"bBD�"���1.f������@�Q���%���^��������3S���SI���8�qzG��]@lӸ��R(�?�P�ϐ^�G�\Ҩ鄃2����m#�zp�ĥyx2����\M\��<�喅_*_���S,�6a���K��[�[̙}�GĿ�B��n9r�}�ot��Wi�~8s�(P��~��;�J��f�a�= `���#���W4������̉��E,/�J��ꍭ��Xa�`�eΧ�E��'�e�
���Ci�`���)�Y��፯�#�޺��TܨTbW�Q$��h���	�gr������L�U<�/�}�J�v�F���8��Zl9�}*}a��f�PN�%��Y�dU �>���, /�� �d�����H!�'fk�ڝ�1��q���0
���o����KAL���Һ�����#����������iE�Gh�Kv�p������HA~a����I���,�5'*���x<N�<�nз�bf�~I�{,����3�L9��BS��X�m�ݑ4e�;����F�3iM?��o�i�T�c{u��'�δ�Yu1�b3qR� v6�.%�,)���>e�v�*��L�� �v�f4@��~xi?�8q,v�������&���Y���4�FL~������k��c���5�c�8|jz����Ӷ>�c�U0g��dK��C���Q7���q�*+0����9�?6�
oco6�	p��=<�%.?��U��J��	r~��m�M�I��ky8�`�0�d} 3�@&��F��l?�U��-�Ҧ��8�^��:���g����DH���-/��Ҫ՟�/��Vke�k�u�q���Y�1�y2|D��}�:y��Sif�Y�p�s�&-}�������#	|���}s���śȸ���D�5��^�d4����zε$*[.�2Yy�V--r�)\�B8d�A��K���eƬ&�Ɓg'= ��T���=q������|�}[ �ڕޑ������0 �J�ѷb�_/o�i0�tl��in��|V�O��!Ѧw����x��/�i�b��[� ��N�Zl<�=��O�,���))!���|/�9m���<�wv<�v�b;�<�l)��<��C��1!UN�8���2�d���o$J*�zr��� (Jc�ú�:M��oi�Đ�z
����� )����P�c�Y=��0(m�~t8��@ +N��8d@!M[ˏIL��E�d�\�I69��1�����s%��r*�ߜU��lI���@6'mT��k���r�i����^Sืc X}�	�Q�ښ��������$���m�����4,���;�]�#��N���-�L^ji�tV�X����`��v)Ke����=���"5��__:="~$�Ȉ�ͼz��T�r��S�����x�Q���qϟa��^.m�'�*��WjK�/�yhI�X>���M���fK"���䑚���JE0Ŭ���[�#>t��׎��cpt<?D`.}/��p3�64� $�V�E�t�]�����r�x#Mg��nN#J7�ެ;��WOSu�'�?�qi�g?�J���ܱ�
0S�	�8Q+�6�U��f\-�T�> Gf��&
�egg�~��m���O׀4'������E���R�/*��D��6��˥F�w�խ�EB����,��,agR��i���ƶN��&$e8��	����۠�[�~�v��y��f��J�v���1Ͱ����6�iP 3���hZ��>��;|��Æ�ڕ�i;�1�K����w`J�e�Z��&?v��Ԣ�r,������&E��@�2�6�5zr�hs0g�ݡ4zE~!;]v���(X�h4�Pkoޚ���EzM�nC�Y��_\��z,,�Kj��E6Č��JX7Ta�D�Y��\
���+Sk�Z�J��/�"�@P0v��<�s�V�=|%��hރ�#Dv���}��?E��Nf�{�8A4��5>ݵʾJ:h�Zl���`�N�nlZ�:A��v�`2�	�����;��-����\�®=��0�@��.�<��`�C�[�Ǳ��&;�K�b��O�=�P�_�!�3�ʬ�=9*3�!��#d��=�5�~�`���*k��3�LA�iW�#����֡tZxۋ��l�p�Wh��qyL��yS�3"��,�~�2g��c��X3ǣW��u��|d�&�{�L���˟l;e� �����+���V�
@�c�`T���z�T���U�7�$�b��
M���o������{[p�h�c�,�<����Ѧ�qD��͞��@�P6��/�.�ˉ��*P0������X��1�l�ʓ8D�J��l(WV�g��71��x���7骆�ǀ�Yw�R*�&�Ϟw���m�eЭr�0 ����:\�Bƛ�2��\��9_��LU0��������s5��eFd�Y�=V �i�E�t�{rW}p�b�tf}�7�_�~���VD-݋��T{|S����q�'i���	��_��=�R�xFG�h���2��A�}���*�Cs�}���\�>�
H@�����#0W��y�740�B�F�79#z�R��c�L���� ���e0
�r�>v����r��~y/��6�ƪ����[OBI�s$����&�A.	?f�����aq��w�6��<�tnf��Tȓ�u�`��Z�L��C���Od�	:(�I�O���]�Ɛ���潯�oٽ���h��n;�gk��n�Q�/�H�O��9�� ���u��9ީ�-$4C�;a����*�Fle�c�%���2�C5NNv]ć)��:K���u���1�ٿP���c����)�M�ڏ������'$X�B��)ʅh��*�$ְJ�����%@).&ˈ�Ǻ��H3�&w��z�Ë�X�x`W};Du�L�U���h���A�q�{���#1������Æ�9OY���y���˥* �I2s�����qQzBO�I��g���<����1*����B �>c,y�\1�*x���X��+�"��������lN��ʦ���-h��͢![��At}�V��� ���qR�١�j�k��f�Ϻ#�n�qx���Ҁ�8;h�H��TR�d�W`KΡ��KN��}����sx����DP���y�?�� 5>�8P>>$a]#D�i�㉉%�g�S�ʻ�:W�J�i��؃�P�P�
f��!e���N�O�=`v�<f,��n�#_�Z5iN��gJ.��������q�%LF�~��P"��-�ꫮP���"�D'�uu<FC>'��P�o�wx����,`�����#��a�햪���וB��h��unY.�HR����$P�$C$���`�g�nZ:y��-4���bx��Do�\��I*�����9�zpKnNA)�Ϧ������=�xOIC9L�"�z)�<^��������/�ndIV��\PMF��m�Q�v��|�b���Mϻ���\ ��*���O��s���� ~-�Q���-T�A@��'�G󦱨�vpx���Y�T�6���� �$RN�k�4��XXm)5� �qv~k#ƞ�Xg2��{0%�����<'�u5�A��b,����ꡧRdP?H��fI��#o�?W���-��: F��0��	ǒ�SZ+�(���n���wN���R�K����i�2d��L�'���'=R���^��oqSJ��@%�Q�% ��<���E�]������{*J�A����Dg�Z[1]�>����=,��BG8[iI]�@ۆ|�����?�䨌��n0�}ڴ,�슲1����9@JP�L&c�k���z�FN�S�ã��3
��̃lh�[{7�ln�{P
�mC�m�y~�&����U#=�
m����8�9��#���ٻ�����}u�W���g̪�:
m%h�	|���_�~��~�>E#A�B�8�B�U�h����'8��gIU�w-�S}=sd�!��L%���,-�ָ���(_
��@���f��oO��g���֑�����H�8�i�e.K䢰�K&"���=�24��\V��Ԍ��Z6�ۣ�P��c�f�3v�p~��_M�^&����l�(�k�Wӝ�����$ل�)�}~gG�eeD�)ϝ++Ưk�R�_Nd���-m��dQ���2$Y^/+#0�\^Ϙ�\B�JJ]���5���7jB�y5`��~�)����,6맣����ÄRHK���.�#_B�l���j���h�zOS(����5��KI�8Ӽ��	2�-p�5�=�)7Kt�h���������C�Nl�O��h�ݡ���1�I��ထY��k���h ���^�Bq��V&J�&�M4y#�����6j�^;$�9�wW�$�o�_���B������U7[�d������� �ۢ�&ȥP�
��14	)<�4��%R3�4��~���e��w��������*u"睙��yO��C�.�(^�4@Dt*퓇8��F�� ]a]!:��ηI��yU!M�|h2Cp��(��P�8��tWZd<�!�0�<��ku_��)��=���n��7�\� �Vw����t:E�6f�r�*D[�2x��Gk�S~�.qh�'�j�Ez�)�q/�� �
��!����������nIL����Q.>0F����l;?]T)���5�i��1��z�QF����2zjO��Ft�xcn�9�&Jj�a|3W�Q��q��g�.q26�t�2E�J��g'Y�L��� �q��R�_����,a�E�Oh��9��& ;�_#��7A�����۟�w/7�����*R:BW�@�uN�; �uk�U�'A],���@�<�ۇ��.�
���|j�z���N��I-R�A����\���s��.^�Y�cgH7��	"/��g6�ʅ:)��]�"0�w����S�F��=)ߗ�l�/;����9�+El�J�&���b-R��GM߀UdfU���t�w��9"����X���T�p����i�I
Hܿ/\j��w�pDh�lDIV���yY�	w�7�jA���&RWq�W���K����]���fY[h)w��&���tx�Pg�;|�,Ӳ�A�����Y�tt�͈�6��?��r��ԃ�YD�@��>����� �<�b�����c�n܄o�m�u���gb�C�Z0���0�&'�c��d���:=KzF�-B-��/v���C���@y ��p4J-�'a���BJ�Ȟ�i�$5A��t^�_�
@I���C?�a�Tu(�YI�H�ke�WYG�I��"J�[��Q�|U:\"�ԏq����8��g���?q����Y6��J
��cT�VƖ�PBzAx�p�K.rd<�<~��������93a��+��Ͼ�CwE��WV���۪�иs��!0h�ʛ � Xr�n����{n�r����<߭Jl�C��S��Vj�U�{�k?R%��H/V�U��Ԓ�x.�m�Q/#���-O��1Ix�7���E��}����Iʙ2�z�Ժ6\���U���]��xӊ]�0��(��	�`�b$�-D��:�~	6�F4#y�w t�
G�7j0���Gc�3!��ϻ��vCr��-�ٗ���9���*�����
r�2����q�|���x�b[=����P4�Nb{�UGe��$�	�5qѰ7��J@yx}v?��v�ٮ[6p��I>�����;l��Ƃ� m�EOiJ�ve<��#���
-Y�����2v8���� �����_
�
#k�5��*�>��M��&㷍�6D�Y��0\���6�cI���j�+���\��� dqe�m� *��S�t�j��q�y���ץ�#�u��T��T��y2?�Q`	�~�*�D[�U�(��s�K�O'����f��knb�PI����=#_��8��ffJ��Mw9��J�hu�:(�����"v���7#6N����2
�F|݀��G��Nv�n�K��Q�j��w��t�'f��diᄃ~�����Z�ED�L�����Y����zN��z/�F�p2Z����'Z}K=�<D��4�gX��m���+�=${{#l�8tg3��]8�.j:����	�d�^��[�/xA�JZ��nY:�n�#�����o索@����|}�'��C.Rcwb��Ӎi��8�������g�Uǂ�9������m�Ĳ�\����Hkˤ~U&�ң��])���/K@q'��澳���+rC�_E߉&�.��0�(/k�3�(@*��GT� .K�'/V�~]bI=�:^��שP+*���?�H��?!����bq1�Z��$�m�zG&]f$���ˮ1�h]rj�U\v%���@�k�]l����#D/DI~��e�;r����j,��͏����}.�*�J����Z�F�n-N��E�425�L��c���łt[�k��$\�0n���g�l(����+��m�Z-Є�{ˏ+�����F�# 9�I�J��ΗD�ꄍ<�
�i�"�,{fy��c|�!���4{��q��$�T���ɗ��~{1�L�#,@5��Z���iy����:�����*_$�dw,�v�̖�#A0�c�X�מT�����o�"�pm{���6����d�ȭ�l�n��� hH`������)b����H����ǯy�N`l�P1G�f���C�2d�����
q�^[�F׽?�D��S�bY��Z�LY��d���n~�̬_^t���j`j��M�����j>b!�q���"'�ֵz�՞,��&�,�)��#�2.i���
E3��X��s����m�ۼ��d*���դ�ߘ�zԇL��9ɜ�噀wp�Q	K�|I<���Ê�RF1Kh����K_�eI��G�e����׻������׭����m�W�P�dG>g��β�#/�:�,�xm.A�wMǁJQY7.	�ј���x	*�����%���7��,�X
�ם��Ėy�P�p��N�N�\5��~Ijь����=�*V�0����d��:����צ�B��� ��-��A=3줖�&�h�-�T#a���Edc�<l�-'��9	Ž����v�S�l��j�s�i,L�V�^(�����8H����}?m*���d�I�F	R�A���hHiK�W�/��i�Ik�Ow�3�)
���-��0������l���4w^C��r�d��!��p�&v��!M{�mY(��D�QS��� g4���yw0����z���0����΍�ǸN������+��H�p2@��4��%HypVu�o0���@�=B�-�p���hP5A��@��4�&��2ĕ�tu�6����x娱s�G��)6�v�g���kb�;����خ~���@��ˋRo���UBfG�7CUm0�E%8�_ouG�����BHɚ6�n��{"U�[cد�i�Q&�d�-<��2 C�yE-<e7�I,���ҧt�!/F�������\pS9���n���U����1)�}"x�0b"5�{�dv��/�H�j�i@a�Is��`����.��oV�8�R����
;(����V�0e�xA��hYb��,~Y+�p�p���$v��`�H��P17��t�zh��++�8K/Ga���@H�v�ExT������5 �4S�G�;MR/�z-�<=V&�v�����5A�a��oA�N����&l��<��O5�5�x��M�}�4t{$���p�>�7=
0�N�D���(Kvsr���{S^��4���ѥ ![���*�@�A��q�<ƚ�[fٲ�����Ѭ)��=�PH��.U!��@%��y5L�{�֢4�|](Y�VHz�1@j@�O'�e�?�i���pNʋ%V�^
��M��n*?�0��}�A4������/J�GƉ#�l�B�X�ܨ��H�g��g���%���(t�ʅH��ȣFS�^(aw|${�J%�J��V�ZV��c�H�<�/�䗎+�*xЯ.��a�2��٘�9l�* �ͻ�塬c���nCp���X7pŷ��
����uً��Y�:}l�w�����J����2v%�`�މJ�َ����5�Y�u�����b��]�] �����"��2��(j�Dz���FUA�Զ��Y��J��g*y�g�������eJ�k6����
��\U�� ��\Z<�����fP'F=��es�Q�����VR��.~�t(�z��R�3A��ٔ{�̗9����Xx��P:cec}�>䂰��hY� �@�[;�p}p��Z����0~㬄�
[����g�<iL����b"ʧQ>�.O��&����%�j��ӎJi. Ң����W1X歏�"�Ӱ��մ����O����gC�)��`�Ğ��VC/�H)�M�mz�=�g�v��~�:&ӏ�ڨxs~��Ĉ��Qi��A�
oQ����H�g·���c����ln�4��H2wq'f��!;a>����Qw౭�v�����t���3�sE�n�M!�,���-�3T,,�l�b���v4%.�s6��a�u ?�3^-���Kp�p���/M�+T���FK�q�7l�� 3n���Y��S��N�z�~��E�ů��ֲR�<�l2�\Ϛ��h�JKw����q��?��>�T#�t-���J�or��_"�a�!�t)� !xj>/�B��%����>ǌw����˅���Y�Hƹ�DkV ����SLA�����x��n`o�}�o�=�.�0�M�Aʼ:哭��g�6��0Vߢ`��8��,�1���hdzlL�}��2n�D~
����]��	Oڒ/w׶����h��Dj@��E�ٗ�љF�+r=������L�s/���d
dO�#��UqQB�%\A�u���d_U:��=�>��\�����qL��Њk����{D�nc+m=���)�o��e�,썂4��ylͼ
'�!t�JQa��,���0�X+V-=�2�΍m���c�������	���	!j[E��Ɣ������*U������ֻ�×�"��(h���4�+���,;뾀sC�*3��ו�'�ǌw�/�e,{m?�l�,�x|���3}=x󍹐 �wQw�׮����)_-��{���.t}��lw�^A��~AOm�Bg(P��G���椲�Q�	Wt��2����h��~�P��>SyA��xn�.� Y�s�f�֚�r��Y�B����^-m�E���]k�y�X��~����v���<�av���.��ue���1�q�+�hZP
�'����� ��:W?�����"�ӈ_��fF?O@n�&�<��#);:�t�,k#��i���p�X:�A\���.�n�H�YA���&�@"pg�D�5Է-hE�����n�P9�rKJZq
�b֩X� %1���m�U��S`l;��t:40��u���0�S&����ҭ�d��z?��{E�qi�\OtM�� ;q�����'Z~F;U���r'�(��P4#�U����s&�����G�V��Ii,�H7�B����
�H�?1�bgS�߹�� ������X��F���}nX}��<a$`̫��� ��#��-�IU����ۍ[	v��j}��wJa�����N��`
<�]\0�h�W�v�m>:�0��F��#m-\`�7�%�aj�<�d(�aw`V��1���fD����L����RHO��Z�+|Xy���XW�+yhe� �bQ�U?�����O��0��X�e�;����+��3�&�Մw��Xi�����O�?@����~� �B�P��7z}�2��cո�N�K������8
��� ,ŵ�{Q'v�����hzzч:�?%��I4��J���F����,��-���w�{��@1�`�s�.��������p�r��O��%A�B4���B�LL��< �A�t���%�s84�m���3~�ހ�J���1@V��
�I��Ԏ����~�	1�J�_�h��f�=Ե�x7h���xlZץ���6���k�h��=���5@�[�����F���*�f('� ���}ӈb���@`!�6��ݿSKn�/�L�3�`��n�rxМ�U�K��B~W	���i�Gz�]P �?U*�$�|��X�G@��Y��:�RS����~|��b�:����������V�<)�X����5� �y�_z�T��"6,�X�%=��1�e��O~}̈��{�hB�W�_9QL������k}���.i��5�G̸� ��n�pwNW(���j}VKV>���_�.h�uc	�>��Ǐ/���s�=b�)�O.G���WK�ey�q�Ȇ֞zX��A�|��WgO����.MG\[ ���?[�/B�PU���%37��2��B?"�]�@p�U���:������ZQb�O�`a�:�����}��`1��ٮ`�?�إ��%��N��r�ؾ��MU���#�Y
�����n���~Ő���;٢�:�/���Y8`b��?,�v�m���f����R��G��B�4'���}2n�Kf�t��#�yo�6H�oG��9t��}���|&$�k�&!� ��, �lG_	T�s
�	_Ǝ���%��<�B����;gt�O�W���Զ��o���œ�,�E�z����Έ�+1㝸�Ķ_�����FT\%�.G0�U,�Ó@v'E'�> �Q�B��?@aMOw�磎 Iǥ&��6�3J����\�Y��)������Y�w&%#�Urj%�EQ��T����T�xX_���@{�ƍ�W�8�;AD�4�ICɿJw9��PÔ��M�V	/.��|�:[(����=���k(H{��V�a��CC]�	���Y:ʲb���
�i���7��׬�ԕs��Ƙ��L~s/N����ZF�yX�
��ij;�.K�K��Nc�7*l��j��Q��hp�K��\d!�U�+��*0{.�*��]*��!�����z���-��[:�u�?�,p'�T'L������l>i�z����jٹ�|�l��47��;�h�*�,m�a��ǵ���B�e�� �%�!�a.ۂ��]<J��Tb����cG�%ߕ'q|zE�:[,��񄾀>'9�	������}f��Wؿj��w�<�B���le%���'j`m8=j8l��e<��M���#�D~c�Ǆ!��3��� ��,|�g]�NF!��ع3R�r�²�!N9�4�uό�9o?ݯr�`�vr���*�h$��/�n����
��M�yKLԚS���!�»�}h�9�yUvz�Б7R�S��x@؂����$���o��J�~t��
e�k$�h��Pm9���<a΢�L���SX���GrK	>�1�P�u!M.;�غ�����>;?3�kz�O���=M ��&�c��+}��%��O^BF��mڄ�w`�hk%��v��"R�����(�P�gAJ0�Nd��8�ʏ;�糘YG�����,�[tU��!�l�؄ϴ�O�o�FWW(P��� Я��aη;W��e|a��	�qQ�l��cO�s����{b���bx=1�N��^�
� ��a���w���u����W���k"�
�}�!����ҧ��&%q@�:#��C���+�q�`��<�T�X�t���2�6z{,��+��.IM��f=�EOr����Q&���8�6�������57�l�x�᧋����/*�;|MY^i;�L����P`�,��.��ҕH�z�+�Q��(�R�_g:R_����K	�.�����Hg/+k4�G��c祩4r3AyY�E3��0Lr/l��0"�RI�Q��A����մi�a��Jb���[��_��s�.J5���=�{ȝ]�1�.� �.�]��$wu�6J�%�͒�nQ �5V4�<���s
��7@��U/�wYwur	�iG`�}0�z�D���Y��mO
����*�Q6.
������Z5�Xd���&wL���n5*B���߁3L�`~/�⿡,��#p+�@���D�G�Q��4����K�	��"bmG��6G��Vr���VG��&iX��/P�O��\#�6=�AJ�[S�(�
JVd��כ�7*LY�h��w��l��tW0wQ*ڔW쐲�yf��-�7^�Y l�O���^C]fms�cq���~'Q�)�[��FF��,��
�L\����>�39g657x��:+k���{�i���7�_�ς�RCx���Z]�O	S�QR�a����WRR5��{P�:�����wz�n=o��.oX���xS���9򎪅�]]�?8�7�X�7�PjN9B3�+UY�Ν��p!�re�	y�*�L��Z-��	��l6��G���:O� @�z:##Js�����	r��3����T��zY��w�o�J��W~��{����*/!�;`	�|?�9������t܁/w�w����G]��K���g��ΆOQc�BǤ5��8�D骧%+<\n¿�WQv̘�G�3e�ߛd��@M_��'�(/Z�p@�	�.2a186q����T���Fi'i���{$_'�z�/�\�?T�B���\�D�(W<�H,iIu�f-��Q�j���D�0���0/Nq�?����'˼�0�D���b��#I�ٵ�H(��g��9��]��t�	�X���8��;>;�:,VY��#cu653�i88�߯+�u<�b���G�@vл�VW��=x�vZIa��H!ݨ�l�k�S�d��j����j"�8B�j�;qPvc8G
D%}A6<�/n�����J>���^�cM!��%ם8m9���6�K�Z��l{t��x�G��u'sp8���K0s��pl�@*��޷"��a���x��y8ɪW���p5���VE�o�hU��;���r�h�&=n媟"�����2<���ܓ$l �y�L?N�iʍhƸ����:Y������M�9��o@��qĠ.55�R�~����\`�S���\s�)̊�r����5����I>�˗�6�61�vB���9aLLT?1�R�����S%"ѩco��-!�f+6��
���~u��ё����C��ș-aכ�8*A��7�#� �:#^��1��Q:�Yېc�mr¥	r�H�P�6u�T��^C��Yn�$t�jr�bǵ�6s�ጯ�����92����3�4��7=.V��#��1�#`#�w��Ȯu�7��Pw�� �����O����4C����_���:
���.�Qy/��������#�	�z������7	:]U�ɱ�]�%Bh�A>�/?֖zV����%P͕����YWez^���~���9�ōRǔ�c���띍�vR2��J���`� ��oĶ��E$���}'C.PtcǄI�6������D3L�\�M�qM��XE4�UnN��
�+�8����yX�]~'�G�v���I]7-�z��6������W��"�/me8����=ޥhh��+�98��-W��s��if��h��Y�O����k$841V��h�xPO��t����]Soΐ�Ԗ����k�p`9�-����O��Ck���9� >���[y_�?���Aͽ�l)��u�l�Y������Lc[�J:
�h��*��z��T�)3�t���`N$-�P�U��v]�䶮���CJ����T���y��޸o�P޼����"�&B/5�CB8q':�bّv��uN��R��M�O���P�#5���2N�^�cW����C�e����]�i��=��fv�	a�Wc��MOa�/.�ݾ��+�Iss~���(���i:���X�=��"1R��� {�;p��"0�k�Y�G�\��b������sM��\��r2'زx;�u���6cH��dZ|�0��jw�jɓ��%��2e�� �u�_\d��"��MG��ԹbΛ�&b�t�@9V
W���9	��<W�u����v�i��b��E��3/��'��藲��y�t�D�	�:����T
8O��F��`[�೿��/����9�����"ITK�A��g'�-P���k<�E]bFo�i��/��p|�tq~�څ܌ߺ�ٍ$v	�L�د���vB�����:u#
8V�RQ�q�Y?0e��w�ʅ�;�y�t�u �}o�r�	���6��^["��h�1�v�ri\� l��D��#��R��}e$���l��(V�P�����N}�m��ڂfQ�x��|�R���t�hm�T�,B_{�,qH��I������>���NyX�����s��+�i2�Xwn��o$���Z��k�¬ʋ����@P�7�,�r������I��Њ!�<�TNΔ�]�Qm��7�re��f��nH��F=s��1�%gP:����{i@E�f��կ�b.JB�9�(.���ȅ��y���ry��C���6�1Z�E�Ʊ�SH�H�ю��|����t��fe+�$.!�1�	��p�ޫ���&,�$/.Bv��5N|!u	���Լ_2Q�9l|l��Di8�m��F��1p��=��������g�o�A��(ݢ	s�����8H������x r!=��p�/Y@%�͒� $�R��Է��4�d[��5�=:j�1���J��J�m-���n�̐��3�+:Q��.�JG$T:�����,|�����g��dZ��A^�b�g]ء?�;�Q��pF�(J�����<�������_kK���8(#S���WX~�V2)��?'������9Orpw�h-�i{�I�t�mU,i<b
#�00,�ÿ/��Ǧ�g���� e��\;\Q�H�WҖ潤��bua~���8��J-W��׮a3�T�P�1~��`��b\JD`���#�saРl�Opj�0�t`U�{��|���K��&?$�ڑ(�ߋ�H����x����Xx1�:��~�f��9<:��Y@S=b]���iy��$��� �婰ع�ۇ1���E���\O���&�dF�����8
���p�ɛ�^��u"~�(�4�R�c�H4���G�.��K�TGQ|�U�@jH�|�i��7զ��R܉/ƫo�i�_J�ޟ���u���|�86n
F&6&ѳ�x�ZT'WB�`[j��,YU�R~�5��;B����'�l�{or䄥���J%,o�-�bX"��1�����I�;���aiI=U�9�emdP��/5��p�m��ς�j_�r�1��!��1z<v�F^�7�s�XӧOS]Qϫ��y`+�s!�쓤R��!���N2�3�,x�@�t��b�I���]dyY���HJ�:��j���/�t8��N�� 
*�c*����OҢZ,����k :ɨ?���1�R�d�������*���7ʠ��h�J���~K ՇWB�և�+<�c�Q=��˔���	yo�x����xSo����!lS��b��S�fY�ڌ��p,�,��$�|�D
k�aB>gB��
�7i�O�� �5C���K'� vi�����ᑳTZ��ע����R���+���k�7�~�ң�.m7�ݳJ����{8����e��At'ʆ!�:3�'�Q;��H^=���y�q�^ϝ���N3�qxW�����
~�!��J����P��!�j![�K��CAV[��X��������V)n�#�����V�3~���m��N�[��.�~��2[�������b�oj�A튐���73�Vrs}<�g�y_H��/Y@ޚ��\��|�gn$��!��;��r^J�3��������#U��60�� TF>��O#`��7>�	�ƽ~.�#�MNvt�Y��5>P$=�6��6U����,�����!��@�[���T��5��5��z��s����w�9DQs����G��v�6�u�z�-�����c��C%p>��R�d-Y �o�)a�2`![]�k+M�&NX)�ĺ�e1"t�� �Q�9&�L�v�H�J�j����ROv�PK�r��7���]�u�o#�� ��:��,~�Gq\^��x���Xe�<�)Q�D#�!�>0Cw���џ��
����~�E�jC�=��3|ֺ#��{��%���K��Vڜ��^��	=��܇?	�sόz�z;0��r]$�ե�W�+%��Y7.����#SV2��,r?Z	H�e�lj�_rK�����n
M���SI����d���/�N�煟쪜�3��37m�^Wfp�3���E�m뗿=�V�V�`4���N!{���0�Z��~.�0	�Bo;։=L�w��Y�m��)=	?w*�k�B��$b̽$�D#����d4�g�$T�JȈ�K��/_\�T�9=���,c
��������Е��Z�yP�]u%��N?w~Oy%*����+��x+:���J֢=G<w��/V'���ߚ2hF�-�!�s�ҿH�"\@~�6�p���+����(9�i�^~@�)�p�;��u�'����ѯ����A�+�H
�`�0���ɥafj����l�|�����w?}~��O��X��*���+���
n�jl	a��׃}�Q��������#�t&�V|6�C]�,V���:;T�)���'�[=+������Vk��c���&?,�=��C�K���}&5��鴩�O��A�G���g�0�V����'U��r���yx^xȗ��x$}w�S7�إ0�������!RĮ���'P�Kom���qZ�_L�*	zTV߀jfʏy�m})c��9��+���^��Ŷ�.�,_����]�/膧���C��$0����@6ƴ�E
��̹)9(��1��ots�Lj?��)RL����J�y��}�Ƅ�dO)>a*�GzWЈ'9�qj����Z!��Y���0J�}\T�{n@�D���}�O���ȯ�w��.�z����`�B��{S�<s�K��j������F]z���o�4�Hٴ1��<ՒJ�?=K�?�Cs0uԡp�`�o��r�WcaJ$�������Iߧ|�����Ǩە���>�	�_uN(uw�8���W�Vi7�m����Ef�����ۼ����NN�`ŀ
����9{Ќ��1c'Xs�`���/�ѫ�.����4�)p�~�;�Œ��h������l�l�t���;7$@�������ۊ�n�sUlǞ�>��TZ���J&��i��SHRL:�e��N���㺍����Q)� ��=H�n-����m��P;_�6GEld&;���@���G-�u�/-q�\�ڱә�������<�i����z-$�0��7�nDq�����Q��4@�Z۔{�쀽f�>Q���{�Cr�ur�=Z�(L��j�6�H��"(��aw��zKM?UCȋNW�hɷ9���k�����C�� }�� �쿴G{�Pߴ�*�t�z������`�X9�j����9~@� 9V>]ީ>%��w|�,jj���i/�����y�K	�4���F*N��H9o��f���G�+޵ʳ��^���s*�ǧ/��N˥_<3�m�4�W �~�,�W�����!�n�:�3�a���%�vjvk�d8+�4fb�Lt�	�r~�]���%D���?�_����d)cߝ���7[�d�n2*�X�.����D��0I�����;+�j#D*���]}α��Z�ڬ7U����o�·�����1RV��Z$�Ǵ��;��%�����ڨ��B<���+ڛ*�p������S�_��+M�?����n��W�O�v�ܨtMۙ *�z�X�1���e�uY ��I�Y���E� sf<ߢ�n�U����c=�%�����*��(���g��ڇ���Ch@��Z��3I�A��m4y��*.���eً�ׄ܄�%XK\�{c���2��?�zR��B��6x�>b�Hɭ�DǪ���K�!�{��I���	�I���&?��%�o�g#���am�S��^K�K�1�
'V3����:�s�ox�Ya�<�6�v�6�#\�ޟ�#�ǖt9g�U��`�hu^sW�=�H��~��rj��6�c^��x�L�K~�=��"rC�L����0�b��py��l}D�>㞟�����&���9�I08�un�:��H������~�ڊ�����dJ�M7<v�껎�/	�ڦ��/|z��+��竈����Ł����� �c���E�W_L\ �;N�]���j�l�����T�a�V���$��2��*3��e|i"}ȟ��O��`�UG���ڧ0��epȞ�O�wJ�9��"�C���@���\��Ws4����'���'Z9{���3Tz�ť��Y�)�c�fՋa�W@����ŉ��k�U�.O�L��.��֜^(���X��3�30|Dt�k���`��	�	�=	�j�2��2P/^�p��/\�$�W���̘N����ꃓK�ɢ�*����V�H)�� z�ه�H``���B�� ��@�Z�M e��N�+-�'���M�'۶IjJ��;s���֣Ɛ�B�3D�@��E�P�ݜϔiB���`�ڦ�fD�F� �B��V���˲�Fx�Y�2���� 7��.UZF�ϑ9���K����qDJ�o�
�׽ow]z�OE�i���j>����A��.h�*1�`��_�|��"�v��k!ƼCK�χ�I�,[&��꾧s0;�wd�H��}HjГHc��c������]>��J�
EtoRIs
�c"�ݒ伳���'1��?�0���~����C��Q���]I��+�nA@#�/�8���AӴ}
��Q`��Dc�X;��?���$�lu�}vwQ\����S:�('�Tb�63$u��0��|6��m��4��ם��"�A��]>����	T����Z�~��F��O���=�����_[�lfo�#�]��!�&�
�/�^�:ދ��T4���Ш�Nƨx	-�o�Tn�;���:"���R6?&�K���/?��9 �s�[L�1О�Nq�wr06~�9���w���T�@�V&%k��*	���k:������$?u$L�:��@/�!���6�����.b5�y������~r|���� `m�!^�w�q�}���������g��O0�c��k15Q�;���D��4�9�AHX�o�o/Oۮ��)�b��1q)&$h|�(1�F���>���CF�E?U���E�2P�A�f�}a?z�,k��|�-i�����G��m:6�.剋ɲ�'����TY�+/�=�)�&m�G� 8T��E�o��3�LZ�3��|0��C��
�v!���# ��rg�.�KqМ�7E${h���7`=�{���4�h����$&��1ξî
����l}������W�<W��	����Ķff�C�e1% DµO�ֱ�?�d���~ak:>�ة��9�Ko�&b�%�l����<�8��MgJ,��l�|�*g^$k5��LYFIs�����4���u�[|ꡙ�@��ߦ�u��JE�ٞ���:�)�DJT`���FS��On�~���%$�kv��1]9}ތd���u��|����]覛�FS�N�SSѽ��&-n���8U(�[ͲM� �8���
�ҥ�����x.<�83��k!����&䨧��gE1����R�7q��Y"%��W����PN�@����3�ڽ�������eT�˖�Z�r�'��'U�k�C����o�V=}z_��l*��ѷ���C� l�r9� �k��&�����X|��fc��4n+ԛq�ڛd�.�R��bܨe'"4 �U��c�m���F+,:QŬ���[M]o4��B?O7����
7��H!&%���ս�[k�x �pNmI7"?�C�2`�R����T0{��'R����%J�*b��z���HFԛ8t}c(���ỏ�}�&��p\.'����[,\�M5@ke��]�I�C5��y���J/Z�<�Z�Y۵��ԛ �i$������q��)�(�j�����S$
�ts��~d�"�Z�h���:-�DR���g��r� wj�V�)�S����~�܀u�m�CA�<�[�	�����AQ�K�|�i{�y�s[yAg���rSz![�f#�@j9[r��U7�&�#�A5��"��|g���۩��z~��:B� ҃_s޼?���A%)�Z�\�46��V��o��oz�Q��]*OK%�?ɚ���$���L��n(�OA&���00g-���w����x�bZ� f@4��n+`I@x� uƺ��=أ8D};�� S>!���hE���8���,!�MUc�XnJ�pU��_�<�����a%m�M4��a�xi��2KL�OX�D��MݑM��|�mJ�Wq�u,�d:�ڛβ�آĽ�HԨ��
���P���0R�⑷Ba����5��=�ZTգX�^؎X@��1�~�%����zz���&�/��byC^TY'0�7������Lu�FE�6�+��ǻ~�k,��W���g^0�w�[�1yU�5!���<i���z�^U��Sw� /��i�c|�q��i�F�3�$��0���]v�_ �N�{�c]PXT���ð���GHi���W��O��!fĘ2��	��ݔڥ����ǧ<-�Ǥ�Z,*z��	s�d3s��
���޽�C�R���<6��Mg�'$������rs'�$�mz,�-�$�7�.I��P�*�&�ce����QT���58zh�p���&��X'sX�'�Nפ6����?&@D�Lʘ��ͮ×�p>ba㒋�L�r�tI.�#���%�VuW#ѷ�E\���?������h!��!�~տ�VPD�y��=��^ʝ6w�xo�������*��g�s���hv���
���]	�G�U�TN|�nB$�������*�����<��Ǿr隭�JH�_�|E�1#�mO� ���#�d��@�ߤǱ|��"�6ŔR�?��+�E�4I���4�<�ݣI��%�ޟ*T���EB�;�a��	������翣��=�'��*�F�d;\�7��nR�{��L�,U�!�^��as�'Z��j���*Uo(O���F�L�j�F�chOF*F/^'y�o�z�!�B8і�~�K!�(Y�;m�0����I���)����(�p+����}@�ܹq��V܉?���)�Yԛ9M	/Z�
�HK�����a�7�!�JX��]���V�5'���&���.?��%F����/O4���p9��Csr8ВVҩ��|y����$��4�8;Ҷ�#�YX�,�#/RUS�\=�B$��k�v<]�?t��\�)������Y�W���,�ZN�V�=iΧ���ؙ��J3�{I����\͍v��(ܙG`C�G^r��"N��
��kjc�8��g��Ȳ0�+�9��t�
uH~u�Fu�L���4�V� ����7g�bP0j_3hHA��;U��눨u��㵥1�# #�w�Z�32�i�:!vx��&����-���C��(D�r�[2gd�� ^��a�Xupn<�Z�x� ��`�E��G�t��
�Dr��*m�<6�l������nh&>�rfF����ջWj��P�`�s��LH���}��/%�/��-ßͮv��5	��7	o���7B�3OtfJ���0��S�"��L��
�?����PN��`<q"^�mF*b�̵h{�L�B���$������x�S�{��,�F�^�К�.���g��qBewkx�S���v$kb��R�K|�BM��@�5M_ǈe�A������-q�1�w�r6�C�}%Zk5�zV?'3���	�ش&_HU��Vd��o��a�!��X�&��M[h� ��5�?�H�B�á����8����Ț�B���=�m�=<�xZ��0;~G΄��{,˼}���]���v����
ʥ�$�3\ކ��0L�kAkY��n{�|R����0I�"5�:#;�v��0%S�J}���rb(g"�W��� ��X↌D��'�%@��6#� %+�T��|��WT@�Ӭa�<[S��Ϡ���V�t=f)���7U��	��P4]�W� wr50[O�ܥǊKL�sכ��m3�(��A���|�3�C�6�Yt�,װVr��+i�C�7�?�ڬ�X�9t�[�'xèjF�����We�4̡�Z�y�,��W?e|�4V�4��}4X�pɷV�t;<s�_[����0���ΘD[7�Z��`�r��yݯ��ºu�]fy-PLJ��;]L�^�:�i�8��'�wa6�Ç�h�W/�>���X�����=FMu.C��S�:�f~�+�e�K��+H�� 8�V��mEs�K��	��4Ő`ҚOt�m��w�6����>��,�[���O��U氎�w���9Q&����r�}��s�;��gl�=�;=����`�*û���ի1h��������H�I��ӥ���0"8�xy����C� �B�[��Qi���?b*e!$E3�MN���]��;Αי�i�F�����5����h\���wm�F/���"��57|"����[uN=���a9�*f�V&�c,�gH������a�Wӌ�M��\�Y�>�]�d'����5��$H��	 ܹ�f����m([4����h��F�SR�~�L��D*<d��X$���:8�mٲP����oe(9_D���b�ml�h�P^۵�%����!�"���怦�m��!A6T�<
���H�BL� �Sg�0a���6���m�٦x�@0�;�/wwA̅;2���τ<�����,�ܑ<��K��<�E�#�m���-�����������fL�KB� C�q�2�Kr�ְ���&jr^��Gn��?�g��3�a1-l� ���P�D[��L7�t��BFjb)��ֈ"f��s��A��D7o�����1|�m�Es�N�-c�պ�s �Z!
���εH/>�cw޼�t�����-x�˚���l��r�����*�"�t�8��$����8�d9��J�NG��qX'�U���*(O�F�t�؟�����H��h]_l$h��j��3l��5}��?�z�z���x%]��̤�����l�w��u2���!���������zhN�^5|�!�F�$@(Y�IC1Ӓ�ĂH_��vj8z��9%�R𿊨��g�9��Qʹ��g[+�#�|vJ���!ңK5��w� e"��h���k��G�U(�����_��N2g�W����7v��#\�%���ܼ��F���G�lm���!�s�bIJm����9���'W�E#�j$�B"��h���ؿ�qZ	9�KܾX�n�~�Έo3�� 7{DW�_�Exg�*T@�d�!|��=����eXv�~b��� �eЛ 'yA������3 2S�rN$#K3Ａũe�:iV>$ô)?�ӒK��2�ԘqM@֥ǸC���`J�-��~xn���[�ό��{����T�S-Y��[y���7뭯S<MX�ÿ�XT����i������ZmV;IiA0�����*^Zع��ł�W!嫗݀�G���w��EK>�@��mAgMF����a����o�~;��	:Ipl+�<�t�_���1fp�K@��\u��&LX��g���W��f�oT�!�M��Z���KϞ߶�J%ʅ�mÓ�ۋ�E=1��1�1f�+�� ��;���Z:�UNL#/^̈[�1d<�I�',��gYr ����2*e?�����|1���G�
i�[A�ĥ�.醐N�1s�*�iN�����5&:�f�Ϊ��)�'2p�����w�0R`sdkyV^;�Z�����H�%g)?h_
��.ĸ��OY0h2������v���c�g��Zj����Z<u��٪���ˤ��1���:�8���r.n�M*�#��X3���΃�pu������o�@�h��N�
��|�y�s��o4��lϰ�Z�D��X���9� ��ݨ^�<+�F�L�e}�y�B_���]�.�Vr�S����Q_�Kȳu�v�h�� <�Q���7���)[Kp}�l��I��'ƞ�A�xЬ�w@�~��!���$�X�X�L\��V�����#{��5�qڒ`Xu5g�I�m����Q�VT@7���I� �Oz�v��؜���h�0:L=c�L��`@İ���&Sv��Z�����$u,���D�N���,�<5C	(�|�Nx���Ox`�f��p@��jc'�X�K7LT�i&�6��Ր1�2��N�?1^KL��X�O8^b"��ʢ~� ��<����L��=��
�5��\��=�4iB����B�s%��O_��~s��/�?D
��,���VȔ�J��W�ĐJ��3~�;�HQ�5�NE�h����0�<���#ѨiEKUǵ+կշw�|jQ8L\[��PSʑ�P�]�"tͱ0��CM����\x�*�ɒ	��
�_-�i+Eඖ�u��P2�5%>P}��)(�ͦzS���KS�S�a��"��b�$��}��-��@�W��'*�%N�4;J���$�*9�UV��g��8�#+_�x��<|�����[yJK�TҿV¯p��a��)`Ć���2ك�'���0����7�wD#J�p�SrX��&�x� �2�7q����Im	:|�A��g���<��'��%"i�o{[��P.�u���������S+���݊G�6k�·e���P�>��$�|5C�Z@�F��uK����>�Or7�s��GJ�Z+�CV4��F�f6��<N$�W s����k ���7Z��*��fOv�����R	��a��|F&Pn�A�C��&���w2�V�9"�{���\R�Ԇ ���鸔�gѼ��g�1$=�N��i179@�zƹ�=��a��ð�kh�)vp�FܑzE�G����H��+�C���-�����wj�}�v�Ѯ��r�`����VǜPU�y_W���_j=�H� ��ep���-j��"�P�|KƄ�)�a�>~B�tHT�*?j����y�3�aI�Ŋ��Y�gɏo�yB���+����CI��pa�|IZ8���S�A]lMl�0P��S���P��?Z��)��|Z�� {R�����kg�+`t��u��He,7+�����+�\Qr�Ť��-�C�WJ��vr��8��OSD��6���J�.���xB<!�%���-��A�R��R�u=6�'q� ��RR�Eǝ�ٸ��e�"�^lk�����<�;Q�x��������lɜꬽ�!4w\��BL&�:~,�S�����K�D�J��QR!n�gXFˑt�[b��)(b|>2�B.[ #���9|Mw�"�����u�x�ǚ��2M&�|��,>DA�����Ѧ�cm�\`O��>f�<� 84thRyLЇԬ&ri+C��H әt`�������P��=4��r������c�a� �#�滓��) 6�dD�em��7�N[�������T_�����-^X�}4瓬^��R�j��_�|1{����1L�)��`b�+�l%;'"��?��,п�aZ�;왁��262�%p��FK���d�(\D�|.61�Bl�̶PY$�����(F�_�K�*�������� @d͵o)ge^�v�-n ��>�AY}�ǆ7��x ���y��%-�Q�Z��U15���C����'F99<���Q����L0\ǎBOU P���?��RU�wo9t��6>�����F���Ƶ|$�`�m$��b�v�f9c���u6� �Dnb��<V1aj��2�d�����.��|"�������|�p�5�D7+/6�����/� ����\��5YIj���?�E5��W�����Z�<�� � g.�.q��1o����8퇕x����8?����氃k��<��3۫0�-=
��D?>���̍�r��5 �r��#5����@t>��7K�hz|hbE!�|�랠�s&<&����޻�a$��#��_/�0�L�I[�/_���%,���^���N�'�F�v�:��A�&�tK��Jrڄ�+(C�֠�%.A]�s��	8-��N��N�]2�h�x�*���j�ڇ?�?��G[o=&$uj�Ђ)�z3�b��]�@�t������5��ְ4�TpkؾA����T�|)�g����q������U�&M3q��_ƞ���YEU�[9}�1��H��=�M��GvB��<]/��q���H�슏��3��o�x1��k�:&�t�h�D�#h
����3��R��BR��j��bռ͊ 5Եz�g��Ѡ���1&/��1%�ONV��z���ʙq�������s���s|�����?"�9Y���ԭ)�28�t.�Ո�h%����&D&w\Q�p#Z�a�Q��@�hfy9[�́
ب��F lq�_������XR�XxЭ�Ƒ�#�ۤ���8I k�>o����-��~}����ޏ���̍�xl8��6�NO��~ C�F2IP��P[�3Հ� ��M��������~38��ݸ�&��?�Y�����6C���t��(ҫ�Ϫ��NJ$-ݖ TC��f���7�E�羲B�牥���?sp�U��G��nUi1��t��sh�7����z�>�Z.���u&\����Z�Q�������P��v1�XS����}��?��k���&�����:�\+r��c_I�j�>��g�Π�Ė$��P�%DI|j���?zYD���U�1>ڥ����W�c? �xQw��J���d�Wy��\U���s�&�^�`�Bv��rX�~CG{φ,�2�DL}�큇=��c��ۛp���k�����8���V^�B���T��F^e���hs�g��0y<��dD����?�2�-�50�圦W���6�E�D?�"p�+�M<�˧����v
�ˍ%���w�/Ԋ�ЏjS�W�g���"|a��q	}�f �y�樤o�j��Ћ{��ej�?��3�
��.A�@��n����5��ش��ڎ5��&e	 p�3���P�r�ؚtNj�2v ��3ԫ+���q�e8M��8ގ��[��Y��R��ؗ���H�.��V7��)!��\.�JlƋ�"q��3���6�6������Ϯ$3�c�u��,����B�H���o��Ҹ��܃��_��l�T7��� ��ˁ�f7��������t	(m%ڗY��;#xK�F\�m��i���b���L�����@��n������^���[�6�V�+��^Z���[��#�� }�O�S��I|X��N	E�9��bH�35���	�7쁵Ρ�̳y^@�_ׅ��T�jXݲb�X�q�8�3���1���a0i8�mB�}i�vq�<>��UZb�b� �$6��?�0}戁\�'�o��aj�6�=k9|����Jh��1�v.	��D��������olY��A�������uk������)���V��z}�mJ�
F�E=&TR0b��o</X�0��"��$WR<W|���êx�ͥ�%L���Ac�4����JP~�\ǵq���΅94������_e�4%��q:t:P�x����א<�����#(] ~Yo���@��"pA�O�~q!�bP���ueYi�H�I��;� <�G��$��:�?0j��Ɛ�Ov+D>(�j��w��*N|vz)7�J+F����b ����ƀ�2�KXSi�.��U��& �4Jn�u���X�,dXN�i�ͲO�G���������ވNZY�v��S�I����,G�8�ߵXۺ������ܐF��"��'�_��]�<�N��z�O5w�J��[s�u�SSi?�6v�j�lv1n�tlghqK^Ƌ��1\z|���[�K���dҋF)�~�f0 �Z8)�����;7����a��sR��#��mV���ɳ�@��I:b�jGu�~;Y�)�Lԝ�EFH�&�/K��́ض�@����`\��X�\�[>AZ���J��$\l��E���P91�"$� -;;����=�ƞ�N�3E�(Hs���Ȁɱ>h���!=��Z�b������bD#�4(��M�L�o��3^@0b�x�bZ+O����C���l��y��M�#L�^��D	�a(U=�h����.Oݕ��e�M��X���9ر���e[���ZQw,(B����1V�y)��`,h��d&���	� 7�X�U�&�?���&�:(�$؏f�:a#��������
���R�~��+�c9b���7���ט]K�9�ƜG~�F\�����Y��#�8��&H�d7���e��f�wbM�%-0�v¥�cTW_=�@{w��ӆq3�����qQ��E�42LP�];st��(��ï�|�8@��MSCl�ɩ�|�A�C�h����P����W�C
I�d�*+�T܄ƌ�)W���w=#�9s8/x9�3��BȆ���O݄ŃFK\P��s�b[AAii���q\ʃ^�<�8�ljG[�J��l��68
F���@�ѿ�Cw2rB���e�>��S�'�_�e���l�y�C�:r9>�C�s_�V�'����ik��ෙ�ߨW
J���uh˰��&��vDj����q���P.B9x�;�(.��~ԧ��l"�?��K��ZWp �#h��M[jBH�s�\����V	$	Z�wsٴ78��.��[Σt��I������������N��ꗿ��2��M0[��Yz�*�1?�)�%D+����p� h�
�OW��b)��S�<�1[�C2��n8��<RhP�`�q��&ߛ�T���*�F��C������9X��b��amO���)�-zѴ������pw,����k��tn����8Q����*���� 3K���rs�
6p铂�Q�A���^���	r=����(@ovsa=��T�R\ʯنCE��>��
#�<Ou43)���`Q�i��z���#=��,�	�-��б����J�{��bIass��"M� Ƙ)��r ��G��Hsx2Z�u�DAd�+�h�*j��7CE4-]�eBԝ�)�� O�d�X��ێ
׽�X��\Af`A�6WƮ씃,pڞ�扃O��
������rt�HhB��$���D����ð`RAw\�d�n!oV:����h�/H���D\��nڥ��ޙ�F"s�V�\��w�,Ў�t�r���IBK��g�Krȳ�(�Vy�i8���4�6�'�K�u}��ce����0��|�C@��lф�c=���ipM­
�>q�G�-�3G�Y�z)z�^��⏂��A�ZcR}T	�ޒ�R�Wfr;��6��g���R�s���'؎���.�N�Q��Q4�o��NC�)��z���/?���#�צ=���AHy��gq��\��cR�m0*	?cb���E���uC��w��Y�w?��uK/�89?8L�N��Kǖ��7J�WAQ�6��B�[�����*�rl~V+�\�;n&�R{Bs�_�!��a{�PF�YY[v'i]N��^6�- �?6:�X�4�$)��Xs�d��UP�p;�3.NI�C�@
�N2s�%��x;2O �࢘��}[�-�?ʯ���n����3d@5��HWZ<V(nw���c;R�TZ����� ��7�H1���a-O=��hl�ɋT�]觌��V6XX�t㉫��id��rO���q�
�BF�g������3P�;Ɉ��ZJ�����譮^�?ڈ�:Z��]�xG���*e �ѷ8�s;��f����a[��N�r��(��-\<��`�9}�U4��/9��������:��	���G�*	,��K��_U�ph�T*
���̖8J�h俪
�C ����`��0[[��$d/F�)�s8�E��!r��T�g \��IA7�M���pſ�C)	5I��)�i;��ָ�C7
� Rͬ��rAcA��m���Q��Vx�a��K+EVLA7Ʈ�6���w�uڝ�c�<�ɸ��[����^��+���l��-_.�(bx\��h�9!�3��'���`=Q�����2�r�e����J�[�^�}[0�Zj9���Y�2
�K}͔4�U��������1TV�a�Z��&�q��bY�`�XA=�d�Shs%�%\�'����A �4� B0_s��,�����ݯ'J�`=i䰫���Kk\���)i\�AZZ�i�UI����/�ڳ)~�4 ��5n��md (4�XW.e���?d�Ք����sy�HܢC�[Df��gE��u9�Ax*̓�*X@--�����*�	��ɦ:ֱ����O��-�y6�=
�m��p�ٞ�u#� �x�h�d������m�q�n1�f$� w?-Q����Ŧk��Cx���=~�&��$�	�<�˔��y�"�Cc��<�����|�x��p�d8�nD����Ll�W"��+�+�!�R�wǈϗW8�uڣ W���nn�z�ddW�����W�gҫQ��>�pj��>��o%�3X5޻����7�`C�>v>�,���������z��)�Z�P��u�Ws�,鷆�`����
�!��=�p	@ڝ��θ_3�<�/E����_qc����l�tD�>zAS�G�P�?h�����w�$��1�|��F���X�Id��eW��YGAbp��4���0���k�qN�H���H�D�OZ�������p<��RY7S����V·x���S�ʲ�\�edf`��f	2"\0�YH�h|�aaX�G��,�J�9 i����MU��F 8��	e�|[ު��\R��0.�	�nk��d8b���s��:��3�kd���l���.�X���O,U2, *n���/�vU[�}�U��-ݵ�x�8@~��[�Z��A�ݼw�دs<��4Wj����>"�U�ױȚɠ4�<4q��`�Β�Q�V����LGG���3����̉6@D}?W�w�W�.�l�p� ��m�ЊaG�g�IS��k�(7����2��-8h��E�ld�6!Vj��[�EE� Ξ���He1I���M��� PU�z��o<9���K��b;+�:6u���~Gh�H�1x"����7�վ��L��1M3Z�.�#�H����N�w��ǮM$���a�C�M��{�w۬=��8���R��%�5�*1��} �
DKh7��*u�}Ke���+�a�W0��Pl�+M�67���/:j��=��|V��\-L�B��Mɡ���)d�Z������ɿ�WJR#k�oQ,녳[5:Vh���,�/�~���i�����5��x��O�%(g,��BO�=b�(0�x��M�wZ-��Öv�J/V	�]����/����s�C٠H���I͜�f��]�Bh*q贈o�׼�R#N����\�7t�X��kp-�:��
Q���r���
,̨	��O��"ξ�N�??��kg���Dk��)�V�^ƿ��� �Q��*�9²�8�H�$�U�c�M���Lx]�	J�!diuP��g����n���e�l�̓�4S��A�n�W�?F���DK}<��v�� y����t�	�_.�����T�uB>L��� N��0ɶrO�:�t��dp���/\Y�L�ކ�)$���j���¸x�z(���z���z?e��|'��������D��7�W {<�� ����'���7��Qr���
����븻�y�Q6�_�!�k	/�g�:z�nb�[�W!5�p������q��u���� D$DaO�%�.���eF��`7\�X�0�މ����:�x�;�|<�ɠ�sN	~�X^��b��N�M���dO��+�9��{#�x�fήio=�_ju������nD�	ـ�V�Ɵ&�}�;�l,�޼*GRu���(f�G}�np=�J��B��3��h�mZ��K��k���YX�؅��&ڰ�wɹp�����%�Ľ4;h5*��c�:v�2�������v%v�D�|!h�U�p���)ze��1��v�rX�{S>x�&8]��ڡ�����$?��+ǸmU[#�Rq�b����XqPI�<�G�D>˕��E_l�7R<�D����إ����e��4��GI��h�(7�ʑL�9�k�b�+�;
��>2��OD+�ܐ$
V	�bP�WaC��;o/�1=A����,�-HM������!3U� ^L���aw�6h�k[��^[�1k�\����uιR�趞��:q�6g��%�Qu��|A̓����R�"����#�
lbr4�(^�ǽ �,�g�j`.+�y�6T9J���#�-D�\���읣csw��H�*i���ޒ��ig{k�S$�MM� �lz�'�U]�b#;]����8���QM�Z+�A�Cـ��SyD�u����e�#���?���'\!Fez-LU(2��{u���[����:(}>�ߝ����nuv�_¡��6�ʟ�U��Src{A(c�I|e�[��g�V�[�xKŻ�mxS����uǂO+`�Sv�Y�뢛=�D���b'K��������t&������|z����I���ۊHlYL-Ki@��:�����e3���K�C( �Mpޙ/�/��d��I�2���&�e�*����-?q�{�X���j1�R�[W8�o�+�n|��6z�������q;�K�+�
����))��(�S`u|�g%��7ξS�#�>��|��s�%y%`!�Q�&��:!�vju���4�{ʉ�<l��; 0�.�i�B��{��X�3vM�Թ��D>3�⪮Ir8��Ib�.�b���+E��lm¦Y28�%'�Ū&'��˛ц]EK�(�ʵȧ©ɘ�K�i�0}j�a}Z�4L�7L�V?ܶȦ���(�/�<x�<�����{�`���%Ƙ��GD Z�2*�y* �{�5����B�I����:A����&�'��D��!3�F�!	������E��rlR/ \c��İ�m��D)��?�����9?�
凂r���?BXe��h���,R�CFhR�	髹.K��ߓD�:?�4���M{d�|���t�
h��\"<�,<�0�  ~�K��N�	���L۞$C+Q��N �Д�h�O[����31�ː3��w��t��j��
@k�Y0a4a1E���h��xώ��d��b�Z%_K�4�z<�Ors1N�k�A����W ��&�W�aR���̔��r嵨 �(����n��Y��|dft.�ޘ| �`�ƾkJ� �
:K�/�8�J��o)unR�At�W� �*C6 ����֐_� oWÃ~�����=i{��k���q �a�H�&׳��Y<xw�ZS2L��!�ƾ�>��HQ��S�����M�΢�r[V5�2�G�P�u�z�h"F�GTi���<�5([���}0��(�a����s����p��0W@@O��)T��r���;�;�sy{:�:$}��ݮn9�������D�p"V�c�8��z�jj��,J�"��q
y�P�d���KYt59@���M^�$vA�}m�MaFq��
�O�:���]Ҭ
P�	���=�爯�5�f2��"l�/ܿ��C��XCݪ�숭b:`睵Y)D�H�>�<M�֝9أ��vk�{l.O��`Wk������qI�mr���w$�Ƴ B��f?�$_��� ߹\>���>�հ���ab��pqjʢ��(�3w�YK�������ƶ*$U7\a���֦?-fpg���s4t6�oj��T���<����X�H�iX��>٬ҍL�Y�xC;t��Ke��o�7��.O��I�]=6۽g�������0q�ݪ'���������f�B�&U&��t�D��r�M�+� �}ީ��m}�x���![�� 喛�"^�#�^���H����7�%QӍS��͇�.Ј;3�c2O�Y��y~ئ�I���NBd��m'j�[6�&o�/FޡQP	\�M62K��z	�$g��:��3]�1�.����+!��ë���pX���xT���r�^�[`w��U(����["�	����"XW��σ��d������-H��V�M����:�Sɺ������"��l-�d�DT]�&9���;�H�o-�RrI'��J�KHN�\n}9��g����~sH�����)�2ē^�N�nEj���G�[ &X���?�SZ�ȿ~�hi���`�'��Ѯ��-��Q?@�ssĀS8�A/)d����˦܁�9F�׹\|@�{.�ɲ��q�p�}<��
�����G�D��u���{��Iz����R=x�/���ڰ�g'����4�㖼z0�AjpO�,����?時k�[�� =���F�Q��M�t�_�k�e'~>h2��I�;������^��P��n��z!?w�<�(��"�w6�À5}��v����4eXw����7#b &|B�F�vaZ��YW�X��ZM<~��|�L�L[] ���Ȅ������<�z�0�.�&�I �
W�Qw����\��D�}^t������C4���ZF��.� �-����b��za���<�ڠ�Tuo�80�m]I �#[�a<�����WC��`-#=�S�������iV{{:�D�E�@��Q�j���qT��#�w�xya��&F*E6�
D���r	_�<�l$t�2��S�Ė�xka�SM����Ҷ8K���0U]dĐI�7�"m��K �Y�:�j*����=\�%C�E����rů�
��J��n��b�T	�iH}���]1��W�^��C	q�)�,aT�;���3�N�Y��!���#9�ġ�R�	Z��2|ti��E���>�Ԅ���E �L�����~l9up������^�ADԏ�ġ�F
J���ǄN�B��.�M����a�=.�̷�A/.����0yw�4��	��̢�����o|*>=�-��]`q~Swc�vf��鵖�:g�B�l��HQ�(o��;�w����oW�t�.i�j5'��ݻ��V ��+���� �t�[:��0���Tj$_ky�N���3W�ҏO�³�n����r%��n׭\/���S�z���-��]�0zr��-e�m���(�S
ys�5S��u��u.���+<B��e*�f
��|T��i!�P�C�Vx �;H����m{"�H��j�6�]�eɓ�G��ϑ���̱�D�����S7�W)�$��!���t����ֿț~��D�a;�&tw���M�%x��h�T�����[W^wu�N�i�v�q��^��\7g��->iqB�Glk�/J��.�H$`�.g����n��m�/!VEU?XMAlzL��+����}@���kz{{[�Y)�5��H;��ĵ�����e�C5�3m��$o�D\��#y	����}��sxBa�4���bmX)
���m!���&�[����Z9+L�9[�^�9h��4�(�̤��p�`�'�'��h�5Rm�kTc����oS���?ش���H�z��y|m�=�V�B
 I�u���d���k��?��Ƣ ױ�$
���7JHʆ9J'S�J�7�ۯ#��J�\�,��hr�bz�x�H�R��d�%s|���n����zs����C�Á��7�9��H���o��T�F�놈x^��A@���3�{�Q�q*�q��}��'F����ۧ�w�_E�*X�����P",��B'���*Qf�z���u�_�8�a�i��R��#��&�fϴk�m_K�,μ[��$a�D+�k��@�yL���֑�[�A#_�p�۷Á�/G�Dl4��\��&Z������$̚��(.�cS�w���#>i�
�2�Vt���FB[�(~*��X����������ZBo�h�+@�Hjt��;tT�}�8���;�ȵ��ś"��E���
���4F�I�F�:���",���l���#&�|DXTPW����!^O��q�Ё=T!(��U00N9C��&�3s�����[��u��8�O�T��
�)9�ͫYĦ<��ӯ���8{�|O:���g��[�Dx�F��<���v�#ba"���dc�P�~O��w0�y�����M���6�ɺx@�P�;w�mD�m=׆>��ҕ꼟����Ն(�
��.|���q��R�Gu��d4}���vH����,��{^�`>$���b��M��Ei$���5�'�� �W:{P1fl��j4��N��380��ּ ٟt�Uϡ�L>���/`RV0pϚ}\�Ќ`������sG���P�����N���d���so߳>>?G|�,,����H`�ν�U���dPA�h5q��~	\�\dr�j��l��oѰ|�f��"��E���ǝ��a�����a��ɀ*� �f�\LN����I�0�����Hk�LS�+�\q6>
a_�m����}ݲ��f3��[�Jxf��C��p�:�I��n�	�5�h~/�H�ѥq�#��h��n�@��_(Jf�@ �V�jH���Koh��;��]�3�<��)�������Q���ZlT���]�G,�z�!�}���Rn�� �)N/����J3����`RWլC��f�қ�j��`*37sO��Ӏ��~}�& ��M��Y��_I�Y]^e�gs��-ޖ�	��v4�YPX��*t��a���.�v6<�a�dR��cuŮ��vψp*ň��76�#�5K	\��\�)�;&���>��<�),���o"�Ǐ
�K��__���I^i�:�
�Nw\2�wS<T��|v��1���L!��cJ|GuI�[l�^��,Ө��W����io�3���/=4xe�S������PXN�`7?�����ǃ�	�.�~Â`����A�d�8�(v�|�4_e��E�V�!�^x�jM�&*'���;���H>rb#M�Q2y�����51�`IJ�Yx�u1�)fX�~���2�ܓ�g��3N ø���~�}e���w{^z��D�h�T'��M?���(��9k�q��y1��&��<��s����EU�y�A�>:ǒ{ih� ���;�·�J�@�E����l�Q*u $D��C�O������X�o{��1�1�&q�n��^]��m���Z8G���,T~`C��#B&R"[��e��7��<�4qѳ�]j�V>0}u���+JH��Yh懪�o!ͷ�k��k6�?P�.�E���"���!��
<(��gE�,)&��slдA焌�gS��c_����Uzbܬ|��]S'�&������b�pG�υp���M�8�F4��!3*yN�r0[�q�ۂ��^?Z��H�"���-��c5�Y���2xȓN�\�)��O�(�Eu��VȦ˵��-�Y��*�N��Q<�K{F�zs�ž�H��� ('�ѡ�4o͘+^��/�!jci��w��uS�ޑ���2Cd�2�	����'�VOD�v$a��V�վr�#�]%�hQw5��ݺz���~=��?/G�����kz�p��>[���j���T]��]Ơ-��ծ��r�L[W-T�.�Δ`��|�te"���7q
�CȖpL�7�W'w�R
E{�qU��:�l� Kg��qP-o�G�ghu�y~�J�)��V��%�}]��-�|jְ�f��|G���z�B]צf�����S�� �6M+7�tU�֬�a����w#���Oe�����4�1��x`<Tc��������h���ꏙ�}�"���&yb�O�
�<��*�.�d����:�uh��ĉ��<.��G���V�*F��FK��b%�Ԫ�p����+��B]�bԭSY ����fE���F�V�7Z#l�VF�=40��;�q�;��m!���f�n��s�y!����o�QY��q�Ht4W���OT�+�5�?�U�(]�ڃ7X$�#:�T��@�ó�DH��I�Zi��+H�����	��Ja�_]�_�h�^4�n��;�k�����C��|[�Fj@E}�u,(Gߨ��:5�f��sZ��4E"��'^I�
��0f���Is�'�E����2'�<�u���n�8��^ILi���������U��(I6���n+c^O_�t�0�af����f�����/�-/X��}<�8�!�F�Z*����N��u�4%��\P���� ��1����f�!��v[�EAL���������f�`%J�����P`���i�������i=�>+�<��qn� Β��
pjɜ��F�h9D���E���g�m�[TZa]���hu�N��
>��\���gq�ƶ������Z�süs��$=�Iq|�9Q� 뙪����_(�g&:{?h��˒�[�qC�N[j�@&'�3wt���I�������+�u����V��믟K����D�K��\��������Ǩ�dE�-�Z��"Ӗ��ML�dnFgn� n�+��ǆ�����S|8�i�B����`��D}��ye�2DR��gj�o�ȲIA�����Z5�a�,��0�T��M>���I�ٓ�g�t�y����+I��Ňk���:�c��G.W+��^]IkW���zR/P��b�چB�n��v�J%��Kޒ���ڔ�{��Lc�:	���wQ�gU�6�)iΉ���c�+0�~2�%�Ka�8ifSuةG �"A>F��H�߸�ڴ�!�B~���D�t4h1ͥ^��W������7s,/<�?&6y��q�ȓ������o_�������˛_�v	�|ށ�/���M�f����M�P��w$m���
;����e-�Ϊ�͚���v���*�놀Xr0+O�[�YM�@�r��p�M�\u2R�|���W�S��2�)�;��U�)���D�G��^ї��g��1)~R�Cؿp㮗R�Ӓ2��Wz�����⚲g0ci�"�v�ĝ
bxO��l����[�d��y��T8�l�@=5����L�eq`��J߰<>]�S�Ա`v��1�D2��"E��oa����ʡ�l�@��泡x>��/ɂ�҉�˧I�&q,��nh8�'����4�1����U�rG!C�sUmd���X]��BK��,iZ�qC5��3+��;�Ӂ�v_�@��"��S|w]>��M��&5F�c	�a�B�0{2*���m���C�yR�M(^1��� �|������rQƓ*��;K��&�^�
����e{z�9���u��|��4�JG�w��X�"_�����a�c�Ҡ�2���;��#Q�\�h�/�ĵ�i#��K<׵m�@Ӻ�Bqx���p.8�s�Zל�%�#�Q®�xU�G���*n�x�6x�0�������);�q�������vOp��B�]5�3_�:w�5�h��b[7��M	���7=qB�Ϟ�c��U� A�h�<�Oj���#�'�
5�,���Fe�*8��Z��7q��@?��L���xq����5t�+ֿ�� ��g�I~v��t�v�i?����$Fo����Fa�"���S�3��������o"�g+S����&�/B����`���!��tu� {�tG����]�Kʟ���R$�&׾��C��܀�ު��"گ~_��&�C//ni{෇�����L���.��,���J!9�O�~΍�ޝ�k����
(�\���s���ua�\RC�0���t4�m�������6[B�wTȃ���ʀ#9�ψv٦4�����^��F\��{� �𲊯0�n	���BGp�	����0�|�/�S�\�MKS���^Kn�+�!$U[xrVZ��1E�ߒi��� �4/�f��Ր��ݩGKm{���ٜe�����7�7wzb�d5�-�b:W�Aw08����s�����enO�b�� ��J�N��T�L}C!�Mh�aZm>.V"��:dF�wK�7"i�̨;ud���N�8�I�-�9����8�l��Q����� �}(�)@lu��q�F�YD�Bf��I�o2 �u=8G"�Χʔ?�o\�Bk����o�����#�a;H�Ǘ��D=��7C7�Xg�)�r]���$v�.}\�~0��3���H�6w�۬<�1�oļ'$�����ô�1�?	�)x!���F�Z����%�$�c<�0�oNt)mr2�� �W�ק��6�o�rG"e�D�j�����
�������l���'Nܯs��,�`�jն{�|֝p��N�FS�h�2����C���5��h�����ا�7U���#0v�c�U\ֻ��X_�m[O����?�@H��t���P��I�+3v�VR�ɀ;��r\1@,���[\`��5� h��B{D�����2I{2$�|�.�	����vM�;���LM��W��:��=��he��7�;����8��6b���0V�o���r�xT��/J�Q���1z�Ӷ{��dzl*�f�kU�`�	_n�}��H��l4ؔ���@�JA��m�-��7���~	�����'^��`|	V<�:�dȡ�Vp>�Yސc"�6���s��Y9�h��f'ǆ�nL'^�Ѧ�-�dG������o�!�Pje�\������2 ���4٠_ 6�|�2�)c[�Zxinۂ����m�Gl��i��W�/��\w�L힢6l���߳ĸ��ⰘP�lh��ym��r@G_6�Ѝv������
9D����ȿv����J��Y�K}@@8	�2Sy���$16���J�>��ߺ�AU}$�M�Q�������O�Q;���!ox/ہ�q֓�S4(�Ě�[����3%q�B��~7X�氤�-���ﮁ�!�+jj��4QX\�c
Q���ȣjh���ʹ����f\�bUK��ywn�lFljp��L�A�������#�u�͒��/�lH��Ϊi���eǦ�A��Tg��=56]��������۟�K^��_����g�_>�����Nѡ(8��W��NQ�{�W��� \h�����	[�Ը%�Io����He�I{j����P�$5���;��J̔��v�"��/�
Q ��i�9�g`a��!�b��ǋ�����$'��Z
�,����X�2o�\o.v=����_O##x�|�sPC'��u����p��X�p�R��BVu��.ɟt	ke�/���0>CRM��s�Z:>��������;�y�����mx:H�,�<?�B��,�ބ�&��m��P<V�����!������faH��|�)��a��X�؄=�����1��Q��HN·���sKI��@�~�=��/x�Jw�O7��J�M9��Oz�?���t#TT���,?.�ؔ_��q�I��£�j��p��^���&�(���U�j)3e�o����!(B�Q���s��G�-`�'-��`����WD0WK���^d�6��y��Ġȕ�;=���H��BKFʹ����x݇_z4�<G}_W�sPv%z:�Ê[���A��5���ɡ�jP�
a��pۂ�M�-��Y�\��1rO�8k��x�Ռ�S��{e�E��	�O9=�T�}��l ��cC��hzh�h�߻K���]wkT�~�� 0�o��h�j
c�Ps�nZD՘ .e��0n�G���gO��}8�dK�x�Y�f�`!����gШ�'=��w��:��ù���SV��Di�̵�mV� �&�R�G�M�\Y��K��K���6jp���Z�յd�B��Hg� W�i����/�q��{�WG�?q���������`��§-h(3w;�6zS:�����
-�,@�����U,tݭ��X)��>ȳB *,�S�{�q��B�ҵ}�/Ԙ���r�0*9�g#��`��6��1�F|뱱���xz���|�Q�n�� 2AâB#����A�uY���F�"of;,�����mE��*����Y�A:���_[�9��B�U�\p`A��iV��~��2���[V#E�_g�.�+s�鷸�lHIu-x��\�r��d�q���1\�N�U<*7?y��Li#�o��b�����bmG�	$V�Y'�և��A��y��(�� ݋��s�S��zyO��@6WaV�)��B	)���2hr��^&S���i�� aX����}�+��QM|g���P���&>M�e�k��]�m����2뒘e_�;�`�8�a�"� �JQ?�Kt�b"����o��T���q�͏a��6&P�4/�T���0	�|q˙Q+���#�6җK�\)���1�&��zr�%myRl�+8�E=�e""S�=�ޙ.�F��e��"�:+���_���	Q|�]��?N'�4���v��cG�βŜ�����,�9�
���58I��h�>�	��|n��]��!㴟����b߱u�hߏ��	���暷|~'&%_Л;" K��$���q1N�ބ/X��	*��4�#!B�D�@[B�t��H�{p4EC�ih�y�֣"�/��~�;r&_=IQb�1�����~��JoQ@��ʰ��_�6�||E$�D���%��{h��w͕P�N���c�x�3c�z�K����he�/C�$�d�LJ��C��E��)I1��Iw\"�>(s� ���ԭ����g�QA{�^��H�<����e��P̐
�P��b���?Ԓ8w�ep9�}o�~4WC�ed�h�u����KR/��ר��P������\�Ï��:y��[�l����k߻���v="�ł�$��"fg,�t�a���D},��сX�Z�9�(�PT��A��cw�p���!&��k�~ka�'�0�����q�\]SH���`<�� ʈ�P��cW��B���%l##�dE�p^��36r0+L�m�x��ċ��}��{� ��Dǎ��7⸡�nMR��4��nT�� ې�݊��ZGy��뗻T�w#@���̇��rPw��0�iȰ8-3z�-�min����/���<G]�����"<�#��Ӈ}�i:��,�G��;gL!��kx*��BE�dpni�t�m)N��V^�������^Go�8�=-�؉W�m��鐢1<P�����\pb{`Q�̒�St�@��@�
�¼��|&��v�o�!5i�t<2�e�FF�֌��P����b�H�g�f�Ih[�x8�L�7��H�Ϛ`�&3�7>iW>�q��7��gK������*ɫtw�T��6�e�m�|�($֫�VV$=��\=�-oQ�����a�Y��X��s^�q��U�D���\�l�xz��NA����]W>2@8`"��3XV������}��\̇��uw��4d�e ���7�֏�=��H)>�c�\a5�y�b���O�t	,�*iE3����!Pz����sO5���čAp)���O�ڎ�VC� b>�71l��,���Ĺb�d�pb�)#g�P�%7�db9�G��<&\&��&�I���~�l%ɣo�����*�q���J%)�4�Ԑ�k�I�>�B~f
[z�y��v�`�E(@o)�߷	�2l|�w�&i�E�B�t┯{ΣŕS%H�خ�fU���K�y��K�4��^"!;Z.�c�r��V 5(�|�����3&x
���o�s��<X�6�JB�J4���伎S�J^��x��~��6�4��̅��8�E{g�́��eo���%f�K��Y�j����˘�۴c��$�Ѹ1�W���3�`h��:��}d�kW���F�Ҷ�3��4�Ec�t���n��?-��`�oΘŲv�dI��W-A�9��?����������è�����)oOlIJ��4�����<f���u�o ����P��D�; ��	X�T��v�6G6�눸�����Iqa^�P���#��5�NU�o�l="*SXL�4O�!%���
E�L>�Q\�m�mܛ'Y��s�TU ��a;����w�ϥ�W��J�������֏��p�>��R����>pӗһ+��	�k/^<��@b���'CJ������E6!JE=��t�8��0nM�)���9˵_B�x=y��c�;e�_@	��W��.�c�О��ޟXmn݊�zZ���H&R]�a>0�����u�
边æß4�x�tJJ&��
;l �5@�QJm��	��!�:�.ԭr㣤P��%,9C�E�ԝ��#����r��%��� ���Y�5��	Ա5ILq���-C[�BO��x5�|�x|����M�ͻ�.��"���u���ĩ�S�����cpy��_,�r6����w�=I���x8�oqu��Hw���h���v�<M0���įʔ�Ӳu��k�ݝr����J8/�%&i�R��,��-!ٷ�m\�;���!����=?t�4s�ÄM�p��d.,?�����f������TGI����l����=�#&�+}Ǽjm�N���$���M��;Ιd��֛�w+~o{v��0m?�]7�esƙ�i�[���ݸ������c�4����6]���mY,a�u���O��UD*ŊcJ�8��<�6��X�*Gi{�¥{T1��>�Xr�銯�h�X'�����+ F�	�	D(��]�r��X�1A��![M�2B�XP�c�����;���6�&�����Sֹ�T|�7��M��!���qx��}���*1L�� ���m��WU�*�U�a\o5��W��ܓ3� ��T,\��Ew��痨�L������c��ΐ���1g���YAqË���T�1��@�zQ?K��J)���:�µ��d����B�����K �B����uƖ�S��=�`���F��]Х��Lh]�[P޿d��&�Z��~�[H�H\t���U���������H��Q��'�D��P=c�n	���l_�����q>�:���3���[����j�%���4bG�3`a���!%������|�}�y,2������q����L�T���-A$�d�%�����l[/�wٰ�i}?��N��+�Z�_�J	B%z��y8m��	jc�. �������QX�]�e`�]��@88�	Iq���R5X�5g��/��T</��KXCDCn4��GQ�f=#����+O�l�ª��Q}��	A\1 -~[�xҮ������,�;3$q�����}�x�eJ�R��i~;W4U-��1���b��F�E��PX��*�+z`B չ��p�;替-�U_W5�1�%��ZG��]qy�3W8ݱ+T}8�kG+���%�|.#Y�T�C�(*���ތ����er���H�`�`��t�k���^=��r(��N*��g��ޤ�P��9u���9�
�ί��
�F]	��`�n̩'+d9�F�,)�]������P�����V��8������2��]:��PŻ����㋪n���-�W�j��u,��ѩej���9K�*ݜ�+�7�m�����٘^����}@׶d��.,xwC��]�Ob�Kf�d����J��ћ(�8�a����bAO�)���l���j��@a���� I�%�&/��b�� Л�H2�^��EJ�p�d�M����(��ҁ �X�Ø�c݄�+S�awei�T��u��Q�QO�9�Y��s��`��5�0D(�ˬ�0��籣I|ëkx<o';��`T�1*��Cq�!�{b�����͉�o�?C�B"�x=�lHn��(��f �2&
,cu�M�� �G-}�;�|���PO(e=:b+�ҥP{w�́�}֒��t�M�-%�,�����}�o���kFAd|����TNZ��l�x�`�.����#�V�JE�J����b��Y�Zp�����6�oޛFJ��t�0�p�y�ŇW�"�H&���\_�3(���(�@y!ߕ���~Uw�y�.�c|2(��'ɻ+ٛ7�<
]����tGu[}܎��e�n�,����z�@��ݟ�X*u��A䵯�t<�g/dB����o�8Rm~�t��)�����8��F�(����#�.'t�P2�i0��ڒ����ÞJ��*[V�d4��EL�ڼH���9ܻƽw�^g�ܭ`���:�&X�L�c!���rt���|�VO^�
�#ה"/�x+o��@^����	��3��#F����!�� ���cRQ�;����8�*Ϗn���N�5z�����BrVaG>g.^���m,ˠ�4���u�rEsƅ�6�mZ�N��$4��?�����|�LH�S3�)� O�aj���=UK�^�L��{����5��Qo��+�6b	姖������S����P�D���Ԋ���	��8"�'�c��~	�iÀ��U��\����~=���m^��B��ڐ��):����w<U��3���&�쿮B�J� b�>Ɔ<����a
�ٿ$��3�bF�M���f�j�]�����\�Ҽ�]p�~�]g}*�)� 55Ƣ��'~Ps��,��]��蚼.��sNò8([��ؖ��˜L��H0fr�9Q!"����Ú�����~M<V��tQRE��{��Ny+ݮ~_o��o.�F�\/����X���S�cV�R�d�X�8S�����iOqǰ��°I��6 ������|����
����bA��"�S����-�l|DN�x5�WW�#��OȞ�v�-�~�ˢ���w��"��0�en�}��=��g�LC�-S�Kn��(�ݗ�&m�t˿��+E�^x��,e�)�ƥ���������ֆ��Y��-��-�.xO��<��^��Gը�8w�N9�[�WA���ܩ�	f�g$A`�A o�*�M3�A_�F��S�/��R�Gص�A�u�~U��lX67&{�$����K���Չ4��(�FO�e����0԰��ثh�KԫK��9�5�;���,�� [R,�#�%�,������I����ղ�*bk���Pi;|&z�sނ�T3�<�7o�Q3�<��4�����GlH3K�|�0WӋ��t6�iG�pD�sVR��6�8N|���;בe��&� .���ym"��768�u�6K�����o[��|�G3��8�{ZӫS�A"G&w���&hH��<^&�̋؞��r�\�ٽ�sBu�̗w��uDbc��3ڱ,�P@7�W����%$t���M���L�����"�1ؔ1Y�"�C���7	�w��� �V�,���rF<�|�P�o_Ԧ�ň3}��]�>����[ݲ;��-p\�J�[��-�6L�v�{! �)��Wόމ�_|����S�N�H��ƈ�p������f�鈋A��7p���p���ld�$���ȫ6'�5&��K�6��1�D�2��ɇ�!H�b��a�N���)D�>=w���?�d��ӳu<VDZ�3���~x���>�"������7G�H��r���\��:��9e���8�9��A���i��	����V0�۸�Vؾ�]�R ��~.]����e�!3"���E^��8VD��0��,�����=XV)�o N�vgA�Z��Ӑլ4�z�g��Ƙ�(�;�-L 
�S�I�����C��KR���v�[��ڜ����*j��$��<�7�_��N�l�W����p�����v��V0�F}���I�ۖ�>pI�� |{���u �Ԑ�g���lI�k+D��7"�u:�d�4�/ꫴ����^���̜r�6؟,BSf�ф�Z�J�u�/=ڷ ������ɣ�H�dxW	�u��y.E���{�P��mUE�V Y���g�P`���߉�C!�`�(�ɻ�u��{ܓ���!Դj��q���;�<�[� s���W��"���R�\`���ҞXm�5nY���
��y�+0�AMp�$w��$S�d�����n�,���}�9�}�"�Czh��ğ�_M �W���f#�đ��?\�­<���g'�,F�2Lf�H����Ld�x@lK�-F�G84 ��i�f#�-&�>�k�GX[��7�Z���~N��1AvT�'�8�l��P���!ʟ��c���~�f������% �r?8�k(*;��r庨c��F�Ml�c��A"��X(�[@�+������n8 f?z���A�5/��5�n����k����hjFz)Vx�lW.K��1��,k�Ɣ��Bj���%}Ͽd�=�~���?�xw��\�k���ѿ���!��v��6��׍��:d��e�:@2_�^��u�!ؗ�V	N�kq��./CE�dσ`w�yI��K�XX��S��N�sxH"��P~���w�3&)"ɍ�5���w@�t#	�E���K��Q-i����QL]�[��i�����������+ػ?
b��7�}.PA�����_�i���Fy���#���i�&;&��~�ϝF΅%�f.uwҟ�i�����'���g];׾�őߚZA>�����-��y/�q\��ّ��6�$�z=.�����K"Yuύ�(��O����´8�@T:I"�3��1�_b��"�b�~D M��;�5�s~0�e_^@>��vd���쏽bC���pJz�p���L�S��i@1��3Ӹb�*���pS�^9������f;UZ?���K��2���l�2��}���&�'bt�$i��+����m�����x�r�}�x��K���K�]J�K��_u&�,��[^*&���|=�����;]�X�Rd��̌_
�/P��k���V}�`��n�/�����h�F�#70��Q�Q+SJ�@+�T���`(�k$vG�^:�r\Y6E����u$���L���Y���7K�=��J#sQ��֝ܫR���~�	�H���z�Ʉ���{%W�>��ǳ��^� kR��� 7T�O�#Ga���+C	��qN.�:�d�	8��lyB�O���;�Sq�ql�E��/�
�N4�"��h&ֵv�����=�ŀ̓ԫ��x?8�|d����d,�� 
J��7*�HS���k# j�Y�錴|�b��y�b8�f
�����B�_Oh�!���.�������0oEy�I8���#Qv@�ZG�t-i�ɰz�S���:��vI9�ZR�(sk�� �^��V��B)��%H@h�g^�H@g8C̆������R��1U"|O��pZ_�<�2=�芞%�#���%%I���x-�6��.���֋�M>�OM��4�����6bٌS�S_������	�|S���/�r��	-@�-��-��+�R2�e���S�Zj3���0�J��Ȇ���I�[�\�:3�����x/۝�!��<N�,����,�����h` ŀՔ�A'�M���6ݜ:�=��wP��ф�"��=Ϊ`����o`Ӽ�&�A
qm,�W�O�������� ��>�l�ːgL+n���^�ܘlShDa�&�QsO�ց����ḧ�dcZ�:�
r`����-�U� p72K
���@9sL]L��+	�n�E�9�����a&8��<gk�=�!��{(�d�發�JT���c!/%���[q�����f$)m�[XM�Q�*��/z/��y�	'�|)��U:R��`�Ux�W/J�9!Br�
k~Z �-��lf��X�
x��b���VeO���|�XJ����4؄���^a���ߊ�Qo^�.v�NS��fW��(��6a
�~��Ƕ���ɐ��T]��z��\�J{���+� �+I��m�e����C�V�kP��,�mk�5�(`��t3��WQ�u���@�J�~�M�E%$�o�s .n�.�������O�1#����Z�*� lB�C��do���g�w(&�!v�Gc��tE��G�F�׼�)Z�g;+G�O���O��0>��,#�Y���	�l��Z�X�y��Q5DI��e�=�G�X	t���Ϧ�6B�0����G%q�(u�h���+�+'o�$��fe����_�iTY��.i����i��_ߚv� ���M�������{ַ��^3� ��������o��6��+�,�gH˝2t�DKP���ؤ��u�Ɩ-9�h���Up��LRY��{Lb���
��g/��������-�.�DϢ=#W��z8�N���pg��3�#���Ȋ�	F�Z{�aY��Ӻ��&�i�4�\���ߓYÐ�Jacs���c��_i�ʂ�Z�@,ۍQ4��\o�#Ef�hm		&���Y����R-�g�Ȁ]�z$o/�Y�N����u����~�����ײ1
*���u��3�E�����>�@q{"�n:oڊqtq4�_�X�(�Pǈ+"�~i�`�Gv�Ux�8m��0V,�ݞ�j�2���H��_$4�����{Pڕ~�C9���h����yq��Oc�i�F}��_jW�ҴaL��f�?�NS%��*�[���5Q�}TƉ�6�#<>s�s�;k�fО����; ��]�zo�Sw|���[��h�q��hn��Bl����ej1G8t9[��SX������r2'i�Fȑ�x�Kk�3ĉPޅ_�{���(1�{bh��f"��Z�Z�Ng�;f�<��0kݴjoz���@�g�[����#�0{�˜� \e��T�������f�k��K�@d"��}�*5�_������s�&�8�vvK��%6��n�}�L���3Au>-���ю{�D؞�V��_7Ɲ�4>&10P�
bi]�d���9z"f��`E�wD�ϸ����6���/��<`��x�fR�,��-O�i�a��*;Gbx	�\�Un�Pk���z"�����:/-�)ك�kĕ%��:l��
�Nj�^J��hƒm�*T�CD�u�y�b���ZrG��� �$��^gf�A|�TB2@��[���:r��Z�R�\���l��*�D�`�*5�J������{@�`�㮙�G�3
��iQ��?;�l�l|HЏ{׌F�t��\ݍ���� ���Cٻ2"�@eP�K;�uʁ��.���Z(��H�X��=�u9I׈�+4��0�4R�-TH�r$��*��x�t�x.q�R���\�D H�Ƀ�����h�٬�\̊���xf���D�2�ȷrb���&�͠����y��ؔ���B�c�r���Q��I���oF.�� ��Oj��-��0TEp/��x�r�ˁ���TK�	[L�>��AE�h)΂(;ݸT�,$c@�}����44ϟj3d�����v�9� ��\ ��$�v�jY>'�<�'��L-�g���/�o�~����Ș�����{Ra���}��y��22c�)�Ҙ
:V�G����ʄ�]��J��)�X��ۣѴДC0��`�����c���*����߹��9t&���d�Ҩ�H���1�R!x��O���a�ʱ�C /n�`���d*�m��\�UARv�r�v�8���m�Nۭ �0�	A��lu�^K%��Z�я��]�%C�����Z=�����6�rGY�2<�p�~�<���G�ē!n��g��%4M6�뀁����z��r}wcӢ&��� ֆ�ȶ�%���y�qP�%�o����@�K�S��ab�1�6�����B~���O���='�|����;G\�h|QlH<��Z/8p�-�sMy�r���8b	��BPs-︓��ި�Zp3t���E��̴//ޖ�a.�NQ��/�א4�]l���j�r�v���($S�����T�z�
������?~*n����#>������#���C��;���fF�&}�e��ZKX,7' e���4�~nq	�S8�lo�f:Z�iј��Ћ��K,f}gD)3�Prt�'����SZ6C�/iZ��2o�\m���a�}��D�[�P�w�w:1�SJ���+�\cLZWC�@åd3�B�;z_"�w�WR
���%�&�O�VU�N����#��3�ƚjw�kʖw�UU�Q��YͺA+C��V��Ӏ��)Q��C����W�������!

�Lm��׊�$��Dw(�˵w)�︚i��~v?ɐ�V��f�	��_&@�/�"��M2MM�Գ�7ƪIݹ�����΄��7��[����&3�(?�-,N��7�V���l뀵���%����ƾ���]���������D�
�7QF�$QRN"	����%�L��z���@'���7�C�<n`������+�,1��v*�y��Wt���D1�ή�8*^�Y����y������x%���� �g�պ=D�8�=,��@P��5���IP�e��0����}��_!��L{���*��X,�8\�%��e'���b��Qļ&�!,��T:2��d�2�|��گ/�E����y��|?t�� >'��b5�����֥�ءQ)�̊jo�4�Z#�����vЈ��}���C�L�� :�n��躻�E�!�-�:<=lvv�&��������9���2O@��u��`�Q�-R	v��5���v���aG�(f��\E�+���5*�AtJ�! ����t\�Y)m��Xx�����	�]���iꏓW�����q�8�	����+D�ru�Q�����M��|�p�D�|l��i mr��ga�Y[E���qn;�3���(�b�#�^o���)Yj�0��H#$P0h�M��n���2����E�!���P��W��]I�Zb0p�t��>��x-U��o7я��'�k����5���a��x�d������Y_o�Z%�k�_������+2z�P�M�K�;�i���q����hb�-k�@�Vf���H����|)>[�SqZ�$��	H��{�s�&v��@��:��^i�;|E$@Esj�c "�Z�y4���F�c�G~�k�.��3,�Ά
�=�$�������*8	tJ�������߇=��,,�b�RIC((ʢ{��cD~'J�N�z�^�Ѯe;0��k�@�o�����t��3���]���m
E��>r�N"Z� ���9������u�B�]�k&�9��@8?>]�.����&�ȏ�Cu�B�]��>��@f^����>�X�+�� ��L� c�2�b;�K[�Rb�؞�5�A�=��T��..hJ�}�!h]��,���o.��R��ku���4tc(�� j��ԃҒ,�2H3;'#�[��Mc��R�<�!T�Ģ�<%؂r�B'�\�YM���1��R������X�Q>�k���'�(23�c2������T&�����w�mn)�5�R�ħ�,��	`t��/�.C����\Qq�Nɚ)���@�"E��웅LU�aeۑ(/�{�Mٞ1�A �xA�9��i\RF~y(Z�䅟��I?G\cs��DȎ·ZKlE���>'�J>��N�`�}6�g%���K��b@�M��+�P�5�xwJشٚ�W4!?N�U���+�������g�_�-g�	��MZ���Wͳ���f:�w�DW.�,Σ+���]����&���ة��GO�dTs��_қJ	rPsB�6_���W�e� cz�ȷ�Sօ�>�Y)M�{t��LO�@��\&�豪1�cW��.��x7I2�i���"�۸�q�[��G�P"�p.v�c �ߘ�M�����(�S���U �e�z��X^���ld�gW�&�~)aA��.o���޶g����m;�*���a؄6P?���^��ϋ���F�F��(:&��D�����,In�ef|�I���6Ҭ<@�}/q�p(T¦Y�F�Ý��6U��m;���4�z�]N5�Q�R�!���pZ�#q�0U�}�x�ɂ$�V�!�*p0�Qn�p����C0����.����Ai�6v"fU��=u�f#�u�|��s�F���������a�B�L��`*x�
�|���튚]:t$L@^D��U�mu�F�!�g�x��H�Iw�:�'cQ��k��%��w�7�����g��O�	�g��%��O�3��B�$�U��{��v�.COY��%�w���ͨ�{�PJ�{�'��Y����:��0� *U�!.�����?s}y�$��z�#�Թ�N��9�2c�k��
j���܉Ǚ��>���*T�~��U�K�b�q1M)�5xS��()�t[~>Z�sOˌ˰{n���
�88�����v�����hu�8q��`U�y��5,hL�6mf9��W��s͈qm�"��ŗ��͉�x�ڲ��
ޒ�j�P�=�Ʌ��qcd"��έn�{����Z�8I�/������J&�)���%(������17��ivx��9p��i� T7�*��8po��gp�/A0�Բ�;��߾c�:K5�E+��@U���hJ��3\Mx�ر�@�ָk~[�ƖB��3�û�Q_�/��Rr��8Q<���<ɟ5���iŨ�ˁ�b��,�D\�2W��A�;myJ��%l�zγ���=QfVq~SZ�\����eCe�
Q1�œ�#=���4���;:(�f�Nx�4�E��3y�m�
�����~��o�ђg��K�S+	��g������#��v��E��P�G�_�l�>(�$��	������&:��� XچÉ+�(<��$�R�i ��H���B��Ky�������v6
+�U=FM|Ĵ�˾|��mXC��LsQ�6��ɴ�'Pl^HTZ���k�G��r)�nG�;���8&��+�I��Q���$�->0ҽ���=xe���Wg�hJ�����O5Û�Of*�aƈy��ҝP��a�ab/�j�[��!!H���>�Z��5���#��#W�Zj�V3����yU��'��4��4Wsw���%�>�6����eބX��^�ꖊ*���y?��Y�I$w~x8{32wt�AHZ���dA-HVU�N��='>��x�1��f��j}ʚ�ӥh��?'��r�Y�>��u� v��?G�qk=��0����~���<sN���aMe{��Ѫ>2�ܾ�ר+Rn�-w����^�X��ʘ/���4�)����F�co�KR����HTђ>�jz���^��妑V(�;h:4��"�0�E���e;~��;:�6zBDF��3G�W�$ҕɼ�GsF���J�=Z:���@_	'�V!�$X� |�+��Q�t3,Np��:�]F���ߓ�
Fpr�22(u��
7��@���,�+�c�A&�QP���F�e���|�)�>+�F�0�1	5Sm>���b�Qџ���&���4) ���ta�H����11'��v���߾ ��c���@B�h����k�wJ3" ɷ��}������m��3ߎ���/�2W����F<�.���yR���3�6xn�N@M6'~�T|gr_�o�j�f
"���V�r�u�����՟�S��W=�H�y�(��D<vI���v|�^�����P��)Z�(����Z�dK�H�;XcF�bS�ʟ��d4v��]���'=k�,���if�΋uV�<��K�o���5���JG<4V�^4	=�p�}��4�c
�װ���b�q��}�%�z�����C��!޿���-���9�m����ʈ��Pq���S#+S��&?�l��֣�	քSG���Sʺ"�|�Srh����f���ЀvI7}����t
A��	�ȭBx�<����fŃ�;�o�� ��q�$t�/u�V&m\��M�:�\�����-�M��{����(��[r
&��\�0�M�+�]�xe�.膚����*��Hz�z2�0�/P������`��>#`o5bפ0���<8N��pw�M���G�$�fi���]�!:�MVֽg��=��i�m����	�OU"�i�h��D�⚤(0�-���(��?n�k������;"k���.�NL�+6�֍�
������g�i�xZ��埕c���ғj��$�����Ǟ��<�4���<�:��?�ٴ�WX�B�%U\�6?tE�ċ3B���]6��A ��T��<��_/_�����5Y����S�T��""��91�f�NiJ\�,��fvMe�Q y|3���E)�}d�>�������YmQv3�r6OD;d�)��g���h�Y�x��<W��鈽!�z_9y��}�'A��� 9{�rXJ�Tὸ)�)X�5�p� ���d�U'-�/_���|�5.N42�NFƛSb=�������OS8��\l��1?|��T)�( ����~	�B��b�<�]SC�@������ �z�K_Aq���Q^@d��m����A7�AMEC�G����a}Fu�K�m9�?��I8��@��1s��t>�Gʥ��=7۶�+�y���_C�%*'����3�����9����|sw�0Dc+�3� ��:_ǝo��#�W'�'��v��Lk1�>.fCbeRR�3iE�-�#�S���*^n@���y#j�W�|����M ��<�
�"�m&�B�Ua9�a�-[E�� ����n"\j��Z ��k"�.Y�7ĴC� R�=]�ĞyjQ�[�N��r*�
���>�<~��B��%��0j��t�)<�	��Fk�Dn�i�J�,��ߕ��&�'�+��_I�gV��y*3*��L�G#Bd:QZ����'�{��pWtu(�	bs�t,s�_na$iT�'����y�ff5�3���Q'���C�Q�"Z5��ڜѱd��g�+�O� �n\<L���FTN
18�I��۶5NiSFV���m�\��@F��Ԯ��;x�>�d��1rj[@�^DZyM�>6� �X��4�lj�\0w5��/���[�&����ȹ�&#b�~�+s����x��Osu�Ybp��hb�g�u"7#��;i�ʙ�_	kx0�J�� �]�:X���3g]��R`4]����;��r�s���F��8�4bo��qr�إ�͊�畹�8#����'�(j�r8P|ȵɩ�@@0��v#%��N��2�y%Vch��F0��ʣʂ�]�Kɯ�Ɔ[X���Q��������%+"E���"�ywJ��{ǲz
3�asI�����`]���Ļ�;���#������.=���d�.2�]�"�s�-Cۨ0�� �`��Ἁi�T�߼�k���'j:�)�������qP�;ɇ��ӗ@L���b��3vX���`����-�C�H������@X���'�k���IƱ}�I a(�g�hޭQ�������y̥G��ڕu�a i���]��C���VO�]��W
�adw�c� �eIH*9m���hسm%̀��}}s����3�.�(\>_�][[��/�C	� ͸<�[��*�PӺ���.���_v��U���B*�k�↍���f���.k2g'��ˢۚs~�YAىxd,T�7�����=PIj�o�}m�a��l�s@s�+�ۆ,-��e�T��	I��8#╮WR���5��'r��<�;f�ۺ�;�㌠ E�7�c���3k 47���$�n
_�!U���z�陵T���uS]��r�>sn�nx�iw��
����U32϶l�)?S����ȣ����D+,�Q������������Q?ּ
v(��Z=
fd���ZI|d%�ۀt;���)ަ��5���������8�D8U9�w�MO1�C�k���0r|xO���R\�TiB�p-�GZ~��C�"�wx��	j_ʇ���.����jm,iI���s}H��3UC����ʷ��ݬ�^�8�P��^y9����ï}��KL�s�Re������;'���t(LPͫɛ����b�[�Ƨn�Z��qe����i��/	��;iܠ>�G�ǈ��m�n�eF�`!�H`�ΉvL��Ҭb8�ڐ��xV�	�]�!�R��04Y'���n���}�#�]݊����~����P��-z��*�Z�~�o��S��`�rO�gW�]��@�հYyZ��ԫ����')��WA����W>+��5j�'Ԛe��0/���
�ǌ���3D�*	}����F�!��3�-��O�7J�j����?� y$(��i�f�$�<�z� Y2��?�S8Wb2�2�bg�I��Sx2�����ՏE���#�N�J��;�Ջ��9������8\��C��s���- P��Ş	���{����{v�L4�e�ήB"����7X���8�ش�=���.�f}�8O�k�C��߯�K����":� �I�z)��)�raՊ�x	%,S�ii��ޫy+�LqO"�!����3K��%~ �b5��eg��a��ENGUE�ۍ��.Ԇ�]xR6/e �p�Ηy�ޡ/���ҏ_�t���� �����q�����6���sΊdG�+C�Zq;�:��(�7v����N_T�;u_f,=�^��10�kG̲tG�?u~Gܑ���!W�<o�
�/y���$���sֿ����X��^]���t��lܼ*?���bs�|�L��o����W��7D#�x[��ZA��3�q��M��D>��⪍'�{'Z' o:���b-��M�f� �I?p['����1 ��i��訫f�	����/�P�U�����Η(�#!�:Oр�TU�r��<�1�"�o�r�2�ʤ�s������6�ekPR�b/�5��ܝ�W�z�3��1Wo����Q��yG��	E{w�v{��h��!˙`��SA7�	*@����>q���v�	��|M~��[�EՈ�^4�	�*B�	��\���Y#^s�C�����£�<S�0��4V��i58~p'lW鸵�o��[�Ğ���"*s�Μ<�n6L�t��Ǥ�-.״\G��fU���_YS����pd�l�{�����K�n�z�I��y���`� /�[�M�"C�>�m�]�� ^�_ �o����j�h��I�\\���l��󌥫�V�c_ �S�R���u�ٸ�^��ߟ�^��._�JYʎ:��H
P����w�ع/�B�����p\��?ԟ���vs�f�Ŀ�[�Sg�>�.�*���&ݯKoB/IJ�-���G��b+~78�؟$�ўt�*��B 
�� ����Z0�ER�������ԝ>�f�6e���!�{�0��F�5N�Z���6���t��gU����_��sR����ru���x�3R\�<T	$e/iV2��*t��8�y#�е�����z�'E���F���8	�SW�����Aw�w2����cLb4�����cL���bO��C���(l��5%���6wJp�)��H��w{�f(Wė�K��u���v���!K
���uk?12�5�L���	A�����i:�.�(ֲ�]�K�[�@e T��.�u�~Z���\��}W 򗤎���Yx�, ���a��3���&�.�P2����L��k��!wEo�͌���!P�of{�S'T�"Kq�1�:�xTy��H���9��&�w�s
�������ú��@ߋ�<�\s��u5�B^+���i~| �U�̾p֚�p�|6��/YCQ9��d�𜘴��|L�lz���OO	�؝�^�����H�̐�*���Dٸ�{��L"�t$�G��I�
$���ՙ>W�<U��C�Μl�U��n�;c� �=5�$(�1��U� {�]�5-�hB��j'6~r�XI�A�'��U�lq^'��&��O�k}���A(� �B=>W`�b, ��|���r�y�R/N�"$�X������Z*׬�'���&���j(��� ˟*(,�Ί�g��^�G!9"f�V�J�o��8������I�$t�q����9dt�M3��^K:u�BiP�{�u�g����,�ycN�A�k]L���"�U��>�Gc����u����Acl�YFP�-9-8D
u��8?P"j�ȯNU��"��ΰߙM����'uQ��	�M~C%.`�/�l?� �C�����s驥ƫ�#�8�6��}�gi�E��$��n�����F��H�Ƀ��Ut������{�N ���|	��= ���"�W�%� �1�w���5W��=��}�%ᥥT�,CB���;7lU$��'�����qQ��Qv�C�*u���!�)������.��٦�X�ό���ES��DȶS
^��\)m�KG!��417 'R�E�
\=����[�F �K�E��h����F���-ث"�� <C������0&��q��o>�" �ᔥ/h���"V�D	�]�.�F�H@��?�`�uf$1��%xk��$[�:3��$m�䓩���!k�7_b��"��IL�H=��J*��T������y}����c2_ws�3D*Qnz��8]'��M@s�J[��/�R�P,xH缿�t)�`���xpe�x���,,xRD�}��\�Vz�V�H�j���yy1
�Ƶ6Q��
�T�ӏ��s/i�v�8��(��@�Ym]�0J���rZ�2���Q&��0���6H�ޣ�7��:x���0�U�Mۗ�X-^P��䁙����5#�V���9�9��zl},;@ܺ��P%`ӵ� _7��WԹ��Ʋw����ar������K���xQ�Jӓ���ET)�?��X����Y�$�AD¸��i�O�a$��w5��$����r�uZ����rQzsI��Ʊp)����V����d�W��|�k�\(\͈y����}>��E���?7Q�B��u]:��9�)L��T(�b�V��rs�aR8Jg��d�ǂ3��u;�<e�<Rg#jۇ5������^�?N�TI����}��R�� �+�:�Fs8�4�' S4_��Џw ��7�mLB�O��)൘�e�.5�ÃdnkAz7��_"���:^�$"��q6��d��Y8��7��j2�#��fP�#M����OwNc��~��=:'�o8F/�g��B>'�?�H�n��x���3���Ea2��$�����:	~.�,�l*���?���7,�Ҟ�5�9츄�(j�6���^��|�tcw�,�BY�����J$�uP��d7h�5�M��fp�G�#�0������E,�y���y���z�| ��,���@#g^�e��ɏ��_�M�ʬ+p)���Rq����@��{�ä铽Z�<c��4%g� P@N����Ez��-x����qfF�<k�*�TTH�N���P�ڴ�$<��q"O��;��&&�4��<G߻���:�u��f��~�[��t�zO~��244��HDJ�9"P榅�	���LJN�,�^�H�U���Ѹ|e���W[Rƃ�6���V�*����pr�g��?����XS;�H�7.Z�X�x}�.W�	d~�)�`;Cv]�WVO;#���^�'�#�3�lW@t̐�3�.@�j�P��.������d��7����/�"�r���& JE�����`9>a�x��[M.��1�]u�zM�9dMI��B070��b��&^���~��vX&�]"!��%�����*�w�,�r��^ډ6�Ls��2�a�/������zef��*�4�F�Yv7Z�d����5��G��*�v�S�fvs��y��N�;M�H��<
 �쫪���J�f�Ez�/�T�G&3�cU�� �G���;�d[�5�����䥥��Vr��*��|�F��7+'
�9x�Z�z<�W_��k�u�[�F�pK��-����`hw���9�f;���q`K��rɇ����vXl	�n��x�F��)Gw��J߄ㆃba�����C��Œ9+��]��5�*K��41�լ�s v���0�8 \Ɨ����$g�����`�SO=�,T@��Lw_:�|`�F>�_��n��*A���itʥ��"e�C�&�y�+ߐ�5(^%����fP�!�B]D�!Dp >h*�k���`j?�DP�������a��1�fj>l[�Uu�S�IkuLx;��m�O����*�^óY���a�@S>��LUA&��S���]�ܕҖ����Cf�zܵ�saU7A����p�*���fh��#��gP�d0è��9�G����ԝ&��b�S���v-�/,8����0�L��8�TC������&����9%a:{�ڸ��n��ǅ�0�^WȄ��i$}ҝ��U�{ߧ�w:<1�eI:{��a~�Z�I����� S��P��G�iqx�]�ӈ_e�xٱ�V}���)m��Ƥ.=Fj08���d�|�!��m`�C�́�O��M]�������A�	G0��"���z!uc,�K5�րɀ�D����2ʡ-��� �����smrXAg��S�A��Y�x��0�� ���B��n-a11Ql�Mh݉�y�&�6�V8� �-��oi��:��v(�@0y�-i��1�f$}�Ŷ����@$1?mN�͇`�'Ҹe������"��2�|'��~�7���M���=;�5���*0�e/�0i���4�ֆ<Q����h����(xm����? ʷ	*��jz׆ݜ��e��z��Kaŭ>ahG�mQ1'�u��fV�(�E�rK�c���s�C�T<!��o!�����۲���1�c?�ˋ�6�s' r�V0�|j�_�ĩ���
��+�E�Z:c��E��r����%Qo�B�7tވڑ����H���|���t�:�����l�^�g��AG!W�RX�@�1şucDZf�R���;8���ke=�_z�&v�~ 5�e��Q�)��Hӓ<++OW�vl�:Hl�\G�e*y@I�!�z��,���,��q�\��%�'�S���W�%!v�����O�么�Y	�̧��t���?p���<B��r�k���tK3k��@�zNp���4�D}Nl��dsT�v��.�.�R��S69���a>�<������aʋ.D�B�����>�/VnW5L$l�����:WX��þ�9+��j�-%����
��MΧy�ي��H������������ӊs�.�X�k�6�r1n��J�)Dd�[X��*�PI�T�=��7�A�\�o��%�{�S��̀��r+����r|��y�����f��QDɎ$��v$���N�
_�כ���;/L��_���xj5�WR�Mj�M]l�=l���2u{���'C��Lj�"��>��0"�<�V`+�b�	^��3�bM��aFɶ�A��^�t��1�"]��.R���RS��y�F�t����}��u���!�t�;���7�p�է�AW}��&�u�u�f�e��z1��'�^��b�;�wBZ>ް_�Ed4?$�ڦ�N�l�^�8�Tn���J�\�F�5��x��W��#4M$5��#B#)"���x��C��u�G�����$γ�.C���SA�$����m�j�p���oe%k�<��-���ب�v�4������/h�!@
�����T���I�3՛%S�H���ȩp��.�p�X�aT0��nԣ�#:&��@Q8��$�M�|$D��_�Dj��e�o���0`<ϒi^(;�����R�֐�YZ|脖7�tEa�����y$2�s(Fd�(e@xq{BZgt�uo󻊌Q�z����5q��3C��c&�z<ly�Yg})���j��~T���2�,���"��X�a��[c���*;]��C~	(OB�HNМ#s3s�܁\l}�8�M�rص�#��a?����3�R��ߖT�"��kF��ui�iݝ�e����8�`�X#�Z�ؑ��T�M�v,�F�Qcm��ԡ��5&�[�8�e�U�u􍹕�X�iQ�W��ż>�y�t;�Z��m�#��;��l��<R�Nߝ�y0����S4T~�k՛Q�g�$p*���_2qX�M��݊�;�#tءY[w��0��yen�^k�-E����P��TZKӆ��l���N�"���z��!��'��#8�����q,(C�IN�A�N������g��U3�F�Kq 3��U��2���9�Ț�A��rS�f�:xf���O�X�6�tU�qH����wz��zbF�Wa.eE)��i��D�X'x���᳽ɦ{n/��-1a�(]H��n��l2����q��«�bC{�8^�8���'�^~�9�Tz4*h�-E/�=v��7����獿]6��	 �Z�X��s��%����^��2����(5���G{-]
��E6IV�����Pm�$@|5�(��4���iN\צ���V�'/�m;�	�wϔ�*O����Q\���77������]��~Y��J�7Fۥ�����hm^ܑL�GL!�4৿2	�F���������$�����H��SBA�$�n�������X�(#�+�����t��#C�7���C���X��F�΀��7w%�*�rJa�eˡ�����?dЋ��<T���Jia���{Fsj��`�A�_�������HJ����$���2[A#��
�0ΐ����$��~��c̹�t\Q��e���|s�+�ʣAR�H]��%Q9�@�N1l�k#/)o>67Yٱ�bD�u�R�H6]B�oļ��wX�E�ӹJ@9������9.jIW/gK�������C!�f�Q)<�$n���&�꺵CGā<����c��vS�Y�a�hxn���
���Kof����5�/��
��ѽ�~ �n3*|���ֻP�w���q7f��� ;V��	��iK�q��}���_ ��V��dRI�,1�|oK����+��(�H",�rC��R;��䚿d�jUX�ܣ?Y*�uq<諪�<V��T���O������%�UD}4&�{�Ɓտ���.fR�Ao��C�}.k���>�u����bD���H?Cx��R�@��4||�ž,3*�%kwѲQ��={��-���g�,�ð�|��x���1�BgM����M�k��jR�	; ��i�gO�ӿѿ�C�(�4ew��؎�jS)��1�V`�|n:o�k�(#�E�S[���vO�W3+dA$a��X�����)ʌo�g=G�[��I��Y��|�CU�ۿ.����>YN�$�'ńǃR�-�~�`z��I�~���:�%��[:㱐�����m��Y+A���E��$���{>e�?z�{�
�ѱQ�<%7P�nD$,��ˠ;'�rD�D��j�E�6�j
�����i�T��l6dg5�{��FJ��zo�ܳ����M�F��Y(n�1%�j%2��1�g��hoH::Bh;�ЈAb��(-?�z����9�����C�PM���(�o�RN��X��th�.�p�[��0y�g�{�1.W�,xQ�mt;���@����:��b�+�n�U��B�k6�����ځ4Ĝf�W��;�8��n�Y�ċ�({�C�X������X���d�[
�e��v=\Ô����él�^��x#%�M�plۼ��J��^LR�@�ʃjH��P>R�W8�����$ZG��S�2�����ե�K.a�H��h;��N.��2CV"�۫���&rP�/�P���p�-d.O6��E<�D�{S�Yd�j����k��e�(��sXl�r*������:ЏW��5��ߓ[�Qp*�"�� ��TH�
zh�ƫPg����b�T�1�mʜ��{X�R���!����fY�g>,dg�7���zr�`A3 ���$����%,��o~<���M�~��I@T{�:�a%C��5�cׄ.1G���K�#*u� l�ą8V��G�
fq'�sY'(#�;���8�����
�i��+t����j����a�݃Z��M}��4�_x�B���0~��+�e�T��Wz�$�4�w��"���>�w�l�'�m��T��`����I�2A�^UGT�&�x��}~�
�-b�R��H$ɕ�ɉ�����BsS:/K&�ն�I�$��죎a>�9�=�\����ExbD��/��6��Kb���o"��8+�LM���������=��~[<�9e��k���[�.�C�.4�4�d9wFB�N*z|��l�VJ2�V)1ڔ��ܩ�|?�K'��jK8M�@��,m3@���a?/)��0M��ռ�{Z�q�|�ߥ�7ȖK������se�����T1qR4���E���|S�v�g�OS�$}Y�Î��|8��"	�����I�a��]�����L`Æ�I'#	�����-��ޖ�2�=.�֮��-s�Dy!(�VC��B��8k�r��,@�7��)E�kz��k��b�S[3V w�Ef�I���;��3�ћ6��!o�h��ܸ�i4�J@q��m:��^��x�L���u���U�xrI�|T';yan���b.Ƴ��Z:��S��G��MlN�'v�D
�SpaAHQh`���/-�>�׏�U6o簍���E6t��lzN�����Bq����EP�M��{M=���?\����F��ب?	�k����`���{��f+���O%P��Ը�b}j��j;,����={>6�.�p�Uik�D\i�W��t�.&�'�~c�Ό�N���"P;Ip�w=�n�>�2��S񺣾����.��g�~�g)U%�a^�cF�>f���ս�	���׬�{YvTr4-��:�p�sKc��'AD��)ۺr��3��L5Q�yU�=���c.�Q��o9�!���p��`7��THmÃ�[�{�XC�6�������G`�޸=�&��u�ߘ	2��=W�?���atY$�>vp�0�t���Ff#|��A�H^SE;��?Z�7�ι��c��� ���h��[�߭�OW��Vv�v0��}@��I���+��)E��p�!/���h1k���8�KU�~��O��[�u�_�T�:���?��6̡�+��:�x�۷!_�}	���ʲ��р�vh���uGO��U�$3�p��.N?�i���ԨC3!��j
����3�llU�#�*� !!g�9�w0��F8l5�`��H�_8��3e�<���_@?-��f��Ϥ5 D�]�X��ܫX�F��#�%D���z
Xg�f��J]ҽ$�;��S����n*�D�k��ח=���Y8�A�AuR���EG��٥�πB�5}\~=�1M �5)�2�U z�����!��L.b=k�u�����}�asQ�.�=��{O��@A>�LW�qGa�1Y��c����7;t8��ʱs��"j��Ǔ�a+�{A΋4j�A ���nI�Xu�O���f��L N�~�d���$��u"y��2��3R�u\H�Oϐ�*��f��I� �&CF����p)��m��p�d)�OĮQ�$t��q��D�I�Y�>�oF#$Ff0�A�Vw�oM˧�b��⨦�O'�#��2ϝ�DR�x"�Z5f�7��2i�R�wbh�|��x�y}�jq�u��.�yKKT�Up��b �!<؏�P�5�B9�Q3a�}�H`�P o���{:(X�R�w�M�@�M1d��4�P@G� |�y�✬�o>�ՎP�����jV�{,I��ǵ�<Qm�.��S��@sR�c����'��A�/_�,n��,���=DC+����Bn�u�dA��;Wӊ����ag��d>(?��ȏ��踹kn�����J����{�
�ρJ+�V2�T={fV�@�3���� K�8e�_��0���Pi�X��lr��yQ�Qt��f&�9��Ĕؾ�w#�h�!�jk%�>����ux!�a�`F�u���#��	5�?�`�e��8�`}S�%��x&��^0h�7�� DpĢ��s_�$����Sin	�!�b��.qrF��J2���qh�l3Ye_�5�o/F��R�g�yZ�a%��,�-!Ր?�f����T��K�KqhdR�-8�����NH
AI���M��w}Y�3\i�lPV7c�\������Ek����
����b'Ć����i��s��t���9�p�)5�F-��؁��/��U�M��Ν7�Ac�k�C��>nCp��}�Xߛꋓ��4S���(�u��ŉ����0:���͟�s�?���=@���V5gF�{<��`dޗ���C�Wn�K��<| ��ƭc�'qt���F
>:%�Cx���5aw��g�{���P����?U�W���eTgִ�!�
FZƶ{U��<TBp��f��޼[�@	kfRT���nK~�33���d4��G�Tp7V���3�U�Cc�m��9��lT"�tݬ:0S�8�>	,���?T>�fd�Gy^�[ũ��ɛ1;�w#�l\秐v���yAG�b��B�R�o�=W����=�O��U�ب%OS�k'��(�������Fg�P�C���݁������֍�;���0Sv�]#ђ��OYfH�7��ع��*���#_}n����k[�ə.n�
X9��l>��ťY�|Z0D�,F��y,�$�wQN�`�����_����l�h"��⼞�=��	C��@���]9��Al�7�?�8ἈWYԖ(�^���l���2ۄp�V H5��(Nk\���Wr�.۞�� �j'��)Εs�_��<�	��q'����T�wێ�(/�i�d��W�nɩ����0����3Rz��
+AN:_N�?k�N/�)44-WE�������_�}��X1�� f$H(L��/�0��;�6-�<��a![�-eI�d�l�8:sb��e�ؔ������.G�\�]!4�4���G�Q�?FZڦ���=�Fs4~K�uH!/�.1�GF�I)�{GYh_
H���k���lY��maK���A��6�p��B(���Pxz��T�i}�7�j�k �X|׽�6v�: ?D.�H��.�P>�	�߷՜���;�D[�I�8�r��8���\����i�܃B�!	�wL@���f,�]'�k��a��:�#2fi�{���ٜ}�-����b�f��#K.=�GØ��.]�d��q1��������QJ�o�P0I����c��Q��>y3�����eS�nC��ab��jy�v����I�iU�%��T�@��]�])�Ƞ�mq�'��Ks ^�v�4Q]��o�v��M��@ }��4
������ro#��I����e��%�d��xd�p�J�)_JNl���%!f)pX�ZK&��N�WHq��Y��$�3nh��S�W>���3�h7rk�)t�-l�s|�\�k������.t���9�z�/m�����_l���q'p�u��w��|S���w[�\E��)���_�ZR��U��a9b��S�f�w"��Y;hK�\�x���ePt������|�9�+G4ӳ�F��eW��}�� �`�6x����9�z�$+������ .��
�	So]%�"�L=����"�b��h�轺�Mݙb�=�)�3"̪H�Y�a�k��7<[�#�j��Huz~7�jEI�Ҁ��"~�]J��QJ@a����� E�sU��c4\r�6����Y�P��4��JD�rxSBl�p��[�+[��Q��1�h)W�)(
�W��
$�mK&k!r��L��<�ZzZ�߉�4����=����^��r�W��Q�L��cϨ�A�VKv�7E�Z�%�ˑ�Fp�JɈ��&��J�w����H�Gx|� �]J�=*���D��C8B��� �7�X��\�J��\�}4G�Wn~J�f�pi�ԛe�'�P�g�E�����ε�R/hf(=� ���w�Xu#�)�{�d�B�P��z70FH>�z|���EǬ�,��{�H3����?Z��)�E웚�N����-�@���4���[<u1� o�|�I%�'�� ԩ�ݡ(S���҄�6K�V�ƌ��E�.8�]���- ~�y8�&�!��5#Z0X
_~j�u��������1��(3<pO�\1�d7�����9$�EcdN6�y~����[��n7�6o�(tr��gr�j��VD3iZݫ�訷&���$ �����V����Wߌ�qB�;`�Ym+�Җ��}44/A`��됖�c`p[�0�R����rfuմ� $���J��`¶���垅 ��#�%��ݸ@��|�I��-�cZ�݁�#��F����5��h���I�^�6���3���u���q��O���
�����p��L=�������
��.Խ�8�㮃�%�����hF��mo*d�@���N Q�k�C�*z�k�=w������&`RL; �o~�$�.b�W�Մ9ґCL|�@Mp0촉M_=�� ���1�qu��-����j��D�64<����R'����ǲI�]`姡i��dÕ{�\��v�.@��Zc��Hu�p.q�H����G��B�-x�AW�{A>}]_�-�ݜe�iI�����h�u�T4�x��{@"�W�
K'"Q�a�����,M-�Ŷ���-9u��!�?l�	��Du++�r�y?��e�%����:se{h4n쫪%��b___/Y$�����ߞmL��ir��z��U/Ϳ2Kn�#8/?;}5ʿ{Y��z��R�i�5]N�-yz	��]�W1"���}���k鿔�*��U�}+x�Q���֛����@�Ƹh4��� �����Q��	"ʲ���A:��Z���@��ED�G0���Q	\�iZGU�=DF�6>�˩�NՍ|����q�c�3�߂4���EW�Q�RF',�tO��2����D�6܌ҿ�xE�:2�xq�����;B��6�q�)�^B�)�B��ŊV�w_��i��(/恏q�D�NY;���0=ife�B�����p�g������.	/*�.��G6���k�]������!={s�3ٴ_��ka��x@)ԓ�
Xx��X�Q2�RjL�z=CL���e\Ώ�jJ1X9�~���w�T\���f	�&ucS{�X'iǶǜ�b�ۦq��"�a�����=w@���>M.=�7�O)�ժ�V��X�A���dgO��	�NM��P)5��Z����Y��L�μ��}w��&�\�J�����V��I%�
������W�h�Ե���Sr��ۂq�u�U����b�x�[bșn����a4!	<$ ��ANe�_���}���@��0�@U�Y�N�N�	��:6���i5�2q�y�+G�|�j����C�I[��p?�X�0�X2qAu�Ozh�;�8V�\_�����"�4S���K�¬4����P�a��TϻPl��[�9q�1).�iË\�������p�-L�>q��0����Ml�K�ں3��(Z��1����
�r����e<�Izn~h~����DQ
{\�= ��E���\����6)L���ѻ�S�r�C $�M�8\h�k�{Z�P2V�jJ� ��X��=I� k�$`�C��<���V����`�xw$��/C0hBbu�����K����*����ˍ�q�V��e�e�+LE ��������=ICTL7��\��#5?����㏟�[,{-�ؠ �k��*��>�����)U_�op�N�nEFzmQalh��ʎm�Q�-&I<0s�ͯ���i0�A������L�����%X�F�V�[���aIb�I�����w^ih��5�x�g�.y�#_��!���;�H_6&�[))��Ҕܷn^_�����$D�N*	6�gN���T"T2�K���Z��O⠠ĩE}U��y/9ݹ���iTyS�N��^p3�܉�02>��&��5�ϩo��&yh̰Ǭ���t87�>>���W�R��L���&��\O(�hT���X��\�]onptKr(@=�i衜��ڙ__������k�d�j���ӆޢ����os�/���q�D�����/a&R�-D�]�.�F�K��S^
��u�0�2S8X�2��x��E�׭[�[Y��/MG.W�0��؟U�Q�DJ�[�<�FX����[�@�61)3�(���� \�]^���r��9��}�D�D]}\��bAU��m�QoE�L���{�|�n�
��D zS�t��;�1i�Wd�1,��L�)�&�B��T���5-*�������i_���d�e��s�������z�B�{S-x�TntP: �����-D�̝\����Dvr���!F�ir��������{�w�x�h����r��� vј�۝�ѓ����`��7�gz�L�M�r�M�̺�=��(�b'1�`�}�ՔV�9]y)��j�|��Ϧ�C�$p� ����{lշP�DT-���N�M�Ɇ3I�>}GSx�(��O;�
G:���� 5mn���=�\��Ihʨ�o��Wݟ�_h�N����@�	�RJ|�c=vl��:�_:ajl���@y���Ժ���}�J���h�Ӧ�,���D\Ly�)c��1��٦u�I��0+���.����Mg3(�}_�����u������bN�9��q�? ���ʒ��u-�40*B��Y�-�ܡ���{nBM2�f�q����b5��Ë9�w��Y���y���3uVA��?,���KBtu���M0@|$Y�t�;���aO�Y��ğ�3��.�k%�h���ql�����rQ�Ā[���i��H�^�+n;n$�H�#<� ��o��������87�í��r�bz�K�2LU�a�$�t�I5J��ؑ����6}[�����9��Y)�Ԟ�.�������#]�i����a8Vg@;q�{Ӻ�j�����|8�o��U&�m�kRW��?��p6v��^L�I;�E?�ǵٲ.g���-%��J4�*is��Z%0������[`�
o��W4\$�kﯡ�#"�ղˮ�b�<9嶜9��P�#�
��sx�L�<A��5	�@�Q���+��%���Z��]W(K�N\�l�Dv>P/C����=ڥ@�e<�/k�0�S�8���jx�d�K�;�ٹI�G�w�nz��r�\��r�.��_t��R���Uv�9~�� b��j}�SNS�rܶT(ԓ������(�k�DJR��<�YvNB��b�>�9Y���U��;x_H���X+�L�>|�����2c�89I�_��lm{+Ʈ�w��?/0��4'�_jyD��m(ݥE��ن�%CG�������C����a�i��b�h`��$��{Ÿ-�����Ab�#���p����W�#�x��F�S�q�qӊ}�$�j�a�{X	��s��R��5�\KtS/YEv',�į���P��&rDD8_ψ�u��r�̜y�	K/���&�U���1��3�ygM�����`wH��q,0�愇�}Q��t������6|���,.�k98˪���&;D]QXlp^q����F�'��{8C$H�6���@�}���4����3�%�wB}��Z��-o�����<H!0��%Y����_��s�ٽ�S�9W������Ӊl�7���잕�ݴ�L*���2LƘkVNq�x��<.��V�9��m���:����	�R��x����,��z��=q|b'�I�)�\�lku����c<Ӻܨ�s7D�+�$�z�O�PI�����z�kk]>�_�N�bCn�u�T,r���z��_ ����a�G����*��:��)t8.~��B5M�oU�
m����v=Z��t�g�ks�Re
ɭvXj��}j�q�:�+g�\���}R���Ti�nƜZ�f�O��P��j�>�������H�P����6�l�т�Ë�jhg����.�2'��V���#TޞG���g�4�J�k����k�t�8QP
*?�>7�:͘��v]��a<���￿7aړ�0�J%M���$��� ��5��h����#�ǌΔW�u��!�^4�wV��	'� Ƃ�ծj�d��6?��;��dG�x��IK��o���D��d�����h�oƙb�а�����Z_����FANШlY�Ipiq��!�I��F���~"��{��-��6E��~���	��J�ځ�5����=��T�kE]<��:�&Js��9:	g�G�5� ���t zK��7�W~Ҧ�v�b�؅��%�9lsTv��&2.�H�F�؂kZSv���>��I�t��U�Į1��o�L�y�yy*�Q��4Dg�S�#���gP�����:H
���7Ms��@�r��+�nUC�D/�<J�����5)�9NȾ�g ���E�ߥ5�5pL�pQ-�2�I��ǖ<��8���};����?�/���.�2/(.�pe��X6���t�X��_pb��bI�����7
b�߭}�V0��HU6&R��D[�CI��.u(]@=
/����׉6��1 )�[gTa���Z�4J�3_���U��_��Aō�d�G�w.�����|���mZV�M��lHǡ����Oz?���%>^�,Zr D��nȧ1H���)JL��m��m�KY�p�H_ONǵ�@�r�_$��ܗ�S�Q|�[�Q�:�Y�
���l<1K�j����i�*��`�Y���^3n60�L(��I8ۿ�}oP������\?y�N�Y9�uEh��m>���w���D�m�����z�� �ɷ�K�5��P���n�6����`��(�ڊd�jj�7�t��ק� �u�c���l�)y<Aa\�T~Bl��5��"M{���j�@�!X�$��N�kڌ3����b�(�u� �44�A�ಯ��`9�:��	�?��%�]fsT/1���w����:P���� вk�����֊�[�y��`�O_�ұ��0Z�N�4�T��a.6�b��oAQ������ �o.ǋ0S�OO�G��t�����t%��C҇K�š�C�F@�W;�h��:�܌�����A
��!�� �0"�Ω0x
�p�b�%��s��R��ROс��8���Fa���..K(��0��}� J����yd0M��0�$��8�Ťw���>�֣V��7+�*s�у�h�M�ؽ'�A>��k��(�\�ڴ��}��<�Y��.�3_O���m�>zZ��,����a�������N�o�;\�8qIn�B�o��	����9�ݵφ*	���ݴ'�_��6��q�l�3
�	�9l�:f7��S�K�D�3O0)W�4Mf8�'��L'	
�M���X���0j	rk��ҷ�63~ !�ۺ�Ҫ��3�s�eҊ�"zՠiI���m-�;)�[�Ku�əq%Pl�?��S���˒��R�(�0$FC�R�
� ߓ���,��N''�o����w͕%�q�/����_Zն���H��Be�}&��>��@/��2��5��\���"���]�Ȋ9��%ɪϬ���)��������.��k�����צhF�Y�%�Ŷ�ڡ��Y���|x�����B��K6���I[���ae�]B�OQ���>E)t��Ą.�
�W��/M���v+�^��3ԸU�?~e�:g��A]�`c7��+q1��'��<A����G�=�iN<��]N��m�"n9s�EIb��v��=F�Y(\�$��m��t��vՒ�a=�q��%	�������-��-)���e��� �X"�Z��Ec��RB1���
6]�md��N�#�M�.=�L��F[9� �swD+�Ͳ.`-b�y�-����U�k���}.'h*� �،6���a��N��*�q���G��[vZ�	��^��m�Z{
A=��PR7���_��Do�y�tM���iۮ�ݫ�/n���Y'6�%C�Ҳ��R�%�v��m\/���P9A�(��1��@�c�VK���q:ܵفG˜��K&qᑄ{}[л�{� ��y�>�D�vL`�����m�	qS�O\�̩j�K�f�J^Nf��dq1���G�	��ݻ� ����>lcٛ��u�T����|B�g*����>m��4����6N�I�݆��mlo�@�\eu�t�	`*'�<)��%/������<����Ew�ٞ���5�<�\|�f�a�:�z;�1��;��r�f���ZC�r8@�u���x��Zr�G�q�3�zR
Nĳ�(�<�y����~�����d��?Q�6���f�����D-�'I�U˝s�4Ոe�P�*Di�d��Q��{�6�o������Zκ��A���dKYe��O"���R��M�/�7Z�X{fݨ�c�e�{�V�<�<G��c����L���M�Ah;�����;�O� y�e� k�
��ĸ ���J�?�w�0��*�rs������Ⱥ��A�*�_<F*"��k�QYp���:�����]��������;|��?� ��:���c�l�B�/��6� 4���ᒖ%��y������u׶|����?qߪb���1���C�]���?o�I��.ܗ�r` h�Z;�β����6��=��x�t��f~����eǘ�ﭢk�	RO����ިa�靓Ԭk`��\�-f2���#�W�>���~Z��#��}d��s�����؎�M*C~"���Co�T�l ��m �c���$�j^M�<�@ym��XH�i�:M�Zj(ݹ��*V7�c�Q|��|9G���V���G�*@�& �fX�$��#�_�Ԯ�w�!:� 1�xH~|#dv�\a�C�˚f����:1�xi��E��#��y��.�V�U ���J�����>��y��>S� ��{��q���HG;�r3<��Mϭ,�v@��MW둣9��)��SP��/�]cs�}��26q�ȫ�;�o�Qĺ��ψ&-Inw�&a��P��6� �� ;�x#D�֡fj琻��F{@dFs�%��G�P� �2ǡMnZrc���Q�Wh3���rQ�¼{���E+����j��GzV��9=�!zA�� ��0�,�yfe�/A�R��]���A�!��4�����qv�������T�����ʡ��SZ��%��=g�2�N�`Mf�ȉ96�%W�\���r�#�|~��:�k��P��s���C��c�x�yqF\��x���jfɜvc�x�E"��]�h�C�i���ɪ��N�үI�+��$���`��Z	��-��{�ݤ����J��o�@=��,��Ƚ���f��$�l��I�DL�]�{�N9�c��cƽS�K!�˕,F�a�@������Ь���O�i�ޭ/ �"������nA�@��pBN��]���a����eg����v/tV?�2Sf6�M33ENn@���?̱[�<��gU
���.�w�a� ���9�P�3��ۏ� ̮
Dl/p撨�[�X�!8��EȞ�PEH���A.@E67��Bg�V�����7�9&��џP�=�I�(a3��*)��I'):V�:.��/�ħ��|�"zdz�"R5%���W��]�Ђ��~c.����}I��ΒĒ!�50��u�k�%��yXU@�OǓ9~Ϯ����<�Q��T�&D� GTT���/�R�g�����n
'�e���)=i�m���Y��NK��0o�g'O��R�'DG�]JtH��M��]�+����*��ɴ��2EK3W�ǽ�@"��=�(�МRn���6_�Ӓ�*ý�L��&(i�׈�cт�(��/�:�����t�P�	�m�`�Dxy@_�������j���Z�pi��%kp�a���-����|���mg��X���f�_�2�x��SBR�^����n���u�İރ/c�G�����%���ǃ�3�>�PĿ��p�Bf�" �)ZX_eX�8x�Fcj��7�Tݓh?k2ᑄ�+X$�1�=J�1�N@�ܙ��Z)c��Zm���V3��e:$
��g�S�������������U��9J�H��]p�=Sa�^0�U�5:\�RM�^p�N�j�z������b�5��s4���+i����Li�ƭ6�]^�Sn�pF�s�ȡ@�{!G�� �KJs �v�e�ԫ���%��V�&DlH�r��2��G>��9���b����p������3���K�(�&��D%�/���=7MWhU��ajϬ��kk^z��'��B��
��49W>ܴ������@g�/Ψ�^+>b�j�(d.֎���wQ���<������d.u��f��:f��Q�g\kaJ�aȘZV6��X�0/AQ&�ϬR
�5���t$n�VKH���N���Fҷ[%%Ζ8j�'_ӧ�+p�,�6}!�e���D ܽ��y{��f^b�F<��&Rp��ׄb��D���>V�X1E��G���ܳ��
[$a����x0��ᆓ��� o���U�|I�&��)'��E���]4	�;7K��@���O�9 0�֖��{QW�e��8�g�D	.KgŁ���$�qi���	�]�۾�㧤W��?�Ք���g�[�v~2�H���$4�l�y:͗>�mќ�-�~z/�Ų����v�"�;d�s�e\���nՍ'q�B�Ϙ�;La�G�_s5T0�����@{^���k4۸�|�{�ysL�a��(���Os��:B��ɴ�&���Z��}pm�;@�'�����R�K�q�� ���F�9rV�P]aO��ͦ���#�o��;��#���]�C��#��H���h��E��$d��
ذ*�)�;"Ug �衘�c�
�>�X����E^U��g�}��qR�<ꊌ�� M�O�v�空w�-�� M��|�]-O�i�"ː~�L��;7��)~ă�j��	����-`��zjP��5d��G�Q"���(\�-�s]0v��,H,��'�� F*���A�� ��7���8���h�_9��Amף7t&^)ע���,�MK+ű�f��X�*��,��i����Fχ���>�J5ܱ��lkbf?>���Ðe�ѽ_�����]���J�9�^3�a���TE{n��FcY��Ҝ]��9�"�o%EJ�e0�D�"Yl�1ooo�Zܻ�\(FN�C���r0�-fs�"'bD�V  �$�\�&�����(�Bu�������w+3�u(c唴B�+�Ԁ���6��`<����LV���{�YY`���Ur�����`T�nS�4'nn�P�D|��w��3�M#4n�&�s6�D�)e�	j��NS��fps��c���q�/	�����=g�������j��5ͼ��;�1>m�*�~֠�pYE�/�p&3�I�X�.�a�������,�͒�H�%mQYR0C�S W�����aʤ�mm��L0ؠ��q�ʿ5��i�(LV
aG_͛~�?�۠��U���n+��W{-W�sNF���\O���)��h��%X�p{q�b�;��=�hsH�����۳�Bf�g���M����+4���\}�Jyﮧ��p�_�ö*])��q�ҁ��e�
5�X>�����]�� �+�ew��P��O��^�@H�.u��މ�6z�߳�O��+n��������[W���)�IsD�q�heHi��%���w�9��'1��:��B`�P�2����4FS�8]$4b0���p�Y+j]X=�A�E�V��Zq����r4J���%�࿫�r�*;Rl�����E~��P���G�p-0ͩ���|��rr�U�f�=��K~�:�(ln��]�V0.��t�p�=�fG�`�!υ�S��˥�T�l��G?��w�+04.
.̗��y���J���Y&�m�Yx������9���٧!�T���!��5����T��ҡ�\����e���s��5�w٬Z)�Hn��VIܿ]�+������67i�͢�<�H� l�>���)���9r�A�~�]�5�[v��ڻ[�\\6k?��S Ȳ�4�q"��a��o;��E=��ñN;�����8�=��lȚ1�ȩz_<.=}��MM�E��8�I�޺�%�Qh4���<�:%E���]��q�����VX^(d��OĨ:�l1��<����ga3
M~3�F���/)�%Ta&� ��JB%�ឨ�G��Ew�}��NV���*@�)�����-����]u]S���m���p!�f0�[]�#����`��EN Uuq��f,���R��X��7ub�0��8�3���:Q�a|���@��!�H�b�h*M���N�I�P�Z[_ʛZ�����?�%����s���P��fD�;1�#Hݛ�Z_-U���&ҷ�+,����W����<���54��w�@�-���y��G�(E��qo7"������~�%qMU�e�|���Njد�j�(��6��z����(2�)�%H�~c>O��pXu���m8�4,OE�sb�r辬����z+�|�6���ٶF �������F�K��T@lp�"���r�mR�]�&���g}��\�B��R�84Zb���#���pMX"8��Q�g;_��.Wm@���ǞT?g���v�aV�^m|����mȌޓ��Ʃ��Z�Z&�j.�Lj��;p(Ζ���~���ދM�j��>px�X��J�8*4e��FEo�`���*0��ت�Ď���()���$!pt���b����� �k6'2��*��L����g�4ܖ<k�;�?�=(�`5�rԡ�3�7~�C���Y���YY���@9�����եQ���Uz>��ы��]ۆw"�C
���e�q<���0��Q���� 0,����;v�^(�ZX�|[��2�)js�z�R_ok�cI���{�����`�����#�jQ7%; ��q�������?]�*|vE/sz[��}� �B��%Ӝ}֫�9�uA3@�796ల[Z��
��ys�l��ß�W�� ^�,_:"D��&d��n�1�/����7͛x@�K��tP4wu�Q��9"]�E�9��+�s�P0 4�}Q��I����?-�i���=�0����Xi6|}��S� @ڎ�AT)V�>c��dD�C���ΌR�ӫ��F�E�o2�0�����r����2w
�V5	P�3�1Ax�)O+E�ia	~��׼H��;6�劉�=In/��� ��q�עǵҜ����1	���q�@�����ÿ,� "��ɻ���tZɋ��׽6?�ݕ��Y�(u��
�#�HnN����`�5�)�cs@�B�=}	��s��.��iC�H�st "����epz~.zD�7��d�@��\Kgl�1m�ᩀ����g
�����-���t%����T̽ ���	�}�n(�!�mux��Z���ł�h�:�]�],,2�Pr��t���A� X��t6�+��]�wf/ٗ���$�?�憦+Ű���t�f*Vѩ��9��}��[���>N���UCbC��Er���ޯ�[?�R�����>��_y������<p=�������\��8�OL^%4ℬ������W�2p)�=�ྦH<�EF�'��=X�����9�K.��9�Р��SG�`�l�kEJ��+
,��~tK���T���55�<��~m�yu,�����z��[u}�5je�Q�ލ����]��5�1G�V�)�\Od����0��n�#D)
#o����)�CA������O�>T���!2��]Rߦ"/깪� \E�pB����v�Wx�s#�W#�L�R�9m+�������ى���em��p�Oݺ�;��^xN���ֶQ4Q#ĉ�D��T���h�mk|b�g�|�i%rc�E�$Ǝ��S�L��ʨ>9����"uX����h�,�����w|�Оz=����fWW������5N@�[M���)�7;n{)$�(E	>G�af������G+���^�R�C������ !�	]<�VY|��]�ȰhE�c~�0`����@��,D����{�k��*���k8��7�,��L�?. �w�]ocm\�Ϩ�' Պ���rB��#RC�(�+�C*��]0gX�k/m��|�xL�k�E�A��0RF�11��~d\Ղ5U���,�NI�2[�*���1��10Y��JS�3.3: yW�FNd����X��ֆw�Z�M;PM#��$
�Z (�G�<~�!�=����^�xd�U�JG����+���O�ɳR�?ҵ�^�x�͗Xth����4*=�~ii��W-��ޗ����S�yKI�p��u��]�f	3���.1�Ꙁ�ik^�@vI��Cε�yoUJbԶ�rh&�&���9CD s�P��)?��8��BSU���������E���d�4�d7�l���~���sR�Q�6����sf���F��B3F���$�/{nDwa%��g`��w�QI� ��o�C���$����a�����.a�b � ��֓�tN��"4Fr��5���S�X��� �]��D}K;� n�&�T?j$/�K۾�1�������Fg"X��+&��� ?-�_�s!eS���M0fF���g=��a���\���zV�D~��<.c��ׯ�i�%�AK�c?ΎT��B�� 2�"�&�j�T�FPE�������y�n�v7����k.��
c�x�t}���?"�.������f6*���n=�m��8�gE���E����K����2�/�D��+a�W���Z�x\�3(ތ�ڝ:B)q�ѓw��63�\���8�~X�+D�jԣDw'(���9��nv=k�8�a
:8��|�}Gx ��C�us�@ٳGO�?bD�+qo� ��p}A��ǉ�Ӝ9�}%a�o))Ͽ������)羸�1����rNZ.%I
�C��5�2�FJj5���+)��V�����8��G:帜ը�\�������in�ٹZ�I��0���|'��d��85�x����5�;�����ߌ"rUМ���0��	/7�$�rbSaѽ�0��uD��2�.ĵZ{'�S��O�<p�'ʯmla�n����YĆ��^d����s��F+9ݙX�]|���N8#�ml�<��o64�g_iI�#��A�rp��f��#��;`�	@��S��Qp�%�ҁ�������:���M��	���~?���c�	=�03.�`��'��h7p�\�lǈd��m:�~�#����n�w3�ь�p�Z$�̍��&�^�s�%�b& �C��`�?y�q�([���"c��劌T"���Rඝ)Hqm��=�t�%޷�Ϝ�"��;u��� +��ئ3CsT���;���W
vrc/M���'b�^�T�z�[�MK�t^�3�q�t��.)u����}}���#1mg)���#�An�{eu�&(8w��� �d�4u~/�4�_��)�oρ.�k����L4�&��������f�ʄ���O�qq���JǅaA�dL-�!���>��G�h���$ΪZz_i���S�u�o]6�;ȁ���-�Oƾ��%ci��i>?%���E���c5L���By5pM$���.��m�2���%����J)0�h$�m_%Vc�:A��*�ؚ�,��,c��!ۮ���3�L�T>��ǿ��x�}F[�l�
���[����cU�J�����,!@JX��VJ҃��}�)0���S]�f��7m8�i�"�H&��q�q [�j�~y�e=�)����)��e�|{S���\�v&�4d�c���9���P�e�D+G[��O�^�[i
*E\�>�4쯲^�FZ�)	l`%}�յK��hfQ%�I��~S��TZ<BW�&��Wj��P���T~��=(��	}ߢ*Z�t���$@�@��跌�K��U��e�����L�l@�� )#ޢ�������Â�h2������d{J�������#���P�yDߋ&ݽ]�]�o�K�g|�IhQ��)��
�{���P�	>8"�?z�)3���������8i��Vo/�p?�~C����P�����k42�׍�L:����>jh+�͎p�ǧ|џ �:;o���Q_�Y�7�0�#�h4c/)�_	g�O髯����yO��Rv/��F��b2)">O�ф�t�q*ܞ�����eP�t�����E��:m��ib����/��F�p뭑�
r�����N��y��lk��SX�j�A�t�	���L�C��A���T�
�M��"P����όxX\'�;��C�0{����ͻ�,��@y�uc�\|�C}xؕ�1k�V�#h��[0��O�k��>I4T�7�&���$�|�(�@�E%_P��i}Ӵ���۝�,V���v����X���u٩,n��;��G�]T��N�"e���RP�1lsDE������G];��zr��+������֜G���j5��i�@PK$�Xqe��c��"���$,���N�t�ƀ~�$Z�Y��ܖ�dc��9�C<���A��D΅i7����ֆ��@a���Y�%.z-^�$��7�^���)еY��(���C��mY��\$�<
��x���dVk%)b3�Ѵ��{��k4��ݳ��%��X�1���*�C��>>
Ӄ3�z�S��?��L5�{&v	���ʏ�Br��k>�Ը���������Jk�N�}5��6�Lhb*��msmy�H�$�R��� �l$ք�w��%��ύ@d�(�0�8�-�ֳ�L5���GB,8��?������B��/����02k�v�/�����Mm�k"��i���XuBp��N.�lkrB���OxcS��ҥ � ���� �n�6UT��C�e�+��#�@�� T���r���K��m%��T?�V�6c��q-0��h�F�ǎ�NQ�NT+�k~�5O=Gaa� ����vS5�c�C����\OG2�(��x��e*��I�^X�5�>�ԥ^ϓײ��aw4?����%�;����k7d  qA������4�DD�yw(�d��t�z�����]�ɣ L��Nh��E+�y�͠䨋�?��?=�>�}���3S��<���7�y��-h���K����Y��� ��?��-�+��ɾ+W�`��HЄ
�@lp��N�(�@��U��fУ�����9:�$B�K$��vϝ-f�3u&Y|�?øګ@~���~��S��.e\�S�����pR�v&��3?�2�B,N�(�m�JVt?�7�M�F�L��L�2.�H�פS���.}�BZKږ��ܿ8��!�a�L�p�8�Vq՘R0U�c���ÐS^�:������:��x`it���c̥ܰ�俋�&5_�:�FFm'�?�����ܩ��9x��>S@O���(� ��O.; �z�̙�a^�KY��_0Ye����d2l&X Z�^^�ǡ���v9y͟D�7r��n$o�_x��ޅ�@s�_+�A1���D|` ��SMܘ���<=Us�-㠋{��,���\X��`���ҽ"����4tJ������[k�mʆ�|a�����a�'�U����ec�sɴH�)D���w�!;m��J�uY��$�d�����9��]�$)LE7�Wn�C݌�~>�V�"���F��ݥ���/���'% 4��O�o^�?�%�8n�Jv5�w=������y�`�K8�vTY{�ڸdy�'�c�A��4�۹I�;�f_�l��nIZ�[��lKǠ��5�O�W�}�|��&lsf�	F�v�W��/W��!C��݂N�]�}�0>����'c�H�϶����m�Ű�
3i��e�� #K�(d�Hc����­�
M���+l^of�^۷_�"$��4h�����*���豋����>d�ה���	h�gM�=N�A�^��o�]O0�����{�=����IJJ]���6�+Ex�N��ق'�87��{�l��>��{�^�~�D�<5���w�V���.kT�����@OW:��{��hr��3�Mʕ
����gu������:5�?4I4���
3��2��i9U8�e�W�4���@j�!�N�|�L�r������e�[}���R�^�#�9�p;F#����F���>w�xG␔y�}�	�K)�%39!<m���63�^+��N&�p���Me#��\}��AM�!Sp�J�Me�7�����s8c<<�$�M�}(dc�z��ɶ��XN��2\]�R��W�啁
����������Rʴv�5 �Ɛ,_R�G
�;�8�-�뜤Sw�P����=�6=V,jөW�;�R��!�C��'��ݓ���j�~t�D,Vi?�l�rݣ`������ Ɛ��6�34��j
,O����+Y�������k��[��V^geU@>����l�g]���g�[0ٷ�������_
^�P��� ��#Lq����[��fy}��C��
�(�W�ț*�x�d��L�2�sOѹ��v��N�f��y7W��|����t�=/�/�����>[�~��x�)��o�$MW���G�[�a ��x
8�$�i�Wn�W������H�����I��������%8z\���S��Z�P�jց���Зg��/G�+K������Α�l��~�`�U�k�7�
�����\ !��#���#X�����WJ�h��e��[6������������/�࢚2|�o�H��Sq��%�!@I�`��KMA��?�7eCo4W�1�D�);	|�(X�(LaY��`�AZҩN6��=�o��T|�1�������w����삑r��ۋR�{͝������7���x�4�شϓv>�mlG�'>�3Ө�Ϩ�(K��\Dlc�b�b�(���l��������Z%�j4�tl}u��.b �g?U _�iX�3a��2o��@ǲ]��F�X��*��ի�I��s�|��J��K�o�-Kʁ��h!�>�̦�}�yF�ݾ6Gr:nFs�VxH
S�v��!܏����}HP�fD!�>~à�{.W}|U	�`	�U.,���SY���lF�thۉ?=��|X�%3�1JI�qX����iDn�v&
�K��C�z��.�b�����s�]Իrv6����$���+Zk���թ?� 5�o�.��l	��pm;7���z��zJ��x�8eU-aME1<^�b��&]G�I�����4u8��Eq�7�y�����%ZG��m���Ka��@A
O{��é�Ӂ�M�So�2.A�ɑ���1���<���!��IJ���/:�0-/���gkC9Jg�Qp�
I�t����f��`��������=��9[��z
S��^���ݪ-￧�"��Ҙ�7!B�w�s�F��iѱ�~�J+#\c�k꧸�V����X>iɉ`���g!r��6�<%��������� �9c��lxH3o�kkG�h�EP5*�D���ʿ�Nu?~�� v����g!�����!�6��.@~��oC�R���0�Fɟ���sj$QV��5U�k�2��V<�EV;6��Uщ�H6xL���o�|��K`'��<1�m���r��p�o]99k7��?�M�z��� e�<�3�˦?/�9����my��᷼X��d q�<���@��N
��U�x�r@���'#J횅Cj0�p�*1`j"�getNX��τk�v�����������(������z$Z�Ѵ�Q,��k��n�;#/EjC�d���9��@
M�c�]n��9�����&m�Yt�B��>���v�^��ö�q"u5��4�(@G�k�9�.�w��F����@�	�P��\E�KZ[�܆7��0'lE!��/��7�-��wר5~�S�fS�a.ؓ�i�Y�K������)H���hv96�L5h���Û�xcF�!9��s�0��#L�i����';�2�I(�s��.2��]:A�x	�!O� �y�;(�̀-L���iI�#-���me(4�0(J�0RG�d>�c�ּ�v� ��M����x�֞�Z?�m�UrhR3�1_�仾����O�t���*���Q����=i�W��s�{<S�������������,Q!*�����Ϋ�)X��J\�es����J &��YR0��xUv��'�|}a���ܖ�ً���M��40?���~b�ؖ��%u)�`©hf+냒OO��L�I@/:4V�$�O���R�\L�⢱���v�U�ʹ�T�Nދ��L��
@C�r@l��V�Y�~�C�@��˸O���Ǆ" � ���.�"�� �|�׻!�Qݾ˝+f�����!�{�ѵl�R2�"s�b���+�0p[=$#@�RsR�A��V�M\ONW޿l��-1��n|uۚP������8��ŉ��\�����x�hs��6@�|p&�g�� [��+>���kg��	�R�]���[-�l2m�P�Jq7t�WXk�ZP<u�O��#UV�fz��Ύ�3۾��7��2��}�2T�x�;�_Zn6�N�7&x���eiύ1M�2ժb�t���tdv�%EwLMHT}yr�F8X������o�ҋ�vNc|� {�	8Nƍr�B1�vK��y!v�Ӭ��b3C0�cUzl�)rY8��t&}�Z�#�=i�i��`�,��ݕ�xB�#�|M��7� =yϝ#Xi����3@��cv�	�uG�7d����U�	ԍ��ݕ���{�h�"�e��`;Y����;(�L�cL�mƮm�*�d+W�@�N�y�˝��^o��g������$j��Ѿw������|u�
E��G⋳�u� �������es]�%&@.G�s��	�$٭�V�u|�D$��2��b(���� �l����o'u�6�O��u�:���6[B��D������+yS�;��7n��s���jQyfn����sR�{�,��4�01��6���O;Ņ��2f*��O��&��8)]��N�x�9���V+�[:�3�[��sǀ���y���k��([b��k�sE��d~Kß2'��h$����Wr��Q5��\3%F z���J�)T�o��I�C
��X����ZFS�3F���F�v��0����q������s�zߗ$�qգM="R����Ȧ�C�Yu>�z@Y6.&�at�r9^�Rk�.�tky�]}��@����{M@����㉽��a�X'~|l�V>�^�+i���W��?W�؝^q|EH��٩l�� -����_e+������e����>�O>�b:jo�r��s?�$�'�d�]s�l~+��N���l�oѐ�64xV��L��Y:2py�
��n�a�n��j5�"	��[og�Us������e�V�Y�M�q�]�\9ħ�d��������ףF�
�7b"���|��d�L]��,�+�{�|A��5����W�p�� ��:c�ףƁ����R���ͧ�g�����ux���k���^�����'/:x~X�#m��;��ى�n`�.8'9I��@�'����0�1y�V3���m��}8�<�U/tN�q�-�Ϧ��R����ɡ�S�bBq4j �8���{�~/�|~����h�a�k���Ȝmb'���Ypx���d���.��P��1L��b+��Y�6^���b����Ŗ�2R6~UV�KVˢ�y���j�C/�����qw��u���-8�H��Z��a�ʝ�)��Ū�O�.i@	�����@���!R��Ew��6�v��9�L���aK�6H�e����r�����Iy�ʊ$)�����~/�R����ޠ�m$���`5O�aP��92��(W�o�O$���I��9�]b���{c"����n��P>TWR��� �C	��>����R��n�HV(jy��nuv���B�Y��kd��4Y��m3� ��(�����l�Ԟ��v���i=��B����JU�����;:���(!�#iK�8���<K��˴�E��T���yE�%����P�M���] ��_qnI�F��|� @�M1a�%�b>�̇Z.yC��t\T�!�1m��D�.����+F0�yY%��6\<�>�L���i�e*�oHꂜ`�����
� ��
+�}�b��H�#��K�gjgT��Sm�`�.��2NZr�x��?E���3Ɯ����ظssJ���K�	��]�w]k��C��C
�0�Xy�_S����b֢��0�rs��g��1���w�H��:��U�Z�3^��V�Z���mojC��n
��S��L���X��] jc6/w	� F/�.���yq���X[W��E��)Cv|0����|���[2Sᴾ�C��M\F��u[W�[Hny��ꪉ��D���s�d��'�0*v����.��"%Xʔ�����B�/*'���a
�r��4��:�TF� ,�x�(�����9�=���(� 3K��@����~C*���FL����p�&�|����H҈��e����Ʃ��
���pP�eR����JF�T hlR�T�7��E�_l|��	�Ø8��rx�.���Ĳ�C�-L�LI8�:	w�h�^5�$�Bx�Z"�c�Ś����Y���T`Q�8�$��LU���P��%�I.Rh׹׳�	aX�7F�֦�B&f�~�c�c�����������r�P�&k���������e��U���V���;�]�<_x�{�&�~� [q�^#A�L�$ ��4�,]*;z���V+�W.��vX]E� 2�W�(5�'��&]JKΟA��5�I����v��Eؑo���!Q�d���_�%%���l��!K�k�ʮb�?26$O��<����
�����+/Dޙ$���gs���AS���[ͩ�	&�q�)���>�j*��9�`�#m
m�Tqv*Ѫ�z���(�p3�1��G��_�ۤ�s-r���G"d�z!k�
������~�IOP�������x�D��k���0�`���!_���-kwh�4M+�#o��d��o%h�ҜB��&Շ4�9���!��5���?l��?�ir���h�W�&��N�� .[���a��6�a�f8�32��2��Ր)�w̿Ne�dq�O?^d�l�E=Ф�u� �5���qe���W	\r��j�ʗu#���}�V�<�vj
���u�|�4��]��� 	Rs�����u �����F��J��|Ŧ'���:Ċ�wK�w+�A9������@���PP럸�όGV�CE��e����{�c����kN��B�t��:)���&��민Wt�>��T��I6a��.�����#I��\xV9��em���F۹���|W`���j�k�.�胸'���4Ȩ�Rj��f^��) 2sWf��?�8��'�&r�z���b�9uPꇱN�$$�8�{��L�ȧ�����%���_�����\�ܕ��nt�R&����?�f�O�����?sr�g���:���h�)d%��pWQ���:��=�m��V*x���^�!A���HN�����
�,߂�ykA?lx*C�qb��j��O�_Ӗ~G��#ynk�dr�Y"�N����Ӯ*W*,�4	{ѹa:�5��W��H��L[|�q1�o4�&3u���9�y�n
��=�aw��4��
�(���87A���Vۋ��u�l��UD?D֗9y��8���].�$�:+Vd��W�b-���02���(�Jࡹ?�85���Ѹ��M� �N�3t���1�<���c�INE�[,�����W3 +5��k�l�	��@zV��&��y�~�_��V�C�����j���@��p�@�X~�o�J5�3uΝ�e ����:��x-|H!Z�Q�n*IXĎps�s��L
ey������aХ������	���T��M�-�h�s�|�Y�b�Z�j�k��\!�z��F룬�?��� ��ϧ WK�+��Ǒ�<���'�a&����F���^x8����P+
0�� �A��p>	�55S�ⅅ�S�U��pf�<:  �%q�J�b�n��k���?�M����F������{� �'԰��*�{�ED.e|U'��^<^'��������䔕�fko��Ǟ��{��1����
ݳ/�=B�ׂˋC �&�I8�dIB�h��/�j�ob�W��v2�����W~����Q����߹*~�b��G�qp !���i�Cr���9.b2�O����`ɫ�l�	(��Sn�*���%�}� 5=i�d(�~͟ߕ����@ر�T/I�m������^��_e���� ���Mq����G�<�Mc5+_��h�7�;>�ك�ď�*�^>�!]q)%� �i�y����J�i���?��ѳ�@�|�+{�`���k�hÀDu�#�������kr�b��U1q8�������Ihr���̧l^K20t7&���ZiM�쀣#'W�ڥh��[�Y��L��۞�1@qdz}����.����23�0uS�;�ESb^�V�Z����^wSw	Q
N`�E��ʑ�N�S�Ѿ��䟆{]�T:UCC}�b�DC�yS��Ї?�$sOZW�IC���vYS\pEf�b���#Jǒ˥0|��k��2.��O�#� �68�$�#������u�E�xt�6��}WOl$�Ϗ �T,���+����r�����W���)a>�/����wK�%��p�?6I���q����"A[�֔���16ѳE���0_oS��� �Ҿ���Աd�z�f@�qCT����m,�j/'!�8/4mۙ��w�^��K���qmd��3�k� m@��SQ��eQ00��V�z�������Ю<c-?�[�.�`��e�P�`Ih�H��=т��ذX&�o�3����n�n)B"%�Q� ُ8�ۥ�X��_<üA�L2�uۿ5,7Gl����_���ӧ`� NT�2�ؽ�WK��1 �ȭø���p��\��ɢq�ɭ���y9pфsM��\ �
̢�*(m���d�yV�T����,��u�rV�Fn�|v�}
f�YW0��h�³(E-�)�]����$ט@WO������}�.z
���������$=��1=���vF�Ń��P��5E8IB�c�� �z���-䌏:��.�NG�3��I]��*�� ɯc�S�bƲ�(�{;zڞ��j�ԅ����YJ>W>CPx�51�+�ߚ�S�M��"���|*^�����t�,x"�ydY��[��ߕ��Pp2��[]���g��������p 
$U�F�W�y������&X5�8�-����+���-7��%�d@�7s��U��0�6�Km�������d�������V�Hav�&�C>XLaP��]P�@��̉�3�\�|��tS֫�F� ��S�qH&�� �MH�AJ���|n}O��6��z�d��`Ge�j�x�A��ߡֿ�!�x�MN'��H��:��� _>-�&��x�{<L���ˊ�]�Xzkz���!�1�S��@��9���/������D�T�Q�&��y����l�یV�e1Z"�	�lª.HG�������;��߼N�m��t&i��8��0%{w�ᱍ��1S�(��	 ��|\�!|��� �$T$w-+��$�A{gO���l} c�����ph8t���|���ў��e�ǖ?��~㜳�s隲Zj�z'����� [�ڏ�χ��pN��q��Q�H��j����a�^��D��CdM����kZGVX�b�Q�:���\����hvE�EOo�
�f��ު�e[z����u~Y/�.B}��	��w�3�y��`��D�K��O]��Sf��>�:��,Q��
�EE~��y#�J�AV�Ĭ
��t-������&kU�0��*e���yA`��r��e[)gU^�h�&�o�]q�r-zU��#�ǽ�n�Zg��p�loԚ����(�u�P���)�c��} ���Q�R~����Oo�{d��5��sR�CuIb���;�n1^���D;%������pJ��Fs>9�����k *�b������Od��?{�!&a�ZV���A���}��
����A��y�B���u��^j�Z��a�q�?���l)M�ƞ�رr��[���<h \0���Ъ�p�.�^q/���)$��0�m�/�Y�S�}LJ�6}E9�G��t�b��^�!0~�AW���{�T��(O�E�5hyĜ���%����;A�k��8�T�dc���@"G�����(�-9M&A�^�r�G
\��cK���	k��Z�+=�S�7�}�+|-(Ru&���������HЏ��KK�-O��0'�k����XU��i=��i;�N{!��ϴK�+w|��"��/,��Ն����ރ9EG��6,������BǠa�}.���kREa�x.�OnbJ`]:(�V���T�S*gn6�{�نU?a3��vHYL�v��E�D
L�f���Aj���΍��[zxk�u�6F��;��������6����@�;C���?c�̚(h��Dz����r���~�����0Y�B>�P9�m�娐��i�3-�ᯥ����3w,-�<?�dk5?G=>p cR� �6�9po��Mp�u���vlo�`����e��3
1�*�j�oQa��k���[�F�42q�C���y���6"K���8+�}e��Q�I�E4�$���حôٯi&�W��.�lx2wpk��w"V�u�0{x59G��&�����QYC}���^�ƌ���s�ej��T�:̏B�Zȕl���Kgv�^��s���p�V�9���uϤ+������E�zg8�9�9 �r6�F�3�;��������g�J�#nK��[������au�IH���6K�˾�S`ih��U��qWʝ�=�jg0����+t�M�"��-��1�i�H���涼�&��(��	�b��&��~b��x!��蛀5�Ǒn�
��������¸��*H2�p��kkTړ�$��j�ܬ�Y�$��b.v���$��r)�o<Bq5OÓ����`��-?� ��2";쮤��:�}�>]��{������j�����6�"�F+�	5wt��g�~#!l���}�I�;��R2�
�R-�<�^���׾O�Tࡐ�_&�|b�6�,������� �i閉S�~֬Kuז?uIudN��i��a�:^�8M���؄U¥��K�нX���E���uH�[��hT�������Z�R�{s'Y0h��,&O�|I��q��f�PdPG�Mzy�Q5n!x��#�����|�Q�pr%-�^�}+dU�J��2��1�聂�y'0sG?;b%�V~�#�Ό�o
m~�d�(-".okS�'xMc��
��v3�ð��v����"*��������0o8�s�^�sZ'f����a�"$�Q�-�/Ÿ?�3<����QKBK�0��� @��p䍊`�뜰G|�j\����E�e�k��)m�4INv����5bPT//���{8?�*	5ը��I��B3-����L�� �����m�
m��%��y�������q��*NyF���S��d�6n�nvOh����2��Yv���@�d�Tt�DڀH1��^gS��aB��+Q� :���R�r�q'] �47う`1��K�ec���Rv�x��k,u���La�i ��!�sZ���p찗;�C���Z��zeָղ�N��'�g�'^�|��!p��t/�[/VG	IK�������cSk��<h��ļ���7�D��Ƣ�thL�"�O�j��{�Lm�g���w��cć(2=��`E4�5l]�C-��Lފ}	N[و�u�脾ޖ��m��G zA|�J̶X�jTcX��7r[9�:ix�"�zx=�����a��yLZ|/#��}���kO ��GH<A��xg`�q|j\1�l	�:�PIC$s���S��&w����򖡰��f(@o?�Gw�2kb���9�H�D~r�vIs|2B�W*�'�}L?u�$�� � �!��MG���k]�;��������EfʮRuڐei�62nD9�BD�G5р�V��?3R���<G�v��>��VsmW�M��vA�	���b�)����7ٴ���X�˥���n���q_��*��l�7A�-bY��7fM�6�"J��O�ǅ�d<&�)�P�g����{P��N's�z��mbn����(�Q������te/�@.g4�E���}����0/�ƕ�ʨ�3�i����_}IH�l�;7ɰ$�r�#t��5M���>��sRN7��
��w��D6�+)N���
�W�5x���:�	e�!6��*��#�q.5U-��(GX2h�ؖ�9�YX�y�a�u�b��qc��,%P���X��y�]Ԫ������p�~����֐�o<�'ٙ��,�3�[o��>��5��Ρ���d�{ſk�f�&l��\�}��簑��A�N�R\��� ��4�ʧ!�OX�fQ�=�l�c���'��>�/�4���ڦ%A�����WkL4�����p�C)U�od)� �k5�7�F[~�֏�42�1fT�v�`>��	-��`�2
e���=w,�ߎ+���N�� "�	緮���fZ�L�X�cp�m ��:������z�0<D��3�B�^l�+�y�jL\.�1eU����J�fJ�_�_q����VRX�S��q�Uռi�b�xU��5��r����M���T�]/wn����v�s��p �wlt�s;XOb/Ҩ�ta��ꝸ"�Z�/jϺ�eeƺ3|d���-��?�3����3nd�h��v��7�"p��N8�eH87HHD[b�Xs[ޫ���-�37��,�[N;.º"���ӹ�f$�!�-�#��*6�4P�=��΅U�F�2��L�)�1za��Y�#�Ϫ�r�Al��E(�?�SMX�Ey��/r|�����5%�u�x�ۡ��?�9S��@E]��m9[Ѽ��ȸ��ϩ��GM�~�E�Y���h�N�(�A����y%O���!Oͷ��ˤ�������xg)�wh�fV�PONӿ�
���VD�[5G:��̩��ы�2�/��� �Lp4-!��ln����X�~�=q&��\N��K��%Ζ@Q�8̉��yw����UL����#�:��g쫔�B�gc��?J�8��"��)$���8����.{F�_k�\�ACie=�+�&ܦ�Xq���U�����f�LYjV+N����n���l��%^w�ϛ�^.�߆��9U}
q�8G���P�`��r��ol�!�p�W$"��b��(7�}�6&�Y
�N����R��� �;�_�����"#���@���<�?�oz���$�'�*n��\��q�e���)��݃�������k�f%�>7qg�`����7�흄�O �T����r�Q �S���%��V���\F��Ru�>�h�֐c�O���Dֶ䯜5]���ԝ"߮�2�2X2rI\��=ě��5�2��,m�yd�PY(	d��-�K�����&�sֶ^.TsLP;d,�#�+�f0H� ��������$>{�a�|D2��t��,XڥJ�(�&4��ƌ%�cq5�+�������4���̧�We�\�/V �n#s����C��ǧ�Ch��`��#���(�EbgK/AP��Z��F:��1���� u�K�@?9V��7=�a�3Ak���K��Jt���Գ��~p�T�Q X�`�]�m���R �5?�u��������x ��:{�r�k]��=|Xb\,<�������-� �+߲D�J��gFј��6�]A�� [�ee���s�X�
 D}�;	7�0���>�344ðH�}��Tlt-)_��y��z7Z�������[���|�\���&[j��C�DLnͼ5�Pa>�\Y�	��ԁ��JSٍ��!�J%�?TKɆ0[4�B!˝b�,|��	�*tS���>��M�Z�o�
��a��:���+^Jvh�=nNR������&á ��YhCq+h�<;4s�B?�1��{_'y�l��gg�0 �U'�{��fB-c�uD�$��Y�y2&��A��>��A��(�oR�Q��!|���w�R�����0f�%���p�8���X�Vdz��Ty]�-sc���C���xl���!�#�� k,����Tb���^�C�Q;�[��=��c�\��$��kS��F��ذ:m�D{�A��Ů�Լ�4��2�	�Ceȧ�8�&��]
J(ii' ��M ��Id5/:x����;dG���B�Z�=��d�3"&�\VL��SP�#\,�3��)yzΰ�a$��L'�\u�s��Q8��0�ĚMd��a�9X�ߔ�E�2ΥC�%�ez<�����L��CB�=���@�I`�W~�g����1 ��J�캧Eߺ��vFWa6��`�Ѷ\ӗ�̶V�A]� �[�V�
�h�lМ���#����K�h_�i��ռl�63�z!
�{��3alQ��g3��D���h���i=���5K����xd�P��{�k7��H	��z����
ؼ��7��oŭ��m�7��⺧�꧱��č��hBZ��Mb�O�l���s��5'���S��qx��H��нD����9�\cn��Oۨk��Ǌ�b%]������w532��N��3�� �k�Շ�k����r�`)/��Z$5�j��}묃��*0���+в
��|禖N�����RpB��+�	�եJ$�5TYK���n�%^����r:�'](�w����� �l�bX'ִlAǛf$�i��,�lf�`�����z:�8��"�IY�̢��z�7��~�B��]�kx�kgxm7���yЛ�=Go�Mb�1)�bT�"�]����L��a�сΩ�D��F�߸O)���( )�\�n��m�{�­֛2�7��Ps�(Kԩ����H[H/��~hYV�Hn�u�[�'Oe�8�OYͫ�D�;ؘ�H�����<@2!��0�h6�����D���4c���m֘@5.��f������_���5��� �����.��1�]�Ct�+��eٶM���U�򚴇$�zMk��6ē�1hX�I	��"=�=�C$$$�YǍ2���##ҵ9�N��,�>��ulciZ�5��ߨ���^~MR=��t�]΀�Ü��K�?jZ�2(���;�X�M�Q9�Y�j2YV9,�ܡ�5�
2&�����Na���3�*�W�j��G͝Գ�n{�?���/q�i�L|×)�O�N.Ϊ���b��=����2s0��X@j) �1o�.�M�Y�gv��a]&�<��f;��v��+�ؗ/�n�->���x̑�M��ߩ���q3E��M�v��F*o
�V���g;򾝤��<2sf<ʆ=c�-��U����3�����P�h�M*��,�ڷ}̪_no8{F��Z��J�5wL��
�w���2Lk���@"�f����QLƐx�S��h�g}є7��F+�F�-P8A
L�1R�&-�	5(=��VdM��"�!Q��([[�o��$�o����(��b�{~�&��D�?c�[�>42K�v��V3W�Ѐb5��:��k�#��!��2���P��	�KHs(���i��f�?x�ܧe}�
������R�:��n%[���?�9*U��|ڥ����
j�֭+�W����8�-��V�B䘲�g���.w,�.�E�;����;-�O|s�a�R��wyem�Ѣg[Z�����m�,��c�C�m���[��� 䢟"�+ND��N�C�?�x�3��������1׌Jަ��:�N���?�e������fx��L�L��C��@?+�����ZQ H�p���bB(Bic|Q�7�u�@z���C�{�
 ��)َ�P;��F�Y���uq�0���������5rz9we��k�'�/BÇ�]IGR+�ݡЩ���+AxG�|ͱ����H��ퟍx4�F� 
�˷�
4��m"�^��+��"��<&�����y�Bq��H�jMdSd8�LSe�R�(%k�����?�!P�`�*�L�^�Ŝ������w�����tg�q��|j?���R,�����]�㓴u��^S f��km��{WB�@!GfG/-��a���������A2�#�2��A\:���=:��ռ`B�t�@��!X��Q���,���R�ў#W|���&Z�m�
�irʈB�X�w�P���\��s$
��?����)��^1��EYv���P>ً���ޢfoN9�HX�QA)8v�!.�Ú����X:aH���2�/f�[���{%p���n�u�}�FP8�2�O��笖��?�$�� �qإ��u���|(�	�.��L�8�ӭ{�̚,���C�������,壖�ء��!�-c#a�	uԛ��n �BJ��«_�Цưl�0P�e��f$%W4{�,�ܰ�*Cᇦ�1�Z3/�Bx��~|��t �	�-қ̀��hն�WJ'	o��S�%!;�<��J�z�Y)���@�%G��l�ބ�\Y��362V���3���k��*����4����.�Zr���I�6����;��gn�D�n��썽敡)I�.l߼%+c�ڦW���9�S��<�ߛ���fB3���.E�'��D)�
[T+vt�z�	xZ�z�c{N����PE|.�^�[P��MO���UFPY�Q�*�&tO�yŨ�=Tz����j��j���B��\w����E\�旤��V��0��������=�@M��@�R����drR:l�K���1:��.z�E/Ӊ�im�	�Cfv� ̯��e%�Hpr}]�wN ����̵R��p|���_KvRK���\P��(͟��9��ٻ\���oķH��5)���w�KY*%i�B�K���έ�ܯ�M�wy�p��n߯��c�kDMg����n�ث"U�d���b����0t r����� ��#�+�&��������Z�q�,dҺr3�Ǯ��/#�g�u��e\;^_g�p�ZdBTTt������>dMWpkbӠ�+���i��>��LK%�G� ?��~E��Fr����S}E��L!�<��s�3r�5����℃)��֭�b ��!9��%l�I��M�T
se`{��p��1�m#��:D�U�jg� �A�YW��1ϡQ|GP�&F+.��OD%W5���T  � �X]�
W�ҼSl��U�Y��l\��{�,8ڂJ`� �G4���y�#S�jʶZ�"[����:f`�4D4�	��zU+��G�M!�p��7���,�)����{%�e4Q��&b��k*�y���l5&0=�J#�P|�Y���6�lG���S� ��j��
e�$��e%�'���>3��txm�j��U�$�f��5�u�GOx��^�Fn�*\�͵?�V��Y���~/YO����i*�1r1@7��L�yDλf�G>`l��&�����Ao>�\V		�nq�σV����I�UcK�=!Zش��/��9��G�e�{�@�9 Y�¯�����E�O%�aǏ��n�����b4��D�a�K����v�>��j�U�c<W�;��$��w���f�.�q���-��	�g%�Ov���1,��?=�K���_�3����I�����O)J��jOպ�@?0�qv��1�Uy�c��%3}I=���j��"�_hÀ�8ġ�wop�Bq��=8�ƻ�Ѷ��Aq��j�M�e�]�>��ٝ6[��|���v��kX�<y�,�22��fΤ=E���2�X��YحC�=���]�P�T�Q��Oqw��ꈿȐ��ܷ�GF$�I��k�hQ�~�Mx�]WZ!8"�2Tb���l�'	4�=w��~|�Y4�xXK̀�6�_��Z*�%qr�;wC�w0��*��bE*����cP�9Ś����'eӝ4�/�ʜ��ke]�BА�lO>_����p�Ғ��P>������UM�������b�,5��>�__,�+�q��jU�-=�1q7��S0.�3O�˪-�*{޼��"�!��J�}ϢG�1׈�p�E����H4�T���mĪo��M־�͓��'~��>W�ž,�i�O@�dO��)��>��_^f�L�@�И��~����dF�,c���H�����*=���s�ni��`uaog��r��5{|��F�-Ԙ�q�*_Y�X��m�)E eX��c�g!_M�&�vL،*ph�௹�1Y�2�+$�����:eZ���>,N����o?�M�&�;�-����TY�g�i�z�S�Poɺ�uSߥ�e�����߳�b�h�K����/9��ƹ�Ϡ�.��� I��,L&��d�H�X��m��^	��Y�}Idt��,�?E��8�7�*�=V~"�M@Jy��0���?x�L����V�ҩn��KɌ�fۤ���h��������5'~w�{i�݇�"�W��`��TrY��mt\p��jx�D���H��&ك�+��f`�1D�LW�X��BN�z��cl]n
��%6g!�%&NfᰗB/�~?M�}I�&ͷ�x��'�4ĨT�s!�z
�z��e���r%�Y��y�o[��&���(�0�<k����Jg�,����M6�U�
�\Y�7(�$�<� ��Y�[���h1�W�>����Qr�'/�J'`�� ��"�dL��W��if����l����Q1�����u���6�kY�P�a�%o|ֹ�]t�e��0)��X�����J�;��D�� 7N�>��Y ��M6�ȯ����c
�66�9 �T�vR&]w��ȥC?��H�F��:K5g�u�Fѕ������`�E��⹴"L���6�*&�0��
�<�t�]��S��ک���Qy�?�E��B��ax]�|��~��ij��sP�>,hwe0ͽ��io0[s����#�f@�x���U��
���>��1�<�gf�xʅ�+}�:�A;ܨ
-�ϒ�R�)��p2Vu��PKE{\qo�,5+�����濛0~��1��"~�l��U��#��D�g��3CC։���o̎�*v��2U��.ʵt�m@�z��	vb�ٹF�3lE����3@k�Zt���SY���9��;Ē��19<Gj���[]�:dd��l�W�V�|k�W�ZY�_����'��ڭ3*���De����q�1�w���8��F�F]�Sįk^��y�~Br�<�|�1	�]}[)v��	��� �>�Tw��="0xo��I+L�^AbV+)��z�Cs����������Q�ƍ��c[`���zxDq<�� ��,�ï��\�o�"վ�ֹ�)��Qſ��aOp�YT�ՙ=��+�*�<��4�� �5-S}:��C��
�<	6��t�sz�U;wV�*gЖ��P=#C;�$ Z�ǙnRִ��QLM�BR��7rh �ͽ�p��n[xؓ��w/?]y�L���8��ܞ��b�w �kv���7w���������1 ���,�����`��K^���U���b�����1������G�륎�9�qђ�1 �6.�UvJ_�>�� �K[3����E~��Rж!������X�,��_M��=A#�X���^��\ ��7#.:�u�/�2̥!'Q�PU�:�t�>�yUn��1g�>�����}ˤ�/rm ��^H���򙹯4�|�`F$�(S&M��&��T�V3�`�B�:��#΁�KX���nWľ�[}����4|K�	���zyd�,����jI�n���=z-v��C�'�bt=��L��_-Tx���̡<.�������G%<�0� �vyN��?�����-h��m~��/��*4c=�F�(7K�n�O0����v��Q[���WŴ�pU0O�=�UϙEVY��y������r��%c��2n�
�I�S�:و7 ����H����,<�+ m2�l�:��g��F�W_�Sq8��	5�q��K��-��G�xK
"j� ��$23v&�1%�*��^z�.��W&-<�?Mo�@�l.�%�q<�d2q�Sm/c�d����U��f�匿|l�E�U6Ӧ�˞j�.>(HE�v��#�䫝����x��Ij����p��ـ���M]�+��.1+U㤀����=�(s<��2Ua�����ef����Hض��fR+�%y�pC���c�B0�o�iH�)��N���5��`b�Ű�JW�UG�]܂��Q�Y��Ο=|�a��o$�7�$��u���W
c��Z�}��/k��!��"��n�?��ɍ-�� �"����`E�9���n�Uy�h��iL��]��6�pG��\ߙ�$���b�sغ���=|@����6('a�r�Lck�Tcw �p�;�<ޫ��ԕl�ϼ�,'[����*�^�
�}!H{�M��5Z�.Nmh��xD��"�XF�y��8�Ch*s<��"@������S� ��/���1�z�����t<kn+Re�p�������;{�&H�;"��q�?^�[���ۺ��'`�����gT����.��G��EP���"�4�Y�BZ`����iM5.��_���U`�1=ۍL�<tÉ4�@)�!$;�����d?��o��Ք.����Ͻ pL�SQuc}1��!y�[���l��W�L�&�g�f�!�x%X;/����a�ht?�?�����S�7���4�kU���%_٬��(0V<4�ɰt�=��D��!3�p?�2?�|VP�x��f3<��Q5��N�ĝT�QQD�dN
��5Y<<R-|}q�?@z�є��W�z�J�v��g��1Tc?f}*��)��Qc�~.FG'����42\��C����DzYŲA�'�u<�d��� #����a�E$#=W'^d��ol���Ӿ����[�VX�E0�� m�$KrF�<H.FP�DZ(N,��Z���~�m��k�j�
$\�3?�O�t��a���c���Iw�1�pҷ_��~	����2��#&�^�f!>M���&$a㍇n���=x��gA�u?ʥ�Xfc���3��5����!n�qp��y6yɑ���ݾ糵c���N���ذ�Y�K���xQ�G�x��$0[f۬/�sC'�=���a�`��ң3��Xk�qY�Ȗ�Xx��Z+�u�L�g��>�,�̮_˱T;��%�Kl��O��Md~�g��C.)���\�8Pƌ,��mw}�|q��������/��ܹm������n"��o�@`,�q"��畚$����8�D�F��n�<[f�Bs��:��Lr�rs@�8��1��=9ӊ��I�-�t��ywg�' wk�������z�`e�a%)���5]n�U�5�R���\�~"�&�	W�fj�|�Q�ą����_G������0C:I3b����;�mΛ��i"d>#�m:C�2\p�W)�k-��6QL��SǬ ��"�%i�PU�h��`P��q���:�tR��)mAs��@����LVI=�>�T_��O�=	*v)�e6G��p����'��v݄�V�������ˀ�����Ng�u��@,T���l'!��<<�*�B�v`(m��R�����;�S;L2V�E�g�H4盺Ⰶ����B=����pnE�}��e�y���'��N��Ӈm���R]��[[�i��Z��R�����|�8I'9�����
\�Y?Ĝ�zM(S��5f7rM�JB �mI2,*�ўd�����qԞ񌘌j���2����/�+PT�ε��*�՗��:')�p��dC��y)Op���MX}.fu	U=�+��r+��:}I�M�QG��/���V/*��c���/���3���G㴲k:`t�:�r:޾a%!Y?�t���ڌa(j�$�$���%K2Qg"���+ v���G�������4����j4�>N�T�	���m�t$�"�ʍ�r!�M���c萗m x潶1|A��z��*R{�"�?��cV�pƯ�~���>:?���{��\g����f�q�)�X!Ɏ-�x����<B���{�.����>���q��z��A��1ș�zj�Ќb�G>%{C�}��c�E�b+� `�L&�4YfP;q��B_�g+�O�@�$`"%)*���N�ا�Q���`�t�/w�H,I�> ��k���<�A���@�V�{�� ?���m�7��b��`��7��q=:a�8��
�=�Tu�H]@~6tWIB�6��`�-	�W������q�!њ�-^���q��>����_v�ǭ�vj�pI�6R?��A3D����9QMK�����&D����d���p}U�	[���O����0A��J����}������Ak߽��1h��""F�v�~W�1}�\U&gq�ڲ_��5��4i]����h��_z1��Ը�4�n��D@cJl+���byߋ6b!l y�=�ΝIk�+��}+�w��Cj8֯\|B:k���+yܛ�����R#�<��*NXJ��Џ�`�A-(K�g�'j��k����.�.����v���}������\��1��㒄Ϳ���b��g����>)����k_��*F�/[v�J��)��+8n��{���C.�8���X�;���gQpB�ja>K( :��wH"%�v���Q;K��\�>C�i��&vk	��v�쩜��"sL�-�M����c�V#��A��Ƶ���պ+�O��7)n�y0���y��h">���m��|��_�������F�tn�k����%Txr���HS��	��5R�0u������X@�*�5|�EZ�dBߛ���#9Y��SF o��Np��ѬJ#�d�y� b�}�l'�b(Q)z�0�g����& �pP��7��j�B���0Dm_sw{)<,�=�*=�m8S4^��Z[��Sƴ�K��ߒdu=F�s���*𡱴���M�#�2������u���?��t��lbZ�@ɒEʨ��kKta����?��d�\<��V\*��Ǒ4�杌;�Y�ʉ��SB����g�J}��;g����ʥ"먰3�?�{0ޡ��G�����ܝl+�)Q�wY\�j��[֬ʹP��f�a�L7ڥ8�M�6 ����V��ʎ�>����I�"@������̔z��̶t0,y�-b�LY]��hEy3-����_x�sj�2�k���|m7`
T�תV�@��[~�ܺk��`u�y����A�/��`S��C{t�g���Ì>0�r��
Hل�H>��rO��>��T���Qb- �@��J'3�&g�:�����c��K"j+�^��άi�V�����f�܌>�-�]P�ᖵ�=sS�_Lo
��s�X��'M
0Bh̃�1���k;fϫ�������=���� &`��B5��(��L�~,�ϗ͘�L]AD�����P��H�g�'�m�N��2���==��m�'��ň^���RA% �l��gxp֔1���8�-�rp����Ĳ[ƃ3Zj�QJt��}�B���*O	nj=-(�@H�{�p->�Ԣ#j�l]D{��iz U�GSԦ�A�z��VU!���>Cd�ɵS�乱4���G&�5�c��6|��Ui�ur�4F����r���%B-�T���b�/�'�?"0������;���|,9I�_���o����a�0���b��	9�E��+p��>K��rx����Ǌ�R%�Ə���Rasz�������Sz��P�^XYE3�S׫�$��p�ι��$��n�J����[{��hTe�e 'Ϳ� ���g��E+�3ȱKA%#r���)�b��8�s@3��g+�5鑸d�u'��oXà?:���!Q݄�$9�e�1� ͵q�t_����F����C�llt��S�n2ۄP䈐�ܒ�(m� �[��!�X(<B���ȥWT5��>�o���8cK��;x��j���+X�������YiT�*�P �B��wp�<ʶ�X31h#M�X�H&��X^,�c���t|}VSoн�  ����P}��W��y9���`��FI����]��3���$�J���$H��g����l���U҅��:��֬���j�����50�͟F �]��&���{���f��0�\0����mK�E�b�}y�h&��AzqB'�$1@ �������F��D�e�3"�h��
�9(����*�Ix?@�t����c�4�i�!���Q��d�?T�+�gcFw���t���ɓ�8��>��&��Aɲ��ǍNץ�3J �J1���gb���� iD�2�4��L��*���Q���a�n�8u�װ��gMi��q��а"�3%pa�<�DV�睆��	FNdb�a�9�Z���z�r]uR՟~�4�/���!B� ����#!�2e����0�������b�i���6� ���;�T�#�PG�p&rh�E5ۑ�`��‫�	����EJ�^���`�l�崧vʃ������:o��}]�O�~��?�?�Z���CJ�
���W���&o�V�
�S�}y����e��D!����Gk�H���S��J�<˥��Չ�ׇ��9r�i�T4�|���J��%��xMH&�]�g�L,�;��.��ΝU[8�xQ�6�������XG�z83��F��x5~؛�2�JW�����{	#Y_H^��qޙD�L��!��X��jțe���Aųo
QF�ǖ��(8����s?�_$��6Yó�ϐ��^�r�G�d�5�	Z�M�z�n���*�c��,u�� [��xR�ف���}m����KX�&2[� �t=?�Qn&�K�6�Ǿk����;�l�1�0��L ��s��I_�.'�){�B�w���L������˦8w�{�܈]q�3���oF�C��1��ۏޔÈ�}�����ԕh���]r�V�/�BM� �Jm#��SR�,j����:4�ۯG�?��� �0�h�^�FX��_���Fv��|�����J9�w�lB��N�c�	��V;�Z%�u�3Xr��g\1��í��Ҟ��?Sz�hǦ:�̛:��) y�e��Ϝ���#e̿l�R2f�֕@��Q�c+��.U�)�2OW�� 9� ?���Q����y��T,�Xw��l��f0���נ��0A"�@�/{݂���\��;���Ĳ$���2^�=ة���� ����tP`����4����ŋ�
�2������v+@��F�O%����9fc�rW���Z/���ݚ����`C��q�oQD�E0��d��Y|��z>��D�j��oy��ގ[� =(����kr�~�~�,�*��'��ry^4'T�����t���\|4�;u�5j����	��bhG��YfZC��[�:�lm쥀F�J�Uܛ˒/��絥�F�	6#��Ε����LOS��-=e��0!���e fH�M��<4�ͬ�Plþ�N0��ؘ�N����4���1�aƲ�5-K��pιQ���Ę|�@��K���k
���@�����k߶�?.��(���	���B������f�͖$|�d"d�_�3V� ص��u�#��t0	�E�\嶦��%����M�!��{rL�ǁt�)}9{�Eӷ+� a��sφ۵��,��W]��09?K�#��o�l�5��죧���q����K�����ı���Ӡ�W�-�`T��șe�<�DK�?�̝��1�u�53�z�u��T�b�>S�|*�(@�%U�p�l*�Z������̆�1�����J ���-.u���"�K�2`�� �yd%~�kW6��H�K��Y4� x�����m��դtV���I6�SJ����r̃e?�D���=ЇJ���[aQ�I=��`d��B��ct� ~jr�5օs9�����B��F�ڥ@@>G���0�10����O�J����=����K⍲����m�)���a�x�Σଖ�1������{r�lW����e-��ʦzd)1j[�<e�����&�H4�o`t3��r;?�`" ٰ��1s6��&�O+�ޓ�)�l��>����3�u��uk��8h�\E���&�i�(��	�hWC78��A��	C��om�L� =��� �"�A�8���y��� �o�n��^e��>�,�L[���������Q�ȟ@FV�L�~)L��2�䉟D\hH�2��t$��E�)p��:�I@���r	�:�A԰!	�"��ۗ��$��c���>pR��
i]�*#A����q��/�0{Ѭ��fqL�*-�,�y�m�oc{���s$k^�7Q�G-��[?�ӱFW�0.�"IcH��cKKo�FR���������Rڕ��$D�䆋��V��4�ʔg�iJF������!�@n����~v5b���0��L;���}g�+��Ң����͑��w3�g�9>�p�� �<�~���I����<Y���Hۥ�Eٮ��ۼ�P����q_�-��p�e���;��훊4Ÿ���"��R�"pk��ΠhX���D�u�f�Xa�wT ,;:�&���
�/P��f�!D]�!�&ғ���dCS��6r�@ʫ����-n`?ܖ��]�����r<W�x��Y��L�ݤ=� c[����mQ��}豌9�����	'��uV�Zw���)B�*+'��F�6V����Ok<������J�����j�TQ����WlUN��4�� Ym�Ȩ���HS�\�%��[e�ǂ�D*IEp�}=za�G#fry�6�҄U�v��)1���*�9oIGk�"�O�"�>=��؛'.3��6��o�j\V ���C����0F$�>�N'8���q��H��Ps?f�`��W�d)BO�6`�WU3��Or������$)��9s-����k�Cb6>�^׎���>CW����{���ǚ�������Bu�����-ݶ;��;i���/��x
�{�ɝ0����c�M=�S~߈l��x�B���3(�C�9�YD����|F�j�-|P|�l3Ic��Ook�V�tR�y���0Ӷk����@��� ��]
��~�Y�;�ʯ�B�2V�I�v����Ƙ�7�@�{�4�un�1k��|�D[/Nny�Ʋ�(�����ē>�|�1ʚ�O��=<Y�%�0WD!�qq��2��ǣ˿��~lC�v�o'�㬂>\��{ 	L %9�b��R�^����~��vp.�uHa2G<���n��"pw����r\�� Ii��_o�ɓ��m�;oYU�1GIL�����m�m�twr��������lt��:#���EL���x�N��_��e�>k7�i@.Q3���IG;������T6�eKG�кi�T}R�"����ݬ�:��|�Og ��/v����4��!�Eç��K��kk��!�b��k熽��~U���~)�fU�'+¦�zڥ�T���/!����^N4I��o��|p�h������g�ϫ7�`QY���f�1���3��ݷ�����F��*�ʁPz����N�7�m}��`֝H��a^\��[m��H�r��ɴ�j;9|�*�O/oB�N7v��Q?R�X�����Y�c-�k��՛w��q�Uvw��tfe��Z��N��8g�s:f����v�$�9~X�L����-)�?{� �����H�-RH|D�L͕�4j������p%	�{M^>8�'���7E�(�02�.�&�b)E���Ш8N{X���ֽ�O��\�jX'�L� ^����B�+	�H�]
F��$���K����늜s8B������s��q��Q��L��ݟ�(�A#zM&-:�A9%��7�����v�*[m�{^4d��>�$�j����[�K�~�J�xrit.�"S�8����&�n0�����`!�
�`�}��kh�}����r3�]:�8 ��x��1��!�|5�:K?Ã��}4�W�ߙ��Mv��I��w�Q�M
�ӭ�����I��oѼ�'oV7X�)ٙɸߞ'���.�ӛ�z�0@%w�엝�p:�W��u!W+���0������ڡ�XH���I�� E[�^�z�u���ܒW�@Ü3��y������� ��qc�ށI�u�]0Vz�O�o���e_l�7�q��k�Ss젤6~}߻�/Br��� ^��-x��	x�~A˸t1;�*+5�0$��dG��޼>c��Ҥ�tǤ�l�z��p����'d�R������i��[��\��Y�ZM��+��`��R%+Kο�;"I�����^��J���T�}�L3��S�9,9S�`������||�s5G�P຃vsH@�0&uG���9�y�<�[���'ҳ���Q�M���vRZm�ԛ��Q�%�J��<��A���<�M���{WF�\�ӂ��	���Vj�""�sW�fa��?����_w���h����|�E�1k�?���ݥ��Rc9�8JUL��z�3L8�|����l\RG�6y����E@@v�v|��)u�8�? ����}�K!yf��S;R%��<e4��bt_vRI�x�x���h$�}�q�J̱�Լ�C�6GJ� Ym�I��Bꁏ��=�\�Ӏc���!-^w�#t�NE���?��ï�?Z�m�xE��"��z�fNx
!��7k�+l���A���M,��I9�+ț�|	ۇ�`��x �٫}�����0���;9����ǐ���Px�\W�^�L�\�DZ�)�^�' Հ�U)=����K�`��	���:�����������^����BY��x�4��I[wdئc�:�[��9�YL"E�����	f�n���o:����!��o��DpD�ɟ���
~���9ױy%������^7�0MS�+��)��E��
�l\�*�Ϊ����lbTҴo��G��gC)�%-g��gϻo�I��P��� ��#�k�_�9�kO���Ɋ����_7T%%�0j��%5��Bٙ!Z_��g���I4�x�r�N���m��Tމό�G���-�ѯ�"��;�ª�t+[`�]Gg��y�0x�65Ѓ��U�+�d�(����1X�2�=ԍ�،�x�����~��X'�����n�߶���I�Q�_>��+q�ֱ��h�`X0�WW�/n�xR��
L\��q l�����NW_ح�^@�w�%5^��"ٶ����{4/��C��D�&��nGu���ݗ�B�O;5+ht��L^���p���iem�׏��E/�S�jM�����$��x<-��_��0 �z�����}&;d�	�0�,
�]T��e�����VFv��,EY�����J��-�h��n?^�����^�*���w䐔Qk��sL�u�Ҹ�Ξ���r�*+�"����i�p�Y�9��gugjh�(u'eŮU�a�X_-_hyK���a�aEz������?Z�q-@a"i�E�$J{��D�P�1��#W@U
���i�E+�����'F!nK�8ƕ�d���eH6w�S�z������,U�X��!ݾ��`u�7'KH��� ��	�qK#|o�Rpl ,��}���l�Gu#�]���8��.��o�7������p�H'6�6Y��<���;&�u�kG���R]Be1�`sxuP	�6����+�y�]�d�pY�hY��1a����� t]Lw
�T뱏�OUӹ��)��`Z0��s�͂D#p����kE1�����d����0��p�
�4�3"�A���Bx��e�V1��TG�	ɘ�٥�$�&w���DL��Q��`V^�s-�
�CA$�����N��p�@;8m��}C�@V���G=���Y�'����䠯��Ǹ�:� �T���xA(txx�y��;��Y�f�[��U�G�r��y��;�a�z����C�a'pu�K�h�%Z'[���G`�{���F�_�[9�h9��{�\�BK�Rܪhf62^{a��)�Nd˲y5<���6P���i,�r��Ԛ(]=��wl$ v�~�k��~.'t#n>i� {�6��r��H)���RS��m�����_�u	�N�I |?�� xJ���x�J��V��Wv?�N�	��jި�����,�ZγQJ�R�Q*'���Kq��5�f������í�2
�{*nń�f��W�r�3(�l�$֝t����g��:b��<��[W�����26m����o�@x7�Da�Bw��r��1/ �v~)����[��Uao�s�Fڶ4G�'�xa�.4`3��8.ۣL&�� �,!+V>^c��μ�h��R�$9�)
\���	���w+ �@h`�^;;�߾Y�36��ߧ��F1�'?޿��cm��*��.�n��zj��< S���>� JdztE*�]m��no�0�'��Mh�+��d���+ 7,7���#�`��	��[�V�+��eB	NDu�(!�k&�)t�x���N��([S? z�ƌ�h"���X8�!{���0Gn)���R�_�7|�5�BE��Ԏv'|�=o�AW��2����P�E�%��b��P0�-GW���-�P�
�H�ۢ��6#O�T.>���*-���b�Z_�7������cw+h���T2���=�-E���*҇�GW�(!�:�j���E�8P���B����������<�u�{KQ�dj�L"��m1��I�ʹ 8s�2�/��P[�*K�N��l9QV�����O��?��	���P������̊���~�B��bNQ.:�z|d���+mhK�W��������d��-yI�����mhe�YG$�Q_ː?	�N&�e����	���_��mI�/���k=p!f}`/"f^5k�Xf�=���F{Q����yN��uC�ѫ��M�>�m��i��]~D��⦉����лC�S
����_dm��ѭ��{������@��pX\�:d��!����2X���R*@���^����To#5`ț�<Ӻ`��̅C���˱p�ސ�f���b}����Ew4�w���P��$���K��^}H)fx�ɧ���'�/��ʹ,H�[�~�����H�bp��V�cQצ/�Ƙ�O�����@1vw�ߑv�� �d���1��!c��8/�N�\ۜb���%6��XbXG��V�JB.�X�c{�A8����A��ӭ��{���� �\.��T�#@�R�D��f�9�ut:U���};.�`�o'�}����&���B�X�T�/��zھ,d�6f��\��l��L��b�Z�X��*Ȉ�$��)�&]��R3��]y�_M�X�=z��3
���>1�Z^�Z��s��:�&�è?�7}��:����G��Ώ�f|��$!�5~��k� ���&�P�Ĺ��y���,Ňx����U��	�G��L_���gD���c��'̘ߣ�f���C1ϵ��w��I�W{�{�ϊ=,�?��߀�Csn$A�ފ�4��ߕoE�=S�u0�ƿ�*ӯ1G�k�~^�~�tB�#I�����
���]H�F�|Fr��2��"�����	�?i�T��1z[�A�C	}�z���B�k�0��c�3��G�5�s�|9uN!�W�~�5��]�R��ݱ�ئ��8��Ǡ��/?� w]Ia��O��\�$�umml������.��9#���s�#�U��>�O�6��UL̾gV�}��g������Y�u��������\*����+s��E���xA~㫹����(qL�@��j���=�t�m�t�����/��|��[EM|Ț���>XǄ������QkJ(�0+A���T��
�s�
�I��ԡg �7kw��2����1���-ْG�Ӊ��aFE��}_����N�P��3\H��Q�P	�\h��h��<�̍�2��' ���4�C�U,=:,�2��$7�"�{U��8j��\/�s�
G��"{�~M@�h�,y��+�&b�Z?�q#���a���YZ~P�wś"2��E�<F������w�K�݁�f��M�����RX�d�j]9�.���/�䅺Hz�ÇȚ�d9���[qEe���on瀗�$Ig������Mogਚ�U8%�����ƫ2	8������/]�;�B��B#��r��-H���3pp�ߔ�'1�L_�1Z I�r�c��N'ܣ�ٝH#&w=���3��xX��S�+�4�}/ԙU���#wږ��R����������K����+8yS�v#H�����bH3��Ds�F�{N~��yַ��Xh|b�CVN������.�[T	��œ��E`�GaT�F͔���{�^Z��_8=�-�p��Κ)�ro���?��C��T'O �e���3jmq����9�sΏBٹ���T8��oS��X��:(��f�s������wn¢��,����-x��=�ޫ.��s}��a���ej��\n�bo��S���	�����ې��|Z�yk�:�YR툇��C��r@�,�E�F>{��@�FS��HKi+�)���.� ]�w0�ċ{r�e��E5O+�s[:iN��.t`Y���^y���G���%U��!X�}yz��7Ω]C�м����J½�o5w8�|������ |Fj��"Q���QgfxG�x��d����3�w�/�����3��oɾ2�V[�8!WȹG����rme[,3hfʀ��n[O�}j��Q�B���;��yg�[�
Bk�vL��-ER�;�wsC�_��-���A�+a�C�d,���Ǳ���
	@P>�����e>a/�����ST�Q��
s�8�x�"��������������ٔ�Ӥ��J�%�;�ꌀ����a���co�4���C^R�kNK#�h�����o�3�(���N�����#}G�̻�pgG���0�Y�[JǈQ+���c �:[3���� Z�*{�E�7=��j8����(��?GR"6�҂� �VL`K�j�+o�T��o&��vs�Zn�`����|��*�xS܁e�K-4�[��Yӫ�? ڲu��I��xO�7H<E�>������Xf��`�}��/|��׍�O�Ҳ���t<YG�w��	&��h����
�5ݹB��`�:;-
JJ,���;�8}�@���V;b����q10��8)��څ���߬�G�PDID=��(����Z|NR}�� �IE�������w��(��i����SZ���9=bDIAhn�'2P�g3[LO 
�#S�
�_m�ԋݎFcr�y�Tn�3����N?�R�Kz�������-F�\<O��r�Zy�*�qJ����8�=�.f�����b�s=f����F\:�Kb�v��ȅ.�N2�ܡ�x�:t����W�{��9�u�����'��7T�|-x��b 
pL����+� ��������AY�;�t!cq��.�@��M <�Ң��Љ�#�i6.�H*�á�Bq���|4')+qO���Z)1~�2�W�[R �W�\�y��F^����Lt.��J[����h�j�IM�D������0W�����e���j�Yj�5��bP"R�ߚ�'wwI[nq<1vgz��t��D��(v���K�){Jq���FH#�b#�IѢ-���3�$�� E4�k�aǴ8��Fi��mfi�>�,j�`C���a1���)���	�(�G��H�3����Ԁ�T� ~.��'QG����sqQo}{���g�dp�����~K\�>�]�eR�<~
��)͹�K��W �g��͆�}�s��|�aF��<!l��~y��5��Tm+�]<���E�o�Β�m6�`5�E�HZ j؄�V�`�(Y�,K����۝��h�"w��c�d���"���ي�H~f3v���z�-�v�R�1R��/�SW����S�9�����m/��'�E	�[|��/�$��\�l$6D�_�h��aIVc�ޥ?� ��R�W���+S��!���KY��<ĕ�S�s�n�K��n"�S$�d��\������"'<-���q�e�Y��>���L�����-�/��e�8���d�_��;�d4."��|�A��5�[[�WH���9(@�5���s���
\n�����c{x5 �lN\ې%(�� ��o���\�j."z����0�%�+dR�(k�(h!<�L��n �݇S֖%�$.�}�:��^��7��W&I�_&4 ���K� �ȁN7����W�Ee$�ȭ���m��a`�����Zb����s*��i�6���+�� ,��.�ɲ�`�.�
g�( B�hc�q��5D"Ϟ���E���ר�=WO���(����O^�lx��6���3sd����G�;�ރ�:�D�(K���Rq����E�<�A@_�ky��*�4d����LД��s�a�UF��1��xH�.��9��Aq����n��_���u^1���;��ZY�����v����ZAa�1��4|�����?�Bo��Vn�����s�K��޽�zZ�m�̶`��C@��&���~������N����"��*\K~�FQ@�>j�����7��c�;t�����(S�v�zKR�@� +Q�"�CDH�1����?�h�e�$�AX���,C�,��1�j`ˍ�&��%�A�*���p@}�<�����U��WR�Ӏ�">�����/�ib�#j��oq��y�?˸��O`����?h�8�7`gP3Õ��j���<@��A��Wƺ���?o��
�D?2��S�9lK�`�����C�o�\����"e�g�k��M��
;�K��Q��pT���Zp�(jCL!�Cd'2��ܧ���R���o� _�zA��Ǭ�-���8�(��r��8���Т��nz�͙��g>x�V�/�@jm_�@/]�L�&��2�Ǆ�vN ?E���7E�����6�o�3(�|�:\��݅`�b"�'�r�@M��ϺY���+0����mF+e=�F(��:�U���Y1?1��)��h^��r�S}j#`��v�V�_���+�/���6k�JE�������T�)�����(������I�*�:�y�:�o��B���qΣ	��<�ٲN�LFJy5��O"�/,�-C}0�n�iԙ	�Ł�Ď�bTռ��S�}��f��w�!R�y���*-���nk��6�P���R��"՘m�.E�9 0(Bu�E�'U�k��=*+g�����É�z�G���Cğ6*h�	�������cJe5�\�c�㗅���Py���(//�J��K�G���i��?շ�e����(�q�~�������$1�9�!�-��n��؍�!
}>p�f*��Kثo���/����;
	�>�M8��C9�����A - F��*�`r�����V^�4cG�8IƖg�ܔF;�F[X��ʻz�^����Q�ݐ�*��}�]9�X9鍝`�,���s���Z\GF��(�y�pv�;�˰_�R���1��薔H�O�jR�@k�Ҙ{y��!�� �8U�H�B�
�	��V�����9u�ݜ%z%���S�͓�1���i�d;�:�!~�}}��A�((�E�Q����'`�=����A�q�㞁\'�b(oοlxp[��}{㦙L�k��c/�Ŗ�:I�Rg����񱺶{��W4�uG��W	N���@�Ű)� �]}�^�cDOw��٘�±�p(�g�/��d��Ci-����0����c�<���mt�� 4�t����E'$�ׂ��� a�ɜ�Q�Y���bv&���ly���� �4�Y��'���	��ຽ��{G[Л?ï"%Zj���zx�a�
�G�a�3�	e�����$��� �v� U��k�)��w��ѷ0%�10y�d�%i8�*�t� U=�2n��B97���:��}��PJ����~�e��<�a�%;�.z#u�����+A�K�@l>5��Hą,#��}Q�:g�qƸ�!���&�C3��>�Ԓ�ざ,���V��,��~�f��W��~}�P��K�����_���{��`i��[�������fzmڦ�K}���ݺ�s�U��?]��9��G#(ˁG���	pv�;��#�"E�k�z���rꖆP��nr�?��ݤ>�����Y��O�u-i����v����j���u�T���]ܽ]��v>RŖ��foR�p��Ij�����+�Tow��5��`K�}�G�²�������\O$��Yޟ8�����a��a��=�}�T �<��������e�q?�����nhʅ�p������'��"& � �e���^�Qb�I^`=Ţ9����>�BR�H/I��1����jc��,rI�KH�巗j�p����鴔��V������4�k�,������à���l�5�e�s����wx�op��]����VK_%�>ֆ|�T�3��sr���x9������z����"��B�g��Y�<����#����gٵX��V����vl��v_pQ���A\ݞfL�M�����u��"�Ж̩̺�~џ�y�4����F
��^�|�LU��w0T�<L�6�f�~Y��E�'��L����gZ��"��7�A�t� �%)7[�/�I;薟�4!��u9��2w�i�P�cG��ָ!�%	-K�P;/�uöm�¸Bc�����CN�n��WFn	���=͎2�
���h/Y�;LD ��[�RI��;>(o5w�k��@g2�钷i@b��}�ӯ�?�S��8�������h��W���w_BEZ-�]	ݬD��t�o��!��5�M��-,Z�z���fꞝ]a��{i��+��|�i3�ԃ����w�qC+���FY� �7\h��8kLBrbjN_��Q4���5�Z3������ܞ�oI<�2VYWbV+�o8z��|�hK��D�+i�0[�8b�ފ~H�z�D��	�����x�x�gt]�5I+tAgBf�q�10�;\rE�1��
)kzl��^4�r��1a5���
�9s��xi���n�i6��WrR��6'��=ޮ��l\�����c�΀,Q�K	�Z�h�	�j�޼@g�)�'�o���ܽ�6<H:I=�+��qi����0�|����̉8Y���#-�x�~oh�Q(Y&����g���>����S��I5�E�hk��lh]s�[��C���k�hp<�V�Wꜱ��C�l��]�LaU'0�|��Z���t��w�ђ.�hØ�������E5�c��y���Xl��T�crL�c߲���+j:t���=�zwOGb��,�8�p���^��˕��Ni�u|�ޯ�z�K/�}�o�N;��{w���X��l9�K� �}�3`]8��
ܾܹ�,��Ir2ё��+�3P�"[�C���P��ZC�+��q�dz�m5
]b8�D�g�p}�[؟�J�]�pw�����U�	�%�~�'G%�h���L�S#H'0AEi�b�l:j��.87R�ǘOFA��]e��V�Ӭ�Q-�"��;(~�����>�����F��uT�=*Q�yȃ�h�[�`�ي��P}UO�t� W��me	nܣ��*E�MzVSi}���X�����<^W.��0s��|K����Z�T��b)�m4��M��*>�s{�od(� I���	��"��܋aH��<�9�v���j:�<��#�~l5Á+�o�[��ؐ��ˮ�`���z�rq$��3�27{�	�}ծYV�r8~��]D�uv~�#��f��9�B�2�C��$8���yBl��W�T� l���ѱ݃!Us���X�e�ϑ���?���0�fb�|� 
}����Q,�E	��w����?���B�D�A�a�C!R4yV}5Bٶ�|1�|���l�����*�;�_���P�W?���F�]���pUh�LĴjB�`����	t���P�����r��y���T��P��S;#�ԙ�#�muqϑ:Zd�N���Y��w^�cӾ���|�l�-{Rؼ���c��]1Aq@��Jgn��p�U�ek}ث��?f��e�,�3pt�ø���ݑ �r�z�:Su+��yŋ���*����b<�V0I��;ґS,�$��dt�����l�غ-��lӬ��麉a{��\�G9�]~bv
|K꬚A�B�H��2���]�U�� �'�(���@�}�����sL|I��=cG��?��)��h>���@Э�	�T~sqTbZc8ݾ��sz��D�JE�iKos�-���[���C����	p٠��-Z�����u��)�� 02��O�� Ѫ�Q�l�z3�=. ҿ����6>ه��K{%��]�3�7�$�$�pq����ZB�8{�
���~&�@-]U�pC���]}^(�G�c�݅�<[������I��G�q�_�-�3yT�9��	�'�Q�9�(8�'�j��2:|���q����6�ͮ�%�ДL2x���`}2S�x&,֎&W��.)��3�/���ׯ���!<T�CТB�<����=���U����o�(ʉ������*C�?E�hq���O���?�\$T�*Ȍʇ�3g�'�"�o��^��9l�H�=���3P�S��@���J*����^B�?[�?|��7���?���I�����r�R~��p	���9Z�(��WuӮ ��g��t��������%p�����pe�����`�[T^ �=?�� "��:�by @̌f��U?�T��֑C��V�2�4��K�vr�f��C�r&i���t��;��V�#�4U�!7g~�R?����b��P��d�7������U�q�����z�&7͸[���@�N��r�0p�9�B�h�b6�S��h|׫@��.��x��ׄ7)B��C��������=x˰�"ڑ=m��tV�~i���Z<��q�iG=������xY�t~�����*��7SϜf����75�=v��8y;l���W�Z ����η~��j| �Ax��9?m4$;+g�YU¶J��Qn��
FE�U7Tz�`N����Ԍ1{{���Ơ�%9��<s"<�W���O�A5c����|5�̈́�%��b���/�Z�6�'�/+H��a`U��fKz�Yr��%-��HZ�T�4��CG���c�/�g���g7���z&�ZX
�f�+]r��Lom�mM����r�[��%u��VUɆ�d������������(�К/>�-���B���:�n�5~��S}�� �;5�����O!_��?!p�o��^������F�S	��AS���,��@��>�F�l��I�lB���)����a?	)�P�*�s�x�X�>�y�i�B��L�ǚ��Mk]/SHZ�-��E,������3��E�/ ��w���:8#\Ć�/��t)�֒�I�i�~���s���;�T�$�3� �fH�F��#Ã.��j�18ڟ|������wl�	��xZ[��F��/����b�mi�p��+�P��f69��i�a�H��n��l����	�iЖ�M��H����K���3��U[C���rug��?j�C��ka�v`�z��yh\�TLQ���h�5�z���K(���K$`�`�'%�j��X�b�k��ҹ�l�}Ab�n��'���{��E���b����8���5��{��D�&Bɱ��i��f��p��I��2�d����g2k����6�y!�:��a@���*9(��?r%2�[��*��L�?)����1�{�j��Ʌ����h�'�7�u����"��4�R�sJ#^�ހ��5P�Ce�	Y�rC��+�uv���ѓ��ܩ�S ���
������A�m_G%H6a��@��H�a�+�X�\#�_��G�*(\1J���1k��6L=\|�Ŷ����Ws����ƒ7	��;�5�G=�ɀ��}�����D:�����i8��B�ma|X��w�:/Z2����� ;k�)nk��.�ק�>�Qa]3�
���r-a��x��
#�\N8;�ʹ_=�ݛ���M���d��U2[��zEz����9i#/����N!C�B����.5�}Ǿ۰�!��	_O��>���Z�L��֖F^ҸхZ9`7�k�r�^1�L#}�t�C,�T�w�X+��>����@7��D���Oyՙǻ8�R'�m�t�S���=+�K�{"�%$id<���j�f0)d\8��S�q����;�1E�rv�}�bG�E�m���'��/������ew�0�w̦�*��,#�Yr��ۜ
��I��q,�Ro���ę�^��du�2C�����-戨���mxp5:}��5щ�'(|�
�;���F|��_�u���6�Mh7U���|r5���x1Y�!v,��m3����!9��1Wc�l����f�0.��#ˡ�"�ZSP��&0��7-`�ƶ�}�J�O�öxq�� ����Ii��n�X�Ny%G��y�_��f ��=���F?K���m�Z��/�V��'��wQ8M������6���Vu�n����pF���Kx�Fu>|�������G�R���ߵ�dS "op��fOL�ڰ��/Ŏ:W��v�%n�7���L��J
�n��lW��sQ��N�PEP�M�lȴ�5��nu�Z꿯{���Ǚ�5	g�g�d���[�G_�v�l�Y�੨*�ZmTdIO�b�_�lk�JQ>�J^�X%SP��W1h���6����~R�e���@ �4��̝.	��k�D�cŻ�U���ƱGr[Eܑ��ly\����PѲ��r=�2z�=)��ϲ�%�@�_�e ��Z��o�jb99-�����Iǆ�#a짮3X��]��V��Q8 í�����(�������A����.�\�S��|�)��i?�H"m}1*L#9��ir�fe!q�r�b�?�2��5\b�0~�׵�\�v�_��ͤ���>m�%�ۿ�^�� �i5�Z�Vْͷ�T��0�tE"�t�7'�q�'e/���/��U����։��D�G(G�� �X����q�.��M�]��!�z8����2zڢ|IEIi|���� j�[�^�z,�E/�eH/�>\"�3F���w�����=ի��L�Yp�hL�C;uuz5�e]�#Pږ�zG��:�'� Vv��Xkͩ����MΡ���.��Ț��t�?��/���������	���_U��"�6f���O�l~9t������?�!ޡ)*~J=f�M���a �G��HMչ���2�����B�����D�y�}��t�F��S�����S��~��j��9; ���*���&��0Kj�������k�"��
_M�:�����ћk태iX;�S�e�I�Ƥ���Z�F�:�C�2�S!����m��p�r���>�D�5G(ƍ`�f ��M�����A+� c�ٽ��V e��il����$���M��<���݋�ب�M�o�IJ���?�Kd�7�a�\㓰f̥׶�V�a��g�ɪ��Qix��Ȓ�`kŚy{��FUEe:a�S5��lغA�]e�W���Z��K%�T�a�q�i �*��3Ͻ�b��8\W������J��^��Ɨ3��̂iC�|6b!�G��d;�\����h����|�� 巘�YAXb�>=��%� �q�9S��w��i�����ֱ��K�+��.����Kx!�tޛ�G�b��V%�F�hZm��W�[��~�H2��4u�=�8��P95�"��p^�>�To?J\ ��v�(}� ��π�uQ�x`gQ�n#��leﳘS�Õ!��ĵ�)ni*4_o`v��1e/f�(�j��5/��"n�4�]^_
�.��w�G8�b�{�R�2:�����l��	#�K�>��}�W5�t����
����t:5������Cm�2���d�#�¥����׏*��m���}4����{���zf�O|���P��	�]H�:�C�@�jԯO'�eS�Ժ��*4�:�3�m��>�b٬�G��+L��J�UC����_�t�0�b�B��y���� $H3�C��S �q9�}�Hݧj_kP������ȹ��\������:�������E��T�����C�c���M=�v�?PH� h�Q�>tF�9Bh-��G�k>E��'y�B�wu�ܕy�2$]fԧ�&#Zak�T7xYhGv�.��mxkg{/�g�;����@��P-Bw	��_t6����3��!�}���{IB](SO ���Y~X������5R�1z�vBBnT�}n|b�3�af���{�}����9��P5��z�ʩ_ũ�x(޸XJ!�.�tFYUai$�q`�6�AN�sWzl�P�N�<M�k��y��-/X������0����E���"��#����N�V?���&u�#�q�7gz)V�w����[_���$����ǈe1��G*���^�ϣ�88��tF����SP�4)���B��m{���ba�h�׍x��@#�"lh��ϭ�+E�z�sM�����U�n�>��V?��U����rb��R4��[�k��f�zK�3���e��Y
kȝ�z,	I;�^$FIT	��*� >N��W�!�--vB����p�#/f�t��Nw�g����t����9�"߼�4V�o^�Q�8���l����9}� h�`/%�{ɡ��7j��A�@ͱUQ�[+<1�ߝ�jnƽJ�\�\�Bb/��Sk�hJY���"���ۇ����� ë)<�;�=�$����Ǐ�G��\c���M��� ��I�v��d<�^�đ #:hѕ������.B�GT�h�ݩ�YY�]U�gJ�Y0��+�e|�y��8V&tj�3�ܨ�w3��/�c��M�|B��џf�p��a���^7���7S�*�eƂ��/��h,œ�F�O���j�
v���,��vBG����H���8�(���%K��#C<�/���5�vɳ�Ū�ZJi7���X�hG�B�,z~��
��o���Ɍ��3/�"jt���8�8���}W:=��a�7��!�:�v݇��ٺ6�Q�<�{�T}F �b/��Td��)�M�.��K��MR�o�_GK���UϴDC�{�-����	�Z,�K��(sTE)ky}9��Ƹ/cB�͕� ���*����Z~���Jg!�H5eg��K��ݹ��p��:���xV���R̢*�v˅S���X
�?Y��(����B 8�l�]y?�HNK����`��(��?�V�>��{�\'M�?e'�#b6#8��0��F,�����jp�<����/U׌y��������'�X���!�a����%��{z�$<�(K�Q�׼�?n�Ji�Y�t6gS�{��[�F��6�cm����
Ff�`v	�xKP2�M?� �(��ih�X�̂#ʽr�� S\�C�́��u�;���3�u�� �X$�8|�&��'����?�#��U��58����� ��ۋ�K�.�t���*���H�/�5b��sB+�`H�q1C^:��jԴ :\1=8s���:�}�3��6�� ԓ�/�ՈF��_Ӻk�ղ]����sJ�w��<1ft�f l�Z�^�P�Iv݌������������h����c��V�簕����	,6C�az7���S�OMC����vGu�+9��i�WvU]�3�b�/"7��|0�6�eu�<j�y��rE!�!�7~p�s����~&��^�2��DW� �׃r�t�9�/V{����4DzͲ?�gbI��z���DA 3��rM�ր[f��y"N�z6s�!V��/I5#R�.��z�
�\̩E�\,�������dQ�"C�t���]x��4�ָ�P�Դ83��ϋ�^ sy|I��:����8~k
 ���<�N:�XG�������kR��_�z�����'
)�h^ԿL��c��@����X�&L��1��{�u�jq�}�-a��PF�RM�*�|�>
���"���U�D�}1?z��@���ߩ�l��L���2� �E��G�1aߨ&J�us�A�b~8w��8�|	��x]4Q�&X ]��<����/�ɶ/!���]� )���w%^����с��� �sgF~�t��
��feش��w���	����3���;��,����	cr�|5 �A�|����`F���Te�`���a2��}���R�3.�-RK����H35HsL�#���6f(pی�t��#�B��f��XuW���_�'-�ڭ.�cU �>���?7���s���n"b�;�����Z��~�#���>(,oj�+!f\&�	z�)�| �o�G|���ע�2��0���0�De㒹E��xFz����Me9;���o�H�gH�,M��]7�3�t �*�^��*���㢬���FT��J=Q�s��ȟD�����"������zK�?������3������j`� ���?!GF����`� (�{���؜�(צ:���4�pH�]@�%�2��H��ݕt���g�C��:P	�8g7obrbdmi�52��_ K3YU��缀7�#'mT���Sbt�@!�Sׄ&RЯ��_�̻�\���3-S�g�_z�@o�~���D����3�����G����	�I|6�z�T&����+'�S2=g>��*8uAoX$��ҟ}R{C��8o�W(/�G����l��E�w��N�l�o�1<ɔn�?S����U;s&�j��B,��Q��¨��1	�^'e]�����Z¡����(4�+�s��2����0���G����%j��Ð1)g��z�N ����_���e��r���[֪$20qtvM9@��偺U$�2��Ai ��#ԴH+Ѧ��ܙ]��iU��<�q�|������f��Ud~��Q?��p@F|��E�1ط@~�y!�����)��w�x����;�����S8�C��pݯ����`|��Ն}42�E�jzFDz����.����I&Bn]�&��n�g�lz����y��p̒�R0���	��exg�E�߭�)� 8�f�+���mU�����X�-E�$La����_���p�ZRw�F���=(�#��\�L\�M�QJi�[���>�GVv�&E5��&!_f�Q!�f�_ )�%�ߵ�Ȓ�9|JL x
b0j��8!���W��?�u�|.�e�ZE<�����{i�~6��9�ãp��v��m�!ީA<�t7�q}����6��"d�29f���=����x����;s���rU"��\���{?��l�Â�����M,ps���2�7��P�x_���s�U�19~M��1cTz��Y�����(i���G\�۝���s�}��-��=ޛ9�ZU��f^桃��t�*��4|z�e����?"�Z�&��{�?��+1t ��{��}���s��h��q�{-�M���Jr#C�l#yd	n�YO<[��v�.���	R����=�w4�˼�	� ��4y�{��f�:P[�'�G6�S����Ξ�\�o���9�h������[M3��s�۲������֟8֠6��z������W'�+��_�����c����w���nT�͖Ϫ-�~?~�d���&���t�=X��~~�n�μ/� �?k�s\A���t�, �a�\H(5�B����W2��7�`EL������4�}��j�V+��I��JgQ��(�!JHp�>[�b6\��A<� �DҠr�G^�Jg���9ܭ�	�fk��鏝��W��`4��2w}*!���R�����a/�2Q\F��d�
I�l�\��KO����G�e� ��/�~uڥ�.8�u���>E���T]�K���l= ���/���Go�V��8CJ*��^d,L��?�`VE�a�@���6`��G"Y���+l.������#�x�<`;~b����)W,>ZmZ��>�dx��:�}A�m��z�%E��j�7°۟�)�ۇ��cM�y ��A�7-��(���{J�������	U,3�vS�lcl?n�G��s~��N��P�s�
��a��<A��E�bҡX#�nq���JsV�3&ӡŗ��^.�W�c�F��ul�8>���o\��$�d ޔc�u����W�9�$��o� w�;u3߽���n$d\w.7�[�inQ��8�rOp���H�*�;܊d�a�� �Z��(iH�j���J��n)��������*��/9j�KD'���[���~� MU�}.�$����Y�J���� Û4�@䉲f;����L��M���6{�-n����ad�0�}�9H��:-�l�W�ݠ�CV���������"<#
=�)�W;qt�G%IN9�wV��(�ŞX�{c���S	vJ⾼G�"Cȿ�|��[�ѤH�^���mY�jG�'�sĿ�r\@Od� 6�Lf*׌>������	t:�8���\�3b���Co&���*sW�	�\�e/Mh�=��!��� BY��1�P��\��X��k�푔=���Y����k�K'7��-/ʹ��84u N���IDl�L�.���� ��>b��1:t@ -Q����G��Veu{B;+��5:��+VF��/rE��g���Ȇh^�#PE�v�t��>�6I)���|�����9JN<���8Pbݧj�4Xɣ�J��z�������R�F~���r��m;ѣ�N���&\��șN�iw�9wN�fO�k�F��W2�+�յ�?�2V�䱬��JL���.}%�Y7�<&���E�~t�wĪ�\sr��$�ėɝw'RIE�K,3����x
r�"�R�=��S�_ʪ��+���zt�X��V,��!쵼���z�����^S�Ų��_�\'f��� �0�=9���f�`��"d�F$E?�t��J�"�������P�j[ֹ��q�]��y�4,��}�˥aѴw6�~%���xȿ�Y��$ktVfR�����8}I��MY�����Z�'������)��&�r���,jK��}ޜ4b\#������[�y��G���B8�B[h��`��?�/;A?>2�f8�\�PO[GI(�FIl͆z(�}�Y���!"���T�]]�uHr�����*�h��\&�b���{y?�FYJ��4CLIJ3P��<S&�L4y���M�/}�Xs���@�����?���}
2@��2o�ip��+b�}M[)����4Ԏ�6yd�h�=�'�H��6�C���<0��#q���� 6��>n�ш��Ǯ	�_�Х׵�ox1%�y��1u�>4:0�GI~(K����i%�TF-�mA�9e��t����%�(R���1�M���*r0v�yb1�A޻vmUv�r��~� L/���&��1r��6_�������@=��l�jv
�ڑϰl\up�ǿ���B��mH�u?��8k�3Am}��B�]=�~��y9�Xj�����Α�U4mzS�"�골Eed�vW%I-�v�L�z$?���;��'�#.�ܭ^�������'1�	%�X����i�y�TQ��d/�U��y��N�;_������t��F��n���3�Dy�oHa���W8�|,a���0�F\aA_<��rsQ-ϻ+��]�R���5N
Pm�˜�--j~�L�%*�oEc��l� %M���~��L4�z�&�E�Y�$�c�QtFU��-A�9?����[D��a��,n��$B�&��^�iBl0�l���m���C����WI�9���. 7��y������E�<��a���7������Bc�r� ���cP���ܳ�y�	.ssZ8�W��"zw_V�Z�+>�������Xa� Ua�S�o�����*l��h9�a���Ʋ(��P8iCl�<xlb���:;���}�,���N���d��u�1T�5e!�M ����_T]Ij A���ݷ��q��,�x�I���(�#����$�#�N�Z��	���������� %no;f����P��¥�V���x-@�����#Fj�{��x��[����`4f�����Q����g1�S"�8�g9
�Pmw��}��\�9xmrMYx�C⽄��~%��V;o,�N��`���˟�������=� 6A���
.�~*ӻ~��+�,=�����Tq��}=n�#�o�-�������*�p�Qe�ֱ@�N��P|N#�#��R;�t�Ο:��u;	沮��j%.��eJ�E��W�����B��H�؟U�ST��,8�:<"0)�:��?�T�����t�vy녟rl�]FKU&����F@��ک$�auk��7&���Y9+�e��	��Y�(X�(�WYc`~��$kb#T'��C�y���bRKvG�?�A,/����h�9\�҇N-��^X��nT��m���t�d��˨��~ɒ�[OåO	+�&&O�g���)Xç�M���2!��)� ���Zc9N������P�be-�HlE��}��ɺ\mR]���*��6l��][(c�߶8?8nl��(�4-s9U
�D���ڢg�:�b}��Na�s��Msj�6���+s/{�vz�UK8��^�LP�Y4��a�HK(j�Pg�>�{F��!��������	/%�A�'���EҞ��&r�%T�)�(�B�6�!�X���>Q�>ݡmX���~�5�B��K?�d�E	{�����3�E';��C��mv�3�޿�m,�)�Ek9Č��s�P�R�RHK����5m'�����-���b�0�F-�ZQ
7!��)yzlί7�?��2+PgF(:=?�V�^�S\o RI�m*ӱF�y,cT9,��߰4]��5����F����)�O9�Vi����$� ���6� 0��+p9�)º�����rA鎥�K��}�愴A !���a�:&��_����x���}��v�j�ҋ���oX?68P��a���� �d[���i��tRy��6�`���ҹ$O�@�+�P�~����ʽ��3Ow]��L79���w�#�_@�hF���y��2��	dz���_
#��ȣ>x�?��K�`�e��e7\�Eۧ�9��Z�{�K:\�����-�N�8n��Jd2����Z,�z ˂�z�yWG�.��&�.�赸)F�[d�B�/˘���$����fog��Gv&�?�f�¹�8Y7��t\��u�e�]��[_l�� ���g���E/��̓ ��U��}��U�HC�3�[HD���b�c�$KV���@��Q�&�罼��+ŗpb���	I���)u !hG��`�щ:�5m (���A	����o�Gm˿�E�e0�T�$��ܘٓ��0��7X��"���¤���GQD�7L�����^�VqpN���+�QlZu���	���σ��^?њ�dc
W��쵀��Sw]�.��ʸ���֧�mlT�7��,�	��S�q:X1y�Lπ�Z�-��VU��~>�k~�s!����T:٢�3�t<Y���q�;�?&�(7������EEH��Kg��Є溟7�&���nȎ�a��D��Sq0ҹ(���'�w�b�n���*x�fh92�>���ǰ"w�#�����!;"�7���{N����O-�tG(6�C쌘�O����cŤ:^I;o��J���m�Q)R�t�?�m��4J�'�%�����ٲ�K`�Ak�1)5����9��@���\wc��3>(�z�SX��Y0h�=�c�����[�5��0.��̩�~ 8���uZ����kv�I�_��*���_떸���k�X��f柯���� 5=�$�z;
^�R�����w�G*b@Չ=�,��h3�Ef�׽��̈́���A�;Y��mr?:� .h�W��Rź�q`&�_`����p�	{��;�;��3�]r9��d-Dw`��h���r[wUm�`K�c��gz#���5�!T�;@��'�f'7j�0+�O�;�+(�c�륇�q;9���Nj����Ы��ݰk|��ϗ���t}l�L¯�x��D�5^o5K���҄��]p%�I��tf��鸝0n�D�A���4ʚ��c^p��>*kZq���Dp+ ^��*]'0�M3O��~�y���[
BaZ������,�� ���vTs��<�0m���d�6����\���1O��x���`��I�2�3i�[.t�=Jر�_~�kF��w�����+�e�d_@�"c U����tÍD��,��r�t=��8R,j��!3J�迄c�-�p�O98x'< ��n�Z�!N���ߢ�Y2��i��îPV�*�Q����М��.\��6;��9>��6�Թ��ҢQ��ؐ�<����Q�g��ʲtm1[��F�%F`^�c�����|G��"�c��]X+zr"X�inIޮJ���b�"ԕ����_{{2�h�|�S2M���[X��l���S�L_\��@!Њ��i��SHo$}�s˛�Pо�B�-��H���$vRk�T{}�{��p�:��a	!,5x�UE���B%q/RC��=^-z�lz��ڪQ�w��:�V�~V�Fy���zq9���=>�
P�K1,�
чҎҭ��}G��wU&�VI�Ճ������	�������q����("�Z�Z֊
�-NE�Æp�8�c��NjB���aҧġKY��  hѐOw��s�۪���&��pTĽ�MF�]�}TqVv4hΡ�gH������Z��M�H�ey#DH>�����H,E�1ugv��h����W��{���������
��� @3������̅K�E����qy���BJ۬�б2��w))h�0�bZY�.iq*�,�V�.�v�ظ ��G��J���(�N��*���6c���_c���Z�b
Z>�>K��%���� 1rMC�͕!;���|$��E�ag��g�Ej.��l�܅�P�&b�' Ӡ�;�ƹ�����YBz
X�|�f�N��KW��m��^��pzW�褈�G�C����s��n;��p�p ex��,�����&�P��� 2^81�����l��N;hG�H�qO�[�訌�p���[X�~�8g�ܒF��둯+R��a_U�a����D&#5 �i�=���]���)���(��V�Zڙ,�h/w*G�=1Q���~�@Ђ�v�(X�c���k2����\Ƅ&����>���1s����s�g�&7���;�d%w�ُ\CM���.��TY����}`J������0>�և�.�7�%��x�a��y����a���g� ���Q�����J�؛�v��L��[.�c����Ql�(b-��������Ƚ^�m��j�M�>�^@� Q�b:G� ѥ��P3�bK�r���x�<�9]�;��&g���%�]�v9���o� l�ۍ|Dc9�a�'tv�%�zO��Z�/��b��$�հ�W�+�c�S>�"~;��^@h����b��0S�-���0�q�\������zSn8uh� B��������0j*&����*����r�_��y��bFYB�Ց��bn?� y5I<�m�����_KL���/ybx�=�o���R�[62�li�
�G�&q���.�邀�*U�k@��m�pr���2r��z�"a��+C3��x�����(;�RQt15��~�֞��X�]�}��f�����n�_�q�~�z �i㽥��_]�k�^�:���g�H|�~�ѿ������!(��cFb�2akp�P)�-�,y��FxC�Dߘ#9�:{G���S�0�%�(tE�p�7��~:N̰5���H�5��u���`��qab��0��u��_�h��6�3�*Hl��7�9��i���n�^V�S9�Љ�֟�[&��GY�֮@��<F[�����O�.���d�KKt5EO��{�P���r�������	\����y۰�yⵀpg�ݜ��V3����x����:�^y�bf��~�9o�M�(C����=��}��Hrf���!-��뽠Z�|����^H���f�f�����}�l��~H�P����ҏ���+�+�j�0�-	>��ҿ����-'��ɜN�0+s�����|<�U��׍�\����%#�E�j'nӱ�+;�KT��<�.�� D���9A{�l7j�n�x�w�����`ӕE��٤��\��B��N�.�$	��J�T���.�$L�15b}�h�|�@���N��p��������CH��k(���'_��Tm2\/���2�����豎8i���T��Ԉc��c����ayWKq({%G�!�p��H��cn�Ǖ��eV�P�v�|���:%�����{�3��.��V��tb�v�Ew��gyܑ�x!]$C��^��c�4b�1� )���H/��-�	0����g6���y'�mB���5�����{�����qCF�|.�"c$����v.pTB,h^e&�V��������!U\3�7(�}�k�>Y�B���D ����h����2�ĉd���g �_�ͥvp�њ����JH񔑤��p���["VR�����)G�)Zvv���L����c���E�� � $&�E2��ASP��;�Y�Yt�=N�(p���^ᑝ�0�?Zy���j�yW�����&��[����<6�#��Nl�Ļ��A=�i=K��{(\�E*]��i�R2ڢ�G�u	9�7�w�r+7O�J��15I_��8�ъcN��b�*A#.�*g�6i��;߹cky�ih3�sVou:��D���o�=>m�z�k+���9y�F�|#�9�K��č4�����-87LRQ1��w��q��^��ϭ�d����ve"
����,�K��-d��̧�� >$*rx�3�Θ�͵���(R;Id]Z���pѪ�2	��/*F�:���,��'�V��b��U�ʭ`��m�k��ԍ٬>Q���P��r�bT�I��y��X�������RL3v��*����s_LS�6IGk����;��/��88��Y~�Uc�d�b��I6���&ڋ^��+��#^_�)���!,���.��ʕ�e\ec��� �\�G�W;���1���5�Qj����@)J"���1m�x$����{ϴ��/�.4�{��|���Hm�5������[�Ȳӑ����#y��A2�Z#$��1V����~"9�ц���o��#Ą��~���c��m��;��^�=E+ҪL�������IA��R*�t�cX��
s)1o{�=���j�KC�u31�З��3Uɒ ��603xi�
���]�l��!���K� ������F�Ԧ&Dz��2I2]���px=�)|mB�:G�'^��#$<�^�� R'�5����,^v&����*��f�uq�� Ky�I���-&D�ԗFb�^ơ�1�}��? <�}Ym��?y��������&ɐ����NfDa9�n����,v}c 5���i'�կ��N�Yj�w��t�Ik����I����k߭2����&����5V��D�X�"�6�/R��w�&�أ�����Xo�����J�风@� )�`��"�i�Xۛg�mQ�)G�1�ߒf�T� �[����«������'�I����Jܯ`����^hi�:��U��A�*�,�W^���%k$?�W~��Pbӳ(;���w�S��2R��R�3����*�M�U7U��E�D�\�Y�����Ţa��8E/�9��Cо��mwdڰ�Ƣ�Pl������C�,��xH\���e�M�'�-H!P@=g0kьM��с|�ݠHV��,M?s!���/���_`�79'��5�~��X��E�Q�8�w��i�SS� ��m!lW�ڽ.kp���Bf�3�IC^�M�7��(F:q,��zL�it��)��:~�Yd՟����"���Iv��m�f�������p⊰�
�H�����*X'Ld"�S�/K�:X=�Poiￎ�����RA���̄��^�c��I��u�4p��lڿc�������zG_-���5����|��v��@����&э��Z?���,f�n���٣7ǐ<|�;D�n�� �`�
b���yQ>���pӓ�K��%�Q\�Bf�ǅ��A/51� �x=�㡛ZW5ޱb�
y��*����-ʻ�K��;澹b�e	o�tQ��<�l����S%��kLc
uoG���t�1ͦ�\"422C�\�nMJR?8�a�
}s����>GG��r�%9�b����t��Nݯ&�R/
�kk�ؙ��
Sn�bI0$�
�k|��)�Q��G�S�����H,�SD��+[y^�ww����F+9L�(�{|A3���<Z�k!�$A����bGE��.#�j�#k+0j�1�&��}c�o�����퐔��1�0����m�~�\jet�;s���a[�iUrL�N���Ún»���b�~�:l:�����k4L�r�׹Y��?�����n��՚R`��6��8t��i8ҕn��<�ǣ�y������*�Kp����tS!��Q���豤����A�[�6Q�i��ƞrI���:�b�|�'�-���/��}i`�;x����EA��
�� &��,l�(_��u9�:/�r�nU,�'�{��v�&"�e�����:���������͛p�j��Pճ��P����ƿJXH'`��~�p?g���0�m�0#n�Ț��J^P�/K�n�S�MM���u�"�%���0�߿�lu���,�0�*R� Po�7�qm���� \���[��CX���''�Y��ڔ}��7xqo"Ň��������=J�#Pk\ �q�����a{-�m���^��U�]����]��jo�1y��2tN)�D�մ�D䯬t� =O��.|��г9��ʇ?�����.����J��hf�wv��1x�4�O�T`[Wj�@A���p��%�UMb*������^�4�/$�aH3�n�5�RH+)@vجl��@А-
�ѮK^���^�5�`_⿷�����B|:�]����!�n���^'v���D�1~x�� �t��EC���1����-�Q>E����l،���4��طb�!ih�,}W�y�eA���K�0��'=uQ��]�N���Ճ� 5"��Z<���<�X�܃�L��jF��F�V����l��/�.2��uZ��<�v
�%�8;��p��cA�D����ٸ*���\��jX���Y��}ݴ��⎭nY����d`<�o�r�E��12j� ���m_1Ӫm�!�n�|���
�AJIx����F�2��o7��� �E�s���#��w�~�_�b��eqJJ�߄�ܵ_�k%�p�ב"�F3 7����z.~���"��/��
y��ta}��|�m��o�A���_���/J:��	��B�E�!a��X�������6֬G-�����W��n��Ճ�H���V,��ry��H/��|�>�E�1�����Yse�3�=e��b���M�N��"LB�� rHO�'��X�[wN�}C��_E�#�W���V�M�6����/@���bW�;?���Sp��LM�|�
	�X�)�yޟ=ܐ�&�Lu�I�z���c�e�c/,>�n�� L��멥R`lF��c�4�����q<�k������Jj΍�,z[OU���\Mn�<1_ut0�,i�2P��H��X��`���5ֻ�d��YIe,��}�0&Q���8��om���!C����@G��+��d\�Q���&;
�0�":�����6�EZ�@r7���t-�/�T�B~���@4��	m�D��MAzG%6�dtA�s�՜�#����r��7�ٷu�?��<��WM�ғ.�\$j�����1�l'ܭ?���G+;��T����F�>�[~��;<f��m�����c_���z&��)��ٶ�{�o�y�:���Kij-���dc���D0Xպ�k]��,5٣�|�ݛ+���e��t��|��)(���� ���/����զ3�.��`t�2:"�&�>��� � �0a�����E���.��A���/���Țk;W�����݈��d[_j�ƻW5n�9�5~�Ӡ����?[�OFs��űe�S��-p� Ʉ_�y�},:����\B$�)��k����w�_��8���w�� (#�\�Q��<lo��Q?�2)c��t��T�]����^C�&�B_;M67�?��K7v"�}�ñ��T|����q:8�������(�y�?_�A_�����;T/m8�[KC�t���g*��Gc�n�.]�3�rrh�+q?3hd$��ާ�&�]5��OCI���8�ro1�`,|���A!;w+����"U�V�YS"��j��Ib}�k��y�I"h�l�����{3�NVU#�J�u� 6�K%�ֽ�z�?��(B	1uC��u�㭁�w}�j<R}�m�d6|��Y���b�ib��|4}OF�-��(\��榴��f����9���W�a}߯y�Ձ�┥/�'��m�(�E��ہ^#�4�ܻ֙P��۫׏�~�:;���U�GY5>%�ݵ�ZT��';+2�+��Il�8khl��$n@�Wg���;`<�B�V��j��'A�=K�/�l �R�Tn5��C�^�Ö�k���f��k����� w�)��p�v΄[,�<�񇑒�p�΍x6p��#��ND��K��D�N�xw�4ܽ�ꦘS`g��2��`|8mY���T&���;�۫��B�Nhsa������3�pje|v�01ǝ��*,��i�r��\�Xu�����ae��5Վ�I)V/5��#����P�M	^��/=zЅ5�^*�:Ɣ�d�뭊=}��ӱ�P�5�%A;?o"�t�[����D����>[�)qga�,�BR����N��5S���pØ�c�&[�=���t�F�@܅�u���[F��%d��N�1~�9���h,�$n0>��Ӂ$��oJ�ܺ�����>\usdѬz6O�\z��x�ay� �)t
2�v�CD�YJ��>	�+mA�D�5];c��� 1�)Nm�/ulJ��E��v��_���R'�C��kv��xRҫI�����jx`��!�$�Ңw|�U61�������m�J�g�jI��E�)� 0��RJ�I���nW��g`O�@8���"C�eۧ
j�8���M��)�\�"$�����$hc������q%�BL�\6�7�`�+^~���.���o#�OӅb@�Um�	��%�s4
�L�=_�`�-���'�F�F�a=�a�4+��\�T̥��Ѣ�*ԩO����G�=V��T��4ƀA �8����"�j^��6��̴߂	zT�A��uF�6��2�K�:-+-0s���i'���X�d�\A��[i&㺐���Xk}uv<���Z({/պN��,���,��=)&��_�([�b=��M@r9*7Â����D�:��B̀r��$k��;����FoYSR� ?�xSw2�Lz����1B�[��:ѐ��24�+������^�QV�Gfc�������{�-��͙�r����#�55X'���FE�"���]2���}���ܺ�;3T�О�@�^��k1�����v[��g�:o*H�]4
�|�pFm��ȒWe<�gc�ԋ@�uV�:�?�'N���b�`�H�ܒ5��־�Җ~q���5����������`/y�f��T踟uOL�:���M�A��M��NEw�OȽ�]�w����jS�k��S����M��7'Ej4be���+9�(�A�R��Ss��SE�[�jQ+���4�=�Ǜ}�6�eTH�B�.��XFt�p��J��4��X��Ʀ�Yq,X����O�0M���xҟ�bN�[&nn��QS1�����((���K��,��Ʋ�1��*	���-�Y"�����g������Ž�;��M��=߀m���Mzab݋�j*�����C�\*��H�ב���8�,�tD�Q(ܒ�d?q�S�lj���+!8�	��D4죘�ս5�l�"���~YQ[��ᨣSNF

�U/�\hڪFV5j�	S,h��!h�A�0#py��C']��3	U��7$`�:6	�&�&P���	"��-��O�ȹU����B�����V$��i��h�\�W�4��D�#�z���JRlv
��ԪͿ�Q�g���8ҝƠ�>��O]z���:����y=Ol�Rf�D�w/��5���5��6V��؋��-�D���F3�v��D�@0G"=�PPo�w�\���z��_y��6R7�@I���;�$9��4�k(߷L��TBj&��#����� :%y�y6I1MDF:TI�C2��a�dg';����j���e��:Ἆ�##[��Kf���?���	��SX�Śׇ(�^mpKNb�����5���?�hjRM��M�g!�m��Fw>%>�qb�d�]��G������i��\㥏Ҳހ�)�RH�+W�ۏt����Sl�j�ד���}����Es}'���j�z?��ʃ�ߙ��� /<���4@��/�D:0�1v=1��0|�Ť������TI�����ݶow���%,V��5T��(s��[�A��k�`�յ�e9f�^�r�R5�E���Β�W(czA$\J:�i57�O`�m �4uSH�c��������⺜�u�P�8.C���Q}:ꤞ��� 1lP�ZѶstn���cM|���tD߄��'K��K��˵���&EW�WS^����J���},Mzn��C&�� cz`�v2w�������͸�@\��y�s@�s`>�>;��/���� �@c,{�������;�i���d��g>X;�N���x�{dŃ���R��C�,�'ۅp��[�	�f�i,
���SX�M��&B�z�`P�,=�k쎙 1��m�N5׉�7f��Aԧ��S�S�v�:���տ��S�:E��O�K)86�)A�S��u�M�S2���f_�FWާ��eύ^O|����}|c�b9ZY:a1C�[�ms�p��TX�-�d����
�s鸚��h�(��}[�2�U���=,��u��Ux������{���m��
X���^`���s�aC��c�'С`�*lH��K�h�FL�Ԗ���	t�f=�]�O��SԑL���<�(��t��p*��Ӣ�*Ϯ��ul9����~O��α� ��ꤏ�@�n$���6mQc��c$2�t��fŧ�����
Z\��N֨���������Bi�7���D��!;P�L/���.��k�;��hN3u�����7P��ƃ�X�/�h%R۽3v�9'�g�����$7��ڵ���M�BG�D�ΤȇZRC��Ț`��ZnEV��U\R�ؗ�H6b�&k_)��g���J��`Ӿ����p�l�Ti0F6�y�ʀ��뮦�g�wX�`�|�5s�J�\��.]�ąb���ҁ-�(����3�I�ir�I;3�P��϶��,G�rLfa���N����o�CA�<Ǆ��r�"	����^7��q����#Y��Ej1%�C8D��upp�!�������ۈ	0'.�I��Nw�<�6���NJ�Ҁ4��ܧ��LѼ�k4� X�e�,-���Y�!��wr�Cq$T&�s@�Q�9���vw熵�>'gÒܥj6LD	�}!_&��G>p�10�������"�Qԩ7���7@!f�J��!7U$_2���jmU��;�WG�����#���r�
ǆ砚���8�n���SY^8/2��*�������/!�@�k�h������Yɽ�{w��%��~18�_)�>��|�_�[��f���a�8jz�xa�F�w������j�9l����j��\Rk���q:/�H�G��!Y��$pFm����Z�C���☋Eil0��Yy����?���
mV ���mי��L71�*�9��"H&t�kP�v貦z6���9�̎�ͳ`�n�� ���V//�nB(l�PW>�	���o>�f�Z��0�켝�9��`#��əyr����w%9�N���$�<n�R��\�y�\�T�1�������J�uQS|�H�p$���*�fN�ə[��Cd�ؘ�(�X�/-{:6�����N��J��p�Nm�f�*k�iɛ
ѝG+�D��r��.h�W��B˔ƛ��*�=�tkt�+�$�tt^v�@��O9���17�VWp�w�8�w��,vNho٩l��E�ִ����i���tQ�W�����/#V��c���� k�ɒ�s+��*D52^ucv��uk�6��d�=Ch�� _o �����˝ ЅJI��>-�'��+��8KbP��ڣ�?En����Bu3�`�@�\O%v)����N���;]x��wX�����(�d��E^����d��@��`t��[U�Dϗ2���y�M����B���~c�8~GS̱<���	%Ϸ�#pL�̦�I�>�#�Sܓ��/�q�?�e�\(���p-��$�a��Na���g�?>���,h�>�u�����dZuҖl��1<� ��>��=��9̚�K�Ç���e��:�O�㜥6��c}� ��?T�b	���_s����@𜖉O�FK;k5Оu��\;L?��R��K ���a�#��?y��y0�k����$����np�E	�TxH��e~���>/�<MF�T�w�B��Ym��U��݇�_��#�*�T�K�,���m�Y؉I`6��n�7#�yjMKDk� �V��Z���`I���Z:,7����tp�`�9����>�r'�%cQ3Qu�
��"y������x��Cs��z���A6����D�7�2ދny-�z2�i�;*J�-�ttiBҽN~��/��ϛ���@$5D��pހõ�E����P�a�2(5����n.u�w����/�?��W���mi~�>{��)�|��K��)��R���m��Z�r�)W9�"�Ό`��'�ۢ_��lzV-Tj����i˱���'˺����+kfYI�R�Υ��\�D���<@R�<�6A����v ��������;�\���w�kɄL��W��2A��<�n���H���+�î\sJ��@(َ����U������?����������0���9Y��6)����3��FqD�@����j-vz!����E˲��8S�p��wQ��j��%,��x��FJz$<�Ԣ.`A"=C�%��4sc�kfa�8d������Vt�T{�9��XRS���l|��
���o�m1�!ё�M�����5�qM��������5����C+�QM,��i�<"͗ҡ�4	�8ؕ�@�b��y�4�9L�gο֨JY��3bF�|޽�4��!j<�I��Q8�{��.^�C��:6*J3��G:�w�e)k��	=5@*taq@�_�R�M5F�)�XhO�(�k��ԧ'�0<���9�����m�W�fz�2d������ž��/�Ԛ8ӝ�y�P)ۿCw&�6���V��w�(`��iReGc��a<������v�D�w2�rA~���Ņ#w��-��O�1�D�.Kڳ
0��K�L�ޘ%\�&SCud��2d���E��e� �#�m�v�<���g
��CBa/I-��_2fb��&z#$�>�١�����|��x�1���������s-%�n0�������_��JSV���̿*�Cd��l�3Aw���U��r��gNCNDP+Fh��vfdĦ&j�P��Yz.������S_��HqIcCx�V6��50�~��r��R�u(�t:	���f��q�8���\�
��J$U��O7
�o�y�L_�㪧 ri��{E\[�ep&afF�����ؖ'��:��S����r9:I�c���A|4�4U農������5��p��]b����~N9�\��h�v�ػe\F�6�/����U������v�z)P0�#B��Y�$�\e���?t���D���$��Y�X��&���zJ�xm&��S�!>�u�3� �������92%M7k;kc�TǪ�Q[�V�4FÑd,�hz1�*����0\�����uJ��������v�S��ry���GGHU�t�6�_MD	�1kR��K��4��S�zHGL���~�/����n7NszĬz`��Ah9�p������;ьr��ay25��z��N�����)B�X����Ud9Vn��7x�Ќ�t#�M=��y�І��f�N^V)�
���k)�X�흩D@)ʶ`3�A$;�K�+A�ۮ��0c�Z���s���^e8G��*��;���k7���ԋ��}W1��V�T��Xʞ���/  �&E�,/`m���Jd��q8hopJ$��ֲ4)|��zK��z1�jd������s	Lv�D(9�XE��nS:;+��O�Ԅ�~P�\���_�gF{�;�!.5�ɶ�O�C�ly����u��_��ڌ��X9�Q�3��h:UV�ԫ[3u�t2݂�]��e�
��?`��np����x�3���G5�#����u�UV��ˏ8��w�`��C���}��6��f7���˜�r3]�>�E�p����
jZ�-���On;�6�O�(���a>[�B�/)�#1�@f�����@����F�x*��u�ͫ���~��0�Ȣ�G���A�G��/$]��6p���GCs��SBU�˦� ��fYZ��8��������.��H�c�@��?1g4����A��En�@4�z���L��IM�$R���6%��8Un]u5��}Q������ݙ�m���mW/^T3Ig3��!꟨��!c:e;�N�j�)����8�n�*I�@�P�O,c������B'�q��Do�b"��!+p�����L�Gn>��<��!��fc�����i�gE������e1Y%
���m��P�rKF�)f`11q����!��kw`Ie��y�&���d��Ϥ�)�f��#)�6x>�4����زZ��;�{�cx�D�d�-�J���v%�J����"Y͔`�n��N�nm|�C䷘���,s�k��n{�A�h4��n"u�5�(�%u[ ږ��gW}x���>���Ƣ�G�7�⛝[�}�k��ml緓��79��x;�ɪ��u �ǫ��I������Φ��`�zg,�����q�(�&_�K���#c�Qj�n
��l̛�joGm�j<�>p�Mr�&)��ɨ�������� :׌�Jc���X�����q���h|�3�T�:Xq�J���*�c->��s��O�˳�5�Dy���2��3��j��N��tV�4T0�p3�XJf�,�x�?� <u�HeU��gIR�2�=�#hEK\e�(Q�>_;�)�;��A�Y^����T�@gy�lr]�Iߔ�Y~4f��>�a��@b���Pf!�\���Or�Mc9X����Q�H�nՍ�M�̋�༲�����R���#��P���,��X�pX��:�ͪea��JFp+$iP�?�)l�`��G�����_��:N<�|��������|�)�z���O�ԄRQ��W����w>$?~^����SR�w�AB��M�p6��]��,�K��iն
ItJ�����~y�w�ԎbWք�+:���}B��,�DR�&��)^OmZUDjd�P��W�'z��!U���3?ڒ�o��B;��ĕ�(��AО�J�[��ð�nס�j���A��H���\;�����e����%�э]6%j�E�з��ݵ����o�q�f$�A�j��t�� ��c�koz4������cC��^'�"��=+��7��eMf֊�H�r�V�:�7�y���\bv{d_���X7t昡73��%�Y�p}�-�QyVW�]P��)3��i�E��a��QP����������2�U�]�Z�HF;���㦼�Ħ�:���A�W��<���c�L������Cw+W�t�X�=�������oɾ�Y�J��56�x�(�ZN��)%\ꫫ����,2�8��)�xf0�u4���|2w��f�y�Kv�G��R��Fq����~�r���oݬ.[F1�u���J�i�u��U��0Q����� ����P��~�z�%�3��N�zׁ{Qi�e���^�]���KU2�����Q�g0^���:�=PW�T�>��'u�M!�NT�x1 ��!E�r�*@C�TMl+
R�7�T�M.�rP��u�h��:t��pc�#��f��G���T�t��dʶM1��K	hj/۳��y�EML�]n4�o���s�V�.i7�!L>��Gي�o(}>�a�l�5Ȏ�D8|�T���	�$n�R�y�v�2�&B�?�2Bˮ��OI*������b�Jb��+r���y̍9�Ҷ�}���.��|��f��y�w�G>��p e1!O�_5C��?������邭ƋCK^���'{��L�Pt��� �s,7���Z#�O��h[�k%ls4���h)�(S%x��#L��b}o����?t�@�����EF�"�7Q�iM���R$w�]�ɪ�"x�F��V;x:v�z�Σ��j��`���£їI}���p`�fYfG��dmב$ Y�%m����ñ�f�C����f�j��:'�Z(�O�ڣ.W��40�b��+�A, -���	]��xe���P�<O����RN�ZTLY���6���i8wQ�_� ~r�
���ە�X*�;^�(�H�(�*��YT,Ǎ66�^�Z�h������I����S �֌3&\�g���H�0d5���.�&��m@���5�	~:�{�[�h/@ӹ��fե��5���u�G*�c�Sꁏ��9��{-�" j'���VU�n<�]u0�[BR@��<�i�?�
���[8=�pH���UZ2���`�SPA�}�����-����~�����ec�p@
<����G�T�#� �+^�'.���ug�K���߼�_|k�/�]D[�vgA1�6?�$|ٸ�;?�_~�}�?"K���J �}:���U����|K*�N���\����\��g�Ԍ��C�Ip~�"��QW���$��Y��N���hK=�]���w�p�E\L�[oz^#O�ju��Wft>E��;�o[�+�E�=:cR��j_���f�Y_U���JZ��0Ǔϭ�`�h�X��NTA�./���M�h8:Z��Wz��P�dZ�-;�C������YF�?������­S ��E<iM-��fC���5ZD6�����L�Ԍ�.F`_O����1�u����G}��.���"��q#��֤��.2@Z�� h�\y���J�y<�9��(���$�td�� c'LM�ę~�s���X��÷��j`���~uX��h��τUe56�	B02Ð��0�6��X���e	Vs���G�R��nS�o�n��X.~��Բ�{���<��~�&��D^ݼ>u00O����}y�y�B��L�ȉ�'�#�HӴ���b��g���P����]��;�i%��4�;���A�� �b�k��z��4��c�#��@/�7߳O�)@���˭!$XW֋�O�mĘG��l�%���"V^��+�[0���
�V�͜hPŒ�(i-�B+HgϬ�F�����0�'>���t��۝R�� ����,��rn�@�amM�O��^0-tHb���$�d/�l^�v1���'T� Z�A��� ��#��`f�����|s�Ϸ=�p�����XU�����l@s��=l�~M�S'ɞ�)xWm?,
q��=CY]'����(�H��AΙMc�,ggp���o�e��"�_R�V��i��������f���}	���XW�Z���?'����P���/ҕ8�)�Q�	��5Ĳ4�?����hڌA0MCl�m�T)YCb4��� ����qK<����Ꮳݚ��d%����[m����3���k4k�|�K���6����^�I��x�ax򷰾�v� ���b}{��S�塱vN
y��{�F��>좑Z��~����1P/O��`3U&������ w�ܦU�ng��	�ce����	��qηh.T��iRg���E�6i32�(@Dy�u�Uy	괈��t}�I�ic)|���e«���ߕ�_qD�*#"�oJ@���k��s��h��غ=\D�)dG�ܘ������c�6{���H�[kj�b��&�*'�{�hf���D��g^S_>�~	���w��6��Ʃ�i�I���F�1:�CwU#���Kį��cӷ���9�T�mN��I�'�p��>[�޹^&�}.$?k0)z�F��$8���g67��n'����i�![�݂���n��>�bK)T��m!��M��U�?/[�P���g�.\ݡ)/���MRWn��$N��Y��H�g����Ò�j��C$�DN�p"�&�b\��Km8�[[Mh胾Ҩ��;�k�>��:�$�A[.[+�=�[�~�"jc�Y�1�d�L_��#eӇ<���KXv��� /2��O�c���ٹ�9޲r>=�a��۬ɸߛT���7�0�����A	�n����=�ޚө����|dg�,m���>�� (δ��
^h��c�f�G�y�@\����A<��B�/�4D`sFث��H~���<l��N �}\x�K�Tp�]E=�hqh�C��ƙ��!!��W��u)/�+�!f��@�nz|����p�"ލwC8%�_�3F�ա�o� &��M�O�3�1VO�֫�S��_��m��󊏭��\r�l�/�0�W��?A��M�p�`BLISGl<~�>N��3�Ց�X�Q���/T��IyVX��� ֿ�#��;q�s����v0��q�����l�exh,uC5�JŹb�F��)���j��~�.obW-�������Uo�Wϝ�O[Z��ђ�Z݈�0�%��0\_�3@�[���r���f}Zm>D�+��D�TQ�}@�jH�\�k�6-�V��ڽi-���*l@+E��1#r3�$5h��s^T�_N�J�߰��xj��Nv.�	e�Zۑ
��N���[��>b~z?kV�V:��XȦ4u&ua��#�4��]�X�:ˁ������P�y����}r���Z.�d7��c��j��3���nN�`]#�b��a���16a��^�D�*y�\��bNT=��雈 OC�k���!Xb����������#$�ƀ���QV���r��/�6��p�W��j�ߒ'=D�-�@l�������p�t�{�}���$j2[cZ�Йb�΋D*{y�X�Nі߀��ȏ(m����"vt�,l�m�ޠ����[�2mYt�j��k[(����I�
f��#%�����?�"�i��S�$q�Y`�A��_�t�(� ����}���K�R�,e�E�p�M��부��A+�$yK�ы��|�ěd��Z���OI�EP�U��\�5xD,��� �C��)�r����O��$})a��\�?ޱx�"9V*I���X>��_��a|��V;\� ��Z]�[�����������B�L�����*�6�LdV��[�a6�	���
�>bN�0n{���y�'CW��%��6�:>Fؼ��,�z ����n��T!m��2�i�w�x�{�KPt7��D*0aו$�o:~(	C�q�E�,���	l<��x�o����N�{��|e����EQ���\�m�e�iqG�\ZjRj���y�g��0Ǧ�>�ʝ�֡�ؔpS�vQT+ )��7���h��a�r�o�^=g��Ne�Z?�Mr�z�)�����?&_��i�@�,�';㐳��7�	k�E��؈�S��o�+���KM��N��|�q/����P�1��4�K�#�йYfJ=s��7MSI������Uɔ�}�D�n�>sa�W���5!�t�Y�r�e��j`2�k�竊@���9�p��ɪ��Te����f�&�
Ȉ���W[����םq,���s.��R���|���F�Z͜J����Y$���QQ�.�5���!�G>�Ŷy��	�0�>!P;W����ʲl�0\�m��·?]Y�eV��q����g���M�?X�1��k���~�-d���0]H�����
�����������"�����X��ص|I�Z(.�_�	������l�i�.�aO>�?L/I)qH���ֺ�ϻ L[�8As�'
Up�����_Y+d�Ԧa�{��KihW,�׳~�DFAk��F�o�t
�.~�Jg%O�����]�K�^g��>��U�ID�X�3��H��g a��>�o�O�Iɲ��?��x&�^<�.����M�M�}��rv�Sbj�J_�?g�����������I)��<���fGHz<pJ��t����N��:��p-����8��- h�1]�[i���h�p��O���7W�M�|z
z�rn��]s����y��W���Si�*�WV2��q��LK�?��!���i��ʂ��8�v�w(h�mb퇠Z���
��&񛤩�a�k͒�\��������qi��BKY+3BƿZ�������6�?�S/������к����;���k=�RZ��y=�>w|w��+����N?�L��T���.gW�t)��1��O�J�{k�/�=�s}�B��7gZS�����[�84���0v�T�,X�tj��n��Y�'�%�9��g�U�jZ9ԁ��3Lj"9�`�R�5}�U�D�ED.�	���]2R���&�|i;R�K�Է� P=�K�`�xJz��W����L`y�B^F�0<�֧�i��E�W��ҽ�S�-�H[Z|��W�o��i�c���c������pDHt�����%G� ɶl1�$)���Z~�[�z�d��/>~|�ߣ����K�O�Z��'ъD�hM��D�.���v'P> �m�_��;��V�[m�*V��O咓1~U��65���lݎj��A��O���Pn��5Ub�GU�q�Ƚ�ʍ+\Rp���r�4��&!9��Q�鶗��sM-�0��P)�?�,#{NIp�9�"��C���F���Ӣ:w(}c�8J�%(m��s5�]�Ң��D���!nд��[A��8Y^���͛r���x�b��Ɣ��eb�)뚷|%�v��_�#p���ɽ3
��~'}~�7�U��n;2���<%�h�ˊrׇn�����8t��ԯ83�|�_QE	Q�a�e,Cq��LJ�CZ;��~�!���U�����z��C���2�-���[.��n��t�qgA��|M@Gd6]>gɶ�B?%�ɡ;b?R��!�g���.�=�i�!J0)���G�f5��x]8��I�aK9|1t�x�J� �%=��ֆ8����$��q�����S����!F
YX4���'���.F|�Qu��!ȟ�Jݮ43u��gXh(ՠ)+��:�{]�mm:��r�L�m���t��M����@��R����o��G	A�'�0:N9���S�#��@W\q
�R[�����`g}mǸUKRObX����:'�9�*������!��3O�J�9{�um�}[�D��ci�o��������n^�D�[,sA�����f�b�4b�'g��*�ef�3g�o�Ȁk�)�nw��|��Ӷ�("Y«nb�9�����iT�r����V��my0;�9�"�<��qy�= ��\ݿ>ɀI���M(>t�$�E[��x�ale�X�iG���VgaJ�з��WL, d������^��?�Vc��Ln����o8Vn^��c�"�d���%�ЦV������=S��zA�����ZZ�?�a}sܳ�z8q�J[Y�#�&Q��{�����7�}�m�,�!�᥸�W牪�yp�g-���,o��(�lĳ���Ρ��y�Ks9{�>|�,�CS��j�q�WN��N*mɬ�+n�gK��HQT\M��v�|��f����\��`��`�,�'H����t��#F0P
@��E������?~��c�t�7��j+RJ\4����c]z��/������n�9:��/���]�?�rM�F� �iu���P�cV;�	�7����	�]0L`����������ņ������*��CKyOL�x�矧�^ۙWW�*�	t:a�j�Յ���{��6���c�������t�ʕU�l��pAz7��0M&�/���%}��)לR���a\����S�QJ[K�.�3v��������A�/'0�� ��	qj2.?�VNN��ɰ7*,�;xR
@Q��3��D���G��*M���,d�^�jEmH˄+��htN�6�4�������������^���"���v	�.��M3]��ڐ2��3�<r�@_���U�h��ݒ�+I��l��e�A�ɷ�}eJnM���J�+�z�M�-+	�E��z	ץjmM�k�gR*טf���1g��+�t�l����՞Bq.%���|��{�^D�Ȫ�2g�j�����ގe6�0�<����Zld)���D	5VJ�l+=?����d52�^ŏ(�gz��x��h))cbt�#�����2�E%7l/�(lEk�bo��T�g���Gl�����'ѿ�gb+ V/�C�Fѥ���`.�1�CI �����P+m����FN,)ђ&����e#ȳHM�����|�*��3�Zq<"*�11al�e.����_�k�]��ޯpK
\�z�!s���9��MKݨ���Aj�݃5�I㌘��:d�х�w:5	��y}H�|Q��t�~/���}�-�ڻ�RLeliƌɡ�`+=|}�y'�pTx��"���3��9���7o��w�}7.�<�%��5Z��(e��e�KƯD-�1�:��.v��.~�������T[��u!�&��`E�doGr �vm1ڸ�<�m���Z52S��*�H�s��)hp� ��h�٣r���>--AF[ݣz8��q/�?A]�����#�7!;�0�%q9��D��H0�/\��S�XN��F;��ݔ��:��J��&��\&̷�n�}������21�r���-� :��s��(�c�;}�a�J��T+6���5�ƞ�>��b#�&lW�H 9��B]�NCaI:�O���'�">3����nDL�.q
�lF���M��+펻����Mۻ�91*�|�vA�$A�>Ѿ`��KolS�Z�%S���H�,_�i�~�¾zx���.o����ʫ?�v���r�U���N�e���
�t)\-��N>���5��w����PE�A`a���s)�g�`J��?Zz��*#�-���L�2�iYسWiDn��%�J�WK�?�nў�E��bƑ}���m���Ar���^�r����y;��B���1B�&d3�LUC��M��Y����B���x0[�"E��F8�~ҽ��S��t�YI����7!a-P�Y��?��?�\�S^لUǑ�S}8U�i*I}[g� �qӣ�#�ј*�<
�0��q�kV��H�z�r(�ڧL��� �����I(8|h8�)1� �'3�K�jL���r`�����/�F6,o���}}@M�������r�O�Q��XT!1�2�m�h�
��v�{u SSJ�,h䇅K�`�ґH��-�R$����P���SIM,���'��-���.ǳ��t<�!?*u��<�i������..��(y�L?� X��V�bߪ�[�ľ��H�����κ?H��bY\����y�?��4rH����g֞�V�l;袘8&���(��L�n^�jx��u��Il��R�8 �2$v�,w��1��å2��i,v�D��a�k̷�S���������i;��L�Q����l��*��Ze`k��e�Něa��2�܊I}�'S�X:��M��F��
�-��W���,�u^����!�-'��Q�q��Z<<�	�(����0���={����%4�~}�p�S0WO�S�S�:̘���A��d\�4]d�H���]��=&��>���85XH�&��:��)Zet��J[R��É���}�^m�1+�w��{ R\�m���T˞Vő�j�0,p�<� ����C�M��K��&!��g�\�����?U�Q�
��E��:+=[qt�� �{�)�0T�a�&дʴ�,U��|�qaw�����Uy
�l��ϋ�#�A�W��#9��8WJl�قA o�i�/�S4vdS	*��f�=^�/�g{�L��\d���W���4(轊Ic�lWIe��4ж�A���N�w�7�qn��?��[�l'�_va�8lo�b�ȵdaO�����8�m~��"�rR�R<�H� �_�
�: 0���ގE:���M�Z�H�-<��L�v�)���!j^�c��� *˫ѿFJ5�<xԜ@JX#�:0\��s.4��6���-ٓ�:qa��-?��l�q�Y�	N-O�&L1�y�� )���q���0\�OlX]�DW�ʋ�,��^�&�v&>�fo�������h?�[A(^��F��� v��,�����p.u-]b�7K�4HoOn�Rb�k4|�!��͡��:�U��>�b����<������^R�V��}�+�yy}����M��V�2�s���~��\�稦+�~�;������H���)������5��.*��.~�r�m�ZZj+W�0������hNƼ	@43�!�?q[�qP��������U�C�ٴ�~�L{L,�˘"�!h�NQ��sÂ��U�C������݁R�]N�+�ՍL�l���DA��Դϖ�F��CSS&��I�ؗ�+��cj���hdh�#ou�(��j�����!�� <R,|����K�$�B�(����[�.�k�:؂����h�¸&��cR����7�zs��}z�u>	+nA����=ܘ"F�.hᔶ��ѸN��>]��V��ԩ� ݬ����F��gX������ ��S0�yQn���Q��#�VIW�
ce:A�M��5ݓ������ȥ-=�"H��Or���a~�]YE�����8�J��n)�@�K'�{�n3��k�P�g3G
 }��]<�Y�ܙZ��.,��r��C��7O0����SګD��(�1������<ď�s�x�Vj���ě+Y��	��u��P�%���GK���Ao 6]���j�f�`��=�y;K5��zV�[��>��4*svlիCO�<�naD����Kr2E�=�/�^J�x��~��=!�� �F
$���}C�Y�C}�Q�:�)��>4���ָW�Mg�=�>���&Zh���R�Z�k��T#2R���Y�^�T��&|�'��z�-��t�
�P�`G���6�@����'�2�$�j���\N�Ȳhbo���p�m]�l(
���NW%����g��E{�3ϝ0�JO��{o&��F��Yv�n�ǿhۓb�a�Y��V���� �L���%G�p�<�<�����Y�����R��O�!�K3��N�乬�̉s�*�9U�')��jV��נ�����!M��n�o�m�����8����8���F�ɕ��(")����x!i9|����G��*����v}����\fD)�pg� 'IV���dc~E�K@k���� �{�H3O�T���A��Q�݀g�_ڃ��.$�A���q�5�W���J��m`���Q�x���(�U|{]Y?�c��K��t�2>�L��z;z�}K2�iP�s��-�)�Gk!��ݓ����P�ed�`,{5Y��w馜�
߃se��TW�2�1;�G䀣��a���`����� �>�KE�}~n��jS��1��5�s��EJ'x6z�pB߆g��sQs
:�g?�#Du<-��b�6U��������q�}�f.-����I P�z���Cd��?k�T]oL�n�.��w�+���~���R��A���\Ҩ�4P�#e?\�m��"j�)	�� "�s�V��fA������f����(������'�Y�:�b2f?���T�Ϸ1���JP��	�X�=�� ə2Z�S�S$��<>ְ�n�Bn�0�0�p*�q7����'�S�9�_�h?�I��#آ�={(���,��|�?)�֩�����ZBz�^2�IT|�C�v;�W�����`�T�.^����}��M�$��T�A�g�=LD��1��C�� �k�0�!Z����!�uFq�ث�o�,�R�:��ӣ�(�)3�F�X0�G�=e:�P]<:���i�i�,w�cKR����IT�#�C5�[����?ݲ�A����2魅��T�4��|�����8}�W"��)��|�.�,��v����i����F8��,�v����9.�l[�rl��I.]�&R��,Ip�rF�h�b�����LaK��£p�����u��t܌`C��^حB�ͷ�z��1v�e0>覦m8v��P�$r%�����.*-�W���0=��C����E�&c3$�=�=r��a��'a�T�f�;��=��;)�9'Z�C���Dю����u���Z�����1;�y���e�,��a�P��~W:?��[��t��C�@�@/.�^K��������z\c��X@y1�W��^4OT���3�.�Ǌ����ˇ͑����璃�\�(����=�(�h����嶂�hY�e��A3�.7]N��R����8�Pz�/����&��_��y�L�:<Xc(&Z(r��q�u�d��i�m�}f�D�S�KO��Ԁ,OD�aq���YbOM&����6�,���SI��7��N#���Q%{�m�}7�ล�k� R��{*z?�#�YMm��i�<�'��@���H��RW����b!���Oq���ݲ�k;���ɩ��l�S�U�Έy��+���w�D��]�.�駜q䍠࿗%Z�C��/�"�(���\&Qk��ۛ[�����&������X<RU`]���7��'
b�s��:2��X�������i�Ai���n�'�����(8r�\���+�_f���ZF9����֩�J΁�D���������e��m� ��T<�ITL�i���RduL�3<�K]�&�K����4��m�Ww:���B$�v��A�ɂ���5��OU����fBg�^.*��V�m"V� qd�����x��yMTcS��l�!	���ZԬ��(�7�A��cH�Y[�{�	rI�� ��߆b0�W��Al��C!_l����F�u�)��mn�cms�P�"�RMFL�!(�O��B�[�~�HLM��{Tbn7���lE���MH_��T=bf#�����q1p_�r�.����b�^KxO��-o��6fu���c
b����Z��0ǟ�0E�-FRf�k�|;l����OG��w��i쵱Ø�#uu�D��l$�6��� �d�t�Ʊ)t�]MwOP@9�pȔ%3���A��s<o_2���f8J���j!rnaj��e�{KV�Q������x��.�6p+�c��~ʰ9u(�N� J�0g����ӕ�\"�lg��( kq|��oV��n�������m�&`\	9m�F�J;�6Y���!�I6����x֬`�i�Y�����'��G�iu>K��֑q1�X���;X�9��L��ڊ��MJN���đ;^��E;����C$��f���s�Ai�9�����4��8��{�	ES �ɏ���� ��n
�	��Vb0tF�oC�1V���������G�1T߈!�pQ@��޴ ��\k�N�C��<�����B��e�0���Y��.�Vň��a,���\8�^Ǘ1a�[��p�~9rdr#�T�{���"�C�G_�v����S����+� ���w|$c�FV�����b�I?FXV|Q	��u�<[�	�����JS����Xѽ\Θ�A����\+ĩ�	j]֏Љ,�E�i��q�<�QD�<RR��߀�n{%���f��T[�\Kp�-n;Ǜ�N�e�b�.���*ޘ'��*[�s=���?f���bw���b��˨�;;�M�������B�Om�o�*��/�|t+�V�%�K@�;�G�W8�1-�:��]� O|�3Vz�p����O<�b��Y�8� qB晐T�⃿ҭJe�D�~�� Wq��fS�����!�i��w3��j}|��(��q�`���u�YO����I"-p���%�J�o��FS�ʊ�]�Ř�-Q�ɶ�?�"�F��;G��K��z��!g�2�Bb
��a�kpK@Rd^��ՓzϻS�i4��M9���C�C������!F���0��؛t������aT:2�{�ְJQ��ئ�ߺ���c�(��؆oa�e�^�l�����Ŵ׉ə#������5X&�C+S�E�N��G���T!K_����#�zd+�6A~�D����nZO�E&���sW����*�,�Ak��+3ߕ�_N#���m$tq��Tz�����N�JG���De(�v��J#�$ mU#���K����`T�T���;���ʋE:к����H,=e�j��9�r",Q��fsΌZ��/��J���{<�i@~���7'�<�*]x� ��"���Q����
���q�q��Xl��D>~�?7��lW��5wUR��i*��T��9�Y��>��Q��|��� Q�����=B����$��!\9>��*:K�M�*~�B��o�����33�N!��g�)7N��]��ޙ�$U������F�t�#�L�����2����/M7/�D��.�$���u���a�Ճ�>�9#�e�*ɣ���o��D�{��C�@7��`�����+
�����!>�)q�j�����7D�$D�$��&�r�aU���:���#�:b��g��Q�����v�0���e'���	�԰��M�I)n+H��x��8F�@�C�7��T�����!�'h��f�,�.럴��7�����#�.�Ĳ�Mdy�ߛF�)wƀ�fH��S*�B�.�+�:�u�Xdvq<�ۦ��Gr�Fп��牼�e=�&.Rd�xh����1T[�ꂞY�=��ʴ�B	��6r~�A���Edx��1�����A�&d!B��V��U_^�L^�p�b���,Q=��7RΓ�r�3�]���݇�7���i��l/ZFJ[? ��� d�F��B�ph$B��p�3[3����ՀϬ>���'~)����l/wK�m 2��qi(��w���6�m,dr��FTS�*�Ũv@����HM��{��Ӽ;K��Z"�����Kfr��G��P�\\�d��V��BL7�{5��e��-�,��s��"���T�������!+�����lJ����j�ڗE�X�8��Q�z(�m���Y���������lF#����'�i_U���7���U��uԽro<��z>� �\���
��Қ�]l��#��`��ÝqC&O�,�*�ǁ�ލ.xhmh���Pk���YJ[@_�T/�C������F`�6���Q��@G�:\�5]1�,�~b���*��?sZ����ѩS�0�JpZ'�`�`��C�=#5�m����٘"q��P-��%[��͐��:�F��!��zQ�!Z:��+g4]0%���ؠ�i�(ѱxQ�z���H��X�����c5����Գ�P1 �n���o��m��߃Na4���jy6T��E31�^�.x3Ɔ*��X���6�����d���-�]/����A��s	IV�W3�\F�]s�zi��u-�"ZPz�+Ow@=e���ES*1�Ƚ'5Otx���f�n�t�݋n���i`�8��R���yS�2��H��c�B ?�X�Yr;�� ���^�R5.�ž��+E�>�j��
�Ť�o��}pho���yܡ�Ҝgàp�Ι��������`��O1iX��ϧ���$�����b���Ps��ʦ���do;&+�Uq���m�@��-Y�Dz�tw��$|JFD�:5��ޓ=A>s�	&n}�(��,Y��J�(���,��T�$n��n�&�."���k��/?
��d���_�a�Ҙ,�' <T��ԁ�	��@�����W��F	*0�7=�0��T����q��H)֨6q�}^̕'×Of,�~�`û#�}{'��:$�kY�,0w��P,�	:f�քX�i�K&�'*��u�5�h�F��<�6�"ۀS�N�ގ�J���kjg�=��g�5KB��W�+��'$�{����E�穅��.k%k7~Ȫؐ{}��s���/+�N�]�p��A5'揸�~�I:��Ӌ�h��~�8s��vu`�.��YM�|�톶%�)�H|,N�N�S�c��l��s�
=\�ܧ<��b�E��Uv��_uM�NZ�(8ű-Rբ�����?G`*�*�E5E�2
b���RH8�s:��v�T;����o���s>��y����뻒\z��Y���Ѯ��^W�qP:>�������x�v�5��-�>d�-t,��F�~�_:�H$/��5��s��NDiT��4�e�:?�E��_���M~Q����݁�,�jd$��V,��)(�o��
(`�k��7_���\��p��B�� X
�ț.5��i��,`���{�L�$Q��H����\�A�Ѳ8�Ѓ�eUfK��NT�@��ˣ��.�X[t_]F�tm�5�"���ڛ��ʟa�so�6�*C�n<k��y���.5�0�i�i ��P�b�y���Aa<�Pzbu��@"��w�&F;NX����t��Z2����/D�U�����O�M,g�љ"g��}�}I\~~�zy��fUs*@�8&���>�(�e���ŋÀ5�SM�)j�ZvZ�l*[���s��..�nNpd�([!�ߺ��ڨy&�{˦�mf9�.@�ӯQ�`uo_=`EFC��mUС�z���։���)�.�.�Jqɖ�.���{,RL�:��J�m�u\�����WY+��Gk�Q��j���TD@�7@-Ħ�9���#�\TSW��}B�~^~��lc?'o����Ha���|���J!��V�"�^?�4��mʾ%�:��т=��L�� �2 ��t92R/���(�z=�nU�R� ���/i1�/o��"P�P�.��E����׃�?i)�=����#��h�WYq�D�����Us����9Ooo/ĳPq����Y$s�{����j��H�V�s��VF�B&B��%ro�{��4��}���`7g�4����G`�@LCrÌ����7�7�HAﮰ����A�����4w�0�^�m� }�"�� �kJ�v�މ��ܛm����o��JC�t+����Ǘ�ʹ\� 5�Dz�7Wa�n�Y/�����`�ÇO��4��	�˪Ҵ�v=��/�A!hy�~������m�31/����j�߳{?�0F��-��qS�����rLm����m��@a�1�� X�dp0�(�?�|0
�u~�ㆆDGTiE�ڊ&�a =E�y�W��oFY'ۥ��1��\�&ӷv!� ��JL0���U���_ɥ*x� ����^a�C=��t���g�+��	#�)3��E� 
-Qn�W��` �}�H��:�R���`+�;}Y*�#�B�^.B�w�,ד��Z��R�4��s����3%�8I�E��@X�k�:M|��*a�c"�F�~�j-��L^����bkѪ�0�|z:_�g(r�_�BS]���q��
���mǻD׈"$rK__ ��ֽ�0���ѹ�?uT�-�=M�$݈ʹw�����8�sQ�+9��9@W��ZBj�*u/C=~��!��$_��B����Ffܿ�]���J�LB@{��� ,�LT��)����'qHQ�iYD��r+gǋ�:s�o�@��}���h��x!x�x�)p�Ud��؈^��F������=�鑃r��m��'^��!���E��3"��I�Z��iƳɒ��3�u���K�i�fm��W�ڳ����+66�|���m £�����Ƃ�'��.6��Cgq9��kZ709/�S�CU�N��=_T+��TT�߅�}�b���%�={��Z�Ë� �@�Lwv�ֱ���@�pjN��K��>W����xg�����˰�'E�"h�r��D��3\w9��R�F����1�R���ᬏ�=&2�pԅ�{�-���ݒ��9?��'�>#�n}!m�|�#��7��#�����xǰ�5Ř���� hS��}"�T����iݔ���ၫX[W��3g��;�;��]=!�/U���ĭ�\Zp�ïL����jp��gK���.������o�� �SW�r�7촢8Ag��?s��-�]DP���.|�"����������������XN���&?�Y*6���v>�zpw'7F$?��˛�;4�G�߶k"-�
�;��t�j���J�;�e�x�`
R!��fA�Ř��0'��,��6�.������^^Ҏ��^��
�i?J��)�67'�Ɩ4,&P���i;���*-�{W��J!>��� �6�j��9E�2a�YwF-�B1(h^�k��H���J꺳������X�1�)Gj|��F2i�e����n�՘"0��{��C��E\w��#��{�
!'L�'�~"�[1���]TRƳ�ǐ� 0zF�'�ǌ���6��b�P�~��
E����o�L�������e����Yj��>��7o�u����l�DMԯ���4�n0��b^���8�{S�sK���e5��dT'EX�$���b���k��D�Yit)5gˤ1zo	��U�������38��2	^BT��g�x��b� ��gQ6��J���ѡ��~��샲/��d���ԝDP�0��,c���.i�
=����I6zE|�Q�ѻ���q�ʃ�6�����`]C��;$����P=)��JJRG�KC�#���/���]����s<�B<u�����	16�KF��1Rl1�5����NL푺�l�-���+J�`s�ڻV1��s����� ����Y���-�c���ǵ��I�c�Jm��GQk$�#���7�帢���f�v�o��wW�ƚ��!�Thk�G�^� e�r�q]>�PYT�s�$FW�(�i)���:Sս��.y��L:c4l�Ҳ�x;�8�Bg�<`����K+����e��S�����> �K�����r�Q*G{����]v�$9��&�e��4�Ӈ��$�����Ȱ���"@�,G����|���sX=�g`ؤ�.�݉ȟ�_�w
�R�`�e�R$� J�^�&�b,0�!�ǟ��l���֊Bɚ��K���#��\�*b��ff�%(mE�6/���N�>Y~�-		́�6�F��]i��m���[9�uf"�p�m����>�>CT+���s[:ݟ�|Ź�<Tc�
ak]��ָ�b����L����J#RC
nIN`����{�X[��\�lZ��K�<'��X��]!�jK�l �3����֬(y�[�M��iȠ2�.3RL2&Ol :�Ұ���##o'H�6U��' ��$4Ƞ6CW|/DL�e5%@ݚ1�mSҰ���Q����e���6�f磖�g�V�� �.��,_5�� ����+��܌J)aKuE��sQ� �1�Cƽ!�5����"!؟��!���/}3���S+wi̡��Ú� ?�������4_6E	����L��8��-v�pox���u	a����F�z[q��`�o�nʸ����Q�P��ơ`d�F��أ�ކ*�c_�^�&Ń��k�p ��R �Af$���As�	O�Wv��v6qK�ՍM�υ�#����}c+G
�u�F���w��d�T��ZB�`�Π^F;�g�B�G�"N��[��]4A����E�$<���9�"ɗٻ�Ŭ���6�kKj��W�[��WJ����
^�ѬX���h�e�̄���-�_[�����S�/PM�B�N�l$�h��v}>u�hl#�mLou,&_����_v{	C8rhZ��Uӂ��V[L
Rn��Մh,����f����6͹�8���R���y%�n�c�́�s�����M'9٬�︘ڂ}���"g�>������(�Ab!��c�5u].��'+��C�E�!�c=}`��_0��%�������D<�8�d\�n淾LBǌp��]�/'���J�,mO�^��}"����$P�ĕ�~P�_[d< �
���>���}e���<���2����Nx����3�zJ����;"49ϧ�C����)0��6Ԭ�������`0e�o�~*資�%(�R�ׂϨeqn �;�����!��*���6p�~n��F�d�5��{k������7�Y/V�%ä�����o8_#���R�!b:�������Z����`b��h8�m�I���	�Q�i�FX�XEЩ�b���7^�Lr�Ʒ|��S[���2��!{�,G���6GI�l��R�}�I��'��<�1K���$�����_����Y#�6cO����?}�C����%(�Lt����\����Ϛ8h���rU{��σw�S��sC�������.���,eӂ��\��}�̵��v{��=:��sF˭��D͏�ǯ a
=�v��jnœ=�x�󭠥n�%��(����Y�(˥�/�e��x2�mx�X��D{B�rc9�����S����R��p�����	�g���7R�х�8���2�'�ʽ��� WP�h�q�JC���K��xCy����oj_2��"����ڒ̑�/bA7+��"ș��gD	��j]�'.��a(�y��U�c�aԅ� ��o]����m�7��l�ú��������-ʩ"F�x�/7������m��ů�4o��/m�O��!��%r�ٷ���poCN�� P��Ǧ����0ד��Ś1so�+�!�aІyL�C$Q���M����[|�K�w	{�ʁ�o�>D]���yo�8�%|`��=x
;"�`��{%t�=�!�
ʔ��;{��=�_����^ܢ\0@X���a2|�(�j��W2���S|�]'߽���;�HtR���2�~��.��eC�l����D���ڷ{�C�pv6����U_Q4�Z���f��I��Y��'�җ9�3���Ne_�&6��ܸ�}�gО���P1���ϙ�	����:5��~��%����Ld'!���6'؄M9��l%և&��0^����L�%��Q�FC92�.��,�:���)��`����r�?�qjq���z�(7u��@����
�2�퓆|�\c���Ⱥ�ި�P�����Җ��<����B:�HU���<��fY�����?�r^^h��$�G���<�9a�����P�X�3�#;����"�,=\oPP:�,"V�JЂ¹&�y�D�/
>����A�^(��P}�6|���b��"%kL��L�1(�h1vgм�a�9���#���nj�l�.|�m���:᯿i��]m��ⷸ��;�P�%讷:��6��֔dxPǨ�,���>R��QŲ���Z-�0Y�P�|�F�h��%8���N�F�6Q�z��+I}��_�����[2˭���#��ނ�6P�:h5��a�u�/<7)�yE�#l���µ�2���߇���)-�8���˝��`��(F�b�!C=���1�n�9�n@S���9a-�G�`���ׄ�@�c�����`^R�����V�	��.�;e��7ܱV�֨�{	�n��A��Q���`����q���5����T�K��L�N+p5c��[W��<U5^�0'T�ɁLm�������]��.�1��c�~�#z��iVE��{��i9���<�iǃo���D�],�� �,� T8y�����0 sb4��3�~�P(�fҰ����s~N�ΠV��C��O�~� U?M�.|B�軺��5|ܿ3���߱Y�1W��u �?\�,�^~mȖ��w��7�,���;-��9�jk�%�4�\���Sw�i�[֐/�ί�>���g��[3(\���2�r	=�p~S��{7�5b}F������fv��(osд�h�:�@�tý��m����5�*�7�foV�V�����g�.�1�hEf��(�\��uƳ�*D�6��<�%E����N�Xy��B�e�$.9�����̩���P9���g�����&���6W�v��NT�ްYB��Fd��̂@��z��N�'��;�4���6�<\.��\Q!2s�]{���t�+ �jI�BG/;vٔ�ꭀ��6Ũ7�#���*޴c�@���['�B=��簈� #q�z�������!H��<n��D~���"��N���]���{�- L�F���w�}���RWF̭�\؝��(�ڢ�dm��YO:ϧ�9�)�����ZI�P�z�'��鍲G��W�,��0NR��
�ˆ�@�r<��t���wT5��B�#�H^
�����D�����Mk}���t�e�"J��nr�L�-���j��!��%I�3�3��l-��ơ{ t;� � �R��V�p(�&a%�M����̱��8�}�*�Eˋ�),�B�}]�Qa����Н��iC��V!/��>[�[��3��of�⯲�cKԺ��@�L��;�y�E���%UfW���y1Ǫ��vZ6&_^,\���*	�/W�S&��0(�$��ԍ� )���E�-֎9y����AA�=x�i��(DJz
��I�w�lS���<�j�L���u�R�2��G.���]��Z9OV�vY���D��z_6��0q8�h��t�S�$�p�^�C�����+�C*]��
룹����ŀ�H�d��D��-��.�q3�Lɇ���=�8� ��0f� ���֌]դAyw�<��aI[��gڰF������a�E��[Sd}�I�O7�[|�t��mh������K0�Զ�3O�Ց�P�<�z[
�4���CR_�Y��>_��D�r��a0�S���E�c�}�a�e���ell.(.S���4��_4�>t���V�e����/��Xl����ĪbW��O�8w$x��*���4���:���Uw����/2Ӯŗ�[��͓������\6���e���0�93^G٣����*G�#�Ԅ���f�szQ���N����7<��]����,�ӃI{KC.�>�����M'�M,:yy��ܮ �����lAR����**�$�q��uJ��� |��~6~�rU���x+��;�u�}���(�S~�H����R�r��9;mqp~4��5�?�ŵ}��R/�'|J��/J~�L1RͶo±e�J�� �Db��>�KvVJ���:?�|��t�Z��K�����W翎��o�����+���.�$y��'ʡ�r��?�����$,���e��X=
�K HYɲZ��R<Y�aC�@�ϗW��L��ƫ�W5@����r�<��X�e�N��2c��W3����׋�qNy�]:f��Ar��y̕�݆E� ��C�5���koB�J�z&+J�og�=�'ӫ��B���H�=p������d��}��T�E�����Ţ�!b�W�1;݋1��k�w�?�&����c�M�,O�|q�H�xwdL_Ԧy��]�&F�U`�6p��4
e���_=?bi4=Ae���r�₨�\�x��#���р�"*��ᔊi�!0hǑC�+m��1�.|D2 �o�Ԑs���k��K]x� �e}W�ښD�X��vϗl*a�_c�����k�;V����d�P��@�4P��)gN���$m`��@o�����Q��x&�V���e~&�ޘV ��P/L8s��r=���nhL9��a�Q,����0�>�p,Ӆ�y���\c4���TD�ZÐt��������ޭ���N��hho��P���I�ǿ��p����
ۈ�M�൱]ͷ��
�`;��F�i�_���H:˨��U���5*MW�D2x�][e����sh��Z-�4������'Z�ʥ�-������(E2!4G?^/�'��p0
��2&܊���#~����&� a����4"!�����;Y����4:[�A��X���'��N(3� ����M�|����]X�Y�c[!\nHX�-I����}��n--�Q"��n�過��m�Ռhd��F�6Ϛމ<���(}�:~t�}������ǯa�IE���,�+ҾU�Q�o������f��W)�
f������؂1�f�?�USb:&�W�Q-�oa���@��h���(�r�W��SN���HY�ؕ����`�Ṕ�p����Z�6���f5�^�o(Uy�N��cR��p%��#�`B4����Y��/m��ct1>
�yll��ul��&���'֬���[�=w��&%7�{=��Q�kd�W#�3�Z�J�a*�P����k�L�W�-�4`���� ��iV���K���b����3�]���)p����7&�dp��B���@�3������Kn��A��'dVW�)�o�WX�{���p�'�����N�BS��W�m���qjM/�˧m����"�l���x�E99���Pe�5���!�����c��k�udT���\^���"��{�2?֗��?���!��m)V��c0�Te�/N������d�Qz��������D����:���Wt.�M�2��V��r4�MP���@l�c@��[���?CA�C�r�0OO(���q���W�b�d�z�;&zy�(��u���m�V~�1@�x)i��l�P9L����\�����D��,�Xi��'u�KVkPI�=1���\�ԭ��@J��QD��S!�7Y�"c֡#��v(x�W��%������^>vKao��,ຣ߶.к}ao��]� ���F�a�-g �[���_v�H��Ka��D��&�hG�;�'�7��L{'�q,���U�@L�9b�o<h#�(�:"x�[aА�Bb[vh����+saG;[�q������xzY�MTP�7k��{�휛�,r��\���w���c�!��]^ir0NJ�C�t�!������̄ȴ�'T�����BdsL[kW��W�a�U��sS�%,�����-V.-���+��Cڄ�od��e9��ae�m,�@�����A�_�!qM(�fb� 6�Km��i�>t�_h�����3��j�o�Z�
���b��N����H���5r�}��Y�xP�L�~Dh��R:j �����%�nNX.T�:p�1�� �p��ٗw�ߋ�e�*?c.jD�"$��VIbrp)9�lP~����ݖ"�<���6�,�WE[�� �8i� >31$)�̻n��x��Qx�C�2 .f��~sm�*�V�)mS=�ru��g��m�pn����y�d��n�lwr?�}@��I�h�K�f�	?v��7�F}�1&��
\��ũ��z0d^�p��N�)���]�A�?ҕ�u�;S=l���#+�o�G�e�����;�j�Q<�M���X����m.�{��m!�,)��l�s�칊O��O�k�6�/���&i��$;�Od��o�83���"H��
_|�qݥۨ
e��r���Z27b��{�s�u0���&�ø+v!��s��;�
E��-m�6�߷k׾�Uc���
�v�o4��pӭL�d�g�\Cś~Iy�����ά�=-(i�I��0�&8gIM�wȦr��V�{�nK��cM~n@���)R��Vn�~폊�1@Ť��-�{�n�N���*�G�#C|�޸�����NM[x�*G������������1-W"�w�Hة��`�)�m�P)� GCT��.�b��Dc�&%���]�T�����S ߙ��3���<�M|j��UV�����2K����)�^O`��my'Pv�#��=��Xܔd�`_�r��\x�外&��hS�6IErI��V��=1���&c˯p�]�J�BE����5�J�]'���j���YhMO�nE���pl��ж�������HUz��7v�����g,S�E_U��\���";��&��1���2�����g%Q'a��۱U���xUف�;�����ۇ.�/��F:��8��{7��M�7j�ML�����u�nq�@F��8�>���x�S� ,���Z�B1���K8X���LTO�$h�,	:\�^;B�?��܅X�����>��G�\��Zl�r���	m�'�\�?\�𫫵��e�QwW�?�`��yaz"S�C��>��G:G%/<[��ZQwx�qT�# 4y;y@`��|������:"�S|�4J;��g��a �$��5h�MS�e9��bp��N���[���;W )�Q��yj[�_�/8�eXm���z���� PR��_��@LoLJ�P�<�0�������^�.����N�dH��E�7������)T�?I��iWM�������]v��]�����������ob�{��`��b�;�X�3g��8b��fq.��R꾕L��^B$�m���}  x��8��"�f�A��M���u-"��`���1,�������{�'��_Ҕ�>P�K^
��w��h�����lpi���n�zc
�,�>��K�B+_vX���c�`��J6�[K� �t;A}ɱ�ߡ��8a��� _y	��^ ��a�>��w[؞��9?\So9���dC8�º�a0�ւt]+�^�m�CM�T7�g��E�94�_O���!�Ź�#ܬ���cyfj�A���p����z��!O�j��,��Q�Z0�*y̬�y؏	���=O��P��C�f���R0��b�X�����y�I&W[Ff�n�+��usq@���9%���d��JX�wG�J�y�3�f�ș�))q	�p���s7Z*f��o��r�+c�\���.�&m��u�����K��}?�1:�j��va.Lg;��o�'�B7�٥�6�U�!�a�:�$������z�H�^]��K@!�����~�3�&9i���� $F�|{(?�ww�] �˕���8� C���W��&����>-qO�Z0ϕ%�Ў�@r�2U�fKZ"͍�d��S
3�0����.n�`�4	� =U��^�V����I��H?I��I�&��d�i���\���#�(F����u*hu�KQ�0�Rk�8�#���cp��c�/~1$��b7�˙�A�``�YLP?�ݙ�v��2z7&7�I���i���f3Q"�kN`O+Dv�?���C��>by�dȱO�L�y艎���&E�6��؅�̔��˿�Ff���|lst`�	�-�`W\3O�ɗ�\r��Q�׿RU'�~������(i��C�yH�&qo�A�#s�I0�lS��Pe�
�U���n�n��X����7�)�AIq ��R���)S��I�$)�t��$	�5Ot����+a��]��T�ׄz+��xu�:�}ܚ2K8&h���l�f�%#ߌe��a��.}$�]H�qd��Af� W�#�TjT|�++��T�)U���Խ�\�[���~|�}!��˛n�s��П�dei���v\y����$��t�X��˕���.�o�C�m$�+�{Uݾ�
V�$�o��f��sc�� 3p�����o(�Eun��li�'�&������N0k�uN���?kqg4�FG��a.�lg���S�{���������PI{TcJH��������hCv"��P���X�N!���AS�����,L�yF�./E 7����T�XdBA�.�R�֎�c聗�-5�o�!�O��ܒY>�k�����f��2�8�����ʹ��0�@ĶEz)���l'�Ĕ�.�IXq��.�!�k�wn=٠[�A5��[��
Y#���[Fo����=�1�i��P�����3�S�=�^Q��0��BJ�X׫.�������w}�;.����,"�Q��AӤpz�V�6�"�ˣ?���X{77f���d�,ɸ��=�'�F������S��ep���A�r)ɏ+FN�hŷEA9'ײ��.�-�>��Y�@!�ҤKX�>>*���
AD�O_�ׅ�=��}[�̀��E��L��(עk�7�x���o��uͱ|Y�4|Z��.�k�!���Q�F��@�6�N|ur�#q�K�"���s�& u�u�!?D���Q� 2�Rk��/�*�;�UJ�ð��uX�{�������hM_G;���&�x��#z���	�=�Ml[�*�`��gml'�b�7��N{��d��K����0�0i��{j���8����y������!��>/o�@.'W�!#*{�;YkE���\*na���OM*᫠=dT�.�Q����!�pJ�v���I��F�4Q��0���=���CK��'�� jģ����������O~�o�S54�9� k�>�X|��x~���Y�CY�p���v�ϩ���-�%�"L�¡.lZI�e�{��U�~��tg�	�Y����Q���{2~Ά�(���EE2��3���1�.��݌ ���D����L���;���zc"F��>�W���%��L}��H�#${�eC��I�Z���Յ�V��|�g�f��ɩf�#��I�J]$>��{ҭ� �X��!�fl�U��aF�B{lk6�o�j��d+>�A_'qj���� t�L)�\̥�Z��OEj�r�2Q�!���X�6>`|>y����������܋%.��J5�}3W��{,m�Wk�v����4��_o�Z%ݱg]av�R�r��p/�jx�}$�l���[$�T��8������ϰЮ2I	K�P�yd���  �e����z�)�ē�cy�~��ݎ�1|O�o�:2���J#v�S����ۘ�/)AZ��G�l-��N�y�}�e>�j��8<���.֪iH�P=�A��&��$��%a�-赓�*���)������������F �7�FM���W7��EK|����U A��%��1l�F�Ic)IE�2��Z�>��K��ڠ�`�\"Eo\��r����QɣK�gZ�V�Z�*�")0�}b'��!�*��k)����'��dā!*5H;��4=���W���Kh8^&�P���j���I���\g���xhQ%�=��`�T��ǃC��(P?�;�g���ɭ��W���@������4���J� ek\�\����t��;�y�w=����q�ُ�Te��D|������x� QF@�lY���^
�Fܤ� �J���,eI�P��7�I��tM��e&�����06G@  )���!�x�E�tl��N��wE�����,��>P/����F�@g�oI��}�Jܸ��Ծ�*�0���zW�A�Fl��������J8Tmqe|56R�ђ�Z:�P#UTx"�KƓ�D> '4�f3�@����(3Zh���
��V��:�h"�Z�LIfڤ���=���	�s8b��6qY.<@d)(Ԃz�`p�~-E�ⵟ��t�"{E����ر�K	LF�Ҩ� ��j��Dg�nv��t�gp�p�jZ/�#����w��b�by�6�����k�h,;�"(�ʼ-l
�G6��A������	�y{�?Ej����k�ڙ�<7�|��P���|������z���(ܶ��_Q�#��Ra�|,�ha��g$ղ8Gv�����@�|�i���k��ރ������q)L����JuI���oM41���O��q��͙�h�P�t��NQv�򏧢r�<��ά7u�Q�p�ǋ�^�����������[��u:�}"xu3�H�:Z�����#��x)=M;%G��@�	U����Z̑ySb���rQ��,���گ�*��X�V���S���\u �;ok'dȧ�槯�r�R�\�E-��!�
^�{�9"��J��4}���l"�o�oؠ�_2WT����䑫��8'���2	�)Fр�P0��":����x����n��i�.��4�����(�Ty��o=h7ίx���u�b�K�xB7aĞS��~�e�ú7�߽K�Tu������c,/�/gG�6�p-�&�2���6�Ã���ÿ�l���.vw��a�sxxr��є��V>D�f��B���;��8���C�yt�,�P���0�p�&o�Җ7�
NT�O�{�WH�oH���pg(g �mf�vG���IIx����&�z���)�O��o|� qn�@�*Q�=.l�������P@�Z�6HJ
;b3�W��<�s r��;f�9mR��A�FՅLj0�|�C�GafC�x�5����1M�������W�F�q�;�s|�����2�by���qS�������_�r����{�$��2��p���Ӭw��Y���S*��������(7Ǔ�3F�҈�aT���mc�/���TJk@��͑a�w�C�}�9�i6�c�2W�\=ʮŞ��H_3Av`!�Э���2˥�<�ɫS�R�]QB>�����V�_�:��1�a�mP�j0�����Ϗ`][g��GwW�6�	�2�<߃F�4��K�g��'�pފ(���\�2��	�q����}�S�c�)�3<|Q�v
�O�ו�_Ǝ�fڜD�]�$���RcO����O�)-����8���z��$@��%�%k�Tk�Z����jnw�aRT��˺��aN�3�cG[~�B�h��CMr�$M�7FzA8-Uӈ�t=��jɥD�<��P�Ϛx �q���%~Uvsf6ǝD�K�>�7������Se<O��2��B���E�즶n��L)�Yк�7=
��7�����E"X�ӖP��+�6��y�當4� 6�h�J�l}n���Þw�����;�e�X�$������ʄ�� ��*�6�%&C�h�)�6�c	E�C�/[�aYP�cޮ�5�Y�J�����!��8bo����tQ�.湷J��>����i���'���E���"���=�U�%ot1� �[&��}�X�+q1�ꦸly3��t!P݉�hI+���o�/oyІ}5��meHl�=�qR֘�����Yt��Oc"x���a�;[ )���Q��a+d�!�*���>��%�i�Rʲ���y~^�o��-�(�%�\>�4�M�߆i{,�t\�&N-H�&��LG�Ѹ�a�ȵ��ǿn<?�����p�BY�4�k�iwֱ녶k>�!ZEO�5-�XrmIkt�X�˻���������(���~���P�(���3��7��E��Me�{���huG/��z���@g�_M��8qW��n(a����Z1�j[(�`�>{�VE�cvdX즥U�ɥ�����C�Yђ��8����ċJ�<�WH/��.��t}�����=sWgY/:����_�:��:�^�W�B��MqO���IK����*����� I&h��=����lQ\+hu��N�;��R����߼�bNZ~��)L��xɭO���Ax�D����f��`��F�6-f$T�n%\��9α_K�t�c�0���wg޲V�ݞ��,�Ŕ/]�j<��S��	���g�1(�s�~�Ћ��:NH�2�;��>�92�Ӛ��V샇YūCOU�ڲ.�mZ(^ؐ�Q���'��Ǔ���9X�ҷD-A��5F�"	=��:�%:���ߊ.�T�@��hr~�����G�D���(�buc��kG���T�)��
}�~��?��
PV��4����ɏj������+�)^�;��u������\�p�mg(3��f ���{�ib<�7|��6���i�0\\�	���m��쵖�_�J/���[�{G廙?@�\��5��/i����/�]��^=����"��?)�q��Ȫ��"ʿnL�b�`��uu�N'6�Z����8|�_lʨ��F��8)r���(ɣf�J� ��H��g����]�B92�~�8����U��)�� �h��gffP��g<yj���%c�J�4K�p��^��Og�QR��!�v����}�jv����i��*S�6�ǡ�Nӊ��V)�{�̕D���2����c�z��(t F�9ϰy}�&�,���V�:c��?4�H(�t��q� s�Ě���sM/d=72�N��/��m�b�.2���?����8��C.�\��#���^�'Ī80�H��T��(����L�*��w����DY���"ܡ4��vI�Xo�I=O�
0��뚻)�7��Y�[���sT�i�q�4Ur�f��P��5�!u�_/�b�N�Ć����+�X���@��!q1o����=��ICF��>G�b�X=��T�Ն�Ց)��2�З=*W;�)�GV���,:)��	��C�b�����Xɏ
��Jt*�v=���q�A�~U T'B'��?������r��%��Oz���kK�l<����@Bo�ޞ)�]�����)m��,�-h"^9o�[��.-Y����ƿ����d���pP ��a�T��R����gүH�pU/B_4�u?���@�)��6{5� ���;� ���΍l&�-�.��.�5�L�n3�y��		fM�ѵ��6�4x^rҶ	��G
�D��%����C�f��y�"��	$o�_a�m��$��.7��������(d+���-���Y/e�^������Ş����a�X���I��*��S7~�[f��wNS]htF���%(߳M��ʾLƚGR�hpr���;)C�x�1|�B��0Dg���#}���l�Q��C����-#���+u�E����>i,L�#즆K�)�� _��QF23ſ4Z~#/��R{M���x��JY�Q��)?���������D������c���a0��6(����Je8U��Km{�&��(_s�I�@� ൩��k~{������$���vd媟��?n�(j�b{Xm杗�l�bB�i� �N���(!�v��UXA�{��$zգ��ލ� �D$����`D�$c`QvA�-�kv�ep7��JɅ6ܕhz�w|�H��CÙ<x����C���i&���4��!���ߒ
��_��]�<7v�B������&W�����Ҧ�p�/�&�O0r���X�n���w�I�@W��Z�h�*t����y����a
�L�D(̀��F�p�y�C�A����dJ]���fP6�o�%�K2��C�s"qE����4lь����h��~�E ��È.ay8�� �{����1=Aq��|�/Ǎw�ս�_��6�_4d��/���c�7e�d�6(��@{l����|�����3V��)����:���^&ND/|��Y��b��/U��A���J�x M����H��IX�ձ��:�3���� d0�����g�;0KC��OYsm[��>�q׆�A�~�x���(����Qd����i��,���n��pT���]�xȖc	�7��2Y�]����C�pp;�6˼��y&�AQJ��ϊ�K��Dv�z�!AaEZ�q/dR����^�Y��ͥ����"5�B~Z��qQ)$����ͼ��^̭ƴ!�c$;j�2�BQ��W�ܲB	$nB��.V�s��c`y��J-]�cE�iK�8c�k�����@N#&s*�}@#�W�O���z9�]ŵ:n���6�iZ�׽g(H\N�]�B�������l:M:!ǅ���c���`QP�qk�Y�u�M�s�!�&j�v�!��a�kd���DߙHHP-~6�����@��!� 0.��������G����$�����`w��w���IN(�YB��<��m�â��4<$��!n膮�ve���2M挳��`��ڋ~JV#���>111d>�����7������<��;�$k�G'`z��dt��Y���K�=�p������,��Ȏ� YZ�GRB�OWB:Q��	k|�1~)������"��J@<��ԉ�M��2ю /F��RFrCz)1�6k�	�>(5�`TQ��v�㟮���������!໋�U7����R#�n����)t/�P ��2�'�7m�P�������Q�G����V�\Ϣ{�!�wN��(�mtH��J��Ý�[3Iu}a5�����Yb7^Qj�4)��lgB\ǿ����S�A�+�s��2���݉xm�MeD�}Np�^�,��bٖ*�����p�eyzgߟ�/����Jw����n�+��S��A$�Is�M���;�]
�~G�eQ����S_�K�����Ђ-'�^�a*�����La�KIU!M�;m����v�1�Zyx*-���J��e�%�|G�p|����9!{��}�}@ܼf �O�Z�W�MWsu]�=)�X|��NV�O�-[��r��ė�3@������!���5P���R������p��W���+$�0�8r��b���j�@v�U��D���/ӽR_/�5#(�\�s�f�y��Q~�������)��lw�Ny��>��z� TwGUFy�1^Q@�/����ȳ[�>Cx{H���EIq�)��Gڙ�l׎�N��r����~�f<��������K� �����a�fNIwE��B��waX��k�R�s(�y	�N�4�����vI�q���$/%�R=�v`K/.<56~A^t � N�ƣ)"���ML������=1�$�'�^�|
`�x+��<2wN"b�c�U*�^�6؞%�����s�d�.���ܡvvCb�4�鳛�tW�RB;����g��⩖�Tgc ���pf�t��Tl�h	,�ۆ��Fb�.�T��"�[�~�������ب����w@e2�#�)՗��u�|3zB"�!���B�m�y��@�����V�=k�t�AM}m�:Z�گ$��8OO����NL�o�,�L�yn$�,�J��ك���\g�%���:P?���qu�+g(�ץ֕�s�7����0È�5^��tS柌�,>��U�\�R��Ϻ�A}v�\*�U�Y�HS�*^�S�z�TC��ԳH�ePӠR�k�m�������Up$QDT���ˊt��������(��Y砝�Ĕ0�6W���m�Y�]a �H����1�鷇��#M�HW�|ɱN�cI����ߕE:�N��noi̕-Ϸ(G�PP��;����p��y�̐ET�ֳTģ�s8�����*� ?κ�1 N
G=���n�$	Uu���N���!�M�2�*�.�_�8�7�+�k�v�CGì	�A����Vis7�0��b�FU��Q
r�$[@�V��i����W�b���O�@,[��Q�G�wu�P2s^=��C�F��WP�A����D�@���/���D�!�<���a��үi~�l0A��=\����th�O䀩w�lǒ^�54e�����A��I�:k�AIl+g�$*��!k�B�Rؕk*E�����T�t��C9(�^
�q&$��=��b[-��T��ʚv��e#F�����h�o&�E�`��n��➢,�r �������]t����ũ����]n�8XmS�A��@��q��Y��,:Q�j�A�<9~{*x�U��5�}S�Mu�i=`�ܩ�>����t΢*P!3�0;�њ�ٹ��Ԫ��s�'.�B�"��Af�s��]�&Np��$ì�k��:7�7���=:0g{�a�i��@�xB�\d֠�r�IW@��N�I��$�6�����{�
�L��)Y-�h��fx~���l|Y�	��(�:Q1a��n2*�|
�a�ߴ��s4TY�P��R"�0�YC�7B���8�j���m�@�5���dcӬ?��ϯo�+4$��מ֍7��2����|m�`غ3b5d�7+'��w=9q�T0�_Y;P<ȿ��r#-˿��g�a��8��9aM�J���Ff3��BM��Q_Z�	�O�f�����������-r{J�';�y��j��4	�FoAM�9+�D�:H���'p�gX}>�(���S���Ci��A�����>ѧ
l\2<"c�w�28�������e���v���D�3�@:eȦn��ρë�������3Sɇo����x�3��P�}|��;MY$}�1`�8);f��7,���#7J.��V{qg8>�W�l�/ӎUڒ��O���Ţ��T|o����|=P.�ȃ�SHD���O�s�O�.+3�gB�(΃�"Ȏ\�({aw�J����Lm�_��C�r���y��"Z�]V�CJ��l �U�0#��5V�ӫ؛V���Sv|u��<�ylV�ZȢ�V��Y*���*`^�Z$���i���T>�����a��nE�^�F�k���r��p���T�Kb���="s�Fe�����"U�vZMd�P|a�'������	�ƮW��c/N�a�:��u��Hє;(u�>�q���.��re��\h���L�����W8�:a�c��??6J:e�1�A�V${-���qFy7F���g�XTE��� 蠄𐲋���U���J�5��OA��Vý���{�4m'��y������n�,9Bt^��W=&\�[�s (S��;"Sy��H�U2K� �t�yigbl�ETK�����c.��$l�+�a��'C�]���y3Z1ׯܜ$��Wh)����j������{�8��&�Z<��+]&M�>��x���`�m��R2Ikn>�-��7T�"d�<!(����z{uL!���+�Y'4C��T�c=/X`��V^3��x�(P���7��Q'���@���T�p��u3�S+���b�1�$�d�[)'4,ey�rx��D*�DI]i����r
R��r�V��L�
9��ɁX��?xM�aP�gY����Hh#��P8n$���S)��#��'-�sW,e��B�!)q�
�H�η[����{P�ޥ�ҳ�D.�B��}�w��qYGK5����(�6'�:$��y*J�@�����7?��� �,[Q�rk�3�	�,�9�]1~��P�)W#�;��Y����ʵʉ��/���q���1��E���A��ݞ
I�2�p�)��������9�l7�E��OH���Rn�<8~F���@��cq�\�>g��k��>�$����q9�7�(�I��Rp��#�>Wr�A�甈�U_;�%�NE��=�4�p���r.k�J91�{G8�*'���#�2v�^�
�F�n|����|j�POzv�#�P�p?��)6!�O�	��U��= �
 $��8?	��-~� ׻���W���;=r�\󒕝=��]�H3���u	Q��bl;G^ �.u���m�O�+�r��훖P�R�a��{kEF���'��:��j^~̟��6eW�f0� 3�f0g�Ŗ0�<��;Puz�+�Q���tu��e�*:C2����XB�Ʊo-��5�d�@sC�!|}��H�@���p9��g�����\��8=�[c�>��-�M�;U\k幄8t�^^���"�/��9ķ� ��n|�֡Tޏ�7��V�d��K8��=��b�6TX����$�+��|n��ࡩ���M~�I�����ɧ��@�ʛ���� �|o����D�f�&���I|)��)�4�;r2
M�{爪Qy�z�o�TS���}�1ƭ'�g
��7�����/���6.ɗyԧ�f�qŏ�l<>u�~O�v%^/ʛG��p3��21h�M�F˯+v$���v��F�<�aH�>W���4�yE\�C)l&>'C-��ʦ��"*��A����_WX�Gd�`��vs~��6�6�*��H���Β9�{���tme	֕^'��-0���E�I���"i����4�<���0��[�*�R�h	)t�ÿ)��$I�����:���9oӾx� ��#�g�7�2lgA���1��,��5cT��W�(S�����_C���)���y)ct�3CZu ���"��Xj+�f;��#nB�7��)��c�=:G�6��L-z�����j�iFT ���P������{����d9���^�|F�h6}�1M.��u�&L���t2z��E�|��jY�D�Ù�qB�$�T�W\D�e� �Z I����o�e��'�����w	|�l6������a�1p�������~�':��Hh�\ 0=@�X-An����͑��Ve�4nHcz� �[�Ez���7�@!�y����m�(��h�&�as�X��j��U���q|)�G�^�h�4&K�g���0$�k�er�P�T5.�3\�����,qAA�LXsxhae�䂋Ĩj�h�r����MO2�T�4�&�n��/u)b�^����\�#yn7�c�r�U���9.��epVA�1Y�a�yj���L8'�.���_�,�P�*���Cb�QRl��ƶ�jd�_�W�h���gP�%`��4����9��6}�'(�nr��B{�-mB�hɝ-0Ά.���9`@��*��],o���	�{>��P�<�l��si\�Kz�0/>��އ�*��1�l|kK
QM����"�8�����A��"e��K�G~�Z��-�Mr�?ϨȳT��+�es�	G&�ֽ�2	��C6x�t��4�O�	k�/�%�3)���m%"�I1Ց����B@�Q�34�3�Q�GN����2`Y���O�\���φI��Rjƞ巓��I��zS	���2-������y#��3�+��R�v�s��5Rn`6K9O���~l�_�l����,��]|h5��|�YX�S
#�d���Ҳw��H��U��I�|��l�}L{���k�'�r���S���'޼x��*�z��? ��r���+B�?i�����J� �/�|���/�~s��X�,�4��>�y��c��>��d�끏���m1��	�u��L!(�~��ڵ�itT�3*|YZ����D��L�x��L������u<N%�:��͝��%YzI���8����F��+���D/��u����c��/�r� e�JE�_I����|�nj���[��� |C�r3���b}'��Y�Be���*P��[�:Ĳ23^�ƦJQ�0ₛc�#W�}�lhp��"ŻW,ޅ�X�mg��,9�T���[qE�V���PC�
3	�S���oo��c�	�?���+���q_-m8��m�v�_����X	��=r ��eNQl�IǣC�Ԫ���3D�1�,�Fvf�Q�v��@i/5Q;���-�-�K�:0�`�֌�e���t��,�+�PS'�FS�m'��^�hv��ӏ���a�!>K���fn�j �$p��Q��=�}� �1�+��뵿5���T�:�1��_�d�b�_�>��s�m�\/j��ف�"��۶��b&��\
�=_��Q=��AKn��i��"1n�����~�v��'ז>d�{�}��p�R��p�S���~0v4@E�	�
A c۝��g�_��qPI���:�<�k�����>�x�yT�y�ղ:��_P��������$�>�H��\f#�>��C e�<�G$v�s��dn(h�CX e��Z�2�G]
{8��v���uS��{%�s2կ5�ZS
s;�����9]T���!�k�O0.��T'�q}�%�楆1��6o+{����FU.�nFҜ�����v��)�֮�����;5ugYi8��0�T^�λ�e0�fpy꘯q9�����٫�nk.�G�)}$��=�rYw�X�:,�+��e��ǈNU���Ծ�ڊ���5pL�J)��Y�.�=@��)�Y����7@�2�j_;n�Qʶ�V�H�0$���%����n�l)��Wj��	��
�1�ℸcj����Ƭ����Z$���+�q������@�>P���F�U��F�GLp�w��>K̘�
_fxz�V/~3���m���N�/�X`��r0 2�6�ό<�gY�Q���^kw�WQu�<��� 5��Π}u_��C5#����@ �(Q�|�6	K?Ъ|��b��ь5E�jZR�;p��'���8�y�Y�D�Xb���狽�)���zL�*�F��^�M�ZS��Ӱ��3k�r����W�F��z��赾�C�	�I�U�O�r���2�fI����A�d�ݝ�q�ifu^Q�f��/�t��v����fZ��Ѣ6��M#��A�����$�����R�^�h��^���NB 2ai"q��P�x={إ.��xg�IJ�8��5/#ǂ��%�׌���{J�#��
�S��O��n�k	q�px$+������T����Y�vI3e<��f�#0��_��3�3��c�:6V�g�ɐk��Q��|F�?y��bc7�_���x�V�CO���gth��^R�Y�8��d8r�eIPJ9>�:s�v�:�g����cIi��<e��8G%.��P���Fr���` G�$�t��M����H5ɞ�����5E�D���Ԗ��Kj����/USe#=����C�sϑ��Q��&^J��ԕ���1�[�+�
���Q�`�V�[f�R��'�$�#�X��$y���,e���MA�m�S5�Ԧe���&\<�y"V߰<�?1�F�����0�Qs�6�O���N:�2�~�m�d�;��^s�ـnh֯ΣD��U�ܔ�D�|�P�ZC�����R��J��T�#�1�eǠ ���.�9<%BZ~�,��\Н�7 �]�KӲ|b���a��H
��l��xR�o�;�%.\ѷlg�>h-���YU�ssE���4K�\���?Ly���pZ��,Tt��	k�H���>�[p�&*�����5_б�M�У�����"P�=*�Gi�N���C�؉��W$�IՒ׏c��[R(��� �4�6���E�#'�͢�~nZ�NM2[v��Ԛ��#�"pU�犇闖ol�������[V�Fj ���?������ǥ�(����m�P�҅I÷g>eDy��/���fń��st5T.����e�w�D3n[��By%�h���hb���!�Q�P�����`�	+��`�.�uLj;5�ٟ#c�*ji[!�n�{�o��<��5�6�at~�b'&�䝖/�P#~Cv�S��ge����Y3�Ga�,��~H}�!x'�8b���N��0���(	�ŷg���葰�z;VXܡ���� �'ڟ��i��V�Q�w���I��U�(%�m_��$5)g�k�;/�$�Ǡ#���i&	H��e|(r������ePwCE�'3o���qV�W��U+4��m �	���BO��Ř�^���A�x�W���$�E(cYiP2�)QN��j�1��t�g�M�9 aUJgbi�x�#ǻ�BR �yp��2��&�߃�#��+;Ol��ԉ�#���卻l�]�-��`�\�wڀ�*(�q�h\ݳ���r�`@"���3�d�e�Lgq��b�R�uP�5�#{�j�r�����xiG���,�C�a����uϡ�?M	�qKn�����lm;��U9�*T��䏡���z4�w��Y_����sgG��ͫ���R����]cѫe������*k�"|Hb�̴��%�|�����A`��%��P��t��4U�W�k��F�N����C��C��;o��^��Jɦ|�=C�O�n��ij>9�9�)��-3)�B�!1�ܫ��2�C�/�`;�l�YF��L��|=T7��>Ƞ�è k��������i5��ǒ���|��I�:��4p�6�M+�x�������h7�?ta�
����Z�Ț�g�K�)���U��>dp�Y��n�����F�O��w?]�ϳ"�ҽ)�Ь�#�å�]q$�l�b���P�laU_u�ˊM%��N�އ����.��(�{���u;Nq��^����q;�fbݹ���e�:�����ѯiy���3B\HG������7���z��N���Y0�q|�A��4��p��Ә��.�k���^�G<� ` d��K�aR�
?V���B��z��2+eUG](��;�F#�%��dQ�KR��IYK�F����+�dV?A��Su��0�d���6��=�Oamw�@AlS�=T�W]��}��V�6w�Ŧ��@n&5��E���E�K�D��D���e�^<`ӧ�1�w_���^��(K�?:}�w�C�Ve�;L��b&��ҋ��3�
O�}��ж�J�<��������?)&���7�]\Фȵ���i�z(W�������(FOm� qt�Ql*֢�l�k�ޅK[8`��Nw�-�Y��7U&X[h����G�@ޭ~�����x~1�q׼������Q�ܵO�1�ӿy��NC�=�$Hu��wʡ(.��,;Y���s�g&���v "f�oX��d��/�\�kD(tKDG�_��ch��X��S�>����A[���Q��i���=β	"w4r��E���	�"�^�eoϙĞ*��[-`��B����٨����?(���J��K8���ۅ�SH�.y2!GA[��X�<�1����G� �`�f���VJ\Q��O{|�O[9ԭ�7�ax*}y�F����;��m���������WR�(��i@]�	�߼s��.�bڲ�¡*�.zçWڊ��A=3���>���Wm8���3R�T�+'�#�\��u�Z�����ỏ@�pwd2�=�g���{

�9���v��E�=
[T��5|�W�Im��KC(��}����Ԭ�����M��D�mX�������eH�`����QI>l�\��쾸'���O�J �˫�M�O$���':fY$� G@��qTO��?�Q��:��ަu���C�Sg��T'�.�V��O!�b��N�Ş�Ԉ�������'�$���'P�85p�O� �{�з�-�LYO�739��Hd�G@A�����"@��C��χ�;�r�_h�Cn�b�VgU޽ �Pշ���^!|����Sͩ�n4srHp��*Gf��<C�[������W50��ܯCrj����Y+� 7�9ש���(5��GY���9�\>��=[&i.���q��f���k�������zevɓ�B���5�D�OY���v�;LK�Mlp9�t.�?��`��V*111�=�B[׋��r�����b�k�ɉ�ekuDm��w5�jHA`���=Nc��=X�K�KpKU^�#y�t^�?;꽤����@�+�2���*�#�s�l2����1�Y� �*�!��h��'O�֬K�!S9�Y���
"N_R���lE���H�Cd%����^�B8ݚh���IۃR�h�-���K���3�#�)��[Ouq��V:��!�؏�[{�(�p2S�7'z�B�'�� ����I�h�5l�L�|�e� ���v��9��8����:ڞvr���� h {�}��_ˮ?��m��^��6wŚ,լ9�CZی�~B�ݾ���$Z�g�ŜTI ��3R�3N4gƔz�獹�'i^�l>���U.����A7'Q|����a�ej)Hf�8����1r���s{��=�\�,Ŋ�G��ԶB@���77̶t��}v�Y��B�ݪ�8/�k���Ӌ���vCS���5�*+ԇ3��k�+o����O�Β$��A}�h:�
�7ɋv��+zB��ʪ�˕�����õWx8N�wR_�G3L��׍o�����f��"y�U���d��˯{yNC�\g��#;��{SF�o�0�\�D����&��ހ�t�EC�,BR�'��\�K��)E�|��
pS���o�h8)�MPa�D4�����Se��n=g#�u��x�Ap�Gr�D�Ǽ���ܼ5��|��H�����:X6�s	]1i�N�$\�v碇�q]�9�H�r9Bw��8���NJ�#`^�g�3!W���t�?�s���$��7�l<M��g���io�ƚq�C��B��*�loH�EN��ώj�	e�=�>B���k��	�U�/!<�#9��s�3�Z�F�a�����n�v㽣�4�rE�бzh�
`t������|��nD�P��o{c�V>�h��E����<{ego_��s�N$���0�Bs�v�Y<�ӏh�*�����j/�汅T���2���B/�7������@�����N.!yI&��Yt.$���a{t�ZΠ.���z�iD-�n;���g/�<	��Cg��|W���Z@L��qfp`��,��=f����*~H���&�k�ZP��q㱯�����X�y�w(�7]#����Fs�\=�J8*j��K���{����g��3Jf�>٦v�g%R)�G�0C�W��Dm5���֨��Z��2gp�C�g)<�f��<2͐Ά�n�a�ePV��7Ef�S�)m�N������JO�ắ��(a�u���7~嗕�bm��8F_���P�>����wCj���R?�e��/���!�m{[g�J�Ff'�����3�7ˍ����ph 'Lk-M��kT�쉷�/���:�c���tE4�7�ш����]�(��o\�I!�7O�_��b�͔W�Hl����Z/���י�!�����<����O?p$T%�%lTs[�7�-��焖Ǔ�2<��Mic�rH�Pb8~S8t�f���<�����4˗���R'���Ps��*�霂��Y��еN;5ס���v9�݆b#�x����ʹݲ��e��&�Ea�K��r8.>��p6;�����If]�;�ў�K��F�� ���+�L�>M���r��6�V�m��0;���js`'��s	i^ӄ�=����)L��fYo���q�bj�Hr|l�gK�3[�u�5zX�<��*�?>���\�N�Z��iZX�o{��뫡�[ݼ�5�����9��O�7�b�o���F�^��aUu�+D�X����a�XcDb[������C��J8jU��B6��pA�
�#¥
hY�^�*V- ������+vr�J*����i�w�߅i�c2���H��U�� Ng�������Vp������K����fsf��yh>�>��6s0��"����_6׼��:n���OY��x��[���3U�iB0� Y��F#k�V!�H��S��Y��/i�.j[i�o��.�L:C�2�zY���q�"*�ܓ�$�����{Z�p3���ڜ�Q�þ�q�)6��r���)�$�"~���|���ʗ�Wc�/��gܠo\���3���p��t���x2�{�:�b��)I���U�z͹>.=Hئ<u�������\��Wuq���)�#]"v͈��N >$r��� ���/x�Ð�'o[��r~���Y���Z��g�GutJ��Ə�&���)�9��j���'P��r������i�}�)���^VO�?�l���\��J���b��B���_�9�~��މ���W�_�M!�����zq���2��J\@�U�'�M�������M,o�����?e;���er@�!��0)tJ8��r��!���:q �?�T���s�����I�7��d���\{�>l#}vgwܤ���+�Q����hT?��p\�t->���ċ�����E�yG�C<��QJ�V�6Ё���D۸J@wO38���ދa����%�2Pn�ɖ�c@�� �FR���^
��n�EX�"��[q�f!�L7����E���J�Gye>�+9�^y�OP�b�|�g8r;`K4³��C��=�W� ����?�3H,�5��\ç\��oA\�V�[�ĕ˞E?�D�i�䴞��mV��1h�웗��a٪JO/|��ޔ1�(cHc��u���	$��-��_e_1�����xD�����!d�2ܿ$2<}����o��_�+N}4gh>����.���������gHo�f&�-�ؾb�tր�7��VT{�" h��.h~�˓�[EDr�o��E�82�IWϰCF������)��(�|�35�X�O�dcU	�3Һ���XB��nJ"�����<�8� 3doJU���.��j�����3Nu偢*�\�������^������
K��h�;��ig�a-#�Esb�쵄�sftо��N�{c������yB�f/���\>�M]����yXUL���	z���x��q��sT���^*��e�KR+�]�d�иYJS�/Ԝl�4�L��=N/� ���0Ո�E�S��E�1Fm��W����A�䧻��F�J��6���3�Xp�8��A)�í,�Ԕ��l)�g]L�{�-����/��B�I�M�H�w��;�5�Kr�y�;d�	�(�ǹ�qɿ�-�v"B�G�qaq#PdCH�$ ոk.N�`�_�K����ۥ�d+�=C���Q8��:��)_���}��Ɨ.cјP
�~�ڄ����I��Ɔ�b��e����:��tr�v�v��� k9�\�?C!�B�m�$H�� ������Q�h�K���48�����"u�����@��dO�; A��MX�|���6zl��ϵ���rmsP% ������V�#b'E��/��(�{�� <����=F�=���B8�ǭ	�)�I&���T*ND�kd(e� ��}p}�E��.���w�� �Ȉ�KU�RX�lb��/�o�"0`�RIy�Vg��ѹ����ȩ�!�夎�71RQ��fYe7�B-Q�H�q�{?�J��9�kģIA�݈I�j�nBb�е�K�m)��:[U��h�q�N3�Q��-��ϥ���W�>U*z�2N�����]��-�:�*$ȡ��Wr5�z�+��6}�i#�vT
Z�fT�2`p��#��_��6V.@L~e�!�b�DuҔ9�8���T'>�8�c6������UNƸ�Kij�քB��^C�$��6�� �n��k2�E��ƪ#��4��'��;��0�X�o-��>"[I8����e`O�h���>aY�;�6RZ$�NB�p��g�����-�,�+I�r'a�R���V��4Q�6^sH��lQ����;�cVb�β��3�=�����,��[��ֻ�Xc.�$�u�Q�Hk�drг�X�
A�6�q*8ª� ޲�Zܤ�|��d�<�F&v��M�"���5z��q��a@��I]�,Iю�;py���ԭ�͑�jn�^���%��z���n{��-�L�(xU��͑���u'�}��Q9*�+g��e����W�4:?){D`�C�Ή��w�
�/��k��a��"Lc�N��W8�� �T#E�E�ߵ�@b�D'(�g��4�'� ���z��t����Kp���3t�=@u�	S�έ�zD�ݼI�K�&<�����^��aU[,�aF�	�����r�����j�)���N����n~Y�H�#��9�Z�Yf>����ݮ�������� Ӿea�r�j�tA�%����I�=��� T*�B"�0qo�����f��t����F~�x�W���4���e6�J�(��+��r|"��S](���O��m���5�BT����'樊�6`*U�!�FءH{Y���قR1e*Z���BsGʍ	����ӫv93Du�J� ��Q���a���o?8|х�2�˔�;�&�����!�����'�>�,��g��#��f�$�}�Y2�ǃM�Fx��\/uI:�Z�U��QVaqy�1���������]���7i�j��bcPhF�Lwx}S��  �ě��i��J��f��V.������V���9����J4Kr5�(��H�pzm���XcWc�-�M�=�%AY���T��2b܃��Q����3�'��_��j��w>^f�y޺�W�0������W�������4��CP�9R�B��- ��w��k%��(WVR�|�r� ,lC�9�H<�\�Y"��N.���!b�?t?:
�i�h��SoQ�]S�5G+#[m�z@W��Z�_�bJ�v}��8��8�!�� ����L����@���%B,ќd�r��˘ɘ	68��L8ba~�"?��>/W#��pM�*��I�kX��j�-LyɸYRڨ�0uK}!�{�~��N��j8:��&Ѫ�r�i䥚��Q9���/�xcf��f}����"�e8f����K�v<��u"'�M�1zxd���7��Ԑ�����/Vi�nL��=��	
t�O�T��.`)8n|�H|��9b|�/케��Y�r!��Zජª�b���୑��(='M��cR��?��zy�בa3F�6I�4Gb9||f��0���5+��_%��Zv%�89�~F�U%e�߶���!���CFN�
���\-KZN��䖯<��3+Sz���\�u�?�����G��^0�E�U��:� ��9�R�����đ�3u���t��H�����x=a��]�7���#2~�-��A�3K��IU��a�7`�J�b���"����h�f�a�b���X���Z4Z�8����]o׌���:!r�xT����peM6�
�nw�l�+�>��V�n���D��`�u�+��4�\�aw6O���@�T���2v��2�g��zg����.Iq#�(������0�m �ʪ16d��ﾛR�n��m�^cyP�ɳJY��5��;J�l&���;�����M!���r�����`�	��f1����P�����!�'�ˑ!����E�DF3���[�(W�ת��͚���o�-:5+�	�[��^���dX��ŇV�kw�SP�H�9��i����Z_d�*��u�z'�����ua���: Z\���"_�_���O�e�ܯc�����[:mq@^�f�u/<VIe.A�T4�P�U�(�e"h����!(�&���/>C%�W�O�7Ԡ��%� �xl���5�ʮ4�H�Ro,��)�A�����S�&���^�����)e11����`g�yi--�����B��G"�-KC?m���M� �Ϯ����0�R0�?���p�+?��1�	O!&������L�,"��B�+�D
�ո?TQ]�Q�R����Ҳ�������, �5��&\ 	��}=�N�Y4(�iΞ���iSTa`n������S��Z�J.*����P���E�����>��<���6�����6���8���]�i�,�4FDb�%����;�X���hgt{�p�@ٲ$�j���&�揎�L���$L��Q���i�^uP�"<���о�ͅ�Xܝ[����e*���t�}K�(�)灜�|lFu,�s(`��>�25�ꥯ���ؽ�d P���t��/(���Sv�c2�k�� ބ�? �E��u㴉�kf5��C�A�Bd�T �����2K�I��+�Q��nh�XM�Ã?��ȾP���k��*����}\} �)Q���~�C#�xI�EZ��[�;�M��d�Z_��zK�ve�)���� d��䱂_�Q�?�\h'��,(�Ye{��f�ⷺl��B=\�;i�0�I�
A|�@��*V�IU��l�[�a)Zo=���@͹�����w�t��׏u���6�e:�ry��2��oq��_��#�=�;����h��H󺽰vEErI��I6���R�^u�`b�Z1�	m��PB|�"V�k��,v�q�ۙ��/у��A���S3�5����4��>?Lka!�'37�E#�W��$r�HMv��� +�Ȃ����&̎����dx��븤Kjq�r��"�"�HU~~>U2�V1�xř�_�U$m�pH���a��ꏠ`�h�F��(�D��4]'P�j �/-j��1�\���V"0�Ӷ-MS� ��M��j��qU��!��jD
`�6�P4M��8p2��QC$��v�vd	�g�J�.ۻ�� P;E�� 5DY.�T3��f]��+i���0�&DL��K/�:C�]��F���GtL@���T��i�m@�jF^9X�0��B%�e�6*x;�I��V@�S��<���.��+㪽�ڧ�j�+L�:h�v�bm�h"xq�YC`>[p�Y��J���iM��W�qM�C4
C�Y�X�6dh�!(X����ӽ}��[�w'�*��O���� ќ�|l���Rx�~�4B�?"�S�y���f$��|I���Om�26e�\��,�b�g�yϏ8���E۷o�� L5�KxƆZ�x�̨���tW��[�Nu��a�>�8��iN(��"=p����M�p���L�u��rFۑ�=Y����"��^��:�Hʀ��,E�J�q��I9��)�+�M���=�f�����`j�q���X����h�J}#]�LW��^�{
�]ɷ�U��\�Ьu�/�pq����YP[|\���9����;*��\E5�R:���lQWj�J�ؘ�U�Cj�|�5�Y6r�,�{i)\�Nփh:֕�\�\堩�py,����U��v=����]��e��_�Z���pDS��1�z �N���	��e��?�������w;�yI6V�8C�-H��� ={�J-W��^�I@O|)�̫�VBEڹ��<:�V���.k-ykv�ӻБ����F���yq ��ȷ��Y�Q|��iK����D���w�� K��Q��;��Є�q&���5[8ÎsT���qJ�M����K���,n�f�����R� I_z��gbTց�f3��廿3� �R`��Yq3~1��JE��a�]���t�LU�^;�6��<��z�)T�
/�¬�u������U094N����:V��_��J�g��=IkraS�o�(%m�S�W΄���l���
9w�$
��5r�6��\��1k�v"NgF�ԉh��)��϶�lA�ԲT����0�4��3� ŋ/:�����|^��$׻^��Y'�/�~}�,�-w$�a\?M��1���l2�V���ڬ�P����G�1�vV~O��]#1���/Ǘ�̿����K���E�r	z�-zCJ�1��B��&���˝?�"Bۘ�܅)r���V�g�x��_���u0U�}������w���i9~g>c��X!48�B�Ff�p�H{ms�a�ʲ��[C�v��'\����>>�����x 'Pv8|�E�	�G�H��4>r��nܖиXΣ��juvت4\��8s7݊!�T�l�j��O���Z�D��ck���.A��O��y%η8iN��Fo�~@A���r��G'�6��{��x�eE��m���y%��J��}��=�|(j����n�]I��SZ�}b��,��]`�&�E?/׊��"����%��P�3M8���w��Ղ��l�{Z�v�E�#�t���y��{��G��N�mShd�{ϗu�ɀr:n���9_�s�W�5ޛF9��� Ąc����g6�6 ��s_�{=M�sͤ,����~2N#��jBk����E�š���������`���n1�z��·ɘ�l�x�RU�p�?Z���2O�>�o�=Mc%�C�d�=T����g�<O��o�C��&�^�{��1"S�)��� �$��B��mڱ�6�3:�6���o �F3I�*A�Q�������C��.$��7DZ}���������܏��ǔ�7�����F7�p'@/��A�o�-]�+�
��/<u,�X�;�H{�Ə8mK�Z��W]p9Q��8_���,���X���VS�^4~�6~�8U!����YrH����W��mz.�BR����-��{F�: ;w������-� x�M1�.B�&�A�x�xg�ӿ *1yZ���С+vL���(KӝM�>l��,-ϴm��oC>��r7G�M/S@��ɚ�
��L��H�i����i}�eL�������x�mԻs��W�W�ZJ�@�D��֝Htw�mF��J/Ȼ[!�.a#�����n�b[����ҳ�.�sR��bM���01LZ��A4�S[�#'�V�O/���
�Q�VN���vA�,�u����̓R��JK�����41yej�t�W�6s��SO�J��-��}��sN�wOCzys �_�m~�n��zD���� ���_����|�Jh��$I�Y��6�
�����р�?�RF��=��<�==�d[Y������ԑ��E����y�f#�Ns�$���9�:%�b��=Ǌ�����!{^g��j��v�"8���?:;�yg��s���C�JE@Oz���ϣ�sE7(#�%��w�&?>udV-#P�{xϼ�R'yD�"�	���X�Od�,5j��8Ol�+Ӟj@���������ZYAgcOB58힍խu��K�J�$�y�%�;o�l��'�;��]O=C��?�K�muq����F>��4��E?v��!F����k�_������p^{H�	m�z����2�E|́KsSfۦt�@�va���W�}�w-�T���'�=}KT���t<�)�0�S5|w�5й���;*1�������'��9���gM����|����+�QX|.&���a��\jm~.e	�����M��������h���[��2�H�q6�%
g˃��`�ȹQNTy��k]Ih��ۨ���V�f����ؑ�#'S�U��9JbTB^�R��#C���gW�?Di��vx
V�Z����	�2t-����j���:��]�҈���ǭ@������-F2�|���-�z�3Ba���?ʵ���h�.wt��@���-x�Hp��`�_����M\*�#9����͖WN�wЖl��ؘQUN6� 3˰'/ho���N-��G�b2�C���&[qoK}�*���"V�f63���85d����`��r"�/�،���A��zMo&3�>w� �c	�����L�ćv�'>
�X�f]0�3�BH�V�nCl�e�e�:�g ���+��Y�>{�5�q����5v�p����=��XB9V��d	�FC��v[ �1쎣^���c�*̻��8����[�}k�S���/�����������&��9���?Uߔf�����1һ���ı�
q;�a������ �e�m�%7�N?u��+8�ٶ�O��g�>��?_H���	ۄ?�F��dT�˻Ze���i��Or���+��T^�i6yj[H2��*�]'�1piz�����*�A
�6�+m�ӉL��5��?x�d|J��9��8�]ܗ�p���#'�^��`ӌ����_�#������2���⹻1�{�*%򄣼Z�0������јZ!m�����m��Kx*Ս�osk�OØӤQ ���D�YG�$��� �G~S��}Ը@�>���'ۃn5���x�g{|$vsLn�dm�i�.�usW?�W������GF \WX ��8Yf
f=��|q`�R!�U�2?Rt4�K�w�~goY��������X{� �_ui�/&�zk��'�T���YFh�*���
�Ҡ\�xv������Ke��������n,�l^�ύ���
�^4fY�ٴd�w,�Y�_�Ӝ������n�2ZG�ˆ�N'ɫB�~�!B+7:$��-��"m��Li�rg�UáJ8�"��`� l�Á)S�7��
͞F��0r�Jb��-�>��.�c��Iv�	�>&�S�F $�Z�e�=���*2�[�O���!�IKl#�����.̬K�%C?ч�b�ɒun^�.�q����.��Q�N��M�2�f��˺���[R�����q�`�G�^51E���Q���ɗ��ĉ <���\ٗ���77]�Hn�>�F�z"��zTiCw�#<Q��G��\��oy:�Ԍ�<����G����r��� t���9�М�q��$��)k��� >g��DNAZA��vgl�*��,�z�Ƈ�+��!c���؇��kM��'��E��m���Y�?���x����kV�9(��3�(�`[>2l�E�G7cm�ۆ+��B��A���%��i�As%|�ZĹv� [��.[d��U	@/μ����pc,ѳ��g�ߞ!���G���+�w���io��ԫ��(��i�8��B� �2�|ܕ=�8)����!F���/S�;���Np�αl�
�_�l_H�?{FG �/l|5�kб�+����،$(�=D������]k�R�9���u��R5��q���6� �Vn4H��[�
���]��:X��s�s�Ǝ�m�y�ܸ&��Y��)}�<�*_a��օP��*_/s�T]6��<�Lg�Q��@X6����
�A
FLg��t����W�zאIކl��l5�E\�vi=.�#�˚Z+�����y1Q�Q�!Z<sE0��jK���@�U��4X;PnѺ �L/Z�S��W���7�}WN���L����I��!���H�~:k�U�5�ܝis=����)~j�+���i*�
d�@I#�6��`��1@XKE�~�<�=/D��D�gQia\T,��h扂�WV%J]E&��M':��~M��7?��^#��Hz�q�O{���MQ�Y��4UnK��`;ٮ�*��ae�w�}t�>�����8q���%!;���#3�����A~�QC�j�Ɵ�
.�m���l��]�т g���]���w�G�SGi΂θ�n�9*	�hN�����͜��t�j	o&�^A����YK�}E��V���j�kD��\6Œ�XĨ�ee+�ܕ q6 � ��_��XQ��x!��̡T΂�1�AD���$���$�8���3IAe���}��UY�h^�2�,�^p~ д7/{P���W�	4�W��Od)<��W����j"{��_�7҈L8�a�E�q,1�WIa���N�G�Kᕶ�#�N˷�1e�r����!c�/�#Nm�hc��t���u�ѳh�H�Sh��rgQ�|bC��B��15�R���?�J�ğ�0�⽐XL�̋�2�>��A��<�� )bA�^��g�.<�&��g��5��9��̉|�0��Wu�c��]������L�9Ti�UW+���.����(�"~I+�~���z�V�{AM_�������E��'LK�po�@�jj�$z�����Koh�����D���n~�qC���_�G���R�f	�Y��U�����<
��j�t�@�����~�&H׻�8bG����z�� �K��>�-�ִ�'���cHS0#�M2�
2(��o`��9ɏ7�TOZ�/�##��d�O��5�R���z�c7�3�ٯD�~��?Ǆw����'~��=-��\��.��1��xY�ó�/Zk�]���H��˥�z+[�AQ�J���o�B���_.Fr��%���$�:-��w�Pz��E%Η'��}ܱI��zN�^�K<>�v���L?�C�{K��R,'!�p�}��p��c�|���9C�@��M��������
����p5��x�0��-~P�Jk2.�pL�>�t��w���7�\�oޱ�r|O\�7kK�L?�s��!��[�y:�ݻ�:ݱ�|�>P���O�|�w�r�)`|�*e��~}�&y�'���� h������:e���,i�|���~#�H��MQUA�VM��t�W��mx_9I&C����}�W����C�=�l��W�7��1{	#�I�a���^!��A�s���
��`�dP4�ΝN����Ы��� ?�y�%��Dϐ&��w��v�az�G(�I�9�W�ψ0��Դ�V�l%����@�=
��!�(����.i�Sf�0Ǆ	�Qa֦>��*I�XP&P�6��Z��4u�M$�/}�$Z�A����Y=�5��I��A������Y 	>;�K���_꺔-��k��gn���rW�B�<�g�!L4:��rYQS��l� ���;vQV����,�C�neP��F�7�|�Ĳ�_�O�PK���dJ�D)S�U5�Y*��0�W�|�;tx�m�1<R����r�	��/����E��j�ƚ�!�{ 9'5X,�ʙ��[�Q�����@�/��P�҇\%o7��0,�D��j��l�԰ئaF_�T8���d�7��|�j}��fψ��ż,�e�+����2����}��1��3P�.��Ki���� Q��<���Woc��%�X����T͏Nl�N����A����e�� =B��3���:�3�����~�%��!jx`�8�1��f��sxx����{��L��ɟ�2��<�`��q�D����Q��ih�c�mP��#x�$:����{S:����U��
��,���Q��,�7�4e�\BY2��p�y,JL��l�nGC6��tZľF�z"o��ge\���[gg��h�~��Om�r�b�K�%^y���>�<~%p��QA��uT��IP�dp-�ami��ӟb�� P�7�F�h�-�%��!^��shПVJ�uY�������钙:�'O͍��Ѓ��C;*�7D�y2.L#C9����4��0��o��>#TTA�/�j� �&fGfb �\��+.4���'�廔�gfC]���k(D�m�Qږ;�T9���{���e/PϤ��g|����t��Yu
����G�g ���#�|�`���n�y)�y��a{�z����y�h:�������ʭ,�6���:��A.l���N�@��f�Y-��~����R��2h>����Y��V��Fj� `#��r^�~���-���l��?7>U+���d4ӂG����:��Tj�����S�FeV�΢�%��IC����T��PH3��r����<���4��J���^�]z��lȾɛy6��T9o7�!#�{�r�Y"JB�2���W����������#1�;ے����5t�7r!��VK[n�:��!�3�,[&&6i����{��V���Ǐ|�p��u�y�aG��s�b ���l�o{��d�_��������r��q�\��\����8C'W2ٟ���Zd�Z�i�e�A�VX4��L��`:��z�yB5ɜ-��D�s�S���Wb��@@�rs�/�h��oFLc�.�z_��N �O:4![9_q�>Tc���O��QN���e=�b�l T>�~3�yf9���o�ݚ��Ԧ1��M"��}��R�������11S�WY�:����*�2#�	�3�_[b�2om�Q1��{1؊�^Guz�ZC|��%̯�q����l1.��u\�����Ҹ���(|���.���s}=>�Sh��e�;H���	�p�Mr�W}
L��q�Ç �@טA|J�X��*�p[�%V��ϐ��~������^�P;�n�T�\�4��o���I��Ӏ���,�sB���r��|VJ�.�]؞���[gιC��,.���x��Įy��u�/0�V]�!r����1��O�=�4��b�4i�
{ZbA?RW F���gz(�	�'L�Zxm��xQ�?��%�]�>\�c��f����Mgp� ��H�O����Фa|�\"9��mX�8@��m.�k=l��p�љw����v؅]{�tGc��à�e�?�.�`L>�з�Jo*���pƬ���N�^�n�ῄ�Y�RL2:���Ԛ�	-��zr��T�����@�7��C�J�Ջ:�R@8�ǩ�[g��Vic��՘���g��6o�|i�I� �&nۤO�L�*������:��H<�G��?'��v��; �"J�]�K��3�y�(?�7�r�8��s�����N���n��֢�ڭWq���!i�*��n �(=*_�p�c Iv}�˲I�����0Tz�/�@�5)4��Xb�m�A��ͼ���Ϗ���
���l~qq�5�؇˶��h@�����^m"�"*��s�{Z����X����ql��Sr���n`�
����#i
7�E���<��n�G3~cQ����-Z���<��S��ϭFdr�L���H=9�<�T�9L�Rz-��} ���K���o3V0��������-�3ōU�(�K7A//���;=��K��2m/��Q�ns\����΋@�?Ey��e@��g!��{�7;�J�d��+�@�M�2�A�A�ύ]	��=���XVST���� hm���A��o}(�ÜO> ,�ο���u���qݩ�� ֵ���
H�X�[���S���-�6'K�;��T�nQF�X��6�3��{�H�(γ;����,ISR�Y��|K��Ӆ�n�|�A��
��� ���C��f��H�Qu:	��6��)s~o�N�s���^���#2��x�X��Ҋm��Rҡ�m@j�:���	 N�|A��?>��Lu�˶����=J�`�{m�ka5X[����A4=�W�-����=
]Da��cr�J]��,��l�-���YQ�y,�A�Z��O�`"@C_��Ecg�Xl��/���f�Kȏ�<�^]��S�ih��%(�ß+�&2<�_��s�$�]c�(��u�-��o��Zn2����Vo_易r�֗u�-(J�T[��0N����⇈�q���˧ƨh�=���_������z��1舜;B,�<pt�#Ư�^���P�,����,��A���(������>�?p��P��\렸P#����1寐��H����C�I��$/"KG��T���X�L���dy$���� Ո�?�U���ZCE焞�~�6^� g1oA��3����� �z(�˻	���Zڞ������7��&5U��ŭWl_a�J��;.��֝�GJlCk��^��aJ��M
+xp��P�w�f�{{�CfI(�?q�v�9��c��UlD���.[��dڥ^͜O�d,�X�3DmL�޷0��]�p�gZ�8�Y�$��m:=6Z�P��dߥ�=����E�"�$l�2x]~��U�cT���(�w^� �w<��cOŇ��'�I�,9�
&�Lu�x����BY����b����GY9�7e�K��}yE�6m��ME!&F�k7������.��	9VX&������NP5�$����C�5JR��ǅ���rZY��A��}� �U+���{E�wr� �g���/�/"��k:T$���*��
5A�Ț�޴h���ӿ�9�f��鶱Jl4�9,z���1�@��F�����?!�N_����qm�n�6�����Ge.y����]-�0��"�*'U���c(29�@ o[��p�,j���17e��Jx����isgyW��X��k@pFJ��6�AM�lw3�	^�~DZ��t�;��)��6���X:�c;�/��I�!?�=�@:%���~��̏�ʃl ����2�B��;�<�$�������~ùQ����כ5'��b�K`�Ca%(������j
�$�*G�D��1sS����v��/d&�`V���4�軄y�;^��U�4T�[�Sn~	j1���F�#�r�!�s�<J�� A�?�NCn�݃1��& ��C����(�-��䃙O���c�7Q��l�Z����{\�E ���p��/\^���fZ�.�� ¹V����N��j����7�t�\G�����G��z�p���1����!r/��~�K����^��)-�g)Y͛k����=�K%�&|:��(�<��z�_����8��;���kb�#�+���i�۸�KS�W�������{��f�䒁�!�.� �&�U����t��3Pn�z%��77l���i ��ժ�:d.Yv�*v,\O�G��F�i�JP�^1q�.��bc �1l�W��pr�~�i�%���]����QQ�!��Q�=A��>*��c��Z�¾�k�ń��!���)Z{�zY�D1
�o�n!A���C�@��	������ڸw��5�-;�~j�L߂o.��L�v-Q8�olG�1��2Xh��$�'�?�F�>��)��.#f�g���o\�M%\��D����d���&ȧ�G���>�\��F���f@���Do����5����Zt�E-I��+fR�AE)efM����d�P��:>=Q��#*+q"���t2-�)��f�?sg!���'K�ri�	}_�X7�Z[J�pj�h
73d�wlm��t�ޜf��s?��wD	1X���N�4���F��(ڻ!ͻ��I��A�v.��)�E�1���~/��NH�8���p �vI�Z��-ꛫEU3i�LMv��YoVQܰߐmeV�d�_��j}urP����p-4P� ���^/|j�$pF,���:����T?/��7G<@�?T��V���9=iT�.��-*�X�j�,�8�25v�]y��"�9��g1���Y5i����@%}ҁͷv� �"7sʲ�(�%�io*��v�6�8hL�6��v+p�Ɋ�2�� �Q|t��횮���c�LSe�)�3уl�2Aeʎ�l;zT�	Bu��"?+�*T������SO�$��v���\F)v�h"5�-ٌΓ�싔�m���ύ�VB<*�a���gz�P��@��'Ը�����i*��rש&��>�JAo���5��b���)��moQ1�oLP��,%4B���t��-�d˪�l��m3��t��$��D]��:B0�@.ۂ;cŮ��5�>Ne�ͭ��a�̘�im�9���Si�Wp����j�>�C�GR�7�*u9��)/f0�m��� ��k@�㨤[ʐ��z2H2J7b��C�
�V���rVE	^]m���cv3�߬hD!���7̉sO]4�j��9���B�3�����d��(h�!l�Wk0#�J�����������-�"������1	�}�v'��~z�u$fs����8�Q��a��ܳu�l����1ے���ee�D�@xv)U,|f���h���q�N�+�����T�6�.vhq(̰�����m���k���7]L�PK݌M�U}2���;���~!���x�`1yp�1��
,�|-�X_z7#{b#�i}W]���nV��e�M�cb�1��U])p49y�%ǳV� 3��Gs?t�v���#ҭ"8�IT��O���=�3�Z�4�:�J<�V��$Q�<��.!����D�d���e�ntiknO�k�����g�D��� ��NU��/
jر�d1�@/�A�f�;�0a����B�yN�����v�q���cw�e�%F���WϖƋ@�����5�XY��]�F
σ^\l��N֯{}�|ˊ����\�C��$�U�v��R�gm�4�4� �R���AI�ǥ��j�hm:y�q%��ȃ�Qm�_����N
@�*�׭�3}�O2�v��)z�� 'fRZ���!���Q��P���?^�Ru��F�Z��ޥ����F��;"L�1�!��wb�%��/T8�a���=�1�����������I�M�o1R7�v=�~�j���	I��t��\��u�S;���|�ɍ��.�w�a�����������p����a���M7P~-+jj��2]�ҭ�}d�C��.6�]Vw}s����=�6��ދ��\���,��m������ ���<�ك�5oP$���z2�b���5�&|����R��0���i�RֳD7�I�c]�n�xѻ6��!!�{x��{gX���Y�(�mUr�
�긭
m"������v6��C��`�����u��u�#G�����{K60(JAN��z+"�Q�=������e~��d�N!�Z�&$+1�K���R� ���LM�L�g{g�v(��E[��S��6@���g]!n�rD��'�%D;����+W��=/^a�>���֩���y���O>��{��0������alm6!y��$���Y@��%������Q{��\��.��>>�{�h'�+���䰇�r�]|�qW��J%^��M����S�CKGe������˝�R��nMx�*g6J������h�da��6~0��k(���y+E���u�4��)�<'|�GH-�t���w�c�r�%���7.:[�}��k�E]VW����h�`��ʔ����x�����Y>����ۍ��J������J=#���`�9i�c��Ap��z׉��U9ӇV�oBH�S���\��`�OE���I�~���sr�^k���؍��޿F�EȰw�@�l$�tD��cu�1�Y�e+4�	uB�\ĵ�Z^Я���X!���ꑓ��o�/��#^�ɸ<�3�i��h���ۧvS0��~�f������x$���-�t�V�c#�j������G���}Ѝ$�'� :(�,+�X̔��A�˹���"������d�.�fj���Xm���Go����'j��-��X�@�W�:��:�d�N���y,�ϕA�p~#M�	����j��-�AV�Z_n:�i'��1�`�"i���.�O���X'�X���x��ԭa��;�z���d�*_�!%{h|�?�!C	MR#$����pPX��G�h��F�7��*���d�= ȗف�m�V�:ߡqd�F���0
�@E��uN�ݮL��T�ws��3��Lg�S�g$
���z����G �$��E�e)���[(�Κ�ԺM%I���������Rpi*�u9���n�t�D";Lݓ0kl�Ғ��>&n��#�� �'�Λ���	��l��R���J���A����V#+x�Vl��cN��Ǵ-J�L0r�ẋV]H���1��8Q�uLԨi3MNA�F�NGC�[������`v�a��hJ�D��0����B����1bu���k%F0�J�ku:)*�N.&u�k�<�k!�i} �\ɰH��L���M"?���ac+Sge���a��KB�f��A�`u���:���L,��#r�a�,R(d���4n��/f�)f(d��b/	i~l�ipv��"�LjB�O:�v[LZ�m�-�B��\gC��<�4�Y�o�3 Y�������ך��l7VtNj�u���Sy#T�Yj�=��%���Zj��+�lJ�Y:lC�ZZ�T5�>"\����Ϯ!8������� 9N������526��4������9�.��0���<T�����I].������3�~�"{'����kn��n�Tu���Z������PM�b�-zZ���O-�Pk����k����"�Fа��	:�h��q�lt�P��/������pl�-ɋ�����?��,�/�+��o�E��1�O�88Wq*��Eq���2���6Ԓ5���B��)�3���������\ �������=��)�@����g��z�������_<��`���鴡�*�������Ӈ����.$��W�pU��=O������1��I�L�es �M�~���T��%auѿ'�DmXc�p��sos@^�="
�¼X�,�g0�����%Bjx��]�p�)�.��	����CLf�OA{)����*i���[&��gyP9�v�jIUب�{^i�@����Z�Pry��Vs������J�z�\�G���`��Ȼ=���i⁾!l�r���d^)�]X����z��R߸��&�� ` �T%/)Ӷ�nFtT��[�y����7��,�0S�f ��l�4?*���Gf�Be�`�J<����>h�V~�{7z犨� r�+GΌÉ��|�}���qD<�����lּnZb[tD�1�{SA.��1��բK�h�Q@�/��ZN	� ��N�\Y���V�|�%��~T��8o�̞�R���}r("� m
�lG��B���.v����,g��[��cgǂ��1N�4��K2V�ϩ㢃�I��g�-���E���A���u��7y1�+�\ɩ�P*OF��T]}��C���Z�
����"8w��n�bTl�LKe�Z1�Tn�KY�=�2�vsNj�ݒ��9/m�mՠ$ܐwF�_M��t%��"�t,��uH���&R�W�tZ�.�����K�E�`!��8���z!�b��ƥ�Ξ6�߬��m�oʘ���S�Z��?�K��:��5甊�D9d1h�W_Q`⽤]�D�q��;rG=
�?
�Q�3~���&��D>@\�Ҕm�\���0�΋De�_ң�S��Qç�������P
[t︻@���ռ���Et����1.�I�5����9��a5:��Po�L�J9iۣ�)ë�ɇ�f����*�-$�"M�ޯ�^�Aa�>�ǾQd�O��%��֤����J���6NB�A�r��g�\F$�)��|A0 �B`wrd���E�g�.��ːy��y�u܂m�!����U��rA.�������N���(q%�uR^��l�jڣ�k�l�8����\AC���̒����L{�8��h�	�C&.�=��"�d
�$Z�J�J�C����E��:=���_�ch�:��|>�U��w�i��%5F�g�X�+H�.Vu��ɖ����u��Jr���H�J8�޶B���+���f���Ό�ط�,7%���&B��Hӭ����PAw@�^A)`�b�&��ˊ���;��i�,ٶ���ꌾ�y�����N,<P��t��@�����e�\J���D��UR�����&Q��h|�d(R>����(����~������>���B�%��r��c�B����麊�֩�𡫊R܀@����gk�'yI����HB�2��i3d�P� ,���)\���!=���L�O[�j�OE �� L�CV0o�6�{
��[[!e
��<�8�%@�i��E�q+��>Ģ5�}6�Ur\��$�U�t:O.ܞ͏�{E����L�c�֩���tԉ���l���s�9�]�+a\'��ӳ��W�~:MZF�ڍ	�6ҥa��<y�1��^Hy�.�@�V�?gC�4^z��){�CЙ��On6�v��ؘ�2Pr�J'ºE8�
�x��v�v�8Ix��|)�k�׋<���'d��8��#��F~��P^,��sv�tմ؊�7�u���e��+�_@T�Azo�r���:A{�hf�M���a��2KȘ%��)�ʓ�MV�U����|TPb5BHp�x�T"p�oAE�_kغ�R�J�2F��\C��Z����=��b��D�9{��rIӂ�����l���/��2X���!Gr�g� �G���٧�
�L,�v��o�T����L���פ\cU��޽�S2�=P�E5���f���73��wˢcXƞ�uo���KB�i1�i����,'�Yr�/}C�U����f]�l`bIa�}�����spfaN(��L⿸1�fJ#��e����m��.-�U�x�1h�q�?�g�^��^2�g��bN��3؈f�Bgp�9{]ܭ05���U-��)}��Ԅ-�ͤ]Rҟ��-X�D8z{X�l��#��	�y�n?�RcJ���p(���]qO~�b�f7�\$V�x#?&}*����R/�5n$��#��E��mZ�1MဓWa��������~H)ԨJ� @+D�)�l%��Q�p�x����?�&�f��ɒ�D�8���y�)q����kO][� d�g��VϬ|Y���?�ݤí��(D���ݾ$ �z�<��EJl^����+x</ޫ�J/^�ށ�~�sd�ޱg��egtp��pP�������qLV�4{��쫁�n[r��7�S�M����S�*y�@^�	�.�[3t�D���qȠ3�4����p3����|�<��ԃɵ)*�A�����,��|)��}*��o@��y0�wQ���/^�Wr��JD��W /󓂭R�r�*�nF|S�V P�%ʋXfw��>�S��$U���% ����M��vl�b{$�Ν����Yω��[KK�d�o��q$#e�Y�Qn��8�"9tXp�K�#�$X��˟�?"�X�v���T47o�>��`3��l ���+�~�ҡ@�����!�{��=گt��ｓ�����<�EPD�� �����ݮc97t�Cbh7�y�l�y��j�[L���a�,�o+�7�*�7o�T��g� ��r�d�?�X{m&�=��е�ج����t�7�z�.}�2�7�Ҫ�:�n��&�JW�/7�(�s��Y��T̨��]o��~S2o+�����J�z,>r�^j<�?��g�{ �k"�Q�4�x?� �#�^Q���#Ȩ�����`d�����K*-�8�a@y�UA�q�WY�ۡ�tmF-(��=\�g�,�����F�Rr��@Y.�e1z'}���^�r�1���]el����w�#Yh�e��h%w�����ې�?�W;��ō4�i�n����y�,a<R��3Q3�OX��v]��h�n�_��MT� ܈��a?+�T������S�.�V�WY(g� ��i]8���W��)��4w_��A2f ._�e�S�R �U~��M������W�'A?[(�q�>*0/�Ҙ���+�8I�؃>%Ȩ��_$��^QK#�����[>$a �o�Vdb��83�n��^����hdG8yn�=�j��Y<._�xlG����?����$��m_�1�Ջ�ܒ��)O���O{�S_=c�0a��)$n�y >kԏl�f�TC=�s��6��jT��o�i�����ѹ��8���&�M�2ϡjԎI�d7�b�>�v�P�7��/��@�ܡ ���矴]�s
gK$�H������ZE�e?�2'l�HeZ�Q����,�[�t�%tW`���"��=��0����:��B�Yi��sI���rS$.��e#��G	���c;�y2D�A�ŲZ̩�y��̉�E�ҰD\�hT�P.hp�����~��87 �]��7�����Sf;�q�9��-�W�#[6��^Ϊ�9m(����K��w�/E��[��=K5]DwWG=;À9�Ea8�&a��w�� ���-iޭ�.��k̰҄�r}� ky90�+朾<4�畐���57�	&I�D�u�[C<f�%��o���^B���b������q���eo�G!�D2����~7��ž������uQ�[�`N5�1@��:�{���=�KS�XW�9}�uݨE�B��ƍj��M�`�鏪Y\lE��۳�_�����0	<���i�WRvtۤ_��2�Ef��{ǎ_Q��Ɖk"�6��۔���/0��vY��z�A$�|�W�״���,:x2�Ii��wEGM>�|��SC��yM�����d��
�j=�CLVRMx�¬^�y\��
�H���q�g���l#M�ź�h",�I�ɂ���L)�K(7�@JdPsĂ�j�[v�+1�����v)0slBA����J��J�����! �A8{�O�(�+�e�т,8�)�h.>?��eM/TN�o�0�(dsֱ�X	c��[Q��Π�\�ML���/�1���M��+J�6~�J�rh;�p/B<v4w+��@ƈS8�����7@�n��Q����;��E���l$F-y��]�^"Ɍ��Z�?�:��Gs%����"VV{���*ɗ�����q�l�����/WK�k�o(�]H���L�kי������_���6KT^����Qx���/(;h���5N���`'c#�"}�!�#��ܫ}-)�,�[`өLR}���_�1"�楶��É�,;��$�#��~6��A���V�)e-x9�q@�D�RG�I�lȭ}O�R��yl��Ĕ�!���=�6#�r 2��Ch>}�a)�m��_�:��ѝ�+��>�&����0\>뭛h��
�o���d(`W���\��Ck:��}�=E�4��i0y7�2�o�m��5�RF���L�x��gu����ѝ����G%LoZ.)���+ ��rLo��nK�c�H��ND�Q:���v"�)����R{|?Mނ��l��n�Oimt%`��U��N�#d'��?��20od
jj�]k����I�~����}\K�,�J�N�7s������tgB�H5[#�Vf
���"nP��l���*��jhT�6MY�Etp?�>z��p���(���*J���v�'�.�]5��g3�G�vdU\a�*tI!��H�nP�O�2���'m��1{���H�7"���F�����!o���픔c,v���d��_��e�\�%q�i!6��11
�*������Ps�#�rM��k�#�ߜ�����M�����G�Q}4�q=�+���a6�2�f
vv���W�j�{�K���ߔǷ;);.���2���}crBkSʒ���Z�siE���}�t:�dU��܉ux�����K�=M2���a���.�]�������&��w�5^�����5�!����~���v�toGZ��/Xּze-Z�2���8�pZm��]_�B�ܔ|��/z�蓒W7�q�`�7�%�ho��If�&�@gX�6��D��%oyV"s�9�xK(������&m��!���p4Y��2m���i&1��(\�9�.;�5kd�>CIV�naݗ� Q�0���9}%E�4�&�ݮ�
I��Q��L�
Β�N^[/���Cx�]^F�ۮS�I�*�!z�G��!���!>_�W��g����mw�J%��4�z ���P��g��*���b[���B��j0��_u� 3l����%��!��b���^t��}����<��Q��
v��i^^]�Ei���X��v�a�{W؃�U�i���[�A�R,)j�$.��!$\h�e����l����Ʊ��@�>�bC_�Xr��.4�l�Ȟ�M*>Zѹ���A�"��tv�P���, �F�`���GG,5d��n���u�:�h�����{��ʘ3A�X4Ė3��H���@k�����7]�ESm��s5��Q� ��#0����r��j-=N�d5ϛ�L�78�����\R�sGP<�jnR�~�������M��,����ٝq�\:As��w~d�C+�g)2�ml�}$ӆ��I�]#�'��
9l�qY�L
7��V n���Uz1G�5[�j���L�S@\������P�3�_���Ԑ��}0�6���&	�)R�,#v#�P,(9YO~�����̬	o�LrD8+K����C(T��<[�kٮ�i	u�Be]��u�j�.C���>D���E�fE�Fq ��"��M"������rB������Y�m,B�H�����I�Nט�j�e[��G��Zb+�b�0���Sտ�7��,��A�0+ �5�IB�)�(w��}ym_�����B^��j�N��u���P=
�n�	+^�����5��·���"-��6^��.ؾ������Y��� H�2c��=���t:
"6U�C��j.o�#h�����!䠚�h�I�  ��l)kNq1���������1N)�;����q	`��"ox7���ޔF�!H=;�nLO��T�:l|Õ�J|&��.�\��Kf㛎�ɟ�Ů��� �:a�!X�0"��R�!�XҸs����m��ܠ����ЭI��c��>)�Ux���.PC��9�=Tg�7ыu�/ ҭ��c�[?[��*�CS�xo���y�p�?�]�A��m����$Y(Z�M��U~���a/����~���e�c�ވ�n������8)
�82wM���ԡ�}(�ԏ,*�r��o-!to<p��:�fu;;�T��@e�ݥ�������G�t��24j�E��ױ�$�Q<-��o(,[fq)�W[�(�x����񼻘�EVY��x��Q!�S�T��g&�P�4�I����ʽ���\���G�Ն8��ep�IREa;f�3+J��HW��@Y�v�Q}�o�e)���4�ìJ���D�'a4�Z���X�3Sqm�6sٻ�@�D�c�c$�!�1&$����<�=��j���� N#����y;I�r�cJ7R����h�r��㚍�M���5�O��`�,��@̨��Z��ȗ+:�,���z�B"��&~sA���K}��2��8D��L��8}��V����a�j��������`�����ٺ�|�Ni�`�Ay���NB.�qYԾ��>Et��+$�R��w�sO�k�J%��Nܔk�Mc��1�9d@Ar^ Zv' 2N��D�w�G�f�ҽ����rn�"ZH�;�N���i>a�Z�]�̄�V(U%�����~ �ܣ���$.�ub?����{��UrLX~Y?�ʬ
bMa^���#�d� ug�ׇ�nʀ��m�l��5g�x8q[�B'Gy}�ث�ڏc���F��S8���o�E�񝍐S������	��WMif��{����b��ܖ�䁍�;UA��?K3�x����Q�IF�}}�HM4OSǊ��+��&�ww$���f�U�tW��3�捞-P[w�R$|�v�a���9�|�S�v< IQ	qZr�eʛ�	��X�����,�����ڠ�0,/�V�u"W���.����;�l�̨K��)S�5�a����%4�Z(��R�G�pQ�/�
��� G�9���P�c7(y�����@�H�[mU�$�!�)ح�u�=��v�v��/�/���н�>9ͶcB�AN�-�V0��3�lÅ�����YI�������'f�Lt�W�!�!�g�-�Ǵ��Kif�����Ʌ� U΅Ĉ�̻k �9���@�a�g�oz�H�Gc	�A�K����#m�[�Mm��d����F`�=?K�`�`���W苃����-���.����|~f��[ 3�w#�t��&a������t�}�wp��4B�Ԡ��q���K:4��MY�S�Ah�a�^�YR3�k&��bD�2>[9��,�[�Bo��#0*��G�����Q���o���-2&�Ⱥ�J3&�M�H=g�SUx�V��B��V/�v�q��D
�-nU(&P�r��%�[i���Zwq�� p7W�"o��	�K���fϹ�G�r�a�BGhЀ��^�ٿ��x�Sx6u�:.C�W�'r�-�����=U~=gk��X���1������^����i�<S���1��9$J�e�!Ϋ�� ������1͸�-�"5����������k&��W�g��g��R���}l�匥oN����4�ݭ,O�t������v�q	w'|���fޤX<c�0
�6-�Q���3:\ĩ0R��Q"!jc!i�����@ /�yS0������Kǋ��Y)�Ȑ�.�h/Y��>ÎNC_& 	1��2Am\���l��[�/���ϟM�e���t�I�͍pt����U�eK�DEE����˰�,O�������!�E��?�:��d$�R��.���� �֮�MT�Ż��<�-h��(Pr#d�?ւ��ʯ�FKTD�lE�e|�����h�Q�m(�
���q������mS��6��{G%�qb��[LW461iCz;�����XT?����{�-;�D��7
��r��$���6�שe���j�4�����+P/Q��"��/_�&����f��#�B��"���|J��\_޴�t�VA�r��ЂY���V�`�z&��B���+�����1z��C���a%ʫ��Qy5�v����1����x��[0??+�=ǵpY���7hس�g�h/9)Nn���+ ;��W���8p�����/�;-${-���h���ɳ�+��$�~e���Z��Pm!��,��̋InFn2�o��w
�$^L�lF7���L}�껨��i���Љ._T�(W�L$��@W�С��dݶ?��h�ٞo&�Bh	2E��Ig�[ �L��=+<��ȋ|���Y�	ǚʔBJ�gstH	��O��\xǃ#L���y�~��t$����H�A"��>��ie9NB��^��$ʚ#c�qN`�b@Y������ko� c�8*��m��ĥk"�bc���k�iBt�WRu_i��0B�C�}�ŭ޲�i��Z���+I�����l��Y`>?���.��d���X~X��Wo�};&_��{��<�8�
('�|1:�q�`A�V�v��"�@��ҷkć� ��̎�%�5f!�G@�Ǝkl�*��`��F'#Jl���*���?rMO���B9��-#�Bd�/^�O!�K���@�':��l���Q�;<&�6���:�	��nw�,�Qnh�ϧ�f�	���_ceazT#�xo1WW83a�;���k����_�)
�~��0�!O�R	�Z��8�{�ۯ��E�a8�Y嘣q�Pja:���\�6���z`&<��-7�tF�4�`�,���d�E�ˬ�D̆VPd��"d�M5om�Г�Gfxd@�HF�HI�z	��Ϗ���\P/x���(�N����Y�Ab �F,�R�$�i�˶�.��8�\���7�)֛��ڲ��è�xWZe���-�b�A�!D��!O,�M�e(��E?\�����%�k�Zn�'F3�bp��;���OӴ�[����؟��q�c@��G�#,=i�L�N��s�K~&��?P�/ǫ���Z �uĲv��t·�H_7��3�({l�z���Y���=HWٶ#f4k�L7�4P˳e�6���z��zW�>�H���0=e�S4i�dh�m�/��\ϳ�p��Da>���+�MG�{ٝ�1���r�	�E��Z�z]�˵�׋�A�v������m)n 6��$�n�g�r�Wn} �Q1+#�8=���/@�X��A��>��u��y�*w��t��#N|�	-�)짃-������tjv��&FKh��|Y �p`2z��$�d���T��X��:������3j-ܨ�ݳ����*w"V;8G@��_���)G6�� b� 6�JDߛ�p���u�)��\��Jp\Bn��q�4�EM��zm�۳W�P&a����d�y���C�r/�Y�Y`o4�c�
�o�,B��V��I6��o�)�i����]�s���L�����%��f9[���<5�k�v��Bz�?#`����cw09{_28|SxI�rF�#jHU��5�VV�;���u�9��I�3���DcP�~�
���+{�`�U�l���X6{�-�$;M
��T����c��gM1W鹦�u�j�+��5th�5�7�q��rMRm�����~He��[�@*9��������b��^ۏ7K�esǹa�p9�IZ9�4k4�#��lGʝ~0�B����\~S��"���pꊍGWa)�r�_C�WJp@%b*�<)�(�����Սa��l�Xot�rA�,�8�sUJ�ˣ�0fe�2�I:Fb�xaM->5�q
&�\�"x��P�"J�ڗmW�wX	Yɇ�BOs�*��p�	g�<� ���f4܏��.x�>���Gؾ���^�>�d�&���väl�5=��aKE�'�;Ҳ.UWL}aRMZ��C5���~w�|JS�����R�N!}j;��F�(5l Aj�߿r����)'|���EM�,f���̈����@�P������K�X�^Ԕ~_��U-������N70x*� +�I�#�&�����F\O����s�M�ۡg���k����c��3�H�e�9	I��	�tyÇ;d6��Xn��cBt9��D0-����'U�Vyd1d���3��&�)v���z4��\EX���xh?�<�8�k{�/�h�*�Z�c$��xPN`��WzИ����]�G�ӿ�qQ���DU�L�]�K�,I9�g��Zr��U�F���eE���p9���67,��-�p���?�����p��
0���ӑ���H
��w7'̓�Wʱ//k�n�o�<�� �S9���6/Y<�w����s�#���e(Bt�?b�-�1g�KJ�X%A!9��"�٩��M�{��$��ޠ\���o�¹������I)��� �9�,�`�%פ:���^P�r�UW��!d~��͑��ѱ�Dp=U��32�SZ��o�iad׹M�0�/���I��yB^������bM�%#�2�����ۚO��Ff� �ye��|,�Q�V6��?�d,�8��'Ϻ�f �)#��n��Ț���!� ��&ʤ��ɣO�=�Yp@�`�~|���}.��PE�ㆧ�.�nR��xnNxK�5�u|3�'�Ɩք��^�	}����t�43<��є���t(���F���@+ݾ�X�[�@@�x��}�/o�|��έ����������
��Ȯ�wݼk>�4�����]��C�k(v�ڥ]�H���ö0�&o��\1��ۮ����l&\)[,/yĻC�g�/#����}��w.��򶝜��s��8_�(n�=�� �dJ5�8�>O�u:�<�W��ba���_��o���v�j�<m��
�n�SM�D��Њ���Y���DY���=�ߦ6����h9ʳ��Cȝ���1DS0
����CSS�0�q�E3{)��A	Ir��� �	,��T�h��wM]�[��<�������
B-��dl9�����-�ϵ��p�&����"��pm�t���V0	�\��D�Ku�� ��c����9�B�4��v����� ����D��z�I��y\ͳFd��_�-F_�LU� ?���VS�f�v]Ua���W�\g�j6N����;b���4q��$�pǟ��%�"�(k�W1Z�`� F�~�5�^�W�}<-�|L�����)i6t�|țg����$�G�7>��J�D��\\# k��]W6���/���x�_�CS(�q��;."��n���bx��50�ML~ځ2p�ܣ��x4���`��P��4�U��hH�d���{Q�?y�pvl��rf�Y�h;�ە��2U���Q`�-f!�.R�+���-de���f�¤�G�P�'��l��T��N-#{�ޛ�}��S�[��T1<�YO�7a�&QB�G���7��r�c��?a�*�
���X�W���Rv;����b�oaĢ.��Q�) � @?DY�C��y��Ž�?��x�ҋG�/�֏��3M@���p����`6:�[�sh��L�2����}l�)��������5��->���P�]�"�}/�uwo}J�Ѩ_����%����ז�oܔo��'��n8� /$G��͒��� FS�MR$w䬠.s�T�Vv��n(eI%
�� �}�;����2���R�qg\�"�����U�!�d��QB�Nw�8��݊D�ٰbJ�\{g.t(ˤ#�,[sՊ���~��x����q�&�	��֩4\�ըW`���_:�AM�jە1z��������(�-b4ԉɨ�Yf�8�X2�ZJFO7�}Ky�w+���J1ص��ΡP/�R�^��+�t�H����^a���p�&RDǐu��S�O?��{Z��:}�
��C���՝����JH��#�\��%��Sp���M�s�GU@�^
a�ls����B3�a�@A���s>��!B�5�n��aX�l��`L,�om�~��}/��������6�He���\���vȖFdF�?��L|PfɊ�1�����d��b�Q�NQ[��s�M�<_�� �e��7_k)��d�����1�~��f����pd�~/\p�ǭ��,dJ��Z��uj&(��ט@P�T�}��e@��C"c�.��/���HDɱ�S=�<g��Ȝ�HR�&�Ϙ��q��^R��wAh�|`VB��8�M��o�S���ж���L��o��PI�h��M&��J--9���]�Ĩ@�H�*�ߕ��B_,1�x�B�Wl�n��-G��1G�!I�_�yS!���cmYq��0 �2�r�ߵ'����$���Q�]Аoi��bӡxf'6Rg�NǮ�Ϩ�	R(��>dz�63�>�sQ�W��h4��qp��T�l�L������>���M��h��N��0����+jŪ����m�B���C�>ޕ��ƍ�"/���K�bP�8_5H=�����s���6��b��|�?!�>�{�^�be�e[�T�&{d�#�[��̠���T�b�N��3TT�b0~�WJ�y�z�Z?���Y�̓��˙|��`ge`N]����\(+�oa�����c;�s���!?�?��0�*f���w�*��B�ǒ���s��L�w9��GbW�ܠ��h�}�����#��vK�M&�fpن�kG�	W�,�$�ۖ'����
�4�\���t{�"�Y&LT���=��"T�.��
�������͔��M�T��f��"Г��<����د����W�=�!�HaD�_Ua~?Kq���!�>���-���J�/���������Q����.�eG/+�tڐO���^�24E0�����]L�������O<��ޮ4$���^�S8�B|\X���]�c���c!k��ʓ>��r�0�ړ��Z�r���e��2��/S����	�Cn�J��ǥpo�G�x�BE����'�q5��B[e9�zNR)3-�͈|��>u�����[oh�"P����ȏ�c�Q�*�ː�ۧ�{G�b�����í�N�y�bp0�CL�j	[��Z57�kK��®�=#��œ� �$�a�H۵�4E��>{h��Im�C_f1y��,\i[���@҆ߛfU���}���B�X��M��<���������1
�d��� W�����M؂L����ă�e�>�)��˚kz�r�4Y���LY�},�Ō ��0����x0�S�mX�Ά²Q�y�ٴ�
�Y,����'H��D�+ͅ�q�Tv�nD�����v#��q��<b����wȃQύD��,'�@�0�gQ���xוUj�����-��r���'r��}A(�vA�=�؊���c���IH7��B7�I���%���P%юv&l�A��	���;�ﳇ[y��N�}_��o��w�'��S�|��~g�c�p��;D�)�_f�s���(:�C9����òi+�H�.�B�5���]��YO���m���p���&x@�q�E����%��I���ft��O��ɓ�o.i[
�#�_2�,��)"�V6�J更�#���	x�u��e�ͨ����m�t𱏍l��s��Ot3�����V��K���G�X�4��3q�y:~����:������8�B]}��]�U���ri�Q�\��ݽ��G��e��k�%)�'T����PĮ\u؂]�F{���	����?���r�gZ'D����3�O-�}���jNR�1��g\r��Rh��\�(8��_:5:�� ������QA�)�bqu���J��s��k(�G�T��������6��WX�G�Z�I�z9�g������_0�YO�Uc�D}���	��y"g�����=��i��W��'����z/�0wN�t�S�5��6�6�4�g�D���Mu�E9���M{��bJ~��=J��Y����F���UJ�8��F�%��}@��,�� j�|AL�FZ��R�&uZ&�.9ҫE���S6������pq���=q2�e����>���I��;�FNT���L��U���Α���ݍ!k�1�HG�����X6`1�rO/	"`L�c6&i��)�T��.�Z&�z�-�U��u�����%

��%��Bǌ1I~!w�wu�==�J���7�gޭ�7��լX��	ض 8�Y,�s�z�ݒ�7�����p�sWT?e��q�����OO�/��A�Ӎ\h#h=w<������n���w�r��M�Z~�����%�ϯ�����c	)�N o��S	W�DѨ%v#�c�C�Ū"�CЗ��8̧n�Ƒ����p�	����H�)��{��sZv�ω>�iWm�H��A~Е��-�m��V_M��ڝ@��|ڴ^�Τ6�k��2���T���I���s�Tm��ap�����$C�ܱ�%`)��	O	ϰ� � q����s�E.�H�g�v�:.	S&
Om�ml��@:.����;@��H�ɣ|bB{���-qy���g���z��p�A2W�GUC����ye�.{f8�>�8d���%	1��p��s]��.�WsT�/�ľ 9��-�jv�A-	��)2��V�?�,����vB������25�Ʉ*%c�f�V�?q4ʙ `*�ߩ�e5�iƕW�̈3�辸n�!�	"搱U?x��GC1j��9��µ���[@G�/�F40݂7uj{��㖙M��'������a�\׺��nf��O�z�7��Q�fp�dQ�0.�N���f��F�$'H��U����4"T�v�yڢ6�F逦�����7��R���C��n�q=b�90%(�K���
��6{�<�@��gGX�b�#�_��SR�Vdi�}A'�)CO)jrC��F���}�^�P���|�Y#�㮴	�8Tʂ̞C	ٳ�9b���`�B8����=I�)���m��u`�{8IAE�������䪁�[9Dْ,�(>�+�)�1�(�>A��*��?y���(�&�9}�>��U��J,>��8�^��(�q+��>?���d���������UxV'��T?L]��S���=���-{ɟ'��2(�`vn�>��n%U����P�:�D�`b�ۂ�M
|ͦצ�/�^/��X�
_��Q6Ik`u
_a|y��j'��'&��ؓ���ގw���5�Ƀo�Ģ.5��
1ЧTE������n�s�Y�ۈR� �����iC�O�8��/��S�ʭ��Q��Fp��S�{�!���o�[����5;�-���f		 ������"�%H��O�"I�l�&Sk��zHY/w�E0>T�az�倩�oֻ2�IZ�QR,H��
h���*w�-�����S[��H�.���SM�>db�G�`����_偆�E���l��R���	�{V��i�x�p��8��?�)[�]�ѷ5��)f\�����+�-���G��R9�����܊�J12U��=�%��C�{�n!n��ɇɯi��W>������)X�+X*Y��/Z3��d0(!���ʮF e��=tw����f����fFQ_+#��ƶ|�
{S� ��ȅ��!�T�-4�����j� �W���F^����c_�D`[��0�G`ށD���gm+�bVt���p��5�*�3xO�����ف&K $N,�9��8�,���������D0�9�hX5�_�c?|���%kp�C �U	�4��i�dt�D�H�J�ٯ¤���k��@�������hX8��n��S��+�*�yĺx��ӒYĐi�L	R�7��˼5��q����<�CR������9�e�܀@��MCd�^x���)n�DR쐪�Y=��9(��0��Zr�G'�d���R�N�~*X?]�:�[�Y��!�/�)�w#�18�r�ϊ(<�!^����T��1e?�eͩ�G�7,*Ϋ�&� �`ƸRi~����}���y��&qT������p=([�z��ɕeDR�s1G"��e;#�������ԫ��%�H?p�g�5v�ȥ�B(6��a5�Lˠ��!��?���D�(���PN[��O��T�b*Ì"UyD��=��0�Ύy�eo��kZ����������y�����|u���#�8���VQ�B
���L/sF��9߲�9C��f-T�罀�m�F;O8�#B�u��C�9#p�����j�7�2��^j���p�Q._��FD�v��T@�)���
��wg3�<�K�m�{j΢� �*FA�U��<�y3�Pi��?R[�{���2l���n~S����#�cz�%��M���KF|�%���I>n���bZ���m쾅���q��Sv{M�+%N;m�̝��G���m����6�ƺg˾d^FR�N��{�晴�	�mm<��548r$/b6~�ӷE;���"{�t��p:<�&q�=d&m��������CCn���f�&���&��	/&C��܏�Fqi�����q��B�P0M��kDt7٘⩫��0˶������k�����$�V�G��E��%5�禣�w��V��bֵ1�������EH��#ņ):�3H��� j�q��R7�ä����H�J�wh;R}��L��������CcϢ�ɸfN���PZaJK��1j�S�_$d����9uX㾲��	Mm�$��il�.3�E~�f��֚Iax�'t��ɮBЅn��3�k�n�5�1�rb���>""�t�rAJ�N����XhX��X��^7�$�B;�A+��~�
�z�^CA ���A�b̐��a�`l'�_]�&Z��wf@�Z�%3B�L>-2o #��b{�9(N;��q}Β1����WΈHi^luY^�~m�q7���6���~�xTߍ�p�m���XwsZ�6�U~�F�z�����"��_M7�:��1�w��5��""F]�9�Ϣ�a=�*�DXzF5��j�ĵ��y|�;���#s8�+dU kfo�V��C_�'��jI0Xu\�j��t��0�^y!�������:�D�ڀ�[�vRn;�y���V���lj���'��ނ\�Y�L3ujb`&Vj
�ѱ?(dpj��#��&Nt%��/��Ry_8��N*��1s��
5�j�|�lԛL�%Q�p�i�x(�)��{��fwvܑ�nǉ���/�q��<N.�.��Թ�X�An�R4x�����/�j����7�Ŀca�̆���f
��¤��|l5{��S��Ft+!�Hh�ψEB�}�f��3�)\�kE��Li��bT���M�Q#7K��Ho�YT~���[W�%0G�2���@%m�_�;�/�?�2�Ѷu�⦎�T���J�q'*�5����_--Vkm��P���3_�� ���s�~!wS� �s�W��7a�/��X$�O�5;@��o�����%4���,�L8�����u�~,�>4�FQlc-�r�m��ʫc����x*�+�yY*��On�����%�O��t٬R9<��n������E��O�p�S���$ ڜ&>f�?(���c=Enc����neQ��:`���Η6q�t'�1l\W�ӯ�uG��]�/G�Uj��n��L\r#���OF������1)��T褝j��I��_����l
�xYM<�RS��A����U@���9	�����<��c*�9yݒ����W|�����4��([a�A}��b�Ū��3���+�/-�y|����E�A7�.û�_�[�)o���Fhԟ_�|��0�6s�܃Uvg
�~��FJ2~hB���F+3ض����ۻ`
����Hm���	N�-VSe��|<d[�ҤSm��fui��D��P�yp@�݊��4�I�b
��	��|JYa��Qp�����}Y�.Бb�.͑u�Vi��:���7�E׼�8)hw2W-�S�K��q���}
���r�d	�@�Vږ�lR�s̱�'���Yo68Q�J��u>Ym�z�|,������g�6�}���?�����̞.Ο�v�Y�,���~a����]���I�`I���i"�Q���PM���9�* >�����e�4�3�嶦�bp�"��}䅿Z����n`��e�D�`&�h`8tz2Y�T �호}�z!#�)��	�Uh��v��A�u�E�
ȝ��Z��x����`��&��F�r��c�e�c�0��C~�4�'|
��)��&۳���i������2Uב�5t%Y�l�&�����ϸ���	=��L�)+F�g9�����ڱF�W�n�~����U8MW�0��W��m2�Ͱ�dh[��?yO�A*��{�.M�M�k��X%����Zm��e)�[�P������0�`ޯ��g���Eh^��Z7r�?����H����LB���O\'dOy�zLn糋e��(>�<#s��������D(��.�l���é�/�s�l����nbL�_so����"�N��B�Q��T:��ot:�eJ�"F��>28MX%]c��aH)��� 5W� f���.G��yF_�O�vY��E!�CH?�
�,ǵ,�|�&��Ӛ�-�QCN�LII�bS3J�]���bvu�8�ms�U�Ɵ��@��th�v��g}���n5��SΈY�:~��o.Y�hFH���A�j�ۘ̋�B����ȷ�F[�*�Me�y&���B������6�\��j�~�qA��%z�0|:ݝ5<NE��S���ᗮ�]��w��.)P��ɱ�^_�M���8�IZzL8DW���M i�8��k��d8^{QH��'�o�蘯��ސ�S2��nAo�[�.�[��~bxt\q��\G����4�V���iT��������IXˠ����^�7ԭ��� [��R�>����졃	�x��F�@]�Y��y�_��8��$	����8}���f��jT��w&�2����@�F(�Sx	[&��YϿ�hZ:�@Jܪgf��������% B�p7i
�!�%)�4�,�Ґ浛"�>�.�߲T�J���'5�ܢ'����/�=�?|���'�bU��;k9j�\"}��	���d�g�.�P�g3��l&x�3za�|�r��L6��_����k��Ր-����_X�]g��%�Hk����ne����"1�[��e`��0�Z�>N&z�p�y�_�,��A���c���>7S{�5����/X*28jQ� �H�2D�6�=Ӑ ��.0]�{�\q:��[x���.s�;K���dNE�C���'�M��Q�m��ý%Z܂�hgt!�%���
Ϋ��(kx9�kkЙ���E��B��'�5x�t6C����2�X�	y%��(Ib]��x�X�ޑ��W��	����:�l&.�Ⱥ�\[4��i��.T��^bV��37��a�G]�O]pH�$��v+�O�$���tB�N���n������[ۆNP��R���
�o�Ѵ��e��'*]�n·u��WF����V��\c���䉉(L�ډ����L�\x7~�,��m4��gb\�ȁ4��`Ӵ3�5��π5�$#�(e'�}�C�fC�m���r��S�I�%ǜ�/�Y��n[	'�bGP���9�[3T��~��/�	�mRġ�`��y����U��7Է"*"z��L}����,�C�
�~>�G�-�F|~aR+���<��ZA2��ٍ���Xhn%b�z$	>\�TR�O[�y�]d�GP��I�4�nھ_ _�:�=�Q�ӹ�`�5�z���u콝�%m[KV��N~�|Fh:F#��s���l`,��6I��&r�%`�%*#hfWV0����f��("��'���A��<�\����Ud]~�z�_�></�As���a�P�ί�����(S�=6���dD�N Ȗ�4�w�]?��aK<VK�A���^+��f}�L�~Qx�������.�덝�l�/k��
� ��x8Q �7=xI	�~8t]o�cM�|��ۡ����<�&@�H8��v��R*T�o��y��Wax�;�8��0J��t��N�*���U�.����p�"Wo5z���g���Xcz�Ɏݾ���W�8�1�]�­�C F�=(m��Fx� ��Ɍ�Y���U�H�,��`�����1"�$<��~:��m�֏îwcs�(v�g����vMʀ	oJ?�-�;��d7�vE�F��k������Q�?��+��(7�rdI�L/�vA�U3	��0,=��w(p�=A"�Yd�T�a�.����(5��:0j#���X`2�I����l���.�7ZD�h^��Q�0�_�}fg�]��He���(p�����H�+�N��� �Y�i����Y�pt�D��I0��˖V��c\��,[���s7$���>��彿�E�"a�� �i����`�p�c�^"3)��x���|c\'��R�+�}��K�p*l;q�]�~�7Λ���$w��VX����+�ְ�B�0h��=�1geX�G7�����D�+৶R�� L��q��Dg�5Jt�"�{5�XQی�M���.O�H�Q�G( 
/�"�@���*����b�w_�T�չ�O]�Ǆ���
��^
T;]>��ge�1z�+�v0�I��h���	�����rD��|��Ǟ2W>U�g|��'�X�f���SvH^�<��m�=}��/���]
���g�c�%SE���
���cӗc�P>ެ�J&��q����㷄y$x@1CQ�*���ġҍD�2�}��\y*���^�1X�Sȉ0���K�1P�cV(�ϙ�A���c@c����JI����aG�a2�^>2������H8V�F�p�-@`��f�^�x�����?��&�<�urR�����9w{�I����� �c�uX�d���N�}�a5�<�����~n4����9�)��ZoWZ������<�2��z趑)Q�URG��46
M`��1��?�3�².���N�+K�|��_�P�޶�.�5͚��7�b_%��K���)@3���(�����LQg�/S��S�5���3; ��Eh	��:�3�_v���i����� @s��0�v��oFc��Ly�$�u�I�MQs\���� X��)G���E%o^���ɀ�?��c������b�`�)�.@����!���S)��;�#��YI(����s?�l�>i���:�O��:��0̩����
kN��_�W+}��b*d�̩Hp��`O�40�{d�G;?+gym
!LS����ōP�|�ԧpj>ڪpy�S$t���-������#������k^#,"����:�d��6�3Oa9~X�O��bLV����� ���z�K[�7w{��R�����y"�Ud��ۊ�>%n�-�a&MM���a��v�u�oH�V|D�D\���[aa�5FS/Sh�!�Po�	B??�E<���ɵ�ہD����c+V�2���x��4@��#�I�$+h���I��㛇�qo�"^B�]��'�(�&Q�6��hϧ%r�y�M�*��f�{�Q 4'V"��n�b'm9 R���-���\�Y���UB)K�Օ&o�xg���<�i횅�q�9x�0ҕ~A���Zl�"����T���sUm�*<�j�xRo��܊�B�&��&��Bl̯��_��#'XCA�m��Z�=0����Y(��]K��ʅk��y]Ȃ����EHt�2�~Bz�k5�I��V��GV٭�.X�&�� � *E�Y�\
��[z�D���y��U:����#a��1�z��_PqП�F�#����Q�.ь�P�5�Tb?ƽ�݁�#k5���?��f�5���b�i�������]� ����!ق���(������������|2�tu�;�:�%�	�Ъ�	w�:?�EK�e�!ppZp����:���T��L�̴���[A�i��G�CP��?SI�W
�]C��jQ�e5���pa��$�O�]�m
#��� �������������Uu�7�T��'���J�[ZVcR�ю��/͋r��!G�?,#����ш���!kQ
ؿ�G@0�p#2Qw�g��D�R�J��΃2�y/2,�7������X�i�t����O��/]����S��X�&#g��lC��ӃB�<�Zԋ�(�~ D��R;+����`:����58i��v�wM�Ϛ�s�Oi9tp��EfZ��r����d��?�J_��{,��Я�Ա��
�/|���Z��Me^z��W��k@*�:�f}O팗}�n!�t�����	�D���o��>�I���C5ʱ��Gmʭ�ۖ�$�>5�5���$~Q ��2 �(%:7V�b�!}W�j�(-f������s�p�M� 	R&Q�����y!�G��l,[8'���mB���*6$�}&���hy��s
I�VS�.
N�,&��o��ӎ{�a� +�՜�Mߥ�m�]!�FI[�I�N?X#�JJ0qQ&v���㔼:��7.s��x�+��`H<D(�q8��q���)��u�n($C�j�@C8r^o�{���@%o!�dTx"�@re�D��m㖘P<�#�1_��lcM�m���ŀ]c,�ys�]@��%K��58O���m`g<8;���D��i�m7M$��@5Ļ�$M��4!��f��W3�DF�^��a^�'m����`�jQ�+�҉L����^�X�"4�7w��U������FT�!�{�˵?�������x���#2�;�2#���[���&W|��VD�U�_�ܦp�P���q�w�A����J��J@W	.#u��mF��uB�YG>��O�ʌ������R�,�~��*���&RNQ�T@t</i!�99�Q����W9�tw�+���HD�"�H��	�[�R{_uC,�u�a����Q�p�j$Ȋ8<��(�r�� N؅����"��ֻ۞�,`�'IģP����j���۱�������~�&�a��^��og-�Z��1�����c_: 0{��c+�0�H�G�A�$�'��_��n���Jס"{��
���<��(;z�����Ks�h���eT=�N�����+�%�&��n�=���˄�&@��~�C������r>��Q>�^��I U�?m�ׅr�"N��Q"TH�
bA��\�ҵ�����qo+�ci F[����-ј��m���Q�<A�WO��?�ʗ��� ��^�W�i��R��D��Rכ�9���s�sߢ���^\Fg�(�b� 6WV>&�â�ZGP��_i7�/�JGq�4_0�U�@1���70F�v8R����@20܁���#=�2��ok���N�]۞�C�c`���A%̣)X=�.������� $�ą�r;j��3��:V�W�f��� �n\��k�8lQ�w���`(��������e]|,ߏ��Y�K�/�ɔ���\$.�	���ioJ��i��K�N���a���*䮓��H�}�'��˕�$������4	+r�>X��ވ<a�v�4nǭ�xdD���t28�~O�g~f�2"868c�b}��!��\>��E7��1v,����y��	%�Aq���#�v���O����É��/1K�2�G�q2�:�u���l���~�V�-��	����\Df7�\ ��ư'���:18�����@{�D�؛ɹ58aMV_��� q���OahN/�ڥ!G-�,��#��Q��qP.�/W�!��)�/�=-{�s��Sr�l�&�^�2��/w��&X#���R��Je�N�V��X�Di������ɀL��ne���l��Z��(��FđJ&�.��.V�
d��3-�w�؞���e�5YL3~�F��AU�F�4�}���.�ziY�Q4��)D��ЎY6j3��� c���ފ��H�ҵ��d��L8��n�c`�!�_n�,�!�A<k�	vB2 U��Ƹ�d4����1.����fuG��,Η'3��9��X��J��Vzr�Ӓ=�z��x*,:�oc��6�>��&X��SZ���AF��@���0�(<���t��0sU�<ط�q��`J��g��OP����\�e	C|��>��j�:[���N���u�x
���0�3�C���&d&ժ�o�%��a�|E_���� "�b��A�C�b��e?��x*�?ߧj�b="۶_ܯڀ�FF��BIuúӐ�2O��i��D��3�m�H���s�Cla�"���a�{LC�^���s�o�U�E��թZ%�I���\X�8��v�c�h�>�9?�:�nt�s����j��7��2�s^�5�s��x"M(i
9v;M�r�b���H6����R�� n&Cd�'�u4�Zٸ�b�x=&�1Ĥ� 1�I̩�����cc�A8�3��U�^��皅˜��D�
b��u�G�/����>�d��9|)zNy�.�$�o��?"6n�.qmr�`�Ypy$]�]d���:�8jB�	��Sd.��UM�c�4`[��K�u�H$�ܼi5�G��
S;a�F��nl/��C��u�@q���-�!��Gyk��� '��}��^�A���b�0�_�䨘�Tn+�e���ш�Ź�0��`�{�1�����'^��P����CE/hc�]�ݪY�ǳp.�vZ��δ������?�ۘ�hT���3� d�_�&*4�O[����f�1�~���Z:����t�]�6�z9ҟr�0h.8�f�-�>x��^s@����)�W<�����Zc���Ec�:0|§�{}��Ҿ�tH{^*�#���Qb
��ؽ����DW�!ڋ�[,Z�
~��煱
�d�abVaF-��o��z|N-���`&9�u������0	8�A ���r��`ij�|�X�]���k&,N�1-�p��;P'z��4g5�3c�Fkj�撤�������Nu=�Kf������iV�Pnh|����wk?:��ى�M��e�6m���[��$Ќ���r ^�j�s�� ��:m��d͕�ᑡ��,�+­�j S��Y�eU�s2����+H�I���=�Bv���^k�:���3~8X񐖇�q��.�pU4�1"O��_f}=s��CѨ����jrh�۽6���Z���_�{잦�'&ڎD�;}����]�5�"�yf�-|4T����3"9'H:kI�6���Ƀ���:�׷n��%��N���ɍ1H1���rL��� ��hS��L�
���ug���e����Hs$��4� }�P�B;]K��Q0����EZ=$=�qC�zY��:����LٙX(^	�`��mw�c��,`9~^��e��+qzr�E�Y�-d-�S��z�=�N�4�t��,��͒iu�-v�m��p.]¸'�t���6���=�`�k`��)C�`qᒩU �@Ÿ#��R�s�*% ��C���0�߻��w����~�x/"Fb$�م�S�O��0@���<��e�Uɧ�m�p%}�g�<�C��>��ԡ��O}Iw�~�ڷ e[���ݞ��1��q�!p�v��k�h��}�e\Dt��k���,�~wQ����%&�,$"�-�e^�T��D9�wQh�3��ײSN�\C�H���+�'��3Zf�4��R↰8)���	�����Vn�c�0@ ��_�r��o�I�@}̩�wul�����yu@�9}Pw�!GǱ^B���Q��UV� CM'���h�}P>��B���6����W�����b�&B�A�6� �?������غ�����,���	��E�Z�+2t*�͏����}��ަp��	�G�����$[?��a��Z�U��o�����'K�->π8��2fJ���+��z�=8g��Țz����q�s�V�;(GN!���谏U�ͥ�ۯ�[�Hy�{m@��_�T=��~������?~ƹnG�a���H�D:��AQ˄ݥ�c���f+��
چvgn�3݇A�GmW�X�U>n�E R㕘�e1�z����X�_���^�_��Y�q�Y�-Ru�qQ(a�0��Dڴ���t� �SH��T@����������=�L�vMW2��8 ��~�b̨�b~����F�|��mϔ)q}W�\��Q��a�3�����.�d���.��'=
��hYQ[�Hi�ޡ(�[YcW������ZyE�=� �-G>��C�=׉"���(�Q��#���թb���t����zc�wߣ*�o�P�&��lu����1.����Z����z�k����q"0�*y3�ji�U7*vR��U�w����r$�îc�?�S.┇H��|=�lT�w������������e�?�p ��C{��v�g�Μą���m��Gт^I-��$q鶉��d9�Oi�"Sk���M�-�/�]E�(��C�^Ck/Ψ��XÁ�T=��e�9�
o���B��M9/Y���J�5�iğ��A���P)���nv��=�ć!u���6�*h����2�Y'�,X���B���nK���2�\���O�b
���;��ݨg���*� ��!���aOi�m��?�ۊ��-Y�1>�F }�d]�^�.�k]q���/���X���|yNM��������tk�AT�Y|�S��(��3r���>M�.�����Z��B�N�4R(����@�	\��K�)��L��drX���U�cH����F�J����nm�����		D�'���y!+��(*o��t`nZ|�+%^e���[�O����`~-M��,l�P�3�S������|\���~nDH0@:�ɳ�+9�����V�Q+���`a.\Q�G��Qo?��<D�L��mWy<l�"��p���'16��73xAߵϰH��ϣ�O_�$�ϐ�����ɑs�0�	�!d����O�c�76��U�:
ޙ<=��Z�&����c:�}��2.���ozOk��M�:��ֵg�򝸽���p��tōR4ٽ&^�.�Kt#���4��0�]8��0"���B�Q�J$;���[��'���,�k*O���R���h�������Պ��(����3�� �)8C9o8���,(:/g,V#�k�������L�����(p��t�8���W!₾0uu�ʬ���rP���8�[{�Bk�z�x�ָ�����������i���]a�]G�ӬM=��ȭ7�QZ�M��,���+��O-B��K�Я~�zn�:�`1�C��:`�4U�c"LӯѨ%A ��:dhƼn�o(O
l�w��3C�.��pP�O�).�lof4u��uY��+�jǀ�J�����ahV �B���f_�����&��tK&4ȱL�*(�-��A��+n�θ���}�>�nm@+��£-qQ.y�[#�:W	$-Z��~|�h�����^6<(&�M$*�A�L�4���=���d.�#��ro\��s?q�?+��ϐp[q�9�f��2Ý ��Imq޳�G$0>�ң��>�����t�x֏���/���=.7^�MW0&��G 2{ڰ�N*���F���e�
Vz�z�R�O�d���c���Π��k��z�D�t��:�^��3�ȫ{ݮ<�
^�'�,�i	�rj�'�XI�y1\�����Y��O��>�\�u�+�f���ʥ�o��i�^^�0���Mǩ�v��̌�c?��
�2*w�|�T[p4PT����	[�ag�������&���a�ά��TG#|�lH�c��(�2��$(�*o=�"r��3��l��]�%�;�6� s�������>���>8��˄t�֌���`�Eyy�E�*�q��_�0�s����9���['9�_��}������T�h�f8Ztc�uN]H���u,ٻ����<��dt5�8� ��	 ���9Cf��f-�6dι��=�u�b�c���z�f_n7�CZ[�wX���6�g�~@+Ϝ�+W�8 ���eT���7-:;�V4�g 5�!n�h��Z�Q̲&��]��]��z��m!� �q�k�o偑��Ը�_rf((#Bkh�y��T!X�@� ]%I�2�~�$��sF��*,Z�޶E��UR�04�E���t���ϋ��864�� ;U��bj'�V�p��v�0���I0y��]��-�WO����v�dT���J=Es���J�o�۳�=Dן�c�x;��C��>�o-�iE�qB�B~\Y���㣽`��ek���. �S^5ħ�=����b�?y�������p?E&}F�+&
:ɭE�(k���*o�r'��.鼒?�ԟW��<�r6��`���L��)��=��Yv�7�<q�{�7�u�2�'�����g���Ù�7�=T���e�W{�0���p���Y��W.FQ�y�yM�&�����X C����F�\����"����չ�0���	}�����m���JG�N�r]l Hڀr�\Ue�S�����	Ov5���O�f�f�'����4�R�e
�UDQue�J93��bk'�h�S���+UK�-�>�'��q����?��뽶�(�;�C�1݄���zF��>�7��F�������Wi��S�� ���pWvD/$)1��k����U<W'C�z�s_�7��Uֹm��y��RG𖇾hF��P3ig���xN61\Υ�	�5Q��<kh��MD��li��i3'؅����,[�hH0|�ŋ[9���uO�������!�@��H#��lٴ�+�J|�`�&?q1խږ��Yg0�*��w��sEm��,?�q� ��b�a�@���1�>]�����c:�{��6�i������>��<�v�鷡�K��5��x�I�a�:ͶR�=}I�V�D��S7KI��R=�CY1��,�7�����j�\��,b��n����?F/���W�ƨu�QNGe�{E�~3(hg�$��ˏ���u�#P����_X|��w�/Od��}�WPq�8�l��MM�ֱ15�����]m>��5���7����m�E �gmc�a6"6Hx�� ]��s��yC\%�5�B���5�Ӯ�sbA%}�j���&$I ��d�2U��筑g��>����28$���ߟ���X�d+�JLap��y��;��ܯ������SV-�D;�*l ��,}<G��/q(K�O��#h�^i�8&��T�Fڻq���B:'�d1u�����/ң����Hb%э&2n�'�?h��3��� Q~_��4�&�p
q��O��\�N�n��o$�!f*��A1�� ��m�T�!�����wL`_쯒<^��%1�d����^
|��R��i���9��y�!c����%��w�2LW@_���A��x=��R�0�����%4wd���v�k%�UD��|�DG�-{��_�~��kV 5?,�W�K)cEY�tA�p�0���z��]���!��v�.��3x�J���^)Ց�ҏF�쨞�n���㕝S^}P� j�bL]��Y}��@h��L��ran��̡K ���а	�["�j/5�9�X�R�	r'�<��u���xHRW0zǜ�k�4m�	j�fك� �0� 5ݲ���8�T��:���8�k ơ@��b�������,|�99�G����� ���>0ٖgֵ{1�V��g�}n�q���Iǋ������O*<��xT�]�ØGok�o D8~�ƫ�W_��M$�I���=�B�_o��9�P��I.;�5�����-����#~�~,�~�c��xx�s���Ԝ�:>��rp�)�jSٵ�A��E��po���P+���%�f�.0G\w�m����p���c��LK�����{˦&'S�:!J[�0�G��lT ����[j+�۲&	;3�n~�g؉�7[l
ņB�u鋑P�8W���ô�S�\8�i�7�w��|� V���Ax�M1���Q��n�b���7���H._,e��G�#�������{�q��v��������������Z,¡0�7�d��wʙ�ֺ<��q����G �C��A��f��)�'w�{��U}cooH��)a����4<�a��"4���4��e��S��݉}@X���`�ό:�6'�!	�қ0�y�6�ˢ'��\�q1����n��#����}V����7k�����G���n\E������K��~�;B9�:��R�@�Z[�
xRoZ\E�f!�A�S����W%H���� t'K��	?�	B��D��0�������#���M?8ZԵ֣R�g��{(�U,h���z�\�!rx�o{' b�w��!:��v6o�J��W[X4l�@1V�!�2,	]�}��l�Ui��1U+b�&�05�[x([����2�3�;.�%�wx���JZ3,}���^��f sE������'%������T�LXNRyf�._;/��4��QH˒��=��B����]�_gH�R1�GK�y��Vy����Ui�=?�c��ZJNb�ЀןX��V4����È���s��IL��`�֚��8R�`��E�fd���2��w��<�{%r*���pbg�C�o4�iW^R�*p��?�0,���#��싕�ƚ�t�I�䒁�R�H�<!_C��B� i64}������Hlk����q��آ@9 Ӌ7������@�t�y�<��$���Xn�Y����MJ�k6�j����C��ȀP.�%��[q����'S`�R��Y_A��p�!.�loAϗ1�1�Z��&wp�Α�^B����Z�l��C�R�`��9��"�R�<~�����Jյ�2Qo��+��d,p_�\jS�('��{D?)�LW���JYT�����3F�[�Fg��( *�P�"+�^o=?l�Q�!�~|:y�^>�����6n7:hǩ��d���[�r��)Wu`�c:m�ti�VN-%K�J/&`Cm�����q���F��_A��"S~�;���:p����s�U6��Đ��i�"�Pq��w���(���X�j�`XG�塈Fj��ʀ 6SA�|Qt�_]!7���p�}�M�=��#74х�#�c�~�$�s�A$p�3��E"t��T64�a]Ģ�]���FT����4ϔ-m����"�Yc"��#�U�ۨ.�5X�Ja�4]�㭭͟I��0~�r)2�:�r��l���>�̇�5��(콦i�J�����TRx����N�ٿwTȥ�5r���L�_�fH�|x��h���u�~�Vz�.��_�K��E����rvM.�Ō V�̮h�F�����v]�HXHƷI���d3���k,{�;p=�N��濮�R��y}mCU<֢�? ��+ˈ�#Õ�ሹ'Y��9MgT�_"a�CA�Ď����j�״|z�=��\|�	WZ�?�+�h�����ł��\Z�.=q��l
 trsύ=h7I}C4�".�p��?��ǐ,���WC��u V�!)��T��/��pqb���~>�U$Ʒ�)�C9%�>��/�s";��c��[���U����vf�5�z����sщ�]�}"����;#�`W�7P����a%b}mKN����ᩁ)��Pώn�}�+��P��=!�8�s�-���Ŕ��/�{X�������ߠ���K��OB7ނ&H�2��ߨ���Fcza����.�r�� m�̪S`A@-�������3@Oؔ�a�as��C^�Ҷ+	`������2P��](Z�?uHN��
;/L;B�}���<@.�R�> �/��TM�˻�J��V��\7�F`�濔ik�b���������>�Y�l��|q^zH�]uT��Δ�6ܝ�8�(a2AX?���!r5#:.̙�$Fb���d|a0w�1&Et�p�2j"^%�㊦\�e2�t�M�9�{�W��=����u;	.�w����LY��d���u��>��܄-�]Z朲�����BsKhQ���I�9�-D��Kn?J�e�ȍ�yH�O<�[AT��]�*�Q���5���c����L��.�{n�h�85up|T��Hӫח������GB�"kȔ��I߳���-2��
��F���\`�pI�"�>t�a�8�l�J���cf��>hJw�vkY�r_@���Zk9��훛eB��Z�(��;A���̷�cM��� �xI|�,�K��Vza���vAG1��*>N�z����H0���scW>���;�-��nҧ�C��ᨱX~����<3�YLl���sB��,on���V/�M��=��9o�H����Z�F3�O	��� ������E!f����������h@�%�l�e!t�R�F�0ne{��~WW��x�<D9iM�ٰ���^�Y
�T
(8���WD��f`st��3�h�q��K@�^�ïO�$`!BHwE���c�M����h�u�ls����*OxrA��� ׇu�ԩ)�V/�"�6.������\������6M*�����aVWMi�i���y;����p�k�t�1ɬ�삨w��q�U5˷+1i�q�X^m�����9	J�}sҬB:��{_�%4���Xy!�T�v���)�6A��H�z~�U�\j��=@\��?���<5��'�7�sB�?)��*��:�� T`�t�$z��,�����Enz��)5�-���:W��r�7Q�@�Tq?���@Q���A5���}�2C�	��PO�TȠ`���>�r�����}�uz��.\�`�a�/�5ŮO�ZMOZY���OH0?��Z]	՟�I�E�)���)e��7 )��� Pd�X~U@|pZ<<�Vao1������8�fOC��5t�}f��l|����N<>�	�<����+�m�z{4�?����q�ǯ5��X���R(٭�)ꄧ`=|_��m�Ѐ9�I��@Ɠ̕�]r_*m&�$@q�;S��<��#��I�}ImB�s��$R'�OHi7�k��x�kz����v�Ln=�lA܂/�R�;樏������	�M��f[�q�5%��;;ĺrc�IiF��t��F��s=~d��<	��}t\��{�|x�0��d(OwG�3b�aPC�Z�y|].�~ٷ��F`<Y�_�9m?�s��2?�ǀ��D�x�!&�N�P�K�C-ϘD��2����hh��)�AhoH�MD�.�a!UgzK��#\U��E�⁑�b]����+{o�8_�K�ƠR�����#<zy3��|��Q���B[�VE�_eC���,+��*��z����ͭL4M��>o�ٴ쉩���8�5p�ʕ\���>�]���[1;�@��"[�J����-�`6.�J�G�w��Fj����/O�(Y�Eh�lF��+��TZAL��І+�\��T%g�1]��5�TsW_5rv�a+�F��3Y�^�Q]$�v�+���?��}�_S���6�b�Y�΋(.���O"Z6�
f��,�*��mJ"�
I������g����H^t�R���`��-U}$v��?AJ '�:-+�α��P��r�ҕ� ����*�/<w�h����C�y;w�EB^H����4�_.ÁZ&�]8��;|�,*�R�H�&��5J�9䈕?e��'!e�7;�W�XvDq��M��p;&&�&0����؛���1�w^�ḥ�Q�^��J��/�H�s�W�8�ۣ/���3*{+�a�]Y��;�#c'��5���:LOy���`��B.��g�Ǖ�_>��
>@�UH�q��z�-LChzs�9�>��=�zw��Qf�2��JF;/ٲ�7�k�"T�����u.�C�'E9���1<(�)~�<�aFS����@d`�r;u�~d&�?���܃�����Ѻhw�T�/�����(K��>��+(����e�@��=��!oO��`i�_���7O
mz�� O9*M�ך\�u����џ��!F�O*�Qo�� ���m j֊�&�<�{��L�B;$��&��?|�;O�r��c��H$�vv��#���L5=߬j�"��x,0�X��.5��7�ϾB�1^��y�	4��}�9���������Y`_��"n�t�3���")hi�O��
̴������ �_%��R��7Ha�fH�x�#�t����n w�[����(�l��iW�ه*7�bcBg���o��D�!n9Ƨ��۹ 駞�#x�\��h�A�:���{��׍i����=h��?L��q�m�ف&t���)jv�<8�cZh�a�V�ܷ#�i�H����BP�HAt�Ď+FA(���d��8���e�4����<�z��׉��I9��%�#��(�J����5b�Ճ,��.�4�����81Ś�WLF��>�(�2V��������/V࿫����0h�h?8�Ȓ踈n��Rk���(�dCXE�p�/���	q����Mu#2p�;)G@��0	��������X�#��Az�v����R��	��eq���(mtbG�����^Q{:�9[컸,h���^���������/�D�y"�����܄C�@��e�	 (�gF�� +�E��lJ��q{=�`s�����k9E@���!H��M����Z#��X��c]�<ٸ���Y]F�ٲ�!.G�Y�>��>r����b�n=�~�Æ��[*�w7��|��J��M�}I�܅eV�]��|	������ '��,{��`��2ɮڟŚ��kJA󓹛��ue�@6j�`�ءn�-Mq���l�,d}Ӈ�V/�#7�&��W#�N�B}]�>�Rh�Y�r�ry�k�vA'
�酞��+�8�z����b���57��������v�H�Z��"j��d�'8���T�il
^��̒XZ(����6���f	X)�4 �H�L"�9�����W��$�K���2)W��5�G�kߢGKމfrrji�pF�����,{
*}�P����X���v���驮�JUp�8�j�W�'�^�-�Y��j'��ߠJ�/�$¤�XF�d�d4K�h�(g��!�T�o;ha��;�	%2Ţ�1�^��=Ŏ�Z��\E~;��.�o���[�J��v΂��h�@�*uZJqK��������>�8��r��]NCm)ge�xc���'A��Gf��0j�qLuH����g� rZ0�����\����<^�s6�9�Vg%޹V/lh��o!�"�:Z�A07��55*��d?��v4�⇘�:�̀��>Ɗ�L�H���$�ǻA|�u(��i�A]�X��aX���66j�5�XG�9I�8�%*/�+�����<����B̈́����-}��-
'á�3��N���u%R�a3����U|X�KYAz��:�}�'i��x�N�8�eXGK�eƱ��jEmd�ؼ������� +�:��u��	 N�$G�����N0MJHzѐ��D�d�l_��R��~�8�(O�n���G&�9�?V�9\������Lmo�~~y�h}jϭ�v��k��}���U����I��	��3X���6���C���W]=�r���+��ź�v!����/L#|~�z�7����lm� �î;��Nc��V�#B�=�_�vo����כ4�A�|Ǖ��e�RS���p��߇ُ��>�&�~�T/H"�P���Txd@��S���t1�LkSy�6,Rb�' ]	�-{�����>p���)��?q�Ŏş~k��Q ���5�����+��m=�3�,���P�0@{5� �M
nU�Q�o� �j��(r^�Q.c�`
>Z�|p�9��Xw�s�X�6���(P�y�� (o�y�.�m'���%�فɀ]��
z�R��J���}N�$"�>j��B��(~	�=ھ߻�ޒ�M��\�6��<�)�usw`5�*�,��Y\�`�6,��U�Aֵ[#=F�.s�������<�7Q>������c���@�nD�|I �:���09��r��	llҝt-�?3�
�F�3�p�����2�e?R�I����ZVK�L~��Jk(�V������1{�I�5ph{H�l��1�P�G�,�6��q_n���y
��ԽwJ
�h�ſ�|T�U?Y.�D�m�ަ��*Lo��x�J��DeowAL���n���%�ghI��%x�!���F*Ӎ�G���+^�9����Z�+\����?�c�gz@���#���&_���1�R���ck��4_����]��u��x����Hz�ȸs?�<K�J
>��~	5dXE�߱^{�.�	�iS�;F '&�p�-�:��OA������Q}����N��z����H��)��xt2,��4�7 F�W��X[��D���^�e���9��G�n�'	����lί�P�w�#6�4۲ͩ߬���+ȃ��X�\��l�U�8��'�[���ބ	:�Q�����6�eo$�75�����{����a��L�2`C޵� ��Raf��s�
�){MK��4Zhr=}��_M�P4���&��\�<lKg|������Qo_�1�r��+f;%p�
k��������F�ʩ�$\�ԓ�/�{^L���}6�8#$\>q��4I�4/�Xp��ө�n�D𡤂|h-�}�G0��33cÜn�S����<zs���mF����E��!p(ѳ���v�:��h>#V�j(�}F3��W�-RJ槁�Xj��2q'�6��'�����m�.��QhH�8�r���FGk�fm��K��c�RǼ�hc�j�K�����[i�q�"���*j"�H��t��?��o��&���k�� ��G�YtG̪�yýT���^� I��W��*�+��vٷ/[�>.e�b:�G.IA+�'՞-�ou"0���~�3�c�x,��츅�RC)[������m9h�Fa�4����+��{o ���x@?��(j�d:3�ν�j�z���&S.n�ϛ�s�e���aY3{?u�f�#��Rp(0�-U���>���s�r ���b�:�-~�QS���n�u�ᱠ��n���äá�K�l�ٺU'�{Ť�B��-�mn��g�%Eâ݈_�D�0�m.�,��J��hRMC��_���E�U��&�C���F�7��������6��:ԅ5}t�5�p)^�T
�}������C�S�rRJ���i�͌�`��}�
���
*���F��.�����%�6�mF-uE�[�����ao=G���/���C�xl�
?j����B���A���� ï 炙�]E��ѠM��y1x�ܽ;�h����~pAHz��8�������� �>���v{M�~����b6o̦'�TT�&�[��r�����i|ŀ!ԟ�A$�-�,d�8��j�0����5�\j����%*G��[=g�/gF�nЎ��mB-�[L+lhiɽ~+��eU��8�8Z���B��3��?��=�5�0��ф�ߢg�����m�}����x�i��<�`ވ���< Ze�y�,(`�3�}(���C{UD�B@M�Ýݐ�'; ;8�O<UQ|M	xo�ޔ��!�>�e�~���@s|{��$���z�g�����SV/���I��Ǵ?�=86�H`�+i�p$�R���An�!�)�P�=�w��I*�u(�Xʆ��.����.П��O�$w�����h�;A�J>��eȟ����L<��3u���-!U�ud�+�ZF�u��2( ����t�A�qKJ�`�h�����}�E�0.�A�+BȤ�x!!J������v1g�p�rF�Z���������\q�L�b��i4�p����=I��� 9m�'�6_�����҂|ҋQL��v˭�����oR�������.�u��r�W��7745J����4�y;,m�����o j7�ډ�@�s h�PGo~a����$��ɋ.��Q�0���,0�!/���@a3�3M8#�Z�d)�cz�h���j!�P��7��5/�ע�W�G���B�[�����6��CS��+�Θ�Z������JY���Q@RtK��g��̑��!�?ݯ�I� WՓm9�T�3�-�k+ ��~�������o��i,
�j?�L1 �F��	�"-<���D�&\��,+�&\��V,��1-#��g'y����-�(y�$\q:5'�hN���V1�v�PF��ግ#tv�h~lDU�Op�j:5٥��6�V`,�߰j��3��$ѡ죃���x>�.��!3��{3j@]�6���9��B ��������*���޴��5����z?z�$r#�u����z戠 ىGNx�	�9�^-�?d�cu?<a��/�}k6�wjQF����Z�rsV�`�����m����S�ǐ;�M�,�*���;PX!S�:��`-j���aƿ:�ƨ��N5k�>,G��?.�o@�gC�`z�&jJ��}�P�y�o��@u�I��*�/�k���9ݟ�p]B'vN���(X �?@9w�b&���W�AF�C�˜c�T����Qe�uh-t*�V�4�������Z��|h\��i�/�7�;�1r��_AbTC[��-����Y�a�RO������-T_jO&���RF�!��1b����R�w� :��;�S�-��磝���ٿ�����"��Jp���T�pى ϻiȩ֗@9N��~�&v鬪M�p��ѭ)w�R1��}��e`w�?�&�^7�s�-�|��u ���`����F~�cN�O�Q�E��!?�Frz�KL׸e�1T���x�^��b�w�*k8�H�3	��Xt�	��+��q�imx8��q�~-fl&��Y��K��4�^��ռh��p;�M��#;��[\D�~�Xĸ ����M�	�ng=u:Tm��}��7 ��Qfvk�]b��ڙ�K�����],�&���h�" �"�<<Ą�#����&$]n����\��0�m��� W��貕�V�U�;uh߅� 3�6��uH�6.��M��-f� ��i)���ÝW#V���H��vԿ��/ӎͥ�_��pA�Kj ����D���Z?�1�����K���i�����+�Y1�s�Fh���S�6@�.5U�դw�%���9w�_��|fˠ.���=�gt�����x�/�ND����pv�]��n
����_G�됅��-y�]+�ף�LO���N�8DX�1ٛū��n�Q]��'��l�]�����cb����!����fuw�D_�k�7�����Ad��2rn��9S�vρrQ��RZ�x=�)�yG�#}�{��L[J|Zj�*5lm8bʕ�DMք�!�)*�ʹ�ng )�,���o��C�_<T�scIk�.ƫ|�aU#�a���Z�(ٷ�����Z���3�KP��l^�D���­����.�4�.3�j ��4	,���3� �X\U�̟��.Ю&�5��D����5Z:e���a�|�Qa�HTI]��)�t��:u�;	D��?P�*�
vBvZ��i\v�q��-����F���~`�0��� �=����+%˙-|_#*)�en%�2j�]Z,����z@ҙ�����;�m�G�
OBaC���j�x���!$T��m�o���Y����;�7;Y���؇�_6."1��mr������4�[K1��K��N�6�r���%\0�\f�~�om9�)`RÒ�Z+C�!=o�1Ox�(m�]�y̞mf�Hf�������g$nB���h�$�^E�Cцa�6�~�pݎhU$�6c�1������\U`��v6Hdx��t�bSl��|qIBS�fj��ZN~(��JJQ�H��Fu+�rc��2ؤ�96�H��\~�V��K��F{��<�l��?�,�=��.H@�㲕�u�S$��"v���+k,�R�%i��)4w��d��x���yǙ�}�|�\�׊*1f?���	��[�U��cf��hq����}�����V���y�Klр�͝�0��6%��Nh3Qq?}CX��_#i�"O\�Âuoq;G����6�&f��O=y)H���wðG��F���A)�:50'J��� ��ǝ�ۅ����25��� ��%$��v\Q�[�]��Ŏ�ߦ�16�k�HZ������,���E|VXaB!ݐ�gAp���|2h����8�b	<jk�ר���/��T���p��2��w)���M�!Mbn����m�=r'�ѳ�u�?�����Nu)�2�\a�v&��C̨$�պݏM2^��QG6�)(��=�|�$7_-�.=��C�W/ɿ�M���Z�N��<�9.��=��`ꏶ!1���5�蜪����Q ��oԤ=Ӱ~@ۿ��L����=����é[O�l�u|�����Pe0���Rf��+�m�dD0��-Tꖓ����ω&���!�Y�	2Vg��t>4����A�󯋅Cm1nih������ۛ?y�ժ_��:xh�4�k��ad��p������ݸ�4�}�-���5�����;o�DJx���4ה� 7x�k���B�2k����ͨ'������1LD��Q��,��6<��y�ӏ�J^#��p�ӊ����y������(�y��B�k��r�r�+��-^��cB������{��R9y>��o�M��R'Z.�a��ꖏXy>�sM6�H=F$m�����*�v������6�2����&ͫ��V��_<�s�=�>��v.L-�ɱ��<�Xp��M��:�;VAhFM7�{��S�H���O����T���
".M�Ћ����j�1�60�2���Ϛݓ�"��3QG_�J�l�@��?gprA�%��=9%G{ C���c�^�8w��l��)%'	�W�RC���/��v��<8ڄ��)�}��л϶�8~ߡ۫Q�?L�慓ʶ�RےUF	ӏΊ�F�Ȝ��V?��o����h�B�IIE�G�9���h�'�bP��r�	�l�$���f�e-|�5����MQJ7C�#�v���S�ޑ�����Zo7� ���w����hq�k_�s��g���L��_YF����������%ݮt�Lb�gaZR��(��j����hG��B�כ�z�1����ZA	�
=˂ͬ�+�˛%9�,�-Щ��y�Sk1���|vV�A�Ms��3��V�^�{ӥ��Og�}�3`c�'�?P�J�~���ӦSA����퉮8��,���L����̅��dHk���ͮ�a�jg.}$s�(A�Jt�7����ʈUo<M[�� �:�����	�F3`m�:�9�Š��z�E�q�+z�ViluOv �+�t�������{���ZFZ�g�2ꯞx6B���n�#N_��k�܆ɤ�Ћ��"�<��$d�J�r<��s�^���2j��*���傋���]�<��F1��������{&zͫ2a���8�r?ɞ78y;����c�����f;DpA�	�"ҹ�ӧ��0y��:<(���<�o&��4([na�~��B�;��l+F�f��;}9��c��
�OH��'�$��� y>�$��#����Mvg,Ъ+�ϙg�p����sxf�^��ߨ����+�c��%`���.6g��D�΁o2�KӒ[s�`ģڞ��$6iye=o�6�@H��#ҪA�0@�"�I�,�PY����?�0&8�Q!1$!� gS�7DS��ª�u��N?t@�[̝��jϣ�?�{z����;ʊ+�"Z�����Ǧ*,��!�Vx�`+��0�Sr]��Z#�:8<w*�0-`1��6t!�a�g%<��W����G2ۑ�ho�B��`�QCD��UOߐ�r勂��~���}*�FD�Mq�в��ۛz`�<��� ;�^2��"�0Q��+�@�bɘ��3oJ�g���te�!0��t�츶�%��S� �C"��EGlkwo�_�h��b
���7B�+$3w;�5j7��P��o�f���o:�Ohu�ܥj%��;�n?;�� *W�񭁐�-�>��V^�D%W�j[6ߞ=fx��ۡņO�L�j3�
��NT�If8�Al~�i�r��Q���[^;lg�a6ҋX�[j�-ֻY�i6%��Q��ܧ�izU��i�OOC���N@�=ы�_�r1aW��ݘO�X�6^Ḟ|�����$��;�B���]$�4���<=�f!�#����T#�m��ťʃh���y��w��h�@6���}p��u�<{���Ȇ/��{C�h�����Ȥp�V��N���<2ZQ鴼(����k�།(Yqz�Q#lQ��,��]�}��=\K�0z0�.|�n��z��,�[�����B�{�~��:t��`VO�(��k�<���k'Kﭩ���s�s�9#�0���������a�a��Ӻ�54�F`���BF[��uϘ�H��!_U���	��!��҈J��<Z��Uq��~W�ݾ�ܺǐv�t#T�b������H|y![����CwXR�ێ.,�����4j�����mxM,&��t'��-	�[�!U���J]�w�f����a�'��ɮ�?��p���0䫈D����'5�vxm,2�,$Q�1�=%z�%���D0��z)�r����^^�K��Q�f���*���i_�=V�d:�/	ν��]�>���Q%�dA/!���y+����k~��bշ�����E!���V��
�V�	GZ2W�`#ˌ��Y�D��ɫx'>��t�� �5F>]�E�}���\�{ZRx��6%+Ƙ�tr���D�G�!QZ?1u���*�*����������>�ޯy�= �h\p�!�a9�ᕩ)%瘤ŅP������	������(-�|w��|5^��h�+x����a? ����ײ�V��[/�9��ͤ����g��w}ر�f|��\�\@q:�&�7r�����:�5�����"6��5|.�����5hĈLz<w��*@ͯF���ge��&1���.&�T_Lĳ��T����x��d:�5���$R
�1��GY�~o�[�����Zف�_*�ά�E�z}m!?Oٯ�:��q#
�@�'�$D�r�� ��
�m��f���`G�-���d\C���t��7N׊:�b�l��dK�H|�obSR������~_�+��{ͱz���s
s�rabdm�x���ק6=װ��ӯAt{���w�]X`�~ ��}h�P����rO6�Og�J�����jJ��h��6��_�+��/
���*=l}`�� w�R]PG^����׹�.����|�{ˈ	�d�����'4��O�`�q���l�4D�`����0���Cg%({�j�>�������*��0�n����]��Q��Ƴ> BL�A����2:h=������Jjy�:��8=1�"*53������cХ�wH��h�(*�<k��9٩���I�,>L��D�נ��~���?��A��	��ȱ��i�w����J{-�;�{�`<
đ��PW賅H���b����	��|7�*bb#ZT�H�잤#Ipz}t\�O��+D�V(��Z�v�E�XFL���7S�h��ST��]h?K�&cdł����7ի��Ԣ�&~�Xr��c;��.y��;g���ȷ��r�#�oGb>�z�0 �o����D��9A������Q2� �%��Y:]�3R��q!��z��7Mp�����(���f�k�����_Ua������V&��ܠ�CŽJ�\u\_ѐm ��+o6�h�"_���tGt��|���l3�4@A=-��3Z�,X��&���@���JR�D[W��+�M^c/�1��H�P�9�|����+��ΏT�Z/�
���Qޗ����X�������5r��>��H�u�F֚��-�g�	��
�D�)�3ř�#�����$},V�K�QPa�עey���>���yz��(('#y&�ԃo�)�(&�g&p
��F���3N�J�a�4���h��擆*Ҷ�)l�]�0p���Z���"eLP��O��X'�����ww���p5�sȔ���w~=B��5hR�Pp�  �����'�f�1n\�)^ax�!�c"g�����w!���T��C���(������P���X��!J?�I?�w�� mٞ$�z�e��&3_E�$A���Oe�(�^x�Ǡ驪�����'GG��3n)�gt5�)&DY�֛z��%�x�|��*Qv!�*n��� ��<���'o�؝�$��=S��������l����T�B��c�|��&'�|Q�����g\��W�I�R
����D}>�T�t���� AYڜ7����d,��D�+;J�NC7�d�]�t��#��a��P�!�ƻ��T�wˮ\,;�.!'���y{���I����e$o' D�L�!I��i�oz���|Ɍupl=�M�.\HU��2��{b$��Pw`��b-=[�Ƶ��H�1(ic��#�� p�<�s�^���7�h��$��N��eO�R3�vcr�m�\}a�n�5�� �� �*fF�Sizd�L0����Lfhgo�Ei`O����.9��!���@�2?*߃���1������_pf�����B���}385���d�0g-����(R#�����_��=�W�nY5uؽ�vv,g,8B�r��צW�^E�(ɓ< 2hj��f����[,6����H&���6%��
���p�k����K�2)C��0�g��3� &R�B��`�3 s]���Nw���
ؼ�@���+� �@L"5�lk�.�	��:��v��r#�FF�8Z~��_lx?�y0�3د�h�}�
��M������9s���yJ�q��SI\%=(��u�4í�J�V��8�-�0czNr��cx��[�kx�UEe��υ���mr�G����{M�����͙O�������e�����/�0!��@��}��t��(G�l�0w���U��=����j�L��'�o��5��~p�|�<�-�̺`�-����T�ùJ�ė5p��8��7L���V�T �	߀�s~�V��S��l;8̎;�	�t��ȥ�x�(��N�RF?H��`m�n��^��'Ԉj8n��K;_���T
�i� �a�"�!�8�M��̟D��0U<���T�Iy�y�� �i��܍ ���BW��Cy�bΒBKuK�+-(x�W�,�]cȓ6w������ �o�"��y��Hs�u)���W ��(�լܘ5����^Iݽ�&�u�L�h>	q�s�|�ۋ�dv���ݶ����N�WD�i�9�/yV�?�9�!q����~�Э]4�t�j�D�9�ݨMa6�t3��
b����-ƙj���绬��Ɇ0�dܳI+����]T-U�v�rp��|Dd���
�>����A��u �����pqOj-MY����N� y��e<�k)&j���ٻi���F2~'�X��(��&U��b3<�P��ipS��/0O�Y6����O�ve��
P@1�";�[�Fƌ�)�r1J��)��$�_5�L��#��dT-B�3\��n��q�{CT����-�`8v�����X�|Bb�D,�SQ�I*x~��Z�0�g6.)@u�׬���2$sT;sy`eo�o�w>�kJ�
�ǫ�Q������zC��."8�QH��*R��T)=7�"V3��IW��d��s�;`ZZa��\=�Y�-M-��5��#U��h5k
8-�����9{_��o�ҭ��1	IC��Fb1Q����~K���S� b�8��#��,Y���<�U��c{�.kذ���n
AnC�;��~�?'��N[b��f�JaWca�0�R��v���~��o��� �ҁ6�����Y��v�݅�:u����!���b��V�MsD��f=1�1��f�����˩ڭ�������F#��SO���*�����Oh i�_�_��)s����*�1�ݹ�TR���'e����ܲ�F���o�6�(S5�i��!m�r�u�P�R�G����4���F&0����y]�l�(���9��B�*ʈFy���Wv|	�Oϣ QKdJ����-FO9n� �GG���Q���<̝�(��r�8 ��@*�)����-�1
��l,K��mc2�ꍇH��K��[*D�?�g'��n?3N5��@sO^P&�����[�(Y�bv����MM�Ƃ�v�d�v�b�����C�`�b@%3]��Cخ����Gq	��{�F��U�m`0gʲ��̗�Ԙ-o��9��iP	7�WG>�_Q`�/B�C�"akkyVD%a�m���B�y�c�l �T��xm�O~��FSB�+�j/�yW0k��sê�#u����@��z�G8����l��a��c�Xo��)蝱�-���n;E��3���u��x~�Ň@��
��5�ҵ������aG���ΠX�9��I��L��_#�!;N��vf�Ῡ�ۯ��r]�.�K�V:�!�H�=7�|k�X>�OY_�p.�S�]�@Z��1�r�|�1o���`+c�iᆇ|�d�&�QO�r��Z��+�i �c�G?��^��ӕ&Kڢ�~�9d(}�����=x�KP��
_��Ծ���Àޠ���:TF��!��f�
_o~%l��`'p���c����r�}��ɭB���[R?ׯ���蘐�xG_�:e�J��>247�J@*��s��3��2�m��0�o;Ri�f�/���af���Ō���Ԫ͊��{�rT�tm8������h��"���~��m>ܜ�����5	��J��΢zw��l�.�M�X�U�8����i%��A �"h\/D��/|ۓ#(_�E���fh	��r���u�'.��K$��Xg�4��9��B3�V�e���e-Eu��Q[�(�hGk�^��S+�<\���V�f]�/뱇���E�Q�|���ӟ�1�(=���M�I�W<��L��y��]�f���b�n�C��!B����
(d���	{0�� ��ޢ̈́�<����&�RFu{�n�{����[sc>���yI����[��<3��|:��ln�*�9i�4�A_�az�7t�Vĵ`�o�����7��JYπD�`���&�Ə���>f��SG��56��"��|[c�#Z��XYf��`í��.SJ���	VEkD٠M���J�����47*?=,wo�V�ش��x�n�n�m_���+���t��f3��d�L$�������j���{�+�l�9aR���,��o�^�!��'��+�K��O}�'���� H�Ǭ���0^�ل�ݤ��=��B$�j�\	"R��zZ�W��p�џ~�Vni��ϵ���������Ty�|j
In*���rT�D��(��O�N�'?��Â>w�BC%M0�~��9)<��KO�;�p#�&����*K�u\��8��6]�M�^�?���g?��z~)g̕���.���L�C��5E/U��C�'�gϵJem#�v���c���4���	��unhq[w�s��M��p�_�qQ��n����l���3wш�6iO\�N7-��u��fޱK3(ݍ,�paY�g"��R�9|n�FC����
�Vg�;�b�]0�6S��f��oqN66���'�/2�nE� ����@�m(c�$-�U�\<�? �ğ#��~�R�v��e������VS)�ɨ��>�_�ปO��ه�(�5[S�x����*�$���#�P�O�^���m�o�ũk��%�\)^D�h�A]_�s/Ik���&ARKN�Z��.yy�;�uV��V��{����I�s�PE�
�B���uhrr�]s�!�x�C�/ɱ��(	����L�I�0�� �wv�P���\_O�ٴn��ܓ4��/�`M�}�3S�"����h*���Dy��^� ;�*p�ύkj��02��*'�>�J��� �!�L�f(��րd	8[0�⧍�ي9�c�,�f�/V�K>H��c+�Z_{p�K�FϠ�ս���+z���eic*�`3�`�@���#v���}knٺ'���jF~�Z�`��n�0��ێ#��a�r"�Jݘv������g����� �_?�y���K �@���2?ù��*GO�k���L7��{�"Ԟ���J_*a���<$�>�&/��5��a�����v�X#�1-�%�#�J�,	ٞa>�uK'�_�*%%��S-�3��Da�@����q19��ka���nS�Z�����X;���{%	���odf4�b8<!J�A2٪.�c�<e��{�6ա������r7��~�l��y2��n�a �'�Դ�e�f-��:d�sG�Qgd5y�E�r?㔊Z�y-vG��/��!H��}Դ��0B�ϴ+r��H�}`�A��2/�� ?t<�xw"�,{(Jr�e@����_�N��m?�VNɤ�^�ym�[,�,A���pZ�^\�_j�T�{=��!G��k/��G��;�[Ti��d���&�k�<-$[���(کx#���h�p��� �3��\#�d햆�hNV��W����b�����+W�����Ѽ�du��tm��6�� O�:�J��:�ҩ���N|��K�3���9�,�!b!��O5ǣS�R�be&]q%�ڨ�t��p�jy����������{^z=���N���7����I�|V��c�M��Q��q���NA�Sx�5�����0��^�f��Y��ܯ<��9A���bOZ��%lzz�~ǐ��&&��;\�0K��ֶz���,_�̈́Sy�v��	���%��W�`y55RZ�����b�.ѥT4p�ҋ�靫��W$��%Y�u�0��������N�&��!�r6w��k8��ŵ�TV�'mYvQ��D�f2��i���_:���Y��Xi��Y`F���Si7Z�n���ju�\Y<iߦn3w�RC�	�)��x�������L�@%s�CFV铤�H�&)�eydV�FC�Iu�'�]��İΠ|��vp$��7���t���9��#���y�'~h@�$�Fuo����Tt�r̍��!V�Lo�䶍5L�ϋ�
?�#XNe��1�g��(�������:��z�sY��3HF緣���X��8{P�����B f�$(���(�m���bd`�0��`V�+WdbH���{4W,����=7}-pk��'kD�f�;;��m k��X�+1�%�~!� �BZM
���C��>�qVWc�W�d�<�Ɨ䣲n[(�ǆD��̴��<�/c��<E8�f��>X">������>�z�������1��&��5,P-{6���+���k�29R�9�z�yǟ?õ�F_��?8�>�^I�<k>�C�;rT9�vc�abLH�O�[�������n/�*wZL &z�:\�/z_�MeH����$,[�z�/u9K�q��L�xø�H��F��%����n�^���! Վ�"�J���D/+.Z+}Ɖw�Myզ�{�ۊ�#f�@M ��������������E{?W��9�\dg	y���s豒���WI82���~䵁W�6�:��Ue��,f���=�}$F�E�0��h�����,�3iv�?�e�8�Ƃz(�Cuhtǒ##IX�{r~���ʻ�]�(�W�*�}��|�p��)�l/,߬j�_��0�*`3���^z����d��������y}
�t�ozt���z.KW�(�_�u�۔3��n�l]�|pE<C�J��L��mUU0��o��q)BZ-ݥ0�\���\4���!\����N�C��s
¨��]h*.2�sϬ&��y�@�z*�yF�q�����������zGEScc[rcz0�_'��[����~U�hL�?�jr.FoY�uY bM���Q{ո�$��Z<P��M�.2�v�=�Ig�&��kY���ط�u�i_�y��]�ԑ�f����[5�dby5I1����<����0�<Ҷ��VR}�T��m�W]�J��d8Wy�H���'�1��^�
j Q��� d/�t����En�е8��tĚ�o&1OL�W�L^�A��
�\ī��(�����vpW���^w8<��2�{�ܟ��n�!KodU�z�iG��ʨ�Mq.�I��˿�dx%uz{�,�.��c��d��%`��}{��&M���?��ǚ�څnEnY��ʊ��7�Lw�+Z��M� 0x�+��q��+��FF�W�/�������u_ ���J�����+,���?�3b&�n����]3t�Sj��ca�8"���䨳Z��㊂)��X��pV���P�����a���ٴ*ك�
[�����
N,~h&�U�gds)���Q���z[\ �!��V�3�f]�R���/���Q���9�_�I�H��m7���0/���i=�<1���1l�Α�$"Vu F�t����+ǥVo�]���#�O���#��ށA0wUB9ى7l��̯#�����ʩ�T�Й�3��3��o�y#-��e�Z�S7�>�6H�z�}>��׃V�❧�j3�˵;wu��yێ�L��@����^�2��K�-	��O��H&[c���Z����Y�M��W�K��-K�p{��]PH�P�=�O�8��?��čіٶ1z�|����N��+�쑡��@�U����y�Ci����¬�l�Vc��$J"��U�2�!�;�LS-�y��R�I@8�J� �x��������]� 8��;�\�U�ȍ�&Y������_���s�Sv����,�;��� �D���o4&���\��i�͵3�L��r6ݣ� ���R��.��+�,�gx�`��܁s��p��-c�Ƞ2���������0�����I�HJ�0� Ȓ�`Ԉ��G�JSQ���]ޠz)ĉ[�0���A�·t׵��/a�Yv�מ�^�@��r�M�����Y�'��zXΟ��<�J�q�1��'jy�FQ�-�c�o�������V����ΡJ��	^��@z�,��Zu��CLd�	����"��ؑ�����n����D�����
�T5�z1����.|M�����SwEA�" �)�G�LzSu�f�:A]tt:x�E��6OO��i�a�#.�vW�-b�_��!���Ë���0�	)s�R<\tv��@k�v��w�=���:̲�3��L���>�ߩ;u���Tn*�O7̗<��]�݊4
T�'�y��m1dC8���eg10[*����C����Xv?���xև��H� ���,��C��2��'����[<l,��.�N_�"8��R��N
�ͤ��$�o�x�tD�aK�}`C�̤.u����U��1�3�j`ߨu�v��7��[��m<�M�m>�'���v�:��$�ml��D��E����R`�e��C?$���kQ��$���q�^��K-W�p�xV���n>٩n:\[�������^���W:�擸/����L�Y�e^RVꊬc���S��f��A�o�)���j*���8A%���&zOk%�x�w�ܡ�和�`��ra=0�	Y.6�+q�ضT��=���Y'M��;w��q �&6�l|X������4�x�*+x������b�" ��04��6��ę		g�R�$���H�LS��KO&qݱ'�j.���K�������'_���:�g���0��H��	������i�#��8B�f�<O�Ù�o�C+-$�ЃDx _3�;�Iu\jtǍ� 8�}ӠHҏ��5)�>VǫYi�"��@y-0����������h�RRY���*�����S�	@&6!�?B%���Y�C3 ���Y��#����B�g�Kk�g�e����P�Z�5md�s��
*&!Y�F��ݝl�3]��w�d$|ǃ[!B+�б/t٪��3*���,<N����{�~�ͤ6)O`>�2����M�E��NLf%~��X�ANQ�C�Hz��F�Dq����Z�wdȂ����R]�D��לa��8i>�k�(��)9�����3���D��}M���ɒ�ܩ,x7~2��|g�_S���n���(ov�*H��[��^Ù��B��_��/{x�hU{���o�"�7��
L(	����]kt���k���*X���VXݠ���BC]�Ig�ÜX{j.�Lr���H*�8
�R_d�����?6�֏5 M%�C��J�f#m��N�VXZޙ��j:�[$�D��X5�N?T	?=<ͬO�2�1����ǡ�̐��9�82++�W��g^B���!(��Cɠ��0���YQ�h�=TW�:Fp��<Y�6	���-�Gnvܒ�:@d%�)����H�t���������H�#A۝2�i$����Hq�f��K�t��B�j�wfְ���Ljd�0��3cOU�)ۀ�Y��34�<0q(?e@����B����8�4R�D,ع�Py~@�*�_}���ɦ)�y@]^S[��G{��Tx�E�zI'����Q�첋��׼/�ۦ}�t�~�)nM����>�=�:;9=�5�o��5��/*Z����`ub,�����Lč�;�v�j�h49%��b���Fg��@�YpE��٠�P�Y�ԕ�g�]���4�C�̮�V&��߶� EY�F�d���H�N>"���F'2^n��~�v�}�U�]2� ��bG-�E�~���B5/6���m�e��eI ��5��7�6Q@X��o<�7���3�)y�@Ϩ��pBW����!`n�<cJ�?��2�V�/o=���2�Fz� ����U�?������Ky��������%��k�`G��t$�>��C0��ڭ�@�t��t��\�{��X����;s�S#U2��p��:5U\�1��sm�*��~�^Y��A X�)`��K�mފ3d���[���y����a��#���?J��ۃ���� ��
W�%�Bֿ����1�>`��\K+�;�m���R=>�4u� �/46]�~�h1}<�x�\(�o�~fBJ%R� �?�E������[�2��9�� ��هL D*v�q���2iqs�ZbxF�)�[�c�e]�3K��	�*9W��g��_��Eǜ�J)�ja,�)���0�-T�e���Tc{'�b���b�9s"���8�n~ԑ��(&)����GN[ <pbk���"�B�ly2��iJ�w�\��@�o�@:j~�F.E_�n����H�=Z넌��=&��$�]��X�[�H��(Z���7]=�����3��&׭b��i!��{Q�Q�E����Q�8��Od�G�LUJ�/X�M_-����S�A�j�8�d)<A
��"H��U?��9�n/w�kcN|!n[3�Ĺ)Q㚋��� J3u�O�rlkyjp�J*ҝH�/�*��R��z	+�s��{�sz2�-�G#�S~}^�4Y`�nf�L�ϗk�]�D1;����N�o^�R�
��;_
iu�љWB=�Qt;_n�5�&�u��45zk�I<�ng��$���3
AbȭcG�K,�&OF
(�5܀#���9%d�&	͟�ϧL��փv:ծ�q"�[�t����O�F�;N�����u<V��k!�6�@���k۾W[�nE���R�M}l�j�a�*�a!{6v5J�z��3N��(�#F���C�G�F-������/��S�_UCܒ�w8;�\�9tf���T�c�ʉ=�����=%�3W�grF��n��)�A���5R�R$Y޺��"�!��@�F�I��W��ڏ�ֱ����ɢw���
km���q�������00,�x�j�j!m>֤�����̾j�1�W 3��3j���Po�Q�B�l�(�60I��jf	��k(�k�r������)X�K�I�ns���^Ϧm!
|־D�<P5��`-H��{� �7%4[\���5�����,~�+��Y�nR�Wό�Y�����F���b�=Y����C+ס���Kv���'�	��܄�_7Y
K[&�pGa0F~��W�j�|;a�)�G�)/6z���=-�Yϣ��b���5�,��*���ÿ��Hj��w��T��ksVLtH��r[��q�H�X ��s��hVE��!���R��A� ����^���qЫ<:#�s!H�K�@>>Mj`��/�ÿ�ן^`l�ͫO3C])����k�U�v�y��e�X��>�e��������Â(�${�t�eY��)�;���P�O��B;�*�!�r'╖qE�����w���A�	(�����'�����?��c�1}6Z �Qɤ�~�}�T0�+F"\��0��{e��ߢMȉ<��d��F����x��~�S�P��o�IM}<I%���Av���c(�X�1/g<���CG����Y����/���{�-����܊�$�ǵcx :�����FNg�?�&в�4��[J!��]���k��S�~��o���|�z4�'�j\76�K��GP4C�6�3���I^A�C�3X(�:p��+ߜ!T���l��B�ˈ��r��OWԚ���7����XS��xʻ��#�AQ4�E!]4m� :�7�<���j�6�	�-�'�N�]�m	<bTR}�]��Oॶ˷�1ֈ��Q 0�~�!�{����U�v�וV��)�f��q5ү������~s7���N�/`��K)|��<[�Lx;+ShQ/�2!��[�l�Q7_UV9ш���˪1�%T�!�J�������(;�/_D-�.u�'�F^oG%�n�	i�?#��~v]���<*nsAS�v�ع�$���&��%�5=&Q�]�3֯�_���� "?�ٔLuR�:�b���l�r����=�>X�]O$I(�5��<FS�pU��?�uP��: 0��tB@�����N�bG��ÐA6�_X|�M��x,�!�짖`5�Ed���U}��B���&�4KG�v�J��^�Ԗ�#v��8��S��<<&"x���솼��)6	���Oa����"�� m�mT�������9�у|z�w�ʲ����0�$�m�����)p-�c����ç;������E
���:��:d��?��6���Np��|��e��~�.t�1�Ğ�^�c�v�Y���8ې���>�!��dZ7pxi̶6�B�s�2�?����ʪb��&Xg��N̐���7�BIWⳇS��O�q�B �Q��J1�&��WJ��ޤr�y�<���y@��]�7=�)�< ����������P_"��a#`E���D�`��DE.�s�$:��Q!����»�GzP�Qvx�D'<�ɿ(#�y�u�x0/�$�m����㐘��%���P��_A�.\G�ӭ�Fp�S�3n��}��w����[w���빮���̋��뻪$C��9� �v�?M��vm�N�;�UZ/�A5�(�����@�K ���<4*u���� 3D�X����6�;(�<�����jT}:��(3��"��I������V�����Qa_��������z?,�1���Ҟ������"@)�ee�^H��/�.�����b��e�ꅁ�,�-"=y�ΒB/-7϶Th*X�~��y�F�\!j�>�ȁ�J!��Q:��6� ;�$j]��U�/OZ@�.�ћ�
�!Q�;�,�<:��cY<���QTi��{<O�Ur�N��a���^� �V�o>�oV�4�+��(7y��BSR/T����I�\xF��A}��9$�>�P�W�	�v���5�B�Sa,71v�~�B1̅����P�>dI�4�E��u�=/l@��dǒ��vr՜���v�P��ẁ�6�o/�X�����Q��}��D�/�Tk>x<������	�c�ټ�w��vI�b3�3���]�\�ׇ�7\���f�Kc
_m�/��Y��N�[/4*ˌ��,b��?B�.�2b1E��n����䍰��\Oc̘�79M�r��BN��$p�,l���N��I!=�� -+�v��;z`�L5�jcH�ͯ�&�ROnGF�c\�^�K�Q�-Է�v{���H��2M�O���Y��y9�
M�Z<rDa z���W�?� �@8XmǌE�t�Ѝ0)|]w������ߨ0����@�Ԑp@IE���ْ$\�U�Ĕ�{�s���*9?�E.�3�z�2߀�lV����,����3#h۩҉y��$�c��nL�~�;`L��K���d�g���x �&���1��ho������	�;_��Ѧ9�jGɜ2�L����NaQ�4wVf��`
�ʖ[sK��ZG�k��H/F����� �ӟGt�����OK}鏪�w�qɿʪ�h@��↉��CϹ�]/��i砓��"��8�ь�nӚ]��x&W�(���. ̻'�����L�l@�F��� VbTUF?�[5�/��8$Y�򪳇~W&/�`�b�1Jj��qB)���fsw ��
E����R#r�~�������S�u���72mCNUDˍ�����	Ǖ��cZ�}��t<:4����z��ښ"�\ו�:wn~����}dJ[���L�Xn�-(�B٪WU�&IE��W���uh�S�(2Q	��.�-�y������d�����yJ=���2x�BL��Y��a(�W^]��$4��<�����nR�A�wp���mC�WI8y��(���_℃�J��� ��~�u3�{������u3,Cr8_�|=Y)�vA�#�yuBh�/pi�/���_����Ȳܕ5=̹�-�d�$s��Mj>����F<d��荣UF<��~��~p�^M�^v�!�J�i�x�OC���Zhv��8�'�� coq�4�V������H�O{U8���:���V��?+'.�v�#sp�)�vk�^�����^-�����z`��D8���X��[�덥z�s�(g�f�n�����"��&1�K�5-q��C����1�=X���R����OsT��@4�DA&C�.kG�K�%u�*a�Jl�Z��}(|����o�/o\	 ��#�d��T3����*�����&|�=o�A�`[8���4J���EaS҇U:�ȡ `����
���!ҕa�pK�QT3�{`<���ж�;f�����[��9.��`�?��N���/�lAt2���V�I���oE�
U]��a���_���)ǽ�b����?�֤8Pڤ|�-*-�q�8g�g��&�ř��-�T�5�MA����LK=ש��7��o9aicN&�߬n[G��i�JU��5ϙ&����V��z��0~���
��av[@��^���`�ι�ٰ��[m���W��%�^�����dc8RZ��@���ti��MR<Ǥ�������ꣶ�2"�6�Bj�u���k�quOB�㺂H�l� {��+�N�m�M �`ʸ����pqqEU~#j����)CM�[!���?�&�B1�Q*�[�\�hH�+Z��é]i�Y�/��8�T���.�u�IMy��"D��2JU�)��񋇁��z{Ź"2j9V���`�/��̞�{.�|T�Õ�u#^�~ ��������ri�#�������ew������g�c�L�>'l��%�p�g�2q7t�OG|D:li�D�7�I?:W%�Q�\����BoU~)V�F�������5��t��F��7��b�.�l�V�Im�A�w�}�<�W��7�ҚZKܬu����l�e|�R�S��]�w�������&�4Gv����p�Y����������u!!��)������(�٭p�O�S��Ǵ*��MX�� ��.��xć����nV��5�
��%MI&��a0b�Ty8�p2����aZ^�O���S���V��'!�u�:ҡ�qh?8 ;�!����Q8��κ��MX�ڌGz�)/�����{`]Q�R� ]t�X͂,#g'���s9A���3����;��|U�C�c��W�p�
�a�G�tA�X{��M���G�����N� _��]~���r<�J�}�艹J雛��ɹ��h���偑D~��ww��#��k����:�M��d��_240_��o��IސD=ªn*D3�:1;�<=�17"&�(f�	�8�y���t�,����d,qE�v�fA�����*��� )��2Bw�-��.Ќ���(���#IhiR^��w��� '�pl���Ƿ��D��2������E\�"Ǎ~� 9�i�؆z�E�?�n}2��������R�6:J�@ (0:E�nt��0��f��V�cO��Ȼ�\�	��������k��n?�A	sp��|�8�O���dD8�g<e�[P�Ҽ�l"�� �7>�,��Ҽ��w;G9���^.v�P���ϔ��?)�§���~�͝7L�S����G�8�B���̄��q�&~����9��`U\�d;�A�RZsE��]��-Oيi�ի@Lzo2�k�S�&%wJ��q~�Ҕ"��6a�x��s>�'%��Ϩ������(1�u���b�}_mUJ��Mo[�dA����򎫡�ǟ���Q��ս"��tڥo��>�O�?��Ox1P�Z�e���Of4��ŗ������J�Zw�\�!���If���Y���XV�':E��w��nH�LL:�ǴT�RJ�߶[�Fst�m�al��R�h��h�����;��FWy��^�>3�7�������z��C	)Dr@$���g������/�4%�삶�u�����6H���Rv�;ņcC�"��J3�T�|����vrZҾPv@����Ŗj�;(��I&�|յ���ݨ��K���ׯ��c��pg��%r,2[�/<�/��YWG|A��8�z�M	n3[��"sM��Ch�X�2�\��@G��+M�T07���#t�f�ϳ�?X�.F��|�ת�	��Eb{��᤾][���q��������7E�.���m��񬢢E��c~(�gB�[��yf�g٢�b��<<aZ�l�"��$O�{ͬ;E��M���@��6QQ4���'Ҷ�t�as�8d�@�}vP��&%�vk˒(����4��R��~�1�d��(������(���%OBN_�/\�d�?̡˅̶pI����������E��5���={�����F(5iF���൘.m��rB�-]5A����l'�K�����'�?�W���a5�	a�4�A�攃��*:6^�G���Ԥ����^\�3��3\����[WG}��"JRq�p�7aP��TS�X�{
1Թݔ��&%�lz~ ��TJگ����{�����L] ����a1�R���N�h��~/�<R��y�o��`���Q��ޗ�ψ����"���^��[��?2j��R��ލд���Q�����\"�O��C5��|Z9zV�v/����Y�[\�ζ�!QT}^"���h$jC��ӹyњ�b0H�Sʝz^�o궍P��}����Wq�:9��5a��~����ZulxoY��RU� ޼���m��B2P��B��M����n���)3
V�i��t�N� D�'Y�v?ȁ<J8�7��9A�����]�y���7�K�������7+bQ���m�8[�2��� �V�7}���S���p��&���	�n���)����J/6N��Xڦ����{[�ȥ�1n%MG�츯��Gإ�1�>R��6�vjV1��J�n�cm!I���ť&I��3�7>���[�7�w`��k�(�n�O�e؏�t� 8���}M,�&��` }@��B������g��P���-�?�%oo�	ٖ�M��Y�%F}�zJ:"'⃃�L�֐�~$m��BB�s-s�>h��e?m�ݔ��Fi�C�P�W�w������J�=� .���;΂Զ�~��Y{Z�G/�t��?[�8�lh���n *X�ihun��ƺVzʔ')�U쩏h�៴1x�0�1uKv+�B�sT��h�\G T�Q���t���I�Umx���870��Į�H�G��n,[��:s��e�"Nn�L`��@έ��Q�>3����p��40i{|R8��W�(C^�F�HX�g+�� �������gA�Ṷ)�g��v5�����9�0!�J�}��;5��Y��Fd˨뮓�Dn�(@ШT���۶����T»�>��(��`�4���Bj��¸ɖ�ߟ�X�b��H5�P��b@<��0A+���%�e:7�/Jp,�j���Py�/x�"�A���T;���`B0��v�A�>:e>ڞ��a3��s^��A��M6�y6\���c�jb~Kލ�Tx��bw���ނ��P��ߏ�J�_�L�P�j���:�����*	a���v��2���횦��P��.Z�Bl$��?l`�G'K�1��Ⴍb́fJ�`3�ަ�#��A/fM5��#͆��T����X(�Es`�e�����Oq8�[�޶y�W���:Ͽ��l��*%�t}}��&�;l�<��Le�9��F*ac>׸x�Q"���5t`!���&���P�;C�`K]���*�_��(g��7�-��αiͮZW�B^��e֊§�Ge9��w�i�l�/IK��e`��I�O~-�h��E@� ��8ݣ!4 qr1���0���`�^��s�|;�=G�c��h�Fo/t=�d�*M�߀����dR�<%qtX�T���B�yZ��g�p��m5d��y�G�ny>�m[ ­x�XKI詾���	vY�A����G��W�{I{;��GY�&�7L)u�`B��률�eA2�k���f������g��w���O?�kJ ��OZ0K-Yh�v�
�T���wd�k����d�6��)�6���0�\!3@7����?�*��]���:�po�Z�����q���{ʐ��� @�/�Mzg�+��ϩbD��[�������6=�̧?�JZO����QQH�:��ҋ�d	�!�$j��wu���d�:On�+)��M]�ˇ`��LECV�e)$*��_�\�mC�M5�ٜ"�S��l�6� mZv(wӼ�\ΐ:8��@���y����nJMT��
�$R1�^)T����T}�H�!5���K�Q�g�v��t;��[tdOt7_L&7.)ƻI
O�YP��`3 �\eV<���%8��;���S4�2wA������ܗ6�`Д���]����ЧU����v�o8�RU�]�<۵�C��9/�Ys����'f��⇲��O2G��͹����F2���৾rČ#�![	դ�2��Nj�}�C�K�mt�xD�#��v�.�'�"��M�kd�%�s����V_�'O �veO�X�.A*��Ҥ��Ï�Z�;T#�����J&����H"�vO�>��{agW��ם���w�xnO��M��i�H�����|r�Ҝ�e���(D)W�7H�޹*�@�������t5�N��8�=W(�ۑ-'�n�����Ɉ!�d��$g̟�K�H�+�yQ]���X�[��w~{adfk�)��v�3].�mb�u�%�O�;HD��+W>yk�H�c�0%�xx+��lY�>�Д(X�[�P��u6�~�H��3���(�gEC��q�����IZ�L-B��bL"�⯂h-�e�D�DC���l�B�3N�u��R)�����*����u�����Z��O�m��0�N�IiLHc󺆕`a�Q�F��+`CM>9F�v�Vj)6[l��J�<���I�k�b���1��wHR����_��gO��{���۶p�H81^|#�V����Q�������V@�dJ�S\�Z-��j�!x���[5ڶ�B?��Cp��{��m�f�g�`+A@$��������q�h�a6od��x��(����2�`�I��F�� .��c�Bd/
���Ѐ�}d����YX2x61���Ygɂ�|
�*s��3�������ȷ�S�"M/I��D����5��۬q��6Z{-���Z?�����2�_�?X5�t�� :X��g`-�.PM
ާ�9���1C*$oNX�um]t��3�J��ރh%�:�u	�5�ly�l����zQ>�ܼ�� (�E�O��t�|�6����9к#[X�p	e5n���FC��=H9�`�et|��~����Vz�\�6�{��@c+yi�z�Y\�}����?�����I�?��V�"�����e�����n`��������>�>��6�"�^�g��M�	�̐ŧ�/]�;O��\������+?_B�1׌�xB\eߊ/)�Я���k�R̬���E/��`A	m�l��ƐG<�lm���o�QO�|������
@��qB��I�ɛ�F��㵁,��N��G [)4���:�ⴒ�����_��]=����HF��j��˸�T�cz�|�{�"!�um����v���1*e@\y�A��'���m�t���X��C�ߐڱϼ�
�#���k ��~�a�`�|A��Q�����z�fy,���j5_u��B�7��Xu���a�����ԃ����C�BS����aA_���� �k��ݿX��[�̡}��~��)�u/ke�҅65".��/�з!�;�8z� B]��Bn��&�P3dH��!�U�#ue�=<
������cf9ym\��*o��j������rydew�N1;��6'��j�������Z=�3=wE���D!Su�t�_�3�Ԛ+�C�>�+�_�n�L q�h�������b�e�mMn9h�`�I������~oY}��"�L�?��_��AC���V�z>o��h�Td�a�c�H9���塏�����j���o n�E��ׄ���WܹaP��}�6��ގF	�A�;F ����>�t5�KL���*B��[��k�>kY�����'������;p˚�XO�HR���k�V�C�u�Ѝ�ӏ&�e�f�/�}( #Lg�
v��GT3	�=��=�K�e��?.����3W%}A���0�=)�E�L�T)����=��_E<0�W�c�c�)|g���\p��iAު%K��LV���u���X�F3�+#��=����y���_�qo�[�&/��f>`G�H?�P	��呍n�VpL���9��RM�|R�E��[��p,��������7~#�6rc�2���n[@�Xv������V�ɏ� "	gh���l"��$�Y�eB��r.��tW���lʥ]LY�:0�W��pq���y�[k:���|�9�r�]u�nd��q�G$��<�tE��Ǯ�C�	�gF��j�����wZ����K>$�o��Yp`o7]�����R�~Σ�i�.��J%�ȹ«5M	ls�M�ټ�>��"a!�V�Ll�#���W�x/�QA#u���<|���P�*M�b9����֐V�b�їf>Nu��@�Vh��&��$��2v�q*w}�{�]�:���]S�;��Z+���
��J��݋�0�iFY�Ӗ.�ٷ؄�<��ɧCi��ޯ���s�u҃��N:Y@��y����is�/�X�m�5�*ط��)сR����kB�❂�uo(��:i!횄�)�/�j,i2�4+�	�����! ̱�w���]]�
��{�F�ӷD��3�ճ�A��X�S
��{x���Ǔ�,���9�R� �3�4g�m�����8�9�hY��1^)�o]1�1�����8�Db��g��{=�	��p�QejX��SO�+����ɣD�i���*�3��-h�9�����u�[Ni��M9p�jfU��8k�(�HRZ�� �+�i��N���,�����S�>��\�F�yI�� 
��&�N�m5b0JN!$���S��$�$�̾8Nl9�C~\P�\�T1����_��Y?X��"�DA&`b��*�J��&�&�^�q�u@1j���[�j������VJ�������o���
��7������r�0a��솷3�~�KW���wrEK��H�o"��'Bv.@`,�PX�n`����x�wA�asf�(N3(��L����� �f�6G��[h�����mg��	�=J�k�G/w�P�lƬ�����G�..ɮ���B�fWgvh�pپ��B���d� x+h��-ҾVj��"c����E��!I��Q">~
I��3��H��}M�i[�wn�܉�X��/��p��������I��9��I�����v�;�>竰�x�߆]��[!L��x����:�kI$G�̐�Y|��7T5��!���3�����s������2�N�▀�7�b�4:�����n���V�o��
i��~ ��|걚4�=�D�=�Sp��)i��Ž�R����(A�H��r#��-��*��Y�	]�b����z�'(xB�_�'c֮�4e�%�!��16�	x��{?'�+Bu�c�ٰ'WO��
7ov���(J�X�O�SQ2SX$:��|"���@h��*��a�p�}� _��{20�&LՁB��<!�� ��a��Yn]�q����n�ϐ���H&�}�lic�u���A��^<v Vb��u��X�C�y�����?�5�@#)����l~��F��n��@<]N�����&��w�8@�W�\F���
w��V'tF�6��,��|:���8����W�k�����0_nv<����No��'й>��Sg�4�Th[p�1��*M\nJ&�N���."�7N1�T.;�#��<���A��\v�Z0
O6M\���~����*́i)���-&�_bd�}c����+���gv�Y����\3���;��_l
�qb����ZC�_��Ɇ�du62|�����m�����e����ǱxP��9�xjn��s,׿���C���� R����}~Y�Mdzi"�'z�etL��#�te���G�k~�JCM��H��7��[����E�/��Y�h���C���Jͯ�5ߘ`'<��್̓�?�Ne����W����<���y�ͷzŨ�l��LL&j�<I����Uj8WV�:�M�ۊ�3�T���j�KJr.%~r[��l$����\%���Oc�"DU=����lnܘU����$���������$�h�ϰ���H<S9�UE���K'�U�	�[gYzy�*ƓP�D��T� ��r�	��`�]ä APu���Vgr<8��̟w��Oܟv(	D��#�R" I�G"CA'*F����1������?��c�,'-}@���HM�����~d��N?]�?\^y �)0ku�5�c,����8Sw&�!��!�"��0��{+��[\�M9�y�����j���\Q?dk��,�C=~nbg��@��8Y��Н�;�̎�D@���Z��UȻ�N��9;H�r7(��D�+P��-�v8��	n3Q�$i�aL�N}��n�����>JRS�pg!3Ʋ�M3�ݽ_N� �>���?%ۺ�Myd w����?�E����!E�7�V���)k�Z��:KԽ���3��x��k������&�(Kl$�R�l�Scle����`^d�qQ�۫KTLL�jnl[��E��Խ�2��>�kʷiF���)�H̆X�rg�?����<���96�\�����p��&w�վ��,��d�o�)� 	G҈,�=P�����J��^w yf������q��������e[���5=u�0��>~����㹖u?���f��J;Kxԙ�����)���6���硡p����f�ED�v���M/��5Hs��.z�"�5�����ϳ�hۢ�&�/�;�Q+g�5<�x���{k��S�^�M���MMY-�k�z��<�j����!�<�7��e� O����е/i�1���l��H�8���ں1Y܉�e���i�e��aƩDܚ�rw�~1��ӫN:�60����l�j]�M�!)��'�ƥ�}����`�}�%+��>�k��L	X�$�aM[���"Tt�7/2�I�{��g*P�u���Ÿ��=í�ʕ�(~�U���>k~��V$�Ѕ���.İ�D
/m��Zu\���n�#��)hM�
�kR�@{�Xyo�w��-�_� ��QRo����0�xT�p|��%F��}^E��������7G��_�cuX2�s��O��-�@�x��R�钃���|g��-���ƙo;z��E;�pf�Kj�R��H�a�m��4�u��i����+�l�Y�sonA�bU��-�DA������o(��%+�:dv�7���~�u�P�D���;�p���������R��X��Vxc���I��t־�j�1��!��6�ϰQ�.!-�x~y�f	A{�.���}|��b�ٽs�↲) ?C0B�}��C�0�|cl(�3����[�qEܱs6r溼o�����,�$� ����6���FF��Xj�gt͕	�\�h8�[[����;�R���%d,����	,L�JI�I����rj�f]H۪�;Y8�B���*wU�tC��*�J����:�d���vع66n��L��G	��`�_�d\�QR#<�tl���j(�=`O���U�FH���x�;j���kd�U�__�	�&�ݮƪuxLeg�D8N�>���b$�� q�V�J�&��1O[�每���K�~��L�csR�+���S���M밶����Qel^��q&���O�?X& (|�\ݰ=�.:��_-r6�/΁�M� �m�SBӽ�\2q�Ea�_Aw����(�=�-B=Y�$+�U���������{�J���ӱiJ)�tN�ٌ���8�)d�6��)S�}t����E"n�1�n3��g4�Z��r���'2#|x���nq�����*��B�~�s�F��T�ωX��2�+����8G(ތ:�.��3U�����g/lُ:����o���+uo�7��8��ԗg�y.���Kۻd�>�����=���!z��C�D��^E�e9z����Cl�K��ۦ�{�T�Yeu�ur�������rA�����B�V)[�~�#����=`:l�c���F$��k�����->Y��Fi��&n9qÿ��n���T�)M0�L��������>���;��;,H%�1s��m��-�d�@�v�҅�xN�\�P��|5�׸���V�aNG�)��ۦ��t���Om����w�����ПN�j����.z��Ӧ#��
:ﶕ����I6�36�N7i�Y���Z_�����.�7�x��O2S%#���[a��<?첳�W�Sr"�����`�ًmI#`�^Ԟ���Gh��k�3�fӝQ�W���ܸ9>{����'E� 6"����`���Մ�:�7)�Itz�ǔ��^<��Aa�B�u_1Ma�X�iv��Xu��P��J`�,:�m��!�o�"��}����p�o�. :	�&�J��q��W��G�:�1��kD���eM�td���\�-��8��'po�����Z�{|r;�I_��Y�;�]ȏ̞�|��U�
l5G�*�I�ޔW�>�5�L�)vG���0[)���1�#d9����5�<)�y.hnR4���cP�V�*:5"^ȚQ'��~�yD�u�޺֐x��ƻlaՕ|���b��`��.��Xݢ��v��˧20,r�G	T�Y@����l��C��ˣ�%����u��{𷔬lq2�%_�L1���Q��r�e�u� �����^3��n�z"�*�zH�C̏��!�$g���!�_��"��u
7��
	)v��Q��>`����Dsi-�QnSiA(�K��)�n��I�g�Vot[�p��<��{ʾ���X ��yJ��7a5A��r��WN��ish[0�+
���Y�9�۲��ꛌp���(|^��z� {��Θ�`��|e�7G��{���o���:/:�k$-�n��fb�ۉQ��2Ҟ���c�Қ���`v��1�*~؅)6Ò�C�x�p������<�L�K����/����Ē��b�O͑�C�]#����&�:AdvﺭU�NB�����3���v��{:�TT�N7��"���&���(ҙt���ɟ���\Ԥ�����VW	�n�ͯ�#ι�eY5#�1�B��Ai"��U��O��������B7[`�9�3*N��(�ZA"����۽�����h�炼ſ�ƿ�C���ϩ		��A��`�VŁY���
3�;?�E:*O��q9��K�o�ƻ�jB��V^u�\����I�t�~D��&h��4&ai�8_sdV�]+yL+��U�#~P8��Ɨ�꣟��i(e��  �?�ݧ�������v�����D,�� �j�\�&�J�Z������ZLq�x��a1��_��WW/��2Gy�q�w�35K����W���qg��B���]/Vp8�:3S :b���y9������=Z��Θ��Ğ��y�IE�bg+����An���4`+���U]���>~E��o)�臖lƨ�<	W�b�5"A�+W9ܺKM0j^��݅bz�D������T�<a�z��d��z3�Avq�=%{�
B�ü�>�7GY��_Ȇ��d��{�;�WEm�:p���'�p��a;���+��X�H�<�{L����+:�o�W�,G*	?'
v1}�6s=�[���H���U�O?�YL���Z=�q�1�J�,z�6F�o��o,���Lk�&/���z	�:���,���s�_�P�Y.��3�f͌W�s+v+u(Ã�˰1��7p���6+�A��u��Z;m�ȩ�!g�I�+Xa�a����!�r/�O^���M�ſc�?cGgeh�a��;
ߨMOqx��腑��a�>�S��������g���d̎��#�`'*����܇P�Դ9R� ��ǀ���2�	�Ft��Ҋ�;��QP�يq��_��)���-I�o�mz\{Lqd�z|Y�oݢ�v�EQ6��h�I�a
�4W���)�7T��t���;�m#l*��`us{