------------------------------------------------------------------------
----
---- This file has been generated the 2020/07/30 - 12:16:26.
---- This file can be used with modelsim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 4.2.1.0.
---- DRM VERSION 4.2.1.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect key_block
Vx7RMC+3yHKOu2C12wDYa9KYj0kaM4JurOZLvC/V7VkTF32Sez+zfW6Exwuejr+cC5T/wc3zenpn
oQ4Jc8N5cC2ImP60pD06QVQeqxuD8330XXSjDXp8dwhpwWK0ecITe2veockxsXFM4Ntp8YSGpso/
Nqp3m2SQvMbIIVcxJbE=

`protect encoding=(enctype="base64", line_length=76, bytes=869344)
`protect data_method="aes128-cbc"
`protect data_block
Wve3N7ulhMIrh9yUhcLBEpSWTz3dS/4kTjD4JrPsUg5r4yqEeWo+ohNUfLLcpe7kc1wa5MKSSOD+
wd3rfnjHCXfW/mqUKOjAxKiTvHFnBZedYC83uZYSHJmlQNaepg44kuS2cmbSGUby9FcvA7Be3iBA
6dFvsY65YW4wQgj0hQh56ZTiA24VwhaY6ak14yj4v0293mW12DX7RXUjjVj5yUXpcuPZxZBnr0y+
AGBMf/8CZKMnLifzopOZiFYG9ztlqrB5zO6l/g+cEfH1CNTKZP4/AKlCOM0/hFwuAbQ5MRvaG7Jh
aJBeu4iqDgg18boggVE13IV5EpHXLMqUA1Sdya+zHgekcWgRRjsrmSmpRvPqmt1VZKhQj2QCuQuC
xgI0uUvkvRvKj04P1u0OrLcTlYMGLMrrS8vjGE4pewhShZNt/lKlslXWdG+J3QdLJMhQT9REnOWd
9xDDu9UB2/EcJS4/a3nlVaBauYai8Crnk3ToOp9iz1+GUHLMJ7BVvVA1zuDdb97ioouvkTqw4dU0
LHWDxn6+N8zqXbvcnTXIX5/eKraMikGCUCaDVhSXR0rofCapRIF5PI0bEDuVLL1OzktkWZVkfFoW
b+h7SFAwU/+JkrAis7dsYSoVK/V3DxXbNxXwsduKIbGCJwnReATH1ZlOl3OaqFpELqEwfhwd+bCx
0qQnJNI9WJhu2M6brT1MUCfkzVI/7dSmwef8JLg8imp+yGOJMlUuCt8FXOMXsGNM1daPkKW0fNzN
0k5FfrbuvfH6Nc4N+8oM3xap0S5nk1AE04ufW6bTExuX1GVxfVnjvaHdASHd1XBMmWGAL9J7Vo4s
U4T25T2bG/VIfumLCLnhLNgoPBflN1CGWEvbb6f1pw97q6RHVSncTn9DG1E5PAsMhM35LyzllWOl
ftShiR5TOGTPfkLEcl+fc/3DOTfoORN5muVICtWt5ZmuEoW6afIJxZIGAAPLY8r8I7wI4XXMZ5MU
qbAPxGH5f0DEN4zxP+9R6U3W13bBINCIQVE1pgbZDAf3ht4Kkeq9hLOL0Yswq/VxP6jBtXrravDc
My0ZEY29+8D5pNv5TzDbg+ucXutI/Rw3v0Pj1NkRKZn7K2J5lLcIGISxZMkMke/FWSKSmtCnsPO/
BheScmSAxm7HaIdcSI0yvPX9zjJQB4JpUicLZ0g+7P/8uLN6f9cTGgFrbQZjehjMO5cYSZst/oPE
hMgU4D4EgeQaFi56vYl6//5IqThN8GE0cTQyz7qLgrXWbtQAtSMJF+Vs9HVIG0c/w+Q4ux6caYJ7
QRluJ2pZCuyQc5n9IDs9laSTjDkQ5PDSdnxY1e217LByKB23kpqXmJy69z3C61Wsmu9ZlVJCB6LF
eT9nYK6SrkzqVDjZdVkYg/lJGr167F1A+UgJzJecq/x9AjyFkcO4rT356FMcXtJnj0kVt8xIgP/Q
D37cs+759ReXwFpVzzHHyq06Z9aHP+HTJOAP6TqKDdf2bbt5I1cjEEQXW9bAvCW5YuplGQMpnzgw
0cwT6ssDM69uuEncDJE1QDJmghcoCAwMj7Iw1zyyOLBlIyq+0OPspaNK+A8WfjeGyoU8gp2PpRBG
2wgpX35lsTpInTYrSgeFZrg3Gz5SnNFFjnQ6q6DXNsT4C90ySnHlfsiXN5/zl2DpnrvE0SuMaA5f
6kuj+ydsnavJNdSDQCgG7u3ILdFOjhIZBADAJ2F9Dikp8vVG8awNpOWumPluUJSo/LoJlxJpm0Bq
jqJkwSAZ9zjyF7WyP0xOB1njFVDd8p62elL270/tCpZvIJKY09kUJmP3brNJfEo5jZhBYSjwC5vc
/Fj/1r6nVnLLvEBfxCwf37Z7UxLSM7XsBUPnu17v5tkuVkxRi/85fba5ztH89km1qOGfjQEJ6wzz
FxraDmxVf6Gv+W0+9zai+/EMByR+GtkroYIW5JcRXN60TyciIPX156PljwgzIu4PSkNHVpWONW8s
5ecX7oKHkYJHC1zjxNNlqoNutXvju23bUfW/2fe0v2xSMQpuGc/tQLbRHRS4SXitWAiQYvcGUw8c
hoq933G5aftc5yNF0+UwN7qPgYtlTtmAXznDZ5wo7Mprc7+aCdSvjw+JERzAcBex9X1vpR/XqzWg
KZgcbfCh6QMxgbeFLsoMQbsi8G21VwXw9ZIsO9x5UIryF7A7GYFJRcg5393cNrysT39d2MCE1Exz
ZitmAjOACNE1Zi+L/VuBf9nqjdkqitBDAeUH+Ethh0r+VTfNePQLJHDWIv5zJAp+/+TNHIQxMtV3
xCNV9RU53zMvZRuojzOGttDOZrs2b69AV9UIrgnwdcvsjxgmEOnuo1dUmAd3NqsnC9n/luJ2ttdu
aKjZuRVdOCqqPr6z/WCI3TYUT3+rBRF34tRqKdOxiKdBUxL4xBtV5bHr9I4+IMpdI8ntA6vK4E1Z
KfEMOqY6jLpsoXuD0MApXgFiK0Cya+rRLeNAdxOM4aSzVglvzo7jxakmsZD4IA36iAtr0BIPOD2c
5EDEBIFGCrOOE1WrWvtH8pauzQ8ZlQuxZHhrkrcmT1NKOzSeSLczpt8uMXeNoxoYSmAqyhx6Rafg
oWwVO4AfyB99UR4KyydHQ/SkMImT9XSqM3DkbjT8xysiUk4ZnOCy0pkDw+W2QV/mAU71dqyW+RCE
HIvDlKdoUP9QwBcaAAsskRgVoP17ZuSP3yEYslB2IE8hH7ZcEihCJ0JZAXy1J9HFXw+b5QwYXKlv
o3g3Apgsd8Wo9SvKhrism8zLklmB+mDtrTarZrK32V1DAj4cpsT4GNbonBGTSDtLpmzvnNHBBeQN
0R8Rh5mUfEVixpo5jkj/GDuG5aAUai3TNo/Z3vQ+LwtNoeFn/S7DekoPhfjZ4latLJmq6fgLsHFX
3QO9mkH+0gnKeanyyv8dqX1MTNYlSULHfN1BJM1qk+nOlgupFOTpZeid+Oiwg/eTxaCaH3XTOP8h
CAV9GjUPpJZKdXZojMcci2J2Ltl1psHKZIumiIvHVLkz/x2qPsyAk42elfloyBzIh0AfsA3gAdeJ
FoXvxanI0X3QGI1DQRIZ/4bj35boL3N+ReYi6Niuc48ZIRDQCLJ2XCiB/oVYayRtbTmdNHC3qX/V
U/IE5cZZJkfrtf9OYO8zV3eC99wHkjpIeGbinRPN+esRJ+7/tIRvNqoPlxpOBfyhj6eB8UZGilFY
yBVL3eW7w5/3FHrs5qEzmEqN9Lb9PzRaR+REyYW4IIw2JDYE2hrUSY17ANAGU/sG+51+A1ZCQYbc
9SeS7N++tOtOChNngjH3c3+a9ZRV2zBz8Okhk/K4H4GrPTxsxe9v00e0pZcgOrsi5p/Mbv/efrz8
d3ZmFhZ5B7DR0RTOTi8objVjpLgcJGwIH/bs5EThF6YFapdm7U9kUkq2uasQZnFFT9X1vugyrg38
tGvudZEUMnBPcSNIhHu5dbVNEuY+uXsyccBQa7qGvmgYiAvoco8HF4v7Qk75o0cqn0v7wpbzndEC
LvgVooshAF+DuHTr2aXKK0HQw3LyudPkSv8wJwaiaBgjhbJsiOtOgd17swGnUUolqpUcHbefF19V
trGsr9qUkxP+Gn1cKZwzzgq7W3B0HEPUcnxFcP72dQlYUc/9ZFfi4VaNeonZDi7G5abdgUNv8Bwn
8E4f/Km4DDPSddX+vlMLWCiZerTe83E1Taz6Evza9IFyueKbqc9NPSsujv91jpfBFxy3cyduOf3c
q64qF4v3oOjcYXyIorElwQEBiY1YNN5FRxOovLRniT/FMrxErQCp57UisR+I+/8AAPTWbrG2r5ad
Gf+SurrPrjv22Bs0g4oOBC40LQyL1DdQHAm38Lp4IJikSSXgXm0BbGpR+4csXVo6QCepHIKTKgmD
PRxdAEmhtQIhmxG+KgfvJ8DeYaycVjGeb1T17blTKPcRGRfKFobYjgyA2JqdG9X+KPrMzZ+rx4og
xWjeWonHC4ai/7HRcPOxaH79luLmET9xAkBCkS/f6TzDa7TyprQnNWcNapO81e/icWPNTWMc2F37
n3x7giIhFzT0QEy1TVDvVfSMATE5rCzkGZ5MYW++b1rawkNaIlevl0CwgOQzP7hQvJVDRz2p+m4N
UPR+SLn/jFmx4DJiokX9LoeqEBUjHFYdinFCozVwgzt1hWMOs3hwb2gT5Vo+7xuGeVu9jgBBiyXw
N0mSGcwpMx4zfXEumv+qVriFybqe9wn8Ht6FXy2Fe2K5rm3P+l8pItXC3G3Dlrwmm1cmHr609YYH
wQ/U4yu8aG97Hw7IS49yLyE8t8e0hSAliV75UdEavj3ywsphWBh54rzYF5UPZZ8K57eTHsR2emrt
euxV2MXAg7m4ItyRAYUF6cczwjZz2mOWErclLWZmK+9p09NGtzaZkPBF+j5YPuaa0aucpRa3xOZg
7GpU66/5pBuploJgf/6rDuzGo8S4Rpb/D4FkMKOGzXIWjcEFXB4wfOI3l0w/DBreuMIPS0DvD81n
BveLePPJnzo6OZ9IDz5xmvj+4U/ogzwBrzckWLs2UJBM+2WxTkHY1VFQTsQ9yfLOZadaeTLCeGkH
EzKer1funOuPUcu0OD9weFTDwY8e2eIZ5huIbExEbp2hKiijhzlDvjVdB2hSvbzUZzppnTzTyH0/
Yvta6J1OKroY7du57dQKDkCX1idVgCPghDRpkatmX7rehwnahDCXedfwXMzVpE6kIxXYJg0bYqh3
p/4HWxMAd9pKsVqdDPpuJRAKqMzplGcb7hX5Lpqn8+8GFV5UoqLF98rICh1x0HM9l9o8McWcbAtm
u943cUVOJf6cmr9iEtr0fbrdpRmAFkr8YQtcWGaETMAV6WkgaR/sHX2wTVkDKs11FI702LiGlcnh
4sODCANba7kG5M3WmabBrbeUtodyOj5AoOFWv60J0wvUYtfj7dN3iem123mc15jtjEr3/UX2zwuL
iUfhTcMWGhE0r/utvOQ9rAA1/ZJ1z8POkynONn0EWRZKSjs2UwpJZvrVAuV/NXCa5/1q+7Y668wy
djwQXNv44AC20wVlCbZj50mxwYuJOMjCR+bUJjo6mmIGsJd3Lpj3N1ep81A5sllzSpNN7b51gh7X
1hEhRT/u27b4srozA26t5L0OhR3uOT+ew+GH0xryISbQAHIyP/sqF8lgLqPz5ht4WdylEQETm4mU
jL/GVNRUzPN86E8HLaUKdsKgN4A1+waXdWDhof4RJJuolHU9N4eeHaqRxtqeyPJd4BXOyCz1TZ75
HD+PtCwphs2XQDIYj02n/JkaINC7M84WWT9HXImVJ9K/+nsj+yPbDJRsfRNrGvQVCyl4T2BcfHnq
sM0a34JMcOsU40CzlQq/ShwtQqilfh7MnL3TjMr0Rjz/wv1UoC/6IRayICn2kPW7pMYd3+TFEeCF
lIWNcIP4qmumk2BdFUS6xtZ6QXd7se7OWu4F/2ai8A34Tvl3xVHiCO8rlzTjYpfCcLi720gF7bLH
1lo/AUPjd7ikUEJqIg8MhlLsbou4ImuzNaAD6q2/9Aipo+6Vn7DGHAcUaqILjjH0WyyrCUX1Nx0f
JMrRRD7mLpQ6HtXkFbe+wzB+ZwyT9S6wMa0S+zBnQgkinjpea1NYZDRVFSJ2KebYqjL1mxnOBy/N
G10w1tcjRTiRnTmSyTlEp0brNH6eqt4Ryf4x8TPgEGJ//DEubnxzhphC/ES+b2Zch/pXd4JvU0Pz
owyIyb+Ul/vNOaX8NPYbJ5QL0mB6OJsC3iK1++f0IlWJgLXQm4yzhHdnhNlY1yrfmu4ibbfE0/DC
RehR739BseDdol4TCr6F+kDPvuvCfkQIIFdy4LaZF+AFtgb/42PH1HiD3xAg93tRZxT31taTERD+
PBdmW+xSZLjzgc1s6SbLPdFZNJUajXfaoANM9cynygOkg3Zn0jTnart4V+X3q8DtaM9dDARb8wke
Bb+poQBCqNpvvZHBaMxO5hGDFYqkSuAIzyz+g2UZ9x2i3AHXJZ4CS5lRebWbQQP3OuB0MGI6ztu9
e1sq4LW8cgHUzolKi5rfgy+cPFD8pfcm9fVDMrHhNuXOv5s1R1XEorPeOG+l/I0xS5bpVR84ZOrZ
dzvZ8HiacyIUbl2T6TmmOnb0B+nRTvwY6VFGhW43vKrmVd2YtxhVxsx+xUSEtAb9hcLuSx/ohYtf
kHAQ2kaoOOsJ4qfb1RzYQeVz/OHYyhTJHJbTe7JGKQAuFbDMf+mCXB+dIoFk+86ZsjVBNar5cwcS
s/Q1/vWYD0Tafs5URYXxSV6lcFK+3Vik//ZhD+0elzF7ajzKngo4IFQdcN2YuGXlfYC3B8QAEmVV
QVX8zMU2E5ZvK6tQQYWhMdKUz+iqiPfAIV81DzxyzuSc3dsY+y8a8KnTnN9FlYYvsn++pAp1QSvz
pKFPoXsDOnX+eTVdReE3wO1KHtpJj7TyKmym1A2ZKOcCU5zB8rsTks1NqLxEhUodmW8HAuJMWGAg
ZuV2TIAg9M5NiKHZH8hJ6dyVM+Zr3GVGob+vAfj8Q7masPzGfpOtUjgN86pnFR/CLL3A36kOFRHb
TO7mH5zGtlX49FQrLDKSG1DVGLtF5HSOqG0WVNahtss8NIamIz0mrmNE1SpHC+1SwpDLzoR2wVOC
ipNE2WrfXZSgfZZSccxtzHo6DK42PXl47Uv7xDJellYzIItEgrhZbbFJRNETsJ2P7C0am0JZwCGQ
V2O1nrYG6vJ4PI8aTvA45ZkhCEAEGoNhpsgeKv3kxkqlTwSUMEblSAkTGauUfOCcKXGS8pVnGSrc
/1jXJlWsnmckwmA1TonyV/OxPFsT0hSPHNb/W9j+RWR7jN5U30EnnpI/O2WAPLyDAky7QQWkdhl4
q6HcVztO4ertwZyynpdy8n+eG7xm+5pzqkYtL2fzZxxJev/A4Bhy9ab5el9fMKn0MUY9Qz3IUFHu
2NAcPDbXmpAKxqJsG8Md2NZf68njAGsTodUmS5zYOAsvp4HxsK2V4XW5tl+JsSTkJdhJ18LSxYrk
575hiBgIVVSl6px2qer5wPHWowhHFWTCEiaXq7UWNLWH+cKa9hNQGZzstYdGNI6ZEUk17iRnPLgS
lVh+h3I9T3RMJjMeerVBbQ1s8gP/3LB0NoHJURgQbt1bZ0sAgm8wsopOlLQFACbmlBBoYLTDy3MF
KYR0yxG5HqGRISwO0DxTZkV/0A+lyUnSxVAbuPnWYnWoibElfgYz2sgAIgSB8cPedMy/BiycOJFR
YN24HaZcFbTZSy2GfAK+8GF5C+m/edP+4ZqfR1morwOw9R8yDAtrIHGxtHxllnO3XLwgLVAOVWE1
mMxGEFW1KzAYD/5qOOih1mxrE/2fxOrDIqlYXQwPN/sUy1X5tddZjF+uXjLCme+h9Sie12h0QV/1
9DngXDNCL4D7Xftu3QqvkVJzE2VUeQJpNj6eCVPH64H77VccX9B5rxM07XOgVMS5hNxMpbWmNRMG
epWeTgjLlm/6UwE3IVf7mj/wY1814D/Cc6ZupKHmRZ9SsGJZNhMAfqjpLCgSq7nF/OADrVgJC5yQ
zG8HeUqj33ChkRN+yqtPNjcwilVaQjOsq3KVjhkM0RW/7/kbXzcxRQNbG+e6u7f0yuHeNiQHfkIl
ncy+rQXhikE5mtAQk1ME8/OWUvwVElEVeiFqz6iqOFuVG4uwNh6qnmHWgI9Vt9WQgpko8gQk8u+y
16Z04vuL70JUXuaYanuftYUAZ8L8DfQ4BaU28cj8cgCxFqxrFqr2XC66ZCII/NNZ+5GSZGmh+Qmp
6S5mbxUo867cNhU7iBYW5phXblm8XEXnrP7hjK6O4bmC8ou5PbptxX+4trSLbOdxgOezMJv+CFfm
J12enrRW37P6iiK0YyZhrBSe7XUjRr09SG49F08/wCVPyFXIJSP+dv+WWlc7IOAPJxpzU7BiJgXB
4l8pBwo/nVQj/QXp/3Xt91RqbWtZp9SfKbDbVyeyYh/IcD7QpHDzF09S5qk/q3Ow7fjp7iamCNYy
nbkwD7jE+OJn8g8qseUxeRdbSFav5wyjibNInlmsPZOPJBeh8ngeMLpcxo5hY8Y1M74CphsUm0oF
ZRl9smrfq9nX/78DBdPTR7TkR+R3tgWtZLrP+FRHO40IYaogCQpq0MRt7oUI1eNm5vMsREu5OKhj
y89z69DZKeJRN+Nl19FD7/7DvE7rsFjCIZtBn7zkpRmprUwYQZzgKl2jqAd3nS2M6lzZHeyjPumI
Ejm1CNWYc/MJ4uB4odtvDyy+Tlaz+qdX9SgLYl6eBxcV+u7PyIPG31lLf39qKXvpDAro8OXU+jYY
brIVPhfedneTegORA9r+9PLZ2ratIlCQrX17SWHVkPjh4/XmuhzwLVVsEnPJAg5g8N4UNcrvxAI9
I6pNeY5xu5XhD3cKdCXhMA5Sg9c3yRuEZupNvs4tIO1fJEQUaJckEbwv4mgacLyC1HsUXEPcRwGm
LEtWkpKenxL1XV/NwlvRjHlNIj0PzEyCMd3Vj69aq0TSHKxkqinCpJuEPRyKDuNhOZS9hOumzc98
VDUkKrWzfpm3HhILVPbpwupXKmX3VYHPNJsOW50dL7nH0gG6mvf+w5veKASiwGqJO2BwbkUizlg/
Kkzs5p/DVHX1HBaT8imKtEWgRUF0rHIA1UdW8nTsZSyMfXCsz6uJdI8bTia/x2Q6izHG56182WqI
1HIJC8XPRoI3Duq0V1BgoQXtkRgfb+rcOuK+fYF+RvmOOf4RNLy3WOkbmrpYV0EhQR6r1LcfTSsT
4Wce/sZcCV0PY6l0tCIGDTGif9ciRL9vo3fu9bU6yMuufiqXAVc0NtXxj++H4ek3BFifrJOHPy6G
Kg8Kdhm1Cve++nviZ0D8JypIJK42N+Vnuheb6Z45AwXrKSg58aBbP+c7VN2gXmzV/NxzNWYdxTSD
r0AcN9FVkP1co/96oh2ULmz29E0pRIxFDYBVJzWVk3o866BbaSNe0CT6YFPF5V6KEhjfHSGI19ob
3Hx42kNbEbKAEmLZ+Hq+BFRPgUHD2cNStEcSAll/QVNs6tXgb23BZteb8nV2gtInPyWkWWNCr8CN
cvHwbmJfqhrU7T7WJwOAplK7ceMrZXd2+W7Ajzn8s6ztDffa2lOSreVQ13ZpIcZuX6q8ao/7Orvp
fBTDkF0NChj0ncQSNh4uTsm/scqpFpci4KToNvlZDMCMfUW8MUulHSkETbVPqIAjD2BV59kiSwLB
++KW+m4oXvFHs+BxjbMKrgo4xtUkE/n67IRY2FtJXF+O6lEvNOuwL1ZyPi4+Fwn0Vl3+sU0N8APG
8icDeFQMKp2A7sFBuXzQQMX2obljviBPsTHrcmkgQz8W1VLAn1OqHHXMoyEfGYNDyeQc8bsmUyWl
dgRLSY6NB/gxFQ5TmeK+ZYKUt0PWbL7p4Rtz9GhiUHCqmFAmmIpN1RPGkfvys8YQTIYBLzGP5B0/
vM4W+MDts/L+qvyxWGW+fRo+m32DBo63m+spKlXp+ySRFbYYt+mdEOvzXkf54s37bFr6v02XW6ic
uRiclsATXwm1X02B/vx71ejzcHL/c4LZWZMd+JkNfN4eLS2b2fNh2/SAWsJJg3RxzVaq8wZRjloi
RxgxqSmfzW6faxSiBS7mBGBHhuJpf4N9KXUu7FiqW0AO7i/z+QIzfkLFxFuBGcs2QAEsQyKqVpIW
IClwQxGa51Y5oMmGf/GZQvTqnR/bh3uSZOgkqBsfb6JKl+AN+Z5MjndkANGxktCzmYeZVG/cwxgR
U4E/PFTu8dFXaLXBYSjiLe3ScHbZQ1zcbqgUtvK8uKew67PxZz79oM+n77jIPKNNRutK/uozVOvB
nkvMH2KK65KyeYYdgkHt4iZmE4kR8YKePjbZF23ljD1A/p+j/K+8BtAdzJS0pZHM5zkUnOh/HtyJ
6ewahldKqpqJTKs7+lmojEAQGxIZ1Sv0OPbtJnRWLzDcDsPHNYNOtMl2KzQRQdoazU4Qs6zK4kUn
D4C+VppprfTSNPFlw+4WWp/p0whRD4d8KyaArJBRoMcv82izLJg883A+l2PWwG8Fw8hEMj0YnhYN
vfIHa2QSPtN7GiL+yDDutPEO08bflfSGIzMlRnwigojG7nsX/J7XspN82sY5/Q+fHZmhggNgbMr6
bI2eA6dG6PQnBpktR1uHViXHl67/fdFcURKkvPPeKXVExBj2qSpWvIIuK0vZeIeaGPxiVP9qidGi
/bKgXGBdGEjkGFhDQpkOt4OeYcWFHvs6IGLxXA0COCNQCJmhCG4s/mybV0sGuaeZ95lqCIvokSFA
rkrhTtPsMAwQ2PqFzR0wywV+7rwfNU7VMtVPOjL9X7RRKhN/JDNPEIO3Ef47HFeLmzceuvgc3PZt
jOCIiq0vdqhKxh0uuDJcwQ31bhwoJCCL6z8vQo/DxClIgMLCan4GdNQ1gaROQkjrj+vMUt14SNl/
zwpI9vGiNyvs8yCXr3q2Bl1i+GHxv2VFRVTXhVPy0DCyWVA27HJhObazSBKmTcQTi1x5R5ghprl1
PxBDHoZKpjKcA3br6Hj8HdzGjl2kvvtqK1mYvuQzEqEFjK/4/r5SElugafRPxKeaTcqeoPSl0HZ+
QqP4sDkmp65WNCoQ8B7te2ZjmGwNZ0V2JgLpF5SMJJkTgTmASKCN7ueru2cio+1QgXVcyN6oxKch
/GCJBje7g9Ilu1E4p61PdmiPN0YzT8udV+df+X1UM0sXo3JZQSWtbAPJLf5mzPVwjFGLfyHMjaEb
5/BufijOc2FuZpC3OMtz41X0lMupqyIawmcI9Sc6UYoWN/h156rayx/OSZWozovZWoVGCeTAu0xz
eYjcAZWwDh9Y/XQj31d5MYjFjl+oMKCKtRciTgzyXlTWqIJyJhytnSDB3k85oYpDs7wXifSkHmXJ
JnZVFHzKAQ1awPHt+IUJD0xRA8wl/maX5IlS6CtJrpysIaZ/0y/13HLyC+LHItC+ssiw0pZUTyEZ
21YMPUJhqhV8lAG8dDIVFyGgGUysGuKaor/AToNaDtxkmZIOZ1khaO7B1HlBpI9D5Rog0DfMcxEe
FBYonQ2FfmXWCNaLbm62Oy3zFsN3AlCqLTGhvhYCzeWNtYabRiogoxZcX3FBEaCeGgx1allz3ttW
Q+9F0r06VDa8ZH6n8EiBkxl8yk0CgMGS9XKWrFnnM5z1TJtHLzNdK3WvOjPV6UPNePu4OSoE1K8h
t72lyaSYkHUmemW+LhmbByv9yQ4XzOATMhEvQmFsg9QmqCFy5BciuJAU58X+Mumyi1EAizLVqHbV
y5H7KV9NgjBGbIjdApBXuCKa9p6+XyIKzMi8NX4cRJfXQr/cQxWrdP9Q/7AW8TZp6kns8VCgrOil
/L2MobNUMGfl3szoumYYnryAoZcGszNrTqAy3GNigl1llCuiuYhdudGsaRLs8Yp8pwDhixDOVO+M
5ZaD+i+Ku8XNJ68qyCa/orEDj0Nfc6dKdf/DWm+psmWHC/sjfJ9bm4IMP9NGTl/hmPOHdgv2JcQQ
eMvjZnRiuLgmrMNixQ6/8BWk6HOJOV0LiomkUqnx3NRo1hmCNiIJ3yVAmqExWikKcGms7LFP3bUt
wWX4pDEyyaOiw0FXAqd5uBtyOvzsMz6B33DVXZ4yirUcNE/KWS3UhNrpVsPp5B+v/sp/eIRuZkrs
YqCUFOnXqhqBV+Le5IKR+WL7mqGNdoezyjCkm188pn0JiW5ZX1DVod3qE0crEkVkh6yg0GldVN9/
wMLys4WEi8qTC9zudg+WdjX7AkZbI9qmSefAIdrIQCZQlChvh7wHXfCh7EZAvICc4d+L3uGirJro
5XwqGH1VLR3CziU7xQooteS9MEM44P0v5rFwQRDvq/0jPIJ/je15SAUnY/ykWFA+Gzi+V2RkOR/y
c4rU6XEIEW6qzJGj3goNYro57KaPMqSeM3EPPPCrn4WLBNNbI6IjQ9LJs8wEzKExSiSWhr71LDML
5aCZ5S8HevWTa3JExLRoK9DHtWXlKVJGFREPSiefrhVbzp+OZTQ3bsM6lBDeQEuwFhfryHLDH248
FQVeo2o8MBNLEqmnn3sHAcTct0Bu+9iXkmImxoA2bPrIJ2QM/kID0OIb6gLNBVcbyUEJfkaYeaJ4
RQrTysO+O/2eEQVmINtnMvp+k90ChuY1tKpbIzTrTbWiQ5ZMlwp3FPBM6Ggrdllm6azZrM+KMiTS
QW5uUHowEczcb93iboa8JBKsnagFLvgSME6WFeHLVsvLZG3J9H0vBcft078KQygHB6BpYA2zXB1w
YvgX5FA35kcct+YecS9gfVbdrltb1xJD1JDqk5fqqfFfB2Wbk0xXEe1+LPcavjAJWd2vwxgxZsrU
MahnrLZnYwYzceRKnWzO1R1r35LKJMcpNoqEgSMEn+P73ETWV61ydKFdEBWC1ErqRiXyRjcMIF5G
S5T02GzkZctPvrePgwz3qlJXs24kN6WgvxbIZZfs3YO44dvKeaccU4cTEBcr2FafPItoaOUh6fwB
KnRw3k1EPXVyyl64Yfv6o79e6nHqCaQy4UFN4hitpnVEnWpO8IQaC9s2R6FnmvPD9iWevhd3OJPE
SmNP1MRuFEmbygRmx2GI/hEftz4KNjtES0yxfLiedRxNqDV05jdiP4PxR3kwvz/n2MN1tSTf+NB1
3r0jZazlHKWVEVQc2CTL813j7Ldldi+SgFkWlAdfontxi1s8OzZg2G8evb9QK8WLe+0dMyRM44Lf
8bDZoNR9GsRR4ysIcX0b3Buii3ejlzBSDtHfLB9VvMxPaNLW8+C6zT3AISh+AND80TbRBJ+4XlFt
ZlJWGAFcNORgxfbxf8+oydIERkN1zrdQbzuJLaKFk8KGUgIemdjpWAg9Mv/a6UnXK1jS5tv/iBgA
YijylSh4jVwzgzAsuOwS940k05OGxdCMwqrC60pf/G0wV2d646m0g4jULwFJQmlZMnNy/g8YasYB
EobsKeskwVOCg7aMbd+Ah+2YEdfg/dV+ygH7fxlzSsI7co7EFy2RKWgJa/Rsl+1qEQlMP8JE0qZI
kTJgIQkdcvQgeH2Jpoy6wRz4hda1pHNfmmz7+JKxh6lRDgwfyXYp5b1d7vxIocKz3Z59LPrdwlTu
R/hrkiawCX9xKfOiZtEdqT0nvuc0s57q3Q1Uq1EuD4qzQhX/I0Cs+XVnljShK0G7pl9SY/bxs3JE
KLAHNsrA8TC1HKO3tbHA09pgZbn/0EXBMw1r2R7rgtG8LuSkW9TK2f9+PE5DWsVopSdHR+LjZnmO
FoXN6WdZVgqX3BV51rra52EZa1qJnwsfVM7hiyQhGajh70FYYHeKapwjpuAQyhV2Vk+lo+Eradym
z+9CGV7ZNGX8VumyYjaCPGcBEIagdZh/qXSfGx2tYkDyDRGULzp/TCxNFRun6fJJknzqukVpJIEW
ti+tbT0goLf3JhZAiXNUp4Gh3DmaI483GwFSjzWB96TiSWhazO/yxJRNaNI3T0WR22oz1ss6bmAm
iLqMsGLEkvSX8xVWenyNbGsBPCNxrG4q1y4txaoGkXbdvqgbU62IbHZ1K/ZMThiclxjGrOznobIm
U5gau+RWKw7K6Ig8/BwOhqjuDh+Ndr6zoPituedz4z6nq/uT0bhqAAvFV8J0B2AV6gIJh9mPTCUO
5dgTePllHWOm0H/XC3RG6sSgZKoPqTVaNlp3lFTq2w6KCK/J5qzBsMszbvEPdEflI1q56o/hIdfA
NL6E9V3LtR3CqlkQPC48vRJHl+2cUZphh2RnqSUArEkvYF1cYUfC/lw+t/OGSTqYXPOMdCdnlWpM
Ze5zjJ4CGAUEfzDA5CoGV3GkV6J7UdPGU0S5zKVGsHO803gNmdW5VYLf7VbpsZrYBgEm0hrgoURB
iR9GCd9s3ivXVnNeRtA2XcDMfUPEBSfsMvv41LTlm0UuvASj/UG0DTHywrA3uyXq5mIujt+P2aoF
uRsXovQNBo0ecR4JtocMV49BDCR8DZIxMe/s4Z38mEId1H6wB0o54chuLyM/zQNh4ELWI6hHZZdX
T0lp0qcESRY88dvnTcFpfM2ErSUo660OIqhCeG4XzB160eaeG8H8q/S5focoWSMahwk5T3VMldu7
bDpPqX4/Ss1KCZjjTqGam0S6WaviWIE6k8k5DZVA8I/VOcCcxjoIhW2mi08foMBpwE6LhnFyFkuS
ilnzyHdHwNbkbQ2WQlPuPfkRQp4eyK76eheZacH/oK+c8z6N32EGMW5W7o0/uX7WLFC+3VvYjGOS
053Ll6fWJo0Gxy7MBjdn4tYLzSuIjteDwl1Tss8vnZmJKhAJ/oF9HUrQ5TiZm8b212iZXyB+eeTS
1su9LEpxweaopo3E/NQUsjF4VfntLUlPltexs0TOrxgyCLvB7prwE8UPf/+TxLOMKaUM49IH45YY
HtEr9WZa+WvpWc5Sb+OZ+QbUkxkgZKRE/tq7v+vfphJDiQPXWniLXAIWATb6BcmGpTuP/QBwfYIV
ClXHoXCbNpBwwhGw0yrUOnXiqdJhQPqBkn2XfoFYhONB86dRwOUdALBtocJJfFx4kQIfdCU0GsLH
fXxuujnMY4CuCRcy12OKD/gBQfSyVJeIGInqe9QBRDuWflFyQ8KBTQup2Vrrz+peT+2VGMwTmMzz
CAMKOdOmiWU7d4+Nd6ymEKFgGmh3nX2MBt2Y8MZZ4FkuMh1QY02jzi8veu99yEAtYFvQT42ax1nT
kFc0SRQolkqscG8wa2GBRJCGmrwBzBO0j3x2rJ2ogcUmdFdYyjgLp9kBe0fpyuEmtb7MOw+bDUkB
lwFa+0ouj4m/wWcTYnUZTgGeNX9zoCjm61K98yfqSFCuNgLtqt7UGfBkcGaYLSn774Xmzhg/u4z/
k4/xYxFY9nSXj6BITwiTZtvyd0QKHd/T2EAtxAN7YAwuAmUcSt0cF5cEptJFlCTLq8g2hUIP2FSO
30koPtgcn23ArgkQTyTYhrzgVl8Xuc11HBfNu4CSKs+LjFl+HB3brRho8t0FILVgvG+bHQwhlXMJ
LvkjM2xsDPfJtcmGFHPc69BXHPsJDOHvqZ/O8X4TYHH+GPOflrK1AJKZAsNpns8L1c4xURQR23BX
IsRfpMgENb74El5ugSDRfMmzKEXgK9Z6TLgfRVQkU0QNE3/Ormq92D7iKtL09K9T83gvtIkJmO/3
xYgmHkG8nUQBgQesuiTfaliAclViChrnhYMsGa1SWubrcoDPKzFyOlPO32//BZr5jmH8zAWBp29n
hZTC3EbF1XZojliUB9f2ZCExbX/a3TOe7jqJpdZwRbDioebCqCob5BL7Lv/pD9nuBHuLFBl+iZPY
v7KI0xHlbNHDgZoQV8Hta/4MuK7M5TygBeuOBoabr1VDMEZ4MYC6co8l2sqR6rW8gDKJsO+e4ju4
fRJcJzmkDzJhlbffp6aL34LbLC08K71THbmykoR4LiAzYMdu/X8XYVTVntfZNtUV1+1yJ9FTO2TE
X+qiAmZslDjwVsoI2ljwMuTwpZzOQR3YwIhZAg+s8/q9V7wyLqcNwYhgrN7T5atdko3PhO5sIaZI
IHhd42D7e1QEpBdYMlPm38vT+RVODiRZIMyYfuHOUXaYf2R1l2UGrOFbnb5coAzdzxwbIXN58+Lc
XmKYvH2R396De+UwnaKkIRgbXy1y2DuiJKsqIa+ez9sZDoPqZRtx1VdcPQ8/RtoxK9VV8Odkshli
BQA9knV+Vkk+i7vKnYSUzs57/U8TqXO//Hj3KHROJFRlmabDTAc0pc+fcgJ8x1149lGyDUAc6PUG
lOLpNYyeLGpmGVGAXEI20XGHa03vqzWZ77yhFtjdWu7QQHnbWSDNYdplfncG5FpfeEo/IVTN2yER
wyCY8nKjV1XknkDEa3zqkV3gdWU5UfdGVbdnOn8TEJdW++uGelrqoEsAJgjgg4i4OvF+J81P/Jpe
JeC/hcFxGB4bh1HhFJz+FoBkgeNTvlG2YxTzYch8qE4coMZfb406/QJZjahR1DwUhqo1xFHENRhv
voBkZuclvty30/w5Z93uZNM/6slcjvscThDGiCizprvkkoHxX4p8n0KAKX4Z5SOwWc5Upbw/iGqK
vElRecp6a0eViu3xtfdaoOsvFg15LJYwoHky4PqZDVBNjtUDA2fFqdUZ8Lgd1UEjxuowLnOyon9M
HcWespZJj14G2lxkpy8HCNKtpFl22vPoHShY7YJKM635MIY4bYv0D3MzteKORPBbPJbfFPAZ8nIo
9l8+CMwpfF7LDpkULtv6DiYejWZnImvpWTNtOZlcT++GLaxhHERkG5cEnKLYA4tAf2+ZhmglU8gR
yNpJ1RMimMVtnaQDdcWWEs1RgF+BbuML6hiOWM9WGK1uMedbfYTD5eGZ/hzGLV/L21rBizD2Lv7t
vI+r5Vv232nGWAK4QkCAvsNarT/VhLh0nKRO5jUFhEl4fqDZa234ajRVzaSNhd4EGClk9PuvWmp0
sGZA4596ALuXjxnWeilYa0Ml/Q84GIToizo62VsVu708aOy9rBCbxfevFmU3GSkcD9kv5WpajHPt
CeVaqus3zckrlw/8WzAybNQ5NQL4nKdtErizMTg1vaBMkG0Zzd7KDZOL7oyLaBgJBI3Xb+vCtmvf
i+HVZnQyd2Brlsms7KlczT0XplpgOvs7higwM98ywHvWtrGWzdOeBGGjB6njCAicm2EI8coUsJKE
FdEcc/FBSWDeiPbWMYihIaLgfok9nSLcl70cYAcRrdZu9AYyy546HKxQm6oqRuEGE5rneOJB+GhS
u8BISwZ043Myr8IOgHF9/YqRbkKuIL6VcaNWugemw4dFc79ik8X2REly+eH8LR1JOAW3Q5Z1/Rn2
or7FfNebiCBgCc72IV4Of81C99f649F+PuarOt1+uo2d4yXvY3OmQ1qkNJZhE9cGqJGO/AL97kD1
31+mKyb6MGoEdf0yq5jcm9uplL8Hy9tJ9pWnAQ3TS5q8WBtpPdParHqqXySCl/hWHGfuc7/HT8Wn
0wlU50JJWlgr6A6S3mju2Ovw+y81O8TzEwtRukHYcFkm8zvwS6lTIuMsVqxM3gTpB73W/jn4Ybrg
OXHjJffxrAWD4MAt9UeX4BXtqc4OhfBWFROsBd8GUJqebCmSYAdnm/3QVu5ErVLS8FEbAAGKbTnJ
dIVzwf5Wi7CDcB5hlX0mFx9TGIUgQZRxdK2u0Y81+ufF+g757U2BtqRWvzSElwG+XzjS9uf22sdT
5RDOJHFvzPWyNoUDk3Jc/xo+76JnVUFV313rMBBnEZdD4qmZkErj5MzIL2l4COSVEjZpepZqcDfr
AoM/hq/1XAP/LioQoZw7CwjFjGNC5XcrU/DyOVT7Woce/oXB71XW+OBCZ8iIRwMWCRd4lf3eP28P
M3j/S2bA5cgvnRitmpu0azk6Dv29boBefbcMx95m3uqS+ei2SkyfVH/Wocv+v9HLTnifPiptUJQG
58QxiIWrnsvml+kgEx0ABrInByuQtIoAb2ib8hs0ovVo6ggm6r1jbkbODzUiz+m93HKrd+Eec3EZ
EJ454W5B0cz4rcxyjUAqrBPVzGhWwQ2T0CiUQFfn5xNcvAXCNgSPs9h1efa82sxSl8Xv6n8bDA5P
fw1FIJyHW9zGqfDxtF28BhTR6Yx8jdmnnMSqYe1JbpxI10weQ24AzwLoK659sb6Y6otT6VY32SXl
dp1GY5LGJGXMP5sb+XJ/kYQ/wxy5X4Bzzs0UN0Hh9YIHdRpRhQC3ncSkRKl9bLmj8F4k7xVbI4zU
BTCBlPFnvVVM8msafeivcz4/QBgtGqWsFhydDUcxLn7NklHbeLiFbguWEp8BdLHbZQpPiDNCnKOF
QVPSGU3p/WqNDCJkw7clNRSihDQ6Zcf7xmDDcjL84QOQrSiIR/reX/YPVIDFxRyWfPVGSP3kipa1
Od6/qHisz5o3UScx9rlyIzBpSfd9JbXLagJjI8uZu7khEvUSA0vP7swMJrMXk9a3LbKt32wAFpdF
DDs0jFUjC6Us7GNAF3W2FkmGzYLgGT08GqPGc4S2qMuf/BMHCWik15OWpaUpNhCH43gerHpWDP+u
yliy24pGEIYgyempTT5qi6ul41CjMzGB4IwCvs1S6sg2TjL8I44t2pxDDdTKYWlVKUucFzFjBlDX
Q0KTAb+bqeTsqe3Uw0CDFhjvXcP1wXw9qd3ITq6nSgs5rJQQ5+wRTTblQDAX8mISFvqD6SHNNUDe
nerZ9GcRPsoMPfnG4Ex9TOShruRJyQnqnTX0N+FGwymijZXfnkLyJ2Eenjvt9fpkdw9OOJ2OKcDZ
M7+WdV/TUToVN6s6oysplF18k9MSMA6fATHo6u+Nkun9Jy2jCOyezTNakqXSPtZZOGeGOFmk8qBv
dJI4jvZZOy1sNep8whkT/l2lRTgEl4OIF+Ifi35Ve+QqM0gh8du7Y98q/3bZUbxJywe8TZ+y7w+q
ojs/v8U24v6iSkMsAkx8qtUuJbjTPUlCi6R3Pmm1n2Dp2dE+/W4VYPcbN/50iKL9os9d18XgktL/
Y+yRX/UfhpbQF8O7IKbLtqmkIKjw0pFR3LAzGqnvkMY7a1AH4sD2WPDN9NQZJy1rOzJ/B99MjPx7
Vk7y2vi22uSKXNX2VLUdZYtlZ88Efar1JPnd9MT84rwbq0zRMHdAGaLQJGZE+75TZrqXsgVmfC6F
5+Mv9hpQivGJeB0PAlZxbjUhSYjAeCaJllekVJn/msu4ljeT65ylCf+/nQt9Ie8unIilhZPlJVDI
D7kPFRGEDvaePyZcuPbeSTT+aRHZB1jSMn4GRImemrsQty3D8lVSbsR+XBTZ1Ma3nRyiQNKwUWDF
bTNoZJq8NdYp9pHla9E0lwgRSi8K0/iS9kNoykuRLl87ym1vLsX1rrmgYNDrW6X1UoHUN2HQUV3b
Izfd1KGSDEpLHmxA8bwBa2o4TH+9kmWcyEm0zoWWTxxxHY03hOnd4JnRIEnH67ZvocIeK5dH2bQS
swCKiszUksV11soQBWCUcFe7E2+mQ+11Rvt3gysnMQhbw5XvARti1UYx4j+VD+WONnompK1ukA0y
G0rt3rwP3dprn+nyWDWdBj4QAjxUwdhsaXFrQtE8ZyRS3+Rs7h5yHK4vhfPeVfaikwBEbA52UBgK
v3xQDqtiXKtqh7CJNinLqQPTH46aSaqceUOPOz3lTtjHoK9uTcIdm0T1dwilRdAvw/GxM5l3w7yy
06Rlbs1lDdlk7x/6n+rjxzPFq5YPVNCs/0GAEnvTealOngrryqDC2aHM0KBzgdSV4S+gj3r6ueXu
fpvyKQqL9xruDp+xSEmYtmkAXSjYkSm2QSbqjLiFdL9XPiDM3YfgIDJ/kTwEY9sN40Qz3++9o1qZ
T4bJDlBYRDp4cbMR1Xe15yaxRwjHg8RyDKJsdwhJd0KAsGus9oOImNafz4PuyRWpwO+hwtPL8T5z
FR7eHmtJ0kP1YQBwtaXSTtvcCs7BPR60vj9CNLHzxnOgrDiUFydBiQOTkBMtms/TsrdLFI44NOwY
ClexI8/o+s26p76uS+1ThBy7O+5XNtAxoORFaJtzlBjsz9rPac+nkPkkyOerZkcTlR9LRSziVRaC
tZn7PZakSRoDwDZTyrxeCSYqdkFDmQp+8uTObwK/+DqgaYI7YhV5OJTkziG82LsL4jqj16JtL0wu
sYCm9Tq8BRmc+prxN9jpKTf4g/3uFAsmlOSSYe8C5vp/CvewD3kdOuA9ENX6fAW8oT+HdXeKVjZ5
tyOf1PmlTBDThr3/MW/4lU6Cl9hJc4xVbQctMHjBlDEs7UIy0QCwvSoJySmE1sBvv2M1rINFUysb
0zJDbljCIIkE+9vwwsMTGp7MIDQqJv2IhVDUYUzyjS92k2KPBdpef7i4uc88Gi58IC64VNoBkHrC
iWPwUlXAbGBN4boC/PzI2sf0XorAWAqkBV9GviZv41gkOpJ1elgg7bY+tJvZqMEkBq6hJ1+HNqp5
Df1G68rwEnUPGxcU5DtunM6V1HlWoiZw5GRz10eCdjwFAmTHBqlIz/2JzNLr712K8UYkAzHQuef5
XbSYDWkucezd5EcQwGjKQH5r47ELDp8Q9n8oTNX1kKk99HrCsQbI3ExaNjlFMzvi7oD0fA+qwaXo
otrIXKtUEm3ukXmJzXZUdB53z8Y3p3PsT3yt9Muf1EE2A7PEhBZl8P9kygK6hraub62vCmJOXLFv
erwCm13fgTTpC7AxPG1/ecIlgiTI/Y/XjHJhX+tDBXG0fSFEw+uJ04ljva3ToOK/ixLVex26PNzi
BXGVZBN+ZR8ChccdaamwO9qKH2beIwy3P8qzLpTUnXYN+EwxPekDc5uAyHLLg62Hp8v3vjonH64J
9lL2N9Cexp5Jt8zMOIX0f41G9LyNklYrrsFfx7CGvwSezHN/j3xxUuguy5VYpwl6hCm9K/jKyOtD
eB54WdnWdPtKUVNDvJcIZK5UDDLzNYbcOeUbu2Y/7EtiM5nBOK3uSh6fceYcS9PpJghjBoF6XZb9
PSYcUEySRFqTqVQ4VDuulc6invVm5lNOH9VbqylmpPTtsbKt+VNJV10MLpGh99/Y4hpLfFSVRJng
9QFgCPgVwqMS0b6V6qCcR1KjGaZyRdusbHbPhp9NuxNyihGBhfqukL1xRAWgB/cBlLKCLrdZJQG0
LfHZIRin8jQmldojZdnODIkSYQxDV45dByYFZoKDbKUbN3dkyrpxkO0webPNECntJZz2mlVn9Tmc
qU79GobIQvH75Yc+HisnbSAqhmFRUarY5zkyILDz5AixKtHvV3CsheFv1bkupovj0ZKl3uRatdsU
+CEAZmBxOlAQq04qejvchzbzzXDTBXY9MpY/kLIx1zkCxBz3yuHzRW98nFuvEMwqO96WVNtVUUT6
c62TbRJUc7FqbVwpW7ygqMgGrDNqjLMK6s48DAExP1C/cB+SvIuV9mAvSuNOJjZmBAL72Ps3vsC9
LojlimJHy/nN+k0GxmPHrE+KjXAkxU7hXwsZqXW7fTPGBxnnfNqfmUEOJkcRkGETi5W5Qp/68mwk
QCwWIRZDYFI47KG5eIg2lu5DQqwUUG2AZBZV9SaIKDGuJ7wxK7utzsWG5abh8i/jgwUfSvjySmKh
VcnOr4Sw25U+LtRAzidT1XzF6cgxTpgu/DJy0CbBdZkf1ybbCM0LPvMpbdfU7WEGg+01suQqpsmC
H4iCCUke4NzN1ZgZUi9cmnCaFaSfRobEqkedwznwsTukoxW1SD+RKvVC2YDsv0aqRdSgpggCZgFK
CfPdtetMt/Ti4fgJIHzurBrgr/NXHl3UCDKSwLCciD1mhpMfreNpwcoCcEwGaFQv1IIv08lnlRfP
IuiUzwNCt60bnH+njW2TnFjDHh1UTSkO9uhTVUTdqCs1JqyiVR2JFufPvnNgnKZs+r59CF09BYCO
LiOlg83qIBZNxhmohZvcbX74URJ84el7+AZp+WO2jvE3bmogCW1xABPnQ7F4mijSatIctEJDGrH8
ABNZg/IWhiaCFfDeNwsS40zI/iu4BWbtnCHnimHxrjtfWsE56W5sFKc3wPJD8lSQHROYuwHp+9ml
lK0Kv0EnvPqpqG/9sTiav7Qx7mxY47m+JxU0SNoHtnis6YWz8zpk1S1zormvh0MC/w9Zj1o1PDMY
WSPiNYM3tc8E/BXlo+pfqDgP2UCg9NuWdoQYV/aOTPFfg/2UcvcDFsoiSlMa2iV76aVAgDrDypDC
+siI7Lp7BU+Mudmi6o0KAnAZ5jy2fK8UndESCFsr6L9yvVTvIAhbvqLgfx5tr99n3L66uVSTTwek
CYcjg/Cj+eyfJuuu1LxsQPhpGqSIM4l+v9KK0lFZ8+dXeCngSvm96dyIzevSWfGOGm9ey8EXmB2F
mf0owjE5um8qW8QaC9D9u+GnjGvvHTD7Gm9HjLk3qrNKLKyOmS3K3+cCxltlda7+b1Gbk5ziEAnR
/+rbmm0Y90K0SALSC6TytFz3DMsXyqZAFSmYNXqawFvujANqa2nbA13ErXCApwGwzgLlQr5LFXgT
aWp+G9mE7YwMj26LhCqGesHswINjOQVfwYfYCTNPzjWI7s6tMzgibCbOKE9InEkansq/kO77H54g
maa1jKKGN4plDsU8aj8ISHTo/YMMq5IW1YwkRy8tQBolkfrUDz+msNXmXZFabQK2+kBkNBmI8ohQ
OuScJD9ufWSetEYAn6XHGYtuOVRG8R8iAVxwz7c+FodzuKQn/oiilx7gGkJ6LJDLU8rNEzit0uVL
84WtfRJnJJJttZvnXV4teEls58iMU2pWoo8DZszRFzVck9OpiwkyeJHQqo2Mmn3vdU4ZbJlulFSr
ryhU2mwsQ1z9Vg9No5kfa+V5xuIXKvuT02M96GWUcX93J9pnU2bQUPrKHImZclXJl1D+piDcQefu
cQpOx95MT23yjH3hn+414DJd6nZT5iu16l4p5ebnw/lEF+SllM/i96Xu/d7bnR9h0abeRYsGN+7Q
8VBNVBiPAyHE461lOUz8CUiN+Y+2ZzYb38/FfCS6uawdrBtvtSjv1THi4WtOg17ZLLhpClZf8r70
yHj+iLsrRzTvLdX+bEbOK6TL2sTaNdQSFdN9rmdwqVrz5WLAwDvQEPdzLlzqeGkN6J/lR9RU50ff
vKZ+yyiwhuInHMEVeoqgZMhB+A0nCD9iV4oYMqR4Sths1TW1E17xoOZNc1VHqXF790uEYdrNy9T6
1pMzoC59gzwhRIH2AA6woKWne0T2oCmOebMzauYR8uGyEVqho3oCZcYfevlEQRK2owQRwbIt39rB
2ZIOKAVloTalv0axqR7AiecSHh5WI1M2XLkUv4GEplWLtYutf9OI1XtvAp7h28H0Odv6LgJFQX8g
IFblEoyfkpkj5mxLfTnkZfXkfM0hbqzBg6umFnxsePEsAhvj82BLx/EftqdfUUHSYUtXdx71IPgT
BDQrXJMwOoAYpAyvfVqa8Pxb/5PN551OkUSsLGTI0yFNkDcIowV/oxAIbtclLGGo/Ha5ecrtjAdM
gRY2kqyiHQso8X3bw+mxxZVHYQvNIgjiAQlDxijdkysAUXAIYWpVwKdDqHhnRmaxBz+KPnF1Wd9i
4sVCC7EJqSplYAzA+6FmEd5slT0Ioh4Pq4BRSxO/49uASSGYV4MqfBhoB3rUdoTxnqZNL6vHbNrR
7ojnHls6mt0FaThimSCk6I6d/IkSUy1UDNyiE5WjnDHKo5gu4c073FWLO9ynf32D47w0t/Dva21T
QMAAgt3wKGgxFU/b+hOok06VEqHwtrO0AG+UtQsFzre4kEYjS+OF34KDAabroH5TAm/5oUUyLcb/
f/8uQiFSIKjDa8YJP3HUP0TxreusuaQaqQRAYs1Ai1Cj1I1jbajuBgPPAn8Cgr5/dYYqXxjpTaku
5eYNiKn6kANov7Pq5+WX+7HbWTkrMoxrBCkkMW5EPuQlbbtzn+Qo3ZNs0cxE1WSmUpESXSR2XTnJ
mdk5k5sXmb3JadP+UMpL/NLtsmzMRJgAiliqgVA4W90Dr8jp12pFeK4+aLYBf9xBDl8KyD/EWluV
CGYjqbuxhS4vsSl0AXMA9Sa18iT38sKPOWCTc2TXjNhEk4DNxPZPmdlTeE+/ckyhfmWTDUQR2LIf
iA+NeDOPcGi7hkkISiP6s7luHbcc+COQCU0bGrsIl7o3ndxTdm0Z7zFd1P+k3SzynlnAMivHFHj7
/9GELybBwlC40QwGWh0b9pEcT0U9/fY3WNIb5tO0ZaPT7+SZQf3IR3jnLA+CB//K3m0/0VLo7TDR
sUMHl1ybiEZcWM5jj+8uRMyg0jE9QSNJT6e2Q/KP7+8MeqHJsX7h3BL4K8a0NUIQUXwyysx6UZsi
00yScqTtuOtaI8GuT7ktHGD8HYzzZVi/zatCbFd7Z6MZonw3Q7JwWI1smV4DuVa2/4UHEdGQsiQj
aRGhEL3mva4a3xnmuSV2WJJ1x3WfQvTlVRmUAkP4dSdC3+r6S2zF7PUUoJbGQDpn9RMHobX8abgZ
H9OhnJDk6KPi227OuvsSDPiLNdEehvCJVP5JzMSoPdsEYgOSzwKTjdZoIGUKOBbjBROn61CuBHSt
qfmlSbvhuhi8qJ+nIY0JCuV4GQLGeOJ3pqJiW2eKMjXzS/56/NYi5dkH5ypgt2U2L1z69LIDnCp6
Gqx1TJLLaU6HiNB15R5SBb5ZbueHp1wX0okweSsWfY3EHYP9YwzshjH3UtrDHdpVdzO3exs9hakX
jijCI4eIeiRhmmZEQYusW+gVdyowJd4ssV0R68FergT5ZdxlF6vaq05AsXOTAhp6JCrjCZfVmEPK
yeu+Waw2/8imCNkkqbmMVzeyKP4ZhTXoYWQxckCwyBeoVUw3D28WUW7S3AzNlttccetuASl8TpHq
j5U2yNW0r7C9oPprh+STePyJIKdXA/Gh9A37eaFJHN67Ap68EBHFOCntuqF5if2HcRBUOWJXcz/I
cIp77QYU22Rs2wAzVGdYIyQGgrPKgK7kkMPMP6g8UowGiJWHT16uzNXHRL7bZIGI15gGJkGOGOCP
Hn30A7BB21i6tKEvvqXI7S1vf6rf9lQajfY2Ww73mrxy4EYYctLFbSuDAqvQieJw0M8FPO3fMh5b
8X2+m8UcOYQbq/84dvHhivNcr3z3Mo3hEbzj5lmU30hxesXkPC1H9ME7LXLuH0CTgHjOhE6mjYCE
cWv6EFNNr9t0BUcybDzRzKvdP/HmF8O4AxkvLvQIaB0OnDPk7D5NnQiRxm+7hFzierOQIpiOkjE3
uE4AT9eu/IInlwpNfPQRb/Vaf76PwvQUx+8qK3Mk/8xYm5ZaBtMxXuY7Z2nYO8Mw0o2mYWTvlomP
RpH2ZTboBllqZ9oqiOIA03eg9SS6RlK8lP4yFlD40x1n7yQV/yJHBNHWZ74YtG+xRQuYrp0eJV6f
F07isZ++fXG+gBSKSw3Q6jwaB0LNgRvKPnTRreULiv5NWVaA2hUyMMxrxj5iOt91naxL81iB9jfw
MoWT1yoADwfhFp1hYIm9GB2vNGo7ocq+gJ1h+0l26hHRsdc6nDsrpb28WyC2ixqL5zYPrgyyFQcx
MKLiPzIDI4OxR2PvyWD6TQXlqEwaG1EHjDVi3him8DdaRVYDBzPGGxz483eTt2ZsgxFu82CadRGs
udX9vQxYjpUTsh/oJNnCnbIZyvhfEx6xIP4PZqu8x3wrUDvSJMcQvS9NowKT5NR6SC51OwoPYhEA
aGPovmYrIPFUMoqfRSyconHphaQW8vXHW9QiLHYaaongGQwtQEU+JSxfui3RCCuVL8Vsn/D12ZaS
B/PQPPDLHxwmFmJY8yWATEHhLCGfAN23juxixEDgfj3L1Zoc2OL0R2wWvLfWDPnn07QUPZlZhI/o
6hyXa0tXEfQYRHFXzIAhhApygp9T+HCHMwgkd6S5Hpa0UI/JxBSLnyGispu0S6SXP8RYWppmXMo0
zxSk56X1isU+d6Faoxl6+edWAPTjBYeWsae02FaGyj88zYDrxDWXwSwP9D5NYRlgaHAnpfpCvrIF
OsdiY6rpJOlbgc+j7V7SpZKkSkIqSEDFhhRP8uc/H4h1yJv+VIm8M+fi15hSmC7LGu/qMRnSLJa9
UD+rR+RlSBZUDHk75IsW5wTSEhFe+cmWIN53HwWc75NNY4IEAHDoMb/XqtC0czVXOVEY/Jq/MZ+K
T7Z6V1lQj1ukyvVE371w5e4W+FYfg/38G0iUFN9qPca4RdCSd+TPwllCnbIL/ZYXIn0Xv/gfCeHe
PLiz8G+iKcSBMxL3508PSQ7/2kGZIh3ZnYeL6377VVP7TDbbNn5ccdf2d44/Cg7awM1pbkhasIij
jkEYcptf1vOGe1mPFsrI1BFznQuB5Lw/wZoY1reS49cPmNm6YRFASKbFUvnvZ4d35NSrKvwoY9vz
ztBCjevSL8WltGDndrBVIsMXgQmCJhkOHIruzcbi8zGQ2lr9nZF3Uq+Mna2D0c2P0vegav7HAmEw
mZjU4arposzFuhArTdL10MSLBQLL62rLw6kA4AG+ltDVFN1ITrPKiXCQ0UUhvpfmZLIiNKl4NJw4
Zi2l8qII52+wjXMWjR2JDOV9U25CFtQFwZq6BJK6DrOBVpSpRFqjBivwqlt+Z/yIYyboG+nQl7hu
ckhjqxCyVM7vnV5kTVnzQll0PqO2pkfUzvNhTG/WooAa/g3k2noYKneMF5FE2j3pNVOGFdFD4vBd
GvnlT/vWFqGZpGXGcUJX5sx7ANVw7YXn/OL5ADteLepcUMAP8SB4UgwIonvzEgMORVVUbdkjLwxJ
njCMRoJtv+MnTdvHVceDmRqZ+0h0A1zduTufzJ3/7szrGR/1cMNn63MVBCJcWg6kBjjpj+ioI3Eo
dd80vZpRiwU8+tTJ8d3I8GZpZHTFInVfE2JzuYNPZJVJeyVZFDrNfuNJiDgpujUw1dkY7QNaWQDc
WigmMiNjR8dw57GtKVuyWoBHQsjxtAUQznH5/+sph/4yetfue+nNuuiCRlsfEQI/lsqKy7DKlUlO
K5bSeuHK/db+4oGZyzgdoM9zv1twv7FCCtYy76lK3bMwB7IrCA8ujrN3CRTsH++fC+GIj57r4IJK
oPAe70VYxHvlrX8Ag4PCySqWPUoieyjVkq9q17JxhUaFQzHhczDlSpniFlkCGzmxPqFvmfGHbicV
UGs1bmaSMdfIiqoH55255Ilj4vUPA5+aWGillBj/zRbNY9D3HJ4BsRGz7NMjJrkx3xcYxO/2N5xp
B447oNIVmtkwIKpPc3GYLk+Iz/Gby81HAModdbkN3QxJZjwXODo51lsdAIxaqv524ZdFNbrQTl8N
WEA2W4OfL7UWJzGSgJVV3h8J+Ehf7oDF4lJdwMAxJmBvqlA8B3+XuRGJKP7+dGLdiY7RYQwBD3hB
vmgqwIC2+kyXfdrY9hllYKplWjfWqllT5Eyj1P7vyn5g3UqiA49BowT1wP0vHCNcvVPseEB+Vd1n
boNFQ9Oh8TGD2dm6aw/3KvnlbxoX3xNDd85gqFNx3OO3SDrHNdUGl9llRPrlFMorS1ssbZy5UWc8
wfwrK4Gg1Dp7ovt23VeNYZT13KqXH6CaTbk3g6Ha/4PHQLc5Nmov1ZXwH9h70/5iXRxE9Ob0nrQY
iCVTKlQBX2Woend0qLUg+iLMR8IO5mMBTmGGdImtqIaPdVvdcU+GIWlDIjyG5OubXfVpBHrpLqOR
er0F3I29HUPMrlyNzwIRySnZ8DdP/eb27UPmG9MBPyDmTRcacalJYWR0FWXY5qPw4hqbgpV/XZlw
a00RE0Y1mDq9pwUjt78AnH8W0owwaAqDFO0nZSdwhBNftuKhd0QGPYXONc4lHZy4h+9yUOn0OwgI
gZwCdMbBa6vfNQH1moN9ynKEaWW6sB9IzB1J6M9bN6aqnEaSxLDKZ8RaVemuMT1CtxpOefn0F+P8
db2XtapbkHtGGduiShHiJP/m8vxg3XX+7187aVvQzpEd8VZb5HwTS3PMpTcdcRdqBweyiy5G6xyA
0JNfgFywIKxxEWVJdkdqbVGu2VaWbfFB54lADJSIul/Yh5vg9kmVZP84al75Uc+3KLTASfbHWYL3
inxojFOhX5eL++pKgtMXj0PWS0fTvgZsoUSzR1K6QWHQuAZq2MHQQypfyPvx5AL3MYqvmV1ctrVp
Z3t09lqColZ5ttHSEhhuTXqvDESS/fQHNQc6p2vCGTa2hBx1jdBBC0v2YiwEpR3yn8VOQbKUflXo
ictSw3leH44Z6Jbahtu2aTUf0vwtKCKft6Wp+OYgz/PIyIIN8ef18j5+9xwEi2nnan7iu8/dOgtH
2gEwxW9b6NcS+hIt4ELXMjq0Tm8+/C7LBHUdfUgOWAuj1+0UDarEARodishFcnFz2OnqsIunVj1h
ucGgzq4dpo/QjMXOy0YbBcP3ELTMIPpSSCz9HpTOXMKSlCoMs7PGVhrITq4ejg3tR1j8fruVNOEf
1w0hTjhaoJJrdYpZzD83Clkk3u2R2NXL5Z5rzkXVMPoKm4fOuDRFoVnmK24VYy08jh2zTuPdnwBB
6FDi5d/4DkapBnwfl9imfYTDvVGlwEeNB7bYUtwKrCZlKxfBrYnyyHtUHkglDKs3ZVw1/mvd6Fo/
zkLQm97OlyVAAcl84869qd7dn698H2wMrbrY6bmE14/ekJMnV0vaTYmq8UtDx8N5sBaQUAtzWeao
NtwTTyRRo9nK0KN9DYfDOx7FeFbX5ZBGb+iMkcZ8mLd3Cm7NIdkyOBmrMLqSJC9OpvDu5Z2n0JN/
njocPlMS/CHrqBc2Te/d96Wd7QcV40pxgkHOE1WXliWI9DYXrmQk4Pl9yk3Da+jmj59dzZ7c2/qo
Y40h5MUhW9YtTvyxPtdJVGVqlXvifygtDqR4QPwjJogoTXzA0fiTcA/vXkIvHMjo4gl6T1jOX9gX
X8MWCNae6V9ZqKfsKTB16ViYFnug8APMWOobtM/4tDIqiz4Vm5bKhgXN8kbxxGg5i68gZEEHMgyE
dRhPGRHrkQwWo9LGvL6O1iLZnSTjECe0zsCs66qYtDBq8ZmZm/KCvTGMynynDTZTVLHG5vVbczkE
57tiK6OXUrekrxhtqp4wGEzsk0M7fp3511ciPoXx/ZoUX9Ak2ItFZzrMWTbjIo/W0g1TE6O40LF+
RiWbCjTWAYU6+jTyGHMbayBKV9Bu0IVtbBlsrSxOlobdYj0/2YNyaXntZneAhU+h7bY9yme/zADU
0hstSlB4C57n3wSWOODr6idDobcoA4eFt1PLlT4r26JVsudmoaRmGSdQEKXvdjusLZMPk4eR0sae
Z0dzmfEKLQ2Af5KzLvE0yggBaKenpmedPlgxc+vBRbN4bEbGPXxu/CVcx/P93w08KcGzcIfGBZRp
CgFr6H3ReJpUAkvE06dohLkCuEHyLR/mFDrw9aV99WlQz5usALJl5oo9XhP95+pTheam4Ft7am0b
V0TA9fBU2AbaJ4SlW3cKbfhmpWVchObVbvwMq74Yz+pj40t0HRl0JO0AMEI+0RyLS6mksyPlq+Xt
/pktITyS/hiPmxiR/fbJE6RWAb2U/bweOOc+UsbFR0TiEFNK9rL/1WROkpvAx6qnLyWNrNJ6A6Pg
TfE8WCWBUvt2ii5rSYeOBgTbhs2SngJcWESX9w17K1C87Cwk6ioHnYXbbrZo1pLEeP829aoYO2up
R0xZ9WH418S+9TpVIB5YoI5sESK3HqRTYAQmoK0+kLGrmZbERR2trTHwvwXJxco/WnZlI1pkdX9Y
zK8XUdy7kn6js5ARphxiUL95R+LLZgbBivjTtBTgaR8oHQ9jiFo6tNm7RSEI2ayfVhIN6wfbmxhM
/Ut4ABo3Jsu3q5o3Zywu8oiA/cCl1b0DbK+ofsSpBLUcGcE25PuajxhcVKPj2EMi6FLC24qukKzo
EuI4bh3rGx+h1kO7xpmIuHnYAGFKmVl1Z9EueJ/hkzKWpmHHJG3fCbvLf5i5FGuQztmBBBR/EUUl
NQ8+eKsHWw0JrEaf/qoBUC9X5xN0KBWVrMrwFYwiI5BOLmZwBFBdk3k52LLWCS2x6RD+xfaAw5xu
aj+KQUUpsGhW/zrPUyYWNeM9dKIHMICZt4BDngrnhC7qb8c/NbMDAptLr5vKCYQ+ABNvhCPtqv6x
sgIkz8sjeOI4C+rnMFqW/CAWxuzv+7OJXF+ywOc/q6DMLqg087Udfrb/9NGlEUBCBmMBXAB5Y7MZ
4NMxvjJF2HXq61jddvkBU77b59164PG7EcY/lGwQzdwbN7kvL+MLka8jnCjlUkQD875kzy3sRfPH
Jz+z66HBG0BtJDioJTr7vN6EdcVSsZEKSKhxPbXtlLsRZq1/p50/LgG4RtU8+pzQLAOYy+eYtCi9
OR/q8uWwX/yvgnMM5cJtWBgBM9sjFGWBSuSh1f5Mixz92OkBx2NFMgfdoBT5F6b5Dt4c7IWasNLW
OMCMGoFmkOTZeZ0tgTLScXiH8+4pwKVjdXEnxjMjo5HyrtFth6MhflHfToGWnYuPKpNunTG35ivy
K01cS3o2RmDZyGY9oHqzHn3WUNe51GnTprah+1fvd2Jg7P4/zszifo9T5+4savTp/IQ9zxHh8rSx
OxkSOUWoA22TQSy6eyqJwHdOhizzhSScreeX+I64sq4a61G+TblMRuRpXuy7XUp0SKqnAsTU7cKF
2ocMeYsiu46yuIJRGQMAfmb2mg3atzdEr3YaqEdFLlXTKM0iSPcQU9qoVzJmAQxuSUnJTMKV43zV
dtjd0ylWZ02byWbvW5SdGCn8/2UxXBVUXLjLyzDF6GOp0fI4sta21PEuhLgJfWkO1V+RnLNTLNO1
2ByXFhOrDuQxWf+TdzVLZAjfFaIbha62mk887FGbfxJvCYfY0PS0jCkZDkDUpZ3vjSSCawAq3pEQ
eXBLOKlF0pedUlqaP1XV4H63786WNZnr+eKilm+G3KAT++4jAnzf8/1r+tmzG6IskWL3w9lK7/me
8xEJk0pEqs4kGEt2ftC1jEGBMx69pc6iUPQeqiuf09O7Fv2FDmJE+MMlb9fIJk/fVzUdBLQoGpl0
LKv8ubAXUipZfE4//HxjbzTD/tMPdIXmieVIO3ucQLi8ZhUqaJrn/cFHSa2SWXGwReVBCbaEZELV
Co+7+Xpqt2Wrjnwtr5BflsUx0Ntbj7cuJmSC+xfIf3X2GuPbz9muV1+UirIHCUp07HkbahpxZcK/
ifVGX3tUjg+IUfXKQCbzn2AdDLgkel0ZGW7wyOW1JDitZRD8OMoH/zqZ+rBU1y+/3uRO+9O+Yt51
O+RTd9X70e7nPd/KtMWq+fpHVZDx02stcIyeG+8ue5F+STuHMjayM86ZdCkL5B7XgqZNOV1UZBd0
m8IDER5DWPEMNNmK0Vcva4o9Ne24ko5YlKucpY6CJ/yqhHPRtgWlP7sV4JzpfPvc3Sc4wsaBwsYR
A82HYr+RHlvaQouC5xi8yNiF0l1c9bGUM5PVNyqbOGu1Scy+cvD2MWMSAzrzzOY3UbUSV1abujOO
lZHXZitzo7sdYVT4+X6M5DLr6C6GNfernNrmJ8dw+J/e/otgWfzH5XFH0hfq03qXv8xWPoZCW95L
nLp2oeQzLuoLTKgS/r9ryySe6qW3r0HteC4IE8YuJvNVPo0wIiJFtGYP8RPkjETWq3rWdivLlsz1
JGXfXQnxknA2x1uSCn78+HJ9kix+/k44NG1Ouq4tRigcm5vHn/QPr2XkUzlAue7QTGxR30RVW+LH
ucrxhShkiRNIto+b5fTFNnLDc5Z6o9du7t6/PRqUYHsUbl/xQs5dnCgMlElJ9Yk1ZCg2yfGLMOpC
8vzciarZvkV/24ge22d0bZw4rutS+N62Kr98A27xwDpzYp9Q9dnTvc9/3CHS2FDFBt0p7Kz+yNsx
y9jlUNhJj6l/DZwasAsYeI7pn+el6yemUQFZ9g4zund+pNyfzK8Kv0Cjo9y+gdkkzHVqZbFj8KMy
sSeAM9WYJgAiqmzCgDG7N3VpZi57HWtz8Bbqi+DXe11/skKybuZOLiV1wd9sm4VpFWylKAIruY5f
gpTa2vU663Dw0nvJxkWbKWv5XoEBtHzMNaeFEZcE+lK2I6i0ZNbfo8Ms1mC5wg3tAkqRgfBOW0T8
qs8TDYx34Icl9RfoNOkCNrL5DQ63z0t2AEUMh7OA5vCPfqrP3+lIPMi/pC8wOWkycx7gDPVRwMWF
rVTREYTgP2uNXdhFWr1pT3b2iw5y0Hb8AVTMj+7PX9+zqQKn+31fRw0l8m5up8oJT5usX94IxNDN
FOn1vvGbawzSgxDrW9nbgtKRNsWVZeOo2cJIbH/nn7iMiwH/93uH+qvKPRxu9vGg+PUuAHx2JEq2
oDy4lI+l9djepLIn3YWiPK6sZPNiJwpJKof8vf4s0YmkHFxqKU/v5UpXj6B9GvzJATTMfcjg8L1P
BvOyAsp6tsPy9LxmzBsEpi7XWUa97PqBQYOoMWlA+KOIWK3gWl5i+AO7v/B0N0LHGBFiY/NLpI9W
B7GuaZxAkZtB/1x+p/P8XGgeepbu2YPAS5NsEC+Q3pwDdxw2asI2fnW0stBaAj0k7EZ4jroblr8y
rXUCc7YXQ0Q3dzuFdKTKejPXWH0bcN59Kw0eYq48ivSzfduxXPMLkBM+wg+NBYn7UOo+8mKrVWwj
fJIENd+AadWOfcXxZg1ji5J8jRTkDoXzbWDDSNuA+m17UPbluuvsfyhawbBHqp7hm5aVs613+vs2
B9YbDj+eST7atKdq1MSqm4pAEGVs/Gmu2+p32TwsMkvACj7Qa8kHbe3j7LZ+O8Ov3v2o0pP8Ghh4
gRBStmR8cC398chxUkq7Q5YutXxm1ALqn72b+fhBTBvprFYinW2gJlWoqE9V4uA96My/XDr8rasj
LBRG4lSi9Frg2p6pJjtA6KTjguXo9A2N0PhXTC9YaO26LSrAWj2SfxEjXHzOv/RkJDNP/VoJ7knL
ROf33znvmZkhP9uQu0Yioe/S1onPHY9/hReYFzpMJ6G/d4M878LGFwLxl2WkAGgroNwzSltUYm+l
KNKjFAtLSFktdSJt6kRuYVYY5Nsx9nvHDvMGDGa761bvhklURRfhfA8u1YnDE2UCnE2iuSeCq2ej
6afpYBxO1NuBlRpb5xnCP7IHIZhT8gUXvKOdhb1H+MFnynL8KG6x1VGIZ5seH3TI4GFOBU/Kx5wK
WpN6VYgN61uB1NX/FEhR7fLiRUJL2gsK7G0VwD9Y1sUIMRsnFmanmKufe/DzhrGlrOQkChomtzNf
gmo6lYk3AW/3eWG70GZJhmXdxw/cNsqDZU5iNeo+OY+QfqAfqOaIWWks58YkAc1EC23kiB7Yb0qJ
of5m+BUQ/g1isGRXj6VWzBp+KP3KhZZLW80IhXUNjiLySdfM7KTg4m+CPNK9/uSzY0lLhhBy2Olr
2anoQ/KevNnMfuLIQp+QFZ3/06th73NTrKXybUDBB7ro5aRlABHoPkazpy19bw6ixAsgRNsDjsWe
KFMidcZEY6DmywRBxRxT2NCH7ntxj2+0nxplt0/DH+GvuLlQ4/F5akwlssdLZFdDPZq3pPhlvL9M
s58lh3p7IZb7xCCwG2sTm8kEHgD0GrDDRogEtCsuxOZJ9aHnVNAyvkUfIYaY2XKAbaCbWK5+a3NK
fEghhPJ6TkxVJoZSyfVTfXMOq/jrbFhMHuYmpf9T9BDkoKG8jHlsNIqzzLEkT2VNXPl+X6ONqcfA
gjG3hepj8OIwN39jv48Ic/msqdrm+QDTIpr16Pvy+L6qSxhrAi1rzrmyi3qO80ZAOeNKmNytiPiJ
A2XbDi2DU/QVFjTS7DKc6mSRJCRwfikNab5wg4QFdF+soYKqBIbsGiVMNMfrSgF9K6/rwF6KzE6S
Wd/lP34JKM8s+eWHYbh4gFfSAn9rnp8UL/+VmtzPEumg8J830IHhJ35uLCkb3uBIKTXmKB9fS1Ri
L8qLW/PoyF5Egfd2BiZo++n6SGar+lm7XRaf8A+Cataji3O8gaNpVZm4YWsMHuHJAUB0Cy3e5gqn
Gh8d8yPM23NMkMyx1edayxubwgQ0IABfKKGcVEdYGRkYIbN812T0P49aF0DBkHTqk4ubrTujcrs8
+V6g0ELkocSEZ+kY5+ScmamRCAgVVHLpE3mI1cce8dAM4DW2H1BlK5vwhTtv9LzKHHlFjsQsWf+T
aQ5XZlJhl4rTB3yalzAA2gK7R1wJll4Ggaf+kaWx2KY+iexStO8H/P+VN3g7OaejIv3uz8sONiBs
I60LITzuBKtiDRd8tTFjQhKZY/qCjZ4J286z1zVg/wd28hBiAjpbtutIkxVfCURK+iIDdiLiFvJM
4c4uTS27ATKaMzn3w7yx6oE3FsBkijRK7n01wWTYybSKxpT7RoHwEClhWEiFEUX4ywCwdHyiuIiP
MUJoMgqZcdsy73xl87JRVJJ7Mvx7XhDyOyqCRXbu35j4o3E63eBwVe6IdypWH+lXTuy8MRQZimBi
OTPGGjsHs1jdw1YnEkNJ6nebiOcrOj97FO4ZviV+KrbL5fDQTIt687o5GhwX1rBrXLKZZIPwBUHE
lJk+NcgZ0PjzgAjOeq36vqtVxgQIRfQZLq0//B45lwcm3Kz10h38zEF5Y7r3cLqX2sd9Sv/QzqvG
yvju7m6RXAFWcgMkpowLsw3Xx7oJeMlLTAnoRWAXuh1n5UQCe2170Ofmxc66rZ7UZWmJ8QCIlZPU
DxcpLgn8aQuZR/Eq+/79yILYW17ku59phEV5QfLSZrFw3Q8ptWy1gjlAZ0WDxwkxPJpXifNJFIdi
NvfbAhirOz6kJR5aM1JI72aLos/TvOMP92zT4S94JWm/m5JWbYLkkICoSx093QqPQ5jYRzs+ykGm
oCaUuBLEmy8pXd9dXwUig1s+wimvkVI++AAocnBd0TKZwoGfJ6YRdbtMXG36sXJ53dVaPUmRL/3k
354Q0OF622dc2rxfDyo5nRC0NzOdwlFLYFek1OhHBPCp//CaGe34xj6PuyDrRp6QUoYvIZKRxCqS
hBIqfQkykjcMWOjSXidRV5l0j33M9AclOTc/endzFvatZ6SF1YUgqzGHz9VT+syu2nVzsHpycSOn
s+aUNhxD4Z45tdGccX/wCFswM0NudaxwQ+J/oo4awTqJ1Co3h0nPlKBUzQH+nXlWLkMDKJW4/e1P
ceqgOupLYyMN02mkiOpfgWTGizvzqr9arUhUU+iK6tM9LoT9kt3+1/NO7UKbl986VkiMAjgtsIf6
qTBasKZSSOxtNGUrAMLxbjJvxGZCafwpBf3AfI7J/MRfZ2bfDlIsUPu0TXwSVMTCJUC7bcU1qd+k
tdaw0Ysh+mk0iPJi1ydFJuxiuH3vxOwbC2ikToBOPKGetXw0nRdIjMIn/DNqteQfW0pigRhiAyAW
xH2lSzYYW473/Q7uc6n4sKJ3cqjkPq5RVk4JSRShfOEbwpU1wjf1F4IfTRwadRsTV/DH83J5V50y
kVtkKmfUESIytGfu/lxJrnHYMS0dYK2iBagnR3xmH2vI/yg2PwRYqMaigitiGPt/DGFfxPtUrJDy
hR4zMbsVIRfnnNzmajJg3FFkSD2Db4fNmSDaSD3BERCx4byTu8Upv4OcbO/lDaQjOKxyRBgIqZG+
3Dqh5chcKpeFyXXjgPOAeT5Ixwa2cyNl4aCSvBd09jLMG6VfeEnvdpr0DZNUAvvqgxfb9Xs6BJ4A
mbKJErqFUKUWSLjVEdMdro8oaLf52UPdRWp2v21eWyxS+UHhWKYVAMiZnKQAUkSBbBoqo0YBJ101
05C6hmpyU4FkpZqbarv+H5zyO8EegCFSjdoxAmFRaufNrJSM2a5TJ/d5p6Q9w5jHjPUsOviQZuQE
CVarXEhWJJDgFq2ZJIJ1kFIu33vrRn0H/P4+ZxHQ1TXAXkNfVb6zag2m8tH8lEjIxzJTMhFodwJq
PT3rpVfJ2nD+Oba5//2F+KORC2Y6axDDLguWUDwDxtBJvVJogPyyvcJooT03pK+Kq5T8YPTf4cKI
ZpYJK8N9NYyiTCsBYjimbWmB58vi9PNxPWmUubgUX9CfW55T7XHaymYt5rB7JJVuvY4ccoLFvWq9
bUC3e0hlIvcJMffC6Qy4pBTt4ETiS9qHrUlWZvjiab/p6rZsLfVkP5SaGQgHSckdCtOZCBwkEgAJ
fsvcLOqNu56JWa/zKDvJihsZJi1PCZMVmrzPUEv9LOduWDI8FYF/cq0wotJW6RcnKHZYcernAOtO
PIDgOkYKQlGgIEMPU6+qDR64ssW4yBAnTf6VCPLSyc2UG1ApdgYcxO32uIZ914Me+HRdlpz96wDf
yaydUHw94ytGsTdCUrFiST59R5ob9NdS8pFuAf9OFsGBXsXsVR/wu1Ii10IbN088cr+JToP7pi+S
lC16P65dyYeC6duxxoOvg0ywkRTjz0gT8UnSDnJVloO8YtYO5dj6YIjQgFOkY+ZsHQ/CKrQqMvVJ
8i6MCTGe6o3y/PxlfF1lKuqU21OQQMEYayBK1u5zUB5EFyAvXgKbkog80vA1xZgvV52QI6cSPU/8
Vp3kmypXe5yiBNoXYDIh3mC72n0m6QFvbCW+g+hcxBCnHtm4VgjLQrKRQX0USuGWfz1KSrxkwifW
kUsqL90u3feA4N95T09UDY7DdM9Iv5rWGCLee/24IbQ7BQnz9V20yOcxUabe5mJmisWIKs/L1phg
/7MbB8RRlY1nY/enFdlR7JgGQx34eXh1b+fUmCcwsOVwlIrvdSR02nAtYktW+mudJFLrokZzeXOE
zn10x1vxqOxkhIhHEs36R0iwryMwvpnsdiEtE7o9oRT0CiNbaEfNaLQ8klqBGHrtopm3hX3PCuA4
CPBjqHvpELLkO31n2SQRDBiwpuYL8tnefSrAottv+dv2DZjdx/QvXaj+UEnp+4P51gLpAXy8LJCL
ysU99HLWb7WjnApOFYAK+9WZXc4TUQOTl9RlW9NIZd8vxCvl+/Kjr9GMyaO4TClyRF828EJCfFa/
TKayLcj7wD6RGv3+eaaibVK0RsK7gPLa9T+rdGFtJH8Mi5a1M69qNz61u+5/weM4lZGwT4eOCaBY
YDpRMt8Hawzjvx8u2ZbSCKZ/KU9CfCn5Az3Tw8etfcpGEYUvFAJslUtwF56jf6Et9wVF9Sd2UiKI
jzt3y9oLCna9tzHOeWUGB6+VP6vqF4tMf0oW6t8Qp+RTM9XmWXT30uiNZ433yvnQACcZz1oBNLXG
Pvg91AUGUwuECvmjfeHYCvFBsbnESdETt98e4KAQDSxpHUH2y4Dy4J/hIttMeOlZtm9NxxmgPCvs
ruE1eLbowBUXexxPAVkwuQTamDj424lslOvjq0en0XGpI9f587EpRzPUE678VC6/zoCOIbDL1CyD
FGckXT+7NIOikYqtdW1opfsXYNKNKbzBLoundoin7h97gCDmCQd9stwXZXX1cpojq5VUXb2zBcQ0
PjYygc1Jh4pBGvp1ZW3JBCXMJhmwIdG6QDtmOOA+rv5h14fzXU47pLoSUIxH5JhPQZTRlRIxJZxK
q8acxAKGvLS6Yq6DpVLZ0HiL2qvEJkPeWTUnjkJpyeDizl7GKhSAXwqd76VAQVsWdoQDg5SYJebY
BsnqkGOyygROAIgo3VoU50IQmCp6tqRTu31fxH8JTRuqrMdJO7GnoRha7j2cN9t4YeDzUOpiKhxh
0vRXqXCVwT+samJQB14VKOMMDQ2sGLRk8hVRo6eEMYQguQeAH3Ro8cgsWb5T/kF+nXL3pQp8Ld/M
F4ruNcw5vn6g6ZAzVp5mIeQTYdQzc9BSgqWK1n8mXyHfTi0aTxPZlbaIYSOeuvxR2kqiebD+Hd/J
b2nrVqci0J2VptPIOkKe+vBAdQ70Upt2kp9cWCbtYA83wZ9uLdqE4CbLhRPuLL2v+y31Wwbalvrb
EF9ZtoBwv2rsW+cckeDQs/gXUwqZEJ72juD+mXddKMjTdHpSh17J8uCPqnUywVHzFmD/vLh14HmF
K5TpbpRZrIdJs+WyDShnVog66AO7vaR6dEX+8wlg9bGug+3f6GNFCfvGu3OD5pBvEJLT4uKFxU0V
J38wosNxiyjsuhh+IzHFI2CYlbIolsxaiMYHOcwBL3k5JOs8w9LvsxrLkYiWJiROFaDpCPslVR3P
2SCCHZTsUFAnlS+wCiiXZesq8V0NwMj0FAS5W9IoUxhciQPLxIy5585QOCLKQEUthSilgo9dz0uq
ZomsisXBOCAUBOLVuxOcIbTvDhQe8caRRfXgjncCL3vxEKdB9ogb3eOUnHzPsT+MsRZTCXHpfwio
Dt6uk9cBWSUsN5lqk9Mr5vJH8zzOmD7i87E2STQPLxEf26nhyQt/3W2kYzdncqwt2CWhlTKf02Bz
bVAOvv61YahtksW7r06ZA0ma9b//2Pt5X70FjeDPrXCi/q8CY3sI6zPY+OtDb14JR09kyw3l0pHk
+81wIIzJJcpK+Xied9vHgV0F/o1jyuJ8W96Ov1Mm9UkfCTxUtJ+OCpuw/jDj91gVrFUxq6B0wzX2
MAma/bNZQdEOXMovEAJr1ifU3cLEb89cGMSLzb0NROa5D7B43YaZiiw2B6oBySSXFTxSL8NIBZJV
D1QBTK/mQ44KSzL6GOLDhJ8Ct7XPdZp0dzfIk0TPhUszmBOOudlWW4m9dbpNtoTMCQlPBPsxWloM
Y2We2fPNNJ3ANXBnZbnK8YbVKT38aEztzlS4yrT51iXvR499CJzVBLaXfB6aMF7jvGYJaJQ5z03Z
FzZT0RxjSNhs4bcjF2QTtT0p/sPbOKV/ESNG/F18YWKZEpn41iAv+r97WFid3P+NYM2LRPJh7Uml
4xJvXrHuBvxFB7kPOp09XkCXLuIx3Lafl03NI1B0k8oz7FM+f8AKVqh1UIR/IUN8p/Hsbvdhgtbi
6hJqvZFtcmIxiUspUmilwgnJQ2vb4hH7k/7edswXWgaa0JqwyfK+KMp10oH1Zn0oR2P8ffCdyoIL
UaMCAP/WW/chNluqYXw8bYUivcH8GncvK9DVIS4FLGTJb9yj2EQ+plRtnzFiuKTUZidR0UIIVf2K
tAfQKQdPBl6HtXAhRhJbhlZ+1b6qRJBf6sVP8YkfxOvXw5jPGpuWfKnM5sR+X0RecuSCtf8y4YaC
Jal60B/ODAfBBLZAIbPtaccY9pqPdtx8FZqR7lcsd44z8Py1tcofgn1XiFSWqosUIlzhwW2eVyvw
ckVSWTfN6Ku30aGt9mz4CihsknYQJOiuGQIIutBV1bjiHZZqQnwYddsEjbE/mHvHDL5P8KkYK4UZ
9aXM3l5qUP0gPAgKq+gxyzJC2bA8cLZGFChJ4KnDIwFTMuntRy8bfJ/Ttu5k1jalDT58wvgm41Tp
pO2SjB7WLKZeHlRJ+8hkRLoPhznaPJPWElcCvvl0z/TZ/Q/3qetptuDJLoGFPgwz7Y4eUlb0HY2K
Gl1zTO0YCUI4kx+chDCsybiZHm1JL2pZKiWJ7poyD6FVKRnl/RDlvcCTDv7rClVIUZMdpFFkK4eq
9LwQ6dvizfB4d/+h/f4Vdt8lrieHWWrvIJwhrS2TdIlbsCnsrMhxXcFftCkWb/yDvfgo/5U8xTqV
myXIAndkzShZmwtO83Cnhsdj2qH+F6He37BCeuUioPYNPAnhgXTImcc0A9MLp1QC914lVHks2vQ9
y15VlC3aVVbDVU7q2dceAp0wCdcDtOpEzN3cCIS9kjlFRoRwRdLFKPuYfKsE8qDIOUxF0lLEHJpU
mF9HD/weOvhWJxK5XFHasnt86kL+h1HMvuCZOn9eeHR3MKhd3QOs8xOqyvOm4dWGvInxdLgI1L/7
6KVVJgFOyRU4SDYdk7mujE2B8hta1m+5tT9vn+7KKGadLoNCzyhltV5MJyWd6I42ZEOdvgq/1Kwn
epcc98WTXDI4CtLgX8dg7nm+M/v/FTO/2ZxpCbOYM3QfEfsql5Jy8DwRNrLv29Bc0rD3tXgzmk6a
mE5i7scMIuNX44vaIASkyHedORdCBfaZ9tVz7bMuv5EwjR7HL449ryC1csJVnbaT2ri8YF47P662
/vd1JMQGfK3LERi2F7GtZ7jH78wN4zDrE8saeJsWGCcbm4MNcWvekEwA5/c79LsEIWs5IotNfwq5
JsZXlXXF2D6Rg56sp2jTPiUFMGNzu4gPhL8rFYeBf32uKnXhndN9we7ljyUU/wynZ8clscZiSBMo
Gy3tri8beSqlFJUmzilqdYza4BVy8JY2ZtwfduuLwGCvrLUw7svtmYnXJk568KfTiXaB0P5AFBQ8
AgtVpfddlGzigAHBSfl2QI/GS3wkCQLhi/qSqzpSVGyQHiAYNZqhEvR5AvY3bGdZhCjWL3Jq6ZvP
poy6rwJe9JLXYcbIIlOoeVSLhtgJHF9EZjZm5tX+dCaiZGGS7xhjm8e/2G0XmD3HZsfNb3Z1ZF5Q
/zprhY87irj9FhnsnYuFYKcPU59YsKev8q5IZT0cFvZm77zUvlr7paSldGIweqw4QAmbq8+ybXJj
C/PeU3/aM0Stk3EVS2ZPsVQUByT/lkISi6NSeE7QT03zciKA3ksqP5layayGkLBjtE0VZRYuxRW3
hxoywwAjkYDvC6JGY4+QrV3gmkZXaZ04kdpf/8smtll8XmyswA4yDdSYqaUDYvAB0Aj5xe2V9EjD
THm532gmqgLhxiFYauqproQ6a76DHU83grHmPiG10b81RG8dcu1z8tRJe3nF6o5Y91KUe3V/PlW1
shJY9G+P+G2p0zQ6U7cT9xepsCoFTSGMBD0I5udb5z1ZbjvgpMbQbA6VbIiyxwQWHcvbLoljm5lc
ye5dzuJzrl0lrexG8Lh4aZHWWyO9T29qciNdgqQoHKZrKcU8aRpsAbrZlLJZUrEevi6fAHrXTNkm
IgzkkH269NGScjQ9pVPCpGAwjsdlncgopD16v1Ehj60gMgHk5UuGP6a2n6PxvWZZhYD73WLZUABf
1yb4+B7QGnnpMi72NaMH9+EuAvdE/H7ilT3+5s640GeTcSzJJ+7GS2ayqviUEEXIbIyK2rUGLbo9
+bViP5WV5OIG/+JN1UjC9y8q4DBN4jFzw3sGQDPqwlBewoYtPns5eBzLaxrDyYtxlyMgwzIFozqJ
2ETiRqctbmYQJtD/NiqJB3tqYHRD/LMHi3Fd6DgObmtBf5dWgJuGv9p1fyHf9ufOAvbqkd0Lz81L
x53RYrGNldl4zck9ZzjvGAOrrdAfaYvCW6nCvl62NQZrSUABh+ESs8f6qtU4aThrbU5N+E3FM8xI
YelIDYH70hifZKZxM1BjaVYog9KshszbsKL8WBXaDzONOn9DFZGL8xPHq/A7CSEHZ0q6DhNP02gb
bYsX3+FOIAeZHulT/RzuQ3V7ywJCAHP4dwDOZHXLoKE+H2Vu2G7Ikg8psFTa/v+vKfQcrC0CL8X1
9Xpt8hmJn8xSK8i3C+mRTY8rzyUii3gRfPahtJxhdeWSWZJ4rhXK6W6iTULbGgLUgPY3bNzwaFJL
0MH/CYcDyUljL9CqkWijdAJpQGLVBTYNsCkXLKAG+Eg+Q5i4GrDCOPKiUDOQmgsCzO6pw0GlwEzd
7BkhzN8uXW57DD94mGRsjqfRm3bwTwtpPrp96PVpZWvB6g7UB+sD/q1z7xeKxVWBHVXBYPUhfDaO
GyJUlRC/5AoUEsnEVXv92AtbPTKhfBVq52Vxmlek4U41kQqvP6Qtsnr7ngF4w4AQExoCTNPDlXnA
apISBJcKrfjb//K8RsAba9MkvzMvrdrGopeghXhQ17u80R09Y8U0NObXtnIkgEpStejvUn5HzRSz
kCz14svSjdN13Wym+J+66O1+uigIAuf4TbLEE+iEdNp9tfO1svvaYfv1sYl0Q1zFP6+SZur1eWk8
4yxOWxSxIAIT42oyJbH2/4pBdPn5Hw4w2dKTX3QQrLz7yEyeB1yKGZRlwhcwszV1BsdV9UX+utdf
3LCJ8bBbEH9nRAflK1fFVCjDINeGdsrsASXbPYLRT682lkMBd12CeQlUx2mqOuAXlgsjxsO3E/Po
KJsEfSxXe8OphkNXzuYU1hoW34VxuJOUcmzI9U3K/a4//WLtEe+BSBWuilowrQ6OF7kkDRvOBVOx
FmL3lxE3WLIHUe0byRZUyKe1RMmvjHQIcWeWVfU9KMmWn3bSN2DU2vC6JDUqsXlMm+2+KYYtDktA
cCTHBFvNI+rO0ocKJ2wOyZORFnrXvGz75FOpd4mcFTi8a2sx7LC0OJb30X0VW+K8KbrIJPWjXElu
W8bikDvccVuyz/I8YInQIjuJ80zG5cQc5cUxCTpkNXO/cxMC571EiWHYmzhNM17PRbI3Zwno1gDM
M9kvk8hPZhhhgpUiJQ66B1czbmnp+VCO1v1OhY6HIFamLOhVFoD/NtkXitlQ58Z80FJ3DtDtxRCT
vX/BRu6et3SRwgeGNCyOwDdmc8bf/Dk3XmcEQCtJMqVRy6MfLN3H9HvWERzwjZoYhVdGrNsnQPxv
IudHvkoUm04V3e/Pb4xNBnvhpdLXc0SoM4CjrvLNpH4R9msPGvImbH/P7vw/bYBn/ck1ia/PL6ji
vXLR42SsqZy/URi9QvsZ67HCiLeZOKnIsUvpVDQuJGVRCVjt2fiTv2NR3hp5URFIZhBiygJuOvqr
OV5IagCCSgrgsG6rHY5Fp92VAtO0DO/GFMhTHLm7PrHMxnUy6sCcj2y+VjRrtsNm0jRxDj6ex27e
9C3wV9/XuIshvifcAJuuUGWZ54//VWlmtf8z9XnlEjpocqrwEtEofo6/lslBbTamB0Q2sHanCDNb
UmLoXjuvTUDj9ywaFjBp9HjYYZCI7EActEVbaGfJ3ppRoYaV3PjIEJyYSvVKOaV535quYax1pxtO
QZTMWwQeQFQFJL/GOTsShtzXip/duthWmbZXlxe8uSLAbVmaLgIAk9NDnrNdSfsQdksinr6PMPvG
5B24onBIe0erZpV38tEauI9l091epmwAFPGkWXOli1uOu3qlFHp2Utcll/zxMAQlMpsCgo+A1eUV
8scDReFEcDUXDUS0X96PsIir4kU0o7vW/6cPaym7betPVimRsOCqfBu8U1bQIqaA6ucBHNlrolvQ
whHYd4P1XBBbtETU4cslEGE5fpQFRtrARU4sGFc9lxqG+X2D1UFUp4I586M9h2/hAdg/WJSEjvvB
8UDvwW7wSKWWlDvkUT4IoURzij8UR3I7TDABp5tBdeos1jIV0cVGuR/e4bGXpAZN4aWAohDDrG9A
hcfah/8yJbK98GSBDTuJcVpkCA69KnCCWKO6VI+TuHybGklSrz939Kp4rPSay7Pmz50q7WyGBfmV
bzn6erLZXgNPnkZKRwvRSQ7ydbpY1CTftSTR8JLJiMEnfTTZFIHoRS0YPOUoFurVPO+IrsTXdVKt
2INuyGxUHoBsrZ8heTUhHYdxZ7MC6REbAUbsHG7oVpvS0Dm2Re4vH3yk3NFZmu9PzUAk79Bo6/Gs
X6VNmFfKKYyfx4aO3OvIrcWtM03kDXyx3XGKqCgfVndEUBLsXufve4lrMbuC7NihKCupvRNh5ygi
S54gFpPpv1QOfp8vG8UR3inVRLY2ZNlAKggTTmh9JWqAGrJ7HpnmVLYq64oeuVwmSK/IjbAUrY1w
US+nGOOKHubhFtLFNcbDhA7ky+uXkD93gIGIv+Fh1x3bJ3PJ6p114VVruZC4DHsFQwV80Ya8ON0D
kozZe4eSZz4BWJmtvWTnBoIt1/3O/fRzSAVFhZYNsSg4mb8GEUXQPRKKLj8np1QyofLtUgEUTbRx
dliRo8jedDD6eoIUshJwKqSqzQQvyjyzvpAb6cPeb65n9aDbeRALmCO1g+q35bQejvswHeoKmW0e
P4F5z1mTF7oFJkxUOTjGT6mXN3p1REEyWABdtSo7m9DzChmdOrdssqX2Vy0GLUnS8JQhBh64/ndN
LxUbSe3UjFwqv+wGS8IdDAGV1eN3dYEv2UIhGcuiKUnKIWIb/+/gVVjq2nGhasCPSGciZUyhf8vR
EYYsrWxUh26m5fNFK3OkeHCzEl+K6/RST30Xse6otDuaHCxzNpTLQjO67OUc9szGeXc3eURijtyk
oKGLCBIkVM/EfTH2kP2OBfD3Fvsm14N+WX0WIfkUNewadb+v/wjBKS/mAekQCcUgvpr4zk02DTCg
aZBS9WdNwi01PVJM09SeHSzRTICbiMSrpecKi8P0gKtjy2caMZtxpDgPxkEVNIFgNIGW/aRvfPCl
dIH6mt9xMvNw7jzD8/i+HQA+G1QQ9AI3/QRpk9b23oIi4uKWF4Xt1MPFCuEKmT40KZ+zk4CcUTUN
XnpuNl8aqky7wLL9eBoAkHNsYWYVjpemP+LNljL4eHyI1XZcBxczagq6YiCubThwzG/zearDMvRi
SuUbsp+BytOnBQmhQuoyyBvFH9Edyn5uW+7CgtQ1qROZoBMmwDyg2VVzUWT85vLgMxexh9oWHg9O
fL64sPBUNK3RfJu/dT23EJr8Rp8v5NwyYM0PHeP5myGlkJ4MAfNFsQTITuRnFLu7xssjY8L8xVQ4
5CkQBSyBXaq50JiXxFbxeZDAneCKXTVlD7fNidYhEoY/zSJybn82H/VbIu+9qPH8ez/LH9bdKCgT
7+3j6y9MMd3mKifVOIIBwiwTZ4ok9WZGU/isdQlwpvvsn6hNnA7iz6tuLapak6rDvIZx5w+GUY39
ElwLliw9sZjtrT4BsgG5IhJNLsDDc/ozfJ5nhBzp0Mmp4BulF6DImoVyI8XClOZUQd68oNDCEhnp
NfAy0csnm3XorYH2xeMXJ/vh/GcXdlhWOUAD3ty0PdSRecJh7ncINO4AwfSeXBTq1A6I9cwShJrL
Em2QlH6JJR65bS3AtDt7iSS0DxPBj3Te1sA/wwjOu3RCD/D7yOBJVg9N5rUHQyHzHxGShY5ggp0i
21U55kFutFghjhfA48iOYl+D1rLFWPVOkdqrc1ZnRwyuvZTdBxiRE5suWM6QfDuj5TS2ojf8KXgB
b7F+VVJMqdMsfsG1E3R4A+HU19o6aKfcmCBc89p6vSNaWUXsDHPv1oUwpyfgCpy+KFPPjbmlde+N
IqFcowpkLAcHjR1LMEkHZ+7GgCfj3j41c232u3p6NLH/7Swv1FrLhJzQH2bTqP19Ofoq1QGoeZMi
g4gfPbF12kx8b34VLJShLmB0jXO2xj6/H5P9/KFbUl3hJhLp81f4xFXijcOOrohyA+5EhKmcUeFm
w1cEYvuYUuH0C/gz8m3lEzU7WOIhjG1nGj6SJ90TGs3iXK7R7BApnYsXAsT7Ft7bDH95cmmTSmi6
jTHSPH/c69W6N8l+7S00CFo06A7w6FnEbIQduIgobUtRZJL0cr4HX199iTTZpQmUwksNRVgGlXu9
8Qk7i70/40e2IGeaekkcp1aTQ9B0Cm/rqDH+OVwHqL7mL+6UUkrOzL59jmELPnn2VEsUlJ3yGaGs
NnLLmI1eb58JWThJCib4nB7K/yOifS0HDO7k2Jay/gNKVjl3/F5h6XKaPeqZ2AsfW3CGWW9HXnOq
ZgeMuFQpK0sLHRp1mNEq+PYLsGKBlhGT9Y87X/rKh63Mloa+zlXvPn0jkKR/eimLE3m7EH/6GKXw
oK2+iJtJGD1UEiINLqaF6QxpwVAc8Hsrv5ezasY1Fo17asH77A2eukAYX4aMzvJkkD2T+CUgx3RH
J6x5JMFCgeS7/aSKkozV7v+Qf6XMMbLcChGv0IV0cNnAo65kFuFhQMqF3k54gg0kUeAOVpnwvMHM
NCPaoXbgk+Pqyki7vYYi1g8BMcEIbPvJc8nzTYln6nxAfBtMRpqZJJ+PWLAIGk2IV7hEuJxklHsd
lAGZ6BAaaOctpz2j0XKbMGavFROSGSTK57BQgd40Uhwqd0fym0sD7REfMs4jClGNWCP3fjA3eE+B
7xQiDbEKfsuRnKDf9fyeYuhgyWQstRzjReeDVaqlYIgtgRElZ55R3qsxA34oTeM/9LrTjxvtA2b3
FlVXzV2B8u94sTzQVRmwJCFMvC/dkbQDZnDz7LI/iSEXEyG7rSi9L+zMxx/Qaz+7wOe6ZGe4YK1D
ML7LXKm4z3xMlHxw7RSIoXZJXUq5GA/J8dyuoaQYkiLifU1Jbs92O2gLK5/ZEEqC1jUBJSR1nk8i
ukV/bVPS2uk+NxZwjjU8N5jC8U7FtxOyXwKy8JhS2wTyv4j8mqlBrKd22YENvwPsa6hBgBpVLSeU
QEmbFPpsXrgo0A0stpb5OUfyHDI+R+XimtWKdTlvcsPHPOeQ/m+RL+dgZzmOIsjKIcx1hqrWGjJE
D5XRgdNJnIl2A9jmoFPStQF4oDGMqTMXitNy8IO1MVHjX4BYVdMwyAOS5N/OGlGFRVwI99NOBelg
99B9vDCzpFdfZDvh/wlGeSduPeOht1xaJuoR0Lmm1lvH2qwSaZtQeY1Uw9+mEt9oKSDYZwtHDj9+
erlSN9U/CexknnXz47EXlKamqUkUQINpEms4HOttuYXQh2OhfT8Te9Tx8iA8sphmwBJixkWfnK1E
Ngipyp+fnUzE40C/W2P+DJhCIc0aaJXwVWskeKeCTWqqDOcu3wcZOo9Lyxx/YpqtqyqA+uZynKbN
vuEpvOM7tzJ0c9kPBTHRU0rCYbppwSPnkpq4fHcxvO0Z4/uQsjIDgvc35zhRH+ZjNssWw5DPe7Mk
W4pATNP1EiI0rCwaEyDleLBWSUbNK7HDaRWOkcF4QH2WKg75P8NwNy5Lc4McbOUhN+Xkp4QqE4ak
4pMtkcsNwqwa2KsW6Kw8lT1r6ykhZ4txEgz93MB0x7/W6/6f9rjaeT1JdW+qEw4fUsUe4zcasPNt
EN5quETtf+VSlL7oysGu/WcDvgZfk4y3wy5bUPdcxsaFWSvXWmlnZ7Mkvht6wXvYHdV7IGrqXLXB
g7659fWrOiwwPVxlLs09pXXhDcdNzFvY6fw1rZoldvbEDzW3znLltpaqM36ywNRzYp9ZAcd4wsGk
zA0dnvkQn2TMB0xEnb/EXzMtsey8plXgcI0fM824pc+W+FjtGgDphIMioe3nq4+EaKZgUr1a2J7e
vBywmgAjvWEIkc9WfHhx5Qpo9HdL/+cIuYeYTm0NZWbBRDCfG5GGXVbmQNM0y5iED8JO6Ab4gMi4
aEdqy8jXkH4h2m7mziwYk51pnjKsBc+m3tJZVSo5nesVvjVdOKdc0pfBmBrJd/uZ3CvsmS1Pq9Cd
PhqhSJbKYDAFA9hc4IvEgmKLh1rNSluu2FT/i4dApFeQhP/NvCcGj64+h/FqPAy5GNoItFTpboqA
D1vKAQ6AneXtSXtha1EMAasJ5Se43BbFOFtQiQ9+8JPwu3TaTkMDmv+S/+Bkn/jn1eduBi6sYKVC
BIr3kfVLRomKadCySjBbeHy6qQg0G3MOwUKmfx5L5gNvJgHZ8bphgwr4yROW6g2S6Ko+TEaM0vKj
XUr63cXsHvHipokOy5kCDSNNNam3dyB72XG7F+PqdukUpcI1ZGgP7j5LKG7sOVfm4IB5aiTw+3GN
zcKuOeZZtmFZa1VDYq8Qqlh2zS9Bo31ZPY6rA3iRermxoxItmEXSZ7SEq+uOuiCcOyb4ixkGO8+s
9yLyXvsdssAhxOIfs0OitAfBIU2Bad9vZBmTwVbKTCpSW/9Bk2y0tuMK48pP86RXd3IfS4t/gPRJ
GiOMxfa2p0OS5yCRvNBUEReHVdXB+wGpwePSsS5pO91LWdNL+TeSxTVwG1GTvgCwP+t+tU0LNDsD
UtRmOe2x5SMXtKx+mY3JJBwLrM0/AG3qYevF+wmLa/S6/ePSxT/Q2Bh0z+2eoeH/whjUchdKaIwy
cbRpyBwsqQQd+1s8+dQl4IOFKemCmIJRqZh8kwLuvuoTfniifQSg17kUz7xr1lQCIB/unqKpEwfV
dSAbzsZI6BnSB+ANU2cjb2GbxndzMO676qde4OhtU5oH1eiuOw1pS/qjXD5Cq5cq9HiP+CVSJEO4
UM38h37sWFfyK0BTklJ1GldjEsMAMo5F+Mf5FioPhIm4XjwzTOQt3Z/z8TVe5gSt7z+WfFC1tw8z
NSsxPmBpMspSqgY8c8b8T0Qbk/4kANGgTW+FONeampSV9DtZxQE1PtX2Kj254q6VpU3oQkqNdLnz
qFu2UPz8IcPNFY0hBN5kVoRxLGX76xb2oKaPP41/HIlLLtjyvOld/B47VB1+H6uImR1BUjOm4/O1
XDZ+YpGmtXQL/6Pq5veqMTE8FI2B91ZUPe1Qc7ul6zznrGIr1T7NAPHRRjBNq5MYeAppfvFlcQ83
ckDfnTCACMVIxWwdmSsDd3Gpu1Iql/eYa96joXVFAa7cn7/5Tjo4Re3R5doPxLsndCYECwGU9ctx
mNyb82MIfWQ5DvRoc/uPhcsD1Z/EB9qe4Bl1TuvdkmykfD4xyZbo9LpvckF0YHHVUnwyhIQ0Fvvf
wwWnJqajJThsyLxFTuQAU/hAIbeGvbgDB4YGOI8hg5NTxiT5g4Os2xj+666Lr2uhTz/asNKHff78
rVhUDfnggSBsXHCyQWJYT1/67ZIUzLpGTsY1z9nrFlSJt3scGjiqUYCJFtpS72N15LatgS4TnsKH
TxiwHCYuCTdjxJC0+8pRG4MaXs1rusuk5D532234hLjXSP2xE0d+gD6RFr1p1wwULcxsM+J5/ZbZ
zR3P4jph17/JpGbMjRmf1ZAK9ZVbEnhus96jGsVclovMh1BRn8FgmkqyImmTGxv8mXxInnjZ/tVC
9sU8+hHATbHgg8yFDgu3oMshNnTVpkvDRmv0d4FGuEXXw93kYuCeX88plzppwaaIqVF4fJx7+vCJ
LBkSTRjd0IgWI5dJS4X1Zwd4WzUa7Zn0ScXaAisiGJFdXivW11XSMqxTS7K2tbSRFCghWmsts0zt
pSawySl5jedwhjgGjwr0/xcmcRT120oTtIT9FTzjIxj+p4kz/8Zl0bqqZb406hkRQ4lQUY5S+5Su
xbt9rTinQhc86K/riKxzFavNfr2BI9JoEfjAumr2Ki/6mcOiW3iPiyDs8qHxIqfkHZy8frPIB3O6
4UA+HXhWGDT8zFbURVSEdfUV3YMmrRvNe0myEah637avn7QOB9Q9ejAEAqt3j++hFp0krjIOn9nF
JFI71j3sN+6y7+8xJIUlDVtfqknvZJHtKG9b6gveNu/NVQeY7Sb6DzA5q2BktCJw+nz5SIJ9AplY
AnvfW4kQBHaytm/Hzx5nnVXbvVPTIo15eK/bR/gXVvt+0fYX1vrPdhpILQflaVMUgTxYRGBRsCKg
k8OYg7enyh3KMeOLpp+xVIVJM4coQkvDwS2OU/4l8Fb/bDdoiwNL6ajPhNun+7QMtGp0YanGe944
RPR8/6/HctpufMqhmqsZ0oaC9lVl8A43WHaO4z56y4Eaxs9tdL3ENqE9VZAGzpSqtcoR1oNzXdI8
8fJ/YOZ6YkItvxVtXoGYfeDh8wSrF3zSMrFdpshJN2F5jkBrAzkG3iJG3m1wK0b5inl5p2x3HC3w
Xn6hHPTf0QAQ+wyAKefYRQIQp4Z6PCKg0OpHSeAc0Gsvbu7lIpYiLZE0dpCG3u7mwp1+6494tUyW
xD72S6DdajeuR2KncwOB9GIvoMN1roHkhjKTPnh00fFpkgimrsXIfEeK8SBjO7vNwDq2bnYVbbya
B+bNGIqJ6MqHeAB6FOpf2IRXcpsIcGGPAXFiB69sdwQDnb+0G8mSl2mRLDlO3Vhs5z9pUAcz4C2x
YmTyylR+aqES55hOYP/wIz8s2nnpGYaxyTGMBSKEqaF9+gvSixhmoZ3dpx72Ibe24LkGUJCQSAWz
YnAQFb0nNSWK5eOGOz5ItHc99lQO15WamB+HN7ogjcC85XOmrO9fsgpYxfyDUUdN6Emjt8/uL2ZR
ncQgNy/pccaTrKED/Nfbzw3N9nETLiJbhqlhsNMk2D6ji5M3hPc0w9B1hiWJpvbwLdiSROizfblM
mUj1YrdY0FNROUvopVTK4N/DTtgtflcFGc/IJEz3qqYy/irho8X5ks2RwuKzabj1ewyCS++dhrDc
1kRAwruOk4aolZQ7FXLcopM2HtgSXQZ1Af1g5D69e3olQmFZpCdFvVhsLIB86vPrFnRad5yUIBos
SY8U1boicvtQpLQCHu6r3ZEehc0ntZuoupzLfzfAwsGuLmsI1sO+BDBEBGdZ1HSuXhfOeRV+wW73
jCLOMId9dQ/Gu0OLaeinMhRKgH6yIxdqU8Gy+KW0dy64vzwoxqg1k/cuLGgvVkz18PbLs4DGIkxb
ySAAaF7ljMhgby7L3sh3tyBJ73CmuNK/VgPq1hG0SxlVQnODRrrcaQjbdTw5mLF5ZznsuCJQNCMD
e+Qe+l0Z/Qh9Mv3KAZJWHx/lgBNdM620JCXmJ7BXtBsGaIc2KMs7eTCzQvmDDlWgKT+8LXwg6JZA
gMcrG9SifPazaiUXPuFZRcUAjvyHVwkDeETlNk6GYwKKR6MT9Zu69VMAZLVQAO5rORzM+4+aC5rE
Gw5FPP6SwuTfu+qok+xrDNsXLEGMZvqOrQ7YASmdhB0xImnvlFBeLZqxEHdk6NQjoOeXoxLedTi8
5oUFU85LqBBe6KOFnDWhsNfgpzmASFybI5Sq4RkT5efWtJ7F0hJYx/bkZCdhVCoU3lFexkPpxr1B
2s6VGq0oPARkal//9LAy0SH5wJ3K6yEfc/hnrIB09BOs0A5BYNbCMk51E0+2i9FEV9WjPCVQUOWB
B7Jwt2qCWLk4EuC2EuNofb30Rx6+HLtckD+6+GiIE/Olu9gP60004+BSD0K50jnQjhaAxdwCer3g
lTloF+8XGoU7p6JVM/9U64GZBaa2R8SL4TBE9Ilf+yqExFLT5uSDh+Er6+NK2ziCs2VZ6/QkEeP1
WUoZXyYfPwDAOljaBJFfDhW93+P1AlglPDs9CH0nxCTeIcHO8Jc2AgBufR5dDbbR5214VGDBcVNO
wK6OJubM2iyR+gT81SW1Oi40WV+wLJh0HleVXfXcc8ynjywMvj4g7rmq4FGUkS/ykh90U+3+vyZ5
I6bW3yMXgXjX69Frl7sdf7rZN7jzhTOgmsiNzTt7r33/05gZ8rxTDQ71ZNoU7TX75RqJMAcqOP1L
1CZlZLq8LtqCJLM7qiTE5MXN4cxghIfi4w35eW6ngPh0+7RwxibWeQJqMkdwYoTHZFz9DDjaM42z
2nGaTabs/JbI0I63SzLLGNP6Sz8Y6akwza3C6InqzUPT0ELytfgcsyJdkyO1MlU+ETlETGhBznWb
XiowgTZ9gDm8ZXcmxwNx2tKLgvc6KOGUJC+KlJRz/FAKYSH3O9pHokidcBNMzNHZaN1zquABlcoG
sWOpFKnnmpOJelNet9C0Jlj0Wz0Ths07+/Gq0STc1ptG7+tafxsB+DqeaMlr80lpGIzLvG3lYxts
kCTEXVaQWwXlQsBqMBcgo2W8vEkMfaiNnmn2Yx0pVctrj4/zJwtj2f1DH9z1otzHWPvUXAM50O6a
2Bpu4AcCPqdqLOt1PTeWqRucUFxGUGP4gSKi4gC3QBXOz0qYR/vEPCLcsCDyaijxZGGM5G738Ddd
c2elgNrr3GlArORXA8+NGDpk0ouG3rsB73EIFwcz9DSfVKz7q6l5EBNDh+L5Se68TcSPXzcH0YhF
FLdEFG+u8rAAkmtNEG5AaBBIJkgIjqu3SzrfPbSeReWSB5sd41jahH/W5Vtiz/hQyvMP6K32szxR
EZZN1CkQ/iL0iv0G47MGVg/GarcoYaa0roAe4fBzPsi3FbpfO3UKEV3nFabw1ubGURQFljqsKuu2
b/WUDY5LiVmat5Zh2K2PUFNaqKuvDh5EYYDo+d8kz3Kbh0K8E+iPFhSC351z+YVECLcF3W6DMgTx
jg03BdNk6r/dxZcIoJg2E6bgq6nef80TS1XXLBZ9ay72nSOGbflftbDpvHnNlXFFlcwJVx40TcQS
eM5vqH9kn5Q2fu7MjaL7awdPGFZIzNoFTMuuTEQQQkY97AJIhi5A3sRJW3SGhvNCdlrZSsUhdCLP
X0r1vn8kVicwYXfoWGTjFdSCnx40GJWPziagBFeXSjxzOt6Q37FPGZJa2zFtX2qKC8ttXPbhv809
w94iTCVberGEjvFmANdegZSp/pYQP2cp/C00qDsGMFfLbaHJrf83HiFiREu443tVjEyv5jb4kMul
PmEsb3gnhIuBJXy0hCnVG6lmL2ONhFUJLXdzIPTGaPcJHDcIGAASkxQEfUG1lupdQ1wvTj5YYiZZ
TifaR4+FdFcfjvznqrKyMuP+fO+QhoiRLbDyCk0y/XALWBI7e8QU2EJYEVAecZdH8mFcbOxiO/7j
3obvmjQkHmH3Ib+5CW+4UbzV0PiRTaxx5V5w1PAPWaieizmAP1aejIhKCYB5GWKlGfB5eAdNvbNk
YazCCmjWC1Bk79gVvNPFor6a95jyOug4HCVLTnYF+lnppPOoT8KUeNnfCD+I+6P/Mgzy+/s1CXD9
c/NAbSgoKYu8NYF15tyTZKEDAzDJWxDBANMVSMjg7kEUok7EUeJpDDBAJRXhYehzIaTu/I7+wRZy
crm7GmBVLINOGMfJ84EP7rmSRqdyP5LMyu5D77jzXuYOW7fE5ojWr6jl1imWLyRH52xJvtNk1k/o
BufeXK9zuOocr5HK5Rnp//JrzLNWp7iAV5dAvEU5TG1F4N+oUBbnM5GKyvYWZwI+qELtz3ILKU8D
wJVrVkyUlQoHb2eYONOzxtu3RwVUX0bAQr2RkKN85DyC4p2LGDmtp3aDUhe2CRFYL7VN3lQQkZ1I
ShXnCuUoVG2XqFvNluWPlT8VjkJxVO1VM7IFdZd66CRBfZG7A/AHlvNaoIv4PWS+f6fS7DNdSVe8
DIVRdaRmMdvze+1zO5rKTcFRzWZ9i5ZkwkstBRxQ6BZJmfw6QplOhP3EhV6HNM+7h5c5CWX06r3w
sQjV0ZO3gY7nW6bFiSoNUQlAGx+DiJMKmbKwxy5eaWn+JPZGhG1QAa1vkY0RgK7yv6M6PD4/pgXo
C+u/kAcsz483iKOFKNkWEniTHhj/XgWoDJ/pbsBvv4BOel0Yt+2uxba8oWHlZgAMvrV3c8kI4Dfh
+GpB2WmNWE/J5tq+pIYtle35t7Fn7xDJV9HCwCTUNTPPClq5T0akZT+rdDAJurgKeGketglrI4Zf
cShR1x77fPFAkAm50t+boz94GM6/IWzoJwBTW+l+z/o4H9wngQSFEDeLnM/18aDn60XzMlr+6uFi
2Oe7tgFhuCd2wOuA1O2wk5IFjm2Y9rcUefPMtuX13bb35ZjfF6RnLwafv+N/l8TBIRXKQkMDfPMU
fzgscE1tz7tFDmrD7QX0S3f/BClhErsFQDt7dZwBaiQV2b3r6fa94NcjWKcviZUYCh2T8QS6db2N
aURFAXnPPD2s1c4gL4NO/sBOb+Qlk8hTZffy23qmWHFJH7gyxVIamtKCOWeu6nPFLVVPDVMzpfXC
hfXObktOpEzxWQzE295KxxilcwGhaNGpjnzRq8DvFgaOZzDkECzUFASDvDYtCWROYxJk/A+y660G
PPmHl0XGN2+8pLefGkCLtxE6LUrdvDa/dlv8W+RTojPrWqI99JjgVHzhxL6WY2J2gwEpSj7G177h
fWcl+GRp8gS3p2mXUHuYIXKYLfH3kF6A5DkR73c8PK8+XUyMLgmX7rCXxo+JQj8243VxchZLoSYp
+Y6BkJI/nKX0zDzmhj8yRMDcDOYdtlm/QrROmPZfhiZudh1+umgbMPpQ3JbnLrY5K0I+GQsmS7l5
/LFG0FEd3SVbHLcMObiFzN2Iha+6JQvyvWlsm4wsKE4CPOrY8buy+qlImEgtgUddnucKF8V+I9Kp
439NVkNONtlmSiXXZAyTF//GgXouhTlmZv8HP3QDal05X45bSwv36yTD9j7hzOMS0mAAhBYD7/5i
3gTrIirKeOX7KCLpdhajZ8HkaHu7oKRuMZFtNOX6LzuxuPFlNEyN7Ihu0PnMWbKDTvoxRyanV/gZ
PryZcWzR07KmN1mPoFS6GCdv9fPSoNKfFuMBhAs5HEUcr0BDtlzrw1Uaa2UmXsaEewvhyuDydwgI
gopE1Erze5UGEx2moSULvgSpKZT8YHckzdh7frKwPGDCK9/7NwsvG2605lzRz7+tK65AFRuWUzPC
ma09i5oyL9g4KsCdVee5oL9GBk5DqNMpPEXOXQT6JjCpgKdGmncSf1IRA5XXywAGW5zKPj6ZXlAX
3/Dl8A/Hu+xn4jWwX6QLJ8N8fE51ufVSI7a06X1ERdq6cVIs8tP026GIC3wTB691TtfkotiJrqtj
9gL7BWV2Hq8+1zC5eBepUhBBsaOGcCgMVGZ0v4CwiJVWcUxC622P19pvwXBPhVJ6ZMSHddMo9Jg7
CFjhFxQWi+0E+mVw5E3ZLXWQpPeYup3VTeP/Lkt/uGBSJ2J3yDTgUSBwd9u/0LHLQ6bB3vQyhnkJ
u1l753bzz+ZGVUS/5DBqW03kPrUKJhVnmjgbFpRk2AyeKu5M8QlguN3y2H2QhMa1ERXuwr9jVo/J
rL7Cd4szfb3KNQ6BC51nPE1/s9dA9GwHPyJwx6Ll8mJjGV93YCl6IKhDpwPPlS+M+zRBBJ41SI45
XuvFpf152q/yz33NdxVRGTaNiIHkO/TiZM7H1dZQbtxBrxBeh7NBzENyGJlXlEVpf2QpysaXCJaT
WI2lsJsbd458kblD1PyaJDUSUJ2ncBT4cO8rPz28PGjfc5fPkjoraTzO5RR+um2GzfFzc5dsglVD
VrjhI5GlDmNAnjMgdp6ZS2yq5BnsmYBPsaRYVlhwOVNfN8jLMUkX8Lnys2d7airAmh/72E/dlz2z
by5XdcnN2ImiM8Mcd41VzlrN4VcdIaSoStNq5Ww9FWAOijN5STvU9binnNbFX1joIWym5ZNOncQK
tdOxgCSds/JqolCAzsV8WhoZOa60KCuaTIRBCyj6IywezQ/16O8dbMFaDmIFX+2q6U5JfXog8fJ3
x2fwl7DT9cDulRyRn4oJ3Ptz+1t0nD7eqKj/mjTnGDb9Nz3fVPtEuFsQFMLteGUfGSPaiftNdqSs
m7e2iKKxhjaxj22ITV3+/3wLRl0HxKrb8D6nz2SQ+XtQmZx40lEl9lFPSnVTstVEikl/eqb0dSvV
ZrZ3jCZVGrpq/wp9uZwyISO3CZxjb0Ue9RvOBPbcWpblwRlcZzXBw+OJqTnFUowhlZdoj2oFPluN
RM8Sfkz3MVp/FjRCJFqzxwGWDn36/Bf32vkOfbuikajsZP0SIlxmQBPYblnutA/bpB1bD+8LlRQN
AcxiEtgSkrYLpxbV4GVO//T70759/kp/T28Uxz3GcmHLZmiX94+Vwh/HV7Q2kH7rFG85CuTJ2Rzx
nzJI/wRrfpfd4Sil+JyhwV6Dv7OW+3VUu9BAAZ4LkO6yzD/VE81Rz1MBbErz125PQ7hXjf63iYVB
Sur/TD0l1M+FYYaE3cZVn5lfKZV1KWfLSLNuScP9OOVItPxTc2crRz06/V8phXWDgF6LV06dVW++
CqjuFkkyD28DlOfjKomu0gXBo/fR8fDcFYqbT9DfYV0b6q/2AEW1WdafSYcXoQw0sjsUh+hsqqnk
IjNeMQ6TylZAssuIquyBAOCbKggG/je8M74ICOZUcgIgF6NXnKf0rc5vU6EpbL35AKAIe2OLY/Oy
kJSy0H3b1njrF31xZjJDrVDyth+fdYeE2L18lh3Z5JoxlkqH4oKSLsUQjtRCANYw2pFqd7jp7023
eLK37nvJKzySFG2UvMlq4GPYinaUhs4P9wuWG66F3IJ3IEbl4YtY2sxPB1XlTBl9FahTkH7VSDyX
Yv66mvQqIfyd8hHdd401hO/COeuxTGTvXogAAmRSpoppJL4ooAjPOdW0eJG03Wqr7vKf6fFAlAOI
J/tLor3yHAhrjt0DnQ6KqWtvv16E7yHL4M6MNFln8Ft4gqGE21mNOlS50hGKJks2BeP2lIbXuRfs
q70v3aHruaHrfIO2b8mUjBVSOpjyOlsXo87DKuCkbS4XpzbJkFv+hMLexppXoxnbJ/lBN1Aga/7C
5gMjZFLEfqBS0Q4yXyN0zH4PJNAcP/tdHicSwzYmYYdyYxXjOEiALmg4LRnT29flYIi4ttJmQPK+
gI75rIy2GEOrN2uxx+EpB041cXWKs1l2EHdkb/hibPb6n5O8cQHoCErkV6P4ar7LlDBs7dvnIxfj
KemTWNc6ojNikFPZJtdHulDwB/GOwQbD7+mVecHiSEp6B2/xX2hIottAq0poHQOOprQNU28PT0Nf
f9J/3iAEmtK6Xcc2GtxaqE2/NUtXbcktGDoUA1ckHlS1D9GcETQZ0S28EKAX12ljmQIidT7ZIiD2
6DCtM1KQnmYPl9WY2CCE5DiM3jJ9VcWZ96+FWKJc7bCw1KUoOiEVDJK4+TrWP0fS1dr0xsjCnHcG
cU7AkW3reAv8WV8/rcfslBu9T7bbr1nUJstnzMEbZc6L+ajw+wtwvAlJXSBgeHoB+SaaPjbSAl6g
3N2Ovkm+3+CQZPsFNNMympM1XOwgPa3xNr6ZcQqA20+tTow6EVLJd1ogmcuKzM9lJa+ua7XQUTQl
sAmPPhIseb7ErHWqKNCzvWnt072UH+Fy4L+aefBOcKgP5A+OEBCBu6bfVXoxAeS7a/nPFYDVWmrc
o+HaRxypUafBCbe1tTH45qtYocOSrSKjII6LfyrY1emgszJZKZ/+4AnKmBQ/1GiUZt0Dr58KoDb/
RoeBf6DB+ZV9HYTr42dGlJ+Pcu33WOCqhLD8gc6LPXXbAC0yIVVRnr6HLCgCmnFiMWJEMUDvur09
B9UFFga9jqHNw29YbvN6I70vqxIUp1nEnVnhr91JcmC/CfV9WmBJLN/kqNYEYr0d5AUwzrc+RO4n
O9YkvWma+aup8DmEoDyCsVvxtdrFuAGu6cBwt7p6lL5W/jkdnkmJH4KSU+BSRVVP+rEJhBtsAJKu
ce6HLJF65P06Pt0okE3Z2gAEQP13H/fNFo8uWNouLHk4rVSXqV3yra3k5bwBsbgCpjg3Y+COHmai
VzL/Wm0aW03W2szEVIQlgbBA6hBbOnVq4ZP5jIEyJ179pTwXMCrGQWmEqGF8hPnXRDfn3qzZF1sg
r9PQU67Pwq2LIbpF7LYVt6XgdFlrKtrSms2zpuoedb31MJqS/KAKPkj3jHqotUe/2F27IS5XsMGm
6bejvgKGqguP7eUrm7mfb3jWyBph0l4Ab1hFUzCmbVge6pVJIDeHcxILMKEVNyGXcV0wWsUakzzB
9zqOhDns4Gkm/u4DzSo0ub3OiVP1X6WOQrB8dlk3vWMXTbDt+W3d50j24M19GgdJdWABLElGHbbl
bfBpxqA8Gn6bTBjlzvNKd+VFTjHt/UaOGTqbU2pm9BAF4np0rlzHSE2V6ktQsoJdLtVAj0YAkbCA
w4k6YNPsiRCyDb5yOnqsUVcm9JD+h2MvdrfSTVq/sTsxUezS7r5ACzYYFMViwdL7z17X4R7Ep7hh
oulptdOQ9Pe1p9sSWSq8VsqXk2CcR6ZjEpL4tVksHr5h58cpQgQKFfisQRdXlZmA/IJD1DuIay5V
y8R2GdJqe1uwHzHe3ftc/UQIEkb8Rm+YZhfN58BEHNUpeC/eNH73XHxauKM9zy+b+4fpYL8xolGN
IJQ9lWK/A6MR3bjGVpTgxVyCXIJwOmUJ328Dz5/Ew11fZgMQIbCUazuyAs9eTyHaqbu4K4lHV1lR
ijsobfWrmLoFB8KISjg0l0AWBbi7SB4+96t8P69Ysu5CV7MRkioCgJcYQMdtGwY/+Sz17ceAFBP6
hmIJxD4mGgdj6T993GD9SxrhFWNFWoboBI8WZXdwY/KMRaYVif65PF+rQA3GFjKLfr4LRqL7hnun
fLHwWqD6/17RWsz806vYtr8isoMH1acgGy1iYNWFXSRLBSA+x20JQfE8ywo+/VoX+FZWqDW+uCIi
u/H24n1nBJn2OVnlNSUHy74C6G05HGtgrI/qZFktxftvEvVtdAjBZ6x/LxMAsPhd39fnSG+Lhpiw
Dv5EC+ZJ8A/U/40qPQtydkk8RIoAZSF6+68VonB9wqmlMudsfepyoAi8haLqfkUqqwpv1haEIjKE
yK56gP4/1+Z8Em3vdC35YoPyg4WpI3q+B2O5Qq26KeTM8h3BXCY2jY1XMVCGzuj6cDQymBX98PkI
UG7bsbaG/9AXY6Ml4bAoO6OaWkSy5u60y2phmwTY2apy8ot3D91QPJp+n/DlmX5mhFseT6AekjWP
/+GEeaV82E1/SFoa7aV1EdDW+qiN5Ct7OEU1bfdlcah2cnhG5WTTR1Xy5Vh4oDnxONgYvBVlRGj4
9rwcSdaQg9tBL0YTyTlprH0PJNNQZTh+xUlrTvlH6FWLIltxgItDxwurUhwdO2IZzH96WhGVJH5c
QCG931PCOwiVBW8rGawi9qrJBiY7C7RzsQ5UX6oEymnqb4hTs6CsEQaXsyDy9+G1wODW/aSkreRs
ce3HR4m80LAa9Fe5F5uWL6+gQjQF097gzi9REtEOvsMpJE4mwrpNmk+/92mDtyPhtW3V/H7Bpcaw
3HX9U2682luKFQt13VKui6PtqqjZxEyl2/Wrjyl3zIw/+Tejo1G49Fy6imKxA9fZhbRA+57n/bCj
EkNyhPZLX1pbAIlsAgGZvnlG48NJoCt4zYV/G8iL/CYeTagwOzftfz0do9B5qeik/9bAGkpr49D6
9hHImix/93Vzp1u6oWBYHtK4WOtlUCANSA906EPfzTDX436BpnErIFZUw/YZad8TEOwtOrOfwmVS
6sab561mITTAUfG9AtTmKOlcjqnny2zpWc8B71L/z3z+TSCGa02ZcGmPTXixCSGeUD6v7dZ61bK1
+gIBtniH8S2FtACBsOKIDMqzdFIK/gvU7pHNmv99v3GppnJ24JxDj7BNVdPi/q95cfvRYl9890HT
0CftpFEMyCF5iTGNLYObyF7u1jsCsM1STEnk4IwRQNJ/+yXzK7u1dumXAlZdZaMyCRQJ6C1Fv/Kj
6AzxgOffLo/npgHQU+EIN49W7Yh+AnAdkcrhfm8Mt6EHf2nvCQPlZTgvcJ1NhAAyVmt0tVWEbvFx
0SkRLrD33BPePze5BMVz/icg/ckfN7xmeV31NtaE/koC6gxUQHWm/wFYcKDBmE13x64dRzCui6I5
MMlTUdKtr7XZF745p66Jjk581u6igzazst0QfpGKyCyRx4OKJwzLOa36uki77Y6NQzHPID83V09n
c5vkZX8XFtbGAJf6MQiGMkCdmsvO+GKkWMHnr/AgHrqf7I52Y+DWBEHzMBCpav4eYKTZyPm1RTS3
luvxWdk86NAQbgFgJzZRyg1gQXvVlG6BUyNFxt9unfkYt/IS267UbNMnT6wldjjvGZfR78w62uMU
aSf7iaPZOEDYaqDKgbyljOTli/vJV0CnNhs7fYFOI0WcNDgMZ16fLsdv0Js5Ra1k8QBLHRHhzspc
07ZSVJ1cJZgLcMESwpdsdDVv6dqEp9nK6/8cEWae0zSEXnommlAZUghy0mZJiW01ZD5fSlhCIFx6
E+dmri7Sdj2wJRFVQudMXMfqkCxebe/yZR2roOVi6Zh1XWFFGYtdJOB3Pu7yBLEY8PyfgYEJpTbY
5hn062n6P4CJPCWfBpbuzGjNyGld//ri74LBZ/AJeFRw51rJZUUeCZIx5XqcruoWEnMmpYDb+p42
c18kgzN7bgZytheICZxOBGo/tpYSeaDnZF8J5OKPRNkUquFByR0Wbsq21T1Ii1NUH7Gbr5UtJ4ZY
nHnHzFrIr2ot5eZO8N0nSmpim3rFd705tbhLI6RHW5YEgfIfc71XTYPDIDlIt73eKhnjI2qlyY3G
tP17ytgnAtltCHQWNoTrYxyE3IXROdgb7CqWzTlcPaIDRQDlIc5ukgTsSv2uw2Ga3JA38pNLjqk3
UdKLizBsAIBTs2bV/GCjNaecb2EE9nelBAQKEZkx0lXqTP9gNgW3QhpJXgVOWHKmD9hnuQ71CO5/
HCfPXWYG3m9/vXE3NwGAsIcnJYFRYhxJLSu/69Q2gkekT/fft3RFLAP3ZsDH/gYi2aJQgiDAsnul
N0H1gpoTGz5SH/y72cNC5p0sqmsll68fWnk77gcTb/BovGBj3Somtz1bvgvwWNiPOg0zZWcIlUmz
4EFnK0Zij9HJ3dIUCRVqghYrpBOdOUGM3OSULiMnAuiWNkGJydjAXhgfqc6jjEA/9pGKf6l9PLRy
RzLDKV0cY5k5L2LPhkjfUJViM7/KRIJmWJwJMQXmcdCo59ihFmJNGigxLgbuNPXSMYszRyZGO9T6
FcvyQVtNunR9Pm4ExWmH5dtQDK3/J6owqHBC0Z/o+4fYjYkbWRjn1IvBOZXvJ8AdHwHFj3G9ePQ8
B5K1NxConZgIXIzN/06iJvVhCV/QBRyD9HZ3JXaorbN/QLyYjMmdEXMWGoxQQUu5FrR0mLzlp5zC
MGsclIXBfFgLp1zV5oo67JyDooGNcMQd7utYE4Dgsz6nG5/sL2Dq6yO64+iHV73EqZbLLSgMeij6
/QVRoFBPZHUVjsbxkg6QiusWVwgy5rArFglomakORuQeAnlqlxXz9qIQv75TnbIuAxnicZrS2Wsn
vameTmwFX0sLEA+eQVYKDloRjxveda49odNrdTq1XO9Qw0eUL8CsythZHnh8XWrE/uuLSRKNCJj8
2ZyHkcA9y7xMR+o1p9Lwd/kSqiBEhRb8/roek0sQXPAdMmCif3tu/kFhYWPV2OAkSoj0OnrWMoDO
LsA0SgHJ4FFlM6JzWXQErx9+3L7ygY0wTSgckgVPYSAbBjf7hLhxCKcvPwpQdI4VgEUT2HVGyURP
rdgZxPKMxti1Aij85+nslE1Ma7rjSFe4Z7pb9oEaTSxJ7DJBl3RNWHy5u++p0djsvHayRL1ONZrE
EN5aS6qEbQoBvl3cV5VHJxFDCUOB6Qbv5UUk0bAJaXD2zqQO4IWvScxAM1Yvc5+JWokDkKJjUCvu
xZlccOaYrE50hzxCJ9mVrfGjbu9ldAlsyrb2pAkCml5xPSzs+sNdjHdzNLANiuVSHIj4/yNMhce3
F/MHNjkF7T7DOy+00mG00N/4M1wCd/0rMJL7Ad2u7VQlatKzcF0fxSn5JQNPFaQ5YYzMIEn+P5Aa
ZKu4OSdmAQXoa3+upEJ8CDvZxzDOQhgPiAdCH6YFIXDy+MbNhZJS7Bni9SDn651UYf+VM9mTd6Wv
cUDhy9aQ9kLm0chg8udTbhQwmyzbuwiomzr+8SCE9cY9BXk4sO8JhVMwv7xNpzq50M5VEv66401Q
qcQ4lI4ibFdt6DhRoncRX9ZdisjIx/f99aGOs3F+Gmpy3ajUDcObNPsxLE7eAKMPUj3mv1wqepZZ
W5tEwOudW2XrdZJEvl4dLOWQ9aPqRYel8ZwP5rlNG6Bt4ksUaIrnvRNmC5EfxfWnOhv6r3DVRyu5
O9i+7Tviu6zN2VJLPTncJBXl0oQX+afDjeVyo/ZbPWtArwVapLSdMbFSBWNrec6psb59XWf43498
gmabL44ghaFw5b7nGLqt+7n6OBP0iYhbmX8+9utRh4JRLu8feQq4xI3ObnF9p3G3K/6vNpygQdKV
q6/+Oen0u+4JOgb6OLx2Lnbpbgj7pdTVg27uEDNmxkQclnV5o4p+Z0XxEA1ysRKYxEqo9ajAfpxi
/Fk0csbE0zG52FL0kjsiNfc3hEebP4a+QCHskZTxjEXuuqRZOXaR62Y5JPuwA5NEAJiFYRXP4CRc
JuX9VHCNrNG+wuYTzjb1wYkYs7kKmIKA8luEtk9vMJqfmhUXbp+aOTJZc2XbGQtdXnXx0WhWx3J/
sO9RgpjRG1Hru54ZbH1s3hp3ziZFOR70SF34b3uPxg9YUfj4Vi754kX7Wtg4KONA8I/zlpgsGgrh
lTgXYZpUQW/H/1rZKNcEh/m7liKJmILfemkCgViMZ0KqXFzXXiZjcyWVGj4Rhf60p9JAZZ0kV2pb
uHODV70a7IoGR+EIq1SJnd2fB46eM1oTQUH488Cta0X0XDPdU5NqZrBnl58iOQe3h+bevusD8lpd
0ubJvmsW3EP9475lxZiprdBx6frFHK/ZXjflwebwAUlAjObuOzDYFGMs8rftWgWh+09Boo9nnjMU
03sYiekz+nYgnf1ywn//6krUFVdaHR0hAXAnkHxF2kL/WSBz6QlkwiRk+H9MzCFXK3aCWH3SaHJl
RS/SN3CPq8nUc5VDxfjNNUVz4fRIASMLyLspMXwBS56Qzm2OGKzGD6iqr96wpc3sD26R3YvwNpAX
G9L9HsSAZsP+j9mMs58tKrySiF94SCzIVPLCsBgAqTz1NJTRTQWzIr3qT2tyjF/lO/G0aEoFwA0m
6kNgG0I7+038QMeNlcNRdQM1zFrMeNsk5+P67TM9oE/h73nZ+YEZ5C6nzqX5gq6LJuSVQ1BVQqAY
3dVmEX8ntCDjBjlwgynwHr+6eB/1m/TvlwExXPH3qkHhU+q2pSwA0zW3mu7VYVadqoPs8Ho+wz5L
FTHZa4O6dsqXkBz5ZtzbAgNfwHnMioC2Cm2oC4IRpq1Dcnr1KoiVsRet57OzBfYdgVxEHAtzvzKc
OvXAM3LDgpgVEk0b3QIl2BC/41oYShFwwhhCvNFBnbYQqRbIvYLmti9BqJRbc0KWD7uF1VShK8l7
2088VPT2oYCRSeQEPh8hlDo+pBQ7bczO9rzeJlLGcg3YV/aF0sZRDQljdEvsCSRrEe1bjHhzbalg
g2SCSoKwuKc0Yb6bg3zSK/zA0o5tU2sMkZXcUlkhizqVZcrIlPzHOYs2fMkMo7fQY1ygsrU838R7
DW88wrL7Phj+u82SsLnenoCT7/6ChTgPzROOJrEr/OzWm5ztOlkAywCO1rgqatbzya1Lf0qFATtq
8VyUxzyuX7FnZbznB/y/GK2qN9Tj0qGH/NOQPEsLPkj/lShZXBGYs+AunoCynIGTESnapc83pk6B
MeDMSCl5KNsreHxwFc1DQtlye1vc7vPEjjLZAUorgR7S5dUkUi3gODKg6iN8k9kGjfnUq3JkEmW5
KIrq2NJtoSJlfG/stR7pqt37nUXGdoHJ7VeOGwIjhtCWR0I7MP06m3aqN5hMmXNChdvbmBneAsdh
4aoyK93dZk/qGUfCuPM+RPfeRKxRaTQFQpao5DlN5hlWvswGGM3LZvderOj10Z7HCG/U2fHhchY1
l1BTWpYk1KkBXuycQsK0cNYZEf9I3ViGlehTHN9kPACEPutava8BQzTewVX/Jwz1W1nwFuzARoGz
quGIONCNlX0aP9VmBmZ4iJIUAIWOdvGqzUps3IYn4wkXDSgL/ncyGW9KOSQtuai8QCsKo6NSvxnG
YcP3rGWmFJUJe9TlPIuY8PRL5CvFIJjrU5ZBsDacvXxV6Usv/OAJg2hlhpLv1RoYSC6PEnzvYxre
gjkUTWnzdL+EWOVBZWP/+C8S4pFgw9IACGQjHPmnM5UsMOBaDr1ZGISO7ji/RoxxdBq6XGABDaWY
KfaDeZ2vO9egDvFwRb7OxlRdRBZRrIxxggNduDmiH5rOPW67Bvt3bZ8UV2rsjK/lQhCdoVJBREF+
NQscsicNjxC3ljYGOkbRpLMPOETvnOahIlNFz69pAeCNRAf/nx1rw0iCRaYkS2Xvp1g+3VNPqQ8V
mMULVknvSf+s6iS6LyrMOEFGta5BmpxacxAAaSW4re/Bnj7a2QEtwgmoIRoxk7CiwGrO+cjfaGs5
L/aN9bfoKpVd5YcpLurhJ7wm/evhVhl74fAZWHJTpOdI6o4etigzOC3JhSCAAQKyU+ryFBZtH967
7UgTPauUb8XxdDXls0RuGetDPxxUVSSXRNteyEPyKShszijOJQQnsyNn25yCk5ONPIwNPwgrdmcw
Gxl5Iex5Y02ENsZ2dNqOEsQaxKTs1f1j2PiEQvaFyUtjooqw5yMv4OtFhL+M2TIpmepoDZeNPAU3
HSrrPBWAAJ5l0ORwS/Z1JZPSK+bS62hHVqTBTINYz9uR5NiBM7m154tHTTg7G+r/6DAd5yla5QWY
yv8qd49s4rcm1lZGTlK7fVC9NomZnzaHvRgdZTCpX8/ilXNaU4GYwgBwJoed3/i5wHYO/zzb5Pyf
okJ357LtnQtAMbZvVQZKkdVVJ/giTFtXS9GlRIP9T636qw7/60VNWBs5v8izTHPWMDJNeLJMez9d
Q/AB5zAqpTiUasMbigAYXt+mE/gLAZmQt85a6LTSOYQTSSbZGHNFHzjkvzrg87MbZQRU1zaCzYV5
wb9PNdAjQ0hWHLPOqot/asYoPqEhRmSWaeJ1HkQfuI9Di4GHqPwtNmH3BNgxaltTEoMVcNLbU971
DbM9SPMHkUGtG0+3mxpPF/DbyMMO3mhTr3Uc85cXGpZbjvDvSGbOV8OVRvzeOAMld2FaOIDt0m/a
hJEkSUWwIyav79alqgmfBaUDA/72c3IIRzVZE6LBih+XR32pNtp1XukM3kEHgwBaaQN0qcaPlut2
16gw17e47RMDcpli6bDUnDJGsltfao8BU+oQaDYHTHWhUhE62TjvfPu2fLZV3DLNRkEiTL5wEIV9
BNRbwNODZdaesLN/OOurs4ftuW0EQAcrZEr/v412kQdjGjHu6DjVVnpynTbUBdRXSly8UsnTQW98
T9S8mifggnqEjPc4/na+8f43JHYDsTUkTXlzTnCfJdalfdkWcCve6DARqSlH9LJ4/5p/PiuYVwRp
H8XBS44WJXNS5qirMRktTGRJaBV2dgG57ZwGTQx82s/NFdbDQ2YStnApBfyDMSPGFE2LWT41sXqJ
bGpG8EfDcmdrHpfYS3Gt+osvhLFFEzEheCbzZV3x2dKC1qz9xgxAnB+M7enfPzQyJWtkor+MlmIY
pdmenQTX4v4D4gnwlu60kYXuQmsHYaC/ZMcOun+S1K2y0DYiVGLbkFIFt3lq4xyp5DQ3Tn/of5N9
gMBcN1oO6JcHQBtUSfqb/t9Od2JOn7xa0/nDdDYYSGmBR8WP4hN5oHt8CBinBxT2r1VlxsouD5j3
u6Uuyp2O33eXRUUbR2JZbR3zlbyTTJ0H9aigcoVE995y9P0M7ilAfalsUrwc1SN+Xq+uxeEF4grG
Y6imlk7tGo0XZMo/w8RZ4jI8UyUgIVXkCtxA6uElwyZzoJnD6GH9leOvXIdBTvgYs+IYC0sEfvOT
POGHiJdgK1bGiRSeG2AL8BiVqTtZCBqrxGAfpJPQJsi4hZ6mp2mG3BvltonNJTahlKlB1ql9HtFL
eTmxYND4dpk8WUlpQUGelRdjMxAPtEjEbNK4+eINwkm44fTAPlcp9CKWiYmy6jaE0spBveoyFahV
8SyDNfLlVCkR38aSRYeZufINwHPZQIb7TkIXYwSkwtVM+/t1UHMViQVCJ5NICTVUwX14jVpAT0Ao
wDYc6PEixUSbAJEi3jrAfpzM+z/vvB5JE77iqxRYtjguJZ94q/+oqDFWQIX7NqLCo0AiVbmvOmhJ
A5Hva/wcofoLtRwWgBlFqaaie098TW4d/5W5HcGns2xAYv8IZ0GvLAOcvtssB3z0Gz/za6q/AH7B
k9gfyyNg/b7Ici37tkFxf4YAXNfxJ4Mrk7r6+Py57pnoeNHh9mFZ2IY+r9Kd9BAPyy7k956pflje
kbgRLxX7U8g3mE8leDt3PxuWVHjmAtEcXHgw/P980ggkts1FFFe6N2P+9DqkGk8+jxmDo77AAUw9
PZCJWfhK9OcAGXaDxPt7cOu1NgnWPx0EKrbzWLti1GFhMLzN/6Rd5sU0/MliQZ9xY7rdMIMUM0F4
BQQT7NoaUILMrSBCcvYrStOP3hghFUGF6OSjLKIAhZfT+lQXR/auJegdCuI2poOHMsAtg3gUpxdL
dn/5bulcUJ0ingU6mRcI+ngbkQ1xEQKdkQHK2OGW1W+pKVVcRVNUooMwI6VJTXQoQDTe8W8FZ4XU
mjYKW2xNB2tuW+TJS1WjAfszqGH8eQzBSeizv7FK9cDHkheEo8fTatH31d/vfcclmu/Os/bt2LK3
RXzEd+O05En/h/81Q0AxMzfTr9MxXr0sCZLmR7oNazp6Ww87mOF4Q88Avr8u36/nS8oCMJpBG2Ve
51wkHpfyucAWtsUiWJgdwJpcXHVR3hULCqh5tMcud/aechEDK1kbdEcG3veJIQlLhRWVLIQ1ZH+V
eyj9Z8EV39LedC3qi63wT367bpuLgTA83Kv6hrl0XEAHPheeUKmCLqd2u5iwZrCe9w/dFoi6CK5v
L3MXH1QWYS1BhzDrfYaW+T6WDD091NvecgiJP4zmvtqT4dEhX1iF+S23rASfKPUEV0+jqB8z+l3P
BxmM/wD0lyHwfKrM5j9byQm999d/N6jGiAnD86ByJcs5HepCLg4XmttFuPkNcXWeNIZZP+E2mk00
UNU7ghrv0K6FYOK+HMmZnub2RrNOMSuIAmgNADwXBRD9BOr8esnAFc+6B0MrVnVCiEcSD/rMFOqs
em9ktzDW6nLEIPsdhRklp1gnR27owLPpfmE5vmxFT766wzEliQnYc+987d94ruMde6l21Ixrdk/t
qXkV/k5WKtbQfqi9SdSzPWTq+TwXX+ivSBqeK1fQyR+rc1SdxNHk3MDnsi6IQyd87Zj5W3sem3f9
9mIqQUQrgOagazyJD8cG4rb2+mZVU2Zaj91vzPHrkTbvOuH2zZOluCA40yFCQXThB27nosKaGT9m
QpYJNW6Dosu489L/nM8w5mnkSVIfrOyNu39m7SkOGmE1o2JoKuIdHjVxFlj9zA2u6kuV0ybESpbL
muVC3ElXPgDZl5VOKJ3+9te0wRS/nedwGjTpS8UbNauDuxKaWLSh7Kl6Zo5dY1/Bs7XlI08Vne+/
tV0sUzBe2gwJFYf+zJIs7ugd3rHyjD8L4fo6kPtupYNmqIaqavDP3gsuioD6FMK4Ef6siMd7ZHxJ
kWtkfwjQLwVZHzUesii4X7gdvn+lQWiBVZsJGKWURHvs7YxqugGE/axD1/W/eonXeYiixhQrj2Eq
OUcSTEH2M+uc0Z4ptOep3sN03QoNO2aydBHu9lwEOPrJ76DKqW/QXuEhOyuah1k+Wlo/UEkTLWlh
8LxJrMzoMUdgGcaXmKKxK4oEcSqoShYez/D3MgD6QsXQbVtP1REG37p95ytT556SF6k2AMJCMt+n
iE9KWI/P6dntOuzl1gwqYhcpSwkz+81zHIVvKImT517VCY+UB1YzNhnyUnS2oNjyntD/ThmgaQcD
oNawqs+KmyxrbogxodOq2vrtzsdF1Ug/gDAGMdsMXR67inAbaEQ2j/SAIw3jMyKl2+jZC0atu8hI
iS1tHxRO613ITl8YE0JoQP12gTEr00VEVWFM0gARe2hC37iYBSJwNp5OB6bRRKyxmlQiU+f3kyfF
H1zK1x/j7rJke5jpOOsskXTgNL859FJCXrKVzgBh8sKRouOeIcDrh90FWyUGQhfbPpMYojlUNUZ5
s1h6pzhXDZeIWGVlFnpZmoPhanXCdUWddyp30izbOXKuoo+ot5bzjI5V+qwaV5XVEDN+V9lA5WMm
Z1F9E84rtDmkgJYZ+qAqUb+7jqTIrNLoorkuJxa7u0t4V1Iukm7Co/UBYuyvM6/HV44DWIw7qAoe
r1XykHgBXdwsitXMd4Q+oHU/XMq6sonTtEetnjgPICol6m0FYE1q/fc0OAFjxiMA9xdNcql01pQ3
8CxSgJ8Ra980kAwP/sLuoXlrIBe8D1D/5JY8Qc9IJOXNPFvCdkwaGrFWgzmE5JJoTXvUFO0MwbOD
yMu8fV1ZnBTY6UEY7hOQ4rOpUvIAKU3huBL9yKWctucy/Tn4YJXLo7RhHPjRQAGQsFPOYqIbs6wp
DG9/M5wKjOl2elEGIQFkEOLpMjFavvG/3BLMI8bvE7GsrhNrbkuoONAPb+KMBBUKQOQx8COMAVCa
NgTomv3BnQsNypmOOEYkIbjv14MRK2vrBLIFWnDpfo7nHPND4tpr74XZ8jqVmVniiWeE/reN++ok
gx+HL1Qs9LUChDjhDM4d1SZLcCEk9JimIAciTzs+GsZsuMEc3YlTORYpP8nQcudewlX/RDM+81s8
2iie5zRJrn0HQNFbsnb+xwPnB5w+ytuXP3TO26Bt630JvLFdy3golirdgc0OclA/vr6YT8BNwd37
jSeHj/TCKp9+XDu/VKBVSAK9BAa/lelUdE4yX9AgzDmy/i7QN5aUySxNJTfZbDf21wy+gWlYF9WH
AsEi27WU8UPJhww802JHyqOf62d3zjXpBBd/axs4/o+XuiZMV+4CTkqeKanLYIv7SIYK1ooRKRyS
XrJ999lgyTERlV13RhfETm4k7Dkk3GAYI5gRc9FoY/vZxrQbvoSDDf+YpKaX0PKYU+TXcopYIHeD
6b0uUifekLjL/NDHA92VcqT6UKWt4pxL+Btp9i+/2LIJ4kwY2kQ0roBBHxHTgvzZEkG1OUGTEgJJ
9gx5soQ2ITxid8lTWZap9Oq5Miw3I9oldBj9ouwiFig4qgS3SQyaWuEDrGqFk4kZcq8dxDJu9QBI
k9yiMJOdCaJXI62XebLCV7WEOY1wWBErRpvXyYqq9SNoVOkv/mNtgGSkxpc5NRyguffCA2wZX+re
VaC8vOaGDYW3Cl5ztqMI3XjWbadhcJA6WmgMzWSkAnanO9Idf4RcIy+CFjczNlWMK13p2WlbvxI5
zwhXP7WYPvfJ2khsKLVCoTr8opaNrcrYvzl0VnaAAOTT+eNz/wqV0E4aKEbaaC3xsqLjfPtawdxu
kNa1WEsUC64qa9TPzLZybhV0fXdg2Ol87IL3EKJxTvyhzKEG99SMd5flPJHwizBBPP+RuU9Ua6BH
Jsp+79YPUfQonCI3iyT8SYFIX2FHUNBVWDW/dnNtjqFKJETh2wo16l9T3OSFdkWKovrIMOD4+Upt
rTymvTb0APBM0o77CGwtu2Tper8KF2OjFaqqyfnk4U6Gq1dDOmHL3+xO6h399wuCAhfnNMjtgpO5
DwZGm/tb4uZhIFfN4x7zpCYtKPjQNkVCUANv1xAfCqbl2pD39VqrleqVoJoXwz5Q5R0146akTC8w
s7FqplEmIQFvRhawYkkfwSQGrvNIdZHPLUo5TOKxwHgC9wqk4DHaheewXUscxFt/OmgaoD+YcXPo
91lFCsUy0FadfPTj7i1ZC6u+aM5jGx6BBw82VkfclcyCDvGZHg7X5l1l96n8r3u1ZADDX+ZpyQpo
XUKg6wuvQR7OQ5UqDmf7dgsN8SIsn2PfrftofV8Jzi8JcdDr/6RoGbp7kWReNOUIJ6HJmIWWc+5u
R1Ji9FOViJdz8KYvij0zDlNmHFzu/RQdKKpmbpeLO7kISptT8skIbdFZsV9EiaX4+xx9xgWy8WlO
IQPXlE0qfEc5Ow3Bnu568wGUA2uEPfcJSJ2nGuQYDg7Ia4lJLEYBK5/m9k9oN/cW6n6HeziS+T6N
WArr3ZASAqBuFE5UyuJ6TLELG4sSWLWW+P/kPGeamcOqKQI2EaFUdKvT8RLr7Qo1Uma813LIvkL8
TS+RI1TD25XVJmUd/dlTOl/BBdk8l04fbD6PxmRxMmlJCM+kpP9qdgR2uFRZ7W8AgWCrZe1kox/5
xZfrhrGkhFyJG7PJVGhUfJFLQI9C0ng+Xuot21iNYWCvZCBg1CJ/pZi0XWuZFARTZHGtqhhsBiTG
HlH2l8LGxRLNdvTfFZUN9Bvqq3n+FIjyQGJFr1jg3Pzpzqk6kF/z9Z/kyadK//iL11qD9YLZpjTw
ZndeuilBLFy6U7cGKwkmNi0hVKrVnKOO6NLFQLLJHIE2y7gyMr7NmJgRyEiHvBRw/dWm8tusmCWS
NBJ2Ct4po2clGMZAwJHGoZ5pal0xUzJFR1+rmydaUZuf+ycla8pMtyGOy5W7pw66MHfMbIFt8msU
uir9jA/xYHUSnpjMGvhXWX7/nGVmsXtxcBUO7xxvHf9hn3x6lDcqyN/WUzxP2O+yWnHRPMwL3gXG
UiKf5Rx9Zp1nn/niQEfx33dvQQNez6gEKcV+pxspFg5b0ql+4MfUS5FWpY+j5DzxudaaxOiUFOuF
5kDaKaYDl/nma6U7I2UVF8f6nFJMsnBeIcGqwLamOOy9Q8JIylwvfpXVCekMK/ctPedUZe/fFVNU
cWkhISGSpyDyyJkAb8WWZS4Ez7MaF8EPBePXUlpu/UYAdw5s0DCKLAgg16sXXqsOhCYM0EFKL24S
51WgEvTVGkG2w8/ryMJzWDfhg6IpvJKJITzn3RruPwqn1OQ7vt7XYM3oIXbb5pod7w8e+5kryvad
RRxD9+Z6ynUSaK6JgInZU7mQ5aGmsV/xf2qGr/LAhjBZjNLK1cuIOC2S6MnXnECuRymY5cikmFOq
tS/uim1SrysmJ1x5+noS1nymF8YyhIz038l3gmLZwEBVRT6x2KLnSlO4qZMi7nreacsT2XU4K2SU
v4g0ZshzB7a7jAXG41JHGNoQMzPQiQrUfWCVgq7m6CeyG6Uen9TTAC7pW+gUHguBK03qYbUK1A8A
TGuvkLKauPljungKlHNHAp0Ez2vbke9RHauWgb6DUE1ALxz5yJznnsG5Q/FPXBsVrVN66o841Pof
/hYQQfebPd0Q6+ve+fDf+8wUORV+KC5SUHuS3GmyD0p2Lkzr2zTcxu8IBEten0Bt8h1igNXdXEyQ
GgXHcT3rTCeRQoZ7Qy5kfnemyOonQpMLnelkEgJBcWXNRuiNJfv252kSBN9AdplB922CD1270dFo
632GksMU365d5xTAFNOCvBM+I+we57OZ2OCe9bkVFnlMUv4AvyG1hG7gwK/nxeB5YFE3ok4GxgxG
8zJyXlkTH0QZ5nzVjyS+x6ulQgOGwP+Opo/C5AK5BCxmYxDXifWxJDWfuyF5NXATdvXZ9jU1t7vk
FmP76NsBKROjD6cj5rAsvbL1FojcxsHnJDwiOX/ZAl9ZM97NbC05BHZzAaqEgVBYQ6bpKlrx9IMF
GbnpOQsM0S4yxqLUcObT7gMSYjyUUTUsVXR058RMP71HaPQTdzSLIsyTlwjSfqCRjYMpibY0mY2b
grXAUOBg34eLC5EO5g1StuTRzoZ3CvYKXPO6/R/YmxmYLzduLBh1Oj/fw+gLehnFeWARO1hKpyI4
HGszMnIl+Q7Mc41dK0PaRWpzO6dYTRHu/5K98LXhWIoqnD661WScqGFvgHWkkF++wuNq6V4dnEZC
Pp+TSit4HVUoz+2cunR5VR6yZBtw6TCaHb1Op9lSa1l59BRR0JRR4bNl3rbLmJN+pSXGmH3lJ6J4
ke71YK9iF1fbD+IKdc0T8UGPT6/aiEeqA1I1xbEKgzTLnxdgSOQ0Fcra3Eo8PnPpH5aiXhbE0Ek5
DqBdEvW7aDiYwJLYL6/uIHchWu0nZjZgs37X10UppihL3sM409/Y4UnXKDH85Dup1rNA4E6VHhn/
HnPbQWpSy5hSus39nKUf6boyNhicyHUjdppE4g8cbsS30xK4vRB6hiua1b0umyCVUHu0rYaIb+cb
9crcZ+urphXst46Htld7rnj3xgvVqc4w5YjwxJmAqIosCpOk44Q2aKZxfip2+ywAj4/cVzd7CfM3
mGH4zC0jmFhrO6aWc/nOeUWPJJF/iKXwpVcL2mYV70Wx2XW407RY6UffqwB8LvlSrMNcIxG3c1rT
76jXM5OpWSUjRjpNpy+gdaDHB49cXyt1uG23pSFb2o9QLJlwW52D2zEQ8ZiyOiCx1j6KvZlJKT31
Gsh9o6jnbK9BKy3fn5a9bOiQ1McLry23muIQ65qHrnn4WtwYP/LiJO24Nw0AL6p+aRI17Sg043wy
Z6UaLTozBV0SKZq6wVeEfXs3CiaEJ+NnGxz7TGsSb3FdWt73Fv80bA07qWnXXpXn1lDX+dMinEz0
l4KWITYKGObdWbybHnZ/FalO8r5b6F2V1yeytgOntBON8kHv/sKeyicGoXlvXwRNhVh1QzQHotIG
YUwqKMURA4VE5KCkLqUvZsPUeg2BYCW1ssv+263LGW/6ZvC99J9XtRWDlU8qsgJGeUekm/20ORj1
Oecw84NboGf8MgomKer5CcR1gHXyYA9OvzVkbkNMe2rmc7HG3qzaSnYpG4igLNPXqrLsmpWkEs55
RWmZih7ggWn3GJP6JVwhorxo+oddO50jeHC2InF4m/OC/yswI3ehNXjzLIZDDH5jWSPchdbZQGTc
pbVg4WSi0KlUsplurnv0FIC563LAvTnNGuTWRENH67qsw5bidAX1YcyxIX3gTm48cDfrlBS6JXRc
R6JxU+wT5Qoi8nm5+kMLYafcDo+F6mafYpe5k4kZ7lYWtScr+cmc06DCLyMgVtmcEfZihWf7sxUg
kV+FEs/jvTBXs7v6gG5UxLTDIZFNUvCHKE6naBQUKaon4KIAfuVRrs2NG3jj7Ky+O8FWcAafMUpk
vG6Z29ZzHY/gtl76ZXurzdESps6xCK6tgQASoeZfGyh5tMUyIjKbGlDTsxPTiR02QUO15f27jfy9
27LLRXMxIWpwfurd2AFDfIiDiRVNDi3X8GLE+YqkIWR8wXS0q2D7ELckdD5oBaPX9+OzqZrJ1IVe
sRNWeGu9xusds/FftRk9rQjcJABnd+v0Pa/EA0KH8XRNnNg9xcpv1tdNPTW/bhnMPGagdPChoK2u
VIwpGr52cFuhzz7+IWpumwNmCF93GXpAb5pVbJkN9f/R3T8uO5VqINx7lr82XVMYqgJL5gMnxXBv
8EK7tUt391ENMiepd+8m32knvCq63UbW1St4P59bZX4LGYLfNCIyrSxl0JB1maUJJsUBBvPN1N5+
HgKyAeWh96Z+T5+dP3zxz1CBMcyUhNyJrpFOqKxRGSgkqHgXccshb50pjpofuRzRLYD8Mdq41RG9
QMZDJLJ3zmBdWUF58avM3BTJT8D4Ctn/bXxlNPnjq8ZFs3cJ8zGcfCC3zHI4S+wgmBrD+YNcWXen
DLtAqg8vDFpj0suiVv8j+iqNv9DBitCRYRjGwl1NhhrvfVIrZQbNYgOkYPZ/SDBv2kRfKIskkA9d
J4D7WUXe7EbkJPl/k1tHxMfGGFy4vJ/M+1eBT1PXmX5zE8TuUqVj9qvHKhpa5exp6K6F188+s8MJ
sfXSXb3/ILrbJQYz8ybma+4ygOIjyGWQ7UQe9oBy6hk1kp71ieaon+BgUlH9nkWfRVh92EdGKKEA
ZULdJyTdRBUmkL45I9ojfPUmg2z5h42L7IbKmicDuXmyGXmRJ3aaIatLLX6ZN+Puf6elom+I7sDD
JsFTTMXsT24tzzrOPH8VfX2n3SsUYxdpOVKXqInQjhmX9cUUQ7jBg23tNnvSO/mJEPn83n/ZVX9j
osfU9M0hYVj4eQr1OM3ehUu+E9omwzms6rhlHtqaf0IVhWVdImZ5CDdWa2KcMvso3gL9/6MKlpeJ
lJGymqLU3ONw7+FgkJXtfuUUU9kpWhBL7ypehEk5a/IqHWO+KIY0bcCFqMRSN4vSXK2MNGiBBuGx
kdzTkPZ7FP0QrtHCny4AEDkt03l47UF3Lccov+gM9qARfBZUD/fJY9RxKSxlkTljTunszneLivjK
h5o00DMb6ya79I2enkZ/QWm+lw108W63h5z04+G5JCPlPnsi3BQpjvG4isS7RRfffkWHqYdFjOlo
qr3cYDCLZCPA89gUqJf0h+2u6uonT8caHE/AqQQd9ehOjNvaaznuMeaVuAeCPGbW92XY3RpowhEW
iZlgKgtFg9bh7SkcGYunQRROUreuWeVTAVG2jP71LBwUhOv1WnCbfXbTICaOl9FS6mYRhlSPyTRM
E+St0NJMX3DISUj1Py5k4ZrdRKka9zildWdoSkb2U507u/GNxSuXQM0urxbyVT7bOChpxEP0yngz
KJOh6mM/Gn33x2deX02+R5ti12SavwsujFvU3tOKNdwxfwZ+i5OAHDRS3/0DxJVqwT34AlS7QvV4
x66B/sq0d8Q46Z5XBfiSUbEilS3cYdMTtNAb/uVmT1XpvsoD+wmvK7aCg+DSU0awmd0LQw0s/Ydl
0yv7ps/RiBVvdDnP+aj+NvSzyec0PGEee3tavycpsqyauSoRpaXQzsXqmRi8Ty/oFNPjNSYrSMQh
HxJ97SNxoN4d+K3Z6FRL/XrJU6ERhoKiFwauCfQQ9ycKu/8ZBKwPbDj8zSxD0Kl3tVdunfQ/TOvl
DM5wHLy/IzR2xrbRGPC7/k4v/ZqJFUHNYriY6lCaY5d7UAoJcUzaIY3ggrg8mMS67t+CtVE39xmH
4u0v0okownHd3/Xe85HLQunWZfXFxu7TPnAi3Ihmuh+lTFc2qQZeVd0JeQT7KBS7GeXKvDD52UXr
ypRrrSXuckZDdqZ9KL7qW9jIv5OktQH9A36tWzF7z6Li2bvYYtIQ+HDJtJheNqZMKEVAUiskcN5f
OX6m7Qz3HArYdrIUsbhX7Da+2L/Yqn71NYpAGnBZwsczaYEFkvX1AhKZAKTfRe+QdplEynptKa5p
MHUTeRwDeND79nOynRJuzaZMdEEvaIQPPQ33QN2rOpZIcmD1/AP47AoGLSoClvteX1BS6bXNb/nw
TXhaeHLwbIQN7HImPPXVFAw9Jl32n8m5hU4pUL9CJxbnMaYaUD45SQMuYQNeg7mcEst/HQ2fk7U5
t255yR2ggZx/M4Q+M2UM343e++uU0qkW+1INQ5/a26zqP6mvT6KRJGxU5gyy2uRuXvypcL2CjJ8+
jjmsm/FHNbrMwTfkyl/5zkeVEE3hn+R4KyWmFrwSp2xTijiVSQf9BNHb/AVvt3MiKS9p46hJ2o4M
sWGKcCFdGuhiI/sZo1XJyHumL8JiQ8S5eLaxA8ac+fVh2CCxvuw7mpwGOwb/RFUoEPnKVQj6YwUz
gKfJQs23204bdZsXWCcQC5oLqCd6gZaQ/5/VctnfmWMPMrau/4F9YjZEO2ryENx5cmazCLLrMjNR
37QtsW/6K5dsDyJAt1CWtYqlD42c26ItFtw9d+79qXhFG+NhePT31qpKbEhb+q008WRf0PZy5/D9
uDaDvP4dQ3VOZMNKmrQ+RctP8jnGM7Cj31OFkQ6t4npXMwdtPWTH4SP/H64GW2IfZCJ44uhxG6/o
RA51xnUf6S+oTqfv5lgDKplzMgzixg2ldEptJV1Lyl7tOozDSmPNtJW8A0TQdzXgyJVUHucgJC4P
SzWY/4B9HjY2z1uabArSPOz8fPmgYBcHpDbTr5eTK+Gj9DG2yocH5WwI0YbZgqjD9uAcHNXr8u9S
I/Lb82SojPJFVS7C2DHrRuMrYoB9MELSm5UNLH5nzd3MZ+lUh4GotNlkSgv7cnMN/Pq0/n6ooOyq
l17wpMc5/TXLzPeXPJzrH01U3HxJKHS21e22b4wyQ06AynlTzPkrLEYcX3P9dh6TZSiNDA3exxbf
3Lopxt1T1ccBNObaAM/EO1lKThMH+GTS2HN0p1qFRXy3lDHy7mpldE8u7nk0SYIsa8XLGQhjMbqR
l5W8S5pEzZF7tAwm9kM/2YjBkUjXERQVNBybeOQy5m9Sgu4JuOcszl5B/z2ne3oR4vgXYC2lh5ts
tOLKWAzgfRsI2xwwuwXFV+2FFQQehRaplSBQJynphk5OPQ4V9zeeLFoRCLFuEZp8+RMKeJJyw4An
mMe0C8bfANEQTVgAnNSD/QxbHix+0tvgEQBiEcNCId1c/hGDKYVhMOY2ecKJ6Q3q8Zv5BLFEoayY
fQQ1qWfXMZSXs9LBNivPbd7cOXF3Xgjmt+zMkTCJeY1iQNiZz+1HoBmhNNzrKuYRGRcIWz74yp31
JcTS45mF84kO6udtXOlsjPJi6ReS+akOT2awlbT5g2vLS8w0QCqWyzP0Jl8Mztaf5Ykm6ODbiKMg
+4SVV87WwsuMpjdIrxLI9POE7XwDmHG77DtBesCqwGvQ+mQeeJNlUwv4jFg1IuPNYSjZHqxFPvuQ
CcEbxKRnhO+PiCEQK3c12fHOw2T5O3lAqqH+EyHTCUQvaRAl8T8osDp244AXXXMOI6IFXGSVs2RS
0arREQermgcQedetNqFOgIQf2vGwXB9NqDZawpQthahvuLjObxnPZhKALqTiNUYHtRGQdP7tSb0h
Y/aR5GD18qGAxX2nnoklqRADPDOrWotb7SGrkdkmLRNd9NpgO2KWe6ThXrSMfNwFA/nk5i49wwRU
5QUtuxMFjqSmZYiUYZPc4qBdbAHlyBJuRqleHoguKRo4oG0EVKaYRHkiJQKz0akTqA+a2ZiyrbZc
z5U/8LBWakRQsKtnLYCsGI17GW/oejzvVpKGS0BqAgTOxvImeIO/vlP9Oe8YfLrO1Fy9424BlPh6
/ac8sDAPOrdYCEsml+wROMmpv588nx24Rro7SbTVSwqUH/KkJKvbbHMIuJGwzFaN66D/KqHVcLEz
Q3kUtp3/VIPgl3PWHFkCxvHijCeq6CIA/HLIBtJ6F1kQtPMSgYNVMpLtO2VtRcAy4J/MaH6LkrDR
0Xcbjeu+HKcP7Mx/AoiCcz3t9r6CcoE3v/MM7MfqO8UnEHvlUTSy4hkMLFQ7j8Ngv7ZCptJUbe2K
5fNiT86usqdvCWCTVD8syxBdhezOq0WIBQKkvSGRnfTluBXIWNSqiH9g74asUiTYidZp9BoSddro
4GcquCRkWYP8mj3FTMAlITa6ByVekJ+8QWaAONmAhM3yKox739mJXy4x6//MadcxmOOOZ2DLDlSs
8A6rmqdSLc67V68pH8lru1bv1xZfgPl+amijXDDWy+esEX2PheUOJUQxeb9AgbixRDpbd31QAVS0
0NOrj7Rr00+55HwwgORcNxqwqkmGi1gcbCZxvqjpJ9QoWnt+KJ4JBqUrHYudoFCSeBZXo2xCwSyz
74Aojo1iqRMBTcO1sB93ifQ/+Ws0nZx+++utpqDOP9iBPRYH237ToI0CfunnKvytEjMsUaK0ygrZ
LE0c45hedsB505FQdf7rs7bgkJyFbUTO5rIffoZ3PRDT1xe4MOapwUzFfV0uMdhJfVT6xTIpIYMw
z7rUEr6/RV7pQtJA8Z8kwip8S8c6SUfr51zG61r1O3SlGDyFdAANzCdGBSjgPV+iJE+w6yFCdiMx
rlalRyM5o0bKE97jBTv0Czn053ijo3hdKxjnxsAnJv14rX2if+m1P80aEZT3Lz+oQ/dtaxb/m7ZV
vxLUYzT/bD+ktY9f8pgJVsWvUU/ztOZqOx9W8/QrIYBlUyGpvzXgHBkUPAE2jrhlZB++YMpj2B2h
7w0dJsOqOUWCvUCXOtHRz16ZY0oacTU8ecvBAiRFTLgyzOTg6Q03jXA3HnDuGdHJpU9kUfwzlHcH
Gi48XfPwWBCrEnoFNsRRjKrHdIq1NKDpHn1iYTW+HklwxFWRjg6Iy/3fNTI+qaNi88SsBIua/ZpX
jWe33kYik5VCNO1dIv+NXXs4o0qwNECRhEZv/VxVlgAiESVcb3mbA9MzpCq4PxEUv+4TQMBq7Bnq
8rNY5LgSKgynSZuoWqC55hBTnaoxPSf2JKVDIcvj7Mb9f2pJ3L7tGsFE0gewcE1U67TSXqkYtIB8
edYf+TEetso89u4LSqxKqKyNR7VSk1JbEhpuUZFxxznHf+GMptrmVXQJsN1HPmlTXe6j7PnK3xXn
w3pDQT+oH1jcwE9J+boExBhauQQMypcbAZbMyCtWqnpU01UDoD48Oqr/gxrjC0BTGufNrigEtM8a
+NGNw8Ib/rbWNAK5qck5eenqV2eUho02wMeZ3X3SXlFQXhZ5YZmS68kjiBIREGrNCy6v4SvomChB
nKww2adBsYy7rbAuZK7J5zDLf8cP+p63pF1qaisuQVQgcHfc3T/t+Gv5gb28lQ8VAgsotUJxhtio
9tWIpZmFBMZ/OwLc1U5heX2ek2DUHQR5/BC5sUfV/1LYU2dKLyKl+Qs+mbvcdm3K5CO8FbzsH/6S
K5vKWXLDC1fG6VqlDHWBr+xDckLWY83iSSjhuaBeDs5deC4QI/JBo+jZih2ZtRVm3UsA0lhggxGY
YqE/suICVHl//v8x+wORFMiPieSvfdUX+QhPsdT9rcSO5uKOOPAOjKpF6UqIFk5dS3s4mYyO1Dg2
QCaW/9LZotEDOU+i4b+hMJYGfALl6dzpD2zwPIaEsY/Dq6dGsKfv6Pgc2jkvwGeSGQAjqlVdE3hQ
gHnwFIQNh4P7Psg1NW5loeDyNOrjODZHP6Cq9kuDXpeGZgx/L8JkEmEmFCKLTxxoa1tRo9FL3Xep
tHNnPaKMSk7ppB6rpw4i1ZojOB8LWJlnik5pgj123/SBFXwlm4Bco/vEWDL7D7QI53mBAKxDzZf5
yeuVOxsYwIGO/iNJfy106Zx7ghbrD5sMk7OWEDmf6P4ERbu6PlIOkX6P5NfzpHUI8nHIlV4JJD0d
NJu5ZcPoqqRSrfoCNk6uAra/pEuLWB2OUSUv2H9rwWLom//PjRAbD2aqAxyA9+BNZVH03aqWg0Xl
ff17Bd5kRhcDDALZIHgCVZjI5SjtV3y4Gshhadu9JL/u1SXV0YSTJmMkd0e8l8POW+xk9TydO7FL
DHb1vJj7enTzqQEJe6mQ46RKVKQKd9ewAkgNCFI391BZuODoYPCyu4RTEkJgliSTrV3vzi/ilSHs
xiFCBE/9SCTmO6Kv7UN7TJposIvIDhtVMGtWTplbj1qwKzlksgaefRZWSQNfd+NOjMf3bD6DwiB/
sCQq0ax2qnm/7qKK4m8wGBqfKf1ZpUxsmh+uXvygEbheO+8+bPCyUnHGL9KOz7McGg2xLxwUfmXX
TZQda2ysYdpsns5aRz7KjrE2gagjWAR3NVIMzIJqD069btMr/upLqQqc3QI48kGV9dYKDEU4HT7B
X6vNdNE7QbuZdmy4D/Q59/Snhe1fOQLyTFe+5Yz/d59hHU+Jc3RtkcLihk5CB6XscXynoVUrC/I9
i2Ma8RVcAIoXbMc/UNZ8mxaJbvHywwqy5azhgc61ADvL3e3R0gCZ4FSLUAsDtQBujAtYB6k2InPh
FxLjpgdnJA4xfF0Ym//PRWYQcoZaBsb/vCmOC1T4BV1npxKNzjMQxgRl2zdpJjf841nLNrp/3VrH
JvoUdW7lDqg9Oi/Ekg3fk0/qWtKnWwn/u7KJMCMB6s1alS+Z0SCY+Jt7Ivefi9ulM7Xoqwfi8kJU
Cd+gWCoGG/NaCw+yrdyHg8VS078TGRCY7C4lSN77MI9SE68/FUFfjpD/nNCYYlSGdXynxEZSdQk/
i0ZXsQJWR3wxE1mCKNarC9wlYo4ZqDmtak3CYLNGdUoyDVS//vpFcyCHsJHoNU9xY0sgwmAPrghT
HYvd81UfoxdFQFhxCYMGPZr9lXTZ7H/xSNd2x/gMZzqBHyw/BKM59x3mYUxx4xozwfNaSDVe4kxw
cxqUBt3r/21x7YJS2dgy5rp6LhbXFH9FEh7zTwWCiEepFyRpmlf1DsSgqbBgnufny9pkhbRo3Tu6
IzeIayjio1q5ltmd6M8GDjL6M0/vsz3WBPjtaLSypfhwSo4XgAqMl9HODeBqr81y1sSa9ZAChujW
M/Zx5RFaN4sABFqFLhUjUhIPGl9d4RK/eSx9s6h/IHlVaCVATpGJ3wPLND9AqpZa9PnwKR8jBwev
YgsoEM+JfSVg9n7Q7CImGsEHyh/oBIeNUMdeKIpCJ5fpynd0LyZWXQmzqCN3y00mxnbobeoLcSun
NRno5UFzOYOtigflQ98vn+4b2xL2eKH2oOBaGjcGxQGBktivACmwANOS3O9BTlgjOV2qUHEvQZ28
m1hX94mpBcX0g4MRaTgiZvr55Pebl/rRunuLyNsaafAxs4TggwsG3MStQHYFKxQ/83JZRmhRH4Ji
fddHzj95CizEHDEMaf3QMkBzQaTlitJYkov2MWG+YICoy4y7Tjv6We+EqGwl7fNnxck4TOkQnhWn
5+lylMImcbUv/18eLPUm1e4QPe2CnrS8Cpbp1877sUD0RB+qklWY1fGcEKYyA53soz9P69rAr1hl
CG0ZjGenYW+pIQWn/7D56XxpTr2MiK1M97T4GqfzwOy4w1NeWcXOGORw53XtuGDwDnJbuyJ05CsC
FQl+R62a046RnbmVN92ZM561S84p0tLgXRhI+Bwm6FlPmJGQSrZLo7k0or6f8ZKM2J01hesLnfu0
hKiWkvFTkgco90dTw0SYldZ5Wk/OJQvkO9jZkryUqvI1YYj0u2kTvMUiuUqVkedhUH9oNbQmxbec
RXHkBTPrQu9ABvbVjBBFHSGz48xYaO1Tu3IwMBK5dcpsDlwamBlkawXWTVSUuLB6LO0N+a0EPunz
5O7o+j6OVDS/XiTIpcigJ/XGOeclXVw48teVdvRiD5lvmWS2E/EK/qMsIoxjLTUgJ7Z1rt7xb/nt
OQbmjoLvgiX8+0kqbaoOLmtG10cK5HMh8wSFNYhDb1dEAh1kq+plncW+qhydZbwzUJ2bOWHvTm3I
wb2GNMRfDn6qgKfaxeSh5jmta+FmxG6ZG5kamdZP8kBbRCALjPRxifKO9kGAsbkcwtMga4H/YVTw
/WVHkYPp2Z3ESdTr1zeaXPEaMFnm+4Nb6fHBUQ2+vwgFkkk+CVsJiGp0MPQ75MouVAPcnw9Ah6/r
Uy4f4wo71OI7GRj/jiqEZn1j1eI5xOhnVwcVkioE72qNjCBKDzIAZNIogb5/f+xtfxDOio57QOah
bC1nOWWqHlu6AXUFp868xH3yX4Nm7UAhvdhHq+WYBu3ctdw1557iNCpSO1L0nTqGyaF3EYQRU5Ch
jEX+uezX3eFhZTlWfQf9QUdiMjBCYhao2Cmk+wwR1uLvWGIhnYQDsJdPm7HcFJ7EJrD/qALzoxqB
PG/k0CKR7JTK0jyE1ApcsmObr7QQv+6zCdrET+Ez51AxrGmQqw6dXscXkb0rw6ckGum4pphKgwnH
PzSb4iXJrkdOzJeLBGGe+cMd3SeBIgha0aGpb3CMpD+Rq69GgXtPOV0+HwaaLvBupC68obxVYaiK
a40ILgfqmd/+8kCiSj5MWO1T4l+xRubh0gMweEdH47xbqgQLtSB2XevBACt6iccvBdlF+8C3XK8j
l7N2Aed58i3CQalKvxFE2jrSTqZQl3glKEWGFqCKZ2MRqVS9Xsg3TaFyNnKCiD3zAx8KFCLKrO6j
MX+8rK2m3CiY25pYrX3u35y8X6sdGZq7fK7sTa9zx1B0sVbWij4p9Fwo4vylNUv2RMpFnMBKJMVT
eiAn1Q6CAKHhEHRfaEfu2awSfeSrHSX5YcukdAqVmUIBQiLgbQXjG+A5JQE8ucykvmYKazNmCyJq
GmAD8ySn6K49MA71fN2OlrfXLcXGW/vp0Z4k1DLZHcp/2BkME/d2qMIGUqb7MbaleDerkqUle6+1
xIo6no/aA8/XV8+3p9YbuiZPCnFtipVDNaJ/5YLB4gxI7rBwrgwvVTrrxs9FgSwfxnQEO8QDYrDM
lPyP4a8IuBgHbIJ/+/bYwi23YZnoc+cTMuw1L+0BgYca4Oqw9qw/0tTCaez5dCXsNaCeY9UGBggT
/0NTsADPYCIZEsyvnVFghc7f8mswK+F9jEFzWvvyIk3pbrDZG/HOMz5PcL4odTaR7ECgvQNFmgbR
xPoPrGMXsAZaotjvd80Kh3tgDY8KPI8SBam3WABuGvfW2i2daxgapkq3tJKsP0wlrynUOTO0rzSe
Tsu6wy0/dB2x7ct6KFfDdpH5AcxpMOVEw5EolMJemgH55bseEhUT+QRjsNKIEVmIAg0yKdzN5p0o
oMXvDd6EKaOC7aqaudVutmtleo+VphtWMUn9vmveCh4U8upb15JDV6FHQ1ifmeUKG/Ufa0OMdYkk
Is/+6EK7zhpKMeYK9VsK96mlS823h77yaLdPy8Um4S8zIIn3CNQSmTIdL/m7Sj2kdBYnb8HTZdvp
wOc13jKMkZYXOef00mSTl28zGzTsn/7Kz1W4MFXQjvJ28RY4gx3TxqeRNPLOAzuc/Nlim6xF8Qs2
EWO+XsL+14rfau2fd1MkR/GVml8KRVxbH9rtnh2aO1/GoGwQV2PHN8uil2tWhIwv/nDR5vpdSxHn
1cr3e4ypOMMpiOuKKU3ebcaMG4HgJZ3eIly4y7ve1z0kl2us50K1uHaNvjD1e+fwUMMRdRQNkQlF
iSDq6+sI0Nld9MwQaO7CGqsjbuOjaCpczk1KRJtKJQzBWSc6bLDWUYVN5vxFZApJp/8MB/YpGnFm
n7vGgdgeaqtVxgvFFUuilzYSE+fql5K07o0hKOhEY4aaJEejNybi2GFMDetp2fz5N3AJPw1LOtfl
qEGzp3xFCTiC2Zq9nNoDK22aa4vxpdX3WDSKCeATvkjh4ret1nD1agQ6ExnENziuj6EU2YM0ic6P
snIl1RfmaaMns+9qu0ZVTD4VpybV7T4M7mY8/Crqi+ZMFH0MIfuDztEftcd3Fh1gd1HZ4z+8yWKA
YV8aaHvapY2DjQejKIk32GXM1CUg+PEKRRaX9c2cdZDG38Ut64UGJoCb4/fbvZsmH2I81NPKPWBL
1w6DdSCtYpmgDkdf4P4ei0LnWX/mNgk+ZUfdaXOPCtVV5B5tSnqqBHCRcrFk4js0081ZJVH2eeW/
xZWGfLLz1JpKmLeRhadhHrR66JCbKhFU/kIzoR81UHBtt/X3DDv7ZB7m6AeAgu+hVAs9pW4p5M65
jwRdFlpn/ehYVpfUgs08pGUL2U4GsGF09fyDvAOu7ARgATsZv/wdtOL8fWi5N5OOiWv7GNAq+EGS
S4vDycIsI+U8Eb3VZoXx1bleXINW3Qekl6d6RZNcRr0ov36xDITjGIRRKF0i6WopaICeC9W8IJkl
tDFoxHnU2SMf+d0aABoUnX4YQWz96zHqs0Ag5dJoKZtSqG8n7eV9/IoeKSpCWzH1TQ02qGEN6Tk9
T6ie9kCNvCWnvg7eg3dmQDNj4WWc5au3EDlj8RRR/sJjgUOv5iru7WGL/GfyZPKLJ1dz8X1SbcUT
LGkf1mx7DkV+DiQPZMIDNpyZnx7bvl6TEad/0pPDMBj+Zk3P896Lw9EkocRYW2OMa+PxKDnSvQ3B
xRCTghKJqvdBnvYV9JUMQLWcNNB6Jn8r0iq0jhqCYdgiNVuQbt/tgTDMSP5+UVBIUKQpmfj19h0f
/nH2cqJP4KzsI+S8RFFYAmyYcjHa7G4seeXRb06TbyznpDkan5rVWg+xB9FAtv960hUG2EZ9R0Kh
y1bgCk+wQEv8F4/4BUtxGV3DXon5E+bjCyhQycZHTtns+ds4WYoZz4i39sNiqDsSvRdDfU76mKBz
QY4BLRUGmjEMNPMHFF5ZsUgwlvLZhGhK+XItenuDQajeO1OAFfSAZNJ2W80COr8LM+b3LX/Y0doL
hpEC4NCE7nTB9/rXm15t+xPMSL4VtGSVg+EttI8OaQ7l7Ol2A4qgd4BbLeRSdhgNIX1zwfgdLVI5
3Zr32WwraBrFPddwu4qBXHfi7dh8Y8htB6zkqRbVG0v5e5S45ZFFfObcoMKWh27YkmSMknXG/b0r
W7QuIlPVL2FEyKXdHK19cCYkQWNlQbJwzeUqliGYKIEVwkZVhHe5qLZuWS+5a6H/R98Qd6hJKI+C
dDj8jY+YCtCLOO8AXyuim06M6bg5m76nSc1PUnlqaWTBsfAZyPn9MD6KLuKELOo5PMtWzRI0m7CP
rSrYfoGO4tlyCuAEoeOkGUGwWS+zI35E7bMhhxSmM3C6RpFKXdO1RDttSAhcML3az8uJlGTebo+C
kNskiiLLv6yBmGW0NWRS+qj/faQ9amj76g14OI6X5HzZxtv3FJMsZTzuFVSSlHU6ZtKjtcVnfPa7
fykSS0Vvyf6udfDr8bEBxRcL09KpXa/IqDH5zsxl5kGIsh8o95/FL/oST8vWg3wcNQ2UPA9BYnhB
sOa/yM3EPgxedcumaDE0BQF7Oq43TCRinMRGwJMM1ySdacV33Lepe4xHWoSmRXZQGr2EBXI7ZORd
VqFs6yCIeK0R0otF1jNMSUchdeKB9Tbg4BqFfdjpH4acwFGftM7n41A+O43veHCIw8+bDVhFzQ32
BS0VNlEY7tPtHtNMxEto4syHvGN+ohZPc3WuvBmau1DZN9XOuiy1RE79DdVpm9L1pNMWQKUlsIKg
ycUdjo+KjReQ8dmBfgMwZMM9HkXb3f7DXfycnOnPcjLV9A9jLzLejGU9JV1j6o+I/LggreTzrw92
3/lbei5Khw3Zkda2kGlEuE9EQxkRMRHIdRoLLdmwvRRuRz/tNL3J+CBTWxjDOko45x/UFH+hYjtT
Td1ke4oFibSsJ+IPmaTPQaH6EEadwwMdSl2Eor2qhTAn6tZNaIUStnYZ5qA8GMRu09aqmRpbtSAH
ifcpZGWW8HKEp2wg/x4Np+3HEE/DdlehGaaf2MrZz0ooOwj6L+gzvlR//GhTnIx5NgA7MrIT9bIm
cT2MVPlWMe1R16buuf3PE2dCcZU9xSPijUr9p5oZOxaRdjCluqOx/hmoMMpCopVBmogmV4Gm3cBx
t7O4v3PLmDYYWebA9sCAfIexwgqTI9uPlZ78qWMppJG6dCS8vVP/+GUbtLiq/wqOgnoAkRVDDKKE
OJxCRdAmGePZzoH5H3bjnhffQwD+oSwrMavdSAlA0nGmt70DqjqxDs+MfvTIxzQhsreUoW1578+2
bQFXU91Xl8hdgAGkE8O4Wb9gEWA2Nf7Dx78iiJXyT0kKPyMg4Ngk90wtbkmGdClN09SvjR0sAmvY
tniQQvAXzu3TDtwvtP4ngWOIfmtB8L74sC1lwe1uHTTQmSKCnTrkIMFZrdONfg0k5nHVkFp/JR83
7i4G7jK6/01HEILpoLFGxZClUtCbSaH/IeyTao2KppXNEd3xvbmd9hCUN3/jyyq349nNPj5ywy9P
w0EtHO10d5ADjbwWk6t+HgZ0eIH/w0Qsv7dvOAXG3VbwXNm/3poM5KCtU4YE9pnipDZ2TDKk9Wyi
oZn+e5XoYV1We5SKHZEHGi2JL+YOKSwBB+2X+YoG6XrW0NGTTFKsQ88zi6dmOFt9Ga9AAiGb7EtX
w5dVSHJR84J/iz1Axz2J7uNiComYBciAeiP6e0+Tepyb+AqJT+yi1gC4fYmofQ4qbp8WnzdWWeid
V9SaTgmedB38fDX0TwkiJG/arKjhPQdiqk1ZMHEkyQbidY/Lcww6zbk/x2Nqz1GOJV50RMzgPDE9
4Zmlyh1Gv28QIHu8BeZ4onqsbhlSvAo2H/jcJe0Splqe9RSlgOXw0llY/6hg+iGMsBEMOKW0vPdO
LU96rLX554i2aWV/fsmzsaNkAoCktr1xOpoBMrh2307s6xsxK1SeBX8X8diQfp50817EODBUfhLh
kUz8sKgbg24VxrW7/6YSz6Kt4dbJBwT7op+Nr7dmJ2kqCalpDt+v0K0WV641YEg9Q+M4lDGbN7P1
8If8wNHtUAAZc9AJDLWj5jzx4KpgMw6yK0lTWE3ZeGxfX2qAtRQR1B8aNHSz9f8Rv61ylbCTAi2o
YIfETUQYyeerWjGJqwJZhfAPoMBnNvchm6pYjMToFrWfis1nOlwsy0JQGNw9TMHG5jgGArEB5MYg
mq2oM1aIXtscJVTLfqBwXWkhUEcecoscdXwXtCyaYAtWEiViOj0SpkoD6qQaNUzIDCYt4Y0wVPtF
xSDrDS3sRzW4JKovsW2nZ9NzAyc0Nl8KRp5JduILfsIHs/AMaRGRDTWK0rTiVowwgwpMcE1aJL7r
IkO/7IpZoMfIYZ8lvHxmvD1svwcx3Zt0p7toSkO9WiX0TmMI6qm15lt9DgtooxyrCDZsix4jM0Z4
M3Q79JYP0Cj4pe/q41lQUG9CyRXrMpmVt/7xUEyCSJdMHiNp15EWxt2o+LOmP2VnGbJd6WMOuW9G
hQ+TiUpwRQzeJCNao87Q617jmuXkNbC8KoVmgBPCBkokoYsjb5W27UY3tFRdXxoAdY6hGh1ZJZTu
RecUcscGQ7ZHW35milWQ817UHM/f7PLN7X6tvtXJjxmTqwQZNeZDRcyCkMsl9ixg51TRuGkwpqfW
hIYeerWUFoa2d2VDjZnSLjapoMG2PD22S3WWAk+AJO7IIAt1kiB5aP3drDtUn4KzEaZKz4FjMOE2
pChbfzTuJODtLipjC6o9m4kX6f7eNhovlBypMfWIVc/0CGFTqu8HlrM80F7XV5+0Uw++c3+n9nq1
Rz+Hb+JkLT8U9swry7JzRi+yLiHfjcJZrB1/TQapb7zNj3OAj5PbU6SgdvxqwGPjueg6dHbIU6hm
p1hZZA0BpsQe0XAcGUpeT6nY/a8fCUnHKm3qd/J1HePwPcAvibmeAi5sFQQpLAt679XMC5xk6Qn6
XsyR5b+XhLA9EhNDePJyQuYB4qgMyo3yg74F3KOuYHrr8Akbhkk0tyRMUj3nXPK7re1t41prn+AP
ZkCmtIl0Rw9qXD01ICCarZtC/RtOCHFDCQKF7XEMENGb0aOrU4Qy8VtrHyhF/n20Yuar7Sjs7vCo
f/6rNolS0pkcPs4JRINQYuc88DcLr656s9HdHp35LofMt9X+6GuihuZ0eAEOcG3m4eiP/U+5gZ/D
zcphcCywloyAV3VkRQwkiYrLctv+UqMii3Qz0Yt6mI9T+9dyNDbvTVvyx7ARlHJJnG09clgG+toM
nc5pKsDvP90lpGWuWSVl6Vv/oBaIaZFT44Z/LwRiMqs29lyXHWunRHo3klC38pb2HfjpmkofTHbY
xcBUW0FppEybX+KlCgwlrr9Z6G60+VuTtej/co83xtI6ebLBj4wpQki2GvC7e92d7zac+tAXyw8E
Bl41EC8iCSH64giYkJkapE0G7kuSnjpGPz9tgfNA4lo0LyECX65znBNZs7iMDw+tbpJFDhxR5cFI
8fkKJ15Y33rBdrky6pvnL6yJYDSNd0isbXq3X7R+nhkc8MJqlqDbYZ+K8RSQ2UImn1QJPt/nQujD
S8IEo0v/fCNKpXwb6r+qF8OENF5Hb53ZznsTD8cydrRrDUZa9BtXh+FPowCvgSQ8r5L8nzEZPxFB
f0FYrAmkQlsMlQ3BEz3sYOgGjnHetcpD8oQjUWyrwXOMkSP7M2Ix8f2OsbyJH1oHpnwFJj1EpqoY
RnDOTMEiYyFOr3P94ScpFzCRCHmJAQgAV8ElQITJko8jI3mG+Ph2mdr/D/53cIGfm2TkLlblIjkq
Br5uFc1EgBq7aeAqc7bepbfRhpqBeDj/Nkg/QkGpxXmxbx/Ba/UN6hmLGwcQHQQN+3oYC/0GehQH
JSLiHaOx7PX6/OcFbXaCUwRN98hA7bsgRIXb1PNXqgGyxWxT7qV46399jS8v17A7NRYopipcv291
ufBG11BtoOEbULtJ94a/lWgaZjaQM+seDmEgXepi8KpNb27YVqWBa6iuDQSxYAWO5drLpGAjWUQq
Nm8MO60ZTIugp7/A3K95djV7dztPLIevXx0XmCRKd1ztW8xYpECA3Rfl/qGGAIsCdsl6xQ6N/3KS
ROXWlq6a4y/Y+rrxpW13g9mxCvEZVUE/Y7nzXfl0b1lrkaiJo89OFJknG8+3Ar7aYQavTgHCpH6s
sxOFY849ZnZYzHAQcvaNjNFIlj9nBFyXX+rbSXQ6pMrtIYyc4kh4OvVFPFZrWGgAdVaiKLCDn0nn
3hr/ZkDSG2qlLBFMR/gIn+FO9ox04vHq2sgajE+mugdprrh/QcpVLsLLpyoBTSLKtcYKp6QsBhVT
VSukheWfXcavdI36Ogrdgaid/5hCVVf5N87lpRiJ8VwmCeFnMILY9TL58dPelLJLMxT0A5IJkff0
EdbKCkk2H00fS1LAK3ovVPnQLUtLVyOcDgOOlR9j7/CGOBlPbs7iwR9i3cRzMrENZ3SdUVqKBRhN
VW5p4H8iGareNcqTDk0W9o+s3N+y75x5P+IUYOq61FEKwKak4zjoB2Cw9kcDUJgW2qQWMIb06sl/
wkHapbHmgpo9oVoSOE/dwDs2PvSe3GWyS9dJtBZWs3iLVVu9yNWlRDCYkB+LH9Wg1KPpDqko2KYa
nsrpnjZbkEOk8lmQUotwQm3u38I4vihwOm6Yw7CudLompn3zOdfZdXJY/s6X7L9AVzIN3R/lnq01
JwM38AaJnq7GXXFcQvsPGPJdOJa+6L0UjS031HB9jp7FWMdXamSzB46u7gEUBsk1x4IRURnwu1Pw
fG1rmu1PavEaEAZIoRKfVRAnCFKlnMSKeGwo+18wHyebGKfnsjdAqZ1/I363vKuK67Q2YDcZxFS1
gySgkkO+xLu4x4f3OZKZIMXo72GeIUVSMxay7bd3iUqoxKyRdAvGLXp0OpG7QA2BDi9Y6TqmsrYV
YR/J0pWa1RoW4acPNEy0rkOfAjWiB06gdZvk9d7V1ByStKyLpzJgY3+yTvM9HbgmyhhVSP4RTqMH
Xd5jUhywd8kT6n5IOLF+WBfbHaTTbyWqF/gOjGFlCMl8i5u3e727F3OsFM0KGt9xc8jRmJ1mbGSQ
cT4i84N2l1r1NdsI4uYxdEOI8NhNFrFtz9qbAdksYX1j6wcyVx2MfZQzDPzxe06d2fo4Kn3jtuyn
kmOP1HErcaQl70hihwEjGAiJ9SNrBvmVN4OEBJdHA3zng2OP2j0IyEBtHuqqOqQeizvxAWsEDvfL
HwXm7mV+MaT27H7lI55M+7AowLYq/nkC7hqh1u5HR6g7FAS/h5sxpaF/hnGLDSfL8p7KAYGF1kTl
XbbTc9K+w52c/ReutJGdDdq5KKSU69lwPqENUqF3yVVMXshUH9WEeX0DUn+bayRTQCbdJx2A6cEI
ilBQCO/d3+Atz/aT0Q2zyOVt93j4ybHy1xEi1AVug6dGbGORWvE4WQBaqHe6dZJL017TNWgO03im
2eYz2T5nnU7JtEqyBXQXyfvnGwP/exFVbnBuEyrz2MaKnr9X92XmQpi4QZ2TZ9Bay7jRHGuMA5Ks
Lv5oDUkYM1rkXYIpb/+nLB36f2L69FSU5/w0sMNd5/04WgJwBgG+BbA+YlpwaRQ71q1k2et0sqNH
GGUFR1zYqB7AhoIgIjj2OtLk2i2unFK71O55D3rLVXojhEjmRuiyrtgG3DLAyKUcBFT7XupAnr9z
BVdr0T91v+akHZOQEf64/Z054R+tDIHKRQCgTEtgtCoCj9AADjHrStPKpBMPRUWBTeXNMfcMvkgt
gAKaSyEBCV1elGyKL+X15y4d6mNQo1vUayg+qDdQ2cP0QImHdyH83N+eCkypGg7OEzRfIWVhJEYb
n6qe4Ly7EEfzSFG8BSrnZ5izzh6bwRuVlGOMNeBogntDx6EsbC1v9Jx50Xpq/HxIizouR95PHtt8
2xMm169GGMn42VEM+4n0nrVUuDkncknUuQimekP8QmJ/UPe34WDXGk3m99SNYJq5TdKq03jJ/dEE
VcXs6K/PxE1kP2EHweYQ9zuKhVdtxgTkYsFV0KLh+XwRYaWbhHND5BfJ9yeBZaH7d0bW2htzNZtG
EOXskt3ftHAkpIogUFNlMzgWXzco6ZfRa9SQ8lHdLrFeOTybw6zq0hUiSHh/YCO9JzEHQXiQlbKD
9SIfcRiiz29Ql7GUzf8cZ5PAkyjmJiK++pFRqVrm98olhZPgaUjnGX0oZmHT5ErgP5LPRCLq0rGW
U+VsuRj5WOog1GkJjURTvzU3pLJ8pZ/XqXCfY3aHYO0Im8N1lQWbjeMs6ll3mhis4eJlxOPTsB+g
9UNZPlqcquQM5CUDy9U5caHX+WrLErTSoCnQowbQlgMMAnqH20SjVd1zBFq/JLmtFgVDYHQDN1dw
xCu3HoYociPBpZ5oPpWwNvr7gGNkO9qvHlmxpgEseOTZcE3ojkPcGPATqamQjrGx7oI9tzIopGxB
MGTBVkhEIcnOW5/NQl0vGCV00SVvahnIew2ujWCyf4baXih3WfXJsKQ1XtOnWNPDpCsZya9Da4pI
VMS1ZunUHbyHNVwYXOc3fu6HbaxR14MsCcytW2HbT2PZx5eEL5Cmj0DcnnkquIop6gumQMGOeC+p
dt9hJYnOQ38sw9Q+6X2NNmfCzQ9/Wn5Cn/6h6l4kYtaOk/bSEfF9rz7zxmPJTy6kmksj6CEQJc0C
tulwf8n8da+FppWqo9EWgDcHylqZlmdAyQYY+tAvLTEELWWx6eLC3aGJquWl+hFAaXjZTrmPrTt4
Xy6kJFcoOZFct61OueafWun/ZBiXw/JtDBb0jWBVWtEiJaO5iPZi9nSLmhiAsNEnjiXnHO6UGN7c
9L2lnI2l2oA2ojDlB25eNaBl1vmQQM5VU4N9GWY6npDvC8epHmOVfyDmcZTdfQkBhGMLlUVeybUI
v0Zvc766QHtooui0DemE6aVePlouN8AS3KEugb1yaHuQ/WTboU9dRsA3TBslNGu5OXIzz0lil/N0
I7bqZ2Vcw3Mq1dHvIH2QpJIQoZN7oQMPdUkdTS+6MioS6Aqp5/J3zxBnmcnGMg6CbgRyv08VH9NQ
Bnkjfe1J27RQBCOScc4nY7U1zfLKyA+x+ZMdq8QifBpvvc+JbSpw28iCG/wAjFgPjMDLUTYfYyXD
wzZCnlbiBQcBBTL1BUT8Z2BPn+/nUV90l3BSSGX6UBJZ/LXti57oe14aK4l4kjWDxeL69CaZOZeb
23+5kbCrtP1Z3RSXRuPBOxt778C5BuVvv69FDkeIFjf4pGAvfJVjSO6mcJ+sDpOHKOvBcqRiyT2F
J2w60JpCGLhunHE8A4tP3Hg8uaXKYYHL7uveshBHJnXdr1S+SDaWRB7q6CrotzwhpitPOnyv4m+t
DwkQxHpLyK5trPqpjlSUaXNHGxOljrgzlWX6VDRfzJjoTgyqPKXzLfNeaEECVHCzeRnGQmnRIQXK
+eNmJPuQiflBiGEJx6U7hwn3bwHnaJfTq13FXXwCLv0G6GC6GHnjeaFmuuS72DhF0iue+oNhKbGh
aq20ZgqVeV7WAjpSBWLH8R3ywsUkaPMFm69FAY7lkayhEaNPpblwFGcx45/Huib+sEspJJxpeAdS
SQgWTVTb4C4k+zGmuboUikLuCEQwaal5VW70ntHoihztSw9Fhd0z0X8iE7+hHTlHFzpQMQ1VT791
wyQb6E6mV6E5Zze9ldM+9dUArPwcW8b5S2xeywNXMQJ8ofEQgcevoPRLw4SisSeUrFIoliUJCSZ4
Ja3RM9AFy6J1+vuK8q8q18JMCjlb1Bs6XV8Mpo2+njyyDUC5ML8mCKkjlPmEfqyikYOLR2X0zPaF
atEnqLVXHNCXZ2aG7QEkHCiezIifgC/PhxL8RYTyWWaEWZYPrOq33qUik+GH1BdzvqUGaJKG3NHk
2HFw4pnjspeO321FxYMTcdtyEXjBAcdYiQi/vIMDLkoc5cI993oXl0PKR35h5FUJYCAZiU5wdyVf
XcERY5KW2wxed3ab4EiXq8wrZNwDSUNYwQhxI2jP9Yip8peKxUs5Mw51gwOLgudcGC3URz8vxjes
ngilMDgs5cBmT0K2leq80B7333jqcfLKpNFsxikn7LP/Jxv9NDpXX+LXA/3F7ocJITSB5aqb9rSm
6ebVEtBf2KtItEp1fml2Qv71D5VcngLSiVRTyGGWF4piSoYGSeBxaCis+VSCKqreRew0HF9hWnkM
ypsoudOoxApzwS5v+Fkfv9wLZ5+P1maxrVRF1jZ+L1Y9+T8pW9XBmmI/eppnWPnmoiAN0sL4/unO
EXpU8cvh96fJBD+gBQWozwmhfR7uP0oUiVX0nAzC3mmG4BjG/0VfxJ/ujnb0yRwS8M8xFlHS1Lz5
WfWALLR803ip0t9mDCvL+PZMpo27hFZk4aLeXi7xfZFcQqAHI8F9FVdqf/EnEtV5AQVqRS9ilOK4
Ir0jZ4vtdMHxhaiWSE2mC3eoyHIGLcundDodHYbxNDKiqCaVSGSwzbh97YQJjTo8ZAVWKARKSRPA
oZ0kT/L23izJcfgdJSEwvgg7yeYo5GtN/BMvL/0KkI2Y0YTNiQxGu4aoLD3N9IV7b3USS1CeuAOb
EBn5CghrY6ba8keYZNnR7UlQA0nyZdMMNgLrONzfVyLCeu/c7ZvxQimmwZ6Jf7LVRsTTcpyiWyq0
ownfYWiDJzTtVdVPH5XFt9CLfQGRwCuISbZqzIOJwBGOy56CICTXj2GGuRUzHvy/JinERqvPbvwX
ODLKO9bzlMghiWdJhM9HXo1Ps02Xm2yGlPnwhqAkvK4fmW6lebhiZjcDbIY/0mOubT4vli9yEFAH
P74YG8AujcAQ4ZLIKAFucjoxXfcZlysgtw0qVjGV1cky2Ht3DjU+AEMMmYMhHr++nXWEbbJDfoXJ
0EMdAGgvSjlDaUMjsMKezu2K75tP8n7JHV5caXANnsCVGXobCVB+F5d+ekH71Nw4gzdAgQKWjLIk
VHVjbI0kqJbSBp4DP8f88hEJ7dLkuwe1LaxCN8IENFdJ8i4iYNcqh/tflJb3P2bIsAWJGv1MHtGk
n+7dRtDdCJyBK41J8hrNtD9D+fS7ZGnFLL6KBQMlSh0qtq5WSWxvb0b5QMOEuS3d39OKaKI3wpfV
jnZdobjl4eWviud6W20AMK0EkSwLQqcGZ1hx1i/NCifCxPo92vxF3TVQ3zM4Y5I2CHJ6cXK2fJCH
ecu3KfirAJT209J7EG/XkqX0c0Em4YHwIvjvhxgVkMAPRHVsMD5sqU0d9vJStczxmBl5X396zgoy
I+jzhknm6D6d/+eVQT0x+l+HH0+x5T4c9lEJF/gk33bEQtt6Wjs6NHZaNmxpJuIBP2JkFMC26liH
mczY6rrGkLWjKeHEphqxNfGxPic3pQdxUCshU79v7/2JrZw3PeNOysno9WnxPHZ5T1vO28cTq2gB
/nsGL9NrW3Bk+eWlgryBv9R+p1/xeVrJDSHoB8KG3aTS2498h3Ay6FXxULqCJ1TFVS+EOw9dhwqK
BXkILmxZCgiOJ6gQC/gxhlMduqp5Xkc1sgwKyRP1dMzenTo8vl3KY0jIbLuwdE0ohIWtTpQi/hPY
acRGep8JK4qidU0mheqFsdBuYS5nx7Oq/mKRCEMt6dX61vBF87SMo2hvL7DEF9EsTCMg/tz+xy7N
Yw1G60J9zm/9x4jtyQFzkrCsM+hs+vZHLtkHTgvr6yH7hS5lLRXMcm0DqjCLNUSpwz/onArTBibB
MVL06nHp+RxIf6kH2MPQPSu75lPet6UqYDCmE7BKs/+y/mek0Ejjf+VYYGlVOI4d/6oJmAGPmKcX
jkqYSMp2minOqBHVbIewFj2LZLkgRXsThiqPTB0tVd0THnZ0uksjwi9Rz46Ry5yqKtniDYcKsaft
wkg2iq2yPCeDLAwzFeQk/EiQj6U8Zp+xYw872+z9t+E1xRIfHOSo5AD7hGw6sAEbMfHwomlO2Ino
T4wnXCK+nYnQBqwCleXuYUI3o7lZ2A50wuKG1va40jE7QwgQEUNoXFNBKrOg4B7Ah3y+xkAfI0Ln
Uismc5TOKVF7zK5tjVMiTpIz77eZ14ShLOhf/r8DkFYUybSMb/s/Ey2Y73A7dSHix1P3oyA4wdcq
hmFCRuQxhbif6YSxNUUKnoyqYMG4L1bqt/ZfxuDcQbEqg0US8CDMdjFQ7X205y16PNQSHKIwpYM0
153nR+3xMo13xO9MWIhrKR1ElD5wCrwV5ZwM9Z+B+6lZ5AIikGm3RBR0FgxDUEhvOgJP9ui3hLnD
O51MYsjiJ5oFuFTIjWri64QFeJGheo3Uvrb0YT39H/W9KkFGX4lD8l0ABDt/2IH+heqw+ZN/Qdfg
Nln59e+1ks4nFyS4GWyJLn9TLJbEEbwftr7AbPRhz9spRtJmAYk9fN8M09GL3d1nG/dl5kBvaC2Z
drjwl4xXF2b+lryqhkUnLV2B1hImM4kkQOTW3MOv/MJoLGvEVsHUVWE3oi/9x40cERmT7vdOY7dO
wvqV70ScvU8+WVRl8wBERBJ6bugNby4iyhv556vzA5VJ3kfgKQOsvGgEI+74c5EdivCdOZZ/2A2g
h6AqvZHKjwFqi1dsgjfajtLI4GKp2RFa5GKgO5fxIl2/Qq/HF6vo5wHjLIKDJNvo4HhtBwyYhYCr
mCyCeToRsgtmT3u4DUabdBVQHS7tf51+EBxOSGgfZzbOe323p+zZrwt2+JmfdJR1AmJoXoj0H6wc
0wcJDMRc4kEoRz7xL9fLVwSQs8q2cG+/Ju13FHGVLJMP0+3EZDhcAxKFRFa6EODqbYfWcY2ksy6p
1du4/MuRf4SRaU6+tSw9y8i9xZaaK2Ao3GFlTdPn3mYSpkqUM2huTheuCie4QMZBqFXPxOPiwlHc
YVMW4I4lJDgTdv9ZKNB6QNbcM+GCrQQD+fQGRz78mxN7a4damS5Q1VvLtt+tBzsZP4/kYioRg5TX
olLcQnXpr3Xh3LYYmOH5NPRxUCJq4KeK5EjUmGxiLGUjDN6460WqAgreObxCiT2Uxm+gTTVxzYVR
RTUyXGa5INKsOMslZln/wbAaUxBsPHFsLzKaTC5LWUzIwH5B/wnCuoWm3BdDe1JEzuEboH8U0FC/
2JcWx4WndMhRCmaKZN0UiKP08/YGY95QbxENvdxx4n2xE5AxPNsHXR6MJtSF1g6YcCz5PfWj0stS
id3S88gONeJBzTfnZoWIPHqE4VQPlOYWBnvxDrA8puTsjhUoCpeprkI/TWe4hG2aL6q4F9K5DYYQ
yDEIzBUahlV0ZHaHrWiYSWHwcmlh21ePuelohnD9LnUuelIFPYbgjdtH/RWAEd/JbfwCkajm3qba
HU9XTJMVe/6jkW2hnMOIDFK7spOS/1SVJ91De4jk1C2UB2K/oPPoT5nMKyLzIeOEa/Gn/a7qx1sm
C2rbMH2w55xa+15k7JMhU+qMxPz6P0h56OSEqZeVvLrdA2fClZRO8WgTHRTtsnA1fI5dKoI+yj8/
auGPe2Pm6SZ9HKIU5X2HeWiJJ544/WcGfJQ9kmc29BrJaCtTEO0EQKwFT52ittEzUNSqoj65s4/z
/vYCzDKvWqkbiahJTSBewS+4mxgZGVE77Cr3PRmhp9b3jqBPACFWLA8TjbwFC2nWWVK7DWxt+lIn
87Qg4njY/ZvK0xH6Yn7ZPS8vTOSmyxpZwgdmuOV8+oODkbz/Y4KOyjzQbHWv05BP0NL64O/hmlaf
RGliLH1x2am6nF2QyYHOFEdtT3NTcxBl9kDLAkyibNxJxRHNsDdtLbrqVBdS8Oj1zFk68vYnugAd
4dR8Lx8Ie+Oj5b52K90ktdHNpqRVJOQa+HoV2+iSH3GJBujMAlpjpvjtLyoJ17FVOf7WvTcBB27W
VADYaX8u/5cURqGbXVIGDcpP+8plok5Hv/Zo0kkZaBbgFVOI5S6ngmHDfoCR5/lFaZwz7kCvx8wK
X32DAf9oCN6oi9O/2bvvjWy0e6nB6i4zUIraiokzJoNqxQcjt6+ug9ikGNQ8Y353EkDDOV8F3Qc+
lgFp6oy0DVIfNtMjQRY66yAM2yG10bsDLkP0vXkCdda2ZO9ka7mhOK1yhb5brXSnVdf2ZpPYILHL
VJ9tqcUNHZzRDe+0kg5DplKlGYd3r0xaTWNgIyKzIyXOORCAdDFYB6mcu7pYPtIBTUyaLUrAp4dP
uPOxTknKa8phJjcZYl5f2anfJAux8VVyhh/uSKm6AyqFd7sGlO7dczOuLzQma1h+cNVpC73MBGhr
fzVLsPnohfsIGy7gb3/xfIgSRVrgk+aUObaIC98/r6h4BsblYCjxVamZyLA3JCvgIBUDvfAT4N4m
WEimMGAEItsNdgZLJDJZCZRZDRQ7y13DEjvBFYpUVji8hyR5cuJHbwcla77M3QN5UurRxid3anDx
J2FsEfOIgg+ZtTDoatXpC4r2zOYB+xzMeEYAVBhN51gemMj++mdxAKaM6+a/3gdVQDOdMs/bfTjv
ZM8Wyh4FigK3UHNKwW/rFY55zN9pbq5VrlCKMBFrX2t49teMsrGkeknGxNjOHgN3svinnlwkEQqZ
up3h8jpptJ1498rZp6BGZrkRfpOsoIJ/PW5chX8vLn/b5gVLAIS/9YNwCAMSPy0h1wlikcxCOqg/
DbYESOFhYgj2KPz1CXzofO0EI+pBEqKhC2yvHUEvWe73Geb0dta5/d8T/H+sVgrs7suR4FDA3Pt+
G0vq5ClSH4qLC9xTmsrbHuD5iwNR1YOeONlm6D3evDUJIE9oaBxFFXroZoqMnWTwCbmLYiNTZz4x
q+dNu3CDRegp8rziZa4GyjoXOhqPVJatUDcpmM9EE4bInduCra8OyZqRcE22bUgDMvSv9QA6e4s3
OqhCybAMJ8LX4kJxdMQdY139TNc5Egmpx+4GiHMTxO1PULUP6J1O4Z3DmuXSpNSQRz1/ZGh4efs6
9IPviZVtk5L8jhPMbS0d/DflqxQBhPfEpQV1KeIgTfjAVmyVgVEb9U71qEm4yBFint4G1dV3qRpA
zFFrvs6NERC/IMID+CTcdw2iaPfc+wvE1wY2kBxLNnFGfP9yPiY3gT8JBe2yv+rNSqCbszihWLXY
L+KvBxLwScmRX/Nj7SdRWSlFChicit5ZPNxmIUUikninBPu+1hzZGXwzDUCMN1KmNyJaPXTslMIE
fobUi1tVLbm94ZYGCU9ie20R9unQPuzMPcU1v4z/0BVQYt05iRBg1+7PQUbq6+IKHpJKewMLBVqG
zNL6MlKHFPuPTydOpfb2oWQyMgGq+j8Z7orE36eh/BBeu5uEq7FZTcp6IQrE3rkLJ2e3vwZEZsLC
xUmA7Zmn+Irx9MvkGEmLTeMN3uZcdArFjmi81TGDReDD71Pb8ku+4tDUvJ3MCSlICDTRrQSte5r7
OMqLvwa9eOv/YlKlH5YP1QHUTLHOUhV3xcHvjdtdpS1JbVVfBNrSdvt9O1AKq7zjdBAJG64+kSl0
IxmfjkXFxAYa+aWGbWwGyp5CqdezjXN1nusEnKtPYujKHGWx4Akdm19VCA/P2iHP8lXNJqqFuEha
pUsYkfMCVol7L/ehSAx3XtKoNVCtgNgDf0JT0016bq4BeY8nmyEeyKeL0zxKR/viowpagcCfw/NB
DgTuslDqZXFkFaaDxRmh5iz8Dg+rAZLyaEQpbqpdmg4JD0rgk8FdoiwqZWAF5dB4BAlnid1ay1Q0
+VLlUb4f4/4hZ0O2arRFNKOtj2tPdqUr2Jo7PkHa0wWm4Iy5RzbfEKfJ/U8o6Y5u/SheLy8DkKpu
Xdl8mp7HECO1BPOSuS9G1/c1tWL9GGXLVjtZGPSUc2bgRO7miJr1gsyJYka8Do7yByZkWMluAJnm
Ogz9vbdaPfnyNfdJNnddXU6EIlNjXapDsMv3G3+rOgDXUvVDltteChYikkpqIYPBwWmi8/gS4nOE
X/Gi5zDCPGcgZAhZ8BLfk6g98+k+juvFGhK97q5KxUwqshL4imY2BwcfiittHik9hr5dt2edZb0Q
Cb15otXZvmobRe5V0Cw2sBiC/ytZNaLWzehQzkxtm0qqWzIanDhWyOfs6k5Bl2RqzVLbyOXYjvQi
l16jmqP/8lDmAtPjkwyl3ut1F7yVIgTzaMOTJAvtFYfyzP3a24SCXVbxIF0kOmXbQNMR/hoVr232
NWjz3Zxzucs4x2gspzfPIg11WHfO3lD0m4oxIv27sme5pR6+rjm2TNbPaL7RMv9TgyB10LY2Wbl+
gozxB4BXIXtEHPkq5qeLEah8T0C7uMF5ybcQkhIJ4gGAY/CNbWcCJVnP3LV8Dt2cS3srMpLWvTA8
2CA1vG4CE2FHGHW7lkkoSmQeqetw1QwwVfwjzbbT6elVxBRChIW2hh6zZxYGFl7Ud6oC5CUSqkYh
q7FT58HWTEYhruMHPzA3cGdpiLdVBKVc6flb2ChoOQspg7PS2t2llRq7PeUU4QkT3CHF6asJEi6v
NVkqK05s7bz9N95NG4bz9HP10kzFBpx7UVT/xeRq7/Bio2inJ0/tfANgMLVPonZ2RCUW2KqbjlLO
LsJ3sJz93HI/p6b+4LdSlyrDThrFK+3N5mni5QFKeXf/a1KNHPlY66puR453Y9SZpkTPk2SFNgUq
NvMav2C/1+Gva1UQ1moyUmjBAgavTTUTC5tcTEGim4/B/hHOo0D320+47M3jMxc63mZrlTWYdI3J
D0lwzQNxLK+7xfgDPkHSM5393oGkfta7aEnLNmfIaChSuz5qfeojF/AclM06wpf3AzmhKbRNp3pe
cyUG9Bdodfe2GKCCKQ51+hZHIiwXmRsCzXPa23tz4OSahgKtcQrQKjXUOwHkLuSH4wtYkHwAyMqj
aUUBnDiwZYeBSAmVKfAmjDeMcrgTq72bUaw1veoky4aTqdfS/UHy0AZ6P5l5hPU9c6Fm6HBUhORw
oLfIDglZhhZMT0QAE5o9khG7ITqjII2ilzdFYUMMlyXbZY43r6Kx76r6O49CtrPERHK0IGI1KMR5
OAdb/93ed/346k2nmW5mwidKuN04Ska5z2Gq6Nb3dpJxM74PfjObLTeXp7oogIxwD8iTOhQiffQo
Dwrure+ZDTLeX061+vGmZ7dPoUCpUdwq4Ll8cXvYTGZdnUbvDQnERbw//ETSVjmAso2n6m4DCOOU
2nbcI64k9BMg7Z62ps1kEQXkrgmAg9AZbQez+Kb6NaoDiIkQvGMNh+UDR62wluLRrH3SRogzvVNV
N161ZxPiCc1y1R48+wdPIRNai1vXAQkgMdBKfwEI4k3kY7nXihYZtJTK7N0P0nQnIQ+seRsUdDtD
kH2EAInIRl6HtQ6Q40iFCY0LDcf94sSD25dPDGcJlYajkPhQN8uWnbKa1VDwrV23YJEhBicganAq
Nibm9FcPla9FJGumjv6wYbrdLBQIfcTE79vpTCXw7TvvbjQjnutNplUMfY9mV4pDQEUnhDcoXuTJ
uYHZXeZj8XJy/FOZtDh6HBoc7tsFpVJwVK6QJ/9hEdF2thT/VHpNgF9F7I8JXonXe3cWPdyM/JPl
d0VMHuA0dQhlQEM1lu0FWT9aP550xyRiRVDXQUfBMWGH/RNmdU8pnAsp+2OIO6Ewz4PaXLUYcoKQ
C2xGgNj3oLRKsmQSlwhhpGs0CCIlffXdSexObM4uGICsIUeRbPaaYVxZjNjX9Y5uUOXr8fBFRQ3o
mTDxgqGYMWO/0JXpvYqez3wGTpwYGbd2cQB2zpkiTToakb/lc9yYovtHXEkLEQldWcmFI+0XkHmD
ZhXOIhEMa1ye3BywznW9Z23HDUen9wJuK+QKCh0+Q/tZFW9zBqw1ttdQCpvAzVLkcKg/5RU9K7Iz
ngPbaObTymtgUgoQSk4IifJYF5q4DFsixJrCP3VbJF5pFgdlZFv/SoXQ+dFAxwdkaRpp45Bddjmz
DctjqMbvqGWW3thEi/GrOnw4Ly6AWR6hMq/lAnKaAAK+jmjG9Xf4UCXCHFyHOCnyhwNANj5OTDoI
HMt8sSTcorWdfAE1rdIwIEy5kDY43lc6T5s/jMKzIZp0mxrF3ijLbcn2+eYLvo1ioIUTgzXcS+em
wrJ6eEk3LfROzTp9zZRxK59Tyn5t2AjJD4/myKXr53819ay05HNuZ6/boe3riItypdxJcebk3k71
KuUpbDkdMbK272x5SaDsZZ2frjW44rMvMqqWg5diQXcF6ORKVDI5b/Ey5dAIO0qh2oD6VAt258Dj
pplvoQWJyyBUHlOH9Vg9G+4Vy+OBvwOrdDORnQWb9qg6JPilQ7AW07A/Hl8ZoakgDw51x7PN/b1B
6RkZp9i8fXVY/PEr2RzkdvBNRU6ql/qOwEMvzKYEYPMk1s9TFEQTK2L3ANFBjn/UgOK9JZMgIRHH
6Z/fiJ3yck0yqmZVzny6kJ6nEN7KhSZ3xFMSYWWwmdKpePUK6nmGY0tS/7QkmzzGnSJJLg/tgvoq
JGQpg17sADcqgMjm1CKg0JL0GRJXiYUVwO4Oum3+ZdaB0lu04z+kgwHzzlz64V8ocCuBcmRAMbIQ
2Q7ToVuD2Qxw3ozSPX4zJqe4hy2W+Psth4VmNj48d9YKanxXF9kmy308ELuzTkbUi/OEJmLTyZlF
6o1vyBf+TLt4yqxU7HAjRAC2xgPvbCpvI7QQXSP1fnGmCuvRD1+yAeuKtLbs0JXl7gsNJSjTnUmo
JSxe8FLvBhphIV3LmzwGa0Zo9x9E/BlUYXKt8DIEzOkfyjO2BctHxOUPt/3HUDrmhCZrgjkoP7f7
+usM92gwoafUz16qnOqG2YgzULMI2Bz8Af81u/FVrCxJlsLymN4+WyaymWfwMmHpJP6AFrsPLho7
22Wk18YYDH7tm/fz4DZMN62sFFmEO3Ml6yIrkLWlkFmcuqNKvTJ4j+FYJRvrdkhKIfejpxUchp3i
TiQGQC8iXB4hHdiraKe198RMnfUrGZ/yIeKNPVpNBjsPwQCuILU1DYVEJ59t2NUqxTiIZrste04O
5NeRv8mhMBTRBbajqYSt0MARYtY7155Gxn/J01kqVkd6gM+PWUpS43IGVpPNNM0dh0+76Y6TEj8l
llzcInP0UxjfM/nc97BZ66Cfv1RNUX3bJNo92jb82YlzvF1rTvgeImBpybJfV/cj8yA/AYwOGy0u
WgJJmMHT0lzvWuenXjwbxH/BEiVT5UjZOJTL1y4/Cmh5PXN6yFKurRxRAFgX24W60gUmvILv2R1N
13BpcvzcEwC3rUlXJQmtvzVQ9SwGs48vbq24Z37zoRibeeVqwyAQ3LcTYUXIGVaWC+2qqzoZ+zR3
MREjNZHvDLeLNM502cSIiV3P3Orv8g8ZNOub6MDNNOgbG8NfrMwqU8rw+soSq2YgINSzysaMf3cn
y0PMFZ66OeQs/g9VzEDpGmwelZHFtYTnmoQvHQyh1VJn3gisiZpU1r125GZcOmpjg6qCIqgO3ECj
Ndi2HNTZox8nCWQDLorQEXqJPrGm2pqM2RgFGL87QgEw5D0J2XoYsm/8/whPvLozJROQtTEtwAfp
RUOpVPNxpgNnTijUwZYajhbqIya/Tnu1JQTup+NTkopIAVKL7qbHqWz6trFCR7xkPQFkbxl14GNI
7tkPyDhX+T4vxae180RfuGwRRw6ansZ7fBGq2QyxtmElUSoRuQjmey6/yfI4IBTiMSBrRI42snyu
YLJhMjjIEyZVJE+EG0Nl+adTI82kARW+DeiCI5mYkxOx2dRZOPxwk1jKuGFq+eNyVDzRxBU3/Ik9
pWvTIKRm0Tpsg7qs7Y/H/02HsKd2VhC7LWhlZhxCYZpbNqKkzt0XCQAXRf2lJ/f5V7in83gy6ck1
uLthrqDbGlbdLs4XFrqnDLLhILpWnqkJNpOFeu2qgvWDXYhb+vD6gSc8aT1BEsaj2S3folJj7cJw
B5L5h921VK/fj0zOpTmZaVoT1RkcbGFvnVchIcXsSJh+N2UKRHu4NyVad+LpabX60Kp6pNTSQhA7
iTws8cqDN2t8UCIiN2i7fYxg/rvAxXtxJeyJ+yx1T3nUfhjLK5nifYPBxsXRHVPZWo88jKSYm0IA
4Disofbb21jJoL5IPFbA3HpU/6/ycYdrhGFpUeLcwLO2l2Fud2+MKrBvWRJAWL6TuCnSVRVW6vjv
Ay/RzcRW8/ckVEqSbElm+SD5PKAewgrpJuavYgBD6pM91RnxIMUI/9K7lnh/qCUy+c7mFhCzGvh/
xaEFisoursJQQEYBn0FaV+hvStymYbvfvVbq1c1xXGU0eavfb0+ava+8DGyl3YW7R2QdB5EYdlyj
Gb7V1RI3U+DQl8dSlPVM8vZbQ7GKAxcpOS+LxS7YjRsaUkRNo+tOko2sUKTfI0rL4+ym0n2wQO1g
8H/N0VIdw+lVVrwvsl3bnTZdkur2b7GY6VzsUgUPplvq8jVVBqu819lRveETkjoBQ6qaFV5V+mlk
w7IK9MK1yyvpCtn5yG160omFQFQA9nXYngxIZT5EfFFtDWhin2e4Y0X/AxcmN/cuZiKsf/p+n3tX
sIZPLwTQw6jBfEWVzHvulb2LvoZff3kKSRSeYXTq5eKsWIeSBHWnEClMoWyJDpyCNuwZ92jdspwD
xEeCZb+3k+uL2iuPPhgLbQvQwMQB7W4klaj5u8C1gl4PLZEy8JFBrlA2Zo1ds+GFsTjwy3fddpeD
fxpItr6vikPHYWt9c1CX/zaL+HF2WUhc8Wz+DDM57/dl/rI6qjEnx04k+8HI7P0QDzxBcdkcwxIb
rEXFgA2h+5FCLLhT0hYC3LbkwKfigdo4xcmMIZfNeeYg04NXTwTKSS56TlWGR39PsXSP+MXQhvHx
53XPK/YM+I3Ci0jSQAQkxxmQq2Y+rXmGUqlBCFW0JKU7AyLyKvEqOAtXJZbPlHtNyqjo45UiS6P7
fiM/JN/zBARuO+ZgEvdQ2S1sdKqzRijEcYe+DQQiQ2+cGmAnbmi4CCCGelWDt4Zq9ah4Ceyw63dx
uSivcR9h1U9KkDnHvMrP6nHTsr8L2jYhsIpZTc8ObL+SsGkvX7799CsQMBOvjYGD7jHOhB5LV5h7
oFuuUXDQirTf+xC5GfAZdz5kLKs2GS2Zj2joLcL7Agq0vr+1PQpTplZPxmwddtPKEzSrhDbxzI+U
EbolhV2cdZBbtbSBXiDe+C7eGIIRiHENWSWt9vJakkAaKqxTvoXVH60PEnEwlbqv162Ad7jQ+flW
vu5N9+HdQyEC9vT5dQ4QRsVKME2ZTQ8QglWdP/nhGI5KNcPIT1+6fDf6/8sgNw3UCBbectcN6Tio
p/z88pRM7rkU8qD35I8xdWNTibR3P3kW4tPUZDYGwJtkW7CgW0rRVLHHATK1WLLHJHVm/kfDNpnG
fHfhBRkuLpBbPiH3nHMrv0T+yPxGWxio7GktOWRuh0Bz3vv2dzXKIooj0xnxRoQ4mZAd7KeasErL
aYzh+YozuVd7ZW+MNGNT6sHiVnmbms/udVYAshOZCdtvrR1+34tNHf5b8dy39a+OsoWjsKhOZzJg
IEWCC11EkwK9Ul0nEUcFuwgtrtch59MaRH8vob1rgLNFZL5G/Mx1kqGC8P0o0i5IKB8DCO7kxinE
QvOQcfNGYxf5Ypa7RGnnnSpfub1GpxmibOnkL9Q+pnHwhWBOy0kzzXxFpnJRNbtROjG7qPmW1+kR
KdN4eyXHkbFI+c8L1x/zaha2T494Vt2/XNrNcGXrpBP/3EZ8bQyQnYgpcy8hr5tsS2RSnvQJ8Zyk
9rvgjtZutxplDDyYjjGvl8AzM+NeNA+ZnOo7WxicpzTezyT0iWOZCeN6Qz9PyOHbHZblHKMQgRPf
2in1K1vhwYavJ1H4K3W6Cu9sAHEVHyAHzFXOht7HFvn/9o3wVN7+NVdiuahcnfyv9bDLG73RNiyN
be33kmxH/ImkGFrO0nz5Eg+iC2M1b38TR7h67W1Y+FiQO5bvm5GK9uvpmqlNEQkQ+yi88Hwrjxkk
lPhpA9SyH5ekC5WTwsnnm6IBaTpIraI7whVseSfKh3CNXR7wBtb5wqU4avTK/FJPYNMh1P8t0X2y
qJmk66WHIEsfWxht4HHLXY5L6zV6PzlG3RrzHYgNyMfgNvMSy7KZ+4n883fJe0OcXTv5i1w5mhxf
Lwvqrj1S5D4iD7IibX09rir0J/7DEnF8bA4u8rogZEqq5ceYzgtYDbBGS7oXNAfYAF6k2JRuLK2p
Urq8oUDNBFmN9Rl8XXDhoKEy0k1X0tCpISoESXn5zp9JR3MabM0Y3anYfY8ohjLKmilzSrhjVb54
jS342HlBo53Dk1H/bnyHzbvmBPAYT9eRE/A/Dg/WLXWG27nIJFbX7EURBHvMPrcmmoOKqVZiFqnV
ePNogEpk90CJeYgZKPYYyCS4tYxVtl/n0hwjg1zHq4zETqUi1t/8SH890+Nag7QQnsjFWLkIRkAW
P6cqB9aAKTORFqYwb/J4My1oFmAnD9yGTL8w0ERxFMkJb/HO+B8DMXcrzwBrLV2R/eTgfDfXMr37
QwaxZCyehUkzfrb77uDFLdK380PDeaWwHMO+BwWWX8CS2QGdqIk53A6WvE/+5bBbM7sFBq4U70mz
XMT2WaJGXvFGfIB51IINiQ2YO66guAAYdywwDPvEIYSX8MwdLwugGCw13FuMTnmvl+CfHRWWExhP
Hwty92pXuO32U6QXLzMPh/pXmOCEEY9Sd/A8Vx/HP0UrqTiUVHZp5veEk0eqklMoQACdHBpIpUDv
16k2qm8aF9d9hH7coGAE0TYJ9NdTx3b1M8KkEe9EH4gsWsESDol16h3LbQ+m20QekCRmyBx8nvzP
VhYW335OeKxUSSF8yHBN3q8L+Hi3mjExxCHaRXJe321LphUz2hOyvLQZlFYU9/yU24TY/D17ZkBi
XLm26ZKeLUyF7qHyZAIP+RSHg0gWR3siK9Cvo2ywtX1ZMXvRiaTJ3JhKrEsObqoTNZhwaFhzxTVE
vgt9txnMnp/jb8PbfZCroXinU/zWkdNSqLK5NqpPLECNu3MwCDM0a9FtaUVG+kOErRTF8WfTW05X
8aJULYz99WbNt+UNNaGpEgHq/g2GxAfnad2Rvsps5jv4oQDfM+8cUTXYkwGhAFC6dY85nCBBkDtc
B8wRuHYox+2W5FuRdRCQjf7QphHIjkVws9tV6JZq18zN/DA+A+IjbqWGKhxO9oQIq9951ijrXDic
Aemt/Kq+yU2kNVkixdRVFu8jo/SoOTmK/ppLz/mrTcymV1olZJe9PftsEw4cV1UalMpJkPSoRHSd
QXtpFeR+mcbBROPo6fkFIinYDIyhqPX69TJVK164C3eADWHE5VuCbyvC6waCIk/VulnPHVEM3z4+
pivq3sw/Gx4i1HCjSnFr78fAtY7SyfjuXSMrIIGeDL6v5EVQTnM9JRk9RcL3dsoc735n8akSj7LB
j5HXNyZ204gxNiYKrvkLVik28yv+mphvzrmfOko56xOuGfRkyRRJJzZUHGWDq2h0hoZSdG4DMYKI
Zo2WMxmUtXy64Xxbr+4O4Jqn1QWB0zThaSdXXIyW2bNWQGQe6V0ALCt2B7jH2+xGP9h9sZ+HxHd3
3WHLcIbUlNLYBBwDaiW62TipIq6lQyqBCBjOtaZkSCXtcY9v8HdYmXaQuH4VI7lrd1P2tiHO75Zz
zrVIStNdDrD5RBiobKjKMXocqMJCAVsmqbxIbsNP7kiFiz+rCPL/2Q/jP0l0mdkr04G+eUz+Q6PI
gNdxOG6DAyE0egbP63V1XJfreHFSrElbVYP850915HpHR/OOY+V6k5AadRFcvNf884/BsjK/GVNg
AT/L7moM3aZ77YVFT3MDCz1PtZNXP+G/Yc2Zr4vgiAI34+Jf5r9H+2WhvMvyEj1GsOmWTFEcajDu
ZhorsAF1DX0XTkcbAOUn/nib2iYr+imbJmCoyG4X0GorXHnCV+AKhwYuTDyrAe3tZIMowobJEiUM
190AmCQRQENzB5TReeM1np4hSEyxgfmgEv8tC3NJ5ib606GUAIuVU0pJJAoAoPHrS9jyJJuTPlrO
/AKTYj8JsD0oPSSJYKLZzgba0XjzW0pzKyaVyx310Tnw7DlABbFdjvtDKEia17bujM5OG5BKSk+b
Da7wihoANtvdJ+2/YDLVkVP3VAwawOWm156KRRGOkjHzEwENYScw1bXAhx1PEiNHhpYGoDrwj2B3
agFOszIU3J4ucO9URwM4gAj19adcnlIjRzN0+Zgo7su9vo5qA3R4rfnCQ8Kfh0fGJ9sGlhSzm28I
/AlZy/GZAjY2fn+CAA1nAqclJ9rDccxJMJ4l/WV2WJJkzb+CoRosHiGb1vL1k5cmGfZg0I6cSSQx
40EsoLJ2/C7Zks3OKgOgqZWuWLdZhVel0+VaU0oGQ16D4SbcpCStdmeQP99E84N5eU1Hjy4L7Xhb
9WGA/c3TPSsyOMW8rr+jFn6Q+D6Z06m9S2Z2/57KqV9LeRPXlFob0GAD6pGptA+1xTpBt5m35Iay
NMpE3dfLVbuaxZcoI2ep8eS8TX0k1L4lKUf+IgWO8cRLxT6JNRlgwmxeVKY4n4IgSPhyXZAp9b1j
Evu9RM1F6+b7uleGAoNITb57PBd0moGwRvvD0adBoXnv5gnEObLn5Hap2xfrPu30nhhjQGlbS3G6
ovEI0joWwfRrQarFX3Sk1r36IZoVP1Jgci8rMoGDK1K41+PBWQ19ZOT7OeNXyn+zGoBowr5YWG+j
AFDhI0nKppiKHTP8e4aC/gsy/C0JQFgY6+wnEIVDUDs+6VQa++GnKrNenGKOehe7/MRmbO/Sysor
KwUmmYgAYIAJiYgiIrkK+XyMeXpTjMEW8E2qvhQfumLaHrwV0/RW7rLnbyQKkiGC7wCHKbDtFPvW
WvinE1slDrJgwWSRBhboIPAxmXYhI9frdkWY5Qtlw+FoEbQZSn5e0XTJ9vsP05+d4obCln5XScpt
+a9sXSgDPpxS0KlFqzf+j+lUr8jAGcs/3A8ExFlIM8/qWYe6b0eTytw7VUeZcAf+H6JTzefLIBW8
H6LOmB/bvJ+vDujSmTa8LdOtA/1qJXJ4Urf9toFrLglYg4c6TPT7UwW8ecn2v3O+K/VbNFSrZUIr
FbQAT2Vw+ecLbdCLPymur9jPPy/sbz1IXpoVxCH+uWzq9Wtg3JBX8g4EhFg1IeHprCc5HQcncjZ/
aOd8ff1O/YJBC432PYTsEubkcwxO0PjsKMeZDbbk59eaUI+uHg0VJGW9PLd4ZWMsNGaphkO0sjq/
eVkpm8++W9MbVRZRNU6SapD13760tmQgtHBS5R4OXobLYxMCs2DhGxK5/mPw64n82r6qoYymy6OZ
bPLyfbNb0r9ECB9/Ydoab6bTtbKVGd1m+5abKkK4KLVta1EWrQ99IlDRIymdym232YWVCkWSCZNS
c5JBZ/3nLalGBs7YbL6Sp1xC2bK6LDVbWf6Wskw/Zutnbz+iog37S7HaREzo/KrGiBkrDqa9BH70
fUwg1eF/HnbAC5+IPhwBCN9k8XASRP6Jnt1g9EyBW8CO2gYbgTTDTgW8P4UDjIUBV06BIud2y6md
N+tiAyPdriB7p6iPwpdWABdoBBJWF/eCW8BSLv3UM+z2BqJ81xpms0jL4xaTEMbH1wET6dWLwYLC
9Iiidn/AybVA/3UxxKU7pkXc/NOoFBIkGVVl10AA+5aYUizqLTHhi4oQHCefzj8p5RsF01uZcE5A
RVce3BJdRs8NzJaAqsocZunAek6B29akjS7QBM7YIbnSMs6yDDiI5lJCRVk+aW73450SowuA1HEP
3aAvQds0zeYrYlIxzWSqv9P9+BwxV2tJri95REoUpZWunNIKr4iiWrX3092XIjnFWuQKsz6Gvx0b
tDMrUrO8cNQYdD/aJM+UqwK70+tEqJ+tNSFqzckQNQMIx+NnCxUrMgMIWiIY+9deqH9cgEMQCh6Z
h1wHPw5J7ZsU8P6f+kq4m/ag+sXtDzOcU6HVWlmQYgxU45E2UafHbJnnK8nY6h2lVg3QCiAMkJ2W
v/4UP6AojUR8JdU/Aat+3Y6amMVHvC1bZ+ab0iYJv9dj38lzGRjIcFdeXGwxrrTiCp8sRWszP6of
PD3vhcMuNSmsT+/Qu0D7gVC0jJYDuNMxdiZtBhpNWKz9QcOx3ZSBcqfVDVQ2GvnNj36P2WTvcNTK
+81DCOZlBQKfzjzVK3lIg3kYmGCs8ZpKb3ItkB5g5GSZhV56rCgawPSLRwJLzJNQgFLxlu9itNkN
YX7bBiEHp3e4zehZ2OQnGbRWHaZrB0VL50nGkU/66PjC2f35MnI8/iryyz2YdkSyz149qGjMOlkt
tPe2qNLRwa++dxIgS5FxQEnFSsbksmUu/G/VMTPVzQVeRl7rLFFncCh1K7s1dM993fPEmyLNMdtr
37LwIJRBX5gA8aSkC21gZkhJ48xmpikwQ9Z1xaGxOD4n1BNdetRtLJnCn1T4+xDolXKd/+RhmoJP
cxURKusfJLYWf4iogoe36apgm8Vj6xg0oUs9k+60BTBJHbhVbR8vHirYP0kyBxI11UF30jXH87Sk
cVrgwX/1K+BNcWuwcZGKDA8gpey93ZdrriXFTw/yfiNdrzV80Dj2NKzTWcHfIhtOdH5Bxbc6gGEy
jATEvcF5tW99MYRtEUgmOz8NKrNSyqvO+CuITgHnlqxZmragcqw+rFMcAeNGt2993oHo4UjzX5qV
cqoCOlx6a4ptPYdXy/xecEm19JyHJ8RZ/1Xjv5fTqYGbIi54pxqT5stL7FSKbbrKuBA3vGBEZcNa
ONPxt5ovgfHcmDMLbQ745iODozOciUwtgq5gUb/DAJH0O5k5Q0qIjnuxPzHAPVMgDYOFcsoYuVCp
Rvx1bzVkrG3ftdtJTpfboa221oYWgeK93WH3l+4WQuJmMY9ur3EpHwmbRJMdJGa0pXNZxeyqvjwB
bwW9vnEKI2yxdqvL+uor0GwTMzUelED9XjZAsH54dLCvhopFTAyFVKvcwQVqB9CBKldq0U6/JJmt
GVNQDc6WCTi/Kx3iJtvtpZnP7RlMm10fPWI6kfXaRrPhYUDRSGZUiOM2Nb6taNVJ2Ijqun/KJmt8
Hl6SrIdw+WkdW/W/1az8x0fBKvBDxLodZwomyEHIGCNfaI1aqZdxF2qFaGtq+TPec2Wc/ypMD63K
ewvsoCmh37zjBfZu4k90gS8q+HgZBiJPe7LiUEVyRxZQJP95rdbFYF9sw3IsClUJwdFWSfIxQcFF
u/+vS0k2QTw/FZia5ZHtn1HAW8v9ksilOuk6HEVjvh/CmayexGF7sMBCCTH7g86QAONSLLjD78fV
6inApx8h824XoFFrBthOZYVFHxXELjTmAPRzZIPrQE8FWeZFR1HLt7Diyn44lMx8CQ4KsElePL1P
TTb3yGXkiWVbWUEtd7klnWvyu37zCZcQPh4Nh69YXdQGi2HkLym5KIYcUC62hXnO5q64UCe1IGqQ
DxQVPhq1ZgJ9A2vYoLBahIat3FF3e11ZTEQRwFzs3XJBAfpVZ4VVeYTRH/hw7kVLV6TM7GmqVG+d
TGw1a2Pgo93qON9KoZWGHPGV5T1ll/wdBdzhmA/N1eUAiCYZ6WrQTJd797eWCGu3vzf7F+AVZfXj
uN72DwtnFKKDmLp61Q+RklRZ9gGPNeE5/18hrqZsqs3bfqP0qLWhIwpxFabRs2gkNXP1EaJiOiAU
kXujLCvDEw4MTqIlL2RlyCgP15JiMjhxnk7pLAIycSYJV/nKSXHmKEdWhKVdE1fhSZbzJDzc/ndI
/asjnzHog7Y9264JGMldjH7W0lVmcrIoovtgtKl5LQjkEWDEda4FsmV/KGknfh33C4hiUt9NU8XZ
uL+SVvYAlu9RqTj70WcCG21svGD0yRJk2Iu1BYaoLpqYLlCxESHsHqWXCI2pTDIbrPZ4onjCFIDa
ZZ8SJfLP3f4MzoH+cIRSagrow92zAlnWpqABZWFPhMb2LLWrV4d1TblHrCQeOkBayMzCrxJMu4dU
ZoXoT8Na8uUyd/dPK4WsweKICtFyaatsmRViU0lbUHi1Z6VV4VAVO8rLSwKvCETBekVN3IbMHEDu
k/XteCPEgChRr7Go5eqtGExaBl530Anl2WRlAyTkaXlz9qboEKrH+k0CxQJDddRCvJCqw/m2IyJN
1mJVgGZw9Pl4WSuiyz0UNS3v1fB490RE40DBMfC4zLuBkXUX1mNx0aUOCjD1mEslVMUiojCgkKGP
DMYMonB46IU5Xsnhk+084gEDK66VvbstdIlskD9qEAuK9aTRT6okuKQXF/yLOz6XzQlmeFzA8NRT
6q1LW2ecs+FfwtFEMvgc9Wk9yXXbiDTsfpqNjJwQ5G/yWNmgbaLw2cJ2h7gFxjNfFgsYi3otXoku
eIkPqfIYmYdJ6T7qut449/zTbd3Qklbge4xiZVhUCM8+hL3wg3Fgj2CXdGWyD9mYTKp4YKYIdzoc
QqGjSk63/3zFIABG7Gs91zNJ9OpaIV38WNwzoaOcUwkg2JyoDcPihDOb0IYTIgu5O/knP6GazKNw
Pm3mNQOByMyqq/gwYQzO/W6E5+eFiZSbv+KMxA2EIxgY0mitBEv43IHcd4zLBxbiog1MZ3kmQFjI
QaDZC6VBR3WV570nle8wP0Fitzgz0rTPu4ZK6zgkaa6tGsPonrcCo1FOCrh5nX2dVvyE/qXIRpvP
UfiY94rPMu8SzYxmY38bltlADMr7cZyH2ZDSj4VrRXK/iSaTGVNHPZv0kKdqOWBBo2bYLaZ55Yp1
3vDosyfgzWJXqUnjnQYWzw7sn/5OF/cgFcxHCz17JGoijNrp1+4mXr4Ca10nnOyMfXkLugS8NNrp
pETz2erS2UYJb2xgDvVTZjx6qFMopEyle3L0WiP+1ZYxvWubV3+GB6lTzGYBI48u2qEYdElicXUG
iaDf16MxJLpGgS9jTau3BlN5xtLS2ietsY463oeAo696naOyUg2nhKec0iKCKXoa5WQak4IKXcx5
HsW7kZOggywVZ5Rp61GbFUZ4apa0ayvYz/tRJLCAurjClnd6gJxJXKBJvQQGW+OS4Xh16Roz0Igr
hfTDctWZ+dZXJW98mpG/cNA3lLDGxQbzIO//nxcTS03glzHHql/psMQw6l6/ZMQ86Vlj54Mo4rvl
oMYRYeXTonMJn0HvWcyVFEJEsdkIR7SLDoVju1vv5Qe7gz48kMQkJUf/dnX6W9vxxxo8kdbZFWXY
ze7q96L/OiZpSKp/+CgRkijl+VcxvRIfPHKKvy+u5iIDCwdfQpxqVrhifLIX5SnOPi5dKBsuLEia
8ZKLndlIFNOu+kVj5NH9B1+hMaLh0xjDu+KMVKaZjZZKRwWGtvM6u94bhCWzZO/H0F+Ch+zz8dCr
aNUr76UoRi+5V/yhXLdyOHRZXA4M/3NEjZXDt20+SlKo8RIYpa++Oem/9IO6amfCyvCMnF/tukKt
zmD4YiWPp6liFfl22J/nY+Eqn9FD2U4xAj200EsUP1eFJBKnzHUK9EuRP5ZzV5di/crQJHV3ctZS
9xVdh9XbtGPY3rdQ4OvAZsGdIarfism2QiO8hoBAGPBntK1YajepQup3E+2nHbdzcFu2jAthZbcN
skXoVn0bz/bJzQvlyOllrwxkWZrWbjZUYDuhN+WlzoEnCsinFIQN+r9D80qmD15B4eXVvHkX6HS2
ZF4J4G3dFY4nz9VJ70yEWGwNdQN8Yk7GMaRwVynt3wLU/ZaR6OvQbDNzmP6/hfFCwL6vfg518xWi
ch7MRLLwWN7v2EYngadXRMpkcaWHS1ZsjNq73R4wgHYNLXU0yi7pBKXuIW78D0aQaWEru5kUwMJ5
W/6v6VlyrHKNW5+GDobMT7x++PH2rST9J0X9R7yh/dfACm6/aKO7IWnUilSgE7ZMvXHngkPWKrVB
IePaP3lj+l4ph1tGNPDXcPhJJVujY26V3PV/YbNaxugXcNHfu7uJ/7lQIrAZ5MlbAdzw5VTsfBbI
Xn90hKCA3XpGNQhzN9m8iGtaOXzG5BuV6zsb7S1CtBeODkRByIonmkEoKrn1UTmr33kZ2Zh48TGH
TfIPcL5HyQTv76CKaYDeSuPFesdEM+ULzvVDr1O3lp2DtjVE5zc+peJOdUkBkVdIMcLQnUY2rqbF
VgAxjXf3zICVzHHAnJfs1wYQobjNi8b+kzBYmGD7hTu7tNMZdANm/086pGF8rhHOafejJfTC/idu
o4pSmf5OZsAXYI+4Xr3lVZXljO5M9p0GOk6BQbINVLTD/P398IFV/7t/tv3WePF2T4HwBWjYSDIe
WHY4tKNoyS1m2JkIrPcx0PEAPrjXatx0CQwYHb+OOIRXTKM91n3OXPf7O2hkrmuskL7rZA/zd4W4
R/w0/sl/H5DcZUf6bcdULhNrXYgxDsLOWpq5u16Ij0kIxU0R9bI+1MdiLo+PKVr9JHe+t1/3+nmk
2gWGhRJkI0mXDIUkpqZREOAGcn7eBQAcnl5XsXF5kiLFoy7caiuGlhxz5Cjcl1/h4U6PIC9LQmGM
3c20g2PXmxORAiqG/rzJFMGH9rreFHKUFGrn9ArG3tl3urTUMu/1JKrsraQkIs8j/wpNY2Uml6YG
SRH4Ardpg4ZZ/9o2DMGTnWXMiBV6SfOAfoRY/K2QCO9bRAKpCLxS5oclIU3FHYGwwpQ0CdNr1o2C
ZZyz2tlxZUEvJRCaYtry/TV7tlrOHcrS34y1Rx6lT8xRp4MKIy5RPE/B0uTfEk/84+WxR4r5MtxG
0CNl5/fWCj6aigUYMbFM6zpAcJKnlyVS3UpvBjPctWODTEBM0Z3iC0G03qeKslACJZrh93KZY71x
tTkOuW+irX4QRafGfAK4v245ggGObp8FvKpXPiJXHM3bjtJ5EK+bZXXkhGgpkQ+Klm5ZKzF3mHQl
cYy8AeZzxCGjS0d9cLMHip/xQMjyHRNAZ8/6P15uCuMkf6eIcQQBRRuhNkO9Et8XUBB4412rg2MM
p13VPw1w3x+YM7qIhpFgm1vXz26V3p//30AgaJ6Bbrjd28kb0n8fPdgcBtPGjKRDjNrSZfajgK71
wqrnQ7Elsu+jisQCpVQPPsaxNJKwx79JNmwNVtczIrcyPvGsrjfK1btWXvaqiNaPc+d8XHyh6LUk
PPdpEB4z8WIlZpdLBYCApCxXCKyuBqb+TCVGZK2oPfJNeY+UfAGQWud/IpIBI/Lu3NWgE66n9BdE
KCKk51truJ7gaRLQNTzY0nL8loUoXSU1yfvRlBMZgIuW91o1g6X91T/7WrXG5hgtys18uqhmTekK
Gldahp0VOTm+G4nxA3hJ8NWTacunkOV3mJ3/e2GaryB2+dXEya9DaExhhw/HVg0W3uhumOFu7BJl
DbTYGWRBcHT6TARz/5Ei8SysDgaX06PK3uGRCBRwoqbNSXdOGyC9+rUk8lv1LHVpcfIEXonrzybF
uYzOxlnbv2z5QuVGgAvKqnhijTAj7AEtcQHIeOU/QtSq5QrCH5l1lPeWrpZZzbisbNND4WXpvSw7
KcWFfq6I3AnBTbD14IGijHE7oxQ84y2IrSUt/9JnoepvkjiptwmMpJOFlu6kv2cXy2eyfbHOZvqh
6EyFzK7TTdALJ4Sv1VmvOcdMn8yNwxp3rNT/QzKKW6QTy0l6ARI0Ic5Ymx2OVt3NloIJYaEyFrsm
JH29NDq9aWRYsQLiy6OzSEmOEuocnchSgrhUFOncHd3qArICawwC/Rq0dUgxwlETgciykT0OlBCe
hUwP4pMxAgt6QT4bSD+NTfOpqlpEFhTyGahPOcMZW4bDGjR2igtED5PSAMCjYIRwTRzJKJ0hZy4Q
4f1Yk5hAVancN/kuWrq08e/BX/41fRljMpklMzh9Ki0b1xhhJeGbL0Ta7Q7w8j6RDgxoi//aS0G9
zYlKjF8JC5LzDIyOfWI9CMz5ItaKMiy+zGm0f7ZTjbShlMyn1E0TH8BpuJkfaGPdMXMUYTHY7eXt
BEkRKQNsUdbGG2Fbo4ABMN040p/5iSaItZ6y/sCmxhUtvCm3360DmQ2TToK8YNwJpA4WDmCLRbiu
m52QCSNdcZOHqbw7SaBmQI9kj/Z9L2rd7a4PAhrqTfh5ZCdkCSXDyaPBDGUArf2SUmGGBqwae8W3
NnqRRF94e0WvId0TIstGDBD24jL+H4Fb1VfGfKQszlIVKyvGM5YVIUtUI3UAPNU1qPO6QORPOK8D
VlKvyUl6ojTMBMDg0ICVmSw0xL1GM3uoGH5729Mi0XtYifDaPAkm074Jek1ryYyWp2AAYtpsQV45
3NabL+GFhvECZLtfGS9B4eX2TKqcq5Vz1bQfUjApRqD+V2JohZ6RgU2KIay22Qsxtin0qwvnNhKZ
9Sji5LEWC4WMgXAODW/iIaHQfenVs/4VpuCS9mJ0XvIrvRqJKrHtE904YGl+Bs1jmjMMLsrcs9K9
WJItF+tJPqLfwY6/MKMgJVsqidMcByg4Yv2e+ZUJbZG1Ow+vUq7KJohItXdAxbxo1HdS0DOYdqwq
v8KgQb/ekxY29kq1s4wHWnmb+dnC0mndyZGC65AiEMCaZS8IaI+kaK4S0eEZUcHgpaRAZi8CYw/k
IT9ynyTK5iL8o5NuHQ/xod5nv9XZTdbzSoG2Lf4OpM6zJbsuhoGx61kVg0rbkH5F68KEVMoMZ2lv
c3/qsvmovV2wIPbUYhPTT1eIfNKkJYJvPq5xL5f/GvQ93ies/VLakmY+RV1nY/u91l1dCJEb7wl9
WJe4A3RTs4Pw5NURu4y0LG6fR5ZO1LqcsadSrj0Ov5iDarsI3BZm6FJa2F+dUNqAm875oCbAWA1z
UsmQoz0bt/Ba5R/TXabmQsMXL99uAizgeBwo6MMHHu3OfYoyXnZIqblnAibZ4igpxOg2qVW2+d8L
dim0w7OTrRuo7CQjAew+n5UhcQ2NcO1YS+9utjBbDLwu00lFOw6bju6v46KxHLKN/+LOEy/+AKKG
ZYzAM/NiJbl22+EXJXLYIyBI178oEZnJ47AUCNXvkfnM4bqqWurTFeydohQ4DLpjgDIDngxjGJK8
203fcH9T9zO1Va+QRECaFIaMD1D9Ccik34S0J53HaaAE/DBzKHWtwSE+kVwndOm84eWV7bEzGpsE
qibix+Vac8wQTPNY+zpwK5XPAs3UXnK4sMgKMMa4lBdIb5ttfVhnuCnE7bCsjD4bTbqwF0ISuf8P
t0yuN/qOh5sZdZ1JENW3ribKp7YT0Rpum8IPQ1XaBWqwy9WZMw5zoRqIagXSiYBJfpqs40hrG1cG
cfEYJuDl3MfetsE0MaqCrOWl6p1dhWr0EDtbyYHchS/prc5yRo0OO0PdlYo6L0rwqQUvTOm4OvmD
fcnPoRU0XaNKe/CrDUSldWqrgSOQjyvFci4V8pPwU2pk/jGT0lC12ZzkddG/U0ciQp+3Eq8Mo3al
7kA4LQKLDV7YL6KyZ3FzYI5Jnh99JxkFOsnvBxdCdQZ5Mo+sQs6LRzuXmZ5/RNA7ee9fddx8gMwW
23dVIYLHnBYijyWDDX0NnNjw9wstc03y52TdtohRKqoBfudaDcd/c9HYR3/zIhROpRubAhkItO35
3wrNZK0J+uVwzog+OAzPmpE5qtqKM1QrBG2mrNFKwlqlwoD+boBbgigMg/b2n2qNuLuAvMhtnogC
LrdTOFqbJZUPr0zXNhTmFonTOrN7esV2Ryt+bdyIkS3Sk/BDozrFsDqmxqC/F6UUcnYobh+z7X24
dYucAzAhY/KNfj64mNMxnAkpQLcExEYe8tJP4H+UB06KYuwDIgPTk+I4KVk6BJ325wyxZMcZEa8q
2QOrzvNDfWAp683H+hp8VHzYliqhvCjDv1Bvq6owi36HrhTXPIBJ7DUPO3eCgYPzFG0lEYJgqoqj
q8ycbZoSWA9QwHXGp/xlgrZAVMbUZuQDAOvgCI/9DOlXts2hXMTp6ccPhBg4K4qTow8afQRXD35j
EHlHVWDwLEByo3zl65HSzuoQbRfp8+GufvtkmcJtel0fz9d7L2uFUr8NvQ7dTNxEukqs/4WGrsdF
KSDzg/YHkOL9Wd6dttQLoPJpXp00QFTo9mMdFiZR70qt7CbidWpL/KpnxHSH6VqZOh1vxt60VwHo
8i045A+MkvTiZtMmyj315p5TSPXBqbJDd5SvEuW1UodGdjdio0jgUR9B+zMWmM+8nlLx1pgRLiaZ
sGsN3n0KExb8OVHXugQKbcEZl7kqVlkHk9JOsI4Xrh5KXgEEOJyUv0VyLusnw07Jk5a6rcH2GYT2
16IteFXw0Pxg57Z9ftzR7B8JAbUVesf9iKhR9nYFuyJQAM49QWUXZEXz5rWNe3CkJ/qrlGsfMfKz
Fq9IPSriuIwwT232KidkE51sWA9lnCXDwseOi2fz7P92fLqwTMzVD4OffwZRF1NBVfYltbIeNG5Z
55AK8hAIIU2rMLB7hY4yTgwW+cNsBQdNGJkD4RJXrOegDqtuxLxMbKiQPhELBYIHyLDKFEY177zP
tUFn15WVlRVkE7iwKJ0qphI9NGkUF264r+MSHWfUiDVcRk5NREi1sV0pa+2SpDuC9E5VInZTKI5/
1v/6IO3aF4eSddl7oOMMhehV4wbGX5XnKpWHhQUdnQhvzV4brTSkD1UL5JX3VmySD5g+LN9by5Jz
UoZf8yMZjf1fc+ZllhP4WgFwZiBifs2zWU8OrzO9Bg241kjtYJrgqPk/QGoFBN3LKtvZy+f//kth
flmp1Jf8PLVulsH1qZgfVt5vvQeYDtrpb8FVXClinYeTHAXBi5I8CbtwE+v+XmAFsYJHF1vqA+Kj
Uver21piCzIAZj2QgsG6Tw+v1opdB0UtxqAnYJRhvZ0JjefCZnSL57PfrWklKQAi2ytFi6+/2YNh
f45HPn2DRL5FBnmEaOLlkkyyen0Kkk6n0YMFfW8gANa1pRoAil46Sd+3IsunKcRYzFqAlc6fo7Bs
R372lxUh4+VhYt5aMn1xu+t/5X6lA6q59XUGNJqdsdQz+hoNx3bevXf5vIQv7DRP90nkTTAVb5jx
JYp1xK7bfAQWPwbwBJBcd9+91Ni77zloxTtc2f/Oa4AuDroe7xsKzv4sp0ZWbT1uGLSpXSjwRPa/
bxlsd6D38wlviBl2LrEdjRvZAlQ6BsM52nYXFC0UlEBTokL4o6uI3aN9YJQ46C4DMEcTgjvV4Ku1
rjZWAmzdEhfb5Aql/k5fg6WRPkDflSahWsG1scp871nvj242KdhPyckM10L2lJv5gTqGFegcA4wm
l6XQ4drAAF7/HIgzYfQ62i4bfU5XHtTBJRlEXx2gjk4UWlN7zg/6XOQRC7vig5wP9lBJk7+Ss+/+
5XHA91xHKWH7N5hPsUE4U0oEJCy5r5rvNFOpVW1phpeJdxqcLwnUEN8hBQill73nvFoy+5s7wlVP
EvPQmGff7GVYje3zakMnXd4FBhztsDOHWXaJ7HrdGpZSDxgtxQOAzlZtWgh7e2NirajNha1pR4y0
XlyTuGur06UTHxOMESX8hZQm2GfKVpvi32aTKqDa0js2va8jQGOCaey3FAYmsPP2O5k7MyI2Pg5/
nNZTV4fGZQrKGgh9sjSO0/93HQZvVD65U8mfxBmC2vcN+uCsAfOZbkaOFfLYAOtPqUcGmZXoKnEU
tQNMwu2dWvV7WNh6U0+GZQ+uomZle3OjyrPBf+PEokvoqADXfkeFP9Uo/l3ECsCPP95J7xjTd5g0
KVU00Ofo2U7MVy4Z2zbYc9HIHZiUdO8c98qqNW5hmIp7JxcGhMyqMuP04lzv1MWwhTRnqLzV9oc7
ILdH4EZmuM6ovMaGbDPnLHmeNTKciGEt/rOUzyliMn4LUWrwoBEk4U5mNV3e/PLN9lnpi0ufobop
eAN308P0uyQWaMB4T4IqN8Qzs7BFteoNpp5rA4PuogMfemaKEuekGcSF/aJLYkT5xPW/ERVsgNPc
bEjngvvwwbi8CcOvT4lXMP5QSCOzaxihd7jDQHfLx/JeSFseNsnc/WIAbjAOq7DGVO+IfEccXOH1
glhdwwwlYOG5Sj8o0eZDIMobae9jzt1Etoj673C5hyunF3u+wJVAVRxtWDSkeocAvb8IfU+gNSC9
flK/FvOpOw1o1ABy66JthmizjxBZnNK/grJP0qsqrJwHJPhh9LqMiE0sP83hEP/TuVoXDrUSFxSE
SKO7SkJJOaoPFX/5wz/OL1Mfa4ymqyLaTvxRSmC5a4QUsx09oVCNkY3mfWsx6ODaPdWNFEk79vDD
6YU2IOwfF0fI8FJ87D25ZkSNSoFs2t7B/QijYbk1JpxvZwcabJi16b7xXlN51InsQpRMkk8nNNep
vKf/DAh/buDabgS88qgM5/MWpjw//0oo3GSUgctR4UH0eaMtQTL8uoCXvxMntjYQVqKft/gM7bE1
/VaYwNeg/GmK7HFj7w2qxfixY7WWIWq7AN9zrSPG6jiWlo2e54WuhYi+Q/8/3hJ+rUlhHrOWSqgN
FCTUz7whdprZLqf/2jixAdtxY3WaNpd5OA+y9vK+D5fEfNFqfJaCaIegItiex1r3u20E15XVqRNh
ootIidqNjz44LYzJb5ic2uywETBt3v4Uz7Pndnqyf0HhnLaPwmDP3vGymiLuJ9HTsiHlBUgAtxGi
p53FzTvFX5EcAuNvmabg115O+yhu4JMDL44im9bHsERcbUnyuPG8bQBjO/NJuQdITWtrtsEcbVtr
OXkICRo3lfhLmbIE+pN+q7bfbisAzbPng6YZhcgZgu3LgLaaRvILb1k19TPbWt971ddPd9SB7BFU
T4XhkIJGZ4nd5iHmjfHRV9CowfL/nOxxzWYzyw/SMK/B3WogWjaCMQuGPQwqh6N1vDs7Zhj6o/WI
bwOc1H+MIMMmDdBjf04kvJ/Nq8B/NikXq2yN2tvT9epSGBJrNGGapLynjODZhPR9Ph509rE4nBel
lRT6OAS4OTYIExEQuCUMUXBhI+jPiPRcGD0ISxTR9O1fn/i7klSOlx9fcPgyPnlodm6k98hYKidq
OuOEXxaT6aBrZfXRxtTqMg84gEvXTifseoDc/O6MXFugOcG7/FdWW+njbR+E7NlGktKy5s7HmFRN
0BgpuWYIMp9KtdIXDH7VUIyMjU/4Im4Cmcs7opvyO4h3HO7uHEkpeYGXifictSSASXPfa1bahCU/
4KAgHQPK15+FfMQshYJp8PaJQOq0hnpg4zoN9BtC5C0LoksSi5LbJlruSeLrSeS4f8S6NHbjrnRA
QZh7E2FueipwRjV8Z5BPLupfx8NKd+qc4RiQVKU84G9Q23tUHVotiohvnwSZxPPCOL6b5uQK3vRX
v//clnevqyzGNuxVkYhtTKUNUqavRqq1qC5BDWml4K6ycy17f7RDQXpoyeSY380ZguaXLFSb/ldh
OQAb1QZWKYSRbIq1fY1LH3OSJir3MP+oi+Ip8OJ1XtEYp8pWWRasJloU0rdOg8ASU6xBjjME0Gv0
rkLO1Zxa8wCLnuAC0VbokB7HBg79S6PzKML6/QbwTtvfMHSB5OUFCTpXCu0mLlSbWlBLj8GzTiaQ
NbGs8/wTEHCXc/7Lls0beJWSXBAb9HMqweCD+mn5gDZsPLZ1ckPAO7Q6sBnIvS4uiKUCW9XDgzwV
ZY7snMPJpyHwEWxF2k7eXqRQapfMHSNvzr28mPNOpisOWOLy50Paqxz+097gUKMSd22i9CjfnOru
cq6jakLrCpqJgKjMP1bv30D3HpcJpOG3M+A1HCpeITAUBw/L6ww3t40PiRLxONdI8JJv93uNkOG3
b27kvf2PaYR4OElV8dElIADxvmsD3HXpJcg3b/DV4O5YPsNguu3RKezHcWkLvi92iMrhpVCQGZq9
WGPOvYa14H1wDGF2OW5cmfMgGW77coO2IbhyZ0D90M0BFQg7Hj9yTzfW27l+iM+SQx20kBVoxcfz
92K3Dky4F46dO40uwZ6Ayt28WahpPnI4Ui5LqdHWp87w23VJ6pB5uP8AhrIXrRQvUmOaYItxBdMb
UwKoirU49K5kTjDqM1ztSBioINZCBTjCktp7N4ZM8NuwpN9Eg4CHJzJQ5+Xsc4LO8Rrly5bIUKEg
83qEbK3IyikfGHpcCcll65dTV/ZW3tjDRVFSQhw+PtUc9orv3vrOPJlr2k6zv111GK5csACQI8YQ
TzW6mL6JhcWSpu/YH31GcwnUjgMXEwzOB2Zuw791Y6ZFNCFQAI426FYEUVb/1YjnClnC15fxO4QU
ymNm5tfz96mMcKQCHl7nWg8O6OP2ZlBCD5tmf+q9xoynN22zGJAOPFdK8AFPgOr9CIVay00lbu8E
dFD8za8mG0FmLmjRVQSE2IVzYSIPSplm3ZSnBA6TWlNBSwpqDQjlNIWK9OaeIpMxS40dwIHr+GDC
OnAv+97Tfr9N4+R0thrMemmrIbsCRLDV3jhAFCkRBxqYhTjolGcfzoTnjRCmyYtuTIfmWgwu1nFQ
WnKSUMBFJpsf9qyXp4txYFbay/5XvVi3BxG+OIoqyQGHzaJVCGcU7vALymx4ODR/wWE0FQmbYAwd
bLENAKT1nNJvEFDC9RLlP7dWx5H92ln45rW+VjFaYEzeEoxrT+RBhqy70LHnQU0371IV1mSjr6s6
cQRe8v4yY/bMIuexfQgE5AVrJ+5e0QerSaccp/NK61FefgO2uZ4RyG+J8rNNmiWgprTvBScCHLJr
z3VVIboqKNgXo0ey7G6p/cpMSpWvKaBsrqorVi1+Xv7GsAtvBxCjqHbDfr4Uxy5G5FmZE06lnzjH
mqJu4ye723kSpoYT0iRnpHE0Joc0tEdcd72SQXcFwPUYNljH6ax27cP6FkdpCa/NSzVWdv2JM65T
yy5khYbPEs5DWaG3loc2y2FfThPHhP7P9rOTNGyL5dRPExCX5+5ZKf5Ij7uWqaa9kDIn8f2jmoEt
u5yiVL9Qmrmkbh7TmfPlR+5lJ3y96/cGQFlMTrfgmmJCnWSVitjtfsMqyug7aZhXm/ppf1xbOmr0
+sGkAov2Z1q5YkqX4vTPgHecNO5O/KT/CLI6O9l49G324fwz693FDje2myJ4ntJG80MMKjyFY9nZ
CM8C2jiTWcWoHDiTwKdvVJmD26Gt3kb/5rB6tZ8Z71sB17d3/c1ml78R8YH4l9qBwmE9CzwXisKd
gMdNLwKqsEHLfiQkSpfxE64r5qBzN11tasOhncmRCgkrXbc+zkkUVuFH/etEf3zqCUiPIjNIFxXj
C1l7BTWkSl6v/+3PL9UZi3MsY3xnyBTMgU5jOop9hEIcPutIoZ1lUAuOnE9AnSt3fYFus3vMP8E+
Q6LG42d4+9Qf/NJjuprNozuaW4htFOnM873dwOiM1FmBcPEXUxfz4Ms4vu/+uXunnJHNDkTM3hDg
rTSXgPgayh1iKRX1r4YXaWo9LbF1YdNeluYbh9iO1uCxhjHuJnC58oUd1prevcDzlKyO5yANNRl0
fovnSCNr0BeUi1trmpwGzSPLCEJkY73dRWt0J2zKSR9jtKNfI24fz9LfzMDDnTz92HNB+4qyDoH4
eiPT7I3io+6pN1yyCXzZa5znqoqr6Ae04pvku4ZxmkSObVsL1sv6bLviso4FZnXcwx7N7s5Py59v
8Fg39mx6iz5xcZ0EHEgcx5K/wxk4YFADci6VVbz2mDfQRDvXIrE2stPGhkJumvctVyBnMGhT8xez
zUJZqtWjkIRHbiPaoR+UwINh7ITdXL7SZojXyx106wL3OGq1VXdE1ninXnj6vXFPGNMI4sz0RA5z
N9ZIhhTttj9DQmxFxv8fv6ngQQCxdRUKXpg7ABTnhDm5HsOLCnm05hLH/6UDa4f1VUjkoKxCNzqn
9cfuzV4BLf+T/neUhY3LPujhw2XBxJac6BlCQSquBDOG05G2S/VHSLPgpwSqVSL/R0Hbptg+s5cI
Elj3M5VFFM80G47Kmu4VplelASeF8klyFq/us1et3Rdk/FI2h9m0RuLVK/+czmrX2hIvvIQI8+O9
7uuyuwvgIFqnV3YGLqNkWXWG1QtM6J2nSZ13evVZNnkfp6qQ9FWOhd1+nF296iAmYm3gXiRvzrpu
qaGIiey9Up7XOC5pL3OE5rRGYO3WB45KsZQuHXIuNJVOo1vb95L7pxBPmx3zFKBtWjj2eAFuBeXI
AcJCi8Uqo5HfbWDUO29YSGH94elQO/5tzg2WBMFwC1McLl2uoyY7PoS/dTk0Nlzc1nMpPn1hOgpA
2DT8QO6VuZScBRAhi1QbCvYgnpoZ/2eGhfXJaivwPFCXk1GKgl6DWri/nsA+BEXZrasCuHJ1n/IJ
k6Hj6CB+xpHO1ZxXpy5q8rYDbs2rRRV90OUvl+zHjLeeyp1PRw4ACbGsBwlKbqaNLF5rM87YWHyC
F4R4Oy/VAjpjsybiEMIeaEajoMFltDVbRJC5eMKXrzTVrgOrqjpf5l02SKZj0A+8sjDAFa2d3054
adDruIpSCHCgM9WvFQKS/Lb3Q56y+OcNB2agsNz7rLQS+U+9jyiaUTxIg+uZokHS8uFoPstF/Hnz
eBwTxOGKn9f1dNEPGGkggvm+VUtmOGOFJEwHWkayvGnTr138QZ5YtbE+LfsI1Bliobrt2d3sX+Ju
5Eu25m4lLCmNncBJ1+FuoWeENIX1M8Ib3wZ2WakjKF4w9BXpFR1F9yZW7J2ppCie4eHy2O7bDKCK
HCXSRhkLJf6CZauK4hnD2AG75ZBzLVM79DUfpLXFleFzAqn54/K9yWJRIxe2gtl4moKhlix7H1/z
BTyICWqfzRfT07EbHzHCrUhNA3zHvzmsHwYGamZKkcjnTqBwdbQI+1V63wJTOh4lgiscsj3d6e8j
s18/wwFkqhFbHVyXptZqT+8faZrY4GQ2WOv1EKI5K9401YqBB8NyiuPtOsdSLZCw7vQxN5u6FQ5T
eE6wC6xMvaJhIlvwIkLVL6U6adFeWeOjVhPxwYdaH0eRxFLN88RJEERHDjLB7EaYnK742RTA8YnC
RYYwN61HuWMqoRA9V/qccf2wr70o5BZVg2UuMhDDrd803PcmKdVNT+Hlvi4QW17AHgePgZ9rqIsX
6M5MxAZywSpec8aDxKgODBkp4FhBWWpBOYgE9aRA0rAKC/HpiCnuJXuj6hyu4BmmbQGzvACWCExn
akpFUNKHWcXfostslTDhGsyeK4hH518V+ejX5rQcGgzxKwDcDGYN+HM8ikZ/hjP6eIAIEV/tD30W
eI7UDbnvUBeQiWYogM3yNMIdOEZPd7D+UyqRh7Ar4zOA6pxnZvQWr9DNtiZ+Z7HtnJoNZr+IxUGM
cPUFWgB4U9X+aEOcK8qIBcvMDeDXtHE1jF5rFCxZVIdY3pM02k0Wv1p3GqVo6X8fl2B22/lxoHCi
vjCXaXHeZNRdfA15GWpl0iLjk818AIOVelD9UMBupK23S+XPp0qSkTyM7bGujDjvLRV0TiY/OfTD
2RtsnlOtcyjC94yLHYsYbXFWC0dYp4NeYJGaorPVT3kZgUpruL6uQj4BCQ4sCAHbbRzmHamFrzAl
j+CdE3iQR3Sehk9CDcxvPrA5ZEI+PHrdWgxrxoCBEKLkhbhVD4SOja6WDV3akxENxkga0WMobj5x
1S+j0vwj0HY+Cwp72idnfCUoLlM+iXgw9f4yJEhbzHDrafLglBTxgcNJaJuBKqN4DqT+/hJ/fYHb
esjh/TaZoqSAq8hS5dTV+s6rbM5Q3kuti/SEtNr+FJ5TADry8pHGofC5ISI/erVfTpV3MeqB+ACo
qzDxbxxWbvovv0y85+ljhn9a7sUhof80sH+TNhqjW5y3jQ70BbLTsZC/jYd3vXcnpWKb5oqoIc8+
cX6pT6WTkr39aLRnaTjH3bDY/24VkNQPTm9I8JZ9Z5RXPixc3YbUnNsMxLGcTh0GnoYPamlg5/wt
TKDnw5QiixvCFo4IYtWDVckOtwDqNKtWotiusQ440tFw7VhoXErglYoWasiPx0fphkaAXTCtt0vE
p/9KlE5+6D98eWOV3aHzG40XBN0g9xJCZlqwhoy97w/NMQq+YzmMl4GWwfaPzn0kMepYFdL0qS3+
eLt0VZFU+bOQedFW3bHBYDMeWbHTx5O8DpB1jDhnhcJoq/5W2A8C1HpsPrMrjC5lXfYSNDpTzimk
4ALlq+8bPoNCl5Dpo0lk6YBYSt3aUeNi/G7An3/fl4UjVi3nXomgwmt8CjP9MlXxzspIhYlPsiHj
pdaRWlT4dfEFvtaO/PxTswQbKrZZlupOoQzZSyeA9HTJvAyb9GDNz45yttki2ISRYmuBynK3pr/D
bOKK0cxHC+CPY2Z92NBjy+PyBp1+Iygn/0geSK4vEayU8kdyCeNSYdLKyZo5q1ap2yOhSq92wuHx
8X4TWY10LFcz/WBTOASgLuQoMg7jtMVRw5RgOwLqSx58BkuE0dKim18dZZlWLVBi4kM/caCxOwPg
EqRnu83dqmK/ege1CQe5YKGNhQxOSMvd/Hkb4cJmHYCjBZdvDVufLmXCK4AwH996KzTchMYqLY35
Uu6sZiA04XmXspniYogHKBrH8e647xW0j3GpEWwjxCZRS5qkdA3qFSFg48iBzoDpJHidTCLVQcR3
3r6iO4McXEiY8I46X1JnYSgEeFsVv5gZmK6Ytdicg8g2Wb8LXG1ED6IbDQ8nZxRFkarhcnKQ4BZ5
LS9xqiPd+3M00YeX9YZXbr/d9IUJSTKqG0aHDgioUM2v/Bs4VyETPiVRLLUbRm71RcVxU2WlQfzB
NvJdhtDiAObxbiPwxJ1pSdysUDHVq4ndtLr0D/XX+AqTkOppOZlk+s3QM1e6curmGtH7DtGXpyjm
fLn+zl4YtYETHcPK8Z+9YtQ0zW3up3NYdpPvaWXnnsem++pDxLA89S0Orsr2rIE0KtTk2olgg837
H85rKNfDsiQevSNxHlAo+x0Pa2KM4NptKe4GOJlohNXVUrIwyRs9FABp+BiWNrn8PO28EGYeRZHO
yV9ghqH9+6BJEdc111mF9WgqBs+s8rMfyVWsMufKSZRkPY/Uqb/rbYvY+zkVus1/Ig9iWal8gHTy
CHTl6bEXYckfITO5GJzS97PZ/oiXkdpeqGlA/JA3FStq5fO/4LpQ+6GZq1WdvL3VjZLBEBDXiy/B
WyiOVtLEr2BkIist71itqQH8WxCGMeRIpCILKDa4HXctPIq8upgZbN2LYZxgofTSPVUHyIO2UpK5
KhgdQ/V6dK/qG0DAwX8lCvsXmdEarSmrNaVshW2ytGD2+JAGrBe0rh1psZ8R/jko/NYe4TW6RL0O
Tz0B5b4vI4Q0I7APDAuBMWgitVnl50mWVB9OfDqrIsKYDN1ZrsNaU/R2t/rOBM56Mo+oZmugS01b
4FH2UfzKlaEDDt9fEaHKBVT1DSTtu9o6+rotLgVUTkFBYyflE3ZKYbHrnoP84tVTkzHzcOKH62mO
6bENnhwmDG2Q71SfxJ1fxOdn2RlRPn4isretp2xk/DsksWhgVFH5dDSgENEceI20JsktUZkMIyyg
lIKb1wJbJnGYZXOG4U+fsJdUIpZjHbTUDZ9CX1Nxk4WRLvT7DQQMy3fULk9fJ9hYD1Xxs/oYZfwI
/35wdw57rzVNjKh6cdM9mcc9mk7MmWvS5ue6geKtYlvX5P0eRX6eSn2YOxH79XRUhIwO0RLQKwsl
4nidzJIHriKicSmCOE4khGBLq026saDV5rNPiHnFp7d28ZOrOoTMZIuGGZbwM+qiUtbUxzPdURuJ
pxqyT12qhcYOCmdcZdfBK88lNNxpcY3kYRWKTtScO80ih9NkiAocVyi1GKBDXADE406WMSfvAdkD
pGen/ptqYCjiaqlE2l0n3Nk014ihrBxhb6ex3f995HFpy3E1FvrANvgdU18zHVXtKKZFeic/Uoaz
5cbagPgkhXPYc1hqPLR/wy/l+pJioFm6r0mnpnIWxFnjIPtQcWmmvGbxImDFpmYKDn/UolJlxm7a
Phj2OsPzIFRShXYVbuxkRPdWQgcXRI7lXOT9w6JgAgf6chOCFo4MWYF6sCTleS6bY+o/KeXmwLsn
b60xJ/T+7FKmS+2huS1U5Nb3FEQxNUut7lNw/3WgY2ghtgIJbl6faULE2i3d1nPhpmvYZam7ZoIG
U4UkGzjGZE7ZauUxK8tk4CrCCFSQoHdzKcaVPiB1NKZ2KbhgoWPm2e5Vn4TFslQDg1733RoUkyzS
A7ALYRzc5VOaQHSy8SG3bRRTgMTXuPuJHStvx19/EjHnqZVf4QMCbs3lMhi8h6QZxRn29Cog8GaW
QOk9iEunWwFWEV0dOrS+VxfcrctFzHh3GEsJHYa9J+bcer/Txcd/r1GGDPed68y01ZN4wF6EjPGN
Efi9MrUZAk7g0ZrgPjPapcSIotZhoKdIZJUW39jCYKPWnBJqwz+4wwbN8qsJMSMQAl9NJXF7GnKn
yXkL0nwDe9zPfHVNxR2LtWLI0HFfEKo3Mg9kBW1Nyz5wpuk/dTtATaAw4fAXoMzogheo23bfeQJq
2RizjwPDVulqOODU5FTPvu+Rm4jXljZXq7X2MeZnIkT5ZjxaQLzDM0/mIqQGg3lPW7rCM7j96klq
+1h05zE4ogMgntL21oEJagzHGtei8L18CyoMckPuoPdktIvlVb/GD9ezWlHVgyAI6CQsiDvSV3Va
z1kWwFVBtH0bH27dT+kq42qmWknRgLReQX65eiRp3lgWq/IGb/93VtzNnSDdtPM3i0CCAMnWniW7
viD1YkqxutiL1+dSb9k76vc/lAIuZoLRPwTYBvDMfwWxX7lAi2VTXbIAj+/4KMse137vQYFvrEGT
BwSkwc7/IuFXINnT6zU4Td1o64GErqtDWXKARgrc4p00KMlGCU9nS93EcVtGr7Ac+RYgumjI1tMq
Nru5a3hy4coV0PzCAXTmPEcDbgVptVvwfJZEx/p9wCUrhIJGTcCcMF98nhmqc/WrMs3Z/YQ7kp8j
mc/9cTS2MS97kXaQ2We8IgwtvbobcLNlvNOYtU+FM+P8bnfEFtwDye6eoQ9no1JtnslR3l93AsNW
HL3lu9Afvz/Ps3VZOfaoW6ytP4uKFfACud41kuAnmo1hGDNn329t8RPIsSYUH9GAXucdG4RqwVh2
CaRZg3aHCtyU6GiBlrjTyIyHv6IYkh2FQB9hZWfsPLnja1w+EO6/fihV8XOVrKp5+Q5OiLdvcKG2
Znlo7cVKEzlV0F7n3ubVfTzJ5lkA0EttX4mBgEmoQ0NZdkQyTaONSjtNhRUR/jbd0sFWtdZMPdd3
wvdO1UkxJq6+4rqPApJ9VPX/TcB3ZAlgVWQoWc1OHqz/o24GmWixFTrtj2lGwyNt0tKAJij87uP7
RkoaFyn3liKafCDlX5JRvQk/Ei18qv2/Fb1FIGI2hR9nkUE6p/Ow6C3lRzXV8QNSOrBWuVECo1fh
lR6k1S4gShPrpXamgpZO5+u9HHKlq5lAMuiEwPGvJ0kqqWSoujXE2aH/Y2lJbjv9vyikmgY/o/jh
hge4wkmRL2bJ9jgy8znoeUif3pmbmsn2MkHgYgzU9/ebdwux4ezoLoIKag8JD6JGTKS9GjXQf0T1
+6a+fSARF/gt/2Lsq7UzeaZUnO/Nj3eg3eHCjfu6sS2jS91h+nqfhDrNiDyp5KhnVsqS86JbAAfO
ur3w3IfceXNekAp3nkF960tl0qDt+hiZ67yOwJ3flEZEYwSIZvGfyUcGkI+QE0iHtdUSvMYMquvz
x9SussNzytV8LS6IXMk6Zf3S/WROYxvslyzsby9VLwKqCOaeP7OBQPqZ75oEYFCd3y8jZ21o97q7
MINNAaUoFGWaxlIsPIH876qKT/nCPCjahK8Dj8fabF36/hPjXODYjrXczby/r83dA2P8vVNR6rSx
Mx23CxqoYNNoBEhOdGGDF59SSmfnCZ7SV8VKFAq7nqu+9/usOVDnlTPbsdmjGCuHTfSiSvqPPPeG
63E6LWB5Ad1EBp+TKPAITUjsKmqZpuaiutrbmMwCCCaeHzP38YfcWebZEERr+2CQ1y0d6sPvJ+Sg
bsHwtXhWZxJt0tsX0tYc6tK32BaGSmdBc81nkIk1Xri16NI6XaZxmK0czGh1u850TEhfpXsPptJ9
RDUUhJQ1KiHt/dpcy4P5PaNU4dp/XDt3UON7yR+zPO+Clw3sirfxFhQYOZoAqK/xe4vJUL7N4rOT
mJigPXHv4VUMmiRm8fkw5dU2EqI9EC8MBET8M9+ZgLiUf4NjuX/PmjaamE6cLNNvqZVd9ipyCTu/
/GcPWPuOT+Df+bWCh5hdw63g0YrfxkQowWLfklMP9oIQtgufejy4+ZFgIytex6t+UPMzcqY1nl4r
3Y9VRHM73KMpcyDXrUckhMXzFClFrviQAmFEszR0KMnRtMwR1ROpi7N3u/phs7oyBG3xcdjoVvCY
hzO8WcikfoFrKGkW+s/awEZ/rAqVm2WgdT7KAw0WG9y8gcEwvuJdfgGwXHvczHcceMLq3puyShWt
Fnyn5B3s3wl++MVgr9CqL2nJQEmVL4utfwhPAF8Qz/0Fh7MC5ZgSjIlOQOB2D/MgySOvpieJHEFT
8ewV4FofZ5zB7Deg5jJdkMZ8rtKsKoAG4QlMI+BbvIpgYNLwBv2z9E0TO7ktRUVH7AbCihszL0ts
eKgKERMujZUctFBU7jkKgZieMQbNq6Lrkc3/EqMj5u6+4WdcdXemO1rLj4mYBrMo8yJu3SgL8/GW
72YHI7717Mh0gJFQ1wyXsCr4ZY2OiNujY71BiQappyqXQtp7pKnJo7JI1aue8kCws7B3iCynfBbc
inihwXvSCm6rOJBBT51GGrFN0+HzPSG5AXJud73MxsSnp6dl5I4f2lW10YPo9Dzt4rcFjdz+6lXE
Vew7ZXrha2D4ul3qGUIFQpE6hCbL0k4q1Xh+FTvgAGu3Ln4wkykmcQ4gSKtN5mp8uTP+PrMBlT87
vTB+mk3GwPyK0wop304mEevg1ZYKya3QdENQtFxCS5+j/i1ul93T/Mquqce0XYhHyiWWPhcqxkWo
wb5gIv0WDXW/HBXOUGRtNqXHh3/3QivtoOjyI/0Xhi6ALc6pAR47cCPkItj7wSlh7hhfvscoG/36
DxkdUyI5rE9tvl3+qj2sZwYy/lXTNob8FO/imIezVsLFJmdjkIM9bD7xJVdNi9q/rmZz0dJMlShA
cNDR/MfPMFcVnvfUoaVZQDDKWeo95Y9pywqu51Jq/m+LSs+Hmx2A8h2qh5YEcmZa76Do048Fqrr/
wN8dTQo03Phu5qKWixU9Y8oxcN7IMSsGLQEHxaX1u1RaMkp/U7um1bGintm1Sr2CfPMGhsBF81Zf
BYDVM7XDqS67rfyKorqmA4Es8922YNvCGQ7sGPPYMaE/IE441FVsWCYAFGRFyoIIM3/ax7atJIu+
Nwn+h+ID/ZQRokM0E5RTjFsfkpRrIGPQpr/0GC6564DPbTJD6A4uVjbrBtHB+BvfXc+JcbDb5Nnq
0KjThWJlISO3n/lwSlV/sr9kSVP6Df+8pj5Aa8m99KFdbXHHk3Z4vJq0517aQypNa/eRDN2vk2KI
QzrnHgbUPgZb0g7DG6U3EVe8nnYSSMEu2Xz56nrPphwjg+EmKfs5UVFkMLFz+wZSkkz8dAQNlBTn
ijNcm7DvhETXbsDcXNu5UF8CBakKzPyM4WLIqK0kGDLXrdRpKY5BkvujBj1iCqWGXBPtnGEbEAtZ
HO/RM0ZSrhE0JRwl/H36Nh/8vJekthoF8X2+4Wx4V5/jHmBA8WM5W43G8lwv7EVXZn443a5uU/yj
RNAdsREWpLJLjtjIqpN7mEQUtWSC9ra2pq2KvCTWxNAFqYfh3dzylLPGVhQwSmcdZhb1ZRTPUFfm
7mozdr+PMuAngNHqeyrkW+Ir2jQhazvdds75Iw5hIRvnpMUrIWk78attff4IL/sMVOXaf8/c/o7d
9xBU0g/tBpVhor8jheu+bbz71LnLMkd6+Ux6kCXI8NZwYW/QAKw9/gY07IiS8uK/jV5rjQmYHUH0
vsRkCUQTzrIGZ3k29M11+rAtW1+fdt9TmbXVCdzSLGWO4kQcM4xQNOQxhl+cOaknGRMqr8EdZQJL
vkZ0IQnejGCUucgbA6LBLSFwGjTzBHi5TZez7B4k5ogs8BlcL6AzUiJLIH3TE9e4iGVAEVUD8IXd
3fuXCBRpfd6TFhZTIQOqtG9yK/gC+D395ut0YU1omDT5Z8FnPq6sYvXmlRgJK/1KG5wzBpLsjE3z
k1TJcG5Cy+tuyxiOxaqZNDve68xv4klHsDctRw0gzlU0wcvhUpepkqhPxpRvNVjzxlOC+MCnzYtf
UcRRMm4j6pZXp39mp1iO8NifB0xNbFpGFqNDu8OHxnKWvs2PmVVmmsYaTYuv565yKUyfzQDA7Xy/
CPf7d/TmVYqXmX5b18zal2uiZ6hC6VLnJy1IMt1bM/T9bmy/uPIRnhRjKjttdAZnWw7Y3LiUPBj+
DnDbHkjolqI4Sa5+zlkb8cG2GCifXXtSBAPpAM5tzEPJ3OoQ7C4Gb8Wo1Lb7aCvSoilBh6BQTNXS
I36e84S3QNoZOOEqrcB6OV3WWPX9ms3fCllukbR5oVrqo98nsjOnsj7U+aJOqk0uS+4nGuxoHbMS
sUXnvyF7OPpY8Wo3LZqt930W1SZsoMDEucqzsUuz3Sk2ce459e3jH8ZodjEtEf5uOsMAehNJwthe
RlErzG3F4zMNTnTJl0vLLj4cFHSnpU5gNZ1c5ARnQZbh5OERv4lLWQACDgBhOlnePok2XtjhcuvQ
KGV5wdqKd9sq6i3raPsCFHqHS6k5ivGLvgP0n3yqBRRIWLmGCAiMcYzvTg00sgfSmpsswzA07Hys
cHmJ4qvjje5Wawwzl6zpCW2k+rAzWFM00G3LgRWVG1DMGIlm5eqiVLhs515PY8PXzsCzphcJNHsR
v4WUAp26sDh2BHqHi7qxTOANJJ9LTtLijNvva4P2cI5INQDJ7jZQYROyJDdAUT4gMQicpeVDXGMj
E1Ababth92hNTg20R8+Op7khoZp17K1cOuX6gr3+jwHQSU1Dh90PO/6ZvO8Fj/S6N2qxMpuBoDm9
TtlIKLM/fyqv3oJ16vO0m12qmfWha1xv1Jhsf5cmG7B5wb4Wf21XAw4+qbNVpmCkiZyP2prdqi02
Y0ZyxkSBloApC9a9s+OL6sQ2qEvA1bgUv83TFUDk1Bs8tMaTFLX3eNPQVWrqmol/KMQRJPGQYUMl
xHcOIFcxey1veuYPhzjMt9KbxUo5U4yVKIRA2h7643Dq+tzTa3oGuq/X4L2+KA5yErCWNFbBLkWo
brDvWSyg3h82iDqilP1on6yAn1dmrn97MBYeSAL4CY43J9K7KAxW4Z2pOHIf3nd7+8txcWAX8Oc6
pr+wsmOZfxOt1Lq6NB6gxU8FitFaIqYAiVMRipncoz0d258FRu925r6MQeWhVPzJ4OzA3GwRpi1G
XzNdJGoPnljkPz5kZXcx/L48AxSs6W6gdjMUms/mLuRwoDxYd1sNJYn8G2n3oXh0/S3g8L3ze0r7
25J6sWBz7Now1cQyjLOnmGzZ6YJ59xeEspXre8DYisOIj+G55RCkQry+GQdIS0ikjh53a8nhxNWX
LbDc4FdXr75tNCfHp4/Cb3gf+DakM6PpnBrxfKkUnwhn1ICycKfuw/v1VhE0hS982yX3Kq8wGgSS
zXIM+4iUSatnR5JjtU8SLotIDHLBGSOqzrEYvAFCvUcZO8imxiWsGOXNZ9CsfXh0S9PEEqzwVzRG
odvDOrR36HPIZDDbdJVVEyuKjSR7YcolkPUq15zK0HgmdmmwbRMSNPtGNa5axeccqRQA31NG2cn2
lvXPQUqeySsONN1uPb2QyFhKwBlQkC3cfpLDotR6uwxXCd/W7u/TBwfMzXBHIl9P1f2bFMc3ZRxI
XwRECHROY6TeDJLiPf0rT4o1sg3wVYV/IUmVIMzyVM6jPrtYdDhmcjqcTo0I2sGZwBuSW4Pia/Wr
hUiVBzTPRMKj+miVmpxaBGZsaU/YsBaR6ZfLzgKp7a17vZPZ4AU1nAxMi8shWAcFRsa16Zc6JyPr
Oqt6zWh2z7RWsLLGdFDIbfLhwvv5+hLJ50OYBv3ApUVeCGWoc8uZkmU5T3OWGyEl5FpZw1QI4yzQ
0GljW64f2uusRMMwuT2A/++L7f+HDsVdUdL1gf/2avlVAFReoDkSU+SZbRR1+VTDpXy1XChukruz
48KE1ekISYavDZXLl03eEKYGThoj3kBNda3KKQxS5kq1XhgLKMkHXON66ETyOAzt4CpKhM0qok/n
RBGbdUmIU4o6NLuXFk0rrxZUj2652X62/9W0wbPCE1Nl6OH4X7QfyecNPP0Ijy2QvZiLRX6yW7MF
6VjoaEqStaIy8VmLlatrxMtn5dXvXoUvWV7cjwprVggz528ML/QFCXfjSABYN0bGT/nc0dBFMFC2
vZOH7csLyF9QU/qC4i0IzqF9ZAomJ8KtibWeFkgOaQ6APu2VfUBzs4XxPsTps3m1ZiUya4+vDUIQ
LfMFEgdR2JFEJr3yJs21uYuTo0LHHZgU4mBI6erFXVnlUtp1sKA+Av/mOObeSmELQ6uFfjRv6Pk1
Ph+10Zol1s77maxyRH2Ul62kCPz3DIWNEtgL3PUVsPrGCcFsWHyro3jBBWoWNU84yzNcelshsBdz
7RmnyKEr4SZK8mpQCTXIjdG6/QawQiNbc0YDim+O7Bn8BxgiTJ8b4Z8OrIu2Ozcyzi3DoqkDttzy
rwXTfJOTQjioonsVHGHWX5miAJgtgFuuagGDF97zqhRbp5NC3QcipveaGOhpWeMSvz3tea0UB7HW
B4r+jmSJkkJl7VgspQFrfglymkAhBCj/eWjxgXxpqcUB52mW68KIIOitc6uJ8u6sB1QskeS+HbOI
xaB4iuGREVRG/P25lIq1tsPg9sohmouK+nm/1r97DI3ar/W7txBKNyooaT95Muu94IFg7PmyFy/4
8VqnBw+R7ZXkMBUeJFGxpQ+B4KVSl/eIBZIEDrd+FtLgEtarGlO5GLrUlJRlWQpioPQMaUpAg8sb
op6+GKQlskJpx+wFmrD0oLdvfdPIEi2Fnl9ErJQsNuMjAwG4z1WVfpChd+mmKUIpGsSuuqGkRTjO
QitOfP2xhaMqrko6f7eV6m9xsKtf32BmNumyuJ7UIZpI7xXW2uMgCAii8aKZAQi/GELG3Q/ve66X
I/TmHefuaQXRjDdx2k89+jWGw8iJ5YPA8RnJAPLEzG6j7NxgYUtqT7NlUP7DGH0MyJQcSNlnShLU
lkfA8gb6BGpudKT42+n67SXiC3g88iTLt6sNWh675gA/vA2VwALgKe0wvlg7hvOkPLZG6ssIi8fZ
dcYK4nykmqI9OhVlMw3Cdr1x4FBxaf0Nbz3azKANDuuXSUIYRwYB37XL4KZqt2DBTPNwRNVGBOFm
dH9EL7SiQ8s1x20deENls216FHdxYUizKaoVHPIScAzRIaTxWfuPktl3LttFaxmgg+PFI2a0oplY
Owkmvs1bMddfK80oUJ9cTH7t6m8HsBKuXB2XbVRGDCoFwrSM7DJ29JhFlt4HEy+N7PYx4Xqh6SER
vnDHoqve2QK6arTmYtal3oTof87XFUXa2B9YUXA9PvGkX0f6lw9L6u/rL9omP/mDaS32ql0k5ZiW
LmnlNaYr0oHk5e1ZqMUMM7ObKBKeJSCm5MoENGW3SVvvB3LCh3X2e+eIl8NEIfRXufjJGXVVg+D9
9QVAz9zC22t95cj6Oo2LMv8McczGJyQm+Bs7WiZZw7lNIrtcM2FB7oRBcOs+1Wf7Lo4ubBU2j6ha
IvmZdkxxAFYGtDRyt19Lq4zG7KxMIKXwk9f6TszV13W5zTV+00SPdPyullDN1gAOMQeeS8VfzwtJ
fvxUfRC4P7DtgzCWyYKf3IVEqspszbRhRK/u3C3MwJCnl/WmahdUZBXVovFWDSIH2qGQ/vdhrSRm
GdWWpB6Ut2V0ILxpn7jOGiGrLinx9mbz8LeefDlADiH1DNplqlYKMrdX+K8svB2wcU4DNmt1b3NY
mt25iKAtDR5M2LsBa8ARLyrdzZtuNEOf21FJtkv/0tfermr++FeEWGzwDatycVaQ+shgdNLBhwQu
viVYuu6CkY8JnNMlR2XrEhsU6eZlk8EQC2NUUixbQqNOMyvbTROvvX4yiVMiJMFOEh5aAwsik5bx
3w4NgCesLPSYpJZAf202fJeE9ixdPk09Yrs1B2MXuIouCywP4Ju27QEp1zrLapLF5HZQC4w3M47A
wZZ3Sc97lW/WFJ6jpB0KEuhXfKJGk5KMqhJJcUS21KT3e9MFswGeMunwysg2OojzFQpQHgY2X5l8
jnZD/GsYoD77/fnkt6pl0xOpFXKlB5jiauD68pybDnmf1qrcaUXMCGXtf5Q1O0kaefyFFCNSq5SK
ymnLIUW5XXgnQ1fq8YET2OG4uKWdMvntx70E6VyY7CEmiURdqC5//MOx6AHK6vWMT/UScVPNARYp
kBZqTyEfe7YdQYGmnWaZD3yaf0r/gbmQbeTlRc4BLqp+42xk6YE4p5f+/rWw+sIume2+8KqzObWo
W8iCUgXovS9DU/N1EcM9hc+PYWCe6TIKHU8V6jSndxKXcNCCRtDCorcebBDOn3TsqfpwLUyZj8Yg
i4QVguJE+SIuoFMcIIadjeIKd5ZBa3Z83UExB0xeZK7XnE4p4vAtV+U3CLJJURh6Wfj6/DBWOqv6
IivrcVMJoi3OH43QDrfI/kDYsJpV9BM44NNGLZq0hUnhHFzuQfeO2lGVwXOoxA1SH9j+df32JlX1
Z+jt7iPAqFwxz0WbgrgawVo2vQBSWS/GliLLtvQRxypfhVbXntgyAoaAAEgTqcFPYMNehjthipnx
uqiZcc9sizCVsID2Mtn6loRsnmbzlfjVwehy8KXguEomc91JIqx81AA1fC/JTabiFidhqqF1zm3J
4rePwN1UpI80X+Cz6t4R2FoWfkR2AIyjua5HzXlzW1rKkvZnRQ+pDERe5P3uvv2aJF/Obt6XUZqE
95guiLZNXv9zGnrQpmVxB3+vJfUNXBRi8/fl5ip2Zn1InjgCu1QLsnBNgWef+IEH7UyKZElCqqNL
0IxWHycZxSpk+D5gqVPDP9ksmzJh+Mvdrm1OyML1Rs4yFo7P2bi1sZ5oLE46XDrLyQtGrYoyHqdv
+jv46uSpFLajo4kPuaTORQNL7zfP6kIJClUVSLEJs9rm5Dj7JLTw271OaEBdxpY/ZLKHgrZlvBSV
6I1q0GJfQyfUni+k3fYVIxrSNskc42HX8NfX1sD93X51Era1yVXsw3puGVfnBE5ZQNNww+y+V/em
9SlgKcRYsAXFheYHXkT7+p1lRa7MZhC2FcclQ3Xt03znYk4YDkqiyg346jaZ4Bi9EaCTJXOroSyK
v8Bi+jFY/cdTjFsb+Qf8qjrrF9kppIckDIbSwqbi9vnGGgwrN1flWuoCrtaiEw7+upM58phGhVsw
DAd2zMbM1BkursvYcz2y3OEFKhm3AIbuPrTXmBMpqJkob7lpG3eKtfkUEakRAr7SgzNHl/aviIsa
CZuQVFYIQZhKG7w+dNZPEpgd2z7beOU/LAGRf9YiI/RcfbXGMJ4bJhOG/EnWklRWTvX2hlg02cOB
RdGN5UJxo9USGPthxbX15wobR1BXkCj5/icgbxHEDqXL6z+Zz8aX3WW4BjSh6aawhHKQLXBhll3r
iv0WakGJSSesSY1s4/F/y6ik/7LCd2vf8cooYufJC0pNJp+2G6iw6CNqDFDCchgJhnNWuzKQvlFy
qWTPPpDnv7mh1j/SHo1G9P2PhMdmXNGjymXziKDyIxehzmjdIv1jC4eEnz4sjOlyFP1BczsuVyd+
m5UzJ442rLG4ClV9z+sygRSYdhPTfP/A3BzLkTVYq4MWC1ZWkp93AyDS2B1WupFKWOECercXdEGn
P+aRuRhtQHJFgoJGubrhSnShpjj7XLV6EfMmtFsFz0thBIzYWEmFPhxiJIvS+BpXzhyEK3vNS5Jk
2knjC9mkXYakRv97nQqUqfSTThP/VNqPLNjaUBXvw5z9POG4trvjFZJ9liiO9fbUraHpD2hxjNaM
mSAVEPncevTiT9BBTO2oN6P3nkQtQ1068uocSCFXyS8/jLHtcCYSY/9lJHTwg2MCbU4ILXvD65Lb
mKtPD1f7FZgpzIsj+GphyXHDdPI5O/KU8l4yS1oHddjzJNi1Yj9LXp40kbrOTKMUWxQ3fShYlOh0
LBvgdlu5l/Qf8udIkT8kfe5QcGCvhDTGWWQEVppw3W6LFyf8y5nR6mjralDULsGXNsNmkgDxZt/p
JUlxap1WPqLtZu/WJ3szX1UHxLCh3fwzNqKroCoulY0zDFOOdGxYQilWVKCePL+RqfiYTRfUFpKi
B3PB1WPXGCTcDABus2rV5mBhYKBqhHFJkwf95Jb+8ar2yxivcUiqFIfaMFZNm5h7AxiQdEiYJMxP
NVXlfeGory3Uo8BYYfpFG0JJ+BJvIHEsdHzKOsJcO/Ja+jaLA95zYxR5F+zjVKbpSKFzunaxrn4Y
JSyhQ/PrtRKwgogyDOwqQXRvO6Rf/2bsigms68r4QQ7j0Eyd3V//OUzZLoSCfK3VFdQHcq31oCav
Fg52ihJq1YWtIzEFgwGclvhdjA/TZaqpGL4FTKv8OAsOht7h/zbZYgDKXt90ICzeeIsBbE0GoEnd
MSwUAx/+/OexoL3fGV4vYDpZwTMUw9BIiDScplO0CCHQe3FX9SmyxngDjviHOfrQvq9z00I482Oi
/RNOSic4lTHc/SgMPxdbzQoSMDnIiFANGM9JniQ9nGfa94PHQ4Shv9diCN9sN0zzIyXjV06vxiOi
rk8qT9XwVKnDRFdm0l+Xc5IgRHOrGTCNyhgdAGd1hLFTGc4CKWP/4OmVSqiHZas8ByUlw+d+aILe
8DRbrval9EeMLCAsxTO4MXiohjA17jTnTOa80WbHARFDTJyQ6afriBC7uTDVxcAE135Ok8fSJLMh
m+g00pYt693oBylE0UnyoAZqRP23fIv0ecQVUzE5+b8+ZSsZXm2aXsXadNGs7H5KN79WJiwdJ0Zz
trmdB5/FIL5DU9mn3pDwpL/ODxuZ6FDRI03bvdrqDSbqrAMAo+cW4lAEcF3aPv1Ro+iwkqkZO9wj
jTytcmyqHvAC2HxYVnT5OvsT3xhMzISPDKBwQYbQOtyE3R4cZPlnLV4Dem9Ewmk9FZikOx/xcV6q
6gJSJtyUuvpfCtn2Vb+/qRdjkMA4t7lM1iTj3GEbMuf8oObgD9qFsabDZDxO+Th5JyIpcod49VFq
hilUrTO7JIyMWMzg1PRkmeYSd1e9OKBxc0X7wAF7XQaWvwKAsDx0FBcZ4C0QvP4sAKgN9HmwZvRD
W7EpH7sXK9ehB6d9oCg6GKG0WnrgOwzxqDv/c7TNqt0ST5LNDiAA2n8uwLbaLSybFmLWXprkss07
CZBAu30XsoXgZi3LMIiCxHHXyiojyMl7EwYG1h/m5xzs2Lj9riAqrBynndJ/e49AK6R8pHRb3BAZ
r5K5uV/iaX2EARbpGnbuYGSuAHi39OxmYbmzpW+2AQ6oSumGOs2StF9xdqU9nlqt14pspIQstlJR
pbrgZy8G+vHYez9gl/YAO5aH2pYjLSpBlmkOWKxGuZGL+B0mRBwifv2zOhC2ulKy6prPfrZcz/F7
BHpgLWUEJ4C89YqMD7r0WYzkX3P/gMXMXjhp45wbSQGErIwfu7JRcTqpbNxBPkUSbRUQ3855XIiL
wFncGk4j9t/pqITTC02PHdDvOkAAkbFUEGWbVAjq5+1Nu6bDKAKS54OtGMELJFPaSIICr/fHcje9
J/EGvFLOjQPg8urFMP6ATIGeGIFKHZD/eRcbGU4qWg3quU4iCIaj1iYp9sJasbMcRfPQ6DIZFtpe
JB+cV7dIOq98XGswNXk1xZUp+bsKKbhZGc6XS08A6gN9sIduI6ce7f5BWPab7U6HrCH5r1FTKofA
pfH+ze0Zj23gubty991nqCVOuflS1V/wmee7TlXcG/2DlSrZoY1hbu7Z5WV7YZYKJOng67M38w4D
/RADr6Gv25m1XtRSX1o9RY4CBRA74AERBD6QzY5ppWzMJqRcZOwdckt9WfQiROFbWOgiWv5HZCt/
zAIY5jmUbckPrEvQ4AmhzBM6i8QVPsP/wWDRr5NMVaYVH7bNaw18gJNTy67Qgka2exyy+h06UzF6
JQj3RGmL9yMUMJ7ve74GHeRYIcW8FoZ4j29DAs1GaJIkeZm+CUcxeX36oJ6WijvfQoF93AXerNFE
GCpCM3LTU/m6sVN6l/5brOR4zcjFX/5I75cAsFI/Z0QTnLt4n1PmXk/tiqn2PMIWs0F18OsT18HS
kuh30HCJe8hkY/KKrBU2eurZrbN2YwJkLTDdL3sXm6nPAfmbtRlKhgnjjH3gVOuyLkLvhfKaQ4qr
1daiM4gLEC4vtpvMxFaGKEQK9AJFSoTKOw+CF6fAoDfAsA1YJD6+zZ0I4TwJV1YUPoyMp7Fop9XO
GecaqYCMppctOUjBNf5q5s1n0/Z/WNEuTznJVzQBdW1haZjvg5TZ+rGL8JApWZVz3zf8t9BfRWZL
v72heKncYYXracvYLUT7Fb5XD9Rny6uT3Aso46nEICO/pzUCi2V54u1cuDgmLuU959qk7vI/mnrI
sQv0MOJGF4fv3owWmGMcVgqH7Z7M3SheamkSz904Ytuxno6hUgE42DOo8XguIwpz/E1rpJG+GfpQ
F+LgZrE6GsgJlEGfKQJf7Iw4PZl/CoUJTAOd4PaXeHfNjFfaSMoWmhx2/i3BFX5TTTeVv0CbEIK/
6GvVTXkMCSM4Gp8xhIE8bihT2OWdR55LANCwkw7SkIhM6QQ/wtqu034ZVf1YD+5SujYQzMBMtZli
quyCbwEO0xIvLCatrQOIN0Fr+omRBOjJ59xHZhS4TlQpPfJXEpsbevyDkG3ZqH9TyaKAIlRy2Ct1
ylzVt8RL5ry8eFum65STjWRHu/7SOGKUWBqWCcB9aQRCVjBMJvK1mTwsp9w/v9NnJx0c5yKv1ZXM
R8MHfq+lNzDBwRx9sFXHMCc9Onh5jORO27kBNeXYriPT8m9XDubuOSy3ZvaP9+HZS8sJmBWuy0nc
OS1+IuyTlOJtZlAEoe32tk6Ff/mx9PmlmXFIOylFylUtKdr9yAvCjNPMW8g/kSchGf6xFz//tnbU
pT+F3wb65E43JQX6LQafzm9Y4SG+6fWzPi+LSbTWa7xD0gPGP324iMEpbtaXgEaes97XDVIe887s
tFVbWBkjOp/xSByrTVcOfLTuThOU/LOepz2AoRIdx1uzBwG+1NUzWaF+MknpaLWxOQVQPUtaTm9D
NZCjsIEE0eH+QxVcx7C8JX3AZUpMRTwk5nC+9thxbnVu+U7tt+aHdvRijZLhOHPsBmesGatOmsGg
ON/XCZKkB3VdcXSM1Ia+4K1O56DadZdciEOhEXjclk9RXvbLdYTu2f9+drf7shUh/xQmRu9nidge
5Z+hjoRE/4ZeiY910sHMx5Yf+9fVjFP0tH1MqSr7vZrK1TBs+9ac5Zaovl0BvPuAEpKIManmA9ib
0ahS1gRv9FHwuH95/Vrq8+IHQPlsf8VDi1gd+SZt3qklNfQjDMk/fnTNT42rvt6FLlGOvSMrItC3
4obT1Q7YmXMJ5GWc70/nLgVstrsyq6rc4S7+PLsyuab5XJn3nEQnqXaYHkSnLcwxXdI4CkUNh0LE
dqgLXBAnXDCJ09oGvt4VzND/aG2YJTWiqppT2OFErG22MEAc8wP270Js86HOjt2Fg6s3Gce2HN3m
rFeUhhfBSc43pwmETpHyqtJfk3S4owzgUO82kZW02Md306fG4IqtkuAAcV4C5NBc6F1c1y58GwDG
mMaQ3nphErWJVlL0Ukozh7zir/zNS/9KUiFdCzU87Bdf19O/VLvBid/in6lWd9uX2ovFjVlnu3QM
5ci13EIu/7QEMLN10e7RKeg7geHHt3bs53qNWyzX3FW+bJs4YZ5lV84nAFwnqYs92Uz/kXaqVmP/
VLnXEpdZo4bfs9IWzE0ewXAO03p4dEe5Q1Khvm+cvxJOgw+RkYFY0RQ4/UN9Rut6sBgBXVOOiqDn
gVI47DVPQHt09lYOXZj3yPq23q/m2S1WCazcT9JvT6wBRbJhJ0lBCVj0q9Km/OctJgil3d14dZT6
UVtnHkQZL45ke2m3FGAJrX7EZoTqvQdO5OzG0HO6atBtcu0xFEfoALMDlgf7xxi1Bm+aFemiQDzR
jpWk2jGhBZsSfXDLaC7xA12zVjGSlVi1PbYRpp0JNApAaNZthljUsx4dlwiWvz0Zh2aC7mnQz6YT
4Bt85YVdZpYBv1JEXa6NaaUhcQR0U34frdkkjjXJePfgeOAHi2RZuwzSE8j0/jREKRR7596pth/f
DOkhPKjld6OlYXFyZKuMPz6CAIZed2u+itJQnD9escSsHzUGywHqMAI9CyhYEwkKYqq+LAqnXdqz
aXc27YqKq+6e1v+d9Hy9FW+SMHfUgzedLN0idwSUZfwXlP+QFxnXU48xBLBsz5DKZyTmgw1G1Ktv
gflTUGgVVZiM99vJbPCyVKKnCaQM2TzsTUac40kI1eUMsWt6bXbut9551lG6HXPlAIIWWAUpMkps
c8V9kfze0xKyVwhNKM/SkSl1VhQezqx6FsMeaWcDgjYTmysusSPDLYymWLZa86r2jbsbBdvnEK11
lhbKI/Ft71WBPBq8K8TIK6eoPnGZTbHXjVuP6A7mM395sKOJV+YPW1igx9Jh9vfNhWtgSCJZLlGU
lchf61Ax/X53ExNc4wNiU1IAzrr6uYb0AGkzm+TST0a3KdOcQ3KU32yMBLseHWOc/bRRo9jyPH5L
HVYRNcVedn46MO5cadqmFq9Pbj8Puk9Bls1E7oYA3gpWyRJ4DuWgj606F6v/e5O0O4brITi3fce4
+54zlSBP83rTZl9nNtXoka7xnJfX7czz9ejCBNx069Mn1p2h7HD0zU8gjP5GylJVeryLYtYjpsk4
+NJAvOsCM0pKCPqgdEC8xtTd1wBXKsPSMfng4vP2dtXq8xPpSpyet9rQ+Aai3N0F5+x5NO08Zjz6
7YhNlQMtRMSqM4P+eeXSvb6/5lIZP65AIouuiUAuoZpTdbClS8EFOUld+lKrhfZMuEAIzGVFUVzg
MUuGPpKFKAhjcIhvEFVqEo2Igd6FKDP9xMopfeCre7UfsIVcV80N2OgXTvRUdf5SFp9FhL81MMgm
+Bu45UGWDqPhQ8SpaLgcmNd47Lh+q8rzTpid12P71/Bv6fDA4A3zrihb3aoYpDH/woVYyl+xnHob
sBwvPnsdvosG+DDAtQ5j/YCcpLeTJCLDUnYCG1hikeA8Uv8na5XdDTtFTpbmwTr8ZXavu306GMyJ
3uhZaWLOuzmNGrcDO2Gz6RyhACLIG5tClwFCjN4iVdFyla+yobezeoAmYmoKuzmc5ufmno5dvnBs
ooXVwAF3FgU3+OtLDNpBn6Mwx7XbAuZOJwvCV593k9NdebY9EsHM+0ujZ+e/xZqRiY1+hkaVYQJz
qfaiQmdDqfoCh1Bw0ogtAblqbTVkQ9iknyjm3tPtYjQ56hnv5SIxP/I8xdZy58yJSPnhDb9FGKTZ
3YW9FfJtM2QQQ1gcAr6qz0DvYo9C2k0Zeb8IH+VeT5KD3qphE193404xwwT9C5uk0w06//+O83M5
JPpZ9lzAJlpgd9AZ/57bDt4PdO36JTVtqJrqOJTvNBU9wEfmiT+OdaWebLjrXv8IanVDWq7ScscL
Wz+6GNxPCuj+oy8/2AzxftvEofjTEGnv8hO6jnAAK4dq/NlBP6uNjf+jylF3qJWpeqrmjiQOidj5
aFaZivJWWovjVDUsrGnAGG5qRRCRMy5xSVmDFeCoE3xG8EdRNlq/GCLYNokQiOOUf9pIn7jW8Vmb
+uXKBr/q9I2WRlfvur5MRV7iHoemXyx7TUrBDhdpPyLC3Rc3JRpfog0IIsMMNOajr3Hgj5chY/S4
uR8Tmbh4tuY1DzIHM4WNi7nQu6URmgBjjFqs5NKul1f+7Y42+rroyxHsbKmyKZ8VWLTCr2BSOGZZ
u/8Eob7BLvyQBLm2fvlGiQx5Zjia7O6kruOyoy5CVDt0bR31DykvXb+Sm0N7IICHysKnkRFdA8fq
2nYdMWw4uJUq36Zv95xxBIQkPkNu+dFMLVi1cscj9kzUXq4jcwKSrI+8OR5wJPH+l6+pLTdqwlGK
mapnXvDvlV9VswMI2A2Js0tc/QYkW56TXUPBQY/9r5X+9eStRpG1sFIrm7BEAXTkKJPBDJftuMr8
tIIurM+Dj+ComVbawcSgS1GEAJ25xnpuAvVTItZU3QFW4/owqv1Smi4uX8UDJR78rONJWaKkAOTy
HAs7iNC0sRc7PhPifVHfSIt8oDqL+HiX8hOXPTmD/lbiofJZ2Pwbf/q4stm8CsTy4ahxbXuNYs3B
yGuDlY+DB1I7fHZqFmthSYeFdR8A+YgDQ7nOAdqDN+HjNlFU8YtBy7FBI2xDGC3PJ1OpDkxyTX+J
pYW0KdCh1edKNykqZ3Pw9h+fJJmmPpIv4eTFwdcynh1z2DfysVDE6awI7SCy8+RtWndQ7kTHU4v9
5HZzSCOWMj2P6QKdFo/6e8r/z9OHzl+30+Itjoz8JFbxvNWlyAafEvQAscSm9e1/2rJg0s1T57QL
pxoygm6NnQJ+5dGrUTNeLiJHegOzeCx5x0PTiEdTlaGRQuKYNLklSxCI+4UBBpHjKq6alHJcKUy5
OPoLZzswSC4EK7Hlo5hiAEK7OKpQC6e3h8HudFkQTgOGroKO864/2uRoyywI0WNnJwv3McaUZA/I
5bXPDDFfBoz/R6V2Bi2JrsMtKI6JJ9CuOCaDQIP9FEZyVqJKdrZf8YymUhSkROsNw41bz6dgwXyk
ATZ8v8cQecvSgj4rxzQs2yUlh0mQdpbZmdIxjeWeeAxE18K3UnnLI30YBTdJVNriDPWev7+zYsOe
oNnpZ57tVQBrZGngf50NuUROBxMvO9gohszROxB4Q2pJ6UHZIexqIPC6Xsei1HPcq17cpcJuwnxO
+zzkVEyitQplLtgxDdybPFiJp1rJSirsG+AQAGzc6u5Ud+hNltBfwfEHM2H6xoowbz33WK11u83u
F6NWfOdvIcZoXAKD1duGZtOXkUCOZ4cFLCKV7/lfiGnxJNYzOatLBTOvD8AI4jaG9IASjKBAbuzM
jRw68iFR3VRikUl7X82jA/Vg/GFMeScRWXB1VgO478MsRfGiAt9Q7ID80UnEm1LyjkeOiR3csQcK
CjlFG6CL2KyI4MGiqSkp7Xh/pQXdB0plvhDrnepgzsLFhQ3eORPdXkH2Qh+S4euSvf9s/aUwllC7
BsFdOrttZRpKj/WVM2jzk7h13Brrlw1+YaZPGkp1DiIuzETU87sxiO9Ca8nKlzOPMSt+dlGBr5em
LHUji22466kde38pJ+8HssPfeQrvanVjyrHW275Y5tjQjX0W43ZjudLCSJmZndbA/z7NxxOpSywf
JmKod8n7ZJEfahrcQe16VTy4G8Uu63tD/gVqSxyIWdT4SbHLUx84s1SAN6wQN3Yb97Q9pjKFudNW
zRckukLXeaNMvqYQJiAyNGLThdx2gZrLuqdyZkh38AKyli989N3s8GHg735Ctum/Gg+tzMmKBY3/
fLx8HqI8JkjdKjwmxAvizXSoQcOGiR4HYr7CsaQW4NmDfs8/2faAZxneIr/Ke6aGUMed2nBtNZhx
E9KduatipSb0FKzG592tohoTnvdpA3wHpv75DmlQU3cf6ZJdMN/oZo53wUZsJN65q7IlSVwUx9Yt
uk3J8/5KKnRpbVdfIFFA38yquzHV/H2042wPJ2gV/vDP9kIGSyy9s40nKPTfDsuYkbFas3D96Iov
YUgT4dmC1BlLzyn1aDXdVSrrZEKwRVN7RkPHlLafpexbGikbhu10a66Qnx9aYVGX7D+I+5lrkgti
DHez+4MAnhCk/bQ/lbSuUuhrb1fRHM6FWJvTs54rWRwky9I9F1l+bIvYLdLnKacnhsyDNKAKxa/w
8YzyKHbrryQelLTB89cxTo2igpD7+z6ZXSJMhlsmQpYF9JfIYHD56cbPWaJoqbcw2/u/tJKI5MuV
fUPD9HRwYIM6xWap1iCHXZMIuHcfI6yYdUabFTT9HTnPp7xRmQOCLLysJpQd6bw4P/JFatO0h9YY
NPJZr22ssNnvC5QuLhreJXsuwqd3YSfFQzgOeDr/UgKaXRuNeyeOahAy7UeFWwk8KSpaQ8QbOHiS
tkslPKVye0LngES8TFyi9TQ5g/Xr4m/3hqI3YRrIbW+W8V4rnCsbLQk3ZQzYLASAIL2cqKixwhuV
R9ShK4g9BEEYX29rf/IdKb+Iic3oZM2PRsrNc0YSndPnu4zDsm3LGbfEGCExrqKgJcAxXQSvqrNj
ofiI4Dlkxjt71GulYIDHC727flyx4LCROf9mwSMz7nmfoYILY+C8KJEBm1Ay7ls5WGo/WQSqEuLz
2QEeGa2RED1bw+6LDG2Eabe4NZYPkUTIjsPPHOZHhDgJpmfkudlQnN1txNNcrkjVF4PC5A71QgIw
4chJifpfI72Xk8cKgwtnrudEJFGwPdi4GwnvE6fGGHgQ3k8T/QQZyt6LbTyOjExTLDVdJWitizr5
2HyAar3YjlpYz2XM2+XXWINqxpTLeCoyIzKb4rvQD1iKnVdEG7OS2+CFbvkzoA21r1bHyutTXogA
FW7HEiq9WEpelO8jpCX6cV+o4+GkcPxdFBscgN+5ZzAE5n4ARa0PjdS0vmtL2QO9dc0Nl8sqZOXY
RTdzZc4qguPkNlP4N+q+XnS92YVroQvP951xKmm3rx1y1WsyEDx6F2rVFgirAEj3aTHuUXL0Gxu0
tCoXlh4vKL3w8z3imRy/R3EVDW4n0qAkw1LYb6RKRfj+gdpWCiVLe5Aod0U2LOaw9/02Ue80W9Ct
dYpTUlfBykZNxMbvQDM1JcibMa8i/IDm7KSbz4dJHqaFDy+PLtDZ2Bfa/n4mqQHCTa2XNw94E91t
m/pERZuN5KAlw6L+jYNjZtonprkLVweX7O1D0LuNDlfrmv5OGu3oldMrkXHCnXjTMol8Fq8h+niT
83q6zKzrCweAsz8mUbuDBeA/wjimIFJNXHGuDSRKx7StB4Aw0rQfLQME8QdQw6iatTMNLQBVKjdi
a3LztpGJI44MwzmzrDx8eAK7RfUpFU2jeNXBSohYXn44ojl/gR9G+bmM1UXAElM9HyNV73pIJ+/Y
qu7Oah4FwO6zvTGz5ghjbLghGJhL8+ewBmVnGExUBqv6Lz1TLY9i7j4tq0OJE9DGYtSR0JiyAOuP
xUNMr5RGEsPmZH1bwHnt+wV/1fODKZpa2mur0SFUYLGHhyLGe7lauLRaGIKczW6GbGrjbcTHR3mH
c9mVYjgj9wTyEI4c1C2J4aHo7GcON8Z1KzOGpc3JYOqsPQETVABB3zWcEKi3u/orag0lWbYUfKer
y1iqrMruYdi18ISgqj1Jk+ndiHWlaEozvz9SBc9iTn06y8kpFP4DEnfSyGobKv3KR6j6bsTRkhI6
hXA3RC69SON2cHeTUGocUd2TYCWOIpd5prIeXXGb2QkWbU5wg1HuxIOzJx6p1IMw1YBrnOluwNVa
0UR24efjp4AnrRJiyMHCmhA1O/onUEfxnMJCtAM3Hks52fQ0vJkYj+bxxH5Sh2GDcZmd6MthqRhS
emurTE27G0OXheW27TCZAdSkRmXmaQJdbVQkt17mBY9Cq11xW5iA6u77LmhzNyCH2fNzSqkQKsaE
VbnXgQ5qs3RaQt3UH0rlNgjy9NVmcMtcHZ1dI0n5vJKDPq/Wu7DzCSLzElWXs4FZ5xBN8qEM+ReL
Yu3z8VGbTA84orw/74vO5DeONOtYZcEq7nxZv8nP004uUYpH+Pwkq2t8voMb4z4tS6NUaxWKE+Ps
J3kAnJPR7VUyVquNrhDhVtQd/rkmS2GUNnZHSPi+eShTaXvp0J19n26u0sbQ3z8YFmanCdj+uTdP
tSw1Cp29pl5zv6nLk8ZSkg9FopivL/Q4lrV2yg5oz9kq3D0UezX43XvsQL6RlAF74jnw51f4BMLU
cL+WD6kOOTdM4w2ORZId6t2EkaL0EVrWSyw2GK7Qsy+EY3rSWxd+fXYtkjXOAo9/S1K5pLv4/WCZ
mnRAp/a+pFBFO6GPpZApTiHxVmX1gk5Mvq1YBMHYQselpDLAGktKUFj50WACx9Xe9qjathYMbGkk
uSnzzRsDFyAErl7BeFXVbRAeOE89BuuC4Se3Zxo8slh34UNcCU+HhjB1tZDzalgvQHE7FzuWPx9W
u8QU68R2OhZjdiHk1IXKP3LxYRPrL1fDNNRtPik/9bELfFrwQofgxwN4dwq+imJyyfNine9rQ6zy
yMAlNlj9DLq+utUmf5yGazJ2RsCTH0gN+DAfrqs5uKQYgd7pOQ5Bx+f78oPXdS7Z16ddlhfKlrzJ
MMXNw4VbPnov18ocewJwTbdmSDQyt3NjrcZ/wiANHwCu4IhhRUPw9T5ptoJk+8ZeAoNi2Ws+9/AN
OO6pi+5s06pVHzfLkdAZvD7/PtiPKHxvUAMGYULmCQAcclKai/tmJFWWJ5xBbSzkRTvu1MRm51oo
LuluQ9Ns25zFTaIqF6yEpNa7ES50al0xXtXVbMBpsBmnSRAC1cz3EKwEDKaKGw1B0H/68kfI+YJ0
1o0wHFI2ZikA1qyTMVxMdGtmijObQJPszz7dvKOoWrS3SOw8d2zJuxz2qSEUxK6nkSI7hS+rP+mo
e3Ir/Zngwhtq+T610wYn3GJ1lCss5CiYmqhFdPq1WTEbsuwP3B+IBcnBa0djGjXzoLW3Eg3/cnCw
JIiN/Lo/IyhSIspFlHDuZtbSb8guGj6XMdIAR97qfouj5/IJoGx+heIj3CTb16PSE7DqYG0L40Rt
ywqfJ1Zy+ENJ/mVETG05kbRrOI3Xyfq14iFA2hDHJGtIwK6WQEOrbTQRucUQeuK+LZKREu17wJ/B
5m6QhrOPZktv3f/AILlPXQ0S62US0yEzU8yiSvxcjtWKE0otEoACqKo1oQFrYxe+kSeHTtN6fptl
ZlVzAHHOvv8eQWiwuR41xzv2fzw0cfayrt89ecYRvn/649Ij3Q1UvaWREYET2ji7lTmsOetwe6Y2
9wE7hwos0dWOin3H/8mIitWNXccm+f4LS/C+trCYttPcuaaIOSJ8K9TozA3eOgUM+zxl12S/EvUx
NLdrF0Dg7QtcD1gt4kGBK5MFJbxX3RozfTy9uarAZbla+OFsoXNz4Kw+V9GNXf//ysplwpkCRSpv
TWtFYSeTJ/KB2y4eTkiw+tqM8qR9XGnGDGJj/0qG4N40M8jbxMxnvxcKfnHbaLjiS9OfGgBXBAlF
X6usCUlvKsBCyccJIDJ4tysp/oiYw4do8VKyWHM1Wuhtd4f9kNV9R4uJNmj5zAj4rUgxpyEKFTVw
oWdEhUMv2v0KyPTef2yUbBpvP/QtGoj0cVZdzZAMrjEgpW2FkIujaY1jA0wg5cj3DA3C9rSu4beJ
UWsYG+jwhEL8i8RI/wnzhJJb0LNEzjhjtfp5aixmSfTZ2U+ZSrnIX7rmqJMKFMFNstktOwLlLx+9
F9LVWiKXTqVwiqxTJYEDPa6EzYSM4SfYJEKBQRs6RI0l6Z4lHISaGPhv9qh11n+YrVY3/k7cecqz
IfUyeW1vRVu0c6Grdkkaf9bxQB9dXX2V7KSKnWYRUiks1yNw51w0ouPEz+1E1YOxhV8W2+dFJlnT
RqfnelhdkYcjHlYllpxJXxGLkHgqY2R9BY+KvM1ox4RRGYt46dAxRAiG0TdpBIog0oos+kmLYO4/
QBznPaPxFDcwH4wbPtvQn3TIjbVJQyyvV6HH7JV+qX15oY3HYXY5vD85gdQo+h6c3xcNKfaEz+Eg
4QSVdkzsDJOfuMX1OlKUcHy4HKcWgZVj0J12p6lo8DM++eE9+VU7xu1EYJlOQxhPhaqUWO/LtgnG
E/JuEBuPalnBbrgr2cgm5r8VsbsyO4o+bPkN+LHCIH7zuMqVXKYXm0i6yVqdBpZjm0lL2dhHSZej
uT4zoH0Wx7g8MAqT0wxtgH7mu8AlOyeqw/21/DCrSNihUzqPVuwmC4jbhsBzIBjOHZHczRXbR8cW
/V3wJfkt/oKnetk2/a31DM9Ic/yPdsGVX9m0RX0zb2THq37C8M0bemjvngVKTu0LninrrilYQ/OG
TheBFBdUK+56CY6ZZOtlgiKFzhi+8F0qd1iPuNKtIUUang44T4ndvRpVkfKn7TgcK0igZs80T4RU
JZzuz2jDgzgekyDqPxLUmt7oznZZv3coidWgQjktaluzABikV/WjE7WSqdCMXYkynCEiBuV6V6kB
1O0NxcphJpLNOPBJuZSutg5TFVTdmWEZMV9WJcPecODjNIIKijq7pSP2Mj4i/u7wGUhgSsUJ6ya8
KJX29MjMzpD284HnS68lBKDmHrnMd5KBoiFOMtht70rMiF8CMwWtChT9ASSxlmBmTogQdaJS2Rd8
m4Cj3RuUcqAy/bQQvYKSVcEFnaZYfQz2KURF5SscV6CaMezB+CtYqctNHACNvXl9oJ4dKKdC+dRe
del5BhEx0rGBovmQHF/VF185JzfHUcvqQ+nWGO9mz1tqeJjvupfzD3ip1uQvPnWH7gLtTHoySbjo
waKAIeOCcu0Y0a9K3cuaoZaih5vnspH/Rxj3cOVxwBf09UXJKkdvmvDpoDnevh4loCOKQr1IyfOK
ZhpUYu+EKAAIEKmuwrbmnugHvbmoHQ7nXUZkMUIn2h4UcLiJ/yaXbty+b8emY4F7fOM6nJYx+LH1
lAG+1Dx9BbCtAv/FePKwQXuYH+vA6EBkiTO2lbxOrxpzX3WDN2/sGk+Mn6zalHIfoFys3uBd/0F+
URltfKNzr+vxCK7UuqI+Uh19cZ8iVsb+e5Ha3+pZVjjLsOXvXx5BSQG3vXg10zUZEbBuJ1Go6gqS
Y6AVszj3xoYGIVe/rddzfCa0wEmb8iFNBZoOisUDrLXybJzzQDz74JfUnTW5cK9FbxKxZlFES4pu
dLFg3t7HdKm3QACI15Oc86tWbXJ7jhXS65cz/wzmS480xP4bx9urfY6KWp+phbfC1mosz8q3iY+U
TWKj7EyBZFolbdlpUrDyOS33nnqNfajilvbhAN1DWMkhmGfaJe2duI71TOMJlQ0P51gnQX3hIDmp
j4/sE5f72/Bd9JHRzmaDDZMF8ci0g3eOxq3HMuCY8dP8TGXOKRtgiI1XCtrMjCLKYxvRmb3T5+TO
qk5aQjJGdzTCHv6EoI02x0A0y9Exd1D8Hl5vTEMtLTWH2/HrHPP0CaPjivaq4tm4Ia+/uN2dtCqb
V9wwqFuh5AEKMgKTZgPRjoMgW2K7zwvHp9uexATybW4454PLApqPGdRTWObDo1utqdo/I8Ph368p
bzPyxvAdzTZFcG/4H4YtXyusR2pB52xK1/jqWUPPRodrO/J9DZwfPntG8yLjI6zxoVKvZEkafUJe
vJTnnzAPVg0xUyGdG/+2SpYIOuB4QZiENxFg2yn+6FD0qf7cTALVXAXrzsP8C2veKeRzLxY1mVCE
RvbC+ZONwY0U/ZOC3mqNht/k8oCWO82jaMznCiiihZawdMNfnXeRwjCFB9q3cpsYWCDFffahCL/Q
5DLldyoHQ2pm/rVnDALpy2ELzGzAhqVOVS6ETwIiJtD98XrVxIhYqPBudUz7nj4/XCMv6A2AW9sL
Kt0PHdyp7v1FaAWx8FL98RvKeaAgViMb9BwuZ7xN0hvoZpQDLtAv3btMQ/OgvZ3QMFnbNqs+yH/o
AOn69iLhjbmSsWqgRpZb0+Kvg7IO31ivyZz3UPN6OdIdpIN7SP73evJVTEgCEjjRYQoaWKvLFrk8
wvBDUZOTWPIAdZrwtOpzATKn/zjGV25dOGuqgTBYT5ptkbbtA5Wk2xbfqD1LoNwZdDSvBl9DEwr1
Pyyuct6uI6uiKAW7pba9DcFB0fkahZLWX02fu+4a706TymwIs/VHQMPedBW/vyWqDNsrwBiCbnBI
sqtrPOTUpyzmNKMIDIymUL9oMrw6LePne5aQ+vQtf/4a+6HJXb0kGs3jh8V7GRdDNWlzwDM4qNs1
bg+JUB7Dm8ScAlmV3YZbal+I+0zslzg8mh94sy3KZMIuuJsOJsVfKRY3IrO7U5Gm9dutm/w+7dw7
xZ0C3Y+OmZON8qLWE58tRMZ60ZT0mwCyVM33lSsR5SEsyl0W3zcqkkBnuoVEwv9cGNIV0PKKsvpM
YGO02hnT1bvK0PyIj0/MmEY3KnJJy2Yuna20aO8GLdi7myJ1AKRpCCQQwM8bnJCidweElm/B+UlQ
4tmOmyh3GXql2cOU2tIzxyvz2HZhEclHDHvl1MyP6uHAyYYJj2Kdnfb7Y1u/qn2e7Ua8tLbuB58W
aIWxmVbXee+PtnSN56JNcAV8s6UeiEDEo6ZBL/z5gb245aV/btg8BnKY6Cswto34TzyO/faJ91GN
tH18I+PyQWBZbs659AKynqNYm2lNy6hOr5dlY7QqVlj5qkDzpucMcsPLkOoVyqBWAzLS2c67JoTt
Z7LM//JPEGcJQ5IFFKauN8HRLz0ow0WPFygVmqE7xy1ErULUR06LpP0yQgKT05RSy8FD4EB1SKZv
Pl7I+fo2O7EzKlVS494WBeYYd23S9mI6ZVDlt62wpKs504n2+as1IuCLMh1ZPS4+CwJg6/PVJ9+R
ZfYuM5Dpmcinzd9LDCjwvdzlGFolfuxCFMNf+mI53g3BVDcFnCXVtPNaAXnhDdgkqx0Ae1k0h2Nr
7SsB8PzE0r9+MBui8p6JAp98MbGmsGlyoKBEWDxgoXDEBoB/mb8Pk4Yxtdlettv/1aizABhsBCyD
OeQp5CxsjV78SAp39yKFtK7p/NTAX3pDh/7Ql/MuW5oYDlmKa7mkFzZ/yn7vktvXWHD9IZDXIw+e
nxrossjvc65WbBUwy2Kw7QYIW4d8poSasF0g/KnA0N5gB/WMF8MjiG/fdv7u4g/c7qi8FuMEWiTg
qB0TeCcqlskJtNSez+OSVbgGBEsJNqgPzK767RxvpaRJUCv+9oBw1wyWy1A29yQo/idoGwefF8Cj
67oOaTY1EvD7QSgYe1NKKJPpeXngDHSPj/b3sPYED4/vslntyVo+TcQ9R1xiPuTxeg3PO8bpBlM2
fbStpnpBeHatmH1DXd6e9NXs9PtENlv0l8sL3hKwujOX44witHSEZhQ7EvzOTVGJLtcLfRstyQGL
0iBJe/0AVdK+8/GTyNzvLP3qDTc68EjN4eeEZveWETMHkrBvYMV2HqI3zQeDSs8GBHDpVoPmAdDm
0bJk++bv1+vMEhnlsWEXrz990T47voPTIoGPx44y8XMbZFDsQ+YUVqTG4127ya5qdt5xfyggiYdk
fuN/ldoy02W3ZCGAbQKMNvu3wfTnidWW+bFodkuPlb5bsGmzFEpILZl7OZI9Z7U4Vz/hl2PehZIu
crUWHCoDBIepAxr1ZNivic6mGCZmz5rmNCyjU3odt8n73QH2dlc3j//zFuPjT7cNtTReTnE8hjzd
rOtljrB69CWVF/1S0rXcFfitSP34JdU/VLMppH8j95PzGNJ24lP9y+tj0Z8GDUu4dwTR7mQ8Fwpi
TaQccYM9YcT+S285OX6hztUyHFslYOhR18+gn+3o9zwvChAeGwB+oCjwDzNXqoX1uJm8wsfW5b/5
wLX3a16l9z6xjd8wUt29Rl1sVsL5ToKMaGbdhqxrqgiUQhoqOY37mLrYBjHABezEzhC/W/tFAxT0
T60vPW9kvqOJotake2+tYZQy8QssGW2QKdFg8JYCcE266RQ53bSv37dk2brCUTKz0o2pEITO/kCu
iTC0sOjspOkPQZ3X+4L9lgAHpAjE79pYoyG+WyfZlVrpw2xzwe4VyMg6Pr4ltSNLnOEXJ5NolYEB
hrdqW9/DpXa7bixL+5Swk591tIilPW+cULuB/JjE6HfuV3aiZkHXBYTEmdKoBb6rjN0yr9tajWUt
CRKOUBiMOG8Z5a3GRzToYhRJMjspB3IK1hv8YS0EDaKIHeO89I2Nj+q3iCfaOzZFhYYWwm+WJ1X4
Lw2WrhAQl3CB6IrJuFVwZrM/GUde9SSSMH7gJvG95w2ic8RN/keeWTjzjSkfAptDcvwSeHacjagQ
KGWXyH7Q3RhYVYk/yWE3iN2+iCzFp2CcdUBxPgnQGSaFzZkc70UlD6M5cEGjWhgxxbjxjmscREuW
USjBay/ExqkBqeP+M6sEXZbN1ERPklszb3TriyPLyoXt+K++F6+TaZu39zUdI516VOUmzQZIgTxU
WX/GN2+r5GTmfcmnijYPZEitv53mOeUMUzCdaNYR6tJosgbvLj6dMZ+SESO2KyBdjClnDl1WDdqR
dUAze9/OJZVzvYK875TI4UukNXCW316HFF9Iar0ucQV8SOrZuEYvjmmM/meQXuDkAbChM5U+tHym
Vqwt9RwBpVwFjmJaJtIesGyooO+jsR89lS8YDx71fSXws0JPCxHTmvJerv3RlpPXE9Yta+t7AQJ5
bzGThlPYaVbZ17/8wbrg72SH2QiBPyD1QnoqMPIMD4/i/WO4j9e58Y6jstZo/5rnMcor7s5LmERk
cOBHAKmf3eJLS+MkU6hcAwvPyuxq7Lx0oPfhl4nKIYOluWd0efYJiu/cm19zkvaW1KgqAO8ibxGn
yllIzgYHh+MlvRlzd/4MBmkgMQTl/tImXk96TeANhOvmEsYXptfSJJmQ/hx9jzoXEIjD3ZCWD3Wp
DGM0xml5RYOAGuIQMadz1lkytC4b3067VWIYapQwo1rjXQCJnE0zfKaz3SLFb1C3CplJINZMzlHO
uvnCxhRdDzbSozqx1LhYM7dy6YuyFsI/9BKnY7NllZBJU12NNMJSjuhHvSptFOCtNmDwsdeAWSqj
LbVk/0Pkmhc8gpPCZFCFtiD4Ep+BQ7QZAJc06cQTHPr+6K/4SI35gD061i/09tnUewd6fKlnl/5j
W7AhcCnnjzKxB9Wf/TAYU7zLvvAEFwlyesl8eWtFbO+qAcSx0Jhstintq6IIkO33RltS/M84FPih
4PB9XgRmIJpUd9JFHvdorlWmn78XR+FZjSDfPpl4Cfn819VEhUcsdl7n+6pFHueBZ306b879sApv
wIqs3XGGCSOYvM7IDvQaC1hUO69mJfCWrBAsq/8MuuzN9dj0JAt99NSJNEpMzcI+c03dvv6yiIhm
PFOkY5meOubG5XA1Iq42RWCGXQfONYJUGtLY6/a9kLSNONS6zTQtIXt/m5Z4HXODZFsN6YWon03G
6QUGqaKTTATQbEOxqyxlSDp/yxx9g7LwDIH9Nys+kisuwnsyis39cwCaLtWV96bD7Zsz5Ibqy5H0
OCnZjx1qCpxKug5nMJWCg8n1HJKw9xvO7TELFfvyq2Aj+/aSrHPEm6vlvu7dlZ+be3i5Nm1R0rLT
990U2I3GuprD5sUdWDd+FWlgOsH4BmwcjL6qX3czg/IORd44rU/es3TqllNo6y0Wg8aOJWb9an4B
ZhFd+dmvILOlE9DFlL12aNIVbSMbK/LZj643SebjKgHAy5UC4o+gVgbcv9O//xmBiUrdGzSzwzAq
K2MkOIJZ/yExZilrJme0/42dAC0sGq4XD8tC0PjOJyd4PxUN4Zw/7H11yilHSaEPM2tQZc5Bs4AO
3tbEuaybimlj4yIIRzwbS1dtE27xEaUviYaEyGDiZa89fQ3mRJeDdDyeiWl+eg4uqxGlBBG128rS
0L2db/8lBDuipAjnpF7s48Z2qDINGM5c6IipBiqeLkEfC9q2zAxsCWMGSdIP2Q9brKIOG7QpHj18
Sc+9UYYWc6FU2hjoIOopwgAVaCuzgvVKqRP8BsgTgeNhf0609kHH97HWEr2cFEfxKHd6hB6EP0zF
dXpIS6EvMgniZQh/jC55q/Vr8jA3Q1Y5oDTKogaeRugvtOWQfyL+EykqkOzDmdF4L0tQHJnP7VmU
IQ2TfXPpEgiFB256+OJJq4idR+QVpEduytEYLX6JaalThvD0tfTLJDYW5SR1HRyMC5ifSpU3acpz
TNGkOQU1m8vrFiE1E1LAQkLzHPq/kaq+zpPhTvcyr83SoDNw6Eu3GPnBWo+clTvK/GAPlWjJMghm
jRrLNfXqCaUabWP0xUzxn7TLJ1USeTm+7TygKO6vc72qIF4ZE8v8P4iDO39dKkk9LVQ+HCNshmir
KxtkY2H5z++VWdJWici1mVcC4gPRi9d1gHY5MK9yOsIi1YvPsf/4Oer3Lcg/GAD5JLlQSRe/mx7W
Q/HcutO+5ZVLHqpqNAQkYHjysthIIATQSNky9TrM8nBkS2AdATmLuyfHILHj/UNBgCbDyNVtcqTb
f480wGbfgqurVSsyS1Hs4u+hQ5oj7DAIczsqjTEg9KNVClmkNkdtradceIhxsmLImLTkFVO82YCm
oxlJT5ornD5ReyXpra4GGs9uGa3lszuBtbw+LESj0BC8/+V8qPYOgXiPgajSUFPyfTiO8Nc47lvO
5kyoAIi1/pgL1y1zUc/Nb5w4MLLV1+882Pe2nim4iphLAwTaNVR7FnKnWFxGukvRJv3ue0FGvEZu
GDL6H4o5CkNnapj03XM5cJGwKRKfncpmxDIlFDrArVlLpDVZok0E4uTtuLcNh4QyMoZkKHD+OPTm
SQK3Dq4tky0B0+05nrtGG/+NJFaJ8PxgLAXB2oScoxN82Dq4OxCx+j9Ngc+sC+cskC+J9AUuylj2
TAflZKyiytTxumr8NakFNuxGkYr+jwYaVTTu2VW4saKSZv48pVLK5GCr6BDnM5MlLocVUeW0mYZn
5JkYVTBGJpxwdQbojKFcZz63NdMW0Xun7I+fSAMByZjIDu3O5sQ74Rxa46Wy77Z1sl6HHIJz8ESK
HrdzLjbgviyBt27/wDV+t7XtO+wY4JPyQaKV308j8c2yr2SJmenZrfeEhcAJ9x9RVa7vIzPEMQQc
w7kvqBU19WTgFZtiwJ2/87ES6hQUfvgzvYG31mTcWH+HOxq18rOlcY86B3n/ULm2b8FTEPWkHjO1
kyzJAW3RmEGpXFZ8m2MDiHClKlMKUewCa5PwA4P/4VAVZCaNG7+Hay/aIMlCKbUrqnLNFdH/KVMA
RjS9KP23y1gBuFvPQ9RrkBjfNK4JTPQUYWj1OuY3p1pVAlAbDZLeEDpHF1foNLbdTJ0KkJfNEQmH
UbPir85Hko2maYWZ+U3Cudxv3IV0hRjvo2mG14LtqLQIsZVvSAKlk1kT9whuWFIMAoEVJaZS1lJ9
MBnVWXWl3JztfYeiIlJN35AFryCv4drbJlemOOjzRGJwwZG5KwarGTPlTMH3DhKs5q6dpgr1UFqQ
xG3rZtUEFP8LLTIRWzyhWzlhFnSebL7Ab11XlBeCfW6Fk3hZyyUGoqRObTDrcPHeM9d+667JhvB9
raeDBOnowuT1bQNV8OIJsh36xsUEFUEpW1ttfvbUZMINf9zyUmkniOhDnlvJCi8yw6A1Ng8XYiuL
w2i/efs5drGLvi9u5taa1Fx0K/o4k2F4ayIBiKjbOlbk2pyyE0fzRQZrJULa4nLCPLJTTKriIPVl
u6QA9f+6X27jMdmFIXeGyXi75HBMaeVozO/ElwFy8PiJGaahTLV8FqAaVD2Rcn/WMGiTSep5bClZ
SdmEZXNFq+jwnpsjThPCErMpFIdmpvB6UcwpMHyuvvpXpZzwKQEK0yqDQWwJ5CXs+UvWkDpj0nuv
VPHDG2qIXpuz8JavACfa2cY2FevVVMs0WBRUVwnfxWNBSbaI1lr8TJ3kfujAW1HvWFCKQhV1YX0g
eisyQQ7/iDQYAG1CNXJWdzhwm6W9xvx8KnDsqqxwNcSyA3StLs4Xec2SwlAmHuGn0fyWx/JfLHSZ
NAFHtkvFIsjiux+EnFblJY0b+8b7J0XrzbpjMCIvmyEi2qc7FPm/BCru1eplwxtdBnqjgAYwX3gC
3H1UCSSZRx93Zuheiqxtt+x4fqOHoxX9hmxid/GM3Uz/8501dpnwWQTV0l/a5no348WlGuUu7LtG
49q+Bq3Lp7PnBWQYrEjmNnMlOgEEYaiYFWkoX7X1Si6w1o4zy7nMs7GcRp/VIFL3SjLm6wKsUH4a
UfVzTLplpzDGpPZlqjcCrAn3cLodEIpHkHGh74HehqS19KazDPtX5z1vhF9MLJLl54PuGv/FJ1zS
n92f+SCfoVB8L661onmx/6laSs6POky4XTD4L8VULQAJFTSgNxzJtxklmTmvf3QUEUVTG+SWBDc1
DwTh59p2eatMY8aScjmcXCDdEjbCEXGRYiuqe8atWsKLvkz0fwejvPXhRZeGXH1XvbGqC11ajFqn
0XYJva4AdNs6VaTdM/sAMj51OrawDeYJ27p5KV9BQ9y4kpDY4GkesMCbIdDHMiOT5ct+kgpmgrhz
yhM8Dq6lvUI9yNhX2tqWSB/kfyIpbBa5EI3XzSOuB1JVBvOtjRkxvB0GJjv9nVGevInXobJEr2a0
+UOcipPJXxyE//Pnrf9FZV/kpr1+3blJQxp7zXkfAcM7TElaUk49bjTPEL6M6iEZBYJcO4XDdLx8
8clmMLgVEOHjIqjqwAty8IQ5zgwQn13ZZ688bDM8E7cjLyYy9R2BrpyzMZOUZyPeruOg0DojAnr8
AEDtKg4OBcXkFlPiUw/oR6u1nAbJjtt4Ve38PHgFUzv5aI31IBaRn6uhsreE3ZtM8jVUZkC6Ex6S
XIyXw6VmkvF63jwVh1OgnIGt3yChu8q+IOb8gCd3tpFjdym/q+WvNf+8Q0+BUmoJU6ltKVnjznea
eEc9iH0dj/mq5llvleNr2zJR6SGSD1NwQdFmRNwqXWOTKPKbogimdt8gGsI6m9UI0hczGlv4aYKY
jA19RwoEkhAME3NXD+8WBwEjB9jkSHS8cwKkyBDtxwSIL2dkXkaqMi/3SqqW97LSsgkFXL7w5Xfi
TDQ4V174xSCGbdurAqmbTd8CHjSSrfQUmr0qq7KcwkVybZhwDDv2WEslHpqKFw0Tv5cMi6WLwdIU
DijAROoPcUG3HtXYR1zD7o5bIKN7lTp3ZYo7ViVtXlZItDQspffotZt6XaG7dE/VteJUNjsVILjH
mYsjIk+8ZRXgfsiGxq3kTlJz/qoYUyWCoLyYGtGCH3fWE6Vu1J6YNkqh1JT+RXNUpu6oKjTWkcGr
DUpwaelXuYUg/xIrsUn0R+7Il3IFaond04rgxmjsirzJmaRrE435YfeF1+93zcq6bChODFztacc7
gSWFjPcxe8EQrpAGo3/a44UxOFP+nFycUA3c27/vFx7hTOTjAhOfcPRSCGlN4PZQ+tRtF753IDj1
1RLy1lX2KcmLSIZZ+DLz8mP6Nmpfn7oaDoKJlI1iEx7AemfSXOXIZHEmMRKQjgWzLLjbT7pgXJUR
g4Y8dTiOhbq+b7MIMOsCC65CM5DozXoTgLBeFBfHC8xULq50BB16xAGZZx8sNQ+glwmHhTRSDf4L
eSCH4kCeiLlzEIFpyOvsXyiItIHpQVhRXU1HjxgiCdvWvL3xHx20rpKgwdAdKSJAB/vehhrAZcbD
gBrDeUzKXdeqnxS1rmHdk51ChTXt2IUd+VatxWGCozLz6XjgPa47meVqWmp4/TQlbSAsGcqBE/Dh
+66PxkTqqhNoFv4LK3EttbyE0kuolF0pHESE+wKch0jbjN2dZAoyzB1iB+Xr7fQ/TEoH0X6D2swT
blE5FfX6LhvovCeuqB8HYrjk9s6MgdLaW/hrsrCoyQce1rR07QOFbhDrxEgB11/+paAlJf8Vt8TG
WWPw9I7ThwzLofoeAzbtmdLtWBSJD2BRvxxpbPznJ6PvD7SQbxOPmejurxPXEDpebJzmybd6duyz
8NNu1I3stCoLYfPCSD6nzjcmWcO+ya7qYsRvsQxnSlgtoypDsH9pqxRre6joD+KFOhmznWObOUAl
dCcCPthHeSMUpFUnYfXsdBg/seJ1OTQiiKquRGDr79o8SRQxE5CtGU7lcehDnvbLXGJbE704KUeC
Onteei8qrvLhnJ4OqXFsZQQg9GP1kqFAnAFYaHO2hp0heQ+ujKNqWC2ISL2hfWKFfTEYYrzrX4Xw
+yBSK1/KsdJg6+A+VhrvsiUjtQEAcD3Z1AMiwkeXv4s9NoeBKXsY0xZof04H7gMLlpJ8I76MkOOj
W1ZaQbVmuCIZDw21wYRu57Kx8lnwEgMRr3Lg4+e5/Yfa4OJ2DxHeGXXu/tZSYD8ULT2lDTr7hwRF
UDI7rVq1wJg9CBFAf+qioe8oVzX+mKjy9S0TuyNPuR1mOfYeAjmo8HIj28Eul/qjQWWn0f6fJRUj
7yia7tZMdBdOd4mWz+IcVio9chJ9hLYoTnXD91mQSu240k0neGRs0rKDHSnqT95FGw/2NfOca3BN
MuuHq34lozyBkkhH/S+8Zgj2qMiY4k//iEOF+gTwSgqMW8EXkLbGjIxQgpYMADRQGXnQyygEzDVJ
4Xk/AmxkkSVX2hPB3Mp80mBezdB/pm7lfpUzvxs59twBiv6yj6BK+0mzS1mYP7qRt9zTxE9+hT+J
Vv/1elrQ8AWNKIqZBcXO0CSYnHZxo4E86qeMzZkOlDn1pHpFaxPd+6Aw98ckVatnrnRsmzdsQ7Z5
iHLMRkO4LknrDXlbeAfbhJUuwsawrnPl1854TH+zJGWB6KS3vrin+BQVKL7CpjB2ddIe++3cnrUJ
jhn/nw+WWyfL8T+g9DpZtp7flmg0yAQLzb0uxgkvkvCnRLGZNKoJBDGTKSatSxLyzwvHmZE50/Vz
WHkiGJL8iNL6ARrutWxPDnQcffiaTVA36UmWO7eLNa9fIR+z3+LXz/qL8q/+vKXOPzeWSkEcqPwu
bpLaG2s7aE14MH/dr4omktUwA6PhPYYd3+dKp23ImJAgMIjXv2Kg15o3U/9uOh4b6DFZyJfk3mMD
dDRA8Knn2Zpg6NHGWQ9MWTqxFdRgAf9QMQseO4eAT3nN5ySTVLQBdIcMR3MEUOO5M55Zzy0fi0co
vxHxdNXgkvAF+I9hgl9ypzjaPQJ2ytmrB62it8/F+/9/YoRnmHxmJGLWQnNY86FHGUzVZ6WjYGak
WznqEl2A2VKIJt/zKAUU6O0YvUNtfuGIJkNgXPWCJdt8zxQ+vrSFlirId9AN3//dBfSjP7YyGe/a
Gbianx6FsN7mVLt9OE5EP8/pvQYLX8txC75wBpNnoYoJdoot8zZzRZtJH+d/HT3Zc/tAEd6wZkn5
WDm2uMgEg9oCZMvohw4iXgx/9rJQDzQX7Dq7uVbj5lrPyCDMWVZFEzOR1ExxIIkiKkXILU9JvBW3
2LqZflYxh4HDO9TgvfkLuqSzXMM6GL257osd42SukDeRVAeiByhY+6Yi5QB9PC4fnEQ0+MapwFv+
fZFhrZrbQKxEOIHcjtuOCUFWil5B20wSLIcZCOM1TySkL13rXA8JHbormxrCXNPoiTOId4JOMqoL
QvZNo5w39izQvn62A7hjmd5tz7Z9KJED/3q+BieakPPpJOM6uTPgTDHvml79BZDPGdMR4pezIHN8
uFZFjjElwNBliBoyGr5DeKesskuJ8pC1oFSnspDS7Qjg8AflAnvD+t180JIh2iY4mj6X1yLMFtZR
g8eijZji4AEFcwk2fRIRBj5vOElOXOrXfhMauRH6SVmJ8NOr2RzxbQrPk00f8c4UrCGwsj/lUiBG
5irCqlyibm7cD5G5fL9WmUc0kNGHMDn/87kdBXSKocAml0Nkb6KuCWerEIpXn/AFYB6UezTRYXXF
SGvwQIHhZYGMnUgbKBdx49diiJyT6p56MuL7RXnaoNtqdAhP4GPAGm4BZs65yBhwzbyolM9/yN/x
4AClPgjQ2UvXFdcXHgLocjF9VHFvcrljgunT0zbdWAF8cLiTGaSGLA3z3Sna5sqZEHYd9xcyDImL
0G75GBlEI8GbJqjInqG3UoYNW/5J0vFKnGoJeMPKLHXIZm2Mx8gfQfGfuQ0UBFMpJkeKIlwjTZrf
OuWxhLOzsR8oLHM4f9i6zUe6OJfmxIHqic9MX9xAl3QziwVch4KyPaGhtYIwqBQz5GTKVPYriTk6
sBA9uNKEzH5L/k8bXPndgCKRnz/pc+rZWPWgqHgrCh5bM8rIeS9TnihsLGFzhpYoBs/HIragZTVr
LyW1LnUJ0GeNwfWpsCThWppzwDAcNg2C+N2xlzfl/gfSoFz4illK5VzNyCgOZIr11LDYaRkdZeos
YZV2JLMC5OBIZsAHjobkMShwwt1p57OReeoi6+L+hrkdKL1lJ5UZnFRQcsZgUw4IcRiV3rhHxcMf
qVnhYEq0vzWLJUpewaFpQL6BAArKnVJlx5EJxr+7VklilqKZnpL5pP4GCaH7S3Dh9MJMdWL+mK4R
e2XoEKn5KSTBungj/CzfpU7l/EMzNpheAN0dxSke+85nxiCYEys2g23g2QupOT6NorUkj52eJLKs
WqAaMolWRrdIxrtvsIkByFRHmbBA1Bqyq2KWTHYf98f44+KUxTvmVDm3Pijbr1CX4VTqLf2h0pWx
RywRYYaKqGx+OUhOvnhhRob2WgxcUTfaOIp+7vQO3i7rczfJUcIvilDZavJe9YmJnKtENv6obVqF
VXh+MBWq+nOJdUbE1ZcGza+GaDp45VAoj5ofE37EnIwBiGeeIL+SdouzonDQulVYY2qn5OiQ9ThN
+oZIxv3DM+ptxz8KwLAy7hQsbVUxE9roa4zAg0okMWHCwPDh1T4kFZKtcDKOVRFSP06OD95jCd0c
0ircR+gJklXAgSpw48nkPJ3VwW1H7yB/zNDXSPRVBfVo/pnEPbHZoyffmE5qMJffSMlg0S/QA539
TqwjrpJ6Acdsus7bP5FqAD4eL/wDAiMAs6E4jo2V91AhR/BHQVwWHb6PrIU7o38tu4mb4DN0PQh/
/aUTCYsyMLQCkXKYU4+xoQIi2DMECNSG1bKlyHj1tsIrqCgFkpfdqM2SFpU6Mhy8UW2vRLNIGIPt
yRVQjAFMh0a8ZKIT/v76GWaYVJ66Y4cFJw7hOOln8rKFWsPOunas1yk3BH2yqizY12Dge9W8mmJV
Jtw7BQjBJ+psKMCu/6ywAlBMi/3JsnP3P8pex3a0oNJx+wfYg5OMmkbIGV+EVXqrBrP9lwLtaZGh
nb4BlrGVxYsdQceiHZziGfKIG5UGx3xmISOai4E/mYgDCIV4yP8J3KHtWJ0GfLKvUehZOzDhKy/m
vDcgkH7xU4rCN2nHhgPDxXYfjxYqrDPYKqsUxfsVo9+4S4LsrIAyp3u0y7lpYllQLqamcVgi7XqJ
f2l+k7Mejv9K4NvKJrtb21eW3ZepNiAbMq8K/gaAo/31oVIAM+r9CMFMt4Gl7dc+h7Zx91APNNow
81EnSijjrOaNbibSQA6yFvw9O7r58+CEzULvsjj+7+6TEV7oxoiD9AwfQ0WCNy8kVlqtWhXG+xyN
jJdoyLEVHC8OPNVGNmGqEHQunU+AGfgnsBFgTrHRv8b1JvDSlbsZ/fQzADPANfo5OmqGC6SqBldc
Dy7i1hWVaXYJcQYn7/09w+oCTKgKnfIbmEndJMzDW6hormd4VfGwQ600X6RdRZoJ+ypkgEEuReAp
ZHk8ImvtBxPtCHIGoSxxv4Z3S2+2adDxwjiz6R33D4xueIamMiLE9pH0XZFqO9FFPYkl2MPYFYuy
PHd5as5uEa0XQoYBV9EMj+29cjymOTGYZZOsh0oSwfsj0fs5yKVV/rU+zDsO99upXETdn9fCxrZo
a6Po26plSNepYkm6Qh6URoo3mG6PE1+/z8PTaXfu80wlRPQsUxG1b042od7CaVqtPNR2nprgsT4/
DDSPXFjlGUp3Ra9nbnYDzbS9OSQcPno7s6PM4RFT7kJ90t1rj3889XD9dBe7cp0y00W52yQiFRW6
wzWCXBNXNSiS7nt/43rtjdtAx9K1yFqRHY65V6PG1uP7182wNa1JDDlacDjJHLWwAl4F48MdAzdG
bD2ugWJYStPEDZO84hU8QRMRzHCYkiKOlEWLCaMQPe8+xgQTOXucAVDRCKuMn8GQ4h87a0ag18j3
K3SqWGZnZDVaWPA399uGNgnZBvgX8pzO6rrwIsuUoBxrnYwqP5QqLtBnwH12Er8pNN8U2mfHqOfr
t4sd8m9VCIPZDdp4z1AWWQyae6eydbb0gRfzCgrHBzqLYfCdxXGaiMam0PYHsTCI75vRSKweND72
wdfyrBJ0wuhdVzD9/3vPJep4G9UBVeVDZKoUWFRjv0ik2wJ7o5Bip+YssnbcKWk8aB6I+8QTbd7U
26MCvj7rTX91kyuJt2F8vObIAbGcMLru2exY2dDvk/GCQt7qO2HBGJci7fKtyI0LtIR5PeqH3cq2
6Z9cqKyp2MGgAHeomADsR01j43kLN31IHk3C9+wI6mQkxD1t98tJIHOP6qhr0nOk5eZy5LxZ4XVH
txUJkidydEM+Kg605INOO+TCHfzG0h/u49nuJtlh5Jx8e4SOT9tTHvda8emYgTslhTRArYoFtFNa
Xx0algKq4AICmBCu+gTbrX0EUGB0HNf36onp1LjUwnJNuPKigcfJlT/oLiXssjQVhUNp7RN/KJ/m
ulOxJFO85hahxjG58EDMY8+0Nf09A+QrtVwevnyMgtKQzHCxr5cDULbMdj2n1AOWLPhVkMzTHoqp
5X8eyXZ0oconzZjMfT6WTwMC0Dh5PAuE3hRrnzqD7+irTI4gNEoSoD2y/1yUok9/NY6s2s3IkHZu
HEYL7tHoOmE4JRRoIkLuGqnNdcGNx4LuPNE7r2xAvsFfq639WugZhTDWTqTWVdXPHiRyZGPQsGyq
ZCrf9Ou7qQnalbrZWnUzzFiGNcLin5NsueHpiYsTChvw3uWXKe0ZcbdcRWMJO9W6qdaOOZ7ZxPFI
c5EM90FbU4YsWw3SIdqjGmXU9wuU1bZh1oNtyfSv/6A3iILTxLNhovzKukpTN2mU3AAct2lsDj9i
hrUimVke4hp2X3BAEtgM9Li234q0dTTQ9DZwlydxpobf587wC8P9l7E7EvjBuVisMR1hdNMLnua6
d0A5XKuGCUvAl6RLldvtv9wguPhC2+LcMb+BYGKo0C2V1MUpo4TbH4ZrTkKYfFThgqqCCJ2GeDzE
q+aXQNRKEgc107fSOyPoT0a5NZqjjG0J0vQvpZOmvN7MTc3lR/LZipQaSwMzJ/FT4ssIJxIGImhv
GjHNcJO+9+XaLGB+r+frIGFzic+uOhz/0VkNDAYqNXVGttXwCtdbL606llWhkFre8vLMNAwF802c
Tu+4uXxwcLxj7ILLfx14dTqoUSE9y0b3tHByrFd4YKp9nCOlP2egVgF1Tzr2YikNXr6reCtnikav
DCvSu43TH4DJJ4gIFMuRDf8tsbZWAIuv88QnbsZaMZYq+TkBpmMmfuoqOar4gOHVPj6wzsQDbUeT
WSYGCyPqjKE/rqhnHG6SWypfOJkBcCxYeq4dYUOyytLbpZzrX35v4vucIYH6YtXUrkzuXnozGkEu
PTZWn7KPpCl24tz/55OqI+eT5bc/u0IxdFHwdXVCDTeKTmulKuHn/ukj7EM8w69xdo5YRKs1MCIL
tB1//sZdfQMR2/FIdLOSnDRLCntu5AS9n8muW+GNJo790s7xHn4XWDZeN1iNVjgM00T3Ae1p01+w
2/oGJaFluaomZNFtnFPq44+NpvOgDuT8uyWela4F47lbetRB+7/nSsoYaslh+QC/WgD2okoAa9gy
8xIzBWlENo46h9YGnadX/6XoMqL52RxKylmYVft3lfAX/Cecuw3HF47lavBwmyiJZzENcXtRjdKo
fop17bJfDfdu3L3ro0JfIkzMyITCU7HN5e8ceLt0tjMQY6HeT8Oza02i9vc5cwqW+gRqf2obU5wF
6m2ymjjpvVmYaq7ouGbb0yu82Z5VRN9DTwMSl6I+HsCmEQqG6KVzDIBmesDQo8IqqR4AOI7vsJyc
NF5CCJDFRJHCAuYu+EjsO4vo7H9lHdNRUmwlm/jnGHfmJdnh2ZKZh+J9gkcD6mqse9dJkNZNF6Rv
feOGSlSAQ7E1H49E/mR2IEzMCWkyWjuhqyIMVZTTW0icm8TJIHW/JRSPyhWUs+rMn9AOOXE3h4/S
7Rbk5aIlZEvkTvdlKh1IGZDi9H0AU6UbkRF8xMPlpgFDW9Dfy3ZsnWRJr4Wt9qZNddLs09UCFT9g
37ynpQ7VPOlUbQ1ehWAaMr+OSZEmjUN8jkYts/xaduZ0DgVLV7Q+NpQBWGM1PSQRkPHf8CWd9vuB
TqigPLMZGjUQV0qphpYYQskeOPSWU2tT8USJ+qnNzU8e7n1ljvvVFRCds+9QAtgF+oSTSDm/S9sE
6SLiGWwG9it2gae5WMWoT73Pi51UCLFW1BGe2pSUT09F0y6tdNo/DxCHh6ZzFznWANGcYzdtLiz3
1FDMlsLCSxmWMVSOzOf8Fn9+4YbHYZktd3kIcINrx9MhQ7AG5aOO57SE/ww8hVxWnk3hzbWqnQnG
iEj8xfnjoZiwaLvAyIzW5PBpiB+d9MF9GdHfrtm4OpOb2aRAtDCvv+Ouj20YM3ap1ti2O1SPBHhw
ptjUHLDSQgT9dTKlsCw4E63W+iuV/txt//MAN0vNa0hZsB0JSU3blfoce8CvxiZLK9WMInJWJZak
rwcghmKJS+xV8kHrYFMwbviVoTWZNegdSFZ5vcQJvEVrjeHhK3VtAhaR50JUzVTeTjlXkHMPGwkJ
dgRIcY62wjnTdIN/gipm659HTuDi7qnsvLWii94RqIYw3gg42uWF4Q7kWN+XhF7ZL+f7tjJknaYF
65P2sLs0gayF2ouOVPCDqyh6UrRJwqMWJ0c9yfnaL+oMnoWqVIgIcJmc7JblnMKuHvWpn3R1H5yb
fp+QckPSB1Td4Mbjo/5qwDL7xa05SvQD4RloKa44oQteYSWNIRl0eCWdcntyFTMhB3GpNF443NnU
6TniyrLgV6BMgHqQdasbRMnXSDg5oZx8mGXZwVfQGfw6jKvo27YpcaykE6Gdi3OL7ruxIkMBrKDa
RlySt5iSxPE2dgxnppU4QCPvpD6ZYCrdCmkEQrohb4n0HK0kJe06zqMeu0ij22wmqVDZRGXy7/yN
3boQ1nN2OdI3iNlP4ornQ2SHxajrmcrBg33ixn1fYph9mL8LwfLXy2k+CSesSnOL6vxkNvdXKPeT
5/v8MRe5O71xLZjb4Sdc3wUekYeWx7hY/Hjc0HXlDB+ForHfNM9PawzPb5PyEquRv+6tSVWClyku
1Ne8ZFxC0HJwzUdBItc+z0G+eOoxnREXg4lQACr+AOdf2s1oGHwGJ0/FNRJz33xszmSSpLv5g/RY
ymoED+fLAx0exx4ZMdsql+22WZurnel89BkDWzN1kjd28M9/pqSbT+VNgNo+dno932ALuOoBlAI+
vEY105gP+0p1GBuLAZ2J6iv9DNadi7kH0GzMEYf9r2OYqbIQT9GVCvlereuWcmJmA5ajdYicsch8
3gRs72OXA+y3DQ/AuZqlvsQcTufDF/lQ8hCSscR47NMoIuH13Ug3hu04d32VQYl6MEjM4PZb24dp
Mq5WbJCBTu9u6fMlb1/pyt9kbC/tr3isUlKl6RYomNqvkgLqzu75gOQ0ISP6sGtdDfaMWpi9Vsou
pNeTdiH56YOWF/jL8VGxZte7NYvRXqtOZ0ZOs+KWArNsUOYrS8axfrB2rcJdJ+NpMryHx6ahYXWe
92O4aYGgTICT71phAuCRWKBNbPC99p86Fmu8uPn0pycCp0T2fjZBjsATwK79AzGJj3Y8nl7bYIYG
i/ckE12yA6Sz1JqbpG0cxqBlsNTzwYKnnJrzlq6u8897WnXck7z2oXnOlBJRj5qkiUQNlYmdlcfR
5rl/CIWhNoLSAEycSAP7pWqN5qlhjakTZjczQRixeyI9VsRaHWpOGVkK+BTTG807SfK08A1JFEWt
vHtWP6dPEE8ybnpi1X7v5QbEITPN9AkzzvjGIidIlUERpq3+6UKHOUkdLGEV+WyK7VK58l2hG9u7
Ro/a9qXsCJaHpqcURi1I7IL2n560vJMo7I5RYoUvNzSk8GRCI0L84rIQyhDCU/wgkYOBnM0qeNef
3iPcKUkj+Acbaw/fWjBdK4C6QQg0Z1QRotK6V2FDXbK4TU/aj+BiwlCjUXS9KSHEYQjDFVJNjYTT
oC77H6qF+fFC7nH8GdB55V+4sk7+uCriBe29qKqjwXm8feVtmDp7pMVhQIs+i5bi+TBqj16voi8E
E/iJQsha90rUBY5TYB2hcmzfRruo/K7SY19g1ph8jTKq+pnP6GEhiKBT6xKvKpM+DFXytSNNtq8M
KwnS9Muqbd5tGNVXTMG0SiyiFTHX7cMnasL0MoTYbHlfNREDFtPiXqF2vbzmD3+jUaUCGoVAOqjB
zTU7RdPG1uYvnxk89soLIrhkYW3iuN8RDfmpzr/3/p1ILNbRX9vzWXpb/chig2G7StlxF9+rc0RD
FxWq/pKMgRgxkCOe/BG5Ke5bkoNLEikPsJgvwo1LtD6Du1X9sQin8auz+p5mBRdFAFolahOFyEgl
bI6tHFqWo+naGHBp6dU2BuvgOF8R35CKqCwM72IfiJuzO3P/t7dQV3D+w20t71w3lTg68nLd1ql3
xkGR/ZGQdXeXHCaQ50ZETN2AKKfAkQ2wdYLh23EVpi+uc1iMfBFeFuh+jI/QSnBgMGpHN51/zqer
Iq4zTEGzRbE+O8IOnHTvjzEa6fU3CBcLY4HTs0ijgptml/0ypPBqKLlbyXkUQ3GRSGwLSw+nlCTI
pJRYedvDn66krEQxFookNyX8YaJeGv3bE3qTOBVzQ7wYH5i98L9CmyJNbxnU+vzq/C83NOLdf3ah
gIX3dfZI5r7oUDEGysGEjlSwJ6ZJdMVt4rrGTywPiojlk/VwGGnn1Htpv9mnm1lmjqs300KPjGUv
IXsRaIhdlngHZ9zkDYXUsQHfAWO6qEIbvQX+L6Xx7L4vYBYQdSOID+pDwcOIh65fc0GznuTQ4eqs
zOvuKyl6vXku8z6SHD3y+jQtO3+80x9Vg8iRBHfZ5RvSCogDpqmMgKCMtzkb6aEOAAfTsuvj59ph
HnsNVtyjcX0+J1zNC3aCQI51shCstTFJdv578XF0+H36cjTZoScH4zC8GP8FP1ivY2M/2K7m3BJW
1FPZCgQGo1ZFQbFjWzIK2ks7zScnmazGOLPlVWwYoIhDpwaQB/qHfrM/ZuOSSPmZmCQ8BKMy1VGd
ZRlLvdB9AdQS+f9mNeh9rHJSVILLaWrPA9YNrhQkkeANen46sTbiv7LCTGqWYAXVywYm+RIfIPlK
AcwAcXQWnprM0SnHOOW8QdY6W91HY6YPzSRej3DChVSIoPJfuWplO7KsC3s93mlL7dWEH69/cbOT
mo8eBv56QmFnmCly2p+fEZhquwAp5aLFtaQPiUCaVejFH7C5qLNG8IraKjxTtYKDMEcAMlwgcwTM
f2Zk6/qAmubpXvKnwAy7fpTFbZy5+SJTwLd1Q10+gyewEu3naTT1mLqkwsos5rX29D0bDZHOuQgS
E/vtqOR7Msg2chx7l4iTxjlIus+Xd1AM7w/ksDgWxqw+8Q5ZcwkF2LNve0MDVEtV9T62xcJZjGkY
P9pP7GTfXsluuGkZDeKqPHd+xbZ1tZz7Z6tEYWCH/8n+8Wwg1jN9cZuYRLfY+Wo4TkPEXTOkKWOS
k6Hg6UI11S/Pi2ac+MbVLH06Q2VGpTCGa1D7I0hdlpzn2HtwzHEN4tou2J80gzusMcLQEHlcEyoH
6jXtXB6psGN3HdyahtuaufTJMCF71dTTdChXReXPJRF+3uXGc9koDXAxtYHzts9EQ5hB7goO8dm0
ca5dEguhONzGj0CChVPgqQYNqZsTNOo3/mM09jmqVPL1iyYKUpFL+WSarB/f+e0Q4vlS0RP3Aavd
rbecvZ3A/J4xzGmJun8ki63ZiNZnI9GGEX2OTgN0GC+RTtUskksK/sShVTd1XA/y5qA3FUOjog/5
2dxC6384xy1sq14NA44pg7OShGKfvC5XuQVe7AX/sJeBme5T6C65I3mOSFGHWg8vdnxWTMFaL7SK
bMYYg7MrOKWKJaGYYpmaqNnlREyx4qDO3ztklZdrOa4dVSrmdxu/l9p/NUyIh3ctz9VEbVqKGE4/
mnQT09SLd5R69oZ8SG8IY+UovH2m99DC8OPpnkGiX47hRGIF/RetKArOx97mo70gx3AWEKkzFydo
f8ZxJv2oJXzTKwD+fuba1YmebyzSdGmTVxMuVS5O6+L3Re/LTWTR8KwT8yZHAU47uwc0C8w+LlSz
5oen5sLJZi8RvnBXaytK4s4fOHnYzh2pUGIK4A7TsqJvK57h6UXHlX7SZxWzTc2du04G0vayCOw/
UFSBe0rqGMoZ9j0aUNrFg4API5bm5+V7AFh/ete7ptGnznwprY2VFHaX5A6Xb6844Uy0Exmw5M4/
5R91EK9nXUIPNF976r9h2xt/yZPPrmCUevZCED4DcNrSNWM1jAPD7udXihC3Nkx9oCywoWGbcwyw
q2tNNunWngpbrJ886Z11PVyOdoFMLTE6cP/9KCcoS0dUCfFHZUgksdrluKfQUKaXF9Bk6TrPIl7h
tOYx7io6wGJlnKIComKGvuERyC8PQM2gYEPpypSQEA2jlybj7BwKYCmpakJOS3OJtMRQOVQwYzBV
RCr0hCO9mgGlhfxG8FWaAQqr/fdC/pvmWea0u5mXUHfzFFmFep5AqgHMkKf23aeahm+4QvALLVn5
M0XfCmBiIM/0nYWB7D/jI07NqK+2oMapz6g8wwQy+Ylb1NO0Eyn5LKuGjIiq/9Zow/CRx7UzY7G6
MWT5HaJHp6z4OjHcVieVpBb+bNu+kxVry0xtyCG6Vj8eqXlhuFG9EP1b852QimtKQwBuHy8m3QtM
0KsATdJOdszueCask4+jl9Ix0+JAGS8X2BuFlP0k+SbDQ9O6XaOkUiNQeFBsttN/HGx+H6NumWeK
sW58aSl8WlGyTYIR6CQ2VSXAIcAXJH4qUNjnqY+U9wb2JTzhzpANOWtfLpGBFk8ARHUryhYMbMaa
OallpI3tkE0bIaDmfkaB8milCvmezlNLzhgQQ8tFGLIfFD3TOmcwGx4YYZKPVwh+veCuyod17EiC
2SHsbYIkq2ls73GRq3ekri6ZUSaSvHvca5LxaAxAMeh13bku0hqMpjJwtpl0YBhMi9SiDTEBedSp
zwVFjuUwwREIL7LOcnX7F8H3jThVT6EdglibBSy0qQIQ6VYA9DvUX2J3jamXbZk1RB9aKRT8fo93
YIdZt/wrtE/h29AEF4ylyH5v7OPXhN41rIWnKwgT/dyvyNrdY6GSl4iQROoUWms0YdK5QVIttjIG
MF+PcrT5EFxenskO2v61yI0MBlZHuxcSW21/S16aEFTvnb7+X/3hfbcbxzZcgownMWiyHyuxdVJM
/qpYWA3wr72xQQA7Ary4L6s0jgkKQhmDN4lx+sl8jGaiP62i5luT9j9/fYZ2ZzNE4T35neGsWBCv
c1MgoL8kIhueZDLPLINHq4yhrxUk7fkSgISPAeEVcxMqMMrsJQVD/PkJYE3bxa2H5+60W9DV9sqY
gtsYUqRGMYdabVz+MOHJiKLan3iE6qe2lNgqhrM8I2JZhraCrJnQI3gbZ0QA5M9DzlUZh6QhGHUm
PF/GZ28LeVdCkWJoqIqPmpK+9iPaZkZGFlOx5DVkOoNVoQqco80etbcLwcpErhNexssyqtKGJmyS
mt6dsDFmCCBElr9O8LIlu9YG2uM7aZ0/mgc6ogW4sI+ndMjd66VksyFQLsNu6JBEgK/zKFCAZh1T
b1EBX+GQY6+78qiC8pAmJ6D449V+JR6pwdphjAzzebMv2d7OSJy0Qt/WJe4QrtXZJ6GDPFULwLS8
ZKfhTAoZF/k+6mn0FibxDX4q8m3DbC3S44K+GWpbYNljRZuSHplcwijuWwVUR4bZYn/SKZ6K75+o
GMkYBSdhyzg+eU1wHlIkWJt5go1RL9DWMsMKqTex7Mv8jYyZJb7QE1yju7A4ZuyvNSCuORDkm9a9
toSo/c3RWQ/o13rJgHzhyLIu8xyu9Fb5/WC32BBo0p0ouQr8SxIPs0GsdoHEWc4wZLoOVJewBmgj
EfOkcupU2cu8DGFlHAiM9sFQjFuH2WHVd+T2muKmU2XpHdahAZVcwMfBtAVIl3UboVCAOD1f8csA
bkqvzmanf00f/PFHxbGCJtP2LCpVEEtZ8Z+RjlX4nhXn16y1Aq2Ocmvk+s61UuVftY33usJg9O0x
Ay60QLIermhR00slKju3J5+9dTBDqNdIExVhTaDwvAUO7BqkGPJE3FSla4O6pu7zpYBD8wWazyqY
AHJDNOUs2yfMwQIcynr2IUIvO+vjmov18WJqAwjm8Fc3VAv9daE72z43OzCQ3rnY4ax8CjJPHqt5
Iw0RNEChoYLfSxDftvIj3M57JG5DXi1T99wrQUFoZODXqqv1f0IdLs2wUap/276+HijC7rNlkF7W
nmhWXMk6YVHPmnXr/BIG/PXGNyQWtzCFfgW5lRnrsVkNLM/kDa7fyDQNY+6XWI7QDo+AgH4v9EZ1
zdcD5TI5fRQrBO/yVn731EmFzED5vgy2PZFQW+xg6fcyoCKvf6vloFScpTiW0STv/K5l5A+jW7hn
Y8T+kDUGNLFiUtZSgU508AWJbN4TNP0nXnEWMydkAlZM/gR9fdvYo7TaATFuIaXXzWgnI2OcDnaw
fNla+uWDhkZ/EO6A6sJD467d7QrbiuMbkgM9IoNaVWNoemh93MUcc0fYS/GKToY54gc754Kxk3LZ
AAUUY1ZgL7NTYgIb9oRBl0BVoz0dfo3Eyzc26wCnOe0Gk5HzW/x5sDDLVr31VP1oiRrJPtRy5owv
bgeAnt8RA9XSyOdC26zmGZTrfJouvSpINQuk/C3WXOt9XH4HgeveMRqSimhjkfsUX/MXroHx3+dt
QTcqK1jM7JNgfqBO66lf+XtDCSkaINcpvDcQes2qHGsnAezWyHZf4TBFYEXbxeYG4aS1pZKsv1gX
OnkZVuiMBzXDkAPrWQFGzW0LEnnMn8dAs4MLTxhHRn+HtvGydMwGI5Vjef8cUVEWHRxxC3tnWAGH
6pmSacVN+eggMiSkDtQI/a22Yl89r6q/d7xQMKM03LBJg0UmGaTVHVdKB6dJxtS9fFFqMuA7uqPQ
GpA964epUkBr/VbBTR6/8RxxdRmLdjj/anDNg+vKcmAIMkAhY18O6nrLs3MZnlZt+UiHbpo0XjlT
fgzJbS2XRdr8ZdsortafQP3OKRc04Fl31GLHINSwqQFkQYm/rkOELczTrJscRpU0YYrHCsmknZRJ
x7sIKIR+rVzCSAdA1mXYgcZCtZ/b964Aqui2zjPwJPAqfwm9X5vvVh1VOEZrshQfn/G+MBa69ZUq
Khcr3dNpC9e/8fmazBdXsLOFoZ9tBSNj9TysA1nO8lhrlWotNN0JEXmHCDfMyxf+XJ7FGrHl7fcY
5Nnlip2UT7reIANtCf+CeVjtFuQmfLELyXr/VpykUpprccWNzTNf5EFNVkmv2HyEa+B3JTl/TQ2K
zAXZjtkO9o79tYDeeUy0ojYPqhaNX2UQTRPIDLSF9/kiaLKGdiEh1+Yh6Z9LtOaBw5LGnRpUy0MD
oxx7v/8DUyOb0ncSNpNTyxoiv2lCt5nLYyA1hbqC84VBLU/GgY2qkCG9Vmq7nwbhnh1LFB+Cq8Fv
JlsP9xMUkfBlQ/eWnEn9Ip4eQZN2cUGJGuvkYGGppTAm3PQMJfeoywUwQ6wv+q2m46AHIVvgAuEO
JpZ4hb/Qr+nlFF+bDh1/mqIvo8Z9PgaKaqSJ5/7Ygyz8iz6DXk7JWUwSVhPAvj77SiChT3pquE8t
elF/g+51fqRCdXpfZcRPrvRpjPjiRnhGTCJuZIgTt/+usnj/XCM3pp0o+fpxWwAxcOo5pgtU7TW0
4qyIZDJfkr1kBzdZf97yoxvndVcbt50379maZijjBxkxBfWKZT4/+h6w7ei8k2grMlEXYJgWzEYc
VNxViRbBZxp7Bq4irknGc88JAj0T+6CUQaKfQNQFwq+aTjymmwZ9S4IKhXYjwBRRpmTgFcPYrwED
GT/0w9iaZf8qOfOyP8tF8pu6zPFG4SVR18GEIDXtJyB1K2ak6TycLoRB0Mh1pqTzYKbk4rQhoTP4
qIH5CmUqHi6458Xbzj6ktzUB7lClnWkTr5L3W7Gx9erxj4lujBeM6YT3Y4jofW10F8i2DznA4h/Q
aeSuggT9faD7bPl1PfXdzGlhUJYPvXkEAVj/2Pli3RYIKCzodzbVoVAGD+FZe7hPYrvAabtjmODH
TG5mMB92qBO+egZ6K5l/Xy4OQU9dtlDiibOza5lTEueWWqYo83u4RmwZT4u/PfPWu/C8I4Smip0b
ZwuFf+dIBfPcp2zC5/JmpGrBP1z1/LLsF7jAqW1OuCUBeEIgWPnjldz6qXK5rge0R0v9mEdPuJfu
ak2pnceKV7OPVSB9a7dYp4Lv5BcRDOmf/p+t7bDTXUnZlbrHUQikGO86XNDEpLLBHu2WXgjtHjoV
caAiUhjHCBEbAOE9IaL9KNRWiPaqJ4VQuRsj+DO3/ISkBeLq4KRLy4tEK43HZkg+gZ+79+WSDGKH
wLi4vjlAqf/DrGUEE0599FgvGe5+UzdI8sIC9vZRRsToQSftN2yG590qlv8s+kuhm1sUPy7E/ovn
62ajNajK/hjgo/UTVObpUEcJVxuVfnF6ZJ4WRQ7TRDfK/a+FwERS/WVA+GkiwEMKejE/sZePrlFc
GQM6j0910VArfpYz0vr8Iq0sUA1fyaQ1NBKRgNAhPvjkvPeomv9lwAUEHg9uTtnecxu9Q0l/++Y8
n+dtJ1XeJqOgKaTmS97UAInI3JbQSMjcMRUsWnNfUM/J/iCNacy2iEML8ZuCeerwiQZAsouyXZy5
X86vCM7LcWYMIg6LElnivEEaILstXT0t9Yjsf2LhWayH/dcXebKaJ/U95WSbJShyxHtLegcU79TR
S5J8LwUM0RkS8J34uJ2AH9MyrAHTuNNVWzPOADxYH4fJPqmh90NAYc0elTfdrTpARJ90b3JqnEJf
RV/Y9ePLLV36IOO6Q8ZxitqFuyU5lvjfgvaA2CQsLg7qnbOUOg1Ggbken2XnY5Zq+dehVcXsboIn
TzBCEyJ4f/1a+dtYIpRcbIaS4LxiohdQMoc+fKql3Qquu3py8SM3jZB5QYFNc8OjHCcDeU2yDb2o
aFw5NrsullsPg4JrnOwUBVq7bNwAs8/DjilyVLuv5CRlasFNQycm2fEa6Ge6WfZbILAcmyJQOQaJ
EISinZrBVaVY8C5F37AeJcMXukSPSq7Wzmn5b8uKRV01rWn3h+4kkVDqEU5qOQVPMlBz6sP8V88I
JnEmP74A8BOQveEo38inlrnNUWNXvXg5G6UAOMlIUpv6Nd0VZ6IpzVOlq2jUAt5Zwu4UmezDIP9H
zaEcnujbYoq/Mrl+gXv+Q/fclZfcoYvErjC3V0hVAoUh06YEpdTNK0seFjqyPwvJZglYBtgUD8cP
hDin6O5iE8raBw9LZITJ51Z3U6XQW3VAQLKpITwPm/2fjsi+5oJmsOTqcuy+xO0P/keRG6fe9pz2
R00op9zs0sDbOP5t2cKcw8wxoU4NqUP7zzilykye8M3Y6JOSHVLwBAGihOdZQlPVYvPULdtI52vj
MKfuhcQf9UJqKojx1eujXl7TFxMWIblog3V4uD6ddBoklVsd3YW1ukxvs7AuaaR2ocTNlllfU+Pu
92ZgxKD6NMT00njuZ8AXQ32inJtx+6dHNzKkzEeP++PJq+gVIbdX0+JPI5fo68i6kgZhogghgbg6
KaIhZEEU86hYHIazLdsjH6N2yl2KtYGITgHvo2De/jjiIkJ1ukCUP2SFaR2abCrHcDs/R0zW9Ezw
paC7i2mGdE81K1sR8QJAODLoc6nVI3zPVsjaI7hSBkEAo4Iee6q4+iROxzOCPC98ZGL9RkJNnKGA
dCcLfsxd4o2k/zXPc0wRpA0oxWi7e0pvlrQJtIpVZrFWPLLZDo7k0Xr6TxjnnGwqzjMrxH39ozTa
QYMpYP7o4Q9gSt93kbZIVuxuyhr/jyfSWXj1gC7dE0SCJEmhZM8N28GckUMKGMUhXR2B87b2b2nI
SfF94gR+mWiEX2ojegnAkjJAoC7mMB1knkTpRCeT332FttEf0TR6m6latIsnpmQ8xk28ov8BnJxP
1ftoyojTeZ1uz78c9e5SOOBjlr4K5G9XQRl4eRU5Li4RlWI4MH8bd4TkrloComlO3EltGQ2C1HVB
wqNXRv4fxyvCfSNkEkdd3mF1MumPazjA7MlhX77QPzkfdNaOSBBVMQJpJ68IVCeQjmRGms19otEw
DEjiPzDlmHWvph9IFiiWjQ9Z6tnYwXdDl4C1yfnSmeyMS/atHhaHHtUSm66iLYlCVu+E3dQQNq3a
QiThUR7jPJst7NeYr/grSRVZ5ZVKzKAp59AhaWWqqHcTgVBtFvxxEOZtNvxkCVZD72UBoR5F6nQI
gTmtSc17qOfSU6AzR5bby1lbPX5hAaSLNRTYOk9+usP7LzU9U23MqHwj0QQWCjx4vvjifXvLJ0fp
URbyjbcyjkWSu+obI9UleRXfGx78RX5qLGWBr78mm3AIUsUnjoWRE1C/VNcEZS2Y1hdqopl/goZk
Rhzb20k3D+oTSZR8f7uaZh2sYqJRbWad1X7xJbqFLIofmo5beSAmOqV3hwX3vJLsdxYE5yw9AN+8
FpDvCtUCJAlFqSHQL5ez3FsxBV3KZqYio/g6SKLwBaikwUjvjC3uc52LyfUJFMlmzEJi6vHt+HSE
BP54e+sQ+phA0ZvLV/ZLsdRbiSPUEKmB+iahFua8mLsooGvo+xcuERKsgvPLk69vX+Ld9yA+TFT8
vYhn6hUfAm63q8K+UuLH2k4HRQx4oVPnrNxDU06vH0+UlusD9Y13U3WlJGf4WVjg1MiJBYUHCs7A
I8qVP0AHtxyPhIa+wbPiEgs8/WHXd9nUW6kduPn+zbifD+S+/C2dl1MX0L67YO9EBKFMIIS6PRqU
GWeFrKKjt14MBSJdwSHSp+B7YUctL+o1PZQFOGmByfYqGYzSaTVJK/S7pjt1+43ybiCvBNfIzoPJ
Fz1LFxv40Q0IBweIEHr+EolirV7tW/n5HQirEOjCOUpjxYrx3bKAyjdgXp/DxlxBxUMEm1UNStmC
quCGdGY6RGfY0y631/pRmUvhAc0URDrFV9gAHu63dylqkTMfb3DF0LtxekoXp7LS4cX993mX62eT
lUrzOvOIfk1oF3G91cqdAOidSeiq3PcGcymTe7IZCiGPFUvbag+Bh6j9gt/7E9zusoCZSll+vOqm
mkjJKk1bV3onSNZMi3raGphnoaVttwtDDpFBbsiYA5IOcnOrhLNzH2Slp4G9faC5VKyaBJ1LmhDi
LMK0RHkYFrztRazcIwtNq49WgW3Mt1f2AOTAeUbp477vQTfYNLr/t/H25ajx4HjzsO4m+SI9tHAG
D8iPsyz2hOfArUVyCfc5vbPIk8M6vBeRTPwOiw1bZRdb5dH/+lKNqn0kj28qhs9M38TyFOzc1b/H
RZPVlgXeydYbI+gwN7cwh23mWHMKYw6+2+DiTpK9qGI4HxHS7pxTSKhM2B5GqQxGq/LhTPPuvqb3
6U0f7Q0Q439DfrEI5dqNQUlfwZDWMYW2502ksWl81cAC/uXbUo0mQ8BNA5wmibRDbQ8GxvR/kN30
7hk86pYbln+XpGABDO9TeFng+wRHG2obZBlWh73fx7IATGU1mjzG7z1MDgIZa+GzhevWB3c4oPBq
KyFgwaAkIYpwwxjfN+PEQvlG6NUVH6ivVEkGcvzsQPllc23ZMUgGw106AChhUuLzxJYqGIQKRF5z
x7aMO7atuP8AxcyS0zT0v7aRnNGo2zOxnztgpZtP6ctj5Rmn5EpX7lMb9Rr4ft18I9jDEtlys1zZ
As6qfN+E2e6NPqghIYYHCNrnvlUu0aB5KHDS54ZMdpCNL9+cViZ8XkabMatxgrScthgtCXmbQRHP
DGMo20RRHO1PgEDkimxgByYIv2H8HQEwoY1X4xoHIUPOKaWHLFbr9uVYV17yvb+d8H6/a/vU1Hc2
sfVYGXsEpHLwvdL33CgotZS7WBWHvIOn2IjECoJe5+5lXo+szakATcLUNtWggOVmFQqxGCcBnDdq
84g5bNSMB9ag01E5LGwKzw9up5+xJuCWJISFolemBBvF7UgLpOL9TnEaxeY8eQOAFG3e7uJwgh16
ETgjzL5GWDkHfkG5AgRqgT4OOVBNqplOaGEiS8phtFbG471W3QPCXj80QVq7nitjKSCsaOInTlpM
k5m9ePJmU4gkwKBfEi2167GknK+uxmfIeZD5DHQNvno2tmfUFN7+sTUR8hcUkVSn7oX/DLzvgEBk
bF2l6bPdnsyJcMP7e/kgRptvlIh/iFoLVnto91+Z1kIMd/BOM+dVCNIXZM/9G5nUceyvlgVP43em
fKV4Dg8wxWARrBNi2LFLyYYbv5vPjJDNKJrXiy59x8VbiW+aWLaCO0RQVBZuV4gsR39mYgKxmc6S
aYRlZgPVwdg2casvy2XjHzMeGTV3YAMBAbxJCjGtE+qlZAtz7hFFyyomKYuD8HiLvXUhN7a1fSmy
I7C9NJtDjk2Rzaet3Bc5bqdND7DhANH0c+S5Exa8oQ6EyjObstS6IWR6MfsGX8k4BYHFeyCJct/X
k7AY5DYTcESCjnQ2p4kNt/2dYnK0stUUbm/t3G8RT6zYeCUmlni1CDQRbcd1t/1b+J2ZUeIRYIoo
KfVb/o2tex+7Rn06BUoSqH3fd6Nq+goEHVxe8QD0QkYfDQLnH77hMTd+722FI7JVFOh/eN8hqnRX
RbzLeUQ5Hptlj3pZv8Och8ubqLtuk1Rtzc3lJTWWIn+e7NukWmaYjnedw00AMp1ZDhiQun7GsA8z
l+b8P00GjrsLh/yzwbzWXPsGeFVDQXa1m+ZBhjFezMOUilnU/bg59q5A6V+TyUOImves2AfeWyB1
yavide/0AR4j5T93OF7erfOThEIV+5+XQw3r+kNcFtxNthx2deSp64DHQsNzChPn3Yr8vEIbs8QK
H6lqX/c46GAwYVX7056BCRbEXwjOUBponXtzQWXMv9ulONvrhdvBhqIkn4hA4JR153D9++OLJDwR
288IVQjKwP5eFyEUi+x80+5g203xh7UrF+/C+mSXtrSeTZBstpsH9q3gku0YvQCNZx0AnrGQ8Iam
gIcYNO6Zhfd31YQLGNiPl4j8tnxhGaxy6npFOsMyPrFXD2BWVZngQpg41u79QV4VHLnKLsTQqWqN
4Uc3+mq9yhAN5FrCZy/znCeWp/ZhLASNbL6CDhkArowiQHhuiUEocVffkmPrOK4EKbk1SpymlIS4
oPtOMFJsVCLqyPBkgEXv118oPwnHxqYQAOkgb06UGL9KzZSQUmu6KrZyWZ6EfdpCqDI8oOqS0t++
Md7XbLX4lmhAM7ULbHWVQW7HDTCNdPF+O9MTmXZXWtsgktvSmF0iVaRuJg/5chgK9lNTRG7NmSue
3aruTdVY9BbFruX9rmt1VanX+oLizgVoyqELnm6LlaiM/KeczgR6g4EQxgT3D3ybu1F8b5Wc8H0v
jIcqAHa4T9OtdRHD5N9qDduYaCI038Rn9DNOwhmBKFAHvRk1F8vizvwsUx6xcDN6eaFhPRLG5Gwd
ZXAFjJ76DSaQopA4djPduuU9+XkIRN3MI626GdyvHsDWs8YUPpaZF51/LrtNfFm4VNIM0gRGFcdG
OtWK2PAG8/UwkPJDWfSP9nXsQeXkrzfVD9Bn5dF194ZryKTs8EePZMYiB3+9r94M4XB20sTbaB3c
u1JnzpxoZf1tikMFhhHtEcqEutlqutISyPCBQP0v4vGxxS9ONrQeDX/AEFK3Dk9hhyzT1LGul2fD
fzwt6MQoO6gkarQYfeBve/Ba7VTXiu6zfl+0Llr2whXfWgJ3CIemRaQGZVTfl8V3/R4gO3mfux1i
TpwpHW/eonNN1EDB36vU7AT1l1WOfarfYHVeNcr0TejjGVzP7Xo3a4RocUzBHj6xGdl/NVvWSzUQ
2H3qGaNJqwws5uTcRXoNNweLi7Pdv9eZ0AwnSMeBo1LVkshL+cQecMK30ah8FzsemPnGOH6eTPAh
iNcHoELG8Pai5+K0+AfPiGlf5jJW8bLGv9WwXHumhHu9Xn1p5FdeiLLWIRLGxmOcQeIX67cmQb3E
dF1iJYHVZbsHaJ0eW6iOtcybZnSPKW7dMmPMI5cHXv1PgWe2d+l3FbkdWWLSv3FMqCFih2qJoVJw
AwWQvLlCVmFG/BXierl1g7cMQr1pa0sZbFesYIZF81+sYjHiVryAud3KavuoPNZEG1R72fSSrUBF
toukc4J2DMpZrmXyjXxxNvjwGhko5p70VTTFiVramD1iHLPnef4/9PM59wboKjzI/ppAHNgMoSJ7
+V7lD3ET1+H/4jO3fB43rlbB6xdC54Az5L0loHDDuCTeivJ7a4hffcqe5FicBf8cK3QWrTTZficB
snJtXUQhaqqqZ2xPBg7XS+KOd1GzGcshLFPyoz47ktmFWtuQhQAw/spT1EM+rTK9xCfEavAdjn2x
P0+nLJo9Ooea5ul5Ho96OedzQMZ40uv/NrT1sPwJaLnKErkhFIZclhnMfmwq+V6fLvTN1w15Ryrs
VKqe+6rwmL9/d37Q4lnXXZ19hGv3NoLM7ciVz1JuXZFflsLsrfx+lZ7KJ3iuMnkEfbzemu5zKQNu
Ua5SaGW8gWfbNa+4Hs3apgLR8N2tyFPornzdoavL27gMs/0phfuDHASVpS7aMJgXFIZ6IrOJqUkK
Xh+hEy5QbC2WiannN4MbCMy99+tiL90q0+HrsBIWO7Zn0zZ1Yu25UShht6PrFYxL3hsN+Y5HLJB5
ZaKF5KShYYbDQl7gQmJBXBnPQttjgAGGlj7NhGBH/y9QpLkC3WtqsV7DHaQm0cGEehjcK5GxYxFY
Yua9/wP2pHrFY60n0O4obB7hSdviYNoDaOD5vaDV4vjzS05z7hTfj99ta4YSbjWBTLEyi6+vtyqp
Xeb0L6fuScx/oJfNWhgH/zYzHJrbI5nRwbaADiz3ii0n/8e3aIZazq3l5OE0ReUH4NmKzc2fnHD0
n2aHrwR39TyWJ5Hajej+e4jgG9RZ0wFPGsADRz+S+7wqBvytt1h1N5rGf+nTjGoxZ8aKT5SaTTYM
RCEdyzq0uLDiAfuXuraiTe6lypkiO0LMlBompIC3n0skjqZgQhFxaaCLkoh998aKKAMgcl8VzBbB
+QgnU/SpezTtj0AIrDJ6dpNACJ98ljWLbzHQ+KPgKxxD5NasqQUS7zCBJ3ejarJTiQkwiYVCtVJG
aoSO2rg7tTb1njql5BW11eFCLEGfMh47zwpHMpeyOLeFC2aYfnitSBeDTiTKdFm1HT3o9jGHEjmb
jd8dz28BLtvak82KKBiT5sKlTQ8a/LGNmsO0Xk3y/87QyLR2Sgjh1W+GmxxQYh4CURalT72qp7zt
BhEYZH76VOJWYnNCRdU1ZcjxRbfll5rFzgbNrBqqK9kPh/vW1pIB4A+GSYhIfd2lOv9BzSNiCqqR
qP6OVNLLcpSyCtXk+CYkdgULUNGPsr6SPGsZ5DofafUX/QYS1IjuGyAOhf8JpyFIbqkn7EjUw3jU
boqFup0CXeD7jEbW/Le4Q5BJM0wF6EseyJ7moI12KoBcBUfnSbe+fLt1hSgpZ5HqtueWh5VbfHRg
+RR8uy39Tlq0WqNo9+/3wKAdzhts63WjAUEvrJmDVwiQGYhQNzNr5yEy3nUjW+Yof8AKNL90AWWs
P8dCSFJom99rlhuF+nXnNPJPGdflLuEgajHdp/GHH0cG4omXN6lzarPc1ix53oQMliTA0w54G9OX
iots3oTN9rJEYb6V/uemS8S9BvK1wyu9ZRmlLncvsIWSmOguzh+1LUqXbnX9/nR7XxOtHTKN1tEy
tYAQT3O3SVoGeB/McWWLY1qDUYvrTff1RmYSXUSq/z+VOBHYfXTtmDiuXO26okY+w7Mfc1KFpr1Z
g7bofDK09Z1e5tPkweFxU4K+ZcCyZ+jkr6LvR8T3pZ/53yRTPUKemtefTla8/8Rn2ZGlMm8pPKe6
DA58jiNK5qpZRXqffvtEu+fYHx+P3mErgsGfi2g/YHzMesNwoMKf9owItXgeWnaim2JQzeE9Xns1
eCoi5T7OIBJjVHOguM3Pg3NEfUMUG4Sx7ZFJc6UQWvgILzVQp5MhmomnbvM0jAyKqkeRGkCaNrUm
xL/xOOF2E5NIv6EGT9qGrlyaea1s5Pn6Fp7wTqVrr1xqtJZQX+gBVYL8O0Xw9j4WqkwJtvzmUcV8
FpAFVo+7aKdTpwGSEygAA6xsFE4/kuMN3T7NnzCqV0KF9lCMnCK7uazLd0ng5U3XT5EyyWiYIr4w
PETDLFAxY9Ei0td+TIX4MTh5l7h5CULpsbcZZVF0/8VDWtbHZ5MyHhCVAcPkYJGsT66GCU+yiuyM
9iS7tHMYrzm9HonOqpF7ZL7DhOB9spcu2kAl/B5g0B2zhFOIPr5ufDLqgvlopQmHfQSU007IyNj8
oPk+sSJslPz+tp1LL4kasxvP9XzC78zT3U7EWwL4SSnRLl7ApaEdsPMdykbBmoEDJsrSU46uVcBB
+G71a645nHN6cp8z0rq1pCuMdTRyVoud4TCroaA+t8br1W9BI2lG44NOPqq+r8SxtBdxNMlkxOTG
qHFhdCwk0c5dgLDwEffPOp+mSv7bujTafpAoNkNJPbxKUsQxVpIrdtpIpNf2Mjm1AnV/y/D43T31
F+xoQxJ4WiLjRbVM7mKvCwm9Gfe2Lxw7397q1AoovfKSk/RZ1t0Qnjd+V2RggBF3ov6t5o8MOySC
Yr4mtF05vpm19HfDIbBRb2icZkElMWy3nJF0yHFnE9ABK8nJIHeWfxpIoJt3Nv+gWqmeGVFQ1CXx
6nlG9E/0d0clVNH3DunpQ4afO1UX3/9jyk1Q6hmfO/m/Fccz9QbXO5EkhExSSrYgjstCkpZHiS/G
+fuNS+WjGOm2+O0vgEYEVM7tttUIXJXMVckIt6WxI+QV4JpEMSW7IuwZOmAO9b1cjigK6gZYi6ZG
6RIPPrh3a2sOH3xLdn6lIrQN51iPgNkQolmYazyn12Au1BSXgMrI2aLDk66IfLvKKBxbL8xVa3yj
SdgCkxEthuRM5daeYHBMjoqEj7eONDsArKY90Td4tIhWdhy3f2OjkEPc70CbuU/OYflCzOjG816u
xhcnN52PDUjk9/bbbX4Z5iINguv70lRWfqfNyABkp/34AJQjSCO4XPbFM+HBe40ELECU5esrsfYP
2becpOLEMMoAC34gbcMc/4SucA59WYMyikkTc3eduqSG9Iq3VITEX5UcIPw5XF16tI8pfVnepI7o
CEYNrdjbyyEZSRtVZUn4bONvTPAc/vFq7hHa6fCy1Lx4LQLDHFgZDs7lJYuTY+geAIalpeF2oPgH
uXekL3ufC75U0oX3mGmaPjfWginbGlnNZEcoSKnXZhj9HPHEnv93qTYEojR4MFa+cGoEV1qGEIAL
rPfAfYfCZs/rsGmCIVmNPAztR5KyW64w3/uz8fv80BLZNqf50o3Jz7sx9h2SwsPbDr1my/XeSQv/
QBGTtEuxx+V/nZpnhAeVzYmIJWeRMmTXN090R0cl9PEOTeVgo9NLcvRflj1krwcY6Jmsqqp5VlW5
nnvalERoZaEVD0czq7n3co9S5A2x4KkzVLKddvvNPzjmeGDYvXA9U/kBAbBZWaVELL/RF3nUM7B7
ZosSV4y5yG7nY/c6Q5aLvZiNOj6Yp51vtv47oZvSWQq3M3pSM0v3PrG86DommdcJj2g3XATIMjRj
tFxmYUzOIUN3EfP9FDhp/IKQJKDUJTM7v4yBhmDD04l7HjOX+X4KAlQpdfA7V1APwml3cUUbY9i1
484vD4092EbxfQnB/wXd9CmoVPJDn14jokN+SfhV5zIsjx8dg5a291/D4e0GXdyXWyTuMbbJVnwY
h0ifymhpNhHkx5b2wBPt3XwWWGfiErharXIeknFslPTjQJhUO+O/aeHQwFF2TQiXvye44CzaOSs4
eiOdSZol5UYrkSJl+j4FTPB3Uigt13MsW3U7fahNz+jE/B1iXDFAhCtBqjJ+NrH4NJ/se5x8PiDw
cDWZXClYDhtfV4ns6h0pROPzrP9ieYxHGrlYUEEqDxbhpZnb2gF0hdnUspU3YVjPPAPYWPbwP/fQ
UKKVLGrLrWuKzMUsnP22IGfKbHDVQKNwyVY9cRMF/6HBufTQLzuoen8mTtUOYfjhLNdACdoNNMLR
1rwfPodvcuxx88E1Q0n1JTTWVFD5H35hgTGMHeeCSe2WHe4AsGKsZGWfsoVKS6GFFrwSTkwOdDS1
5o46EIL305Kvnktw6gxaDu2JQ/ZjU4lrDXcULRLmVQ0QHZDlag2ljQaJbnKZADnDIJDrs5SGuVwY
1RH8FunFSSWl5nIUuOesYokSdZW69SaMWyIjN+4QGVjSugJ9Oa0rQKWacRc2REcy35Qr1NWSeW8j
2x8y43lPURdqYuLXWCeycxQxnP4zoVmfYyu2jVt8U2Q3qZFkpw/RqpU8QiMuGkk9uhaWcN1oew3P
0ImOA0cLysE/OlY5ZG9EubbMeoma2yulbF7TE4qfKnshoIC5rAcPdLVLD6yzStptbe/gHTMS5WNx
VDwxW4GScJBuUz/nxttjZPaeNAuXM/dIduSRnoh1wTcTYwds785esqb/ABh3elQySnwaULzv9ToD
F7AXoSCTDw3mKH9mDNMVjzbOJ8I/Dg+qmjuORcAjPuEEFK3tTlt0weT8Nv90CL+j65U+QLbWyqhG
S0qIFfWQnRcyoG70rmzORkdbuY4eq1Ocg3MdAVw8VUL+PJ5nnHi4Hz+MxjSjSOMCuLIgR/zde2nm
qIttnQl6zYiviPqGVlhOD52nYOJxAVwDyH20+LcQrGIVnWmCHTRR6NblRA1Gpz1raR3K/aLSqAaE
ijJkKz5v0LLC8cy47FFDvO+oLUay/RKgzmuduBjACnkVgHuzuW+ERmAcXrXYqAPj5uj/VcqCgGcA
ua276FtwEaH4iYFPvvAGBoTLmCB6IAY1w/lFwizwnSPB8ruoBs4RQN3ph1k3um6ix5fDZiU+SB0d
hPrSBkbtN2mDZ8DOVphkErSMSv1hUOzph1TUVSv8pdIlnyIgEnaddLRmHXMDyUWKNpk+//1UaLX0
wmZMqrq3zgVw2oL0Sc7aRg/0IAXIiNe5xVTOOcawSm3FGDU2AsWhwVl54lKo4K26WQiHQbcMYIJR
zgV1Xmvcdf+1N/gATOZNqCxu7kiuVhPv34sam3SYYnLVbBP09CyWZexmS7IX4id+xWYC7Hb7WpE9
xVhCtjW9ra7wrcC24QebeGpekH5YaaFuLLYYj68DFCcYKpzyZDFtH2+RYHawpeT2+m5ra2SWZzcP
+VIRIN+lyiaL8aiB/deaAH5NI+4GKkTpQ7QoywPlmmPo0ElU6dlMFogZ1N9RVKmT6uuClK6f2Fx3
iI3HqKzrLAHCzbKd0OjpqahYO/tIpLqUr9RHhHhYK5ZK9Eh+SnHMKXhvqgBgeWfQq4+WMPNL5Que
3HxeJ1WU97J27iH9iy6F7ybJrfJHYh12z/FO3A1TZ2iPTopxkcItJS7nslmGR2Zp7Gs5PWvBTUvM
HrhEWcAGo0niD8RSzd/ZLXlTZjDsxu6qDRI5mfazMIDrageTDQGl31xsW/pINWcK+OLrOcxkTZc2
2iz3IpMVzKUryjnQzSbYrJhCYuYw1PTjTH50hV0+vHVmhe0Nbd/CfLc4nzMl7oGxVXYx6MMzVZ+P
qsTsX+UBHZ+PrdowVjW4EgOFBNhvyLKqm3Y3qCesJWzzUWtI0TAY9uzxkznTmKCmN+AFDlF2baXw
2ENxNcbaSEpxUmCT5LCVjM/GKLsT3u42OK0+gTqXaPEpVmqOvKU8ra+4pqL573KhTUuWh271rYKN
wyrLs2znyBZ3XWJILJ4mqzAXSl7RZ76aW6eRrgvsWz/YichjdILR1yiaElSD/NO8utu2Zpth4oBe
pxDSVjFg5zvTnK/gygV7uo1XpLvZgz7svTcsCPNSnSegaB2deqLk1f7BZKGx+Oz9GXj5udBKlxe+
6hqzZQRSF5A5Pm+5CKvOb1DGCxWud/oYY7hKgrpHlbwXOVznuit4uB/SeFKE5+RuhHXCud5ye8yK
xtRwDSQ2zlcvbXcSdMBojP8VB+VmAhGJbRrmMe70XK9PYPaJrSfL3phqGph1SznG5FIQvJV0rY3a
x4Tvz6I30Mi38F1qjx5SAZzkRtXlmqv2XrNdWkJ27mYcXNMqGAFv4zshvXxhoBsdqZYHhdPKeuc4
cit9CWkZMIrI4D2GHWvwynoPi+ywenMTCtUNvw6RveCyYlw00hXRygr186rdZuzKmFiMONnE1Cwp
mfxtGkWsjTzChqtIYN5hkvqI/64gUOmTAZW4R51cKGa3CBtELImFa8cG4qTd5V3HvLf4BkVU/aZO
aPJ3NepDjs3Rz7CdyLOYdiJWPaDGfez32no30wuLuNRkPJ3olcpND0o4qXKtj+WmQSKk9lN5+orX
XDQSS6OMpK7d942yRkzZ4X3wpnc4M0VyGNjCjmH35neOhg9+irVlGJTy4bUbUEwVvVGP89wuv78F
caCyEl8alFUK4RP3sQDVUmWU8ctwuZ7NfDCSiMvrzbGqrSdDS/hioRI1G5xG9nXQkOHX2ANncdjQ
qeoUKuFJTpsgpp0V9EZJR2EBBE/AFtcmGH6MBa7d2swa4BU0ObOr4OYrLTKTJf2HVgHh9UXUkQuB
4Hqyw0qvgUnR8YUZUfOoAUnyUfF1WnYhkIypL8qpGmDBvdC0ez/DdCSo0gm4OQCWTe6G5798MnlX
62Pm9XDQPfuqW+LouNpHMj3z8m7Lx3ebtMM9nayehYvEcn0Zjpp5gvOejnZwLOHWfZFm/8A/QUyj
Qk63mY6tTbngBT7Jv0LMvTJ8QfxizQcU7vDaAF05R96s3of6ZD74xiPL/PhODJanadqmQDBC0jUr
avkJCP+RU6ArcPAfuV5VapmCFUX0S9ujO0aGSDiEbF8K5t/8IakYk5QS7dUnN3xzuj+QaLA6hFj4
0ygMJf8Au5cM6kGa3TbV1SlRo6tBWKBto/R/M+tygYbkzm4Q53P/l9fa9XROIfkpvX2aJoquaEkF
OI+cCAlDnoU+WL2u1sCg1NT+x/lQVLEE+iBjrtxKZB+xahiyTh+AyXC3xjeb4t6oj17dKv2Kmp4V
QV6CmqNcUnipCTZYuW+aGxNQuCCCAa3Aky8Wz8MM57elKcrxaBSh9AJlLQsFgEt2NmNuCLD2SYQ6
mxnaan9bNAjJ550nHfDuQamVS9ARDRvtTrbjK1yOFxqo4P8Ql4yo3Lol9SvbkIKQEN+97nIf8b8t
O9NwQWXMUkqA0tMYFsVKitV2zMCL9UIPkpbL9urrQyUod+h/fl9nVobr4DUVSM9wdrB2hmIK2QtM
jJCzRsbWqsHoooKC56eIUzNxpqw9ros+dJ9i2GLvKieq+UfbdwHkKAsROEKru0jAX9L5QkI43BNR
4rj2vMdEo3rocvN9MvuSoX7l6q4SzFg2tCofJ173vKeEc9Y7oqH0NhNjGESCqPI/hMHq5m5BrKmY
0rYyx5eJw/OXZ0rvRZs9+8rLzM4BCDpvegjRsV63F1EPZcv0ODeukzpyWwp7mT+pb5doU7CZdCDK
r5UOPYRWvRmkwbTne0Z1/24dPSeBYWNmk/VNEk0xKDZochWo9OGY0YnYP2cCIi7rhRSHblkfakjU
dvaaZ68US4tCAqa1r9bESg+VypxZpqwU8gaTtR+ml0OYs2ASw6wTZPZb50mGNKLUDbgncj/r7SOt
jp1qRTTReKWirAb6L6yqXzSOYul4GEItQZKUTpklZOi0c413i7cvd+LF8Qmhu/fA3zpci3YW+4MQ
AYYBqXcKfgNL9ym5v2NRgSGe1KIv/eR9KNTgFpi9MbHnO/pSKIi7NrXH5lPpZCZkKNM/Sz9rX9N6
Bv7nLwUtHDwE302lGekGU77IrkS6GgICaTXQtUXIWmcL1HtKbQTd7Ow7hGEZTkW+2u6OBjq7xKsY
iNM2XHVD2edaO6t78GPVxkcmuwOpdz8jFLYjff7cePi0xNCwwQqKnHQIDpVOPTWLjJPoKrCSC7Vv
Z6rdYQCM3hT7BGEmd42MtnK8JUVSQroIj2tSMAHuOGN/uww04h6yBr1t1tSpsrZEUBim4xVMLp/l
4AMUA6C1hZfB0LAW5lIZkCH+08XW3fs1B/HycELDRvZi0sWwIIie7HKApMao9SYkvK6fhFBJLdod
7sVKVx7x8u888Pw9nQHSVfLCziX/9obzNZIElR3vfJ8XIWXiCGmAN0z595KLX79nlpGPsraKOP5l
y+7gOJJS95FdpjqhbS02scCv4YqG7/01qYmCeaGlZ/ZjYTFekRKqBa9tQepWNC61N/qY6HPPUPEr
QB70DWAQQifP4NkHTnxMLrWP7RX+OqDZ7T1o8MLviJ+Guk46zqEAmrOo3euaY1cC0hEUEfa8LOR6
JxDaRQiecka+djl4eWOYUlI/mljDWrrfrETeTJWR+7Ze7zwzVKRshKeYSi/SI3v75uU8qzo0aT+Y
3C7Fl6vOM0OTiZ6P8tGAtc5F24if5s2lpsuaFNV95ZcvCXnioMludPEFX/PkOLJSMKWGLYVPn/6r
c98gVRFJOG0KKGCZ6IlszuHGHxs0XYmiKwftQCYQ+0404ywk2yVky0K3nLGnbkle7sA++zU5MunM
sZuhvN9R0P2CnDKaMtgZ7whji9Yd8l4sZKDxJQeEccsyl7ujMyOpBucX9vB5T99zK2VWW2cNDtcI
KqfrmP8WOPG66fwh7T3J+Iy6K5tr/36GklRKuicXBmfctLwcj0ng0Wn18vH8TymqTzMYp4YSEJt8
keAXrBm+riJQHElzRs+K1Q9sSjr9PAQ/K4+OeWpFYuQS5hbfe3znqqzKLO7rDxwo4TkSZfDp+KbN
KPxErDdPmeNwO0jV6ZrHf3MTa6ntW76doZSeOgzG9N+i3PST8ysOq9M3kE6ucu+ibR6J6oOO3+Fl
GVI8razTxcV7EEFKV9xCL3Q2XXfLvnot8ULktTtJIL/M8uFsx8mOLO7GK0hj2LzGTfmxEjpQisiB
ErZZXQ0PieS9JdlrNiaqeufe5EJ2tZBiQuMyVCUXGAev6uRAwpepx0EH0fMFhSbFdW1Mfn7l1yWJ
KCTPacUmLOLcqFlS4zHXe39J1JyIpk7b/QrEaI5CrtMOi6ZvF8OqBABd8kGnLVWuf7azgTO73KNm
Q8kO0XWRBDhaS0ybBmc+40FmU7ifWpGkfN5p20ySj0GILoUusMFOdwcJ/k50zuDPpx1/mPfPGiLm
ncc/B6/wPv7pobR/yFHhxtQQsSxTAlEJrl93RvMS6Bsf6+V7hgQmOMURT6EYrv6IfEysn1rr5F1z
J1npw0MbWVH2YpRUNs0mAi07uzlj/m6ilkfAZmBfmSM4J6GtDCxz4WYNihBjwgmrFAqIcXS4Iq5U
cbOCP/7L5rKqv5GlncAa1tpXyfQxxKvycBq9jFl/0Ds8nkjP6eWIY+s71D5zzbt8rDGEu6MCd+U/
03DjBL1ehjTGdJ9C2lCY4x+11TrI4Kdp/sR+MTdKpdDOx29mEPCn7g2XosfXLuAOl1MzuV0iPkKY
Z+q+B+Syvgy0Tmuxg0qfklvN3bnw2/ujIIYDpMYCoZFfxNoFOFjzfucsRbBkNl8D+znTS1J6XEqe
O9231wOUOa2RP1LxE0pNsV751JOQdOqyx5vAw4G9YqIleQ4RP4GliikQDYebe3PU8l3t69zQe40d
UPiqvleSG6G8kJygo2Lpe/Me8Y1Ci4z9ZRha/YSv/ItcXwasTKFpyF41NNFRvkMdXln6fExgm89N
UYeT+imaep5caI34FdjId7q7pXvl2HC8du1Nu7BtFRd+ptRG4UL6ZSQCwvpjw9E9uQ71K3u5gQDj
kX2woW1DRT07haYdKtYYD0sSBcEArzbVSXksq6CrQUvCZ5E6H8MqNFBSfcPQngaJCFELw8l5VCTc
wTWMgLdZeaHMju+Z6nJPvUXo5dbgUECd5w0bOTdKayvFT9dMe0DEYIv+uD9DoMoGwG7uIoaSYMuI
rgVHWVnXf25h2pvEmonz+YJe+xEncYiqk7Ehio4ERAcNi6PLXhoyObWBfMFIAXc7AZrhdleL4A7L
lTRCuQiva0ifUVYZkh80s3ZUu+Gv6GPUMcWshGr80IPhn+Kph9QDaFLEN4gLYpQ3PMdiLd0XM8MK
sCpFxewVRVgGLw1Z4n6muHjFcS3x2x8n6ru9FlWmBK6Nr99zsCM7k3OuRLFmBqgbG1uoDiGYrmkZ
zBh6c85AsgPBTNydJzU0XxZS1A+7Vw0dQ3WZ9RMuFI5gFOmK4c9CgbFwLj3XM55ZiPa0C8M6uv5U
IEhd8SbnZmsfuypi07R9I5U0Vrx4oxe/GRx1uj7yClaJ9MM+kPA39M+zCLgWDZqmg0mFcM7YDdPT
gSuhgxpXcc+tY0FfeLjHzks3DfvDy9YhJvyrjENpDcEE2Sy93LYPFx3QO/0zDKwt/rei496IpVi/
2N6irMbHjipixvQO+y2mBvaJZ06Ck080BBPkZh/qIbD8C0vy8pvBP6/fpFwtjW/LKtoysbfCIdXf
/HNzUwh604Mbm7iER46lvzp+d18EThiNlCc1LrR9TFwtjWSxWhOCtwNW284lLKoyvfHPDICHZOuG
yhRPx1cdtEzpXaz+MGQF+GlwQgz8PxB5XZpXl5t0LjD45Xwo/+Li2PX8rJF+2u5LWupgSetBn/Hv
9/vDkaFeWh8mL6Z+JhIvHTYW6RR0/znbol19quxv17YCx2cWCxSjERKD/oezivXgKVPtAJlvRq9s
dvEY6MOztkdv8V5Mn6BWNrrgOjOf7yK4wc7KZcJHRVS+bIm01KUxgEosyS++foygHlshF6BrLWNi
7HW8RuHLDfkV1ZjDFm6FQLKLXh5/IAgnG9vXlk31EyhEY/p0dlVEojs6yNek5LDQ0n0TezPH68g8
P95V0OLVyhLn85CwMgjum+PXYmrYGdaSh9qd978ODl6ZM3siouHVQXr88scpfNtjIeRW3uASI5tP
EhoQdfNuzTy70iTtGjnbUrBJVdw27rPSyD2d5fYFtieMLt34YM6pXjp8uLjbGC9f61b36ilXReSC
sjoRs3bMqRiaKtQVQHbrPabIvM/YuGbdrEjuC2g9tGz9UNbB8Vgiugwwlwnmwcufbu6h4olRN4WN
dG5QHZd1vv3Bp7Q7CKReJiNd8M2qBtxLtlkC/ywitv7/8260fuv5dLXztIQTqWT/8szQN8yGfQSB
E+zTeDPo6UZ8QPqiZZoueq0HsYVM8aRujqWN87r7I/joNs6HEYnnrqHxwvf3RsHvvvqBuWHdAqeq
6LIhPL6rhuBFj4sd6lL1Zo6m5N0K+56NIYd2cIxkBv0Qe49m3hPkqFaDRa4YZNKL/A/wNweUUejd
3TBtnHa7bqSf5xoNS5ePawJakqS652tQz9otKFH3wzjQuDvBeGTqWwRFnEiX+QWIcddpkRCw2RjY
WrRtmoQI8+D/0zvnGsTmBeSrfdMTTCK43B/xr75AQXGPcyboB6MG7omTsrqbEEuW0LBliAqrXu2E
L2ejoSBu6A00nmGehh7vJAA3tIHMskMYIftcRdzuD1p/l+5gM9PkOwV4sipODKpAD9j/7TlrKiuh
BG7+JnrQkmgpNTWgQY0pgq3yjGkDniOVbFdKiC7xpInP3kCB8RWwQmqb3TkbpHwYrTGnwhy5/qRo
niV9/iLmt8mmsvEc/BIfbytsDnLaeLtgB90fXvw1k0xb4m2BIiY8lnrIauai0Fqhsktrx9bFuonW
t7/XzubLfRgM8pFhfySeaxCy7qx5bLLmUNuifQkQHG3TQjKDHDhkFfaI0m5p+oxBTWNxjOjRIZ6v
L5B9aE1GSrrsg4/EVwCFJ6nKhAJRr1lcsNhkN+reouONK0trq2nLWwcdFNzW2wbyNY17F+xOBYOR
mQKq87uR069Tz7pLTu3X17s0IOcfhCXF2reB0FSpi/nBDiGrqKVXYzYkiqrYzktkl8ICbExTd1gU
xHnvRJwGSd1hlsgmnKCCov/mgBTc4Stwo0t2CtOoy4MvAsXN/4ieb9lWWdxs3XWZF3J4geSZ/4tQ
wSeG4dLd7ADp20PcQQyB2oyG8Zn+onIM4vfDiyaTM1/iXpRgUzT25YdFhsylzyV32NVOxg13hSIH
ghB42eNETGirQbgdI6T8KkZsFSjjf7VAmuizSPP2Bpuk8g0anqY+hlRHLHawmEsM/8PkrMr3cH5a
wJnv1vq+cfi3wEDLIb6fZERyiClXU7VCHIdv6GBupfluESVNCqP7chAIHOqXvrK+ENXGaC+ejgYY
cPXs7/BOa3nZsp5RrXPwmONYzmlgluwKERZTYn60ywFzfaKs7LOM4DxMV2xl3IgDzXKdJuscstop
Y2t1deMxLZPxxUb9ooGyXmc5gVi+xNFldcfpIHqk19OnVYv1hOIgVF7Wx/XtrCct/KZ9VwzEOKrH
QdKnFeVcCdbj3HPkB63q8YRv1WekLGYkekxfjZzIeQQgJXrUPFYY3oMHGQC4tCwKwq8IDv+NZyBT
+7XNTr3wQgWUO0CzMvzoSWOkRHAw9D2x57gGpudKRxmYFyWYReMy10nkmWJQdOn8v/e5d3q99YEJ
4woM3Fuczvd2rJKE3wXCccMUfRoU6fxZz7igQ9ZVGtyhz8ymZFm+Kqmz/sjtTv8HVFPuqlQZBAX1
bPwGNqUCPkkwdxs9A7hpRg52/CTTSgxkPylveWnjv90pUnW9Z4pvZF2W2OwuDU311rpXN0/OEJOY
rEQB8rgLPtndW8txMUg2E6VjkLlR+zNgC7foI1ndxq3KGSCHXaeQ3Phqyg4R9FQ74cclParZMtze
kTMhJQeWhxdnwfKXsU9YaTGEn3YVEjANZhx6o4Gfm1uv+6HhEj8UTFQwHDly7sY1qzcluahm2dwU
BKVcnuvc1sFNfAzRGYMzu32fnLt3+LXHHq625gdqa/V7j0eCbvEKEPgAnhyyOv6UtwqsAECpMR1A
E9JO7mVXvyPEvDkHej/o4rvmf+FEV2JTP6989rJ9TbQurbKbqs5e0Qb0P+ZkgbSJwLlCoB2sDWoW
5rs/6NCHeKYxGj4Z7GsgbQIEKMgg7p4jth5lZiHnKHIlOwdd+aND2mjCCYj342Z67gozrbyJ56AX
PEVeD8+031MOK9VWPTNK3XX19fwIbDVM+40TD5/2lCEfXx1wSTtBTN7ifoAXgyWPeP9BapkzoErG
X+H2oUdSB7/3iH5pJrkxN338UiMP1t7tbAd61da05wOUmvDIKBApgCFXe3mJHlNzMviV6VcKlpkO
rGTLJN+DGm9vAEpM0sqAIemyWhYJe9p4ZcIzlbIS9g3GzZlYm9A+MfJHkggtMKbVrWPIQLhiN+jv
c+sY6sUpNk3eFUIX8JJ8Kubn3kYjXc8EQPJO8iMFK2gseXwRj6zhwxHj2zmHF3fQQX9bTPblID+T
a1KhwZp1zLx4cJ8mbANGo5Rdi4dP2IOmLeXEdOpVMPRh/BzW62Bqu/XOenYpi1EOmN85oCZnkmr3
ng30UkV0jv1yAJcrEyKcwhZVwKlky/BgQoIXErJxsKwbmsEdNtIJn8sx8Y/Ih7GJTgBYHpNiV3MY
JwdQP1Cto7DOJr52dIzWDpsYf3hwP40dcUlT67UPlAE4kQ9vEjgy7ZSAZ0uvAZKnnV5b4gqM9ck6
KNeG/oTizND3hiC5od/gaYoDoFAhAdwaGY7wg1cyNmjwSvp87cEiOzG8PGndQDnN5f+MHE18diwp
0YUuHtb9kByyTrhqdXMhxYM6aukxhi1J4anQmualAYrEczONImJW5MrTf/u2OznWRRqlV21PtqyH
eZJ1Ig6b166kqEiJ+YvS+rOATgIo+2XHq/PcLhQw3+1DYKh/+mlYY/J8HRDDqtB93bH/GZfhF3wj
vQhhAFyncehj9R4+CzopoZyW+kqBNZkkfQivODVT2a61etzicMwbREl0vzwjUsLm2vzdBEHbyHdW
93zdxsK7+s49CPBrho7+IQutD7j9MLaDRP5eJS7c1wR+qCdYsXUPtKhX0pIxXPO8dwGI9XmLBunn
GkuQCMW3axgxUqWt/Dcz9ZnLFISrJPAdjpzUH9VII3vcGFCGhx6KUwhtJnRl/scHFT6EdzdGugN3
uJLC1Wwdzpi/jiYJrP3I5BI8VxiLEvM47jynW/SEwzEOq8tVGLzGoZ42r14qcZiHbYK/4eit0bGY
hyPD2lUN7RaUWQxFuZ6ICKYXnol3a8zUSmROtE1XvgNmNZrpbgO7I3YkZxopwlMH8kTjHRHVIuag
uldQsW3bu/Gx5nYsfW5H97EXHGkZH9Pt9Hur3U+2QPvGfbMlG09IVu+oTI+NtAWSdcrC5LM0JJ1m
6VGPQC+J0k4vgNMD2Wr4DfL8cLLxJT7gkcJXIPfN9nzt2KorVDRpqO+KtvJMOlnq6VutwWxFp4+T
N0iJXDldPgyCsyHWvFQ88evIotdDFYsWXmLN43rLwZK64r7PX6+xd/VNPSrWxylDUriQEzJ4RfYu
j2hFwaK9MSPkRpOmVKZ19njc5tP36d/ujYXBWhBdTSUj5xFu0lOSwtvw80N3/NsRlJP6VDfRw35N
YpkfjtQj5U3XDMsNVGc5qOFGBLPDoAPogDoO44VV+kus60anmXw+2ujoFr65097mWZt4DdxUotcn
VddrVMrDG3SslJq6zuWm9V5KdvVAn9Isn5AzZ512S5KlxKkIxUID1O4ldaUgtV5HeAg53g9Dyfrf
U8NsEXr07xg9GZsCco91L4Yi1hbDhzuj4bYT7dM/ERDBbt/UYsn3IY92yZj1Ip9MLSeM5KiilZHz
tn7zYnf2znMejbE8Gua3GYCdmAtac4ZsneDplT+a6Pj2op0ItsLznwNKAkxxvazKxcgqkF788jqX
YDx5ZRyd+3qX4goui+bDFby8ynifm5QUwpAiPG24hugrsI5g+NHlYa2/8E8mDxMwFRo173j7OFX+
VcqeBZivNpy2t8xuNEothhlvSCQXvMpcZwBZzXOpohh/l275W1e21OqPpOKTA8CCX8RGj9YFOJqG
lxoojqWQQRAfg55D058/hjKRdiWZfWMzjDrqWe7CNi6pwiWVoIR2Gcgr/E4HMvjRkqCPNNVukcLG
50t7EuSh72rmPNs43I7jiH/9QWgcXdmzEZcTh4ZThylmbfI2okN6fuzvfN1u4mMupL4xPKyp+uBY
HiWvMeUqv7RCsWGSAjPVX/hsJ352jXRFY1LbMzmOHeJ/9W3aOJZfQQnHuUUH6XRuFRjWCwc1HeN2
woN8BK3jkCxWaV2cglAiJbhKSSEEwAjx0UfpL9K4Dx7Clgbv1qYB0Ahb0//1FYvzceuyrylq/yKR
DgBs5PUnFZ2x5fhCIpYuwG1hx4RyO4+CxiZPMzGoQDsXz+sebUvMEJ8WfGBdxzaTYXl1NKUD2MOc
yOhSk4OZoz2YnmwmyXxObCleiO42BJmiSCFhxfzk7iYqgSSM1b2ICh85UxtTNbzgf8Ov1gRSbyvR
G3R6LJjCX0W4owIymbalN6FB4AT2J60rjvb8vyIW9xwD6CoowWquggVZO/QJaEV2e1+6R/nLFnpo
YsZ8TDyJS0bZJMHejFZuJoU80+Pt7tJSxKdRBVrdinT4OVPbICKBJkrqs6RB7AR8TztBht6ni8Xw
ktUQ6dooBYvo05LGamhKpc0NcBDL7v9foakSuxXBaIIRhBdjpqRMNcJGigALkYl/qt3m8ZtGvgYA
zoTxk44oEjODtQ+tPK462na/Z4Kv/Zshe15iI74bKdd6V2fj/UXrMA8+FX+GQN9tAbgUkDghLSk3
IMv6C1DdDQ45UoazyqFDH2gVROdda/gZ3aoDOSs7kFq5txqp14bGmZJwb9MipeD71LDMbW74PJ0M
d4O2fVI+I7Sr1ww1/rVgWDzIWrbg5LKJVblM+BMhVxPKRqTqHdm7l0bNnaKyFN6vKLr5tvKnFVQh
6BdRJE/zvbatVLEsoXU+JzkCuP1waATq4T8DkXTRih4Nlujx5mkpqAdpaGqXk5LeuIiyJHmnrXvM
O2nqiSQF9xerVVAOXl4PFCKQU0J1+5KM+mp+ge1byzv7Df7b4tUMKOhsqjWNflN5VrMLOOsmJd4s
Otl6HqgNIkSJoB/WfBOIrJSt8C5E+SnaFYPNwB/BA0OFTzfuEXEg78P0iKd/9LTOPt5U5h+PjrLL
tTAqZ/WpnPDx5qGncUsz5rsHcUY7zsWHRWdmdV0JWIpepj4ZfjG3HnLQcRXoPTZ5zx1KlJSEE8ml
uoT1c6d1/bhFJFGGNjZVJOqJiHhvHT4s4vum64sdfJGOH8Dso9NMBZnd2EluySj0U6e5AX4TRN4x
EX/BdD/7151y/JmhSwULtpmRaYusyr7kei+rnMk4xe0DnINBL+qn+uq5Dw0eob9vmjZ0wq5inZYq
q2PpcMG5ywDuNmiDc8FMxMx87jbrQ4RoCPfxEnJUWP1nP4eF++zuMrbqYX6ydzPONJRPyTfj6uul
FVALuTUU28yzBdftSE15q6/SgnU25SoHgZuBsdeX4qt3Frmmf8HFWjDTJumLITkIfotPUkorq62g
TNc1VPuQpTahDabRP6kybbd0XV9zq286gATN3fM4ZAQmz8SW3/omIxnTiQ01Mcrq7s4p7Ah376Mx
GQQvKH4FZHIIUNim4ht+KEsOnWwbtoZGI3qWa6JdO6g1ISQhnZF7i2IX8f+VhKg+njCpkQK9iupD
fqDt2Q8euvL7RCiUuVEqBmJ8DlcR3cu/CK5LL5/oWTmX6kJQ2w3VJFOahVFWRn8MNcVFgerBgikz
yJsZzQ2oWxB0kPNWDv/jnKJTd2WLFhzzCAzq8S+uZoV2LvnJsRm0qxnJo88agDQh5gFicql6d9Jh
m+cpvrmEsnQ3CTLgNREBmffWuuDARlbslTKn48mTNTgMng4SwBcSRuM9em9HIQNs7rB9zHnzQeHz
B7fYgCVTdRpRk+v6G07gZ4BtjDJnGdX0R8cViyM4L8+FiYj5BsF08hLpNjDo07sPLPTvWTvgtu+q
MbWzsz70dTSqFex3Euey/hmaPe5xPFdAbz0zdC88yqsOn3DntKoWzh8Y5IGeDo9cAcYGNoW3bUX7
lmZPI7iocPtGktZqUKBpMdeZBrQDwBNMT9Hf+FNVjqzOcuGYQpB21vOfPW/+KkCQ13fbCbsffUZX
aUjsFQaWGzoQvAkTFcvG/6+ckXU4txAO8xKtasjZHeYpZV+BPFenU4Gb70p6VrMN9H2iPgtFgfLn
+zW4jT4jSc/mtIQw5PrGuSrWaP4SRSx678E5v7Q3k+pbOtMLxANCYL95aVBBjffqEJXtEXpH+PVA
8hXBlY8xHJvTa+Fu8+a7CgMVhv+e3w3NU/Yikq7gKwb8xug+39da5iUiwjFlJSuW2Xfeut+gmIBj
nelkjAfcOoCOQ4rmmtAW2v+rBl7NETb26C9XNWQ9+qbhJR+pVWGjenupO6SXBilCZv9KQ8VNPogu
ETtXgNuoLaGlo4x1Qapn9kokGUG3UtSxeoIKMsiQ7Ex6uWzm6f5v8wb9+ARYDe735L1Roa1cLgWU
7rXn629Zbw8N8a45eZKPEaCq4qPGjtczkdCmvPv4WtgEGemWJnUj1ZAyDIQT9op6YEOsqizaWxHW
ve2cuPCw0LH3mq68lAr8GSLWDMt6oNL4dvFr/7FUpk1MaIXuy+DnCkEG93CUQ9F6zXMcAsTOWf7P
8++j0OaNcxxzL/zpenCPHim4hkarBAauytCaCYs3qryiRD6rP5QxnMedjHCVpW3InTbTpVZvbF8o
QHF9GDkCQMVBII0dMKEZ+22VXxN8sbUAvD/MOGeXgsw/eqPp1G1LMvfciqwbDNvD6NLHQFoJIUXu
cilfycrcU2b+bCqlFc8G2P7VfyA4aM5Pewzu2cioDO1JkrmL/E7kf5FUMMhQW4KPE9GgenO966Lm
/eC55fZlbykDNIyp5WoXZn29vh9Nuv+IARLqWlFw2RecR93Cx5umKagCDVJkPX5qDLcNonl3j0+q
3INEjw4rcPVDc7sPLUwTUXz9JmkcfR+VRP+PFKsvJDlBxZ7SwTfJUM2ZFoMNLuuJ4mxcUpHzMYw7
jAhxY2DtjvAjI66CRn6N0fzxa6NpsgrqDxNdgeuUZP5kOtP9M47Ot8qHOH/T+eoV3SVYDBz4gcn5
NynQ0B6jLerdO88hQMFbbP8DTznxJfqvHfNvD27w7oyWh+b4+5fkMXvBfsjfigcJgbGfQVtne8+V
eQSjJFAyAivpUTA6GD/xrK8G32iRG5LLgKfyv4/UzdiCBSaRNF/S/t7CBaQvhwWn8t/xn7GKFGW1
32g6kNn9SNQcbyjVBT3ev9TlgRZudEeseRJGtLcY7jkMBDsjF01opBVfuYHk3uXYoX2j5ppVvJNI
1Acej4zBAlOF8Tq/SowtM8bf07eNmNCP7foNMwrdsyIYOBkDkkVWEuFL2yvXX5FzZ/RllZej95v6
ZIUZhxoNac894fNqGiedQqcQWWNL+Zt6TNRI3hhjd+L4fszyLmAR1LVV64EKVhKY2UAe6ftkxlCb
BJ1DxD8Br828O+MF2g1M6/lOhrz58yZXaOdB7TMODLIllXmJ+DBxC8GgIs1YLfKOIIjImQR/2/cG
+wDc/tnLnEuVtLspsDmFhX6wo7X9t2gPLiRr9PjpEej5Oi7CY4YudcAINehJw/A4TumcKysailzX
CJaHTTbYlrNP+1fVu9bjJytGx+XhJmqvZ0k+yd1ZocgDdnJEt07OmUd4MDAB2pnBfCU5DHfibIq/
xGE7HQz5N7ahWmSRENG9Qnj9QOY/oomeZjWhqwUvNpR8rUrBhAsJqIMJOk2e69XGmH4ZF+R+0KQI
XpLhQRygWm5wpYUmiSWmfgmdsgyMAnN6BC1VskZI8BjGPB/L0dwH9n5/tPX1e51PKt08ZpaACR5d
rooo3SmbARQa2yRVmrjfFawVaKadlYIP/bF9GPcaUenBrG5kuo36z5ysF6+DTnBmlVuVmAwMLLNQ
L+1UNsMcc0feeLlALvLWZCiVdZYB3/QI/yegnQUhk81kQkIsYEZtWNDJopzeaSxUYS5ElFJKTjck
UnWs0SFS4zDCqPfNWfk6u/7vd+39NY8UwYDHbcgX4KZtqoe6mzdounsL7LtcQEhrT/HibqVwZidV
7IK5gnyQSPuxt2FCoW3MqjKTx3yLY7cZlisaG9rYiNgZfy4NwbGPD+wZ5qQdd4JgfIVXYjg63yCv
DWJwFvWvYLOClouVpsV4vmaYASkACW/kAbAcWHFIxaPtnydg42FSawsNBaobHE+I5mxoYhpIPPvL
XxvLIg4apmcE/mgiblsXyE+52ZZmwIPxz0hMnD7ocPQfrbewkHIkN6BVaCqBUtL5y5Yfomh4bNj6
YgBgQOLwAoLrlFRrDEYsHOxRVhlOySfIWY26Y/oeA4gF1E7MJxqXlLPdgRe/SFT5byk4bLZvrsdu
VxwZMVLXvDyQYz7u0W+izfj5erOwlZM6s6/+GCiCtc8lulPhOoWOh83F4OCqEgE6SsCzLAtXVOLW
s4lyTV4dB7uxAv8oFxMYlP8Ziguv+AA+qMYCD1p0IxNp4ZhYG1YzRX/eGEAhlHgWaQi2y/k2ozlX
s8To/iY4AxERDS5LcBAXOon+g5IV+VRKdCWhG+cwqTj4Ctcje6hBcltDX546LtrNcYfaJPzycRqb
8PNUkHfiqJzb1MSNzAmo7gha7hBt+pCy2zeuOPE/BsuqYYmWkKmAnweMz8rFTePwgifAvfALC6b2
Qh7fRcRbR+kxp0jcn6m5amlJ1FDMaDk2hMq+hPyrbIWn1sHLxQ1JAPOlES+OJ8je43QveqmoNwzz
CUNkCIKT9CGzQ1DDjYG3Xqj+Y+50qirn8DzHVIUBcdRrZZir0964QHHeTp2JVgOlUGcTTJFf9tOh
WW3KKFgXsN9y28IDWwVMWYfMpwaFgc36pKyxjU6OzuaNSaA8S9Jhs1duEWGVwKRIYUfdKutgZ1J8
8w5CW0/Nbu5pnQkOt6zfGpE7r0+/Xg9KCRbbDf/8mGK8s6Wile5KCf+XzRG1myN5zmF/rNyd3xrb
s7B8SaeNboZwsKb9uub5+FvFHraDrjnihSCBHGjkMd79jiZTU1LEXPU5kZGi6kZ6K+ngwDQYlZ8T
3+oFebSXBQ6RNtz6plKh8vpPzCjY+MYbt2O74Xpn3qEe3XRl9RKAtvcEOU7O3tRXA0BNHOyfVdjI
/ciHF13JKm0DL/TT1q2iAqoGPOzXlty7gOVTJYntdtiCKW287bCmTKbIaL+q43/MqPaZp2G9IwT4
ZOyDi7+eCVk8/fWjN9uo546utzCjcSX3xBMp7wErjfsuBpq85yeXdQE4ynuSzAQ87UQRM65V3MCu
11NFvOavcFf5u7uXbiJCpaNoe6ufqWEO0ZdxUBAHRfLTK7JeQweCQ0jB/apAdyDL8oxgsXfQbLYR
u7Nc6MxUa4yhGJGpnGx9jGTa1sDNy+6QDMiPuNJAgK5y6keFhGrgiRz37YiFB89n2dUWP2kLYLg1
XeXxP/d7EtqIw7kMyLU9A3UXVcLswoLB/mQzS1laTqVGiZ/6HvmedtJCJ1PBDVnqTp1qTk9qZa5G
s5Mrama/FSQ9lnEyrV5xPXgRC/hCkrYcxgNRW3q/d+6Q1Jptw8q86tpU0dM307sXMD2r7Lr9uM5p
GEKjdgC1fRrqjCvIgD3K32DfX+oeF8uWLtZojjlFraR3S4DVSW2VDRU9O/A+nS2/0G5c9TYfNbO+
flLXuVcwxOesyPePzmIycAnT+lvWSxCqQhTljPaRh1AYrT+SvvtJF9nenBkSQvo4bAbLNKkiRkGw
KKgommdPJ8qUflXVvkJaTCIdLgjxkDIROdAMwWRllfuCscDilz0lVWmnMVzmIyHv2R/53XgRl6Hl
6JU5y7kILrDfE7YjLZmUyIutQ0EH4ZxND+sirOHPusUHtnUjoXH0sDB8XcFpzTDD0wsNXe4o5NIl
5ggrbTQRFnAQoH/tMoMB3o69sAFkZNjI9cB5feElK5OmS7kmyx/ed2JypFFZG9kBvFiY+eFgRIbL
DWJ0EmlHhzSJLedfxi1bwuU4eJImUitw69e6VNMXUsQFkJxxmBfVvU9iPMs67OaaQMHUypn8GbuL
dYQ7a9dAeObwP8EMgMsgymFN9Ul2jDdgBwETt/qrGQubpyxtC5lhS96RgIdTbkVuJv48cY2sSnRl
cxCz2pR+KndIuopzP55h+8sn1HnFKViXrVgbAaWF+AErG3I063ZSl4CClH4Lnk1cWf141NzNKSNx
vn/b5AD1m98sdUj5FD73UvafawLApKp7r2pW7jBRgp9wizgaSAbsphMtgGOFIfw9vvpaywCqPf6h
z2FQNhvILh+F/t44eOhWDg2JUaF3I864v6LeQAdidRTesUf3Mcbly/oSke9lYqDnvycD+e7rSZAP
lUyk5Aqg9/oT98XbYfGYN4aExmyOFtFYP3WWuUSmJxeQa0cSaCSupjpdWrZGa2WpoKoZ/6lxO7Oh
jy6yqOKUnU7djX++FdM6HU1JH/8PMbRoiTaIixpXxb65K6+l+hvba9kA9R0kiYbFuUm2SJ0eUjcl
7hiKw5UX8sjzTpHP9Lv4n+bzjL2+U0uOa9kfMw5SLm3+RjVi3XXyN5fuWudkIPH0yC2dx+fWtdSW
orTEm5TMHjQmkflTBlHtbgd78rAU7siHWlo1/bxLrRSbKcBsnPWLAxg36SH4BQFSk+hH2QhLcN4y
sbNvM/9sHSIYAw16TqpoQXBqsKCyqLkk7ASt/79c5xtAI1FNes8Yo4N8gmOS/WT/HyiS+EiZAKfn
B1lcLeMef9WXHTdRpl9j8UNw9v5FBVKKx/PV4kM689TeUehavZTlgp+1aw1kE7u4nZr+bweW56XM
nygW/ZaEsZx2OPHEWPdxF4aujCcrOcpTj4/yNf09h/up28kl7Akv9/5q79dUJ6mMClH6HyZ0CJE/
QypEBCfEQxT/rmp+CxJ7tZxzy0VP0dwvsN/bGz2HOCkmZVSFHN5eLB4MTxBUz7IzCRElh5lN3Csg
2ea9o5tVY3u/l4rD8BZni7B+JOZ3tP6fa+lIAL7E6GLjZPz8NqPIKF8ZiDXpJQrU3xHsV3j5ZLjB
nZ4KuiJzmirAB43nwwnVIPHHETAhz7CFSdWtW6Fo/12nskrpqV82fjuT+1ok0RP32fOj92S9lL7j
RwgMzphKUBRfFMZnJ6u43bUdqDawODqSb3y17QwWbQtkXMFCQk/iPAGczv3v6Jr3pqFDvqfEGoYw
BStvkH8btMPWfnftVH9AvCOw/gWzFeZGO0TvoRFn4jqdtqHYi449RvHXJh1hSK4Dp0/0cMf6nAG/
NsO02Z/ttLAVOY8vLxMYInmn+AiffUpIHc01AW+TeJ5ySV8Jl1iXE/vnwGg0Tkaf8gARqqeQqD71
WGSCk9X1RCZL06aQrJFf9JaUbpL288lWIMIO/X4Tqxdy374JlFxICMJewPtUlAO/tTAIA5KmckXm
xnOAhSnNiXZyzuk7Qu/2Gl+2D0U+hzmTpFgFgPLjX52kG9avWBgzGjUjKslZFkzOnp3UU/Qa0IFt
x3aag/tWQOCDQxtKBgaJW0m6fbAc5dxAbnPbrPqWZ3hE0h+ZgcQbkAYqGu7Y6moRflJe52BvrrvE
59OGvMmYbRTBVs/YAe4j/WYmLPjxDmRDKoowKI/g7XPCOeVwoiqdSxlSA+2mgipsYKEBw5vM3xlq
TXNjaAiJM0wgDwM/pOjWe5KWICS3H9lBakQ0zWK8K7OjfmZg0IQXGpfjsHLsofTD18T2/5L7q9LJ
TueC15TUkJsEX3b0zPA5hXADU8N5pv0r1NefEPk9RYEJpAxPICyAm7/uAa12w/DQc8IXKqDmwocB
Nzh7+nd4dYm4ayrdRRG1b3k35/UdKoLQ/XBh6KcNFQPb97SNnO9Ihf0Nk87Em5yg3JwtiWhh4pL8
ixS49TmYo9qQr2eOf5GzGzS5pLKe1IxqutbZq4KSdVYRArNttjjqd5F/F4SjqxulL5hUBE7cJhGy
ZShJt1insil33mX20gMdx5QyDRw68Bn+AToN7tNvkh7xluKwWO1yii87CKDl3+3XAjwryofOJREh
cbtcczRwZsP1DijOvvoedWvePWwI6hjWhinKFLAOSOZluV8GKufIsDwpgkOgmt4vAHMFBgP88d3x
e3TFoke0DIhN9N182M/8RvftBZnYzkwS7N85akU/uf7c34S9T75vDORfXSAhE3bZ/Z3AHZ6kopIs
p8nmMHctP9Fq5/BglLP9KyxTcl/r9S4FWSATCanrAUFFyXBJfrMoc3pgGIpAQLBnL7nwVHwprqVL
NZmyz3e+xgdqa3qZDrERPbJAcPGXaGfEkGrMdZ+/yHcXo2iYSd9C/ga/DlCCptMJv/iY3oFeeKOd
PNCKUJo69qrsTKBG82xqGML3aSdbUpA5Om7wOd/Xv1WZgHsGP3tpACRp5dI3BKN/Fi+vpho6WVqZ
52ofP/PPiv9ySn1iMJdgWZy/uFbTsi6PyqCu0ZNprt6NuKu2tGTWaZuM0L0/pMwyxr8mi3liCcUb
y88yJ621GnnE7WUsQk3r59njVPesiDUObbP/SzgLS//O8JlARCmbftAZlhceV3kT+uvA+F0TAOuh
M7Jg73GNAwXS6m2u+nqb18gJkcMBR8s0732mcurkxl5loltKZMtcGu6M9HnvSF1pgjYi0PNmBuDn
rWEabX81FfmlLvDgp2KQobIrBY7x4H2NCLRJgTxrcpFvFX97vW4NxdtXZ0vroyWWJOn0ty1wrafG
rDBWQ/qOL2EipV3J8G28apGMkjn2jOul62xSK34eaoWCS66gxoq/UEOKoR7aoRDoECgo92a+1O1w
9JGyJgCZ8OYUSw9MsJb1hIriD7NbrRT2Sk9X7BEOogKwhjSNPypoeaVuBFxlPJjyRmsmELdZ5ZuS
09RB2kO5AVeUFQbd7ppifTa2H6yrnoAZE4QN5u+Qw7bohGfXx4NDzQl6m6iPcKPwW/mvhdBFguR1
bgCL7+LulXFszbyy6OBc3YjXK+ZGIT6SWT0OGeBggjP/52rylNRk7lJHtYLPEAKl7oAjj7Z0Dn8m
JfIzxx1gNYkvnoYOUAaqrTr3452ZqzkGXoBU90s+qLZfllujJ+cpDY0Ex/ghIUaB45cxd3fPzytS
BpBbF8y0jNv0YXgWHIO4GRQYmOIZuO2B5tJP7zq54tdjCXKvpn9s7l4YL8i5raY3wDJTvleGRuMN
SsItb/C1Lqd/Qgw6E561IomAgsMDZn8H7EHYYtNZGEet+XMTPZqTQlV5p3Q6novuicP7vWKyWy6+
F5HCzCy4F+WPg4LVQl88xzZizIYlAGMh1542jMiHzLUDB3U18Ox5ZsGCVQsERjezs83UilfSMeYc
JXpaS1UZsbHmt5VwS7We5hWkRQps3gWD6XGDbqYDJoSy4YPIiCt5BaFmdxNDheydcpp2F5tvaXaQ
VVcBhxRe5f2d9bQTPP4TE2tsoWfyATiKrISpuASiIqzJ6DbQzrIx8Ghd9iAnF7svwyPDv1hi6MNi
UjdQVFfNknEsT5gUjv8w8Yi7HUt3sx84quu/khoEPnGhW8V9YdB0Mngul+Ca7HusxQKHjOh6sHlp
WcmLmhsuWvMmvdJWiUp998fP7G3CtECqAz8FAOVptibv540kHkOGyu/eF6352mtDkQM2Jc5iR3fO
+gNdzzkaw3+6MNTNRHiVF8IstpmHkQAjKulFyDdp6X+EROPR8UxHbGMuRAG/2XLm9fyCmLT0BaWn
MKKsvrzhAga/ogLqcz25WPYHSSWIUUxOOkyFndKSjCNbamwC5y+iKY/ITWgme19Gw4GFZrPjXNJC
3zqmKDC846MOR1OohDPWjdApywkpBRKNyKWuCM60awDB5cDC/PS+/c+7kwbU6I+j2T7ILVocdkKn
xGlJim73cHZFeFxDnGVjHvvDapbLZs9mMy7tLoGDQMzs6XHecAg4rE8ZC0QzVHiiUvvW7Mm/omTl
siKEVsgioPvruwwirs2Yx2zh1zxuVdxP4zKYiNTsoPPd/0ncDHJU1X1hBU0CTZllNmmjKt+yitng
sdpDsQuB9H6rjwtUx/o8opT6PnKOwFYO0QzQs4C+MoGOcvcQG6fOTcDnm/bwPTFyV/aOAih352Ma
sAv0XEJXH6bu9HHibdIx0AJViOu8Bn3nlEpZ0NJNg322uEgNlguRKylESTlxo7I1Q7Hp+JY9TFeB
eXCz+F0BO5qxK6a7707tu3tERDlkk+36pGotRjD4zJRlTMSRXqnQrUD7+NQQLM0vWijY68ngVZEq
ll7jpAY7i0qB8Qw2BIDq/v/pvTA3C0KMUgzJqe8iPasXHQCaAcXUpyZwjjDqtQVoX4wB47g6ZV/y
eStFM/5ZQRzrPfC/k8Sl2Qp5U437C24DCXqzsjM/BBQXD7BJhoNHJ/X3Wk3K8OUR0TPwUCwIOR+d
7sKn7O0H6ERTxozHaG/erqhpi0KvZrgjRMBNxj68fnAZ0BdNUkjBCenulCffJPcYEycmAqDL1wwO
Clzh8ehPc1ecJbBGYPHDkjCdJHXJtegEACRjAiBXriZEuPzzZxLie/6j8mBJlFM8CfXpnAJe4NvU
eU1LqNUrLvEJSt8kEdVhaY6+HNZkGlhFlqWxvdEynN4nXvs2O/X2VgzC0Gy4U1bcqxgw/80nY7+3
kG02xeg6rIMh1eLRU7eEWEdq+mqozR4hBxfUb4p7AD0joRqbzybTk4J3hkjDDMUmDZNYoeHARj8c
Gg8qKlgazADAMMeMi0+qeIr8q9lPqpr/DRLkaokuEJwf8+KqBQH+YerWiJWhwRlnuOqtrmN7ZC/U
eJFCQWhxdZKOioWk855NATkZYTsKCIdqpcE+E+z2mm3w7SPl0CE15GBNfjJAKf7iFByg3rW+DgDu
229aB8ve47XeJPk9rRx0uvjLnkRv1SHMvpBZaN9t8uKNVpKApzImbZeGUJ6cRLZR78VMqfektcAH
1M6Z0h7X5nBtQY54TZQIiLqfM44cy7OLUMNo5VVtUkER774rbQD7EpR1yy2uXXyYGgoyYsM79leU
DGnjNtFMpuVmrEXumsnMYaoPrpAUDPZc5YcKlQCAZK8zKMOc37VtsGOrRgNbzT79O1mtIJc3GzV/
VkwopBQ+gpfdH5TOXvM7b0reHMyYZToaYJfnHan/RFCjW22ph5qMnFZB83NaQC4w8LyYYEBq0R5b
J9YBJjEdPSMzCooQNo10rIL47eMsAUIV4mtoXski4xRbX6R7+KKj2PlDHtT8Wy8Bk9x5OJdYOwdg
OJa9j27IeJJX/4NSFLMQK3gefd60hJf3oFI7bc/GC69i2JjN/Wl2d/xqVgCnN7t6HrjN8vIFSQg4
p5EJc1ElV18OEkuBaC1DWnfTX/VATCPCi9rdFInDYGJVP29aWDk0Gg9ZHcKf9GNgZXyU/KEnKwmA
G8uEvyoj9i583qzwOmAgFo1eh9K1Rd3+PrDJVr9D+oYOx3497l2tneDWMdCVpEerQ5OaPX373LCs
Bon2dNJZA6JewZ64CV1rKCBpHpxlRqu7+eA24tYQnbFjqVHsOebLfkCAls2C92SkZVCYJJPFsX7B
B51lxSxl/qXINk0DIo+Fd8Hc2bqrRvYz4WHfBDemkaf2OQA3cPnlYgYmdjBPyuFebJgbCs6Fvskm
SFWDfAUFGCTeJ3li9PwXWQ+PPQXDRIdEglfYyFr0m0N/gwxErUzsIm+LGdsKV4dx2BhmQ9RBqvr/
OahUtaW/R5JIbJmiBB+3TTWLXOHV1p6T7ejdLRsMiwE9fITzu1vEatJ0Bt2JV0y0/3x4uCfTrSGD
mtAWtjD/r77Dn2OiM8jYr4pTZZo8Ntyr0rzE8tkJ/GQV1y/YYt78hozPgwNTOHW7CXtRR2ct4G2c
KCsmdoWqF7j0XCCUNO3js11ptwN/J8dWd22u5qQUdAhpUK28W/HR9+hxXGAyizhhuzUP8wm0KTKC
fWFBcGrvKQoGPIZUF2UGKAgaptoBmkuwMC9LnvTNwfcv2nwj1Ec0V1KsuV31Z1uRq0pxMSPej3zB
Vq7uVS0aj3Qy97GbkY3Bb9/qh1BWS6PpRBI0KBCKaAkuqbt+ZbDlhLjCrBRHryuEmBNsCt2CLyUZ
JBWooKEkV+7s7gob6YdRj1aK5lNByiTv3bMQ52XupZCG8cFo/BnQA5bQ2aWfyGUYftEbA9dNJrIG
Wgbu8Z4JBToeAnx4P6S1w5Kx2JgQEvBzyMNwdYSnfnPNO1KrlECrroUUkTDGGIMtMA4Crinuli5B
1PajlGu/5gM9LLbGY/M5nRuZvc9aCtyxHdQbiMPvJV3uQfliGRaSBTKa0z7EXu7JzJiZU0uc7LLP
tha+YmVITT2uTPL7z8DIEK/DVfwCxqL2ypUVQzhd/gVm2JhUklX+IY3q06PM4TL4Py1mrlM16ggK
zJkvaCE62Ne6/ikYC3isVkn6arbCnfZJd39IoRceJUwpS1mlMKGzPLjF0PuVcbHyViRSLtSbMq0K
EXOsLjtLcpIIP5ioZKfYcClpgFB4Yjp/aZNHXiwKHl2DigHHqobrLdYhI13TdG1VAEVswzZhW0lF
IfA3GFSIEe+DMpNDwlOEreuorVrniacVe5tljXMCodtywf493kw6EEJsiNrfyiLSkk0qyhWDMjJM
OZKPoenEZYq7swcCUdOd2Bcts9C9R938x+vwU1ycVXbGWTHQpolbzPzbfnGyXQu7E7BqLcAxdJ48
PfUR/KIbTzjFtK9kdHEPWOA0a+4H+cR/mA84bpTpFi2UqYEPa5f/vQyLHMaRIORSn9kGG/eoSIk5
tO3Z7BiJwyG72/vQMnfBd2DTuEhE9VjPLO1p9t7UBWyyYwEHcgyoqAFbpk7QY+0pNrdMucOmk1Eb
81V2xQ/BosOKP4c5s/QOwiMPgFBk74a9TGzE6G1ZmnUJblwXR1/v+41coidUWjizpvtNg2t4LEOe
7i6iqS2EXkGtc6R782SiEzZ+aXRrMVNqvF2dwf4w2Ox+XFAt0CBgy/Uty1L1pMbYgBrfysenN6zy
b0+neVNWyHreBXpwaGMdguWvTX1U3JP5e0CmSrrPQVvtFO/4ofdiAMoESGiROk3drnbRY3VVs8K0
ve3aiAR1LNcLNFCQW/sMwHyVP7f0wOlOkFL6dZeLw2EoyROHZaaaP3qrSI3If9ER9z6xGGEl3G1R
r6bLJMIMmK+cAURmoTNeO0IvD4vXPzO2CAZedSm5AaBZRxfOGQ9ehPLymwhoDlbuwg+uDLhx1k0P
nJiKqrD3fmDulnPcdWWd//neCmlhdePRr/2SG5aqYdoQrzjwh4BB1gncJTf5/+zvEgHHSudEKzHo
tPAq1vUL3hAz/gU0R9VzAKRnwjBIeZFQ5dU9pFNfYjCTaWeq02cCv4IIAX+GUBsk/jM5b/c/Vl5C
QGxj1IDf1MOAtnQCn1tLJBDSm0Xd9CMz2ehTroByRAgUf4SC8xQNcx3QNr78ezHELcKz5f5M+2qR
XmljyfCdRLvh+1WMAkWjsw8bePY0h5Bp+JE//J5PLvgOuwPRsU6yXl+gvvLkvR+exI3RhZq4EdzH
W4446NqTmVvjt0IQDYTLJkXTXP2SPmeqK/0A29quwy+YhfCTZdamwVdXGvKHkmbOzdwwL4mb/+G3
OBpUQzBugkjQ9b6/uL5OGpdoXUjULrODoITL8gkAQ6wcU1mK6jufSbTkhI0uBbxWn9WkjjAB+W8+
HI1lOLZ+pz22KNPtZ/EqOe2TyixXUcomFvY+h4c+72TDRH17G+/LIx8EhzuLh5/lJemFQ8FePEe2
fEGpl3Ref/kIplbwJ+EJEHUSoSuZP2F/oz6CoT2HgVTk+C9gC4CW4p5zMoxXX9232QFRQfqdBx/u
22H1beZ1b/zx2JMWsNn8tTtnB29wLeB2lN7nhg+6PjHw41r4ic2+cUvnXlbTrG7iJBMD6JXvVsxz
fosjdMcjE1IWgds/rpybfxBA4RGWMQg62LXlD236PoKxHznXHY9TORDVY5L9yAV3H2d/4kZsN72m
KSs7g1EVT6fE9AnOmdxZPHfIGlhhxneN0TGpjKDmEXd4vvdp1HIoQoi+J6bHOgJMiUxiGid+gPim
gWvKQWenSfZlRUP89myGSZ8qPDpJ8Qfgrk1SCyUmQYpwHXJlUSvDTVg5MLNyx1IXxKtsdi7SVgrl
+mP+KmFZlD1hVddffcjOqWuyr6uS4vDQJOpMtQhD2hcJxyHZVDvU66/aRU7862Zlyx4Ybq+hWyoc
tU55rarKCp2lrnGs4UMwnYf7Ojh+8V3YIxDX3pctwVcLXwocVMkwpr9a3S8DGSKw0cCdhbCEMV+d
kAwiZ+FehU7VTSWKSV6iJEybK8YzoqcuiLO9tszoSvLxp2CnOZohhaBKdGYXG0McSoUzNbpdBIL7
QOhUlPZXR9PzN8fu0q8Lb6KFNRNL5MuSXu7D03GHLfkWMdhpBNd3ObbGk0tgosexb26ONyH9yTrP
yKLWVIOIS2polZFCVqudCuyGFEpCC8GGeprNj8y6nTgFGSeyk0C3n3Bl3vXrIS1c2SI9o3K5evNX
daIpP4vimjeVFYCQImRBLOMKCK+jz5x6LArWGDV0V/E5fd8qR/7N4YzTJVzEGwEqYqG9Dx9IBtva
+zwHIywylVziZqopTo+Gp9lqfs0Yz9dyWWw7T3Tvj40bEZxw5Z6n8/nAcm/J7cv/+OpQ+1g0ozpF
iDo4njigC/HQzInb4ISLk0bWZNF+mErPi/OyI0DKDWR3dYCi1icj83gUGyI1hnJdAlyoyGnZlz9/
HC0nsChFve1rhrdWcroleZsIad+yUhNjrRQgPqwws4L7dWX2cDxGscliRUSsasKlZWBKreMXqbl9
m98+1rU/Ug3JKYUgP7BSNc3YIiDT5WnOnMXtMz4bSbf1T+YdOcnjAIenGvvTDJhiWE3OKjT/WUH/
vzwB23Uic4G01eKZVazz+jR1oHkuMluWb836lY3kIrZxuoEa/JyLngMbcspKfKrZc3MqGavYDjG6
afskGBSqIvNJMIq/8dZjM1l2YPhXywR9dc4F8S/MXzZNbA9y5X1O3lkNEl/O5QPw/joLZQJjrXqr
57BoLKqU/sLowyAiVSsA70BvqD/hmferl2IyJrRNcOedx1iD+dpnKb5/C9+jqKXnN0GGOY8HrlvE
RmoX0CnSYzu1UkeYltQ3MVg/5s9NqnLBZ9CvFbQhOaY2K8aPMx2wrOs3yVw8hmQ7SGHzb1qhfMtc
Va/9AeUIQY4bz0/sbcXjTgkoTU9LHY+a1PaQyhN9wVI799vN6l7THKkPLt5gE1ATcdlyR43CsQtn
jsjnA6UImdWaE0IIm66W+zmycqcpOsW+1kh+K14AzB3t7CFd0VifTNhua2ZQnjkeh5ufvWacz694
0y6BcZAf0hDJQVXg8NFrfAm2pdTFbM2ALhX3BE1PPFxOQ5wXI3V6FVIEhMn5X041/xfODicauBJb
BkL2Zp1J7IXhZPYvVma5XXkqPgNq/k89UlxUKktbFDpmIfLSp1rr7byjXyGKsnxfl5MgWLbeDbNi
uaTasb/Hydyg0t2yZBfrhpgcEXd4IeiP9N6sgvS0/nYK2nVFwSTnrAIL/cPJxzuEJwGozbnysR5L
iS1DISTcq1gehcn9FudQ05A1mQUM16WLGkor7cxPFx7bcdy09vV8RzMPdGbrrbTQ3TO50zWLxDel
/39/843wLjaFG5n6xcAgV1qvOP2xOQWDCSPPwj7cMo3k82AlErG4ixiS/PU2fvmIa/i5kOVXW4BD
Jygz6R3ySg0ujwafJYrPono4lUUqZjSOee9VPC8EyZalVA6BTheyF4DkHgbHDWDL2Y07VZKFCh9z
rQnmxCsz4pB/9B8B3vW1IWjKSN76NU+Q2JwlEvB1BUHKGNrK2gIOa63B3bWldfcggpVlR34gBczc
td2yxhJC9VIe+H2il/SKAIIi+OXztWpsr/nQmUFNJk2jC/qk7GE+5T5lvUPldQLUYqP3bdHg+i+P
mS6MCZ3oMTau9wuStHLw6xfH3Sf3p20qTGO5PQYmLB0DFq4rZxD9N5iQ6RYoljxHvbZNI9A2LKof
SlUtYeO6C59myYN2uDd28bwz7ney4D3N7K3QkCBtS3J69EWdRni2pVHyKHy87IOT+Qb+N0Gdcu5o
iveMOpQmPLKN2cP07H1rMdCwmNk+HpevP5OeuAW1rzLh8jjCneluHCKDx/pQWGrpHxo40nUuiekn
ObnMLNYdOIojP4KbadeTfPNNXCo4iMsUhunLv23+fHRgOYFdYt9592kik8dmDFu5R09k6uQrEDZn
ZTalEhbQOW8+fwqQEd0sRdIZxLp+b/Pjj9b+wR7IVARBC82YneFWGq9bmXMwAdxTOIfWjKNDfgGv
X44xfdOV8lbIUTL1l1JN7SZsd2d2GShZHURJbgMtK4Pk5es7FA19TXmxDdmsurhjw/Oor0rdxxWq
n1TnvlraA5GkS+YsffMobT1yYrZcLr6JY+Qvb0LO5+XrqHp0alYjPEY973d0n/b65bWFLoeWOJJ0
YD8zMJLqbOp8uD3+RYAOnO86w0nGeHgMNQPowyJbE0BP3fNdYqL4szF/kl3vAHCMXxG+5D1HxsfL
PdC0B2ijXPoRlhWJ7Ho9P15VhzzNBV1prDB3lDs3gpQJqnaHFRgrjKl9Ndl+vE+ptta/PEsDsIS2
BaulW2Wb3RjLEy1h476hC9cqCrdB9W//Tet2qmiFDY0zLTi86dGuHIzVJ7zfjKLF3W7Q/8nFJ28n
aYTs+rIdea9iJ7RsjGsEeLRWYjfF2c3YBXkJ6PP1zuVO2ilPnVg+xoWg+BMt1RpD98HfTV0Pw72X
2O6ct9QzJIMREsDKebZcar7LcLwNaxZS/g0xm7JHW/UwNrze7jj7nf6tGOZ8kzPyOSDWMPGUWcrr
ZlfnUHzicnjXpWBRuZcPFRcaonzqwKZfF7umZJFFuttWYkvXy/SprpCKb3ovyjk4r7IWZ+UyiTp8
xbEAkbtscWNKF3bgimfFE54jrDUTqSQljAWVOibtznPrv8+OLoR8QWUbjo5C/CBN35mexxajgsLG
IuHF0VJ4RLg5fp2LVypPJcRBV1N7HwDip5iEf1Ii1tP9HTERqwDQeAuWpWZr7AUhd52OeOkRtVYd
TVBswaf65fVPc+GsUmrN5zvmV8+xNAITNXamLxhDH+W7va3xwgwaAkRRyVtNBcyCM807b47CwZIM
6a6rPkQvl+fTZ6BkIhQcTAXQABSYYxLAjbR5qExfxH2544My7QvFjgNtxyx+G0J+QZzJ26SvPP1c
f09dOseV9Z0kHfXtvrnmhGe4NI1kwCGCMIJvGwhaROwL7vGVNoXzB+7GFXrh9VlukAor8CjUmyhe
9MAxhqZ3uCPkdiW2aF99sOoRjeyputt+pnkb1JCnPYX4hyvG/5rNg/w1w9DU8gkARYPKpp+OECD2
k0TSCOouUmQS6E02klz+rIHns7uHd3MsKSVMWzI13zj6sL1Kpts65PkyiZ34JjPc49sNBB77kuqr
vuGHRiC1eDOUNA7pLzq6TmSMNJnOv6C620QAIZcwDhjL2i2D//r766FI39lTRFsLTDsR/LWJ3KfX
9MDNj4OWftaNCHPZbn8hcqzKCKPnAdUrsq44l+yw4byj736rK3N4VZKzPGOMkyFndKlpiZDNotMQ
BJyua/6Cc98foILQvfzwn5NaSc+A8RDQ1UychrRJxIUGs+muBzIrCPWFNBuxwVKetULdPXlVq84B
GIsuS4VKJb2AqEbmDadl0kdcIAGtokaIXxjYqoozaePyp/7nGrPlEEzaxmPRsYNKr9NmbyIqCXoS
KVF1w5BREcbb+8Ni6u0/Q5nU7QV4DXqNv989piZ/VFBhf17HzVAeFQ1I5K4w8ykyW1vM+D0fho2X
EeFKGuUa5pLFFWlE2UgLUINKEAkyZBOgYlpbWzFW7btYtWAiHVYPFG5HtF+W/4LYffXs6zYB/rKP
szvbPSDm3xz+6vJRCZtr6C2GMG6y8VFmsr1SC8KuuYN968pz6en0TepqUUD1D9cGQGad1QHGYWW8
zNjySxmQ3HSvR1LpZk5rrk2LKRVrXOU7qpJxgLx0Vjqk2Wyu1wQZoBVt/SrtA/A04nHGxj+IALKb
5353fdlUV2QioaKMqIMmjU3g3WOlWWxAPwv+VU5OHNTKimnxj2xw0JAY3w6exR7hPAWrZ3vFEipM
/Bv3LrPpyxXid3iJGJvsPJBaIXJM7qIoY4QxmqoFAp1v43c2DmAdJwvyoSBCfZzImO4Qn7DyUGn6
o0z3t2yTgCacyaSWgtPDaRCI7rXGFu91+VzU3jva6ro573sdpZF+c8L3KrUXB5PUPC4sT2TBWzmB
2lXVOQkbHPHO9XaxXuIS+cr/6Og1FjSU7oPePqgWteTHtPNVyiRmvUnXEwFwOlr30m489ZiBBm0m
pNx3L1wkv+0pCyga5i02NZHFfjAqaXf/12AMlU6IMmrl0DNn8YZMPBMjrMRkmr7wxydas3IkL0eE
hJfJgb1a9j7fhniSTmn+8VHIgXUvpXpenlsTbiiZIGXCi5/Nm9rR48C6fvS198srl5NBLOmintAW
tmX5cqk5hUqLNSevV6RtqbFNb1fsPRgHZO7WEcV4iUgOAxdDF4iQSMsj6U3usUnyf7SF2BywvYhM
IaZbOTStWLGhQK7X+GHbsQrkvPlyo/H+FDRH2c7QH1ueSLRuzQrJP6Oq7ajai+dFOUb1trv5N7vQ
Y+rwYUu/QSstR4vYxg/wnj6tFkHsCr0xxBXzZXUq7R5EMRVPGlpy0ahUOGa+o27kq27OrpyLp/Ic
ayI+bNEx14S8mYXPdMXfNtN35Y6QKs4m8GJrIt5HDB2KjPvg7f6JaI4dSxXpqtWcDNrVbLp4x/I3
VUydxol7QrwJQEFzvPr6gQIj+xu88JKqNU2njRpY685UnkPSlu3cPMhzJy7UIgvZNY/JG58ljq18
rvKXeR1Cd+Do0VVydOmX8R2lRXpba0PeigwZ5oamHyw8bfxH/IqbFsLXoYRDltXgQRz/J8V2ZG7+
F4mPSMJ+QjVOXUcDOjT08/OV58CXszYRFoKQroBiIxOPq+AdL35RttyPUG+pII9j8aD7FbLtxlBT
/xIJkdei1jExmsYkdHtprERTzIZXR+CGnlpBsfVW+1a2BTA7HpOLlMllC/GRGN+ocDdS/6VAMe2y
cHSc8sUd0jwI4+knRlYEe0975GdxiHUWpK+lnbC6U5o4zNWc56Awy6fvR48yZADUwf4A4pSR39t1
nrXi5yEwr574HQwGz+7mP17uxx+XDnb/TtDoqjdzsBX9KldB2iOOFdWtfgcE99Bb+azTIAVUwycB
JaOyiek8hby6G3ZXIRSOWhvFnfmTCC6Cj1Tdi7Rhb3dzQocivArTG4vQRJl17Qhd2MABt3h656Xd
1p7PIMy9LH2HRh39ClSgq6GN/H5j2Bt29RJ1WnddiRA7vZICH1T0jrP4/d5rb/ZdNIQsXFsXJRaA
SPckfDYh80cL+9hCL6H+i9uFPW2XY8J2hc8VSvDmZtnDvCy9SCPoN3IwSwHKk7h/rtBZNAKA35fC
xM/3y4bmrnto1SRfXL7M4xonQVWRTElcH/+VpapG7Y1xzo4khNysYL71EB0iE7xh/24z/5Dn2rYC
cT0/8YZhlYQiDc/PHpOBsDutLRzWgq1ojPGFlzeNBxmupelWck+gF80rR6v8y+G6M3GBLwT7HB7k
mz2BP/LZbZY6HQEtZmEwseHw7CQY/Oj5BkLGrz0EkUDx9rM5Rg2wY8caNSEPtV4l81r+Qk8/qlO+
V2XEn6zWZ8GRU+CPWwZRNtjxesgU2iTcs+unl3fbfDgBTw1qMPvNibDEwB1O8LDMXW/5GwS5CQdt
ogiCTE0i/RkBTD96CSViy1Qx5zCXSSeEE0b6YCe4bcr0yERNHovlTs1jgsw2HKuK8e7hxS/b0+6x
q3vxGIyCF7AQklNvjrDrJdiHjulc+K5U4PnCSkzqRE/gJR35YXjrirxlxfzOOZHfiqyTgOy0mHNJ
rcNkP+TYKldpCGdaWjUBC0KP6raiZdmYG+UpPjbIgl2DiUiSmPr63MJlWyHdXMQiN19s9r2YgJm4
NQfPH1XZiuKhsS2EOy1jTTXdZFgbtI8JMavwFQ7MjPxyGgGCAMzBbmhEbUQ+ugBtTLO6L/vgzUWv
y1ohH8kfquT4DZXQJKlYB0/myF7gzzhqIakaBBNedbTbuzVl0sPZK1Hifm9o71n6Xuzg86rzuXV/
4tG1m3j7BT91j5XxRXr1cP8KdQAIEw+p2AByt3A8rYp92J4JU0R5VtLcmAaQSXxZvGzt0nICyqF9
WBHo820fp4vsg6qjR4PUKljKKRa1dtHjqI1eVeADwSu9EkBf0f81JbxhPc2OMZoqqCnacebS/fey
IdRjLgJPG7HBsmjZ9/TgYqnvnWA237IstUtKT1qfJ9CCgqypvasGzTwNlxfkz3S8g6MSW6oF+Ouf
10f+YpAZNhHzEjh4+ofRWpzfGaUpTjC53xHVp3SWw/TAn5vwleCCHcjnDxG2lYJ/hMR+cCkW4jC7
rvhwZJZw4VrO3wS6rCaKoL8P2GMcwQF6b3KhwzHi8OelatcuTROMfNn5QXPvlg1LEvhUR66oE2CO
XEKAXT0vDeDUuUZFg72jX4873st8H8r0iF7g9BhDw9Pa7QmgONtVgxUeTlKUfudEyLyc1vlHVLYh
t51qpTbXh3dw6ZgaZsRn8L7FF4YFctZuoM2lIutYnwPNkxEo92Q8UhqshPi5s7dVa/Hdv5EZ+Fcf
YsIOJRrGJfF4SUk0Xe7PfUgKfdQcrxhzv4m0lLHY1bTgQywY9XH3FTej5unsGPx2UgSv00SY6nH6
Pd14bGexlSi8mkPInHQjd2MqiWWq1xoVMfiCDyUqSRILcnl++LOEtMbUoR1HluQyt2zuJVHvpogV
HlgX4TaLv8/UGfx3CCldh1DhEU+i38pG912VoMcLFPmqw7ibqKzMY5ilpRM9i9QtY3vsvRtsCKkE
VBTq6UUYYbMLMvKTOcXilNIKi1P654u+iWFcYAdZpRzbPIYXEyOXiaThhgQxboRWyZJcS46bPTtl
QDjo4jmjGAOO0b7G8kh7uW8UkoTAySuysZomz5nJ0dWCZFoBSNPGoWwdBrW2iJ13wdHRn3xfAyu8
mFGt0JZj9Jic2bvV+o90bRdEILUUVEBoOdrKlIJTmbJqVro0GeS5RthNVKtvsZNJDIq8pAbOwkwO
SE7Fhy4i66O7fbDFAl+zYpK/nuz1qQXOBFIq20xv8bK11iD6vVZP81TblqwjnGNHjmaGeJKX8nVe
daUeAphFDkrNjOdJLdyQFQ69rlXF0O74QeIiujfrcOnB0WdqnlMN9boIyK/gq5F3WguNN8XFEWNW
VfdIXR1m0bkwdglWiHP87sYXp0aJ3TtbG/r+NJ8G42QkPdzLboBg8yySXZytJsRfVsGediclTAAl
wchsrGXIyMEB7AOFC0ZFR5pgV0d3HVd8s+F691TChCyVnTGk3i63GKx+QhHbwkTPW+R3wRUW70m2
IPpZxRvLDErLR5UWc04vZtT4mszZkX3IQHqI6EMzrPUKvdCAFhSdugqtqvpzGAqyDZ6CpHrvyUtV
eVkNi3u0E9l08zuvwt457C3lL0qEyybkxYCHAeizF/WalDFr3zv3eeHuNeNHuw+/WM++iGocIo+l
1Zx9HG3BCsEQWI2Qp8VrBxEUc8e3wqIQZCmpEpD8MfAqDnUbpDXtAv5h/POSKfljVmTFxatbadgT
jtxnxXJhdOGT3jyUJceDpOr1942111JemklrH+WYmNJPrnJY0cyXrj4f1Q2fJ2KFVF6/YHLr6rBr
G/t8ijnZFkSuyI+J7jZinb8mTJIvpf3qZPRS1LcbNGcEKcppiylBWjJUq94EmGaFmzpepXaByuFr
NETZvjy+gOA9u615Q9+Sn0Eps+i3S+FIReD9C233hzJKiO2v6I5cMlaTb/3NkZyfwjY5ZsHPMvB2
agI03p1Dtpdl2Qu9TOej29raKJ//l1/tK3bBENHoq110I4JFec+oDVmTc2BDopsRFojF2ozOoTy9
XdzGO01w9F5hs1pA0SAQqBynkkJ/L2Uv6S2LUfNkBjSJakUeDEXrJZPWGTh+J4rjEc/cQBR1YF4q
a/hHvN+btb8XGB9Z6ZQVC0LGWcBgZQQC5roXLq4Lqyu3qHX24CLoCx9BZnyy9wc7b5a2cKP68VHn
snqDoBywOb0QfWZWpPu/oMFfKlboX8HmC27udYy2DLRub3RPKcV13qfSTQJdeYemXFcBib8Kj9BV
8001gOxQ6WEwYn1QGIrT1CyxDGCbvEpFv2qx2eQyluQsEKvcnt3HwtKwRFPCyYFoxvucBN4lYvi+
sLGSWEpCdOWcaTtsLhwjEbjhOu7RFKK5tdveabdY+Sqg0V9UWhtArBbo+BtmpSn8xUzt6EGLMv89
HHw61r83VsDHU0aVaFaWedhpjk1hKDVZ8Boz2iBudgiBU5tZnXC4FCBO6prcx9X/PqKpiBCYBRF1
SBInfx2cWeuGwGJrcsk4zLdQmO3ZFAusScMFng/p3VZeBba6IPqbAH+Y7GzPX6T+yKpXQ2zCX6fF
B6c0MqoANUI6hhVZRqNhcJkDW512w1wGyVQ6OdzlVbvqQb3f6kBbb4ujyKigkd7HOe6nWM6u4PG/
E0T9kvo93I/cFWLxamTtMKMdxbBjcOO3OdbwUZSNqb2XM1rcqCZ9ASrt1HrtHPxtmedV5abLToPq
pJ/qaaM3mfh26DxKLyX3rRFuxPZGh4tYGjZPOo/saNEaLPfE6fhuPue//XdLOcyH3Z8VWSbyPwit
ie8pbxE8fwsNujipgTfSVuZef4dd6phcHybeJavlBjOO390kwmFPonIli7Pz4bHwYjEjfT/hQqf3
XulbUXVjgmwoKg188HIadbTRYe0a/S/x7a1+5n3n+8amU/VXo7YewZlB8Xjnqb20CCkJGbw8ZeeF
8XpFbcrkubWLspwFlQphOvv08TF5MK1d0BB9eSmX64p8kalZUE4073vH3MQO7yCPSL6qqVwrfcjw
51HlYYwW7ZmMw0ygfWB3QOHTOdLkSD5HwwomTAkqW+G64lmRAkZvkOBVslQTQ2ZScXnr2nM4T1dS
K40FVBD80FNAA7a6AvTjLFNcCJ9WJrhR9KCfYG6jxaYKakSdE5I2ZWJE/5JiYRai33xoZxx8PfNb
mwIyU3RhUDkpnDxU4N7UmWvEkdx7PkyeblHRJTv5YC7pexfcqLIlVUAawzj4REXdIgq+cVSCZJa5
+Pber7d8MB4IkxuAaXuH/Rk4c4BhzAp9KI54HQHRgjiueJqgRF47pXtRLcjRhZ2VX7mVp0g0FP3n
THZzrwVShPQNBeHXMahWWYGfVHH+WrZgCVNUPOyEpLXS7YnhvCogzh6toc00D5gO00mI2Zjfox1A
F7UtZ1dzVprCs6rgeVzLpCG8gWyPuf/EEYAMZpuctlc5oW9XFjsrR43rlGnwVH/51YO7eE/e00CE
uKKXvP8CrGQlx4xfFUQel1rb63verT1v2CFGVlODiWGwZyuRfm+POcU90JtYqox51rHOtZc1CRMX
40fQkKjsy3h/AnmUGsJnXcuyFKsDtlRCHjolmkkr+icyPM+eF8B6ml3JI1tCBBqyRy7bw0m/KIsp
Mq5WJu73/DDyFmRazbiQjsN4Fc+XivW7zpLBNm8rXHW++NWHfTqgHfninR2g+kg95we8IFy3RWaO
RwLeySM11U3uC6jDibe7Y616oYDoTyadYl3CPOUKjjZIPdiuKBH7TjmDf2YlGAPk0bfPp6byxJk0
twtJUeMcZ/LcDu3ne73UrX99bXfYnP3jNOrzb2+qx7tY3pOpG2EaqzeYGb6e1mPnFPu3y+ABulvG
metB1Loixp9ezanCpsZ6jWO0Opawz7f7qPxlqUrwanUlGWuXXm/6X9EX/e6GFQu2vSM+JoeeFReF
yChhJ+cJiUmLcaEmO0Bw/4LwUvbL5KUKYvItx+XbJ1PG8VrRnejB/QUBBGgrfX4RPPNdQopPxfMz
TeFa9/eryTBYLNv/7v67dsyCAMv+67AvkCkPcD3mnx0ysPjRnoFYocn3D5sIg55GKMAzwe+r3glY
2FHGwczAYb+x3Rqg4Q+8vkzlpuxgLRGE4YecueKmJa1pciy4AsA/00WOg5q0iNeICYunzkplXJM2
XJaSxuN77q4QrOOC6OliXMg3PtPTB41TrFofTAIkzA75WmzXtcUHEY0mZ8spQxdIty3yELvrrrSZ
hVZOoS5vizNwRfZkJeWghfqzn+anHH8Uus4H7vNAbGqLDuBSMdmMh0CK73nbD2fIqwqDOYQSZg92
oG7KS5SFpezwFdMXEiEB+joU16NcO/5mnhQs5mO0XL1KaIAze523dd/PHaN0xsg3OHeg4CQvLq+5
g22cTx0epDY6SqVn/k4VsQ7ZaPuqRC5uWAcsGlz8xQ9vmZwxFDgM9lP8bfzBUzMG4X9RF51tDaYE
1ALFTF9fqm1vi2sgsNJIPDl89YBjQEYsdhs+IML9QCtocdjR/zfG7YE+A0NjpeZutOXLJIyYDi/j
GIJ5NeaZF8HNrENiPW86GpElRx26j6jNYHYclOex7InBekTt3tG/567TOzk3jbP9p/Ig48+XBRma
d7aWWoRgegg0Urs8be+ldP7U4K9Qbqrx/2kDuDBXueOv7KDFYTcUjoM+LSI/70LxWS4HN54CM+iP
PtFfvXXwFx+BjcqAFwyXkEghvbWfCr5dqv4u7nXM5cJo5K62QOPq0xLZk2rXpuE/93YVNdSVT7NT
YyPdRDmqhdi4glG5dbTmEX5z/vNKJq2IGxjF7zrNl9qPjOLm4CqsCCyFrbhJLDczQgTDhWkLaelt
n1SO0sFHBfb1eb1phyTBmpI8U5w2qMxqTIBiuktCQXqdaACvRI24Mvwl9KlxBArxp988i3t77Ap7
chj9Nr2hv/5h3J341ZTSeDrw9uVUoq5nkpv8zlOF4wW8619nUU4odSDerAKsQwhAF12XMz4Dm2dq
03wup3xl6dith1hmFASei8Rwzyackal+FqxanNE4X7z/GeBbkr/n8f88UjsEX9vIRwPFpNlyzLOT
6/ZTV0Orrvwy0u9YQmXgOsTR9VV4XnxtfUjpjMiBjZqoKVz1mUC+tfpGeOG2wRqCNEMqgtn/70Cs
UWOZiGTa6vdPEHobEqvwfujFiKooMvqz+an9VeYUJXBCR77Ybrm5WOg4nT+BC9xm4UqupYRmqOFs
GGDCQ2l48tQiJY8By5AC28YI0hT80mTFMO+yGBNDg5aM5e/DvSlP7NsUoURJomzTVJsC0CMWqARH
CERRcTb6bLbkWAwHxPHO5+fifA2jBOZ1+irG6vOxqNAIHMU7F7ncJU4NETd36vhk6/AgRbpcSeXA
zoyxS/nB1WbOHLbLnbD1bSF14cpvk4Z+hbvsf2LMgEN2Tc7mxqa+c8uxP+QK3FapUiyyPSa7HQmv
4iz5rYh9gKHtJfSrKs0sqnEAMORcp0yfArwHoYYHTr/Jyd3EakGA7q9fvtIVxd8WoAOQZgAIr1Qs
YxToFfmiJFF1niUAFgiS1BiUR6otA9RnFPTwClYSwUhZaLPUTlPTu+vxiJ71Qk+j/87mLW/XY0tR
cZlk5KyzcEz9UEUUy3X2Vm2JP1Ai7FZ60PnUI6P5mlD96IYkckvHQBIClaL2M88BDIRCx12Y3BqN
5JWLSD925Fv1pHHHfSF3enLmYYwRrNBCOgikOBTyFGr/tjhKS7TbysDztDkzJIkPzR1wGGGmGIbx
Gp/3ZwQ6PplkZSkwMiN3PpbYp6uM+qN9lr75abC4OlxgfDkxPQSnRKNztIj2QrBXM8E1vtfUzkKu
gtClzJmfTouxYa73L3Yoo5nqSZ4csFT4LBI31GyK4nzkXbOlextAqvNOiW4X0MFvMOyBVitdRpz2
siHmKN1yMUsHWXWWt4gsRgG8hc2FmYHD8Bf070PVoIe/zotvkvqL/E3gktIrzsiOmnXAn4gU4UgV
cqsUz2ASHky81I7nJWGvjq9Br6IcFAQ8OoToEwqBOTji/lxpAZ314suAtqfKjnGhLBGQ1XgQ5sz2
C1D2GLRmj11CXV01PJzD9OLPSVmeEo/XQW1EBE4eu4Ox/cxUOSagVu5Icow0k7kpaAEPBQ4xFC5k
Dv7fEyigvgtdXo8QdeCPiH0SFlmSWQA0aqlIoDEKvwciJSCbnPCximprFLgL6hOTyIAiCIMlLjJh
lk3ohi7wWreupOVPvOXZCi0o+psmQFo5HO2WP5P9cKmkTi7ZDt/JEoys0Q1IJju1NxW8/RLyWUyN
UhKZnvkrgVpLpPTvQVKUovBkM+LAipq0Iv58FgpuuUP4HwABFo14bJBI6gt3n8gG1acCyMZPVAJQ
QW02uL61qW7kTQSLyjzFnaL/mcZ2G32j5xf8uKBANyJNTewY/V7tSyUunz+oqQE5vaBrfyDMAbeU
y28YH+v64QC78pWFtUSg9hXGZiILAvtRZ20gSPHb8aeWp7LZmOnzJeMDr7S058JxbOQxY5zOn84w
PazPKhgVdyidRB5J7UqkAuhBKgpv+jn5ZhPHMz3qOSWatZihwGCQebEV/M7VrmD/++kxKLCzH1rA
tz6xBuhzMnw4vD5K0BcNqwzscRyozdsAUwN9FbR0HklOLi1GXTv/q2CKizT4C+X92dIvX5hyjPD5
eDDzSGVs57Y2/piriThLBk1p2wurblB2V18WGg+PcEmI99u2IhGYODAwe5Z2/HF+K4mJrtCyw/vN
PCua2e4CKXHmracS2m8FOsdDtyeGbOWFa6tIc/Xv9ozGiqHabAP+vrNGwvqMpYs+ZMV43XBD6+R1
1gH5sOCKJMPlNuV1eN/Gnusf9AU9KJr14ArDlF5zwTuiUuUjGFy6zv1ntRaU+FpzapneDggznOxl
VJOJYAH16MySds/u5KXLea0ToyP50AEo0zZgZsNQ5MBFQZRcfuvLHGTn8np56QxdrVYjtjSgGet2
ISBuBpT2IzpXMwtOJx3CsIaxandbI4Er7V2dUXOA9q4CsrcysH0yjzUs8qjNzAeeaWp7OzBl3hCM
X7FrgsqOSDjS2CTknCf5y1deCw11j+BkAg2v3ZzZIDCNr+Ufu3aluzvppovg54VTU9RT3R3T/Zd7
eGqTBPShmHdG+P6DX82zRNLl+BOnn5hLusngQdPurFOM4t1CI1axykG1GCwriTnogGax4G7s0+C+
97YdtRucDH6C11mM49YmBn94B6rM1i+rBR0WSDP4jAtev9gPlSP2Y6wbXddvd60boQ4U7nwm4Kra
fE91iWaA/tdbFq4cQrCg6baz+Dl2MzCFh3qfvkpBaZkV1YLUwdbXCLLW/v8iarBCHlgR5pgZla7M
WoXp02Xu48WgXgSRD6zUseBqZSxMppkIHqwOnd+/9Is9a2/eWrJ2gZJObu6fhBJDudlBJ75LCp6z
/9tyeruo3AIF5OLp8dr++wMgsWCnAJNAX4oLtDx4kwar+FpSdgg48DNeyGthV6g+GxPZmmp3i0ID
G5JTv/LyWohsxSXa0Zpxpb3RWC/j2rFZuCuzpnEt3Wcfn18g91FsdBsozmfDMPg0xckKkkiUX6ME
aaCbFXZJsjq/FfuEgg8VjtPeoUEnT2yhvo48U0Hn0AlTOeMtHtXtqJxrXgQ90iJCRlWWiFQZyL7n
vleMno0W69YBiknYmNomXlE9qcBcBDiTH+y6s+0EE8v4UE6SfK6SpFhHsAEERRX8A/hTZ2/pMG6b
2liq33FvobmpfvJORmYwjnXJIMfPs//Da+iT+8Vnh51n12XM1c5o95lN8efhdaATi4+agftWw+td
ziTa+//q3NnnY/L1AjkyFA5sizq1KiqtZPfHjDbahg+Fs8d+Tc6zVuk5SyUUf1ueNh16pa/VEc5I
lt8YnBInYvh7dx5xMw6SAk3Zow4muMILG+4OWgAcfy83O0cxpRsQhmvPdC7RcVA3iQOqn1F0B8xj
B9pEh1gwjPH+lC2IxQdALiP5VcwbAIfq4HZxYj7Ji5j+H29tHmihxnPhMF+MbbYfl6cMdIJgy/mT
IkLBwb3tJuHw1bgBrvfYJSdD7PZHhHtfWuT8h0MCNMZtSaG5JXpZta6PYFXi56kp6ov01KNTJJuV
4hU05R3gPW3H3+vNlmz77f0qmf7Wlj88t9dE2aK3EPm8NRel3+tnNpbOCEX15G1f/Wv689DX3+Qf
hPESHebhOZ8hB1egGc/PpWDZqqsZkF8uvLDhU6UgTZ0oilcJbi6qRwOOOHjMw+H+DhG6H5m6wVSc
umf6hDzy7zTvkCQO2KZS+lq2Zl0I9b1x/Hj6c/D7BeFFVlFSFmSw/SJ88vztqnJ7RTy8EYUTMSaR
AmeezZ6djZMAwVwOmiLCrFrDD8JpgQd+MqP8vgcSEB+Zh6MvLpcHQgdqGqe/JoJ2qDwXtF9o8cb3
dCuPc0MkYFfaAvI8fajn3XqFfRybjyK3Glrbo8f6obJUWV8QSqQC7CZxNMAS5pcmOlq08+iYBQ2T
YFgR5c8UwTtnCT+rvvNlHHyTVtjQxyi4+CJ9VAl6krVjXu3fQNJIJmQC+UVhYaf3VN7J8U9rui7j
q7jVeVg0Lzpp69XQegesCLyIsDnegFK1e/Fozx+gP6IVYEFmbvndNvm4ZGpemZN7W621lhCk8g+e
xrOmhxrSilk+vbGEdq1sL2si/w0VNWTMJC5qssAPcsY2s21nXlQag2OQh5ebkQnP2ECqX9X8Cm9q
PS3wg1iNh8/5Er5iaNZ8EosG/8+SuF0i13G8n8TQx+/mN6H1eSE4tWMzd+P9IT23ke0Pe/waU6Zu
oEvBigo4c4u7Nm6elsZQU6kspKUeIa5Uj6qFNB9GPTdEr7mWu5nmiqSKIlLZGU8wKA5WzLxqkTuO
2nD03F/ki0elXoeHqx6IOLK+bTkq/Ps326CzLOL1dyuGRF7eqo4scOxETQuHCzjGXLme3F4WCbwy
NkuZMcLC8T7NcuCgqKtnfEyUpbtRgXdQxagQ9qQ5fecpxC/5fplokrmjTDYDJzg/vOaSGTefhSMe
A5nLo87dl4/fe+o9QfEUNy2OJyF7GhmUEh183EVHPupbn0DRa2RgTzcu6YBC3+bdhBnsMru1bAz3
d+xn8ftk0ajspT5cJk17x5SalaBia3qIZkLByaOyNITkdOzU7ArXm+/K3STLokWS/ITvJPZ8HDWB
sEnkuQTcj9igPxx4mDHMf/shwR7nO47TwQ+yDZgOoO1zACUiWZAXtpnZELYLYyCLq8KAg1WWLiFF
2BfFRU1TG1XSS/NSRKV6Y+wO07fG385OB9td/JYm9p8nknVReQArEfTkeOZfPzAxTiEVd0TjbSGE
6KtXowQozZ53lZf4+oC0xQ3tk0hhkuinu0C5PbeFyGYhS1LWj1WSG1XBXCcTzXjWUGh7hGrKpeVm
iAfekZEuIcF4PPbQgWT1Qnbk6VWX3ph+kCb9QB4WX8JHpvLx+V17ELwZPAe5Gbs8HkrLXa2miWzz
YxycANn/schG8NAaQjqr3PWRcFDI/kkFukC9Z8oqWy2kdfeSTzoqW83Qmiy9lCnH3Kt0v7TZf3Cd
PZagRPLzYF2t5qjuxkflhy5xNRd44kGzA66rcYjVi45TVtdrjdKgcYhrtqoMph4nki1Y7Zx3ZOdm
AhTafuWUr+2j7dFNIal+QUEgXjmtqQBc442SXr8ywLF8eFoi1DAlys8XOfz9sN7DxH+jUxSkosxX
0jdSj+nYTXs45syl6E9iUPAaz+2D1gFqWNNjNi+JxD/uV6HWdoHvhSbhT0sdN28uHK6bFYaEglvV
beYn9MrSLvkIbidD2dyx0ncr5bDpqfWbE+XBcTYuYSffgA8JdyhKk/wj6Cq8+IKOK0/kR3gguIhb
8halY/lqqHy6h446TZ5nn4AFvffFUX/dgonqvSUjUXvZlPXa3GGr7xt9RxUwP8eFl3SQeFZ5ROBK
tNeNOZZWOYV3+Sq/A105itiwzSTVHaCaE4qKBXML2Ei3b4CtkSkiUP2xduW0U/vOcXsKRKVTR7Ye
2twXEV2yLbcyyLSLL+Io0twE6fvgObaDAT7tiuEhwBcm/RHMNzn/ZXjZAGwBNfnpS+lh8qfJi3rR
ExaY3lMI0kQGmQLws7bWnEObMwLauGnnOSZiHKMswZcgxmXO/QdHIUq4lrDb65BTfDK24qaen/qS
D5jo8c/EPm6gEH6K3WIhq6MwwfXPsAJ2BxtKdmrPFvRDdECJ2vfRdGzee0jj7cFOIezSmOu6KG/c
dNNjhjhNKTONUrAzioHmaKZj88MwHUT9qLD5c3oHwek87cd0X/6RBizDYdi2pbNWPOcivMCB4nSl
MyrEdYAcQEeUV0TqtoeDp9QQCmMAwVOXmUvErEkm13OgaLq4tPn0B+8Y+qNPpJ/SR/AZEb8ppsUt
joxL/6nWxOobgOnlv+QAQyEj6Cg5MnVkII6jlkxJV/Ua/CgHlFmeLvn/go2JvABZDSiViBORGNB2
Yah0B5TDPumrVPBEAfk4QiN/lFx/cGJw9cJO54GBhqSehggoicJ0oLcdUReRsQNaNR1jsKiN22O6
yKiLhOxrNkSZ0sxygxv22pZRf7Hge5+Ztv/ewHgpl8NMGlO4tHuOtRupImK8ipxNwzt4bKssJj2g
aacx5Ob4MggCFM/NKRLi1juqUyXaUeMvfLa9yPb1lrN1+byMQbGcnG/cZYgJi57X0l5XaP/LGjXt
Lvg2xO/xsCNm+SZHH9Vb1p8mT3A0etv0StjH8JtVsTfebO3AGgk3ezCdxL13xF/xkgGB5ZcEQRd8
VOyveyXjKnjj294OULDyifWbjLF3AsnyrV2gJKlXFBFckowdCK12nATbgzZqcsV0Oln4tEKQdPSS
GJYOroADz40ei31DG5cHaPGmTGNS/RCFtZziMMfJGBN539HIAHqJ1P1avTdbzKGBot++BeEl+FYT
07Q2n4Tkm9ZFmnWx9Vsxodb0lEJCUi/PWcvb2+Hg/b2n7vH9BmtHsDnx6O5i23cEUYXWfYCHdSb/
9GPZ6Pv0m5IATI77ER5G0j6zZkNogwNW43eptAtY8ZpLTNQ49Gb2aM0uU4qFMzIsrm4hOB7nI+fz
rB5S6V9cicdmBZ5DtB8xfnfiaDLdrGCmiMi9y1RSFYPFQ3IOF2bwZEnSE7snOMcW+DkQIDvFk7Q1
CUOW7eezWtYa49z7fI16gEfwwVseKEVNmCg9BsKmAdzD5cq1sAn7W7GFr1wuqkPcI3UW1P5b5yw2
tqP/vL7+wCsmUC3tSnrlT7tIDdtHBNg9VdoGW0krIhWTDb99Xv0gm5S2LXCZ30Ihjibt30jjP+DJ
OUH5vY4mHtJIUFu6aZytblT4W4nUD9I9jHS6r5wsiiIBeMSkOTh2o3t58HD9DtZZAiMFRVOCYBps
o6Q6kWtlIbfsDw3MHyhSGn7+80JAqG6mKUT9gypH6cOwoE1jdaXa2oK3xLuxDCzBTPzTUoLRh2jf
vUl+fn/Z6yb7LcimxaIUCBfunMqnd5DTDDfKiDIpjJOSyt6/zk0qv7O4+AhfRxma98owLGntepvN
210O+9E6uYOqJj1QkffRXXeHyeZfiTn++rXpbtkxieCXLj8Z3uXHK4U5Ayp//2ljg5aXzYWnKRpa
Vsp6RzsayFTgUY/aC/Lae5Ah1zFXxNroJ1LU/pnwMNN8r6foEogsfE6wrOtRsIey9GqmjVZmRggy
wnf/qJyJl5KtqDNNG7lMc61mb/pCAPe2lcSepWVpUgd0UjcEqoEJSqoYMRAB5LgnyTvixZX5Xf6Y
ZtuAhH7ZkdHTcNY24Xru/fcAmappWf5ifJpExRPI39L7GLnTOoJxKynJZCRZnzR/bHEIppiu+kMn
eW1/63vY5Qi47d9RKd6+eeNKT7VdZKHSFxyPqD57sEVWRPIBo3ARvUYryPQ0tHbF2Dxe3Iwy5vSI
rIU6BWM1544lmQN5NsWNwXS7fmizNQkNbBoSWhFeuXhlPYhDAdPs+Gg9zS/DjysaS9HuRIl1vnox
kCTr5kpmBfnlqcLvj7ectCBU/vReRkEtePbbXn17yJSB2ppY1Q/L/wV3BiFT4Z4lS42O6REDKNPu
DdgUUIZz3Wf4LsA9wt/b/+3IQ7LExwsfpLjTLIHv5sSm8fjx3UJLUHlEus/ii8nxor0vvrCIAvC1
9x2YGSPq85Ts+h41IKdYmbqpgQVNJK/7DD7n6j8n/rdNo3u0nHWB5MGPeXAAQsiHpEdMin5xiwq2
3uoUwSPVqc0ce8wqaflTMf8Liw/shxNE0yua8vpy0sdyZQySQhwKfToeRkmx0IcEFQ5qupzMHLvL
I4Ld4OIFXF2msz5FjzTdxYEsDslwgN95H6XIHsNEMy02XeVsMOYDF5uaylkaXnxdpr5frVBTER0U
Cv77BW75yu0jXPN3UTUO6C7AVxKLQCeVonZEtVBCVhH8ZPwLmi7VFcoJvsynwRTFzfykGw+0uAgX
HlGPpOIdBwWrzcwva8vpgt1XqQdTkE/MhFde7B1NqCIOyM8TtREHu/RT8kfw+PRvwd/fW8kjGk7e
sbvd/SRhvIIXq21IAkUE4XfI2glPZAKlhAnJcLe7fXptbNk/onLFQLoozBXt1iTOZ9tahTIw+XFL
h3nA4qz2QqBI6rZ2/IM36CrNmDooCoAaUzKmsSYh0o94RKBqvh5tqOak/bCWnSjxDyZijF383RTL
4vVNlnEtVSXIlLXP9QFl7m2ibX9tbTJSNrfCyI5vg5SIAHU9lp9sbXlCtLjbuZPuNJNcp4JluFfL
7KMnc61rwuSuK+w2rpN35CnqrPq9Grr+jDJiGao+YHgf3FgyzR2RClEI7IyQSEC6lE1jpvPPOuU5
R11BLkXZYgLGv5O931VY2jl45lIuRZLqAD4tuio2bQZAHsKF6l0OZAwrTktT6XP5KfpanhcU+p4i
NJzvEC/N8qqIw5kR/8DjhV+IUloFQmRJSDcMAyXk3uSVotkjlnyYinz4IUUPP5ccTpus7YRFiaJ3
Iix6O9aSl8iGR40BV2wBir68+hxpwLjWx8D4rAkYHWtD7YJNQgteCDMLFSLx8xsmaJMWeo7Orox7
jIkmYKbz2S3wZgIiTaN96+7y9O5WJnJTJuTP5sSOQ8e2XqWYV0GQEhvj/frVQqTDokQXbu2GcPB9
6rK1zX5d2hFZNE+yaDZnPupxbgIU7CyyVGry3Yw+EgTny0Khpt92JxUhrReeVB4qmE29QAn1sXg9
bPvnuCHKdvPCs52Kx0Pay8XqNn7c2MpNzO/6Mgt8wmUDvCy9dfkfVt+OTs7waWIkOYCesq4lcLNn
iR8JvK0xuKBt6lLgLDZXsXLuCIhDchMPEH98BiyK16XAIGIEVhyOe5l7NEvEQmbhmh7cpoAVVLMA
oTnGZ8b5OILrTly2DFmDT3S/5uOd7o3COBGkqbLnII8BmSaJzsdmx0teF2w1EM8guC9gws0qPhKg
rXw3nJTrZHd35Nv62+SzbsynsZi2xGKI/RqL9JzxMncLpJxKYRj7dLYioiISbiPZSUmyUj945HVy
tKRBoE9dBSnc/G+cEuZQA+edrsznmGXMgjMq3INmZRAmifDqYfmLXFCwQgtjiSdc7MAK7KmdjCQM
Hkm/qjDkF5s0Mc7e0r1udOIHr6F2pQnTHLerXoXVAVdpSfa96eZ4BT1bXEIrUQnF5C2HpAwzAq5S
orJFqMkutT+h50FC+LrZpiFYKynJrD7Gvy00We7ZvDaKR1LQmEtvsaO3SlmvLCSZWSW+UFE5R4yw
HNc/M+ehIAygQAsGgqIdyaABEqeqtsZAoJ6RSkJZ1BifQ/U8u68lDBV0sSI9HSBW9CCmbM+z53hj
mYVMtk7SALcfUvk4lCecJnLHac6qDOKzxN62vbxfVkGGwy0BatXQ4b7e6FDhfbXX+57FP5Vr9yRL
x2M1X+wodOs4H6FyeNAG9OV0qV6iz2WHn9gj+2hI2ERoEnCnQH1H5Wt1pfQtHH0xEjHoMV6wf79l
8/0yhk9oli9cMYbA6iNMEcGdTiAILthE7nfgzvl71PTfROXMK2L3ANL0Af/6f1Z2kcZ9vZ+H0YiV
+awTfa8dm/RYmdRfgo8SqeVXABQMKQl6pF5DhY3Ucpp16ZT88GZPjEnEEsGfud8T2xIEJfT8kIPS
ukn/e/BATbPzV9cwJVoMUK8CH3UreWwwYmM3dcavd2Z5u1g8bxtHOgi/ZPbWlCAHA6Rdt6TAk9cK
DhNCYEe3b/Wla+D8hAfX2VJ63Z2NhdFaBDKIpVKFOS7z3hA6lVSZfhq1Kw9+yWb1guKPj7JGI2aV
ys3GgSJdqlafLtiw0WSpaz3KKT8+YtZ6mvsMDeQkSJypmeVJM14aTW0yEiZnOHnNpyBIJXytZW19
XTJLLTJiQoz0NtdPelG04rWveZ0b49pbodlKUegzPzGW0MCVxkinsB7FzKdj2MIoZPZRQOYgQz5r
PXE+PeB1bRUcPrjhDBX3eddfYN525hNZ7ZpM6cTSYj/qV6KbZ7YOwUdNNzLB3wv2r8wmoGvxRuY7
u/U7saPKCZRlh/wp7W3lpvBJFmd1JL7kKljwYpf1KHGBEefvyduo7Jc6RZ2fvpYCdJZdp8CBBQqZ
7y4vxJY1WzRj+709cNqgkIeWsfTXQhfM416saqjJvIbaWvGIUUTiVAG29mJ/joFzOw9U/L7853Y2
XZZBCAX0aYf8rdjBQ+PN7mqGCARw/VCw1sXV1G4dGYkeggPTAZID1suu/GB4qElhYhuI8dKRQKeg
gaYFORyLM1gX3rRZtvBddo+1gmDBR0spe4KtFOzfiqUeAPYN5d+At8vWvnQk5KNPrgeptRMdjswB
wakmfBlA9WIUbkbHYzbsbhq+9KcYliDWeYYmDOHFIvYj1oHOPp3tIn0b476CuBsQWc0S4aXug5LI
w/f74GhXuR9M/p66z+bort9btrLzHuM6+O8UUY1H6hyXaqtBwhX4eXvDPNMj613t1z+w9i8qIjSH
Qi/dMuNUXhXLqcdMWGZZJKn/0J+XSBGWzJ+UN67KmjdC14IiQD5OOejvj2hhYLd6CUDLKQ8Evwwo
KrGr12DiwjhrNG01bVd/Efu2eePMAzaOeJ/FktAWnJtnHX0YLAxEu5lW1SeyWzthd69ha4we4Nwo
T7p3GThcmDusn2y5+DA4XmJ84di1GlTtPZ1z+xf+2Zy3zUhw0R4G3NZF/9o+T5FMMDYI3hNxjwfV
S6meFQAA0GEBzqS+bOYUMw2V3IvQisqQpKIxA82zsGLlzjuho5lXXhA/09yDWzd1ekDqxQU6BU8B
ZwY/qSHYuAe6w7wAzz7Ke3k69UYF6icxll3Oyg3WRzx7ovCLyKuooEv7u0eiugT2zu5Q5ndAS9qf
nU9BfCUBH90Bc9jSro8JdXTXh2tTLFD948jmBBauSCBUvC6YKG+HHeCYJy0o1KgyUfrfemF81bGx
LZGCy5fnQtv0qRWV91FAlDSasPam2M0fJMHqgirsX64MJwemceLiHnUOwpy19I+bsPW36oq+HWOe
eafYghEVTVQurMxT4kAZtD4+aNcWjywdwafnoZyRXx7sXCehW3m3TYdEr4ycpR7365m9Zc/iba0+
jn2TwkaULkVmYQQ6v9C+FXf076fpagFI5TYcZ5Zatt6j5iYaTzc9X7glSHFDetUQ9WVItQ4luVyR
DRnNXFqbO6+KSzh3UPLO+E1y7AkGuDQ+u2y/GoKra6dQg3xxLRqur9SZDTA5OpQicr5zb5+59HYz
5ZMPYVohQiXlTVqLgCm67iZKCzfFnbhGXhwiogzs+CuvwxwjrR7efiaKDQq+q/zIaL76U71ARYk6
1pq24tfl3n7QnM5vd3lYzIGCs92h9Umji7Or5zkdYayoAkIsE9wHVZN3WfAUseFXVhZBRpXyDfKA
i7qSS4TTe6W816HMtbo+htKWi33hRIX5h+A8pVaKScvEeE3Au31cVjRnDjUyrxErEd6bOmtIAxhe
X2TXQmHaxSLcaCXgTIs1rabMj0YWW04HvrgjBBBcrNIZHDo48MkAQbR5neZdftBfeQ0yXpQmsjCZ
Wfbgw2oR9Kz8+eNTB+RDkzlfO2XXS27fwUgM3ZX8muJnV0UcMJLuz5Jm5wmzUy1szK99J+9byKKl
4uwnvtgAG7UNDG81CiwedrtJ53/IAybbcDzDBft451I4eyi0oVV0sRUl9uobNjNaHJ08zVxwHQQQ
ijylthhm0xwP/1aqBJpNo2BcjoZywdHwrPiwNAhFziXYbVEZ7rR4M6tvqjzxcriNJes/TIBR8Mzy
RvpAgS01ChwsIW3Oqm41X6hQp6tMI9FFEwE+2V26aCtyurqPM7Px6mUSX/Et/d1mpBym5sPV53u8
bgyBe6BbdfftrKttmVg8/fysPcyT6vr6SinEAf8Os/fNhga6C+aZRlTZlreodnHzj+khJYncrcmi
rAc+yxsn6cCp3U4YP7tXS/P+UXYULxHpHk0TzM563th+TyDYctLn4K8bXRXRFtbxc1nsxkM1vOoK
aF5suMnHAutzUikPlovEo3bILK3qSymXznEnUSVp3c2Yae43aLGDDCZsYtE2vU47k3W+elqOj+4S
JT2wSywenL2rfg0pLkMKTTeL49eXLVbgvxMWK+8GeDZXAWHSObLk3TNTJJqHwUUlPDu4uVU9LcBK
BfCA95EIZAkIVsyajHywuOhYTSx6ixX8hUvyMmvVNw7lvQeL/mVlHF3895gw1Zfhsp3PgYDvLGkG
7T9BtgPQvjJiOtkOug68fReaqzn9uIxMjRsi1ZYHB0LkSXs0z1OU92NmRENQbUlfdoVRPpEmnQHV
H2o+r/nFc7VW+uBat2fkaNxmfng2VMq4fF+rRvFdygoBbVSwe77y5Tq/HNkT0i5+bxdmDEZl4B08
wODoJCyFIVKDATiurcDNVdFBgTW1AoGQ4J3TykH2X49FrX9cXcDS/KPaWkq3UmMz3DmX9kb1t8+1
34zmxA//pWXqNZKYOFM/1Rq0xka0AcFsx3VfM9U3jWgPW2UJrHEFwwuUY75UY6tAvo6I44qbD5qD
bLB6fEyLKNB/Wb/UphkEEE8gofGf2iOwHhrAGXB3wDNSMKuRofRqq8TpArx+u3Sc2qJryXq4pn2e
kegF2oy4Be0HCHPrimrqaBNBnsBJV0Xm+SQBeIPGQEcSvnN+x/2PPfFrw543fleFF2l0U23aTKvk
1ZmbQ2u1Q7p02Tqpuw1W0RJnMEuFPZyKpVSk68w2Q2dqRqu2qNTrquBazowQV+P68uFJUJWNmbF4
Z9Z5g0nTDebPWn9pGvqM4zQOlkR4DFo2RROtCZd9Rn+ocpc88PrvxV7rfZTBKnabuLW3wKYSMEiU
Al5tY5HDEGhgERrPcJzd4beveHkrTHpTcDsKkFkFX3lSrh+9EAtbNGWa8P9BPvOAQFTenqjJs66F
m7Jwvp++0OlP2V6ZNhhHkkcmouLnU/rTxZksMO+wIoETqg6WYbRdq8xNCtoMKZMNDGO8XNtcM4KZ
0nELO072/dVkZ8f1iAl27dcfx1s7CN8oD7pEy6sZrWZc6k5R5zw8nLC7EBcg5ikmLgNxeH9+MF5n
7AX+JJdHGU2BjKHehP+TAc0Q8Jp+DCsdh8IFbC8UScM5C9aP3x80QB9DtJUwHVwEdOGRh0KEWs1r
06+ZE81MqacwELQbDGCBoqvZe6GpSCgZIefzrnJZz6AHt6SDbAxQCkkXo38tU3nuE2VcGulVyzDR
GKkN4DYyvVDjVpQAaFApE803gVBy9q5yyG2V5TMr6cWZ+R6/dP7FdmVObJpKRj9yET1uja90dXRo
8zoiAR2RPiVhcNDcLsNTzpHH4aJ53AxGowPz0DewHmhdD8Vr1RG0CD6DEdnKwYBXdeSrWK6ojUjR
X+6XdK1XjukKKL8yMMfXt0ngO/5YymsTzDKl1vMliehs8S1DxgouWGeV0T3SoHKzMTUHPznLMlRD
WkEk5HaywyvAtQxMCm1jhzvOToxygsGL9CzXrNGyaqLoznhAn5sm6DxyeEtLh26TfDs7d89+xXxQ
5e3uhOzYjFTZsiyNLaKfc8/Rpbi031Y42DieokD9BP8PvWA3j7LgDNGc+36yTTjICRznvfrYkR3S
aWKnD0ULhrMrG11Wx6ZONPgfwWIYR68HKTJ90MA6g3JQD2AwMqrD+Qopka8WanqeH9ZN22ZV/mDA
tnIONw9Slbkjcpm0vYOV544w6G9xROG0Qi3I9wxSTW0jHZqok127B745kKsGgGTy+Eb+ujsPlU7N
88HbMYK8fiGjbErDThAS3Hw/QOTQA8K/a0z/3UUyg2LhvvjfQNa+1or+hmqvvAhm+GXI019/40jm
zPbMTCDEemKWgVOUGWjsuhrIAp7pAGB2EyX/E4othcx6nF0rjdiFEhnQjZlHNU94dMcO0RyzuJcf
COx59ydsy9Ykppyejdxv2QLMCtwZxN2c+T7JKnAjy/RJCDMYRf6hFpya9suyMvseohyds8+XAboA
4m5FnwtBxlmEXpHiuKuFAgvJUQv1dA3uQ+Y80Mz6IO/Pa8wGswv1u1ndhgX0suno7iS56civW0P3
EbYC7qk7lZlgAA0gqEt36hxNjYaGPA/BY0uPFyTxgo5f1v8R5OvCz8THYoxrI8vIlqU7srSIDwJZ
WjO+p2J9SqpMVSU8bTwaTh4t6HidcFDwmkmiuFc0x5H+sw4MuuUpN6ITfyHlwK1+60H+0yw5M59w
InV61lqlBubkFxGRtxugE/c3nm+uEGI4Bi6LVmWznB79AmmRC0tigcHHJTEShvvXUlne7gfESnbO
Xpf7MwmuQMzJG75P2tkfJMyvrwawbFc7iF7q2ytaOh9uu4R+etijauDmgU6sriT0xCoAxSxpQDw+
dOc/BCMUDBeF6K92HnympJRq0/PAshrWnacgl/rYtFTBT7YJMC/sHb7ckBopDjqIKeaJ/Kvpz2e2
m9gYgEqqcjiS7n5Pl5B0/iaAG8ncnuKubiB7anqvVvywMr1ndvOPbBMxwAtr0oO1NWBAYN3BdLzo
MZW1t7xCHcxK5fKPKp4plPvvR7HKoSVp1JgJFm/Z3EEWOdWlffdvAIn4J7AyXZsZMaWaeFaUv9Y/
zqtnmZlOY8Fvia+1Ign1EHMePZSMMedY7wehcAEBMlSUOufOIYN/WXjuowtGM09g0CahAAGvcYId
pct0ctExcSbYJeB2z7zKF40JO7RtJQ8M7doD5I5FFali9wQIva5lsEPs6VFxfjzFwEHyxcTEGFxo
Ttz2QDoQvKoqpZ2YVChZSd7EI56NbbkyUlaRvFDYUX/XnGjaluhS6L5XhE/qFc3oQrXTTV4SpJSN
WztqO2oQdl8vP+ybW4ID/I80jXT4ES2H88QdAGkebT3Dmpex8t6Lo0CT5sBU4xO5QSlR18Z42Tme
h0JA7c0uBeW5uBfqirsAhG9iAg8H++v6YvqsKiMSfRXmCs5iSha+ucFuXGlyhNj3sbQB1d4iFKbD
muWlpC0t0VT87LDocn9SW8zXlSzM5ExaRW5TzD6AfiZW9IvAPGZ1bKYR0GdefifL5RcX/U7sfhla
CrcxEqweEs7ppu1iI7InpuXlgZUCVm7StWhU6uUKbIgnY67RQLZUvgxV17iPOsO+P+TA1E23kXn+
DzX8VUjNnTyfH3xNu5O8YYAtIU8fzxDEKtRh6hAN2EmaGskgXC5W9rve0pjQo9SK3nBSElSNgWDl
JYsmF8rjJXL2bQ/lZMgFkT08TFSnB+TJWQDaHGFM/sHt23AmUVbI0nHfO8X+u8op/d5xR8ps5M6z
skPGt87dG5crp1BF2nmHNZJT6GHIqdoQ/u8oAegU1mx1DPnJDOed4HDae64oqofV8D418LPxFsbP
R2RBf+bVBkPl5ViC8J6lyq/LyLZT3t1aaOp7ml4lWGgH+QdFbL9nRK7P5tQR3OxHnUgJZG8dWxry
kdHIowofgwMMu8IPlMCSV3cPcDQaK5hsVK5iOz7o42s6UG2dRdZc2+CMG0Xcdy/a+GQQjnPpE11x
IYMFoLYnce+Je/R340icShoQCkv0YE2qbdyUzTLFT0TwYnyw8Gzm98IhHb7jn4+kxt5YOs1rAVl9
AWAQ062/WlbGoDNuEi0J7sY3nnUEt4QWVwGekgVha4FiZ4jhh9t2oiGkA6J/16/vzNhTXQ2eXcDe
DXvdpy8vi48FouG4kOw9QBdcj205YDcYZFE/4hjQ0YjvJvkkYF2ZMbbPz1/DIindZinULGjSE9YU
9SJIC7LzmoT6teOKbowYVPn83oJC/W/rDhEmKCYziEQ+5zjbjVkIctNY471w9LtW1Z438uhpWf96
etpmlJiaZoHlib4sreBWuI1RGAj6IDqwAm9zwiU1RfK+9Mll/DjmQMf2sZWkqgdEedvB3R92cSSY
OqBCD8/1oJBwgQpnf3rPfIpmvKLP14qyNczIlwUrPcynkUWiwWzQat2OG+T23FvonpwJeJG4o3xJ
Tif1sRy3CnEOBbm9J7kttzGxRFVgzZoJkXP9w8ydx2N+WfZ3ySrTb2ZC6rNEtd2e8n8eO635whrC
mW4dytCHIQy71xPI2BACcIuxxb5B3ae1u6yaGu5U4QL5nG8F/VUwX2wakNc+iYW//8VKkCUUt3Hq
OJ0D5v3bAUrnqZn0F04l58zgo/N6hdRfU44SJFuVYZvrqrsuiezZCw0VMUdpo9w69o40NVRcIXtc
nAewyDw0+Ci9lsbn8YuVGYsqotBCb8nkRIkrjSyYEo2gOsbR1yLr1iBOCbGaKBI3OoflHFEzaPKk
vUvTffw2K86kv04NWDx7Hg0PbwQoQKC0Tu5u2IVcwWILtua4y19cpon8cYVANKUFBRsinQlp3YlR
tMQvZjT8E3F9Sp0Ds5qI6vY0ITkzilwUVhFXV4dmtaJ71rbWrEEdsRFytcifXGkdDKlbrNLtBFs7
LgijDrVVvxAdTjaq/C/jJWAE4dycZe/+wdyDdO7RBleel4iyT/apKq79105o7F+zi+0gi7rQkcXY
tYK9cRrI4t3+57Hmu/VCCBU7+XTVafpgqcVZRYvRaHg2hH3voGpJ3Pc505pCoqy/8q7We4XN+LLc
R2l4DAAXltAj+iIUhL8BUcNOMOsUM/H2XWV7yBrPEwFGtO13ZaGQnusOr9Xo4KaWfK2i3yrilZN0
dMHZt/DiE20+D7kXGzaTX1FFCTAzOOa4RaqSBWBMmdi1fNTCU0197PbHlV3tZkO3xCPqev3trCH+
4Aa+lc6AjXVG3BvYBGt5uQXc2ckSfaHxKFviOpS2MAhJLbs7Hxn4PEgNCbDAIF1+izYfRz6ICFSG
YkcYJzDZIVp92gs5ojorjKs0mXH9YC6Zi8NbIcTvWNwjPxl9b5rkMGw5zo3Hpk+6zrKcqOThW83m
vHDvHUDmyn0GrMp/lg6A81GvwkO4bcW5StYsXQPjqUPt/PHNhdMfjuPhIG5i51s6KikYcGUIXKe8
BeHqr3mZGVaBMGwoYgx6rXuCIlE5OaaLL4S6qCc4b0WFYTlTdRfqH/Vi4yaSLMS68Q9z0t8bKeYB
up+9riEo3/oe5qT5CIC7Q36cE3MPYk334yRE8DYMhMG5+1nNVzsTAJIsD9/ms30O/q/ChSbp13O9
ffPcu2jRFn7Np5SPBIGxk5wt6/bXVQ9H1krmAe/OhFF0ih4DUlu/luGdJ5396me423Dwg/Nd0svS
aX3OIzkLmNF29nIOrp18ZrO3QOve3xoyYN5fTgJiAy3udV1hXYGDCIz7Mn6EKldtsPHNvOR/AHEG
VPMLtb155Sbx2ZPRRdrrjg4GNokRLsyxsaQd5uNSYqx1xmB/QSXshhbbkLs+MPLBu6KGbzn+Ajnf
MJNBP/RytjiVceWq/HXQtXoh7zntY9COqBvk6HQEQi9r2TCDy6NtaWfLB9hKQuh9jeLkvoDpt5Rj
mR/BIDr/jzdwWNMbxb5rQ6bqtv9cZBR7gd3yHU4P/72vNxV9FtNbX94VA6bl+Ul1St97WTrRVQUH
cWqua+q6q25Nkvi3J3AQrjey6Bbhnh889JXPpgTkG+1+82YOR13ODN6GLOiATQV8rslXSsOBLTGu
oYe2p9lEcW2K4c9SoSsaihvtYGVSKXL/hY8fr/qGMntVrgfrmfuwIABc0hy4E9HRRJ60SaIovp75
LhhE+Jr8iUYlbfK2Q+hRDektBhFAK+weyoOjh2O08Z8DINA39T2Ll0ThGCHn7ZZcEirbJzi3vWYd
2bZBwz5kl8lIIYByYNnjs4a3zhLWVYNWdq3eKM6GeTwpjWWV+zRXllEt/pPmzDhk2Bth0MU3Q1nv
+IXJyWF+r1y9xNwHXoDqRChY+T43VthJrEvGeYJ+5pfvqz9sOuAkugeG2dXhXLRvVwMyS5Kp5KSQ
Vd8cPUOFB4Hm/1d2QbWqm+Ryl0FqBKDExMClThAr+BG8YHE0cYCLtUHdpv7Yd4dvKBSUwdnQ9oWZ
GQYC3zLe/ZdbsiuE+e3su70Qih1vSDRvM5/eYPWGekSnBcN78jk5XWV4M+ApYiritV/5RXSc6gRj
0wOffF3pVnj7aalEHRi2RlMxgb/UguSoPjujsTrP1UnFM9sjcKJGnlSAUrpz1A1yjPNm6NCTGdsS
jADZPrPvBiD3IP11p6oMaTGx2jws3rsPOpvjl0ewwqw6vlBPae0a128y8DrphM8DoX5G6CODYlZs
yWUyhDW2OQqifpJinPJ5jtFJ1JSB5bRFd4eXTk7GkXf/iV+mEvuicxGx3GtYDCvJHPmYa64cO1hO
cnjAn2xw89uAYZra8NAPbwvgqYYshNVTG+PKIO5rtg+XJlLiEq/pyCk9ktP1Z+hP+KFGBsT/MLI4
Al8/6m/XM+o3gjtmpLovPu9k1gMHAnNGIgyUYcM1Ur9LxmMGj3dZ/tztzjjZX/Di5B9wQDb/OP4M
6v4bW9v9IUiLl+J55U3ZvHblAtqUP6bXgAxJEflpvhM4/R/SoZIMqcJLdyFLMXVe29jqBq2FgSvL
wP1VvoZ2J6vjRS47HRxuvxEeI1hcAk9rxVzjgTY6MQpu4cpuOlXoKvxRXinaVDAVsh3ATg/ERSfn
et2ie2uTQk8ncQaHXVB8wD2fLisLRtkZuir1GlpimnrKSUgKskCHQzt/OGcBvqnZgDArWGijQrrt
CdClRQV/Akh+8yIWgLpJCfHsqmudiCW0E3INC4s/qkLRSlDnRBY0utWcfIoHBXSZD5Tzioox93bB
wh61bWGemVitSl2oCYBTiPqiNnFxb0HdLSXn9Ofjc43JA2B+cDQEb7qxmA7+AqeUP6UXp6sMprIX
MRpHABe5DGN2o33OUYz8WuF0xTq0JGa+EGvGo07m1GaQYmbEmyDUxPKQZKc3oVjIK2JiLXT3StHq
6o3ips1AOrlGRtcUm4GRb9F2AK7yuXbTzLL/cFLqwyF/+GFAe+H7+szw1m0tdRmk2bkObuJJJVWK
0NyUM7pd4X7JFbG65WDEn6bPDQNVqUUw8eI43t1qkcPwm5Z+LBNmrFpqG0Hl5bR8BACyO33IVEWI
hoi2dhK9nBE2yjOu3e3QEvAkWZsD56q1Qyt062JWxV/bzS1Gtk2qYPZmUBZRy+lEOTYLWdLKpdI4
Zyg4rMUXTidJsCqjxfexxnL9+tPZkqaKlbmh/rUAfX9lkdVtXXoOqZ/sxsYa75ozjK0PfV+mNOaV
42X8Fm2OAqxiBBDBQSaciZyuKqDrlEnZR3Op4I/LAiXSMFQ6+RwtDgghuct2t43mxS50wDnrATGq
UEMMS+OdtFQTfjtI7MrCxvIFCfa0KXPlaI7dwIEJSxLqj5o9GugISqHz3vETOF8KmmpQrHwTXdF4
GzK9dOoEEuPopFVjNtjeYJayWpRbiZeUxir+L2/1ODlTrugPkDSoUJPqS57WPd8N6kQzVtJ3vDUY
E/4LckDOqoeQKDiu1Nu2tcGU58/xG2UCxWPxRN50gYlU4sNb+o76hfiNuWq1WD6JDlIogd+EcIG1
i2jC42RosD1Dhu4+cNUGZPdW4I2AdZ8cNKxYANsuXMFM0azpzy1HdsMlqd7WQJAaaxFn5rPm7iCr
w9Y0sf/qNIDI2G6iSjNRn161k4/im/imh8JPYnwE97zp9lEzauhlfJgAa9pJrx6SKAy6YEpuaN8D
4eroFJZGrK4XSjE72iDzOaaJ0uXR92PuxvZ12Tp6/rZftmrV9BPF9Suu9cZjQ2IPXlFsZPvpkQj7
5VgbutxUf+AxTOXDiNOpn4W8ksNO8hALrNyQ9/p0jNwxs2UHWW6ZpvgIkxZfcF734SwbzVoYWFMy
gCyVz+rjtzEsTYiinvgSU+jwhCrT9bvNQJaObCqK6C6WZHwv1u8PQ5vAXEM4kxBSXuNe89JOuKhJ
Xth/tRY/1w+uGXXzppZ8bSvkq6bcXs6BqS0WlZNUhTbYxhCd2T/EMEf6LmLLeXfcGOMHVeQlGCBi
Ykpeigt/ZyYwhRE0ICKHtRTJJXdT+9StQmgzRtxFCaQIX7GJpd5EG3NCn08Hc/zpUF6NH8NZn4YQ
OG/dwj2HlM8yf+zXQT3E53oa/zpWIxn0PBsQVSxNe1rEirNhElfvj2XpSqa/IiOjkHRI67xTlDkO
BuF1MCGw/FXwLQ94ijTdsK1U0Niu4iFC+vpADjQJzt72Ohwu3JoxBDcwYLaQEs81IfoGsgmec2OO
DmFc4QILeS/rkiFI05TkdkVZQs2KVIzIPWRhrEZjs90Q85Aj4VYMkVQyTq9ao1L/wdyNmS/joUfC
a8ItevOPLJf3VJ20cjjFU0eyPBXtgrTYtG8QVuNtCEgG29lvHdwCZjTKeuZ+nKub9AYn47YB7QS9
BCrs+TIdjMQ9TvzM50IQIkJpl8YAL8c4i/SbkzVzUVsDlE6JcDSL/OhAHr1fUlpFwtCm1BWKkVCX
9Xe6+kaFyM6x0ckMMDeVVPhd87zv6O8ldS41Cvr8+kSoyxddyzvyZbnKyCwhD7EtD1lL5g6UCyHx
U5lLzLZUASZffhpX4KpSeFBcWgGdOwuCHQZSrtMNAYNPrfuXhYSYmXdg7Wg9t/FYkbkicKODi3W6
4Fox30nSNLAFjcUfXwq0dTAl3s9Z8B1rCZ1eXUgklhYjV34xIovizJ5uUQ2hMRnXdh+Ii9vBXJXg
V4Q0zU6QkJP2iVCIG7Gv/DGYVFJd3XdVXdWOMhPJumOCNlAG2MEPnektazdd+bvdS4mM49Mo7clb
EBMwt8IYfkoekuWofTRrwgJ+oeyHogHFdKWDdUuUXnQMX5SN8HJHiYq84pEYCgbJJDREl9uZ9F0r
HfVBkZtdDPYv8GA+BDm7GLGiMjKf6Z9jESZyypMILc05BA6ugajR6AS49rAQaqxL2wT9dDaJvHCI
MmWoNhD0SNQIC72SKxL+aCPgh510xauLsZDYGr1lGHy4CJR0DzC0//IQD2l1kbzmbKf11yYrc4W0
StGFr5cmRrlWB90WafzLrpc5/PVvUJUFWUK3Z6q/JHoqdUPRzPuy2CPYptlVHbeReEUQKTq6DUPX
+KT6KFZuAmCeGYFsXtvtv2BmvDg9rKOycinCV44P9tXqkrd1JIzpz0j6mFZRIpY1yLBtgxZ3WV1S
NVn5SxKEFtiGdctXI4hPijfx38sYr0g+MVOY3jaJFettOowllk1wA34dozSJZhATKvc5j/Jlep8h
Nn7ooTf01tXmtJFp6gSQ2AUoJ4jOHGEADT9ncIZ2TgTpJU335343EeeX4vtwGGpGj41H0hBjR5kt
lkb69CrY48x7x1nxi/ix2lQFRdWH48Df+iDN8JLLd4Imt6vJk/FyyE9OkJEZMgzoEBWHDFZhwnWk
N6kOvoqGNRy0ATHfTYkdUIXIDjgL/Zi80vE2EodQTn+Sr7NoDX4P20Aw2FVDcLvsMORlUXzPhnk6
ZOg0iwenTvs5bmtO+i5dYc/KL0K1R/t/obEgLFVkIu35QhjTikB0kfc/4B4zFnZwy5o3FDj+QI2s
JnBED49NXQ4Z1XsyzQ5MZe0F3zuPzKCrBMBBJlkHNMwe4VLRLxYBEJYnEldSu0GxlVvXrSa2mDoj
lORz6VdRUrCqaIC5fwilWxpQjYU07H4uwrxcUV9smxkT3/O/JGfdYXzzIlV0xOhOj7kVB92QdB3E
BFgboBh/KKfsT8KkJ/HAN1Tw3OWoM+IEdJnQD/6ETXQioY+EaKFmsFNrfO3d+IdZyCzTsScotKRt
8a7DNyieJusi+ZWfrB4/M/ftnMsZympY7KxF5oL97YedPrGu9lrL4sAwBhyUcsDl1y1WBUg+GBYJ
0YFwyfS2Ajh89A+K88uxbVCZjURgxqprEtU0E1y3rYKdvOvs1sQZ/ikuoQvlcShff2a2BKQlvzEb
lY8fSzZX1+8hdbqG/w5na+cqj3Lae209Hk1ab4w9Cy/UqZ1FWpxdkzpX/J84jvqYJJD8MUGp7zRB
JouUHQZcnSEfia4h+ZeIcUkT4V4H0Ovf1OTahOFasQTT8rbn6rOR9yzxWxS0F/3e6+4zMKcgaXYH
IgCqYb69YbIqC4/MhrtyDSkz8+GVIZ28jhbk7AdNcUq1Sgp7K7lw9oOwUOOZaAUeppji+2jyAKko
tJPvTY0w4SYq6iz8mwYxsOsnJBMLWkpSVosBZ/kedcNVhym5KPN4E8iVQr+XCp8C0BcIeVhqncrs
Nt9kGTGdNqcS24b5M2WocE3/4rALCJy36HbNvEQmL2+WrXareOlw58836hdhkgAEtxpl3973cr4G
OKctlvVtbcXKfdHiLgZvvxAcC4uxujXNPv/+01M9S6NTbkPCWkK1hj11kl9kUgap3Xp2zdbbciLU
Szi1dgkr+U5Bg8rZyFUABCj+bWdIFWKHzKMoVtvmM7Y4MmPQuT49xFfHc4ehLJ2+m5Y+9ODwY/qk
N58lNbFQPYn+ocRZscMtjX6M96MCcVDtLVJf+cKFUUdOWzkUD5J2t+mwQFL0Lv5sQH5ZQec7KD39
4ZCxP32x3YjUzyl+Id5rxJeYC9PhKx7IVvGYp1cflmHu//AqQmyUuLh7SSt789TMdDnfpy8X/x67
yc9vVhEfwwAxHCIWh6U+NKg9iM4Q2GkrwF46ZC+eKp0TINIX2zyH2zNnGiVm90gsgoI6Jzr/yms5
jLUhrZHYpnTaRC81T+Ownz4JN+N5dSzbw73+6Ewrg8XdhhU1xzmx88tcjRUkyUlErdf7vq+3bAka
He6sFHUZI/4zmgcZhRXa51hNrS3nCoWM3kZEdxEd2lkpr9cwGujs7Ob2kcCmy0h+uPsLvyLfdALn
OykpKNlJFDlziPHrnzsvQvnqLruXm1DmeDA22ycq3ge1ltLLyJBzD9ZYvoe2eDI/4hzkcHLxG7Ut
ZftqDOLiic32TeBQ7CcEVgz7AALt/pELeDRik9oC+GEM/evvgsPE56kG4a+fbUSBWtaWZ/2pazWo
3nmQLmiNhxQXfXqnDitr0zGhP7hQQ/cLEXXUGXhDidul9EnntR74XbabmLp1Nrk3wC9VsaRLEOXi
hZu5bsame4remdyfqdxPFxPN2VJnzyVuGppPuQNWyecOwDDQlzAj3TmFeZzlrkbaj+VWiaxIKhOp
qJ5+RGrdyZJjureqM/lZHimr+ZN/KHPFeOtKTSJgaCuyAiAp6DqPJkVUYmPXcFS+WxEnASSw6wS1
hsShUywVfAkXebrM6qViPjB4353XCgBK3qilsLPTgg+XZZ0oVijTLrjZCq2khgEdnXLaRliT5Xk1
4RC+LKX7dUY0JWBj1rQYgBCH5hyc1Qj6bwduxuoCgfiDlfzQrb2XKEL/1MAbrDEJK7xQrtffy8nf
DUa710X8+q3Gj6svfYvBBVDiZInIi1RNQ74UvCKfh/CG31tiR34hmUaU3gpn77SypDIifSBs/lke
UAS7vAJkw4KHa9/PXDaJkRwG2BAz8Et+4esUq/GxYX1rej0ZeYLdz406GXcQGOl9YKwjGgRpYAQK
54amGXpqvulO5tlaMNm2lJRo3c07hafugHgtR7onyJwPoZeyfvfSGsxCUAQAg59ObrNvK0zPpeDX
MgTKYZYbP9JpNRLPgUNmmt0GjUc7ogsqUcCaUUK1g5npoUhQsevSjrlU+bKkJ4O22237GovlhUt1
VVnI8pe50mKPtqElqynhDuM1Ev1X/vzZmVaoTJ4N5u07ysHtVCisdnZ2810C2HjR277r/IKq7SAc
giTW/4bLeREQJjFj7DuRYrlNflNOlTeVUFKXWHQ504tSc/rpmzlZWz/Vo023PvUPdWkKL/1wOaVk
ngOKLj5CDgwGZ2PBcteLMxvZk684sap4T189QiDSdUFBzOhf71h3hLg4vrtSCVpOcNZl5gFnpujX
OLdSDErJpNWd+m9bOEJcSfdvs2qSNyLl02ZgdFexf91MYUdUBvN+w7Nc4tDrE63E1ymXe8IQQh4P
azdRGF0S0J5UMDnJ3GyF9o0tSCxrNZly2Ty3KsgoC9EM+AdJRUtMiGxc0NpF+tiVtopcvr3jYdoG
aa/Mr80IcXo1Zpa0X8qmqW6/cO/mcHzWUpGXl0ECtfIydXWEpoPdSWbgLkWsxRq7Nw+KbGU5Ulgs
SfZggmkvIT8vlaYXJjkNPnFeiQxe5xtyO0HzCwn6blmxW4/IZG0/CJqNo9OtdvJuSg1elRW9KYdE
ZLQpqEI3cD2HSPmQIfoVHXsS94Q9RrN4qWTLzgDYAC8bck9F0y6bwApuqlbX8wt3fJagb8pPBZU+
JYaNkzS/XAREYs8JRXcCZRWpsl6330j35nhDU4nqmigoGXWgqzgrPXI8SS7udJBnukZgk2Ik/cnu
YFImibaUxLvCQ/9TE0pvm9obLT5GAiTBZl0gjut16rWJ261fYy24dxrPAauHzvKyWFS5LZbPPGrO
C8GepSEREFd+CzmW8WGijGMCB54WdieTPj2T8xaNQyF2DXTRGWigYiW2UCQ+geQ+kSZPZ8MWSyPD
ShzI00A6LP33JpQX5rIcSyBm78+sPUSA19fH6osejvaQ7j4bczTwWv0zqWdE27x6ZCcwiNvY3K9f
bxAaZzExLisEPeimhGwvIeI3FkMZ0b8P9BjeY8QhbVONXLqSorP2YH3ReH66RSetmemnZ9MaCpmG
UMQrboclyLyPsvWqhGZaDCWSrCW/cAiR4CKY8mATpjdXGKLdSG9n2hepyGNSAzJHJx23BUBXXiIv
Z/CDFXkrqeY+hRMBD4/SrkXJm/PpL8/1hTngRO0Tf62Z4QLO9K+cm2z+LPXtRkwWMhoL5UxCr3Fj
jYiQCRdF7qfJNV421Wh+7Suf2kd3X7gJ9aqPSgio/5UQC3WItTauhzcuUgWMIlTJHfkEaBtjJNku
JAIkS3Gmh/ddnSkM2ibwHvxhaKARM9BdxljdEHR4NyRhJtzuNjzAGoQj/mJR+azM6j/YdJf0vyB3
cW2qNhETVH5xIuI+lZx9vAhToFD1DZsKCqMU7GYi6gKuRwzG88+qaMlSQvl0jJJxJnsRyS6fBIQt
VjxZsNjV0e5huA3ibtIRU3qyzw39L2dmt6poJOxrayGDXQZ4gEJGPvbNmdp7gvSqtQs/pE+1um6F
rx+FT2vAIQkJhjadOKJFdqu4eJ6GouMur3rfR6skA76CSwbwCh9X90/Bi9Prx0Umf/PivB6snquA
fmwmtkMU2cLSEjCeSCCKJ+QFxFn3zEeOZbdWMJEYsaDz5Tz+gM1trd6ZYGruAiUwmnY3yDy+bizb
O7hQuZ8pAm5lTTtloTFEDV8vcydH+BIt3KRSY8No333LtEwvfCbooWX+FxJcIoSe4T8+JbmHnAR2
0IybU/fj3PxDKF9XG9kTOqkAOLMtoJ3GOGdLtDSAHzWWIFTepVHfyruXg5sSbPXd9FQz0KSvFS3G
70Ctu1mN5n+sEpnjAGZN82NA2qXKBrgwu0C3V/XAiDhpIpuKmWRcJZ/APFUp8hmiHT0SWGKTTLE+
0u3iXNeLvDLn/rodN8xsxy603HYMkuhqOiwXh9KnO4FDRiMvoiBixvtSdnTVREhrJ1C0NpZmqa35
PoAKP+cVY4Z5RWH2ytOozfjI1QUOHZ1kh2fQWEpk2F8MDqR1/ayY5s4hMkH1l9+ESytlbugoNvDr
bgCcTe8A/K1JYoCG+VbH2hGjaN8xXlANe3o3mU6qXAlWzjoSZe9I4era1YOrQsdu100uhbQL2HtL
AACglNhOMmL6mtrxsNV2z0IqX5PhkDiQD8ovfoO1Ynobxqa8DL9j1mPZqOCg2UOiaBGZut9hu1M7
+xBmQKqfabOYt+NlpurWOf/2GTd+loZjh7saZcyFy2jJOl1JcQi9lpLQOB4EK06yg0KaXOOB9o7Q
uHMOmelP++/Qv6RcTv/FFEDvwZeK4VCfOh2W38txcXACl2GXPbkIrkG5Gh4LFnYTuSyzvDANfIFA
A7GuP1xD/GIWoubEUQ+ZuzaxxRw8BJvnQyCbQTnxgTl/L3eZqvhri6wVjFnjPsOkR8S2ZCMEQql5
kQPln9MX6U0zesug0BGydG0EHSNZVDb5XHKVJltDiEPGqfkxd2/BbV+G7/gfhw6h8bjbWCSNIsyS
H5gus3KxtUnzXKcJbWOM+FwThBSNofKCSJbuU1gpdjsog8MBcOqrDxFPpmK1vG+hTCQqa0sJnVTq
EtlNNhwWvDVAN6mD5BjtX+cuaL6Xdo9OJ4og4hEB1ejvgokvlx/rFomKebLLu/xKLA8NMEgTYnbV
Hg/cHFq64iEO2PEOcDfm7rVmqXtreh14E3zOCJZ5YUEbegSyiAdmYoF4VrFTuifoV3s7NacSa1Q+
DLj4VFqE0r6pIIK/kiRLT4b+vjtM/uMnUl/XzMa0oIe+dRN+MFKsLqKdmkZPhL5UUY2XJnWqY7ug
AOPqbW7RAfrqaOm/oIZ2gtn9Cum20ue4iE4HvrVouIBEAOm++eX8FNdT+I5+oEtIObsWKhgdnADe
INLcGJiTppm1PX4KFTvgX+dwDi0IlxV4E8NydDwVpL6HvLlTxSkZupue9MP3V/iwc79fUKcs8T5+
ixLmy3TPs9uI/wVGm1uH1S/0bXmuk0nudvdECumDbfn3R5E3nOjnGV4lLhX+rjC3dA4/2AfjoVsu
1Xr2JRFy4sHD419b8rLYnnqFeFTiXrmDQ2FEawcanQdZzI523oZDy28N/NkQFi7os0OlvNMh8AH/
SC/t91V5aRYn21nk0qQqQPrNFyH6vACQWBohoUDPvx/o9OyOVnRdIt2pfAuHj31+auv8hMoDnnBc
gM6rmvpzLGEaw/z9eTs0kCBu3B6oVmNK+ZEt6EtWn5uZ1efMTj5Zp6CRSQ9a69/uDesP+uCPOht8
bzo7y/FoNJffvvAmBaLkSo/kvx9KewznE0Yg3Sv9Qx0wYX4gT2AnFB8Q7bN9dh0baR8n92kcINB7
VeGj6Hxf0uW1jGoa3vpFJU9EwXWmWbJWfn+F7aS+NkEimErKvud3JeXZl20Y6+C9HSoc4rxMEnZG
tEDvPtQL6+8x2nm+jAY/lVLELBKFL3tQBFCyU6hai89F6r85x0FpgkrearWtqKY8OjJnjzw1UYci
ZNQdBK0WsBTwXbXg4P+/NzxYlq8b8eQgeWo7N/HL1cl6DAP6D1j+EHt/TKG6cYlJ+f7dGhsa2dGL
faMbNDt6VVW9Jjpn4YI+pyFCUaIb9ZySQ0jCwl0Lyg+FSfKPNwadQkVd+a9RQ5qKSGNUOexJNg8O
RaT10e6/1pb1jyQuEAfyO2Cesni0iGBiqTi7qZZABNDLyGUH1Ael6pmjeuk+y3O8Y/d+PJMmIWRD
+kXuPvFQ7GeoR5mCj7eB1sWu9xvnk+dYVWu4lbu8oFhNmT7ubYu+MXb4+gqF3fvyv7Iuf2INh02I
X5Jcf3x/lT6XixBG67EgLSGY6hANweJW5uG8nk46ff70f9dHKCpVipXgR0zUzygu/56656m0/q8X
qg5XTksfSb8sATezbYAM3a6PY8D54D97paE9kBl/p2LwfBztqcCtIYjJEnZGV1wpeps+sgzuxxJn
N6gTHmYVeMqphkOmKphdCtwGWsYxq1uwvSPT6IVjm7P1SkygW3vLKKU0vcDXJNvBPX6Lbk4vtubE
D9uM6xU1cg8lRizO1ESRf3f6WVgIzhULw8JUOYGXAuBw2oProQP0gdqTB+sp7T+oYnmTgCciMUqi
nIaYfF2wemVvOeQr5io/vDZB36GQWIdLvS4UP/PLs20D47IrN9r+XzmoSEPDZvTHAdxwpO1eu/7V
Cly+2MDNveRRCfWnvpUdTx+VHxIQfHrxbHjATtdE9gZ9htQBavAw6Ej5hzCHA2D6uzZ5xgqozY9+
TnHWsGOst5+C4inPM/flpVX3VRdc+qqJ038HCAI3tPv57ERsBrivZnx+WGMLOvjDCzXI3lHMQljI
3x3WmAH6A5pwewuSLmRNooaBkXN5Ed+aPfggfRl9UMPnJPi7bBBPpD7bPww7mdGKnPhi4s8qK28M
hMVI3lg7WqcCEz7/1XWZ4h5PIF0KW/OZJqKQS2eQuwr+xQZpnQHoPE4QNlAfAQ/5Q7VAsZQbHqfV
f5N3FFqQQTcoDCeu7irE+jeejjut5LcoOVppITd4/SoiorfSrVdbe1adT1keiBKAmVqq4k9UWgyR
jV/uNy5PP9xke10e062ikYT5/LYnOK0qxL/8GZHC01MtP8X20SAYJa6Cw3B9VChSrPcvEF4TddAg
f48NCpi7hNnSutzhH7bHPNM5cNUYoiKNKjnp5BuLmvQ2aZkmv3wtQ79EcDCTAFN1NQpByH0RaWvV
N5n6g2PTXjgCZj1ABXTgR0EWdPvWVOaPvWaXN4tWYCUujf3VSlxXDuoapOi+N8LkJlbFAz0ejIum
M1ZRBjL/26sAmSN+2PzJZxGK0WCwydkRQBS+e2YL4gVFG3euGdN2VGOBNpwBuSQbor/aHSfqTyln
mpPy/wwI9Nb1rCSSfQEo3UTq8cPru5aYoRyFolSBNxA+wRABbPeJdTwqQN3hk8b9FoKsk0O+Qgkx
7Xdb60MayjhNYPTZbKQh7sV1NxSHctBYHx6aUSpqX1MpWcMIjWyOe3YVZjkrKig/4BtD9HqOH7YA
XZNdb72VFfBc5FsQ+UJLekEhZOtItwLNhENqzoOvvDMkPYTU51EEQ5KHPUrlYkrtx1B63aoa+fy2
N7AjJeaEQzo0Q+9ZfM+8N3AHKORHOg+nOJczjDoWkjfTHG1AfQY9j3GDhpY/EMWorZTKOCOeN8k4
O2LSrzks1o5AHtulELuAg/RPGIyda4h0miKuXcqDz9TZKQqbUvFQm+rr/tse5WFO97AWkz6ZJC0w
9x7nMX1lzbvJwn71M1Qj8EY/fKjRq2CkAdEhttPgh6e+SLsQHFecSSRcAGUr84x16ZyOe0ib/sOL
3yh2lm+n5fpZrzn69hw6+rSCtL2PUo3iMmoVU4P+T6IfRwUTDRv7uh0+m9uyYmaribmY88xH3ghE
zuZsaxDRHOYunsqPPVgWybNKcmFU0c7U+cSGrz+xRtnFMQzb1GUnmz+1r3VZ9YuFW0dmg2idHmbF
JQ7ZWEd3OHPQ/3azQBFO1m5UOOBcGZMgZbb9sWYM7PokhSacoR3JhlB8zGB9hlyzka8KZY2mQ7rK
B7ww2HXsLUPYuXxdVUOkhIVqQpKu+fBv+QCx+KKj9h33CUFnpFmDV5V9W2W9V2QyQ8D2x8EOU7uN
6fTRfNua1Y0NUjnXgMdAulTYSd/Qp4LQ3TfgOSpgyl2dwZWR6bs3Qk0F6tPLzRTy3rKWMjw9Hswq
y9y1E9S2pt6U1Q84eolJT9B9MjueeQf/wOcxxRXO7n2PG7rve07hJalAK9E6FV5cfydXF0hRaxv0
9ZrdcvQ1mYqdZxZJxiH/p1q6u94Mu1wFeZDtTvqBxwM1R77MPjP5f1eyX9zkNUflN5TRqsjZ/Ly0
CAcJPqUCC+U9GhB9i8zXCxGYdaJ+45T81ctoY6pbtF1wa3fwQwTIaThPf6Jnu+WOubWqhA8OjI6n
YvZLzLsJa70YqCGxdouq6Xkz44kQ24LOUqkKH0U4gkPV8iOCGHUSKBdGKRBZK4TpWo91HKFNwu3C
3KeEfRymWo7OrvZV8mQp/CefYvjqtYDRw1pl0C8GD4maoGYbMGVBci8HPBcasqlnkvSHKxS+fefR
nxdNdURjRw/B9woWEVHhs0H5f4AeBffNG7kA3k2M+bOG7soCFsTTdkaPg/tn+OMUlGVganltUlWb
jXtn2dvqNVHjZrH4JvMHNZV32wWE7mILYwh40L5gqw/Q9jpVME6JeleJj7fFrJ4BQT0RI4ndY1c9
q8VSwLJZ7OSnYWJtJolN9aLDFcGYgR4qToqnPdBgUzuP9VqYiTzMxJAyJKaJPXETv+mtAHk1NIji
qG4ELnXuLfUVplIzrgkYvFiwtP6mso3k03DqXcD4IjGacY7G4OTMXM7O/TMQVHYr3oO97zva0KXT
WUXbd2HkKU/ydKj+XW9ErnFbgj16BUXyyl/U9pKhUX+UPKNp4vXaeE5DMcAHxG42kYxfcerfph/8
bfEI0pBS+7WQMQAwF32VjauKHAUQf2lgQuIAkebjdlDha6EkR+PugIafGKl/sstB61hGB+ycoXsG
7yfWYr5dmo4aDgG0Vk23YR2GYjifKXH5KMdODp3jqoM6i994ZX4CJ6rfh4+SkRzoO0DUbA+GTMOC
bQaWD4cKnasg5DsDym4yQxNJOqmEMIRvQZzNTA1CoQ+wxPJ9DS6kSOdHZz3Elpic30MdfDiM4uvd
T+8F0vnA5PLPrmsM+WNgTjvlJsCHLxBhTt+Z2qUOX2tdMswkk8zGX1r/RMusHS7Q6CnYYpxWNpBS
fqnrBBsH/GxF5aOh1HrC+L3AO0I4qrG7H7RnfPeRO2HJMh5RyGm5ystuZX4fQbzyrPX0FMfICWef
xtX8z7lwRNhs3ZT/Rrf5MeaVBoiC28FT/OauSCxoSNanROxwrbxF3+42osT73t0ZPkWdI90MOd/r
fOwDebfAYFjc+uWkhmMzpe0vnuYX7EVb/LTaWuodGpL1poS3fYl5gsCyE+IOxdFXoG262eifPQ0R
Vd+IFYu3Xzwgvz800rD2hfZGET0Pa8zpu/JFf9ic9Fx8VfZsXIBN/zEC9AjRDM0D1CpZ9yuvl4zr
0S9gSVmrB5DOuWDGGqGyxL4KFU5EcM/p95zfU2RqX91WnSQ1L8EcGqInyO8CxpRJEOE5huKQ0QMj
asl5h8tycuai1OnPK4rR1eVzqpiQPcTuSaVprb2JBTo7gScHH0QmpXObBsky40+/+XXcQ+UY0jrG
nfkQhWk6wljsGJtNd5byCdFAwrniu5Z0D3b/bSe3YAagW1iMEGYose/qndxRhwyhP710OlDnEf8u
5a6KkQ60dJMWLutJ6/P+6aNiX7XliZG6h7ox7XrW9ea33+0Cv/ijtONbM0/HvTjwKdDQY2CYhYwQ
fZH/W8vdIfTEML4Wo5nOw7BwSvMFsb2lzcylXkXUUNsdGLsZFRSy0tX0U+rbZqmdqQ6QLCNL8XMe
hbnJtosig55aVQxddzzxmeEyyS52b5FNEh6xkMdiFRLMPVWlTajuxwvDs/IEyMs3pC80Upi2AUWQ
nkM1pIcW401620RAueDgTmkLp4LWgMddvVOd0xVu6KY+UuL22v/a/qKLykzVbNm8vwd06skqPXyf
Y6uK6StQZ5xC9ZBnPrImKpKFjpFMKlzI2D4Akjuj2ED1HEdY6pSdOpJAejvCRDfrfDYN2VJzMsL0
DX22FSH8o45pydOwdgDNQgGDknWhy0UacpsAVYL7rkjhew/7fbdLRMlr+Ytq450jiH8eX5b0b0LA
ffutORQ4ukDTmEC4HuMI+YXllEPBVaWBqnserQgCY2UQukM6RA8/C7kveSOSykalNJZCnXAa9wFZ
SS67KIqUVV7of1P5iFTyPsEB7HPSKDW7Sn9LGD1dOCSE2KlC5gy2PHt1hp/wOB/X7tRpjfh6f9IK
X0ivoYjWm6/La6c1GRLYm8iUDGZP124ptVutEpbgg/H85ZFzyHEQ/lOcusUH6uRnqWlOTNpVzxLZ
5BlmBTsgf+crz9p5syfqgEIsJUJKL2f1lfWBc7LPCBq8aO25uDT1h/uTJjaANmsiYCu6MZPne3MZ
oNs85/FydC9x8fygcHcdO1X8O/Itnze8zewL4POONf7eJjUbGTrMJpov08DwT5gq/FMdKZd9e4Xm
c3U/WQAhdNxSpsfkJFxeFL3qV6AgmFDekS6j36EWZ+mmVDP7xDk5mUo+GxH6L2/0oRQARjmM/Bc0
8gszdTIqFZrpLzUmXO48OS10dChpRxHQWqseIlfO86lYdmlGEBpS+McAZmSOwH5V+FTEnEO2w4Fb
gT89pcsD2AQW3c3Efm2L/yQ4Ji0u4trIgo4YduJfn9/32B4bdpvCyRxFFzdGSMOv0kLK+Qp4bLpj
o/TXM6Ha7xc7Xw2KM0w7GyvQXikza3DkZy0UY/qzkpl3qYLfyJX4x34YKQerRbKIk868PQSHFkdW
FZmJ63QD+3Yit7iOBPWG11jbUChPlmNPrLFfoNa7Aeel9Y0sDurCF+HfkQucL7CP8eEPtFReXxtk
iGQkNHf8ZPt6Gem8TQdPctAOZULkx3Wucvt14PAQUGRzVpE2Wzlk0jgSluFCafmvtXkWx8gT9uLE
6CdRUPv7+QPmmiOdcbHUmfFSm9dGiM6+z+QBP4v0Z14IjYm+ByZutZcuhoCLKf4VlJvf/nFh1S6u
ljTtMO9naT2heJQytIP8QGlwwWe6JCP21sr1DK0qqPnXlISRBZTocMQDkv5GA11Q5v5PMhyrx+rK
e96Mq0a95NLtKgzXviJYSDSrtR3kkz5j3/BCab0opOpaBTyMB3f0k3K3N8eFK0s7fw0mEJt4U2Se
uiwitlFjQe9QBB7v7uSAASAfnt1we1NGIrscdI/EKPyPzs4xDiVlMnLiRtNKc2bSRquLZqkTn7Wf
P9wxbcBOCPf6SZONPauIjq3mqS5ghkmORbtKb+qD4CW9T+vbyXL1QFQ2hxUmvoUpAGFLZ/TbE4tG
ec95GHiB0OoKmaH42K5VLhYLlpGddK159VNmhyYFr2eH7OSZdO/4hHEyiSuT8H+r2PdNw6HmTFkd
2ERz1e8KTJOGJo7unmG6XSKFos31pM5vKBLbGZhL0edJTPKJw7tmyOh7F3VWJx+AzNMSyz8y8Nfd
8PNuk7WdmghFOwlIvNZcqTRBz5S9pZD9k02tAdGzFn+N+i4vUPvoECeFyfL5PGTPYRjf61QDo1am
asz8z4Mf1ckhStUsZeb737bjlpWJCvXpKcjRn+hcqlepEK33aQ+xLiund+HOxcyU/TPGsEytSm3i
CdR5LaDKSEWMJIya8iLXnfmjwaJgphG5hSt22aibl+U0yFaNf/eSx+eIfTQBrmPa3xSyEKVolfU7
QwW/2buaRG18YlPeeRHmhN20eo/1jsxArE278Yls6x8ejBSmvrYXpWlWktaKzc4bzJ/a9Uis5EAk
HnVISeoqxxrHogKOgyPnMWpkuoEWDqwSWHOjeoBcvCnpiToTPjrZwMF56QRS7p7CadRjV4bBeyfd
4uVYeW4bphoyknc1fyGGu1dSJWwai3FTo4z7mit3GgP84M8uVCq0lzQttnftHFMX+v7oylVs9uBI
EBap4AwrUR4sj/0qpc4FZMsj+bRdnonf5aRVoq6szY4HI/8TVcCt4theyZzHj2X79oG5ey/F0odZ
KGD2vFuBfa0QGEYwJwoT4UlH/Y38YnxPspMG/UyXR+4qF4d39cp/sO6+qXcL50qWQOUIGQTZ07Pq
8sFIY2NwA9ohQE+0j2+pLbHLRMLRLZPz2A/aIVfodTQmZubxlA5obW40mhDAg17cBsUmkK77gsoE
n+eUHAma/+UdWhUuFztqUbqdkq9Wg95RX2vuucFTFGJtW5oWcTR8k12N+3oTu7fMAGfbnE3NY9P7
pjb4fm8Ux+AbZw8Sb8jJn5zkQnF7SnZAIDmlpFEONEAAfZKCEfha5DRybGVYuZwEUmOJaqKr06O4
wEpUn0/4KZt3qUdH1oiOa3nmk/k5hW09HfTo3BrmycuIjhplhnFBlca9EcHTQdcLOfsiPdI23PZy
rbIo41YoB4nH7VVbgy6s9aAiCaEM/Q9ONJNjuiEebGEeL61JfRWdZOQuH28z3i6ESUR3bt5cOKAT
tEKyYdILqmi9oaladUvt89oJqjvOPFRpgE+JVqWlRDh7RWhiryrVW/dnHF3YAb3z71l7y3WfTM56
mVQaCGTf00lstlZ3MnsSYJPSYFuzO1s+MKtt+KLnvmeszlB/JUIVPTaOwngsUMcLr8+g18EJ2eXT
PtM4qJk7cKWCYx4L1a/zAvio3v6fsThUmFdFG8YXDbx2bLzqxUtTH8fZrAvi9Euquppcki/8Xo7D
aUQkBfT5wg7VXDCHZRztDJyxErT3EHKjuiXH958gOxuGE+INB9tJJR7Lx8PyDxHzFO4hobY6FAgX
guBA0DpXsRFPuuiJ8uBbgh69wUwl+WpYM5/kk2XOjfRu8swIRThmok5kTpOF74Fc4RZDssA6LGom
I/Hj7XlX1rzsP3PLS07H3zm92tPMbMdVsQ7mNWkxhAesVYI5JFLoXCH41TUXIu2FUuJhp4JU9tEb
iN0mBKgZ15a7zzxS2Et+NxiYt1HUgCur8ljYKjF28EPxuX8X+CZDaHlTlpSFZE4tajUy/gJE62qY
DK162e3BkA+G9/5f4D8W3SrxfxPexigzpvfvZCOpxgHlzjuRg1/uSjZosdPwfYq/K2kt99AIV3vE
Y8oHBnpSQdCUo8RUeRj4DSra6FFnSmXx23aAp4eeCeuLx80qZo/6nD9NVsVwUZ+kuRbMEpPshe7g
1Svf/FaNNLzuddtzJNsUJkEfyA4JxaZsInv7ydydF+a7sB+yQjeBQRaBXzku3bupxsG7iO7x/Nop
Rp8ZIPCuDtrlIjEeeEFJBd67L47hSqcOeNLHF144NV+8z9g5JwyIs/vsqGeDE/XWLCW3O7j1uaqS
AGFJFluRA3Cbn1/A5otTRRDnfEhf4IUlq0wzciRgWiY+ETRa0We9gFN++WQPznNmfIHnMwgCjXEf
Q3UgUSmy+9WNCFR9pQFVoKP/tj7JTbYHBBU3X5HVD+puE+4haiTXdd+kl/VxRKMdY5lKtdNHNjis
sgcXgu5Vv5mOno4Lw+nsYKbzcCUgBeadwVJsB+yDjvYe9rpfDAYkYIDvO+ATHvENM7qHSAscwrOV
OhnpMeeltwAbsshuo/aTQKEcNXN7DqdMC6NY8sjwoZ1KV8beB5+Ztt7Wkyk8qdkxbT3R10c73l9i
id04QnbvXuRdZFLm1237ULXyJPMQXuyvrO1r4Wc4Pc9Utw/BvvdDykOk9FHaXWEXRj0W8bHA0KZG
YyzLbEXf/UBYBb50n5jRu6RS3MY0Hc7xZP+0EhUNCCrp5J5ASNcGTjifFiWBqwemgr6XhL6KSd+Z
gKadGKA28Xl+jt6WYoFma6GCZ29l8KwHYuW6+7i6BamQ2KXalBQo77uxCFD8b2X3Mdu0aQVjBPT7
6AVTSXfuWWsPAZ5GTaGiekimaqYZGKR9Wn88Fqgxg726rhWypM9mWhhx5YVmQD6OFFlErW7rw8Vi
mQvRPUWz6eX1c/vdGKYYvgBxutxUHNp1cPI9Nf5G+hmJLmlpSaOKGa8ZkRoClUiA8Gk1fOIzfnaC
0lLKNOk+qxH3/Poov3bCbsHz6c8uEqxXhLNeIjET8tBirVfC4zf5SQrAslCiFNfM2zavxyTwvk4s
OtqH2SAj9jwACYEQSVg5uZyqwXYkJKbO9VFLniMpHso4LsDMekt9DgbM/BKygl/dhFmGu5JSXD2Z
FU0mVogS9fjg5e7Uf7ekNB2GJKTIjwOTOEI/AQ8eM97GwTVK7eSQ6XeCvTuOhqgr6Rl+m/7sZ6vU
zYA/p5qBksggkDC9EOCv0zcftBzadLusV6JDjdgdqhgjVNwwJbjhg9dr4q1Kd7eXNzRMh5UtGUFE
2PeHX8pt4YNT2ikUYVLAj3pyPklunyhP/gcu2B/dKXsO8KOB7sP5wlkLcdP8S19AxOw3tDTdWLZ/
MtSGvTuZIomaQ6bUymIIVoW5gNEt5rLjVWajYKN7eR6hKPNKDTDoBUrneiYN7GqntMmt6wBcLAfV
Ndj5TEHq5JZrnIp1MFLE03UMGVGDeSrmGH+Fs19kDeNACoK8Rmf/tyGNuG0LS2sj+1XkDqSGnyEj
iToEA1/np293fWWjBe4d/FzWClsGOLmXo5uv0Wop8GsbU+dauhxzLpk5/tzABtXBrc40zcfSWBvy
OGR8X1RcI9aGYogknv1vjccJCboIAvym1r7APAgBHoiCs6x4wpiCv/oRvFnUkoX2Nu8am6BVx1xQ
D0eC9nccaIs+d4INfwBrJWLOcxWxv/2gI25ncgtnZMLhJs0Q9NzpApM316Kax3ockB2PIqUVI3I/
3FtBUPfTCYWbp3sgs0CcTO5f4UJcpOZjqzwwI3+rL2napMBmEymSvPHhTJ8tVXkf4JNbQlcw/azg
KK2jK0vuLm/Sb2dNhu3n7uhGsUuI1jgaMMdPhWvSXbT1uqaMlgUeaMhnhsSU8sUUESkjY8e7gNHy
LhpiD03JgZu+qdPMd6Hf97sU7mYlH2tgNa6APdnDHVdETp/jTRaC8IRWTUVo5QcUmt7t8XLO+2mm
v+GvrL2A3WCG6TBNDDxuCb8a1mNP8LBn36SEt2HHqH1E4nApy8RzR8Gc1hEkVBmRyERJ5Xlq3uy/
tXwCqN1U6WbmeZilon4z5NH0Akk7hEMMyRyR7NlCZVFPEeQX+/KSkRuP/ojQjIMgSdITHo/LfIa/
oHKMFRcwmKw9p3bQWU79HheVZxwfsTWo1EXXcYYjhUBxH+Ue83jkUMPEhPx0k/+JaJb1Zl11CX6D
hBO3oVLONPIQnLspbiRkLH521SYPVkSE1uSdCwWm0wWsBt+vTz9oUCazpxpIDYCbYElXXn1BfL1g
Z7mRgmcouNzZn+VMDoLGUGZzFbPgeIRaIq3g3NrfrMh8i+bbhQS4OxCXWV3v3EcifjGyjojYoiti
DDLKytVyLTCsHgnYQsEpR24iqEzjjs1+7vaJM/VUNJ6pG7Di3K6A0x9t3t0fZc/WXB911h6dnul+
X8IfBoKlsRj69mGuf3V07Oq8w2yOeKYlh+ofzIG4hmzZ2943KHc1PXq/BlLqe+7swmuQpRcfg6O6
qUjGpx63ICOSj4SmVamr+pIGDOsAL9lrc1ru1Cl9Q5PYC7zRYzEbG0rOXoziA/hCNiQuqQKpTkJg
L7WeBcfn/USf3guWgZSP2Q453XwkCdBz3YAFoj9q0zfmGcP0gfEZXNS9G5slXx9ZcPlA+YGk0MMY
bdkEZ/G9fgD2BTx6dDblzSaUZWbTtGzmkrvJH/2GrGHRloROWmZYOR32Xa1wVNQ3XEJB3NgjyNME
IfBlOqBm0b+KWuaXtFsV/pkObCEsB6BEpwHf7jDP1gI6aKuJvRlzVRi+tZjzSLs+kqz9VyrYa/yz
hwWon99DFJIp6hnz1xmXaj7YLpYAKYcplW2FEVVJghh5MtAtMGuuOmuQVao0MO1IOvTvv97G6pvt
InrwbKlQzNLlc58Jl0mbWhsZzN/DeFtmH7Ovf+be3O/avoNOSTDvzGTU9s9czlK3W8u3AjhiW0Xr
NglrPdDuZ7hMpdrfEa25Fpt4Ohnj6BNJBaJJGN0Kl8a0ZpmFoXIqMiDHoXWMpwYeiFmdZiz1suUy
EDhdpM+ss0C58r4OJkzDM86oTbLPBoVAj7KawzwEQGSV2qSYqJp0kPIU6qnoUHSv1nX9kOyrLlwr
79heQDrZiCLkupxHUNbENACpqcVpwUwFF9qjUkfKhQHBoers/YjAc0ChtRq79C6IULPLT+VuoXOe
BurwErOTkW04nzjGZVGBTFKVPkYc2dXgrJ8IryDEMbh/IuBln2i7Vq4Gi+BDgJoae9w+4+7MD+La
IqIu+KzmPbISf/KxuEUy6X/+mCrq+hAnKnQnEj2vwT3DEK5+5jaMNgqNJo4l1EgApzslYB0KZtzw
UFidqJdNwWAuHkB21dMoiyWU5eDVX7xrbNyEGgh6w9sJuHfBj/b0fkxsEU5iSqIl/jXfEUKb6yCn
EboGm+myoF+NcE07es/w7jtYVckHGbhnrba3VmDbX/ec+9f0iYGQ1JZTe1QyI2lVzn804Z1FLtrb
twA0/3GoHfTRPGDSDaj1A4gQ/LKVeq/Yh3hucHv0rHWS9G45gBAW3o7sbyTT0R6/hBN1x/ElAKKn
o9Qa3nqV69hJoEbOwUuBuvC0JU2Dit9PRoO5hcfgz1ltMI3zSGzNhzsGRHXOh/h3hffCBxlEwlCi
35lB+jkjKd2JMe9SuVApS4V/9gv62ly7Om9kJWgleDXjej1/aY+/wDoR5IC/z7SLP9xduVl2BeYN
l151WfGNHvTvPFrjW9WkC2/YEt1Vbc2p3lqAcBk/eQiFE1KtAwpDejoss9sSjEfOB9958tcHGxot
mEah7lFakt+sy+cjet488h8cYAe2f+qpNBwprWYSmOC2Anxe62/tGF6kBSwGnlxDKO/FVOrq0ODy
syS5Fwn6ynLDSPHoLNJBBmPK/ovBdrzaDqPp3ws0goZIH0ai/B4hPv5bChpIqbLaHJRj42oGFWa+
hHzP+HLp15rmeBF8epQWHDEvat4Exm5fLXrND1yRm0Za9bLBU0W1cIiBXCT2VBJny+/Xj0MQ+uAo
Nk+MgCTqXUenGEuQx+/HjGLsfFNBHtdObx13EAirxjNsDYTl53xFuC0FsvxNxWjTUvpNFK9SL1eu
E5rv86fvqWCJlQ3EK4nZMp9DqtSWq56WWNY/ElWODJG+kykZbH5akDszBxzrL3ejjtWt7AyZphdi
BOLbyogPUdNc01Cxp+hc/vcM+yd4BjlwZhjw5Qxq1GHQiFJqADyRbeJhxBY50VdpLbsSNwa+XeI4
eX2JydTk0+11R2VrWFUFn+c/IFgUwsenbv7cycGhhaiomzv9ALfozUH2pPIU+Om7hb+0kxsi5/jG
1gKTZvrQyXYGaFg8d/UbheM+d3b88AJ7UPtCQGE2bwyAe3hqS+i0CeQa/e47otijRn+VI2kJ9KS3
ZzjTGCkDshl8S8JWXgLORokw+cjk2sP56NuzR77bUo7zkmhQPg+LoHNVHoymKMqZfcDblu6OY5Wp
6vGuUosn2N8KhYXQXvPNN+1Bqe9wBrLOTMoJG6+6go6cqU9qL4+n1373z735jn6BnCPwhvUBIwHU
pTeKpO5wNfcP9hkoFrvd6Pfa5PtE4QNgr8wR4f12QdAKI0fQGVdpZKBKq+keZKygQTDdKjqhWDjA
Fh/x3FwkAZ3TLwuTcOqNzNeoA8AeWWnCDS7Y9y0uS+1bgpRiPkV+0YCikreujEwQHv7NK2DmfyAy
y+TJ6NEa4CkqsNMiTWN1vELhaMlWTIV1iD00R1SJ64gIs2ZypZZIaSf6ut/0Zpn0JSsJPafNVEXc
hjuOaUvBxdHyk1LCw9rUGQ9JhsYM2ZuyamhE3pyMn+UymOSGrd2wKESKfNrfWHZ/kV4mHyhTmQxr
EDdt5T2+xRlQHrIqNiGJ2fUIWmQNlFii26bHUAqvsNqpOKQJF4NWhpVbLOdV9ChDcMHU+f7ANseM
hLbkTNdwSkujwz2XgeMMRjvs12ZHRECgoCwfc3+UQMJQH3ZQ7BHH5AnJNrbGwJEg1We5EiFKOesv
xRJUxNod9rYqcbK3NVAj7ClcXmysPL3BMPOETizPEhcvVNLlUY+HjK1Y95Sky3w43jqjMrTKiNAv
Vr0ihYzwzwhInKWBr9pkTdzyXFIu2qPhxOwrGmlznqvdOcnDrk5PZw3RUNLRAOhBiFWQKyBXom3Z
DjPCYX+ObJ2dRu+U8advYvRMUpVeCyd4le8lwYKsV83PGywtU9pXpDM7z+ByRJ2a/1DmT53pPrSM
BL1EMI+G7KcvVL0oj7skGK523prF3nZD0/yFD7ARey0l9w5TJ4FXZYlYDG7u0c/R4VgosWkcP7rw
vuCcqYhqycz9cAqUYLkWPG5e2CwREso1uVbjKCsnUpUW+inTO3JgiSyIl+bRiOjZsegKRujqTyJv
pQ/4OLwTIcEcKbLIxmnvzP9Pn544wrQY/eh+Jq8n8nr3ScfU0k+/NEfUgfVYIXHCWVeYaukrOclD
y8UD05DEP8PYyJBtbIdoIGEQiB3sbxU5sR3zKlFuvauRkDkXaSIVGU9xw7Y05HojL7FSjyb2OVnE
abIho70zZ4dUEqTIzVY/2AixmkUorcuV7P7iwHzpLVV6YKIHsYKaXYtC8CcKyv0m9NJGBvJ8xjuz
JUq341Yi8eTrOtWhe6w4b6XHrltcr4HezUkL5mrRQFiBGzgFO34niQt+SnMPu8fvJ4IEx4Mx4HzI
eajH1LhQWuaX5i3fB27CHdLJy3venNLQZO3ZPO/qU8MSAJmRAUQkgjc46ovnaPsnzmkuf+uXnllb
d1vHhifxpBlXJtH3oeK1xz8t9f1pjVPZbuiHBfEckg9HueinPnYiC/NYrl4ti0Ng6WgED8ruchVT
zQPEYZD93Lah/2vKWOjXAS53k1ZKUEImUyEQkukIBR+5+lUxTBESYkZ53h/KGHyBr77fUp+yOLjb
rtnctxaf5Hz2ocC/pqbl9Hg2MB4QHUjOjmxctu1V0SZGqBxs/vMfv6I3oMG1hCieKQsAp6J72ox0
KL8O9Y+HeX0JWS5zUFoGRJ1z387vze4wjKyeOG9iqawz/7hvFmSLCeGjs9LGSV5P/UslnonVqZlU
ChAU5Z7GkN5T19g4V6R4Z+bsvSXW5IcREIfQXefyKkVHzFJnnvPSyyUDaPMFzYAV5JI5CgSTGxKF
gEDYJcp79KO4HattSqBj0e5B+xnfeAGqe3g1NnlDu+8nPhmpjz1+bmAS9fXx7wPoWt/XkfjO7VZo
OSAdT7XBzgSdNKVsQ5J1tY03y9+9fforzgfqqBslMJl6wGkJHNByw/5mDOD5yof4q6ojHd1TmLmW
tb7U5jlhBFZBOJCMB6IvP8opQJ/AMFehb97//OUKQZJwS0T9KfaSCXxr6rESMmRVT70YQF6IvsZS
IiMpY7kToAFiqicky+3ucQhQxizYzGC73nrmZUPcPzsxv/wnBffPPx6LHMeG/rM6U5NMfmG6jctx
bdfoE1qSQQ7js59XxbNFZlJmJ68ozT+c4Bed6YGz1ntianWOYgCQ3rjWJCdRVsoSZM/TuFNCA+3a
pcvjEscCnIXqdYD3KNRJ+6VHg46Bh2psEgu/hmDhC5DwYL9rVLXC2DEo1crshym/lKkEj4LWAulv
oP/+qrJZQM9fP2rg2MRQNDR05rMDenU+caowK12Z9VbS7MFzSceIbOMZIjhd9pGLabRacC0C15tk
z9UlVX29xs9ZQoof+YNmmZ5BZHx8hR4gRzVr0iq0UOXP+jaHxK+jggJ6iK2kwqXhVPteOQztPWyV
EKmavx6tLo6WnVeE/iU7arzcDt3c0alSA1B1yDiWVbfwuaNn4aZbd2HW+7xF4Dm9ZoMNP1uJv2Rl
/QmRCl1S1uOLuNoG2g2jzJDZXAd/mo8XA2AzIyKFg8E9KC+qk2puZaRKZxYZn5Rq592aIPmq+322
daEa2CM6RACFNqAZuqvwWVUIpFqIxU38DTly2t7uXSM1XSIwADlRPk/NgEB7GxtqAe+Btdw5nVv9
RivPYbHWUJSeaJIM0iwBIzXkb6L3PaU3bUYqJdQjJq+Iv42888fzfshMnylcGm5tJJinPZweRXks
28JO9KoWwbpZwaVbwxQKq1pugnOu8rITPeV8mVgb71ikmSPpS9zIWSe6jbdcgEC/KwmiYTzxC648
k92CCajWNxlPYAOzhym9y2RWrynkA51JBzjPnwSZtmjODbB5ux7lm6vDl3tHcjwsmpZzWT6Xf5z5
8bJ8SyJyWMRpLvZSxzdXFhgvgWnhnybZ/hLe/CdbQDEzb/VyKEjOOLHAXYSglFLd6KhgRP6TEelJ
gwWJylhlZztIlo3K7WzhiaEJ9sVzAcGxz6KMlqfDEk+DJ6a3rMoT2ugFgEyNM1Dz8NGungHlwTk8
Govd/6CEO4iPp0vgslezFPvlGp/FbdOMJu74ueXmlS13chIFNebJ74lOD/Ltl9g06yZBZP9Dqct5
l1rfrkX5iD++JTz/JmdhVFir10nyzS8Xv1DHBDstj21iVYdM464LTKrFLBWSrkI81uDCspv3psy+
LB9l17rNjl8BU7E8zhlFjQnnY84R6G/d/RtMIyjf5pr5dM24XcmZM8BGi6t7tuq6WPi9bkMTsneW
oPJqB3kUn0+DJCyY8p9Zk1+cp7usDfVi+Db+NHlHFStZ8f1U9XAsV2L0GvboXKPS167K1evZmweQ
AnMfUJruA2IE/PB8rseFNZVt1LYxPIPZNSo2Eh6YIWQ7goc2bmfcERJ19SErS7YTAYID3Jjlg0gv
K0Y5baSt3gvGJWtlvTiMJfnj+O9/752XWuPH26r5Mr5oGRQkja1Kb7kYqQcGh7Dy0gr00eKLn9x+
1TU8nxAJ2K2r1DJV5a0i/rFAS7s7DuZtW+jKKUkISjrxiu8W5VSaArz10Ev2ixoUVHzWYpBh7SNY
JEQJdKwsRoa1k7hG0aV2mepV+aDLQVSfmLM9BPukI6jcy8QsRK+q4yY6LN3JycSNt7xlYfKG4qr/
Lks0g4ulN58RHYpglt8Elbs4o0C3A9ToXt1UBUjscVgBng7sF6cPa+x6Y8Int+PFuEya7eAYfK45
KXZebifRXb6RTgC0vEQUxfSYeK9GtZxEdiAcLYzqtBW0NJHnJgzDw62OSuRurx8wEYCg+VbkqIdz
f4CmXhjTzegHKwCdaqzrz1vEoy+VrFcGTyuidwNGX+An+Clzi15Go16oYYvLPnY5MtTHgIeZjBzO
NPnuZirfnzpluh9tJXDOmSjRbbO6Xz/FmS12N2MhccrKtLXYg0rim2RLHtFqI648Xgx7J+PnZ+yx
RtQVrY499gRZ1GQ4YZuuxnpfwtXmBClzusL3kp/GNHUhc2dC2CFWcJevBejZWNsxgPFAMH6E6nR6
mkfCCWuJ5gSDjPRXHJE5zRdXTZUd7kQ0iGMehSH9naLkfua4uxQaB+7azBCUch8T+blDAMykasOs
OtRd+HzC23BHk3XKk6nizmnvZYym+9yJ3DvychRL7gPlHCt9RajEpbFqOuNsVOOoN7pIfNQRDUYx
zlyGZ8IDvX3B3bVi4Hr2weMH1yutEqUXhJIo4cd0VP9ves3YtlbaaYwRRxyNM6ujhDnqgwS0s12w
TF8kCPVUfU1F7Qjs+Jse5a7rFIwL0angnHLsDbwe4djsROz0zBDwnVexLSqziVghVV+kwXDF1Aym
gbAO6+d8ZriO8GdNGXZ6Hbwv0PzKvSDpDaxw8AS87wqak0RqwRVEG83Wd+6pn4ivIdYtdl4H98QL
QSpS8+7Wso8n855H045TZiDQ+Ia53AYHGrXWned1+fJzvg730LH0fVEB/PFZH4fJw3ULvR3ItPKo
uTBZBLn3G2yVzeb7SoIhtw6PTy0wmGSXWC7WVEl1Hmb5xAxtBwgCtDEispBQAGsEPv9WrfRGxPa8
SPwZRqxhSu7bCkj/jRuYijsI8s1XHGEv6GAqBLueeBNEI5H7XCfUBEFH+eEVxxAZAHoIYE89+3E6
EEJPUtvE7EZP86WkqzpphPrtUr5Qicnyds7Lo4cKe/H11Ab6bNUvEP+eFYS2+gElqoRHeqS6tkta
UtAbv+fMmMkXDXx5OipJUiPdifm2KA3FvHaorYasOcZGSUl2EDE/tRNoMFW7ZNOipSOmUoWXxnwm
yCXuMkW2J8TvOisLeStSgSgn1N8zxlq9/+F3End9UAKMFicx4lFtSkMZX85DeKSt9+JgGtb1LDmC
/BF05pjKvBGRe6rbUqf54hL9r0xTTwN8ETAE3lnAQB8dU82z/qg5+NTsbu4Jflqq4lpUjoE8YZ2E
mqjekoQkXrvril8IKpVmKIQHhKgcJEJ+bdCt+/SxLBwq0wt7YlkQKvVEumpL4xqxb6HUvUmzj5+v
zgbI5Vkb5T7V/Pvkbd72S6m4FjzwCr81GIhrhqwrc8ZVAwq2Ynw97BsNnBtrUOc6zrBsHoADIZYv
BtZ2+6GUVcejbIsrYJnaFZOkgdXdAQ20zinJWlzhRuSWrR6C5XzouSc5F9h3bm0EzFBhcYI8vSNj
OHlbuFttTr1NUgzE32TTMExghWXKlTotLfraiY7YwjKGio17Alt9HDrMHb48YUhW+lt1yvyy1aNH
jIkSbp/S2N9JhFP+eDtPqRUNtJF++hmyJnjKLyvqF1fHHqcnSTYgsFmHP1JbFUFnvPllwhkcd4J7
30uALUxnDnDBmtApitRvmz6XftLKsL/9GN9Y7eMaZf8wFvKJWT626ohdljk8fvYJSDM14SwV2jl5
YlZwLwqYTM//eBeC4IKQNg3BC8pe2l8pJLyensMoq+UY7BAuZ9Ome3OsM+yH0dGCy2AbS5lEkktM
/0c54+OiPq+IjZQ2iCfqLwf/366mqhDEV0XYZn+i4FwW02rvCMdurfYhsJwIFzPWdShu3Rr9XAKu
cVQSz+YJtL3gfEq74EPABUid8cudc2y5091/3NMf7g0ndd19ayol2GQXGvmSzZNWST+dUW9JUqwZ
xIV+TFOSKg624UllVJJ8HTDegOm2XNvwb67EV+LgV/T0JeAcizmar8Q3BLu5QH0gfYetzpkvbDjz
A3X0qKntzkyPlPL0wbDY9kcoaWir78xYvUWeRmoYxgg7C6X6EIa8t6CxVt2RO+KLVrJ/CMJoW8A4
vAea+d0HjfYaBVowRRx+gF54mA17EQeg9nIC9wjxy71yTMYAb9q5K4PanquUEdjstXgni6oimdX6
7ZTJpdFPGCMv33FNdRYDPCLRFLXYoytEkSg3QUrDqSL6WvHn+UhSgjiVpsB0+fbM53jKfuvOYW/y
K/0eoG1D/pdniPXsdy1FGHXoKAHz+mjrstBvAlt2AetZecurOzCU6HYYwPQ7Orvv+M67RPpqEw3d
FbLwJb2dSxCiSd7ZMec/hrDnbN6xMewcuCUHXNyWeS057RvZ1Uuw4Lmkjl8qMxnl7D6S9J/o87RN
5+d/QGP5+UtujIRYZmdLVFac3QVhDa3aaqEAI2YB9RJCKiV/J/T7Hm/H9o9zqv2dqm2TVvWpZGsW
JUETcc6/XYGbBRNUQ3hpbzT2A06xkXiKLdMac350yvDLoRp/qp+QyuRz9ba5/a3kzFG/jLP5ptJZ
zKkXaPZujKkIO72IxfJsU1L6Itkg2IUzyENUE027NPOOckHFOqCOYlLfDTxr30zDJ6lKrmuYjqLb
h9ozv+3tV4bL2kE9eLXZGvD/j2yRFZQQF54H/5x/nRB0vJvvKK2JIMKciKWzKhGo3VHwVgsdgsND
Apr68XUj4tFVd5mnn6WtaCBVwzlXiTmc2AUC/11antVBrcowYf8Be1T/06sxDZFidCP3gWLEhsYK
H18241uMk/js8Ms2hls51zniPVmkCaTn8r+6wFmuj681LqeStN3fYWYoCLG2nRhuPU8mDgiBu6xw
S2z7f2HF254sNmpijyScg5ZFI7Mbk/MInnIoHg1erzsGTYdCX6wS1+MSO7LK8BIP5beTThm7/v71
nEq6p4EudY/0q9zDMvAnoTbl3k9oOHUtY8j1AIakRHQXI6HBXYIYC0WV+bSe+rTXsJzTk7nfio6c
RZ0U2I0klahCXodcEGo4e7pawBllkoV8FPztJnabxXerWCcdmmK3De42LQVgqkNqbDPhhEvFZ374
FGrT3PjcJVZNDHlf4GY0Js+jFCPMYxNplo8mP/0SSxc1KWd4DB4h3nyYGvcbrmG81X71fCu8Tj6P
WbCu0xBguwC4Zp+hUY+kCZPvqic41kGRliMXquhvhmOFBmaRDKT5TwdLnlc0QbNRbrjZnEst2O0A
cDPxe3tok3tZuWGFtQ0fGSMKIWWuaz1ydVdFwbozEcMcgMiJdAwmS638s+2lhg9ntecnHsiQMW2n
5okS19ZTR6pLOMGuiHjk+RvvVmL8WVNq0kuqPSQ+G/7FU6VfvAq2xDD4bwn/GQzH4BpXKN99aeih
mXqr96bnF9REvwexh2G+wz4X7iSDI/InUzSQWA+UepxN4YEM2SGi5ICJNtR/lyerr4usvYFbOR2Y
eX4Q2cnOz8H0FOPQL9Dv1JJll5996yPIP1cKZ11B8DBK1Q/AY1J8XvcjS4xJhiUwFGmrjtFqI0pt
kWe8IJ3QS868/9GoaEaeRtk86Qdr69qdZ/TUZPXcjJPUpugwTrqBjlwBXKJ/BGE3MTTMA7GyaP8L
fPizt/+XmtriNNiKJTmRc7bkkRwiUBTC62EEgCg6p4MWou9wHzB5L5f5tYdpMfQDCrfzTllaUpLM
5tcmUBTKEbQ5INVudJ6VXKekD3VF5PkzLFK42/YkOan9i6avJzrTAYANfdYZgBLUnuy8Qf9J2VGv
ohLPBrTS8bzXad3RbNyo0hr9+BDZ+FPeuQH5iHViUxk78nLMcBmiXutHRMSdpPqtCl77w6TM0K22
0tj74XgcJZc/myFjF/ZeA4LgGrTEWBGEk4ovNXObQTiojom2iNw7zX6orOTsukzLFCOvfbAlY8eO
anallGdRtE4vyJhtDPliCiMLlbsrrskJcmI3XXPKfDzF76aqNnGmaGJBEHinJ8Eq0nFu7EOMuSoD
WoFyBdvUunvK0yHD9PYaxD4wqbSgEnn803Qn/UHqUWltMeCTNy7pl0GeGBT84J6BxV8Nx7OgcA/q
gbHcc+fULqEpAkMWIPCtLy5JTz8nblAP9mQkuFjectD4tuvfKx8rxA6GdAJoWFJAvqvKlh528T3R
xBQwx8WrJIM89t5VIq4/4MyRRkcNKkAG8OaQ7rOAneDWLPFvQ5M/y8hc5TLhdrfCvFYYGTvAKrWd
fewpr1UIXlYZXVFULNpn8CQv6UxBInxyGVp0WokVBIDgGJjIzpkYSMAYkJ9v1m1LcnDZ9E3cKrNr
MqRFzFb+JZAd/kUCu7SjE7hIWYky4cn4oLXLDhtpcRQU9OUbhuPmED2/Y21ZQD8QN8LWC8IGdVm0
rbgxhbCIZxvmgXO1Or6CkDN3OpKTXBtW80BEpR7tNY8fxloIV9Wf8FZbU7TL/q57Yg0KKNZ09WDI
9GoT7Y06HqIjldZ8Z/Ze/8YWnCGBZfoRIcXMd8y197L3J2Kh4DW1N00aYsKlv4yREkxqOnXQp0AZ
/M0qH/MbfxP+zEvDH00FDGOW76A/qCXZ8FEIMPhNIlsd32XCpp9idQUrQMYTMXDM/YLN1sK5SSqD
oVFR0F0Gr20KCshNUXN+xF5uQ0Bzst0wRdRq9qtCyFtF1llMzVaqOBlRuqpIUiAg+h0+UOgFolH7
quJ593e4lmTi17ormNfDSoYc2c39slK9mmFOZV+EZM8najJNzgkczWTdfZcOHhgBRn3cPvH/UcTD
mynkpRD+1dT/xAzg5ye3WwfwGFpHe573nyUSsrQtEOUOUP5zK4egn7SF8yFj4Ezj8l1sAkcsbndx
vObDyGxK6pVIIC7N9EwgUxle4J56MWT11DaGzyeQ5cRQjRQIgRKgYTf9Nw+S2GnyZJLXB6Mdpkro
yPJGEsFh6WKzOlGvk2GLj4/d1VIrN6L6W7gD5k4zpLZxnWhzIOfMoVAdsi3iANBQZe6GK0E4QK1Z
+7fE2xSenY+3a1XzAxL3b6Tikd9aphSHE15L2wUvOWyo/Kc5rPTVWBjJohcrMiav2KzSJsoMApHq
3B7S5lhn+tJYMsmFLnngK4aYqdPy7+owd4Psl1NE0JqGB+K3f51e8AhZbBY7W42vWXsNQlvZyB+A
hpW52bpKiwTlLr0oCJ3L3fsiQZq/v71dVO/UTNDJeo0Z/BNyhnSbuRjRqJqYynSV0cEaz+2AbTj3
6SfU+DBbm/sRaC3/X3CAXXagWiYhtSUjOmocD9JpPkoPC6bcNIaTruEqPzoUDY45roBARN+q+Cm1
8NIdu9aiTINep0mzntYtFuDlwCfBSoJyavtxFO2evKgGbWeqgIkEAkxO/D28c8YA6U6VaDBM95pD
VJXSt62xOb9fF7B5Mr+0sX0+xsv/D+NHL911ek3Uo/cfyuSkco4wABHUYnmDh+lyBSz3a4gvoF84
4rwH3TdONK6nsHJKpsDXjyDJzlQwjGnjS07dxH8sNbeEL5lrlqfEBZJ5FwgfmWtUQDS9Pmm1lw25
t6S0+JAwmtyGASTGp0M9bDJt1YpujOv7doQg6f92l6n3WdF1R4o5FJwEk66lL1XHFYz6+DqwYOXu
zRCi3iMXwTLC3aQ3S+Gc/Gjk+iEkwqxXbkeqyaC9aAE6exYTHipEBEEb3IIvFHJhoPSBqF2kBiSp
C8qHV+j9vVSwfKiUAHHsd16JtGy0RhsMHmcIcpec3/IfF51TytXal2YSbqvy/Y5dZmnXxmHq4+mu
j5RAHvFa1tPaGVPavl0lHwYQ+IRrlonYi1XQ/W0mB4HzFplivyV6a5b1985Iv9s6s+MSyWEmzwik
uCu/wvayzoGOeFJnto8dunnWL7xocG5WolozJpiiFkzPZwIkB3NWkvplqPRK5UqDov9FDPmJFUR0
1dAnC3vfAZcNxz7FuwPiXFAzxpJ9z4ktkleC5gQV/RCiVPEcuENFlvECE6MZOCoLSophZ4yZr4OM
mvUuCCmzxwMmY+UPcA1Yyz6Xra/5DKoNxm3xlAUyy0dL4XUc0qQDElzRUH+ftT+shpm2T31l8ZFL
s+v5YcRlYWwSdvHZby++TZZbabnfClUynmdDMYxdqgBNY5y2zBB4ozCH3az+eENBWuUwOyaXxhz6
xQPM+4JgD1ayrpZ90JIMVCL2oDkIssIgUarMFlMRAXYBgNseUQcOLhVtpqEmaJfA9mi/EreD1t5g
lWcS1CAwABIEoU7qtLTjbTEIH8e1+rglvhD8HUjIyqycmhK/AIoo7LXUgHyGXfnVGWsv2YbxONGi
tnbmMDjXVVuwmRddQBbXK/VipiMkbMtLfXV+RcksVcmzNhrAWFS7n01b3R+Wb41vY0iuOic9Wi22
jGMD/3JNvju5ZDs1DV7dmEffZO+0sYPhNS5DaImA2r/k+IsRtK5FUfUrHviJeExZgz+djgiAATY0
C4CbvuICMd+Sr6KjZfOkugd3ArLx7STWd8N8iydRWuPmRx9Ku51wOT5AzAm052p2IKRsDhIq8Vc3
TtPE2EFu0qzPMXdCQ3VTdDcL0Hg+5KlCBfq56/JxlW0ZbbBy/qAnQHbHOo446HcNjEFKI5mW8yJ3
2TJfJhwXgl2kkpbNyQIeFBi9sxmgX5NpDqBLmfdB1OlzheCarbC44srahsNczARIJJbIp2zfa+G/
7LHuC3maH0U1VamP71uQRs4Cyn1vf8JfoHUkwvLq4L7hAZs2nC54jR5V2B+eRawf/vfZlLSJcoey
VmZ6kxPGuXWLdQMk7wGnYkcXhtaQhU3gqqCeCIQvY2HwAXxFEvFByWwr5p0vdL+/eu3m6EzmbiOI
oaZLpegl7evLYJzN5UeX0zdjvx67CfJtVAFZFIStn3DrR4fqbiu+U3wzzYqXjghtJcrFMA4E+vMj
wa1uqWHjWkmpRsmsJzH0TjceaHa+IybcUvQVXTZPspZFFdwHfjDHgSG1s8nCVv2MrUsYGZSTPLb5
4qtBiZApFOlxanPDkHcjzqJMwJbP5uNvublaL95khFtSAw7lGJ6VOpcUac+vBjV0gVLXyln6e/r+
HBVapEo/MOCP+3wcQ9//OTdLtymqM/InSZaKpoSfqUTdj793iWDt8EK3i7osbuCAHp4xJHC+rbhL
0crxAXdrqKnaGwVld9gAkTkguOUC2Kr9RCJMRKdFexK6KN+1RByrSF58HOAXNuuNlhot/R1VJcwH
qgxntPqosq+4wQW+8iuENvx6roLFJQYmTrS1FHSdUWOCaxXp50WfH8vQOEEYm5L2cfMY3a/KntWf
xOMwN94A38U2WPgGatMOZ81islS22IkwziD0AfDUaV2ysWdyalu7kmJMLEUafcXcw77NxF9hTjRj
PlmdITA1mevCOeDOJnwqg659xHMSybLPpeuReNlvjkO7wVkRJaGu3jI8Opgsnk4uh4iLUwB3KTiF
T6vgXlQUaxrnKdvWEhQUQNXWdInqMxGeqoSkT+tephnmhjHv3pzC0maW15XrQD1CUjHnEBbXAEv2
SKCJkICAhmFyO5GRF4FKx63nuJfqv+QH1A4e+ANY/3KW3QozEI4zJe1dx3XeQkx4kACbdDtd+AAi
Anu/jJMUU6oaw4EQsPxy/EnLQpoH5eEU3+wdIsVwgl+jcZC8WqvCBcr5K2bAXz7ZbK6QzI2LAXyF
ws5VF+6qDzK9e0ary6KKMYwLwI/tYLb6tY7UV0yLDm5E5a6tJWzx+6mTESDTQvqsgSLIVOSKeRTA
fWOJzXuD8BR+3qnAqnL9qYuNkgJ3jWL4LIzlaFG6/KGo9QEYOKW9zqmOWv5nFNg/LZrhDJgwEPAa
90GO6aRFoMQ0XxkXfArglctBk3ADSrXGpjaHjXZyk7DlMj+QVPGHK0F+M7iWZzYD2AY26REDnYyE
cArUTqYWxIF1QlGJPjYbWtPdxMLgWhaPvBM2S8bgtV0gQq/SFTSD5YJktV3+SFGskKelyLYsh5pL
M8tzLeSkYyjTa8fhZfNxUBXz0yzIrsR0uMP7aR6yo99AGrnSENcjAirD+mZymcTeaahSglsV7K1o
8PdqwvFTO/rO/NlbS8J9mEmVGJmD7WURlIw9b88L8wiI7l9Ng/FuomTvYD9mw4yjekQuyK2BygUU
z7czXGPYCsAshjcKLEMF5C6M4rIBJNdAJYX1iuIFefRCiGd8JQtvlCQpdF425V2CPXwvWdlDZCqy
dRSW+y3YtkZLRHiwUJZLnlXCVkSCf8masy5r/vPuwvXsizfFjVxdC0NK/uIYlvIh/+JoeIuwcVFJ
oRGwAtLf8D/+YWPMOq646SoQx1pNLCY9ZVAdw0aBmRAjyGr7tQ4JAjUqWNzNYe2Kx19XE+X6hhvX
rpTFEQgcQ57kY6H9XEor78UUSrFazDMA8SLwFCAtXcYYnos//dRFm4jdzp2QWQOKUjF2F/e4DaSL
DOvnQK/n4AKQmV0VHQwIKm3gjZjAAwAWlJxJuTSpixn9ux3TgJQKaPs5fEKENGn6V4jh6aVUsLPc
tCQOiJaZ8hsasfGqpczCeLG82lXrKVOISSsXK1Iuwzq5hFH4X9yrj3SEJAOFTy6eqJETxUgETdwi
jyBp7G0JpthP/RwUJc7Kj3w4kG0Bdfvaxit5XmrMeWMmETOHiQjpZ3JTC2KIgoO77CP+WRUjcUv5
V5OCG67gP1WaxQympspVlENr5FCwni3JL6KTRi1l+3K3ZgOaiP/MMPrsSyNG79dGl0pb8fDC8Zai
vy7XqeGSayDxlxoX4QEkFBXPKPQW+bo/BypSq8T7NrZ5bnEXUs88vtKTb/MfLGBXMPU1zayetYtM
GDNGnBBS/nPzb0LTlncSwGDDDCuTSl/XRzMPgM21oYG825h2I/urUiG558ikXu1QiObKU2/rhhE1
rV+s3qOgyh+Bt4yiVOXoWBJ+SK+YfyCBmlkQwcuCfOLKjS3q6w45XQauuAmSbNmCki1xpFCedvuy
khEixG4ApRmqMHPr5klfJmT1H+z0U/JnHJ+vpEJ6CFQc/OrVO+pTFH8aHin/zypgoBH4JR//DIGU
DHsBV1T1HylDk/jbON098Em04X5UdisEbj0UKZevtCqaUJuq4Q2tbA8qsbgbOxbTGF3wEWK7VW8s
tMMHnQILsY7u/pbDsubrM+areyqIKoQ3cJCvWfYsFqe3vkDNZWLc91ko13vHisCDm0jHdZNdae4h
4URR3+aDlvYw3QoWF5HJY9Z1MkLsiS25GIsNu8F8Q2cDsTGxxiU1voaacaQIY53VM8z5qQOyagWz
+xEYAgiEvwFTCVwFieptudEgZqeWt0jztXoek2zBl6AbXDmdhhnAYpZ9yFe5AaMF7vrXm9NB3fp4
2ehv99ZOrrr7teo2wzvq1NAUHQwTCx3qZjW39uD/1Ui47+5gu1sIOYcgiHpcTMRVR3lksp6SmJQb
kJyl8LOkC8o/WamUUz9ujVLBz2+dBN8uW8enVEQAE3+XZhdNpyJnlPA6poDSYWwit9nCUNckxQLx
wca9fkQxD0xHSh4U6+CL7a4GGQSo+YrKmVGiSVOG53VKWr14cr1TdOyNc6DJ9C+GE5sMcaieVUrP
H32+1Lyqy8Unktx1zVliDAqG7qqJt77BRBaUvoFsj35/szYjLZlT1tyki+VBGrjO4e0AwqbowfkZ
l4eLnRyMq90bpIT9HsPmgnTIk7HtJj9dTxyq0hxipZSiACTy+DaEwHnhqi7EcFTnl2dk1JiYtpEO
jQ9/Rt49Q+fgIHBR4gkfxB8/T6vhtH+MYgnSEeISacxpM6zDpPURCNttVn2J4YxrZUD7b3Zi7dp7
O+CNUttPBMtWlfeK+W9I1HEEp7YGoDvRBOpJqdunyvhG9kmdgFegKANnrSCaGyuoZ3gSjcYmVC41
drV9tAWOgyErNjNVXyM43SrMVqQiqe8iEuxzkzxbBa9xvK6dOwfRVz16E5M/M1lsuPGVNBwydrRe
vyYBqeJ7VvhSbrd3A09+C7Lq42IRVV7biyQwBxXHHHp6egMrYc1ruWMljIZMgTfDIi5/rHKzuosm
4dt0yEeAJDAhd+mGvSCM/zf7jTBytc/78t6Y8Y+YX0y1I5i5dBiXF5zhR8az35y2/khPbJNxAleM
QsKKFYp8nlLa47X0DsGB6LYiXka+P4frv3eNG3gRDbpD4+hEc0l7miyYIBuQDU0gdD7vOnDcCpoe
i/xzLi/nQRNbMoBG/QvvUfqaIgMmCXmK0hlIhvktmka1zbBBJHApHVuiX4jTtbXiRwMRSYtMkiM3
S0Xvok5MlzAOWpa5dcnemvOYFxyxILrLm3Q/miqJln/oggTcfyUeKdATUu875c4tufhSun5MRI/W
AUjoZV21lxhPNmDM75Y2Jkx1io7SdFLseolquWXmzc87a5JmCOI7iunxckuUN+bwNEdZoVR7H/pd
TqLuMOg/Lrisr+9qBwFrfOC9Y+WLgz8CqA2JsC2v/wHD3LQqUBn03rRR2AelK+MA7C50KUgeJskq
HxaGO0R9holgWYZBUcjDfWbhSOeUMkRq5GJIgAX7xu7uWtg/kgstDf9pjtp2cs/WraH9OdHmGsBl
UOSrTWktNDm6g2I1ivYWEMBfPH8xnaEXf3xP/LqgEPR5O+y0P98SRe+5xHf/tlYT2CztIRmVsJU0
ZD8wtLwZ2KbgULClOkGWI3m+3r59AjnhUNi9KqZCLILbFD6hEko06E9dUb5lUxl9xLJQlSdQbj67
JRw9KXfRfJGIkrZfx0yGY4OddnhSm4mJD9kMMhPqOATo1ypYDAQF4nIFhM+n+rX6jFaCmlSF1enH
gWQ4VuHrwK3cjsnpf6htDp4A4wfNAht5bM8+3+y6fJTEFeBRPD/KDZ2LezD/pLL5yMFTAATGiLK8
aTxqDN5GQlRpsSQw6Ykpv02CJuSz0c7aJgYqbkgOnEwbbQOIga8Dh2tC0weXk8nyywcQsq7KI3Jb
JqRo2hOhTlfbJAqtEEvSYc0OccZFGPqSE1pd7yF0kxFXuKkfEPqU7KMvkm/fp7ZdXtQb2nIhleVR
wuITkAtfk8uM1kR0xXw7wYi9vK+DBRh++5rDFDUYYs+t3SKxix7w/btkGR+QxVhgh7X4J/BGEJBO
b/q5GAnvGdwjHV58j1Uu3IoLg+0GsMYGIdkwI+BWqgsbDoDZlSzWWYlnAWvwCLfjGRx5pnL5M0Gc
Mh3Tk9NctfWYtxrVH/ChyawhOhQQ1vzsP8XBo1q620igfOTstwYN2b359yAwjxK6UpOmGrc9/aFW
mwgu2o/4FcE4Ll0j5p41q9OmnU6KZ+JNKl48Ri8SNZ/CI77GA73fIndYR9Xani36iwQhRd3ApEgi
BWDJ/3ENwo3bDIPgYTA2vM/+s9lmKf+Txriww3e66YNa9gA2HiU0KOIdRgz+znu2BracxFa5Q6Rv
tJLMsLcRt+dGkDoMQveHILwUcJn+rdCNt0nlBdIiQBUsbEy4WwFGlpIcVYUzEDORINy3eLjZCKdU
t2QNxTalnTgW8q426YaBHmSuwLRZjG1ylnIzGECJly9mo4M4gPknl4mQm7FOlmynM5n6owaZ4Gg0
yUJ8q97KodKPBmHgk0bZjWtLuaWYtpD2BXv45RotKs6AlRx+qmxQbfyLf2ZRDzDgW9iJ5uSX3AnN
mSoRtT3/KV4az7s9D7Z+osOTCG/5oRlNw5VoS6TaCVMGE21vXGy+7i2l3jk51hzzSitIlh7CV0Se
wtqAZ0XrUF95D/cHHe7jHczmn4frE1y7KfNAzVVBxn2Lz187Lq81fK3FOBUJcsOsX9YSE5+CM+Kj
eqaVrWTazG8SYzbLQmbvyQjCnNSlTfZrJLIkQQluDA2Xz8verEuw4fs5OLSipb5tG3AfaxyBGQjJ
6+8jMcU/8slzyWja/zXw38zuJmEIZ7GlQdkmmgKtQT9iKQ57gkqQEFZSz9qNgzCl5Q/yYeKIc4PQ
a13UmGfTtlU1mSwwMkSBOeDzIRgDwOJ2dzWjNcISdL8jpk1gEnW2dn2TfpaPHchVeXI9c00rZviM
Ip2temAlbL9X1io/sBQOg30VPeFcuQPgIprxFaBGSoptbYmbhXGPlFYs6jG7xDg4kcX9driXNMNY
QZd3qhWs3jF/TCSUlU5D9teaZzG2guQBCC7JRckVKr8nKUDqJt9G03sngdHW58YONlKJMyVYe+MK
2piXAfrNVKo6CjBH7KLrHqc3BkNL3MlU4BMwDjtiSt4p7rBIK+pR7j5g/oAzi+gULsQ7N5+1bYbZ
Dv60NYTI0QXnJFe9fM2njSp8fGP45buuXAYT99s5CvBSP9pKzqtLWpafedp8gMKDiVlyJdlZe6sk
SJQmvcQTZCn2cccpEMJzVtApyCpwtWpkBFPwpNLkn52JgSuxSrEJ+++bxj88RTgwQnJvbr5/14hC
7YaTUx5D0fLxIQXRYDaOAN7GgkOamAHDcSl5jmSoIo2z94Qb6x3eu1I0uy0Rq6YSOrKg8nPi1arK
hRZ42ESfV8MiCbFGXBK/wKJxGkGlwyvOGLH7udO4VTMW3eVGj5b6TM23gsV2zklxlXiMAmn4dq9A
o1NZsgkBeXxEU/yslPpXqOJCDzfYvDyuGiQl7ZNH+CafxhY185oU/IOLdhlmN3aucCrtsXYbAwix
XIDEE52ZXgeRgHqvtxHJFNLRQqGGA+1KlPdn22JbicM2q/ThYzd6QS3iAnPKPAMlLIRT9ZCuCijF
7UBEkbzg8OUV4QE5Rih2LJrA16LRRbOsc1Dp0drkel7u75B8c3gLwWrs3SKYzN8zrSJbWzfzQpwl
S0oi9ZT2kdav3sKSTV2eGfitHrCWtZF1xtzCWVFuOgz2MxLtGSQjqR2FsHAtavsNTH28Blj9TdXS
Dv4Og5JDaQm9DqQJ3R9Qooxauq7E78pl+tBHI5JyMyurMS20SIc7S2nT4k56IJqAtsT5bOCNPN3O
IHx0MS7lT7qpPj8HpgIsGn/j0nKqW6wtt9e6MGiwkuUYIDGgcHhRZ8+NJr6RMtxTa+rvajB1Xp7u
ZwukjhqdXua9H5cMA2cLvxObyXpIYBEEWMOOuV6AnZusyYaQr0LK0DokmoSbuqcufkaN/9zcCXzr
hK5FIv/IzN9uZU4e0rguwOr/itm9jDA3aC3eXJXf4WGTQjbGhuz+n/MDrY8gPwwAjQwDkJlx0MMT
Z/87l37ycz7oVIk4/PE1hhhUoiJqeoFBBAySWTU3/67I+GPCvdh+5W31mmfMNkoVpVJXWopVIQih
uA4WqHZDMj9PkXKWxCzjD2KDKSwMrlWNETuJD3o4z5cTnT6C760BqLIrlW0O02nZmhVt8rcdC2oM
mAR8CHwI5cAx2YDKU6URZV2cW3UU/OK1BGn1Ekav13JB4hvBfkzNElPtK+/bnnX+k3ngEPKvLErm
d1u/LP0uv4ESUm7icwZZ/4DeCLcAX+AgJZLUT0bFDn1d/G1hJmJIrYnb6qlLw2Ojovy+TW+GFnRH
i1n4U6W/BY1KM2giZz+zTbJG16su2BP6jJdn/MDCWH9GagEJwQ5jSb+7NbWZ1wqQpe1oMSm+LML3
dvDp7ouK4jVMtX0wTs2JEGOJHq1VGQZHkm8/WYfcJTeGTvDGFPI4i8CrhpBmsghoOtg1+USrlr4c
ofIpghJyNxrwQIqH5mPlQHOmGXelCkdGF0Ldd6Ki9bNOgwLCNOlhw1hdWXhJbQ+lbvRSaiNYF6HE
TUmzRs9nKfgXMigpnSF9IHk3JY9s5masB/xxBp/SG4Diqehqvr1yFEA7Zau3tXTTvY66TpXYWUcU
09gFPKovvyQuxOgd588hWKPKZKDVZHhnoSTR9PvzPr0TDi+InSgwMrq+htgPYOCERUZNfQGkkz0C
eBo/8NjKSIP8bb6ubQFYzMEvPIb7sAfyaX3qIeUnZESk+IBHOBr0jScqxa1sl97AJ2P5GDWudSio
q0AEC1iZ31Lbrc4AbvRvip0vC2o/gNh9xxOQxBKMv+nSTyk0ml8pqA3Iz1j6w+nhLYQVRm6NqnCY
KkLsgaYjdoQHYFzC7PtwewVkmx2Om2REswreXrNtwYi+J+KdpiTdHybtiLp/uYSfbyufb0EzI8ug
zvoCHwbCRbZMarmkloJCo+tLSc6B9yM3d4XmjYB0ZpiGaNxbvCP/G+5QbzapUYg1xO3i9j/ubibs
iXUEMf7ymnq4RfX8ipOXGMAFO+gftro9wWU/s8kQf8icLQF3UBJfdTGby9DZXaSQHZnhWcej473o
Sw0UddIRwoNqeoiUfHzo5JtgE4yOMnckpo353HF/tLrjslD7Lw2WfwzYvqCtI773QpI1UF0GFoJB
utDfRTU4jq1S1VNPYSGG0DDjNjBRN67wiOQKnF6uhIhH4KhkT84aQn5oeV4rDRVY+ETj8w+qiGIJ
Gufn0v0N6/pmwsy606mt4Jffb8FOThjOaLxgyYp9s3e9ZIx2djKN2DF5lLPHZcfE9ilqlTT3nG5j
47JIHOcSNWzM/qtF8IF9XMHCdEPxQ6oDZyCbPtzbmCKpdoWqyibjuFfLxULJ773//rWbuVfwrhTY
poflT+2DOsOSCKg4EFcK+GVg/ndxkTz2yU4lTmL6QVz0X2WxR6UxtHeCd1cX2uOah6peUu0a3gYb
Mf6x6RKwTxdNFKP15/mTot3cMEvZT9Q+oWipD72OmQjaEadMSw1SGnzn3qNmVgRp7aFQC5TSJrcf
IsWoCIYII9HZZF+yvMCL71PVqFAnFPUSFX+pvlVHJoj7IZhmvW223YEARHQkHtUgRXd3uhXR0rlP
vOj5ZvMcCdRZxz0JZ1s7rlnxE8kFyQNcWeHrsY2jmLz4JcfDirSl1Ifxt/yLSOUWGNJBx0mPCLs4
93IhmWgY6/6HS6taa7Se8AZCC5DnKq0TyYk3S5hcgoo/PPAA9NXRMVUlRfdLEH0YWXDtMB/8dkeH
rMDWpVS0oCtWjymEdBj3ast8YMVCCF+NAxno1okaPPJnX/fIXEzWbC1jPBfciZUccqRWp3Au1l7R
C2Ca+u+mordUoC99tzyWbqRgo8eWSlkj0vKW3QhLxzvFYxjhQs5TVyNeHUcOv4bac4f5la4sEDl2
kOTRaXbTzduKqEe7k5Chncf4CM0OVQD+CSV7bi2sHEfr9li8mbACKp4OK3IX5ZBaTzLUJHe0nPmN
W4VvL2NJg9spceaDQQjT9zAQBK8idi3P2yO2LNGzAvDt4JAYIXGEFvzuHLBAUbwovi+0l/FcNfgc
oIxJNFs7M+SeWeviGnKqVLG4xvW8JEXIlSIr/1C55PboBCwkQZSEAEgpH5K6vcjFhut81ul5SNE9
9Evz9+QFHBSBNOM3h2MVr2J/Er/Ugopr+XCca2oEPnykZfTmZbb3RLgBd6ZRM4EuS+EZINTq5o0l
2sLSZuDY/xIVbAE6WcJe7cdYzt/qh21s8apBKl5BA8L/5zR9v70vUJ0iCA8nMr+8FmA3jJvmspX0
pCRfkDQeeN0QMfXAV5XfRUpi8sO/0bjVLUDgc2UKVjGqLnSgOFzpVLVEZRWTRLdvMOTulX75xU3G
XQgeMXAK9x+IUiclOuPflhH9Q0MdOs1jCy+oqrbKMFzPD49t9rF38TQWtr+TA8lab1iQVs3qJt77
v2mpV//HMFK4BE5Udb0aUjoqbDeiY/L7ncjSoN5CMljYBEG44ByM9JCbSxxjTddyKLnyHC/hD+60
zlY0zV2M7Bkh20gPMZAHBiFnD8mfar1w2FhOoDA92nSjYoBxYdV6eiLtxnWRdM7gSbAyac/ba5Kk
fVG//9RJwaYU5DdX5tFKMuN8O9P6+bbImj2x7DctjCjZJznPh8AL8LHc3x0C8rHbE8FhITyyusY5
zJug5O8+KYmhzpn/+HYORQAkHgABEa7TLm7VG/9yUsbUUIZJhezu7aI+i9IfL8sUclOBhZY2gQZY
SVJZz/bpHgZexKg6fpOUVOl7GTP9hkzdE6qZxdJOESLkNPZanvkjuWeJFfIt1P4jSRM+VE1qOuId
OLFkQ2Vyjxf7PX9zkAed6pPbHhXMbd+KE+3ZZaAn4CQXWV6CqLAJXir739nP3oUu6Uli0Ws2M7oI
rvh9ENgmAVyXpfQyFKrSQz1OrdhGE5LqxDhKHV9so29Sipr86HXWZ+ibyzb+B//uCSdSgn4LFxNx
3Erl2H7xDerABUC2p4+fq3JQvgIfsPq0+AmXe8oevmdqgTsA3srT/Fv2a2aExyqixYybGRlLclLb
5OF6lEU965Ivmr4y1SnA9adL0Kdga5M10vvD1zQ+2/+RynYholCOqlElZ/XHd8/moByqwMcRe2wM
Dznke1KAtdJxRb7m4dgqJNI9l7vcSu+eErnTxGMCge8noCW4ChgJ18LjF0wC7S6In91h6yHix7XA
SpQ0FoDKLtaA69vl/NoJ7tVfs45L8szQcswVRnyLT0v247iTZaDpwNcK6PahC9xgqU4cBlvA2R3A
NtPP3ZpRFQig3NgwPPtkILZpt92sEzHiwO+12s1UHqo4jaQquhUu2uNYzeBXjbN7+9jgED74rJ/d
Ad7A/WcrZh+8BH/Ke8KErIbVMdEFFcSW3nZiQvw4Qb/VWxoOoD81xCFkTTMejHtUnOlOIufwXVhw
8zt5WaHRRa/C7GZ2Z1ZyMdarKhiAAK/dmnrcBPN2kv0JEPYnM6Q9KvGDAvplzJBzVRdQUvdo8NKn
ce36R6pe04xC8JRdy5mt0sX4TdsnF5H7Lva3CaMCeZwSeDINEgOSm5WpvxT8cPFMTc9ixcVKgcD6
/X++tO0kErgXp+o5NqEXsDsNsopeoidzuD1x7KaPi08RDZAIuLjb6OLdU9OE8Ri1Pi4jW8QClmB1
SI1HGft+UQvqj+LUhvvX2kG3Y9GdR+JygE3GUz+heQavzzMr66U7y4LuWnozNZmsiGdXNS/rtAA9
sniA8xrsa562BUS37RR1MWxaNNb2nDV/vWlk09lZWzAvN33cxYJViEQd/Cn/pa7qxfQYqq/lBTcZ
kFHisNCfPz/mfWpYXvFPBFgvt/WGuTGNVSd1wtahbiiWMAtls1jITsSP5Ll/y9YZ42vrMgvq3tfw
LO6E85ePsTrwHLzpYvgQ+BqossJNw0Cy/fYVXKYOsixrBoj2x3wrRer2ZB8HVU6UeZgdRrRuuuDb
ojUU9zHrYWvATssvK2HsJ1LHC0GM7iA6bzOw6XYXGM2lTX4NY+goctUM8iZEz19LzO64QZmb8nXL
MuZuG9pFFN0a6apkEae3q0h0CEr3Fq6EOmFdh2W0wR+RloGfMFyYCZgXCBYKUMJ4r3UyWHCwAGN5
A3SOqf1joZO0ZCVrXcziG+Bl+9gGwKeJwGlvSyRWRWonsJZz6dcojJ8YNxBEEe7afKFqTPYjJSa6
L9gTXTbbwxE64D2EaCuqRK0RsnaoG7QPvLY0NQWW1q9qL0qmblwqRV4BWTPQDHALxD9CCHl+HY1Q
KBCzifGLKZzJWTP3lZBtWuZHA9mdX+BqY5lJ5sMddkl4oUW+DbUs6YokAtNr+IWdylxApTMF8SOC
yw691ENGD4fjD+FMvP5/8RwRVx6lzmUViXWhjVluVsFTqQVa76h/4pls63imJTjwjw2BSfCIhqQ4
jspH/GxA1G9PHVw3LdbjTdORgl9kGFpS0zKuLd97ZEKFxcsqy2+TLYrdkwmFmMv8jLWoy2jwEKm6
nHZHC2VpxdTUdq6NWNzaEkKN5XoVZQ9xSh5VpX13QjFOhttiWPqLDTOKlAGvYfa1aozHNLZsSdye
Zjlcnw4OqIvRhgX6MDdOscxhubtuWNts41TavWpySgimacwKMY0Dq8NOPeb3FNhos1J+4CQ83D1n
YStoDR6SyluSb0gk6PR8s5t2VLZ8OJRv8dgNi1wTb7XxOHUNy8GPrtSr06gP6Wba7J696ri9uk4r
8ejiBWozqt4HQ+bSpCvbDLI8RCzEGH2e0S596YUHJj8ub+SSs6hAmYuj/+IQgzJxDWbIvItmZEM+
/B98TKCH8gtqYWIOkZ2N+btpUomErpvHo85HzV/5fVpWZ6KZewi1OQNF7RIZ606MMIhgN+gztMS+
PqtYaDNQowkGUBTz0BXF63WS2JXZzMrrLDrAkzpaAW21M2yes7/tQFymYJBtbpWVOFxXiArt7ScC
2YHlSmwDP2XwLHnyTeEyBYhWyDYq6JOtN+91Urj5aR7Qv4++83PFoiEFgA8PKu6RPTXXDH8QiJKF
c2F2H8n/stGaSOQT2Fd0Rs/fBAMlEIyWw+R9wORgGh2P3FZV1z7Zmr9tZ3gY0YhxFYIRJURbQowQ
VhU7XHR4B7nvYj8TLf2pJAjyCnk6FI/9lOQ0/1hynL+KI3xWNGxIFHvS8oSIo/WlfgqG5JWlaLoC
7SEDueVhXhLcQ1TBuUOg91yUCZP0SUEr92vmDpLxmXIk80JIZ4KphICa7zI00jM9jAFJVqcCMJDT
LjS47VghMalVMF98Dbhk0OyT4tEEqRoStQPUacU9NqIBKtv466WTxcNxYFTcpN10qg0CGuohLnqY
lN936wJHv+CqBeSHnGYb26CkML/YNpWi2CooZIpVN/HyWBtt7YJejsnozkVT8nyp6GoK1LCwwEPN
7vV8S1Fp2b1h9VYH2pe/zW6gV8wJHz8xKnStb6QopFsJ0SZSz4c16zfVhtt6mQse9dwQ76H8wGA5
YPco9eN2uIVCdEblTBvX4aLxg+tuecv1P3+x/aKQrjYhIIkOHsA5+gZJnDScFqDLCt1Ojs4v5xBa
eAGeq65LhgTjZxOaj+P6x9y8/mPR3NFQVhvdyDVcAqvheXxNWzEDF2iN0x+zcNkpSED+e6s7jWcu
U6U0DmOBtmH7Yea2Bo6J16/Mw8eTNEdkBSeZyapvY3ru0LZsXSRZ0eSOUCT/yryyjn7jbuZ+BRef
ReChTOZchGxy1mnYnMhwXdpNhfQvJuQ6AWlaJvQMzcUca6wHBnTseR/60Ut/Wal2XnqabbwO+Qjj
XbC1/uUBj+kezncJ/jB90T3qYO2Xa6hEPDTfnAV6FbN1k3evYZPYInj1Yxuqw6wbs+61rg7jz3Yk
vMXxwd8Igo8WwSh0GXgID1HhOxCEEpkxEuVI0Gjc36TvICy6tPa6ldTV3gxYySGlgr5FIWi8zSJn
xSBtqArbjTCL2EpsO8I4ETN7cGWb+qQEshj9II/dXP5C3RH0V3jX5djZwQrFrc0l86y1y60ScXdt
zSNyKo98/hbKrKRYJxdBCAnxcIuvsQpKSJTB9p1aE3VuJ/hKRHDtFPDbs5FiJgNM5Mwd+dEkqiBr
YlNTH+P+De0U9pTVbfa67C7H6dgI1JPNhoaw/wGUQphnAl4eXlYVUwozw8EBkuNj8ILwe/JKNY/p
JhvcVAxwRHO0WwzGeESV0e9tr5gWYWuN0yW725TrEOjfd8Yx0enhbzCEd8Yf3su1MOWsH5SMRiGA
AWSk9p8xBjiQQX9VkkbQ4b4JQ7S40lBeD0+trgwNMr3ME0mF90riaQZyuzKO8d+gIsD37Qt4cJNC
nrqlpbb9Q7l7M/or6OVWhgbS3ddjwNbxdo440zQwLOpdy4bX3R/mFvqYDRU7urfMcHTeB+TJ2lUY
vqN0OXfkZ0kbYOuGO61PyJyjlVHfiTp1WvDMgqhTA7fQ9a/eXbOBV63zYerHMm8uLriYnBgQgqEq
TfwVsKnum0/zyvwlp6v2aspfHFpyh3Nh4McCLeMaf6HxYd166GRO2f6AP3X8y9l0/oAyArtBvP/o
8R5Xuv0fd6g+vRpHo+cXj2G1c0jBIzWxXiLkDohXAXGxZ5+wKSZtvji+dnEuz/pfHA1Vu6sO4bFR
ePmvnd0yrYwuVS/GlbE6ZBe0/EJGEwn8o//Pi2gue+mHwbCA0LXJoWySG+ZTzZvVO8xsvyyNv9ov
HJs0IxX1GTSuD1pON1QXL/SVEcRQglLR9t0x2CYa0GLiNDosk3EyrV9UX8CIzb+/Oa6gG6DA2SMb
lHAx9Ubv3bzciKGY72/CavAfletrHUBo27FvsBNrkIQIRoNLaDJhR1RxY1fVrcT312wJxofBEyFk
Ef+sCV2SwIalnlBkwFtJ1Nps9YLrrEf+tkSYtjd6331+7oWOl5tVBFzlHN3EaXPumrCXFAr8PWNV
RFdSi2xVHf/KZfK9cuZdbOHlJZZCKujHU9//DfnuEm89XBT4fbij1siDYF1dlnmaWmJqdKZisIbc
NXANJ9E9CJ67sF7BdffdKUd5DfzLKC6I6s4m9xyrxGQ0V3XZrR/K5CNh2pmfE0cvxCfARkqShD9L
JrFvgpfY9vXXRPrdRyIWwPL8DCaVhIM1H9hDd/dLyseOOwh9DyviKLrF0Rjz+pXbEmmB3ej7P8ZN
EixW/DKCDc9SMA8LW37j+dGlY1gTh6I6M3nvPysGpNSdks7xKBsstCnQ94ryAig/KaGNN0SHE9ZX
bnQsip9Dxs1GhwEt0N/Uc5jIu1t3u/XyNcpe1t64VlR/P9xACx5rs6rl0dVLjDee9RODQYR3DkhT
UKKQuJWBA5TMiv3BhWhD1PQwyeoAPEn6fwdNPWfabzsxbCoWUg3Lb/zc/UwJhO+vWYzvhUGBb42c
b17hC6Wqn6FzWypnN0HZR2sKgLAWEILxkTajDrpn5hDFlCtsou3pc9kb8Jb2mHWTWVfM6Myjg6BR
aqFbW5M4rY59VH+Ag9qkjYDr+sjY0oH0PYwVSCy3QRAVlU6K4pMamxi+YM7gGaCDZ497r7UQW+AG
Z6qRcH3rUq4a9wRZDts/gl+MMAb+bFxAYGmb2x7IwixYd6kWPITPUVCeb/mlgtc1XvzYYxB74+8j
FPQsOgoLuOfRg1m6W06gBOCpANdByKvdyzn02BNviGptQn0WDKpukL6w7P3e92HuRP8pW4Y9nHQA
ZTWLSRsLr9V2CesfPLLyv6nt00o5dnAQxxtNCyLB7A/ZEiHyfk0TPdBbaxhlVaSRY+GuVkMQuuJJ
R6WatfoYWKEyPPG8f+OJclPopDLT6n6XGDDUqttkNMvfQ7yGaFDUFsinnrdNcLHXPiEcc4Ul8FLa
J5/6rD74kifaJW7V47kflRldgZ2jVPyD8Nwc2kP/o7hWTUyJvxyxzrIU3HtDbCn4x6h+gav5DYP7
5gXeKCi5v/lj5i0yByrK+l2+mImgFxTGFpAt4nCZYMi4RhuV7O3FSONSbB8Q4Z/EdpK/G1i+4Fox
U6r10PqncWDqh68qm0XMXkauS/B7QllQe0VbxlOm2rJ3qlh4PVZZezlx+NGjjqtS2BZCkNKbz59f
3shOGndioXXKa9ZVxrbyh0oCpK3+GgTPe6fvlMwpUUBCJJdWw4v/TKIfD5RZOZT/m29XUb0WcD5l
b2SGghEUXtWGwk04C8vriS8mgAi+nYeTenjmoE66cNYATLqupwawvfYtA4jtup0r6qY70S9u3Pzf
JLTHIPhTcw7WAy+4Ohojlut/UHQFtZQkXoI9svvWmgRDk7rfMkGfi6UT/C23vbV2FKox2SFRgs/R
H/pJCcxyv99AGhq8iSFtVNV7zxi9rUWyqL8hoWmAeLFE6RPo/RBtG+7G186/BpvS/HGqa2z0Go1l
g1VjfKEIwrrGiGqLpMO0kwLxpIWcbcstzWp3KcChmyTXe0xuQ/4tsLzn8pXHXs7WWZMscejB7N/u
43Avq8AGvYHn/A5VtgB28lPs2CvnQniii22AlD1YnWPZP+LggfC1WsXYVuf7H/RmReFwfEaKS/Iv
dHKxC5ZlLdJQ6BhF21O8CiTU3w5WBO64Rc18hPgSGcUPUIfqtutQp1NMk5VaDjBogd362Mmf+8eK
d4d5/KAMgtidJw4NwnFEmmIOIcDR6vh+1l4u0guOYOuREcfBmAG2m1vbpLUy2+DMfNQWM1GUMAD7
/k0r2XgM9UihYQxnKPhvpRABENRXlL8W3z+4GxWfD7gfOAqu64JYG1vnk26RIv/bAKPWv9nOzuFm
wvCqD4/WzKdLY1mPHzoqy0iiIKDcAqR+g8uJu4DxkzRhQiaTnbh+uanrh5EVZaSQ+SXbQAeDMjJr
bIvSA0WORK/+zB8U5viLUSuVITWI54ZAX6MfYZCSvkn9OrI3bLP/TY7EAFXULaphqr3sIFCLkTHH
bIf6R5W76MtVn8RVageiNpFqcNW5WpT8PtcGgj34rAP2BEOyVKci3sEimTHGh+ujgObdgcGaKACe
qBEqSs3FYjtuutJ/BsfunIzlEEmCnKy6jXGoFEFUviFJG8ByF5HwNHsXNCP5tV+PZt/MMUIUiiCr
V3PjHmSasy2FoOG2CvY2+/9/BOvXi/yd5XeyDb2V2AnwFGhgRoRQm3xyDWKS0TE0Jie7r1HHrlwa
Dxyj30BSz4cdsiF9pKV/Pvqo9ZD7BiXGm3qwFBh6W4+8qgl1lYysw75pTl7emV7FCyz8WdsJgiOa
1SYEBbEQNfTXr3dHx56KTxC0sqT0ziV1FKHsaj38ghrw8sfyTs8WMt5qIvA06wqWzynCRKl395jr
UOdIAIBV1sh0awILQIVgUgYi55PQODgPmDit2gEhG6FpplvZ9WHNtxFiNFS2dqkb6z3jZGAl58PD
36pdxJD2A6YMckIxjzZQZfajUd7X1vYfmDorO4R2Bd8VfKmBAwnDr7GKXLoo70Um8dkT9+gWWurf
jOZxaQnL6usLLtJBPXxZaHPvLoSCOeGgMzVl9fqEYOxD1fz3zgcNUAxCT2W4dFVeXKdh9VlQq8Ah
MbtVz9uMlSDXQcWGcnvm1s3doz7F8ltFn5NQlxtKKtv1qwMgxZA9CGLTO3cttzBYYqYcGut7RRu8
nAeAUlo0bXZA8i+Oy7Q4+4pziMqrzsMu7P2tSaLrZk05LlTy1PJ91+CUPU7w/MRxU2kvG3fHZgZC
bMLnUOd4Dp6PDmlaJbftwXsGUfCFuOJCk+dLXoEEuY0y6+yVjnDrRps6SZSma+mXBzTbgSvKxfR/
q6YSkmNKUQr9JXM3AFEWYvDd6t3aD2sAjzvt7qae8Js1lCi3f7OwjkNsMNslq25Wl/xzl6+JZlRP
iS+hBEhhRBuTaaBPiPy6+X8lRxE+xR/RMRT7kbG5HKrCqj0CEZJZOLpO1IsjW4CX90ALrBp97gLq
gHCm6p5OBzXyHg3aK7B+3H2hdbXO3rY/r9BUYNuel0vn5FF9R+vLAGO/uIfsOZrNzTUgltDbR4n4
+p7xe8dqNqvRCbja5v4xeIlBwpLztng5eVhmKuFeqwjo5+K6hrhIYe8EJsMgLn4XCCIXgqJsql+D
yNF9uBFy4v2n5p9h+Du3OT2LrAHAailvQu5qftFOxsaubWlX9IyqAMbaxy9+Fl7arJnkNi/eVlTb
hez393+TUM95F18mxIet0+cUn6CrFNBrabimo48wZ60p/LEGe04rNcyKF/RSkuwe4WV6AL4c/8uk
FDZrZhkz4jN8KZ2iyF+Fhoc1jpq6KnhinmsWLCSBcifpng78o6G65YH/vnGVKSWQr2o1CZ523csk
amDEycyqvjyWmqv0lrO+uxjQjz0Y9gpph4aIFQO1g2zOr5IK3VQjpEgW6CIR3Fut84i7iObfwjDd
D8Mgp6Vhf+rf8zl7mFQqP8pfy+4UUs4gaUAbzWGLZ+Zh1osvjA/85cUocsKsPgrYK62bqfi7/W4w
FKAQnUi9qkBpJdSjnQpznL3xyXQTZUFgju4boQ0G9i+RWDwdMzh0gbBkyPNRKnwysQztPMuhMxlr
BNUcGoSUiw64OgOODmaoRmHiH/agRr10B1C/vHnkbxqP4MgLOEg++mPap+/SQZeEwrrwbRrrwsNI
kFaOTehs+/rZ+tOv6ZoKUqhbA+vIw5fFj7Ps1E/n1sw20W+2kFjeMoWtX3h420v+ZE2p1dNUT3Dw
JrSyygdS7j5j0MCD5kvnFAOhThB6tMXAYBbThwfAMQ2YpvonAcNPpKbToeDKoCFjThtspe2474+4
pZA547DzSH0yom3ioeyLtpqxcgwAB0RcVJad40PCCdHyAUP6Tdpj87UgBOz8bjpJxT8hLEvFQQd2
hiCwxWQ43Xv1FS9uYgp80vTjvqC/bXNiSIoHzkP6DjmH1xDtX01JHFntIpLbXmxgdK3Fs72Fg8X2
lMCzRSienxYbRJxjNDoWuZvP1mYNwQF4S2zq76Hl7TNbqlfTGQ5A4BnXsGf7xEhAkUt9/TajJ+gR
P7JP7VpYxIdZcwOZq1I3tSOvR7Giuhdj6Ups2z2CHgyPzhVW4OcJigIvgNXTXW5x/40T+Meka9+N
RPGrAaE5Pl/5QH+r2n+khM/CD+ucxbTtOKeWD3l2wrCWGV4KGQZojG6CKDFUPywe2Cv6Oq/Y7KcH
K3s8YtgP8Qwuu00TDEQjUBgQA/m7tX6t6m3vdulW6xvOF3S5xZgMx0JbcIQMkA84CaRxFe0+e9vZ
CCrT4BJcVwLmQfLmb1+LTKAbliSdXKaOPC0k0r+UvSN5gyELxYPaLzS49VNiCDwACvTp7nIn0Bw8
Fi99Lnb0O19E2Zx917UuSZ0biAX7nCOXZd9OZf0/5on9CYLaau2Ho6AB6onMbvV9UOqP07vqkQFu
xi1a4fflB+cfBoqZIKurBR9o1x7RG0mdvrAJ2uxDwrBAyB4Dtg8NUpheIPNMJVijt83fqIyEyVOa
PUyWznGf+c6+saR1p0Ii9Up3JyIEPMECGOmdKsC5qFwCEIQoliAjgSi6WaFs/xMnmE7yMBiUI2zK
PKHewFeE7X5mc1m0mRv60FGCmh1cfuFQjUOoKYV4e6ma8HTVYtSIetPf1p84Vm/B4PbvnwqS7xIo
/99EY0qNc3NZR+A2c+7QavHRQkAypxNeXzGs8kNhET3zRYAzg0Pt+tK6dVokDEUngybZ8pPKVcxX
YNrNbwGWQhXnmqx0gi/uqajtzFbhQS6HpWpjnSNYmT3znjDaSYczSzEGryMZgxOkpU49gmgMz+4K
ga8WCOJFRZz0ZKIavlSHydAJi6yVQIzJU0Bma0VhgbrjfdkiOl3v+G7vG7gDRpVkySkwavvcLX2T
MWbiut3/ZoUTLCb8YOIzzNHt/zmiA5qbvJEmAvaSjNMUAZkrCcwdGD+mggLuBcYynKZmUAMDmJ28
oYctWZnheLqtHXfwhV+jeDxv+aDf3E1G/0tUl5oHTWrKanm1qMCf2bGWH5h2QXx1abkU6KUY2mau
9DO8Xv//u8nCeogAgC5BDVhLrTh/Ry6GEINUhX7sqEa7+nlSwsHrj47oTNSuPnDcIGIZoB2V2/sr
nZd2RzY1TBDLhn6Da4wuVcpfqigA7NkUxR3WJj4qy+GwxYRs3IbTbw0sok7BW29XzaP12HnKzeKB
92AIliyzvOwsI4puz0rK3FB7RN1AR2bLeI3tkRSjfJYji1cSPk8LXLZ8ezFgfpS8CktNWcgEJ/jN
NlHkvBIdCJyz+SiglB8QvZA6VCHWD/V5oa6Pw0MhrUK58XMInsluke+quDd+v07K8640PICTGa7T
1rqjn9uunK7JooeeSGMit1cz/39cg7mbbY4Jo1LTWsxUoiHxFnXROo8iIPWvq338TK7pZiQ4r63h
aDCyrtL5Y2TfZV6lMdtsgY5ZS49F251ThdaMS28lZtUDpZPmZkHZsjk+5lsrtS7Wul/aBlMmAbaa
OfQ+Vwf14cYbKoAdnbTRvmYdSis7pLLUCFAZWnjDYdw9KMOJO0b0syzaBjXVPp7zDzfSG20/8N2c
7Abx4FmHrfQ5ez9HKLTa8fUt8Kzs4L7PfknXZKR8vFE9UK1xsSWVybjujZXUne8w2IyGOXnJjKsK
1GrNoVXfI+j0p8/5//gDCINbwAp62rnqIFAW6IAK1vj7fkpNJjyzJ93YsHEhewcdaAAIq/4exQw4
oj1Yb7A/sJC8dTUtnD1sDIJbYkN0I/KM8+jcmNmCA133fSY7gobf5PMDhqceVqnWbRxmm24dT6EB
ix4FhwSmp6XHvi3qVzzagWaocGFw26y+CyHII2zcY2ZaYCKEkhrx8MHUVCWDK4GDCqCjtKN+j4J7
rSDSPsUazU9pvQnDvKReOv7eNFXIXEQeaHfTHZ16Gvh2/e81gkmjLU4Bjnp3KwmD9FZ8vl78j9pS
k6XcvJ9Ys3v1UED9amO44VIqgL7GE5EgGV/p8iSb7Gs5BCBPaRBMh2raBl4kh7yOPVW5OBtJkZI0
t+zHGbwi2X/i5Ri34kYXqAZSa3/s3+gG10N31+1ugkCmyz3ssORbV6iJKEb7Yx03MmvVaJvrsRm7
OWpAIpT2Z45UiwhhzDGJ4m2P4ltWciGBVDwy4KS0ZNj5zbH8kkZ6DwT9CVrYuDkgA99qPQMdWjd+
FWG/m0hBkZ18xJKhd709ivUZJVFKvlSVL2gWctQdiL+/L6NzgIiS4Po+Qeu9+zVhQo53FXuBGVe3
x4JcO511nn/s18h4F68zfd8x9T/qFwlHgAXvozb/n8kD1LOzYGockwcWUpMK59RGwVV8kQ8NFPJN
HgRdECx80XsYunh+51fgtZACRbp6l5CWLhCT1lzbFBavPvRXKb/aLNFtUmrNc9oT3jRaGI+89LST
MbFrXMkEZh7vaORUaMCvKkVr3Z0uaLNPXV/nnT8vMJ1lcydVZQcCD74VetXrwLJmn5dfHJ+A8w+1
HXqw2VSZJvc/YAFspFa+i3EnfxZwbsQjgyIAzl6Jaoc45yp9xktrklL4Ld8CiQxWmTIWc3YHHGMq
QmtA+K3LZ0R3onC3YHo/r94OInWHZC2RvLtGhppCD5zsTdwraXUofzY9GBSqcjU1Ag27udiN7uNe
Ex7abeUMbYZQIMMGbYwSNtemkf363aCmeHRtlX6hvV979eTFh+oi5IoC69pr90kRvWtQQRjWew5L
eVig0v1VxwsD+wObvFdKLwjSAvXl/p98J5kW8lD6WKMNceB/8I/UdIYHhoDBcm/U7T1QhYjKMMAb
pteZ1TsJt3VNLpMtnbfOeiqd54BC5/APvBCHhIl5IwRcVq0l9I5RwnbDfvkHFxkQrx4L6u40HrD0
jQH5gAiZBbbxOnSgUOYNI9K5ay3eVSDI9mZs3oJiax81YyWuK3TypQuT/u/1sxjaKkMFD9/zOuYO
kLlBz3K2DsCrO/1vxr1htSLKNGQP24ZAoeY0PI+y/HlO5AE8Bze3Nb1x9mlKe+UZKzqeDHWoSMLu
qu8T9sfia8E0/jG73M9kD3mjztZFMHJGNVJRNynqPi4/vM/BgZN182R02J5t4uAxzyNoOWDExIuv
hnxm0dAxlJYR44YX/BkHNZbuSXmAgeAap89/J9BmE6hgdiJBQfUVTDHY86T2H/vhgN4h5J/16CkL
b78gqEnfHbe2hw5UEHX4ppIGdUPja14aKixbdneaqDygS7254hIBerqE+hLvQxROMZxY/5jB2s/D
tC/jVaCZHjQqaPKifkUY5Wlm7bZsdZcVQez+ZVxW5hj1UTrmUYkpaHJOP5Y6Jt5dKMBWOfIB9rNT
EMkNiV/CyazNjXQgbPkaQEdS3x7eSN+sOtEW5ukJmPk1yJ+ZszHeA7Jv6w9O/L/MzY7keyHvoOf7
W+0TGNAhSutQ66KNgtobqV+UZhGHC+2TS8+18AL4SXWu1IBSmfD4lxsKclmKgbo01Gx+01YNLjA8
iw5/VDGT3CAhGItUBs9QzQSv+dU4u7XZVai5KNcl/hphecsgpJ80Xjqp/sUVhYHgPLI4tkDYwaXZ
OZXPAui5MZKHPgk/WqqHKNGMplqsTSn9b6R+6VunyRUu4ZbcdG2S1XWuTUcYyaaIzfqru0osJ2ci
JUYXnthrZBmPA7cnbtBJsjHmaimLBluY7vo2vBM/uBnaIvkBlNKw+P4AsRtnFHnLIqkx7PDEoHKr
3A7cn4t0etSNsO6NHmsKJdikI0b/7IbA7BmiVEFFMbojGs1wQBI2Mlu8p2w/JXGKsiUDdnd7YY1M
4RGuLvT4c/C4biCTxC55A63u98UM6IQDgDhvRwJ4ekT5Yv+iOdLjpEqjzNAR/Ok9VLhIUnLILjFr
iAPqUrGOb5SlAHkqmAEULUJTL249mhoibmcpYxTNPmZZ29onfiNAwqJkUfiucIh98B5/RYq+HNFS
s2VMyy6MXpw0AhggZEJeV4674Duu3JqVADEWoN3UoNmROTx/X5wu+SmJIvMoWbw/OmDd6qUuwCSU
R7+oDPMVJBwTy1lsEsOkTE5d1ekPUQZq7uTx/iC8+1KpY6oLwsNRYXlEX0d5wUkoP4Fp1ic+EuFy
PgLIrg5KUlVc0Pr6hj3RBA50FqLGEReOnd1THUSmJOA0vDtPqcOvHuBsdFWBjLyy8WbyVbafzCsZ
mMvVazxqdrszslrZTr+8TlbMI67o6lKAgLAhL+HWg1n/bGwnWzLBVfyHKVQtauDOHBtp/XtRiY5T
8/ho/PG30sFsjw3hnfRyCfN5IiIfohsj6R0tYJo3U3+b1gNlVxLNAtms/aWngTr/u3CNOSozSjVm
I4CYrBVWgqOA0OasqT3tVYclyJu/Z9i2k1Ju9fuF4c8Zs70ocHfuYUK9DFmY6xjtDWmqVZpm8rk+
GXa96IOg2u3zJlRNYJM55Keq95ahg46HP6llCKJID0vl2LcArwW1h2McY7kLrmxKahLRplfUQ4bQ
eHRpl17TYvDUgjXJxhFF2qJpXbTIu2anHuBrwENvSr9X2LdyiSBIS6e5PBvfbjPSPm076WelRT9N
To+tCQWf5MzHcPi5wp7+7K2UM3thI5JwkKnftFXCdSrB8WnZp+HcdeD5ME5RRIvvKoOSAaLyJqLH
vLvzWpFq6r+VDrzVGDpoobKPDkRmO5bNcM3jQEjAmdexz9uFuCrVR3G6KupHJ530S5B6zSw7vzEN
26owpZjvkEJ5p7MU3iNq/9ZnRdCfl8vqblJMH3uEVWuJOms2GEpReb5rF/erDTJ9MfLQGTAC6TC4
aWKDSTb5TrKJGGiC0xnBqAda9AlS7oMouySMqFDhEftXjSWSwWzvo5s/2WkMCOWIAEFikZMepTF3
4A4IejeaP33qcJ/abZTweHZgvvgHZNzHzt0ddCTbanKvpDF6u/J6CHEeJpFn0mYvK//gOZrkd1E4
sRFBE4zjm56+ZyMeGjjY7rU0SJLX2pCVI/rgPPTxGwbVu6Y+bQjUp8sO01QWLz9BOEw5qh3nOG3C
NOc/SAsY4kt+JZZz/CZmyiBdoej9UUTmt2+qn+DTmoBsO+ZY81C+QvAFfE32M3II7IAURSMsHsoo
PZzFGcep2FMyaoTx11dDREZ7NV2gzCnmLAtJpgKfLFERQW4PhmplK12m3bRnVcIaUzBO14lxnnkE
eiQN4HsO+hO5q/eOCNAg0cj7xKfFWYcrptZXjYFFopiY11KmoBdEnG98xibky3zlxQTibv/hAJNM
g3M8Xzf7XFlpml2g++0V3VCp6qsh2IzVtrLFRrseAczi7aIsKnfQg4YtFB179o8Y3Z+I4sXG+xSx
EJWprs1UcDQ8V1UEuQgA/nDhQ5cG+pTWEzd2woO9/XtAPpOWniK7CbHzCJ0aZfulVv3gnBPpcRDR
j4+FeVhQS0AkAqU/TTfUrXRRxuaziiqqCLINSetqyV6hBFluhyFPPhgOUO8tbcDNa6Jdvy/S2tg0
SWkiCRO/k4O3Bm7/2MvjuMfMEA5hgzIOR5/vISSmYy8SySeLcuSQN/7FDn9u6/172BBx04YD0Rwc
zpS0RXyFyx5f9oeOryJ4qV1N/8nPLcbV3elTtd9q4TlY/zKOwdTpZkUZ6pyeNd9+tz27zu3HO9W/
sO8uFUoCcHEPLR4a3BtV6g9FJ9Sc4Qx5U93VjEpr4/NAzWmgvkXiuIgP5oSOjr/4XyK36M4uaCSP
DvwTaumL+L9qVLTs1AQvxS6uT42O4XNT4fdgGxXCm00mZ7GAIu8a5XyYkuTt7MQHEeDcPdbFM6B9
h12H7ljrP8D92s2zS8oOhrY600JAcm0/kV/5NndV8rQzQYBWl/0XlqORpv4FmhTPpgplLM79xWCT
50hf4dHD49m65OemZ4QaoXN5X7PPd4GqB9CjHdbXFo8p8mq+hVk+KWIEefTE5nIphkxVk0jXHcid
4JRctrn6IzkyYhAWnj7D/9lhevyziu5Yn8zSY9JOhBjSNbKZ99MKFCSoO5ZLNkYKZJgKN8XC63Hu
tiFHazXpxfPxaTaKpHpjSPPrhQwEm7LShQim8FOyQTtlGsoTxIszbxiTX0jt1eJGKC6g5FqGq7qz
8L1WqaHyZ5ta82EMNu0BPdOFGqQPgJAyymMMoafBsXNsFaigi3tdj5YrYu/DT/QkAvgp3YzR+jv+
G4W9J8LpK6EPonOibGD0wCba4bckp3BKU7cd8pnrU13y9SrdlEXTH/YwVgwtItLMJUBcQKjbdGlO
WHqNoYrJ760qVhh3ucWmSy5/krr2m4KWUAd/7aTSxGc1uWfuGwWOp//9FTmXoenGkpFK/F4ucRjF
hWLNq6185dpu+4LtwuSklFluI66VVBoZkxyX3caND7zpau3LScE654c9cL3pqOU85LHXbZEtb6Rg
YqM/Lm0MXH/moFRNGp972hxislTxj8mDt4NPPXEdl6FrtNNrNnRRDXWxEc/OB7AZfk/97iqWut+5
tdb1Lo64eEIeGzb5v1IcMiciG9lFPxLwwcrpGAX4USUnGCq4ORKx0E7liuYB8NzMoZINhHxdw8KJ
2A5tqL/AbYJJOUfyc4Xl0Vr4AUkYCs5nO6E1mPqKfygrpxcV0B1Wtencj1iXtAxAkkDVZSGxDPxm
33PNc3RGSILbkLtvj0fC6xWxO7marKFNMrMuS0qd3jbip8MFLUQo/vZ9eYZJsHKAl/j80le1WjRE
qQX65PWLwpH0yb4V53d5x37xFsEeKvCg1fZMErfH12+MJJck/SISbZ5YiE2hMdDk579TPY10vBs1
Eq5swSqx5Qy449phzrOVH0eJj/CuLCNzLFhr6yUFMGLdeNqLHjcUyI8TGvtO/B0euuhy5WD9JHEn
bxJ/g6BHkOo0lYGZVbgLA4m9uaefaOJDzAW/s5FrhfWnSb+U9OXstPQQv8j4dgCUhxWIDXdkeOpt
B+FU4D5FL+J+p4osErYIX1FZCYDlPawQq4l10kRqk8a/Ux2Ky6Bey9fhD7Mep3cQQaX6+xO94Roh
Qr3etF6vFt99pKUbOPW7VQwA9Ie3TCp8VQPEGUbCm3UWYy8Js0XwE/loPjDXYwJNVNQT28qmei5U
FsqZ4WFWdJBUH0X5GOmshknPh+SQjUCHUNeehygsLecIW75c0mzbKXoZzW9oEKPQSseGakyNfO2W
0shSytuPr75xns9HiWKyMerM2B+1WyPiUmRSZKO2DOJnd2k0MEwZB7lQrdQ6xnbcAPvpBu5AoKzP
SXs8BNJ5KVPv5Kt00gv8thjz8cQD95bmW22KCqshIwsOOtYODghjEe5JBhdjMjPPOZwZwhtmFNXB
8ezI69Pf7nB7svOw3WElHjpaRR5Zp2GeDZottwhTvmiUUo8EmuUUALkg6wDAAKEn7qDnreEr1ki0
gJNNcGJcLoMMpQGSUMXuMAUZoxcm6m6d6rwWQL7GDTLVD/wNzpOLJCwi2fQkHj15gGDjeAp8rpdU
m3ibAX8mlkLS0iu3py0vSpsw3r7wVwOx/mlimiCzTM5zAMEaObYFXvZyJM0pnlMvfb+1aoDsVaZK
L0EnnBp/eAxtxIIFAg6C0dj1Ffq7QcBc2jdKXxbok8h0jdgy4SzVi6tkr0QA1YtL9M3sDJqxkcTm
/1AMFfk9QaMrQL76IUQrWZK2mVqgeZG/JjED3PWHtktl3A8JqH8ct2dy8nvoPejkaPKPhQ8nBUDJ
IcI1xQfT+kyb7+gbC+iFdy+bH9DFELraUAL3zjD8Q5pLdGqL+4fGXUBzghwL+Vabym1w9V6w38XO
yIYdVD93rvv2QpWM9KaLrdm/akvwOsCkkRl23tu24bO5yoRiareoiv9sT6hPZ5UBV/qHyQTMX8iJ
Mxyh28JLWJox6tlIATpSZEjUPFWMOg1U1QNWnsQEwD9CGB0D6kExtqWAq7AKYoVJrD7/5NIa7AZ1
eO5U3DMLsOJuIHI3nya69SNXEgo8gJjcArAa+krJfEtGvwRaCZQJKbJN0Vw/BD2utpKNTQvfKYUI
PXhFYtCTu+8UEjdx7I9cADqHA6izBRxj4A+2jHYX5Veoq8vDFoof1WtNb7rhpXUGMs8qetx2b6G3
GrJHd49vIHOHEZi7DVJ9Xq0ZHx+Y93gqQpfhN0ESuG3WTUqeEPqAAoCNi18U2OCSQYRaHLIYl+la
WTiRVx+DzJ5WOEjggDgiL5kpPiGbcyDuX96avUejgn1QA7pTOQaMsINvdqkxPNaBVSGPXshsEQMA
+oN72ecEuS6oV3QnY5hvqzcMRAdDwZld6L2JJyw8rGM9eHufEkBk3b2PfBFcjtmNUIUW6MZJS6ou
y9aeBbjjtHkRHgpUqYHokof9WbUp34LaPYpH1qcjk2NKFpkLLfOcnitFfAelvPoCD5mDzHOy0Z+h
wm+hW3MGHMXxnA+lip7x9hL7tTwVaLIaPSxDMkBg7MCMlsBd4j5mV2XDbkRniO456yNqgEjF2M0h
BPQ83Aht2JYoSDH0i66v8+FXeiVax39dOd8ZC0XXeJuvv8sMwrgWflhC7IMDEioMI7m88nb7IyQv
lJnGOLCZO4D8kV7kyXag4KUciwWef0CzwiMvjVNyxspeze985Nb5G5upnAMNogqxq1/x7B33Z/Zu
Lcu+MoNQL4PbYp88XNYkhfLht2upBx+7m4NkCiz6G9jIRCC1zQEoUVl3L7P6HtB6FuBr/DaYEM3l
xV0BBd+7HhG+BLdfuglXm4WYsn+jVS7G2aQdWQ30EL+iS1PDLB2nxfxcBYSgVgoq3/0t4/XEpFLi
BEKLWbdeTf4GEuAwhU7K8JFPzSbXcnlNQMtNSpDMbMJjDfGl/fHzZL7S1BSJe4vWJizKLxA1M3T1
WN69RpmAQLTaVk4IAml8am17/w7mW5vjFQIcAFNoynvg9igJB9kk+vz20OTk9vxvcNim6mZSLh/m
z5pbpBL4Q6BDQThe+HdDNLn6ls3kMb6gMVm4mTgKZjUGhmkq/JnyWvd0eRmK7+tnt3A9YVNDpHsa
qqM4XVSyDhKnudmyXvSAl+7ePwuPv6Be2LWkta9v4m/ODoIWxhdKPa/Gjry7Qs64w8NGOThw6Yma
QAYAJW8DCVhl2di+dJFhkEzabNlgBSIyO3xNMaaOxEMjjLDNK56BDCFRReGQH4EqdTLlrjoqBF4x
10iwNiwNVmdyr8Pst7gawGkOeeXVIwzUtk4UB5H5BAddY7nK5w7EzkL1b+WKmGBD+oyKO4eUu7AD
nEyVNe8kXd5N9qWr2FywtqZoMFxQhCWbW7bU1019NjixHyAkkEK6PGjdWEcBIjUrh1yjuZ6eOp24
QAtdcWIKp2EYpZlKxShk/aBhnHGj0Tb2uTJIoN8Vrd0ahwybameYVSF3Kn9TIZL9VPBBCkD2tZuR
NjmkVwsm8kcQRuS0wy2YpGxzVjM9D79i2kL5TEkR9aXFrxA/nz1ywV4kM+cfwFOlAA5UIDvKr8k4
LnbqZ7ioJBipA128xyKVtCFQFvbp8AofcNVsf0fZF517vkVvuavkPz9ZsTOA7CUM73r5GApL+cYe
eAVa2h7HPZ/8oI0esSWqiNcV4nwu1pkKVFbZ81c71wcCDFieQAUn/96QHo8XYULFQuJABN+GvJkd
SBo0YwPKYw4j48pFEttk2D2tXHHNtwvdBNHh5qI5Lb/tpXx9nelO2ecCznShYsGXSFTx9mMPGdQs
gshfsDimGQyYg0/lsEOi8GGDxQHgFgN3cG5LEvOjQZ4tgvt95WfJK+UliAZdUaA8klV4o6Z8uVzf
VAGs3YXasG/vzNF8nNcnmPJzZeCuocXuApplpCDDabHpUkvQxaeiGfp/idA0U2lY7+9cS17cMrmo
x3eTLa6NODrSrRDCKEpPM7xVfJVgzEa/O9eCAub+13FIz84Bd7EC4Bpu4fssEKEe8hN4Yepqmou6
G4TY9zd21JJC5LWHPz0KLGL/Y8zzJ0lBUKugxitSbVQKlKshSbiVtU/KjXMioEuX9mSGnNoCuvYS
ooPIvBox0SaIWUNz2BQja0+tUE9tUN+4rSfIjlwRs9dCck+5dh2dGz1RSjmbexzmD05a3cRS6GOj
9buGNIKhydkdjbO0IpxIpDP+8GYWDxbXLlP0oxRNr4xqUV0xWQH3qSTs0fdXPLNGO6VKHqdisP5s
zg3OO7ZCGtGvYa7Ja7iLETjW0b0Dp5YNfR+c7Dn1ypPIucG8H/4X9x1858t5e//+dvvMynXTq6Zo
puR6fqXlHQzH5w+B8AiRF6AtxF4EROofrdtDDXQ/2RRmuF26V3ISY41WSoj6DU68oQmL8eXv9oHt
1yZZmNEGTjO5P/s1N3i6yPJmCprHGdsgQ3i6bESvtFrbpVyINOzAJqgaQNhxiYb8c8ygTNQtOud6
i75PRZOvSlMveINklr3V9JlpLQYfhd/irYfe7Q2w9NrTCdxBc8RdcP0EYi4zZI95nsNSyYHG1DiS
GiQCDlO6F+TzvsIi1y7dCd5BSY5eKpHIz9ahavincyRdmx8RMIl6oIO6tY1HyK4bfM5pd5uIYYqv
Lon/5L1IqD+59JNu8k+Ck775vlpEn/Bk7+qngAQMQijqqMaTGsUBYjBraJ/vFaVke6IkN8uuQtCB
p/V89l0KmTWHo2+T3mt32daL5hZuHMeOIDOEaNutOvzCWCcOD6VGnzUwooAgWN0OFJARnhQynfgn
h0aT8AWCK6qmkRhMgzaz0h7lo9qN+5Oro8ng02qyqduBx43AIjP5zHR4CzWv06SOK4U6OS5JkQ4J
w5mIpAXBlVhb+/NCivXjxrhZpVZN+nkHvev8XpBHmq7HeVF3Pb2WZ9yjudEM91G2tO70M2cIV+n2
XInti+8CQ3UWZbOSBurhgn/TwcJ5e0Wo7OogJDzqhrLpAt2qguQuxoCngYKRiTaVigwNpvZwyBFt
wdcVloyRm8BYR31bRJA6XMHJ8/T7xRHr24sfW36agqr8vzrM4co1LxzVKizcsP216ptB6xbj7VIe
KiB3LTMCZ2ysn2U1+8nrpyWHvY6gUq5baZBsQ9RRK0vO70wAUQDoLhXJrm7R3JETzadt70dAlAHO
i6Z6RpX00hAVImS7tv9yHfJSradruxbn0noDrgwdDRnqpoK/EwYPIdFJwoNO9VciZmI4DKqFs5e0
VzmDjzPkskuZTbDa3ThkCUVxx+lYuFxtKkjpaTj54r/vbHxK+A0kET0yFyZthL98RcjR3s6lBheE
85sVdNRmUE7wanVGwnK3hBvVaKFcj8xFB44iH0a+RS4cyyd2grOEbLMZMggRyI73T5mbpVwHckJa
4FI9z9rjwFWtyN8LVTPl2o8hn9OX5BJx51QyZ482kYshJJphOoLhSQ3XbIrd8EV339itbs0RyBI7
rCqCkElG53AxwZM4ducfoLs/YN2/FqvgJZwcgyYsSsHYmKqvuP65vetlwk2xry7vpjHjGN1cYHbm
/6v63fsiIJxxcOPNIXVMvt4n/YsM3y1OkXR99vgirKtffmmDMXhT+3CgJ//COmURK/thGQTpv6gt
Es/y4sHTjVpqQ1G3pz+aN5JdrcCQkin5CdpdATYGFkifb4FRIjyfxwZh+au1NXYL42AkmR2i/8Es
KpKWfA06R4gSFRUvUKi1OC/mxrxj3CnU6299PIDX59efYqlsI7jqubtZ26EdLLVRMIsxbephZKaT
yBKxok+2dV68H7vY1co+z9Pahqf9v9ryuNJx0NdS5w6GCO6+kwkMhCUAuz2J4q4brPI0YU3WEIKR
S9KEjvnm4eebQZ6+Xj/afWwahS3oGT8qy5z8pxHDxp+YwiHhl/rFCryvwnj+bc53V8LUjNtJudtM
pOreU5MJ2HKzjfzvihfLE/hxvXNHAqvGgQ8K7v/++L2PiPrmgHQ8mO3C5UptD+VqvmH/IZhBgXP1
nOq6AO97KVOZnuWsPKoOrZfwQpB0WFsGaYkkZERpC+oc8Tx7JTZU4Bty1eex3GtdIe6YdPmn5hp4
szGavAZ9hYsLjLswqCFsMAuceQ9fbxt7yyx1MIsbZbfQc3D6V3gYWFolbICV3QO33rMfWEYhTS2v
DU9mj9Qo/ElbFGtrPm7+e1xBMd14q8uIo4A7GwC39PDbcUA1TecHMKfh3fJy9dxjRaaw2CvkgJYp
UtqOuCnHzNZ83dKBrsYuLpGp5a1uU6LBPqW/44twn1hrj6Tw5D5ebXMR3DYKnBf8sPpB/wUh6TRH
kU7W+usTl2z5zjXs8twnU2gtjPD43ror/yFJZGN7yVReNEUyJBdZNw1rax1LlwrOnKR6lrIaX57T
Db1z2OKHtoAZt70PJkH/pT2KIxqB90sQ8i9xj9dlegf4M1ASUoPTSn7FU5l0zOaEehbZoKtuIiBj
Rv/guIU3CehCDPI9wI3gCgYNiTlW+BxTa/J0qQ7+Etta+wgywZ5BLoxL/HH+I+3C3Aw9nsHxqY1u
dL8KDO7b0qZ282nOkLGjLRwnR3RyGFrRSTkxp4fJ6fy1R+0BpOKqWyamSCJnYqFRqcU/N7xIk7wj
udxhndxOoRpQz7+B14l168WqAyRqATNT0N6DdpTU1w9iIdHDNWskav8k7wK55Sa1vPuPRP4fG0wa
6/KiEElqQ9G8yj/nDFZNx3KI3TPu47oxEu7Q15/QiRIbbUbaVLzs2OkadKSmZkqlPQE+Wvjqb5c8
cKOlF9e5Nhh7V9x6LiDxF0fUSVDURxpnguRIl73QiOwZjtgLk00Z98leQHjdoG7xo5BwALMytkfO
HZjK2plc/uGekf5VufO6N903SfuJt1M0qykZzAg/bl8dyMTAhh+H9adN9Ps4bqyuCOxvdOzpIJiM
p0rAI/QIgL7C5ky6RJPFESIbgdv8WuIkwHEDxbcO16x57RXQHpuiaTbz/rb+rfaROyq2S45aJ3Lg
QZ5sMrx8Ls+y3lD5iSA9pOc1XEMjY/7NfJZVYL1k9ZzrFpRuXSHP5CSkd98dAZ6c3V7xQxEkB1gU
atEruklXHh559ZUm2QPU/IeQF11yZWMSkjQBzvc3VFct3UImpPbqtR93g8p3HYPIqX+Vm50RVa38
Vh5i+atqWZbTcqsJ5h2zR+6cFOGwXLMfoLHj0OSXaR1eevcWZi3H2zqMBsW6T65wl1awEpTGCtA7
1jto9tjVjEjvs6Q1FLFrWkKz6JZL+kv06DwLy+4pUMfdjLPJc4AV/AS6EMPIQAQU0WJDCpWCSCbR
NqDiYExVRy6jWvI8T8Al9DhuABXBdYr9lhm2vsT+iuUKOEygNvKxYQCfxCLw7/QNE1kcRWlP9oeM
3m8jMR0Ayw3/45UeZwPaRhZNJoQmw8wwpkHk5uAtEOQ4Gj3umgux+9012OD5Wvj2Ts2SIwjmPOJP
DEgGzyrT+cA+1ndVuoNMjntSwKeCUNtAKw8lZ6Mv2QHHy1+rh+GeIbDUi2ox0pM9PgxYIaWfLSiX
fIzrUGFuFxLBysCHlMXjVaYloBDLYT8d+CVtoCf64wzLAI7t0bjyG2qMlsoTTUYIpNvEkAAeOVvv
ULyOYSx+sinUg/jL2zq1/T8KPMo1fJz9z+D1vwwC2V9eiBhS7SRKhuT3sAvB8at75S7x22m8KQ48
1iSQEOFoyZgzfxGefHBRLpafSvTGV2hIP+Zo0AHyJ2u0VkO4uj74PKBZ+/OSGTRcW4ftQXNe+Kfk
hltlMSqlM8H/IPx36LMxnh43HvwcpREeuWFWAWbQRBeNnzgeWFrjMqy9QOMow8hZp6Gins6HljTt
IxQJhZ7UWnifPivVcDUdBfca3e3nmf0U+3oEl2sIdcWnYwyopJuUVTzogzV0HmZxmUtzu4a99LXX
sYCsS8dzVf/LjKWwdQwj/JNPoGZYVIYbye0ZW9lhhjOaUq/tK6VDS69bVLHuXp/VuoO/LiwRLys4
NBAYXtMJTywoPBI3dPfurt/G2WoPX8zzl3DlrVApB0S5OWcVRwsMGLD8DvzMkTXZV7gnp9iTp5TQ
cbqPlwuYYaU2a94pHFhcGXltk5BQ3f8G+rm236OxQIVBnAAeAL68l9bWkT4PcGFcCoVCDYivyrAY
YCJOtkK8fuZPv1jNgBXt+ZBfsDo66Bh43DCS7Ou8jGJBl29QfqeuUauLe2fEkCTLxH+YFAx4Khmp
I/D3AZo6cvOwzUu+2uNPhqIZoOrI5YUbo59DZcrnlkjiLkpkX6Fen1qZNOO5tG66lsam+wUSIsnA
geqe/ZzsROuV6acduYTbtDfAD2DiKlaBtov6KwHVQtCBP0dCP0olNmguYpd6tQitDkPOfpoktZjv
oTwK3jr/p7xfPeDDM/KPVbTijt1o4VYZ6f0THWoEcwKUyqudn7wS7oGz4CTWNnyyT3seLr3+89Q7
a92syvZHX0wTbzc+IfhX+X5FdtD5FXqUSpm1/DQ3kGej/PGYW+4vMnrblAPJ4gy7nGLgWKg6ngVT
mSuB+CalrDOD7Xy3s+7bNYI7npgmm6O3NnWx1BTejwGgtP6+DDeR7DPcUSp0TwnQwh4bHx2/cAvU
XIjCq0Oy0f2JRzdQHBKYP8r8COTpiKhEe37aKQxAkpowcXvt2UUmZ7gdoehKw4OrGT9G9pfjLP/8
YG1QsMM2hsWJXvGO3W6aTb52ZgyMK0xbl4qi3I+f6lYVY2Bd53ncy8RZNIOjee9ltWs9r3iCpV0j
YGHDR/tdcQcEGTErdszpGn6f53RTOmmPKB1aiXw6pP3mp17W1jSGA3xkpELQP7oesMLvAiXD3z5N
CY00eo+ygbpVSvZ8iuJX50DOYDptHxCqmT5hmeu4u1Q9sdBsiSq/GXNSBbULXQshC2AFC2Altifk
ajdFIGwBXKVWPecC9yHkbAYX+iEVro3ovVD0zgJ5chVJA5Bw4tjz8b+IYEJfv5BG8oC1NI5I4i2y
6jBtpm1TRTjCyIZMBbVYXTUHG4rOLZwOVGOLbTLdRr3qOMFv9Xw0auAYksafJ+d0scOURwftYfN0
FbmtFOuP1PhkMjd0G4Z5nuyog1+X3lNYGhZEmacU4/RGYxE8j+9aP9WRZKJ4BGvekqEJArw7NT1z
hBWziVnxxmtp1tpQzCYgq1s+77oKj5qF04T3fSsE8pDTzEWzRK/2hDJtKRYDLt+kHsKYdJHpcnXE
P6tKMFEci/WsNY6cseX+x1n70IvwCssAoWTNLz0R55be+SGsMWkOq3GZDsI219FH4iKTONRx5PtU
DBqXY2PdJ2XYN178B0iSDa2L3npBYgNP9A5N421vspC/nEGNxS6OHx97JQmbDWpT0TMGSOa6qtzd
7PsOdH6Rkhes61Nf3oVTl8nWbG2/lQOmbd9lO3OrnG6HiaHdSS6po6vup4VRSAcB26iwK838IYHF
w7bkNw4VpWHtEGlWoQp8AZn+GeJfvv1aOBbnhdkH1EulvAhdL+ESSc0Lp14Bu9OtZAMPg4CGHY54
4wDoOj/3OTzU7DSLIKjynQsusJl+fm8lepQDagHEKgRU0PpUOz1Lci0K0BHZuhabYtW5OgefHoST
bUE1mAJ4Y1d3uxSpuuRcSfLOKI2tH83OzYCJRUiltQs37cAVXyzKDHFCKBD9x3GF2vAPA/tMQEH1
MfeX+6nqzQqiT61ZXzL57Ib4k0LE2Bgr0pPrNUujIYco2JkNjZchsj+/xzD2aK+kgUhsZCeXObY/
RErDFnPoSOPFDOiX5Mg3gp6PsrnnimQojZqWcyR+E4Yf7LnTHBVOLfFOfbMT7cSimziEr3u/Wzad
qy8anuE74YdYGFGIjL6R7sYPkjxKspPhcOKIJ+9Zu1bE3QyiowA7Qp+JvNurSF+iH5nd79oeciKI
bNcL01LUxxrE+sNci0zw9/flVFNFUwTkxH73C+U2ZIMZexRD8hbLxmbtsKDByJdrZiIx1PUzjVOd
IKDVAxeOq/f8v+mJFGE0zXO85M0M/o6YuVyORzOKQvyB8+mUFGxZ8ZuqlGCxLMwRMKdgg6ULK5D5
aT3RW7xOTSWFM1uPPez7hpMaQUt3Vd5kujQdr8mxBoTvc8fy+nhL6LQrnQq7oZRMxiqXdU+hKnIg
AovVkY4614GVSmwdfkTxBGOuJI4oHaUcQza5vWdUd4FdJeCtBds1x89VgSuAzKR9+gK/dD8+tS+7
26LGZnbZCTzKx0QVN+b7rtgbWbIGNtQ9bsQOxktrr1/t+6mZ+3lbSodOiSDouW/TjT0vUm6furl4
l9/x7QnSPKZORZqKlDfhamVjrq6YJj/rYOVZuGkFQ+NjWzMtebpsogMKE0mhPq0D97QQqmA9Co0Z
5nuxSuhhalOx+TtBJY4fx2te7OMZr9SzI9wuvcoIcWKznbbqIiG6VCcKlaiYYyk1ZEUT6qn1ASJa
ztbdEn24TZujAD8G5sdCU588OLlF/7k2pclPAfrnrwgHii3kJItEF90ofl54qeaGiYkGju//U3vm
Dfk2vy2dCuWyVq7LYxuJAs10Cs0bJt/8Ydlu0AAd/mDm2S4V5rp/KKmcRxzbNDqZEksfi9MRgxK2
msbPMJAP2BPBxNk+TaAPSQfM7NMpz3ijmVNPz13g+VWIOy3pmjISRfGWAj8DVuMsygzr8saDn3ut
RkfUfm7BKx5Q/2V2i8y8QBUfvEloa6UWsHGRbmXYK2rGG6I+CexzAaNeMdTfHzGT0lh0LCKZdf99
pHwN+XvlhnJqxhNAb3GQX74B1KzYyltxkDvWqXR22PEKdcPyE0rwrh04QiV5TClhQ9sOUfAYmqoF
XgHMgUEBi/vbDOYQexV6BIUM5qVFnKUpk+kcfVCCoOiAq/r7HithteuO6kPCAgGDYSS/PAenOSqP
MmnFuRM9Mk9RShFah/nFG+dSrJba5nBBQCgYdpOJxkT/1iVxWBhBURi2MepoSz9PFUYEI8s0KFRR
mNu+xK85FfLBALLx/AjiyVL4eozF95rWMhTLSrLw3EiVAGVIXnETyjEptaCGlZhnHwf+kaibykiZ
4GMXw/trU1558boU/7RV6agA23J5POSYWynJPdb73nwbLhRCPob99G5vyNMHz8f5dcNPy5xs6N0m
YuPhwSNGCnHwjhGD/2de7fzLk56pbS2LkQ0Fbqi3Vvc/UvtO/eB8lngeBIPZfowh7YUAOeJVS1EV
3UixgH43idJFOBE6DWr4LuUUKFV1edVTskX6lXom0dqqPB0/ivAzsjE6ROg6ToDi1GSrOmo5Bza0
sZevdHK9OurijgFo4/2IvXp8xK/l14rn4NXf1yMPO0gafU01I5EZOU0Q8ZjCNeMBidxgGb53Pj/b
q/yqRKJnbxW/kP06w7HhesBsGtkA7/z/6OX8KIcaUig8Cfx7LfrTkLt0h7Fvi6M2Bf7HQW2SrvUX
TYm7rK4yhuBhy/PTLj2pMSp/H5J9sCIGl7zSJqktIO27d3U53HB4hVuPxZwBUOp1ruFkQyqLmwD+
w4iZeq700aszhnpeqsQcRszVtFi2f+0WfTy8Hmv03EL+F4Iv2TSbWY94I23PbMHHydUxwlAQsYT7
xwh1Uim7jLgGRNyqljdZTp6d55lbTz8XRoDX2yWeqMmqlYLEgQDrTrHP3O8WHQZu1g9tGNfv5Iv5
85DCwdD3kSwmVWYdnM5kfL1lDOvICGxSkD8V7HOEIVvHicz0r2iATlFBeV9rNbXtdXfsqHjcI4th
EXvfCdXTQLFSdWOd9WQonZ+rReuvy1yPloaiBvjE6w1UCvvwRl2g7bY+oftdQmntpsHV5Hy9E01G
5OLP5TEwB4oMDNVhjeDCHcg+Sb0gNKneqYcHsR8V7MEPrqvm0xF/JR+vRWuZZI3wc6iEs5cce8JC
KQOb33xBWo9h0k/4g+i+9sjav67C4bU2PChSXHNmmQmAa+KyeDNW588udunM2VrtFjEnGFDthetx
JQWW3+HxJWNaQPIrjC0ll6x+xWEWPf9kN2bi1Nwe+nEt/fKQU5qE9yHRzn7T9HAEbEp6SizM+ucT
WEZdFh20m4hWt5DOORgmZGbCLoO7d8UWUWt11obd8KTr2UVuWv8dZuSNoiyIZ0bS98wKxz0QGEQW
fQEYsdMWLldh+8YLAD8P/1/3vDCQvySpdhb5YBIx+6m8wPHeufOuZgTNoylYuf0z/hLw9kbu8+pF
nsjzgPvVIL92sKDqu3LmN7LxI6MELmIfZSB3QqX7mncg3z06ol8UbRTGVOFeEIsN4dhKwc2rCYdn
Km+TrNIQVL7Zxwb0G6JUtpRvTMy2Mdbwpasji8tIr94u5B9CBZLNx0L8kdLVhYvAh7p4Kc5kYr04
GjycO+SqGp6biMk2al39n8hxLng/vjctae9bocVO1bg9kzo+G/Myf4d5KYT4XGZXIGjv60IVjfom
MBZxsE5oZ74rturg5ZOZRS1rbJs1kNunSh0HRnsg3wz/n5SlZ/NcRNQ8F869Sj3rCH8EHd3ik0Cr
ChcgWCZAWTa1pRLkNTX51axx0cFJECb4JscvHgU6WYqO5JWlXk4oWLl9ju0cDKPpI/+ad4mhuqNC
3M3A2abZYCRU2COXNJSW2d2Ux9tSD+k0Y/iGtD23M4gwAFCa8H7EUezLlWdSdpHlFeBylJc7PHPB
cNKW/HRpAZfJjSiR5hvckAlH5U0AyMLo3LAWse08wsfgvcivpIy9u+mQrSpJgXtlfVC1xH6Nx3ji
a8iJJvXQtYmJ8UjdM6HGd5zH6381EdxghtnezneEonsiXnmXlv50RVOq+hmyvKL6XBS3JH6NhisU
BBQz6y/a+FB/h/h5gkK8u7FDQULW7VJdbByJ1ByA0zQxTGzYyStv7rM4GDIUH6xNTkFh8PCnGT1m
tqSzBt2mQrQMIhiw9ifo6FJp00wE+ySqNiCY8Cfl+Ff0zCy6vv1MeXz4mJbJUE/vzTRJOQd3CFnw
Csn3+9VMeTHGOw5Vo9BCT+etc3XD5ceygs55mz99EGNhW55JioLcHq6U+irCTTFHvPFDD2E14V/N
atmk/cooOO1UkWH1JqvYVAx1voIlGHAPcwnafZ+ZEU3B7nxmoP2DRRag4LUj1M5W7lgWODJd23H3
EPclYApsFKPBPr7839FZL4R+K4BlLriy/2eGpvyjm1b2MWGekBXY/T2r8dy6WRlrQ8l/U63qzunp
r9RdlNwXOJHH2TtpnLCa++K4KxxZTrmRrqQPSVwlp13MAR3c+9hVKphSog1qtk6egYou2w9AAEcX
PQrt3TwaoTsc/+m7I6OqKAuQG3/ewMrvX9VHuQQciUezZAPzAsV67IT0TPIFSoK0WzOFr4XFtRFI
SI0ysN/VBY32E6ZD0ymusM2B+1VyTRm24ReaStqyH1pdVi1nmXtv+pmBmvwA+bO6Cmn2YzgEi6j8
DQgAFfSSHdE35Y3334yR3F46B4Y1mt/sEYvG7B75+LMpXc5JIqsX2dC2F5+DmIZhxDvrR6muspkJ
db7H1NOuBFLhP3cXgjvHW+azGrd3/+JFQhCdROCGZ81mJ6dVE31gONmASLP5pvwX5GXVM2L18F66
qm9R0f0xkuiY1G5TtV0skmf9cnxS6fwOe+INLO2O5+Uh841GFZA2nDZwiQZSJoeDNFIRrRw+suUo
iiCIPMByXGj2qlqbBG8NWLk79hqEf0pX9nXfVIemIluGcVu1S5JTtgi9+DNeQGrsBxXWdF+ae/4t
FCMOeXuzn5f640OGVrNSJyZOxB71Tj7jl9VE9MNX371q2LhSPbQjL8XUFctVfRNw1YX0JYgnxtCi
xVILjtpeJtNugTI8erAEULI2J+eUSPVxPqV3L4LONk4vChI+takN+2MqCX4wINjFKMhBFosikO+c
mDK0lNr7Y1F1lHa4Aewh8HxrUhqtxFrXRTDsO61AdOJUdx70Hn3ijX6qUVLqcK+prypAQgERhes4
uVVuVaysdvBDkOtxrOt/CuJG+EVGMXaAN01UAGPom/FyjnMsLF2i4z8kGEpIl9zv9Gh8HFZsBiJr
2IL4mjRbSxPmYjPd6yW+PgtOeJm2YyQ1oYgh57fTb1YozcsvPvjLKu307eM0Vct71WqlkBrvyrAi
INaW53l/qIGdYVviKSB1ICmjXF/80O3T93lgqcuYrnp7iMXgIzVnCOb0BzS+nUJsU8na/bq9Bt5D
8J0gkd4K+hedpTNaOU51Ijqb/lMrLa76ax0UICy32Vl92dV7rFyXJBLW+HbJ134Iixj5SoZ+A3pm
9E92EbpPLOTFE2VLSRh2VKWEhBCIRWj/xofPcrsN3vRPCL4RRnKcFcoFrjSYN7q9uYgfsNiJbqZN
G3ywSwyyf7MtTpZi+H9WsoJSmWqpXOTOnPtnA8xHj+mKdC3udDRRDwWzGOXLAB/mBFj/PIj4iJat
2hMUBSmdRqqTIBkMLGfNxSQVzNpVkeb9PxKXizexaZ4oXjBEktT+CNPm4NxG1ACVlyVxEM8KJFrO
HWD+2vd/KIqXlocbvfqyNpjkdqqSPd8d3kyCjy9b7dSzis3TEVD4vuJgJGwwjyvQNUxotbjU1Jew
BmQ4ORoqhmN1jaogGF2DrQs4SlArUIoUaxMuzEOkR//RHEN1xuhqqPeFqnWJYW5FRNSpLnaG3uT8
fGVYiw04I5z11UtdGYKCPzL5ANYXhfAlI+nT+Z0SGmKf28sDOH8e3gcaeO24rmNSns3hQvXI8A0F
a8mdsH5MOwBgUogEk96PvnHBaC/ybgm9esi/QhCZeR2gNfnGJk3+QnwXAIW6F1d925Af5uohHpLJ
N8KAFikXppXlls67RhgMAwTg2s/98BaUNXS6qFMDdgOK9NrPMFBetmBPJq4G0bRHA60MNIPc8HYI
541Meq7m4LkfqKwdUUzXdlGDZDd7fapd7YaqfVuzq3hZyiTtUbHLA3Xbni9ioFLRWZNwRu9GJV0r
2x1kZxlwaxWXeEClf9wWAPmprPtaqFT0FY0sjMZ6bnBUONWVzqa6tPg/nF0JJXVARjH8mB/XqCCX
bNy5JXC/u4GTOg8iz/vNdDxq1xyteJMZlz6vQ+iV/PHb6BNRbApBFxo50SqwOx4GZ4pURcoL766u
5g14aAgZCBgWAwmoGt/r1bYhMa+I+OY0YltDvhJaA+AfUHz2RBSF1HvWWxapc0vS/V/L2bSkuqDq
8WE6pgjxaf4XY2HZKQbOiHp3vbiYIox532baQMcOipX0f4uB6pBGpPPTCkmendR39ct0mAo8KWc1
nSQbg1x2llAaW4/SR6ykubFgNTyawBQ9Xqqowe7pu2z+/ta3mOjdDIuxS4edCxgYCRP2gejMPn28
/7VomRVjxEiVjbTT718zJpExgcj7vtjbhXtXJBIQF01KvhNhnaIDRuLWAGx3xv8edb1k93sQiqsj
nkPb7p8j5xAs4go2G1rzJOnkP4jlFjwa04S2CSSFovuHWFsBqjcEBELjUxDBxh3WZTK8QmV+y0J3
gfJ5IVMnOj3ONoT1G+c+ynJxdL87K31EuLk8msUXm0xK+Qz3X8v5pDRoJuHOuG7F2QfZt0Vmikz1
BPEGI44jUDYrRLCeZgTplJhsrrG2IZUsa+DnE0R5AsFJI7WZNCYjy1hrcsqH8nlKr7vNEj1EO3Rs
dbEOPVhdqSf1QZfgE9CFFdbBymJyAG5n+pZjfEN/jZj3uwLz4/H+uqe6W41pO+zV+AsPK8oLh5AZ
wIPv/v9qu33HTpOv/2+t+Xnp2DoJ4PfpMHlrcehl1rYR0wEh4/cdh9G4A49lIfyK6N5fFYDumtYv
CB9xmHK0UJ6yzaWFy9kpT+GfgC2b7wExNm+gquci4GPrmav1Y7f1xLtwBxJf3Ff04/EsbRYVeCGF
75eWd0qfJ0pZ3rn8GSkQmgyiI6tbltOdZF2AtGjVEofWRW08yc5fiBlCkfhpYxDcxPceZs1j4lrU
PD2R9RhkfSCYVTvS+kWrXtE8kZVy5mGVxEqRR8ZQB3oOR+s6W3ZWP5cFUxD+JOsA43OmhSe4uc/T
9s8lD+iu2ba3YIU34cNXNsJCwYpLVPoZk7DW0+q/19czQIoZUqKaaLoH/VJQvIGek113wu+oGdYK
qxp541HjILHoh64NPYH2FG9VJ4n2RKnLgC1H9h2hsu3fVFdeu6m1M3l0JDHFm/5tbqHUoAQWYH6K
4FjRGhnZATVStZ08NRWB698i4xQzdQrI5KGmvdCcilgDl3dPkZYQM3YZaBeiR/bqdGxtXyrGXK9q
Z4QuHS6pqa6k3DT4eF+SXdmRhlZL5m4epWacFqc9MG6p6n98zLihFcYWSk6cMuJfO3GWNpn2N3j4
ruacLNHrNdf/TABVALhdyIRn6/igNtIQf8metyuboLt2EBAJ2m0vZ6JD6d+lm19CLV+ojkLfDIUH
ytu5slTlaVfF+Oh+wXugwQgeh4rW+CEO8oBzfDbk0CT6IpZhcWcWkyRUfQsdAG2LbuQJgkg4C+JY
ZCeYpY4e7zUgzrogO3Xd8Ln7SO0f8qdHbRTNneKCdv/AQHcSwGAT2IGDqV+o6QgZjmC5n5znTNk+
0VksC9aHv6pHjv/aKYysUzBGiJgmHqs+ezbUN6akUvIOnnwKyx/Hz168uiKLEDmeY0JlM3l92fM9
yJaYzliFKpQn6WOpHH05YrfSJuGFCQJJ/CN9D9fyDDCTqhwaJlXTmr9i9ZPzRmpPV/HUYi1KKtV2
4lX0iYyWwzHOQEaFegrbHlrZxhy4QzPU8Cmb2pYWy0qRsvAzER1++l1ZltVwiGq6AOsQy16nzlyo
5BCTf54yjyUimO3IoIkkjhzGEVG+o+gu++/nk6gXk3TeUOABjSpCMBK62QursbrSPBLnfKuj3O9n
wu3TTDkZCUNeRwXr/+HkJD9BLJr4GoAp4cuv8+VCMrthoQHfdA8Q/1mgN71ybA8/CcoMLXXMmOEu
AstxR91OvLQ7YoI9U/dWOZDvJ0Ykc31RlDIjVxFrtnqKpZdJBj4cq2dJ6XkwaoOX/jhpVbUtoV7X
v3SRuAZotoRXbEY2mznFezBnNhl9BtvNa4lZYr9hVrnojlkINNlU6rb+w2kTIcQothU//F+OThRW
TuPh5F21mS4m4bL0/oiJ6+GEmDn2nyQY1aWmv1TTabE6os7nkdy24IWVM5IjZud3TVzI7vh7P4US
+MIQBB23/72NrWu3XT5q5aiz4MvAry6sRL6USDtQROCgnlIiERdxos/uu44LtgFH3sqWPLz7hRZR
cCI1OhL57XfINi02lYsHKVRmMCYERTCFsH5uu2Dm1PplDNlRLZHNIWfys7e7ryJVryicr8NE3VlG
5g0U4E9b8blKF05wI67lFpmzZehhACQamfc0WGdQt6VBJyfsg/s9xbmwp0+oT1JKRk4LXqgwZBJf
hXiRLMyWIE1KIymCoWonNaBCz/J4nEJebJrKswOcyp7xP3vqEUxvu2vrNdRxqiaSP3jZvPML68Y2
5g/hk6HHmNL+vXVSsLUhZoqq53aj7PwC1ItbmSoRkTkf8WCu8T0Gc0JcZyycOy+VjbQsPhj66O27
8V29g9yxSWdt68xj8KnfUxnZ5UdT3YjYf/I4rlxn6ztZuAUTPZ0i3hSIegI5X5uxnOQ8pOmwwZGz
uFVjl5IycGyDxagTy+Mla2Vebw6BDP0T4lKP/+URIq7txkutUBVswG7y1Zgp3DoToNPbYh7fFHT6
8cUPNW+aO9KQqJ5dHDlmislpKPLn8EKTnMzu9u9GhICJcvhbh/gPDCqTR2DM8Ok2DoLNKr54DRw1
4DRNRtqlbdUp+WLnKtrU9x5BQu8eIgyibv2SrrNHWEZVO8Rb3FXTVz3eF47ScJOeZOuJH2lReNfQ
qu4ySDmcWdLOIXKDxBYRL3BY49fjh8hF6Tj8H47Dvl58YqxSWPN7k6toJm0Wf2mVWqD/POOqEK0V
5Tcz5bJiTGAXnkU82JwkhJTJFWioOyk8ELQd5MGyT839zLesWyZdOVNcY7zXm2vqj4ucfOgN0V8o
1ATeVD6GZFVmamcqGVuiEedgHpm0TgBJ0PbsNLb+Im+13/xPZjAo0aa2KCOTv7fl782s7yG41L8y
n4L8N0yDyF6Kqn+qomLV9pctV1P34WUmLSfKigi7RVD0IInkjr+RMAR+8RRjNGsInILYyR2QSf3m
DY/CzjHbTN2EzbyoC52O5vvJHxY1bGnlAtzJLNvImB2SxQXgOL2rQhXEgYqT3XyijEpfRe751oxN
XoB2Sc2WI7S6kT/vHd12JvhxhlF3xz2i9B34nfQdGAMlWetBZ6b7BOEDDUzPkF2D1WH/epJC2rqW
ovcHCHAwTxqljKAGtNVdwx4TeSNC9NB3RVt9y9CQ++p6BcYGCN2YahTsaxDKtQ25yi7/Y2kHbMwC
FBnmO32RbpQLXS99pK20oAGprMelcJ+xn+TiH+OV1tUWK9nE09BlsVufNr3r1oauL802jgcakyJ7
Q4s6jBzhwP5Y8TUnc6tiXYoONumsemYy9nA0rsyfBvF2M5wBZNidrZUey/uWrxxaKyDSoVZHG6Wr
2uplKqs7yop35fQxTWQGpVSYoI5zsJSeTS4WNTwWpw1hDX9+9MBU9eqnHyQHLzh8rPtCg7RgdUyk
fZJyi4COvcTgKIcuTW+LrIYMMDlZmCJrOz2oQqcs+szPlw1x9hKM6skXoiDNqjRRSSps6TSF98Et
28W+F8r1kgaGTFUJg08SGbOvo3naSenmgtk+HSfDhg39beeg3xvPOXr4vrUdxAuE5chGIiNqppzN
C+mNA1EL8CIU1UpmtDUDxmMNzLSojP0rnncHNOtqyYCXGbECoWO2Q0bV+yx//gwh6zdhVAWZu5WQ
34dCyL4Y6R9zkDShV+1Z+rOD9C79+DSWAzi1ZvnWt0NWGbpplHWmfoGA/h/fb4lAdDeo1pmECP6v
GDkUn8Tt2jFW6FDWgRRe86r0l5/uY4JGm3PgORF85QIZ2lnpZKya3dO3nJ4ENGdZYJ81T4dCwLgW
3/3w5+CxFVFCvmRTAtrXmfZkacCxvWA5sXbSGdoELwhjwc+FFDEUxmwyYvnTnQBnW4/xqowD/42d
sgbj7/WIAtLgVLUuXwTV5SvbH4Yn1wEpsGwWXyYW4JQWQENBPe8SVbdsRclBtvBLXG4o/TG4JvG/
qe5Qc5Qa0d6QWmVLDwjAHw/fCnO+kbhQ7YcZ5ivan+Ct3knW+d+1LXNzGl1WkSRLa8zHnt3D8a3x
9NI4WXzQ/DhugdsgjQBm23foCwBOVMQPZxMjioJkDDWbTaK4F75yIxjQlvdUdop2M77BZ/HbIlHR
5iJDZqaukSyt+YsCH0G5nsOf7nWMSJf8L048oZ0gDWacp+wOfZJfKYXPNdWyfLN3V3lA8wZMLin6
jJy5KhlUk2Jb7gJHzd6vYy2escn8eAeK7zkV4vLYmPZPHPr3QPZQQSD7Z4Xd2wELQHvWHJG2QozC
WPVe5Iv5yi7JkTizq5UwFh5J5t9JqfIquaLAhlgU82VOB61A+cw6tvs6KRUADiowNuv4MOjFVDh9
rKunXKAQhd+uyJjLx8AJnon3LtmJietAp7jCVURS1cEj1dsRt+qEIbxu/DJrRDWtJUTlKWav47dL
DxM1Z3C2xJqt+04SlEojVL/6jV9Fz1ZoDkoxw5TUhPhhKhmatGv9gYyM+vuipA4pquNziXhQ6Xdo
sh80Mt2YYhmuIAHCYQdo0GfRDtTSU+9ZfcNEkXaxMHs/9Mh+JyRgu7xrrWha/y8gmnLINqlEWVYV
Jt2FXT6RxWRHJXWDMS/YM2I92qYqiNPIwK0VDAN8n1khBP7mSEpAKOEjX7MzlnyoM5xJ9dVd4rcI
Wfb9AJCKNDRyUsYQHJN2+82DwhtSvFLlYinzdI7ctZKgkuFxzOp584PphtFUbk6lg8MwPvwJ75NX
8vUGJtMQQAZH/ZfJ/i4ZLFowIXaAVCCze5EhR9yfeD+5V5Ed29QHi6vouvFW9Y6QKy5dVs4AXd62
U/MeoKWskPM2IxmfydEwGKteNsl77kBNsEfyPKBaPWC14wO20X1dFoBZ6sV0vkzaPAqnEGAMaBQX
6ba9b0hGS2VJUaDC+HnyCR/+OfaXMdnLiZAZSebqD5szVZtsX6Vn8vW41QS0SFPqQrTWX33Tr0WW
mGu/ZV+PIz96408CNmDb8rIwIQB3/MDi2L9UskcKu1RAYm0HVamWBKO0+TJxHyej5cqX3MubOlOC
DPRWwTljTUfF1XxT1/kZT8dDNZspxM/WDJrol3KiqpQBe1n0z8X0zlRW+og9diC/gTTsQG7cQ+Ot
sLVsfh+YZt0gKkkuo84d7x2nyn7b4hUVhIWj/9Wy+jsvrmHzxNs3GbzOPSVAx3DSCElAQJYBRyL+
Qh8OukwONQa9lnGOFhatvS557Pxiflin2vJUUTw7bU5NmsBjEgvC6Of5BiekxZcNajxh+Kc+5LwK
8P8gl0mIJ1gGATyAbRbQcXRXMpkwqfqKJCiP9h+/DNFwOSOli+FM1km4fsdROPdceIdYl/97VL7e
2gjCdjCUFsyuZiAu/drXi6hWJjI/bu+Zi3qbvpdJjh8U9tGWb+MjS6hWs4efaHC/x5upI+vnF42/
/CY3X7H0+iA9W6R0Y7pE/z3EfLqZwe3YiUNADaDBJuS1c2NbOPzknDeQmE47IsKOa0FzoJGS59fJ
BU6poLWscfi/a+8rvUQFikdG8o9pa4C456fbUaLllQFxjmS2/f4afIsZFNJldfgezFBhtsag/ue6
+rRV1MsjBIh8LbY7zYH4SALofDBBdaC0b/wnFu7DF4Gamogkd3H2rnD4h0QxeJJjsW8kiB302Tm4
c1uoef8VpkMstHb9366CsoXGx8lBnbSfz89MeH3nfx8WBGqwj02WL4Oiq0Dtmf9XdFD77tKBQ7/g
BMwCcpPa1mqCdyt9pcmk1IzOH621lDOsMg0q3hndukxwHfYJHYXsIL1h4PD/vWNeO7AwufcAEKmd
H/3kCpto5/Pc662O2S88rHCZE5k+espeGstrZeOjq8uiAnw0fldNJ/zFK3wuimXti6B2nCSlWf+1
9yZEN5fHiDq8PrknELObQ2ZwttlDqzxvOHkjxBfBRvf9vgTabk9TQ07+KqbAZKpiCgFbtbJS96UO
ofdAe/gOvOXBnDwJH5Yq+5nat25pLFwXtz2GDnpxss4AaCPAVppllzRrGQm/1k+drle+rkDc5qoX
vbS6WMbClJZhfW/c7NWUnl0dobI20reUEdF6mTPFdrBl4uUrl5kQ7flB2lJILHNxEHpYCXzUTB+s
n0oZLmWz7XgMnIebmwJWwKlU4M2MD81aEJApLgR9es4Q3nUkYLJ00z90E4lcuit/z4ynkzMBorGz
8liyQ6ae1/G3KYQIAJg4ffnSHKAqiNuo2565Mn7IXt3SdUbIn+tTQC+qJTbXz3qVBS2hiOo3rSmY
0tRYOf/2AldZyiXtxvBB0MsufEoVDRC5l5hoTBhRPZeh+N4/1ErIIPBOdE+XNqyfMdTg1kl6Q3Vb
og1U4l3QljmK9LwSksXixlMaaS/Q5sth2PMnsyoM7m1qtbn12Dc7zQvJ/LIBW7KgbD3T8GgDfpYp
fLub6ht81iVT/uTgSk3UFedgwjw3oVAAX9oV38ycImPISuJuIgBVHKZZcd9Rb0s5fpQRc8wGMjsV
/wTr8dTbpm7Hbdbdh1RPiyc0AmaruwJmPSlsPNcaTYR5oLuy7kBSCa0v2HdTdRx7CAN3wISyoX0B
ivHpYOTfXepIYGI/ReOEqtX/ALTTw7+4lmO7k5s25l9TP5BsbGej+DKzCFuINNt48H4vtswyVnjy
GGi+Is8UuYh4DA22/uUL+dWN3X5D34btp31SY/wLfPvw9G7n4ESLmziUh2KVUjPDh0mdRwOx9pNS
cIEx5lQuHV7YB6tBxU2WnJdXY80A24BX8s8j2HOEs56LiYMT5v9RWVsFZzZ0Mo9vGCtVgeBb0m1H
Eto19mzXcrMYL5zxXAuPeCtKHqA7jEJvPpn+qOqNbc8et52Hi6UnXUAflGztS9EIukYF/8A+pvH4
WqRQNomtfAwTaS/qnXNVr0Jn+oLjS9EaHErl20wPqulDCzPRpO9QZ6lxedJEt3sUN9/xHtC3jft3
kj29G771YdLTkZ0RlTkLnr+//eYmM9bM1DSb8WzKY7j66GLGgKFYDdrtcTFh8X5nMYrhAGsX4OTf
Hmnt1ZN8oJKALMpz9nbXEg/rZdaVKVONnw7MRKf5IsyJ77LkCXCO1zikVCpBST+yFcqW4f/+AOa/
m5MbOcN5mMFxx2reMlI9gdjrqjpYgKcwg9YujBLPtRoePicMQXd9R3WO9RVz8u1h+KafYuA4EAbE
V0cB2Jn7bXLAUWYrPwrlHW/PX8JmwarZAP3eJyV/5vDiC9GFb+fbNFPeBLQxlSVUK2qlytv2to1N
pj58BP814beGTP7mfb4fmbn911PI1V+mTPhZkUAsDrk5pC8ZBvDe8voQwLCiejNsQxuGzfv3sdU6
tAMfAO0/602UkaPG66lQNjr/4oSjm8kjkO5d7winJoC+7xWYbe9X28KitvgeKg7MelUJRkeLvjSL
xz5yxVxuzGmmKwv70FeQsrZqVXa6Zpmxz4RqtaxLD3U3owMZIHyrsbwbu5LaOz+EbVqUhhKvnw7A
Qb6CfFt7AuWQbj9zvlYXrr1G/lvB7k5q6UTbMZJTOuVfjiEWyHj//w42SH/GlAr7VQu0/jjCs6Il
yYbRCsykHODyQT/4FBUhEIKC7PRHUtJX8gp2h5yRsnQM9+Ewu+377Oid10SuKHD8sXvrpcv2Kwvl
/R98gR8Mg3pliYTSwJ38caXjd10Px5RhhOltzZ+Gqh4AMbtfOlPvUiytrK6ERnv8UJ5rcmW4MEUb
0HjT11SliYu3ECE3JtHmv5tO+7sOcaCCtDI6TtlgNUp2AVPyvBT6w3gxOgeGbc/MO039w6OpEcuO
LYo7548eKMcTJjXrHFC7/6IJjkrY2XKrBTbSiDAJQNDbtaHt/mFRj/+aumhs9KlbtShR0wup5W19
hI2rpl5K/HulbTAWfh9GXPdaN1YoASfdcwmu1mOk8r81h9t16fgZeDMxONk7nqv/l4B+U/BR3z2B
JzVTZNpMd/iwNi6Y7LsbQizrQ/Rh1Wim+mhzays9PD5OySXLM7CruaItKwq7qcseko84vwvrF/vI
qNaWacnL6XqEM5z+E7DqpfUMSTJxxc1IKr1TfVr426bA3ABdfiyfMdCbZdwghC08xPg1E/ka7iPX
rQkF05jGwPdIycLZrguBmSVySGMNjG2b/DRiilCMmqtrPYih8oJsSnliWp5NsP9J9MSZY04o651C
zs/Wx8SaoZddCyYkgsbh2HhfSpAO9RO1Rw6wSR62Yt1ZaYUGZN6M5TlpupqIpHYgPOSANc+nEsFt
nQ9Wt4WuseUCXTa2x3lpPUj5338Tlz8Qm7Jg1l9UFMGOyxJrybUQHvu3tmUydF13unFHApNsdjS2
lpQc0OJpm/iOEKIvGzaoiEL2E1pT9zkhMt7+mLHfbhd0A2/MUTrraSwnzQorIZCkS4uMXqWI3CW4
/O+75/a9wP17CG4X343mzrYDfVlzYpkE6eDjj7f2iBgEW9i5jdxe2rOCdpyVBCNPM13kuClfzu0p
dpJLpxe4GZsCSecjL2Ifx70rHSby/WjtZjm3FOPBn+IGnPSlWW6FvPEAqUy5rnzm2v4LT5ieFo9P
WD5YV77Fhc6cgEMFgD4LAB01kY6GZLungx5eKktjG62aW320oya0E2ZStfbP49zLoajJr5PjLV+q
YRvrEjwdF+KY9qKheRoL2ECWPzouh4BF+Nl3ICvlbuOAhloDXOSmwdDIYgSIYajCevsxg9YaSRu/
kN6L8uVeOybye+CT5rBdrhKOJJaJD2Kfeu3aqI4q7wlMOVYleM0thBwYqOoVEErS3cUEOOBPAXmg
SZJJ96/6vpOBI4OY9GP9AWEsrcMtKYgUn0a4OpXZ0K6eq7qUJOx/wz1Gf5i8H4TsGwMetmNN5aNy
EIMWFDH6gCi58kXhZPSB2EMMWk7bAK5piRe/xBIm4SM10K5neoP+mY3N5imvhw1zbnjeelLvDaPb
ETKl5mpPAyaAxhE+IFQBZPW9EQmDb84Ss4MWEkZOsU+8FbyGYXBrfnq+TxDufEQP10fpZe92tcVk
bcHX/Crz3hQ/DUnNcD9yjHOgosvj7fnAMt6rK2BDXFvvG0ldqLnCjccjb1G87UUErsfOlJkYARUD
NNPK0NsR30/v6YhWoY9fT0wflg1Ck5BBJYJNifcjxq+hlTwavsWqGdkF8vWRmpeO9WAAPI6bqpSc
CcpM5h1HqRFAec2tnvsT+MoyuSeMr3Ywv+FMQPWBUBWnoSz4bL3ZVRDSEZpzZd6vy+EwrO64gQyT
5bjH9WgswlvXrLO4VCLguytYz9sgB1tKCCPPxCz1PMlPg0J2CCx+x0Ss1C/TDeIT2hVfo6w5ZPmL
QmXFVDR6J/0GKrmuGqnDMi6+s/kVPSk+HoAcAMzGbOvBAtaYH8n/f43u1iFb3Ll9gCocEGkZ5E6V
0YMOm3TGsgtTLZQ90Cjy9Zqx+stGSLKQ8WvuTdI4vIcItQYYei4wsM7l8JY/Or5i709pQjbNUf9I
SC2HXh1bXyR706eeoGWrO+vLFhOgyr1CIquy+RxQ4juU8e9XZs7tVno7Lodf6vVnG+mE4PBSL9j1
YwstIkyFbktbV5EqYZ1FEdEH5AP+5/oDZwydc4sur9M1sbci3qM8ggv1d8QbhM5oRI1/vcqQiU7n
cL5SU5EvaynofVfuprqAFxPQ+nWrnSiWZF/kchjgDkAV2RbXgvZiVfvwXNTXx+LJgTWAX+WygkKh
MEq0fSsNhTTs55qFgf1bk90tcpRpBN66s0NUgTgcFfW1JttIGoAzkVBnGwBK20Br0bR58A9WYpoz
Hlj5XD9SY4D4vKrRdjA+Bczt/BwU51qa9UPXzP9reNYXZ044n1stwt7uCZOV7WdUXEzTBYPqSH9m
qlHv0SgK4l8bFOgYlwoss4wWPkmd/0KBdczidVo6p2XZnM2Dn6CX0dZhkLQW32hAiBdgcSuEQwy/
7jvXHn1spkx3Y6Ycz5zS3X+Aug6OoUxGP245uZ5O5P5p/bs0yIjUlDLOOBFf44AyPOl7zaEcOtGM
2JaGyxT+e6h8ZuG6MZEkxKkWBR59L8kPkjgC5kxHLHXOiOI8D5TYBTWptvv3Z6plVsIseSc8iFQ5
etC0wjTCazhiSccOBhU25uhF6SEv65qlSMNnTZGI5QeQwQJkH+e6EC7xMaZghQxvZpbnHV7cqfaO
cXZRz5EjYWTZGNnF5yOcVz31SgACRmuFbwvPeLhVhZFBa9u2IcFSnDAn1R3/38gilBi2y0z0NrAA
LqhhX0nnRa8KyvOZWTE3+qIuhfpPU2eCcijkydkth/a/Ts5zHOxeueFqpX6xTeiGWCwyJq+oqCRA
zWptc/NKihYPA3M3MjufmPZ6ctI8CpcLj/ucEJtlu41fLnR9GohRlbW7EDYB8EIZ9Es2zW9hd2Aj
HlVGvj507qdh5qe0WL1TnjqVzsjGdIGp9I9Jc3m1vTcF1LH7+IKOUXR3xPtUD+w2EA+wX/ULGmKb
Zo9KFHdOqfPwxrXn/d3dj2tvHfAAjhpJOCSb1zaWZbYf3+56iuAzOgcKec86uA5uJvnFKUtuxcYO
TZcbb6Gd3UnRxbhRgo+fp/pCE6yNqDjmZ5QJnkQ48tmK3uZsJQEgX/OgiW5WT23V1vcwLqA5LHvr
CfVDSgwvnRpo2jsW7p5R5XTBLoKw2+sgStCz4cvu3X56V5MLRMXWrVKaihs8V1NWugBBrwT7WoZ3
6Vv3JFlLQghYb1my+6eJSvdXxUkhnDU9LW6JahgRAsLTuttenuSBt9PpYbRqCtqhqO6fEjFRHcrS
d4izBhRw3nQrbqjJ/Py4IuyTjPLCOmsY0AgvNN5MC8zAVNKD9w3qFQji0ts5+SKLysQvLa7cngem
+FRfVou6paMPS/W/Z56wokFZ9UZsMkNO//5xrxksevvDXX7nNdEz4Yl8tv34sm1LEyGBTGufIFUO
6td3KNNW4t55t++x84go3TOEAtBoPGWMYXQt/NupUk4fYI3KiqtGM/1yHz7JNEb9IHPew8IkvvrL
wRHJ51DleOF/H8ETwgSyx0VvTsl4SPrkML3ibhTCXuaoe+UvfvIITw1SkAjcd3obQb9/XbdXIk4L
ftWPBVm+r8K4w9i/lXIQMlU19x9qMl7d571cF/dHoHNWqEWIdovuvc8AQe5j19ZOMH17Fo36xCwJ
TUgy2EoxGYj19o8fHOyfplGN3OMOU9PgRQu+Snv/jv8r8yCMU04R6yPpBXkkQU8EmwhEUzQsjbNF
YpOoylj+mL4AXx+4uWhJy5P/ZpraqlHmkXDwEUiW03DEkPCV5zSE4MJJqSbofCUy0Or4Ln55MOJ3
2XCIZ/5Ch3W53mS2QHCVmP+/S2+YehfkcJsXUb2HbYv9ny0aASopdYE7Ox5Aq7MrMtmqlk0iYOgz
TQt4qGJycRK7nXd2oRfM7TkFJINuk9c24hqojUNbDkO16h0zB0c0WbqkH6M7kUhGYeKO4h0xMZqK
NRksdBNap/B+H1QC878OTA10ljBWbi9tKegVe5QqMfFh8Pvvz3YaqbTrTyZqpY5vBoLFfRYqAMD0
BfTjiVBKBI16jltlX54B1vNSmFXlTNBisxRnO4O/MYGkLgrayrztkhoCkEZ+6QR0tEtrU9mwOsM4
3LAP4Jglkxz5fZ6CYh+ub8PAbpQavBklKtdiVVpaBoKEmqU/shZ/WRPpG2vOO1ROgqLqkiaM35+u
ThT1d4FI0yI/8Kfa/baaqePu6aL/mZULuV1ZLw6J5LOdH/FzRJPGz/cuiDLRFMLP+nPitWCFm3Cq
fWET98YiwPRVpXLF/UaXiJSXgvO0elL3hQBjT1rGK1gaj/wyD9CENwI2deBxLMP+R7fz2GeFt5/f
yCkMKG481qjOlDMtxV0B2wuK4hBeCwDKPOr7smj2KEbBewmlfhCvr5eyF8K1gKXDlPg6dz4p+UGL
h93efdArJVFVskpoEA76sZOwykrFlUHuydE/hB31D84M+t4qAw9qA3Gi+vKmcdDYC0k2CS+mLLWH
78dfOQv225VTPDCavTD6ycN5eNnCuA/BdxrEj4R/flCmVa6H/N5MHP52BRGu/OaNOuIpWT6IcGxv
wYyZ4ysak6+A8crzSJftayuC5UWcLuuY7/fVW8L/7/bI2MuztoGjuOoPk3y9JimaGy9pgbvSD6fG
fXhU7tQkYXBJXl5NelM2VSDGbQJjTk4j9mQ4XzAoNO6tXKt827YRxMgH5aIJnFok5OTijf5tF2tN
tpNuvrQfouFH0sJ71j+yiCxm20p2TKZFhnedULidbqG4FrbhG7y9zXVM5UJqhQXhTwRvklNt89Wc
qwz9gCIO9m+pyMUwnDFOstyptnJxVicd2m70FuV3gEKStJc3o0VdUqmBDl6KL4SMMJAzeZUtYqsw
oxGIeTDm4W9+ggaPUogh/oviPXttboWAUS8CRHrstEJZC6CHPFJtqfBgRG3OahUuZpbekECy5lR4
rkSy/LIQb8BB33hmYkG5UYM4Ll1qf8dEi2Dy+YwMbzg0ZCT4ge/RFSPdT7F14BUnxYBHRz1JUET3
cEHCSP+D5wa2GhSh+kPUAflSJHRWsS6JcP0LIoXPPNNK64xzpeO0ikugrN6Ok+v+FJdELxp0lEom
ceHQkGWShG/XYv9lUB/Ne5SDubq3ORB59uFeid3rqQwkicTfSHPihAvEsmr4zM8X0J9uYypc8YJH
dAO6qhjBVqnynizt1e9c2SBw4O+nfIQ9190aoK23W6ptHfG8Ea0tp0WXQOBYG477z5+0j8BP3z4Z
CbQRt/We5s4jGkqyme1f++31OhkmOz+cg22WU3Yx82wbnYAO+DGHIT10NsvFYcXOvD8KAPisdjwK
jZII8TCTAOpEdfaVcu0sxdJ1pbLP+1RmsyUNLk3MM++OF2x4P64PWrv3wr5qP9vvoLSvRYOGvLxR
NGb/xbEd9m0jpLMxzLVEhEY3LAVivxuV7wQ3Z27HMm9d6qUg3WO+msjDThwm5YbuUHd7j2GOuulC
hUMhWvUM954MEU6yFYVA/Y1FMzCRa25v3AOAcdJjvD99qjkJg+qayE7gEBRc/maahBRhJRoq3za3
omJ6sCwkoaYAdbsVeZ/tFCQlnuPj/pF0fNNL2Tc9a+VyWnvgGCZQr4a0FI91IO+VO07ruclPqzdm
Ex1Vl2Jkxl1EEtXg5Fq3yLj/QHSsuZpOsOYbqsdb3TMaEeVTCOl9cL01TSaLVJOFvfTiT+HTtqlw
FDJ3CjaJoGBg+IOxLi0F8UrsY59yary9N0nn7hQhU9dBRv0/zbj3rge0d0FmP1lZyQpcGrxDO0me
3TJUO0QVW7Av0HxPFqcUFpfnH1JEOLQJm9FrF3wqsUWmhAMrqYZITDXi2EBPq0tNF02Suy7GrF0g
rocByfMRrU/GC6hBDw4DyHeT6PUCQiIX7bLxpyfWGC9kGVQ0rppgW7jpdBSywHEZiifAR4PUzP3U
IcaP0SnzdsbTQ5rKhvtokekB73uyfh81VeTJjtQCCYoA8Zy3l4uSJtlS0AJ3Qkhg8ZsKF0tGCWUb
PGNDT4BKokp8eBN5YiU17c3EwsEnabZhQ8Yh/CrQVvElAsbNFiOwOHl4tTZS7X5InCLzwRRBU4TI
+CgwzqNm63qNRG+m6XteV/Fl+PpinSmG6iRAvFBnVtJ3QyvbpTmI32DuuchCahUJ50JLeYQ+zKwx
RMuV8GMqD0iB1+DKuVGziPYQHvCWw26Lv5J2eRhiY7MUIJjvLUB6rSHtFTPD8YKjLWNpV4ElamNI
sxwfdOPUe3bg6vut12sP65G9kw2DafI8PNt36BAgoubCM2X+8TYdZpjr1IgEIwjumphYfosj3UX9
O8ypauKfXyQytk2g9GB2Bq9X3Bc+HJpWIwaVWnF+yWMS2LG85NSq1CchA0f6HNywGKomNfGSbp6j
IT6ELjxG2lzyK+2l7nZde/OKq16ARV4W+bD93XE1RCFX1ztqPqCbO+hEgmO4UKAYPQQnhu0XFmGQ
OqTsSqHTU+SMar4sUkAZHXl9+d+XcmdnKaIv6tJw0L5/pHnXmCJO0aTvtrUNONN2yjGl+HYw1t6c
K2dTlKAymbH4P7nyRi4wtCzSh4WNMIgzZIrmDweZKTvV+iq8XGOplyMegx3E3VXh7eRa+SXt+jJ1
ZHFNgwPTl7zRAMum2d1SO1UYjENOyhmssZy6EApcRF85m/7DK1vcyUn0JXvHHFVkWadL2nrY5NZw
N1ild8nhI5erPzJfAwCre8nrixdlnBtA4q0+ZOgMlMZobSD7yJ+tJyLIDxSHqorv/VKQpxJuQsP+
UaGinLR0cydxB6hCO5YNpuhv+2MnY9t9LWso2VJGxnPspC7ZcPdpX9g1pqQZ+6yUXiNhOeAx5BCL
A9iz6s+MvIMqIzAQJ9L8gYompMAJdPVesDzu4vXnSOvHYo+x+cbWAA9GZaexVYKJ9q3soGyJsTuq
o9BcZDEkoRkpwXi+AEekN6TaMimKCkZ9gbDQ00Ufuf9rN4B9K8hrgQjKNDL2tHm5qv6ZooITT7/o
08G1D24t2FKXDA5RE9rN9tuk4ELRZouytWdCUdtu1RkIvMUArUU96aMp8jtHTMNOwkgKGgKobK06
EdoydJ3y9XLSZzYu56r9Zai8yTOby+RBtYPqWaQFDeCebfXi/0kod2Z9wxF00u/bcU/5/FbXDXyq
cDMAMsIjz3nBbH/OBesZNyUw4Cj7Lr6CimvaH/LCn6WfUwO5mSpf5QredwLKCrVjS7lvrugEh32J
eDgzp/P5zZMTN0a22WExlEM64gnaSjvDhj8teU/rEj297Zy72wHhy/7kNDnku5xycxzFo5QG8z1c
j3qqyQN6lVtcfmY8xXbbhfv3QpmwMKyaBbJTlDal1NPAzYOlUB7YIEk/NUFkI63AP0zpu5NfWM9G
80dOYem3o495f/YIuhA73qT45N8hbMJrwqv2/REp1o0NgsLzb8mMFVi4H0ofBWDsfgo4tyG32fW5
mvi6MvQjuXSUG9WN72OxJUnVhyjK620TKxehYI8lwLGs23WBGhGJ2ZxXygvmQw/ggNkuT1yxxWYk
ncdf5hdieAnjPTPbHrls4L4dFT9mfHMS2G0+H6K22nUlHUdmclO5KpCCgkBCRvFo5ShSJ8Lo+0ro
5l0eox/0AJzKTZxIo9D5XfB2Q4YKSC70KuySL5fvtCG20QZWWHHJpr2WhnDYZvDpVb2zy+9bjvGd
KFVyM8oDYUbEC/SH0US+mrLv+yh6PvozYu99FVEJAjHDPGlG4a9wrhk/1nYRDZKNETp3JfDWTneF
NDuvsGdLzfCD+VJ1BFYc+o3/aTdBUGZ7+JXDPj3OPoq2mInr/mFiJsUAtYzrhrAygxy/cVNxqWTR
I6MczLBugeSQA/fGRHgzLR99F5L0/eZp+7eH6WnQRbJRzVmDNFls1QcPNXuL572B9EvDucpL7tDa
rHB8/KTtXwcmT0EGbQDW22AsKX4NW3TQggQcKkPAyJ+IHt/bC9he+wT39jKKZKLBljLCmPzZUXoW
+x5mXzAy94XyPp1H965CwbbbwOQjpiN2gm64Cb0VcrclILeKeH/w3jnEiUsL58016OLLI7//z0Qe
PsZSq53/A9mKxF+y2dnvdYbQtCgWficvc0jY+ClhsfocoV5bH1ReWcY4EWiyLwbEpmsXs5UZQRn5
7PAEZAP9R7uEwrso0cfkab7W2Yn1L0HZhZfocEbyS5vpPIGhZjfdaBU27b02gUoX1BOgsgU20LJx
IXTnjf/NyBQe9gG/75FMJcdb4cwvD0vIVsQOAz1qkWHjhp0jUr21/kI/FRv4C2+iwWzdspSYSJJ/
W9ZMcE2Rr/+MehjTwQ2nKo/yK8OWU9H+4rI5jKePKajNfv0fTSiku2oxxCufORd+rAFLqF1AzPDM
KFMUzaIc1O0VKZqVNEB4V4+09UM4DEq69lZv2C1oMNXuY7eLO146YTZR0SOmswfaVNgY1fa27hMp
gZ9eAaV788Gc/IEcQZSNVDoojob4Y8H2S5XOEb9azyZrHu9uifUW+HWSy/3g23Jo/7CnXBGYkPkF
rK+A3Aa0dySmfhjShIoG3kltGshyux7wL8QgR4SNGg8tKh9RTQ53lU9RBVBLcaDkmPReZiePAEEb
r5pLd6sXu/vCsNj9wLcyAfWkQqKUVx9oB13zpOiaUIRfNxLFZN9SSMm/OooYl2smmF8a37IDSwBx
5rrNAkjyg6onRXLBQvQCVu8Vc5MZg2nCkayZLMzbcdBreU6YeWI7vTigq7m+OgqxG3pYROI+N2ie
8ztr18eFEW7u0mVdS/7vEP/mNk7vi4qEfgtew/ZM9PYGbYnbH/oeNCwIxiBqDbKCedT5NsdeB37P
owLmAngYFz1PhGRy/+FU1nFhs+LTMq7Ios+rn435oCo1DNuUPZJIEYkSH0j9pvACPRwy1ITy6J+p
4zCa4mk97PZUSov066avVXgKLoVTwM8X9f6vIUT5DdG5eFf510kUSz9U+xNfGhR3eT6ORF0J3+KE
8nJHZbT6HwDLxXt345/Qh4jWxqpBwooj1ZE+93PFmhIciSxXkpaoMMJ49AISsbh2SPDrra4/p9++
jmrtDsUsf30fBpxrSrbglkkW78ejUryhNgZPjSxi3bbFZiZOAgf/jRB6pZfpYyJQBaFc+FXuOId2
0E8B24tRZz5gIgYAzAQ74Zf0pmChrxRW6XDdIZCzNORcYxzm38h6q4eC7DzfL7jrgbFzb4fVMIdk
TVgGAXBEqqg9v7bk49Bom77YgdxhVXfoJ+smQG9uROrqzpxrBGHN8AP558utlvKRhFK/vMTWu1dq
y9DjTb2haOkJ0Rqcx2zfSrB8mpC19yIVgcTWkLJ2rFHSRyqYX3wtEJ7pWujTMo/qzZbmyh5bNIXE
/YoGGYNcbVy5e5JNOHPs1ZDL7eHH6Ck8Gr1C7wSuWdwqSLkBFxvYL5tKBo2vhHMuQTFog1AVNmwL
qTw8tZTBRxgpFG3bRefRPl8PFM/p36eImXhkicNBJRA4T2c/yCbNjsxhrGjAu9Jcp3RTxOuXfp4L
CZiFjXqZf39LO5Ay/eGnYfI4PUtFEkIiPF6wg0rcQNC+Dfe6Ur8VX9cHtk2aqcKMcEaDxrukvDg3
gnlRYs+fvQ5K2KQta/YnQZ+3ERvft/lYO6dC5TuNL+vMOTza8i5QThXTA386WqaW7PPHwXF6h4u9
DtJx6TENRkx5VOX8RCM+eO2eXoERAnhKjnASGL60v+DdyeKbzFdhkc5qw0h+Nb7ja62B+fGp1G7s
XQLeGywuSRCK/hf60zb5zeHcTEihLdoGgSIzxX+dAhlhDSA/k9TFQqG1ZkdcBiedw5G3DN3jvXzD
QLncR+OVJxRnlSvQwRxKRZGC7+hsrbytHhG9M+Ca0PahhFINyHjJVkXHuY2tZal1KO7WdjFUFVrl
Akk/9D5WoX7idtftMesBfTATNo+dxmK2TnQXXqxtBF7L/NQFY1Bb0IsCPFgDUaEH6/6qJY1dh7YD
yu6fXhWetg87DqCu4IOKJY7VM24jm10AH9P92zL32htdmuO9g95cBgmjJZwqAtQ47knzLNPuTNAF
wuycYEsFgOOwin2ztEzAdV1hmt4EKTLffS/kE7wUhjw5QjapnBf+0RbVYFaI16DfYOWa1ss9DgtV
1e/2Yc4BSDjATG+vph5n2lMRV8zxeicadBy43OLW5x9Uqj1qZPRoNZQByhoQ4TW2yC59sbewvFwl
deJchTdaLbRi9iR3vZiT5VFUJO/jh/cwBblwm0iI7m9jT1XPlen159nfW1lpF5tshR3AMfQtU4u9
x0qYRbHp3BCEh68ucvYG2xsgdxG5jfadaHhzSTVgElehFnZk7mT3F3xfyua+CG4wflALaIknyGJs
NSEJTOStbOh47mOVeoIHpUSaJOIrLIxa9z4Y4l/VdSYBQIKKH3Ule1AdM5ZEj2ar2O5xYDs9pD4d
x1VBnfHGgMZVpJJyI5uVt9dKCQdKkumKm7lmBBXcZu+8PtG8bieZw6dlanryZyixDfyb2akXmByW
nohJUGc9O1T6zetaeca2a2WCG3z3eDqQlB1Vjp5w2/Y98bdHS6fqwsg8f6Cr8/o28wzVp4miCKPq
/Jx3oZrGUXHsYmxGXhuDbjQ/hpPwHTisHo51o+AtSrUA1qgQ93Ft/5WwfPhYxq5dU/O3pvia13W4
ay/ooRmzRElE+9bVXAiQRztLVmgtoz1Cv8OW4gh3kPpgpwktcQhpwin/Bwagwq/W9W0dyFjoXXVE
rMghaSJ/eXOBVcMUlFHbtk5/04HTNe0oRAe+Dwp2felJ3itNxVoj/80AAbqj+P4gQ72Ow/YIBpQd
QTVCTeOC0plRXG0God8XN0pq7FgOz5OdpOr0Huq/4CVQQgvWTDr64c91j5tcjzvf7xrPAmmfa3de
byMUmTaoQe8ucaSwY0fyVYuQGCzmsRHaS69AYvjCLAlbixy6r3NtBYxF7Sml4ipBYaWR6KgU2G2y
nOLUQ1OZh0Ol3zbQXLpfIDt8NcElYU4Q0yFgGgAT0nKGMViUcxIswkx6+jmnRkEzE7gJDgJXsK8s
B4cE2S1ToFoO7F5TEowNT0POTNRLtbyT4PLvLu3wUwf86UChjWVs9k7UiFVLK/khrS4hmC9tpsim
EAksyZts1pARgSoNHhIg6ex+KigFPtQ3GbwZbySNdN8MOkT0r3+blMc6Xux3TWLdbIJaN0T1n2XP
YbNO37VbDXHl4HQ2mhCd5gK9rNnz8GTi++3IcSQsbysygkrl1RFae3CglEboj1kjcgvK1CfA7vAS
eL/Gd7lMV6zJxg3RC8wAWDAXdEccMn9pos6wAxtVz/P30xmIezeyb6+DtZf0WIdlZhJFuSoLyROQ
8xV4di6DEcSMDbKCjS3basiBjn9ulwlyBUmq2vDidMSKP3UziMKIG7PiSK+fEQTK/eNvwmE0AkVh
pc7Irny0iEakNAN5jxS5vrOU/w9RMh6rGCNGZUmbXq9Z+9joKbLmQxe56BYdD/Y4Wv43MbmzXRF3
aklmxpn+qhmoljP8+9OwWPtBn45J2RbDTL5dpEQXTX1RZhPdzjQaPoP5blyKf2vUkkZpK/NXGuIT
laXNG8jQTYCz9czshH4OB/hH33+eJu54xyCopAPRpinH0xzDJILi5pzd52CpTwGiKBdjhqGlvDNu
AJQVLqg871RsAH+7rddfmBfApUAkHbW3fmdSb3nuRdeb0ipwODns6j0i+wlMFY8u1m7q9WsbXI6g
xyWchExz6C78aAuYY0tiPNF9zaNWToKpbFkCt4vnwk7Y8b17a4/6JIz5WVcK/rVz4ky+mu/kPAWD
QVCpdzesk95ljP1bEqpraHu7KDfK3dwQQLxwlpp/aWuwrobc29Z9VfBI0NSQVDLwczth4ptdLuGR
x4PAoHoE3lbv3AEis9F/ddAaTbQh987VxDSvHO+qcyYAdhk9GOSyj9F9hiAGoc3RR+6+UK037BKl
ikr6+sK6glZ9JTs8n7rVjQWVaO+0XZcoBTAOlQ0VrrTlp6868s+t5FvgINvzaCM3CwSady0sS29F
dUUg+IER/tscYaFRf0M5Q2zioyWTsl86br2xsPCxSLXafQqqPF+CTNfx9tJdXa8R5KqZehQkUzSQ
D1PPbRu80O8BuMML43O4Oy1vf6Nk/++fai/pNikHsNtt53GWz380ghxCYlWGfrRGy7IJ0zDOHBia
MaGt1wihzj2XUD4mey6nRMmUFaNO8MuzmWEmTW21Y1qsjOCunJHJkaSWtCr9V3IHHypvB0a8y+CS
MWfgKN8GYL58jTE6r6jgMWzu3+AJ1joC3Mfur5ZoHpVUSSi6tMF/xdB+bZuXe3LLJoqwGKd258nC
pcP5VOZ3VocpN05Oq+Ysnc+JxUHVoJc97Xak9/UFSoIp9Jm8NtVGCst/44cukGl9psCaJ0mD8G1e
QCALmrNZA7784GMpsxlZxoKPGuzFmXi1ggIV+qNFuFUe39OXwYtzyAgE6UTOKYkboBHYkRPtsrlq
8gVpE4ZuNX+q4EwriZjvIdLKh9s04Vl0mP6PfZmMQAZH8/0mzPxMbVsVNBrIuM3dq6lUF4aEzdvz
tEMg+cgzQsrgy/VMWbncOvoeduU0NrFjcFRZvSrDWrpr7jBQKfPhuiAuPxqUaIoOGTNtGOn65saq
rAMd5U0m6ePKeW9skGPhcP2xU3XWGkOq1aO+tBpp1SX71WvoVSqQ2cosrfOp+zRCpcRX4XP5A0Mt
kCf7TEHOtxOtQfoDGHdUoBNGPyGVCuAodin5Mb6ku+zOoHAbYrvzPQxqd1atA76H358cRc8uJPjw
VUlS18KXv4Yct2+O/gEj+oqpywjKO4dFBjVrTqyToNP/AXb66szexw27rMj5KbkLJq6+pU2htN3o
cUFoKsor1EOYsL+P8iJXhf31/+1XGsvmjnoOeWyo75XvRP2JsGoXpQGVE/kNtcoml+KWb0OM3w8S
bklhnjAydVHSKhU+0F/laoA6Eqcx1UCIRn8iFS/rkYbhpW8a9AlMPJnbrrOyYx/Z2yyt8btcy9Z9
EJFu30m84HZGv+E/AO/Q78GBS6rHHNDqDfS4hcNtUlm3rQMtehY5n6fYVQSP7awZCcaWRHDfiebv
XB/ut46dWZVX5FuXKit4f8nTk60k9ky/U/fOb9ep3WdbzmYXr4iX00jtvrVrYieC38WKNw/glCF/
eICVeG+1G53Mht53xVHX90KvC5KOiwh8HZ/N9myltJJ9doJbJVT7eCuDldkU21r7Xq9FJSp0QUZt
XAYED0KYKfNoljdhrkzsuDfRZjJ0aMB69BD37NUqG9l1pwS5AWvb4ahPUI8I30+p1T7BhvMcGJzW
CBk93ek+kQSgksCUO6VcdkvsTPYzmQAlCAJoJWFPclSpKatzgb5ldJM4MJymq5Ypcw9LMO1qYi+i
dhvNoCb4ozAV0J7/6DnygloaQFmU2sPpgV9TsXjYQVFB41SlpUEgmeRjBQviRidN3OeC6EkrthFW
kQNNBfrHXaHQTF+CV5ipp2lhyiiAVamj78Ro1/QuB2kbVdQOJIfERR0SHFv1oleo3bzFAv9i4Qun
4vwJtJdXfEeoIrmUa1NrVRMzK3+5r7uuhjF1pRrlYDZG77dIyHTOe6UHa1CRSLRs9GPBe7Lv+Vno
ZrHBUuFA8RRz3ZGrlleX+3sPJJn2MtkUUvrmy5ezK+bMWem0+QXoO3L7RnqPCsmy9Px6Fu7rtrpR
dcIItu6ZxCNw2qFRcR3QbJ9Qw7TdhhJa0dqRHnakvou+Qjr8IFNxjXPI+VMSWW0GtS69BLbbFmT+
YZmPiLvs/SV8n8gGvCQ9PjK1Ql4f2KclwfpQyz9NqzHg8jPP7CvN49XlujVPc6xaoe6Y1EOTMAFf
weDEk+GPmWLEtqtfa0g3jBtudrgKrWwRKpD7hBzbjiW7nyhvMwyKIwxiYS4BnKgEu7V2zEeiKmgt
hLbihEQk2Nw/5OVSBzoZ4PusVRgJq9F3qCBQyacAJrqumHjX36LO6mlPliMPjx9Ye/EfJ4363Yma
n9ha5MwiuKBcFtFP1fWtY+r2ISNPhELVt3egGSC36lFLD1JpLvYbTJN2V7pQ+yALv4mqtlptbrif
QYxzpwe+ilJJfveRpAymEzTYzdttL5FQaz94Nob311soHmdMu0UABmpjDRR+QUKfQaslrYguo7JM
et7q4sQNLi8fWDQcIbVi+xE4ID5U7td4O6UHkPVO1EMhFaPBjEwwKPVlw0k22ezQnjzvECqLH+Ct
780cs1yWLr2zCW7ccS8C9DU7Zjod2X/FhUF0NuqKz7p1Rw2X5E4mq5gbErnOtoi2qBjj8Lv2xpaX
HFY8y8XFS6mKy9cyxpRop5oSIV2NVLGZmbIvCIY1cw/vBzl3+OBq/zpi5xgvS6QXvMigtnXCAi4a
Jk8fZuDcLwRQsjCZMGhanVxiBtyUB6WWsuOcqgxv4ThtNfd8HHWYm4kD4h0QX+2YNXuDAybCEDjP
z6QCpHQgznWFv2qpk84pK5Kdgva9cWRl5No6VXULnq7ys1pEFH4FI0tAj0xfmGhDxReMJnNTeacM
Gk3vitEpyIkxvEXgDtUG11WhNKwJULEUK3EiZGKL5tIaWru17LB4aXyz/mI58BvPqoLVT+/xIed+
IJdts4t8fQ24/apV4ejJm/K7FwdbVe+XmnTnmd2QXzqaVi6BS5Zu5Gjn6iRDz5LX6GBv78FqlHp0
UNKMgfRcYELO+gHBq9jC5E2t5hhk4BUtmVGlm1VVEOfcJYcsfCZ8UL5eD39OoCoF+VhO96ugixIF
MTScEjbsDvcsHwOlVxc0MvAqGHMcFzzNk8wEpyX3Rlmv0PNoy7fwKFBfpcdS7tIw9WlBBNKL0Qkk
lozXqRSJS4WYOP9FAvOJlLoMXLMBg4H5CA5rDZJRcAIJ9jO9nD3BgGyI4ooEr18yooOVDTPEA4wr
1jR5GrRgZCFvVEoLnd66FH2KQSyfJQqB3HwvJVdr2X9tFqx5TkkbhbV1lyQ6wKnwn5PkfD9AwHzk
wJfqzE4rfET1MujljDuWWb358vw7yjnoZXW8/mBBAmYFuKZhBRGcy0q1tRbK6UJRoyNQ9fjsUZPB
tIPDl48TtQ4Tog74Kg74PR4H2E3oZyPoYkteL5j1BvC4nAZ1Ez/iE2yh/ZUAJxxrJ3OZBM8EXRlm
mdSQMdy5Dumg8afQGaH4Cn7oZQLk2zoFJyStijQmCuGa3TqIlShheERoPOdR6Ov1ELfdNytwTt8w
j5xajcDDzEfCAiarbp4uw4IgqAXqNZbrxg4818sYgHr3Qx/spDXHL7oVjMm+JYh31PEaG51VLQUm
csaYt8Qq453Yz65fFSG7DQnwwButa14MiYPBFTh1gAknVYyqxm0ZUpbFBSy+vkmYKnpGE0ZX+JSS
6hl9JV0mcZAYECFbuB46jd7noHS2RTyZirrgNBUcKvTlHBzYHjAppnZVUMi/RksZiZ7zsvYM6F16
Z8dV1/mp0R1evs94vy6DWcyd91effrbIcRu/wHTyag7q0AvpR0nyDMP/LJiSLu0QL/gjFXRL4W1j
SUKr1OiHzsQujns76X9xUK6/J5epkN/sA7O094BgDxG5CqmeQDhBJUXDEB23SzZhc6FhT29EXJli
E8kPhAwLvZVMkJTOYoWqIRbd2tykAatjSNtF8atOrRKFKTomX0VbcrR9a7PRqWfk/cKxQNAWK1/X
Zy/hSS+9Yf8aS6AeB5BQTsIxmbHEdnAT68N6IH2I1A1brAJO6DzIF/rZnAzuB+9WZGB2l4BLyf4R
BMiKo+PHPZM9v7E9e3j2TOP3stqitoAFyOlBUPDlXALJ/GTlttukLURTUZbN3PXjLXlvBEj3gyua
AGpXi8FVTDMyRb7mNBYnpr7PdPn68dDUlURJSy3MUDLK1WjyOBG1IDaAFt4f7cVHdA0vd52VQu1g
QU8EcwIAN/x4I6Ga9xmkIIKJ284MQ35cUHIpjuSQH/Dj88DImrkf+uep6OLJNNV1IHUwlJZFFDqB
v2kwABl2/lql+INGSKvC714ZAjtosFkpbTF2uLIy06LifLEVN5HUvYfMxyjcDO4YERXuB11bmNop
4sB8HXhPOYBpsqUvR+sHenidRB31ooTkPiQFeSL5dFvy5ZZ10pjVp71HPNlRXUcXyjzu0n8+qeHH
xvuj5UBfYTepSlxw6fdLvyPjdg0t9o0TdLB+7fHwCYu6YS1rFlQGuWye311348L4D26xsbVosI0C
HFAz8Yp1n3+HKm6pFLPI7T7lUiXn4IdPYQlVZyQZpmDHu+yeinEq+lJim+C0IXLqbBVyqjYKjexA
UJVY5a4z8aHdlz/TEe9HHwKXUwb7mBztA8DzKIFp5jGz0SjUq4HV0jsgE/K0AT1FaAvKUUnANHen
4CZtbAtwRE6gw4bvNygENQh2PtTxxMIIZU2kSJRPLcbxVM+wQI4cLxUf7L1QaZP6fcDvjuhJFTnx
HnNXUJQpscIyrFvDL8FHV1x6IsWj48doJt/+9at+pEqPVe7HoedkHEu923fRFSuV/SsT6JYCEecO
YFzRHVeyAtowmHMj8/HD0GajhaGgxPT38Afacd8g8TVUv8Svj9prfP1cO/V9rTLlIfxJEvApKxLu
qvJN11TOLB5sd5qGjmcCyz42qz9Kpc+gxX6bAv+NbYFapw0WyOPtAcWgmKMCn/AwEdo7U54sG/BE
5v3BHqhX5O/CydY3Wx4g39AMZkklGE8T9o5+KXG7SUfYEP++yxbx2P8xar3gtMMPhZscBY7aHhxQ
ZC8J6ECD+Rxh+JMfP4xHDcK5SZOxqzvUvMSizMbZxJKRrkXnKqxtPWSjmzp6JB4qUI7h7PAHQxO+
ngKhhTp5TXCbo2uC9nu6dZRYyTrDft44Y4U0UmOYhox5gjWERQ+IsbpWXjZu2MuX6dxxe7MdKJjA
ux89D0n2Iwe6OqhE4ybSpFsJI+zftEFmfM8hbJW3GDaCjMlJG7wniqCXJa0iX9NQhd1emInfevst
udyPSiAkKCDf604wY8Gtdn8UHsrOL59VjC6mHXEAab02hrDTzw6CEWJkWwF7cmk0YGc2/R38Tr/q
2g3bLnH1N4/TOY7+XT/7zVgTLiOoj7Wik3rdiyysfDoDXrXXg3P0HfXaEULkLPliyFH+UFI0DKBZ
SN0bvY77fKN2wqHypUETubTgr/p36ZP4giKMDl4P3jKjqc+IsRWsp5sx8/GigdOZy+E3Fqib3KVA
N8mRWi4Bb7R6hUY3Pum7toe316iBIKVYOBTkOIU9yGxAc4PySZYYC2wk/zqGAKLr7bPMTz/y1VK2
3FNog/B7OLIH5V57GX7wmaPoduJwSOr89bpPxg5LZFTuLupeXKqmerIBmTdo1QefU0mEN681wccI
Qc89UJbYuiailRzpvKaxj2Lk4eUsuqppZZXA4+qCh40YqDJnp42vxC3c2coUjlZyd+k49j999mzd
geFm2ppa3F2A4mQ9V2xTX3ltpM73QcIVHIuF7K/D2WQkVT4ADPtd7QtzkANvXMIPBKHF6bDn93u+
0dceYjxwfvPGsUUjWbw4m9ENZpUGRNzov91jRsRZNEZW3ufm4SQZseeHE8pwzSsYIzzZOoYqPphM
XUGC8UrV8g3mYLu1LsGHs6I8L5DoPa3C83px5kL2Soz8klZhTA90YX3zjuAUR4Rjvxw6GyZbyUxd
AU8lPxdksSDHj9SqA2Su8yBrJqvlGvHw4AKLWFPLpDEXM2D9VRluFpuPw2bwWR+ZsD94laTo5OsG
E4tVAYhwScXD0cDo6L0N4gLXPqjdlETEfRmIbn0HyyNGLP3Yy4n6gDB0o0736F43z4pFoXJ0zWty
uLOHKWuyXD762yiOLlzdetT+OE0e9F/1gZARUUeFcmXoZVZ/AuNVC2cUe5LWr3kkxlHouvtSn/i7
mlSN6ACsiv/kD9DRm1O5y4zLGyYCvjlYNin0flWpxlVHtQ9kJ/ebfx00m6ss2khM0nQaMs493cke
Uo+Sp9Q1QWV0sb0VmYQkrROurlG7Gbp7xTwLEKd6xLqb58/oT2FwKvz+4zTkLF11z0i70rU8McMi
SUw1TNQUmvu0ijUF0+SJ+PBIOLOycnCmjpSssfZjPnucsgYPSpT0ExONTsLL4YCwq9+Me+VBonkP
jA9WRmZ3FzvhiyVcN6V+nXXBe/yDsHGb1kqAByzLEvjM4v76a0RmZMCeXneh/SOHW+BO9BupRgXy
z5AVnMg0qG998TcCi3o52FNrjdseRL19mOyFb89Jl8XN3lDKTDmt2ax+wS3WCvNW4ARkoI486OYS
IqKxyUvVZGHdlrnl9L0ei8UKXi+pS2wmZ4KXDUvkilzjbrpxb9GKiPQ70kZC473otis/Qyb85lbZ
4QGiL39B71GU6T4CxPnW9phCZz1RiN9B2Rt9VhWEnzXRcB0y14KOs8daG+q0t6Dy1GGBtjk2r3Vi
HpJnTo0ZJUDUzrdrXObNsrhoeqvUtiFsBEtZ5pPhpMZnBf44JgYr6GcboYww8NxLlneS4gQCgnp9
tSfqdPgOODgP9nxoYy6aHGKdZ8g9PG2+BXzJEBMFSopYFhbFWe3JpxCfdYV1SBJVajmJ+KcIETg6
Sd9NV4sGFkDP+DkXtkxW9sbm72XVCtaq/cy0W0Kxr6usvxUjhApvK8KK7wRVGpvRJ+kRwNHbJPNb
G0tX+IqSP42xjom4dQo67MdMjCj+Kpt2wxGNHKSkHgIwRJWVnFjkoMNYfN7J/mFpr068lOtQqtN0
yzpQC1RXjRlmSZiLxJyR/53xILXfyIeSWq4fjWVERYgantNiiRvCajAJ9fGpv7XZQ1/xJAg3FV0F
gK7wKgDSXCcH45vnucN7aOIdbnOngYwOfSCczbVk8frttZi5WuIkUMCGXGkgUOFYeBN0IrfMVUpX
qhQISQYpA5FubADFESRVrPHTw/tHjM5QNXS7EuORu0vIFpU8o2f9fUOGbHYCuxJWyfwLmYdxZz83
QbO+sprSXPQwQGA7POEuxQrCmoKa5Zqp8zKiMPAArLDPbp7tsC9vJDp4F2jxk9hurqC0TNQQMgML
IfZxEPZuF67YRtkYRKTKdogDYy/EW6TR0A19l193KfHM4IOb/ewCqI4N2QvgumvrFt/cvZ8QE6xg
kem/lu7B1ZrT7V7RK2TuTkzlREuGoP5i45OxIEK4NUqS0OeRd25R1R0YFEVQafXnObjtA3wmxj6x
LKhMNPVcJyYU1fU9m0SQFzGvIftcIlj+By+Q4vgtf/5ubF38Mmqy0JQEbDdxLJWYnHpfQ2Vw2j4a
ASGn77PLpmu54oayXU6nB2yS8T/RkCsnXFlu5sfaMAiCpu446aOkzczBc08oBTBjL/adTIBDWXmy
WUyILI5mmo3kkiQaAdpvDFBnAgU091eqE9+Ul5AMyJCjw7ksmNoaKLV1cI/b7oEYf9TaPGAI33X4
i+WjwDuFk2ts5054C4SyvZn+Xeb2j2BYfcvkqCJOJwXjVMEMD5Q4z1W9IRbd+VBbBVdFiDzLn0EQ
JbmHZkwQ0E3F2HRcyu2a9+eYc2UWB8YnDNw6gOpKW9jvWjqJ5AmOB8kHZt1hh9KxbEoQm0Q0mhhh
Jphf2wiHoK/ZoF47Xw31m1HgMByDIo2YVNE5jQ1UCM3WPGJt/g3CmBiophmKwZWnP9kRJje+PEu3
y8rqKnPoTxq1Wgnsk+OwyZTLj3YrzA+WshLuUERrwq4/dvh62x/OaGt8XnouiJ7A7ofcT1IGfGV1
pOcXKGHJ8L+bi0qvJMxyg/C3JUyTaykcpY4+aOeCxXi/Lb6QPxrdk0VwGPu+dHl4n4a/ipVSnu58
S2VSjfiKAY/BV6rPsa8OFrQI7gNsyLzSYjUeWWeiqcMws/7KKYQkPO23AQ/gjDbIud8m7N/75Xa5
UwuZIdV3uzRS0BS6BQ6lRMv8DAWDIDB0cUNb6bezsmTP1ZlaXgDwZU18zXJ6kqza1U7wt4KE7EFa
MaNmyNnaHt/jK2s5vNBXjC+NnMvlr4IiSQ7+RCA6lbzjH2/kQVzuuEScE5GXBRH1+x/B9BQobpFA
vhFcn6WPma6E2m9KyCxd2BJxLL7Yy6YTD+UiQRzQQJHe3xuy0SR1lxEl7JMdJp0s1vGhGzt4L6Wr
IN5eAU00K938MO2rRlhkLG1S3ISyfnkES7ckBbHUeTUp9i3mTsinK5kEDmnfvdsoQEXCUZc+VaQV
m63AEit1aInY9cbPicB5ZcRkfp0QZDSsdyaqJWoJMlGtg9Umd1xP5EOqFz/RhOhYdTQMeCLf6/ad
wt3YXfasn1SYHdSej7RGZ8xqiCtbyR0aq6Dii8aEa6paJ5V5c6Bxc2i141L5eX2I0H9AmTJYtVAw
luDYLV8sIoqrhNO7DvQhzSvEUeG9EaVQoR09HqNfD+CLEP/jLx4rqyItlSgFhYHOoxRhZUqwuwRC
im9ZIrybYF8PxIad6pA4gpZw4Wa0kzm5wkyepidCUrIHdItk0+5yfkkwImVpeh++Wrsl2gPUz020
/tKSxY54mGT67c+MqJ2N3lBWu9V8bJEcpGyrOWdKeISl0W7JT1fkZoakzrqxCWuPZ09RBvSSyGE9
+4AS7/5EmlOxqP5gW+lPa+PQLd61nCAYGHTb+e39D5GnnnTRtt4l00MniBfZyn/elDxG7zDoJFgh
Nul0ThohgOSqkyBP94v9ls8/6mr4Ao1nP7c3eyJioxE3eo3J3DSlCfd/d36qz1ATqo6uo3si7uBp
P0uiWD4nplGDYVVmT7KdxRHMsEC9fmG0BkllVeGBcyWQqE71J4O3doJvq7tgtOKz0FPxfeWRBC+h
qNVeXzb1d9nfLzOu1JKZ54lFBaTYM8I0l9IY11JXruUQn1NXuImk2p70iBcyNLhrrn5owAJUX1t2
F+5//jtc/ZjXUrfQiJcilpUwCVHdQeH9EPIRcbMiL8ehUP5QgEihjJKs4BE5jnjSE8zOgxib7bvo
UJ6NBq5Dg3Y4k/KvpQXBkdwAU8oiiZxJhMbO6qgyroRdm7jAmNYat9sikKGhMGCUG1paOx/hcO3n
AsMJDY9AvPHy5n0leGRhK1bdFCLMNMSAcMeNRS5RpdfXRoEcu51RIn404jv+SQo5kaEijIEf/dh8
aZ0nPlmxS3yKXQIvRc6mqVHZI+TWDOSSkcamPr04+K3H4cbWD22xaWIFn96z5CqCxmFJq/YpP8Zh
YN0pEMFuVi9YfDpsP7mbH+6oQ1nJfjwXkt8wp1wOe2RRmF/7vb4NtH135LVxrLZI4hoqDM4rzL17
YafPkSaIko4+P2CtuiMGjuEY19RiXoTRj0iTTXHHKNZgDMSHotZ65ZMa9atGYMwc4JuX3F56UQHb
wQOcPkW7hspSObUztANmhQ4if2OLvIs+Cvp76ynMjW3uX0doZCGlwZev8kxJjjtV2lC6apN7iGWa
YSeVZfwsn0CVTZW8m4GabobLLH6M36oXrG+PwrxdZHnd6pNxkxUm04AsTN31lIJ8GnNSHkXNtsLK
2EXtvkC+vLdR3/g9QbQeEVPjIa3NgdjJwLTzgsxe2kBgLVRsPOOTi8juTqTQqKouORsNChMATBul
gL25hqwoYjsXmOzUN44TxDVHnzK/R3ZNWQ6Zh/rPScBIbUbFwcg5k9TaEEmYI4gPDosUG753Tdt+
ZIp4/DZrgGjL2hNcit7VDLosDSN70rGXAp+HIoA+NJWHABryGByW4Ty/+niW8nDf330VZPawHnB8
mSWWXNiW23I/Do5G/vXmHXQyva4TTyJxfSakH13qHbQzJ9ARMrD0ZM2zvA8rGyv6tdp4acwBnSXU
a42RT21GuWYOieWFmXit+2y0HiihoNc5sU8BVL3rnqNxgxstLKej1Zatc5tLNCp5BadIurL/7EvI
e+9EWQ1KTI+5hnpyI7/WcvnU4zRGFAxbkuEwy3A8+ey+9KgaSl7QoGVTez6EDI3LftXXlA2S1b72
ik5VdyLUfibo7ON8S5qDZ3AE+Z7M77snx7X4n2v6eMmP6WGlDKQibZM8cemajIImZmEZfZOhzr9t
oJFfMhd9Rab63ld+VLfjma0P0QUChf1k33dGbpJ179nHzWnteT2+gNlOT1BXnoY2XMMV7E2XIue+
SIqhQWnKoOlEDvVuOyAwsb6QPYKaDqx2v5+JZipvAUpwsody4tsPZUsjne8l9gVu7wKlyn0b8FOQ
CS8vwVcSixsykcYnCx+GXVph3SNWr1ka/atCZhkHHgiKLAnt6vL1KDRg6KcdjPaVGwVmLj3uNwly
8yxByQvDHYlEGFPxegSDySVTpjiXT+WPsOM4BcmlaLzTxNZQ6QAA8wW75FbErLsaRi0ta9odDWx4
WfOw2NXI+NQ18tSE8f4s30MhaDNxjtfn7ttOSC8MdUo09i4lIDs/bzX3kUd2VYamzPU/4gaf5ZxF
Ua5joceaOReRQgA9hKYYHU3r4vPDF1X50AtKRucSryMQBtk6oC6Fl6Jjztyn3yzqgP0BOhxbpv0o
oSxnkzp2/uUjNI7YFahqjSh227s644xOUbmUGbYPKf9K5Or1W50GDQrlASAEPv82HmwzkqkK1xGF
+AJ94Nbrpq60LfCRHkYZew9SL17hYWxxfVK3RL0DFXmEylzaHXup9SlEdt3qlC6Nqwzdw0bGE18Z
DMCIAErJmq4OqBbrYUxMHVwlVGhSd9vBXoAwGpLE+Fz4KUjgz4C+7ciBjV94nIUrGsnnuuOyLOZ6
b3hSKpTwwnI4O+hyzWtWbcW8ekwASCyws+kclxxY3Vg5hZvne6c19+Y4OdB6ixfEjF431mpbBkwZ
Tq9r7fWxFA2ETjKGbH5p1XJvHcrYVSCHMYd4TdBum/VEr+voEL5YlfOJPF11I34LZliylJ5GQ5sq
i2PQ4lkJxlTKnfjncjcpUq/2ocsPfxQ7Nue5JDQGY+fBneDrPXYS1OEYfBZud64BMeDezNUQC1hp
dj59cBbsoNY6k+5XkUfIKT+KinJDFKYaJ2T/yhAq9IGIV9DFR1fNQOP2PvNQVfma93LljLPQCZDO
t+9gZTkgII9swAhjIhItiiSkZXFJk6UXOtdAfozqL/2v54Qd1HUkBgG4gnBMouxaXagb8pgYxKbZ
3VQegmkQ7P8M0Rngq11BV+i88ptXd+2k/5rZzlZ1qKBl0eufVYNU/No757SZ2w+4lKl2qP//ZvbU
28tkrqOcpK+ySA/8HXdC0ct1jqC6+44m3Om1lZU5ZUAuqG6+DmF+RXWL1B8Oe1m9Y/jf5kQwVj0O
DKFDDe4p2dVHrrApNquRYLNH+5/1kh5VF2KWyuBOqKOzxe2aDEet5EMVRATlTeKL6EInu7GRMVRJ
fgRK5Xg6ad6ZtE/9wuN2l7XLxOXZyARNThDZM+1FRUVKUQbv/Ba2Y51Lolva7/mOO7LyNEoNu7cD
pRiLePjVFVhCVSTjbUK8fGCQK5JZkDmGiAjSSgLxR1mOvbyouPnfdhYFU9cQZpr1VA7lzKdY5A9O
oDCLpuhL7+TKddziCH3I7uwJvqe5IsfBwc5lUamWTfVPvzd9fxCIFGEFGwwuNmC4lDBr1lDF3/C5
ITrmOXBPCulpqJD+etAmT7P3nw+BoXtz3J2ead66Vm2Yz8MA4HviDDNJFgkY5MxOIITPRDjMmttj
GQGVMoCGrRYTVeyJ1I56qh/SX3FZAzlagpnQSRQG4FsWBTuUp/TilP4sZOalwe2yEL8iCkT/6aeb
eCA341NkonPgx5m/vXLGJxFJWivznYP4LoOQ77wErL1mDtGRNGs/cg9ICJcj2W3H7u5NjeqDoYho
1KyqrOHaGD065T63RJVoofCoKHYRkH9dpR0J4Gnl8a/rlYcJDDYdu72VdYV8vi1uRsZQ4pexfRXh
D7lsnvPW/rzNzgACD+1xzk1ItNdeleRTuU9LlPdu1An4d5Lb8ACNu17QrycYBXI1updRj4KeVpsK
yetr2TPk599veE4doGxuWP4vdd3I2jKjVPZkiwtDYDVRU1eqymh/RfnFxosVuoEyfFgB2CCC/nf7
Dr4TmFbi3XDkLFnN3c5opYZvfwh7Cd99sB9WzEgKkNYg+kW71Ca5saz81QdpAksAVndv1KJuaaor
fxbDzUjiDZWdRM1h6tlJBauebbRDVAFfnv6432me+3Z39D8iu2bleeWX52DgF7z+bbL/Cu8qC7mu
63jDwLVNpPyRY5aUyaQCE9KOOVq+IEDdk8Sxu3eu6EoRtglEZvzXpdW4u8rFAL+93ZvzqeZXGK4P
WH0YOEOXFFyGvQ+WCZC5Xk4HhpnVeF1xsC8h50/CmngL2cCGCnRl4l9EAYLfz3v8LbskjowISTac
L0t1fsXQnUfMNspwFQQ0ZULyPcW74sTkPp+RQGCoPAs9Nw96yDNSkcKGU8oN261mfuHAssP+2JMK
R56dpI3HxcAOXFb8abdH4l2wapP0ntUZfXLZgSnaBftyI+434v7vGgVD4suukrYPkrF6nsAfy/PF
yTxF6r++7LdX2vGwFLo4prr1C4iy0PgHlPXG+gpp5M0msxscc9M30pIpEhSNbvPo51+1WGjDkxI2
jt98bPcIhMyrHq6xMcYuvqMnA4NS6iMccqyClkuzkWAzqYToScXXwyK69UfWuFNeKighJ4bkJ13E
LMNoumkNaC5B3IJCFHqOfBUywl4I5yp1/EuRoifPiSzn97BM2bNjC65qBxadnj17ceQ7D1zCsv0w
/fPYmaPSH3RC5I3dqvRRkqMvpsjRz8nuAaPxYgPBuCgxHLsHw31fnhMQ5hoOoZu9CEe9dmo1+c2m
g3an7/yqY1Kns3aiL0ijXHF3l3lfDulQ3G/T5AnKkYuq+1C94HfjTdXwOE9qKnPce7XEh2d5tVxg
qJdQYD5wh8NNpX3Rt7wPmVgQlj2V32OwGDjvgdHYacbY4zHjmXZRLIyNzVBZ2AJ768civWbnKutM
y6OGrzSxdLPDIr9jKRmXDfhR9tWA5GOdvCka7PU+G1lqFX983joRnI6rUrBAlLZFDxnwx05tP060
jybgCN4oV+nemklBZLLT8uyyXc5lavqFbfs7QgbnlJiskHxE8Zrvx+pJNaREWl4qjiuaQa65uJGm
/tStvG6vz7i3MpNsbJJjx6WjM0/IH+u/YmJrMLYkb01xC2PoOJTvQG6H9lZjnVlIrj261UnfncNb
jKtAs6ZbetRmOxQoAFHmqTWONmnWMjoJgjxmbT7fmPgYWVZytZyOrw8SFje9heVE7fYsmAiwhPHf
yHQJUxgXIc//+YN/i5KaH7LfNnualw/3CP1iZpf2pkap+GUTWcIQy3yTiCLYh/YHauuQVymIdFE5
iMxsYX64Yb+yGC22QFNDb5px8rPVk4eLu22lq1CyhiuHDy9pi2x4R+1hTF7ekLqtqREaUd+X3gJ2
mxdZXRzbk8Eezr0kgHaq4uJEDy05D+9Ujd/fEUFd3Ea94kcem9T+1nqV/YmJCHe5xvbrQ3pY4YzE
3CM6vk7jvazhWE9pncok5aRTQ+QRKiXTcYRvdVVg5qZmVJ7YMJ1GdwyHPWEBiBOK3fMMFFdGVv0G
Zi1WxiwTTEdju6G3kwbNXI/izwhy8zpHc20WGfToSlqeTD07qRM7ZVcWIM0xqKTZ/FaJ5hiqZZMQ
+1Y7T51h+4HIibKA3km3/2t/GMzaHaZkg6EKvc4LDO3VCnRSvoEjUhVHjBn5SPA8/IP6CA9D9p2+
+yrONeRQhSKzwLKC7sszeeBbc1awtXSG3pyXlX+BPNYdtlPUV0p9e6KmoAk6kfJReT7uvRnIe01d
TttuwCCDTGqKWHNRIitsnWNJN/PKtTET2bfZeQNFih+v1dMlzg6A4K6OGMWJLkOP7vgghbtppczF
ipwPcmGOjUYsP58Vk8wgzFyvc3aMFljLgQZMskyekqMBYoL/JqlzMh3Bs1PWJ4mUvuUUlvd4c7rv
7sbQ6fX415JAkW10YW7ESHAtqJcxguVLd4LNmSWvMhtJi9/VVz3H4hXt6qPnTFZVyGu0ExYmbTNa
eKiXoOlxVssD00pWB/s0YREP0o7dJwrQYjbZuhkLzzssZrFRHtMET1V1Jvb/a+E3qZZZvLosT6Er
GrObRgte5P/xWTm3erNuzCvVTkPXqMdqBtq0T4NvRC4zV3o0WQdjdYGmJvWoHskMBOxvzqvKbCTi
lA1FAVe6cyMmy1yWvA52HTsJajFhYPFANurCevJFwNx3FbEA7jwm7qY5Ihdg++C+eLV4neI1V1oS
a60oqE6OEideqOeVXkjzpw51Uw6/2IpAGHffB3pQYxmspBWoVSek4V/1FtW5EfN+2ENMYeE6RvVL
mu6uUfYe+S6vx2c2OrmJLsqYkZ/icSm/KJeHway67j68oJ+Ry5VLuShSUJYG58mQSZFPn6AO5bAm
dxCo2xiAMh/1Kr/QZj5TJw/NqjbgyCKOlFQp0KvPPtPza7Y3DIWvZO4CK8KkQvZOOqxU3pRhB+FB
Yt5U74lyONCHoHBVxTKDCEr4H2Lxx5Yhi8o2EuNe8RY5l8GABZZT52RLbKGqkZAXvccSuzzHQQlC
3USxr6GIALl4dtoRJ+npyaMpTAhey50eN26aEtt214bEhE575yi3SGPqVQf5CWyaJ7rfpF1M/Exh
Gzwx463l0LpNNHpVrfj0hb0Z1wQFLcY09wQosQvuadOIPYgQdFjzQ+3GJf/rbOL+rEtlG0nIES9D
ceoB7Enh94J08mI/4z/M0RdIaWAoXAd+9JwOOTuplKXj+40ZvPjHH4tHY75lVAOGU+FJk9RT49ch
JlRgnKsqqOjtq21xR/LnSQqvCuFjQOIOkPxurilfk2sV4XnsIVBaj0NS7p+aJfN6sZTx01GXobpC
8fSjSBrhTlin93dsAWMOZQUZMrC/jOulaC7aLBeL0Dj/vTVh4k0bCRG8MUkewziXR+3EyRQ4onEn
+7j3akhUe8KVPTG3snHcN+8FL0HLqH2dRMRD27B14qqaEV9EXQSESpufvOmqjkX+GqbBsCTYZVrx
AsIjVWBw3/jqGyUa16Vw3//Pu1tUcAP6f0js7bn3luB3JJWKAwgTZqcGRWzhT0qA8HHd21esm2Bo
JJ6JYvT/mCf2HuXBrk+T8xTYjXRLo/z8+CuD/ilz8s++LuEkf4qSpNdVcYKjYdrJy3/m++/ZmYv4
Lb9GoG3LYBj9NkXk88RGl1Lf5Q3D4z03l5AX9W490n0s8yswWgrRv6v+sXn+ZHYBOl2OpocmmDi/
FN5yJCFsdhKnfq+J6Va9Of89D5Piai26B2J1TtSJLNZQVsjYG0Ddasitr1ymCvImY8NGhTdFImvf
CPrXfrfF/RSruQw8lGOjicGx9hkm5HfQeZodXew5McVNPJ1KPtgPzFldnaPNUYdNfkYrgAvPimFl
7/zNQbUaNFaSL6bGxpKQEUlBmJ7oo6/XmKLjl1Vih+cZvnv0SaAsyIidgNTNhfeEsfR6cRp7lcL6
9OtKii8th4tQ0QKcW0T1jxq4GXtJ8LNVhKGuRNAJixgqXCt/FTfqnuEiQ4p3vyAdbo8oatNk5dMa
526ezD5SD9Bo2xWo/kQD9QgpLAkjSuxHbEZgrwKwNmFJMCPx6dIIPkcwmFfxVEp978esUJV8US0A
IwCVXYfBRoyhk3sEEZ2auKcy3kAYr/0m7XgcXH28uhlewL9ic5xaU6uLxRvuKx0THYw9vdSXVQEF
BUwP+qVEUeGzO4NIb9GrZveUGmR3Fj7UpAX/UZuCrsdsX+xqzICdiM2P9tgw7M+AK6J9wUCAf78G
ehXHFLpgGTyKvRe6E9wJCYw6Q4Dpa/Ab7JP+uiAslbOBaQAeWFjS6wR68lkT7jx6lCAJSgADyIqp
kXDmkjICSuHfGbWrIv2AdXGw624QTZJ/oH5slkEoJOa1ToZInFvN3AuqtI7ajcpgzyDyEPyrNige
sr1Sf/tBBOFAwjBzaOzxyA+KDbHOPbpg9O4HezNBM5sTkpQ3Y8+NZlYSVD0Rg2joRybKv4MYRG5V
B22EV4wBQa/ymt0zX/NNPZKx2e1AOFh6k77C1f7TFoHeeVe4ydZqsTCI6u/b1YZMD74NJ2sZjmjZ
UsxkNCX1sRaeYl2Or2qi2UXFyLU5WSZU3x3raiwjDHux79hqjQdBlFTqM3TK2TDgXVfiGqiZr1PN
92wBucGYW0+991klLtjc37K3Z+OsYVLL9f/mcCbXQKGBkKSUo3KoI/G/h7XQJT7Jf+eP2YrZwQPG
ifZbfNqcyGpRX8jGCV/jGsIYoYWl3a2PGiC740JSv+btO2RsmoFbpO4s5ssCebCn4B2DnRnbIrPa
Oume3iDkM45Jv2linR1bl4dDOb/D6MCn/h+6fI4J3K63NajM9CPwHG7+pW4usyprYeSV2V/g3p3z
aaV7aApHWjWQDHrheyIH3ixgwjVDw5rF0TGdgLW/QNhjcpeJQ+XmvhFro0dtlEL5r1wz9AgmzsZd
R2qGX/Qoy+hP4ikOe/Xo5AgKDNYNSyN8g1nQiULMh7ANVdR0N63+xu5U6aiKn3xQ0EBgty5WWhwU
8rwSBrnpQMWhmGCpRIU02n2xErdF2d6mVFYD2vKA6bCErdiPLdcb5bI7zoe1CGc7Eul32jxlUEPI
zepNEB6TOCefgMpm94IRn2IJRGyo4dtLTR1j66cqmEkPYwh08nWC9GdFIwY0fHcOg+nBCOWxXOen
jkOEOPovwgfzwKF1dqAK0Zac+M2UfWf/PjB1GM/1VqHHFGScrYSIZJXaZF6gr59gInUomLODU3LZ
HUgvp7Iyd4DyiIDw4Eb5+qD96bcLKSMpokVT1rxYGk67VC8ashxB9XV2yLjWIBt2eGw7jCtO6sa9
y7Ipb0fTX2AS3sDEajXXnj6NzPpxkS8m86o3QbsVi2jTBXQPwjZ4OmboU0SUMPJQkl9DJECeHSx5
SrrCCdS9Fbrz5nrqMbjQW9i+FqtZwkYuUshDmY3uMypiYIjQYxt2X7p1yr95qpt8FpmIf8MRE9jz
Jud9WBSkdcponN0BjtuoHFx7+c65mOh5dChqs5o3bqhHBTD8GqADhnJgIUXnFSNTk1uBp7Vr1sqa
QQA7iqYEoaegoPvD4ykhzmhZNUkBkId9krV0wCKd5M5RrFY0PHHCoMMWeQ7Ca6AktUjPHInV26af
PhuS2psRg1cQW7id8BpHyb5Eyttxe9kS9yboT9VrtzzVhaHBJV/4hZFYJtJE5pc9EOBvigJCWVNZ
IFNGOIJOk2Pq5lfpZXRbFnfP3cfycGFSX6ka4IjdaMWUTLVmxvt90EJVEPK6xLx1/RQljQS+bITy
KCPN7HH8ikYwzR4kuXb7HkLi2Bs4tQuQLdrjTK+TdtBmSoI6VH2cDpVDzcbWQTFPFbKb5+CUJ4SM
v0rgkOSTPGQxJi/qHs5NVMQ/t4uX3iqVGMbtSZzkl15aE+UDgkqG9A2YpX0Dji6VHcMIT46q3Jx6
GLIlJK89jxB2+nSb18GCn3L82t18Q92RMuMkc7XTCJCo8znZyMLS3EejMqPasy4ySOMi2IAg0Fez
zmb7eSXMfxhbWK/U9LfjCi1POvJ+Nm7HOt79JRNjftTqGF/L0UMp0xsSp75jZhQvwEOZOEOvWG1F
qIi9JrHgq73/tb9/nzUF5pmHxBOFci2+eqc7X86cGJDz3mCnTTK1GYcx+zp2Muxy5FohDd7wBqoc
0QfqktU2WSBjqlh66duFdogvjS6/9t16vOCpeKv04TVG9BlFtavfBzigYMDWuujcCdABlTECLLzT
yUBM8VwYiMba0pcRdSnVRk1V2PkjX8LUTRQH+3vWfu7fk03sQz4SciUQgj6s/IN8CyIdD0KGKcNx
OxTg/CPDOcMWbpMpB3iA5KubaLoZZBHSgaUt5eioav109gQl+8YKUa7U0PjMnZ9jKDlDMtKxrfWo
jfAwzWRD6OZZVuQt6wleH8rycmjtjrAQq0/8uUKjr/mXH/i9+VBai0fgY5seKnYPYVMSUcD6KH6W
gLkjJHo4yahdH3ANNY47v25guCDp1lDgVcn7ZlsAjULrqChkQoEcT21MRYLCKaC56+0+Me8lVhOd
maCgQQ7ZhB1tQuK9W78F6zhf+jQlUJKU9+KkOX6kSL8xe90I3oUm4YAwMdzQXohk8XsRdjZwW6z7
Fd7W4tD1R2PcRXcNhZQYMpONGynSoUwTg1vw15kenBglRndNt6AZV2OPg0mmr3qMeUeZDzR7azqm
P13TkfOcxpbRfg66gPyvIdy99yb0FVrc4R8URBK5DkU3Z9TZZW2pCWJYT3CzYzNYFmAGGNgXcRDb
nH23FtH9XHplHey2aIe8YvbgD/BlLbfxY43fhNsNtu6OJdHEbfOqNsdKi+RwL8cgRmeHtJoD09nr
XBxxTT3EoHHTZ/04anRdh7u20Lqd/qTf7ugpB+IIocQD04g9ORyE+haKOIJ+rArLOPVWLaxehKS5
cINPq8j+9tvpgiCmjPrvGwz9lNjRmMeqiRTmT+qPiFf2xdkuGYkvx4TLUSciOi6MEm9hYbb4MGX/
M15i4YgCjKgWac/WLNE/ys4eD6R0GqvOHQpUFduqmTTvtCUK2b0NGEBMGlkXsdTj6KNfxeYQTQwD
UEaPDN+It92Rrh1KC8Y18QiecJkUZXAiIWg6ORS/4cTDBSHEWt9acg13bRr3zJGCsC4BiHMS0vw6
ElSgq0hiNU+tKnJjHowI3prYNEXyti/TpV9nfJFhwb9tzlu8ttCQp+rpEdlomm7/N111SxGN2bHM
zLm6Dil5KwPtHzme6z6nrSXp3dOPbdoZkKC24TEJLEgA14BPA2Lwtkq6jpElX0DIUUFMvLwjzlRh
UeYfeBSbyuqErspPQHVL71y487+oAwhuz0VJ0L+ozzG6Qq9KwDPld+WrM5a7d8R8cmFrzs8ymMr6
wtKxIzn8f46surJ8/kNtPcNYILh7B8H+uKlx6Fn9Et7CT85+tRG0X8F5MxVgmgVIw2vEynQj9pq5
30jyRfSN5Y+m1zgSMgkHFSxx+VORXUoAKLcuQBtqpU+5NlaPZxjerUWBO47o1AOVuiFH5uzTATg7
Lv03AYQb1Q6LRLtwj8rrychS3wU1CKiOUhplUvt+/qOl+QGuuI6LnjunpwoP7K48cXt+8sJBg7zG
yVDmsiy6D2SsM/MuqbRghAzUqzAIs06CeG7s21HjynEUZJjRlLblDB1ctSOQM2K2uU652AVw6XqZ
wtL9iLyWwY7KJsw2RT3KYinCmhb66TxhfoHNFRuZQJ2+3kJIUL/WvS8MEnp5uWWz4BxvM3JHx0HA
2d6bXwwIwgC7ru1U8n0wJk1T+KCoBd/ttOWgWCznwdIP0nzx9AwnfhWOz0/h/iAba2UbKTdW7H2W
F8xP2vjPhfzEiOipQiflpZ26t4n1VY5aKbcu6NdFxNR7H8gLTAEP/ps1MD0DVREwHU9fQNr0lTAp
W8qdpCXvxo8OkY3c6yPN2/jGZ8xpNHa5sKzG75wzU8574mZaDGOJPjPc5lPHZ2kh+YXgDZJ0+9qc
+PKNmxyuJH2hjrLSTu0Y2PTzBERyR8Cp8WlMhsmT+6M9pR7VFDCIpnUDH+xTsKIkMEmFbtsUV74i
1myLYmLDtGdI55KCxgyp6A8QgWeReVSYmcPSfgR/B2cGY6QjG8KI5t+vuDludwpewxiUbI5haJ3z
XUtR9ysOerFupIDls1x8wJfxgsfU0n1hZXDnw/8S17tGMcRhaoahZgQmjJJIvaMjm138kylyZ5NN
jLZ79gglsIR37xuk93APjy6E6pqR9zoXomxZNn6GIQH7HOE1TtGNljrPgd3M2guXbSrdx+fFaIYP
yH2+QNHBcLXsGwES7XMnMg3Kz7rR5Uv8rzKOlDcXWV8nD3Heic8ykN9Ycm8WrwM+WyyjydovmBM2
24MktX5Sh7bii0EajVwiYO43h+GZeRFTRDcclKD5aWAZnhMsiJhjHz8a6/H9NGkgmXFx56onVSh7
3adZEaH4Bh/q712YX9lBqDOqAWjpD5UpoPYCnbSctDDDmyq9YoST3/tt4hTe9lXdEsKKqPzdZ2k1
5mDTQhkYCHXGCc/QUI3jDTWKG40IyV/0hrAs5HPKuEAAsDg8hAKTD/orMANAUoW9xCxdEj0qiLSl
wIKLfzWjjy1t0oqMtsJH0FnHLUMQGZgKO9qMUjxfclKcelq9AuUn0C2mmGaF7lIOI6tgWS07bCVt
nz0362YDRnyZNuAubAqXP7uX3Pm8Pr3R3xl7M09DXZMz43mZKs098cg2tkQ/f181Kcjvcr1zUk+M
L/kRss14NTYGdAN9L+pwBz5fE4WHlpQI+HAqcoNDb5LlFoQn/GNl8QEy3N2l1lEFmNlU/q6d/PjB
AFIUE2AtDO9wNb0xsEwaNQu7FUszoBWWWuZPnvkjfZdFCAhBcZO0kwYiwf1YPGRRcNMlb9qNesFI
20H/sYTKbnefnsIzafZ+slHZPMHSqx3pr69u+HpkcfvaJFplQD6F9U+C91wD6IhtunFKVXpoEWKf
h0fst98aWWDLXMedWAIjQAoa78Vk7w1Dij32o1y9vGzHQwmNaIq9RdOBQOqSGZnG4bZvADESeO8q
m7ocoGGnPVo94ihPBZat8I7CSuyvMdKqStE8Z9CKHg/Y5L4Wq/0IALATFq1izKjfg+gkuAKntExA
0si0I0p8ILX/7e079ixvKBY0qENSXiWArQhHZfWc85Nuu4mqRI+0YVwvqznfqifddwIbxh7xDLZY
w4/yjN0MPebcJ2SLvmILkGzXIl9yCjzhgz5Q3+DA6l/7pXWea240W1c536OsnAl+1ba6dx0W5jG3
rLR4PYnVWARmfEggcwSOH/pVqO0MrtfhZDd8W62oFUMbeNtDJRvnXmTRaZRKccYb1++iJ4QyEI67
Vhl7lZJb8ryucGZv7upFcZs9uIe7xaWm0wS+QrnMBZH3nKxAvFc9wrgB1fvlOaeIpQZmfEMLjojW
WFMN+eLxW89mJ1lrQMiRqbIGBV26eIpr9CtjWZc5fTTgfJDBjE8Iuk0zwePlWO5oMU6rzGNsVXou
dgsyU4NupPFyovC7zQLfW/IYUWoK3v/Gam169H+lQ3y9m1oTlkBBrakMBw+6UnS18atGLcFPvpBn
E97SXQcUd3wKHyNBCJqHFK3nLFObX0d5PiG6NQ1uACrcq4ETGDlX4w7X+MZqnIKSc3zAPYWwPXy0
KR96YtMeFoq8fgtYWCmrIuIx9j3WcoumHmeAELgKBndX4TeQnb83Ljp3Ya6u9/HDID4kvcJbEwuw
bMDWV4ynaHkhwNekfS1cbRJn5FdAR9TUT8jnREZXJ7WA5q8HYGyjSJHxfPjckTKSjnrPeRF1aHhp
Ir+AjenW+CrFwRgac0MZPFDwc5aEu1EkQKUP3ZKPJuDF9Rimx/9MIdweRheoY+v4Q8o9cxwMRe2E
FdfpKQV0zSO+9Pjm/B3lhk/pazkyO9vX1EnZQvEa3xmo7T6oHOBP9eAzhc0lGRY1YqkiWs+dYoZ7
892Zlvrdt7KdutJwuCB/Wljpw/IyZ2NMhhB5wt5nr9TBg23jylsWgQ8i4ZSXmhUdeM42oS8YTn0c
M/sD0mP3yM+L1BC7qLSqhRycprCNsbqN6mXvGq+rvp5506lpzHP3ujohRnc5ITfa5Bjry9VlwrIN
x/KfJfoG7Uqg+bFykpoDX+0qwtBToz7mdXq0UpXCB8O6zIRVDlNJbov77aqtNAWqyG63FD24ECCw
EpHSb6C5J/MaZgIb3hcV5kqZeNwV7J+747fhzUl4lm8GCP4XnFE/tbyBgbC3isBYrFltuf/fCG2X
Arxhn5HDqOGsVbS3hPfOkYknr4ufRCr5AdTOQFabAQA1LKPEbD2gfZdY+zy8L7LGHO9VgN3bs4of
Rx2yjE+g+aTAzoHSXS1+ssr5bGM6QUB8XgGrZPjnUX6c9aO96SdHanfqSmy1ofHx5Epo/d0VMNpZ
qWBqnrgh92xa/x6MzDX3c7dOK0gEjWEu/FcuWwIG7kzAGlv49USO7fBqE1AfbWdXiCV5GTtEfMhH
tFJ6iDIbn1NujMG1sWjfxusfEmoq3VLP6J285M3wHvwuymjpa2s98WKn85YdHfaUBssXY0ny7Y5F
L24txB1a+0wINrRW9iUsL8r5cbxkfaq3YMhMBneVlZd0TkpKmJMB1n83VSIwDiTT0TiY83D7d8ua
9h0PLOqBNbGiD6kvuRPizmFAJvGMkGsTkuCP6U1EuF/xx3uJhIr5mMN5cqAhK1FreFOQ7T26wA0O
ojh0ZgKPzXRTkc9d8PKDHZzwar/UOVUbNlEdk0cTJh+wkzVgk29NWqsHFtAIa3LmhWP6wVhcd4ML
aeLUGEP/1+RcPp0edeJy7o9F26sQTYTNFQQZE2XWnUpyvilZTg1NZSE0OljiCmabIN7MMv7JiknM
Grp2JeIRp/2+F3tjE4cqDFh1qe1Yv4tlNuM0hkDe0mxMK4Jv5/bFRoHxBSEY+4pS3PQxijziN5um
1yR7n41QUb7YBRl0SrkSrj+DYUUgZr1EI6Z6tN+bJfQcxoCtZC13hXzEg2RBmWPJt5t2soqpl5f5
zyV4IY5ZDj3nKs8aEG8ZWfRZHY/NBKXG5UhrPoBHUz8cT1olVSTSGK1BkeCIbPhFe101o2d2Mpg4
owV42BtjhdAGHtP4Ce9xWsSOvDP/a+h6zTPVzYs8lW7ESmFntd9SRitF9gvovKH8r3KElsfhU52G
fi3+p/mqA7WI4JEED9M3rMny1NYYQAj7j3btVm0NNt5bgfV2DaOAnUKstZGG+t2GBislE7bbMjrG
Ak+LSTGv2+tlXlevJQX6eH+dC0CopnFmpDN+QgyxCgHxcwTPUdwZcQv+2JGZY7lPGy2WcO6Mtyf4
jp/56LwQ4FzeaKGJUJvBtDc7cSKRPHcbr1FUELbQIMiF1WLmY+xb3dNgyAitkVKHwXywZgrA4Zr4
URtuao/esM0cYhvu1JmaAWJtVM8yt8m/XzBWT3yy88myd/SrCRQX9cmeepwqmaQRUlj9teN/XfT0
/iIw0mqghM/bqCw+30LwtK2htO7xOUaiOfM40ZRhhoXh7U5tUS8nCDWObFacMC637wWAN7a1MVWj
iX53t1wbYnTYCmpoE2jNswQu5pK/5Mcssz9e+uhCLJQ63G0Vna4q+guRjhiUsFO7g/3R/gk+znhI
0ZEwl3wn4U0XmviEN4TAJ5Sk1nnGNNCWTRD1FqQPNCmvBdPr6LySJOsdP0qIsO2Ccs910zv7jtrX
Ewv32ux2yM0o4jcsoCOONRVxVb85tF6G42ua2e9IPIsJibG1d07y1IZUfsI+S6IgKiOeZP4i9lvG
R42KSR1RvjuEQadPobzuQH7bd9kjIYmzp1B5fvemv/8RxGQ+mku25k+TAsAcQawm18yJhsFlKhr7
axvICYy76XMv/VEuRf2ElJLQM5xZ5wyzupRYcgbN337zywb8BYxxGABfC0yk9XkN5F1vpDeNuIme
heHMPlE8TmNxtGME/InGbeE0uI/T/kYAI2dQUqIt7ELH8aZVoP3/YPmGXRIGIQTLW36+OkJhGDcj
F0scDm/SdMN9bY8pMgngQGJ+nODEbWC3qb084JWjOczXj9YwyJMooik7k9gfRnOY53yITL/Ycmlt
XMk2Bguz2k0DYvnW/3etq7Z5MrFJB9OPUVUjv+PustR6XYEJ07KUqGu4KGxEvtW/mQWlPEEwSvcl
g2BooGdAGZIXlkupaNGUpXVai9AWqao9hh/CQbN7jd9Iu2Q/QQMHgqLXm1W3sHxQWQy11v2J0s4o
GpNK/JpIC2JFyptwF9SlkE6J05sNoYD/9Yb5ixxFJ23Y4skom/V6ogm71qTPFrvrWkBaS/3m+NpJ
1bzXcYvZxIvcOlDtLkbgVMdjyCGcDG9PFCLDB9Se1kaL+ybzLMNNXsisgXvJ5n0qr5owJ5fbXcaG
iT95MgSdFvk55DJX1l0OnB/QLxgkKmg3oEgOtq2MzAHBUFXwNwnFG6xF+dh2AVQmPl//sWm/VNH9
Qw6Ji5ob92zxKePJxAJtP6HYiBDzpfdfFbtx6tzKg3TCHIZ6/F3kP8TGbhj+tzFvAkZPr/ZlAKa2
xKrkCi2rikqVJVBI132+rma+RXv63M7qOMYY7jfSYUMT4/ERkM3O8IAdUf+VDWkLI5IwglM7fX5X
MYj7rKY2pMs0/5AfQNbNTzgn4uJyYROFCriQ6gifTB6rUXIx/h3rWvrxG/OYajAqyQKeeOd6MFhf
99B35MxYNqlqxlhg8d42kmYRuRzn9e2lPjj/E9iX2PW1vx5tdzEHXwcSKvJXZ/QCgJ19lqPUcNVP
+6VcG8P3lr2LiWN4U80QjTHVhDlQrNP2fdxZKCjEfyNL9FvdqymQnpMXjtfwCXxF95Oou4wQ3L5z
wRYRzz39UdFkWEH1FFfE3BUokf1pkJgpMojBzKAG8giGtq2FyNarTBvFioNgz9xatCxr/TGd5RwR
IiE350rJ+SrpfNZwSBj0HXnTijfZStIgv4Bw68nxcwUsI2TuXdFgqyNU1//UPmBEsi6e2ZgVZ8xa
ApSi/aj2Iv7F+zujNDiszhHb0RkdHJjQDL/6KvQ6g6LLlHUrSysM+IniFAqEaiZfV9yFIcI4qrFk
drHlashAUgnzFJG54JyvwyiG9awSAMm7o94dJMn8SMmd3PqqhUVte8O1CBApykSiQoPO+K81yNGE
QbBYu2mBFqGbmxsagXV8+ujnAwnJeoG23YZ0q3WnQ9eA67GMWHO14xkJ/dizeXNh/FeUCvOFlLc7
wjpCWUWbSDRPgBVp11lfd1vmmwygboxbvrVjV/JLSgWWyFKNB7j+4trJKAlXV5IclBrpOOfxGIMV
Tz+KgFxp5jrUqy9jYlZ143ShSa/2a37YVb9tuEkCSJMpkkXK2Tg/7Kx+OQrxJPkNxBe6PNmwtOiK
AZDjMSQ9zFCGmdIdfqtDvtz1tApCX9gcjsI6MZX9jrTLdBoUxgLi+OrExzh9G3CDP4JG30P/vZ/s
c/XekmhtTmfGD45Ar4t5HA3rHouLhpf/LeDkpn2j1y8AorC+auL7y36xbKvic/QOAI6qBe8PKL7j
JoNBnd0cvHlH4u3NmbqahixtBmw8MD6cVKf6wUIGcKPR8flD8YtSs22OBJCXKZ4un6itkS5EWXq2
V1xLUhEBi70TcEMvkTK8k5n4cyrwhBCBOQozhW+kfKr1B+acN/DNtl0zxtS+0uMjAcpIheDd66hy
Dfcbiyxzk3iiYRwmTlptZTzeHmeTfYnW3dkjMQHv0Ful009B+Xl4qduWsyv+TpMytqkYf4S+CwwU
PiQG3rugvB0QxznqPTkNyWH1kLg2CMpidmEH08MUgnZxjUiwlX2ZTl4a24hFU4EPiYUXDaHq7bez
7I34tozIHWiJDcRaLPTCaVUaz0OuDIzKrfyPnrCy3d7qgsgdErBLvMJtae2afqr4DTTxg0IeDQUD
8JT8Z0KDmyw4yofafuzKAChJJB4L/Z3mdI3cgNtEncP5k8km3STPX2dDb4A3cONWPJFFmeciC1+7
qV+1OsdnrOpEKJfw7SbI0s4LTvp3zuJY2UEaI33AdG8NE3uHAI4knXtwWpqKPQ/mL3Bm1hmWKpHR
oFbYsWnibe/hOVGjhIaNo7uEYQ0vwqOqQbPcalCl1YO4xRGhNd4eZJ5XI9UwRgCoPrFrHBEvecuw
tLVDoQCoLaV3TmreBRMXy5x+eN8XVzYgyw8W9kogwlFiYMw/Pt/jnhO3of8iAQjMB7qu3zaJsTQv
q0tKA+gQLcya/D9yZB4XwCM9TrS/oebfC1WxKZAIb1/84jWYhLo1mZFqSLmgG/PAjxxh9araEAz1
SMjIC7fND1SvcU9XRkF3oefrwQe8+2iZm91O+vWv9KeFyFCMPAQGqf1FNr/l5UppQHjsz7OJbr57
+/wVxexkKR43doVa78RL6R77Ts1/+WRhVBx397zw6e2bUN2XeLNLbhS5at5lhrVCkDJY1M0KFZ7o
1/glUq7pmKyWGt4iP8jiRqX2EnXr6hLZpeHKc3u0kJkUgkx/6AOxXAX40iZ3DkC66esB3xisPzJP
6Z9rnhoV60MIRhdrW56uSM/a7r3kM8Jsxbzhrrq993FT8p+C9oZetOH4ce77JuGr4UXS/Ik/91gh
GMdi0lF9pcl+Gm6YrxO7jzyXsVInALUr+5vPOo9h06tfxrNeAggt9RLUVyn0xr7CjM6XjpefnE++
oGE5c3w/tPWNq3wqaLJUuqIf8PWikJZWRKA9Suv0gJcwjaDEd51fgSzJ8XFA6QiCROC4/nc3yvc/
ZGtoioVembWffLOPpJhpZ11aU3ZANznct3MfGxbul4UUVjiZ8kU5Y9lRH/Xuwtno0/gNzuLpQQ28
Sb8+E0MtIyqgljxrasx+UScv9QQhwMhgTJCzUQw3MnimelWrIqmNZ4YSYR5u40iX0aVPLyiFRP7G
6H/GT0enH6mE9IYHRWwiIMFC0wy6mNIC5MUTkfprHEYgFumF4881kNj2HLCIGrn/VfbsiuDLK2MD
ouPuIPFHWKTAZOd3AmY7o7XNhu2nnpM17NHtBtTf9WnxvOUKJ89VpRlhtR8+TBdjZOxsL46G6b6W
j+BenXP5eYJrMnOL7sX3A/hifFKKg80VacKsFPR2jfYsnKW9PzPt2Z02trwVpszeAlQmBl50Q5L4
V5lBntrVxeTelOwyS1hfWondMfANZmC4wKyRoKJ3lPcsapl3sKoHRr66HO/f9HyrNplfQyNBPcAJ
b2PLNh0mbBfeTrv+q8QnZpsp5+JbH95UBazI+H6S03w4bEE72gGdsjNHyk6n//hid3TEDWb6xLNj
cKx3iyy0geoofufynrR1U0JXRrSzGYGZf2o+cqKn9oufMbR7WGkoBI3gDybBOLczFCWPFG+b1TYP
cgzbkg7cDdx2NDDP15kM1Iv3L6NNMCx1GiHkZPbWAtbOIbNZJNcmn4cZqzsQFpKVT53+LDzxPLZk
i3fmy14ztHohy650/bUVZzr8gzgycYpiwa6yRefXLV3bnLXnk4tDL1+XbEF1wnOLKaDdxDrJxJ5b
MXKmR4nt3XfZ7yDn/7kLgM5AhBCppcOq43jYhf1PMUQ0SClrdtreFAjZ8H2WO4JfDBxyWKa2kpIo
bm4a05Po51G+KJ2bYjYqy53PYLnCNytrdYhb83VQxbgxVN+xZI1/yhRAZf7aQ1/1vCfbgiW9vT7k
adEnKjPRHEUTG9fXl/bR/VEts+ADWEiQQZjNaZQJRpQgZULt0BuI632MEzC8UtTkr/WoSIIvfD6M
0bAacdFT8T3gQE8XvSOGEtI1TtPyUf7/boZf0nDjxaeYi9JsDu+LiRYEZpWwkPa593c14agg4oxC
mBBeEF+vrpQWOgyN1fkny+Oox/Xu4rNwfVfTgO0JAzEDraKx3zH36b70OBL30KCduplGIVUytQhv
FZTW3LBRLignSB0CV2cDACR5DA7lbaUWfptQ3O7Wf4yGy3FMF0iDXF5RWGUwBn7czL0WV+U7Xr1V
NdxOt6z+gucG8C7R5OGXh1lZArF1qeqdkJ5yDX3Ptivu8aM004rjVuZ0PheoayrQJu09ePQetWdN
86nnoQGfPWq5SGeo8TslTROhpf5YfvlTbuq8Evj04RH4HNzfnxv4pvB3QQXg/XPDlMzrT6vLz0XL
RapzvfMIiOFUckAQEg7XFV6zVpxPGcv8Mptj9DDfZCRlvelWBqBleM9U3FP3lwFerXS99A8l+eUT
RoCTPQQu2v8CmpM7lAfoeP31r89oCOuOWwJZBDxJif0mc8VuGF/C5MYXAOECt+uGreG5CoQOOUNP
/9tlIM4J6k6EMLGIp8j2BGGvgqkxLeT54CUkW/p1GDkKR4wvMKkIRG9GOObAOtVQCT0jNmS6fLng
OF3JICH2deObGUjb2uI0HGwmHIyRGl2sduqG2oqClPIgrHBtQz/gkM8i3OZnWaLKsiXQOb+1fra7
3aUP+hADtgFELAqOBpo7FEhjNrTvtYLE9oLO4Co2JPl4Z+TE7xWMgl2j4P9z8qVShLtvs90fD8V4
ZBxMV1PZzp3/7JJT3cHyBztFbySsFys0G192i04/yv6WUmecoDvnBK9lKvYQsCcmNLpWlMSoi1BM
EMiaa9KzO8sRDCRYyqsNhJnLadczJdPGtIiyqUYyMOXNpyOJwXOwqRGbNGSxMJZOytYgP+t0dW3I
b0RUMTskR2WVamLKB+TCk2Lf1ezSYsxGD3kM0E34X+qrlsRQwgTFrctyjaqGpWzW8HTn5UldCIAm
/p0bVdwpa+EPmXmZjW6wflsHDn3x14QwAxuCNEkRXzIsTtaztKIoGasl2Ri6ka5+JSJw/s9mL8f5
m3RzqSsA8FrtDYZq0j7df4GBvyViuQ9gtW2LeoN8blJNCHN1hngMIyaoaY8o9l1VUNPeutuBEy7Q
qCNJ+TgwLRMHardhLbg4vNJVgKx0MDZ+f0sSLNkNdmcOFqcXp8xyO6Zdv0OPwzdtFBhU11+u5GmG
lMT/EfLO6xCd0dXRzz/FwiYoElcww/5Lrotav5+OQP/2mrylUJ80WT4Vu1mwslskIMLk5ttFxmAp
9OjE+doNBJafFW3aNk2OOTfXebQcDH+VYA66PCepGyRCcfNytjjCZnO5+Q7jXpd/AgnmYd3PSmHi
FeHp6FczVEXKmIrd+V9i9A7NDtyers4xfonXV1wzwdhOx9pkfX7dxjOtnfL60KR17s4IfDo+ByBF
qG8eMIrT8MVymfmla/3Xr0k6pgKiEk5SlUzpl4IUjvMDFwJk9qnVRSJpzUx5+DD6hT7KOG51Kn7v
5Qq+EI4HoFBAoDsl3zWNiFJBIQdThxP42xP/Z8fzK0ZeVMKzaVpFI2ZPVSKHtCfaGqZKR+y0HAaf
CiYJ8MUamOUOE52HJ2hEZzOy4gWXMtq5fRihDDOJUTtRUvuHvvJRJmEfuuPNHT+XWfZjfjWigATj
9WMIMOIsZJUIWZ+hgFiU3CHE/0CTjEVOySbgVrj1EFSgcT2Z4cqw7XFej7KgW915VF3y+hx/Mo3P
xSt2ArUX2of5/jaNw40JxjlMnQ4iytCtguEEBWhHqqOOGqbIt0fFnzAaUpcCo9BqDlj9hJPiXjjh
qjXFQKLM9LHZjyQQVN0tpSTugMf6vQeXheWX8nJSVBDGNbaC+jrqaJ0CnWGfclXX7m9NlCqopbLN
5PQuqWmJAzmFweaQup5cNYKwC9B58I1Ls3aF9kmlgObeqJABB5Et6EpiBJuoQZu9g5XlBVuQ/lNI
zc+tUgPGazBL7LG1COJP0XrkXhvz4xvL5FRFaGUBC/1AxIJR0Z4p+zlzi/Ep1VCsW+/HeUxNd8F/
6cDTNB6MACuao20ZiLuNLKMjyJFJQoF+N24tNVhfXL15kmpDUb9gp9hqOx0HZriEM8Hzh+TCrqwE
ePVloBbgaUeC9b1BfC6XA3eKb+0Y8IXrJdt97ZvPEpsAsUZMvDm8awzPrrozIxUXz1Ql6OSoYOYH
CGCZyhuwTJqvbyHB9JDfAByJqrFCPOmz61TbJ8sT/5y4aSOr3BBYfUR38GuG9IQ5DdDXiD45gP9z
q2VO29dNn6/aZ09GTMCc8vbn+XCNLXu5icq3Xq50j58F23FKGoA6W0JK1FsD1aCfmGoWVngv9cP8
dNEFgUCSZ2ngCCHkSvIebJ4J3Q1oPyNj18rp8l2CvwM1JaJSAqBEt8WWUn8CCadBdmb+DxOdLskX
vnKjG4/eIBCXT1Sb9SuUYmd+RdrKGykyOyUDGaNLv+5QUyi7blSvlJbvUvvrKtzAXAuuBxAx1wNn
0ceEc2cUfb1oBLvImlOOiy2ZsIg2EJjMjQ9HV6Lp/0/UBoYJYc74yK2Bmyv4Xe8PKVIfYFyhoL21
HQI3zuF1jruIGLhMSbNRHpBRlf9g3MpXvGz/tiYUb0A9oD8mD9Yqpr8/vOftdvRLBnWit+JD3vv+
7gd05G16ATbUp1DA8deZcRtIkMZVgF4dsf0iTrER94nkSln46IB8x/PS3lO8m4jarjTR+tY0B2/6
NBt6YVklQAYNM16MfupyEVrHGSFl9rAvSQTCLcVKdMEPG0EbX4l6A8XeQu80BCzVfZgtS5MKKwXp
DnuaL9eowFof0trs5MZhK6AugrwTUJ+EqlV7Kz7NcV1Cd2R9Ed5az0RUHZi9SfFtrupIS5xTo8+8
DzlIxxp8pu2Cv1OMLqjlhUmqWbB7Hv023oz8o8nH6TdJdjPyANrcKkGR7V8H004W5J92T0ZzofjL
cQqMVVE5Zzr391U4WizUOxRYsNu1wtRBqdiJvDJ+gUbaj8Kulo5Hi2CcnoNyzZEopXxDHJGZQyyc
Ewxv7BFvJVUgjwzryNuKAnIvlDDxRDjGQPZlrVIZz4521WZOZBGPGGFsXpM32+cuaN1Y5+s4/maw
zqOkd2MWnJGjwe0L9fCAucQ+f5ozx7i2CVuWw0u9M2WBV0FbYqilCaHIHocnm1/+TEl2fa1fJ/mR
n0oGbYmDOgPBRlzedAh+BK2rS5cTp/iPe5vqAZ3VaLaxSrA8bJcvyaqKrwE6cGmB1jT+rBqYy/o2
ReD8L2T89+cAh4jCF6XArLkJbUDaKANUVQ58cotwhQa5fSZpQBypZH8hLcpZeJteKDtogaTnCCRs
QuYX14VCVSYS14y64nlOcaAuVud0EMJsSAGrZZFEjH7KxEhYq8L1ntBLBofSPvwu+BmuTUXKuU4S
AM7NDX3NhPKEvdUQZ1s9IFxo/7sU+yEqJeYjfaQxLgKQgFI+TSVivYizxxj1JtQcFNKdAH67gzIQ
ke+9ipknt9SEkYVktiRen5OvkKqezhyf+9nHkmrCWPKnzrocwFasHGBA6xoG1o9xTp1K6nEbdklc
Jyl/jZ5NlKMEnNmhbfnaeyfnhgdfA9nfO4EeKMc2VATwhsObn+l3dnkaZaghyPkxjRMfWUYpnOQU
LGAEVpUMRXCnc7Qeim0vyavgBugTFZNY6A0P0eB09IGgfO4Qmtj1SlWsgzeKfRblrx6+LeFf60Gu
NzvdkB8cYKX2tx0u4+w6vc6Ws6HLYsofHdBfHTtziuwdNvM6M18T5ErC4/q1zTLEwM4fHbbnqIiE
z0TQ6qyRHQN4wAnW5/PCw3fCef4ql9nSwtRjmJoHaVypeJHmAKQGcpLl3gPp/AqeJKBE6yTZtr8K
2/oNv1sRQP8laNkRsqilnqUxzYi1QJq7+g0V7dAYtubsleu8tsIuhhzenoiyZfMTamMLfQjLp/Yh
id4zYeAWw/k0VQLN9bptkRd3Be0Ffn+z5PHPsoen5bTie/DrZ9MLPAKJJ5w+qRN/tZAtnbK76ZBa
J+yG0WKHJvUqQDv5PylQD3D3qAzOsE+Bwg7Y+02+uKT1yrtZRqShprbtMLufi6y++kHHeI3Apw3w
J2vlnAm485giQrnDVEFoBt4lGQU3TjQGmJfZl6wZvzjo5o0BsSo48dNJJ8nwolpt5JLnDH0GfEwn
jXOmpwsJl/rDCHD/1BCSK9wfJAlkcSGt1EIxnQMudQaZnx4dQxjX7IZvo+m13fzI6bOZGzSoEpfp
tBJleLlZABNE6clmyA7BIKiviSn+qg1MRlK5V7WhhsqcCOkrDQ8gh08gFnYAWVrHNziIUIjaFSvf
17CAImNDY4ss8WRRYp6TA2834ToWWmJnM3lZRgQBKGuV1ARhwq6+2511ozFZRm6IVjhDOyPhWulj
e9aA2q7ikM6pilRRBgqtB+7BjZ2uz1AbjTD8O0LSIuTfZaSQLX55bDR1CsilzY/yTMeUluwoPXnN
gxMkd/9+l+fNSC8ncQbGaHLdd0L14qpsNdJWTuzMC8LYVEcYkdGw0zfMXTygf5PF0LmmRB8OQ5O5
0fOqQhATBh7YedjXwqYOLoq2eFeWo1nXvSpyMv/Pef0QST07aGLEuz6qVacYLQcwwHfN5S3ow80y
kT5TnJcWEUAq8azHDgiE3VjKH1j+USqXTwD9YZQgvBdu+hGE1zWj6XoGMV4c9Ff+EvGP7HFaKjGO
NQXaS2NUJBUWPpkPSJXvkU28KEfhW2qVCF4jnKb0xvR/0y95y6wSoh0JmgASqRlqGAWz2G3uICpm
xnwfYfhaU2nBrCEwYP91yKeDYbyc/Z7iPqlCAMFWomceL9dHtk1OZzLYEVznrdZ/tdnuuFq73Yff
pFvExm/xDPGjlZYfecbBwc2O8NJtCUAj+IY3Hk6Ooo/FRkexPeYzKcuU5bJtwsMEeHCI4AjJVsU4
LsD8APiiJk8lbax2MvF9dvCwpP3guCeBCnwhEWuTtEHZ/Ci2fc6Yj/bDh8S0NgfAfiBKwZHgv7MA
Wwg279YBAJ2eRhM+B5SZdstvMmgRp9YDDCas6apN6PhpPlVZuox+QlbkH4xVjTMUFXFejOKBtpJe
RdNQLoLsfUiDZYXt/5yjkS0wpvvkcdx9vO2NMJP7CYAyRcKiz220X8THydaUyIss/OKLrFiEcKuW
rqG50XhfZHtCteDGWpWWVshd4XggqsK5xGGfh5U1epwibpqrupkKeQ2AFa1Sj0u+gGqGbSEvwBvs
OeupJArpRzM/3SdqoVMFvwHIY1neY0phzHb68yPglMsCAygMi3gqMzQx1lQ5471GjoZAQFTX+oWW
8QtfgZHrdDnD5k2AUif+w9IwgRX+4U0YxBBsqNqvQ5HC47HrihJTHPllrCIO/+mPvGlMxdOseq67
qCwZxLqLa0Y0MikMBMnPCnpr38zIPYUbbBJmstKJJczQXrfTGSjHbpxzgjUjRe++ZprsM1z9621K
OBx048z5tUL9QnCeRYe0cnqCB66zAKI4qAoAfp2C+mjK3xcQexW7xQOgBKwloxToMvJKkx0JGkHw
mjK01r1Fgeava2lslkHEWnHlknWqMXu7a0kRu/MZnGWpubJFiv63NWV3A0un1yc0TmzKc9BJo635
0kBGKahnvvuJnblBXjoyjt+djRar2naiLnKh428//jY+7bcb9T4A/853TGn2BtMXCLoT4FpKvMky
ThyWUCGRmMlOrwqKpT08VN78zNHXTE+KUvpvFdZcs1mgygjPkHfaE3TJUzIFeEsTnZ9hhA7Zi4Rw
yU4amPCWueIf50OCh2cv/8hPzMsWaXJMLr2g9ewyPQzILsYJLns8ypWaeuSYkjUVUqCkZ7o4/JKh
gD4N5CNzgbiMw/IsRYtDDbZPJIHSLqiUE6jPvU30q9TMxtHhQ3xOsE5IKwBIgW77cKqgSBpR73ol
qvaQTIwddTkMKKSaytYQPyD7tNimDbjl45phNOe84vvt76o/GIfBPqUvs3EXjQWo8lIy7+GXtdqr
Mc222WQXQk87Vf36WQ2DOMNNOX3ng9cOOzbi/aNbg1mHqwwcxieWQ07FbVuG/LuXKcXJhDbBVwwh
JkqBzx0/GKbJKoXauJ7IxLPObd7fuFrKvHKlb02NaEkSyaNF5dgytLMrlz54txvyizvIwf0829TU
mszo9U/WPkOViffcGYj09zLdg2nbs4kh7Dpg19rA7nRJTTeSmHjHhYJFto4Rt0yttOCfC03i7+ya
NqwK/cqKn7JuTCyUkYIgOU4PGxJ/X+kef6DmiPO/vNzfj3aduOBStvQZPSBzDfbaiLcSOfsz6xxc
BnrzsEfy+uVY2ScVOB8w3VyyuLru3hW0mWDRecheUVHX3x0XtcHOaZwn6qEgogNIHrvWnnh5u9zT
vEc1muwtLTUhrOVs7KC08IYFMWg8VYI8lDaXSTqj+BI70D2F6I5FeaI7mh3PIuyTQluQnjJyj3WD
rE/ywDOp85oOBTAYx2xMKxvRwQtEFhE6f/553ZUMk2KHpF7++hkRVnQcXu2todlmEyfYzZfJ6pAj
ugUx2bpF/1poBjMkoNj2pVv+HJuR4aZv4AMZIt0Bpe11jLM2arA2zLwm6iRwz5ftL4jUbVhtTfC4
IvS9xlB4e4zjL31TtfRI9jst+gQb089imf3ttnhSAts8S7LhWguCI9e7Khms81mMI6mOLMatGL3M
oU3WoHDkeDFXNHEwwt378WQ4VgiBxQrxPNwiGGXSUzghRmjxTxf1+X+kloBtPIDnScsIhXaIl3pO
AdQTx6Vxg9VCGVedf8YPjGJOrSmLoCOqCgYKTBIsVZiVzG949F5hTfinKhkhog0ZZGaODH+NrCFf
xnO7cJxlNptGmaoPzIOFbVTTXEUY+gJBXXr7vVlyoe62TN0kA4tcCfvk+TzWGCvr+ZsgGK0J0WC3
P4GGPpVycuzAnOdsaDQfxdG/PvTcGWMqjExiOmqIIMbwSc5TFn9HC916H9qb84cYuvhTg+Gv180+
mX/VTNrpN6/oeEfCthhpkh9K44Plyu//gmjrFE/yRjBO3urv4sQPT/YMzxe4t95zKMqaBVBgXMKp
7u2RuGZPprNitknH+bBvbKAVWk8tICZ0fPR5yCTTGijZP9TCyzUt+LrOpOeVfTOa6wsFWklhEzK5
C357BqyVN9sY7lq8G+ouOjUALG5bMErFW5BmhG6QqtHcMMuHxqPrIcCNt8p/s4jEzJOek6jNjz5V
UYTNwMMFCCnBYaGpaQ7AhEyh2uX6sExyf78NRY6Y0o7DqXd1EfpS6wq0PPTakKlKxQzVdcWIg7cc
bek8grqqW1DqpGw8DAXcxfxvYr7embUxirWf07Iotvg5K4cQyK3NqxRYVyNDl4fnHaveggUSbe8I
X35WwMJvkmHmoXvRim9U0IZ8aSxqxP64ZVGJQHUKtIrc/V7vq9wZXMGuRb6rTGTXssd4v8ARVFgt
ycabahfoW7gW4Ng/K699mkfaOijehfnHKVnYw8TBDxwPTP63RxSWnphHn5AuThKAnoICvMowp3et
zeuYgC9JiSIBQV4oDemNEZPUo0e5rIXq9PbxTRN9uc2JsuQA3tnjPnyu9zm9SWz1lggBeECd3H0N
K8KmQP8KE9+7qwZOrRiTkZAdoQQxBucPo8Zfm/Xu/tM7xiuLo+IKesnvPNN6h2vuQxDVn0/Sxo3J
4r+Id9Yz5LgfKVjiJgRWaViGwn0rYe/cdLE4U7n3JYtlYHVt7CCxHHf4Bn5SDKsvjD7Jvne4AgSj
X1nSjRw7/Vd4Gp7I709kHay4ZxL2myfDkF/7Rns/tRcNhdg9jeD4GpkZtuyphKuakM6ngxpZj2Co
f4bkv3GGl/r+r5+FnLRueRgCWstX9trRFgR3aw375Ft1sGCINs69ifYUL9ZPkbGAGyYRTBYeMa4F
gppB3IYSg0KKRNREZca0k2BOhcLZho3ZcY5/DvuRh1PRoXBuguuVnLgcTNWaNoL8HBkMHE/RPI6h
QqsoWu0huPGY6BhP2qUAez00N0C25j3DatGRvj9z2ypbtq5r1kB1nUfpNaTzGwEMTDOJfH0RTNpn
0FlZHo/8HJcExATHADgst3B2UoVfqVwjKb076G9Sb/kIkA7i5EMMh/cqREHEbxud3Ns25w50zhOh
Gup/EBSI4mu5h/v5wIkn+9m03GwSuOME/SIhhWZTUq2RtI2V7g9f7vB5rCa9+ww+PZ1Rymva5AXc
dQByb0QZYnlBC7gXR5EriwaLQBTMk8Yvr3nnzI8UmnPH33/EB4SYm3/ulmPUCdKU6GskLteJkAaT
zqkXj/ie59ERMJdVrsibzH4Mp8yJjcmCsPIxKOkh6MWzzybFmjRBJHSoTTQgIqkJ9R3FAltLXndK
S1XlZ1GNZCcLeBR7Hmhb6yhCLEZvN/accMP2CeEUVNC+aWCIFAdWuDQKC6q+Hq4XU/03o8Iiri9T
SrY18K4kRFEHLqDbPEKAAcpKIwoevxg1ZLs1NYq3fBzuxbJaI0HUJtyeiVhiRHa+1QXlym7FETjE
Zb4p4mFfr6SD3EKY9dSitosOlq7SsCiI7K2OqbvSY29c2bUWrafl47ZhMnEt/mpujtFyht78DS6U
UeqcrnyEtM7THipfxoee57jV/bebfLsuz4EOly0nu3++tIkYTx1Jh87ym+S5OhMVI+onSDGhIocM
Nj1ZgSGRxsn4F7YHJqZdwET6GsZ/oDoOwfFhU6ZGUjqDQgtNkQR9KTXvJPoFZ9hjY8iFV9oj/W6x
/8d+cz0O97QBIBBNM0Jj4yphnRXeBqoY+9sxvi0oEUPY0s9yEpV0esinx7i851MkwktPMZzjOxUB
vPTepOVp9elcudSv2Gw/upmJv8H/rifqG2hLSs9wG9cTU+cCo5ZhofL2yLttpmFPXwEoYA7cED9H
dWofay57ks8jGPkDZ7FUDERG9fgocdd2XXfPVIj5oFi3aGKTJvCAI2YJbskAjpSOdbTYmfhxqYYe
hYR04YK7+Mq4iTZddAw98qy1iUDOh2ci/QMn2v45RX1PQ5x2lyjhbOiH5xIHEFm3K5PUt8HsE2Hy
d/a3GdxLnLiq/RdPekpPUhrjmmGxpsuN1iV11VWqCfh3EaSUlXfVmZdPdO/HqhPLS9vXE7rNQsjG
NJ2HiNgamC9sn8xJpewl1zvcAs6DD9sUmHn/m24lPwClPn4Cn4h7v0H6Q5mrTq0A55NrHJK1zeYE
fEC7vLD414zBl1nfODygvdUSYYgRdNBdfgM29J1wECobtVKSYK/T5Au7jrL/c7Na1OPEEn6kXJ7/
5zJlxFk71X1c4YSEU+f2dg+lOwwxEy0UllkGX/L6aLGuBGe8DQzV0srvhCPXWTrHsWrMP1Rirh/T
1EiE+uHCRaccSXn65hjzI4HKi5/VGyN4gK03sPtsQBxvGAFX4eCbb/clS4uyjCGa63ksoVlwNQYY
BWynd5bl0yl0plqiYeghu/vbLqPSULyoQ1GeyFUaKEOqAAgCORZZ4FCORDhhkSF53XfVqxpK7myy
zXJyLNQ/ua0XHeQJ9l6cysbiMxBFm9TXWDGx+R1Ri6g1rVqK5A776uF957H+1KKQezBHN8YeL9FK
QNN7BLZH1DCoguOwU24bO9mMuaqWC1aQhyzVa2nKYduZR/ZurQsqWV1ytyyL5RJm4/BzXizxovw8
mGK3N/ib7cneH5X8wtIHBBFq0hcsSYd5kgVkWSzrS7VGL97C3/GC0NdjF0nK0/qTIPO2cP5I34+S
5GaLxWO9uM9lT9JSnaldy1d6u5DssVvSybyX5XzZzVRSjPB/Si1Gh/usd65BKViCZBy9+HlLcbKB
MrrBE7WcYj80Pq8WSsSaeRDeZE0pyCQUqsU4hF2yh70z3DXehzGXBHnD4ti5BCpCqD59KxnxUZ5V
PCVeVrNYhQuA8jm/0+3GyOmHsKoUWFbqks1j9/fq38JcLPgvTJBMNqeejNuyyReAk4bYB04KM4hl
wYesF9qBuJvWqBNtH/LQng0GJgwDY8a+kFl2eaSlTgzAWohN7h6jxwazUBPJ1lwVIe2vmx+3rFso
Q1fzz3ANjTWIr0+KAqOW2fN7oANEI25W9z9g+n1LI23Ze/F6h1VoS8SsU0DF6nKxsexkY6EEtJH8
T1LXu8Vkf9qe92icmyoQrw/BM0doaU8qngr2rLjUSxe1sJX4et7u3E62xi6i4LfNgRm4eX2mIQb2
8Z22fc3FLy4StNfnIxeNvWg5M4OLdOiYYSPXGfYD+0kocLr6WPGEWyUIhsnazk/FWVfAOmtk8iXG
nW3UxYeUbdiMO+NiIfW4gMI4Lf898KdIcASu/4kCuQGwkgW8bKsGrRGeuqI7sC9aB9SdDBkvtxjl
oaZMdaosXB4sebME9PYQM/TxQH6RdFMsLmfxCFGkXCg4mewfZN8WR8C1SM/v9lEorx5XOmFhPTTg
WiLa6a8s5n+uKECHRmMtRpQuAAFL+hlJzBO/3C8vCuIEGfh6ZW1ya5D9Q/iCjtfJGVwlc4HRYQnw
RUl12y8+0A3R0AzAqM5tynQMcMHmEyBb02VyK99OD94HkrKhHpFkrmXStvEKpOuLTZxr82qh1gIM
cTsN6f1SixyCQXBBgb8Nwh7hB7A3dk1oVrOtzQqsseqx2zklo42yq4WVnmGwoluHkmPeuomlArZn
vWG1sFjwAb+L37sxjNpRcmffppojh2lh9WUGkZOuq+f5RRWtr6sYC+vKuGOM83UYxJrz3+fryGDk
r1tLHf7s0i7F/u38kgtu8neHdy0vQjx7HkUhFc5XqY8uNI/N1nj/esgmYHZQ3h4x/KoIsZXZZPxP
AG4VZJrmAXgJRSwufhMAgHJjIziZQHAmlq4tAfudSr6pjqnNfcedJtMGR8CySuKNVNaQegQQzsA/
dOZv5shBqBCf1QqrFbydDyPoE4XT4vsAlqkHdDhIqx6buI/itLaM28DXE7N3EhICG7r0dXLUx7vM
euovFgiJrFcl+FAXLlW9GkWbHTydBN5cfb+YJDugkOARwqnenDptUJkkInZLRo4lUyjkh4KCs1GL
r1Q4L9bLH+mo+AGp7b1gkXMJt0luvY6N0r6zYrfGvdWeQIGUX3hDvjUSAQJOSqZHVAPefGJEasN8
OXAmrQbse5nhgLa3u4wlPOfpiOcUIuxmhR/hb0P4oalsUJKT1weHZd4/TSkfA71+je0V3SuuXE6C
cMpcx5TnvlycSdvRdVy/CYfhFBQR/L/6sBGrQ8fPD/3AoA6Zq6LUC4oA6wI8A64uENnc3qhFjs9c
oYGFwC7HE0tjmX3sQ9bWnvTdi9kR2u2VtE6NSU6UqWpCzT0Jw1CDAieuXPYXOq8OGFq4HQc8yCrZ
3UbW6vqFP98ceg7i98CQ7MdUSAhiS1/3xJ6YVll5Es3j5gBPvz5zlayXFdLj5LDWJxhL0/dW3pTp
1KytIAXfToqgoeKPv+rg36On7/Oc7DeqPw+z0EYOeblwFGZknxyMnxu9/9R2+baXSRxM37w7mkPR
Sr83bLkpFFsQ/umx47xQUf7nMII7w8VMmh8ZKi8qxPP1Kh4Oh51pJvMMdLhbQhDZPkJHFkTdm6xR
SW8qR7cC0QSk3+1c60l8NMmzXkR7ua2pmtt7ZfKo11oQPPtcXP36GE3EIC+ULhBIpvI+EUtt1wtg
JS3D7agJMAmV2c20jfOrlfqV7wwFPXKwrBOh5cvAO+EQUxxwHG5AbzWevZ1dbsqROsdxlKb5+Oli
mUzTrowVBLWYvaECOYTl2WqjhSYtUI352c64+1wIPW/x/vt7VkwOZio+CJnS1i02KhJGqdF6Oyrg
t12ZeaJ3PdgzlmwSH0twIqVkb9kH2ZlN2M+5aPRn1LLMuAq1Mbjwhsxf2WhSC8QUl1JHLntM7+Qt
npPbFbb/Li9e7FjoPMXGmaJsOhc5x4eIVRlf/xDYry/ix8DRKPZmOpRBs0YK+Gwn2TKrJpZALmot
YtOlA0j/heeGBdWcs1VuR6BHgs9zE2Wn+enIDjxrO/URThU5YPt2S0x8qws2ryc7y5UW3UGO1Q6V
BOVDFiGWsB/FIUbmNFbsORZrTkxJ0t9pPIUhQFRNa80wsCObzCHmrgmmoxyQlVN4/vsJ51+rc5Q8
/rL4S7n3d4/eDVh4iwlpoJqnF5C4luzDzFofzgKRH1NpZ5PilA1kEQNiBTZlOMHk/bSG3oXe0/i/
VBfANxuUBDFwubBs8qaRlbQ1WsUwJYfONfexsXQmblGGR7L+cDMWew7BqeHs2fVPd0tGQZgsnrRe
HkdBjLzQGDsVFrN8DnO/5CFwDw8QOg6KqdjVcnx65pjc/tK1lnPqPBDvn27W+o/dWsvL4oIa6X6P
TnnFng7ct+Ca/8CXpnr4W28oHOfFysqTEeF9aqF32R8lJO9Zs3TF29lrqcAyqvWg1SP6fZGmO6qQ
aGjmMeC4/97toZxQ+9ZrhXuZ/UcnQk6Ctk656QJzH4nvj6MkEQ9abugyAfBuxXEyxTvLdYFJcKZd
r/ZeH3cucCXOXcvF2t2yUP0Xr3GI/4Z8qjieXD5Wt7X2G6kPN7F2h95uGQ7MWZtpHCI/HGK3tpjK
YxJBedoocSMaJ2NIub8HJ/ALJcG1T52xHgDjjxFFUTMWl4I+C49zhZCNAGV4ylGxlqJbiAau7M8L
vqFTRVQonRKd2pGUaztiOYTVEGnSa6oGaDt67B74Nsf3qrtl3mUN0C0dTEAvtSvSCt9ulgmULfcr
ohI96feTaFXtEJJGv38e6aaQX2eewKS63i/8zKeBzRVyfpnXB/FNUkEq3J8IvxUnzfNgWmHXVdMP
eBIPRf+C2STC2r3aQvTt7e3gzfW/qvKaY9dfIh/hxwadWO+R8Y4O97JgK4yXzUg/RPLmRPrHDYdt
9p5GKYI97eAgRUvE67a+8JSYGGxS82tXvauE5p9AEUN1DJx16UOJAMol3/SK+cGeElbteAwF2rcw
PGLhB07bVZV3ipSPHo8NNqHhqnIq0SIoh1PWPvI9LBwKcyJUKzL8BO7advAk44n2tCPGbGIy7zB1
FPuRdramTN3jGlLQuoFhxnWP4ygpP54ZGO776PyrHreLOB/nqhxGIIbiHYxKJuNQ9hryghRVopMg
cpnezgMhAfmSiyoD5ccCE5bXs6wPMn6SFprISbt9bOlZU2HVFxouE6WzFbvwrFhGhwJmo4M7TMJ6
EJKp0YiJVHGBjyeRebQ63yOM8W85EsElpvgW7Cq+vwQjKZI2Jzj+EtgBM9QSwaFHT/CoPm2gxlKy
qOh/PAnkYzotQQ126ScJuwPqDjyqer7kAYYY4OPoXLH7p1ig1UqULKCgjfUpoDx7sw6BzvQsQQqD
9APINzMgRj0mdRrWwQXM5YNhVAhwoiHNvIqQ7pyg/TIIY6eORB3A+Gp0fjwJ3uXOVQh3bq8aNNON
aoAgVBvEZ8Ji9DN336LySxwGhnJK1NA8+/NKneDiKhG45wr79lF0jMThR2glvUPSwbLgOFbptiIe
3MpoJDjXOK8Poxzwzig7U91KFR2s6LvQPtAX5SBpAhU0VEG6rjzcuC56kl5Nnc0BdtklBtK/xqsh
4GzecJh4u1iYcp/HwOlHunJDDRn2Pdivj4H8SYSidcxoiRn4td4Rc1DV4BeI2Vse41PT4hRJYUzi
3bwBnnRyxuTkRaJc1/pPnYpFFh/3LimXu0QgUbODhHbvWJUx0cIbQO6fLAAy+1/NTFX+BDJnAxAz
0Kf5ZZ1GC+lPfOdyBEemophjQTgPExm9mKRkoZJ7Ogd0FUFB8ZBYuPxi6RqPWoDrlGgmDfdmwGTX
FCvG2y2d5BNhgUPMtN/YQsmvmOJZ19xokMhnNoKldP1XvZLk7zDLsQ6BCc13N2aYXuZcN0kfqh8b
XWRoE+rzO3psI1Bz68Y1QFuOdECiHX+xPr+qPr40nrtu8utXkhMJWCcjJ+7z/Y1lsN7XX5fIwovf
IMzDKXgcJ0Zh9swNXaUhOPMogdxWvAAvzBesI0Phj/5aHJzNehV55ULmRTwbBveCz/bGXGCHdQm8
732CGlZI6SqCbExdPCxmc8oy/kXL2gN0DeBPQtC269EJCR1dhieXH7xc9NPLut4p8L3TB8Fw/+9O
lcb4ZFjTbCJOWrRCFwiiIvcVbpWqoFyoCmTmRabhFjhpz/p4WGdOUuokeuF6oqFPv7j60E5MwPIC
t6SClqjaQbCjuLtA/XjC421b4yOwQwu/qzrHZB8NuimB7xAsXoiEowjO4rv5Q5nxk9VEvEgFacPW
G42r8XGk0dTfi5xZ/PdckCv3wF9XBwvrfLp7ErOWAsWjm04CA+Jj/mLkNyh04759wMe9ah2jxhDT
m1z9KtCnZcCUikxsaQrIT0Gpy44mm4FnIxmEDXEGQpEKDF2EfUay88h7RUZmLalhI9KLFOlXFZl/
/pFwNpTvmG3k+JJvCrBTCkTTgAo+uOqOh2X1lPIk8s+sEt34fjUGUIrPacFSts36vuWRrNcnIXSu
jFIs6K8tOYcLZom4seWBTZ59ArciTVcqdD61EeZWXSSZy9dXKIQfos/1KEyi8U7SHsFuTF1TWp1Z
an/+MiL1aOvCtPbI2+ve/tJh2fpUSknx1M1/yIGNbEvsKMTdr1Pthf8ZXAM1+7C3nY/nVMuJkVvI
IatVqsX9cB1JpWtehlFCxyXT21QLv8vFfHaDZ94gZKOuu8ybHd7N3cMf5HeHFBLONmmCU1+iZwql
fKa74OaRZbjStkXzV/9dcoXxX0w14dIVEOKeyuKCadTYqPG6x5IYvBoneuueXl7+TXyf7QmK6zaB
Edr+N6j0Qj7kuzpPc0qy7ioB/3NF8USMj7E54mHSutzfSPZhzVQPuAO2o1phmXdcT1ZYXPWMcnry
1wMEYBRBmtAqRovtrvvxkcoVw1/eFMZ/STqaVS1xT1Ox7wVbtVsnzafE5bm5BadYCh9zoElExUWr
xrMBUBJXKJhaeCbu8cY98dNX6vXwg2WDzGtCS69LPvb37W+qxCGb0fd9J2geQ7aeT/MgoIu8W86j
QpNBRkkMHgt0ebxVacgG09yWy3AhXJSnVP7XeJ4GIuvMHKu9Imm3SCiotApkUXCvo59P3gpqvweX
WVvhgTTQfS4hhab43JIvcKYe/Q5Oa/xbnxubqWJUUP4od42MtGnm1GykhpCw1lBgH0JVCWG8fDxd
VWF5idZ/S2UAALp6d9h4n3U3KIjroq2CHMczTafpIrYS1cd3KqEsiCYsfTZJB5iToBsk5z2TNEdF
cEOhrCd6dy22OegS54rttow4MpmM6fymTidzFSmX9Y+19StxVD+rFRcmJlzu27pB47KSph04Ni7X
kPrph65TEerD7JHERlGiWG4g+Qn/axdA45T7LiV1OwTmnQJmsW1WDnSbTqWq09Kg8hxFgS/ObT99
i2qUPbKd2eSldMWCsfvAQTeZQiDtAkHKlpPi6VualaOUz9LeBoujq8GAglyBY5dgmUik0KOhLlt+
lbUZ4cUFDqBUrjYxWkpzMaaL0tOiT6HgF7sSdw6v9WeNlQD0mn4MHh1cw1gCHedyBxrPyuXqMF/P
cf4e9XSJVr4qBx3KRcMEOGGUk2N+4xq5iLYPki+Dka1+7q8bvIYXRYfJHyWlB8ciSbY17fuwLo1R
VQpV14h9fruH8P0UPiKKZogGJxMwtX9zDyRAlAUo/3zeSpDdr6Mr15BAZCWzRWNL1y/j1hEN5AbJ
CuD9ULbQiP0K5NJc9MMRDe1M7ra7eHI17KOhLQhzJL2foLrDWvPvmjAdiGd7Z+pElVxod9pOQidh
s89Ni9lsCER6Fss+W8I065O7J5Wb9HTYshOLUuLCmhjo81MFOfguj58s0XBwM5lKUVws5EwvriGe
R1fyhxwxJ1WEMSi3kgW/QJ5Deu4Q2ItbKX1B8xERtayzyqD3OSH8ho27N+1KJfVS6YqMqib7hcIx
vmpsLBc2AYxG2cQg8JV/CfRlcIHJPILOHZUt/TP6j/FWEgeqD3sUzSxDfesz6PJp1/ZDpRwSEyv0
U4PFd4a1Nmtm53kM9EuCAFzwm6TUidF1xroAudVCv5dtg7DJElsrIqRqNNEPpVMt+8nwepFesJHZ
xccwiktMxYFv1thR2cWFhkdT3MzGmhEUpAikgAAN49jD3x0xRQkY9aPJ0eQkuvGM0iUOUzX4AHRm
nbeSJMIrp2iGi0gD77rYus6FKfxcp1m8kW2bNKA5QOfB0Ylwrf20z9L/R9FTnNQmARfuime98CX/
ZeTJ/2eKcB+hua7jo589+1iY950VoOWIaapXyWXyugm4/zfPA9VxgSnKNOv9UsILqm3phmPMjV6A
K7FnDY7XjWaTXvMBdmLMbJBjjrZsNXIS9525cUFMBWDSy+Af5aVsbkRUG1Ka5wK+UPMU99zibo3s
kqjB5ULmBzIoxXi0I658JlYkBCM0F4IOBsI/SqJWkteHc1HPd/tUjcky8FShjMo6GLkgkoebLVQ0
jFHSrDLEFO7KW/zJcJoPkOKE+S6UVGdyMHSE215IJ2/KXi75DzvPAR5uEObXnCDKIDaB4pQYr58i
Lv4yhaXBDKOIQxPRvr5ETcJ2PXftmyJzBCOFBKqU5ZV8Ta8JyfyoVDO8GWP3nGGRyUn+SN4P27/5
E7R7o9qfh9kvtVNhVBpwXqo4Z8zlSi1ziTWjdSJe4/261tioPqRsrr8TwdC2qzd3NuKJ6zLU8T17
OItyEikhzIH6TXh7BjKcbx5FZgdbi/Un+oZjOZINwagTrFRB4p2gJEWKVxJru0wdgEP5pkK5J6KS
L8ZJjpx2N53TziiIt9YtQcNZb2kti4oDA5nFINS1CFyLs0jcZYHKpzKJC0daoTq6mloAFBB7/ZWx
u9krLWe+8GqB6nTLGlyn7IHLG/k9MNyjTlBpOk6n3gvJ3V/lmnAC8QenMW1hM4t/XornG0e9B5IB
BPRVak+wsDht3H9b551JAfcovZ4FkpDsRCEIG68ARhY54yKkQoSPTAL35KpMVLeaVt4lflvNc9fN
UcEWPyrG11AZq0gtpPAfUR5ne7XDKku90c+6OWCEsuQ4q3B7iDkpc1Ig8+gvjtDU3AdgoCbq7DzZ
IzdPFvQsaxgR3OelGxcpyP63xQOy+AlA3xrmhxOAwNdxlKQKQIpk3xRucx3QLyCQKNOn/ahIBBgK
cAIOMxDtD9SQCFyYgx5MP4yXBsM3Bd4Qh7Q9Y4zd8pD1OKcSjQ9vS2sUv4kH02ZLorlMmOgmkNbt
aAZ6Tz1dizUZd6JqiDjjwjTMJ4GqRPxh/7cc/yKA8YDNP6bE0AXj2T6JZEF2Q02I+7KJJF7TEiar
94hoYYIiNMtyLDZBKZiE1Zmkf/kYYLgZt4lN4qGcHJOH1iXuR/2hMNbGkyiCdiDkq+APcn40UWYl
VJnW080RvYmnof3pR6MGQzap23sOUAH56jFIQDlKtcrizotjVxuVTGNcqTEgZKjQpNTBQX/UfCmH
Q6M1mvNsWq5Cq/9N1sKiUXjCIxk/8eIezPn16bItyWAaLgKrq+v0Tp5A5iuIjCynJGpflnwqUi5z
ZxXkx0IWl49GZgEX1nhVqTC0hfmAke8CBwfcH8eAQob8dh43SOtZzW8oY4yQhW2ciPJ4tg2NeHTa
vR4i6ZfxzEF+VtaiGGqwzUlW48dZV8SgZ/V8B6BsalrTrRy0qapEsjEmLSboo2jEUo3/klPlNaGx
tASCKHRUn3Ld4lprK/kjjcDDCzATf1Q+t4U9D95892P7gi5TH/F8B4zhL+CXfTjBLAF80YGoLNM6
hacRHAY7eMYwJUX1rzD6IiKXF9m2FHS76Sc+4BdH9YcogjwJM5P/zj6dRuenvsilHGjARnTetB2R
IjGjLbcigjRxo235adERejMlyb+u+2vUVtZh8/EhZMOs8fuFcsrO+wZdbO5gj23wpunGQTWWDwYa
klU6J9MZDedFiqvzcGVLIeISmRYjJTJx/5X8W78IDd+NMskUmFXDdXbP7OTqeeyKeV3M8sldBsYE
h7sZV/0mELdDwJ/TOME7NpSTeNnQdgmYqgM0hYk1q9NxStLke1hHT+bQiFr0f41agxWWrhZmdVl3
HHRZf1caTDNQhMceCXO3R3cImivLAjlDb6UPZAWPk1dBYMqIz+sqOtsj75BqxOo/NtLjFJ5xIWy8
vNr4hkI38JHG9zJ0kKug2YcxIZnEpqoVRFWey0oZbEXlm/HyWMipaAd/ZT73Zonxmu+XtDZIa5Cq
IDdMXUHttmrfOQetM4ZxunhWbl2s3tDpkUKNzfxFmZnwaghwLsRRBVQKWQERXxZUuKcUp95KDCBF
zvP1ciINrW3FmtdXP252SI1wByI6lXaov+BPXwPZYwPJuPFV6wxUIKkWnCaM6hPeMDkTwQq00O9g
prafW6z7COrnIq+zpkTHoB4FFi6fvHIdbPDQH1oXG90Ue1L1Nu9/4xwBrXu51+Eltyk7RFrjJmGu
ky+AoUU+d//Y6aqWgjMdIJtCJDeqIeqByS6n6ong2DTmd1qV9m3VeWqb/8DK4ehAHkVSTIT6GPNu
Aq/WDiENoiSP/4eXiW1XM4MpW8LrTTN66k1CdULksT8ykHTtnYvA/lQcJI2jfLZ6KfY7nksS6EAr
MV5kBgaeAuf4EECE8Ix6hyFYyQhqpeeZyxKJ9VMznfAMikYLDLdnsNr8ObmTxHumt2FgEhAm3e+t
WiYaBoPwu2X8/LYdR4nK3H2PLTr9+z7u9Z4Sm98Gnq6aLDo6CRgfTJJpUWaIBj3w57J3gPxNFFy1
+0jqAXYCo3rUOcXVQcY2LwjoGN4bV1SlxBrG9i1wnsZRdZQp0772qy/zjS3ONpudk6I1anaBQ58y
Lnv2jO44qyknVGlwO10o/OmTLz0iV/4U9gzgFE/jKXuFCsd/Q4I0QPatMxp7TC+TFjqmo3IIDz9G
QBFvodtZEwl47sxJL/u4ewXELByA7TBumpVgLbdS2IdOttx2rTz99UTcY8UZR8VxTQQj4LJ7Upyn
ySmg04eAEuFFLhiNltmR+IdzyrCXB5RmfPgn+yxmEEJqNlfjhwnM0j5pUkZR39gl5Iwb+3qzda06
W4RRvyrhF0/nfH3UDoP417j2m8VKl9oSGU/ofnkAsoHC+8GFVoY/mrc43Vh4Sl/F0HLW0tvb4gbr
KiziBizTOzBoGqasjZ30aOCB9SzaYxONLgZdE4On+I6GdyhYZlBWLmPYQSVM6dBBMc7xybwLyZrK
wsMcgI4PR5I6b+xT9+TZZh9r/I/s0rwSIxsPrdwvWU16bZkWQO6Mm5Hugs0t312AIEsl6xx8JQ+b
1Tm/RDPvm5530Y+TLGisCCTDlqIQSfZdPzuwROEBAwkba6RL1AyCPD900JxjFmYr3aNqlJb/Y1Lg
9TMigHoShcIGxUZjZhvya20Tcz9I6NTdyTFoI96+eh7xA6GhotfRfrPCCiEKqghu4rOtW9PO1iNE
vB/XKa+pxIHdrn6m1CLBXciCWo0nDX0HapW0HC2TLPh94IbSOItZAQUiRLEIOj7qthFkHKeupYYk
adZtBP/Au9G4Ftd7Zm2ylFxPK3KPFyAU/7MNRKzSVyJzw8LFNrz3fyIuxZQxbvgwsfN0JLwGYxdu
Yxo10cRBOw4JXyJzOaK801+lBBPZH5avv4omm8l6jyK15TUlj+Oqhi+Sd+zX4I4nPPmR/41+bWQK
A5HXCoiRLRnUqwnNvclLG+wPNRC23LqKYeLEcyPxKXQ5qNn9oATylARCQDtw+2O5gtRjnkaqc76e
hRB0iXyRs/NN72VncfrAKHXhslSei5rcFhk7CTTmWiZM49PVnMtlfAcdxog7XT0uXdQytpwuvPhw
Xp3RdRFcwWPZTsaQTIy+G5HkQCIN/Yb+98AkgPyNEaKIX9RmeEphr90io59YZwZ7f58MRCZNPe6G
cttIGFmlIAforLvtwwDPLyc9PDJ/+8kurznFOrmFMmVdIEzLidvj52R1hD1eDMjOgV14L0PrDzq0
B7c6mvJ3JMcoqCU5MC3cmgkBb8vEkyUoMVtdVT/Dvfl5qy5DiD41ZaMnBXsjlt11KAZmkBbB6AGW
InqVKl5AmU/tUqWHL7T+PB0KUnfSNOzWjwQCR/8vKOaajcHtooOQmqqJ2ilUvL9Ld6tbX/9JX6m9
VgxQPbrANrVTkiOMSm0PIum6Ek09iT1p8x8DxDy+cvQpIwO775wUKImU1L+likos0Dt0VALMSvO2
kAKYFLubHKi09DoDhvTwkmcID0SM9ie0JM0SC3kfbA7IMGuJU3rmBv3j2CBx+bVYRL3xd9q0jTgk
NUlyrCRsjhbZ6csmE2Kt+ErAUNP28DrGM7utw7HTD2w2OBawgXdJv+zxzHk1zWaSLC7X+a0P1/z5
TyTUc2AFSEoMfR8U0xqfz06F/zWKSwh9UbbyD0eXjr/gnn3XOtugXk7/8o7fxx+xIHguNDE7yXbs
a1XkMcrTBB5Icrq9oBD6UUJHYjgq2b2i/9NsH2Oa60l2snGDfTZY+4nYGTcI2MiLQTl859uUPKe6
o+TLg80idgRBf2A76tvJvkVs1fP0Pey7FXYTrS1mCZ4QpF9gklOuHG4EtW4Y63lf/GFn83zCCaC3
kSdQQr0AwuzD/lGNjJwf6S1GbsA0H3YerkPIqiNO9QyoEYErn2zruPcDtD3Kb0txqYWtteVvorpt
z1kLuuLrkYakPhk4AxXRb8ymfD2VNSf1M6tOIG93QqKAfxm+X8SrY3BRzDZTsWl9m8sXfK/vVpj5
vo5DFu0FwU3QSNhz33ew47buPJiMqRyYpwFrZWIoPmxCXNIOglITcX8TFKdn+fsIu5oOFDB05mAv
r6+Af1lufwA8Y1gcushINOBR0trsPgvNHAUCWvuX8qGpr9OfLscTy6m3J7P30vwwSXqcU6edgTDw
T4P+PYQwVADCQsfIlYm35LIgqzPZv31MTh7sf2vER4TXl8c1M6AZNTS4kB6V0AnZRS5itf97wM/Q
RuTqP6YEgD/5Wxu19wIwJqeUOjnH7mzs4xDqWfnheq1EWP9MNGyfyL+D/H0pwzBAERi4TRbWE7i5
usUhgsp3EUT4F5hz8RwkxCZxthpiQDSVvuC2xEkU620qCfN73Df8nW7MWksy0wTLGRezegY19ITD
rp+v9D+BczCsqfdyRwTrsECuxykexJlHMXbtDE/IAaXkfL4BdhqRw0LPL1/lJIQvK7KgD4c4giek
EBv6Co0cnIzjBmBN9WpnA4dVsmK1lXmbNXTmmxVIXLNT7kCvLH7dY2kEC5EjsWjreN/5e8+fNraF
5l9pap/G733Hn+MvtobCW1SjmCloxIhcP0L3uCteBXUU6Kz/ZuwLqT2MXyeGe32vZT0PJAAyOJMd
W3m2qqyk6OPNGSF7qvLKup0OF0T5YYerBsbhas8KShw6FC+ZpVdIhuBcck5hvEf9WzrfTI67+A1l
ebe84yszBp6QDpxET0PSAT+dlKecY/Q2lKi9Ks3oPprOskngrGAmAeDFaYDlD/YCo3PUlbEVk0i4
w4IInQeakqP+3e2yRmnMOO8JYykgNRXmb7PNJHNSzfhmCQnAnaeix4NG8PhVI01YUNfMkb5MiZJm
4JSZe8G74+dcXSnDOVEO1/dzecZMiOcV8f+HvW+zbrivf6Hnwit9epSiZ+ONXTDvoJM+/2e4/Kzo
EZevb7ESyrYRPjOGKpfoJddAjNEfaix5242MGsK6k6PWQgholCYmwTeWRLBRSC0wbsvsZIwF1Hjl
cAX7QiE9wUWPzIf7jPmoQze5oTc+jv5m40mdKidoHtW06pFnykclKeUBMU86lwstHwJg9sWiWVYJ
zKXWPgEupq6FQqlsI7MZ0xUrYfOvYKvhf2JEMDXnRSM39kctdkHJbkqxyFPr55pEKgVluNTi5PZV
y2E2zMVsfBRV7ZtwKIv+YYKE0CvAjbGnZJUJ8BMdHn5TderlUb2lbvAlFONUVMIJcYo8mURzsMuS
JKVfgQJ+uCDoewM29o2pMv64S1/dqZRJ8WIBQvhgBYdexL1RRdu1wLwqavklvJNEa/cb0+mecGJ7
L8NW6/gxls2FP0M/nJ0TtJ3IxcvbS0sZ3plY2P8g+ZK5Vm1Rma8oYHkPfcLdsTeiRTuVXdvileWP
YuysspJGIwSLj5QrZt6Ps1cV/+qvivbYQDh8egnmuaAlADOtTbhfMsM6DnyskKrb++qPTp9bvvSz
0ZnssRXmdHJVQ/bNY+QYocSvDRKxcW1eZqt7o/F9B/XnRUMxhPu0VXa4h81FURPFWf8h5FHeCh3c
34HLT43LOMqHlyZiq21JXkc4Ia5j+ZAVkUnQCzbiGRBbaKdsmSyEIbogaPEAK1qpsKr5FImiN26K
PSJn7663UmIjcjH+I2dCgBQIrzVM0gIAyGPiHf6pkHbCRoUGM/XaErvIQPEvjT41qg/kvXPA+Ja8
dS2rIOa2p843BDTC5usI9gZ7fojWTVw82eH20AhIgXJZe6bJRCM9dYBbFlsYuI2G9p/Cm6JSZ93C
PrNLlZJk8ADoQ1p9byEX1fP1yTBJqqJAk7apBIe2+lUbsXt47apXq9F5sV2ikLcpvExaLBGVPtNc
9oR40A5iNCRoKSIkN2FKjyBiT8kJY+WflzHWK6E9SomAAEPJmBZPSV612YW4B+KhYbIB0hQAcYQj
YnPvfLrS09r/dZiSa0xzEq5E9BPOIoC/A7HpG5q/FQmd5YT2gA6pGzM576ImLXrRV4C5ZWkr6NPU
s5DlZRtMxivu+EYi/0WjrDpSFtlnG3cyb3954zjbZWC028GQRNeymNc7DlJSAwq9glmBMmgpFhCs
ks+0Rdi9JoNCtR4IWE6v12oMeKUNJ3djNGyCnPWdr+QVZtBG+ECX+ABbtqJj4WLgPaMnigsj0AGj
WFmshDm3+ArNGsFElj33kUMFbnlhSsKDn1GrE2BO0nrN9nKDe501HyBguvMg5wOqLN2o4kz76BiB
+50eWUBdqQNHfejFLHTdoptXBMOUQsvCnwi8wMJoTKDBoqHXZuyByQhaSE+eNu71AcKFD6nLNq+H
W+s00uiJM5jOR/4cRrboNbz7CsVlIz2TURrBxHtJHK6MXy+EYM4Z7OwtGBHGHJniE+M4O08PlUGf
4npgTwSb/TIL7EN1H4oFz3QaAA96vZK5uNdu3f4boXd9EOh4C/Tg1lLmt/cNrc+KYSm7l/P2h9fQ
taeeXZSLAMlfoG7pCyxff740ocdIXna6ERfvl+TWHJlij2dbyRWr7c6npwn19g0LkOPl/gaA4gSe
5yBk758bFX8pRF1ps1o5jbSw3iMA4GyXQGSgYsPIJ3hgJDxfCGNgr5OE/BhrZ1xpPmLz/9XcIqRq
KuSiaRJycfEPMWyPJguby+F3wJoI60vu5Ta6l7qDrtO+ZQCrwLnbGSf+yK9N53nXl9mbi5pNw2GH
OTyS6btUCKTJlhM+6mEIYUKIle02YFcU4rE1VG47HAWthHP2rHneA6DTC0gWjxq13P+hZl5hnhdY
GyrKCWxApWGV0kscA9o6zh6szeiFudyWHGJfeRdr4t/YsvIMzdfu10XlKsdymaJ2Vg/zwr77Bm9V
YYPc+Mrq3s8CC1TD5egxKrgG9dGTb/4coyR+7PH9vUDUxBlZ0Ol2pBzmfH4dR6h0kzxUzo9pD0o0
3xRgy95rUCU/q9es3RQs4mwMgQIS44ICQNEwaWkH6QeSFuJF5S1g0RYNzM8W7qTqrIt/2vJjPT3k
RSjaD4xiN7yASq3MYQeJ9TUBy0N1HjK9KGK4RhewRr78YizIa99B0y1X9kS/qrqPPFj68ccscKK5
h/83WNVbQAt1acr8tMEIXgA9qrmsy80NrZeUg22FTm32EUmgyrihXYMPJNUZAapHrLcnr9/ejMcY
5zLqkB51p4HVTKVzWxLxjxIB7DXEVFlmRpKYkvVSGjyu4ls98dt4Zd5njF8Vr5kXMz8jmHER1VqJ
dEX1n0XFs6momkDA+YZxElat8fo1yIruMHRY9BL22GrzD3S94Vc/oGhBK2bl/LN9fAqe4DUmRMsv
sFpyVy5kotYOPnLoL0+Z1PwnwcvcGo3weTQ6ctxnnp4ZwDHRUxz5OwD/ZE6tQ9L+3g3yMMlM7DhT
gI7gk1MJM8LnmyMm92OTm5Vre7v2tG5O7KvSmjhVc06fE+4A+2h/H+Q7WOIRwYnNQJOv+Y90+ZxI
rhvo5qBMTbHDByYBB0/aHGZK63C6pPqni7GjiXnaKee+yv3oAaTPo+vXq0uXwNuDRy0jIq1EhPRM
JcTzqXrLL8R3OpvQb5PHRmZaKfuQDMcyws8YMoTJQeMsd7N8AsT2CWEhks2BoES6Rab0IMSRF2L1
aHBnk7kAsnlD/V/BaU2EwI5oBck1jaEHJFszeMM8WIChPO8oEn2yEo4UZA9bC596bRzl0obGun2/
0vwLL2lLBBbWfAnpW6BRNids1UE6rjNNaHunO3yoFSpI43RkQUUhBIocpRKkrJk8RYpCZx4JTDgL
BTumH5XGLkRs8/bBLOZKZslvDMoeQHSaL6ztmHPAqHe0cXrY/B/EWlwxxpqfPMuEjPlLuwvpV4cX
ykfU7rhAVVghrV0fz4yrbgG6KU8yjbhnCVeLBbd/DOmw5YyiTcGY/ulePVXFwkRntbRrWoeIXek9
2+6GMYzEnNAylwumaIp+ZQ57jh3zs4hCn28Mdjs7AQeBqTeJyPYKjBBzVpYmRdkAIgJigpxb5kwK
tdzowA+TEICIXn4/e3xNCDtlUeIbxow9TzlXvpQy048u3tAQwqGZtr2+TTbaRgytVzrMAUj3wGgP
4p9KFW48q8sWMRMpewbBkhycp+Ra30AR93fml2XPYDcK6RlDLhfSjRsZ78UvyNcIqDUNR6Y4Jhm/
H9ZKRP23I4xHg1uv5En+3yLeOBkZ3k9+FB83UAYAZjvYD/4Bg542yvPoT6+1QB7Wodsee3ZEvIqW
yyo3MZ477tGG5w1alFvEFetDiLyrfsweHA+zoYohzGS72tllKLSsG50cwtdZ2A1a4IhdAyOnqr39
BC8mEEPe8EaAPlq6J11ZC6oi+j4ORsmHZNlC8TJ2cAy90BqdRthpdgCDDyOdI8S5Eev79dLz1yjg
9apJ0u3rIzc56K9CNGk2cbNegSGL6eWxk2VNvYDGFHp7aDi68dafHVLo1q1e4cQHX9f7qpoGmTsb
H1eYj5YNDsqVccZOVRBFjviUqcMln8bLdei8h/mhl3JCRJ17IGETJ8dyVqrkPLWAyHGr3G2eryB0
CjDkJ4Q0skptH+AGl9tBNl9gEiefISkjLRcr7jkwm/1rarotB+j0OWorhEhdLZMz0bsiJrN24KyU
EGclgizaNSQaIAdaldPNCOc79GMt1tA5dbQnaMEsC70Vk8HEFnbODfwEVoxDGNNhEnL74scM4xQv
5Ryy2NbbFqH/uEaFXBEUZkAE1RZxqB5C+MvEz+Di6Ji0SFmE+XGehzlENI3x/39vwMh+JSPn1y+e
InCB8adMeoEiiela+yrb6XFv48pOx92Ds8WHd94WH5yneEbsbxoceX9FnHutr/4NLQ5B33KXjA2r
JmAKWhHDtZ5N1oGt9DAIZNYJfmMjFAKjT4CjnTz0SMdn2/T9IjS1DnpVIJmS65WgNxlBtSk4pv3A
n8p6fIO5ev/v07HdAM6HCgeBKhY3fCwZZEE9C5aIbATjnPYml8R9LWelR4e73dPjCKjyeBsi5lhf
d+d/Q1aQabq0vjaRk5thYppKDow6snrbvYLiwcqGUipmrzpyYTJVJz/HZKp28mi9gwoIT9W7ShLW
FE8zBnlCtHkf1Jg3G670Xq6FaTamlBgHaCwu3XCYKIfwWq6z/1XpXevxWHblUh4lGyu54EwSkMKN
GIf+PAVuZc02gzp03hq1ftiANXS4wBNXgWeJqjWswCAehUeBiyrNXkXPt4y5qem0UdEhnGRteAwa
5GLjd473VDG2vw7uC2UDCt0hjpw3YmKo1BNUYCyO/KOSVwES7ecwJh9DLOn7wbHUfBxqfqIYzY30
F29ldILzg3Cq1Ug9K6k3vxFYTlI2W56bkCUNVfPr2BnIkeyqWreeI4/CXfIBs0aREPG+ykowDDhE
yGZ2ZqoTjvCaqsbvK/i5op8yDC0i7gUYgdzCHq/C6NNrOc+qDj1kU+YOsMhRPC+cCVKAe3LBDEkS
CPjCR6jGA8xXIKyzFOn1XfrZYLdccyCjiYmblYX3oOXKk7e6lAF8uwe6aQIGWnlDFRXdlcU8EILT
Suk/jpj5oilKsoe9PANm5/S2UP4JzkMmh5usc1ir/HQy0WBv20KXcQgHoI9jRbJWhpGmP+FwUQL4
xwxz690E3EV0KgQBxAeyW5ZhStSMT8YR5hkdoXFAoCcvBRXijlse5Ba3p/nRkidNNY36gjMStMXU
NHw++Knxy51Xhh9PVpV9cxhpZXdTewE9ogpNs25ajqdpN9ODgKmwnCD9oZ3UJtHZBzr5lRJtEb8Z
p4G+VnyjG13KgbA2H2Nz174XHRuOjoZk2AF9RIe7XwJ0ZVd5+h/OA40lFvCZ1DQi499U0eCkOhP7
ofU4WXn/hO+C13TUKJVvuW2PUANkw6w7N3I1Cii6HRHMqBy/s/sXI1NV/hvZBA40tdHflTSE8vxG
Lh2MyYWyMN6rJqG6VU5agL52s41IheuVInmt5jXcyFUqWQ9e0WfU0aA9HZPIThbVbYWhS8Ozgvj4
Kgccr8NrDdJyClYkCVTilvxOQ1wxZtcZAQ4MMUsIgn7WN51BoohmeQIy955O6srH8otUxHoau6fw
F3n6nv6VAzcSIFm4+DBFNCEmZLOlNeJwM+KgCqpdjNjsGF3XNHfXlcW56X09Vu5hhVxwEHbyoa+9
+U6afNkkGp4X8REHM4yMTZrUwGrGtW8KAOMEZZCMGLzNvm1iO9l9heFXUyvXoB+wwx/ZO4u0G6BZ
0reAj63uvMQOsHL1N7Wou93sL2Z4vnGAO49E/FVbkh/IqCL0B9jr02lQg698tjIsllk3SkCpiswK
9wAb236fvaJQC89QAh6Xp47SJ+ogfbMII8XuP6WogfWAm/Y/tsIkazTN9Ny2tNfWb0kzdlbP/lL0
6WghPF51Ul8YVNBHwu8UiWF4B8riMcvKyYZKlPvB0quxzBT7oWV61jKwcey5cVIPKDbvQtSOgu2X
DrnS6h5NH/J1PC/yq4jNgnaUcz/pJp4tN1NkLI+YNhNw44BC0hQ88RMskmRChLazW03Jtx6FnGHv
9KowkcC7PARXhjfknqqXiezpMO4ZzddW5Xxv2ozjlGEew+8GCfG0pGwOeMgACINUQ+7jAANmLT1z
6DUbKhHlvp/s0uhYFqsC5P25wkcE3M/qaU/BOglFI83+n2fFNAUybOO3Q3L5OWsw7psF9tyaHsM/
tuWTxlhWgoFLimsCxACSGu4g9eN/6akypDK8kRmo6GCgxnMZzPTQDRnXxWSgXc+u1IV9sIYNUZwr
ugk6udOrHKzM24XkeWss5gIH4rAKfqQxwqrO9YPnkzVwIEnICs986XQBYLXJOWRpzRmdvq9ipSyQ
cQXZnGU8ELJepRNpRnweOFE3c9xbJrMf6F0X1Jv/414T3xZLsmOnzA6FTFwoMrBZXmxEF6RJXbM/
5hiBhFwjrIC2JOriBX0a/ztCx9JBDVws9jlTvTLEDHa1UUCfNrbyeK3PufYFX64LK+hZ+zfpMcy8
pmlqBxCUAMHFvZ3ff/35h6tEtRiHro0MU+XZY/pYW8MBvuWnpuZDJPIMobi5Bvq0LJAuLnoEBPIi
Q0gFBp5e5F71tXd1vfpk6OJQCVi4Y3ynEZBrVuk1wHz7j8uYZ2mRBTm3DiWELcEUeIT5oJlI8S9u
LIaj8Ceri+y6Lc4J9maS4LJPMH9eXH93DjZa9ltZJxbGkHybK+c2RlkuQA6cuN+lG0SLSRUsYrPM
gsZu5yv6ZXQhvTaGCKxVpj/qSiEk/OOabEFUISi2Wd/pKqTckm3nhFUkfDc33LFW5rT140UiLzFi
fqeBCin4CMBzSvhMidjJ4GeUZzDM8LpG6xOINZC3Yo5Nzmtl0O6pDJ7Z57AOzZYu7WZhqPyxpIYK
nfjwwlVcgzbI2SISx3aleiE3UXDpzuJkXpNr/H4fkfD0woccSy35W1TslNB325CPagG2RuTSygE0
w/gDtNKXbrWY0s0n6+Phr4ccWT2Vj+qXMc2Jouacw52A8iQXhm38hplIC1LqdnSOaxihUH3vec0H
BGpV3tTKcXa91YvP6JAcThO6rVQem4QlfDwPA1Jz4amWQMLiFp2hqFXRDRB74ij0pVluvlNbk+MY
z5f/SsLOxoI6i4vpjB7PJmwX/0cYvITzMYMzezsRJCKCpOoPFOEHZIv8rooBg4v5D/WRuguXKLF4
vf0tV2uMhzmX6X/USuJpHnASeZtfpqQYXd6szo7hv0p4GbmKlfovkoY5qdoyDThdb2VJil74LN5/
oYkTXlgu1de0HeyWwkxtP3aWwTWJVmZt/XuqlL8hMHpl6/xoxxIsnci+2gBVWYaSTLzcnE3qU6kX
uQ8Ot8ySVM4LSqmm+6na+ptkju0oPuh63/ANJuGHqHlmVIQXvKglhVwEoZaQx749AYz6ZIJnvG64
2gpo4f+g5mtqZvesjHaZiUJ63mfYpOfo5EXs7vEHSWRhdczwF6L5YHJuKfAySwgNT6vRFhHPSoC8
ed2BeQ/mv4Qfsx8CdKZwpfcOu+SuEs4/2d9J6cAgkZEoPN0jg+8J8e9eyKBl16Yb80C6cJhzVH/U
KTGR+3S9gCwASQx5IP2b7FBuzlPUHbjVFJTlzGAFwfboxOLHVX5DZpHo4DzwX7OliIhLbX5n2o6J
yxDCWZ1Gu2e+HPK4kHh5uuAXEYWmevq49qRt6hyW1zJWlEmi1bZcHMbWb0p/4TivYYG7CHznBTt7
/LRrd/tjXyVNQrkpxzCXJRnEcuwr7FUyYivxKAhWMEZdYVrETcCNbUQHdk2kWhxhUQ+PKp4ORPud
lw37g94FtP/lDMbmZE3HkDlS7l3grybt4jUGrWckeIBpuDSQXXXR75BPLKWHvxgaphE6wp20Yyfj
eZbMqA44vmdraGj+0DruhLlyvj14xgpzLOjyhZ60Rga4+KMVYSxTKwvXzytpZFe6AYRLcplOEyzu
3yRBsbEpMHATCWVhDpNCIXpO5WXkPNM9h+WiMYgCUGDSexJeB2aI1S/XfgftQ2fjtMUU5ilzZhal
F4Y3gqYhA7OuU017AAkYGnWnIJFEmCnShYX1i+qzWGd7u3P/hZNs4A3cu2pU1t9VmUlpecWisvy4
p3giu/tSl2wNwOjkPX0CcJjJk8PPpFbWeQd4X4RoJurLcSr0/X2bJBsMFAwYJHWIEmdpbbwR8zje
AqLuSEKDCRcMFAbJUWLxCJ1Sm6i8y2eVAXoHEJu2kiz2Jxpea12TCYhDXcaYBOgAX7+49yHkoCE0
JVhL0TZfLICJ+wu/5vDf1UGS5DwnilyjRBJ0Pgi0l89enbQcPc4veJYdkPgLfB5hHjdYOlYG7Htd
OqJ3wIuQEYrSPR5B9zjdalKaWG4Yih8nImJjeKnJaMUCjTXaPlXLYM45U1RlYhmwkfrTHDCPkbc1
5TV7TlOqqe6w5D07UIHegm6xXWuRaqWjxe7kK0Le1oTNf6cALY5Ok1J4DXpZ/1eFVFbanvvH2/gp
I+hIPtHkiz0xV7vRVUBsuJ+aP8JYjiEupU6pur3YGix6vQdbXf5ksAdUw/G+43N1P+w+WTGhedz/
tNT2xXx9e435SbYmgJhBiYHllTbvhtCK22pYNDhv2vjK8eHNHn4WEjSlN4FGrLFIDlBvWcCh2Imf
C4S548NoQYKD4iuAL4sm5wzA62hmlRKkiTQV+u6OzHf3CtK08JqxXkpgqTUtn84wZ3+Hv1pF8OT9
9VsZbE4AJgwRkGNxrtxrhPYxU1/XZzX5bnjynm7Kq4Km0u0iOSsu6dAwZPsp00AV28TwTxt2gPyf
E24iDax+Iglnru9Lup0Chf8gIUYIgPvm+BhrRQ/TqEjen98fh8hB/4zMP0jyjksEdQtVRaUkIZ4w
CgBc8++99FdFy4VSwV30oMbX27puPbhzIr7QFc3r0zJH/F+KgLyDTKc+NLEXBU+Wrq0b8yfPYJrn
WU+juXXGBj+TuMbA/Jb9i0iAvYaiaC5Wy31vM+yZsIZG7S5B9pgvKfXhPqTBCyApuY5a8VVdCftD
k7y8s/S7oSHr40qfh8pi8gQ+Ei8GoH15vB6oVVkeT5nDxYImdtKeZx5Lu6MdoRR2qV38LuJN80Kr
dkttW0qV2Hi0ojccR/VCXQMLMS813KTJ1xmNOIdi6yQJ9EYPbKg6bVWIDIc69J/dr+XbQhFNK84L
7mp93obsdyotzSFdQhvQQHznyMFbOOA5+liwJKwO1FKXbje9mHC2BKEnx68/3d2RZy1fpvwAJpPo
q1AoFquPRnimkSXholB/RUqyG/NAHHVLlY6hCOXwg3leZiLe8j30bIxrqcAwCdGxsBTKzJxW6xX+
MzDkW0lPeeiHfedHzDas9DH6WMLVCfs0z9ODSXuyE7Ns7uE/C1sgZIXM6RlEyCMTZ6vriOE8JqSI
vadyWAFPy+rypxxAopCGN4a+HBs3ptnsEuVPWfWCNVczY2pGxgG4iB61azbLBCl5g2BtdK0zF36e
2DMx5g1oHVntG1UimpsDV2J7LXLNc7GJqJK7KjtVD0mCdQMVbeRgI3/t2iUXY5E7xX5jj1w6XVQ2
dxP/NIMfjNOaX7RTHWNyU+08wlpY0pxVW6HzR0/EQsZn3ZnZQSM5qHmZ6G1xHOI0+m2EGBYo3eLM
4faUzXcYOjtuM/JxrJnsyGYgmMqxNu1p+gAKh4FXH0rLylBplHHThr/J5WSY6x6NuCyC9Kie2H0X
UvBl0KhxjNcRgpf33PydKoFRX8XJJb2ndFLFuwmhICkjQVDouqYu4HzX3/q8msnUvUzBWkDLJh5n
cKjDteeFaoIoT4tOc9NEheGvueqMWl7fkjpPiByoO5VEE5afG80la3Q9JGPR8MFYwD0ybgD+tjvX
H2MyWbnD6VaMTEEsqpVLpWcuxnQp9wGTPdhnFt+XTaaCyrQjDDsQm4GVDhsb9Qo+xDPd+MPuS8i1
rwGVc2k7CSMcvTYG4VeWPQgAxoyGcq+H5A6kKehCJd3EmVbJdNrSq7kdNlPEHUPKwE5kH31Icm+e
AnHRJdZrb19P/EkEcz2zxwlx02D+HTmolF9gb+M6FA2EqoUQidtsJ7ARc9xqdbdI7J5uWLSaF7sZ
5/Q44EKh5EcTP9IgErkF493IwBUn6094VhptBQNkeKH8mQv7YuITmFMEBxZlDq541FKacbyNaSZT
hTzn/5PZLp/HjJMRLTHWqQP5ElQKU9NaSZ+15xlCvFHCRYQ05VjtOijH5nTkJn57Z3YbFjgHpfIA
dza8g3yDtax9CByADS9l6VCwbkd+a+RElowBmaHzHx0GuHavN/dTped+71E67m0wrcSGbgGKHz5b
3OfPbUf8LYLyBaVWFmwawDOAfq7or4gMGOK/bSnpKilvzLcOyUyAVRV1b/Q3kmO0DdHevLEeQ9Sg
hkpzteTegUIuU8iQH2ZSqhmtn7ra+h2S5zmzJJgkMBpIWGaMWlzCdy4LAiBNgSqRcdWhH/Az/fCH
yZgoqxCmttkdZTC51OdEnFXeon1Y6aWri1snKHgROjh+3G9jGsY8r3gOIHRHLF2NOd+YWxbQQwt6
m7/CBDFfx/3Qo+c6H9+v044UHDwDjFQIdSYViS3d5OshYjGxKpn7mR8kiP99SeAUBG7nOl5FCThz
sdY8kPkOVtp7axqm/4XDwFWEO7H+EHd9ucprk9EXXdVo50yl5QYRXuWS3kzCYPYJ6p/Awy+yZEUW
ulOr9QnYYqWdBCWFSsfrBR4v/aaWwdgXwOeoY8EaR+z+PVt1AS+qkRck2APyl23NkwT3zlsI/r8T
p4mDsUrFj+XFF4UIVNx0XMgW5j8YWC23W/yf3lS/ZxBIWyCdPwMTiAttpZwefv1XaL0SnT1g2jkK
spXBPeLH5rN2NMYdTzEiywjAMZM+ak0Dgyq3dgX9aZcexqJFQ56QKPgLW2/KeetUZgybHCQuTxnq
hnxoIEN/rrIIOqLTQllZCXPkDGp8mWrZnH63eBGypli16SoAOGuud1AdsYLGghQtobR2SuuBJazo
71Dw9X7k3wGUpopzODwjPTay1snjgm3GTivFpcT9x+XHbbqz1ZqY1KcI7txgECRSHQt3Y5jImcyP
J2CGl14LLkuzXVc7NdTaEhfJZmfvaltRtKu7KDybSTc39+HVvjjPfMu8XkppBKADKVlqdeq6+owR
v7Xx+40VvLcdxCRjDMbWRVvOrS5FF+E8FhTI3zb6fRxV1dvEztOoU4Kk9mtQwVgb1wFQ6t9Rb1tW
gCWHBjESlku/aNijADfxVW434abaCdFJXlEKPSVjXYMblJpVmTo1VBxZd8gXjcatdqlP5/5zOu6I
k1hW3+Oo7gTisKYGglDFjwLp6yhCRQ02XG9casXqKVmSDRzspAY7YHc+WOKaaZTImZtc8sWy6BPl
LrFpzcn1DBMkwsK7KCI8YwZrtt/lD5tAT2Y8ea6YWEUG0zLv9zY5jyucnOVZXIFPS6FXSYxkkBR0
XuuH8r9egyj/8Gw0Boj+SS28wf0JxVkXdc0X2Qg/HGQpYCkpEaPHehkgTsTzvZCU33/Y3XeQNqbv
M13jc/cJePO0GUqOLrh9UcD70Zfr+33J3W+YkEwVxwdi0UXIEXV9pPYZzCjLeYnD1WYaq8IGfKPj
L9booB4IT5iNoAwD+OHxFgmxnCD6WpUClx5TKx5F1TbZMs+98uyBiwFVhILm+a2ZJMurt6GsT/6M
8PY8x9pewrqeiRXmPFi1PRqigX2ysMWz5iSs/oasQe+zQUpVNJ7w/HDLRB1jweSwvRT9PMU7jMYX
K0CswU7djQ6JA/X17kIwEqULP8ChScjUmkJvO/PfrF1qXm2eiYRubF3HpdWGoXrtt0Udo2kqJa9g
GjAO7sMOHQPEZzCpIPXTDwYQ4eqqDvmo4KoZIA0NDDUStIFAuEiQud1syaJ7b0PDZuBDXPuxJZ21
zjlTi2FgaRNhvuK0cHSw0XWPtwOIUfUl1G0xah5DCUwXXr2iH7HzBLgB/HcHt/XaXSkyGOu8xnIW
P03c7yFJp18IZPWrgXZ8qjEoqLwojEMK/gAe10CKHWq6vJjv5/668TISSb97f9uM5Rc3GQ/Erxg0
hm6VfAdbKdz1ruBKVKM4ymKXMPSFouCFsQJzy12yrzvP2dZRlNUimD8nhZZfRpHY9kuh0XJQIRqt
cTEqukUmVEeMG3AmZq4mW67RBp42+diV6hn3pEz86JQ9lX8mjCxNU6foyaoE+iIlLOuq3slQEA7B
AnE0NgR8kz/Zv8Y3BStxqJC4Z9+yN8ZkIdQsil38fKPEMM8CstZh3uBkte3qFfHJ8pE/1JTGi3ge
vvdvahlL+0akkdhawYgh0nnQ7VvGi1adtW7jygVJPzB9lxuT1QXVPORKwNyI3Z00NTqDtBFHVvBW
60ceTWhxio7gMsQ1chv+8Uk/E3akI8rTF6BDEXZalHIp8k6BBzN2ev3Kj3WhTndrSJ3tb9HLLNZG
D6oJln+SmCcXXpXAEobzx7OU9s3GlAcYIdUkG8pXRZLWLiVtOt1/SH+AxOjTWSubOQj1JC+ffUoG
inkOVHMo2eJhH+4p47UqzoSr2xtsMo8VcPkbXaAJ83c/+sZzDoZubVkjVIz31aIuehOb8TI6sVsM
EVnb7KA403W0vVhD8rDTNjeLXT6k7sgCfB6wxfIkFuMdTonqC21vFv109QywtGUw143LzG24sl+0
eQCGXre9i3ux4QENW4O7Mc4cs2TMTUL3VYO4VsiZ8hFQreJh28fQjfQzlvCpwDd1RPi18rDPYbP2
GkdGmnohJVswDjezque3ibTjABF7IEGMg9hcmnKaIw+yL2dLmsI6zeqTbJ6HvlhgL1FhHcIo1zmp
Xrokb6dkjsw9tr5md6lOevKrHV3ZxYYjOExlnQkPwq6IwOv9yNUNAxSsaPTyuFJtzLpMs0h4bYnO
9XEXDLP8dNtgVw9cMXvBMW9qO9hb+HZkQyOI3GbSi/hk0SiRv8IDMNWI39wiPS/w+HL3cEftNMqM
SRTbSgZpWoLv70C8eJ3UhJl5NwxRyxnfJjj3RVASKtMktBs082pypECZFuJLFVJyvpoT2qHoYI2n
UZMooubZVV+bKARpNd+G53jU1gQUy+u34S4N89ZhogeBv6lb7xEi2EukymmevULQPRQ3q64f6Yzj
vfe/dgfXpy/p6y4hLSNzQj9DKimNvU15P66s8/a7fGGnDF5d+7AasQy51HSAP1ZvBMdHjNyhojui
b6frRH57QJ7I5CaWVpH6t9ulQxQieAUCHcdv8Df03SvhXsxTq0YcIr5S+fx1vFDzLOSI7XNgjGfr
gS4UvI6/DalOT2qsLoAa3bQEzQgWiMJOkw8UfyAEZIPvgTwx0TQ4Rnb9D6/k5IHao080rbLjnz94
VmB0eLFSrnDUMYq2wgPyWK7set5qYCsM37mUFlXVmXAH7hvuANszcshdYzFdsLdPHnmIDFpsdpF9
zMkKQ9SBEo+a4oJcD8M1surWdPKv6JN7j+dUg40GGO/Pxyf6KCupzqCUmYfJ9lhaY0I3fl6Awuzx
GkYAFB/5mGGm78OBLImv+9NjXDGjDYdCWNuV3dtx72eqb8atxSKRKMbESxSrFiMKqZ7GeZ8mx6Lr
GFuBKrp21R8aCIwF16WIsAc0ZnP/ffGK2gJrPSo0B5wgoC1Y+30l+PEAQBPI7Dt88sUlEfpCFF8r
zf/E4+ir/rQLbVJk0BW1r5eDvnHW6LLh/VqXSxMXuhdWrQ71ujZAOt9iIi07fi7suMMwickLikI3
Pn8zZmt2C+HiBT7PZqZkSxTDUAK35Thz+rrqJ5JHUpsMyhHRsjdLXSC+X4nt0sLfWOFWPhmSIPa9
RSxOrTw2KOeRQFRLMpuFX0UKOOat2GGhhE2td98u3TiXcMAUNLWhGmZa8kHgVUngQ8k02iHuYtPh
9/URl+p7CP7JgTy5bxiyfXgxV9ni6P7FlTmw0tlrf3Gu80wodG8E2nea9wQ9zSOO8ie0iE+8MlQb
KId1jaGt5gYceIFX3g4vlsTxQiYHxSC9qz6dKXgHRLayJBZpYXMQuqXzfSU1WvycTTkSx55hjs5x
OUtAY50iMAViGORwuu/oc1NfUBolwhOIMd3W+8iU5PKbPTAgcrtlnQvmoFFW7kRr3yjV+NXwoIFG
nHVlh5RKdg0JxkFCYv8DQccVg67Jt2oncLNtRac1Cmv1A1EknpW1F4BjpgiuGqp1HImdfPwC1MqW
SKIwYNato40U+4GOopA88LwocUEOUsVs1Mc1uSMNNsQfRNS7fwgvH2GJfTB6HgE302fwxkNv5oMk
fERvFDQ47NF9cs3WOGxJivWVnussELGat4rBeoACE3gQC0bQzW3Lt6RK2jt1TPFVH9+B2JV4epF/
kV6/KUF96yA7q/UX13GxxSLUnUn6Umrx0jWuqV2K3q/508z0rG1ypS60cf64EVblTVOFzbJhuZO4
D9DaZyxlQ9EJIh/KQl/L9U3As0MK89uAL0cxYXRmHAaVwzs+fk1D4ld/FoZC5yC2oUaax+KnV4jx
Ogc5JCKhWwiN0OslTJEBAjrvLfb/v/3auhuQgF5FNhbmr7S7wS3rWPzmvCv39tVKUNxl2DlnpG5r
T3oeNmGxpPAS6rZpFHaaraisxcPERjLXy0Nr2vjtaIVMDT4YG0Ovfx83TnhxUpsrks06lyofvdgN
X8HR0BTns6dFm+cVE6gzDHnjPAf+y0VPevb8S6W88M/dUGIx6Bxb9EGFGlQ+l/l1Fz79iXJJf1iN
KfBNmj9fKtg7GnFb/66csly3O2msxWgP2YsGckvC5hUsoGZ97JiLuD7qfoPHCD0yqAO/P9Abbtom
GvuADq8lWBC6za9hNRv/NkOqiMQjq5gmNJ8I5ZC6vuW50hVebf1dHPtjE8KoH/A2k1kHilgZ/a9/
02Gw8kuJd0m/tNTJ6lfOo20zG0C9D3QNSnotDpr4gfVAkLSkLyHybPNDTSE81dyfkTMNsLToPjBD
bmQP5+9F/HfhamAczfrNeavwIXhx/X6jPsQXBCY9nYrqEC8xTLBlhbNhBIlmzyv2tQBeBO8zUDAO
aUWxYSxNpDmzPWcCMNpnVgi5jOrBYUefdpm/LBT/tq/vEGqIOCe7kuzig0bUshwkFMhp4liA51aA
gFRnVbDnRE3MWlZjWR5n3/1TUpetWqFDAqscvM0j8MbiADkwyWV/aCoRsHVo8km53rRZqlKKy6zr
RwGlFNwevWbROs+Iz26gZJnCL8C9aj3pCQgbC+ZqNC5ZNnXh8mgtFYUW56am6JsfhyFAl2o/Oyyc
4Y8IaQX8THhi546RkjpNRk1WTDILNQY+9/eX5Up01nVmZu2yYO7jt6Mrpf46x331DqHZQLkfxGxH
WZzHVDoChlrFKSUuAUIwh9KQ2Dkz/NdlsgvttTMBwwK2JBvPvhTrR9tF8l8shzvawsrydasZzxO4
Ere5+DeAsI+MTz0R9mM9cx0XUJSKXdQd0JRkdYRWnFmCvX7keDdpT72/eMuNkErROYFmq0fUnF6W
qvd6tKYT8hEU3QjpfavlSmULWxDtTjE6dNJ1H4Bg2TvG6zB4lUdrAR/J7c+BmQWHRqQ4ggq2v+X8
PD6DEGHMSMK7vp+Z/ClEAkOG96u4K9s8Fmr443e3/V5IbsII0B/kHvUuKoDYRZ7AsmOGQLOswZVo
uZmvVHjmHUkjuXDbYhF+YA8S4mYo62Ul4HIdqfrnDxjVmWq2sDZn85EcxNO1e0S84RrJnDp5s4Ho
IhQCnx6FyGY+dAbcQJD1GIAycvpGobpBHxDTeoynXteoeR1IZdbiqHbtlEovM6e2VXtQuphgSqI+
dZzMm4s7muuh4FKo2Mw41LLwuKEm/6SLFT2mP0A8KJpBt1K0D5iiYuk7H1NGLzHFaNGLYQ/+Uv+T
tTJIlY4EfcdRybld61r4Q/mjuKCkWP2xfTQgy4+l011Z70s5NqvFr/9c619eD1TJK7FGQ1qe/s5d
0e2S3U5sWacWboHGXj4IEwNVKMMdr9xKQaAq94VqJE+s03IWIiQaRTSXLlcI/5h6jLXdLjg32L0t
/U2dcR48DWbqVMsP2y9UHpE/1GHU0/W9nN6yDy5V4iS2bQh/ltLHV9a5jxXkiumvQUjyd7JUxDyj
XZ3TCevIJMQpYRXQVq8WJS2worLqetiy/2pLxAG64Z2HGSkfo7e4aPocfuWAIb0nfsMjESsr4Jxn
HYn36W1BW9+rSpH0ti0euHhRGKB6rPHfZwrKF4Aq2X+loNn1YScVekvGUQpXkdNb0I9SvDL56dyT
usoYzOpWA49w2rlaUskIXVhedz1k0oBNd6dFpQqaLcyi18zdjGBW8vlYDAxYQhPaPuD8GmMFHDDi
6yxtJPJbnJi2MTxgqoO0QsghKZUG/ns/TFHi40XFuozEURkx607/2KvvlddcUnOY71QW+kHb5ExY
AoMb2r7J9kaV+txUZsahpjko9/DA/RWQQmVx9VBNxVPKtcMuOBYFoVxPf5lB8xfla0eowF6ggHUo
GuhpEYw3TP+FI7/FtsxG3j+p0PhcEKIHHUC4VICLKvjPYtZt0/ftnKbNomKkNRcmRPjHQiUkiZZb
fxLHcButDrdZ6vfr0db5EX2HebJR9wA9yuF7RQG8cubkyhzCQQlWziszhKX/rLAX+I/Al+EgZvaC
KmJXmkloDcnEs04+k6xQSfDr9ntKu1qyivId1qII1kqhnppSAhx51jk0sKxto/vt3JIs3q7Hmhfu
Os3jVq/HxbAvZVYry2ewwcbHLmpa2LU99GXI6CTKPO3OvItmQ7NHror4M60CcFS0AYaOogoA+n5D
Ber3k9kBq9EDXABfBAWvKz9z0a1VSQq5/kE8KPZXtlGQiShvwvai/4Wcu8rJNxnFzPrK9cHx0msa
psMwmOUw4i4Kz1toP2TX4DIdS5lPbxG+XlXVOsfuLnkLsiovVNU/T38gDtFWLj2JnB5QjGIBNNU0
sbyzsvG9OdU6lLJJPH4y5Kz7z45a9YCwndouIqyhajy+B+S5D8XCm3WyzbLl18JBqylSJwHaCp3i
Jt07DB10s/iLuzvvlC4W+lUhmhxqukBjMWJlMPmZZdsmySb2qNfxMmqMwMbUsmPBYTLMjTKqvse7
DbT3bMJ68EVWXQrRnNharEYIWv7FrTX37pMMuvbU2wbjTnRKN1nFOnRDx0AcTbfFcCslTFsNLL00
J2MV9+/25Bnrfn7EXr2gG7VaX0k2itDgsGRcTxsyvy98fn06uOyyXSrmCNc+9EiB4jic/aLF3Oiz
O6C4NlKjGO6WgwyxAkJg6K6zIDOAFdrOcCMLKn9qauxHE1vRNn5+YXpWoQFy0C0Iv7Sobjy4/3Op
Ec2ClRpdFgR9lFWU3PoM6r00+yMl7nSt4BJRpXUug25yPur/P80sYmEfoWXCEUXQCZatVPO6RNeh
o/+HU8Y5CZ2k+azRNKRurQ+7ozeXeUHQZIYgKNUHTZfPk1mt/xWNuxNGok2luEyTtwY+2Qzn7CIw
LymBFepr1xdbLbhAbeYjVJGMYp8M95LvVjhwVDoq0hph7+ePNnH2MLCwAQtjRiaecvhhqdwGW5Cs
JecWcu+ydo8Hl0Wg6b3gPVpb6PyGUGUAoy4PJ6NKzghqxLlpH4nk1jk6MnYrV4drHa8F+wr0a2MC
Djg3bdVFHcJnungcxcdQtpgreOpMbUFM6Wxh5qzjtoY+XtzTeIRuifsAPrmXYeJQ8q42e0abA2FZ
aV59KlLLtEoZ3goqo9BNhaPJvyJo/RZQsvf2Ammj/cHPMt5PJhbkcFDg2QehzpltZ/zeFSRjvgxb
dJcwzA9Hv7AIztbnLQ/Q4G6UknYtbe3xdTHqhMSNS6nVcVpWp5w+yO5uoAeFpH6efha5caKSg10w
jD34tB2kIPeEQ5h8Sbcg88TnYgFY940Ddn0KlYo4gGUkPDqxf8OQWsO71RO0bwEojektfxwgmR17
UzlTsrk/MXw6OY6BZV7+2mE5H05AwOI0Eprr2SQbdrOODHxgnOkoFJc4+BTSvyljiR+1mIPm68pi
fpFFyBWNVbTcBnv1ycAPBSpWd3mZ5gYkhrms3EdrVhPaj3B8MYN0rdbKWmr4VXllyWmvObuisrsW
YXMyLMYmWQeVpj8J8XrdZopKVDnwdwZz0ibpNtNi5tX2NvKLAnMcfB7pv+YFDkq2T+3eRD8wHPp8
ixi1R8fm2lnWlYz12mjwIsmsk9EuG6Wuky5NYQbhZCfJ/9bEElmT4uEiz+Ew4hEig929m6D5oF3b
kUi3VPj3pBT7ApU01H7vzlUENKeuzFaJZEhDPrhYMXWbKILr6eA7OKTY7Z/Z76r4A9cue2sj76Yq
osNJXAIRImm2JFqIeuyhNkw50Gsti3fS0SjXihQNQKU7+xeU69qMCdSZCZbizdmeS+FV3FbLZl8y
1TTClsGl7Vqeri9y8kCQpywbdSwJmIzLEggFpLl8vKuUYcwSdGcg5+XmMrpsSbXdUZvhPxpCw2jx
8SVymw4Z0KQGSrvHunde5rILUyVIZ7JaLgutO3zNz+MeFUnG4TwTpjlts/RWGrlVbQjPffa3C8ds
X1JX7JCGk6oYSafsCL2jo0bBP1AKWgK8ql40dZL1bO7snO+xc1Ab2ixIKcjHxoseOoq0hz6VuhPx
FgQVzte6AI+e9D+/55HxSsUPrwFXPW2x67LDq02k2H9M5pmSP6JqUSISEh+B/PU7i+EL0+UeUsrq
HLZozGFexIfE1UEZ7NeDCEB+iqTWWNExFZGo+WKPzoUp2Kfn16V4fPd8bSqGUE+JYk+VJAeYAJvU
2Xbww+x8pXaWWRFIALSvnypkJCaTPsvtkg6z33PQbeBJUE3Z6a/P89hq2v/UBjABzneuLuZ6Nk1G
ApVarI4zu/8usVdCp91DVs8/q8cnNovNAj7OJD0BTmqnoZT5BEkjnfgU5VarRH7oCaqsO7LVZGtB
amS94o1CzjCr7/TyXdpDYPEa99yS3BZ5L+Z2HKuUkvMitYNlsSJM/lcV1yGE9ctnTr5kBbzmRy5W
6nxELqROn1PUWUWSCLZz94ls8DMp/6GNVg1VQONG+bfBR6PXqn+cLlmtvD7qjlGmVhmuWQaIKAH0
cqsznPAhTf5J66xFKeuUFplCIWpipsj8bYGmgl143BV6VLJYpwd05A9IFg0vCN8MuzDGw8QI1ffD
Tf9Z1noC4bh0iq7DSUcESnHbRNanGrierI0lagHKOndldVcUU7oFCJ7VBoBNrfLUCGMtmN0Wqmzj
xzALdUg/jBX+Bs3XrDCCYeU9qdHHxkS7o9usWDubTDnyqWs6SFCnn704uLAJ0eZ4EBBZp84xdFs2
gfZXy3khsN7kyIQI+fyPIKXbEqP0F/kW7UIzwkbri4JyPnT8o7Pf+oVPAX8Y2IK+kiv8b6j2vy7i
hz7CS1arnO0tN9YRtBo9l/OFIFff2D/MIF3jrOQ6fm1hvOpo8W5inYlDPfqASa6w/P9qOB9dOKiA
enTFACCe9OoFvZCkPwHfRMrk/oHJOBt5uO1+xkShCxVeADN+DZCQYscb/DE0bMii69QxHC8E/kqt
YMzq/sQimSNRg2rTCwUjDmdGDJ2O1Uq3746OUQ6udxvVEVUSmFIelLhacXFteQPEsMYi0PFCpEuS
YsnqjtsB6YcaEa6p8kJVl9Pcv44SHplSNVbaO2VKCpubz0lS0OjGjywpwVyWLXHJ8DA1fZ/4Eykw
8ADw4Py/+NhN2I3twyEeQHY1CQh6KvQVGp5GGa7JHRXEH6rOR2GtjFcJH2mR0sXYV5rgReBanN0k
A2cYL6nKtnHyBIjz8EqQ3UEjkhbZKbM69jWEMqX/mKrH0/TFI72zMeRGIjrBXnnlLxbgMAe/e3rK
Y8l1vVk04g/TfMJFF/GfHLRarf23lS6pdRIiKgHBvGP7f78gPea6JdJ4X8+VpovAf9xfsOHbPpM6
oSw/qJiRU0BWAvFmkdC60wktQV6TlWyi01vBq4pMp0vIik4VwjFsQ6Ckm3xdQeMHOdGXwp/Ns33h
Rqn41jB4KORklNDzZoKAJUBM+P/vTh1RvZ+wP9kO2BNZAn/z3QGIdPCCS4HB3+xATaKkXsdPhUxl
fgpD2xvyO9CpU/hoJcYADiMMtq3deg4IGV/30Y0TvDELn5Dgl5scGb1qqsHkmnBrQzkGiLQPm6ko
2FBzp20L/gSHAnBeVtQw88fAm/9zKKmUDJ1NJ+BdyzpRNCfXLqYA2BpTLMz1HZp05WoaEyZughGA
VX4tkKFUesP8OvCW9NdwEZHdR2VvecwbTLJ4vO5vOmWfKmqObhZ1Wq11ULrJ2cpxHnm3729Myhb9
n+ZSaJtBo1pbvebniRsY4/PUsmHIzbGgR1vSsaIPgZr3++5/XZenaxhQpEWgnvkEjwSDzhdkQ3LU
T0VZkL5vlG/1D4SeKrD6n4SINRMzppeO+YWUH9bpASm3l3dkY0Uqxh9FtcpcKBDN9F1W2DUCcsCy
UPBHcFAlw2fIp9D7Nlj7e1/nbd4qqiVbN3kLFaaEXDz4xxfhxQnCk3MZ5GPnfG+GNY1aRsLwb1t3
zTjSrEJu5fkhAXSKeCHJK2G8Rs6bODnDv4zazrZhTe4DkNf31QxWHkCfABvdebkveKZuT+1ABqxF
nnx5ODd66176/aOEhIh2QMZoJ0j+8ReY3yKMDyIyZeeY1R0xzH6BYgUy62OYDUn2FU9EuzB4jiyi
mXPxa48IV6UnEZZSMACV6N3crhwXx3W10SoFJQCIL39L+qaIEbXJIkMKLqnawLl1jlVzZM4IeqxY
YmFkz5sl2gGx2EiuJ2NMiiPjkqPC2CiVamYDUF7TeqRctXE1fhJDcSWKkNzIEGalU+iLd+YgDyRc
qMMS1pKwuDGL765KNZ5VkZMt3hwLRWKDVDM7wHorhNzaPxLlz8fn2s5qr9OmmKY5zrpBapZX7BKr
DdB7T349t38b07cvl9FxqMn+LVwmCZ15Xex1gQpDH7UR2CiE3BXntA11EnJj5pAHAIZBWovGzZtg
GsuFuO6ndFvN282du2+fdPLWACYpLvthf9Xftb0h3MRXb1kKjZmpjnSCLLlN8QyexILPLpvCoDmx
CUPqqjf+trvUJaG5u1v2pgJNlGD0j4P/7WpfETahNS8RhKrKbgNcFs9qb63tzXM9dXM19T2g/3D6
uiVeXzC9jgbTgSs7WbxU8zkGO0MLK6CKFHZkF/GJ+tyzUsw26Ga99JZCekMRnYLryYhbc0n33oyq
y+z3AbLdJXQtA399djc3KQ6iUR+SuGGtGneUD9RN//NX2nWgGlXR/OwxV2/G05naf19kM0Bv0jip
H1QGKFKyZ3ame3TAdHrbulvbpvqQMGEDZE9quMBBPOAxHqOnrw2kkJAFv01czGgbGaJhD0pSULZ3
iPCk+N47o6z0KrtjoBF3gCgiKR9wf1mmkZC3Auq4Nna1QJLvsV5XYOKBBvpiWI8NqDHHCF24oCC+
uxyCqriRW8D6J3SC5VvRYWaSkVncz2pyZcNazYm97k8d2i842WrHIdXWTEZsJ6chaV/PlA6Ioh3i
vIpYGAP2PA17rZbXWe2htgoDtYbK1uVp2OdMzLe+PJyAXXZl3C4BDvDaFwya87TW9TcZGCkkK2fz
FFnXuxTUggJHUMWrp8i7Z7AKdahc+xv2pJVktSlIdUIuCw6Ddhbs6P328g/AK7fgp9ynSqS4IPLg
tfILylHBcAFxjCLAtA3JLz3O5PGbISvj/ca4he2B60ADaqi6z2NNbEvEGSj1eHFiL0jPvGhqXsah
C0uKUL7dzNrfxwDq/tBOehq3ADhloUYwVrxTSTNo0ZK/aBWadCKh0vL5o41iL9IBf0n6XG2kEjIG
Aq4219pUZ1aXzFXl580RJZxi6AhhgToG91Qj/Rd9xFqfxc3+J6CdP5MT6cEd/Olmv7otR7zanJE+
UX0oanjGO15XuyZw2BEcb9TXzgT0i+7+xT10GxILtOs2ad2DD6CPsFVMWPM3e60MFrc18tMppklp
85C86PyKXhWtjsdxWE1dI4BCZmPJ9eydKFUMS7QGzviTmhXrbkq2h/oHrSy8EgY9D7iJnqkN1up6
vjo3LmH5I3Ho11NpG8WwDTSStxE++Uawy26h6+Yxx6WzpqHS2bQD/BnhMh7l1lwj4znT14LwN+L6
tcmrDwrdKsiHHxjoOAv5XOye6D8C851Uz3gobJWU7eEPkRP2ikAhmN5XySDno3zD3k88XoOjgJ3m
U2Bvximj4Mwbh6suna+XSvgtcZnP3fXNCxvYkkOY7I3HjMkh/rmWPARb6+Y+jUmBIO5hox8zudCp
cHk6RVOP4YwvTofKi1nic/zEPYnvs+k0EHQ7gyjH61mXuoielRPre0POkvENqJHH1ZVhyxvHVb6u
Y5errwzuh5tdMqJH/zDIyVGKJJuwluF/KLYfdMb/T+ofHjQLdo56g6+YmcZTbgKLuB2JcKTn7x+A
sbA7wQzwOOuRcA9l0NmqKGlnkjfUSsEW5+wDXyXbSIwOH3eqETbsusUAaT/u2b6JV7jDE5L9n32/
dmcSDt5MV0+dMS6XWg4j7RN2byDh8ymVbpcczULOCWwr2KJooNTJCIUa94ufKlEjuQhys6oa6f5c
Zj1BEwtqRQRQPT3Pw+Zt11fDzhkB7L7Kxhh3mRAsWcm0w4d2a5bk/ti0tJK7ZXdQocOBcSjXfGol
PGttiCEwdENVygzWMXsfehmAOwUaEtfSVJ2KyjCZYHJ0KzVJ8pUa1nJGBxv4NEGTjuJDEkxyYX67
LYIqgm+q+rquoCEZdaaJ7ITzbIus33TfoJJyIUrXpWd90mDD7DFEVVJTeISNGdU0Eot0wavUY7l6
V8tgTPkvscHMVGqM5pT0r4Nda1IFAXsOPnwc09GOTUpnr4wt+R3hhB5wuFR2pablHr/MtztyX6JM
FFbmYmm/6GkalfGbm9Bdsl8/PUxlSA3wSP9G7lpi3w/xOfrSvvNtaIcDNyyAiCtWT0Ocftiy/LLz
b7cIBrgsFhkqGxYXvSO+1DEkqpxCyMKXnn9Dmnd0f9JyhnAdBmqPUXI7QNw6EKnlbqlx43J8nz2S
pMEPR3qoCz4AvS6Iwhxlwo44JV8vwY3eZ0GyiMeE/zrPl4C8wS/YLAYMbQYmPqcI01qMM1TbQUND
FXMw0R4euUFjgO7So3rFDyHwGbM996KSxT1GheUuJHgkZZeeq9IiJjeDYOQYJe4cay0Qj5ymY5qh
dvrNX7hvY3/O995MT2X2Wu9qXljEw9GQmE+KcVLMXH9HYeEv2J4Yvr55IrCw4Z26j3xplYIOY1tE
95JMP1y43raYEP8yeV+1wzn09RLFdzzwSAmoFb8LnniQtZisBdNb+fc7CP1TbPdaiTg7eyF6SvdU
yOq3KurlUCGLWU4jU1MNhiMpoSsmI3DsF2L1wV+NFB6auCoYDTLHvu1xn1nCvlQ10ODArIbm6Ukn
Wv3RLf96yuQ1X+wn1LTT5aUrgxnltg8tsmhkdT4ZlGQx0KvdUYqZGCajbWU1wGdn3HqYWbkjmw5h
4BVN+SEM7YC9Q6Mo61qqU80Rz2eIo8i5MGlnY8F8Y0Iz12IjYnL/fPSJ9v0rziFAugUwWp+6GHd0
ZNPQqrZ80sNLpA2+96xlKrTQmMsC0WlAu3dY7vIk+llpbLsV6TJ0CTJxM9fBWK1D6i5sxRkS+9o3
OB2C34rEE2yPAZ9i+oAtdRqaqICrBkAn4Y57STvETe1iUC0m4GMjmfMDUDbW4h6EIYg1lfAOw2wn
tPvcJxZFSL0GbP7wgfhHOI1wqpoF9hAbDNxGrvos5By5xEx/eBeuG/hCYg23tjI0HTa5sJ3Z0MkM
kZokjfUA9RoD/EFjoD3gNUoE1fyfUC9Zf0kuFTQ6hD/nFz1tKxWbck83/j4Zv1+CfW3zLSSoOtNv
z1ddNXfOEVHcnuUShmcmC3Py64Ui8IrJD5AVRqKh6mdcYyS55CaK64vu4uIhfM2PkPgpILXkZyTj
11O88TIzH1XJsrhm1TbYGOh2g/XZQbKvDY0+aHER3wo7RCzDuAf+WBgnpI5vuU9zIMeg21f9SXhG
W84nV7JoB3jaL2Xdm2WM5skFq52ikjrfhpboaIZzQOcGMeRk1X7++hZza+etn9431NUcuwLLcy5R
3FpcnyKm3k0ddsTFksxPrY/W6qbxmeHarYxbRjgh2MCRN8VXcbX0+LHdRPahSllr7QUDUIK1eYYl
h59vvGJxNW0qXyDbYaHq3KgOZTdpk+iFn0mjG5Cv8R+UKup1PZXeeDDDkgJ3UImMum7Ci15zwH0o
KX4MhVDJoJQl5rS/NgtNz+PTdwhZCsxnOhi/4GoD5BoJw8OTW7ntdDpvpOeZ3j3xcUCg9JUNYUrY
mDyu7+fgMCYQ4M5tr2lguA0NTZeHAft0dKgGW7pwV0myOA4bukZQGgp3bXmQscyawKmmjU4zcveH
KyvoI3/xZBbes4V8jfiRnHRKfKtPZNyJCaR48g4Xkaw53fb2e9ErxtME88DQTLE6p9pt9Ow2LxqC
VVvw8XWKqoyqfwylQZFICLuaCXrq/qWFocl/g/C22btLaSmtWBB6syo3EMUHZj1ve7FOyMlTFyB5
JMKac9W0ilfreTBrkngq00ncUFTedU2mekMDrqdrw1LxfPKKaWwomIPOLnPShtlMx6IUqFOcLpA3
xn9A9y8MdCbS+wEK+5UM+tqlgkYCMJxlc9V/iUWCbaiMm/0fSRMIx7w94vmDyi93xQMpWsoSoIY7
7oz+zsOdiTeoVEGZhXx2pLwGZl4j3XCmc7CXjIIT14cb/h1vNtUHO2zfEWp9uNJySHajaVzy/lNO
UQ0V3JbF4n5acD/SyWkQ86wfRhyYr74HofT7I0tGwkCm5PiY3nbmlCpbOoTWrSOmmzE0FMzKvNk0
vqnfgbr+M0ykhGFGZa79txq+KmyubUwheKnkAL6VRbh9x2vc9S7xT3QYn/UhK1d1yRtIzeqInkf+
ne/6wQfbW/RGjtI5UaQ0Mo2LLTQWBcCHeovx187DlBqyyDj2USYBE/0/l54eSAwto0SQpEYDz98i
8bP80EMjsttvLYOhBPkeDijhtdP3ADhcfLAH0EqTtjAjZ3jCun4aoo+9Vn/BuoC1WSvwVlA92F7I
Uzr68EMAYamq7XYlXfVZqk0W8HXPIYOH5T65yhnnJhVql4t9Y2e332eUQARP3lK2kjQCC4Wa+6XF
9Cx7fLH5f6JBMuTWOZci+6UtIvYlJ6742ocgDI9acROBZ9EYyIEOLJxg5Tr8cSeO9NALIbylogrR
nyN2mMOh4ohErDfQDBsUfKdVhE/3rW40gnU34q2S+IGZUlLN1b/oIeUqlgfs0bHlj9DNzkxhEQNv
jJ0yehSlWXidtxUSvKMQxTQoMBqPMRh6cicULdT0I6/iSFdV7nMTsQUZwD9z8DJ9tF9loCAITK0i
5kYgkneZQS1TARVEjZRU6+0ECUibb9KESfADOce2xvxcOnFH60dVVoZXBDI0XHFWLhGt6UwYYeNB
eWaKZUAFnAk4FLHR1uzWClnZMla2Hhqi3c9aAp+0LcVOOfNJKHpRrMH1ACTMhEm7oeT9zOLibNSA
09KQFFyC4UK1VMkZeIEhQNfHEZ+R7T2BCo82CeQwjirHyShe2PzZGn8ggNnuBPeAZ7zbNcydpZwh
SJkgrmk105C6w9QgNyiyPRWlsPoou1G9w+M6kgEGyTjQayeQCEClsmDUbjbDh4lYW3ek+Y93D639
RQNBr/7z8HHsdZPJCPPQhwt7aDE94PCbiMjvM1ZUfzcMzK0M4CcFLBZyUp/b302LFUGeYF0NrunG
ekilVqlyEQvmPeZsGH0oXrQ+siDBSu1EdwIyJ73ueSXtgZ6LfAajpiLDW6w0OsVKoBKu+zN3cp1U
qlNb/PJZpxHH4YQcIxpvQf0KHZxJsNnAuNTdQUfWN9kGsc+YssBjgRfR2Ux+NhBmuyhNRBNMAdXN
helMVzcraqj5yv4FNFFgCVFsafij4Nwf9ttw4Uu5SvTdofmqqYMTA0Y5r2jtNYbxgpxUETzWPswO
nXxY4flrUfiNhWsLYX2aCai8MjunIKndeASvP11udO069XuLNw72ctf/2VRL5x9Lp946daevLhZf
AwA24M/QB2hNr59KuDAwb8V4691k3MUDgmkaKgd5OIQrcOTm0eUl1z8tGf8oIUigBhhZhV+MqkIR
B6T1Ok+sX9rmPu8uiFQ3GwA7nOIbcZ+YqDziTP71gQkYu9dJmmxn8wRo5Xel6noehQDK3tEjDgxm
GYuWG855Z9taZVZMne4sHxDsBvCCnMe2W9+vk5fVyB3qlRRwF1aGpwsUtZq09HcrPAaA3uJ5wR12
koLhqlH2QPci/S4Nqat2ruDun2T+RhZWNOmwfCTPepizxJ5lYX0Gx7YrJy1Dh/dwOhtB63Yl4tEo
SwykIiHsnA7xkTgTRGNuW8c5hTy9EivLySxSXWO7PYYW4Z/2zz2Nu39O0H8/aHRt+QD0M6LdZ2+P
+TqDGgljRkzJC8VrjZRRGxg2QnsuTyNOyXd8WYMjuQWuChwtLg1Ba/vxTwi996RIkHGVrX0hOKtR
9g+ZEYYuGjmwTYXQRRfnOq8PnQAq6NYFZifKS/sE5y1cZH311qWJm4RLgZjjQGzZZl8JtZjYd2FW
s6G8PVWp+0hd72P6sbw8HLX8e+Jp2RGSqXVjT6Scz/umQ/xrmNs9JMeQsU1jHZGNX7jO+U9CPpTs
cNDDJ/q38eEq9pUbC+Hqx2cFtYjRmPMogS+5ixwRRgU/eZDXRA+Ob7hQcIwXqU5rnuA+rYBZqmH5
CPHK3jkfAJGa0N86z7YF4LnTBYOr0PMbC/jq2XFWcaFYwdIPf8w4C/e/UaNonUEuZNYUblOTTQHi
WoaJVYt/+4lPPOBcwuQHyBnMnZmyOp5lB3OMNaH9BTV6LgHfj+5XcZinnkjC4AU2ZnuuxtlHy3QC
PdpzL8vawCLV0xtigjo2Yu7GSzL2ls7VAVH/dGniCoIo8B2dTG24dp3YOFNyEPWGCUOrwsCBM0Dp
lJzi/piYXHi8o2y1IcxCk9hJIhCcZon5aUB2QH3xDgiS24uoKme1zYJO1BWj5oCM4khDVDdb7YLt
4XgDhYe8lEBIEIOVsicNiGILJlPP4IWks+dJNlKBCvAvPWnpOLTDZf+teRRYFY3dh8xzhdkWBUGb
m+s7zXJqzIEXa+NRhfPxWZhLxpMJMBE2VrkqVbGRGzdQn7skARVacZ64Tehz8oh4eJTHnJzn7Hbs
2B7YUB5KoN/zCXBAD7S5vvwOx783+NzC8N80VSaznClXhsS8GgeABECHYASuVO4bTpsgPrp50+CR
sI+89KTvUkrG6Prg47JOkZDGvBmKoSnPlXgJbGKJEJG6dSQ2aoiRjW2vobSTI32Xf3HU6MrQyzPb
GdVYZFZsRetVou0qSHyN8G05STW3rJih6mX6yxGbjjBQ8XJyec2xGzh+unaJXncXj/pHfqDJLSqG
HJFuJi2cEEoQF3GHjBTrgOHD48nAQlmRCMVuPM5HFJkfCRVMZIOIvCZQSn4T4JgJz1elhpwJva4h
RtgMiexVLyO9kQx/ZVXB3u3HReFIfqPuNls4IKTqtC0z+NiEGz38BYlfLMkrFUjDrue/LJsd0Uw7
Ik1ptf7zqdfluNCJaMC9tWxeror7vJGAfEj/+zCxCR/GjJJpBJnBOCVP8d5TF6jhyEvxzKoCxmJ3
lTGRU0GGalVI52ACSCe4RpoQLdittcU+5WxtqFrTLlvtXGGX7yrWm1jlVeTNWQfs2pcTjVeF/PdS
Wi7P7I3DHSa2LBEQU/QCFruffMSSieTN2MVJxcsipqWO5xSSmt+lJJF7hmaZX1TbpJC7+hD0uEMk
swZdmSH3U7B+zNiEIzGw+X3K2K4q6D+ao0X/hoaj5FbclhKg5kLLZCwOjEX5/mjrGkazSvoaYVEu
/5qoCI3Saip6Dxxj+flwOhUIKulAQd2E0yHVOpqCB42lt5YhFznGXu44bmjR4JMcmALeSq8RyRP/
3yjb2cAyjpk+tN57yCl/kLFLrI+/G3RcTUJhtPdjjXvur3lqBbrh3QrpBl4NENwu9lijRzzanQjP
TOC6qT0Le1339LnOeKni3LYdIuJCkUp61oP8ABUZ17dlSSrinCzqwyMvDqtd/Bq1GZ0svMjiarNX
19+XqjPkDKAs0/Ri6gz2dwNROti9Sf73Ei4xub938r6zcS2K8Iq5B7D01J5Sdu4Ca0A9nIzjMv0o
3FTMgrPhgeAcf1Gg2SV4/joXmDX2OKDWlvpqw8MaXqQkTB5xiwPWusncRcMcZ/fB4QpOZ7zLymb4
m60QoGYEJqbUIrDiuc0+b/OwqUazLXDWFu4Bwx1IGdyRLGYx0+9EtrhIONeKWCoWbosa1h/XaILw
/MHE4hwN0o2cNOV1PbzOcoA3/Xa4wz/VbmdGqQ6hlqeqigUknnqq8E4AgR3LvcpJLnukO52UqoZW
c1B68iTmRphhrLao4yg0NOFCFV0PK+xE3DjV5OSxwHo3+piZaCyeUJ+iAxAv8OuLXBbgwBnUHoQU
Mxz+P74PYwrXMUGHYTYhLb0CWbP1l4o7h0TOpLOprzQM2E8zGstcFhk1aFSQqYRAZdiLYlt3oLKD
M8dXy9gxR3zWgXDrodsmFoGR1V4xdiuWSHYbMGJ8kvm9tXzI1UeV+OBuNR9RydTuUrlHTI2JdEv8
KLAmHsme0tmPQS1wI5lgNg3CrHkaTzIkxEiLIG/6blPari+u3mS3CTFS/brFCJwyOUOc7gsX/biF
ox1ByTUsMDk+ooH9rklnVocMZJBiYbfPqH69BKQGHjidcazsxgyaVI5+4uRKCxDmCLAvQfi6Anc1
GxyCF+FXHsZuuyaQ/Qdk/5df/9Alcxwokv6rscfm2q7ZXZiaBaHmhtO/9LVY0gDrnZ/KgpfTqPmh
+B6tKhty1wx8yWpUgBP92uE0QVJlsGs+++/H6SN6ICCAoEXKep8Icdh13EnfjLY19iiyi2363X99
bA+bOZLnv/SbyWML35o4FwS63kixDtdMNTl5s4B5LgPBRrQxexN+yAF110Yc56n4YeumLMIiQTgz
cQHzcGZVr40/q2gf42t7ypkCd3/L2JkspDOe6ulsZSqNHVPDRVHR8l7J/FpeXaExeMViLpn/N96q
jEhA049l7Oxx4+wgGmSGwfpINspBo7ABJQdbsVOudduAt65vmjYXEZIqiu3PHBmef8RtrazJZJOP
y7ejUAIqCU8XfJW3QXWwu/FWIrxUmdjenwftR6VhJ1dFBALbkq4ot7n0OkC96q69N7L73F+1QJhR
/kEsXudnRC5rJICvsrmpXYrmgHzVyQhQlFYad5Fo2j3Mu2q7O2eyQlFkdl1rDy4BLWVWFE3E0Zf/
uyJRFyYsqHW6x1coZ12rejlQlQy2kzwo2octgxb6rJ+eOFg+8luNrTkw2obHkWM11ZIggqcfU5Eq
jV1asPDjPy5+8Ul609O0DeXEaC9GFEcXsuQ4/EHQgrD0QUapNr31VjojO19CBlI0Y7Bn34cZ34xu
8EDG8jfrz2QrNBBSMMSMT5nUg5D0lCtKpCF8hN/24xx/vk7gMJfByttXnxcfQTvMmNQdjbur4vrs
Sg6lWl1vnjZk2uJNQYSPiumitHo7GDXZfvhYqaKisg+LO+UrRsGUhwLEV7mMi4gyRIP98TSr5yj/
n8vmhIUojtnl5lh3nrmcXXFaC27Jbhl8uaO+zIM0GGm8P3mLp3oT0Y53tt7AYcYxFbOGaa5hdoYs
Iixz01I8vKrmSzhVZauxZjCdfMXDC+arI41YNtEh2Xq8UiL7H6YplTHD1UA71gBKmaZAEVHMX6LE
My/qttUa4ibi+1E3K246bPMG7nlO1Ixd+UI4N06IamZPeYUemAuB3SoeZ2mYZuVyFGoEmck3mWsR
5ca+CqOSi1Yfkarqg2V+Zk7a1OwIo2+YYNSsuNd3j3r4DTbvRIzmSiLUgtRPPZTq8VbXkkfjnFqm
LJLaPSC1xSQW5CnACu7L8KaAW8tAhaSRksA1V5GNQB5NH6WzUUCjtk2+nH/szFP1tcFghIKoQg/Q
zgYjXKDeUGUtDpBWUD25HkbK1yLwV0vlGHcl3+jgNUwvHZxKu7n2qu31t/Casv0K2B+N6tnbTdka
sR35gZCIKMLSVNhMsvbyHwe+MYC9g1Ug36T/YJZGCdib00+WIAwQOiUHrWMIJYsqn7D13gi/UWhL
HlN5iEw9Dxn5Ld1U/uiIq+ryN557SP68n/Sk9bfenZhSpzehipbCH0Q5WbtNwGfoWS0dj09xfa/6
C5z6Ml1B/A5UP+q7a1ba/5jQ9B1txrh/jseICxMMCmiD7hflAh7yQSmuW6RC5qmFQBBJcnRxPkzp
vN7eTQZAIfFWfXfvW7S8KTUjexCk2B6yYXfud521ISVjro3TRxqxnrLboDX65fVBtEitkxQd4Jxa
nAp3lOAVo1NePkRXCGI9e8NXhs0uCEOLDa6eHCupdG00BdFPSsB3VaHgqZCod1W3Lq2e9qpAm+XH
bhRuc1fHalt7L6TGr3/FNQ+CyiuhARBkHoYVwcCEMsMPDIGDz9VsjS0YCoPnGeGjs6C8kWWwydSH
KYmtiJnwLRPE4WF0W6bYsZBSOUOM/jiCkUjjebQdZ/v4vY1ezgM/qFLrd7tWU/rY19URDohazuG6
yQ1XilTc8/9kKZnK+Q7cvXddIyE5Cgt/eX6C3feeEuuh++S3wqxpkhumjtokBSm5+H6jzjUHmWXC
DyL3NIjlCWnOxOrkdGlZhuAFlrAOrgS6zKVPY/fe4C9CriHkoXjDzmz64WwL8qfQLNXMzzHMwdrM
JfUOROPOAhqB2o20uUW5JkJ7upEwPKbfVhgf7V6uSYdTG8ElTB9LzR9aZwr9yoAH8L6gc+SCWKnt
7KWrIj8L5PfakTKtK3gVuzggzLTEEgqHqf9JmvXBv4wiZZTxhFXqoVOX8B70AR9S2dyN6++Yb1VP
A9WBiyrM7gmKKVSZcH+KIXe8ej4EXAMaQ+XB2RgQGwB78c4YnjbgrrsDrJ5k6xZTbg4l0MFB9URo
GdxJU8Fc5eMI++Y2NQppKl0/EEpVF96SGYx1viUB79G6XnVP15w9Osp/LjndwcJPUsxXfZ8V9ZVe
WprXxwNPUAXtT1B+93NMnvr/2Q4ygmrFyp+/snrr/NlZhkBLQTpFt7oWaLxBkpUM5YfYex4HVb5P
jtVZOhwX2YrJiwduH2y5CO123r5ADE/1IkXBNYHR07Za7/Ytt430oENiRAF8Bh/hAXybE3Wl9Bmn
4MuWnkjeNW/BzjsnyHjbnYMzLf8MVZ6wjBEgeJT3zaTmgcPIs7YaOdKRBL/Q3Ehhm5nuaYt2Jv7Y
/Ana/GQqPa/GuLeB0/a3GdsNEpDuKMiWxk7sUPGEvsK6Jz3OXMl8J7O9p595C53pNFzwe+4LdFJC
2dVV9k3mNTgm5lEc9eE1jeddAn8+qfQOHWeg45De49wI0AdbtMygBd1zA6bTgs+LYBxnm0KHFB1t
ey+LvWzxFXUM8JqdohpE7NCLsjkC+TyNj0Oq/Fau18+VseuCxmQVk2GF92VVKsB8toVj9mOV5Wgq
gflZ8jc/gWlWy/AsQu1yJMEa7mXe8oPJCPkz2kOM2fMpBXhT1d3nYDN8ZHVdbFAE3Qgo32IVAv4F
+f1hUThEfVyIOk18k3xq0fPDrkB+sTEK9F6zzE6d5PD2ODLJpG1Xd/7+9Nd+FDLo/JCQmkCdxbXN
faIpQOfry1IBIqfRdhRXNgx93GI31lbDF5lId7edZ7kfoPLhR53Es6ssoxliKT69WKhkw18VD/fG
GNCHbjr1vfPqR0jOgIPgzh0KM74RpQGRB1tmvYkrKXtOxMZ/Td109L/v6UbktonAU06/Eu5dqvHr
Q+resIPtOvjVj6GksgPz3zJEK9JYyMduTtyATrVfI30Yo6yySABlHJEe/ECf0rgr5Udk/4mocoph
gKcmGQTCkmzzDiQN3wRTxrdIQMCp551aBqYUHA+nRBp931HQjVqWvA+iIzomvAtzG6I2RKHUZ9LJ
GgJg/GEYNCAqrndJFCnW6JXfSrXhPBZZ8mlnKZs/ZIUyJ1KSFSQ5fw8SYYTBeNaAY9medheiubos
5gYpqKMZMIy3ftS/+Y8z01eJxyOzKCkvQzPjEmtRnPAw3Vz53vCVLXZcVlEf1yrqW/lZ3+lGJdr9
DaEpNHxc5Bc1EKMjRTW1uNDrSKC2rTDEOjRahj+HDmAiEKyKBcQ6luAM0zYf4A1KMXC47t9uIv9+
95amTC9X0gwk3c85roCqaisyKnkyVxJkQKAliGcJmTHHHUKlVOAXsqoG7jLJZ32/CHXuegYqEbOT
PK9LxuIiWM7D7CvbHUqTj3pfdkcxz4pR8F7O+BkFg0PNAVux+jpSCDfyXH5Vz5z8V5BzdzEqrtk0
TeN74nWuVxZ4iTnFmSAp2Pb9vkcdCoQ2sPXV4UhqO2BqPEpYIRUcWAnMxOOvRDVzaX81obASJ4F3
0qqqL9OT7xQ5pV34YCTRKEU6xSZ8ztme+RgVC3rJnvtA1ZtSCRrDBW5x7LLgrWqRSXVjYVOPBjFd
LwV0kvgX8LML5bG4xMVEG0CODnVvTRh/UWSj+TRo5PC3EZ0vsvHvfK41R4BFo7Y+gnwyaW7sizG3
0XxAz5r/4DuxSDPH9gtQIvS2J0OaDLQZHI8nYj7V9SGf4CZzSn4ttHKNUnbamIZmvk9o6ai0PlLs
3zaX82x3+nZQDx21CWb+YREP4ypRUBYb4BmKFt8RYlZehdbopKx5TEtNgm7VOCbjLozKWA+pr7BD
QrfBo6mFF48O/YBWgbSijxryR3ytYNxxfGZB9wUgaEUIksc7UWKTdw4X3/sPnqac8r6J/YOP/FkN
8Pgl9OeihbfIeLXxr6TcigYS06JKqJyyQS4j1EXHq43C/76+zDzp2Sq/Zc5SFBMedRSsBoFalVDT
HunSltamofLUhiphRgACsR14059ZQvsFy2IL7620Zpg4s2V6XQn2rCQnL/SgNexVJ5tjmKc09B7d
6gSOKL/HNEkFPTZbspPd8adlYk7TMxht0izYSYt0g7cKgKAb6qdPaO33Z1MrUtqTBvDoe9qon0pg
F6go7Et2XamKF93pj0MoQ+kThaeW5CqNalkAUzaVsnXEL7iw+06zIg4PEPm/Qt81ibTkrFIzDofj
4INkfhfItjqiBKalhwqRwEZsqf53C6i74v3x+WjRbcFlc+/bfIki2F2MTwuYvZpeMH0fULlgmYS2
PleLdYuyIjSmKH98T/mt/H45b8bkFaU3RrMNyiyZ73xM49Bfro07GPl3HhXOVB4P0MbqCqBYm3ID
BurzCvh1eJ6oVSJZ6ykkONWdxMjz3JM3U0rGqZGMELElcOz6TsgzYAotqZfaOIetV51rkL7Vg7AR
HWWpVHiopTOA4bD2SY3bxRY5TxZvnP92GeVlOsD4vvPj38H5oL6Yt8N2f1IWPPOmFN6ashdrN43i
9po3sTsOvCgdX2vOlULUcqrGC5dFJd77l3bK6fqOaj6bCoiT43gWJTX5YYWfL69Wa75FyAj8w8Nk
RKDzVVcZb8gTIRMCvhLnfIaW9jS2iFy4PrOlfZ96uYf3hDq51pKEc/9Wm8ZLgRc1uGbU5952Z6pk
Dk2S0qAicMeQJIvj0jopkHs7CxHZCQdZXyZBolGL0KAiKq3VrQDY1+Vu9ay0LbuHpyJrVdzm+IqO
wNbqlo0kGBuZUwT96WcjLeXc6PxY0rE2JFAHJifDlXnddE1o1yyL/FjhajwmjuQHSwrSTb26VHJk
Wu9Er3ijHaAzs5XldeNqsgb3rpZx7155mbVODs3o+iKu4D2q0fOizn7CvhpJEkemqOssnwV5iLR9
YxDqGEhr2AfejfT6tk0AnDAaXDXwA8GmJ4Dt4utDrZIhFnNWxqSx3NmnZDmfox4RBrUzHW+CLSlS
q5f68Skd4XuKda7QZ/H8BwDdiuJvGMsBi6i9UJ0XO86nE33VO3KvsuJYElzVDmLRsaVGKsQOB/1t
hZP6qAdhN0yajUwmuyqULNibk2eySUcw8kd+1XtKT60yLVRm9sTwkrA1NG3xnFCyIeWDxCF49ZMX
PLJLPQkrCMlvB+9h8uX9dqtEaFBJCxPdmfQdcl0gIuf5YBcUSjESEzKgvMoIhs0q1Ln80vvY84/M
+ZP7d49k79QpQZI4w7OTQLX/4aaxomc/Uk2NIFeiVYbpv8YGA6gfzHDeNzCd7ztd4UWhfV+vkUJn
/xHMd/qB6wwXsmVkXilKptOz03P8osNP9uAktR8ZQDWtllbq5rigcf+9oI/lqDaAUATYltO5hUvp
0QbDdWUImaMVqZ19o1OAvyqL+3rzCGE/FH9v+aloAbprUUeQukYnknanA0sbfzcJSFMPVGZJyGTI
pZPm88hZQsLuNfDlr4FkR6cDDMb20/MBDofNOpHsveSAO++ceJH+eEn0JrykLsdwUxxjYfentUpc
Ro6/aSVzVqA6BVsEEPW5NpvHoZwHDYIoZS2oiF1RBVqvKx4ygUIkxy21AxP1JUYngOcNTs8szk5i
tT29UhChzd9esZzLhjVNvZ2CaxSiI4c+wYM47yVkVJDWL1lB6xlGEri686hry2+l3sHlR6nvaTk5
FuId0HDOWS7iXpW0V7qhkxFcj5ky0QvYKg02f4qLGt+dSNiNEk3UmQjcpLo+A8o15KCtPsLNAFv0
wZbArkKxHphJQDelhydw5E9f4mMVB1tGIFf5ahEulH4Kbz7u0hHJ0xwDYsixyQZwMNuHL6TjsQAV
ytFf5b7o+FbOocl2m2C7jwmMfSsARelyHiwssd+QrFvPLFeUnTfR/vomiXk+uQn1UTRleVKUyORt
eqM6NsJrh7j7zYSPV2GamMbp1/IDmTHHgWarxuSwt9iIO24aHbXF+RSoHp+qRcTY1e4PoMmGI/Vw
Uk+XN/9fzPzhj3elHqEZKUPbAnTNJmZR/Kv9b6ayaKN247UkmX2dN67rvvBMNvtgW0eSovR2Mgp6
7FFXKy13FWG0C6IEarWlmAM1Z0RTJljSMf5Aa2UvfLz2RQmlS+A5LAYz1yk6f7BQp5NDMFEta3V8
XKMjxWaVQTDJzl+bWkXLXIW9waTezPOpRGxHu1FF97ar3KCqvh+1hEOgxo0AHeB99kRJ7rEf28B5
bA5pA5R84Whucd1qKhS9UbgIeMYx27BPhFY0ux275hElNLFvOqfov68H+wmxtIleDTjjie+V2DHG
iZJdGZmTvjZxWLTHnGPInCxKlP2B8iCmg7GOW3Hx51UpZwPkdZtO/6xcL0UKlF0cfSlugAYsLHs5
UKzDPI4p5T08cvdB8fPxD1MMocmr2WDAB3PteXX4Z7Gwc7ZtMf3F3kvYjM0BT7y96065xCRKlBhQ
VNpoTdtn6mEm7ErSbMuqjniAsDrzdVduAE8ehteXHXL3aos+qLmQc1zqABv/u59ZvI8cAFBmMjCV
SGrwUsSCK4XDnEWfgD1QaRG0Av5rCHxKyfd1uBU/S8fCUB7oycq/SInvFUUf5RB19oeWIXWtFSiu
33lWpa7IQ60O4QXNrCkDX+e3vWTKEGe5xDPmks6UlOmm4iMtTzb+dABa63UBY63l5mC12Xawpzs4
hw0J0pdCIBKn6R/WORthE+QBACsnggDpzTde8I08ZOlMoLOVdP6KzPFlaNZJq3v2MS/XimKTgVfH
fTxwpdx2bZyzJmNHsAx/Qf4sRzjCMqmLlWEE5mnMU8MkjaifBQxbOgtqWHAjs5Akk5JhGygx741E
OwX+FGZYkdGkyicbKZdzHM0c9xkc2W6RSlnuXPXCqVzyUolmGf4UB5zgG8hTsVgaT3vVEPFv5U3x
BqutCrQ1qzlP3kZpqAXvVhhdkyUvQi/CFHjQW15i1GUmJEXU4hrniZnFDZTNrny8gHYZ3BCJu3/U
XCYh574S6cXkwuRpK2ylEOungwBh+X8XNIvQ4UUdOVoNf6/b+PDsPZ0BsyMQlIgqg+O5a2SMWgg6
DkfmdYJXoBwqV/VgFfa+yQf/D0tA5opLzINzEYNnM/2g0Tve2GXJHrQODNuddk/bsFm5kpOdkEgS
hm3KYQIE9npaqD7F9DFHXkhdZ24/VZbSC3iAUYSz6pxBhG5QSe+Uh81Q6gzqKgg+HFu/NPwNGfTn
y2y6cgY98mPQeZAg+BRx4YkVUsoCc3eUrxcUCnwABh5p7RzSXe3Ay4VnuqKzTHPwa2TL0mAHerwG
Flv1F4iTL+9zx+sOEMyk2X18/pOW/1zYCRNpoq42bhu0K06qHvf9FJYK2J+NTnW0RWA43iEiwbJW
VQPsL0sE9qNAdzHd2OHOvmjCe0h4AOpvPT/K1pUqOeMctxKi8tlEb25OpfZh6FvTQa2ftfuMNqGw
O139Wyr7ADJ6AeVb0L4EDX91p6ToeM9t7uqM/rr1eaL03KAunO5FFht1kcg+7Fr0ciHOP7FNXSjz
s3AIsAEosPwqdk99i/Hwn+I/5vWPE/UzPThluIqKAOU6mB+Ki2yX6EeZuQaFPQ5LD+sSWaGEjalX
VyeNvrutaWLoJCb4e5E5kuhthq1+3OW/MWngD7T8MFj1h9G44Gwtea/UFrJe2BQ6PlZQ7cxiZLqG
a3TaTHIHZnthTVIVfVmk+2fVdBQsIddJeF0bXxaKP8bictkHAmMc8jJnb5JEpmaTBVcvPH9o6cSo
lMoDszcZbmPt+9hCTZ4wANe/ayX26Aa6NGWuXCDrEQsX1OIE7+4WmmTbp8G8BikN1WJkoRHPpjD8
L5GDeLE1aKlmSjqkY0me7fFcLC8VWQDi3otksH2WSCV7mBe9Ub66oCswqapkBVWk7bnb0EDV0wX9
5m5gM/reYc5SKUFsIKlHNnqJSut4aAuntRd5yjkZD/u2ch4KqbJNyht9g1EzpCbLN1rG5itzRLnq
swRKk+yKPyaIdcvGpAvrqY9DqWghDQDYvAg9SmL8PSszMnBTlp3Xkot1PshsdH4S3RER3cBKPpyd
WNh6lvaxqKWts+Ne0hdoyhh3Ibqh4Cj2+uQxSbO1ae52NTyTZoow69RsKAw5v4yDJZn1zu5E1zyg
4aOzxJfMOsrD/huVCQkMICaEhYIgeZtCP9uQCD1tUs4xIhVwI2U3cD8ApOpnlqL7j62omVcdnvRD
fURP+d7MBgah2a3ysTdI7L17NGCqmAOGgu/aKQ2CQbCEWBp0gF+m38p3oMEYwX2LVLayMRkR6TRT
iYVJndY2zPBFhJdgzyG9dN0maheX/w6i/Js2qDGrvSeEUh/ho+xIWLJNrnoVBUapUn37dLEVjhQw
bdgBt1UfbyOyTVpXBDvbbMrAHysIsalM/OmMIz4rrYvj59Hh4e8HQEwmIpA2wCh5CcnOthjQXCdg
kQgbd4e9OEghyNTXP6HAay/e9aCms1yVmqjt40eCMPBxNXI9ckX1HwnqxI/hRhbgrR2JiqES/Bew
c0qRLO9smoSb6I2c0wNVsBYVkJg5tyjYhc3MBg6sdbMOtSGHTDk6UrRekn7ws7G2tfJpYFZz33t+
sY9EGdMTp1PROcGjABpLkgZfJkqHt8p8M3+JBuVJw52Igj45TN5+nj+rmRosGW2gTRq7BWCTM0kl
YlnEZnLPgBVDwJ96IQgEsHZ4+ksv2rHEcG6+9E2eZ8xCbkkBoLykoUBXN5nGqkEfQvJLF/2Agvje
DN1wXxaiVgbJw/APKYu6ouShddksJvTdgUzPej8REKlwv54793M0bUONh9n7suUmqHtjfYSPVa/y
fl01/0L0XI8m0NuH/5P7cShCuGlQgcNIwLkk5w2BcZ18SQEhB0XPTplfLGdK0oWJzdCBRISuBC/B
hPMro/jkSqQxRzIOykmJuJRAXaeYNd8Fp8mrMhiWVREmlpxJ/nxrXIx1zopT0tegV/RAiNwqQCR0
OAv2Sbu6AhcsuPRpQBypOE0xxX/9K0Zb7XUtewxMDknJlYbYao+zYmYETtHDBoLF0iqeA57Yf07m
7etCZcckFbtPTRamjSzEjBLL42j2XTNwpEALFMClioYUT4ct6iazr76RaVeYSoAupV4zYmVH6Lzs
ATuKk4gVCPUzwFEt41P5t0UPuI3rupEvystPxzB/P70HCaHFoBxvGfPiIOfWTsrZ5oURjNzDrb0g
KGlgztjYkHv9MaMEF2O07Zu92ExDWm4rg3K4ju8zx0xmujlQGx7mq8s8/iP0mCH63oD5Rrx+IE5z
IywJnou9i0OEzaJcOBOJYTZgRYnjkBq2KxT5aFSHye0cW+02ZCxa2l/WpI6SzFv9P1bQfN2Gebkl
z/snOMayu0dRNt/9axAd1HFN2KGDcPRCEg0aSOXD/8XWJDCdiHpchyca8jRXzKntYBYnj3Y3/Tsa
CBMTLdRTf65GrN2wHL/1z1edg452DmExQeYIJZNgjSJw2Rn8zFm4wrWlB7hHWw++UUFKyTIJhKAl
J0lYiWR+Y/dCFngb6HQr1Is/thDoGeUEKXecjBH+M4upiqDoCn0Maq4/N343FmrfArhJ/qWX1YM+
A1SV345nl0BaRz0tkaDlFRBKQLBDvbiqiu8fhUQIsEJhNCqmKIOUfGJXUUiNvOk90rlw8MELXcPX
V8iCIgbijCwfGeggbacdxUD05oIlqaDOVBrHQKhVhesNJdiZtHlrRt8k3uZqQ/r+aEnwhKYNXSgm
XdS3HeyZvZEmEdcz4iMaWSIAPL/Z3ROyjVZzPvy6GX9vAyViM1t7D90Oy0ebnaH6QFB4wD0DKcPN
eXmgPJd2XBDdMpTWGD3lP7MzHI87ZvZBLiyc8732j7dxJgzq2Z03nUeSb6uzrXzW7BwG4S00xALo
sJFprPub2R4aC4K7yPISWP0RaXXMyxKRCwX6J8qXQjJ+wEHIZtSLyv7v2aXmbh3yiSqUIwF1pHRZ
uFOPXn1rtjl9pWulFGiYutoT9256x75ZWQfeU4r/Jp3q/yZhiAvqp0UMCqatMuqalnMJjKIODq0s
Cs4toMWF6yuaDgwFqfm3BoQQLdvV/IN9Xn6hiuxCGYYxpTywGLlU7Aw8UtMReHWEroLd6YsvyMAa
z38cNjluPA3JtSRJ/iGE114hMFld4pDlU4En7MqvMrXNye6vixeQAxad7ZFS5zd/imeJHpKEP2Bf
q+xmAyR38ThhTD+AjJGyDZ0mo+IvNa9r/DGQ2nWgvf1G1ai6qT/Rtxw9+fLe0oTuKIMvGHxCboMN
KOdU98pKRnmCUnDlNY5KH6Kn8II+PmywizOh9xsYowUlhTtKNBERuzgiMEsLQ2waE9QH2jA87ELp
LX/bKPjjlpdg2WYfhniMvC6CB3Ei9uQPj86lXtRmBRWsPk8ZJyZBN9ltlhajnOij02LHhQWELbat
coSD7Hs+iIeNIdpTbBivJuXhl6NyWaSNqe/tmXcM0Czn4/cM/HPaX/H9PlyutcOPAvbu9MBEj4wH
X9sMYo2wmDlKg+1K9qgFP2kIFr4Gy8KTA3rPv0an/wq+doDd6FcYVdtJHEGx9G/fZJem3lKVMAeH
vPpq75rs+0L2RoN9x/pc4jGcWYBv8gYzMJqVc5bJYuDwRFV18iH5iqbfwGPQ07OxR2+lDZi46U2e
tnYWOgK5UgVG1gtIXUdAvNuhfUiRLMPJuVZbm27XQhf54AJUdBvPzM+9ZawT9s0hFuns02gxjlk2
p6VyG1boVpvom/FyOUFI0VUgEaFIv/MK8Elkkla1u6UW7KUSOTsmrjnSyHUDx6mEK9r7gLjhNB7T
5cnM3KoBUg6c7hF+J6beAMqMBb3yISnArYm6rJsF+ke2sHWHZHXTHocPl10URX66ZoyEcN0wbnsL
5d8V80XEQLlmrcBJCYX+/p0Vntlf/uK/bc+aEODysypWPjPqXFe3VgzK9nS1b5cuHS0bBekPHyQg
wfU8yXxrqgI30E3LV57NLswCmeV9oXD/31fRHV3BubT8s8UaauItQFV768Nmt5Gggg1RtJ7fvIPA
1x73M/Fr0ys1X4d4HZ7bX71sQ7bJ/ItCBioHQgROzHd5ayZS9x4ZJgyp9+N6cM1Fa67Z38Hpo8y2
RVh3NbCXVyQoZdO+OL2w1XBgt7XmlT5uxZuhAJQ80hfZAubLu1N4RtTK9ZzhoO/QULeLL/0fW2gP
b6GSChkUAQUuvtrgObbEZAsWBfrmcX2JDI0eNFy+tOZu1QcB78cmn2BC1HALPfuGhqOVmBtLUZ2E
UVhmPartFITwyzgiWUwaR/OBf7TVG4MwQHF0wlCWFLMwv66Ht7meMUU5uZZ0B2W5ngCJy/QxLzKi
nm3p9N4+Nkpb+UuxmN8HSlkBFQJjWHT8LiHeD3ejKCpg84OY6pV8LlVxQCGdKRDkDjDPq1KV0rRo
cPF4R2k1I4P4+ZuHge46j/f/rp0F9JksfsAFtX5CrvDopoPtqi5J+kX4Pdzy77AMkGvpc7dPErmq
4EHzzByhXvUiaZzJPPSU4m6Jc7BdahH0cQ0jVjf335kc18j9K9NzGHGUWfcYrDkQQ8efWlrQyObJ
L+Fqbt3KxOsYyMyiQ40iqolnOXxtFNQPWuQm4LRslvEMVzhGjy761O9TQa5x9AJZF5Nv3Uw/qfjS
gYc4rCzvDQRpWLbNdXFzpK0kIgw0/s85zlHg0T+wOPx3TQOxMeiRjencFv0PhNg4RASR2ootROIP
/fsV/wnx71Owj0kR0typzd6AK88nblFfxQZYeAW8zpHBf0I9mtMXMpjAJ0MnQ9oe3oPofiNmFdz4
L4JaqgPD4b5c42JNOatqpVz/PhLJ7rkqcFHHugD0bw1dAjF+0U+1Lz6aFe8CkypkuiPuGRfZx/UA
GAie0GlUh/IfSGI7/WZcWtMtV7zXn1YcTn7raxi/ip3mAjLYsTTFPfoubSNEXC1MYcjOwtYApnWi
CHefMTWaWAz1C6/MPvO9hifKNzcu80KrgboCi52dseXhKHciczFEVyKvs7rBm+Qej4xNTm3Prw90
rGDgA43DXE/yaQ65ZjnO0+U9WC1hQss+Ws3OGdu9KbhG5mnbCI3JhbiTwPRWlFrBAUoakU/XJnam
pbyqWOsEiYKclTNSwBjSHMjdPHmlzBOXPBmwYu6WG0sEnm829XIgODdMD4q+NwJILs1x8NBdnDty
bM75uHikmTtRHxtwRRD5BT4cDeKo6HeNvzixCx8f7j0W+AuUuFdE987N7RuNzbzpncVl0kHVg6Ba
IPg5GFc1tp+5QDf4WtlxMmtug2t2AyZMX1x5EB80IZuwdCNojB1r9T2j0SRIaVo4TSmL3TKOIn9K
ThHlx27ne8vIIbifmlHgfMe4zsBzr+mR5kMtIoV5cJ80ND4tAGElZckynwKaSYDLAteREOOx0SON
l7GmQJ/mmOprp/q2xaZMkH9QbQmCArTvReP+cSFAr9ofC+d6yeItHo7f/sxXFC7mLIZQ6GlENBOn
aqEfg7bJNeOZzqnQmFMUxc0Lf17ZMBtTrHGe7CyB2pWtpnRs/ckhpdq8gZM/Jtdrk2V+tNZOavWd
afgOHA1Ib+S7zpEzKFSunjE9RHW9DbwNMofLdxwT24rkNUOUie77Bc1vmmF3z+1TBC0CTg7nTdgg
b6n+GeOwHNnNi5TWu+a9Y7JWsBSYRdQaYmsVs5cmkKOQXfXMnHOjEGahqUcsWjxWPv+/n+LGMxA2
X6sF4vofOn/Fxv0d+3/K5klm441Sde6i9XFBwDw1I65FaqDU9SkltT2kX1YjApJ5a5xa3fe5CtHE
sY7bGz5i2NvMzMlL2xTHVr/5LY/KOE+Y3IgZ29loKtol/etEjr579uXr0uUO89FhOq/I7vfflxcq
trNTFselzt0ll8qGINbGyzrJISsIqvbBGyRHoWh8TH3dvaMg5p1Q5kvulwSpD+TacaxRo965bCbG
n+8fi2vkAXupCJ8T2sRN1aoIMBBWdS45swPNKLdMLhnDyQRhvWrQ+XOAshc5DYtu3OmmuzXaumdz
ksnNdw3sTSUwGuYvaBSU/WvfImrdqo7gJ4nik66N6EaWiuhEVcodo4T/m9tBnGNzavhH58OijNl8
3a7ErGO8TFfokS2VvXm+V2I/rUdrozYsxVyU6730cUXJna7SLDf5grTwfyultMHpPuXpiVFuuDfj
90FNF3LveWObnHBGY7U4CNnTM2FBatZL6pPVifg+IpyV1GZDjtv24GOF1SniTLHn1MrSyPY3SaIo
rMJbkp6MXg/ZpYvotEJQ0Zf/v+lHtQSnR4vn/J9ulwM4XedYhOHqkXdTHv8hUX1wMphzE3Xq+ORm
IR79WU9F4Rvi7fqnwRhwIBSduaqHJ617gtvb2EViYNKv6rlcJWwapUeORtPF/OjsDUJur9X6OoHx
VLojNWPwO83MhE58oEOWrTYcISOjobyHkQuisCPZmhHg0ge/g9spkqVFpqsaqno2jL35pc+5CWT2
Oc4bv84R+2c22u828HGH144tspQD1rMhIMJPULJ/6d9AjwvASGqTpMvJXG62uC+6VySd5yKRgDch
Xai/CR9YpgklApCjaFxACjSbfc1pxpCOCBxz8LpKe0EoC9JH4poCN54Xf3kdyL08GwBLvRfB4FeH
rxIIlaUBcuM3byr9dt3gvjv7TneHyXqlOL4aVC2wUt9SaAXHhbiZfbF+O2lZz4k1zGgNsmEguLzR
0rZIspFbkDtgFjLOhsbF052nnxzDxff34zawY/LVHMozFBDNGYJUQUwCg8h0/m534Xk2VqJsMXje
StZjep/Kkd4afDgPJ3B0PRSrZYyuWqwae2u7VjKpiZ8ADbxwJPnBnGCFR/bxk87koEaEDsCratts
gRg44PKg4FNcJeQ2vkmCuFPwB5rIetcJ+BMqtftaDc7T3lPv9Y/9dUUKBsOD4rkaCGZop4+4hg0z
LHBBmqi00vk5yjbNJ9mzJPKqErm8tcFy6PyfBbzPVzrUrSlJ9bchQWubOGv952IosApYlVjlmk67
Dxw98Cba+3tEnVC6v+mu6mZjMm14kUDMuscE1VbdY/wfdw4F2ZV2tRfQ8vGVuQEA3mQJeL2Rjam/
ZOIpQ32tL1ZuRPqNULeMSQJDJcBPiWAIpt7fIUe4g1FuRzOHapGR8yGT6BWmePMEbVUhwXoOhsYa
+PNpO9KtL2QxoWV3HWoAc88SZ/Rijcw6NNnV+93LwKTBhYN0120IglWnlxaXZ/9D83x/La8q7K3F
FYRS5lp8sleZziI2G5iv4pFE31e8QGpToTi5fqdEc13mPWWVITIPbKtz2slKgSHa2Y6pSli2ZfE3
68/c4vMpOj5tGXOCbMmsfSHJrRf94wqhi4kjMqvFCSNtskC8L/e7KUiIS0k0lfJAv5Ap30Hil5UG
FBxwkcNla47RwtRP6vytdkJD+TFQcSCNsBJnbzgkxvYENx5dhG9TEdhPMQWhFtBt5K7Xh/gLJXcc
P2F+ymFpDYuGwha7KHwV5PtQ3GWHQYErNjJD0V+plWAc0B4lx83+3V3I6kkzWSItFOVeQ7h3yGqK
vJ+XCA7WNd9/LpOEvlCDfQgPiyQHj/zIGh1OFYUmf96gqZeeIKH7TMia+RrF6TA0CCk8+OpjkoHL
vJNyhihHZHfsKBv/RxEHY1UoLCvWWErB5U5RPyITlU40V/4j0tTN55oTSSy1w6sT5PI4A9xt/8qe
LhZmy/+6AyO8YrfhfOdBvzNXtFVs8TNvZJtuYgO6AfmhPRmjYaiEGsyWY6sDb9tXPJ47sFck9RWb
ZfuvNBrSuV+U03LNtPHK4bguI5sBWk7E2ksfeCEQNOpDQfdw3q900W5yM94Q4a/X/tLvFii0Uj3D
WWQkBQSIIRGtB6n8VWtuDtBKvynm+OQu1wDNIYmkuv1SayIAJhkg9gEv2rn7dqC9O+k5ENyAhcU6
XImU7VzayFHoQnkfpJ64anC7ZFW+V1UlmvMPLn32k4TdsipvlJ1bqrrBCe/pdBAAAmYzj2ZiWdX/
rr32tUohTMrlfTYLbDU9sOxlbB9la7WYOl+dTNqDPYAG5bxul6EkI1WcTEJnzlsY/qmd9joCUvl5
kY5rJOQBQD3sL0powEH/WduCsMYz+Ci21v3Ox3bkP5ADfsdgh9oGbnv4KGVxiosh/Any5m9gRsAJ
uvdbX4W71lwxXmMyfgbx1gwgwltXQzLsNEESXgLt5hd0oN+BwnYozSkpc6L0LTN//X2WDsrRHiT5
UQ3LDmNsdEJpq37X3P1Hf98WdsjNnO307y+CLbJ48euqq+pqDtz5FF3Kfd/CpUIaDenMQ9723Ce6
uaCSvQfeQ9FfBFqqAHZpLD9QK2QQ7G49PF2uc3zgjEIuVIrZgphjPjpLFNviGADZ9BjsPtawi3Vh
S9eJY1u0seerdLPZXz/ri1K1uhkG9nIdMmSm2V0mamhJiMUG8RJQzlEkQudqLk/BA7Eu7wya2w5s
/Pb/1m7p14aRCOYMD72mHLQn7zZyTaG7nVjlqtmHH4NSkoMBI7Gbky7VEmNLtGls3YT9EFU4xAeT
Zw/FwdY8tRDhYMzoh7HoTn1tutA0alFOSc0dXEcXMlYPBmtcEgWIUEptY+MccqZjjYH0l4emG5gd
PGX7NBawmSA+Re88e6RIajKUrMM6jNMQAeXaV4LMruRfkhgK0onvCZKHFzueCAGrdCJCY9Sx1yny
bA9hFFz7ysuQfKMBHuJxaMT7iHWpRfJwNwA4XWHLiAbgAz78fedtMh1fjrzPrQELyXn1HG5o2jNl
NEB8ud85Ob/PTURk4mdyH+9m83NFFtU8MziaewogLxceg6TVK4C4Fkehfrw+9VK9mEBq/UnBfXdz
SwTahUqbhv/WgQC7H/aePqXom+PY0JgfBFzC3FZ94Axqd44EK0uCzPU9iNS/CokOgu1s+ZGDBAoU
13WVKfqXf/e/Nq9rYMN8EGLdVxug7petCJzej/fM1tDKRuUOLTtBGgzj1rZm1yBvE8d6U/qDPr/A
iwZ3e9RxCvclKwGk6zAzqQ7iXTQibPDl1amTG8RSHuKLTO7eC6q9/56nfNBoQDjPTbA6ZGN6iuPi
HFGORqICPxByyvoWHUBq4albSqCrlKMqUQXizUDEt/75f6VMPu63GQGD//Tj+3LDW8vIJgC6ZzUt
Wqc1V193varCHr7tm1HYIpfyMgKkl89LYgO8qLn3ZKwPn7j/8ZPMNR1HAAwfQiGKjlgZ68zuli5Q
adU5ny+hKBK5EGcj9SxN23M4sHG1i8TQQq1ejEHY/sTtQncltR6pkikRcPzqGPXtPRAY3kFV810J
sXGpo8YSmEfs0HXhasgEr7hwC+sNcSuhxQOPRiAO/LQ0T5PLPkYceoLLYlWPscrrIT+X5lcuZdcT
0MoUJw27d7AwvLrWJOeOZzk34lp2u47MWH3HiZXGs0taMwt4K00eS8W8vyohhZ3oddoimM4ybiU/
Vuq0mEcIvXKrU8Kgh+lCeKGC8K+FraorSklZC1s0vvgdTM3Yn5g3q6cImx+XyRaoxN0y6zZ/oIpr
6tOmhlidQsDM2nQyuG2TvikaBDXE1U+JBC33Wd5qZ2ZwI0motcGbsIE4zxXa+NJ3BDffDmFUyolf
Y3NIlW0z1aWaj9+2UETxNqeFtwRlcBekz4rTg8JcSt0t2l9ChRvUgmzIIQbxjuN4ME6cY0RJqwh7
/V5fb19E1YnvWQBrm74QkmFwO0U5S7x2FsS4s5cfRyk7Jpc6d/+cOJdAE0+vK64LBL6lGwhav01T
2QqBHLiD4vngwkovGIZZjwzzTzwzYzv072UJQ1WPtSkhPXJCbja2ecmBeZvB028Nrg2Tzv/kG8r9
crIjsZS8iVSWvIkNTpH6mC7zUVlbITgDDtdU0vy3klxP8aWPV17oSTR4yrowyUS6UUol4K4R31A1
gS1xlauDZqrPDPaCT/EAJzla8qjqHtAKv/zqQLVQR+J6ch0D38BTy+/4mwBvhxoN42pkaB2DCkV3
BscwNrI13HW3yX87iOwCvTqFddH8zaEiDw8U8lRebYyN5JkeufL1vnkELqMKcZ8Tj1oRhRN3nP8g
9zJkhivllemD/0gJsKZwbToG8lJnuzU07i2jipqNrKAJHlhMPaaot2Ts48NGfHWmBtT/GQ0jVAU/
ucy81n4642BaWTK8+q106wuOJ1sl9gRRs4siKB7X33VD0wtEipmSp3xjecc0U9F+1VF6utBPYIFd
coYurEFarHB+qXAxL0JozMtKQ+3GkcG7Z1CcOcKwjtvg9Q6Jps7ebnZSCMjIj1yAt2eq7wli8vs0
EIjgBNKnpMqcVZyoTt3fwiQvfMjv109r36HRuR3+bN0w4ctUyA7ox+t9XuCdAvQo9D8Bpna90odW
idS78a9yLknyA2a1x5VbDBI+nF8RRlxXLt4CVjLNrAgpJ9INQ8T+XLeu6rmtOFV4i/tekCrt/PXi
E02WGx7kuoolwyY/F/S2nmlL5sFmL0zYYJ9XZHJKynfr35iyJijl2PsvWhrqUsHW8nIBCrjwT5jr
f3IFJid7rNElUjffvw8a8d17q4yx6TOtktutA3MmxbLOJs7RRFLPFHCRDJYpILCnj9K6hvlAeS2p
195XTPBBaZZyD1SHEw85TLQZG3L3A6RQmb/rLKMfXduHp7tunegPgXwJXuePsPMpg44rr37FmSY/
yv3s5Okga1YmSJrp5C6KJXfhq+lyJGgT5kPe25isqfb9fM1IwSC8MC5VBqiLUMWgXHlG1QX4f45R
mBn4zEulqRn2/XXzQ5HrPhMHd8UlgTilHQoYmOAGo0Y4aC8Su1+ufk3KzXid9VC+NYSCicXSp+tU
zrZM6Z52EaeEo+Kka+wk1C1g058j/Se+5p12aJ70mFDCVRKTK3ViL+ag6GeFoFgr1Co5c793VRjC
9JlwWb2WrJO3OCw8Fb1cg/gTUyNLL3QA+/CpCx0PszV+9uBugYWlbk8JhJC8AXa4WyMhl6GBawIu
IX4AKS9E7C0UpR57EXrBzFueVFTAq2oLBi2R+llfBww/zYzEXCH/7/h1oRqgIhPhToMa4kBvdqTU
Rx9Rv3NmsvpJwlFVwVOh1pjTolSzckfsiiaT7s7K0eMTqqQwtV/UC2kbHi7qidv+PkmmNOHmdCdY
SSkgTEEHYdnX1oXzGcFeLgRmMl33NJPzSRKsBEkwPKBQfPyQexEEDwHmqtySSSD8VyopHaQVWyRE
vt33KF1QPEEIP3sTHg/F4XuXDSHE3NbwrInQxi/M7kzmki+tin+EMoEBlMiZxujL3lSsvI4eQym9
Xy0lOhi0lYBU2I5oLBhFZAVX0h9FJl44XvYjLFPDDEn6l5+9raI+GJ0QM7VEKlGNS32Fm7CMhw4s
5NoLT2LMm2YQ7iWfCk2Vd+fvVTeSajO9uDokiD/iMQl4fCV/ds/gaMJtP8pBmZaor9zWfUXddx9q
wHnYsbu/IXUvEZnioan+rsynyhFH02i2GQn2Mi2byKxRkWCJaNsphU908hhjODMtikrqVsTHixKR
fAGDcnGs2O4ORAWuMSZHhJckAVqkQKv7p3hB5714pGvbUELyEq7SBJ7v2E8XN/TQaMLhO0v84GTU
P3gx37CMbNEtJ+MHxjyBewX9n+guGIBzvBe4oOp3vL9ieIROKLjPyHaMldeZzAXdtr6Xk4+zgPSo
1Yr/O7++QcMTpvXxADjbYS5K4qur8cE5CRmjmVlg6FcJe14+BzrpFAhsbsBt5gfyp0TNffEh4bOw
DXF7ye0x8C1O75U9rT3pHIAI5dFRROHMwFo6XCF2CeIb3kgl9ljuSBgCJwNkgEsvq/40bCSACUYJ
r21Ngun/xFVDp2McneIe9umCokfAYle/jWwSVEfgGRhN5jWI43nGUhcCHWLZcq4So+aev18MQCSD
XNkbhYDPjGFt3TgXr5ZfaSZ87IGqfYBP2vtr3Dmc41C1sq62GJ15RAPDnbKjhRP7JmwgRvm2eBQ9
k2bChxFn+mCovLe7wt5DjVAFFuBxbkUnTC41XpcZIl4xE7xnGitzIUJjTxEqpTmO7a2pv2lmlx5A
PDoMUhOpCBMw0xgEf+7teeGLaCLWEz/zuIznZ2mW2vgw9mUd/H8Jwtr7lZnwv1AyEdaAjX7JvxnZ
XslxXWpElWQFLhLiXHq35xeDELvyLRWa+YufEF9wBJbTgVCRXFANjMZeAKLakSbECnK1zgE+wnCr
XwAfbf0IQiU1TlNIhJhm7K6qeWRrZzXAeQenff8Xkct1NwtQavP8fTe++NXIYeRWy96GqH/i5/6z
hlNHJzw1S9lGeaiVvwA6O8YvfZAdXER2qGQfKHBvbko75ZUhWNurY/3Xl1Zok5j2s9AXSEeI2rMI
bNnOEQaNzskQpfmY5XB+fX/ab7Fcky7fjrn6OhIiLgDaPh2K0/nzBxlntP5eTgomY+PlxniY1UpL
zL2ZqafZom7pNXS3cBVg1cHgFZTWtLG2sbWFG/L3rrfmhWwjdhMm53vs2rDjF898/NMw56g0twQ8
qpRS+txag3AlwDMwIQS07kdfJfO/u7liVf2dkuFFYkr6nlpTbUo4T9as/FprZhlLx47n8ACBQRBA
KTQREohe0e/UHmUApqSUpLCiBrO1436XEdEFg4LsXSdVeUE3REDubdbVXgcz4ga148c7MMH6PlZN
pTSd2ucbmEeKlUJeLglIX5PNCJY1r/G+SuA03hPusAV+7gJ8wXoiVkGh7rkctUi/RibRRK4wCefj
JOcfmDc1N+CJiAFAG4p0BN3zUSRWyHd7tOG4hzsA1+34Ijg6S/4Vnh4XiEdc22fcYaF60aHW8HZj
QkYkCoZ+71agVxmwsnzyUre+mHcR9ukzCQrp/kezc08p6FjY93f7dO4jnQ5gUhhdj3jawpC0rXSY
+6ffilQiH/p42f4OmXW72tz4xGhDjSDvB++D4gHBSgpnGwq9txq1/+NfniFE1nYVlT6O6y0sZuSr
RPoo274ayhpahdmJ31FQV21RFzmk0m7TMFQf+1bLKcPK6gxAklP61km0qGXoR32UwPWul3lI7Ycx
0vhMMuiIcdue/tganwmWqrsHS5eicqiKPi5QUnxc0w56vQs0e4+wKFNEyaXrsXxGmx9JVZOSDbSz
jsChKgnvQNKFvuhb0inS62djx+/NbO0/TVLBcnMWyDgOmEFr1KwSLcC0R3gcvaqZ9X9rclGVRzQc
0ELqqrkwZwEAOGyATd29Qpzc/3L/KEOJN+M8IdTjJasovBw+nV7pDzTJtbi1XjQDQkK/8N+GqHsJ
vkEDigNq9iZHqh5dLg+GT8ePWPVQo2qkFV86mfO7MUMDu7ah7zgGKa885xqQfL/ZDeEdCBqVq7Mn
Z6OnE2xbyzcO6WzkaORkvqZz4CJAaQxR3CRKt4MYH7Vup9a0H2BIaPZ1fU+YhoAIHNrRJiNlUkcE
sn/G3vV/d+AyHpoSM4/TEVYM21CPSQPK8tU5443QYnuTBW7zCBJJYHCo1TlpyNKHFNQuVRU3pi/L
HA6lX/MSNUt/FSPNMHutb0qWfRFC25ZGWqL+CwpwqVmHXeGz2htXJa5G03GW+SB16HNVFPM92pnD
lSkdS/Vh4t6lJ7chibNYBfUA5AjGvm0315kgLwaJU/6ULeM/+0gSUlweifZz5n1ijedOyxnsjl9Y
GY6+g5FUSgRc1EGICbeDut8AP3uwoTbzbELyHA+Pn6nlCqz/NQD2eWGJfLuok7sfO2iT/Vh8/qYr
KbuEzMIasKqplakmGLNbIvwm7vfEMhU7NkjFRBBukb6KPAG2JLw5nLNXbVgUALwPQxgnFf3g8O8u
hqW3ske2JE5CTYB+wlvkXJbiDUUcHcnAM38gjcuizSK21zyf8aWz7ULPeA+DoN/8oGavf9X2eDp3
uBmz3VnDZy/wkd296BqlHnl5ugktzfZffxR2QiBw8q16RZr6G/fTwj5m5bfsXKBalHTd1YdH2DrI
+Md4FU6x3FLw6g1NzC7OByTpqaA67OI6LFdwPrFHDYCiCJd0KZN0k43fDHdFv2OMWPGhC8yX42f3
zweVPL4DDomvlKG266iKXbpL5OZwDGYDDD65yA3U7A4I/TYTxm7FVzBu+LsU9JuyAVxjBQhZNQoZ
tdyMhe3vzl+L5L5UvH69OSWZOPXa7sybQpKmcblfO3EltxKRcjREILC6ikMX2iXj+j4+Zmk3ohNn
ugCNndibfl7o4gSt02A6RJpC3Smf0Zt7bBsLQkJOJPda9IZjE6Rm2l02YbHXaa3mh2sgbD4rs5nm
5ej97GNZAs1OXQY+V02fOb5jzBLRBfRm1tnNV+7LF4xQB/hfFGBj+akMMJ1RIlIndwNx+gO3608D
sJt/86rmnFRiR++RacjG0kZos1SWMONmuz/vmZiuOa5/c26vxcAhEat+I2Y4lOeRVQPRJiUtwwa6
ASzWfNtQD+AY+i9uJp2Ybz3ksiv2n3GBnt5OLRE9g4ARobf47KJMroAil3h9CIzyt7gRlQ+4JR+i
Gm7kRkyQeD+KHtncJgYQuG8U5ibM9qllwPiEViZwDKnh/PL/lDlZyimfZFRKXzL7w7g4IYxGY8PB
ai+aH9JYAKys7W4gkU6nKMosn2ABXIQQahh+Z7iNs4aiOfWMpsdTENgLFEFrl8DN95c0itiEpMRK
r0C9s8bxnIn6uKoJoQAzu0bewvkmSf/wGX+KQBBEi6BLY7hKKZkdBw/y7sj6p2banZxkYZzuSuN1
sxyFdTfdCE0CzfAY+4FLX8QP9G2FgKNIVfOVtSMRnn3HTfqzl755mKTsYGyjXpEZZisjBmF5b5iT
J812IUi5nK0CO6beb6yVaw9Ibu9vN7dJonaqXmrAHNEwgeb/MEai+U4xuqx2Oqu8vh+ZzDklQht/
zRQZKLDPZ5EtsooMl78KJfwVmOkmhC4hJjNsVIHdYlxiPs3BZTlsOP9JLdO4aoWf/SrzlSZgkLFj
cg3WU07/eaB5pAuMbDsDYpSyhopamvrT9k8M/XAf15fY6rQk04o/0+RF360O/Lr8vt8jTzaPbYjZ
h0AZcE6YvtlCrd+ymWFWLs7ZaHuB/QsmnUx76CAXN9DUfaP3ntMrkqKi5xwBZRE3LG3PexEUINxe
lei7rQ9jxGLvVTdznXu7u3fr8TyfAvsgqiaSMf2KN0SaLP2lQdf1nNYeDQXdM+9aSKM6IJnCUTLs
VxoVH14oXeZcBdTCkecS/fcWvBzOXXWXMZa92fknptMUJN+aBis5lHD91lbu+VwtPb7vwYmvUywG
//Kok2FQbvX+MaUZfwV31BPBPFWb2ZRLBa4M7Uj8QqRJLQeuZbF3+DDJQs/EbEH7BJsgEqt7LGEH
nEmpdDqFRfr4D+ae/IsfgGUHp+UTFur0gESeNVaT2J3B7aK5Fvd9XVjQjJeLpImA9cUnfC3VGbUh
goHC+F/1E5Nb18Mm1iqZH37iba8E+Ye4JIO0ylWNOKJp2PVuSGnGO6wjutCWAdVAfmr0/avnXb7u
imYMH7atW+HZ1HktuFazvAPVD/caiX09CiaiglMeo12Xby98CISAUwOxfxm0Hkj4d9EhXbPJsyv8
4IJN71myx0GyN39x3tKocU3/m/uucYFeOGQYjm2e3KR0EuDPBBMrObeT+yKK0yEqnEZ5fpm37KYQ
KjxX0DTnVKDF5CZPs/OPzyEBHbrD0drAgm1SB5AIxGMVgT1FA3KgalamsFnSZEPhkZfVlA+MrTFn
8ZdJsmS7ImFND23dGhE0lBANKjptS3zdoLvJIyWz12mZ+DpCAm9jfPBDJbAvaiz+BnibsGyODgOW
vIyqq0L8IWVxxJIhVOKTiVACQUecUO6ZRq+IB16XKoDkomGpLHwPKtfWhH1E0An9sJRlXaz8Wo5x
X4nc00wNOoWv4aJ6sSctn+BQVE6UOl2eBU8iSUOn09n2HaIBTH/8VhaOQ4XTKYSjsgcQt2hHWQK0
fKYbgtq1qCzha6RyOlNfhHFY55fjSbE8RbI1R1wOxHGYJvkRKh5Kvk/QjdnCwb1n1UMjsWxqf8/K
ayVun5iBTRgq4TfAPrrTP27CoV/5OUd+KacaxPTeTwCZGnBJIZ7FyPTufhadTeliwHvNcVRrpmzP
lBA5gxTI9Jb+EkAcbwMw9Tgs1960Djoj/d68NB3shpM3z0Cn0tPkamzAN1uoG0WMNH9aDa7EjFww
MpdikDU4LrqhzYu+xP/zpiKBAEsKoFaLrFebZmFFtEFTmKnFT2Y9WRgKos7W8ZeBqvBru/MA9PFA
/n14GNE39XYCWpyEvbxIsXcmPuGOcR+f0V+/F/l09r73nKGwdKpFE1d7zrY1C2vvXLZox6GVAu0W
RkvphMEH+ZXstdtFJmN91Fu3tajdP/+sF0q9UAoklF3W3Ux3kz/tFC1cko/MhNBXQq/qTeUQr+FZ
qIAjDVxEAZjt01h/5bCionlHoRDAOqOjGoZWpq+4cV251kmk861MsuV4KifaEOivlVJu13OfdJXh
7o8AQJZfQHCji0fgonNxEH3pbnZWS6K7AhGOSw5spKnF15hkMwf/efIdz6uOJ6278wf7QrV0rkPh
5RwO29g8rKGfhbJo4HJ+etk+rLr1VXcMSUordYGgZqRRxoXHolk7BDOnFi2QYzhnRXXBXG4ErdZN
d6Ly3GQF12TU6uaG5Kz+3N4Syl16foTPPgtHlPWUSJxnoy7UoDxndviTycp/vpRMnkAl+NjVLuW6
y8gPcpoFiWt3MaSFa9X1zLGAcaaN6MYNGN8sswbysgJlDtCLAn71acROVvhYj4wSCHlHCzty9d5o
yUpcuxaD42szlSBdAQklAU+jGpfb2cyZnP+OqBdDfjk8rtEH81TGWVvjJBOooFPysX/BhIgY63ev
qt6+PeL5Ku+H0X12R77N2G9Jvvdnfb0Z7T6zM5g0cCqJ4N2qti+XB4xA2IrkkDkUfjfp5POuKziF
NRm8+9wSSq0qXtuuFvzsruT/6qYHcw0xDMXasNRbN6w1joRPk82sNE2W9Hcgny4RYohl1djqcu3+
DwmJaT8EwwMzQE590KXCrpy7eHMItZ29OrA2OW9Rz3cZy/JckCGqcuh0px7raECOR5m29CAzTEhm
/Jgw90fDnfBP029MqBw1LstQnhr9aHNxIrOOY7pEsCnNhASuIaI6brbYSlnrXwEetFahcQPbXYEZ
gKmvfKuEfCE99jAa9E/U6QQk0emaJZ5y0pjXrkmVdZhJvWSV3+Ho5xDOIa8nlfFjpLX98hv16VW+
ILDIl4tYjGMWOfFPHEabzAKkDxOgVWzKpJcNp73x2+HEcvahyP3dmzmk2oa8V10CNvdVRhMV0mQR
4axMrBjqiQpQfWPemuI+6NnCjk0TXWq0VHn128oHIiD7MRurBcZvx5PkMrraT9yJrbnVrHfMnIyx
KdU9S/J4KRxAwzOwUGbB5S0/PvUAQUrq8b2YXwmVcELqAsaDhQaLD4Jx+/rZyPpPbqXboMIOVtEr
rbimbbqszh2vOai8c0CZf3SAGjhvv+mT4LsN9FM5ZjkklUkfW2ySdb/rxTJ2UASNPmbnStvq6Rbw
XwokOXBUYA4GeHJFFk0UTwYPVSmVMkAulCDXkCQyLp4AkwqhamPblpjKHxlFiB2N4t2bN8UDLLkr
UeOtYF8eaKxF0koQ8MCpVMGAEgwSlHfhGVP8HEj20wT/szTjMHJFbdGIAJihKonD50m8usH3idwc
FGYB/gSUf4C9vNBmSHc1Fjt6LRRL6dGHHej3+bjcynZ3EzoNtnk7TuuAUPPofiV3dKFzk6H0JOba
B399n2JPXfaBfnowrqqOvWMi96cSqBwJO+gyOZJkDMRcNkhydVDhCYDfYS+7GLU0MHNbmN5wrTqS
HddrUVFn4LnL78/wIvuzmKIpo8wrF3roF5KW52jynyV+3oDhdpwEaNOaOasJU9g8zSt3WTw6lMCN
lpzZ1kMhOAmaT5UmOUPgxthJj379VrKztkjms57sjcII1dclFWcUc7qM+qwwZEeVx3OszKQvRlVi
ncN/WR9wblK12PJvaltWxY8TWcCkFafphU10d9+W62tqw1YqtWlAAfNCCFq2Q96PfKkOrn2Laa2o
HLKP4j2LmjLFnO8GygD6ujwBimfEL4N+lkIWtU/IaDav6d0Ra9oWR3uJSy3sXkiuIo+DaDe5pAlC
88IvT4iQTFH6/AgBM0HCkVv3lr75GoNjF/80djLppeAOYjou7yDgizOoAvWopX9Ml1UJxSMECHfh
yN8uuBnFwKh14bqP8WftMyqdT3uV/7BWxlUe8TMp8qCP1Urvjvm259tli2GxZUhPlpvPcKmmuwLW
F71HO79goBCMLOXOaTwo9JGiUL6s7Sm37gsKcKo6e1xneeq0CcsRWZ9zmceTGTu9yTCpZyKb6C2I
k7LxthrqLI8q5OH4UAVQ+u2dZ+8GfQV8oR9Maiwdz3D98GwXqLpF2gqM4JlgAFjzk+iYxxfLvilm
twWrSBDYAwDmykpbTGXv+ttGgJi5nYU3L91Hr9477ytyArOPQvNr5oKA7gZPQJzvgt9ruaomsAtX
nTHhq+heqBuo/4kHSVUHqHqD9SZNoFdLKLa8Uo/R+vlga18tV9L7ENwWNsj+tfqEUR6izoA2Va+d
rYghkc4XkNwtKeyfSXt25BiNQtBdYnYSN2qCAi7Cc+9FiwVsrBbvwcLEVE4AIw/CaHNJjlmBQpXG
MJjiUOSj5fYubf34DfbesqKHoeYk4KdPR+eUe6xlxHsJdVaT8r+VEP4jp61zU1Fxhtgfg10/ShKY
hHYN7Zm2xUd0e0b37va42BThk84T1IL/56oA2p189pyzV6qjpARIzBfbpoLrIHAGuEHzkBz13Zjt
oiMcUDLhsay684oCwpiuIr6GZgv1hF6e4mtrua1RttHyO/Ha59C1G0VMwj1ACa4ZbcaOVJDDKRoC
KlCxwQosgz520mT9aJrNT+UPpZa4jMc5It89xzrAuplyFBka3SYJCeW2chBA+JUWyjrLvsRRd9cE
O0JkA1yIQWw01/sYy3LCoH7L27AnY1Svbt995R0NaVg/m4LNyyX/np1WdI2Yjv6/UwCJGUoi2bZl
G8XF7geOiCeJBuJBLKkFmkEOYJGfmWlrhBO67fbgqtTtWHbk9xIkkelhhrJtiysTCrtDKpA5I/lT
QxBvcHQPrlH1t820iNovzTho6rYDNu8Y8mQfM70Bb+lTJAMhFOjScAXsD5KRcDgwsL24/A6OqSae
seZMq+IEgvK5RpBkWyyHEmQ1hD2Ba/0WJDOUgfARm/gHghX5L5K2VKEnQjIrP3oG8pAgluiQDqIT
0GrwEJVj4TYqVs9OnHRqtfbK3WGrqWKIALRWT6eMzDrDcVrWhLcFdtEH49IdihIJi2co3hXC3lm0
b9k1K0BbBBARZOKSiTj1nM32evRVV31QBFi+OzPSWT8NQDitv6w5O/AcVs2rjYpcxN4hnulsvPmo
QebNZ4QrjzGllSpiYhE07Uc+8cOg03MX+6Vg9HDDFCalOaHF9XRSHUDTsHheVj2mUSIfbpZYmzIc
y46mVTdcdugKoY6GcWTNNOHYdHEbvVDEq0IQ8xtdd7Z9fvxP+vh9HXYwKEIh4XOasU1VdYKy5SdF
mxJUQWHqaPndqAzxOvwZBKwpfsyM6TDbhai9fTr8IuwLR7vdQq3vYEI1J+VGGY1aIZX1Im/dPaJ4
D+H8MbFgAIfithlqBVksuBJDG8TGh19klJiomtARF8iV6Azp9gEzXnrzL9yS45EJ4C5lnv+VLh1f
g7xVevT97o8mz4Vdz+DeOfsxV+z5szPaXNr97Po3L8v7q2xfMDYS147Q0Lin1HvK/98hQB5JtVnO
umDNXa5X2Qovre2BTZiSJdvLm7IaIAKTD6Pq92lFnKM4ie9z3FgPv7eWGQ7MgFX9BDcEF88Ns+CR
9r4x957w1kTmjVMC9OFvmeZY3VLhb9Tu8/bP2A3LV8XHxuWoD0+Q1/Pyr/4oZdWSFK5XllOjbVNk
EORpBPd48DI9SiYQmJhp46AK57SJ5xr6R4FqkcLQGqr79BBEp02LImEoLP5d8lh6XvXMMw1HvHsy
P/p86Wcrl9D6h2Ds+LsVGScEgvh+qvgL4DVH0GKX4zAfrWLWlyxMrtA4ffhydTsRqrrAHO/+DyZm
Nhtsvex+eDLyhT4+LE7ayTg9pxzo3nT1u5QyexqO8tHoEF6sB3h2f0ztw1v1k/gFJ2gENW+6qubm
c1v9rpnj3gtpJP6D5QqKEUd24gIgu0J+9SkoRncRIMQTkR4besrZ37KcRo587hQQNLKzy4lZQ6oS
cRtrD0JLpV+BuD2wLQ5hRT5ef4HJ4rvnKfm2dZTcVbSqQ7nUU2rA8n3jFq+bbZyForiiDDYPVEw+
Uc+PljzMd2J9pgxpydpsDqZER7jpkceoTC9ZM+9hOaq0BFFQSYN9SYoMsGTZuvsboU/ymMYj+rqI
PuFBXaukjIsTY+qHHqbymd9MkosoUoA1Uqc7zxoHPbya/IH9TtkrvkMzAmcjegBSxQS39J4L2CnX
0yBiZzcDiQY+bjHc4DUpgdCKTK6iG0KoBajM3YLdGSzUwF6A+5C0H5BrsCsBYm7VZqYs3+F9e/af
30DKZDHSfaC4vZTNf2BRgLVaw9ICau25LjYBD5ddA+uxRm2TcIZZ1SQ/4/q8hX509eq8mUj7ujO8
R4zu5n25nhTabexQltzMwSMTKcAQbOTTfZ1Jp5G9AOafPe+Be77MC6tGMHHP4GFbTT75uk381gLD
ltMikUXQQTziweFUF7kD367ZXFWE6fz8OtRnHH/7x/tQZ1qUG9D7aUBkOalEechq2vZx6p2jkP9T
C67jS6kSmn2WSv+mcZCLOjUdDKvEf114JhTDHXnouA7CGd6cqipY8Zwn0L+bgEwZi2xDRWbETJAY
El61uFTL5vHYTm9yh1v/2OhA8OfiSIXXRxfXNTPeHklo2J4Pr+nwfMj+Mq42/TJAy7sJcduP34W3
HrvTd4L5Prq1XUnYE5T6iKqJGQAtGIMbrZ0TpHK+I+m1JZ0JHfogo7sSK46KTif+OuTX7OyHOipn
k4m2QgbYw3ph/l/6bak0M9tLszF80vTas8UHB42D6rmUzxwXM3Qxh5jooTVfWDS4kmAb49WyI56V
zuZeM4RggGNL7XURV+YDDmnuRw0ZbcOK9w4mVEYgDoRiE3cW6Lvv6UkEvPOK5qsljklvyksp/E9/
ChydmcR1VKQEq19gffRfiTI+buy2PJCFRMf111HhSWHkMTkETahC7RdHC9KOXGI3n6+GOMqKT2ZA
zQKsgZ4wrs7VjbKPaDzq2Ri2vzfar6hCn0YbWUYWttMsbl/bPdlgsVRgFjNdja0rRxl7XCsXT2b8
caWT/LKYRB5ZxwXK6W8mOybXdsNCr3GDJvwALo4LuuPLpOQYLDNJIFZgyKB3vZpvYR+K0ons2wc+
gQvAtWJCm7FvQMVjhhM+Dr/r97z6aFMInrV2MqJYPoGldju6LAwIjj37nrFboBqRZohllzdvfFjH
5Ih5uNuyqUDkuXQHney0/9mQ12W3GZ7pqSrovySpKiM3EWIipaFHkQQM5LgeML8kEZeFzxB64VFq
aGHadSDE8E/9zd8N3ESUknnuUyNniqFZEhNJ9acoFmOvodTu70G+NPti7njQ/6scuvQlJ3JpqO90
4pH423Tv1m2uZZP/EsBtGCvsz4Aho1WNqYF60ruT2hln8cYgBXj1B4pT3BPMe0vzCVw7WuHZ/dSd
UANwi8Bbqt8xJ1b8TXxPEDT9w0Qp/4srFzhG6ITxWKoxR1iwidAd4Q9ewXN2e8K3RM3kYBKZup1X
KSBZDUiZJMgTu430CC8K76Tv7viVCkgkpzbHfWKPva0cCnqrEhqT/aiuMqR6jxmtf01y6FUfkbOA
MVFi0e2lSkrUQlDm7CLfCWzm1PwByMO4A0vGIISTOJINCOTlAGIfMSEZMGBoxD3BVGI+2OxNRaq6
cjLPXm2dp9bF+2SAbmeZ8VGG5H9sW0WrKlCTDkUc1VtbKzB+y89cPsxJ/qXpyTmMDiSKBaECCzv3
DedNun0dQ+xzyeagOe2u2U6BPZxUBo3z+7eHPhJ36WmsuMBWB71SCQpZFSFqd9taKePtKPshs380
T7EUiEg/BuhRWsw6IRO0hrU/S08B3nt1/TsEjmailN4MqNiuvm+gPgdUxLI6+rEnGBotpLht1In6
qovpJylNsznSfCmnLYVChECSR8JK1VGkZ/h9FzAeQlwWOuygCxPqnV5IHSPu9ChlYaX6Nwlkyp62
R+Fnjjx/3KW3pQExf+19vqB6l6nFptepBWc/j8I5wqQDxK20//WxePDBeqyvG1PTtXGS1uo7cf6h
ZaU6sjNbVNR6nVDHrtaNwL/yneW+yZ2EE3RNUYABZaKL3Kq0ismmmhmm4uh0gbQnKT7BmiXucBFq
4aNqNa7QnIVERGNgsydn1ZdXB7XonyXV+lQtY7WmQyv6F13ww0vFJMgo/OzoKScQY+yiQ+gicGbo
rLNRumfBSixyR5ejq6WbF/Oozi/1AXF+B1+WCThFZH7pAFe0eTaf+mxu2h38aIIMVVPB2jTe6c5t
av6/47o1fwIr+CFBCcPVzMGNuP3QlftMWakhiQL+hJsf9xd8JmnMneMhOhutE8fPvHUCIncMkJbK
IgAvipT3gzuFKSFO7MPxgDTvkFmgyhfkw/uctdkY27Q93q61dR4uVn+VCzuQaPsPD2g9kTUIiGRH
l2zXi0WLJ/50Lv4PBZHxVuET4efuTsyAd0JP0hW47VufDZFy95I6FQk5c3MSsf5F6Omh+C9tPEsk
1H688L41FD/sj2l+w3aKJU4RqQ7bCSDCcv1UGcoWAicapr9dAwIASorcRRT+Q2WOhR6JoNmQjmxo
FipKxnPM6D3FFFVOP8A7DL4kZO6jIJokRk+4GtEoPDK/4EwwK8mcJlz8f84isSDoa9jWA8XT4ifV
8Q8PmpMDXUqT//aspfnIbgBebMcOxHG6NHdajq7Fy1VhwZYQ6t1dpxXzcZT8bZsAFd/bm252Uu3W
Fk9siGZqEKZK5AKeSPY9VPyS33SGCHIc5hdDBCALRXyqjHq5GuzabDaSmqNtjL5yWlggMIhzfBbI
HfwtDyaLEkAK3vX3awdNbfjDJQX40S/YgOGuvoWotxL8LfS7e7y48evRARFIw90GTzbyezkywPlz
7dZLCA8Ze1ptsbB0ZNlMH18Q62Jk7vFmzK/QsN7JokOYnTFKlCWIuWpp5/Ck6yWgWmTbIo0XOSRC
1W0TKUKMAjYWtpdQpyt9kTwzdMgAu/lmVP16yeKGybHWSMdDZHfjiUn94xV6AEdSFWt81raAkL8l
SY/z2BOAOb5CWy8TC2ljsFZ3TSxzalZ8MlT4M3GQb0FpVz5DkygVKDhVDifjfxSqSKXNAvC9Yw6k
StDTRC8ODbuOJRbd9KnWRbO/0ELB7D15SFVjzhXLQF3Z4QT2Ml5LUfHvu6ZZ6SVRqqCOE44rdMZ5
flgWafz7eUsSji2ro0DxeqDGxxtcoTL1ytMb3UF7DuPZuNki9sUnnqHRgGFYWoMj35nX4tuyTmWu
S/iQev3U7tKLVh4MNaW212Qiu8+VR2AcyLnnnxJgY+D3L3WarkKhVFg/W2NCkdm9L5Lcmg1pevqE
F9zkJxTle4Eoklrrx2Qk+bRaM+p6SE6MGtATOtnVixdo20kC60a18PDT487KE7jrzRd9jgo0pfRs
X0LQB0PzSpCh/ZSHRl9YiK0kZkFAMFKDLrUYvPzhfu3b+3qdzL8ryRlN7drIdlQeo8GEQW1dU54I
eEPyXGAR3Y+zdN0Hb1WwPSSU1xy5ZSWU3+Zs7kEAq2vusr1QuIjdyql773s7lBXUCrm/Da8huHAG
4B3GovI2TT8K+gdEB4icOK/NlpktxqnDm7QmDIlzD4EmQXg1ICGe86EX5OmQZAj+EWnCjkrxS7HK
8LmwPImz/h+ZoGDRVkz+1nnc6oqwCr+Vbko7vo8CAKC+YB+ytgzgvbuaUdu9JrfOXw00//GI0u0B
2zNFTp1U5jJieBXEe4+3PGnGBW6sSRHN4QgyKLfwuAxvilw1fVf851kPJd9SiDHTrtPilozgwRYM
QrfhijG37K/tcvHXgJgciO4B5IcREHEBYMWwTbPu/HAxSZ2NB61BNzprh3BZDkrG0CesJwFaPj7+
eUb+dXMaduSNu2bg4ECBE42OpqnLkrfAYUPp7+9IniLc3MvU074mzLe6H/CqYgRpSOMRPMGL/w94
Kie6Ady+mdXxwbIKaRePE65sFyxXLr0DRUcYvKcG5rjEgBvV8BXS/Kn8fyhcq/iF3UgnQAnx59ll
TfXxiWgYUFLFISimB88eUasrxUggH/8Xc7vRwA9W88crcMw4+VF3Y387iRkiQOzKfjGci58raNHE
DiIzIp75vsR17EdPNl40mYCKoe/rQteRFhH6lCA59lrpkmvASWce1EZ2zmlGVMaJVpPgMPjjI39q
AZjn4tKsawHTEHuADsXXDiZG0EyUQ7fqadcyGVtgSmA/+y7c5zp4Rbuq+A0jvqxCY72WNDLiOd75
A00vIuJVfLTz58lot3xPNLjKMJGFOvtaPEX1pG7B34OVRB02n5Oqy3Gi/R16h1osfCQ5BmNFsUc5
ghlE69Nhc94pWkfLiQfGMZk1XLboTt4kQY+RlSTmVtwkSUXiKC5lLbnJNtoCMZvjMUjiFN7GZofL
HRLJKh061EqRUd8lhYBxOL39R+ynUhLeafV36ff1aLBFJW9D4IFSkC0+jK6dM13fiLlAtCkEbD4W
kTHMluM/v3rybJqKLSWxzOzXwwxZrSeeWO8vBbhi/J743t8pSH00ClOv11Ur/gCRjCSfou/THW2k
7KniFwqrtQM3XmlL1YSFrWaFR/rT4M8o8yDXw8ywLYKvOrP8KmqfGNCqK2UKPOjZ1DUUqCPhxg3y
2wC49w/3y7f0d9yIkJdkLmXE/x91QkkBEn+MiMfLUPTygo1omuad2wQolDv++gF0m6vDCkxZ6pMi
U5iDeKs/LvdGfgcMMNMHe4gr3v/maJrhcGiCsLTTl01fHGe6c+0brBgU6Aov/mcCYlzAcBUm5OT2
8KUa4miZ1ahsjrdEawqBDNvbTeinibfYvmNqL5FL+Scx8wnVZTKpfn9lCZWIPRGly2KrZViVQAeI
86+/B19cIDMLfXmrkuoNbygFHxLWN2sk3gBkbEOZRQHQohrnSCfevBO0saB+YJExCVBeyG8W8IkK
2NF8iUMqnImOoQq6A3LUu2Q6Se3MeReJ+rfz61KaPz+4clgP3nGXeecKVTR4V8S3VCQvV9u+xGHE
tahAu1OOI/SRawEa2/kAgom2H/LlLq+QEzHx2Mu5+G5fualkB4dSbQcy4a9LOMvMsvbcKcHwBzXN
Gh2SOapkcTubfXVWpOeJjLE6S/HKhlzA8m97jgq9XIynkgSjK9FAgxJckivI7mUBB6xhmJtFqgrO
GqmQS3o2wQ39+sUMFoPXIU/k+22pnionWZdVxWh9L529MtfWPJEGWxx5taCWSMVm0U3SgYbJqzAO
aMGFVBKK4uw/fHa9sitKjhyZf6eqoa9W5UqMOWaDlLCW8yMQzeMqbNLgDo3cW5VlmxnbnsKZHbbZ
Hyy9vfHXY7Ve+CTb3RfsimVD6wsm/bkyI889+LAyIwB14E1t05f/llolBlQ9kR6aOurwHNEFQy8k
BkEnVzM59LU46FrZjmyXK0YizUkc4/RO4o0xYw3lpvd68+l1Vc1wISE2pDk3ilPPjZQs5y6jrWyp
jHK3m9RqwFwuXbTS+uf0IMuDVzwzDG+CgXr+CbB1nhGjUSmxL0NbAqvMrnZ68mMx26a0RO21FBUW
S8IjR8blORp3inzX9R3mydiaGFo3pVzgOQRMobFxBHilGUHdt9/3mhnC8ekAqcDU6tIz5f4m/dDw
rKJTyuuehXZ0YQQvJd4AFvjKr9cGogn2910+pmS1udD0whQKZLRyIBMAwhLaGMzzaG2M6ESNGuB3
use/iDiuy1AJh5c1NIj2T6xExlVZmYUj7/VFOoficIX5PJ6nX9AWbKNW/6SoPx16X4+9jdRPNTVZ
oJ3rWoed5cXxHh9JKM2vySU4DVjczXP8xsgaqfmzQESgHmB0Pod1Ufqunq6kRqJG4W58xOf2dA+v
41fgfGTdQeXGeNYGFjGSw1is3KPVma7MdUtZ2l9H+2B+jFitVKj2VTyMwZRTB39gm9Xm3IPG8rkc
n/YXwm5nDopAaaO3IECTNIlH+4sR9RbeIA6zxQUJrScDYCie+Pdhd0pUGTi/NV5+7IOPL+vziiaH
Zgc9b/NAsgGWtPuBwvRQ+uTLqacUJY631Uo5kRNS018TsDZy4sx9C0vWoX7YT7z1210DmnygtePV
/Hi2aSdwr52+9ZwfCrzBvvzuNk6CdnIItsSLIU3cBl693clCsUtKR/r7ijCLQQglc2lz3Wb0BLwG
O7ldBxUJTmZSsRl+hjTRK6fdL+zA4Y5MfzO8Tomix6Nisz3snbsBZHxg4yCFInTay9uWs5wUKjKt
9YROdUoaVFx5HxkaFTHfWwloiF3tDhCNJ2ONIga/DIAEhwrnX7h222NXj17/vCzxYNS8dFbGyxrZ
bWeyjEWf0KJxVIWTprzCudItRMO4pQ/9BI8YN4316nAI9C0J8LsQpXQUNm+qxsUCUnmfOITLGCf/
HUuELkAxW7OUiE6z9z/Ejr+xHBPk2VC0E9XliPjvIBEIJMAX769mBNFZU1dgcMUeQBkxxbyxr1Y6
/cS3qG7oh8eQJ5sl78OKf/vsY9vVmIuVaHyde6CRHCObP0EJqz5cTBpfZR1cUe7lS67mPqyeZ/SE
h+o8GigXItzj5rqJTuC1RWXDnbfyHW2B/TBwC3pEMRKK2LuJCJrsHdzW/jCst05jQqr6znrF9Vn7
03smExL5NemDgawfQmttORhdIVr9duL04iQCnKtbG1Yx7MeLnIymKol3wie64mjqmfDC87p+ygTX
QIOQai1zbPkjlDUVkuZNwtlQR6viy4Qs89p/UyVDLUYn/I1J975v1CioFRXS7CG2W5iZHWr4ex0O
VXsIlTfYFP0x5ZGv2LNr2ywQWrrBAOtZY9x2PREQ18NPamuGOjD5sARK/dWnS9LkdIbtS+H/EZmQ
PRORFgD0YbTqqrJJ76Jgglv8LM5INW3a28veAP4AJuIDhto0Dr1PFwlvOyMa/RiXj34yS8Urw1Zi
c/bUJ1/xHQK21euxfYJbSy1J2mAx9DkXYzqFB6i8q5eyAVl6xX9G6iqJfnQ2yVhZu3g84HWjjYnD
I1d5jdmpbX7c6TfLiK8grtKCPChuk5hYCEjPhmOrR0ZIXDhoNHCz3u1vGLZLw933ez5BE2AUuRBN
GTQy9PWqasnGvcha1G3Po1Y4hSbW6SCamhQTyFhFLmRZsg2YOADvxEfgc1IurgBB65JOHJdEiiZB
+dKB7fb9eZJ9e34PNjt10XaRKo2VXFHZ6iXhoWjAtQJFdAg9ZURv+0VTak+755izOjcHiNzAiojA
u5w9nttq+5Dmso07XYVfeAeXA2cYDB9MG4Dl0VpCk5Gzkun5VM2jZY1CQYZMOKM0OuAoRCRbD8eP
kY2U8uqQW2w1jK9EC+eJ7wqUIS1cm0vte4WrHWUqMmBbCdJ9ubxUHlD35qthcRNfKyRToVotFqO6
5OEvKx3AhHCfMAs5+gYLFzF7GrIAwYxWd2on7zohq4lDBy7jyBpeU0HAJk1ttFTQRTC5nyk33eMG
/DjHVueLMRYC7aedsLUbuIAHq0ZCOiA5bzfbyx7/TuKdRGUmk2KzQwY29puWFUuRiYRrihK40bEK
xXXer7jQWBDj8GTLxioxRZWlI830gPwRANsKRMTYCWk7TUGhXjHuLGmw9wB5W9UQ6nl6OntbG2+K
jHeaRiUGkLrwjPc0oM0Osi9S2y5tjpQcSbyAXukndnmJRXCcW7fErRC/+TRyu6zHWCB8xzI82D2a
voinPXvsfEQn+iI9ow6L/19imBgVpPQ8yOv1F5EEAh6AZDno/CzD/Jxhv3YxTNERoFadJJcUcsJz
wXMrmlBL9Khmq2ToYTiA7wjzKOIWN8iCCKowaJ9b+6kPAhk7aexYHFLbp2FofSXfVi8S3bkbgytS
5yXW44c0HdwuPyFwJ9MWr2vsbo0H81yRyjhtP1QPXv0xSBA8G1J/62HQSyZb1WuiEZW8ytpZdRhn
tfaqK00ZZgzPdrIBABQAHtM8WpaCPJJbqBTwBQaPCjnpk2Hq+R6GL+2gaZvm4tg5GSzow9KohnxA
f2BUVu2Y3XDuC9n7XRvBtPZ2UXQN39+gFtipjm48k4swBbilF5mMqnqlWkW+XJyx6zg2UuVmHcpn
U48ZUtnGOfL5QwmlzQojAY5Ct5rFVwVqOsqwT9IJzTJJKx0lpF02DImQ57nd/R7CWxzDpSuUkmLr
pmv2fIv3WIxy2K0ospsAxB+1QorpVqj+YTt9HIAMHDHoe34PEKMQ3gnPhLrvuBRjcKW7uVKtRcIx
RqYkeAT0Xp6DW+7tqFSjkPK/eqM5GhTXnPUiB+V9D2pwN0fSLLfKbnTekha0YgdjPht3bIqu51YA
Pehft5igPp8FYj30A4O+JDl49gEgHkoXzXhcciLOfZM2+YAymHmFiXBYLMacZc3S6xRhjzRxpmE1
nBgxOYUC7/H/dlEnhWAthA1KLUZh+Od5Z5UyRjZ3SiHk+GSI0ubfbeBOqLNXYz/xsZeY6ZZFpO8H
U4zM174lIzj6isuWKW8HZJ19bJQVk9RbNSXtOtSKLgdK+ocN5rSoWprhb5bYg6xAfLttxrAiYenA
aUzBURzUaMo7O2jyLwEZlU/sdGv698f6oh4kVHY7okolmcI0dUcK7weAWWak6D4eRueHRBCsNQzU
um1dkrzdT8tMEEQxAhfwx8NbZowfyGaaV4vSlS/W3uIAGCjUqLupSDBd0mLtexcICO7o+u1RZf/z
LZPbINi/QJWui7cYsJPkcl4otE6iHLruDA2a5lR0B/8TUg17k6/exuwWpSrUEh2RBn1ANZZF6VPk
GcrfMCwAeq4FsamIOWVG81/RnqQGQqskaZx1nooaZO+jcZXpu3eayQnsMlY43LpagUvaOjW1GozJ
OFzGLkrP+f55XgSaKWLNET4xmsVhL7q4WIc2N6BdsWeSFe2+1g5iE+rftiW1/grNABLvkiIGZaSp
uBA/3YJ/pzQyZElnnUgcMA9uK0Dzc8SeHxa6GxzqxBQfgR4i14IUU5TGTwndNzOL3HgGhOCmH7oJ
MUKeQBHkBnZtt5Uo6IRawXyrqgaaZ9wcFbr+S5aAXsHrAam7kx2sMRAhguEdMCHmpbzZvwY+QIke
OJfDKlwerJH47eIyMsqrzpYUKzzwCx0cTKyTL25kPdOwrahTCCWELBN7jWl1LzP2L17FztbS7p56
9sFehs3kwVZISqIKexAbkzyhGvepPPIM7yQFCGErJXhtyiAuZC4bIF1gwbPnCR2w55h6XWlo4Iu6
ptwo5x5y7CPTmanCf5a5ure+0/dhzbEzbBs4Ya/FZ9xGH1LvR0OY93c1LrrZGxVvF9581/Mnu+UG
EYTqOrFGfXiLYcZC6KtXMs1lpQbNH4gs4mj6kpWxC6tQ2+RnA4o28v6j5q4HfmlMe1r3bA2kYQle
3BgoSmGNIs3ldSCglTAOEIWCukALSEYMtdzkHHhmffaQlpDdDpmOhdKc2KjgKMAiOCihIfDupGE9
1X/sRQ4xWE/W26br6RRmrDwqQRxVSIL07imwNseElp0pxP6lETORrYGUScn7EfMSiag1LR+Act7z
N3yYeaL/9qudSAthfoOo16hpzHMi3g0m1CuywruenfkxVygK0XwwriYbRUPd1Cahof6MpS6G8bKP
1qox0AOpJbYOCc7VRWfjHV5ucHfGU86Qm9eXBMbC1errhnMfa6q9mSECCsuK2BzMlrfdNWGesLqX
6zwDWtiYRJ1avDyd3pB5SvPupvLCM5jUrEn7LWDNAVs/ATFjs++AlaOHrp5etHwbDHdKL0NQVz1d
BqqgYadhlPPZ3n48zLqc3ik5hNUb33cUOHH3LpMMTGIi6QuXK/ijXlat2UisMAwg6jtavR8M/bzi
/xs52XK1I/FF7rwl2v0Hwvl1+jpYEUpi6K7i/G7KSrToB/EY/dxqmYlWRJjNzyON5OYyec6A1vfG
4lUDZywK/CJWpXn+Locp0FDXJN2rBPHNXS/gckiYbdCBgHh2O2uN4mLZQzEiLJSIeuNT89E9r9u0
inLrmVGNFk6T1eUUDCam3JLQba9+C4Ao4fGjd3nWPmVVO01G4PChW0yYGL3FQIL5hOBxBLzc4r7G
DVEKsmQOEq2JywXnBPOVr9nNyKtAO4EwKdi7BUI2Z/hqH8hUqxBh6suB91m3NzdyB83Hr9xyaXRh
3W/BLeP9JjIakkMmATIh5gFW1ycrMQcFFAw9eTg45/oqtTjLZZjbo3g/hXObqnakcN74UfHcixFu
n64WGehzfmf3bKbtwQCfLT3xjha7Z6/0hHFF/Cs5dA7Xahp19Q6hrmy1lJxkEU4JZyn7pQEHUFrn
7132x7Cjq4Jfa3S0nJwbFR1I74kxkiBg/qozv2Lo75ta9gv5FTa87uCjQ9Ef4uscOZVZFJ6/YUdv
kGxBEYCvCtCaAufxB1uOpjkBkR8Tn0v+MbWnd16pKLg+Qt8OnENSGg5NHYCGipW+VW+Q0KJiBL3H
NZ2jTcyXA4mE7KCZmXpqfbG+by75S5sLeZjsWDBgieQOvtgjlGyZwOzxvvVtXLrpH2Vvy5azt9rf
0d/RSdo5X0R2SNDdnLRvtAwXox/DG5LKw48CJmgJxR+Spl+6MxoZ1sJI+HPGia9v1mt+xXtoXV7Q
+XpM408CgxWT/afWczUfnMVetqjZQov7dq4aA5V20M1CMn9GiP+V9thQInoi8B4PyJgkCxbtR1zh
5YMkZBKcARrHBHKAkav9TSU9CTW9c8RmUBh9cbqO40fp0nKMXMBoiwC0IJn+fnHmr+o2BgV7TDCN
3y+/tPuehOAXZmmhhOWNJphCl/2IrEfbpj8bWNcbsV5JWRSMh3YOr800qBiy6eTKq4LM/gadE3HU
UlXYO2dxGmbkkdnYBIKv1aY5RPHSAb3Co0yuBZFbg2G9asF1kjpueQ66dvGrfHLZGcnppc4JcKMX
a2rXdV3srrgzn1+ijJNodmXjmZ8FpUzNgCO+LrYQb1sEpOZ81zGMNNh2XRGohfHi1keb0sHItCw+
MuzgtiJ6B8YQrXSCIL3eXh8dccqgcoXTJZwcj/nl0SJxkNCiCUKMRMBcGLCwS43gQpT5LhOf5L8J
U8LDkTHuAZs9NgRH1ASgdCAECF3cCB4mAyDM8QegtWuAOCQDKUjyeNu9Wia13Aor1e87zDblHsgI
Q/uRx+yfwi1HPycwdMDVpjj7N8NpoN3uKZ8Z7vO5DR3Fbmy7un4xc9F2+n7kSLj7/RQViYbFIHxi
zt9Lq5ezRoIqYEyugf/SQUZUC+zNOPpgy5unQYTJ2W5NzZ/m9DcxywvF6NWdgfrc3ffA2/pL2Hp0
FXcI/nvfHuM23eXrANhEJfXBVHe7nZ+KvIM8lnsmtwpDgXTsvWv4COkwLPwjiM+ROBpbqNl4W9t3
hlaXGK2T4DrMb0scjjXwm0gm1AkuWgQf1iY0mjVIKpCZaVN090oZL3D2JtwinLQRTIOn0ARwWJiH
u8jcSDM70V9K4x8NDupnQA9E5srJn6xTI09tsTOyBsy6hnV4H1lFCjttRdhIj5ptopLKG21Tfx0I
1LKtmpcbL0mf8KreduenJhOWV7vyUKsRNvNkV94+J1Rc0ZjeJ0uVBCpgyjkQ88tQqQNkzzcetjI4
75Z9XKayypVtak5ICXmTIYWk+0OPBugAwI42wq2FECNPG2rcW5QhnUdozXN7HP7HfzbvfV0l9/Xr
aOjchEUH7Ovf7l30ZL3gVC3myVYqsANGafBRJ35yLx7IA4RDPViNi94YTyAPvF0i2kk+2bJoG8t/
6MEPN/sJk4yyn6jJiVlZDBRZntli3tRddKwQ48OplQ+GzkbdKCeVVEdz5WZvaIZ3bFgVmhvGF9kI
vxNSD6ot2qpL5Tpylc+HVjaWiMY3KAwhJ9ZPL/BZTyX9v+er046/snLXkFK1v67RU+CPL7aoT9xA
T4JfmGHyfR9/BMFXef7EZMwDcRqSB2DdrsqaIapaH7kkMOQv5KmfDwofjHAkg6q9X6YIHAvarvRA
sGDa9tD3oMjaGAWa2ouXdmBG9bW2r0uyIsf9OTVChJsQdkQ60XWROkihPQnf319gvoxBnRwnyIHg
CrQ4p8sBpsLTDB75sVCrQ6tnwN/R7kBLhGLfEEBzTji7o8ysyxHNA/ozPROmddkosdt1zSnKf+4F
xGMvfirGuL3honOlYsByRPXMcfdOOnOzmQhRvTsMiON7uzjlZcDpT6XvJpTGLNbWrTlFTSV9Sw5b
fK6bp0Qaj5TX+2aFAITM0KynTTZy4MQjfyZlVCMyd/swLcQSLggByPXgvBLCwn1TqWWY+5JTw7vf
OiYbjrIfQXFioay3sUdbZYdyqYDktOGHihiOB1rUyGBuGrKPs7hJNZqczgTuObazCfzKtIH41Lj/
UKXTXPfyscvFEWAgok7wS5HP5Y+t88Cw9i+Sdl3uRkhWsCyxCsgBAbTXlOLqMGUYV3WZ1f2j0K2v
GT1wn19i7gwJwp+c7IVe62cJya2gD8LnXDyhKgF28d/MjvxqQKBDxVN5qFKODNI9WQujpkNLjdb7
P99Kel4S9Z6wBtsWheB/Sdgu7/UGYgkr/1xy132tby1u/StruLWrD6P4vkTaAJ75FYlvmbN9GMdI
hXfuMNvQzGwevSHQB2X69q6EpsM53Tbf3qD+FcWA2n4Z9qI6e07ErqCrdeXKaCDMHHIHIVh+7WYs
Q4o8JAYZ3LNv3bmQ4jwr/UBTgG6fScoDfzDyHJtDgNEIXNG1Sr5k7aiTKTivWRGzDi5cZf2Ap4gF
QN+pOk/ERYxSyFDjYb7gSvfLyG5oKgHo6qCM2U+F8dxvfQXqALJ98Z5m0xj+KDraXnl/lUAv5gqS
WWfrSbCkLnmZn6/paQZtMVxSp2e+YW3uL4Q0c7FjojRNANq4i5pDijvqqY2bcOwFBzcvBHhmir82
fXJOaNC2vd1PVhpPNoj7eCoc136LrBox2JRmlXJ6JaGiaoWQdHXyr/3JSWqhassLAv0WuzQPtXHy
sK1sU8XB38L9jaMNoLWq+772X2NoJDayQoq+y8nvrtjnxuQbC7Xs1wFBiXZhaMj6KTxfwyN73OMS
K4MvyVoGSgyxSv4Oe+4HJxxH+LboW0i3ukJLs/WZIW6LwMhHfAsHIQ+LqgvSrCvQiDL67HLq6YoL
D5zCTuvDJdRNJ0gd8fR6J92t0HPaKFryer2L3NUx+iwosQDy7EfbBin1Ul71yJuAphud8YXk0ozb
Lxahk5Uq2wlaeF/3oLaiTRJCrrVJos9pKvQA+kAl8Lslm5qawJv7Lnsj06Pc0zUQULgywKHjEsp/
jWITZa6ew4KNJF7c3dEOmlC3QHEG+UsNL3wxgwr2fu/u3sFhgxlWsxpVAbtV2eEA1dKA4pAyI1UK
v5c3ijYxS4ixyCgtJmIXv960VHVxkSrNIROmLF7MCo7NK0dtVn45PiRtvs9Ql6GwW3ttDNCeGFd7
IJ46u7T2agqYDH73aQbyAw3EzHiWKTBCXpcnLoHKwoHd440m2inWLEkm2SFhuvNTZBT5I3v71ZSZ
V47WJmT2Wm6Jc1ATn5ebulgcoyt4N/1zsPxeqN18McMjzp2mEoa81Mp6Fb5U96Kwy5M4XWgJz6lj
FEYzBXMOknDrUx4mgNboxiZ92wNmxsvbwbG5mp9cU6puGz9DYJmREaUgp09FX+aZlO9x61UPpM7T
kOSnMyMA9Bu6RjgarSU0rO9gX3Fe2Ifqgr45bdVEDY9xUJ1IzmT8hSmVFN5wqKpYPbmwynzgH67a
eEKMSHJ4KLpOOrbAsvSVttraeKkwaklBcdWiE5xpRqF2gLNrAEbuEfXcNu0VB8ueasyTMSiFzDrp
emSWzzpIDVmT/0/g1QRgJiLMMdnjYs5jLQ8KG7DIbcIWsLd4EAq5g2fD01cXQw/00pYKSSaDX11t
ifFtiiw3G+iHa7pMQM+Hgtqw1W2/63IfDEMHgPcU75SpjYUWyHbPb47kcx103E2unEKaQXEvLSsl
FsDJ3MCDjUQsCLNi/zXd+/NsokB4NdnnpGpLf+Ulgk+W/wEeCFpD8tTx4pr+wbH5/Kc8OwO4qUl7
dbCfi9V43HvcTlk3kX5kHcnWz/+0OHcYlUX62HGhAx4BXDKl3bo5QwNwETIDWLvUZ2gd3vJgEmN2
1mZxnG6/oM4OmNjfmXoayVhXiWJZcgT31fFG3HKtqnmoARZTk5/ukcJkKQjmMpntLz2kYz1aHXXM
Hbc5Tu0sj010gg5haQes/y3eh8dv38O816TvMlqTZ35uu0C9OmZv5DtdbTO1V9wrnWU66/t8QO9l
KcKzaIKf0iDt32E7Gohz3jkOAVxE0kDCTeXsueSxG5Jr5mTCswLLlvOjOV+iCogVwhfyc4celPx6
ohPCkTV8D1C8nWGMIs3n8TIcpL2RLtkR7lFOQdUrwCQDql6Ay9BUZz4HmX20Lgtcj2WJfsch3f6+
x5GTGVNHfRNXImK9velqZPhF/7t9fom0QVoVxTTJ/7Ye5cpw6gp3A/UFlUN/IjiuUavol4+eRvtb
gSrjkMhOJdeY5SCsD9rftrDloZ3lSsivVU8OKbmfVcFSBjQ/21XXVqgM+8Xym3nD96zpq5yelm/S
LDhju+YO1aQTzPbxXLwkAwqg9YR1N8pRd4K1WtwiZD/hRBqb1RlhB6+23Sp5RurGKagEffNlOkqw
oNQpJd0ClP4sJRjpbssPEWPnXO+VK7A7phi4SkLrOHjVp6A6/ibqpknzCEsKa2KlZb331lyxjkb0
9w14tCQmvuCs9Z15keHv8xnBazCEgG/qWWRuAATz9XQe+2Lkjuw8P1/ZzIcI60shvWnbivraLH9J
n3Fk3y4ai5QkHji5meVKg5R+jFbC5yKeOQS1oRolga1B7YGhDtF+yyVw3joi46D8SmX9kyKw9RPQ
pvN/m8Kfs9x1WExZyD4w458Bc9wfD/8//SALIc1mgG1qPznfNh4iQpBqrvSu1s8bCeFjxy9XQovU
ncz4NE2l1tVDSgCCKVWftrQUxlqJz4jxCMG3gagZbJgKeNtxktGLiTfGnnWDI9PSKWLji4KDP/Vk
22i/il443wrUh8dWkCbfsHZrvRsISlk3HqfuDlMI2gEzhJb8JURNv+OJLo+wiJfnKKSo5MhqZP+/
p/AK+hhGqwesWQsfnmLpv02jycdEgf1BXA3D6m/w5GCcEo5NvjFBAZtShNnWNFRURORoxXU/IZqw
aWV8S/55X1xCm+7kYPwNU/YeoXHve2duqTj9spCtZLbBMwlZ+jJJmdkUOyrOay61aV3uWB75cRcD
ejmSKl12CuTd7PbnjoQ+5IPG/HctHq9A2ln73KdmArqUpdoPSq722Ih54M8PbyxQ4+YSWS5Ystjd
9gsn0F99M2MVykSasqqPWrRuQblfzpj7H2F5U1fEM4Mc9uA80JxmdfIrleXS0BNEoQmkDfc8qR/X
VxluGw8SgP72+ogHIqPk9ABQeRL7xjkNb+5j7kQOWMOkxYMq2Thh6dKvaCkr+fqB9SzsZz+nkd28
FEvh9PWR80rCxrQrGRQx48LfrE9nq+A4N80UJ2dUYuMAMT/aWpnbvEMJeNLA+QwpNoA5imJwH2Gh
xhN6G4Q/N7VrNeTUhKPne22+lY+IfdHOiiOb6LxS1a8/K/wKTAKojAU6MunwEL+hzUaIYmAeRNxE
nrMJgPyw6H65SqWgTM4vGFGAvJUpskDL+7DL3QYmGIbWSxQPfN9ttsAMfNO0fAkXQ/QZUpH/6r6W
wYr5IBraPDnHwlH8hg1RNej1RKxAK5Ssp4T0SyAcCD52O8j4jtzOK0BfBgMQNw/pfV0Q/we30u5O
tpvOrBpN+O178+H48K4YYfcUQGLVZiKaK7q7qhnL4R1EIPRfR6CSpdywGSgLDZviqwK/N9TwVNBQ
OWFwJtxrUqazzofKxCZ0acahwXissdGZJpIU8PAADQ9oDUsCO1uGVhwj3EQZ6NqKO+1HqDVTUYn3
SEZJrPFvsyq0OoRslHZgtobKS0Jqn4sT1gtTtk33x6oTfS+/1O+8wgSAmFucTW5NHNkB6RWVc8gJ
p58R1/9nqJNsh10A/I9b6aGbMpI0CkpbAuExr5E2JWzIfPMUHQ4lFGG91HY6mcOgMrM6GNB/Ecz0
0nAu1t/6AbmXfr9VT9GFpdA/S/Dq1klaRicQBINj8yAi+zBDWsFKednYXhNFgM/upcCNUWVAsjpg
m48IyZ5cN2g6tMYZO3b/djQBw3lvzzvfAi9LtIdhYO6dW2dmRUosCssL8Gd+y6yBChzVW14ueMNm
SaXZbgqZV27iMMLjFc9ugk/UULM7S1a5Ck8CzwOnvSUTtTIy/kw2UyEcYpf5QVxT1kgwkTNHXwW+
uo3vCzBgYWHAdCKpbfSvbeBNjRlXVe7+oGtbajfOdh5Gh7HMJEdgFDhFOIu65ccXTIfK19bWYm87
FeN4wSh7kZS+NQ2odPZ+D4VJDFvKZ1uUnA+BctOl+2gEYfzaPZMlLq80OLNPHB1KaGI7SsabhWIA
TV7kZ/TtJx0QdoVglVsJp4ThoaeJWeV5H/pbv+ULbmfhDH3Fe6uYAaLFmQnpu0DOO/A3MDZNvVKS
FgD+/HgqnzqqPumEH5EikWqiLw4sB5SdO02SmokmWmwJxjNjD4Qi1gzukYMfooR250vbRuGk3va/
DLzl/9tZMh3cqOHR10MH/ejSTXg9vgddDT0/A1xqPDnLr5hp5ypfYvaHWoGCB236NBK0sT4OGvXg
ogy/+uJpHuKjo8K3+oKhcoMntlAyB9soj9S7GrZ8ypDXk4RbliIHpBaILmbP7yTK3JCLBIzw8a8I
S5zLkgvr0u31jFncNfgTXyaHwRGu/iT4r94Va/ZSuPD+m4VPvRYtxWz/K/v91m2nfDvedn75DcQR
hYI7XdfuepNCQjlS5Mdl1/swFLZHN7RMfSSeIVHwthfsQBR5Y0JQ4oVLrNk+9omQi3KLu5BO/DBi
Eac+oQXgir5k5ixx+tmAtku2lizULKyvVrnkHocsQ3WGlDgncs7hsqFnf/nDphLhC13lW6DMf8c/
T2q1VcFDf/YhXWXWbSwXfP32GKqaX1W0YbglqNxH8B5Y3LwiNq37lLYTzAJdKMp8M5KlN8C5M7rJ
ixAGVE336qdQNz245HKmdqtHpojoxl2y66QgkaJ2XeTbaNGHfnVTHgpTunaJ4jVWXO6sA9yZU5yE
VHGPJanJtNS8YDyzS7gXIrXswtk7rLcJff4eKA7kcde6hnh96/nmGGdl4ncpSfGN6airbPxzxIeU
ifeW0JzlEOLPxGQQdfeUl+sNqSNDOyv3g0pATtH5ukwf1N2VLLkJHgcURVHpquu+NIKxdOwdcf9D
Boadobr3XldtznQCjgjJiWPwnc177jPYy6EoTlZ3NSSItvXunqMm6hNuoFOqY3+EetKXPTPArIzW
RpfPOw2T4325NW4VK5xovtg4ueryK7mGHlEpvkTTf68dyDzJCtfiCED09cxxrCIDECnzSUdu8CLF
AnoeD8sCsG1ADzx9BIjHdqQevoLmIHxF9pwB8pnC9zYhVEj47h9T92jw/9r5gJc5jZ03Zqhxqwed
72W6hWBmaaHhAkltUixX5NQbqgopZjwPjttGlwpq8XmLxCesQkzoIUcIFHl6pZCQjR0bomfGDpkU
feDncEd4nQNYU1sJ9/4n4HwqTZnQpS6VPc79labgRzHnGNQPeF/O/7bf0ri2mDEuSsKvVsswk6Qu
33i8kCKIf87kEiAmTo2VOgkYjjYDqLTiMu/29KdJtNHs5o3JG2/a6+RSvk+bsZFcgvio3zB1WIqD
u2CdRE0gaGqsv+rlZTg7bhVlWLeio9rxIrflFDZcMmxxLvRMB0U9vGFSpVcE1g2ZzMhiqP6a55tH
9YD1g2kw5iyW+jJ20yvzvePPseB6IPS3CLaSZEtfFxNeW/ZCGXnqozoqAPmmvsiZwFtQa+Wb91ca
YsdXxKx72l2AGhCfTR8O4OgFslsAMTn2qmwj9tetJ3eaeCIY8cC66t7Ql6LLEx9wSomfoVichIHW
OJWMWZaNDPygBlr8FrcL46wDEvIbTjrr4ESdttJY748Rprax0cNs+z9T58oqlz4C45+kaUN3tb4x
ETP2E+lzebSD/Gr7/1imT0eUfDhfvZFJwVkbzH2mhX9zqwQhZF9p3KoP0XT9YWcZP26WWql4k5ue
cTllsY2lJjYkojMLWhPn9Vaw6+ITPm8SlB0jv+WOweL7BMCsuZcOuh8mtFAyebwM+rR1ju4YZyBL
M3s2FgVR40hj8aIe8Rgggp8mZSzAOlPSZV2H4OwsyXKjfhrtmOUIKvjRhqqn0YIGzXBuqyiKtTIq
GsZP9/G5cl9b0fzI7+haeXipec9150LciOMkHeWjUR05NIMkh7vRVWSiLoOrp6TTZqPG/CnhySoA
t9anv/nObwUkq1zOp9ie2+WJGIq9352t6ShklXK3/1s28ZJxsxMrACXJYGV30vMLzMb3PFDu2XHq
AYmjzE9IY+cf4k0d17j+c/m+mqx/DhXhFV8c/yVCejm4qgTIsclEcVvesNdLKoADxBjKD4Mv/4K6
rwdqANmExI2IBKhrV7Rk2qbbuuv+m2YQ8gw+bwpsrAyK2ZD6WZy815CEPrq2Y0fnf8l8jCQL18ug
Ydt0h7P1xNYQrqgZFFFWvsgJpHDtaqWkZ087JY7BNi5GmXggGGNTv7P5WdKFZKcet1g9Zo9LHEZ8
ClV76Y2o72BdbI9ptl70rb1ZdRqficR4LPg+OL+7iaOgk/UGVttBK0CRDZYl91l8W3/NsgZEH1vc
YxYHUibGG42xNgwtdaHgzr1uQ4TfXP/07kwtEIC5Adj/9edtGytQdYG/gkB0Oz18AcIuHDMwLber
2nIU2YTIsn3fm5hvQZvFXTX7cRYYlq1Zf/k6kcYlmh/kKWv1MAmWJChpwMx4Dx5r302M1T6vmHIk
Sij8ieI0XDIS776RizTFWep7kERRbGUyeynyCQflJ9H/jNQl9hymphTaBSpSNB3u2hsRdZiZNZrx
QdEchb2Dc/XhRL+Zmdz0GjDCHSva6KsWFVlZqZ3Lgix0EfJYOBEhxI0qs/Y1FRmIVGXf6jzhkIZV
c4G+So3VR5fH4IxrS12H7DjUplRNqGB9QvNEPqfzpmdAsJ42FzGgcM3e3rsYSjPc+Ar8EU5YB8f5
J6/gPoOT++tWTTr6ADTFL5LrE4vOoqP5slqiL0VhXkULfVaJvPcx2WURiVMY7Kynw+6u/Gq8Lh7+
JcEJ3ZlXjVHbvuFoBU+irAeS11tSAHMXmKNOCHcCZ4AOvu/onwbKniOhlkrL88QfKRkpWZ9A22Em
o6LLQei6nMUky8TRvvM1qBAGspOJTF5A5r6TmioiRMA2QBWXFknOemPs7iFhdtGd4ADJnBqVrctM
m7TuHwym2c+yduY20a8P5OAiBQS5ShUSfV/JdjJtYxFzPUhY8gnvtyB345gJa0aGspAnFghJ1StH
irPHtWvfMcsyFMii8Fzz1j/3tq9lbTup8jWOjxQyPHOQYmunm0sc4/chhJIkqMxiISgWeqq05XCO
OETPp0LQygWSzvxgMxrB7FN3fB3uc3uDaRcURy8vQTsG5F5BVZ87b5g0D8ci+J30s65yRHm/e21N
3HIarlk6r0TiKSkQhLXMmPiJH5xXSOl62FQ62wsPpNxoUw4JWeZmit/xCAmybvTGDcrMBTPt3YdC
o4RMJCpAhbsF+iSfuJUuAki6Pc5xhfeNmXIigkX8NpXPa2J+zCL1AbFevkUdO4bn9C5wx/nLgO5x
H3XzRX+8oMvsXyWvnb98e9ef0KZcYETXBkZqny8Ps8osUXof1vqW65hDFr6i018vpt6pwx2BGsEt
qc7veVe4Dlmye4c1bdDbRSYXBGH6XB7Fhtl2TLGdRguahRT4lTZkfy3M6d3ZljLP5vkRTyECvO3O
8f4D803CH8apjqjOHMO29rFMbpNSAjuc/gNlnmJ8N+erFgOCWz2buIMvo0aqp28zKNg1dSZnu+Bj
5+75uvTQvQL4AmL9MjbCQEVShVGVHHn8u65qXkb4xghwkioJHzhk6x9anLhi92+1nWokd4UgNAHZ
+4zh7GttZ1Is/d1Oz74jR2Jh1XkvcqEZ7VuwMKzk2aoPCeLFRiXnA7Ljx1sd2WoNZguVeuOzOoSN
K1JlLggTWtdEfhTikva86LPhwuD6+oppXgTgFiWhzbLmm42eC0XxUpVcR18f/7UvthEh65+jLOTS
LCPmBwpad236PvLz61cQQhBGbpsK0nSWkq6ZhRZGC8cIo3ZElWrcRfFdqkkXpNAfKg8ZJFBemSUS
k0rnFUIWpY5+qpD4x5LYBbPknx7KTtAbPbYJbV8yWfPr6LO2/xDM1JGFm57SZaQVqbWeWTUzZT4t
1/ecDgEr+u/I3w4AWkX9ZJGDezdgJks62/P2pCr3ZBWAdjHdRx2W4PNMRq8giXz7GUwC2aR0jXCC
S6ANIHVhkqxBsv6C8zHhDUF+Hb+kVbam2VAR+0QhXYeRytOClAwjLT1YDcby81ybXS/TSUuMO/eL
jNLfnrYwnaJtZiek9q0H6ws+RrKGBf3HdajqTozy/2cDlQ5xNdkC2EFmHwMvieiZ5yNJVBKEAgI2
QgtxFgparjONB2n/+X0FSZHg2BgwzxB8xA0FlSLGw6/5wAr6R9rYqOiKaEoVunYiFxu9lmpcO4+y
200YHK7RA4srjCEiqY/gHM6MUy0OOBIC7/pNPiMIN1/cxSH91dFk5fS8j4ghyS/5vL9OjePtrXFv
yl10ZJJYBIuFck0EeV9v4wFe7oiqJSYj9H0c3aoAG7K0FcafYrbnM2OfZziyvxWzMpyLzzFhOnd2
gDTnn95yjg1A4DgxZ2/ROkyFxE79pkfZNsyp/A8SVRGTYGFmBfnqp8CBnBrpXwnrTiJ+hMZdx9CM
zIb/WqP84ggqfXxaBWoz1lHMSEhlfIE6UWacTVNJXFB6mAD7UNuQxND0eAJtcKCU736WfFiDCyFm
stlGxCxt7MXEQum6he7QWwRgqiVEJCjqyLuqFbdWV9QAqSYlOkSEXEL11pXmXyQ19uCIypXT0JOl
bJbGylx7mJC5nLQI6HGhFc6hCyqTmKc7I5QV5N3mfP83FB9107Wyu0l7b82ZZvMLc6RFgCXc8Jxp
zg43WENdeY9/tzYpRPqlQeCnHWj9xhzD0RfMEZy5jE8Yn/iEw6bF5khWexHu8xFumB5Utp4mw2G2
3rFDYMmm6HcSJtwdTayhL10tPVEgG5zzgOpmiDh9M++MQlrWqSP0nbzpbFoCzxJxfKRpnw9BUflW
LBMX105gdbumVjdvNrwc4EyDWNDJZEJVt/oJo1jOcIrYaFn+fbR4Qj98DdrRP4QDpVCVWdMxFxC+
lFH7/2ucTs3iq3XsKVdxyKAqOytrg3kp9jvMT/qaeTuIzsE5zRJok+k+sDwZgGINyQ8Ka1m0pMRR
CaubkjFuB+mrPpKWMxMh0R5n39gLUku9U7H1NSGqAT40G5pVBvRh8NBOYP/XolWVcqdOTwDrRVzd
QcC14rs9tgtXBDWD4eEdWY8TM2oUBItiTBCLaf+m/oDHRIfhn19RodU39SaEZRfHVwWRcjGHdwy+
8iMk7lqdq5kqbt/ZM68lRKt4C7SI9Z+gs5XshZ7oi+U/h25YxhMSmTq6H3/eJwEpRc4Tnl8ZSkhF
fTbH7e4LsPRG+w4Pwiv3pEziMILw6/rHqOJjrec4NPI7WAsXLHu6Efd+9yrmv01DDmO8SL8UQi+u
g87dWEAXa/NAwi2mX+V0hikSg4zLtcriEPBFijFHbSGm5bEO1EJ5+nlzGSatNX9CZ9e7g5ms4TDR
Ueu062Y7H15ZSyA7yL+XLFtUHsUcqBtuVJaTA4rz2L+O7rE4HpuU0KriiY4b3bSlxBoagPRHyM22
DGpdaOxr47Foysv637hvaY2Y5dVTJY+0cDnQRPv/w8GTL9OK3py2vbs4Pi2vOZ9Zm6eKmzMxUQ7t
+zkUvhR10GweBX/1hEeQYJaWjDo7PM6IBSMPNsQsl+LGHm1CtFML53GMgMQcysSLW+xtVJFRcjmg
2ptzD9qsF7AMPchmShCRdHSX6lHArdIvCvCSTuyNlJ4UiSptie0ItlwulxUjha3NDW+GUm0t8P+4
JjWtFHkgB4wtK1cHQEqGqiVp+svJ2Xlye87bdWxOJqwRDnGaZ9W93kM91k3RaWHn+cLKdX+6/VOs
et8DjHxwRivfWHFxtC//QlEaU7/XknYkgtpUzl+8DXkhELvIE8nDnHQL89fQgQ3eSNsmuRczzIPX
8OntE3l9vLkO/oqoMoa5Mqn9GQknQ2vb7vQeXNpcqRLiwaeP/t1PoavT0jsJwtVRjjerS+3HldEr
XOpQlwfhG1xbJyXq/3TvdBxum4avpRnlMfyTmEFkGJH8T3phEbqkYjXgevPb+6aPPFxhNcU2NLOU
7UqOLbNJf3BHkPkqlHZNRWT6poN+ZHWgXp9UjWfVofq2pODAKDnDXJPCSJhwLP/iyA06YGwKddZL
z96TPcZO60Fo73xuJ2qyqoeI9OE2YTHzMJFNoAAop8xxi9P9wyb0s9Ie6emP4KBAQX7xoT3Ck2HY
/XuYz4fWX8qXGE7Y4PoyHcgXeB6HheLSZjHN4apJ3RyuyHC/BGB5Sv/zhksuGESl7kJmugvQJrlC
+tKIPJHwoij30WS7C7caKAkeFVaugQrmsvKcurIZA5pUFRWqnLlD8b7rulTdMpUFyEp1pkZSrIyv
gGPyjhiX7paE7A2UWjTadmjQI7DuGMniNRDHlwZQfP3YixayKzl0ZTaAYy/Fzd+QNZT3w/d6btAy
QvFppx+IQuIbjdnvit2Q/w7V+d0ot3oCBKpC5EPpjSoa0bnV957ORazNYfn5oppz7j5WkYgGvaU0
bJy3r7rKMF1dxqQU7ri5Ets7p040SIzkhWWyQlOyvtIEPBKIR/iipCyfEk09OjFwG4gsdrHJnTec
VUz5MBqHx161AA7uRlFLShC3odPV88Suy2rCZFKnZOnCD7C1XqcxQze7bLHxqFeMdKICLLQrZWXN
ly3yKzyJPPPVf3BZs8Mi3YRGOhxCm8zwKgP1ongqPNBbCH2VjVOqLnXdyypImMRxGtSMEGcBb+Co
b264zPj6Qcq3YUauukhE8G7wXeKvu93ZCcJFsxBIcVSa5+kiT7ghoT7JP0LqsTIvYh8WI7C62/DV
lP8pUw2cO0yWy6S/gBCCxG/BNH8Kafnn93sYcjZAmUlSaPJ3aX2xTqFpO/9GHumKwopNrsby3Ece
fG2yzTzLELdOwQokO8ErZd1JvkQq51ryko+Da6NOPGBgmrReg7wiDYhIq+SNWgevNE4NxxlIoBod
N+3ntUG5ddLGzS+4jkMMoaaA783GoseFEyJfIF1GQq/8bVWGcPWFMf73ILmgVIyUUo3JdZQrTGpp
H6ppw60nhkctpcwfiBxkD27nRx667JN1XSPUR/7ofxxO8LCRzdwPJjmP+C0oTww9d4Gjz6I1NHsj
ehVrCkziIzcIx0VgEE2ZZwYi600C/U6Df9df0P6lWFFskd5H2eS2ovMGEiqMi/iBUBtXq0ytKbDi
t/JH9/Ot7G41z5IGG4tbgu0oKjT9j+A9c4Bq4sNjGlX+Uyn6mSYzz8UGRz70bQlrrA5cJMX1RERR
J/YxPpdRmjGECm4dxC2hNQt6EdQ+L3kP0sejmyDoV7n7MRVmE327xjM5YBuHewwiJ9d81zBcR7Uu
suXbQs27iDAiAXIdgl15ELZW7uYPOlJ2nWd+uQkqjmJe6Q8jdU0BK1oPATnyF0yajhbYh69frAnG
hPlHHANnRezhhqCkiR68bzOKol3V0kjHor0/AqZzeX+hnmnOpZ75Q+YpWC9D0yClxAXp7aRVZRY/
ZBdCJJUi3yqoILF3J1nBQYp+96Q1O7VmSXPhXjzmqjthCQ6oJVyrZsOW+kpgHsr6JiMVR/GT+0wB
HBuJul1Zk0rdBbrBGGXW+2Rk8aVZ2vo2J+FPYzuWucn+em5yBXsYGKLf7Xp1N4wDwJ+1llAj00Mr
Jx7250fg/YtVlpf6zxPqddK8qgpr5Ka3kpxNolCp1MVc4MA82SViLKWnh0StpBLgDhMUYN6jQ5hP
22xErj62kK0A46MEc0Qf4rxWuSAD3NpglcnSoRTCUVBTG09hVOsKpqLR4STLAOzhnK2xDSHRf06Q
1Dv92VLbKHL5xFOA8PPk2WueOcrVwknDAt37QFpVdjjjGxkwl0O7lXn49NHSRkYQtcJhj7bwspqq
7GF0SjJfmyEWVfti0xi8YHnb9N0wBVHmavU6OyuiZeSxsN6URgqL4HrNfnv/QKBcyLuqox3/QehH
jObrc7Xl2gEjKjJ2Oqs1w3oIel3eWIzoJpc1YTElxa1j9P3J+mMXXD8FVjhjGWw5xU/J/4qsz6ec
YrmPyvsLE1J9sgyx3v9ZQSwfyz+zsyqfCace9xFI1kFpkT5S2A6szsqCmfB7lo+0t+SZxQwKJ6yA
S85LStwwJDeWHC9OTMchZK8B9FXMrnTFZxPzSUzexbsNMI/rjVAtNyM5sLU0HmT9/LO/8M/DpqhV
YUfk1uGECCfR36Ri4uji0jM8/CBq7QcxaTFRG/g03I9q0S9Gl8NUWCDAHUEaT5DS/szEEZtlq1Zl
nphSG8bI4VNn+yLKvQrgWw1UnOceC0l06azDRbtvJrkN90TKjE3HCGV2ZRgtj/YnL0uPYehAXd2Y
ufJEEAxTOEqNNlxVIAKS6rmD3SnRUFksNFM4BY4b+/vSA4wPhW+xxcsRTJV4qUaPKbu7zFvpAuVc
HBDIwgbyXcEUSOriFtYzB9ARFmLyiMpAmWfUghnuc4qjaCPBdD+SaldnFHMOEHxu2RUEBbZEs8cu
JiSkzisKgGGyLP6Nw1c4gTNvTQSxaQLoHQoKJarYtS8WTVhONiPRTHw01Y8Wd0GVDC3Pu8zXeLkd
sO2ID+MM3hNn6/upyLIb76mZhXCGOnCcFdt0II5NpuwLKxAQLWu5s896dSMmkS5JH11c4Zt00HsO
KKf/wzUzI6gYWR4RVyCPYo7HWAoCXf6gnHoLv+LsmgiTXgv620ZZ8bjpF4wW/oa2xD3Veu0dTNze
+w8fVRggij5KLP4CRhh6fFK1aXIEsxEzdLtFKV8EvLEkO2M5mW6YhHkok0uMWogeuxVHquHio4u3
6917ar/B8wlcB+HtVoFzO5pxBtfrYfdcEjfjkm++ONj1OXZx2/B4f1u78Pq3vYMtSWqTDwvVIw3d
odjNsXJHehVv+xXme/DPKOOF6tiR3aACC+qMWFuQjYdn2a98oGn2nWOIdRlZO+H9qrm9UuUQ9tIQ
wJRwTrZLR+Cqdntk0RtKGqcov5gpyB7QzFqaeODhRgVlLWmAPJL8RqQWeP7uB666HMCmX9CsTH9+
c2wWak9EyWP/na707nMXdN9Uiw2WBE8q8P1n0khpyzdKd/Aufi1P8LFwr+q+5KprrDBLkyXwv8SK
jLn3L2rUVRGZi3a3r8K//LXVlRmdFUIXdRkgDmqRX4egk6mM02H8V2vinJNc1vb545jHYSLFlDNE
GfMg3S3Pv9c/Y6w5dpMvMdWVuNT7xoqsA/Nn2aCyeTVviHEpQYG5agAUIczaMW8/2iLkdTo9zVfu
YwemEYNWp9DHVo8awwD9EKz9WBkGO0Dt1lZTL8fbUwrZ20mVPlRMbufbp+qzH+HIBhVkRHw1ZrAF
u2bTMGEp5rqGc48Cz9kXMftwveFtnkFdaD5Ae0NIp258EFr5/8GNEDxzrqFi2mzMAk9NVtFXDZ0D
wius/ZdOdwPkfd4+8Z9VT9Sc18oMMHVs4hn/IksUcpWkh9hobzituyYwZHrYPkH5UdnjjgxUfUWH
UjpaAfXoT/BM17RjxBnnUloYNLdweJmnUcqU3s/0AzLlBGuSYoGLLZakGn8NPHMMcMT4+YHJqkGp
ti7KdBLZqfkhUwIs6WWAlwcqFrxlLBRnpRdXyuiqtTahisOqVcKWPqaOt/B9xpOSlmdddUGdSyrC
A1o9pxNOaAfvjs7MGV+ghtD3KwZ4Pv2FVGcJu/Qs4zhbBh0I7haQNhB/FiC2oOK65CGfS0ZRcHKh
7lJ0qNsRVzoIyj7uKua2ruu+gnqYdso/eI9kK9bYVBL7Kf3xHTMd2ZLar26PfnmqEX6yB5JAYiUB
oaJF59sk8q81Rq3juxG8IUyXsEx2kSHx9ma4TGDSxh0xwyV2K8E1+/tWHr9ZDUtjLUsQRQE8vvUx
zt2bnUEhFz3ix0c+DnaEpgF3f4lM28cetDP/ThGLwdVdRwQL0dpBuw7ye+fZb3z/o+5R72B+mpZ9
1zXOOxcDwUnxwFahQ7cO1wgKj6eS65dVtaEWZOHnnPem3JBz6rWpSPAYyYajOFji8LCbkaQX6U3i
ifSeA11ZCVwpQ3t3A2Sz+VfNIHxhgdKEQ1rECOifUWbPwozIZ1uuIZnOGIrr0a81nS7iZ8G2BBMB
Pwjlke3xAY+nevokW3As9Q6UIigWomUbG8YlnLQ0Dqwutzjk56ZtPZN5orGqew+Yu/qFTLolqT/w
5BlqQz8fhSGB3zspcO2KYMEA/7EKrCBwwXprbP+B5amNv1Bf/aeY4OvXwXm0TyZmBtxkQwv4DsiQ
QkUsSnIn4amCBgKL7+/MjzdaP22+AaQ+1TeCzMjQDTfMjS9N9gl3KszB2ZYZiPJwbaR3sxYVf4vJ
xMoOyegMq3s+rLn86juVhna3AY7Tpb8q6PaX+OrrGTddkb5HnjBtPJ5ybl0YYGliYt2mWB4cswVT
1PBgDfGzEI13PCgv69Cg0dhONYZ1ZNITeQuMTiX6wO1QStfjvUyJDy3n+PTyrZ1huMcxU5QfxY8J
2gg4V1qlwlkFRwaO0a6vHLi2OfLS02j0gbEopI3f2CZ1aB04Yn8c3wdpVAfcnXrMCSZd7eglUr0z
XaW5W95LaykopHgz//QMk/ptKiSo9+3s2hRsp2t0Qp0CEIksco06fLoLM8IS1zD/Zqzi3rFhRa21
M5JxOqpDCpBBvOGGvfv0/Z6TrJtH1i2cwWtR7dp9EhCDJ316E0Mwa5PJJ60MdFsUnIt8kEp7GJp0
S/WwkE/3bvZP36fqMtuKDuvkioVKem1SLzZ4faRycwfFLhFELpbIGLEkjHbvpQyaKicfNUHsMzj+
/1zD/TZOnNRiyEEexFx0MRBeRzAfZDCcCynlubKIk2z5HCBnHqQaL0UhRfr2+Zgyk6iAdEzvtvIY
A1XJvFH5kLHRSRiTmK0+Zx8Jn/fjr1fLp+1d58EGsTpc47yUuA2qMS4OalrKlecTH6pWEKdluP+F
s1okP/4hR6tRQXtbowKarJCoN7ReQNPPJ1hCjBh9iN0NZq7rWLpFcQbzzixhSTM6ij3Fspff3Tjf
udeOu0iYNKGxZxwPlz/8JyQT8f2nLJti5cJLQefXC3HxNvLeJV5cFATiMZPxvqiDSiW2EG3L+9pd
HofYtxoaVaXi3k6REpLG/9zacKVdSARvCCM9OwWkMo89SS2Xb2NDCmN3Fg4SL3ssN3PSYrm2nhaF
VieISA5iIqWoEu91nwWJw5m4Mw8ZKiKyt0FAVrpUABw4Z42Sj3gFf3TUY1aNfcEgiS95KaINwoqS
HFBtf2p/t+w7fFvUysXngPwf/kAbRtya7ukeiQR6/xE9kEI9umBlq6HAKlV7mkBwOKxglF0uFaeT
kzuFCe6uetJ3H+vK6dUJtmz60+8rUKz3vi2Bdftt6pp08XNjpFJ6p2bIjPE2TpQd1rwAMGuPzf/Z
DBFbfVVoDzvHxpIBzPylvQxBGL3ip7f1JMdmPa+MZYj8rJFHVJQ9XSjlplfvKyZD0F6Wxp/TUJFq
0t+eRkwifr3/ZBBS5S/H0JOM+ml+34JkOoFAQzOW9iD4r/J7a6lgbq+f63KeCeAC2RMVQcnPQkvG
Cc5YsXiyzENPjtcm99vkbNs3AeD5I2GmcyMiyPsZ7A2IF7IT8oSnOBly5WpJhFxHIYgaDsVOak4M
RqyK+0f+6nZM1Exg26r3fnIXxhAzbJ2RIv/9pXl0/LpnzeJuXT/VpK0WCsBUCThMKR47KjwNHVq9
4b/OfInUVsi42AJcIa+8dv/vsVePcu+pCAGMzauUUT7FVYa+BTUqAb3bMr9PyTQV/S/XnnCX112f
O2yV6oaKjkfMGdT357YFvwim/eIbSSjtk3CDAIlcLw8Kf1SLK5buzo4tDlxO0JrlHROXuMmKDlUm
26uPiS0oBecUGsPwO3ep4WLKF4pRvgIpcwd0uKNDObSLw5GB4b7jOy5wdIN5FP2W0zkEu++qus1A
zLYIM4T7PY85uyIWF+OvScLA31mDmN6qbQd4hNu87eY8BTrIVJWIA6nzgZE9FrQVLM+3Og6/zXyH
0zaLlKN/PXH28aS8L44/8npDoIrRM46mqXbxbPyFWifkG/axQugwlzwvvogIgrLf3nN7DH26xpbI
GWdrGslgnpoWdqwsJgpJDE79uTrcRXMfmz5OTFX0v28sO6i5RblZtbGoT+ViddAzjgkc6NuwWlpv
i2A0nnYaCx/TMreYeBSU39k6kz+dXK0TQ/JhJI9qKHjOLEU6sSyAslhlqjauErwRHAYZAXfwE+BF
OTKQacxzB+1mdrMXOx+5+k92uoxvLO4UkkbM9FUAuBd5u3daldePWtfkYcikNBG5wEyCjSPS8H4t
5ZyIP7df2lp0n32XT+qV3c1qbTmqT06INFjymUMMBA6tQ3vbAo9MuCbDlH5Px0KCqX19jVs/Djf7
OfR/d2dbrMdlgngbTQOvzWrkZn0ioiKuDKFONDag+j0MkYSxsPUMzcNvu84xDcUyj9XTva+mTKyP
tZQqB1FBu4ODxXA+5BBhATXSD2MoxNNyJuWUOJ/64Cn7VSHpk0y7EzrdjV6vkswYH6Dfssi7cM0c
PBY2uxqBcfyf1KHE6txfbkg2sA7nKwZjCGl8lC7YipKssGYvRIV9TL0vyVjNZ0uA+w6P2neVYN+B
tXWwDuHSTxcButJ8XTeekl4lm9/LhiA5H3EkqzylZ6Tpp+drOudhzXye2eoA0YNBFPrSYm+izlRB
62qwO7WXC/Wry88Pel70AeQ4kjbKdC+4bZkwldYtMT7iomOvD6O/Xazd8Z2pNZDQtZfhcCadvdrd
gOwiaB2Roljorpep5ESWOUyzqhgktwBkXVL1akTYcnRmqAVTDM0VEt9viv3qnuSFGd/1qUJQ/0Ln
lOpkREADhjg8tE46N1jXP0Os08isxOroYKk+blZVQay60NfIQhfjgG5NtGqAhl2WSTvK7otWbO44
dLybO8F9ChzawCd1CRdBqev7hG88zOjSpot7YP4hVmOJgo3WDq6LUaEREIgU0xgFUUQ3b1lwll7R
jBEDJ/oQY3rMDShqNv+Vm+NUyPKmmMJgceH9IfGLbtEKbYUdGBlf9zXghNGYoNBQ+xzJgOAHfoDD
5T+MzuNwNNbiaDBbmdkODR+h2mFwAa0EaBgv990TACAtp4lxrRU1dz/u0p3106qanKHqA3i3jWpm
P6ZmwiGmqN4jc3ofthEhQq6tsJ37WkjHzcRxtN2erWtKNYij4w0XMI3bg4myY1hWOrb+CdaMufRk
KkTSyXAu3ZcARSisedAhy1bzmJOROPOLrF2TKntUSh/l59TV8soKyM5zjTD270djsSWNYF5d9/Ul
ytY8gxTlNbrteFzobz+toWbYaQT9MGiWfwt/y+AnuK97VtcTUPCLhA5SLKjWoIDA5gUb2PkR8ETp
t1oFnZnrrGSe+N1MP5AqCG/rejVPqI2ZvaRKClFdp4tOy2WZHQrn2YvwHoA7e8//UAK89uaHTv1/
wP0qKoFtrLbY/BJel+1O/S1zFpBEUuN/6BGXC2W/HhZoRtPNlHGIfr2XQgtZCvioZrUka0YJXeSp
1zfAATNANOmSGLLLFwjWhR/cDWCRCI37HdkK864VnJ0BJv5ZUs0HhuFkpdwXjIprFo74PdG8wYYk
qDcmp/2QIh+XOains8ATuCvF6DUN1khzcZdYVnoqWV2QOJsHImigvZyAr7h1so8XWItMT6sZMzl+
8KJuNO0GHWmSGP0QCFDi72l2DnbGnB/xr0gGkysUriz8GkjSrFv42vmJuPBk8h+3SXKDH5c5KtdJ
YWnD+OtKMx8KKoHj/c/YOaCCzp+Y+U18wXEXmp5sRPMusHOCN8beyDuGNcf+LlOyMrmlQB9/GfJc
SKaX2y/mpg24q+v4HwrgUavkOwqayjLtyIgf+J1hlpM1BOI/7T6L+Dh9h9iZAGi7XvO9IGl46Aua
ZTFzuQR7O61a00d9UqhE2QKwIpj+HgWjIRFkDbPpLZb8DatYEyVOWid6jHTlo5lpXBIFpilws49B
fkg/f67yrOagTdzYr+YtEHt0iFO7gQLCRO+BH7W14rDpZYeu0DVzX8pXDP6xrDp60hpPrsduJ6lg
NGb0CL2xetWjy+6VuY3/06blyExa/qkC+zXgcsKgnDJC7rW5TdVZTGtzeNTAsDR+hcY5+pbl2SP5
Re0yju4tyfuHeuFdE041KUbFUGLBNRj71wFoFvIIQIWBUd8J8txpzD11cBvEctjv4IoRFq0iwi5c
sPC5YnkzPcTMVgrSdGy1QnUGR+tQd7g6nXMVn6ADZzC09mul2xyYDfV9miN3+gm30jalZBx4Yh9v
w0zgNFgjvP4ylKlVN+qb/a2/aOO5A+yTbptLzYNsdIwzF/z7wNkPqgIxVQzilDtipDv0IFtFko7v
oo8RrEHunqKjIhgC3S7EA3U0DysxE2L75VYPhhcuBOkeQEvd3nnMuxja2dp78GPhOfA/J9gc530H
288q3gqZKCckDc5kDLQlu40zl9A3pFd2RGV4ZfUMnOYLo3KVzF6eZYRkgqK7k1nn4j8etBgWFdeR
PQpPnb4/0h6lTYiBnw+IUkKUlQsWyT+01tcQPF+rSuE6jG05cbPlOu1AmFuWAAadsFXo8rV63Q/2
5SaxkpuEG2T+fB0lHauC42ZHrpRctzKwr0FRGuhdw5SlprSumIIZJffS0GwzW3QDlfsl3UDZxT3H
O4m0+kQVv2qb1iJHT3HqrnekpLOwKTl0NsOAzXuipfueglxW+BMHQ1NiZpaGGWmQOzk4QGaBJ5+y
REmbyfQbvpsuOqNTzKWesQp6pN9f/+ohNEoD60w5AywCSCc+phhF91ywjkbf051IxVcVnI0OI9CE
MDNgtc2KWTWfW7V1OeE7Dmlg5LyUApebWLlROk5ybpQgdknqdVyPWLSqjkxRUeE2I0c6K4OG4g9Q
oneS33WI9d81meXb36INwYufJEkeJMu5GMJ/7Wh8SF6VaEXLHlQR66DmWCwJnlV6418pl9YGzm5k
HZY14ptAL6Z68YkNZHAQoPWMhUPibVF9ai2nndxr9OARb2c5juyr3lrQ2yDEPKkNeGxrE6HjjDc/
Rhkf0gw7g72OtTx9QJKeO7tlxP5FhfkESG2eM9tX0KPahN4xszZYP/nyIrSyZCS0rDrGFSEC8Rpp
ReIurQtfhA8D3v+YKSwqYCuBh/YL87i4DSkbTADTcdDIWiGOGqTPipohvBLicIvioV3xraTtsx/Y
zu2++f6XhAIuHKNC43lg79OqCEw66XG59fu0VYYCleFt5EE6PnnRVbuZEtRrivP6/pM2JJ8Zi/9q
+ZysA8ZkTGNgWnnrXwg8naPWXs2wFLtHdcoSOeAW14dBshNU2TVumh9lMM9dhd5cocE0B8tm+G5Q
zzgeo2CtTPzbEw4QFgkzpvZ74QczK8PIsbdKmNmbv7gg8spHmz4uhQJZujb4WDhfVlH5w2vQLyYU
NthJN9bxHPmZvxb7bkDlFIz1MpU1DS2OLPR7+9Owy8ewUu84aKxFD9pcm4AlpdQMucdsbp5ijEoD
xjsXPvpikSfAomD1nq1K+gbAUFRJD2xTJymcWmpWrMOTC2kXjIpGg2gNv8KNieCWjctkso5PQ1+2
k9hlwJLSc3noBIa4GibBiWvWNYxHu+hrniW2yQYZawk0YW2aN3EyVC70O2qKU5lUZ+e8QArOEDZz
oztITgv4SXWK0fQ/h2oeZiaHdgtZt0e/5cCwZPyv3CTpP2Y9YsHhDB8z0Pefc1//AWpbZpIGxIPG
9O2ERFlJa5gBDBvk+RGhmlapV5TsCfQrS3b4N1rbHI03tTGTZY9OhG2do25oHrsjRZTA/oViOq8f
5aD/fBYBs3anSqL5b5A4PUn/shJPdI/bKH8DIx0bAQw4yhLq85mLiS771DZQu/4VJ6tjCCjdj6Jq
tDwYp+m4pXdvgtehrhgkJhqct/vqlnyfvkxQjLfBEbsGD622npgBo2QGKnmAzaDjhbX+H+18aNrm
/MZEkt8O2FkPdOA/cOq9WSJyqLLAzDdLynwzzAf6kM5txCGrjx8UoTBVkX6215IA78KGYewUGnYu
jPEd3jbvtjY1vHXLR4p0qaTCDB1dfqlyBODhDZ7m6zNesnFcix5KhRop3GwpoGVJDkdjWL9vbnau
CxgPUHiX9PN8UM+hnH6QPLgTOyFeHptee+WMWYSu1OCilclop3D/QAgLN4f7nAIsaU7fhLTvpC7N
gswWeJcINdWSbgbqKn1+xYobZ2qGzj3EBauMajsTys0tOZDIHh/G3gvqnn+daun04lhVyPpMcVMR
FCHd68KIj0IPZkN83zWjwTv1+rKvvtZwwM6xdQT9gNewvQ47NGLpT5JVj3hWWtf/RGRXwV4o4HM1
yZveAmDH0IAgcOpxhtxWnLzxk8puy9GnNenItEo77zkkfh8l7VN1CCLSO3ZIhAAfO907q2tmy6JQ
jnpW31JNRVRVTlQ1SJvov7q8VgrR5iOoyKcLOtm5q7f2nK7dgLqPPNtSGqp91Mz+XV3U66vxQLVm
6dgDP8c7aOixWk0BMNCFDW3ja662h+nUhqkPN0Z0j23Dsyop8dI6KiS6oMrVY887WTq2PouvAfeH
1MbD5eA/aTUXBOMLS7cTSFwkhFIvslbYGsNgMxR+aNtnkpFPu2M6/k4ZH2vfUN8VT+X0n3YU+SbT
//k8kWwBvDXolzobCTVZPNeUQgQlcci5eujeAOWjyCYh29RXWVtLHA2hw10fbU6S+xlzwWNOpvFU
mTfHJzaw7lSQ6aQQWM/pMJG7AOzDnP40mV1Td/1YrEMfEL5tf21dFQsp1po5b8D0TjlEZ5h67D7l
MOVeguItx/dLVK94efXfa8z3E+9/M2z9zTfcVy2D0bwEiTWvg9F4VLXuK8eyZF2xNyRjQJRQKC3G
EgYV4TqUPBxOfsEv8NRFVKkhY+5kfga4b/Kgi3beVFfQ9+boeiN9bmdt+RM+j61SmVWI/+Odyvn4
LT0cxieM9DDYccbUnxO3WwgJBMpUZdXehaK68yoAWmiaSeoOmioJ+vk30MbbWmF7i0Uzvds4s0p+
KUIOA7IT7hKxQ3B5vL7HaNtbZHx5mBNEB9drCXOww2QDHgmi94JNXeUYbLx4iN4fJqH5PZkMCj5G
7yFqyoMLA0BmRRMC+vmEGB3b7BvDeI5zUXq5tUesuMTeLRvccgSxru7zuRlYYtB6YYXdItK0r9tC
NiNMGMX5xiriWBz5CpMGa2vfIakWtFrJ0y4TbUFXzYndsqPN1+jC25m2lGmEo9d3EwSk0QKRXHPV
G34HAIDm+B/ISOlZVx2hDNOMyWxhmlMUSWgRHAZ+3ZenZI/BcFDy6Rra0rzks1EcrdodTJiJmrfB
xPpAHiJYcrMk1GoJhCOcFrwctErPHnCVGmPEh+thjiwmPd/iDMEOe04+g2yRSVdVMzbgHnK/6kJR
cNPh3CKkXJnBreHvtLyezfX+vMeqpoXH4QRJH5ItThvWKtaf5DmLVuLE+ToLy9gQM1tw37b++ejd
oTCw7OWhk8cCpO5e/mAJGMEwPE6UbVxMpyGyhoV1YoUJi7/p3wJQ1vkBAXoWGYP98vB8rBYO6Yci
/gOu8Bm7KHXeEsQE0JVq9q8zvXBPuN+Rj2vzu3c+xvi4ONd56FdsEtqr9Kf4tqZdu/htTVpMxQnt
5NgeB6QC8mIEgj3nWIRO/+XrybiOHoL0j3ykO4+baVSH1CUMrdoRRHq/yMKTk/SASTu4EgWsL0S3
fu/VeQ1rmEvmJvJXTe+0v+lMAnFOdrVFsg09oDJTQ9XMea8ZXejEnnjASci46xI0HHu8BD/K53kW
4QgfW/hd0K/9gkkk8yhjCQVNR8OTZd+dkUM1q/MOZvf+uB6PI0NOloNXAJ/qV9KDc7Mg6mRX9NvP
R29CFa0yAt5C/VE8JmknE4pNKDR/GeW7blt8akNHGkFoSQ0PkxgkIQaGAho6g7oMOuzsxI5IoCOd
mZ8+Pzj/MRds3d4yI+L99JwSK5e+GhiJh09HxrjQC/TYG8yC679GhrYe0lqlfnZybF+9Zt6xxBUe
/2cCUvbkFgNbH0MN04RAg6sXUaKl9VuUqlsEAtHl+2Q3cEJYGzevLAaff6Ql0x2j873VdOQwb6ua
Z4zZKsM/TM5dQqSp+xbt1BIIRXIgejyywHW5e1Xt9/1R1iyFrXJ97QsYMnA9oqTFSPKxxVtI/tVF
MvheHwrk889sKN36FuUJvZHlNAOHDrKcSJOr3fuOnc9ahT0afhVGyyEZ0FpTkeXsEAa7acaNwqci
NnCI0NITj+uXJGIlOA68Dc3++LfUR4uTfKqIbptdO0l9zfJIX6ww34yB2K1x8kxCkJatIoDV9q44
KPgJjZLSq72PSVfGe8V9+U3w+sgqRhBSmW/BAGq6+NNKevVZ7Vlu0uIXjOWNUF9T3MEoYyd/szLX
x6KERNm27Wqj+hbuWC8WGrX+MMTVT0lLNiItvax2zD4c5m/H+zyT/lHGplED2aKFmZWOdF7FWpcB
m84P/x4mO+sASTp2rgfV0FcAmxgxBxV6WKMMAgX/7MqvY5Zl8NjZ1gyTAAKkbJixEZzMU0GYs9ye
NyexV6VQEeUIqPRg8UpEmMPLkn5G+eX5W1BDtTeA0rWDP+mzVcYqz72D/nK4+7XU0mZ1yk9IqFLG
drXUugh8EaI5gsiFO2VJayOKibqQp+7jkm71Ce0tKtMLf9FEilk/ulHe4sAAnOg8OwsJCkzLNKzZ
nNW06AE3xU5nplvxxNvsvncIwnkQ1Dl3yfeUNyFjSoUkMctg/RyCPEjCkVYcj6i9fDHNaNAMYvGJ
AbjtjU2f6i1tJP1rQJrcAypCm2f1KkHjsbnJa82QugXwCTUi9nZMSoRVDwrv7yQYo4fwfTT+OydY
/pU4Ad4Q6BAn92Haj8kuC2hnelb4zqtX1J89NyJmgqvLxHTBeZAgRQMTtnAtwRvXMnAtcUapYwYk
4YkhAYTpYotZlx4k8kIFxs73covTYRWNInA7GHWly2JmP/rbrHV4SCm+o2GZzda05fSYpNzbicL5
F/5EMCv9F78JamKMRrykROZ9JdsShZmEtyQP9JLH8cbnoMvEK/yQ7PzlosyKWXci5M22vgCPCMMf
+vhSHq+0ZdOyJkXF0aNeWBIWT8zTxB29Ov2e9VW0eX4HdEOHjnidxCI/uPnT2S4t1GCFcZLnu1uB
vILXCXIAjliH2jLv7vl31jzLZRHMfnV1JGBFzFZv9NE31eCLjnsn4tBeNJy9V99EStsnRR5pLdif
ym4pbXaeX8KNSl6kj4Ne6EnUJNKzX9Af+2VE9zfHHJRKumefaDgvOp3i1dZHuldCPAS4OgpZadLP
TqeUuYVJ007nmWWoD6mgHrQyLSuYYC+4ZogrWd4A2rWBKBBuSgBLKANoVtd1Wz58E3B9d2ojkkTI
tHjh3ejSKf4ta5b1NXodE07of4IwsXHvay5iIZ61KVz/MJRHsXXIZ0jfCbLtsT1/EXcw94ez7Yjf
vO64RfHauUKpE3DmlmftlyV3To31y7RAZ19hhPD61uH/tv84xwyMfDm2C8LNLisAqZMfhb6RKNTm
B8L1aRkzqx+/6CgIEe7l9xgOBMKYAGbNGtLetJn5dGXbQZwRotsDFqAf4w5tqaNNq0DirDCXKUMd
Rn8qiJ47DS4t5+HrAFVdfK07g9ZaOM6V8mrMmsN2mXR4N16xGftLyfeReW/XwPQItF7RpjIsfbj4
biAeru7/kqQvZddD75aMVWH7LzMWlJtOYBfq0CupE4iOXlqBH3T0EkB99s1REiDEMjPH3CSFf1dH
tUk5m39R2VGjFy1vl81HF+4+aQlkKCnBK2Cl15tefuQ5j8CrpFfOVLW52VIFpCqzEh6u7hVAeE+B
oKxIvPRvYC51ME15TTYaGqMS+HltAdDbwaHtV8X+mys/wlwDc7qWaiGF/7MIbzXXHJ7t/jB3JtCH
bmer0n6hEE/1W9uS/m5jgHhYIXAdiubx6MsBDlCWOMtlD1L7AY7d+SAllQiQE/BzVPTzLulz0OeV
Arz+Ddy/Ea5uER1jC1KQyYEfqHt7I1pleDmtTKWO9gDVWDbUUSaLk5qbYYBXZ3JOPlqfyQQx+c0/
vV8m1/jqurbE1RQOzB9A7XdZMjGa7/c6YFVGzbSXwEjABuUyv83a+gc3MnOrPpPxOJnTA8tX/rol
cnx3YWkyX017MbUXMshQgxBI7MKaY4ywd+lWsVDqOJ6NtAvRHfbPWE8Mc0TtEnqMEYYfoCGPIYhw
Vty1FR5kePoRglPAj+qxV1ssdcXbrriXlZt30Y+Ax+F0SmJ/6moHR0+7DtpjYu8XalEtxJ8R7glU
a5Zm3HN9kaT7ThONAWTvQ3thcdP5Xkn4RPIIPm7TEjiX4MnUY0w4xVQtmVJxxPxMKPGl++N+gdr2
aJ4hwBf9TB0ELz3oupW2AvMHP7NPqkdiw/co5idr5YefhnEzf9Ja+vtSCqjsuzlJJtzVUcAP6JZv
x7zCa6aTAmTbijnj2Oh0rubk+a8BXFiBkjySFEZPxGhYKg2jWp0iUfwEesZv/S3p9RkfXV60wiaz
EpqoiT8Wr93w86bn+L+oPAEl/EVxsIyd7qHV0GkzZd3KOhtGLiRIehna9sLDEJWEcYcK8JRX6hbr
mlXD4nItoQJ6BDd6zgzawR1QyAqJAVxxO3cgCs2V8Jkjsc9Ic8+IgPFCDh6tTfdsOHxBBiXVDOx9
HXsX3ZHCVATuYLzY60SsnZsFTgZnBYrK3d42pQ/Xz4PV+BV6VzYo+O0SDNj73YLkJX7iwNWeuvx5
0pdyxxidORHEFNXsF1ozXGqD2tpNsJHMkPSh7MEAsE7m39vyfgAUn/lHtp/MMS21uOwIfVhNMbzf
EIklDJAtgfi0IkoOVRIqpgioBAQAKdcqTPIhvAr+8UW2D0UfbBO7hV/GT48KT2E77zrPDnQn0sW2
EGjYxr3VYifkMylFCaE60rOUkHHtKjbIDHsd/ELJ8/Kg9LfxE7gcUIjtvOQbX5slnIr5ZG4Y5UM8
2r8IO/zrJTShfcP2h+LKcNGl3PK7DJb/kbC+MDVxGfjQVUY5DMREwFkxtfhs5H+bjZLX6gH340jx
pp6K0fFmNaf6xNU3nouWTvaze0YlFYRkeT7ki7DssuK00Kcq2HwzaQuhtbP+lu9LzMaw27o7I/0M
F4srWJB5+t7kXb1om3EM3jEJEH79rm+aPjzPIEaRkHc/Z/qt3eHlOmUByH0WNAAsqEAqKJ+BHYHn
ydMUHcorKEbYK7yEPxc0vhN/62kWxJF/1w/lFdIKKty9FenYiMlAKvQk/7IHdscufACifwl9e+Ke
rhKB9wzI36Mf3GjS9yFazVEbzoQLob8RARm7lx+BDX6O7WyHi+SYLscREz935z6efzhbDiked2fB
RXJjFf1EdFAYRrlbJKaqJFgkKdppwpPFSS9tnesZ70q7bUNYZrPCrIFLdgUnKBYKyhD+fG3qi2ho
k9JRMvA8o6DsJyfEcpmN8QHQd1V5xtfCZ5SL0ds9SFI4yhmCSNQqw0dBwXG29j26F8jHZAUR8OQu
PzALKOeNSeiJ9UAE4YJ4vZ/uTq+Wkv8G829DqA9wwB5AgaEUtCsY2bkNg73heyYLIwS0MPyVUYai
tHfYPCKDat3hnPQlg91eQKS/Yq8Sb/gW/ToULNq/+AM2z0RRGcw3Tk1B8Cdr0984/+epIO8Q2386
gzqYFCeMDc4P61ZupYjyrCjmofo9sOqH/SkYkfVAkQmbpkJ3Q6G1GDN2e+xs8epIoEK0Ytt5phCW
rBDtkK9fgOTjb/9rnJgIARN0NEdjzM/InsEusRC2kdePWpHMMAuIPQGxmqr8hSnBi5LaHHggnA5J
Q/pOlxSLLPGseU+l+KxLt0o458s7qANmmWgFUAJYHVMT6/ULoXOcrOFjjgSa6H5UtWJTTj07fMb/
ZoCC+wzAVjGH3yyi8LFrFWAfoUZQ4mdeHmr+UncozZFeLf4hyNRH7sYhNMq6kSxtDKBgvi/sfvIo
qGYMll5YvNysiC5mHpq6BUXnsJTcnMCm/nHHCe12GMj65adhQawbu1Fy9aqSgZCfnxoA6xKJQ2Qy
tfAE4dnEJBsNi6h1cl6P7k+7AgzDSkIuughs5Oig1KTjxTU++gP1IC4Qb2cSASS0IJp1pOzNbi/q
JUBUKMM5e+qTQ7utGsF8zSnsqVfZbdg/xNu/9iB7vNhzGqA/k1UBk5BZHPixgkMcwrXtq5FlCU+H
6kaS1dkwG6aJesN1t33h5D2GG2ID5AM75obera50pdFkBa4SpEHXkIOVmSFJ7iwFHK/YMlWCg9Ob
WakrDdI4TVvIwtEESwrjpQ3LML/xSlPBkeYQXyElNK3sE0s54hNqK/fvGkGafxifNh+9SJms9ITq
orlxItur5/IwoomiWyO9mFLYZSQKy5W0BpaPjRm2iqIGz4UkzMjiw3NvQZxl2Jw6nGY7ndK+tk9I
nnSdPgpRHmo6PPuKTBupK0VTViHjkOfV+aTeeckBkDq3GmSnX0oEQuDXxwAfc9joyDLaAA/vEvKf
p2aZzRBZBw0rktU/ZQuh5+ArSiX3aWdgwUQYs8j7U+hKu77Y3AcYl3UM9JlcWr6WT3Qx6KBSzsaA
JsmnMiZwoYaIgiJSdJcfEn9Pll9clc1h1c/Ji1KYAmcfE2J1tLoHEH8A9QRO5EQ652aLsqqHEadz
pSAQqIH0U2uX+cFQh3Ee7daTFYwh6mMGKRtwHcLJfenFIgoaG3tQKthEzBmdvME3qB4de+kapgem
k8Ph1zihoySUH23kFZ1QmRjV4aF6wWzU+kgJt+qiTvS691y+B5Hg4dWcawNNa6st5lkp0xAR1TGv
NWWz9qov3SpsyqAiRGJdtfip6Ij0IsK4Wc/NLwTfyx8qvigHHpl1IC6mjEfpeSdF0EOBXbhUd3lc
Y3HH4NdNC3yBLYhJxLJPL/JuCPtgBAr2qJH4iIowMmnNGlPx7JRdk4XNiVnr0wRO6TfJfcVWT513
IMnw2qs51X/JxNvMR7SdJZpsj+MTqouvbjEcZ9OKRTiT0SPi+3RmtXE5PLx5mt+OdWWwcrtbRpWz
bpI433TeyJib/2Rh+hr4BNXUTW7tInene5bG8e1b340aTSGWPmJA3ccZZVGdSjkzgmt2/JOaAt6a
5gqr1zvowhl5JFEGnheVOENRSplHB5r+mCsjzt7HfXVIsv0+SsnBDtqtbDwEusSPGYoiU83GtaAU
rYjPSPd/H9PPD2Vg0FZDjY+YXOErNBmCHyqOTfWBEwzGbOHalgB+jq+ovU8elqLjj0/T9gmAJHfR
v/ETC2NQbi95b8wxTQuT6+M68FMLVEc9HVLqwIujq0vBe83UpavNYpsN5xQdTPZj260B77pF9c72
OygilleaqKIgHHxQsGxEYKHKIuzJbwXvjNWwlDCm8p4hpO0puoYTGsN4paE/KcD/om7BAM0QvS0+
lErqlSwxqJaM8Y8OH2wlsh13o69epAD48h0n//5b0EmwZSW44sfo0dKX+HNcsSDIgka0HTXmm+LN
h/r1joxXEdt0t45lWJtmZ34qYMUreks2f7nV5hRDFvlxuSjWuRwr/6MLTlwgOcqd+UZD9w1o2/nN
I0nSv+sD2Rwi8sZi7HVxKUq7z5nnIiOcov0+kZk3nFh5tjcNuHTj/UgtvnfU8IhI7iieRLxDU50q
lfP3PhaceCSURMPJEwEjyrSEBc3vgACAHDY78bAhnwlel8BuI0V++yuxM3O7JfMiS6IS5PyiLumM
OvE5iSf41785IqB945iJ+4WDkzuPwKKRFx5Y+b93EccHje7YxezmTUZJd2lBqk9y8UpsvJ7rN8D6
iLWJMATNKWGZvSmVaoIlW1a4Lfa5SmrtlLKaVCabxqRP4y8j2D29HhaNIUFwwZKjFb8gkq7UHOgk
h1Kei1V7RCt/eI3YiN4ty4pr6FTw65S/K5oFIZyoEtFEp1irKAX5dJUSmU7mB8eJ3CrDDXbDq7KP
CP+e0HaUMMZ2zg3RQOgiXUMQIFd2mmz36VqhI/gvo36Zehx1oM8HJDqKKejskO0z0fmLvVgp/UsF
8r2iHE9LyKCNo6hvVWcdYWraiqya9Y6RyD8smBA+NelKq4eWSur0CE+ZG76gvl1Aebwls7T5HGGZ
UHhId+rHmW3/QsVVtkMMzpx4CLuI/r63eTJmLykCFdwLzRl2jqiib8jsL/yM+wGOfPakH1DaagF7
he+2H+URYodQPvw48DHqXLLWrTbr5Uy47ZCSH1IIf++Od7PIlQj1VbaFkR7H1f4wY/e0/uXiLV7l
Hg3gFvFxl5xjakaDgz6v+nMnOpu4JT4A/CD1a/Q8ymYqdythI9bC+0NzYMPB2TcHRLJSR9ngkrfq
ASV8ZeTvb5SCy+ae/nvUkbd2e7+zZ2wcuGHt3kOMDKOey21IfV1xW2IxHPiIA4HqBQsIHEShXThH
gQVJU3oBK45lWkbp2VWvGaHFWUOLmMHNDyqTNtrNfooTfrjdn+IgEyOUoYFIu+mTMT3D/VHZ25ms
BmfYcXUi+gBU2f7AaQmQCurQNTQzhY337wkgEiaiH8Hd1LnP+DeI8k32l+BhJ41o7ovJX3+8rJra
Yinu+q3QXZ7G1IBnBpDhrM8u7IQDI/f5FuAKa/JtZgXuzyD1WJiHQUDiexDhXjWZouudYs85JQwK
8Ucg4bXrqF8dYeb309Nl/q4OESiEyGUoX+QAbHIaLBervNCAdkaU4bMCEdtnwVcFJ2M4ulq18+KT
0LtN9JcZij1+Lw7cP709DwVG4E8hKrm0/Ecq/XPOvnfoyGXcuBrIGbmhDBKRDnaT/JoWRYI8f5zU
ru/wd83cTti1zYOCgMuIeP9kp6gUG3tcVhh3mT3tPH6XgEViMrbdU65rE6j/SqdqJLvVdVq3EkDO
BW8ZRSHY/RFbvX+FbB6lNkcXVNXLyEWJttu7qX8/90EMsV3wi/sANDiRWcaHKjZFZ9NVZNPy50oy
AgSQFGTJeYw0fSE2sxbMFNWgdDEhgMMBJuZ9KiGBYhXwo5Aq1T6I7HRQmpz+WyZTTk/de2t91A4j
QNhkhKpLYvwZu+Ox65Irx65ENFWkV489GtznQy4io5td8Vg8I+UjWAZq9jrbisxf92e6XjvJyKu9
yXmC+qfGpjbb1Hd0U2Ia3oenEnrkGqEbQgJga+sre+/Xl7aNEg7MhaQ+5OCNZ35o1Z4hSpcddLYF
n47S1QF5ZBbc4d8c4MI8AmaR/4BfIVPpeYvuKATIKvZ7/7A/OWJ3YUKa2Y505vazjbK5fLRzn3Bq
RRE3rnbGULQ/8reOUlCML5tOBZkadRUzBVLlbAJz/6uTFb41twTC+ptwBgOi+Cnzrru7em0PI+Az
OXWC7NtgqXzBfglIr52Td13CEPnUTvXGfBPXnxfzvU2j4JyQKOKYfln3cRVUJiAAEKi69eN/8QZE
0WWl7bmSSx6FJDYKsOJoEnzSpGjdO63Rd/BOhG0dLmwZcHY6tXNAMCjWSUAHZdWAKby0GT4YYhlC
4/vDhq/4NHT0G4R3+EG71krakJFShFLgCYiIQz1mGBBPyhkm+EgKZSpAnv+vJyUzMy9yLYW8tj/k
9GnjuurlbE+EF2edHEPEfFFsLcVujMhfClIBgmuTCEXQJMAj8O7SZ/eXeor1iBoGV0f8sppT+2xd
2ORGHO8Ld3yX7z1/csEquYGqJkM6uHu9GfWupt+BZ0WIAWRWPj76fatftZzqsJFYyT2dQeGDoaMR
2dUfBQ9EKUGN6z/vDB3bpP4MuowmMRfaMC6xsWOHj8am7j/PafkkLVXI4yE1LAV245DG7VJjQNZq
ovUcvTesrP3QtC9TEO05uQ0zlcnd+CCJHURt8YpjXCHvElesWMtRIMYRxiV+bDZjgTqwM9xIHy4z
bsbzN5ci1LHeMYYL+5d+SrzN6tRk2wKXZBsjuWZH2NzRqsuc48w8s88EtRZCPicoayuVtVXB6uRa
UBD4u1lEwP7BUknxyQpz61lq3LSQ0wZwtkwmRWLoyOGI0ylK2T+lN0tyon0TVasEa1YfviqxHK8Z
28sJey6L8TywYGOn+ycF+foNRYADA21EloY0N9UKUaciwzdAkAylGNOJPFczGVbrZPmXjXwhJJfS
tnf/xjNd0LwoqkQQAZUo7zFQWaPcO3DzcpiYLt44ecmbcFtnCPtwsWbLR5+ZnJ8spCSLccUvJLJ5
lvTvo+1fLGRB5cLno0dTHtDmtoHOiTRn1gNTt6QtJJ/6Q448ReNlApYMwIQhWGkRH4U8nUTTstbf
4QU5tubA1ejSE6jrQiXdiX19bHyFZ+jvslkFqGUeM6T7wIFwEfj5nnU3tUqZpUMvl9LZfzU5CJ5k
rB343N20O3c87sxA0MPvb+8aB7zCTvbbl/ElVSOX0ybqPu/iD5GZsUCGGH28nAVJ43HMM0o5Krsd
DyCYTtCpD3XNpc49iZ6qlQmdJGj4wCaHOLXyNFTzlGlkQrSBtYvG1o0OzxlP0oHYFj3QA+9555UU
EpCaBhMemu/v4Wfz8D2f6ZuB+YGZBr+d7Y1Wuj7HfOeBF+xk+ucCvDarlUIrJo4GrF8evHLBql6W
ryE0mFWY9niIY1tEJGKGgvyfKlnYsxtOlr1vQyiTb5EdqVl8ZdUDnHP/xL3oz3KbLN8kyK4+VVod
keySwcJaf1ZiEI9MOlNp0gqODiDmrec2PNRbLK5u94nlqIiQmPFLbRY7mILZ1AS9WhQ3dmas+Cp+
7gUMZO8l9PgdVPZpGmS1xKDKGW/iS8f6sBw3awNtSaYiDMqCxgsDMGy927PTSRq0w3nXywC0+P+G
PnLXZJOiAhDSGJ71EbesIYF3sN7UZ/Jtop3fJLbvq//8AIoIzhoCCgauVeVyt/Ttm7wZSEExQ9Vv
BAxCJXHRH4Hz8+BToqCGuuAJK4KNhOtSVkuiYBy1JUBtqUfBtfRgQSFRKMbgXYhjQMSgMyT2T/bm
cmXKe3TWPckuSUPCAIHlUDJSmqyHvhO1quI7zpFIILASZ+p7CDSMkmqodCsfwc/BX7Dv1944Vcsz
zdv0QIfysPD8eWgAgMiIfplLBM4Uwh1vpZEfv82WOGUFnqirjdaXPepQ5dp/FTFyhja09JIRwiVn
JyEsC8ZGzhzosfzKlPPO35+6VhWCfDwzAMOWYTEGydblDiNJVi+mgkftksol1dfpEqYHBPoz+/kB
gGkZC5K8JXdQz9csFSXXQhjwdkBr1i0OVv7R2me7YYzgeUmta49l01tt2jR8NZailLeVh++kxQmf
m0cId5+W7FRuazAzdg/J2/GCRYrHaBaoTTgmIfocplt9M59q3+k8OYorKs6OMi/cYaNyugKuPf0+
HWYHg1G9AIeJKwYRgy2qiDThhAkEDmEBzXtmVJH6h/OWiK2BdMcyKXD1wwLxU++2sQCzxjXakqXO
K2vWC8+OWGDoWj/jkOkS26v9o+768tNvjUoz0zrGpU4rleXTOjjqa+qXPEE8IoSFI6vbFz5FhEWZ
53rIL5+42y9Yak+C0196XF/3vCHd/AkjwbuYRdFyMqTkMOrdD/8bAY3a5b8hJDDh9IVq6FjxzxY4
sJRXfDsH0+iQ1TkexRXs+9mEO/KmlXmkgz8yf7btCt0ZKYTVdlctsQhSBTCW8+6id01uHRj4lBgi
npOD5bZ0thMQpXwLNk/vtr5FDSN7vTKayBzBwAqm7LWzsr9OsYSgvqf5TtuQIpqqo42dCZZ0vrGk
NVAXY4G9pYkx1WSpAFznTmlXHTpfdPHewfKZO9mQrk8khaxVSQNwbN5ab/s5bNtFA/voq8MDnX0Y
D3F1YwuNmofvnNbNz6T6JfvHkXYG8zNv/f5sIPcfvPxbVQWQS8qxXLX/kan77ggvLM7PTozpEutW
8rF9yqF+EvDzZe9rQbISFFw3s8oyhe/3FZ4ZtKNCNfes/CpXWG3tr8AqS+PYP5rRrUUIJmxGMlDR
sWaV0apzjmJ7YKlJPC3wxWjroTX4G7iG0n0/mlpHBMB4c/b2vdIVFwCQAQ90kxplBeX0bvoFp6wX
75gNVYEcqTjoUWtPsKUESs2AZFhVWI6xEalJ1kgHN4JT5RQ68BCchtY9DNScf/t2ChCQpMjNC+au
pNv09R4RGOzC2ESHGHoU/hpwe2hTOr/rf2qXFwFOjk+NWhIE3WwnpqawMqhEpCwejauOTOEo6Lvs
kn3husphZCtxOyKpuxUNQoNUGnmfYm/Nn7zDSdgLN5afr2X4fytDweEf+4R501aqWS9diLZf9XgR
qwCxpAP1L9g911030A8FN8axLULm6iGT4qMLo2cxDMD3EwyguUyTCn26rbZledh4wV7UQBU6+yDt
bQx8piVbdsPtQfnLPKv2FF7EDqvqZHHMYyZOFvwESTrVxOy+Ng48NcE6r4518neoNA1rlIgBeSjF
QaOVM1xSQAkp7NbjRNy1DlIhVsHv8gYPeyW25+ajBtQWrjIswXAItsGf22jdSMM9rGslGW3otlEd
CbX7BxjySsemOlnIpUiMpbQxgudVWzp3jLaPuX5fAET3GPdjqbkZsBiM+wg+J+28iTKUnPTSNlSw
34cwFn29+c3BLsmV/jbkbK8i6F0ZGSBEpoX2j+3ew4+aD5PIH3jD57C3T9d1pWsdTgunuI6V9SSg
gZ2NjxcSGpFP570MxuDCDHS5NngOIJae8i+IQp0YtnRaA9pEB0dWQzr0BDFbPcPzftkjLWlkK1yN
SsgHh3N2/Z14hmXaQYD024ctGEYYOFCB3ACbvrGNV9Pmb4XY39qhwirail5X6FDG9/vaxkeaYQCm
BFkIhQXhS3CwSoDMmrHtVR3RDQXSE4bZI9Rt7q8SEqcDkOwSIZu6mPGD6mltf1Hxu+hk9kgWVwt/
jq+werzaCEEOER79Ih9jioOZj0ETUdeWwLrnPq1PHri1D0e3A9CA3ifeFLqDkIzTqn1Aj7ARb0zS
6z4SkIRAuzp5fNsWa0eNFPlg7JeZtK0Uu0TxaarZ2jPlj8hVxoC16EWKlLTDq5fT+r1srFuDCE/k
4AqDx775C7mDZwJvQ3S0/zs4439okzV55jw0tg0W+qP/F/DWFw4pxgPTpHRp+M6tmah1yIBzNQac
MRkG2ZGDZc9nO0jIVZbnE0NOMioQQ97SvzaJPAiykSi8QOpkrnlspWzZpfONW2bakQrSwQGUK6mH
37P8pcCfRAVh8lZtbA2w62oGCAUuJymaUvDZpoBV/QAu3s99bWmFVrpU1722j+yKgrw6M0+4Civs
1m2qxcploOHrxI4tMm4LLY4qj3vYoiUARepXdDbOKn0b2IEW8EIgFeVkS2F5S428SxkaSjN60nHH
Vvm1ffD+qizPxcgsINYMiWxkjeblEZmR29WEEUYhmdjAkej733VOGbJQWRMp5Q8Qxj4ow8eSM5KQ
LSZlng3B1T2c3WL7xd5Ky5Wu7kUA+Elt2V6fN65V/4Tmm4QGYbv2LeYPsMbpvCqz5HdMrJ/0Ol9Y
9TSyeih4taLegWIlib7API32w6QGLIbKnx9TCcIWBzyOCx32/j5nZ/aTBiLI1T6ZO1SfRJgHnev2
IBdd22Jtmzkgurx8MmUrMzGYqr7u2g5O8x5xWLjHe+n/U/tQGW4xadIKBwSh7wcyxBCtobMKGTFU
2CmG29zERzg00a2AaQ8yMbFgKhKz25FxOb/L9Jsp5YH6Nw9gKa5ofaemDietOqjigJbvkNlM2ikz
bYfUm2PyJnDRUCci9DK9wVutHIAsuQDxkd068vZh6iEF7JVUdVnrAm0x7NyWj6FmQkvsrOKJ/Ui0
o0uuI3uVpMpfcj2Zazr++aOoAPdgmlU6johwlupaU+OPxhhgqfTKC0iVjmLMR0tkEaWwphuxaC19
TUJ5p9gQzNJ+gsPpHFFKTSEEY5+DwngjasoG4Lxbdv5SuD1VrHoKul9UznBVDgs6hfJgUhCLPz8G
1Iyxrtf1zz0F8joyJEa3/C0BmEPPMmnG25+C8sml8uaC1wdaoJMt7s6Fp+7TF/FwTCZCQr1/kIvG
Zi5mj3HzDWdpWnJMlEFM3HacGRAb9edUjSxxsU68KynWa7rE738LSHYN6KpGyT9APns5qgCYFoT3
9ftfIMA62ToSrqaC1wDGMNmEb+dT3Pd3UDaq66FW7wGnOcVVkmLhCAfb7eG01aBn02iZuoE0p9PD
3NQ0AJgtTTJgQtz2+w/F1ymiiuHhzcuTZkBX3DLm6x90/4m6CTaQAQhOuQiKco5MNvqKDC+f++oG
kYKuAUhAQWSCAmImc6UtTLQFJmm+/tMfFXsUkTNjK7kIw1e6C1a7g5mNv4ntFgpbwZoPr4Ybsdpz
2uRDwVC6Bl3x3e6dxvZmsIWqJQSXnLMx8ImZRH4jhHVHQbZ7a67jTiiu17JjFyCbM1PQs6IShz5G
65ql9UICGkT/FR30YmjDJcyOlBEoHMlX2/iYFYJKSn3EJBqtv4PdaD/ch7EcKqHx/F0ON8p4gW6O
5e8loRougEQJLJ6MT2Z1Ml2BW3zwHcH/HHAw3frKnHnyPAMUB9QJo6iZjN7Gn3rguzL4Z/v42POh
b8GsysP0pLtsnF8FKvGaqi9bIfwoGIwu9PYHLfWUBKY3D872TeKbF1NNc3LDJHANxk2kRb6w30zh
zHXBi/5t7z5MqPyZUy0AW2a/zyyGCzohNhzKfM9c9rEC3PRYFvV0EUvgb7a85cWpkFKSynaDmlHO
kEEQ1n+D0dvCtvsinDNCd+PgVZSCLsDWAtsVUNliuZuOQfuOnqAMlJvDq/l4sT2YXcWyPViu20CP
wTMoaU89sySPIf+a8iJCyswP6IyT9iuOdzfRIyuN2VOWLfUO7IJsql+Bv5jCnKuBJCzMJYZu8nQE
70QTPy7zNSxtJwtzzlPdOHxftbJDvxxQpBvaxTFQqHnA8F55PFlcEIlua+kWIbWv+G+ovzKewTgA
cY6/YljapDtR8+tBD/MVRof/qQZYrdcX1vNrieK4gurMpiARFYDNUunu24hOSh+/QMNHImLrwiEB
+BbP+VVgIgYY2GrKl1P4bbZ/dk87CTudebMbAiuUwvrenAojST+VQhGH+9FrksRelqhom8U6hS30
cyj5t4ZzfViSFRi8/S9IzDeqmXnmx1gkzdPArdG7tH6nBAkQ7sQoAfIxvMvSwycTp0WdpECMBBrb
CXUhuC0AQaS0yDPgDmlD7bbBZM4oyy4OAxARtlJ7X9/T1KbdXVWWx5R2ZM/TL5OCC4cw926S9OQs
RT0HEY///FM9s1ZK08PeyDBvisxXS4JBg3pYCyPUPV7+bZ71m1XX5F7DAHna8fQmAa50Hc4zFgla
axFEO5HMh4LTNAxkVuNsXGAvBz3UQekSXBt85MV72Oj82CtA9Isuo4EASB/Fup+RIMuPWSjXykBU
WfmnQrhgKtZ948rfmWFfUYu6bGdZnqP0feqGqbRa04/UKNz7whuzzcnOlJpATOjAjwipV3u0ooFe
0+PbE5pMvVUcS4mDdjOfkuXHDlSvaQ5dh7fi/sY0OO3lDaRbWOtny7rQHhWrvCryvB/vOsSfRMr0
+T47Y+fo2mGgpaIBgJwUBGLXcOM0ot97IeJHfavN0cpK4XpzuoqBqMNwc0175R0k8wD80i+EO/is
5OrTCJZRoVbex/13RLGoi/liTbC5av/cnNXM1veXwfyoYLYpM9VJlwNQs+j/VdrW6eLy/DAMedG6
VTfH/drptdla2r42JFzIrrwNdHjlfASz8InT9tdZFbhw6dHEk318Q56ZBRMsUGApbYDtlt57PYSw
pdCjjb2EqN0gUqbUo1nxFeZ+loz8/J6FLAp7lWHxZt+MgSJBqq6UJ2reFX8dWQsgZiYhu71181/i
kfrlcgfu5f4XSArBn+BchmMmdmHfwY5xYbafgaUg+ws/8vl8M7/fHEXkjsU/DU5ggZNemG5to5yf
+A8y6ul5Hx6vYwATtjx3yZF3cPkNUtSh+0IBUQaq8M0x9L+EC8oum7DBcYfCHp/yBEIY0FEfjPIo
T3xooTQXzMxIK4GRQWOietboU5tZKttAA1Ag1wpdXsMy3q/XgPFYLxV2e98H2cRuRG9Mndib4g++
xhY82eAfex4tTUkwr3kuTXB7NEU7ipRXWxRGNB3bUg8f1JiapNuWuwlSfDb9OW+ymQQlYI4XWHyg
EgJY3hNhRNh54X/25zZKhUUn6ZtB0Bb1S9MzK3+u8sfiD+6cdSRZKScOurWCcXqPSmtTJl8GRuXZ
+OHlNMiljIjx3XhNkJyL2HyIqrknBcMt9Y4+CQTKq8L2+GaemwQazqu2VgewMugvezUMAtAtYAk2
M2Ll47hp+z0yAMJnYmFCb+z3hLkSB+/wAK0rM2Lkl6z7Ep6P6YsKjMgvLl28Y7tJfVRurCOzNjs7
rnQiOKsuavwWKLcw1Mrek0GHrfucHGMHREzWQYq3q5qcPQYgoixXebCt7DRKhQiSJvjMSbr8Rf0d
6urtohIFwwTMOhKmIpUID1oE3jS/CH7SZkcjoL8D9hbkoYURBYJ5yzcgwfAPvrcKS3iOazHGLdDl
XWtIGigMKyOX+k5Kf6yHALuJpHVLBd1/OZw75X2sOCx5crFiSfhchNKiV6/+W0iWOy4tebp1kJiE
YcZBO74GWmL67zSgSTzHe/siBc4OZPQ2JUN+zuWJYzKqxoD41olMBd99vZop/hyVhJ/2kF1ilQOX
w+5KSfAcu4bYbeIlafkQy1Ji1SzC11b/JmA03l29BVsu3VhcQnpJBZVqOEa5dKgLvjBtENhFOI9F
Q7FaSClVBXh/O9l/5pEU86mL7noPwbYiwh7sIEJqfTfO6jegA7goJs7kQNjOh+JtSBQ2D3UWXjRN
g1gJxYDVtyzOSv7rY4wEEkynhNa6FeDca7bQ9nW96zaZQXbseCJNGSBjG1ZIWqACNP1bhsvt7l7E
Awi1meAGTiPHW/Hw6KLb2wZGbeZlcjdQHIWgmSkYq47Fyi9F6cF655obOcu01ds7I3XMguN2LCIL
bJi22M3Wi084Azef0BOMNGcR/X3BYCkTlZkvQ6OwQ3EI1ANm3mW1Y2op6JfHO2nquZ7OdaaOfQBE
9gNgJrdRB9Fslt+JdrD2G8enhjK0KJKA+xlP/MQvjYOzuh2rsXx1W0d79WbDcuQjYyvip+ysaJep
IYFhLw6NLiTBt2F2Y4CWcCl/qNMo6Ei+PV/g6lHJAQLdZrHFz1IIwW/rBBpStp+ZVTIzvX2G2SwM
kY2V48m3EcQJwIXi+IuPPv5AlVGzY93J+O8uuOR46iqxz2Dh0o3iqwX1iW3SA4foyGUtscTIQM25
WvU50V5oCQo4X1XAGwXjSEe9fauCa5oVffgs+EfzxDGu+ydyLUjtZaI27J7B800mg542FL5s3Jz0
BEbtHi92JJBYBLvShCbJPIGdMcf0H/kgliQnx3gNp2qbNCVT5vuIx1NEkeqWYqK+kJNJ9j+kqK6M
qEAnUx0iH54IXKRKF+u4sVIUm9THcGBYUmL5iwTbBv5bL0R0imYc52I+tyBJseokbyVTozt1mdPf
SnYYqAbX3DC2bVEXBzJp//KuYT0TMnpoPCuvsAR6NlLzjWmRML71SNXAP62CQPUSkyramXJ7KCZC
Pr2tqPvFjXfUy+kwWnH9OzvbhvFqVSD2rZBFkqlsju3QAdioLGGsdq4TM/qw3lui1uZ81lTMQShl
Dn3oqE5spmMdeOS/0J8l90c3o06muzoDe1iVXp4XWV9SOHtfkvMGwViPcGFXvbOS+84WWITMqUzf
dgKeRftmghIOQXPISjNPZsJXMR9I6RknImMuEQAv8/IOqWp0oO9vzIt9/HNtCTYwHlFBzWwcpXx6
pryPSlPcW8CssyYHg5kh1PWQan8BnkHp3e+D0gQYQVYtLpu3bjwt067WXwbo/BT4YF8hkCqYp7wv
FP3Ibi6cC7x6yM//FjorE8ZW0dzfMJ0Z/7NmgWp+JDaGCaPqAntF4IE4JTJSlMh3jSfFAWPHE1Nu
Odunhkp/UDF6cRbIzur+XdjYDpC+/UULKRhEcx4M8JfzrWUE3WeZSlSyDClEs+69i/9zpJXQp5UO
68bWEbvkuVSSGXIBx6LQV/AzWzWrTE3ajgpubgz+R1z6yw8MQoX5StJ/g//1jOPIpGWO19bGTfQj
m+6reF4twCRiI3F4veNfXQFkfvZH/lYdqeFefRAzhB8VUW5ko3AEtTDAij02j5uAsTA44ypQ3+jD
35gAcASc7tN0PvbQI/n+NHOZVl2lrOw27p4wCsQ8bl/51SPXerMEB71oObAcD8RCB3/OwwcDh965
Uz7T3bPpEq5nH9rkwAiKQIsmKU/Md/mX5KM9IUC7t3MS0gZ6Y+zSHR0BMlSADzxQqJsT+QNq2B8a
TT3+tvzb6A/kC5Tt5Tp3OxBRkedn5E7op3qc72HWNf4ZveBaJ3iMrJHQ4VR86PQAgZEusOV1aLfT
Q9mUSsUDlyTAcOV5TAI6HYBMxic0Lo1E4knlccEhyCaHkVFzzHim3ixLHE6aECeVyazB3DEgoi9r
y3VbFTEkOPDyupgVjwzP1xe97lsnRQTkSFQCyB9CeZNYq1vQshungJlo60KwnvP+su8kFrRco/RL
u44KH9DBLyzPyqvo/MgNGfhrcndftPZOQZKpjSBzufzneBE0BOCBmLWR6PhoQjsggwtGgsl471xR
VatiPh3Qbk/+sLopZXGXSU/dCa07YA+H1gZ3iME/4qpprbGr7uLFUlbgnjHeMoRdHLH7dW0Aypx5
ZfRX9FWpvFkFrGnNE9VQ0UAFjFiLrvhjuYBFjKKq6xAIc4ZgY3DI8ZMLjoIEw7urtALW65IiiM0R
lFC/7ZBOtFJILAod0FFAGW5n/YJSpt3KWutAa6tYN+Unk5AgWsUFp3UxWaRyZn3uscggL3HIHmrW
BKGwi/qg0CJsUG1jR704M+7W8rOl1AWilWp7ea8ERwgG6Ehnpt11Y3FS0ImfLhyjo8hQbpbmJpf9
1OCd0k3iYyyEe+luGuBQ6qP3+q5coi3Gu7CJM1R/xbCYsjTnbeXExHhYtOXvlEzUIo1RwhciUbDb
R8q+VgYIvRkOeiQo8ydsMs38GxB/KeR2iUgqC5p4KGjiy93pIQbo5IutDtwlMgM0RmGBSTmdCf2C
F2a1914WBNr0GbllTCZM7YK29zosgV+KF0+smAMVcZBp3Vkp/YQsA1+OAKJaQmNMjipoc9fyuR+0
wtrr5FRPRPZ+uG6RV48CVaHTnWpaViVqsOpwmoLkZIEfh5dr3HIrEg4yr2XQkBRAs6EHdXci4OUZ
Oydl77Y+h6QGC+NZnFd7FKyJiIqV8pVHvSOJoKv3CV/yzyxYDf7236pZMDS/FJB1fLwhiDT3vRrd
eCuJZX0VhPnXv7kGvO02nrgE1+W1DDUmMRBXS9Da3TPa/08lt1AmZ1vEm9L2NUojwiBuzQsQYyp2
u76MqZ9zRbPRaBtb8EUqULsQp31AyXlhYoYhrjTsNXPqI3UnsM5vBsqtWMRDvPvpsePqDCJmlLmW
GxRtq4ZW1v+D/Zv5HZXAiIRXWpENKKr2vYthA0zM1CyBqtxhzDFTQKT1mW8CjZdj4CGI8IL2i7p+
nvhHkVuYOHkXmsOkFIE9e3GOQUm4PgwyLdZKl4BjqFImv8/DbWeDYi9GCEwX1iqCsXyqkYi5iy2D
48phGKE6WJQWWxHZhDBnF+Ai/gIeLTzYtXSp4v/ERob+JXFomjY/IkdMg5PmxHXz+HD4zlsZBOYe
3CYHFN6FWHcfFcmbY3vC/I5gYaNvldg1WcAyFCJgjGerMVxVkunRi2DvlsLMQjD3Sb7ctLzE3PEL
zzSm8Dg4XmQMAYnCC9hI2lARUbXXU/gSZS8XmtgeSVgfOeHjZMNYusbXUKdyXvJsCgCh6Qoyyy2c
G0HOLEMbquV4ySZ/DTuUIBh+YXb6zim/N8i4eyrYPTujXX5fextNB9D8NFV99hiSN4pVZx0vmTnN
AQtCHRDE7jCP4BSFBSgBXFU7chvSBF4gzRUWGxu34hduRjkWw6PXQmeqyutcuMGBrXm7EllPaI3a
4u1HXXjdIFYxrikmFbJauhhtqkwBDOwQho4EZBfNYCEdlGE93YOHPZQNGembARtb+5uPDuzvm7nG
aBUjb9xPty77MIFztx1hPMir82bMDd5hY9EgOC4y1hJ81deMapXmrQmzWomNseNX28MmD+aT4hvi
KW+0vXCmMynv8FSNX1f6e9vBIaVMmaCSl1VB03F4H+BopLrBgqx34l3H4potJI+YP1ao+4sPmyO7
mCiibGDg1QcLG1nTbe2NQ3IVjKLJAo6CgKIhH6qcNbUqhcbPBlUYn25NELx2gyQQS7No26OAYla8
NnBlQ9VSFPkIEDGL2Dd6n+7KPQDpJzHEyqpzUsWwQjiRW0mLIw+N9a3FKlhqLnSfB5TWCPw1BbQx
SlJxa/q5O9DPgUdGVMgX9mQd0i3KJneXSzhAizUxAdCk62uHlHBs+uYXIVc0c9ozx0wKFMzp843O
rkeu9zhImxDHtVVEVFyBYxQYnt9AeFZfPpAUDy5tLV6sCYobViByNOZMWrYwXy7xIeiaR16MQUaB
4lq++WhdymFqPPR1lOHc5ZpHGICiCVGPZQgR79HFdvoyqj99FUV4Kaav8SflHOX7cfXWzd6BQEG/
nyhsqbY2ce2ltaHlTNYdAMgRTLWdHsqpVJ3g7gVlp9qkjBg1LDGgAzRqqZbD68cLCM2tpvztdphD
CHB7cm/01hwufHyJejGaw1XYhqQUqTlQ4RfLhRCqwdAjCbqPEVO1Wl6DK5YDllXaUFIUGfXB8FZC
5vM6fgrRLFuIEtnEzmskgdSPw0XbHIVzLA3KsGXkXQKW8h7lROMwBXYvy2uQvX2NyJR+DJdXG9vX
cJfPjOacJmfGKjFZs3j1WdGjPnzcgABx7gEzPrU3Y0KIAzzf5flaWcqIuEphzbCDcBbvp5OGs9Iu
pFdMUqK8FZwqkWx3R3TRit7mTh3ehur93aSS05w7aRv8TXSVhLl9ccJzHQhoErXPSkCKICbBLvP7
GIvBMr6SbVvIwWeOtuU9S1tDJOFF0K/ssXnXj6xiJnIfl5vAKa3mFIcx/7dqvi7FIIfXmbYvd4CF
626+aL7b7IcsjpvgXWPzEQTriRl702gDBqUkDCX0nw8RpUKJQU1kmeY91O3gov2t02DmqFn1BgqK
e9uVWbwtAn6Uja1zjaLXFE/ksFRra8fbAJf3T/uCtAqgct7sqAzT1NS2h0iA7YAG9pQdol2fGmcx
LFpmCVJxZXYGivDVS4bbPGI7QK2PTuRE7NhvUB9fubUglgiPX1uXTfNhv3B4oQVG4YdBgRDWBzaG
juAN0+hxATh5iEfZR9Ed2Gb4i6/Jvk9aMiIQDPtd528tZ1w/Wk4kHh58Ghk/UWnyVHky4npE9skd
Ow+gKWA8alYN+wma5CBIXoEG+ZaG+136scWeS5AzGq+h+DKaJ23CdUhNEkW9fiWDzS22NHTh2YIc
khcnVvw1u5XNdmS6d8Etb8Bc8eG4RPXpd6S9Vh/ivIW925UYc2i/jCovkC4pg/ljJNawld73Cp1k
noKZP7lXmTR46psoIP7b8byLKJCk/i4xCsWi5tSmGnsdKAyr5nG5IhDrbvYUbsgRXJSiqYfFLJhR
wPPGhOhQYGbAxeSwhOBXWfgaHD8iWA3CFh2mrt0OpxPFPoyf1SaObjhQXmtWlI15FDqqhEhr3OzK
VrTtedCvU9TVA1cfxbmfcfupBF4p1TrRII3BNRnBeCQ7TjVgTF4in4tWWBK3xGdTm6YU4zXUDD6D
ALWeTjvXXZoOxDubF9vvX0olVpoZhCNhq0ztcb8+8LaxOZsuVwj7BiStj8LlSz1B5yGBLCCDTb3B
rXA1xG3Elw5MFAMt56WRz27tC9QW3achOfqeruOt8VmekETMqAmWkiyWiY1DuflIDj0Zq+62e4Ox
M4oPrChkDVh8TfTdFRDL/EP4QFX4m+EOXP/4uq1hAhZmIhC7k9bWvOcO7SuRzyKcdECi98qYM1X4
KcT1c1kIgO7RPRaWKjFFWHANjWuNyUORp1rWu7gVGfT4upzwR0t6kp0ytE3+7Mbvq0AHuWQu8UvT
0IorkazBCt+d3kVlBId4YqFc2H7MDyy+riEI0XM1KTLLM1cyD/Zok/hXF6bzXgi+4WGmrhmEzO5H
2ITY6UnvukK8+eHM/mHHGxJ9g9rvrkiXMHNawVetCy9VG9KA4bfVmMnC+EonA4V6oxtOuen4v+mB
au4LAbGxResovf+F4fO1R4OPATCKmh2lixdE6aNObrx+Aun2UkUfPwwQ9XDl4iDPT3MwknEqpwJC
Q8CaDkDkaPe/mKFDPVOCqj5lRO8OkI5vAXLdEYGwzrYS9FXuRAtT14zTE6av+w/57/ArfF9Dcy+c
qywecds/3tTkYeC49tZWW6UPL7+k67LDmU4Yb7NL7FyTyUJcPh1PRsrVUh+P7EXJNilh1t2RcxAz
XYCgPqXRqHLMoGtSWaKxB0Rxj5DliQXFYKRIhZ2iNyx184HikGCWt/K8lR8ctyzR8rYO5lvr7Db0
8ZK5nZ9S2nidpHHruLMV7Bt07OB6oNNcZROBNpSxtxgEPzsZtaodBaFd/goWRVsIp5WEzZ2C+zzq
ZeKnweKzmxAAfHGdhV7/AxZpXpsWy9sjAzcGAEKhpbK9tKpZbITXSu+qf+S0X8lAs6omoBpmIQL1
BY7xuygsl/K6H9lC1JQoFO5LHGendd1gQJi8kZXrQBAWL+P1zYems0Dk2VG6zq9Qq2aZo+R3Sf34
9sj8+dW08R64nPLIXw/EnFiFRK2IaZjKks+Vt9uehKbahH/x6XegC6Z75aRNrD9wK7yhVo0tE0uv
Dka4gLrVxXtgrY7fs6AR2fAm7dPzOn948Pln1KfsaGJvOAQ32H6aG7StuZv+jpNZclVG0cVl6nZI
XcDbTsFiJwgfkIsK7Kj7J/Q/ZwiC0sDS7LJolIajrbMsHnx1sk4AsB25oe5oTU7BZb4vY0ZcgA83
NoZr/dqUBUQ0JHOBYhhuWxGtEjY3CKl8Fi1RjCT0zK/IyOiEhMDBqpeyXEQr+77UHtg+KX/61Ycm
fcfZ85CjJHQQnAlhGvf8IJEssRJiPF6qwCSZGUbKBfcEwjQgE34tZXauQ/iSOSatP5qOzHxVkUDk
LlC+kNzM+ijvI0gcrUqAIGcgu7OPOXCCuP4eeXPs/3i8b2QmNSiwMlyI0IzVHh+OSeXOSqGxt0bF
wyrtPMtrl3chqXEwfQ0AI3+kgSA7Q9a08gxkhjy7eD9b6P+Wur8ExCgXkgGNZpaJthtJsanUpfmC
8vqdZeD91SKpb7fr9zuhA/fZXwXkZvJfJEntveUsYICigweKCU/zNc4BWaXQE3zWwtiOhcK+31RB
VSEb9fqOywRo7obsxrhklmWX1JUwDpEdYyYJjr5De/iDZaJGgTt4IZhI26dcx//G2NTqfXoN1GO9
JcmFewd2IGq20BvJP3n+09oVxfivfrQB0pgj9YrphAwdF61nm8OdMt9go0vDLQft9dmGTn3GP7dp
UzoQKJNXZW0sRs83J8f6IBBEqU5Oz/8wlZUof81cd4TqHcOhyzvRM+X89dLfKC0UtPkowa269hxT
COStTHCK+Hu8xO+LYRZ5Ps8FAblAprcyb6T4aOPEEPDpOFUrO33xy2dl2PizijT8fSxY5cs396ee
qI+JlsZogQtAsfwzk6aHnbRh54HEFFWsCw/T1YiPi0EDoxMzyj6u3MvgiG0+LQLY8HG68QBESbys
r/qQq5CsoE+g07Oczcb2G1XXh7996nM6+LsA0nEYOi21CrPzs1AZV80J5XIHV7ROfuP4yhq1hG6t
yotbWDCvI1HbiwkZRl+XosTvtxyBB+uFVZGPBocQ62a53ZuKl4Gy3mG3ufr4pFJmVilK2tgoifNh
tH4CTgkcOKCRzeukYiRPI6ykect8sdSzvqHl9mtK2pmKrbqwFqlmC63gInLQI6gdyAYnq3/Jk0iD
qqQQErnq0NQFXwek1uauuA/SMZ1yKCn7AJLl07JJhqC3IPyHKn0fEt8ziLrF3pG60AbdMuwQTn+b
64yFg80WVZm9TyMerXau+h9sbdRg4VP253S0VgjLrmUttmAR6zaBVNkPfCNezk7tOpL7FRtdE+6k
TAgqw76ik7T9OjYehmSJveX8x6LhjgljihKh8SCV7P+6+ekRPGW9gg6nYUpBmF/1PEyvQf2x9Y3X
ybxMCFwFBgsMVpfTGWvrm8t7kelh1DJ6Bulr7mFSNBl9o2DfyTYDAeBFt4h8lGlGSPrE8mm8TKVF
aOZmP/hXlBPnw7lJ1ip6Vs1XO7tyhAqNLhhCjchOw1VDiS7DYRqApEd5qdJ9uC4Z9oavMqNHQB5v
Nk316mmQoQu3xnrMtfMrzJj/9tACSIpC24nENr0IA7L5+6+oHztkGzWUJDijDxtSluXJzbB+sJVI
At7XOJr+I1eyKILvAo0+nzMx8zvBiaDk3zjy/xg6GWz9gag+WtHJieGdCij0/4NGYsBbW1WihuNR
IdLBDSsDhbOMudNmHr68PybQc/cQ8wWey4BFmDKb2jBDHJuORKLTbCDEH2YdUPa/nHsODSLoj0IT
OoueDQgai6LXXbHKSgs0Jh/r4sTleJHAsgyLiYpj73qXHw6Rk0lAZ0+X0QTJBB120Ctmz8ayfYSm
lDsE+Pg6SDe4XaGLA5E7B7EzcWVNOs6cvfcM7j2KUyNXFanESFeWf0i7S4SzlbLs24RJtjbgI280
8AE7I83/Cs+lkrwwULX2KhNxEezPJ9KkLt2/2yDVUInrgfduDeF9ba0Slmsd5yTalddpyJT7KmyB
tLFxSDVTZtJfN4UvQsEHVpPmKupPg1ueTQvTIPVR+AzPxdbFTIBxbxlVXOyiE/f2zhv6O4yWW7bj
5zL4o8R8/DgzuedRpK2eYG3rHJ39eZSpjGuY687Z+ojbRe2x3CoXiGkqX6y+pbRZ4vM/e1SzngIL
5SASdr9a49ppe4yd2DV5PUsrvDncOY61JjnVAuVNA7Gd2EEYGofDufMPOpZTGqbXZ5Zik/WTxLXx
ALoX7Q15Eudmg2mxCFLS7viS69aSj6OVYwVv4XRLrKwn0ffQ9NGZyHqgoIja6Qs8glByezBgsPRG
ndrqsc9usxNr6bOPDwZ6RmKutFEWCBBrlcJAv1DeQ/uwgMg9XBrXedTQKXT5IGDViPCo9cj2ekp9
5xOESMt8qFsCw/OXBtdceFoGhnkyk6hTufYGbzAxATj6ZzyLzZibHmbjc2vfHwnWIBDwBHXyZjHC
AUktzIhF3/vu/ko4paZIjH8dZg6uWlt4NRa8SgjnIqzOYMvZ/PwwTMvYKLlOYoiWOFu3uVce0e6Q
5eyjbSaUJyFlYWL85Du6wMPKvwRAryta8I1Jx05mqk+vtUtuETXamvdaXyXHS8ECFjLFs42Cr3jk
nX33oAFHDnK4/V2gyHqHyN2DoRe3LOJNHACm3ZqYSpHB/oGKfWO+SPf4eZPOfFIJhQddwQyenmHE
dvT0VvQPCmVvqSgVXU6isvjhgGB+hloVZs85JO16ZAhmh3I3ar44EHBFPzHEQUPG7Zrw7wfUT2VR
KDd7C3+sl31SxiFdhivGDwOzsK6nI7FES1iPI7GQ5+AXz6/syfaDadfa6dk66Z3xqlfH5ZxeLemk
0FUDW/MfXQHeXqCMe9zDKdSJdbqcThyrQJDSCbDXEtAy+dCyp3cnKS6vdvb/gyDr6s2dkXlk5kDr
z0ytB5+PKGnc4i6kAfSHVtmqrAZGE/df+JE47ASpU9pShxChnJjgBFPyRyjenidqFgzybomss4vj
7VhWXtViUjw3h64nLGQ1Gli1Sp+MOBlytfhcmOqSI4CwTV9/mLf2cOO6LYUuFsOEbMW0ZMt6/qfW
yWRPIrI4TMFLg48mNonQXDvApeS/fn6k39lMzzXSuwX5GTig4+LJsKtwIDKoeogUaAuaErd+zGzR
AXGPg133cvzZ0sgGc8gLYYCpRvPcYie7duie8YoFAtJbJ868Dvwn5k/0Dpib19Bb+SN4FPmIKenX
LJggZKz9mPlk7AJYVLZdVkE1GlRbCdKLh5SU42h6Ke6OSb15OGeDT0fB5rmw5NrROol0QIEAKJnB
ZErhIXQFxHS3y3omEr5fVzBpc4FDQ4sPCLIcP3iG0n1+PH5GmlbKKsz0j/Cac/7g9f2SPWz8w8dJ
vOozrs3blrpUEH/eFSpYHTIGYdUhhcnVKPXL7W8tk+pzr30ccEH0vsxIHKFb8Nb35AT1zFvTcWHx
1tjVGr3mj07rzabklbOG55WJCiOmBcUnmWJuaA6rTFIBDN7NQrc8RYHPVHCsL1VZc8Rny3fRR21P
vpFLP38J1kNdaznYNFboeDjWMYBfHWlWIjKDjhYrHCP67ryfripU3STkAgyHrnlPFPuOaPCA7AFK
xPwXewHyaCiybIye/WnREvtRPfIqTt74BK92ugOfcJW/rd6n/snfc9SwyZdGajuwbN3GAMEIWPCM
kwvI0YLewh5hhPvYdVO+YrKTMD2GgU9ab5+JxQcqykwdj/wDc2GfAjbrm3nbpB0ldaNEVrh27c+Q
d122UFadxFFhZfkrukTcLJLcnZrJMQTFJuerZqk6X2lsWGnzEdawbnR2wlaRvM7/kMKGAe6cOqlj
hhFpdv38KFInvtvYgOZ/1x1GjiYeTKDakSyHlZiM79d6s+duBwTuF2GTsNoWkFoLKqwJEpGxL72x
hx/reg4cywNKrJCQlb5e4S4EwEHpVgMWma15kxzua76FHNt+OM9/Ns9PN3Pr7rAGPViaRr6X2Cg/
Jj0WEr3U42HWBGjKqRc62buQBFazZ4Lt3vgiquCz7d7VjGvgKUASUeNcJjMKJNdy+j5fo2LPrKr/
GCxksOj1ozWSxxk7kVOYxF4Zkd+A++abiIB4H6IvMMxDsn6ZOFYFI9tQwHCn8LVFboyE7pSrOfFm
/kbSljJSKS1dMjPgWIH+4Jqv128qiTEfMtAqm2KfvEtk4hQv43zsBPg71j6kx2QD9qUjsOvCDIU2
WNPoFgfzUbNBz1/cuQ0lx5N4w1Bu0dpUwxmFuhooLymfzIWuu/paJHHRsHR0egNN/Niv5n+qKiP3
jRbh6mo7JhRL1pvEks/e5fFvS1HrTeGftWasKBbNSAGpNK9Ku1fqVwRWdPUEC49Texm8Q5DuNEWx
090XMKvRqF+cwKtBRY7xaAg1Vf0EzcCKPrvufmmeJVLpXdFD1Pt8xr8S57GgQW239OnyT15JtbHo
RwiuRIcxXxsnNtQ+/nG/9Y4PSoI/8H96rvQqBIvZPmms71/YvRps7XO3p8seHQKd6fuAI6Oawsmo
G/zcXviUrHjVxesCCZjgZlDJP59Dm2XNdfi1YNmYPhUDChg6Gf5ft7rc98IsVBP06MTTugHHE+Ky
UM9PlzBeDcwy5m1dU6dUHd3MovGX+U5mf/7sn9nd7RQK0CmDt9soP6BueH88IHAdRI92CcJZDEIh
hfJxH/se3wM6wOAiX/xBls/56V8N6fCl9hnSPdi70PBDrWIOWeL8Y7thy8OO8fPSrmgEInO02wBy
xGetIf6KPfDIKL2Fzf8gvyMMUYaiK5QFXRxx1POKKKTDeyRffpCSVDNqtOuwmNK7Lb8Egqmikdn/
CrhBz3LWWwcwCULOGJD/YsJnzEmgyj+Hzu4NMti+q8L+SuVHTpdLq0XbvAcE/v9VG+4crzLd8smY
WdNXLhcmWfIwMspuEncqKhddwb5CxRM4/4bBVnsZaCMMmgedgiRwmB/nALWGCCi8q/J117m7N1ln
oVelH6B33vbqGbiAK7f/2ihbVUZ/cHBBLD8cnUhj827Fk8URAw2XLZ2JL9B3x8UzLJk8UFY04mh+
ItAl1nhtey6II2QBkbp78VPXHT/bsq4Znj8AIXXWJ2pubkG/RnWJwzU4nSM7gUVbRnLF0v5o0DVI
mT8qcxqSm+rcLRFd9dBffxRPY1SVngCc0SP8CoNwF2ZDuCd3PkfoYL5ipc6PeZEniDQQoBmTErvM
9S2ZFoqEJehkHf1GL3cRgbstiAg5+Fa3tTsyjcXCY31hEQzkMxwLZSt0kepgCmEXP2yo0+qtkocv
KnS5TUvgKtDLBanA/44hiNM1z5lCSrU32w4BV6hPSJQN4J+w1flSNyLeErtkoWbhAEknPdtCXFyg
4K4l4oupeNNTLpU4V+4ukdXafI+lLUzt/m5OBdPI/3cr3tJfqB6DiCOH8fKTrrGymAzDayyLhERr
8Zaa+V0bGUpll3rm+EmJ8BhBie/Rlijatf0O50becpdJuqZwyuJuLvCONimu39zaWPgTDaWFaBm3
fsmG7x4yZ731/15S2V+819bn+U3CZBML0Yxx8hEp567jShhMalK7+0TdD98FLWDxml0jYA9iyWJZ
2A84GGuxpu4aKO6D1EXfbfip+xwkFqVyX7RW2wdbt2+IkHJLlGtpMQmY3GJjNWG9NuigfnbiuRWY
d3V40vKcZ5ULmKhKpI+h08qre+NiWjdkd8CDLh8gXaj/1trsKe1Bl7k6oNFqAijjQwGYQp8kUXch
BOC7xDaU9Q6iLb0gG/V9RzEyrvg9Ehslk2RpyAlRLMVYMq5IEr5FYAwNAXF2TWRD3J+yJhUQoHnC
2OVfCkJwUQxGp/dcxJThC1GFELxMpN0sBrdD6M1tAC8WcU6vTq1SX/W+aKcMl6q9GlAEow7JeSxB
94ibNjlqTw4XbpHj/rPlnrhOHW/W1I5rPv3OQIDVBgiRa7WO51tTuSm+zHugVERqKyJA7R3GrHUj
aRkwxl3lrZsa7F0Yiw8j6o7lIpRWd9rUO4EguFpwgHPqOkjZ2Z7MzqsIIMcNLAaqsxxJGhum/KO6
WkS7PBeb92zYvPWOUmoBXbecEMxGYEkzmqW+aSuicDqX/3nH7qzDbTOW0U1NpXe7W3L/RvriCxLw
DCinWzIbhE9dFdA3hNhyveIDzyiODzaJarS+KKjmdIPxI4+7GsGcPIiYUnVbHb+GABuifyb5JoWr
hCV0RUjwoILw3ovkar1rSeiEfO+rCeuSygq2uiwCIEIhcu0BFm48xve9XpQ8i81yNwM8gM81qqXF
/a/43MTy1gTk7gXZiAg8cP3JCPC69RvZGPLd0PVI3jWQAAz89SAvPCuT242pkui0l0vW3LYup8Tn
R0RlKaVrIoafhR9Pw4Tz8lfvfyDG3wRFViuxetDDcJzZ15A2DNRCKls5+JZVe2L0ZDMhvnrCjF5l
0ZX7PgdtmiDeCHu9EU5S8/TvOuhduq0/TRoznvTzaiue74DAl5g2KU6v0l186XwoP163QemThLv2
Trw8m+8giT4H6ZwY7zw6pAxydNGs+k4e2t7DfBs7efZYO1iyJfU2kmcNNPa2ZK+GNa6ENYJ6haha
I4LQrgcIxYl7MsoPTzpuH4dxnryqbIfOWuM6xDGGPTVKm03PEGER4xyxTtwTHQk6fJJxjykY7tuh
7tozndSQaX/YKqBqxJ2Mj73ZPm05+EWeW8bPoRjDVjXlcs15bRxEn8FxotZN8oBd2knU7RPqrF2a
ImABje4r79FhYnvSNAXrI4naXyJJCDF0vQ26Tekl9N2eMdeQFSFeZ1lnONzhTm5WSFDzvVCtwkbX
uIeDM8HewGqoX+J0JdIFzfaos6oD8LHC8/6owKyCSApVWSWaqOXZrWbJxS38H8npRZA9ymPah2mH
NahKk4+qgLVoAH3m1b+gFOCuFPCEMSNvIRKBQFpcEY10/ulV4pCkN6qKz3Rt6cKPTBybKOJgTpkW
ISRsK8alFyRtOP36TquRxKNP/afRaUgGQzyzWC7il3PSz9ONg2xSQUd5iJWufW8b6IM7RxOVKW1t
kzi1cQKbmFsOGp2blVq7tt+mGGvGtRSSDtai8zabYqAcgIqk2nwkl3H3PDG8OyrTy9EPz1SbOitG
iBUcELX2zsmG+IpHmJ/5QJ1wpokHOyh51OQurFvWZaYK8f3nWVjw+GXYA+VFSXmKPKVslOfYsgyO
vrXsmq1ad6e4bwMEK+iRtheN+Yp+0xLI1JJJKOJ3bXvcCaDKPymeeLqF2JgatN2oEiBd7rBdyI9v
gerHrFLQUet0qGxZV6xFtORPvsg2X5VpdUBNV7keaMUAhD7ufd3DRS4VEkno/DiktVQxX8j+FrTe
MdjVraODMX81nhct4217dlqJ0fWW9PCicvNxNssZAKE4xWus6wbsFlNKs5TUO7o4PqlG/7MbKa0f
eQBH3+9P5abN8m08G77v+MkGjVgPUmBfGItD/FWgNLgAqBLYGb93yOwE4Uh4RFmvDHGSwwUyl2tM
k9mWxwy/Ok79mi/Ps5Xph39uMpWs1L9PlZWEXAXhlvbc3hF8cSuYYtc276R9oGun1XHzxc0CAtTy
7NYRcIbizRh2dhQNa347Zfey1FEVPicrd6SiYRdtEpeispMrmjmUATb+6gQmI33qFEluRBDqvs5s
a194HEwUIdU35lqAC9f+mSlCI4t/j2pIMKq02SmneSB+A6iQNsnGbnWVMxPmsAILVlRZ/TP9QeB9
lW41ThD/CRyuddc33oaxdIERgRF310cdFEj6dn5L8ffV6gZYMSWPWbg9Rm4gCqx6a7cr0ueiL1cs
6BnixYUoT1E9jkkQcVXZAwvDlQEkUcEFRqm1DFoFaqYxZ9hIanWaAmHjvYAYg40tWIGMfY0E42vC
ZJn62Ps0g/4hTCrZVC/TXVoliN3+SFqNyD0/RFy/IMDFFUR+Yk8iqrIVCgBf7+RM0O7HkxBYWPpX
y7BtsosjFb1rvGpW/AYJ/y0b+rYkbnfpheARCox8PaeLm9YODdsEvNDeEfD3rZeigL4IX94I/PpX
fxmxGVNof/tOd6oNCuvZnpCMaDdoqGyhp7Bcj2CjJre3Kcff1sowkqfroTs1fQzZN00ZhmkPlltg
VcyHDkDlHFA8Z+ThQE9Cg3oUd2/RbS1gKv4NFqBzawh8ZWoc4DaQFHv5OC439FaRIDyRyNiI0v2W
hQGlFxiuQxd0TqNpCbtj57VCZrUIXCBNtvGhOvqje6NrkB0eX9aRth7gBfcYkpGEYOa3V1LAwbWO
2I9y+EuOyypjXUeLu8VTcetx6oFdc8YE5jqnpUvq7wK9vdJKbd6iPT8AnkfPtzj5nbC07vuHbS8V
gvtMKqW/aQmBZSAZwuHci6cyHfc7IkMpOHtASJaK0zLjIiWuTQwuV74i9BNnAKBYDJjb69kbodzp
kXgqb4th69ghMO0KStDR+1gnIacF0mwNXxTHhu7vGhpVANWKhHJ2cM8y7MXpuv76L5U8NH4VY+ju
+rFz4K9nRi46IaNI3vkMHBzSZ5BHKxRQ9J5zAemgj5sCqtrCX62Y/WwCIf9cHVnl9SSUB1FnGkJD
AAqNrLudVC5uYoDdD/hexjQtuRV95m6/veq7YX/mQQm/4QqC5Yce64GJhwIWDQtEaKhcyd/qnj/y
KXZLVVKHlutYXt6PUM6RKp6L7iYAetrAuLdbNvmOECmUr9JJ0UQBf1owwScYA/v8o5MGc8OleUQQ
+tDrt4gaEjrzbgoUE4Z9ouUCOc6BJgeiGMi5T8TySVKlAda6trC/qugdkGPugbxwPBuX6BjBWIAy
e7yI3vrJj4Ke+C8cvPUuwZKPx1C3GZXzsQrwid1nYViHIoDRJqP9dCJKaHHGI4jvvl6hkP/LxlGI
PN3M78+IolQnkS+Z3yWV1aiqUfnAkeqguZHRITNW4ndUIFacxHAI38wVGYG59AXO+/3ANKaUPB4h
Zv0KXt1Kjy4OunldHYswF1eSz1ItjCZf6bSHmfFSjH1A3po4uwNdTyF9H+MF6iERrk2i+Ex8nOwS
eQy1UhfVKTMTcvYeYoyG8YKDun5HhthX6/HRgG1ClreYH5vKf5olSPMqdHuKKJ9PNk4XldrQz5Mp
cUa0C5XlOmnLaw2Er0Krjii9QnCeMianxqJp8TOv7IoDy0QFv1p1j15q2UDGihkzIspV2kCmtAWw
/dnGHtFdR8bpIGFvHW8cNK43xIl7kBs05wbV+JnL+qw11PWPT7X+Oby1Ng6T06M2qn4gaqtYrhQU
O/4hktKlHQrFYF/4LWL4ZzZhIhURhzq0bvRoqiX9qeCtog/6gFwIUzpylAR5FWj8LfxbaBBfu06+
9MuVcmvxD1HPvoYJhi4n7LIagyfRqDR01lYg0UAd9n3xuz91Rn/bR4BisM1RsivLnvxQEpw9AI6f
hrVvubFd78Eo+wjr57y5rraFs4ZAcWqN1F28zA3RFkaMJEjI1LcF3H2dYkDldkMPanA1XTbCvBjx
fGAgPNKApi4hWHl6Mu240ARw+lGIT+45ptilbkKfnnpQrn6pYx2LMtm+m5kBfagSVCZdP+OeA6gY
vXmYz3CriV/6s3iJ4keFtF94WLgwsioWe1podXUvWqz1U543hO3FF4qoALYl+laYU/gdCstKRwIK
G9Uw3qgKZihCimuOqSYZ56MzQ55RFNWbjjfLH0L0vMmBYBUXFfHG0tlHGCEOzsshhZe5/9cwuYI6
DWEUK6F1kh2flGFsr8gEA2AO1YBGzmQ2uTLf7cEny22MH/xwr4UgnFK5mukz73OORUKCBDL0aW+d
GloYm5JD4aDjzjZ1mMmo6172nHZZUN8/3SsUkRgbc9iZGtbDIYiqzjSz4COTGPTFTVVu4reW/mTU
3WfuE/W+PLfEJceD/JIweryqB0z8KHGFBWX6msoWeQMuK/uFnuCQMZwYcn2LcoLl6xdRJUCnGVPC
shKWS5S0c2rduNb+e/v9Isfmj9y+jMZY2cGabRa6xhKKTpncH6PNebdqbdBbObVGhhAEtDQvVFOT
Xooczn+sfRBCeSmpXRGhLUo1PsHsHRd1iAInRlQ4PuT3EDWz3DB9m0cwg0EhViu9iKsx+q2iJei/
g9ZfQjtohBUrTePz747/ksW5m2VWmW2sny66tz3ripf+SpFi/wtRraPQEVKPQCrY/c9SYesG02c6
hHosGIcFiOjJwDfQyNJvWF57lPrfl5tEDqCyZ1Yg9wfhCWuoEUF7BpOwSpfV4cMRD0Ngbw/qFnbX
tn2R6O8F0tqC690ty6F8W2GyoroBl9dkMi3fV0syFKIA9TtM/Y9mMPTQgrs/Av4lGGp/KSA2afpp
EIPBj0qTefB7MEkKai+GQ1eD7DY9UGB6z2UDGsEfEr8cvrbbnclTzFOFO8sJ7HtWU0uGLODA9oys
/J/eQ+0nzT6xJsavtcAqyNLh2a2nz6yTE4XInf6hAfyDmh0w5PWJbFCFSabY/nsPoASXYq2SctrV
peDMktd8KIo3vjBnLVuWJsqhXOTLzBwFNI8kRdw/PUdmGRGHuRsjSUmjkU53m9cIEsGGtydc7DTd
J1C6pTYmdW5Pn556S0aI252bPsekwRBYwm3owstoLTqRklBR4tujJAOhRVMzBsXmtHZJDrQ0uLVa
iZ3XPVq+DVxnyWk8mUfxhSYlevbCB0ZP3vshdnhW9+Pa3P7q8NA4Y0oWgXoredegL/gzOw5iq/S/
6cLHvPpmHjXIjoJgLp5i/YnnizwlybTd5Up6/jlm98wEM7esYpp4yhDwmnscS5rK29VQPWj+jGri
tdv1kQoPmZS17eHaz7uyVuawRSFhE/FH6sb5dEBJlzU6ZGnLUXScAzxY3+PNWYNJpx49H5gPqiRC
v+5LKIDINhrr2LUOpw8U7brWqPk2VXAR/Prch9n/kIGkPmwKq1R2CbHP2drZ65c2yXcaw6f4ub+N
AB5NsZUwfbRbiruKUprsYQwydnrd32kamFoEv6rQnOpznnnGrqB9Ef2ymvcjdMvK8skGWVH1TAy/
LXRBORlyKj4lvnrJIm0Gwm4xLKc5rxSWC8iwfjmVraaEt8+BqeC+LjsI3eIot2M6IJKofV/zPGS8
ssFVje2U/D0CfWRmzpKkZxlwFmkGMsb5ukRSdqRI+E5AD707HIEKpkSoyH4k3cZxzQn8oL2EvY4k
77swmbL3jr22k6U/hS1oM1WvkBb8day82Mu+Ld/b0Kuccfm4rcUVFA1Pa5PYRAMTwbVmC1BJ/nvP
P7Mi4YBsHFhBKRHdu5GLdzv1IE3vcg3O75MbqX145fzrbwLM41rZZEupHkv8K6zoHlGrWiQa8Z77
1+0YoeRs/G+kT2bDfDFyvePqwfq5qwiDHaq4oKzsef+5Pk5drni3mlPGNukn7ryUYgcSCvUOdJMM
hUz7fzNIqFObdnRsVWBj5Jj1FSZvpSEn/aqBbZghz5nXIv8ExFU55U80/FELNaBoLqmgP0qtdOrl
1ZvvKiE8UTbiygwCsEuTLGQsCVPxrkkZwuMXH22+PK54IoaJ1aHIf4jDw0ILa5GNhdffGx+2Kk10
cxHEwzBJt8G+Jw9sSXK3au5Rd+jKV1HournomlBmNvWs7usXDgRVkV2lr2FUW3ARWKLq6eM4thlG
t4mIegdzj2sK6p4Z++wxonWK4iyJ6LojDCqXdD35OCEMY6THaOgNZSohkHmog6guV1PtkINR7b4w
FTQpVzrlH8Mb7dMH0KpQ6T/KhdmnC+X2m2YSH6fzIY5qW9KlgDr5+tvNhDguHjWB62K/Rqd+HClN
BaZI/y5FQcy8GjJ6soo+TYtxPGLr+LcoPKOcjODcI5KV+eNkV9trXQ4J7rz3o/Y3oYDOKvK6LIMd
Hnre1p+0ZUaMroitVFDaq7dh5DuWWz0OKRJ6aWA84rmJjYhloTOo6IA6SlfsTO4sHPJzmy2Qu+XS
R983C0/E+COnlt+xUOO6ls54Z4qoYs8CIDM/SaaiGrCS20RW6W9bwchdDOtj7h1cZk2BVt1bIRSd
biH7n944X0vS69H5JoR3Rc93ottqw1gxRf4MIovcELOod2F8yFgHKoXx1a4DUoKHMvm8Xl9HHOqA
m1cUtV+6c7jBUYcvTzRRZybxyAzdvoPSomT1Fr5mp88TZrgKP4dgKU4OKTguFCZ331ZqJW6cSzl/
4kE11ZKuZsoq60dJ3HsOxb1cywOe/W5TsRTsQKm/QxdPBm8QuMDpj3ciLclMXBed1HfUVUIxeapb
hAdqZ6U4GGnJP14ume5zje5/fQVPNTQ4BnqmPZcfSS55n+ox5G7miCxuwzU/5rUWrRkAsAz4uRl7
OlWs+S2GKWRMn7NQ96KIY625iH+zXLS3je6sowS1rzwtnFT6bMq0zJoALBAAYtyBTBLKlPasfzCr
gGMhXHC7ffG7NO6npl7dKlyYw41tt7TG1iOYEYwjzcrSYHTAK7FR2wEDNwtcMjtmprae+yxUd4s4
SaW8lqVpH5iWETJfjlREAM6lee8eehBt/FkhF+mdpwAfPx1rlfpUb/Rdh4+CzRKrmIl+imzDDZ7r
L9BWfecYI6QjrC1okFbruRhTjcw3ZZhARr1yfRZmrQUK7H7BO6RVs6dGP/jSe0eqWkCaA+Ug189T
Y8fdjBPgcgdpMEUxVVWVp0qWRWtPSa+HYRqMmLrPLL1RgRuNo8Xtql/YPC/5GPxNKYbZ6SmlC4e3
G7+1KWVVBnlhT41JYImnhdJ/W38OkwnswYAhmIy9f/L+bhJC3LP0I/7DQS/bFeSQVtq4+N3YWdhu
fCYpfrBbIKXCTGb2/LaN0iBtD+75V/0E0iYDF7+ZF5UHO4Qlf5vMRvmCDw16g7p1JpDw0s0YVnVu
y8AK0O4Mto+BuOLwu4Ob1UQcIeCqTAcVOwtm4XWT5pS6W+U6lwWsAEmOKZjuE1lZPSaAwBvP/xH+
kxfniBcx6+lF8NBTSaqATbVZungmRAEIu/ip7oLro86pbK1mvBHL0cOTC7ihOLg/RqEHlWTsfjSj
GLIED5IZAAR2LPUmdIHPQxNLCfunLSJpu6hYHZQotY7m1OR9eG5lHSTwHPREhFnbMzbgJq+Vcst5
BtCpRgv5HwL5MhQFwp8ajN6klhS2ei4iVx2ubCAcLMak72F7NYI62U6B0hzbdDRVSBYjtWzINAwR
lvU65OauCGB3ct4ZYF1nXY/6PzYhaCQB07tnRyzI+idrdEgQmCrNCMeGZUJ/IMon+pf7nduvb21m
7lexwxr2q7T0Apwe0/a1+8cKAZV+kXizxx0nqE4tTdXBrbM/CHS7PrfnT/kTjwFBjqxfgrfMSYWP
5e0bS2yAEywqoXnndyNygQP6Q8yO0c2hFnGU1wm3AE1+4GaFmTgqs0X9D6IYAS6Yp19V+kDnhB3t
sZQ6e0tfFcfmLNl2bOwf226zQefEGAx11dPmVC6xUeedrIr8B6ogOnXJq90IFDTARBNlnCyPtXXc
91xlq74zJy6qYASYmo/L9v/nJq0C8yMSFBzMr/8pI5pD9eUw6e/lIkc0Yvhhp1Q3xafBuWLZ14lm
UD7L1hTRt4ZbAA1wngzJyBXkwXtEw1uDqlQs+la99R8Ss/8WMW+nrw3hF8onyDhERaIDAucILSu7
+3K/AoNG7RIoSBm086++tysT4+nW58fepn9cSxx5hd47nXxqXmia6ArRgzorFHUw92mi21iVP4sa
CtTYaiXjywld1vOIOddnqPQUK723w0Zx9hcHx6cLttKK1iX3WzhVclCf63p7eWNCwhTtqUn/R5RI
2y8swHn/sFA+ii56Z8eAEuOoyoxfM9k5ms9V0y23+QagNlX4cxMLyEYPjcmUN6qNwqQwkNLbQ845
d+Udx9fqVv8JNjKoQJ9QS3L7BozN6tY8nkQiOgQPL19wD5OCE3oka/CPUrwLxnsuPy8PJE4vJG6M
WhJi7DA4UhG/g5C75O75O6ZuobrIbig4i423U1hSLmQnIbMX1sIly6Em2qmLpE2oYWcG0Neh+hP7
hKIpWhfUuk4jomXzMZtdKPXf+JMcCJXIrHk9b8LNRSs/5AZzjjLnvP3gYITsGTz/u36GE3gGChs0
NVbZaO4e99W9udy3sWr2LFbii1gSZxgfDZgWkL7FcGsukSOw73yuEUuz8UKRDu4mWwvuBCOjEaog
qRPdKeOSzSxWUILJ+LXtBDKjazcNin8mT7X3NWIfX3P6NY7QYxdEBask0DQ3W4mWiN9PQNjMi12e
kKnqyZPMfA2BMYwUX5K5YXSobY5rkJbE/JVTE6g0Xg/WVWqU3YgcnXL7Be3NTbPSARpNf7X5Qk5c
ah1Tv0kaGhxMn59Iw2atHLylrLGg+F86pbQnyFGfuipMlshW7mC9KPzcwQnEHj3BLq8YK0ZTfF38
U3zFZdvk3mkpGlWjQxjp1NBgwouHzN4QSlwg6lj12utco84vY3qgkSUl1OX1MdWxme8P7csQcMsy
16tGqDiG3d48MgYWj4I9AFuAz4xGr7p0OmamNCgiHnPomVeUXrtlBKJBbQBc9wJeJgXR3We4yiU2
p89vvSGdzc0OvcybIXx0y56OZY8Ky5bYGG2L4R2fvZl/B4RJ5o5smTHPmTXIcj0MFqd+H8ksKSQn
PUib60kKoLFRI11APpI07XwluPKcy1tkFSIn0Cg4vSf/30CgSY0ab7QPEuvNppYzHae+KjADnShj
tk99ROWEr02WBVWHa3PONt6w+EjrdCUyB4r/NBEAaqm8ybHZfRH8/SmxM2OtEA+4//RGqdOUtVZE
PJ+Ixi6rqnRjvS+w9LysrsRtu+NInR55tVTv6abZkgoKC/obaT2eYAaveAgA4CwyPTHjWq0k/2MR
YR8TlWdULgnzgoCGfkM6bTJUi6msF0i5C1P3mElvgoiXD48JI0f9dBT5BU13ztGC0t5XJDkZKOcE
a4w0b3/7JLIV/xSOwsfAZEtyMfw5Jn9bT0iN7hJ/J+Xrgadm+QFncLZvKsIjJB711D877cJGXBsK
mIWVvnl7KiFPn/hZ4UJkXx8js34yQGcKSUAYI6v6EGoPbs8GrunffGid0mKDhxKrnhpYPs5ZPtii
vcPXcwAAZ9TnZav24uopW2TfwG5iC2+pOV3Dn+65SiK75RVrT/Z1TVcBRt3vC/MZyUdTtS/u72Lw
YSCMcieIu3WgBU4MGbUkEBIYxDDILqeNeq1RBOvH935bL2OEtlb2XyyQWW/lDB5Pxowj+qeoByrV
0gOPT8OaCNjm4NkVKdxO+EkmZVj0Tx8gLd5NpKz/bBSUFyKatAlfjzZzf7go+6ORffcZ7E28sVar
31xFX6AU5KyG51xKVxxWPxkITZpPrYnFlSR/rDW1TkFxbcdVJZug9C+fW3+Ayjx8L79SRqGp2iTB
EmG4dK37JaiYrBhmnpn8B8aEykm/MRrXNrysqBNV1FXu8rtc9b+Iz3GvH1SuuoZ+RcHbnSd6s3Qd
OcUJU8VFngruclAYrwdtrVUArPaVykzwBqn2EcdO7nNwKbhbXbgRPNGcq1Uguw2zc9LLIZAV7M1f
lQk905/V9phUtXDPAEx1pFropG1hDdIXArhNOZC4TpTtupsyjyWKlOGPjkU51bBGpfm07Q9xCmko
GEeHToA8E2P7/7YB29U5SRaPEGUJ3q0hQ3E6CYAThSSewWELrthkQSSTzkKccvpwsdv5g7ypAz5R
Zh86/oPI8IO/CS1LSfpb4F1lrHeCGFK5OwMaIlCsrNIpDyjb6kb8IEHZqntvI57Z6AvMMxQPVaQb
LB+T1iXHExE4ve7HEXVZ4hQ694AqHp4/Yuuo9TQyJxMy5LvUDv1sTkL/dULlnZt2dQFiGx5CL0sX
fxyPLyoAYwgcOx5PDNd3gKjXewf2cJy6OX3cH9g+FCrsgrELJbO4W8PbzJYLe1cYIOtoqcUSZdl/
ALRCPiHt/sYy+5dCtZrMGghxtjxk7O43/9nWQa2+IDeF16/zBAWMAxDgOtAqu1xO3GbksVJLtUsL
hb+Tfv661PhKt9R8BNtzxPGFoqPzWqyChJa1sj0Awti7xfc1w00AL0NmAq/SxOo4dfbL4QsgjhF/
I7ZkyO1CSo5JL3VOYhTZzM3GaBflzKh2yRA8nc66OIm62vGwY4R4Jb9nWPikmiWqawWq5VVRdEf2
i6OjgwXi1tt/IITBZL12Ghdl9/81iLh1X4/Hc2EY/a1asyBFuU1eSGGZEfUtzajrWePUouNB7dXi
Wibi0g1BREp4QLd+QFjylij9gT4Xq1RR6vVKjbl57TPiFA9LAa69u2oqb6VN2nOsn8s+KRAXQjd9
hLEaEI85M94EyAHLPxVPpNFV95TRSWCWFKhEUTqSWL3ciIKh0pVUx0nxgGMVTOLY2YkHHXoGGXnU
ZKFroRPiT3qkps603bxElRydIjbX524lf9qGn6blGADZtQu+p94VP9SsIHqbIU6SYkX5CpL2//qr
kMS4mzfEDP702KUcUw/EIB+QNJyfbRenvafnH0zGiSimV670O3RUYgfq3q3pCj/YhfX6wI+nGKVV
YrRm4QfiKC0Ynhkk3/sM/fM++bFAsVIlNzkjWFuS8OC4FpYdexmNLhdsxxpRz+CupCOqms6YWPP7
4Bljn96x0m8ZIBlI8EZ2aio3Bt94amiJs82jKayB/pb8i8pFmT13ZqdYLDLuqB9pdKOcEgXkWBrf
w3Y/Mtnfdabopc2CeDhZqHLgmYQUm9Pb0mNCumw6bt7Ym7VSk+SyXQ+lj9BaTHB8CBn8JD5qT/Xf
jhPkW/h22VWPK071KdiOCgb9mWZeKMBUG5bZS1cd9KhO1C6ggY+mvQUqc04GfdnyrOx0sXtgsCqq
Z//NObXAme0R0fpTtoNS3HAjfHsyLios5TS/HFF0puMqkgHyE/cd9qtSWl1to53EDEghan0chuMn
EiKTTgBbjlmaMTqdmcO7QHmiVGnE7RfnA1CmbF1zE1/bOwaAGNJbgkyA/NLNVtCq5O9CAV69kKZz
5O32bh+NE+70qUBcFXfW6rX2XXw+bdb7rTuyW2rdW+lvte8tSWrKFf/meJ0ips5Sxaf66dXs2BfF
k67F2FP3duTvqseVzRxF6m129WSuJ/8Ac7OX2CfZHvjXbYx9N5W6K9/71lzcMVioD7cKeTmZ4dIk
EJU5bfzCmAyH9wY/PTGlQwPs+pvuHo89ms2/wezeeoWuvS3fnL3nHLFflSlABoF+oFIP0XRd/Aiu
kPndDdxZ02Ok9b+UpO717B5BGBhKUf2p8HvRyaYUFEL5LS+tbvx0V4XhS06RFeiGehhr550UQHJW
PwEsZn6xKgzyOKGAFLuVGGwlE5vRM6Lqm0Vs6eAOskzF6SEo0IVZOz1IzLZrC1Qp4AlIE+YQnqCx
R+GLu+zwSjSAT7iLtc+Wjj+qMvSHxIH14Z+7PUft2F5QLPstfK0/I75p7ZP//rzCwbevwpqGmrl+
sgnpPgp3WcE0y5Hd+nbN1JeWZ/wN+tcJitwHPzD9al1EDrMGkbWdvcS6ym4vdoY1xYHlVPM5zrj5
UIXs9qbh1dXuRxGR1YhLjqdJaqoKYhJtT9HMafkKsbKHeICed/lJ/N+qGwFMplRm7B1lTqqnXPdU
pwBG1akBFuP++Yc8pposvjIPY/9HNWLRZVuwq9FFtOsiRNzoBVq/1ktuKtCqSPxUyu599zqigFkn
5GW4GYDU+t/yNzjLQYmqX2y1C6ite+mnXgUtPsFetIxzy5tNnXFAf2mm/pbNOsgV++FaAi/vPNAX
ezxycm5jM4Yo2g+44mDosl/sCl9VW2JfBeB2Oz+pLMr4i4qNr2T8PyGqqzzGrCsKicN1/RoeYpT4
509khy/VKehjAucYu0DrhsKzg/kpch9xe5UbEcaCJre+MiUBUmreJN3t6/1fqd44fthdZiG/lDtG
UX77iBywpmf+/AF5sWSt9PR1KPVAkzUkaawkADmpDKl/AbZG0Frm/FMuyl+/RsLctHHwpFT/h7Lw
+Uq28+ojGunQHxwAt/ORRCmdL/RlI6YHBNDIQACSl0bMP6yJQT943iwlMo6nHsV9lHk7yDsa2FOm
ZQbmAIHEklYL95D2c8JN8tMJp0gjmIyzzXgCbJJyaDcYw753XaU83u65WPQD2UZFPd3/M/SgxyJB
zAI0RTPYUqnc4mZtywkoq4lCjbTrQdzClpN8svV7IaogZO6XeTiZaLK15LhOYtqTtWA1jwjFEMrx
AZF3GmQCMxRHt1vlqNOqYO9t/yHFSuEfFkFu7LRxnc4+1zTpIFt//dJ5gm4nCnIWgsiXimUGKRfl
rAcdue92FQO9MfNxEy7Uou/spvxRgCZy6vGZfEuDT8MQvuZ6NnlbiK2niVTOmxDSqJBP6i0rx3em
Plm8Wcl2yYIMNeLatElEZChcnxYJt0KzTUDke4YREscUOqn8pqKKGT1a2qmpwkV8dl3R2m0wmCUF
VdjpzaqiNk9fpG2uQcsQxtghlkWssBvusYE+l5KDJjS/2NJIcYalxamNPGeQFSP6/sYxcAjBeB7Z
Lb9wcRGTQX53KqTFhLBUNGYCYlByC8rIaVlr3Ry9m4YqOllxX5M+XSMOxwGJg5jFr7vKB67ZK+Ou
LsL8mOTy4UlySBI2z1MNISEfYn3PcQgNmWbwkAioSlPRfhAtYFEoMuz3ozzW+9c8H9cT4cA7tNb+
naxqA3NppImPXU2+SoAzw6SUVEVnM4uO/BVlXhIwFjYBIlJFultjcwd2v02pCRRNtGvd0sM8Or3Y
7QmKoJYMLhWdhZu/8X1V6mmYAIA4w0ynqYixhMDUFqhS2i9F5CQtGyz1JnSAsQ3NXvZTIoPgcias
/KQU0bZdC3m37HBVQ4aq0nEy4KmQjdvVtoD4r7io1trf6aEj1PWVX7niuBlHL5aJkVZkVFpOEcNJ
7DYMoedCQ3fGfX+Z/J+M97sF9hUHeB76ZOKyiCUGVyupvWdcC/vgjFHXvqa4DpzJbYmfic8OrVws
G49xN0FNxNXpef8XcUJkCXQrbY71D/FLsMubqW5lPqjSTS48pr86MYf3dOw68TBQ6+sQ2DL2JJ8Z
b+k0UgaD8L0LgUrgb7kwLKQG9o2TiI7cJnGX3xLaQs7mJdifQ5u0ytxNFz50Mw2WnQG2dCeyW4ho
2NRDKL9F4YQGGlHtxBvQJFG98aWEfc55SkSIfDETJvO/DmD2cnl3cbode/4jBliOqloofcZNEFSa
2sLvqBN7lCl+RDghKGImK5AGUcvm5fU8t9MnVnHzLxr3UrxpNlMOHsysr9R5TEBe25kYX4lFY2Td
E51TIOIw7XagxCQxcqS94OBB4kEJtWEOdPQW/D2KJTL+1txc8D8N2AlrenIrEYkFMUDJPqxwqMgB
uYLd6L5M+XZmrKircBPSmmIqDHW+Gs6j8QnfukAuXANOPydHcWlpm117bmKfen2JsczqBN7yYxxO
xq9ulDds+MAVfy0K5cG9rl5Ceax7uSqa+00LCOj6BTURBfYu8uATpAR/cjJAk1VUdoowmVXQQS6h
VLr4zoGwYjv/uGOmVXGh/UcBLkYZfg2bF6oSjqSArVHnCGeYPwuKGoQcpQBIv1roJNupNDPL+JLf
//CTl3Z3bO9NM8ClIuwN6+rIWzRq8iVgfZQLBIxKydFR0hVkoW+yHZS3V/PBL/+SXu8hgFMFnm8z
xywcmOii0O+0jCjVao6BfSYOujfWmksq0C6/T3tX1+0z8kFHTUPz0uEaL6WgqRLD5aHhkLRKBJHK
ftnd+3n6/A0sDLbAt2lYuqmmeOIPw+kGZrnQKhy4N4kF0tchQTc7RTjQGoPUJhObfnWa9UJgEsW4
VHh6le5aIy0ySanJU8UeTqouEB3X0bVcsqU1mcUDUfzopaPxwO9obkA2XhYufjDl7qGLyvPuXubw
Eusq1Ihmh0201qSO4i4ltRSSh5DTJJ0T62Ul/LLNKwvw81tw8CsgVJ9A6GixPu/zfIySxf7PCaiX
cawEZJ47lbaQAFYljt0EkniwtOIcnDzS1lmzHTUA43RzLpWPfINlQg1SFFSJMpKMhFjfUOokXW4i
HXVF6RuNxGewfgw4xH6VVWPQOm1wbgD2OAYE5Qdhyfgh78QNseSgqySqKRl8Xz3r2EzogDW4EcJz
tLSu5KCaOVTXcatwVuVjeZdqI2w/v8akj8avqng1H8p1aaWyoXFKMDJP0V61WfoENCmMBogC4M0G
LGKxrOCuy94RgpusXQGYVUWje36Pvk1w4b6BoAtHTE6OY1TaL/qIfErXSZsQhN/yJhN7t9oiJbpB
wHlZOOdfjBqAZZNrYg3HXuNcSNtGQV/6AMEsM+oX9CH7QWl0kZyJalsk3Zz5hHU6WSuHJ6evcs5n
p+idjKr0P4xpfKVDbCVTR/tSN0XBhSdSOpmIfOLsKhQ8Qo+x09yWA7vQSyj3ExDbkjftw/7W+kyJ
4riEp7Xewi5eYBqRe53oRtRgmdiM8MJYb5gcz3fWYWZCWl5cg+h4SN2e+WfhsUnsvcPAmGS5otZx
Bdab6oLqgY59ehwbJnDIUBC5d+dvvPHoe3V9fIiVcr4cWVda55YrCyMCUdbgR0tqkodp42XqzJ8m
LMuCkZOcaZAc70RmSiNyCJ7haKXC2z0whTiVDX86YLvK7YobqqtYE4cyWXnwqXsvVbivBPtsC0kv
Kc73c8pXHGvvc5RjjnVi+3VtgeT8WgDx1J0ShrHpWG7q9xsKu77xhDD7cVlsFEPtMLjgwFvA8YvX
d/zeqNQBtFTSUZszjZIndzQJLX+X/FgUeeOjQkCKCpH2lY/pu4SCiS8T/qXoDjj4euD80rJE62BL
85hD1l4Ikt+HSUhRK1GgRV23Dy5kRD+dnhw4rF1FRvILePCYe8i9t2mq0AuENT36B/BvCp85BAPW
ckVSiSV/LJUnxPP44fTUzS3oeu8lMdTf+oSdyzWMJ8Vrfx5ammq05W7Gev3wLbyc1zj8WZ/hAh3z
zazxQXnVRR7dWbyhLCkGvX6rowtanHRmgA+843YL8d0tWyZf3/XO2Ux/3VrKCTm+7tBnxisLutQ7
K1bD43vcrg7JO0noPvb4krsz6oASWStO4/5dAMJOBDDKIXc2nSXAKQW/D6S08mOlAxaj8iNRv7jv
nId3jFiKeyT7NVD9rxMWaC/D9fKKRI6Rlp5y7YD9KmvhX0yxZLyEIpz627RbhlkV1SJ9hWPmM/Mf
lUx1OzrDdGV74ItppKNCqstFWNTwB/dRSH54+GWOHQMLSgyqtcbUdCdJD8PHvAaa2Qq3A/Y0FqvT
3zg8svjL4qy94523Xi6XUn4B6JzEICuAO7WuTWwa9AW1Mc47WduzPZtJXEslxzzkNcbaMKvwcvTf
fIYK91atB4o6/ZDXCMm6lWka446vpQr58qQiKCYMYlKaRIa4rEFFbEkTmoR3n1JE0OtBFf4FH6Sx
qvaIo8rp7v2ZgmTuSn2wPE2KJqZVX8+T1ER7SSbszsjUgP9Az1WHwMnscJhJAdptk08LjlfhiOfP
aCox1pGXBnY1l39J5DZTs7COxDNFEp9YsSVxc6aWgH2Bw8WbL5Waq5pC1GZU2hxAa1vFANMopDzE
ll7mKcVRlWx92/ROKu4hhK9r6Dg5AbZ+PWbkPKcnyCTpNmY1qJI4p2k36SC2oQV942EGcCnBwcHO
cNgGm/T5jWuC80Njc7L/g2ZoLyXyZMRF6ZmPe2vwPyU5qQJjt8zgnr0w1qId/o5v7wa+YDN3zNUu
7M9kD0XAQMLx3DAOIprCkGDmQGquw4n4nCiDT7SV6sV6hpItm3eDt9XZXBujJKDCJO33biX9hPix
uRZWqkvD3ZxNwZR4t9hSHYKxHChPhXUlj6g7ejNTcGHIVu5OHyExb2zzeEgawP/m1Q1gzNfKComo
y2gJr1NyDSngfL1oifo9IftXjp/M488H5IyHzzAT7rgnsqEPUpdhpeqSdm3hIKnpHM5/89qVJsg1
ZFVsbjMeBhB728UaY3WUyVI7aOK2521d6EaMibGkVGOOAEVjWjrSHJeZO823a3jF9ISv5lNs5eQ7
x2aB9aDSgabYd89bK5HvrmEfkEaEPL6xCy9GXslG19QyS4k8YnMl8NXgZlMg60OCESG1gAKH0B/H
dwjHs6x2gaDj4RwzjCfiUKrpXxTcnUtSrvQC0kqLr4+CFeN1m+yuW923GaS5jV3bWNYuIzFdrbsw
9fpJ+21qj+q4PYf3B4zbOdnhjhNNhxy7HTo7zffvaIaCE22JEkz0Ky4ly4W8pQjE0OKwkgzoqAbu
ecuhxqqyDM/ztqNcYbpNJT0hO/maYhmNClFpzfb2LjkV5ETME3Aq8u2Q/7V+o647h34WNLCXLk7B
5IchF11h2kIQe3k20IQBbbifs10jnNIFVbrY+0i5a7zfK5Txa5CH6NJTP8y/MLHcmAQBByZQdOcW
D6mYC5YxpBy2XPy0w0juUxmr2DIPA7VKJRecknoL1vuuoynXXJW90OM6ylPCmA7RyrZToXV+D7jb
rUnK47bY10ohuS0QeYDX/NReYmd49KFRG/aP1hpLBeDdEgQYLmUovVMpAjikO5WnQArmAXXWgbb3
EytukFh//Js5nRX5t2lOIGE3YxVRCbip9mr3E+tH2b4CTBEDSmXqLLDAbMtwN8aC1Heb8YRBRG1O
Zu9bKsK3OiRrZ92mX6R8kFHJqWEnMMk/7BvXEM5yzNLTWnWVsNYDkmjpN/6kvVRCKMnmMFtuM3Tx
54HsSiQ1I4wTTk65QvKKv5eE5DkicfSyuaGFmVCyNudHoGQRGKwIsDv/M6ttC+5kTlrKKpOrYABU
KLhPmzNeIFsjdUZFoIsHNkivIZ8PNvMMsGXCzlYbPNjhLk465Mus67+LryA7TsclAMRQsh7FxdDR
2YuH/B1fH+4p7NkFrfPKe/FMNJlnrPbTjC4p1Vd+mLKTxEAk0EaTEE375JTPaqg2ft/N8NRmtFu8
Lgxcf+e9YQwpDyZgIhsK7oT/WMOw0iy+E66/0P/L/wL+qXcEgqj+H24MdhdAZiNG+8a/STX/Q0i2
NAOhh+kkzs3zxNfk12lsRt+Mf0IxnaWXdekqXBYMLlAwYpTDt+K7X9hy6lK212gBo0jueGzAHxrV
j/2cars9fyV6PKJLRbKsGrrkmbCtrV3zr46+AXb7DtVJlZmFAuyluL1pKL7116yNQ4QVcktYEG+V
l+KoEl7Z+t6u3G2eJ42eRCM8efgC+zhn54Is12aNLTZ7vZUhl2bXrhR59hUBkYCAZjcOEKayplB5
JZ+DvJjO7e3sdmCVe807srT2e9E1NWlBzIR1eZLOv5N8+p4UJwRBl/jxwlbM2TQ08OuPQR0V4lel
lQqavty5hYjwQHWx1HiPLuXBCeKW8/ZKl3YfcbPsji7w1VVF0NOLKHchfHYi7Yqre8GEx+edccF9
gOf9qqffKKFb43kjOCLzZC3UTLJo80sNDtMkjtzbqiNyC7gH8XyImTzFOboUvJQVfWp71hNdltEz
G8m/sa52mmLGSRnz51TMYriBUP1yi/prKYYkfpe/CNYJbqrg1Ma+NqF9ESO8heSZbLHLk3LTZXRe
vhmQawEjv3x2/7ds0ucPJ0ekCNCYsjp0peKX0Mxf8rjZVh5pKSZEU6A5F5XCKw07UPwB4lFfpf8H
lPQsjYoXL206ksilhy1pd0CnikXmqEMvS3SRMhsZYIlDyKMpmOjNolmEjwePKp+3FKjv3jJBvXym
iBGsRL19ieEklLmJnymqpj9SsFa5nBFYDwaGoCSOH6tIM4CZ2QGXy9i9Bwl9ILjM3gTBCRMOugyd
PqUmBKZ/GGpWAj4ZhKx2ZbFmyAaBsGD4qkH3kyp5Ej0EPidq2uB44rRStBUCAUPFQf/oOC9C/PMb
AxSvoBL6IrRfSg1J16NUS0DOBSwBzy4OyEPvdM/byvCh1uEwMbJcrrztmEUJgPGcNOPr1e6lHUsz
+H2qUPVyjzawTT4X4zuW8Ao9HiHY6GqtLVfSUVN1HPzKACpVrxEJxxVuqBZOTMnwcxTPVM+GzKHI
l8O8+tzj8vKX8+T23aPyfl8QJopfr9ViT1OIqSTKvBwtjRFp8w4psc7kNBPvTJBnM5PTyZnoA6ZO
2ws7vEXsormIdgEbYRyTkWPyyahwYoNIMym67jpHWbwjOS5RnJ1n6owKvgeFWC8StoKZdgkjxQUw
kXWAW5GD+ksQkwIvjefmJPvrQfCWFCKHI7dZEVnNWom73gIZvZXYb0P3mNS6XBSqqJWe7XU+eHxy
lJwKLkqiEL1l5big/73ymXDWhq86GIW6fo7YrOfYz/ksJVV/NXydmNmDx//JHRVSmJfqMLJ4KGef
aUaq7F6MSXkQjUYOnvPY4hLhWuTUDiL6PoPrE0Y9JaoIarMTtUW6Q2DkzeMDk1f847j99bS1fHaM
Hes6tTKEn23zfLjtITlhLc+g6WwA3dxxlolIiqUgiwVmFwjXcYY+rGgZZMDzc4Lb+yIAShtcxOP9
GzDa7S6o64GNKufm2aSW+O77qtb7g2+IT+HpEtzqjZN9BvdEb6p9XqjCAAJxIyDEtYi2k6JVUHQc
DnhkBZsTNJ+Ul8jKMIoP7GzH8y5LTvdwuGHHoUOJVEAjnJQnJ1qmtAjuudMXoxTnZvarPgGD2W6o
I1brnZkh4RHi5ZHQmwudygdWA4l0tQF9qOOu2rJDe6JlW5R6pfMEAkzTB6y3r5yAB8Mt9ZLKjWTo
zXhoCqg4PKLyn8dtOgOHakKBGAdKN1wCWTz54TcBv0JJiAIEopY6/iqkTsKArSX93swj8UN5JPZr
XYQK8JfR0GZRtP2tDbC+drKp8pvKZMcLER07x6S0P9G7C04/PYvoe9++0X0xQVYUFPVJnMcotD+l
oABON1YrhbsgUHXuTFEWNQXXteFonQtpKg6IF8vJJFIuCZOOvPV49qqPofsW/v0au5U7/feaoXCa
bNAX6pIMEdOHpOyiLXsu/18+EWzInUrOxyZjyExX37qqzhgpv9Pw2x58QOqAMETJ3cClTQKCc+no
6NBNsNIwdep0AJp+36BAuVky2/3ZfGzVt6gm+YOYVa8CkTF0zVOVtTkC1At9vOJQ09B/NETPeZyG
VqM0mAmKaezOSoe8kd8X4Q1KTlhne6LFC54zIvXW99TRFl4bnNvx6TqWg4A2RmBarPUoDfOx+1kS
B4rTUK3F/6Z4GQPd+ldoaARAEjX20mAlumMLvmvGIk4wpdlgguCDndcxBIQOIr6Y8a5Zw/8qW5ZE
GVer7lQFM+TKqUAU7io0XV0lsk5XOk1/zBYRYEA2bzra4PkN2tsDlQmbW142NfYROY8UpLehPNGt
i0PEJXCqePBEwAkfVI8Y+FqqFuoku0MapSEBYrzQWrtXfrHzH7TnwdN5jTGI8kcyecsxSu3KfrvX
SbCFyFnPvygbuH8BXZlhNQSUbfb8bbeTb7q1V5SXlVpyjc3h8+GEEKNOLV5308RPIJm1ukmqVefO
E+Gk46NuHZYswEGaQlQWgZWt8E5gUK0oj4E3xsl1yNTabmkUIjZRdTV58gwxl6EzcBQS/2OwELjV
VtB3TRGRDy3iZEAsccEptSldGq/GjhdfNWJ9Al+LDACK2KFPNyXbOQzWfD+aRKyZrGjEc7KVvoub
wrXpUa8E5aakiRUIr6C+GNaSmrfvvOQrQIf0FHLFOmJzrbAyGlVLLOw/ETZINy/0aPL9nu+ARxfg
MI7ks8itigxrtbbTGmy9EDJOeMwgI3jjEoe2in9zVcuSODVcrT1Rv7Uka7Yt/t/E4pMGcY/IL2TJ
TO2/M5e0DbVNYWKYnSTMlottJL7vNPIgtAuCFj3YxstqGApWlvEzBnhCld79iq2LlEPNEwaUXjIt
Xf+O7IMSpvYL/AktPoSn92kdWD99XrXL8ElnQYi6eK3IFn/RG8VUtY/B9g3Ipy60I9BZ4F1vq8Lo
gIQ6Npr2kmg00U9tIRsOwcVUgI1djyr8ToPu5/8ESx4s7qM+7rEW2Icwjj9piKh2vxeXEQpzS8Kx
y+hLJgFlXaAstuaDRkFsG/UKL8auDe1Q4Jt/CDhQAtb/0drgnKONwdsdK06StO7j22wRi781pfsL
vYjjf2ZIZoIQll3G9pqOQco0hSmoRvZ4mKmFMuYG63/3DYzrLzz7MH+pkNcrHnOVvdvpKdDgFpEK
MjSSHUQcOuScOexq8Mok1oF2LRzTYxEOHkydmdf3cZEBXCvnjc7iYKMdmp4UzlO/RtddKC8Oh8CQ
pck77lL137mqX8aRQrlvKUwxcTJGetays8Fm244hZNScqC4A5uDuGbb2rOGkdS6OGSfqN6cFrchn
ajAZQN+nTew38OrA7BlRiKg31VaekvCvoc5nwORKALkDx9KWSpQKXdJ3XYhmE6DAp9o0q+CPC/0n
a1qXde9F0sQX3WEco2++xGsnbnT2rHmBXAao/fCqRATrMgqW+O7yySCMJn2j3/iFrNXLhGADxi+m
/q5dToTmXS8AULi9TZAT5AaZssR+2LgiaWBzy9tWjJQsjFBsIM5xXFSUtswPf2F4Xc5qbzdbLcwI
mK54cJgM40VJBPLpp6FgoboblR7AC++EPYe2OH5JZ3EC9cVhS5vpiRCOpGzD8uSdE8wPHv5FMEwy
FQYe4MTZJ/qxu56BhwitN8jOTtHgjaWlkxLJtrYw8rJq0JFovdkYy16fAfGEdc8IOUVSmSR0GFpx
x8C8515ISofes4uNgEgrVEl31XpNvUWDwlnNSvv9GkX2wba425HHjAhPJ4qpD7/D436PEi2QSGRJ
OiiNS0zGCC/RVTXMUhR8cezdRfBQIvoTezP74fjpM7dBBtBwyl1JClgFZEyNio09NJO6VjhKcpy1
wnTkBzqHfnrcJ+s/GXj4tmtG4/5gn2AM5m9JNZOW6GbmWKl9w+Hp3UDrTYewnVcRinmKyliK0/Tb
mZrScKL2t8c70RTc4FqSFpjg52WSeduU9T+XFN8zsybQ3gmqj5pHk9LqyB9MCIddMGRfy5nS2ZXB
blMsbhXIh+2opPYz5tI9uqzr8t0+QVJ4XAvG1PVlnvA0LjK+oVWeGyvR7XN6JY4lbei3fUzWJBvy
oPSaP2nKKm9siR4EIkcW3FN+eOV3J/qn2UhlcDaiIpZjbB6E6H77zxg5WcqYKBkPFkeVovgdZwPa
8dgBFh68Yt3oYuKdNTnynOlkTuxnGVvUaOAD7roLmGHvdAm8RFvVZ6OOKjDuYPkXNhUKfB2gVoBq
DhxrqSaOiciSFaOB9ZHuCT0Yk3Kl+Yx+D6hXUlOHvvxe7H1VRl39XR0qF8GRdOU44+q0sZbQFwYK
L8CA8AUsyqu4Y0YGWgxj17ITkmaDF91TH7iHL18R7mmLDp7H5g/U+ZikWCHLXbdg1sw+kXcUy6vn
M0PT+d6/yTrjZE5IQnoOwFJehRLcCQ1b5KdZti2CscO63zAovCAnHoNjbD19SHHSSzFtEVrmCqKd
R88jMztVeIt3BPx2ZnW0sMjiVs23Ow862JplNbbJ0cMULel2IrMs9t4SR6lVwQWnSGQufE8QEwTJ
7FFWKG1Stcczto7Rm0fFJYbh3Cz66B8VvEGQHhQ4Otk8J9ITLqDfjL5OtAsFHPQUvVZLXy99qaum
N5XfGluH/4nBd6Cjg8SI/AEBBW3aTaUeTgOOyXl04zaG5iGKWUxQeMz2Hv4rtSaXBD3CQ9BozzI3
4ujMx1Kks2aIzCOcwNJLFhGoTlkTHr/R6rTcSLScCuLoxnEdkleVB0t+0R0UPQQcDpH1+zMEKNOz
5y8nPPlPqdTI10OECMJoIjHhx1VyHzdj+n6u3YwPF7Fhrmc/yfmJISy1htYN7sJL+swfgNp5Q3gX
wPFMLjJSjKYrE/EE6YQn1VQmH96MC6Jc/mEK6u7JeJAlX35OFCoSAa/Q8cQdrZ47FwVaNanfqnkS
U6z5QzxrqybGm5/I0g+g9Toxf2tTwFbxJWIBQcBsWMCX0xklwpuwXEcqSldp3KqmYBewJv2FEyWK
rpPWnuH++GCRiIsGo5Iyebwkjeza4xGpIATg5LRhQ5/ErnYpEsRUsUtlwY009a/lxR5rqttteHOX
NELt/jYIYIfan72VR8dfodMeX00Iu+C+a56b5gdDBs9ZeFkfkM3EFz6VPMBuKS833l8Bz22AZuB5
LOmR4xh/YuGUfMvSKlVlEyOJpFn8fb+0qrRPHqrfDV1ZQsP+BcvwmIAwc/mE1YAVyIOptwfFOoKf
/eb62sO8kmyFWoZwOApS+6spiba64Je0lkcbQ+cgteaDLy2eK63v1KpETWkI4Z1PXOjez8wi5lpK
9zoSxxP1N0IcuMaJstEUufgTC9TbHvbtoGUh88fU8caKW4dVWq2eq/1EAuS149zm8vu1eA2ABWxn
SU0cFgoTHT7AEdQYI76CiBWPH0yH6Jb0GDJpUCa8oS2xfrDYzheWcKjtMtvl8vl8L5epdCDcSL30
CLSI205c2ZZ9I1edcaAYE6F2zGTHwsf0iRMx6AE+x9k/CjrgfTnMg+8N0E8e2Te99JxbUHpjiTL2
AHZ4m45qK82u4rHpxt39HCh++6QqhFlnN3pwv4Xqa4guiTXirnPOFkmljGStU/UQQyDxVrT3yom7
YvcvgtOf8u07mdZlpl5PLSnFWKaPujp3Gmxf6dF4p1eTMg/RNUo/1irQ4cjSGEYeenNijOTN1qlj
8pqb242dGOIqe5v5EMP0vPn7my0eyG/7HQidLgsxYLDRWL0mmYU9gCmD4pSNv2xh3YSVU8FKYQBR
SfWamSo49pvBKrqXFpFw7NnKNLnigIbUCKB97afVMPW/EPQe2xgHNpaXVdQzGXpfciIVQ9+rZa3J
6WmMbrZQwTHomnqc04K4qGwTmFC+eKwvaI6vSinNl7B1HwPrJUdbcCj5+E6lOyfvYg6iz1s5WM0E
v9+eQT/yadjHWF8yQpoS7A/qMtNqRgiiqhe2QoEhqzdAXW6qQ2MvcO0FmwiIm9TKQ7F/ZegqlFx6
YRLerCGct4iVxIznnylFyhjroRONVzzFUJgi1DdJS1JdSry9Dz7RpqJQN7lYbM94/YbmryoRIbKE
er9tCBSlQ87upobSOSaHzYw5+XZVvy3GqOsmMn52Q/DpedP2HfSUnm/uA0qiyBYnQqskIx7RsfiT
7dCGT7c/Hc1kATUMLB0NlStwo+oHP2Vvw70KjGdV8wuNTSy9JZ+U6LxiLhw+btlM0TNgDc5tTH15
nub/kinc0ouc6GbRHA5j73ZDDDCdXjri7M2+HwGkl7AG/Ne48OasiZB6Kre/sDd/Oef3sBjT1O9l
DhqFovjjKYWygmlalpzKmyDdQXqen4zJ9bqv8qIdVCLzFidmwOyRrcJ9njs9KVnrKWYGnkseeAb+
l04/lItqFbzcdo+VTMu5ZEXQCiChNPcaCm2j7OG5Vy1NvdDz647uvrs8bDSxvt/S5HzT6WXTDsze
XwyIBPTkM8+MS1677AR3VIv1xA3/MK1Njc3xxYdY/ljXyQUEeJnbhXRxR3xRep6StCpUzBscI2mH
UWLrkltoSAqlFzxJenHvaQ3va8l9NrfaZYFmvOE4RuKxDIOttqHytFCWXYkNwUSerjQ7Vuu4ki/R
ulzbepVX5zju6V+mqbAvAsDITnnRcEa7B99hWn5Yj1uyL6nkd+WfTBBZ40RDB3C+f7ikJq1IbkQl
cHohkI56h1m8h8xh1OzEI2rgCBIsYi/s9ceFOyjAc4VRcB8Me/Kn4k5oTkvUjdQKXDpi6wiAfZ2F
igxDx6lfZaZNtrzCESEWpisKYcyPDsaU7M+tzqNMExaV7+btxv+jNfLkv0Vli35u1QrK9IhUdi8Q
3BHlsom5eOa9sbGDEZJjeHjji/v8xKCcbafUwWRpXq1qperlzQJMGTbOI4TWsEeSXp0lQXM9nNLu
qMez9utDaI1DOFMdxBwS0deHa+MWMuBCmbk9VLTXi8cx/L156TBERZzjRin9f+y8RCxZ4vii1xo4
m3U14w5cOGXxIquXyJxEjvDX7b0bFh7WDa3fgtvMKr+SsnPfT3uNfGbIYzPGLuGWf+Mv86xOVEwh
urDFcU1fiVUyaYbpwSYz4srQKh2aA3937cciHbmYgaSOMvO7/LCV+oNekmwf7+mK8+4z82VDxhfU
0nqSUDbrFctwNc84TjHhlvm4DVWEpIHUmyOIiBKAZBZ9RXzwt/HuqrFEGNJGMF8Io9f7fbdoGgE4
shz+By/aAtiCRZEbA+cBUoOpv8HUcWc6l1Vj1XCKGkXrQQmgAMaCyAVNs/UucWr9L3EMLkS9eLBv
MyU1sxUdgtfl0FEw49ephF9ooUTpi4KN8GI9GsACVDh2BG5KxCCMphAJfjDA6meDGC9T89dgtwpk
5OZFlqOekfHtQ78wUE0gX4Rh7XzLM08QR0IzjpUgbkiIcLMM8+G4jotlvHldRj3z2KvgMXD33emv
LgSL+vYV03mDoEn68s/kjy/JBZUwjpFkKq4L71aNA+pwLqj4TViIdlNwZnmPo1zL9/kdYc5H0bZc
BxvdKJ9+gkev7m4VZQaWx4pEyDDOQzUjv0eGFMTJMow+gCq6bh8zEvqpfNOFelIV627zjEXIygf4
ObH/kSaTVax7wbpGbV+9tCmfsbvd92AvnN2C+Uzqvm0SWMNTVGHT+K2/IQG5OvLBjZRdm0SjFGER
0ASwoAC7qvROcW7aVQxC+qiVyTHNRj5DoqKd7pV+fpPgDlWODCKROgIeEnBOApYnUBZEW7goXgvv
kVtXAkyTOoqk1yRMD+wpaeqvsO4X04N3KGmnmxR70Ndvdkq67KvyZXmSsEVh5aCBF0BMeIMkIt+5
Mws6jmq1jvFSjoW5CAM3TlvLb/9tQMLEID/bKAFqTHtbT3nSAioOAMuB7+ZsARxbkgHw2PLwl0mJ
BRkrHxO50DeCZQFo0J9jtno5ukCyL9vrRW4NRP+lzQc2B7ijM2uSh/se+DSH+o728z8heLPxIPfv
ic4q+kazdhEh8iEk8FzYK4Tui4oMbcfxpk1b+n7x+eK2hP/PdOwwMzjFLz/SD62qCRq9LGKB7o5h
YdSMBI5Wq7j26dta0uEwzVQCoRAPLuWkc+KqLgWVi9+zmwSdfhfpbL89gKjkmPqYOrki3+70j26d
M+ItXuujYg+Dc3XSH9334TqOjBmkDbKnD+Fpbd/Q+ZOcvhMGyV60Hj8VeyqMC5kic+Lh/n1Jclrf
RGIipgD1ZpbzMSlTJuIs1//3/XcP59d3LDwbD44DEt/kE6OLm1u8qVwBpDY+Q7sabvOMN4tYTePs
rqZDBV4UDan6CE6gBO+yulxjfxNHWTIcPL4XzWeSU4OlOH31189PIb7vkDqMC0Y/SAHqvOzQ6aOI
ScKovQyvP1U4k08MEMRk+28EG8bmzEd+GYreyiETxadvilMVSbz7E7jhzgea20GECRGtMpjzRorL
cGSscsCWrM3Mft43UyXzBUOvU+wDBq/iNX1UdEg650bMrUmgiXbErDw3qCtLaCU3YA70f/s9nElW
zaZCfoi/7qmv7MxcuWK825AwnvUgjXL5tpJFgdMRNu5iM6caYx3BQLer4jnKRfRTw4pM4gOAGCzs
zMb8DfRXJqCi49OUOjxPwI06xfrzQ3xfRDHPnIo4JMjYkf4WQkpgzXD3Iyykb0u9gYl0CUU/9M5w
CdBD3heDHPF5I9HAB4s/XY5pZWkeHAQ7BNlY3cYpE8kkulCwmkCNL5x/0iBA2RNVxtzcLwExw2FV
XTWEvR5sz0NpMdm/vtzG1FgcdBq7D41lGHe78FlzqYxjV75F6zMKGNAXEgd6CmyvGiNcZezRunSa
EmtNdccKo3o5xLtmYdS1+7HNJLYymiFI4vRiXFOkYaEQhr7vtW/EEND0CCUy+Cli1yuY0TvLcPNz
26rVmFk3vNTeGkkEkJKPJ66/ILQL+C/h9ns9NR0Rwc9Xcw9JtZNnKY8IzpRqHZ7f5LeMmeblqKIE
Vrih7LO4yW3LMtUsl2OlyQh+EO2rfPx8dtm1n3j/Y1INbaARQoXiksOXBcfLP1AAXwgC2buSBmif
El263kwaJ18mat8+N4pulaIYumGy4Glw7R4XcGh3RJ5lspfQBocDCnNMGCQybD4x7STfT28Qbhoa
8t/0YDSLd8c2uIEUOy/Cml0I1WH6v+BePSrlJOuxHNYPTm4tA9NSgOvBfX28SAr1HDWStqIv+BSa
5NqWelqFUuDMLbq5amKDkTPsXR+ecu/UDlEh8w1hqO+DNVXQPJc8woLIbqVCJbFDPNlnfoa8JZHZ
UBNT8KKGXZAWX4hTFWKcIrQCiY/KjaiG5+4ply5HXC9YZBd3OZuXPcCaS9Tzqc4iXzk/JcI2zN6g
bEFZQX2KhPzav2k770X1oJX00HUF2dXkkSfRfEDSdm9fp00NTHyXwXzf/Ezziw9qmZ8LDt7aNX0G
pE5+F1tKSYPh8yxucemR5iTm6ooORtETi3opeuVI4OfifVsQOyI3SWgA+XwkhGV/EXUuo4KJyHa5
02e3TKosXJg6ek3tESR50xUY+r2tBMjCKmQtXCJlIJV49pxr+fdNEEnXRx7N8v2z8aOo1YU8sSqy
qqaceUx8II4jtCZw/43MBts/QcrP0ovPcS1EhgVKBj6zy4svtRBIydU8UeuKVMzCVvLW+GMPYvcc
gVUCTNIAFIkrQoqfTWJXZAtYZN/nt6ATZaqgZTYkW5S1KrMSkkTIMPONqgpX3Mqy3HB/gvYwYjnf
VHA1T+W8r961MbzNPSUVT2AnXD78l8BZp7kYOK3vfuEgtveqHJ5Qne8D7LsA58xquL6C4my/gaRJ
X5grw4aMEzaX/XCTms3wWnHTchyZF8+eulcmP4ChHTcb4/YfuUA5zS5l7OJTA41Yaz2C4QkB+SAj
nCi0YNGw1fiukxZo4EYsRea0J7BGosLmTksZ87HaqTmRpgj1jI34QBJty2KkA1NR4Ve2tRvk7m8w
qhZSstfUROy+FH7Q9D1T5BlE81wIbBg5mYvkSPHLCndhMQuCg7Uz7sVVc/r/J9rWnAGNHo0M+SHc
NH0WxlQruHE5LNPfQ/PCNgpLcdWJWkBD+RPTk1JifuL0pvpcCvgFPw0odoglbeMQns0yT/b4ozoQ
vs4bc2q2wNG6zsfR0QoVW/q7g+2PnUoa8pHLik3hw0+Q5OwCCjDDUYhhM/4GYeep9sNeFcCIO3HM
8hPIhSby2O04EAoSw4aRClbsXZcjoemst07cT1t43OKA8JqfNrtzg0v37hPjsQB6FrjAGSrsC7eu
/hG9m761qr23W0ddCZUwiBaGM1N9lXqb1Uv+zNtKfRR+ADP4z39eZV2EVoz4badFcxYUPnIojjCs
ACEmug9bKAEdako5OuLRo+wTA9fr6syd5+wGgOEP8MVrcsM13ySYWcxvMMYo7CpU6rzf7rqLNLJ4
dnzUz6UGhVXvbTZ70hjdjuh2zeWotkHVAjf3FfJGZWjJHtHFq3HQZj16IbDhv5i7egPraWIUv+50
+ilTRH+uB0MNWOmCPRnYqB08r7Xq6xSbzuDoloTqFoMRihku4i4Lh8cVFa84PunA1sk9xIlsjQMp
jkqXFf3uRcQEaZY9vPO4S/T4/G2BcKB/l5swbnHEswPSwBOVRvrN43pLKvOxPyRYFDyDG4YUJ+v+
7KYkshBwhOtyS2QkgfSVrUgFcebswM0hUj/uQ+S3CGer1Mk8xrTL4ZV6URyBRU3zJvuIDKnQwazQ
wnVHeGFFgG4kkTW9GnmQYnAZkGgdoPpk6lTrt/7GuKu5avpM+BivqTGz9GiLUzc+yNkmrRCD3Hcf
wiKJx8jKhRKbtqF2NspXYeoWJbqAwxK76euckAH3BACIh7vM6R+grN+x/Lvt7oaA7yADeOH12oGY
QMWWTu/4yYaxPyvUV34w5CoXncOpZrjXcoYgZGloSw4llThsCjw0wRrJUldTT8b+lPG42miXwHjW
NlDP6lKIeAxsFFTRfthrbiNyJQP7vpL341vNWbKwEdDfEN6b+sYJMHuelkCCshj/NBAJJ8J3tYvo
yLtrT3AqLQPPriwTG+LKF6F0xzKhVfi/bGFz+u55E6Xo3KoAfiJQiEeyWZPx8+KWdlLZA4h9Gy3s
sb00ygSZsE8MdutO484AjrazOZ8oBybwqNkIxKeCO5cwhkd5Ghq6cbIm4CXVWnwXnVfqOTDYSI4V
d9sgyzDRLeB1TBOwWgLh/nbsygRHNMmO0G/ak1lEWPl2TvxWQUobyBpVU9jkQ5DWx2BwVbhX+XKX
dLEeBzwGe+7E6rFp5d4zWxRcfG7mQeXfIwLqoOdlSMEqM1M+4DiDPndjlv9koWOZhqIy4hXI9mK/
8ozJP9Di596tkzwVrIuZWdixnqSZNAWzU5KLJ9dX8LN6SjSyqYXkp8C7GRtObR8/G/L2CCrYWWFl
IihBA9a38m++eyZ3zCS5+TddHB5cP5Gta4Oivlc/qmxrs4un/VSuMmPywAWceIsbStardo5LK8al
H0ZSahYeZXJ1GaOMDB3AHkoA/O5vC0QCm7ofYxwXbzJGFb/QkwaezovjNjJuGux/otuSQznZ9t4s
w3PTGn03iAW2zyN6Nkg5K2zzELIIjjlSgWI63dfPU3F5yAaYz2TQSJvaPYU6qadncxStSjxCH0OS
oH//oL3WlsAqgoF5wkt4MQki0XQ8QqUPcZCsQv2mP/WZclT1XBb3rxnL7ZJ3Gnh+PFAtYlmJlD7R
c9jUy/PFVvoVZe3aQ91oerP/Px5XU5Fj2y0g4CoIhOe8c9SlRGuLk7b0L6r8JvdJeTQrjhFPUwsT
6AopSIxCsZtaSUV2qt/xSASVq03ZsQwafmhcrPs9pr1BKeMkJAdV4Bc/xFPyqZnvO/svQlwsoeYl
8QJoNlloWrTqAEARTjL5tpnpDvSp7pFXbl2iXZLFBemyEl5dOFJFg6ij6Iy/YfPVjqFD5hAQSyO5
VKCoTHx+Z7fcrmLDCD9lbCrNLoz0dxla+dtnUq1qdYcO5r8MCOrKphOQQcIwwnMb91pej3d2ZAJS
gZUED3SZF6Uu3vftOaFaeonf6ZGdtKS83SIDQjiuKjYDapxegEAY27BddgXWhrXR7xsV5O+RrLhP
acE+YZeXTSMX6Z6bjGZ25/Gg1vFpBCJUKaF43E2Up/iUSeY8ogCH1YSamKhQkz3fYxhaSMZ33SO6
1lBIqbb9Oa4f2KQVTUjjaBVJMmgDh+cZWZzTZ95OHPqCcFVlqRmYtwwb4tcRQcrWisKwlc30tbQm
ic/Nl4bxWeb9BwMhozifS5mnwEqbqNps/PfyoT2UCsDSbDuHz8QkNBlpF5Vofqcq931Ka0L+TGCy
yKq2DV8nDwVBT/PEhyjBYD8CdEnHWj95lAlmucrsoEbfcoHdNv8zE47YOZe9rXPC8HUXIIcGtmj3
bCWI5iIUTObIV5SS7AnZ0Sah2Mu162rUHKgcmqCTYiruBEqvNf8i7jRgCFiL6nt0ev1OFPN9rEx2
3MAfY8i4O1hOgbMQNfw0lA0Ex43oRVQADYS/2p9b5FrwuU7n7VOp4tx7+ipdg+EXxt+Wusv3dRFg
cJ1ZSGvRorhbS7rv1vXtnJhnoWZSjQpQXWdKTOgX9QYJ6RlpM3tHh8XmwVopKH0yQc4wWAqFZBCW
4PIopVNJdjhpwhTt9emllgTUgii2MAr6wpdjV1iN5jSkl7MpVtjt3xc7HtCretUBkr3FWIcMj0NQ
rHBFkdeL/A352sAJu+5yToKMZMI05cKfUd2ezi58pygyMqISmECtJkCNuuPxJKAErfoVJFCFIh3z
0cutnzBae1s2S2lHWZhVrYyXQ7j+Y0e/Gc8nO0ZYJ8kA1UfTtNrbVPHRI0FQYWBJi4XbcDa+HHN1
jyocm9Af42yvXUULYToKbMHWA6gy57bIBeecEu7gW8K+TrB3spjsn2LfMaCRkApgZ8muB8xcV5Fz
2MyTrabHs3zzxVC57rBqA0oZ4hh1KwwirseoAzZJ7iZbn8LVfVg/3fFUM0jdVJNcPsvRreVq+8h6
d40qDDcGshoTWBPLWN776A3z6m6/TCIdAELjB8VK3zCvOACluKXuzAfJrVxo3cRqCi4cROmfviht
2A7AcBbwEF03vdIahBzNE5ylEQPvQL0FezwXKDhC3NilqQy/PueY+7Lgn580IJArZloODOtdLR7e
u/jzNjZvJkrwX2PRJb76y+cIwVc+bHaGbOF4+lcg5MTAwQim3oyplBPc4QOukeG5bx8WwXE9mKRK
K9KiFHgMCNamDKHh5tHsjhw3VqRzV55W1w++VxNuvYOqUOpYYj1O9N9ceS2/NRp70XJ6MCsWf56N
UzTzNm9hSbNN4QI4Z8GLv/W+gH9x9oxlg+JshVl0SdvVkmTED37lGoxQJpt9JPEubXGdONK0XEOl
n38Z1h3WYwDfLUY01ySCp2zTr7hMoYPm011ETEILATl/aa67nCgbQ1OsiLECtEg2qaggbjvhTl6U
jU7myIuZdDTy4V/peD8s5Zu0Yg5axx3ZcFTCf885fz/yvZWsiaDTPwzfyvB9i//FCYJdh1agdehb
OHyhTeGi+haThjtE2PiCXhHfBOEfSQiUa3W5yWBRg2ZIvAuB9GW0dGsFPpHcDw3zSSn8Cuws+dRH
g+mg1INEp6fEmND953I3yTiXWv4hk7pzkatfog+guTKmvONLlJkxDZGam8MOg5kj6SFvtFwbmRjc
D7uVE61R1FSTNFUnxpA6xGiqzNurHDyeBXmfpLaIvg3P5s/PjoNh3elu0EAiOsHsJQJydX94NWH3
yz8DpLDshfGw5ELFqLV8ga1jebBiUkSOpXWpkkdFUetAL858XQEIjpn61x2cyMHRxq1uksyPBbgx
A5hLy3luK9ebLyXTL1MHwRRXI5nxqNlzjmk8kZ0dMZdF0l6TPo0gTNhFlChgJtKjKlSkWvDDPxD9
dx/VmAjn1ovDI1FlUDx6EWYnnjJ3dC2AsaeOqQk2GcmXoa+KhTmS5wUx17dX7LV6hCPecSwx7278
p0RiGJCBopLEEA79ruAH7Y+tv7RXQuOsfGqDS9B0GTiirG+/Oc7fm1nmIxuKqS0esHwZSeGyKmD2
rLDsQSvkWZf0R2Hu27XPBNA199YU2Oee1r+1DIVcH7xm3q4LXf+YoRHFdm1R6P/mlCFOKtmnfQnx
OqWe871T5xlEQdp7k92IHy4h4G2WcpXpAdU0m4HPhOkBHuLz9WaGUju+QL0B8aw3pMrBIBnYN0ZZ
3I6KIWcVYwYL5SrkBm0KKZd2Pm5gpVvvhMdEbYMtTZVwTf7m1rx8nFbkQKOX9zzhYYySZyWTPz0I
iEW1EZeidmphEYD8c5cZk9rIQBXKmVjjkSA2IUaBq7cq5N6OVZ4b1UR8zGIx71hOzFBpLegQfwbh
W0xdQ90PszX+q8TutZqw2MjjAfjReQHe2F0kHQu7JViVRqXwHcAbRp5yR+bWqSxHL5DlcHqgVRQK
5gq9grWSRLNEUt13WWTAwdk4zEe+7fuZ6zQhZ6oF278oEdZYHBz+XWlKLjPNzSAQ+01/HsO0uutC
7MXxNG3V5oRkcPc3T3jtITnVI56k9WJUZRQBUO3es+/VnESMVDMWGXs56INx7OluKWCob4kYWiQS
1fyWCNOwI++Yqw5W6p6wrLnaIWP/rChYDTQXysaNPVkYEMBHYqXUZoh6bZrc/ilJx0cf4luZzCAw
Il3uOswyAR8NEnpvsu73ARVKqeUTe22qOJ3g+iKJQOO6PiFqCOpaQl4kNNQkKVM5YLdIPgtjlZpO
pdQPu4Ubyxn2zaaM06pIiVqoJdLAOuMnU7T1zL4NbJ05t+NhbIxoa9b4ubwtKvJuGdnypl9Qv+94
20H3hqVuUlIMqfnonUNaY+DC2p2Uc1xBgefrihLmjCsQos2Ml/iK/s9QbZflCaWUY3eoi6LyCX5o
udVS8as3Efduw92Swgrp4G5NRw0k3Iqw1DySQTPyCv89EbrblsE7I8M0zpfjHvH9s+TYDKNBCjBs
XkxdTiANvwo+EUx79b6KqbNpE0Crbs51ys/2DMQ4HjvJRfDc85nBRO5WsE9zps+b2m+XTT73oYAC
DA0FKIBCEeSJouosPUcF7N40tbhNZ4TYeWrmtwvwCa9C7N5R1Gf07EAd2+37dwg9S2FEro5qqPkq
s1tRScghk/HO1deSZLNDlibvCXhpxnbX995Ec/SC3LPqFuWFJf2986yFDG+GjSipY5SXyXIAFpWr
Gm6kUZy0lFcNfr/VWa66CDDk/QzZX81BuKD/bDSbsTXo0xDha+qQ/ubsh0Gia/z7oaDoBe0NaKLh
Qj0aY5EJu6IHoWQYL/H/tcvOFKfctLadflQyxQ0LHgQo3S3xYYLcxJvJZvzI5CoiXJAQPTJ2Ta9F
hwB+AQzCnS40Ur7Y6aoJgymvV7YQQudbp1JRhI8MnPDpag+NjzqIasbUsM3dRjW7IOxst9t/1WTC
K2q6gjMw13N303MHx9ISjw1OinKmj3LqkTIY6sBLWbETPtjf1UGyUu7wWHLdyQJOJATgDYJ25O2H
PPbPc/uD3XYCvEeVyL5Fov7bqcYnFj2mU3vD53EhVbCx00Uy0FmDHthZ/iLXZkpnohAdUEfs6B3l
Bk+zaKN22eEN2utvLwSgw3kSZZtXDpNguUHXsWFRyaJ1cTBVY5g4oWqX9ho7pihuKJLrLm+t4plu
yydPjYSkx7QQM8UGhT3FtIzQcVqFL+WxsS2RUWP1e//PZSlNRyH+1Ug5vIRwL1fT5/nBm6EEkJWc
+yoQy6J1Pc+Is0HiLrUJ6FEAdB2jy0gThqU8CZPjL3AUmRONG8OC+nAROPHSghjyZLccRQFZP4Ck
mwqv65zsJj8PeAYUemmKrpoVKsHzL4q8h9p1TFMHWtINaGMpmVSCJtNwsY34u2XGfuM7+i0IzjDO
HbBvBb/YxhYiG95uQYGoUXl1GKRLjuf8tq8X1ZwdzPiMPKJGVOPVIUifjwZKt/QQVPXVAA+9JxsJ
B834AiGIUZwESJ4sGzlkiDK8eI0/xFYHSFdrUjXEHq8DGshyRFuCNSXroQWN9kJ5sHpp/W2SEEOv
NX19BQSlBuY7KZdKjQqZCx3Qm5TgFuNS/BvwxUyZQfNVnCXJy0/8ayhPvc7M+eCApIIoEa6BaUvD
v9qbD2tyC/iR99aw8x8l8Di8WVG5ybyCSnnexWMPc3OfUPK2yFsmCHeNyAM4F4D883heU7ILX3JL
zyc3JPXB0Dc4MsLfydjHUl+WqPDic8K6X65d8zi/xYoOdAOBPj8pcKCU7NtK+LHkUcd8IM0BSUAl
KMboNHQvFyQouvADYBjDcaUh9gqFUcsyoF4qFnxD4VVD8BArHwFtGQm+yTDWviysG0hnW8aOxs58
QRf2rCmN/DyHmO4ge/YarbjfhQCMACbAC37W2Kve+oJX7MnWlbYqb+2y6Qk+sK3gLWoCJoV8KW/L
zZFeOfs2thhQ2CO/ROIkvPSvyZGEZ3BslxOEEf+PWsEEq/SW8EfSu4KyzQysYr6kVsFuvx+jTD3F
ERjLhze+O8p5P55LIP0SRaCjpZKAyJ9Eg9PPIx04gEIVvViGRx01YHfwGG945mK74RMrVAjUu9r1
8DiAGE3nGaFk7hPQXqpVJ+q9Ay6djuUpBtds40KHuVoSRiBWoqmjy5rMInMOSdF1BTvuvOp46YJK
ZMQwgm6Um7ZnWKzKw+2aBK+4ybnrtb0RxacLFA19GPDhppirB7I4MnCoSJzJsYTJD+myljAGO9km
Be5bpHcypRAvL44TLBp8AgqAwFNd2DCwcR7WHVmTBtjoERjFk8cMoxA1b4PPGB0BNtGAVJAMhZOc
wb+J4czC1LutH8K6RxG2nGkWTLAVd8paxXptBtlcmQ4kL8xOn9pXamKdfOHyGVYG+bEyujKZ3b6d
+MQl+AAjj49dSYR8/JeCLvrJDgmPRrXi2hbr30PxMmK497pt4Xec+mfgqa4byK+7cA4KtY0DQdzu
kSly3816NqeJIGGZ3QTxNi8CNShwajlJ7u+wFkeQgjr4n1RV17VHHe0RkYhOrGkBN8hOTdc/rZpC
TbzQfL34lHypKFk2Supw0jR8DvFbxg7OIpQuiw+Lw74FqThaW+Ug9SrevRX0Np/rTwY+yEfM/t8H
EWim86kX84OgEXCNqDM/gLfAFR465rVqwWYeFvBoTvPY5fpoEDuIyKALFvB/h1jaEEupnvZxFe/4
KAIgM8jC41gCdiqU2DW33+GIpNFjd2SphUg9ORvxaKAkftyRDGFn8DHAVHjhD3HN6fV9x/VYBBCG
jyFk7N57p3DfKUGNV3Yoib8+gi36dmu/n4YSxcnGG6bTT98W2LfHyruEI1+adUNYjYyvimHMWolz
PZAQRdl6BSeJihn52OgJFg+oj9sKb2oJt5x5xgQ55a0J6ZYZLomKyIu+nwRwvqHIRIBmdZO2lVdH
VL8nPockXuIw6yxn+ixDaH76PcDLj7dBJKcZKhOry3Al28PT4UUbdTDAA88U7kG+p2rpsTvYsTcl
Ny/r254ltraIk3J1q8JLY75aC99zflLPp0pHKfdtUvhej/iL217dRCUD+HYAF+KQEcsWlgj6xcbM
CIQXbm1ML9d067o3C7s1OUIE4VwagVkGlHo5I0Puc6MG8XDOFmB7+FMy+hattVHg2cFSz2LIbd/j
qcnc6DvOjuxpz+V29WyIMPoiapB8rBr/xyBkXn/HDoW+H0mHNuf7BtFm9++wWfraZQMvKb8J86ce
pjlYnVoTYOKHFNpZkTVdU7X/loUZ7W+IVidXQ9X+aN8FgkDRF20kd7w/x5jzHYYHHnw9S4sb1aFr
he3AHqwHhrwp1RcFjhVRHlUlsyTCS12HZPYo4225EB9xYZ8nZKkjSCEATPdkdJpYhelbbyKfGGOB
pBB+6viiMGH0LxcJWz8PK6P70Q9kcJqbzHRkuETG0FGPKRv8J3P1mGu0I4DBja+WqfKwSYhdyA1G
Pgra0tjvc+rh4tpV+ImFwQOC0osQZQIB+dfuX9985pYTXlxuMv+OS+55xxgARnTwzX2kza910wio
iHpldzscV4dHJhuCm/6IVo00x/yV1MsGq2kpDnw8/SU1YmkxFWOEel9sQ8JM0W9zRKijildcUfU9
YAtEDeY+lTYmNSj5lu450894GyMHzCeYa/m17akHl8/jsKmdv3l+U5HUES1QcYG2SbQ69Pt4ut5T
/EGwU9G7LlTB/orH8Alr5t3RuoXcTgliwJg8PFg3vPyatVRN9iDuPAu1YAU6ZcFRh+FghWqe9WsX
AhLW4RHxRJic8FnluEzeQ+X0N6M2d7dObkbRg5dgyIgXRCQe0/QAguyaipYoPkJYoWLBYQT4y531
ucV3DQeG5+R6VMBO8HWipoWjXWmePcLlIh+j7UMjrKZXsh+tvjcE+Qi12UMbXbNk0IJK0JHKG7ac
101ZxBcv0yEKu5sHE4ZIUTXzIQan1+PoredoXaZ56v68d/wBFAs3d8VpeHj7LAit0McXkTXYHYBa
UI1v4SvhJTTLWH1SFyCMPjy8BQl2x5qd9RC9wMi4akaQXh+Oqvr4eb4130tRHJEIseYvtCtpxkkI
AicKIoXItk4ZBVuvsWqY+pB6cEpm/UzbLkK7JZpJt3VaC+udThMIFaLPWm7gy0iBrSlDzYSfhrak
b+yHPII+r20F0G6CQSl5iNLPS17y2teG7vzTBL0YxLdJh5TIzOORMlrC51rGLmvpFC5ROsn58JzY
wADm+t8rw6pBsmN3oXjE03lSGMx4dh7oC+QeGKmBF/6J0sYmET7A1ITTlSpIDpgQfEBZIkUqLM4V
p2Oc9YK9x0YSUyBfVbKJlBTH4a+jS1HCgoAdlQF/3zigeWBeSiZ8OjY7/QK7nSaVh2+GuITeQksg
xVuh/Umffb/ZXdFNIpd5m+gSQEmLmPPPWV9pDER5BRVeNvhaEj2sIXhC+1cxjejODPvhMFDdqB4Z
WWqrasR3BNDQKhtMIfH/mfKRu/YZ91vy3GnIb9IIuyzuRvVdYLGAlsrsgAY/fPLa5H0bXh4M5eJe
vr5KfO/nuzXGWnji6WXit6xtelryyWeB51DhfU0fNFG7wBoQhu9nEcRCuTJhwn1PpkR3lWxnmyiG
tch7U2qQBibw2sgxbUjBsGBqb0rNV4fFN9jMouYYE0iFVFfpQAFctkRR/RtHsdszzi71peOF32t7
vENE81QlERnUPl99Eq5OKWn8Q70XRBIzXxubWTwuGwhswLm4XXjR8dZdr42imwktoSyEcoEBlgsv
LWBNBfwOlCD2CTfncDrWJ97WHvd9ZttdLEsQoNbdBjOfD4SWKx9B0To3N+rS4iu+cEq6EAE3M+5N
qqn3+8R7Fi93I7CL/eS9wz2/hB0C0Hw3nS5uBPhrscqmaLnwPub98k3r4ICJo9n5BzS6Kp5FeH8X
T+3MySR4cmonYDWHlnN+CLGPz/TsgfdNpHgCO+wYLRfsygGlf8SB63yyWFu4nk8brmaqz5l1pfEH
+YioNMMKX1/e4AbnRoh0KuQRGwWooqUL+m3xklD85zhmcQ3T3wwKoL0wceuvYjxx/EyCtQaAwK62
qTeO/dDxsoJisB3Ts4iSnL0r2yAyqC+/5fl6wbdOlGdur+Vod9hwI23cIfSDzDj6RU3DbAPVgQK8
KuXdj4VsUEsHBoNzbJCs2bA+a4oEbINPmRrgtMbnXIHyPw4VGVmxNUvkU70rt1DLLOTti+JzhS8l
hoEhw+etaKoaaBLI6fEtCotM+fWEcIGn0T31s7coGRuMeNufyC2spKKQF7tfN7fBdSF/Dva/gYsp
viZvFL+Sw8wcqxDlWq7yczEbpwQ/vhsYvBfq4reR7Jq8bKh5QB1SiPtaMiINdYi7jyMnU4Pv7mAd
YndfhpF/32fgh1uxo+w4STcKxoQ4nZ00aDPX8GR5LgEzEriXqxuEvGHP4wsFWINDgB/bo1woneo3
/ybFwMISfEalh60swi9oPe5gqE+w+Q8oURRfa2UJ0V+5Lroi4cjAB+Lu5tIPLGcjfOYEWvxoaOaT
q9O29VgEIFA+4bWwQ0cGtlzCIb/W6NhrtMG/lbGqVv80r7G70OBt9gId/4P6UnzeOKCnYK1bof1k
NVD5fvckIhcWSbAVjyAguyUXfqarsh3fW5PcEZaVd0KbO9l4KLzug/JBMaypGLBFcTkXVmXx13Dt
kiHZDVsDG9rRpMxrq0MxWoIBMVQaLM/JN9Wm0hYT99GQDNnEwzh09NnKuVrCD0ELiWkKTYDpymZS
Y/1Yjf2xfTUhQLZ2JXLSdStl7GL6uZY9CxMj9CAb3LqOENuFrLV5Y8UgEfT0KFUQtRZ8HNsiI6mX
6K+vHWCbolNO2NFIRqKLEIrs1UnKuc9d96Os9tHbPvNEEkEGoh0N7SPj1gGFPS7myToAwfxFpru3
fSOioUadaqk/GTgfqdHjEWx3V3arBnbiyOWH9Epum5/Q019cW7Vj4ZUHmhkvqMwOVKDnDiRm7Gml
HHSS1QWUX7ydyy+ySBWpy+4phBxobqNeezGfufcFBxEX8Jd5QH84DbnRO1JbfJn6KsDYjNqW7e5P
I+7Wgx6ONlzm/5PEjneRT3Ms/lUXtngLiBHJ/gjxdMu0x34kWQTm8FecODYPJXQKVe2xTGKpFLas
B6mVyc2mwKLWg9pcCKnsIGZhb253sR6miw/k5YNZu92GNMXHjCW3mKW/DPBOpHkIfghSQMLskU/x
bDt6jOGNwKg+ce9fJ0eG2qAIqlCp5RwVC9/xx8F9aPwrQqk98DNS4Yhz58hPxSihmsrXPYDQqXzL
bag52G9X2N4FEkGpeIeHj8ByqBI0NGz5hxkpWsKST1iK2uZL4rNuYup+4f0ivnjYYD2CEk/x+PYz
DRHkdOuCgn4vhORCbjXj5UENsRCTmX0T1nfp42oOzTtBHAkIOsXS8t5RCkvqMQIjmnw6XFOQuaWT
qZZksJS2qKc9zUVQVDQxrDhgkD2xV8T7G0qrYTjBMwT6v7Sqnq9UPBwSlD6vdJ/g0WDupmrNhofp
GJ+9Vl2+xV7qvLCeTpx5OlX8EniclY/xcAN4fOWHIf618flxtj5ZcYawedI7NT3dXMxj0S7JNOGF
TcXBiZGGBMGBaYC0nc99JFzIuIaAvwpw8ogFy6antP4EETLeqccjXv+VCdi3kSsqn5QRqLqwbbQz
ASLV5hp8Ef/sUbL5c6136XPCwXHgXDEjOQUiB9lYW+jqAfyogPk/ePkyD3LN4CF3gkKAZf+GNd9S
wt5SVMyNwWOYDr5ZAQgKd9Afbu/ZE5eYOKRvPVaxiXGMVVlI9/h6ULJYATsVUNHP9eKhBKuFglta
Cp/G51no5u5VsuSJTl9bSNPCLnZS/5KHX31HMVIQUuIqcNSxen7Yp1tMZ3LGuFQbkwE7ccI8K6B0
aGwshKtKPAKcQZSTgthVpW4ZUYbH2O+3XR47IjfLZmSN2wbJRR66uyNcHPmPDnq6PpJfQOTiwldC
YD/HTFnHPFkq90U1GixmbhtSwPYULo3ND0jbaj07nnMfQ+XxZNHLDHFJ+1puXK1US62aoWSjV5TE
yKnZz85OIiAAzqjulU8/MjzGWrz53F8rvoNZ/pbxcwXp/x2q9t7RqLuXbwLLv5ET68I+d3RZ5Jx2
Iy3xIJynKVgPXm/ao4rdlb7ovuKzIBOnu6Yl8EOZwm6R8Nn4d38BxS0T737jlcO2sk1zIzp20j7M
xDW2kqegGV0u414uA2+B6w9bKTk5qs6dD1HSHsmut5gc/mQfLAAeWNSKWYkQft3/Mnp7e3Tb3dpa
9YAeBYiIM6gcsfTiTi+zJr7F0+FIh9rqyXcC+rkZ0waHbzqkSRbOX3Jtp7Ch5pypD5oMRpHZet33
w8uqsDBIijog+wr9fNXgCJM1ajOZ856qwa3DHGP8B2fi2JUyDkeN8f/8G605yPE8wlXkJmkoQI8t
M3SrYYYZj7ZFsldVLZFbELVtMUIHRMuTpJy1/xUJMZw5+SfPFnGwuguXmzBtRSOcmnkTTGblSkZB
PGpzxw52Ez0KChEHGQpxzhPVPExfrOqWJlXUzc32ELpux7pG4woJPpagBuuOarGArHL8/vZmV/g3
9MARmm1N64q6cjEVTyq9PTk+olNWXJ7asUtYagFmvQj2UO6psordLwp0DYSVFd0T7vKHsc05vet1
YIn2lTP36W+e6DqqakzLOWgTVH8iKL0IxAttyq0L5WwKGT9lP6YutpsMPKMs1qJ+rGxQFqd5+MMV
nLsH0xVivzkbyQlhsB1KnCNfeeixwPBImNLd7Qb5HOV+t1jQDF673hTI00Vlfb1qMZxN4OlN2GvJ
Zvb/rlkz26cMdIJ0VT7PdlBDMpgxOF5bl6yVYdoaVSxg/8Pn6INvh4zHjA6ZipJ45ym0rvMKcn4M
AhemaILAaWpmD6LNZfQ3Nl7ShfRiS5yY5dqwOdPV6jtdvGEGjJz1sfIK4R293BgA7GQ0Lj4vKn6y
deZ5Ex7NPuIt0v2rNK59yE4nhc17sX1PMTWJABTLkYk0M/2Ac/Sdliraggs3c4KM5EmMdsBy+r+P
P5xT1ATEMH7dk6frd8P0sD0JPSqMhJZNVDXFoIeqnsA3+lxlLNnGyAwZr6+R8Pg4dX9oYnF4rHGX
hK5RTNjMwpfPNFYrZVDiSHIrIFg9lXvfLRPlgzR9jR0QzAescqP62fPnZE87n0Gg3eWH8bLdiapI
U9zI3agGyOBfdbHFRQt9MBSgm5/1eTbzcbWxo/LTAsf2rfjSfuEakzXGwvoPUBKABWjv3NPP4N93
BDvXQLVhKiSEK6otTeMjMmZR2AQJRJwxynkbcE0Iitu5SrIucvtlSthsUGO6yCXq1ylMVCQvzaYc
qNGlfkINNiLfHPL+XVipQ9Hj5JJgYt1nf92LW3rqlbBVrTRH9qeZ63eayypBYVfLARgDuOgZYOlh
WloVWqSsrKrC5g53+9BWQCLZ5fzTOGPkyvUgP7UpDD+HiNH8IcpBNctRMwkqwinr91NYjcCPDH9o
9Ew7uPxJfLRxDWDbrhiLIBabPjpXSoz+2iKvvznX7tFytrOnBdvVrQ8SbGR2lLnMmRIhba6lMT0y
ZIGJPjjwFeL8wsoMvl1psMYIsAY2d4JDVLPEf+JmMWGPJaRXPzVazJ47/+87M2B45uFGo5beWrto
CvNcynIrlHlEjlr/C4OCGdiVLC7QpmUKy0Q8bJIA2EP1xm+xPUp6o8nCYGwwuf+SmkKNVqqnaOEY
nzbHX6+NQXvF+DCAiSPpcrskcrvIz19kSVcjjF4diO2v3XEILBOC5xadXGw5T5KXjPeRy/ohTca9
ib2vXkihtcfnOgPcdFO7hJQ7B13DJGl/JV8Az/5CLmgKtt8muYNPa5aLCEBbKm+hSPTEXEXP0Yor
ZO89e5F1LAlxESWR5+ik6n6SHmuCKk9NTh9wDjaFIXPmjv45CCeuV4LaezRIIZI2wu0/dqMTE/uc
yaTjnO9liEuMrJRPHFP3wDSNq/IJo1Fvy0AnixygeD2cVIFW66omZgafK4yXh1/K8bHFXyZhglmX
nQiwoILxLtfSukHWgtuWL6h8eOmTmSRwWkeQaPa8cYrMMl/kdqWtqLTKy3yqPuXgPghCzNHRLfrS
mCq1ly3zKmpD6MJHpgMb3U8yt0shY8pJ1GlCKozKRhauRAzbRZwbJCnl2ofsQhH/x3oVeP1G74OL
tg0mmFhN/HfusBSZDmyVYLz159OWweUAKAqvSxvatesu+YHdaSYvo25+Jhx9t8GuFRVcBOcAy1Oj
dpRvkt7yMHsFio12ewHBZkzjJ5gXq7JrRb/2JJKRyeYrtGk/a9VAZQg6MYwdkGeklA94oyB7kqr7
o2ls6jT6BTosbAV9+yZw2wM38I3ZK8HFfyK/2g3dcdu7e67InCOeRP/huHRm1kF1tK5cp1/c1x75
bZYbGg7k3lcqHzwC8wPchIRZTjs4xghXHB7/6mQx6gsKgj/EtGzOAgJEbrGM05t03NJ0kP9b57hE
PaZHNzbhuQbw7MKkrEwtjkhfTQHqUy6kvee31s9T86gxQLRqkl930jzCxeJ+5YbPboDPkQbONOuu
AsDvj3RiFA1sI7Ctp09GcehdNpu1FhRq+4QRSeoVNdc1dOHS7ZR3lKUIyZ6hYtAC53my5FQup+wJ
PDkTIk7lXP/AbecOyrGNHD/7Cf3bDnsVvQpXELzV9f0Dv/aMGacvBhmnz6qEbYi+l2T8Q+1cIIEf
cK2HyWg7jiVO/BTzs9VbGO6WD9/l98psYEVn08FiY+IphbrqQ3DlatJqvqluS8SfcDv6N53fEZqa
RFYOrHColIuy8BhQEYeJ6hFPuNd3BXHmI6MZLfqRin5fyYRZKuZ57Do4gDXnOY8yP4/0DrKpIUul
yjoOp/r1mkCTnp4cdmhnrtTj9JhB+mTg/Sj1cEgTOZUtCz5T+vc1mGW4O4GTVk5A88RUaID9SWW9
9SZ4VvNnj3H3F+v061JIUU2w1T/Qm7iZ4P1R+xg5YB9RdZ6wrUKZ2Y4Cj+nL+er7507tE2jQAMkU
DKJWlnCC7CeIMx84tAoKR3MftLtX/4kOWklDQM+0OGrDSvNHn6doai9+kpVMtYb7/iYI7e7FTV7e
15TQ6QAcWnqrGrsVWNmZp0rxaHMbqPOw0sDZFoBHChZzjemv3hC3j2mQzS1fZHhuEgPp7D84Lkp9
pojTko/NPwTpJN3neuroZNRHbklbKBbtyir6S+uw1NdchGX+KqORVYEEmXrZtJ8KyyYsoW9qoT2Q
DN260Ek3U9E9DgaQ5/cNwg/jMIXJfk/miayUt71V8C4LXigCAS4ZjgysHHo/Q0P30Ck7qsUtpBlP
brS6S5kjTU4ABneuJGfpF63bKULdJiQiebtVtoMMP3+XfKPSGefy3FNcj5ez1SekoxNdK6ms2iRV
I9LOiqe2/sxGcimseQW6IbSycNHavufnvB8tK+fEgbGehfyBVK0gCOXYMCcyCMCOLp+UKb4GZhcc
brTHqnKlPIdckxcjts8DEm8iiU9nl7U/aVvuLAClOdnmn9Gl8ocy1bvvtNxMjULFCPtBBG9zhPLi
9EDdR0FH1CG70riBHOgCqYKz+YUcORz/dzmmztpA5BN2l2hm7rKpWceauvC9TPXQT40xwBZ27J8Y
VbL6fwVcznOab0nkkk26hmEsGS5/HbT8n6VOZm+tBIaO8uEeF6OOLuZmvhEO8Ados7ThPmIix+o+
H7LXKu2pfEq/RitmXO4w0QGMA1d0/tiPuS6v74WmY8WG9VLgSQbQjg2HEgkVX5J3NlbNrcIBBcPG
arhebvJAElRB31v4HztEGpVOOSoZ1iqLI4EoLiX/c18YoOKOUTLAABaGOXq6QL0Jj8HAflnN7zjU
vUF7ejnAJc2U5V2+xSry21KzQe+am8GNgBjiS4SCZiXOcYKXjYEWaiijUQpmDXrCSxYQBOhFW6LK
/UFHKYm1PeAe9x/WflrobaIM8GTR4zw7sWK761KJjgE5hvODiYoR8thxxw+bj7oYj9Phk4q+LAUD
Ym0TGE0gKzKxSGoH2Pgz5FqO1kHg+snxEMGUCqKiu/CWhqlDCCzNDg0TBjW1+EA3jRVl8pGIt8F+
gA1EoTEnVC74pxlkF49jJcQlBDXkhg56bRuqX/uA06bkytMjBzH39pwTB+bPJ96eWoq9Xzycx8GZ
gwTVxSg1PYGap8hEzklJeRYr7GqiFxkMSc5HHL6C9tnWXvVjM+fVThgupVk2ziDT/GK9ZoAJb8t8
ZF1q4muf6PCV+J1zsSZgw+H7+htKv3QNOyOlPytVLbcL0zibnfFZ1ZEWVEI1Gx8RgKQi/pXKtlix
QfxE40PNE7Yr5wzR5IVIRV2q75SXat2x/WI0ecetXUyfSF1WtrIl18Pj1uxz5WukjjTuJppNY/jE
JO8jToibSFk4Wldnm9AUQRWT8ohFTcLX9JdfjrNo/OQafct/gAD3zJk5Dc7XYB8TDjxamK4+fFTk
t5YLhcwZAsxuwcKWprUJ4jzamohyqyM1ADLaOYe8kGysVt8tp0k3by2Q5BkfVn963y3AaRw1Q96l
2d8L7T8OOdfmgNOBz5QISxyKOcHHMDXu62x/hxPTi+An/dIwl1pYnAwNWwQQCKerw+5VgNi2Ixok
GeIXEgeRu6kZ0ocQ7MUE2ksiBs8mDjAXF5BzvIqWtxmZmUHvV6aIvB3K1QQ0LfHgAXcHC01YVPFQ
mfI8Inp6ZSGhp94MlvCd/MxLCPnMp5ONlo4s1MmzcoGOaoiGjqBITDgpEU08Y2miOA1qfpqUtfng
kXANZWkd1snEHTUyIwpAvo+g5HiMdHWCNu/e287k2LAxovMgbWgb9JpqvQ/s6FjM4JQ5+PWnxSj1
UARMInOVWVG/SMNUyRPumS0z7Bj2UBUuDOwX/f6pmc1KRGS5sIHlt3jeasScj80jHZVSnKFfQteS
IMlcOR9fLkt9VPjOLKpH0cU81gNS+RgikFzfKe3k+LOx6mh9CNjd0FGeAFEYrOX+3ve6WuJEKzcG
xFJtbBZcbSUb2n9S2dkHQhg9hcms3QVuQJJQYQYNeqGhbawW8cZRoRXAeQRuAOxLLC+5Px1HPkL9
ewyFZbwlyvVNUyJogIYN4CK522/Bslcki4x+TW47ujrE3KlF27q/frz6pSspavq1KqyOoSMuqMGt
UJe+YDXAdg26c4esg3rt2m1HsfBGFubgL0fNQ/D3rlLTEECsgC4EmobU6JyEcKNbuFwyCxk7NEDl
j6HspJgR8Ukz7Ejf3h9RXCSN08PF3hTmzUFak+TIgYJlThMcbEEyHp3Qtg4vHYGa8mO7JaiCa9ti
tIWloM7LdjKdNwZ0LLbbK5sW0LG5R/AdwhgWDkH8ehHMIgTSRLzVjxMobeXzKhcgaX/I/tyDNzb1
f3JBriMBn+EeslVfNY3B4N/jM0CfdDUIBzj0OgqioWBAHMSz5dQ/kEHW8/G7iONr1oECPTdTPsDX
1mqCAhyE/WbZ38CA/ckC5Ktjjg4Q2XU4AZSUpW156p8Ihk+YsqvJf4aDCW9D4e7wzvTHv7UxcPWT
/ObuinnYCR6hXP8o+zf2bcyvkYIxVNMCM3hvfxD/kIakixov/fxnYOGAtfk86w2BDMNARsBoJLvt
td+NvGl9K6fHLK2TK2Jg/NBpBD0kX0Ot/LBcqhyA2s8cX4vVuL8MOYWik4biMjoEkwOUq/2/UHP/
DnnlhAzN+RqTLLZ/dZwAdm+oCtFaXxq+Ox2zqGBGrxeYGTDzZR3mgYAuQV8XeD6n08v5IRh0d+0F
1mdcsvLZA0FBYGaRivb8Bsw9o/ubFgF07a9Dz5oWfy8D6W+qWrXsP6SoiosBJCMGcKHFCXjxgrvk
4AcZWb05Aj8u5bJjAiD+9IX9XaUraokHfXRzUGdXuix76Q01AgjnG4RcvEkpdyXQ+pdT8Kko/mID
7GG/7CMBSEuV63ExTSoX5urcDqzVewsybYssWfVfw3QZcKktr7KuP/OB0oh9nB873j6aqm/raW/C
4CHDmFwsKU2l4cikOEV/8jdDnaH8uzWDHj180yGn2oiV7eF2jLZY13wt05JRCy+6XCMDABrkI3D6
iV/nwuwnDy9ugp5GWIE+DPsp32TLnZjuHodINyQbMERvE7eS0NclMcWsBLqkGean2cG+aFjyFg0u
PJAFgGqW+Rb3hSc+5lqmyBHT9QtXRr55dPf5t3Pz1j0QWGOLS5gJFjIBVLKwvB5i4usykR2L903V
uD4dyBx/F0PFnnwUfR9jeujXlQs/tDf8YbUh0wAIq9cRkCS4JDJnvnyR+nBbr9ZEVvN+M3DVzy0b
rh5ekBZCu3mSHaYipZSjHtUWpCjAwIe9jWdEnJRFDtios6uuzDYqvYZmQl7BWWVhhUqFIUfm0BpP
kziwUpt5BbqdZxkICZDF4rr5yAWNyCbwHup6MuRG0aNdrZNEtw9KdXOZEGPxSSByeScqqEJA7Frd
pTbPBpQhWr7N3IZdfSMMsOxTbAZK7A/bXLhSvuUt9JZcMLNrek0+LXEMU2bG1qs+6kEtWb5k5a3i
14AgRAvGSsRtnIAix1V37vvr+5Xh7+kZTf6hfNfXStcHUD8uJb5INPWiDvzx/BC5Pdld7xFdlOZA
tV/NyqIMP/zxX7QawFO7GQ57DBT0oFDTH3KRZAV7zj2FTs7TPCLOKjHhnX0acb5xFbslHj7QGzUt
gFnkcAyHM9j+PEQ1bmc0lahfZDUs3EB0z8r7drdJ51Qy4dsv01iRTzM+cwAzAJZnpuJPMcPbqq9q
VsrotNpX9U37lHbfdgtmwKzldCyapMaz/Yf+g0mF9fpnAqd316fs0UFJ/xlTDFAmanciyaTPAowM
Yfa1opm9KUQnpFVrI89uJ1At9YmI/Up+f9ak4z+wSHhQeKBnP1uszzQBM2NbsnnyGUfkIzziZpmf
unU5FXvuZ8ZHDh8zLmNNG4ymmxvFrBuqoZ5HnyCQitzsPdg4KPeLfYry2bPBsFx52ouE6rxPA5Z8
8/wn0ODeB1Za3HYc/xmIlDS0Y2atHeGq4nbKj0xoDMdNP9P6q2X94r/VD4ra/Zgz0uXLP6h5QY0/
50nMZwJsQcJQS1WQNzNaQqij9Ikyza0s2fhn/q3LGrqoLJCfAS+2jycH31d3dcU6qQyhlaksx07o
K/igEuAcYjN/iwi2CKXwfSM4OMl8JVKyQUz8lPzKEmmUJV/0wSpGtzq1JjxUgWnvyx7yYugs299O
WXofM9xhefg/2NBp1i4oJJL4/3XoYtwS0VzAQU1dycSoRXeG2AmcxZauWQrPLYm3boyKoK+RmN7n
jhSJfBxiv8RJHxiQbqGRXyj8KZ6lpzKbItkfMWdU8Q3dzsHYpSjSgYaCUOaHL84VPtO46KlGHDXU
dLfGRSNs5IbQdK9H9mLTpk3Rh0P/K+Jw91X8UvDp2cj0MFTjg6KEfC3BkUhMJQHcsWRLQOWVWsh+
yhquKpjHxordiqNI2wBVuYfT53lIqwTGT3+45uFiPlzP/9mIuSHpJJHe8X4yjnLJU2SezyQ6x0J3
jJ5ik7tAwS7XaZ82cf/Be6eESi9uJ+UMgTZnDp8ym83ahEFlFyqx5vS6ZsPCWsrqTvrcSd1dtqCp
h6eQ7Ee5iEfAn65ihvx1Pq+Te3YT50HN9mVsCvUrDyiBLw/e3AT7xOpmI9icpcn8MDcD1m62Uol1
51TiuK+HdsF5mqKlzLxfzBemplTDO9j1xatR/p3hcF0OaadIL4azTVnM7Wb3BuO/RUGxiw+55fdg
MEX5Q75E+gevRXjomMsdiGUBKNbkP+nutoT3khgHRNVUGuP3xw2OvltdBfVwnCS7ZBRDrl4iBAJx
e7tKMDgwzhw5te36PkDJZzmBjBKVS+Hjm7lyc2zW9wc2vOqATMvMBDkv4kKy9vgMq+kSoayeAR4I
4yliWFKVC2qAnuKZ70Y5FaBzZQC0aGct0+8eWrWi6YThhKz41rAFHjgibdhfceCd9k+y3kIp1Ux7
sV27kJvhcxBVa/1JXGL2f1PDzi7NONxASqeqNOSt9zSL+is+MDdS+aRoUk8ChO0B6goOXyBP895i
9xGSEnzbI+ItM1APVmuKPb8SjVcxg9WATZVbdnwj7YiL3jUD/FgaQpSVbH6vNU0Sj7rW0JvjR3pV
/HMLvFUtMqJ6NJbDA0qdJJlMVNWNJWxY88AJR0tO4A8WmTqfsuu5NAmvV53V7xwxn++gesJNTGVq
LpJHb4/kHzlYA0s9J9Yq0NVmoCXUdszv4UCpiu1eeK6ZOzz9I5BFAcQ6+x5p9A+LlGNBr90+8J4G
vNCkKqRyU8nyr6xjZ1sxlsZJpFgkbqAZlSHbDxTa7zWNeYzen5E+FMkZO4vVfZ2UaFdiHCRSJZjw
mIWkmdAfqW35oS2tklxGQJN3kw/Z4texpvf25jFHrqJeQyhHnWXnZNrLiMB3Z0AOZWm63kBnPRFz
T+DhhUgWRnwlOZ3qTCl+ytYKUD4jGtzJDNdwueOafaAmxOi+jb6eJN8/siMK7em4r9R6cDbrUsPf
Q98kIX7XM4FYLkvOWV2nu4Iiz373Q5iB7hJfbAXLGpDTSyPV8AFTG1BObAe9Y4084XU4VpIinBDH
gN8M3+oiHIT6LOoFyEnS7gvBv6NOZzEbnPQ52aup2/M+cZZ3qMz+nHqCF9Ow0bcKVDbsfgvqIhRD
Bmrpj8Xg56whGNviuOCumtlViT+uJnG4F39Xl29kV5QifaQnqugr2FJGipCQmun4xfQAHuOYDIPQ
zMELLV3kRLG/dbSur4bpKUTftoWq6npE3t7l1aq/ac3dbKExbO13P53uAYVRYls5NhCHHOt3DKYc
NHBHM7Xr06ARWXsGI8fAVllowI5Rk794EC7OlT7HxLbxl4nhKV5nAQB3EVqXU1tr/+nly+yLkOU9
nwXLqH+l70JPQkJqJNmppKGaHzc2cdnmetaBeapkqt345ybJx6Vyv1rGpkx8u6eseVrABmxVOrhf
TVE+IWaSTUD1QUxR3sRIwbkQQZHZt+Nal7R1xSl4B6KalWTmUpwCn1AqCr6VjywUIdEZ3d/d71TX
v0yvBCif4vsVYkODjYNF9TLYx3ZoSeq66Ncut66WeBjmtrpAxg1a9XydTWDfDHbEiz0/03KKRIxi
s7kAzp2JJCg+jawZ9j5gVQXIK6pjDdhNf8997i/DDlJc5TLk8/Cbuc5DisBgBpJDSYWISckpMHY3
7uAileHLv6zST4auofdMAcz5CO2pSZFRZCikMf85zBzkD6hSHvsdUslIbF6v/fD80nWl/JHi1ubx
gtLo4R+xRJaWL83yUJsPr/kHf5KSire9ysvUQIlESHCYWlpid/8+RtXK5/laBAGQ0wsY9tXVD8nI
d+zGdlNm4yaSqbJwOPLcz7URPu+anmqPcU8UTi06cMW6FQO9dgoylBvmm0018XKWHNGP/sQLHsr2
gKiYvPVQ8nCrFoGVR7eWXjqILytvXkKrresh3isAJP8oxLXZyOgnFDQjMo9n8OKZPCSqfPoqvdGJ
j/zGoCVLfDaxyQBkticKptE3wlDg7CQChyJDRNusQardyjlkmwtW4LsKbBa15snuKTPNusyKsATr
ETH7NFMn9vdVfaax8wbhRIdn+V1/YvvBg6qoNWTjt3iJsRh5WhrKlGwR1KnogHn1YM4skZmYVDnr
h3BAKkBigPQ4eQxxnHeJhH2HodDjESqLaqugUbIj3nPqCkMdwtvUYzCYyfHbSQRChluPQeTNCDYd
X1yfkMGt4dzkdaQYjjyYbWnWIbwZ6izkvsQdi/HWl+eVOFCz/kD13GYJ6RM0T9fqpgRxhTWRfsXu
aSUrIz7XPQbW+3j5Ls1RYW0xriyV3A8z8vDMVTMQ/myiFYWF1g114g3LEZ3ID+IDO5TwG2jwat2d
RqmAgr5DFxaUqtsVYXpbZjEuL8VtZbLLnxYVwrQtnFU1S8KI0QuVA7GapBHriFIg0oFAfDHgIEGj
i+UuvXACiISM2ZKpyVvP7ZTkFcZKeIWLUaP07rJuyj4/EijCUdmSf2PcuPADqRwTssylhP+peykr
80cSf2r2LCOwdyXvqODd2P1HtuEUyc0DjPS6y9kqspAF1XQxz/cQgxy4Wquq7frmbugvK1qZ/izv
awawIZFWXax2ZrEe5VA21seBAYi/Odz8eExDblJeYHA4sW4Z5kFCvVdQezVQcIm+35K0uBC8HCMk
6xXDsagrFCk5kMvgA3PLIGq1KzUoOhAJSLiOwvFVANDO715kCvli2SS4PBTS0rBjpOJOakLpq9Xy
KrSD7uQgLuRkYiaFcL43YUs7TCQHkS19CdIAXG84vAbydMWP4zfAMauJ3Pa1yQ4iWkcdKXrkhaf4
1UfNQINTRLE7cU0bnlwgLnnvt/CpXe1be4g4l5lAsEj+XYKpSEXPe7RBIt9AMZJMJGRwjpkXgXC8
ghXq/9dopzN+99E/HPONVSw+uj8MsEM0whvrB8tVbmtsxm5L1qA3snhoWFttWiGHubLMLRqaLWjA
BRp9NSQFCfNkp7hzrriJ5HWA8J0C0EqaWT6+Pq9/BNWa09V2zMES4VglGPYmlqx2zPAHqYKczmQ8
KVa9JPISLx/5DDScnE6ndbIqZCD7tV/WDAKYSNdkxhJ49GI7Yv2whllIj/otlHoXs3Mvt99AwoXz
eP4AECBjpNYaUUIYi1ukT4hAtygUUO6IfxWJnwPNN5KQ+/iugyCxdzSEzM9H7ezCsjNSNYvEZWny
ciQJNU7DbpM/RSHMw3PSpi4Q3LYBci947340TH12SM14D5LHXazWSoejnsF6D9wE2M5A+WH/3tru
dmSKAC/nv4xwgWOzv0PJ0Zm6MJSEVX/Xiu/rB2xmPYxlsc64wFhI+mAlfmaPkgoqLRscSWo6U4a0
ibcId9AmskyD1BuDkkU6H+SQus3nxlbkRORHzICkbxDV/Wr2VZsCGnlRiWfNaTubnCOfuJVqn2oU
ZCBQUEPkCoMeoTkb948bxANAKgvb9R7FtdLqQ21tu1hp3ZaSSPJJLeJB6dhGBGW6Hdx9vhJOSyP0
RaxmpEyiwixLOSBZwUCEpdSYewJYIxbMqwmCkUWgaF0QRNJgnbPLc/p1X0PZdJ7lAqSbtvC5isdh
WRQKHsCt0bjSN033gJFw2oKAsgy2MbO3GjxsTNNJ4Q+YKimPXpAlIy2dY7C/jFNREwVhs4+S9ZqW
jo9JzZefTikEUGlCkP6lKtlg32ufymemKu3NJ9vWNfWNGGUtGD34atiiBev4ejtGpfPxHk4ImjPh
RtthpL+zc7e11BWq/BtANCRJOYNjUQyDZIP37IQKEIthPlOCrkIQiu1WBJ1hUGnfhJj/5e2FSAwQ
1A6GJiJwnMLgc0kOF/zOnnbxxwV2MRs9PK3WVNOlpVJDLAJ79kvL+5e9Cfww3htaD5t8jePTKYjV
Tl+9XRR9YEkE+wrDYekzGZtQYstDc2K0Kdfk80TfyVLbwiAhJJQ7UqGYA0tMgaILLbev+WS+5hqT
U50R31Vi9aXMTdG6KJzz5RrI0Uv56Ig9L1IvXXAE4WWG+smgTo8SKnVqm3G25FPZ22J3ship5Anh
3rQQchoK8KSs3EftnF3G7i6YnlfiyfKt1Z9xtb0Y5LJMrAi0/az8/ukEdtrsgrmRqXxbXLjt4RaU
7kFc4XxiyLgHsiDw5WyTbhJnujK2QqQQgHpvBzTWdOtC9NubZAFM79L7bmYEgqtUwjmlWqO4KikE
VzAioMLlfb1Mba9br4rTK4nLHoNS1DAtbs3HNCEclNrWCHQITcXt/T9GTOxEs8okTUsgVMVGaaa8
XZ4mw2HSrBdEG6qYhe+Roz6/pv8zgjkTBQnF8htFpaw7oWyb075+wZdXL7s4Vtl8thXGTdKwEKFA
/hw51oDz5dd3TRBbWSvgOcMLvrFW722BZ9b6oivnJEdNu9eyrpOXXnBo/flrIIj/W5KAaF3DuP/C
MvsIKDb8Gi6FwG+QHGK88yV63WvHNwXW3hW6yYhOsfJyZUoFpKL+o/W8xSYDqC+Y/doiqo7MZ6MA
3VlOpR6BASBfrlBTXnn8vKl7Y6ABBExbIOGZndSYDfIdWFuPeMrcsIYdUU8ECXEClgaCwcdR1fDm
MjHF/z7wIEuSueAIM/1cr1bOfLxTvomgFmhd4Gt0E8On2EBCDhFrtqGL5WGCG2HASppx6+lym8h3
K3hx/9d813L+wsYPeM0Kcphsss+RX80MQA8se6Pt/wGxdUAxOEbhjZZ/u1MmQ3ijuM7wFRGSAivC
Zc0sDQitwS5hf/jzTrGSeksTYOv8lqhqXVFBWSJbl97/dK+E4+HTyoMcy+fUndhi72g3PS1HZGxQ
Jc19NtXoLNxxp8KzidU9xykPIyCYwUKNccicpFANDiwfkiZqLwAyRUmS7H1VJbIN0MViUiB0DOPm
0X9SV8jUhpsqHajVADXuXgPc5zwkl+NOTbu9zydzGzOmlJglx/36uJDgbyMZu4W9XypW+DsJUs3w
qknmuiWRoJ9a9lg5CBHT01Gjzvp5FdoOePD8TBn6kt8ItMN8Z6JuMv0oAxELgFkIxQ85/vlfaSrN
JDaXHkxvouFcTd9k34S/2KgdDx3WUojmewndEnFViKVkav+20/goY9PTHZhO7m8IJ30o281SFxfx
n12iiB5K6fLiSQAEgEC0lSsF5QfKr2UNjkLs29UlWNSlh3Uo6qvp08EoEZy+sEEtexL2oqa9aeJq
lCx53UXWeHoq4ibVLV1BbzuzdCic0qupRC/JiBsF3Io7lwux8OnsMWzLAD8c5jD9ySF3+f02wR3j
9OarFC4+Vg3Hbp2asdnVK/OPwGeWLqfpjqKpMliMjXqN079a0Faf2zBCSA7HhRGHGYJUnCGfiS6X
YfK20BSsVhoMyRZnezoBJYIgiC4E8DBunf107TYfRmSk4/cEJX0bmsMVZHFLEYRsM7r4cd3O/TTu
4yldZBGz5229j9ghCBEl5+jbzdFQXI+4vSXJrrdo+B5tplGcRAQNjeBCXTIZdtiYHq7oqg8N2YMQ
hybxZokmjTUMGD20yO/EAb0I3Dou2/yIKKiORNIolxjBaV1C+QC1UE59kxZYDSkrjobuQSd/wj/G
Pni/v3UD+xEAz1ULPfEhVmQKfd9Hc/SsExIRvcXV6Pn5A3Q8F8NlaLjQbhODlep0wAx41ZaW9ihZ
WhqB8umeuX/oJBIwafGwub53QYhmaNW9Yf8vu/vRXOata+FcWNip/LhRjYHqZPe5WihS/r5iZAvY
PLdOtHGLtZLGe+zJq95y0g5wh5TTP12Nxnl81X5SPVm2TFeumyKBry9sDUtkSchnnmVyjLXdMlak
t0NfVzXso31TMslXqdhxM3HjALXFyDdN87SNrAPwvxuqvwbIZErT0Au3nOK0IP/Ycg2tfXMxpQk/
ICC3ofDgEcUaikdWjU4rWtqyz8kMUli6Ta8I9ujqT9A7ro5yY9aDK2O/eUj3w1J93Kyq4o3uK622
0FGgdpKoHnrjYb7s/AmBdyVWfjSH8lKxgRtC0D3TgLDvvLTQH1/AarNCVMtrbnRtBCvGGjfolHjR
IdueVMSI1G4L0CfHdeAXMB6CkCuK2VGoVelXPN0ZnZ/1JlUWe+DbGTL5gD1prUlnoj0SlbvWYd89
+hAMUV4tm/dh+SsXJC+z+tUQuKkmzB0k/bhtBtptVaQvPyblPyEUZfjhrEgtv+J4ukWi43p4AqVl
PeE6jeBeRhJ51nNaQhhvsBD3NbRgd6g3+G4JJHKa/dKkoSlJKDZUPGt6+5J0QEXmhO97n/DLYH/d
m/rB7syLcZr87GmeF07BoBZBuCK3NpQXg7iVn2dZ8oOJoKMRyWv2WSZNu/UdigKAmanSkvemoHsf
1bkVoSGyruvULpOz3LQvFsgh5qt8ini3To3uZ9Pi8vWpgzvZlQbmKlkFHY4ZEsHJDW3FsqE+OUdL
26+1Wn9P1u8Sw0kTMejpco5qvsS9tLht54SxMCsjXuTf6y2mRYr/iTTe0AyfHRWplgKu0JLzrY4Q
msHlc5lPz8mDa02rIU78YqefF2xhhhje4Z+ifsu0V7WibpjrhyA3V55dwAKd9SOqHmaOJIVH2kzW
Y7+ADXuCnAF8VT3I8myLoxPawHpJkVAQqc4IAMttBPBHldidap3kFuce5rvhJvdXKmt2E2gx536w
ayE24vrj3brkCdRWJ3R3s4/P/NmLaf/wRcqjP7R3A5vYwDqYdFTjnawbEd29xwBJRckyd0TcGvkq
nIAwovIPIQ17Qk5bRB5cI7ttF/ktUiqvSocmFe7/hP/K+Me/E9bmPadUSprCmdNAm4/cNo3xZv+p
P8+91utIHet4Ebxa4tlZHssPsBelCl/PjKPYRtJEZ0pogSE0B2CUv4mHRPFpifGaoiYgrbVuhuuf
2m6fh9I5eT7YvdWmbCHl4o5h+lax9uuWIIhCX4BHlOLY2mMOTigM52qGw5JXEhuvBGnY+WGRhwkH
L0czJlYYmHqqazdzUQwNhUgkfhXengk9sTuSvBvcJXV4lL0ocrQt4OB5EcERXshk/vitLAq5/I61
DVBTLOo1i0DY5IKswjmuadAE3IQE0J8cuejUX01vAXND8ssU2p30GQhZrvWYjQmnnqYGgFKqh+XG
UIhDy0GiN4EZM+CpXYIzqEEgwuWSShiit5nNdzK4o+bo06Mqxh/LAL8OWedNF1S4RDAuxHk+b07s
AeEp/dPJbRYP7mDu0RLnrKAbxyh+PyIHyNdX94ByrOfALQ5iQLkuac5Ch90tE/iC13b4PexA7kot
RSYPSBfJLu/cBKZYhnYaOyA//764us2oxd+KNJfUhgXY+XFbAdz2aoiaxmHQQMsbcp4IKrrq2byA
d/4ZNFdiaGJFrwWjHvLYeSjW5+s/RhtvozGRL7gjHZwwInYBofd0dWwKCbt5izGqfV7TXz1ayl4p
Bj24x6/hRkN6OsNdbxsYhNO+B0NU+7NQhPcap1V7GoC3+CuiEvnuwbBIa+nsxNCeH5hhVW5P8Zy2
oXrR7/ekmQE5fRdTnaM9jIXK+Fc5lzi0+rATRrBrf+TYLjOTr5wlfFIvl/W2LpQZ/XRdQXMkwraA
hTJU+wBstax6tOekf4bZFUukp06QqoUtEAW/SvpKLRdknBSYITnMdosFFLMacOnYcrxwA3hUL+qF
8z/iPC1VDAvpMJ/ZPPrKwdv0kJM5Em6eEvWawAm6rCKY6OcAV46y3c7jlzo1uI7dScIhiI0LjS0/
z0k96HXkVtXCaLvFlr6ACx1QWn4Chmk6JWxKlyrrwdgCrGY57QWm9hDu3mgrbRZVngwkMoMCdNjc
c4EyWQFxzEJ89LAVQ8+yTy3N3TF9bunHtbX8lqiYkneeKh+0am6TsIDGfHt6aZm5k9RalvnbhvFR
N7fmB1XBLPK5t9zivaWmlMeyLa+6hRXKwYy3xTc9opU7retf/TiPYWO/qvdIEnucg+9Lc+HLpEiE
GWmx0XEvbDDUgFamReu0MsFjMFUPTfA/cxRcKh55+gZoTR6NCdQQlu47t0MRngnTxUy0YXngoNoO
77Oe2OMIbBiJPh89LC0fGrr4eKx79tigwNuyCHmhOW+JDAzr+TttVkPc333Ceda/mmImj5EuU0GV
Uc4iU6vAHowR4u437eyUnLl9dTUz0atpinXZArJJ5uuYmUO00atyOO/1knLCOaSCMy4bDTqkvNFp
+APQ+9tr4YqyrhDlyWlRbJT92FbJkTwpy6BibM4Qk0cJe9GYYMG7MFWbZTl2jP7gGoBjUgg+50Go
EJcc8SJsrZtcS+rSb7VCjOhvYXq/rqOHzFesCkw4s29vVkjF3iMxUjIShqlgeaD8JvisOan4L+m4
pY8FRK4x7X30AFrKpAHbAhFa2u5+UsTtkFMVlehjr++EQ6/RLORbf3osh5DepvhwZjHpUr2OA+dJ
e9x18jUPXgkZlPIqHXhx/unEl+iu3+/rvd203nXLnU2hjREvjaUXJKQsIuwD1jSKpkrsHm/8o0eQ
NE6cyMxEV2h8BORVfzNZQiaFH7d2DQa+dVjUwn9FrSljjVs5SOrWj0h2OURT6NsfMAZ3bBJlzmrv
XC4XyqxUfv8M9AR6h21Qcq5p0aWVuU/rN9ngo/nRDVSYkHfNHi0cXfpqIAXaEVfWeTobukS1/ii0
cA1OrKi2F8oDhlrcSLnNtT2w2GO6lBqBWhtfYIsQwMHx+Yeqxx+/7hNgCsK25PEqMeEbOG4JYZ4l
l/J9wrrFwegZPYyRr2GLPxVomNAdawPvrGN3sCBJw1h+94o6TIz8O+svHbGY1GUgrXnqLQ6bSZ51
8sxlFAk+TWkc37gP+qJwssDoJXpkVtdJ7lCozoLfgoDUXktIp/0zka221S0QWIrGNDb5Kj9oZG0X
0zMfuadQvFGj3SxqLiObK77XhvCvdyW0keyKKmYoYtb/eMYFC9TUTh6g76D9X8Lp4Ot76MsgIMZG
SyqM9tgmZCMBdB6lYpv5hVCGB2SG+m+ZzkWzfQbVd3iUxJ7g9NGEzY/ItKVqS7EtklaMLfSjvVuj
bzVXKTANt78Pbra6tOaWC3z7iGnVz/mJtHHfSG+o3fYwm+2+KR8683X5GfnEAajFzVPp5C29XYp9
NVsrldFoXtE1u/cCHu40yviFy+WBlo2Md+4cVz9hzGhdBZU2oqMgzq5xBdufG4HsXfc0YHZAqe/L
jFkW7XQT2UaRuu9q7wa5/Tmvwy9gd8S6k4asf59YkyDaNWq6XgpoMENWNUVICGcCQBj7BRFsVK0o
ejyQvEryxN3iBTlrYIPoIkliVwVUljLLxiKRbD/I7gt0RAFWnd1u5mw+7EZiGG+X8RN15AENTxHz
R4D7qmskj0BJZvlYu7jwIKLSbjlUBaOAZa92vb+9PmfPPw2459z+nqqWnp8bnqpVuLNM2p8Ripdc
pfm4uhxwvS8rH6DJpnJ3zMxKZk1bpQ//OisZJv66lMTh8+qPYO6FLF0bLOaPKklmxvPl1F9aTpUJ
WAS5yhFCLYxfKUDXrxPddIsFgphuZldztQj+rDtjDANltfXGoJJOtkhqy6pdsvR/OvwX9pCrxO+e
zh+5J7DrnmIm8qZ2z2VD2HTMZQK5+u30TuXhx7FXFsI1/Nimsq14C98khSetajWGCRXNzJ2PcSAi
ee+1cLu4VS7U3Jn2FA4EVsaRnGSpHE79ble4xVheJ0t4SjdgOAb5nrTUNwCaYnrdJaaxGqIu+MH7
REuyYl9nAGyz4zLughG8yxW1/oB0ejhbjZMRFtmos0+Ry//oO5md8ntvn5Y6LiYWQj8iM68Sa8Dn
Q9awgn+GAtO/FMtFAfds0ytOYB5L+PLXN/fMSoagqMVo/dqjNLjSx0/nwouJtxnetvQjPw6f/NDw
Ov0bJEWGI3xP//L30MMAXX2fZMU7LA5N4jnUFuCiCrUMP4L1TuAGl/0FjPp11Vbgf20BSTGjVFy6
uHLKPymfqJP8sVVj3kskyb+fM0hxkR52i1qwksdpeX5GYh6rTTvEIIG1hQ+v7+zcp/yG+ZfhZP37
Aq9AwF9QAIadv/Ihgs7Y+SA0LFpU8Zx/r66IJhTZakuHgdDcyFE3Ymt5sbfn/ZC1znd4OsEk1j3D
ZSYBM7aR1x2l/A2/qiPcv7HK5gW6G9VKDUGlY1cexR24oIFAvs3qI5tZe6mL8SGbyjrYfEEtgipI
0GXqG6unlMooxH+3EVTDZIxMkChZM3qjH8QwT/PSj8YtjjBSnxBcn/WdBZWlariQwvcDSwVeU/Bw
llNfXdjRn/u66i3E0QgXD9JuqXmt2o6aR0/BpHE8MHVCkfnlnWZQMNRiVUoZRF4hfYMMH7ByBoRn
VnO69MDwlYZN7VTGccFLnXpR0l7INb5a3TGVaGXDz1J8QltSalN0J4ic+sXz3xdR+KxSEkcmct+U
wuPZ7J2assnQTzXM0+iuIFXRtaHrF4fBfP+h2iLuem9wwyrQRl+kTZ6+VSpAmdsqGwcoYjC3z4pt
J9c35lZ7rzd8dATdTKgDUsReO7q5qokRnf3s+/89WNXokLEzqA1LIZTeX9nNJk/FJE9aOcjlGwPW
GutOZine1CLuuU1rmZ2KM5xX56PPaofwzpZTEEh8E10RZ+LKJRMJSd2NNHG/vkIxsq/KbQ2L1hay
7Zt+VoqKUcvwgDVuImBBiiTrG/Lu9RPIDpQZAKJWl3s+Kx+GJeiPN9drdoZKuaVtz0S4VZqfoPMi
+GAdIkkz45UCN+9q93ES38ZMlk4DpmQKIRDAeFa19gpHnx61vmoiXEiIVc3B5pL6kIgPUYAWFTLX
2XMYiYi9vAf3r2cP+OC8Cpuuivl4CiYOKhyFChE2sVHMIDEIyvvMKLwKZ2TiNIsJU3LUMPcTJ+IR
12qMxj539py9R6weUwRTLy6k8p/RdfNV0GiBxFpOP6qvyY/WfOalgqaT4J9qDiVSFCiAlXwDv+Nb
cVljOIbAXQe++rnWEDSvcanrkgPPiDTHKIDHY9rxPwj4ieY4MUg89FrSRNUYwtTSxFfL5boFZUn3
F8oA6ET14quaqF1WPNLH5bpalvhO/Ybi4WSI8fEsTmIBhIHMN4yx7I5t47ieKmjjg2zzc/hJt5d4
3OQUfce2UFj7aeUkn83izS9XTcNodMG++pc5XKGU1vCWImDd+W5vqGfraPk5VEf0kDQUlcRnZJdp
r1o9sTJpur/wGnGwEIlUe/Mb6yVg+iNjd8NyI9lapMdnUAMtClr8CQHoUmSuoj/3Klx21cZbgp1J
kamqZxOrnxP/MX4Fy5PDLzTc+td/S0vDPOqZ919JfTaYOZMgQa0wrUdifg9tpfC1tZzSTZpCLy5O
rvvlPYIiR1rVGgDSYG+Pb57pgBUWRjGWnLn394UHGZwG/qy8Nt6R/NtAVvcCVufU74OubgGWZdgE
200rWpUHUq7DHA19RmSG6NEQ94XvE7/YgO2cep50JYr7NVXNMD0a5h+NUAXEn/nASEVoFOSGzqjo
FJMjS4ypsLKnFpT0GiiZeHyZMEBAFQaZDsk+8MKMo+GaEHYHLbyLzVaqZf0WmawGuM6IhU3rZr+U
DsGHGS1fpWEn1N3tiLu+3jT015ebIi4o0y0E0LXxqx6Ow1pYgZo16pUtQIBSadudt5dGF0O7dACx
MCb6hg+27jWZh4AKJ8iVj8kWESVM/QRbjuOwOgyjkf9rH7Wcxt6bDPVZJ6Vst256O7ND0pfxcglj
Pn4ChP5h9B/bnp9tauOhHOgw/QqjNHGfac2JlytG4bUK+ewYmIEtxG7c3ZVIbx4L3ETVnktxSWPO
rO/+DF9W+kk8IXVZQCkVgw1KblXTeE2CWAccm3ENXECUggXkA1FaUd4MnME50Wv/FsSUFHwc0P3I
peFqzuEGjb0szs1wwkjlXlwJhyR7ekQ32QCp2kX94nS1RseGzBakpcDxt4KJZ6DyfozRTGtgLztn
ffRPEcynu3jbDYKDGdN0wogMZYTepCQsxffjMG3o2vjmqftCZopUqBV1T9v9Gf8OVsRCDP74i8QH
VFpZ/G5XjhHqCxJl2gsjJda0sdsiec37CTh6Un1qQjInC+qIkIfhLnB0ltGYAWha/UPXko061wbT
Q8RWdY0vROVzogsZF94E/H3MJOotBMzMFrMlpUp2GkRemXzt1/5ChjtrmV/I/541JdeB7LAaKce0
KLZqFY5gBupvqEVopQl9oUs9HpnNkevnGToFxgIZfXNayTsckQj/qe51kzb+QOM0R6zpIA+POF/n
z1mLT29WWqLsb7jJaBvsDCdPslW8kjnKKduT1m9qymaarD2/OTU9MYjRCzG/GljAPjvQyl3N8j7X
8+vTrBJ/4qoq4aTejsVHiZKqavSVRJQQ1bUrFOa1fGLA533d64nv2WFwAXQocQAtYlROcgUkdrsW
vcRQY5Kl5wKWXnKbBVBcCJwyj01w7G8rtKPWkJkHn0P4Zz2Q+8zeWD0/kgefwKqsc/XH2FePAu3L
+tA0Gz5QflqhuXikCIFCIcfmOZSaIhjJkUIaED6PlUbT7BJfDAVel7jtAePGrkJbtPr3qzAZ4iNR
rvhnKV3di7Jdzlwepa4JpDYVr61OwfzPjLhmxVrHUgp++p/d0mzYH1asrOek2DQgmufjo4n0ssxa
PRoOGfodUN4gy8nCpbZLJw5yBotSfa5JCM+iJr4U+s/5AdhrZFF9/x/lHVra0uC5oeZ3sgtCIwKN
GfSxtoNKrprmim4KbgYJy+lZ2wALLS1PHkrBPYvqXpfPrxbtv9lvwGUDXI47B2kMY0pUJ/bu9fAk
XOfGfT3Le81VIK/+NCHsPVhOtwPTJYAS0iWb5nlqzaWmukRIi3g+V4/Y6m/A6MIg/enCqfWdjBbI
v5w1bvI9/f2CiQGeMLsz04UiCBn2hdPmaRdiSskjImRz0zKjZgoym4tBdFo6BV4s/v+D81IslKzH
ubVqT+W5Sc8xy1vxsZO2g9Yq7tIc2kl2ttlb6THRvVMkmIpgc8zrgxXpgRiXLKrzC/kw6W4ikbmu
jQhypNWTbxkm98Wo246W0OF2rwWgArX8p7O0DXCRO5UISFpiPflcR2uPsiVt8w2IiYsmms/eN3K2
027CZvW0aPnkCr9u6ipUpF8+PjUin6RpwTsKOZ8+qp7ZvJuKksnpAzE8YRhtoh8UoKLjCTTaJLOV
19NCgh1W+hw7EizCXuQ/Ji62oaqi9rlU+EedooaDMqWBcEoiBrn8/S9Px+Gjh4jeAHkp3tw4IJBQ
dcfRq8yNkxXvjoqj2ktZBarO/tJhNaZ1NKFJSXZ7NBgWB5ZjSZ1kzNcO0Ms+/UXaytjjnv0AVGEa
zkhW2uGBjWJy8SxwYRm5TlAR4w3KEc2luU7CQz4Zg83sZmGsf+tzH6fDpah3nSIhEzCwhwwuFzUi
HOfOd7I/jrB4xWSCUhU+HKQp+Vj/6BfJ3dn7i0eBFK/lPOT5KzGIm7ESicm/jlAtk0KU2/EHOlcW
QEAbd8sxi1xbD1udQi3nQTCvUsfD7Jty9rYOE39ai0t1oO+vbtKWdEOqClYST21igGcq9mTYBzAc
lsZ/L/Slr5ERyJbruLkPq9NSStidpl0CyWNdS1v8k8kpSQ4xrAd9PRybZwaxCh9M/p8gl8qU+ySu
1Pti9Gls3lJ4365qTJ8g2lEPiq3iQ+D4TbixhtKBuGoGppbayizFQ6IyJvyuanM3w2Plx8MzXHtY
2ZnRLbFqbfmbx7EoS+0u82EER8ETwP8jJ8si4NqfMqx7VGalNSjC4+AHGZ5xKYAp6cN7LyhpFqjF
Navfq8tJo1ULH5uXQNEx1ANb0OOFy5Vwe9t4/t9fyFeCDXWdKHmSJAcJqxGR070JF21ALLMwh2E7
2dr3W9mGdU0tTGUl1m8faIXTZBi7e+zkJmUWHoHJrc7UTeKocUOoLBh69VhSm7ntO36JP8zoL3GQ
2Te8erFJoly51pvDE0l23ngf9OSY4YJ9wep7boNdpEtQubzUpDKMv1mHS70i1eTtMFYVipcD76KN
EVB4MM0+JjqQ2Fx5qGiAnqhDv4P/0aPhFsqQacTlbTDpNfR4D1b7BBOUXNS+eoM0VdUeehT22qBd
joL/3BK0aRWC4o+hqQlNKRY1oTKDDgMgo4DgNR0gWoBSa8MTJ6tX8nno3VD/YZ4CQ5iZ7PNWYp7n
R2wC/0IrxYx/fDg/vvx/hlKuFr8B3o8K1N4Hutqy2Pe4DAiQ5yH1pVXORgeQI0oIq88nY0VmEGz8
QTThl0I7NQ0ryAwldTNQjll5on39kUYsZdI1x2MT3Aw5Rf9C4/OLn6vhaouqOnZXryx8oHdnRGOZ
RBisQ13oRelp2NAZrXE3meTvxbw6MQjGWp0B6g7GzrE6sXt9YAamOt7XmJ51bXGIvf/zUuV7kVg1
xytKh1YpARP6Ptwna4kGidns9WYh+8IPl93C09aJDrFy+iOp02VPdBOjNVJddojcgDwNPca9hzF3
ya9Yz38eZ1+m3Nn9YMZZ1NJ/PcsWsEMw03cxhbCn8c8cC5KMRVuZ3HnqqjjM6JXOsyrO4HnZVwOe
q9XCvL4PMc8ckuGORH06pyDq1N+NXqbETcjkX7JyvwdRZlJV9tOHUvLxwebsSYBU+rDOfY1slo8O
WWV18ra8VkLlgfo7bNGAQJlu9ehZcRt5JVtqbTUFO5nzRo817qwHRkY0XjKGITpcJhGYukzFBC7y
dwEDSZAzMqOAq/f1gAtdFu8nQz+q2A5CaV2C5cGOQMUhlrMdczgwCLZnky4x744p20wjyW7gwrU+
1bdJCtXUOAPArxbLCFn83JjOdQImLeAYSzV775+2Zos8gWiH4pLV691hX8hHgIqy/CyrZls+ZO/K
Tldh72w0xT9L4CMrNSY3mFAXL/z2gtj/PYJtMs1ZgmuHeZM4fntK0JHawKUiuhb0P9O7LBnPaOba
Vwo3fT3GD7Pq/b/Da1yaJBfN85eqVaS7NgmDgn0J9OPaakhIDUt4uagMsERt8Hhr3NyGdVIVDCVx
oBx7zkr+zVFi/b5qWCB3AMvOgwdpvveqpkEyRyMhSDOiGEash01Pt/EjZohmnzyCPefKd7MevRsa
8SDL2nwox0acRcYT+9n59CjoxVTUl3Q8xRogE1DbpQX/KR8+2zim7pbmiDk7zM3KHIQEEvJlr9fM
ChCGhI1Tm/nuXjeMBQ9fjtr6pYuMHsT9PgK0FB+2KmfqNZJfu9EH87OjA456SdZmrT+o3WTai0cJ
RZzizo2VAxL5/+ijyf+4C9D7K891xEqwhBxtOcv5aF+4MQSKuqHWMJmW/+V4APJeBt4ElAm7zwnF
e8vlN87jp1S2Q7QokDNlE3MY4GG+JzKi3gCDqNZyR3debyP2Ut4Xab6APb847V/UAxNEB8EcNtyb
KmPinGkGtMdYzb4ssbMPU70++yi0PD1bTdQUlSQbj/2+M6cNnIyPIi/86QOQDRjdMYOLxY7cZVzV
LA5cOU37odZjQrTdFPbw6w4S6jypXtQIt9KGjBgRRnoJz3nCSplxseXe5uVYsiTlixIwc7mSFjMJ
xooYz2QIOj4s6z5BzDtxPfyflUu6+zoG6vpDY5Lt8njdu4ilz4z7YKS49w1QKTkzvTTMcQx1U/Xu
4uWG/ZXvcSmM8nAIVMGtCOrFSzKacynh1Snfmnne4U7Iw0bkis57guwjPOYy3cIvr10jY/WbJ9M+
o+1KBARWwxY2/NnfrNG/bvkp2a1zq4u3cTdRX4fZfFs+7SD+WU2BWyMnqKFExqGDqFy2nAFAtE53
sar/eVk+zUDhQc1/qK32Ylfc13TBLGkYgDUHvZp5zYFgv/v4Ld9BUs6cM4QEjHCt6D8rp1Xu1AL8
Z0uPu9b0fks2n4SZvJzxYNPEHH1iulEmnn5C24U+kbKLP5vspmDcaO82GuwrMJuTf3AHK/Yo1yiJ
WfhnVaK/b8v7DmF4Lml2KwEjZ/IelgcNhzYOQb75yE1GCLmyFnQ5f3McEnWBKXh9gwkKUBirec67
pBkbkbe045/xMqzrHzvUUUGW9ThLMmS+E1RL5WAYEH/TLTLVbMO3+xNDsTfy/2th0cHtNaXzVQQt
voeHRFW87VCYYuY+Z8SICh/yQnAe0c8VDptWGghDv0xjjh1lJ3SX0niMTKKMs1v+vqvGgBWQGutn
iamXN6ZAEKzRWIeWN19XzBs+0NmxBYg3plvQIK6EZdtrJWvF4nwjz9h7nNqzRXB6H76phwGq1w3W
BRjh3EXn+fb5ZVPtD6r5RkUi1QpkAZNdZzKrSyX5wgQ7PHeJ00UiTbmhKGilwA/NaS0AGH1LTcKu
Hhb10ZsUB0RalLZSMOo5E/1L+VFhyZ2bWVsVUGzHntC/VaU/B9onXg7vNw4Z0AVPPybwUWgIhyYR
oQhQMYzDps5av4UyvE9KuaWO7LDt4KqVENvVWYV76P3Ykh1JNLLBvuAESNRyk+tY55YLpb+72quu
XzvbcExG4USMHUP8uNyPocT0fL5FSt0xb4TfENBZDzsXZUx5AZhlF75Bi8YvRnJ6hMFyJsa/NH5p
8LhlD+6EGbuw3XtrwNnVZd4+dDBq1WlCYwNtBSyFRXHs8SJ65Vuw2rfNCkn5WgksAkwJ4D3XJVXr
w3C+wfh8EEeS8IPgisrz6Z/vFTnOFrParNXqoIPILc2ysSUcRGSZbE5+XjfMwTiOoSP6xEEv9nz3
Xxxpb3zwe21FC5QnXcFBZqN4cxm7kreFygThJgqrK0crCbUG2iZHAlJeGk7xM+FzMBfKFhldbE8g
TL494mTrbKYsMVcNqvYd5K1aT+0vW0GwTSdCtM0G20ejlwkHvtW8KeteMsac9Xdzzgik+3NkI+XZ
X4yTDqEuFMVxRYr010e7tUQ7kdCMCCTYi0mAFTK7FyKa1I8gj999HzYoSuQgRkty7k8td4lBFOoZ
Jq+65qxWi/Y7ilGl9QOc2gWCTRwwmm0kcgWzaduSOZBmWBLkwdFCT0a2cABjwhjMX5bllm7csdiz
hRy9yE4KqBtLKVpr3fnysj2VdVgrVwBefMQRfkrdEbwU0eklcE7ye/dXGNtNt/Gon3i0lvXwIBf4
bjGXKd/m03b361/eG/c8W4/2VRr1WS70d9vSBzT1NfB/iU1cHcXUgcwMNKCBZvx5ijtDAOz4ldjk
ZF3OMx2rpbtf4/OW//cDapufazR40tUqsDJWPdtthNCiAvYNsGvmOS5OiWktTt69LeyiwmywtGiw
XdJ41GFve7cwmpQY0EmbhM/EVb40UiNxcmWn/vgrtEDvHUPO7NCdyYv1BWX9rPAI9Lmr9V50Atk2
3hBNwRJ8JE+BcR6S2SuIFgi2ABOsH3OM707DAeyAprNvTHszKQBKHayXd+Ow81vKnoc1U2qAV2xv
RCLhSfoSIUXF4iUgz9NDjwnREUpNzPizWBC32BcFw0aTG8zvTCaTg9bTGTAvsAFR8kD645QrEbdv
ZdtK7pRmcdLKd26oX7F1ObsrJQeOTt7xid6ZlN+xjnXX72F4sfmwGtrrrv9undECQYWuol0cnIQi
vnnv0GSd/V3YkHRJuwgn9GZjQlgClxbWhPf4BNiQjCVQ+r/CTj2cV7WZVb9jIDD0Rimu+zBw+zol
0eJPkY9jhAlbMu9L5xNZzT+WZqkWzlip4Cx+83pLq7pqD5MRu2EqfN00wmY7RBs/GNTJd3iJP1xI
N1dDNjUCFo2pTyFYrLQjQ2Oh6Tyy9porKuMIMIQImpgESX2BmFaICmsIKDKzAoIn3r3TnVyh+UMY
pwUBu383VoOb/EXd/la9AdDa5IsTkkJ4fgJ68MyGoHr9dZZJ9g3+AykezeS7r7V+EmdJfDTCu6+f
e2VCtJTUYRfKaZgrksspSe41U7DxKg/RD+JCxzNhdVpcfKoScANa8dT3pat3KgXDkMfkL5Q4ZE/g
VnhD8zIjejCAuPXnT4FCQAtuN4croUFpRanD4hvW3k20HUjaGigoJJxKUVwkPQy4pMfQRufGEUlJ
O2VfYW9mSGskYDzFCEQ0PosEm2JV5RifJUvbm7iKrmQ5uxeHfvTtetMvP2JhJ8BIqkR4Mrlgq4bt
v4gYAuaeF2bl+N/ieIR5ZunQ7CJBtQd9+AgliChT8Gry6MXz2IYQsbm2ducHin8ZEyIwMEZm+SnZ
/oI/fmrW4P43kkcsCN1oLo531q+NEuR3nMvT82IV/j0sUb2oRVZ8AIOvTQa5qqEoxXVGXmkJffnp
KBMOEn8+kD7j9p8WwepBFtvA3gg5R0XGnHQrn1F/QfhaXpVKU/QxQkgRxQsg34mVysxfzSZRFw1f
/JNfBCC/gsMbQSMtMju48scuvhF05fgfkCFeuNYwZ2J7ckC5fliytyv90Aoz1OxlaKi7CAtfFbux
G6wcpT96+R6xhmfi3I2k6xvrpfVvWvg91KliXnahlm7j2QnmxHl/3DbL0sZafZv1XyVgdKAGa0Xe
rW29kaGzMzttP5vOhvCwrOfHe6LXhqc/fHHQWCa3wUyRnGwdqFPXQn3RZDhxZw4xSaEXOEKncl3+
RSO9Fji00hhNxfRYhVc1kwsIIM4oS9RqCVAWmESlhBK+qGMAermGQgf88Imhr1iY3E8Jv2TiONVe
Ibyk/jLRiujzaMpmK0nLJMwGRIA1GulL0tHAPngaQ9ljHKAa/1/ZS+71Wd12ltaZAOhrShBt18fg
GBlAswZ8tScF7KmxCErJyZwXxMBhXRwWAiB44XDOQzF03K7RQ09jOiG1vkpPc+0Hei/ui+85E6Tb
H+qpoa+FAOzIQasR/JxDI5NKOWngAqdJ/Q2GIBJOAzA2po2lFiAN2D07Y1MTUVcdf8tSYPCkJ3U1
lcNPz7wHVAV4/j8sHv78aDpzC1G2hadOTtMQ7oZ5YTalzBnZSrLidYrDAHiq/mOu3d5bBnjABi2v
BcCBYU3SEV7r9rwZDJ+fAzGL0XkQ/1z0tNDgqEtJP/Nd6MM++XTmGXfGnsqKd8Vy9KQWk3/bpGaB
HJV9AwniavJFwda3HM3heJjL7IZ7miLnQmdkf5qcVzSQKhazIDLCp6/ZIgXtDgVaQ7Vhrjbahcub
ZAZGAi+EMCIVQoPIr9+ttZp8uxcwzw0jiprftTxrkqd2K5bRGsIf4T58HZe3Zd1LWGggOF0HU1zw
vJ0Ja8FKjBZVWWlcEYm7nwAQ9xQRMdeR0oYI4GYyMRtIO+efC5sv0K3TNVlPHN9LynrFSVXiXSeM
CedszSsOV5tx/RQMz8b1LkK01XQIr4d2/03/HRdde8eQB/GTz7g3y1CB066qxBtrZVUlVqOZSTiZ
OPp1XycEujLLplCSeHhQputUEsybY0Y76pQm5E3BFkff5yU41spZt6pA8DKtC0CpAiBFGwuh1tvV
oHvqwmDdHQn+4i4HMDcVjdHsJC+g0UIQg9uefwINAHMS/KIgyZeamqr/+SJNPKj2L7zBJnySwuZe
eqOXRqptr1myfMAng6bDGnA/GUtvEZvhh9vaR7DB1hvc+18BZyQEiaBun3mkBZ02qtDK11qs57dH
VLofe8fBCL4Wa2lrj6/7clMA1/hGK60c9IIza8XTH7/Xgewh7Yvyce6fIflit9IXoJCE4/a40E9z
c6pyyRtAUiLSCIHKR1LUPU59F/aDmux1A2Ylg/tjMNgcxIsLxH3yaSvOiYZ+AMOGG/VIYtZRZ8Iy
BHLlSvBk9LoPZfglSSglrJCXfLTy9bI2tpc8uZlG7jPHVr9RRSkf5CxvKA0v+6tF2eEIc0NrfTo0
XGuupKfKJyNBcFdEvlQTjQUlXM7T6BVQqs8bd5mOt1JnY+c2IDY4vJN4Q50GurwMH9TzLmf5d4S7
T2TZx82zznx7kzUxT1qqMTobuHBl2rwzNeQaQYa1OuQqVn5m+vt03+2FYIdU68rA3/27ZHIjQDkc
+odBkxR4/8aDWGva6GeBRKhvRsOOhLuUGP0SGl+27pnTe3MVMP9QDkzUFVGRcKQF5WzT2I2xDSnE
ezrGjFB+JhqdFrqVN0cpkpkpbgiErJ4STU7iP/gy7fi6U1Ig9vZPh4Af2qEEUvvR0eWbqC+0QF9G
pWRpUDIuNaF3B8vNA6RvhFGESkbX+BgQjI0zczPm+vWvxt7+D9V5eyweQZY68aFchJKt6nAuKKL6
obRcnpoWZMrDba0umeBIuizTuwcYxVzVP1M4JjUyEKSXmTfxCERqyzR3hZRUQIZ4XLA51rSOy5y0
tpz3QPLJxIZ+0u0Go+HNsqRdL+GfWwqZSTLJHoB8mZJ/4Qhk5EcOei69hvAjViyFALe2uIYHSvxF
TrsEWrxnoAWT7e+EcOpwh9PKaUsG0qp9OUGkJGjzj5Gu4cWt1BNFRN6lP+BwDcMrln+TUF1zX2ZE
3ZGtyDhM6pCjVciMRlCl418Hd7tOnAXlue632IwaH7n5k/HsRX+qtOCN7mcGyqiSse5FloY50p6g
H/mQTa5gBjRwcEvP1UQlGKimInrlmPEBnYd0t5WFn66OL/8GSntyZwqbwggppnb0IdEGB5TinlnR
BkgOgxdU3vyBV5dpYUHNaYSFGF0Be6Zme0oSwMkwehO+dcqiX/vDPq5O6O62bFLRue3kRQSHWmvu
rHPhYSNVvEGqCEyc3nvYi6oL5Do7HPN2PTo42HXaoEPm0vRZy+VxFE/B+0n3gn8DoCuP51WuhfsT
lSSmp7DAV2Q0r1PVhZxexbkO71pbcAXxTtUOd9iTQec81m0EhqRoYcSIlKHh7g3RhS0hOMQB7GoP
bABqg0hUUxYDCVStOt1JlFpoc9J/rjmDA99bRWcXI5kgwpqKZd4olarg71BQhRaswYWTEIFpg+nO
l47gaaGElu9XF08G9nlwLpkJAA991bMfoRknelFvSzHuw3Q6hCGS4DikO60WUXl8XBHZrVVrLFnk
2R1qpllLxQZ6pL4OtRvWL1HopREtbAbxgLihwUdFGu2lgfJ59yIbU2DiSVPDcSWdV+SIK+jJQ0qm
zaL6LVe9Vp0nKaDBTYFM1Xm5OYIfRCq4xTluXE0yzH14fElfjWYiKx55DU45LtNuHhE5qkyz97nX
69rTIv3/BfhnJ95xgDfm0g6swQ+pGWa+e4tA1W9VmbcpC09Xr0ar9NMG2I3n9GViXD0x3ECmMzC/
oWVlHY5h63dfD4vnlkWdqcElqJf8l9lbx6sgYHm6Rwe2oPLyxpm8OX1aOp9zyBNkFWo+nuV3YIk1
jwXni5QY5VzkQxx7GPw/Iw6hnkQOMFuYSsbfd4iw9406/7iHadi9oVJAuRutb6UFnoHbP39m92ZO
AcMJFm6hrv3VsDm4O0dJwgjm4YVjCCNq2BvMLI5dtPCH+tyYHAIc64iHotpu+dEpXuxKhGHOg44I
shemRy4Dz0WIiOTV3z904tuOqETuXTvtgGMeUTvpJcBnqrC3Jnww2k/sfu4adhl+J0he2IeW8g2S
/yCg6K3SNgzA0pb9SVKd4fd/OSSHYoVaY6py/M/vzLeK2yKXafe0KqUGcdwxRWXlc8a0z5U4VTyb
WBjqiovQqmr9xrNvJc5EDkxNggWM2dIZ55MiR1WpJ+6G4VyeUn5oMDeSfmYXy2qhAxSfhoxYoEn8
0JUI28a0Y+u4+VBcAjhdePH6MNE0GxgiKH+1dY66NfCHOPlmEfI38qPV9MFGVb70tMS9BQA5/xqc
onAvp9H4ru5+p/hy76bCF2dmwFESGuFTjd1C8hPgyfIdv21R6q7KNVyty23x2RTQB0jxQDxyS02o
G0SFowjwZlUicTI79EwkfaG7sOlHtuKkrSJJ4syGkeNC2H/bdsR+LYU+GGGClLDnAW3jo2TDjSXu
tJFDwYZewKllzz8rfRnXhTQumBg0UmBmP7ToBw9jhjSnBR3sayhej/iVCYrWdQYGnMh1tKbkQdnT
SjlMrfvSF74fTQCYs3yyQBkDZR6i6qlyA2NSxlyRFWTp4BlHSn1wqUobjdcAePjg9R0fHi+5mZo4
AhokIY5tCVpLW5LRRAAdEMbvdtv1yWQIblyfV33uBEM/Ezd/NSGo7CGQ8luY6ovs/BWAmkw03u6F
/EXf5m9twD/toZ0o4vuTnx1+YUd7hQNdr26FlAEPzfQcNwU6AayUHHK+UVX1/JIvM/tMf0D9vFnm
atXgelAd6ckOz03XK6F20IbekYTFFQq+m9a/O0/gg6jtLTkIV/8USzHJFjB4y8/wK09iPKN5cIwY
O4OMVEDkL85lwjqqYleGYr3VZvQASw914kJEcEQhfNobmk0mxbDXLEDSuHG7zXx11xhyCJy6sTdN
rT/cLFCIhQg3Gz+xK90hb0cya+HDGGwH4Q9IrS+K3ReL+i2crMtwfN+PhC/HKgn8G3kim7ddRNU7
8ZMpc50ghNg3XCL5sU7Hx1eb5F+csCFQTdCJXJzyW2NCzxWbEg3gjiRShfvKGvfaEtNLWmidRX0v
7Vsvni25U4rimjecTNqjHnvB46ls2fFoQpju5si0X0v3/8xZ4WAGiOqnAxLJBx5XkpeOSF/PtqOU
6a0dh2tb4/0CSXkrAR0dcaNyJUXtIE8Ynu2V35ckLVcAzxqtYb/h+r8U9+c9IzE123pqzCwhKwy8
ZL44bIVMuMt/JjYKA4C8gtg8wpzt5F5jWrexMFwcGS6npoW6q0G9AARsWuW4lyFNjn0DrYgDZtKl
5MbJBu3xQw8MwH0kl89g+I9SuKUYrxRuP9qReJ32UyXpZdkiZIm/Yd8a4zjwKLyYFbh/L+OXSGcz
+qLa1HLG2cqRuo2gaRQ1Lf9ElPmJNqln82/uESJK5LHT5xHh6cgW+XLgluSpnYz+jFh/F5recd6N
p9hqwztkxWDUpP4LmnUVT0ByEp2By/Ci84wGh4NQpAvZLwu5LnUT+VZepEpPuiZNv/EP7Aef347u
tNkNLpiGj0CLQZ7gTcDteId4irhmq86uMp3LJWI8MIyoJo9K4picKkKM0oIok7fZStK2jvNlg40P
IyY6/NI+Rvss2ui6rZCyR/pjCvILObaP7BslHMTKWwLMQsvOHDXzMebWgAo4ECUN6OLM9mcK6Snp
/9oloHs8rld7VzDbxEuM9cBWlegaqjdbktgfod3LEDQgcXotAn7qlnQl8Fmez+nw11LrxzZtb9aC
SlWe8NHCr46ALRhaUNB4giDj5keosiZWXFMHh+9tB54iQ/IuCp0Elc8MvKeCWe8y0kfe6mCNzTlP
vMUq0l9NGtRZLDflSqm7LUFhT5ckzJu3RdJ9oua111Ci0z/HBTVPfytCn4tW9ACLGVfAVlDb+B2u
CYHTmQ3+yjdjlp4iathS2lL1UxNFJK3CqjAd5H8Nw34KVfEt9OIgIT2abJvZkti0rjcd9fToT71x
6je3XD4pvh//UAwEHpHHeVT99VnU4TTnR5YXOk3yNqXLZZuIQw/8gz9aar9nbym8FoDfzTRNwbSg
c4BDrP+HmDJ8Csydj/yEvuo2uZAzl4zKjW7/1F7+YpzkmC/0olTCV1Dhz5+FEwsKukvE2f0CWvKB
dVPhTNa1x/sd5h+/IPacf6enxTbMJee/SHYAd7eVEXiiVXj+G8fjYnB9hRO8E6JOs/hRMcvd87oU
2GlRZuX/uUVUe4lLsO+bQowbEEnXkX2e9goDaZrMgPFhmmuYSNOhLCv/gceEDtxFq2fT11gPbQPK
91gxnehrAUlcTCCiEMlH7JNwXn7bCriQxuyFJPFHLI6uU+BpOWGhzYA9/MmMmozqOa+HyVULm5zK
wq3Ylo6rEpLIm03MzE4fd81HA7L121RTFaINBhu9oZoL67T9ITwUP4MB/6xvcElqBB+LPUNhldS6
PQ/iSe1LuYruqPF3ld+/czw+rp9o3nVDX4xEKIB16s6hoLwVOU5scgH21heaDUyCGH9PrrAF0XvQ
w+Yka+V0+zs++NsUFl5tD0TSaaohWAJkxTYBjKNyBhAxW7P+iq1t+3qPFNR8EMKm2C8tA6dZ6YOn
PTnCgNxRn7fF4qpTuIEO2kPV4AUFGQtxa6Ynaq1A3ONzNJE7DqsqPHcItiI3DYST+W5lK0PmYtxu
p3LR+jNLzKaEcZJqK/XCIb++1Iy0HaWy7fXaTcxqLgkA1I7g1zhXmmGLc9ydgnIRZuSXLlDvCuBL
9UmhKcwNcog7f4MLC79niF4KTBEW8kAfIcQYWuRI6w6Fw/jv+zT+Xu1/mFI4uWX6Z+x64MDMKSxH
TWDgaV06dj0x557VKnEsORG0+NIWPC9tNV6JRJE9V/cqO7N7nGO9TsfcIfRz0WDc1GFHXW3jsqTq
GBRMy5TOijnRA/OY06VMxHUAyVBAVHsdSOB9t5jMofonFc5Fi9ahvS+1CB2CDw6RADDAe1t9tbKh
fxPlB89PFcBVhYYaH+gucUtfknMkF5UYpD+9stryPnriq49z2dSt8pz5GQrkTokxsVU9ps78MyLQ
vE9aICdWI0Yxhsa9WMQnvPPeKpqSJAx7H9TPCYPY/14t+sr43TBzGdZFtmKo7l6LizCLZUdtJgjq
LOrJ+Cb99IH93kYieIihVVavt003eILs4gAfM1L6wsZglwo+9WsLUb9RNbRqg4PP79Ekmyyx8rs2
wjHlzu2n7ddqKr3l33LLAwN0aht8QBAazqHZDSPz4sNNLdd1i6n09oCsFl0WqV7eiWFnLl7+uP+b
mJ6iZ6ZEzh0PX43q/aUtDqq/OLsV/codDlUQwxeXYH5Ek+WbchyxPT5ls6RccKtifCDaGVl17Gbk
dqMsrHklXLTwqxiNNF/+mj9oeqTNH6ejALRoBoinATfidaqmXFv/EgcUh/9AyiPYyJlmXithil5y
zxbgLBJz5po/XUhcIhVqh/OvIxTVLiY9j7+Sf8yOCcHX1kus0a/KzrSwNegwl3pRarmxC/mHFA0Z
NNr4YzTmMyrdag5HEQ+b+8NxDlh1bx7NZvlDIEJ5EAPJdS8cAMQ907ZfbqGghl8quj5r43IEttSo
WEq3mrBtYlNN7Ik1gcqgITS8MQLoyZPGDdd6GGgwHerEgktC0uxUQmmp7oYs5/749ZfXfeOjom/I
AZCWVyWzGkyu1XKndvZqMKR1YhX0IApVxCRTuMpUz5xQo3c0HGghC+XoBZIRH7qc5b72S1EqqYJb
hsuQ3czYJvQeHj+oAsK8wAtmGn7M8sH3dYzRnkPMl8L5+g0oP4A7a+stz0KpqlHANkjFFE5YyvW1
oXO3LGvLC4OnIRJX/RWscnGtn+109scLpXUJ6t3XWBHpIhdXig+IOzKkHEmWPOmhoJIOkCE72IjS
ebChKGheYBb9i/tg0HyCRhjKpTMx/AtcJoHnEyo2hNZ3H4E+cqVMrFurJQ26R4eahIJ5tDDv/5jo
C2QgaWGBbEGA1dwGUyG3NPkJAXz4GtQAil2Wg6I6oK7hl6z442IhPiDTmRu+DexHy/TgdnI1mINz
Fh8/9H5txAzDQvA0aTQZg/K9OIyAqOpKRVKUIyNUd8FgnET0Eal+PTS416G89mi4+aQ3yJZkfA6L
b7qFZAq4yZy07vhsj+Iwqj/Sy8LAVrgdLZkvTaWa0cTPjsJ36VzXQLoEOC1+wz2vkk88MZXkKKzw
gHy2+YASEOeeXHEBB7uT57d6FKimC4hdeSHupAyrdON9sJnMY4pB9TIzQCvldhRumIyHdbb/18XH
PoZSGhyF/4wsWckxMnV3K8wnCHEMDsN4bT6VX7yOWi3V3Zyrqas4fN2YksS/f/NwAmX7DnGRIhjZ
ArwVDuYJpqu+CneAMveXMX0NqeBO/JWImhyA7UPX8yZq9ai4uax5bYZ2T5tO23ZiH0Y5oLu4DXeF
g2pjVua3OrW4v7/EFr9+hXevq6cXhUmNzGxUyfDPjEQa0nV6kcVs97/+5oSssvv04dhjYKDTwpBX
mZquDMvNxTUSfuCrQIDASws7cbhu+DJ5C6okxdiNBet9MOa1JYutMndFV6AFaXJ67uo66IY3w4+p
obhUu2nh70ohk/pShsi8oVj95kQo+M9KIA44qGmWcXTYgF/9fYeWvgd+5UdIa1jHZOuzQfFc4Oeu
pVWfd/YSwpqXZ7/9t8GwaaxhcyNDfm0KfBv7xrgEUBWw9zL1eA8D3xzRE0V6fnvR1oRDlNzjkM2r
PzM26zEYZ5M5AENbBfxuX6mQHmqrPkW3dtIVyI+bidYLV2c9CCAEb0taqtgZZ0TjyftGB60qFzn9
dORKGaDJgIols30iD57r9MQqNWPs4NW5+6kyZSguCPoXp+CB6U0F78JyPkLbR6zaz6tyNTPcpdCa
O0Jd/tpn+Wm2lBZLvxxPn9YrJit1zSG6D0A6xUnCM6zwR07VVmZQFuya6Cw/UMkDmdyvspjb6dxW
TfWX/BfgqGHZkXD13OQ+fErYt7Nx98OObDYrvnqJydY7WPVlEMz338sA/DDzmkoDbWSeE4cDtFoO
ZNUyoqJY3nuluuIcGFglnRsqR0KXddg7cUHrC0jrk6SQwPjg772b+v5kS9CYMq4ewv5ysp14Hr7/
UIonIQbneyEHg6ME3WWh6c/aD7MicPSLfYKHtHehayeOlLUj6+/1HSO5FszHDv15h5K4QPY8mzMl
cZiqYZBKmpEsMUfqQ6ViKihwy8YdU7jMEe83lQDmxRPp/znvAjFX12hvVXIp10j4AQJE9yWE3kTi
kJ4yUiw4JNo9ysxQofrSlEYmEgkBQevwGDSzLd96jEzSRmHxylvseh3OLHQXw5Bn8+1L02emow+G
PkppKgJ7Quhw1ydgLRzyz/BvdXtAF0oDamnfRkkUHcnI5YYWBP8DlSv6gBxw3phthqeDrv/Jq9vL
xoi7JYCTF6n4Ubg+jp/e0GUPHKdUAVkk1GW4++l7WIYL1hkEfdw+y8bPqqCnoT8ydZvODcB7K/JA
Uy7Lg9J05HhL0WMAwzDT6nKqLvTOYay91oe2CKKAGbxHJHn1/5FQuDYX+3snF6pe9u8Uplm43qzP
E0FxAEHMTPgT6jtqkXNE0Pka6RXsD6jDaYNXp9YI6yn1s+4qYJTm3mIo/E+H2UCqLhzS9+T8OxgM
YxHhUkKpvUT2qdCvKK9xV3Fseg+uSR2nFouBDSPiQbB8anWzSjDAHYN4pWH/pa/mT3BtzEZq2v00
7qw4jgQkjqlkSVyUPXBaQprC9V0FhVZHCFZCXk9VMDMDlFQMxCVGUu2s9RvdF/H3ekMV/CTyIMVM
6rNKJjjnxcpH392MMNbWUfVPv4Gn/bUnLGukm/zz6uJeoEoLo+gjfS2OCFRU2hpSwCWr3/0UL+oc
ljBaF6Mpg4yxQSIEbadhtG4Cixi95NHdZnNJUlpbocuBxHwEiTqeZT6+x3hJIbB+Uz6QKes8RA4j
p/cdt8U2e2rJdAzw95QrVS6lTQBAcuM+CTVt0nzTties5CWoUFxJki9OVFI2BgmgUwV+7HM3pxuw
lJX7Rkw/M+oiWx82wYOrwoR9GYoOUt9dUsD6vs0D6Nf/Vg6L/1kKqs2cJSyc+1cuxBD/ZnnPsj5p
nm7bOB9MXEWNYLDtmy/752/lAaFGRhBky9nWyjAavU933T9ntAa7AB9W3NnnnFj5mdnVDHXfMfTS
C+L6KKevKi3jqQlS5oCc2ZD5ZUtZSveqQDiHOH8H+yTcMycLzsG1olY7sJSxO54xm65W+KIpE1E+
L+5I5j3Jlu4JJQg5WKxdoUxZ72oLxPk43PCxp5cerqMW+EIamzUZQp2Fm9mT5QNfXtnTeDS8YhKm
mnaiRpPuoa8ZB6DflUnFlo6b30qcQ3RyiVORFWFlKxhOj+PR/fMehu29ppPMqjX0UvCkV9YmQ26s
Wq7/uWl+ftj5KHSFxI0XZNU1NvBonuIH68YKrzuLIvPWBUWNxxraOMB72k+T0WlhgC8DPBh3n/jt
2Iaj13AIRpY33t7UA2rAZn9ylV5HprRBgPSdL6qu0lmaWNhAWSJgSyvpZvfkAi6TwQr/MmSClOk2
9LgnURHCZlDH/BdRWEvKBgv13aUeqjlFdou9+v9BR0SI1nZTa4mfUzMz1UV9Urgckq5Z0MLIyx1k
Cp65EVbjDk+p1nDzoKMA6Dc2xZTsKZm7QJWzCM4LsycGqlvifv3WcjdUC0J0LhWKWIc0pPS9gojY
gAgwNBqrhja141Zvy7ZVMpYpKiDmr0Rzo5eskEDDC0x67fuqoN7K+fp/UnWU4ErtKCMG+KsQtCvv
7xKU2QaYB1g+Glxbx6+G2FYNKZUCTeOK3qXyqUFUAl73tNe37y8tV65NA0xlAohEHM3HoX1vYbfd
7sqK6GhZLjZi3qPlqEAb8PdFbVt85BYnAFGpGdBkkSavMFlXzdwlc+gc5Gto2/bkVgkFTKOGV6Hq
zmeFQVhzxLqxP8kiRnmZ65V4ovwhwo76cz3mnSpGFZ+VjK6MHVssjDiPdWgu6HQpHLwUZaQSw8KK
VmRdXjvgqc12jChMy9rqC8nvMTkShALUXTcOOnp24P/h70xiL0XXeyhfmtu8/5Bk+K8eyLRa8K6F
H/FoXwbUSZetvHVcFiHL7U+8hoOtWbGrY2WUKpYasOb6BILKQ1HYJaHWsMKab2Vvu7+m5ejuXmXN
8V1WZoYhik2woWbjnPH/MzcRAMTqnjJ/ua1CmEigtwe+/G2IXVp4pOqEYqiDF+11S/r6b+fiYwOy
Iw2d0KAcQAXCJsBzLOsu2Bqd/syn3S4KHAURKETwvoRz655KeeNt1Ht+HunUmgcV00rNcRKuQH0d
92TI1g5DdzTTltxExaSQybJWm0bOCoiFCRRfngMTdiKqu2md+SbP2KkULctWZ5TmO5f2cYgLF+xw
/tbla7GZQUkLjoVnapXGsbQcH8ALi0e4TXFbgkt5ET/MmFt7ekuP9EdCTofSnE3+4tECflClFvqc
ulU+lajul2vF3HnhOrqzF+0RgRwnxU0flVJHh0TED+n7oxLmPMSk9I2bLV6WiK2IyE7VpJcs1mhd
MavnPL27/k/2sBKb0ldK7oY1OMeqFLfqVYq9I40dSphMP2Zy14TOgNS/ISkOSvex4PlMAR/IkXGz
FwPfKfeuM3WwiRCt5bLFjIGB7z344Vx6XJ0yHzukN4OYMC+xdIbH5co/QyS3Z9DoL2dz1Mop0WAb
HSSTh0iUotRA11k+lbBl+Y5EUG/8tZ+LYfATamiLtXj96HaaBF9i2z7M3FB000iWepLwlp8xpg+n
rW17p65HcScrFxQwJZ9+iP7KOI3DAwq6cuRbMXWEPA7xBB3xC/OGqgLnGcrcmVCVFfdebXTR6Oh8
OK46Gy0r9NYw4VIQ0z51UsK/PqS6NhZmGDPrCbXhLMIWjz9PDePfcNPNZ1+2vxoldkqizOr+i/vd
V5v9H4orRLNy2eQd22vI92nHksaw4Zg2fhX3GAWINWh0AEO1fGj7l4cC/bm6DtifKIRz5hkuZ+b8
IwfLPSjSMIlZ6RsU9UBnG0PN1b93EPFhKIU3B9vhQtQKC7phi+9l3waZ3NDIEFmlRDZPvJxoBU8y
uElPyAS1sPI1CkMaIQmYqQJizyd7ksU8uqWQjo0TaGbl7+XxaWz+fcLuInib/3N2N8FUXfR14Bs8
nrz4JdEstg31tMCMJnH8dTqjtIqa0jUqEUXNh15MrNxOpL6GubV9IhCQu6DAVbIxGrm1ex14RTIp
89TWW9qTWc9lGfcYgDvgxFHrIyN7bYCEEbHPg93rh732pNa/R2v4zRZwg1rNTF4KErlTiOJtFvxe
+nXyjvEB3r/41Rg8ocUoZ2HwfHrUrMaY/rCU4D8Rfg5C9fGmXwThY/F7SYtE5ECjUp8kde3UKUB+
mvnldNKV0Inou64PZjkJ1+ChwEKTrPrGvJs4www63UkUZmGPduPuHxPJl8RQHgccXFMGrs7aQbVN
RkTQMAptRXzT3NpKCKEA2epEkhTSIfST96X65a8x6m1Djqg7uW75OKUVd50XDF/DNZt6QX22wVKL
LM7albQ9J0NftbUkg109T6+sM4xhijI8SA87cx/Rdj1gqKNjlHXDqhqBuja+CRI6A0kMOSxuudtr
EEvNpOz9kdHl6Zz+N4av0E0XLuv+xxxLgpaMwJWyuD341kF3CKMtsgVvqzyS+0alDu0HktPdd9b7
oRguCiyhkTWwfG+hYvH1YYx9v4GRIXGyj905J/BWf76DwvqnnF2uCVY24elFL1ZT++9OTlKgp32e
5MZSvyx6JBsnzBUJHFeRk5mfvtlLVBF4eokKvkVhpL9IEdVYnNLMs4DMat9QQGfN4Icz+T50+bVl
GA/kY6B2nFn7Ksj6lbyGCuWbIyqewOdsn2kvDJrbsRBt6IQh7MyaHTQAAjly68LinOMOVZdfBwyH
Q8d7Zn5ZfMho4ofI9fqpMq6bxUDhQaptOK1JFmPJyoS9Sz767mLGQ+3GwyyJre9ln790e0BIZBzM
1CuoAcIeawlcph96FREJu993nNCUae/hjrTGE4X8o517ePf8xDVpf+vpWibH04XcKY/W0+I5YV7R
mJmx7VhqcmSm64L6SeR70NEzeFzKywchvKaWn1TkaR3wsnH+StflLpda+EQcjFGoEcTJB31pTaE7
dHUlu4GMj9hJXNJCdKuFtLGGz6TXz1GsepTb70I//cl0HbptqvzBzXdfcwd7crZqodaQuh6eL3qU
PT3aNgo6UMwEWBOk8tTZXKmQ6RDNlh9+CIp0uKzd77XR/IrSjfOFkvI913bJ0dzwrjzDFwJhx4Zw
PZiNa8tuKGhuS1az1CWhNnOzyktQWppiLYGn06BpK/YBw8d/RecKhlaKa5/W2m0OHEN4gWjs2E2n
jths6rS4EIF4z8os/sj1k5/Y6xF2VJY6PTGWVvMCuMJHjCXXJPLnDvdeZwLtDNDVhIvSnVPA5/Wx
vocLjhemLShXxnPD1NzCIVV2O3KW8orzC+NqpwT5Ju3mkPSelfrtXx53iKY0a5oP0BskcYzUL/5J
AQMEwgvuT0pSM7FdWMxPuyIn8aQqOJdrOgLu1/iF5qWMRkqLLrZGlRnXUZofHWJYy5NXS6cjyLxi
cAR+RasLJOQy/BwDWdUvCe7st2BIy2RabFmTQ50IeNIMWHmli/SdOPyVCSZR/6odmSP2rg3V5tSc
gyMpUnJEoyH46potZCKG8nf3R0GaVtAKvGKUHXuRPyHJHtuBxavdqVodhDOaUaw7iRXD7zEnbVdV
5ZWXIS53INH2OQn2sQd3/LJaZI6BvyP+co7ugFVAXoXfIc93TNGPsxO64SimTDRUesJzje34mgft
X1cI9eJkzJgmOl0FA8fG6HOHjMtIBDsEAs1NZihTMlqUSZfJowea7rRZDqwBAO2/ni2zJPkXBgqv
3QSf0DiwG1RoHZEJqoGpceHqjOvahpzJutS3mc7dz2EB4wNyFHFrXg9ZzBk5pOCDwomEM0bNmIux
Xb+E//VnpuL9XjCiDJmotLbppVdCOlWXSOOBCYBzcGaVAC2lX9fVkO7tE4bTOeRsqVRWcPaaoUwA
j6biRxpN2AtqSFCFuZNSjKtQBIGUk4sR7BU5Wye3AfrF3EBGriW9ceY+xQLt2w5eps92Z9FGMW6a
pPtwOdxj6nwQ3SMVmzr0Sb0olg+EQv3HOxWh/LL8DMEXhq7IJ21CyOhVxF7j4++txZzDZdysYjiF
HOek9gVvIqLj98x8KSLGaogcS16hll8QAzt46ksjose+ab7qak8oNzHnMakYgk0IDRI5Ms1qMyUk
i4WCv/rQ73xiGoR9GbyDZiyur6AmrhDDZoAbJ0wfhjBoTJPdv/4MCjHNfrF+ZOTciYEnCHXcK+Rk
P3HBZRoY5JR+6+vDi6h04ppenF2Hnm742lb7AdJD9V7s4GQs3jXOCM5QXXjusacDj/1iIdiTD94i
vFNlBSpU8K3cCanZrJlJXKuxg5fPVjrNNldiCkIXPyTGZkaDavLSHmx5gYPExLaHy5jmoY55s+WG
WPyzkvHOsPUdoc6Xe7MyfZybYQPf9Uq3vWwIsbVIsSRbQtGctnAk97G5W3EFpCISa9aqPBaqmN5T
3x6/5NQRce7Tv+i+RaFye5ACqTPIOe2+nKGPXfUZlZqd8lnQe+9JibOKmmVbhyE+0QiwFap8bTe9
akeq1ikozi7fSrDO/Zfe9byO1g1vhr2iaHiBC6SSptbeN51BPtH+LxxxUfErEIqZI31INpJTCAPk
K4uuPOAnfwi2x9x1kORD8BWJ01gimRKdWHP5d2DRfxxkPTQYa7bTvMclw7Ahq4KeegC+vCmK326K
koy9gaic63xLmMjEbzv9lljfHvOORmxDwqyOEtmb2DAqUTIgEyBt0B04L29AOSmZ0JZlZ+vN3WOb
4IvJegHhPLGFhD6aP5uR5qNbt6SkHer/ix6wVNvB+JhfvB8KQDp810G6dgaTHj8vqRP5bpnmMA7x
zXpv/7HmwAtKC/quThk3paLGx/TAUxjQb52P3XpIOtupiVO3MmIH0bBsAlosbFzLDERVxk7Vo2kt
amnPeCEpg6s6/fNioDFpkhmGoWhkgRZ+iLey6AhtnRtsXyr7OAOUpjwKeiYz3bA0UsBRp/lWuS/C
MIh9pGT+uaIWxqzODH0Px5Cpx/JZaUS/C3atjYjieSvDvZnvai/UaGDMcgxqq9f7oRuUREjedaWK
bP4VOa/pJKhmKgIWsKVGpdM8d6l5DTu8wSo2RG6tkfIlyww96Bi3QTxbPNJT/OX0pZ+eEzHyXaOY
zr6vbUvV+Q9Vc+4seTBqF+LvKP9wupIAI1Qpt05aLPDploqrw8Cbj3aWjSdcgtv7OKB6d+S2V1AH
uclFEb41GwV9mexGCgswKTor86t7U5abbiMpTAxVa6xEXva5SVJi6wgr9X1QwydQ/7OLZuJEOlLH
/8zZ1R1ML979mNmnctH0GKlA1B/JTTSrEGkxMhvbJAV1XiAS5Uw7deS1bHrkFNCo52pZD4JwzVN6
oNjfUYQQewAGqd/6Dca1Vr9yVEJihaj9ybuaidDqPqzHUPZbIdBGvbikDWYjNimN+jbYd/TEav1J
Ras6mWAkCMn54CNqU1lIuSLlOnT+r0kh/JcLjTlMD0trB0vQBjaXQIx3vMJJIW9CkwKtq1OLLitE
TpJ37Xcxf8LLy7eAG1C+S1Jd+UXhJmO0zC/m9OPDe4hrLYuiOnTJvt7yy/5Ll41VsEnbH906HVa7
tlMYd677RIoHcqtYHgQRa2P4ck2nK6BPUCmVkNmO9xBy4hfYN5RB+Cyn2/wDmCvcjEUzzI2gbff/
Iq7KlrCS1cQB1Fh9Wf4rRPsb2GiRR/Ah/cPanGv7IeQYr0PjsjU2y5IeJbWJxhz+hebDhqdxiziH
S9reeLx57mYz9gcp9vQx10XCvZHtpUu+TaxAziWs7JeqtvqDov8W7Ks1VY41N39N5w4QItwsDjCb
kBRxl0g0gj2kqiJWuJz0leO1BuZBpnfmDoon2ZnpRMQv08jG/U5HyKKOi4nYLKCgjaPCBVneyK8E
BhbbZTNWGawGMdMMxCh6uLQo72F25xVm1b5gZ+2hAaDDitC9Uyn0VyfuQAC8jdRS+eZ+icYNlCKt
CGLW5PCCDqZ2zblRnZsRidatantofwYKxVqxeMcPyclfZq5+5SJDRMo3SPxrwM3wHPFQpn1FTAyg
oX0YRQhKd5O8KZl7bg/gA7+at5aDTZM8djFMMR0dnx3WagJDEXc4iriomORbK30txHk+ZXpDgvGS
pmUubYa47obJ7EnDlIQf15iOYanXACnbGur/hAY5di74Xl0vOwXxdwA/99rjHG1DL9INF5rOFjdu
NRrB1Dze4BmbQCCXCQNoexT8n5S9rIF8OCcC8GN7Bqjfxbc7px3nTsKLyIkod1mNKhB6kORluqzz
0NPDGT0BR6UGKJtfOmblRl0+cBz+2rFsby88B0KZIWe/NU3LRiaTwH76gUcclbH+BuYEdZRCyJhu
JHfJk59lIbF0/ns+faI2Ac+ifkZeLqBX8SDnZlMjHTgdBPooxxJGCIA/hLFIY20FoIOUvYIdDD6y
twFZmmzMcdCP4ErIkniFSW1uW8XlFXQ50gx/w85fmwtWg3fdxLZF/KoUselvHsW+6UKdV1h2Zq7j
vm7YAJXS+99e7dAUflcKLuAFuafrVixIDkQ4yO8GEuv8R8a5WS/J4zG/nwabfYrY6yjpsQ//EAEp
J56M6zm/jhnacK2yBDchIjJkCDv6bssA0xvHvunyuKBPXP23rdFzZpcyTm3LfOcAo2S22Rob42wP
FiilJVyAMRy3pBc+cCS6/pzUWoeHleAor/dy0G/mV/QRffiHn/rODARhPkOZteftlkIXXzV8wAw6
JFHzGGdpAPjOQ5vXMSXahpVbHs4hz93WivrMzNcrBI9EECKfSD1U0s+41WJcTvuEUh2EFeEN571o
8lsr7ANLOyIEZ3bQE8It6/jCIaFTHUaHh1vYUvaVag+nmrahB+qLVh0+oBQWbQ7qV97JY25if01M
ltUjnCd6UeCoVXboE+eCPEHEdqdsCCFiR7OA9snRHtk2SgsDnc0IQi5wi8eRAzkYmHfrKYF9Daid
pR/Fbj6MYUtiiR9iSAZtH+rLlp3F2LMxyhOtB+EtnLqPFIvqCkThBfOXTI86ZNsUojwUr3Ro4m/3
mH1lbi1jbRi+h99Y8RFheuDpoFiG3jtyZeJHj30g/v650Lvhcn0VzeiMJbepfI/MxEbIojnTT/ts
3JmpssJFnqksE/Ad5aiuZKKlosWwJxtqD4O18Ifcd1o2Or3on/8VvT2gTlchKHcoaJlaJtWqQIth
XR6gpHcI/2mu9kkutqQsKAF/fZvCVSlCwMTWtWaH1ZTer03UXnY4fYVmixp05KqDqgbn+f06gKQO
AYzOCTXNUlaYL1evCPD1dj6yVRi5w7hLjqIu/gcqDsuWbC8yYAZG2RUqDlCDefjiOSpZFlQ3Pvoy
7RqmzdXuJA+Tt/7LX6dAhMW4uhb0JaZVEpUUXOSMXf3TcAb5ISmLioti6wISetImqMvOn+uSdmvA
Yo5j2cLPemstVjSlli1Soj9HGwav+J7NLvSTu/YVUJ6Nv2s8YJODnqo6Ai4tX4EANZaktTtdUBgC
Ukqe/ngJLcxgReFO648r9h44K5sX/lk5XKtob8Or8HUJxo7knVThHrzAOk0/3HqAX4miIBDlslql
CtXarPDTOcl6JPjOteiqqVwD55InoVNs01WUmumgWHcyk9OEQlYo8tCR/zN5bO1XP9ZSW0rXFe0O
2QF/jnFtH8Hbj2WZUmb/ZZuBzeA3Yqxm82XG3ocsYoTzhWvA7WcDZ+16rDNhobVPF96ojViBkLUr
5hj96lnC2hJBj9a1Bic9Skh14zVavDwbpVJKTVXGP34nsGua3gFbLdeGtFtbluX0Sh+A5LAzIhIP
yjuTU2zNchukBaNIxv1i4aScQJYgNnU87DXiW6X2gnQx41V1RFND0/6QoW++4N5IEYKgp6ywWniT
iRvYm2of/QfruTm79JmiD+A6QZcUX3+SsfIPDuu2ieUM2wE5ZJaXdjtz9THzPFjSRD4nFJ/SvuAX
yjXZ2SkmQSYJXUnLxEzT8BtKUNv0VM1WJGXCJhwemK8d5Kvc4vx64pEjMExGV+3XIlzfUxxyVdnO
BuKxSBNUTFRw8E0Umq7SHmobkCoqd17E6jfqoG6rETFwsXeOcZG+/XmH9258I+YJIwEAChQkRcAk
WGc4QPPIzG5j35Oxigtl9dvAtwZK3tRBXk7oOqJkaHcY4xU+3QGh21zXOTtzqCnDiYs/Z/o53AqZ
/DO2cyjzW0vRkMPJf6TuPb2h361N3v2lEmbbDrkDE6/23KNZtWHE1uTsZ7sT2ttt1GHqb1c0yt0N
d/hvxkxwQ8V0EkA91jzgyVyg/z9BWhozwQbxr1ltkTeq45W3dQV+BWOCO4ev+AHFiKVjFxZXYwRl
zCWE5eI7LPR3qY3A/08FBblWxk28LXYiikdTedrYolCH/0O4BiOyZTEuJWN21vpvC6A2OvpmshXn
FumrLFAiUweviWH4H4Y8YxwurV1tIVb7BSTXs+t20oKLirXro9W8s3GDQqnMO6S0g45ngkNbBGPN
5dDN72EThj9Pdyy5SgkYG3XMXLQcHr3hRlxsW7V26n9C/zhsDoumlt0JKZxg7nlcDRaWD0dcrln7
0p95NR1bgC0Ur/2XFyP/pvK2tbJpprAsrURHCsvGvEK+fNclc6eqAXsQY5ff76RLVdih660NYf6r
wq5kYjEyL57e2WSY44hwk/8QISZkhlbh9xKkOwH1cQPBup+alWFkjunCXYF/Y/y5RQAnk4KJ1uuf
weEro9EPSJ2oVQy2DFaMSm+shc15Z/CvDH83phx7uXS9eh0C1LpMEmiSRH/E8qirOF7HeiW4kSQb
9CNlAkyHV1cXoE8FvnX8v8pjTF8LoQsCYa9RPrZfc9ckOeZZy6a7/Bl5XaNxSB7wKJ8cbfToz3JH
h7YJTFXJ6ftgRnXRjJeH3LoF5tduINjn1didZWv04PLllNTk7RZyJdQMMv10S/XlWpALnf5h40Tm
/Ew3VApO5M7+RHqOrOXVyjuB8NDY4ga5Ke/I79A3Tx/u2NXJOnyi/Olk2TS2SazKUkl5gxxO/QBo
W4rfmQJu8oDcUOWEqfYc8VVkz0Vq/OZi/DFW1amdySoyvtCo5VyGg04VtGjmZafNCafe59Vi5EXe
p1Ee98dYi1V/rCJY4MdDelcgMyt8NZzX5lEvIaoc4dpiQ3e52uNiDIpy5Of7ID1gnjjqZAFzHEKT
MUf6Oea/3ZwkKyHaNv8eHkCDGahovcNRNehEtpR7Rw+S1QcuhlN+s/5cl7hqemogDAktIbU3MbFc
TiayM4eZxhjq3s+hgkioC+PNoBbl2IX0Tu6oKCdFeIcKPEV1+L3kjUhstLb9PPgXiWsqNWEEostL
2oZ7oKnuWLGaYu8eCswQbA+yiHNdQnBBI08V8+61JlwKF5Z/NG2j2ThIn1LifN6Mhyi7q47m8m4w
vR1LSIcUVrs9V/oHYGuIe1ynbH2jnbB1K+GJJ03C1RcxXxsPs+2PH8eWXdWe8UK6feqT4i2Snvta
/PyvsZggwXNZI8r16lGGrgo3yuDCHEvu9x0we8kZfb2rKhvGAq6OkWDvKoaxqvPDHdquFldqXSab
61GhVrLZsxQOnzDz9BOD3xlW7O5av2gHSYQXJHQ9svxwMP24OF3SJg0ayoVxjXoXOqV+w5nXUfaK
yPb1IxkcB+PayamEo5nGB/DND5uvQI38IMOEOXkHmiZX9IKBrG753t7tJ7EafhZoqkOk24jPAzjR
Q1A5N5F2VYk2v698Fka8UrXVZ36Nya8lm8jd+bM0nLC+miS+t3Ez7k1+pH0ICXJnZpOV5qrsNMSy
pF//bk1Xy3W8nYcAylqFEy1zZS4z7kA2jpM2v1YYpvfaa8RSemTLaaS6DibaOkpvm1w2i5S8BMot
F6VzUgTj5HYyM8EDN+hAcspdBtJrB/spm9E5t8YFrm5Za2MDRiwAgqkioQZ25s1jaqd8tgC2blE/
hGX6gZ1RkQKYnyCrU3L6mGca8dM0jOQWcaF4p34gCFLJJ8KsWD3npKgtTJxKleSlkNIs54zUQNOB
dmajj+7CtJX1JXTvfqOcykLHzPxakRdQGM3PXPQf5z5mKSEkUSOGjCuM7rIpoM1gXL7bQ/Ygt97g
XKKs23Cj6jv70T8BeF9l0OAHfPReRah3qrRXhXvfuX3q4G255w8hzAyu7E3QqOPzTbsj5dNIkBhr
vc/SA+sx0zZrksxZ5LMeu0OOXtBqsvmtECeuTn+htJcoNHJ2kqPzsnsJ/zJzuwEXe+6XNxRjRMa0
BxbdZuFB3bV8K1zvcQEURY5gmVZGudRetx6INymBm/ncmSOTlacs9s8pyVHG3LYDd2dRbF+6kAyq
+qiotUX7yF/VkHpDfHj9Od8ANNLzpIgXfY15vGbCVh5yU5DRbnbeL8koYAkQjRSnybJRbn5et7MC
cb7UMkvuIJSvrO+0apP1JEVZQBl00au9rGd719spDfgHA/G5dBDZGrnJu3Ht19RXfratqTvsinyj
HWgsowodCMb027t+mUf1lia0OEb2sNmTk7Ox4mX2TSAPf5aUtmqK1y3S5hvG2G+DSb9RRpFQKyNZ
eAGhKoiUvWXhmAyDqQi7zA+hZ1YK+PUhUgEluZNUZMk8EIom+6WA4yaTpNZfVy+V8jwpfBK1cBaq
N4J5XEIkVCU4JaNc6Z9yMMbFb6GTns0pAnWaUr67hKYqZ+0hWjn3ZoztUdQG7CB6NJL0u4rnwj/n
3M9qliX3P/NonJ4UQMT7nW4nDcozVeZiu+1YKX8aTeP/RuQ9/nzRt55H1tTf0Hxtv1dQTb2kRl13
KY8XF1z/3UQjre04+V8PLe4aFmNy+BceerPH8duRsIVOlhGaMTY/OjEtBHgV0fjr83vyvit73NW4
3t83A3VGrgQ+MolYEFUUheYmgTqUK4031LvHVJBim0FjraxsUyQ11I1PsLvkudwY8ZC8HyEcCnqD
jXbkm22XVzc1jskjHEU8eauPj4pilGeV8MGUQ3T6sjaxRlqxeiY9Jm8+VxCzuDSfuO2fmw4qruva
Ql15T74CtgDlm6WVNWamjW3FzLpSUxZJ9mwT6r+u9x6VQEczjceIobCGBjpBhv/1iBEvd361TuOu
zByAhomt+nBTA3XC7Vz5x1Qp7OTsLdECMR/76oaTp3P5jPh2L4p7ISkcIu1K6c9luRBViKy6SFAp
WHxupOqkUtJhXmZ2d+9YOUAtdJX5z8WaFG2mne2UIAFbzogkTiHuS30kg3scAzu7MeLwgdLet+dx
Y7yWK9eyQpgS/SD02USyaEIqKu/ECRcTwJdb4Nt8fwzlKsRDsbcRS65UIm0calFTyXGHw8Skz0c+
fuYtpFQ+NH6Pk7w19sLFx8dHvZ3DkzCdc+4UsFW8BhLkt8KeL7qtSZhVyV9al8jJoe+UeVDJT2Zs
2IL0D1ZNzoSWzLr7uRAZUspBiTR8HlFfZIG7u7fD09/cppitysWTRqDGOlqMu1G9lEpuzKAb6mVl
I9X1vyh+5xPSFNR8rMwk5qh1UsbIrwRAGDbi3V1Jcczea1AGIdHJgE135YvIZzl1PlJ+Q+oYusvu
6xc33AEsFJtrNHfueJIxwwzkiO3xA2BIbE/7cb6CQsWYYh9zy0D2GZNMVGyGemI+Mq+gLKAz4sak
Z37kYY1DqXTUzIsOPfKjISDuUqFeF3APEL1zZfxOS8OmXJgmmrh4KAVc/MAxGjvOaCrnQ6Fu5zgI
WrmX7QbpU6WC1HvsmYnAjb9wJFJr4pvpn6lzacYeEBrMds/d2QCTcR7wipPMOvD6a0GQ6L4ChslY
wyPSoJAkz/cu42Hg415NTB8s4dblrJi+rSpNMAT28f/0FEU19P91/JermkDK9KtIV51e+WRQWB+g
3w2SccjAKIVlJu9GlcTQO/Q+O3NsRylQnzkwfMo5L62+9dmHQDiHazSr611iI81pAS31/fzkPUZY
d1PKYLaOcxKft8I8zWMIJA886QOxv/uWL3LQ5sTh74UTJDhvOaqeBPn9tMh2Jm4878sNYP/rau/O
ST7xPKv7jld3tj5q/kq9iyn3rJOQTfTEslsY88XOQLgMEsdJ3TwLt0P7B/pZutBPgqH/9YQep9np
clrZ4scUKFbyVn1ZfV0VguuNjwDML3nh9OxYQECLR8Kjh4bYFO/VEdGxPkGLSXAy7CGRjMH1Zk39
A8kGKt0wterxetoXpzi2EZKQ+0BDEglFtbMkmqmZasAMZXAHhiW/qDjWlWsATg9ANh2bEWKIFaGq
vijOtZw/bD2JEt2e8Xo4cDuw+X9VuDVrFyiXQuPp0HBNV0GOOEc0DU82WimDIVCubYz+b/jb1iGY
8sgfcv6iVqLENXLtjHWx6MMKdmVYbVHytlcD/0DF6TqcvpupqysYZdu8BR1mn3BUeahqwM89MTGw
5eXNttriqE2LIoef8XbmdlGtzUDyELLv0k6+80u67bL7Sf/Nt6n+pap7/zPL2HTrUavdc6N8zCx9
XkdqlfrGq2h20CdS4QqUEFQS5pNL1pGC6ZZWrHM71wtTQ2bQ/Xb0pZQ+Hkmu1mBWHOZLgjsxwvC2
6+y542M6oLoEAth5LxLjGZ+f2S6zffxoPYSEvCZdF4yYZF2vMvsHnW0KpDPCYb/wU/ypCAhSLZdK
KE7u17vSIUswnmZaWbjQbTMFh8ueh1mh4N4y7A8ZSNHmgR3tFdaYGFGiQY21QDwDduZlb/uRDESZ
1AiRUwPswuPnVb0iHVUO9X0676XCnMbAqkAWFzuPeOfY42of3XjeTk+aHu1rpGVoGuge9RQrHVrW
AXfvEGIYxZ3xbgq4cGn85qrYkRqcGgnPDdZQJ53uKFCX78BNUt3Z9gYdCAXvra5RQktpY0NwQQt8
TrvcvIH5ahGxouMG7GfQuNclymNzh7QAenXxU7haKeXV7bKasi2YMVtHiKRGNKUmQzqfcvGBDWP7
rSNKGN6tw8RDc8tw6cVhvqwQ1yhATXjcwuP7x+sataNAYMffsdWHYRMYkFfXTBcvYQkOmk7ogJQC
BYmShMFcnh4TnI1QuXnoh+EEsm8F+w21eJvOMyEPZNI/WEbJUQtdpazSfR+yNLOmFlEkNwwtmTKy
q3oT5+T89MtgeGmkTAqNdfTraGYMqJGOjP3fGebF9HoQgF0dS1FpAIBAQsxLkaPh068tKM1WWH9V
nyN/nS8rM9Xc0K+cK+Zd8SUBzfbCXG1N+ellFtMgVcVaKWbPjqmlzqtAxrxvZ+5Rh8maaJnxeyvB
8NTc7gcJF5g/rVG1Z4fuDIvnvbGNQwXBu5QB3BFMReGpeP/H7sZbp9ZV7o/plzSrSXRfxUznXxnp
L7gD1hiKOxhUOEPWen5LFhUBxsnYe+qw4zIu0yOMvzY2oP56LE05Tck5mUnHUFmA2U63a2giI6xY
aB9Wr5L/OZoP2+ORTOMA9FY+q2jkZIWXjoEZvGWn5H/gRXZpP4528cERe4ez4wOl8kGSKd5KLWmL
SdlOU0e/IbssgZ+ymcDmMgECd2/744fruDbseMjsiYEG5D/8R1Vg93DZnFEMWyI3iznOi5fLI02c
F//8efaUR/UFgq4dQ1taoNFREwEluIRYp34Mq4cYv8C63JFLr2vic9yvlLmWWwh65VmvpDZicDdD
/r/RQ9Uo1kNY7WvrljfvyLc7+FVy9uOC9mqnpdmCh7WuMT/jbhe0R2fVqNb8DpcLDveb7xNTPUn7
PhRByLUusWcudfKIzGFG5Xakr+rXVWCs7tSAx5iA5JiDEsfsJyp3R5RFCdkeGxyjgktpI/6RXApV
Q1qUqVvWpLnRZswBFNWOzvH1LzOheSw8MIQwqlaA1JxJdsHWOxLh5icwjCMMCVqlYQeiFSxRojSp
yeqF03azGASvP4h7yVPM/MfdMjUl2X6m8J5EXNPkcJaW+lFUg/D+f1Nmv9QkdrQR/Od3686cwzsN
udhR/3eemNiS0qanNI8RWVNpxjsn2XtbAcb/8LglbB6vt5OuTcw67oerSz9W5PnHskNQrx4sWdDz
vqpHFeEYXVZuLYhycUXE+kUalJthm0lk9uXBkAFeS48hWzwRCADKV91Gbg5/tLCyAYC5njfJLdTu
B7U64S2XCntdoi7VFsqzxyaFbJPCDjarHC6Derf3lQTAESGU1/2ed7ZBu1pMoeBfH176RtUh4n06
G1UPGs+RPuJsl9fXqC53cImEhm4C6nnWv8AVZWSHjEwwUqMqCtW9pHCTYfD58WmDKfc8csPLzu3R
6AFlmp3uscRKWaAFM1jks2klxdUmv3tLvIVtmCOhPOupP9OrCAM+nDI/zlPzj3nAgoq5uqYXCUrK
Nj3E2tOOMH8u6eR6xdTNhUht1iHsfXBEBjR5WMTpcDoxo5Li1q6e+UdAv8KAA5aduXW51VQNmf9G
gM8K8BSnE3Jbh+OjxcaylZhHGp12CYnTD/q/UKxmL9l5E10RexQk+WwbvAkGaZ218RgH5sMhHPEW
tgb0jD5bxePqPe8DhzKssW78L7wlYOvOLnBeZI0vRg5aASJI9Ylk7LKsmmXDXo7wCSipX0sZlm6s
aX8dNIkIYW+Xn+/UhcFR3xhoYKQXgouZMy6FVa+jZViIo3BGhTipZWphEL7jOg6L5KGLTJuWytYe
PgeRkMGY90qfrrfiS7lEycs9YfSOWwSVJfP9p4QTIJ7pbxf3shK6OVOm6aSP/0KL96OT/QUU1+ll
Ucf+RKfg4mNAlSFbDWG1IO350MIlW0p52LS8qnRQ/bfpEhFKqBvYcTkkMPQniJlJxKO4tvFPeQzb
LxQgzf26To9F4xlZH35fT+ajUFbubV782eTkPif6Z9kJjyKYW/NRdHvJfTWJjK2aL0rbTlvuC8s/
NCD5WtjSJDFv8isE1wv5s+1VXnNcSjHHXKOil+zC7oAkQLw5FjwGd+TplLi+eEBOQ4DI12uYQM9/
O/0Z8xOPtQKrC6WaQDKHZPvSttEKlVgrGbZx1CoJqUUhx4Ja8wGdm+242Z8gCTRu2aeDROibm+/f
v8vtDTqaLNalIQcQg3KLPCg0AO0R/6DQAyNYISTc6WbTuEoCcbWsdOvi9x9DChSGvCCW6aWauiNL
RKGu7+MnxNs6PjIELddCFiWsiLY78hYXNy/ORa7DujlxR1H6B0JYjBJI/yCoQIJ+kerquxa+gu03
VbQ09sL4QRTy+EOiKqbg+VAg3wrzkaUfXsgipdoouZH5rNnAi4hHIAisEddh23HhWa5EdtS8Hd2W
mxkXj3GR+pOkeEzBxBDUGlZ7PE5yuS4uq9n2ZVPLspf0sALukaK7rX1ZLaSDXdCCHNT26LR3qWCj
0BFABfXAP7VzUUuMaZiwOICDTvxHy+MaZgaRadQIu7NkOuYpWnKOb0ZU5v1dBafptr6HloXsde3s
8zgoXsLCxsBu2ZUZHOT7E0v5ntQGbX4v17lIcIG6bcZBnmJMbMGu1Rw2Mx6PYY92wuW6yY23vpve
g7kEbeIGs513CnnQmygV1v67hBYIKAXopthKS437PMR1GxGsttqpHSrWbx0W1tS36PRA0A4stWFF
cPWvUNzHd3e4cS6Z+/eVwMf/CoJN9ESbja9u6GUfQi2/KE2YDKBA7h7RHDEWeeP2tlAfp61RRo1l
eZls9BgxlaRqpqmmPRZ4OpzanTu9Y94UgMrandid6KUOGvrI76zFnX3mI0Xn57NvkOpnmL9nL2qC
L9py2kzueozTkyo+3n3B0S1E6xQypeaCZPTd+zNQ81blCjJBUNS8kDubG92nbHwQYD9L3mqyPV2Z
gTV4nNNAh3dm57iRpzlH1dkBVV3UeGTtLZFRkUHVqwR+8G1Rvkph0G9JdVunL8LJc/r7qHKF+BaJ
TlH6I/1evahk6MzrFUs6AqjxIdQmNd8R9CK1Ii274fBSZ0EyICzrFun8O4fB12KI+ojBDzXZnIFN
GIj+M99BDvlAVWIDoHYNhbH6plscmEfD0R/bEAjz62cNXx9WwdZ//hwDMmRLDiBFjDWMSi+zBZYw
GmksNNkg7EiOi2Jxj6jxAxiYRvIJ1SXNcmmSjeaaKN7plKJkKcg6FILcJFLR1ODoY4IreiHYoE5C
mGaivkYlSx7G046oH4HnNiVGBlPWvfD9vQTwrivzMIcGYGT4giwIdJwnxxk6TGnuZ/iSIZTKsow4
0jCuavxX8Qr/FZNcivypiJUFWtqgESbH3Xac5phRIBDdUT9QksXtN35bLlms5a4W5NxOQ3aye7Uk
EEVFxJ1TyxFgYARnfQvjAVylyOcv1hLbSugAWBoXxt/HdGz1fFk3b9diF2anFp3oQzEDCVFnu6yZ
Z77w5/fKOyJ1wPLvfxxU+YQWabmM6wwM3tK104n+ruV84OT9NAadymqoXUx//QbzClJpxL/ZK6Rh
bqcOlN1m3FPlzw1CAjfBskOPqbgCAAkc/0tYF55kGolisBBHZmcYRCAX7Xs/Pw7NWqIehRoYFctc
TNxb+77DAXXDNbDRbsdBk1W8VeEa2+XjaltU1l3lC7qdWuVbL68iD15u2UXHo956MewF5BjwnzFr
IsBEWWu1Lmv2F48jf3dxswBmphYZV9SbqbnaMnO3BmH3uQFotvgC+zGBGb9L+dkk/2AxrLxSjEtW
z9c1yyw4tDv9K8vVkDL2B8xFNrgJypsvDZLpUNST+KafUUeC+yXYrKmC3o7WXymq6BF6HzKsAy+l
DP6npCHg5GzyYguQyGGhgWoSBDYe/cdLIX5tLAawZ8BaoF2pcAY75evDL8ywh4rxHiA2yJgjYg9Y
TTGmeK4AioZyMDSOiNoMHmo6QxxfGBNANHQCIc6FRm7ssvB8xzLaTKJWBnn9MmOQN3yruUQqUb3P
HM3/sQ+u8c3fZ59GhUpzsnNMFU8cvNrXh7ZhuFcr1QKhj/QE7IGqbRP42V0noyOkjTwsiWwF5RHV
SOteqnm3G3M6jPaSGezYGlKyT53ac+DOC090uN1yyIS0q2E4IE21SyT7r+xHQwMtQKmqLUHGFjoV
9mMRKMRjctQh8jkDVsRZGYCSDsUw+G6lyqdOmGFf4BA/o9szLdHQb11hzQfPyuo60NdTI3Z+H0wL
60LIwO9mvK5w72sY2nj4RPCMqs7RQaMjFivCKHSf29u4q9biBjaLpcSamsgd1OY8w+qeZl28sYAg
qykfDYkuAI1LVfKTRhWKn2BCGfZJO08F7EX408oA5ZPeMtCv2nPDNEkkhPujY1DfH5WiGkYGs+/X
p0h2PBBDSDbhzKsNUH0S+9Oi+Hn1m/Gi4V5/MWQJmI6vdsMj+vPd5dtNCV++N32x9FuvBFpRYWUO
v2hdyPGQnXVyKqSKEgLCkgSndYC/InJV/bURxuVt/SQe7dLzHuFpeQjyfIhJrZ3BLOJMBWN63zOS
F3vpcla0aAvnVGwtQ8zUR0v3N3NMCCj4PJnwQE5i4b2bmYDjJgu5zvO83+enciD2CI+KgOvTwijP
AYiYYnWTcDW0sp7UPwbyjPjgeKxfjTYIWGV0QQJFU3UZBmdiqWV7Lh8sKKLaY/H6IAVSTR6tDXnj
N+xPHzokN4Im6m3Y+IPQFqEczoC+jL8tcH7QTJFsK8IpbAmTUrv+Y4UROIOmMkYCqjZqb2TrnEbS
PiEj3Qm9PmC+x1wjpNVDsEJUfl6+WSO09SFa/GFkJzP/F0zUAUejuBA/gjE9XLU0Nf5IH6HWySD6
gRbQl8d603drTZnD8Ha8zBbgt5S7sjjdRpe40clFuTmwA/OFLveG7BGL3r+KsiKvWsXhyaCXkvDI
JLVof4B+/5rKMzPcFpYFPsvlTPZpUZws+mThO25OdyL5jsb/B13Br4TK7XpBP0SxX9PRbYQdiPQ3
gbknoVi0YZVyx4VSqcVIP1aD18j225AzBj3ZsvInKPLS4JsA1zhjb+Qo0zX/z1RZ1NRvxkKqHmk7
Xkhkt9mIn5R5MfbWrkzPRLIvhLN6AXsmgY5fdFjKd0+mo5IRuwuPCnF+0qxWVWQoOo8as3l8oNTU
Lb5f+5kU1vgDYN4+PhDrJH4oVcxxGm2iEk25MNRP/H1DoR00JDGMFZCeMCD1Ylc8XWMKytouti0t
Bj/s/BaadjwEsDLHvGkx6fHzDH6UMoOSpNxIXr4Yvhm5SuhMQqEpbKr80ijD/mscu50f4StYAgbp
ge+FTF3urLVad9KPS5QDrAPwndQI+kEx50mYsmPoJ6+UJlkISWjurK2WmsIc7ssvnT4fOK7/VjD3
PcnALPzbU1QPPpE7DgmHh4BvINFzLA3YsgIiWBWipIqYeqWetbaddeLl/Z7DhNima0e5+AyeUB28
DFzFDuymrx3K3m51b92O4KKlj1SmcUqTIC+9Bk36MB89Fc6VMsZAZXfPsigVjn7pFMxHC2qv5LmJ
ufZoIo97J3ta8aDm8LFQj7rdBBjElkOsw5dyEsjm7y60Ryo0lG72lQn/doZEkbUjcnndI84e6J3b
99TVCPubefuZ1PlCAR1IOzC6rthlLH6z+YUX84Mo+LVbX5bgw/vRazyBOgHglrAEpxUeXjsWl7EX
nmZLpKIbtjQF685rcyL2l3iUpFLsP9MyxS4enJNan7aLEnmuuzfjSEXM7dMxdAyGBanEmnymb3Vs
/OJxL2l0sBDzYOqYCoqnk+Bpqve8hID7eNNc9eqTiP593gdeMnuHVRVuMu+WoU7vgqoC8lAOgUKt
k1AnRs0hdUFqWkdStOyslBt5v3uPTJMMuxBwR4Nfr/xJCOhxgNKutqg5m6J+5Z2N23L8dl8Z2L1h
mladphZT8fZRcznVelv8/l5rW6CEwOZHc1m971krv19TWuIoQTK6siWXX5kEY3uOsLcEDBWfyFik
kE8PEqyuq/UkPx0Tv6fkrqksAhKRVx4hk4XztNe3eDzXJE5eKYno0ZHsz4ENRz53FsV/r0MBNvvh
73ls3GYaGGBmtwUmGtVxJAgQlyIzPfQXPhYkKbNFtZmLVaxrWWZCEJq0OmutBnntu7vb56LPAT1B
S1mEhlkLq9ds3Tkn5RdUYkp05D2e0HYZvhS/aVUtpRW8awS+kAzbrRR9Ucw7+nNeOdPt0PxQzPeU
Wma/GSfG0jAi6XkS4SCVbt8zX/EiPDKPgsbotCo22S1vlWCoUcXTj+9A8DJ3sq8kPyw+le4Wxulw
SvemklOhuF03qWfhXeUm0Z8I0FoQK2/KOqoOdzYAwkuTCvJts3nitIT3KO8ewRb7eCh8VrJTx4B5
PVrh7YVKtxCEa4W1g5JaMKn7CyHE7SsyW0VrBrfzr0ColZtObvG2k7VZ2wVPuEe7qvcJjerIpV3j
NleaNJS/yqj8S9qDUjmf1jvhDCv6teUk/v1fpVvseQ10+GXM8w3FSf54OQcV9i0vJ4SW1MkDjjcV
1oMDfKIDNo2zzh4sKXx8a6lEhUidSpumzgzlHAwHS8t3mj9dRVhFyZYjazE3XziiHxVWy+xIr50P
tc1dSxD92Zovy1qLEMozY2MLxDbuzYq5yGgdE3YBX7UuTq2zAxJGJUD1ZVTQQuBkz37l0Rc+X7PZ
xOlGh3c1ajA4DF2sHj3EkBC6BipbRe20PoHhXsl+/mLo/HgNQbLxmqdACNXSdZOS7fwUkKPnodPj
DuFs7fsji05fXhgbeDDYubSmpp9lVaLBEukleU5rT+5GalpeOsZilvLlxe4xKnD6gtls6NRu0hAb
+aq+PLyuTOMV0QALSGB6baTfeZcpCPpUBu6DpKFewWubrXL7vrNNU50hUPXFg2Z9rutxajf7ZSaw
c94bK5AUHU2oUbzvcICycH2J0ol3Oqpwyv4AYVbazujcAFSNKQ0agWbvAazmqeMST+3kEmK4gzpi
YEa7Hg1FB81pPBCOFa5+2PHyLDGuOX4EcMzB0VWD9gdfXMRLVBoKBWXls2Od6yxg+HQ7+KelS8e4
8esSe6vkUflwmd6+95MyButlPp4tmccXqGXgcS4JvazzS4BJCu7Jn9KigxvWJZ1/eIednrm01VS4
yqZizs46LhWW1CV/WBFKgHr46ZoyIhGGQdWwx07AGXhmt3JyT2jiU5BVsFUWfYwvkErhypahSUxF
DIFWIOgpc+W4GFtHAzbRE0HdNrCNQ/rDBuCb00vAFLIdyMhIe34A0V0Me+7KSec0rxvTI/VLOF61
yL+fw1jdBvUbpGeXBhAk6sa5LApzn7YCubCq/zbSv2luuDKlfWZo8oGTiLpYdf7ieQI/gwq+PC/X
RDoJ5dZgsDoK9ISR2jwTmi6dcNFku9rrWrSxufDC+tKZ9y8XcGHTBuypmDZYOn3rA/RRuCDXkuRu
VlrdDB/zGTJbFVYdb09CjZid671nnJmAdatNwqP6ngkGyJLqlYdKaXcY63ptvo8ieDprw4bdHvRK
uSCB3dCRVNAcEU4wzli+QLQGhcK+fOjSO7VUHuhXsJ8Nnc9nTWA0Yu3BfpzhS2/xJT4XPS43U6Q9
Fszim4jbik3haVXA1vVfCccV1G+jSDfW7rbUr7u2FGWPKIjYZdrxZLFXukQ9/9dpnzmxqJoBLj3S
HharELgI/NLSrM4j2XduuiPtuVGLwTbcBNOwYeZSQBiG636GPROekWT1Ey42PRzGx6O0jGAqDTwG
a8RvgpByiESa0nBZBggrn+YXM4SZOP/cArYcfXC44ptB9UB2p0O9nLnDmWWzkSLjkSIwz/af1TXn
oGF1LRPVYhYwRGGY2foqmawBR3qf4YMbSto90/e5OvBqmxx8QllvuC29Ysg+PcglWSh7F3+ffIh7
fZEDGOoFSIoi3sdijG1r0zym3fhUdb24zSXvjhykfEW5uQ6lfb32g4P/CuBE2ctlnnxIufzGPayI
0paQ3K/TNeg0qs8SydbAb75hhTZCODmG5qgW0UjUSgo4bhMNeAtEARzl31PiVlD72aWxbO3bP7/z
BxKJ9Y3S/Zvsl87zutgMa6p6gu3z1tSYh74sitUxpqUOgGhvj1UW7mn5E0QtyXn8ZxM6/PF7GEsQ
5cT3Z9QkvGBHI0gi0Ml+VphdpF1Pa0Esj026iyBb3wiZpfOZT+8WjNWIfZOCM9UWn2XP90jque6G
1pNg39mJgde1uUBNE7/RSWW8C9CpcNZ2QrHYaGB8qA1r9FDWfNivgIPmlP1A5EzRIL4e0YWPtCpL
O3t3U3KbVbDeKwvKar8DFaUhAfeMjtrLQZ1qmMc3RArktiUw1WSoPQECE0Sg3ECL1b/AzP5BxcEv
WZRunAi4mmmlyYZ75uO7lf0eTqUrvlRnNkixyPKYuRDzHr2r5zpM8TpIJfoEQE1173AXKT47YZRA
Rpydq4/nXhcuTIrm1jmc6y9vy1p7ep6j2pOBTYkhxUcZ8sq8LiJg5ZiQJTsIuINOAJ7yd1p1M8xU
P+BETcJqXg0BUexL1qvSDmR8iR5HDU2M3I+6A3HrM/msQdXR6WH1NtiZ9ipRaxJNAC5B+qul96hW
rR+e3UptvmyKllxJ8eU/pOUy7VTdcbyFZ4hPkyu/KifNlHL/D7dXzbYqEG2izsNxPiAxJUXcdjDl
RZx6Wiuj4ex+VyA57P3IpZiSowudrq/pUITabzgTyVJUJWE59OSj9Nm1YOHHUH4hlUM0VL3kQdfg
sP3A5TyKj/nWhKoFjx6HhyeW50zQ9MiXZNWP5jgcuhu/zrIe44CmVtMBY7eJP0VAoxq5fgl93LbF
8Ga1MA93JwB5Y7RFCQfGlPkkf7IN+4L0LdQKqVKKf3e//BOu63+/IafbfSMu5ncwQ3fPYiGRil6P
EZgrh+VEKPieUuqyaD4NUcxbFzJAbGEfC9yZJnfXbUUKN9WO9AoA8IoXGfM+nexy6bZQySrFpHLw
geleSds2LTMjOrVsuWvcQyHGNOOkHug34Q0I9BrNWLHyOwnr0kxlANuj1w8egs2bsJ4ZJewI4/Ms
v78E7517n0mSG2efM6k92LD0DQ7MuuFtz/1Wi2tKqBAcA5geMtufYDwsgHING5PXAW+NRS0fixNB
/ZVhFFHUU1aArvut9Zqo5aXB9pR1QRBWSxq2F1dGcDCTuFZ2wW/Hphuq71eEtv/1xnzlWVMhfpnQ
ihSd4vbJpBmHj65IqwdTHeF1X+SPW/1C0GlWsJyEqDdroG6umobO4kw62FWxtCpW0FvyKELLp62r
uB7qQTEZ2rb99U01lKBQ8MM4Ksxu5r20PI68LBYqwCpfszzT+oXQZjO3pTOuGiqWswoYYnD0kGRu
8iJJid7esOtl8KP2EQiBIEk13FLLFggWW8uwPrEOK/K0kASE6PU7wLbAHX01aOcTfv4Z8Q1F4H+q
nsTrKRJB4wamTImvFzcC5ZDLEmCoa0gUgj35RVYD/BhN2CsTth88VVpmHblhylEPA7EDMPaS941K
DnQ4zeBwoFm861bOuzadu+RoIUmGzBS/e6ATKmUYBq+Zen3k31AAYCBhsmWwwd9FT1SnDDvz3vAI
5i3CK4rgTIdZS/Zs8uD0KWu4sSQhP0fzR1loCTwWFzJ3GVk0g7C7jJj1EXdzFOCC2IhRJntKo2jQ
aXyS2AiPyr4B3AqX8QvjQ2hBO/2nyRGY7dYSpU0qWU7scU1aNkjAoHEKifdA7aQNCAyc+/OAucLz
EPqySjYRlqbkN9ihI+EljruwcfNuJJQNshxXOrstOzbSkvnomxKhytsV6kg1zW7nT5NtNHuaASWa
TPxvDzFgib7Q4e0aApxZZQp90wwksBfZmdUJvJPTyXYa+HEDNEiHLEvNkgNLDF16Qn0rn9srmT9+
W7WTZ7CPF1xaD0ZD8PntVLKJGFAr1dlmZuosjUeGt8wxE1oQ8ML+cn56d/xOGztANUxcjiJ/jXDK
ULtZJFnR+z/+Q1hXqs/hSH+Ymz0wBIles7sN3gU9mjBkqahHFD3HsAIuemrvthTvUU0mhI8LwUgs
gWo+kjCL85KO+QzQGAr7Vku8oWv8LdHQ38B5+BAG9Bbssw8hRpgoEIr10/Y5+5tyHnSBRxkumfk0
TgRaV+gHfnnr7AJnrMbOT8nAjP9VHzKpMnUCpMimhHLiEIm/GqeDcrQ/7SsLpDgHbBDolhu6kgVk
EarEkVQBUjJStaFAQFdTofYfqQpzBYl/k4a2siVHv+DHVqSBSl4Whp5f51UNzdvEWE2QjyNYZjpq
qjyaXL/GasAgkxl/mZJhjnx4D0FAz5ek2hONrn5IfBV2tWR5iUrgfxBzeQ7hqAPYcSb6VA7Kt8Gh
GKKdbJ+/DnTV8gGXZAiXO0DBuoPOI+froBvkynpOIoSyjVSrv2s9CY+MtSEtp/YuV3gBr6g9j/9d
g5uKvnJGf3Uth8nAyO8YZShEHnivoo90TBRz5s7rN1Uhll5gdHvpJfZeqEu6+qK7OINFQHUegIsE
h4fi5BhagwJb31oeyoYUTN8CJzCsHauyVgZZn4ybJevnE3KThm2XR74jV0FsfteHooSC2f/OA/b1
v9INg6/SoXhcGwPJNQpkoiRju6P9NLbG2sR388/0bMway4VWIfxRUpsb02W8z2mMnyuXZEu5MrCq
z3MIoPURcd/wGGP65sc3vW6fixePKDo6M5TN550rZPx6s2FFkS3oCq2M31jWHOViopBoYLVMVawr
XG5JOF4UuPN3TspaIr9uk8KgCAGQZDQO6pWnLDr810uZ/49gjqrkoJY34GSLehepDevG5EXg2FmV
AT4WJ8udrJhxb/kVkcc/6tTiIRyHkFs4nq9fiRAAolqPKHIUno6l9zbve97m1+YHX1lPjpgGKdhv
eKoO/eo7xCCRu7nMudVQi+ZJ4YIxMjOZPCGf6R8WmrE0jm4pEL690fKnsl09F/NDW6wBBXudFujB
HaOVw0WHVy0uZ8H6irhxHauobZdajnc+/qDlGaZtlxtyZ7HUna/U1iUZTV/7Mo9nxBPRDx0vZB87
CSXqvbljzMwzNQRa4TU8lbeCSSaRKeGT+fRlnxrj7gqA1QzMP8VGePpRo4oWfYAlb9Itvz7qCWMc
QVmxk/avEYjavGsMmndGc/LjPa+wgguCPMIzNVJ9kOxx45WyHrpx3Jt9jfhwdiJpWjTwWZesaZVg
gdzgMKSPKiIlHZPy0pr0gZEUoh8giiEK6R3nYLY2eWo9MM2CxHRDOqMirSjIsnvWdzCYJNz4nBVo
jgwN8zmwfyPd+J5A/lxU0rwXLx07fjZ7Ngrsle5czyqeTyct6MtdUPE1jURJXszZXMANByWUXqaz
xFuT1sdq8OBtt7QWnmIsr6I7puLtcy2GN8PG7XcshUYpgRZ6GHVnpz1aUPekTR9aWSpVGIEVuLLE
2+zqpSPcser0dwlGYFASyLBdCXiIgSW0HM94zSjr3qjHyB4fL/Wl6sE6hti0PNY95d+UVSWimNGe
9ZpAWjSMSRuLf0GFcy6E7shWBXhKVOA155NPUUvZawVhIg2vrdYM7tTK6AtkI0tsCmCj+54pnx0+
xFy+6/wkP99m11JSg22kcwkpGxdnPhBAw3/S9j+cNi4E02/FTKcY2DweIUbtaFSETeKh8IZ7Eddd
+OYx3PmhUZPLTPVQSwDhpa/GYqzUVtS/PTigAy+/6I3zXvOlSggVc4P8pva6eQdDP1mSOHCoIx0B
HBIfZQgq42akLlmR5vMSrmI38mRhgYjRgxHEd86iQNoxHtSVCH03NJHN00lC32hi0geJsu+TjZ58
GcLM2DMPK8m+fg4CysJeLhxg+qRVCWC2AZRAFB2tWLiPt2kUMpg+V66vrDxgc6XLbXqIw6G0dWD0
p/vfBRu7x8lkKBZDRN1fcvje05z+lrhwTG3Ed71Sob8OQ0z/zysGDeggjMS739YCJ/DrSdYwzopl
q9I9mh1NVt1ddmXVv4F8PgdFSqmxBMl+d6BEbmXJNfopE41cH0SoZClgWznOFsmzkJGjkDi0aHGr
t2m6nbbjJor/yvdq9n+gX8VJ9T2YBEOeyyeY4N+w7ucsJnHfXPNqonfCa0I05LeiUAkyFugGyKbT
DISbLCUAgJI2WDQ7u+dZI1atRkDFcg4DBzUDFK6ZMxRRc3DEVUulKuyoHb2XBriWoZLtlrL2DQ0j
WmDomh4FOWc1NdPY5IXxJCTvE7y9AKELnJXGuAusDLIKmdkWwvs1dqeGdTfNUAT0/ae+ntZqOW+6
c0DUpeIi4D6AI9q94IcsSPnqdKAUNXoJd0yIAW3wxH9y5LJbbPt/DhgALVg99oa//4kvjNFoSOZY
Xh+nt0QmLns1S5sSbCEMD/TTartNWN7sBaLcvSKNRqYl6GelJiHGWJxyh3M2Iwp2b4gVcmtIhvA4
VMAKF+aCWyGwW/joVIE45Eq6SN1knmKI0qUBaxtIG7i7wNzYdNa4sOSpoA0Fl65ifwsIAltO7zyW
k8SiHpUrJAslNAyvAlTrzQIvXoTgpcj9xAKWbbsoJ0JCSZWr6F7bEW7HGdZ9d8ReXAYIPTcpRy0J
6JNhhiS/3cke78iAqjKiw+3Q0MMzCCk4onbK8wkRyu73FeH7PN0/0EcKXKyqOBLk6f14HSRv6xNJ
w5kJUrx+JvHWte9VWy6NjzWEf0cPFp+kIfAip8xJqyMPjtF3l2Nqh7ebtNiM05a1nfHuHnVzoz+D
D94ExKzpFiGLiatpYAZAOiAUTfgAx/4LnNUgSx6jkyjxiTcFwkvRX1uUVwvUY4bv0yxKokdY4Jt+
J2XtVJkAEe7TtHqWI8SQ3W7s5QZLIW98mAOTkSmx1CW8BR24srSlL/HXSjgpsRxDR7aZTwOMNNmr
t3XmZfD7QHQjiM4wPCzfxytZZrAj2GR3ho0b0ReWy947/oRFRHGBulwoMX0RKULGARF44hxmf0ZC
ADVfEwXZd00hCf8C19Spm+ZuWvXhvtxPR/92QOMWHvxtBOL9ImH8ykT7KVYQDf0Z8UtQ0thNyTXw
MSZYM7bSViiMoA7rIQ6qtUjNQzX5N7TCGuFFWg0/VeJpoiJH0OyxIOsw2vgkgdPV+djboHFhSuJ1
LhKS2bqHEkln9LmzuDU5AS42t4TV2SOUs9WCiV0uKr+DTnMckUc7YHSK1MccEIi5W1Rh7QONZNWS
2Lt9NeiPJBiw64oFtLW8y1cghiXgAvJ56zN1BWQ8aA5geN/aE6aTsaYZ4S92m4epnl9e6LxG3VeL
30KZvotnEB8uq8MM9sMKI1nfn6EbUDTB0QKyFtwF4cIYWeXiJjgRPf/xNB6fn3NyCxB0a/ahe7dM
+5lAZ7WC7+VzSyMU/O7dGMCVY3In60qASTVOosz3Ev1W7VluNcxcjz0B+8OhiLyV4GcqipPmClrO
DevrQouoPBZPRv0QifqfsPIUiwKxey2L4MY1NRtPUJjaDma7wMO4NwslWt9+UT3xFGll9r3gwNiH
AVmBegkz4SZmsJiq5I/VieYrX56DiMR/ZwT/eSyRPLTA3dPi1JOLWXo4wvUqPQb4Kyyxgz4hEJhw
Tb7N6IhDOgFgTGDnL5oQmec6/wmYVGfIW1Iq8xXJg1zyVdUAjFJnQq1MSKZ/EqOcbWh9KCm4KpY8
+BTACJyyPih+wXUsUslH0n+7XAyWNRq4B9mTptTykopZ7BBXINcG7qWvr2OTJygXC8pfuKdIDv/V
++1ZX8NwsZR/4oamROgBOGxcc7Na1+e30dAZ2LA3373acPNJH1YbOs3knqvmig5hQeJVo5620SF2
uhp4p9850GbeMFG1tDYFTaUhEBkGuNmu5RG/jZ+JC9HxdiqNWdSlw5QRNjwFVrJ1KMrxAj5kCep5
RU+IYJfAz4R573OFWgYE3WydO8z/7+0BaC3gK6HyU7Jgfcz0zawR3KMbxCaQjNm5S72+0cTvImlk
ngkCqBXtOeSGrSpnqOn3mt3BXAN1AM3up/ziurMMwqVYVPGfBXbcoonWtlVMjzh7LD0jx2oCYas6
75Pn5nGbuKH5PHqXvA0kg03AmuE/qML0Ac1EkaOlj7dUWfrr4JtEMc9IO6yEsKh0RYK58cm4thBt
WaiPjiYzvATQdGcoBGqWUMcspEGaSvRVROJvEhV+LOEtcYV4SFXg+juOlKQNy3YIxXTBaAUSm2lp
k9nYVJ9UxKI7aej+QY2tELG7rMe1p3qYemmACLsdgLwJuGpCA5axzEbDiD6KxoEyU5Ea3bbaOu8A
if6zSekN76WAkR6bATeqLk06HyWm9XX8TGxwcADX3K2NXngGcaQuFipBs1eI3qJ6Zl7iRfNwJAC/
0MrOwT8ZzxChexitXoVpRm+7VAp18NomTVGDUe3Tvqvp2yi+2AeerKcmho8q0IMqerLB2qsFnhNN
yU8U8ZJtngRDdV4kgU3thmyguNd88PeNeKU/jt9TJFYKDnqZi0r30WBzC56r2cPZ+lMQKKhS9u35
H4Ylo3GYxGtnJ9sZ/uO/1Z3tP1zDkcujrojV7lhaIaRsjvjMY3M1eP8rXTNRSm2Rmevu/VCzw/ky
SXbm0PQ87koWsYE9oWPrNfvqS0AkESxc6B3eYqgXSYMaICP2TqRsBZOa4/Iu+wXaq4p/TraGPNqi
IsO4lmfDq53rxpJW2rw6bQ/nyzSwejdwGSZYkUlr8xUSTSBz+3RuyEIVa/D6Cp1tXWQW+Ezo4Yh/
nxqUs64vfUT/jDztWOWbyn5IwHsV8Tq/qf5GWIY75DjOhs/OIOi2wpRG3gP/cQrew8p0QqWrBSQy
EQ8bcFzOVKA5d5U/H13iuxG6Jml5oIQSqM1Qyl2gQYzwKkmZVS/grX1ChzzywiiDbu93L0bywpem
OOzA73EkSLFOfyUh78GVEcENltaZ+3ZEN3b5i+qNPOgb9JTPXhoIETP6T/EjnpALBai8DppuDu41
OTx7N+HTOM+wKTafTVfCVJxcGLSF2Co785kQzxAKyaJgTnCki2HPleisiSOEgdYwWPn2loLZH958
nOSK6viH52eCP3WrDW+ZHaTRvySR8PrQP4DkM/FUx/t7GvYDKa16I7Zxh1Zpe8WEgyzzKZQ8yKVj
bdJtfBooaVS+W+Tmb9jP7bgTJWCcZjpSG5hSb5oZSToILNdUtmWzTKwVf7Gkr/3Sr8O4VEVK2zpR
ZF70G6GqxeA5aXVC5oY2Kd5BwxcPM1LoColLLthwxC0wRMOO07j7qPO4/j8aF1Df9QfxpVThCEcK
7mdR3ZwEH5rHBNECN6HGQ3ql09ylEWhtY8rEAMlKSMSGohjGTdDonpDVRIcHnRY3zLrBvhspkBs3
Zu5rZViaccyseQBElDEmbM2WRD5XTl7MXbylmriLk+O3kne4J+pFVKmKWzC3L96iumeqwML97yUr
5wBUyB/0H9ijxtPUbksuswdYpl3T+M1qmKXlcuta6AgCeHnOXCR7reI4xmn96wW4PxDvuDGtfErB
CH0mGPrE7rxxlZ5LRJtNAvJfkvuvT0adg7gB/OL8da/H3OtymYJcEgsoAyp1TufVUYdLoFWC+4bA
c0kecUW3vW4vQe4EVoqOJd7/AVNIJ+8SQH+86D0P43ijAz6tlYWjkrAt8kb6vhUlmb0gFtbRCvGF
h2s5Epr6zGvk2C2hrKU4ajD90OpOLPAMt5G2xeyCIxsDgJKJFc2qlfInw02HTGKwNvvlF6gOySXO
KfQOvGSgRAdbOPjAlybDjV6wJPFWVfxLwJ6issUHWUsJlNrPYyNSKAuhxw4KnA4Acc/AgS/puamw
7nEI4B2mGm/JF8eXFG/dxtzmh5s3NKU11QzXBhcpEsUUOoc204iRLblcMe9WRCDca/m4/164P9XS
Tcbfnw3pkhVtegOC+cgbJVsGS9Y28olYUVT/GRcHP4A/II0UtugW1zjY64INvOgKmkWzKp3Lus2T
M6qFpe+MrxzES5e4D8OWhivaWFJYvbDpMztkvXh4/JU/DzGZoOZEAV/6OvgObWEO56F7A0dnhE4L
GwVInvU4fCFo2yCd1K9djH8WTmjxEZDZfY2+lsLkhSS4Q35uY1RKv3P/j/wd5+0tetSxhFcDdHDs
l/rfJcdhq8DTamSMPciZVzeMWbOMNPY5psmodl66/B+Abcd+6G6k5AMUMO+aGzlE1Zz6Z7ut6Bic
BP5V+EARwHgGweSY/fwfb9Z2Szqe1REe+Sqn8stesQzSocUQnriMq11PVesx8lvd7n/3TkDeCLFb
25HojkRBV7eFuc3Z0affICV9QYGtsDoAM+uOGtuOk9mRBCAWkzE1pWRpvzUJ4zq8SHqkwbx60EYQ
DgsGfoCna3wZpGTRFIkNP2JWnodrfMRECUd2jNk2D+ouTmn2ZDw3hlpwtf7iC3Qxd6DfCdczOTDp
8/1Z+R8VpGpubjN0jxwSe6L0TzwJpKX2Hx6V20GuMd29v88VrkJ5o90aeFWGG4gwwVNNNpGWiyL6
moAtL0tVTUzSzSCI3hbCF68OdaUW9fGsoAIZvaYdpErxi+XVYSDpLg4s4n6Yc2ohb1YZEuz8EwoZ
MgDNPsM1cYf56nGmPNFkknccu3W1ZDqLoQHp16LSYOBZhqTMSYKrFyWNgWwjEhxqSqnjALvgt+RY
uNGNn5s7VHsH3JWaSWEMKxORfm0NAhSFD3+0iKrehlt1MGwmG6yiITCRiELuRrl7dW9uVDlMREX6
dsNdLNrOfPipCsttdhky+6LJo8sF3aLIUnQS/Ghgp7lISYdcZ2ZfuTd5UHSY0rzjrq7vxs9T/NCX
j7jC7YqcpQa7nVLgZOsT4285RteZ3f9DJk3/qPpMCeYueLoxrnZQyzaIL/CK95AU41j7yHZ5rT/e
ap66aYaQ3nr2rJEqBjMJsb/YoCLp6LpDQg/JeXwUuOzspxbx4WVAQTNviESJ9Rc3DJpiKVZno/W6
zbBa8gNNX1KL1AtoBnyK7u4l8bT+2ZtBB1IGKbH2S1bQ3bX+saRfOPCR7NQGlaWCTNUMqfU4+dTN
si+ogCjTTjq2PmAkVBX9KEeBEwN+OHGfSNPRiALGH7gDKTA3PdgzVZPIcCc1Zxt3pfZ3fw6MH+dj
wOHW3uPt8ii3o6/ybYJKMpfzz0YMip0IU5+UyGmvyToDXMKa6N7hVfy6ufS87TgjVnqNoZjgpIn+
8vk61OZ8wAbe1QxIOB5ylCKG4+J74CIFLsaLOfe+iwOMiwC7DlJG2RN6Q+xzAUAcHpzKhgH7RAk2
onyOZosoYIdWy41IaP2Y0PeoXXV+ZUyeruomGRT55H+UoZ0KwShsk21upfCZa5TOarS7YGhfrj5y
+OkXnBAlwsieYsXOYV4F3dDNaRAlP/oELxu8kjSaQpFpKcfBEHAI5Vz2xbQf7WsI6cF2bwCRmg5Q
QWwHIm2ys7OE/e66Q2uaX5u2DUyIcItBTxRZo2M/0X/xo8XJyOcLuUTKUeOKwiWfTr8ZfXQki4GS
0KO6rIxR/j9tvykSDXl8K7sWpbBDbBnjSclwcGx6JPMVq7NPrdVR6Ja8AClWGqLeEHU4kMP81TZn
qIwDGF29EFAmMl9LaX7qMzo1hEW/pi7v+kPe7W5MpgZRurhTVa5VYKOy+RadSGG1PFi4E0vbrz8G
qBvAkgOYR1biLD2YOuZSB83jY02BEl3QgcjZxhKEzQHRacmdSaaigKQTXONjatqI8gxYBaNyBXtW
4Jjiti/QgEu7+7t9/OSySBtBXjnPRfXvS0jigZ/9NdhCpBDHwwanYQ40wzA8Cd9DmPiyeaxuiYys
/hNGLo/d+z4GIUbacJuk5atymqs8F/B0mej/bJH38iMDi/mTUvl4GUgbnqgZhdxmONmAdagzPMVm
FscN7YEg2tIQ53Qpv48YBp8xwEOgwmGCS0uJpgw7zXeF+9CS/T5ZQPurl7vrXcpoRQx6VCPpxHud
XHLKIj2dynV3mdKWW9vy7mS1jaFduOUqt9UHFNJLRWAYzNCVfLC4D0kLfpYDhkrmr/fvlB1UIWqj
CPPtM32Tb6leaOcDe5pnQ0hcRE1sx0NhiVTDmz54mlJzYBTtv6gfx2XlIxpZbJ6DVyyXU7hMVIms
eQFiBWHFc/cGmS4UgEcMxIyXudIPci2HQk0e2EbGabLqBvKaQbITJdoKlUuXsxn7tvoTxXeOPtX4
eB5uQdd5Qs/+qj6vRx5uh9CxOIM3zcr/TrzjXTNluGRj68gynToHfGJdxSXKowsUMVPPUB+YBeKg
cP3vu9NrgBny8ZnjHC0hhCtFM1HhbEmeWhxFN+RETJyNNF50mjwoq0Ti3vq10whjNssQR8WbFSNj
FqpBrO+fIlk7lnuj3cWIfdYGA7f8bvh1U8dwS9hPSsJezWk0fmVcRemeZrWGNXB48dwYiM5nO+eB
VJFxhWII6PPcentFoeLYE+KbGghxj2UeN/G3M1e5bDLIrsAXIuLr22RJcoPU+1KOq5WwOs6pk3uq
Lm855OPB013dTJKn8ykLFyrj949tOqSRq2NxcJzGuOu2T8iHjuMxhUO9+4EBFpBRZM8EUrRHf2ay
fYKj8/1wkNsn+ZE49A3Pff4F2Grn4KgF7Gi0xGEH/6vU4EvwmDKD4+odrvNMMz9/dYXD0jwIr16N
A9wPbfuuXCqrJxrqyLo85HfOCuLb3DkWN6MI82oGGxF3pPrg2j5opd4zfJJc/4ra3NQAiWI1R3/1
T1rrIZpY+XfOCmx9VFCHw1MpXhrDXEcolDS03Sod1LyskYjOKDymdkM+LOiY71hp/wUO3OrBSo4p
JloyUHxVFIo4s9aLqzPkPc6EeasmjgCHRouTmlQlD4ki8rOkr4CaTnCE90XKYnfTgntcmHLt8UHD
Mi5XRLW0+x2zyDJ9L8wVKNbEOc6PD/ODh6NwGuJfssFbtQG8dH/SXg8oc93/UmkiFpVGzIyqnHAD
3o1COBBlxdoomPmYNq1lWDMHBRaRDQoa0p1ykPnXaplagKICRjmNsU9yOCb5jO7AAKt64RKuvRKl
CD+klAE/mvcskhpigvG+p8qL7WnXdYHreXga3p/0YzJWMp5SfTSUJsj6b49xgLL4NfrrtoQ1BQgC
cNfpM0SgI3r3sm+rygRfsOVU6Y5X6jjmw1vbGchr5y2PuoRNTQMQpFwoUnhudX2vSxCXi02gizS9
CYIPv271paCVekk6EPEshLjXd7ayNMwVB2Kyl5+flFiAekVU5ybDyLuv6jf6gK9xfMw8ORgY81xv
j7mjFMQ9fGOMCaItHkzDMxPz40eZ8e5+5l3zNx1bk//m9PGAPDO4gXE8/qkSACfoh3MdDMjJODwt
beLV0T5JQBI79vrqeNcnZqRYthucXrQTwx+MUg5qWG+l5QA+/tRiWz085VPMAhL+3ox7yAn4i8tb
LDGNK/Xx/K9xkXhJ8aOQmFxGoP2OE6GEjmF/2Rcg1+4gnyVJhWbPWshQ/SeXpiDe9+v2gI+1iS/A
jAl4+ToWzpSqEoCgTTiMTZH+v3wYoyWAJTPkbh5Wwgxe6kcGIoYallZ025q3XdgwvfroANDI7wYX
P6GIRSpgDG/1v7Je6mYYPXjVYiZ069y0D2amiBdiZ0XFafYh4T9IJoSwqC2tRk5QTVVYcsBiJONP
QL5ZFh5CX7kdriWjr7iyjrxTaBoKCz8abNN/4oFY8CxFpb9QpPT12sNX8VYu5E0OFSG0BCHn/Rjb
2YE9flXDFeXUY0+2ID9W55oIk/0+iMq9m/Q1ayx53qsnkU8M9KkfmbmKgr4gxjOH3Up7uWlU3E5Y
T9XidMtqbB/Kt+G6JoUiC0m+rZEVNQ435BCgVVsAyuRXD9rGfEsBDdLFUTJu3Jwe7W1FklZpUP3v
0RKPyvZHlTrCe8E0RhQU0ByOQUQIsgA7Qv4qD8dww/vMA3Uf9vSdND9xvrIfCBrPRGtZXuLrbObB
RO2bFDiJVAv/b4RLuyfQNvVw1MO9ToNxPJTg5hO+qzLEjS9nwA9jL0eTZbE03DGEyzx4Ml5+OZB4
y61zrGuZ1CtX0oRFe65KuMgevvIQwowh/vmbkSPL85rSrMvOH1buBpaZKo+AwI0rPPlGilMircdL
rEjDIddm3wKesc13WGXht+E97M4qJDkBMD3ID+427LB5foAaKUwJQIVgJFvU/OhZtfFfADhZuz9Q
Kw8RlyIR1Mp/kkzYXCgMjoH33M6XPr649USYjg+pNO2LQmKcMjwaWnsHwejGGaFEYZgOH5bK0jcH
qZlfWwNICbgYEJGw8tSuY0rBaZCFZTtbJZLzuhkGpv5oPiVekj5VkcLc0bZ7YPsLdMVt7JLw+wUr
sPklw9fJt1ksuBvIXKdthbAPFhL1AWTF1isMJz5BXXGiNwcm3P+53jqEFtgHyggqVJ0U6SZ/0Ns9
aGEUE+f880+5kyoUeL0UOe7rO0jYiCjKGQ3edIJHzK4jz3vwIb+kYzBtIUnX/oNQk4Q7WCxHxrIV
kl3HPV9qBwm9xanNRU9vmP09UPpqrLiSFBgMRYg1xqKUxYvaR5iOhJi5HvBApnJM76VQ+BzdRhC6
6zWgC5X5IMyoi3AOPN5f68v+6BeXRryVo23mZ/hT9i/bsWoeQ/cT/UZQnwjy7UVRHKRRYXYw7qqO
YXmMa7bDUUZmP7V3ixDkowkdDzRv3+I6RoWpQ4QUTks2CzKKZRVAnJzFdrc00hjzSnf7aLN0qc41
yVJOoxkEavvHsvrAqODOa6MrBxTFufq1am34sPmHbxYG0quXvdzsdh2Ih4IO5bXP72x8SoF9u+w8
h98btBpWm6k3v6Ry925o+P3KXXgfJ4UVadIJ5QvxKkFM3fxYIr6UREm94DNRJXZ7uD6DiePsvQe9
iOy7ANuUcUuBHYfJxtTtwsCdrdFpmW2B2zNmBRsuLEXlWBl5fRmdgBcwPuad6NCwCxCPI8jg5bcQ
m618oieYWECmB8JrhPd81Ey4yVk5ld1uI0U8ZLB3UX2cD8wEQjIBUeZZSV+dJrXO6pr2Xcumvdaq
SUDBr7yFvNGCN3G9GFFkk0hKjf8WJoJPGZ7QnRBqZmE61JGeif3ZhvhMnD0L6OkitmEpp/KLuu6f
PMfhAbZEFi9lPskaiJ7NDp3loeXSrhRuabLi46NE2DKB2lKLaTYc268sJ3ry4/2EKa4itNTO1drE
2s8z7lFqtYgV+ZbevFWKxDBU51ySj5OdBvqgeATylxQo7LNCMbDAfe+G/YchpwQ8goVzOfHPLVLU
Sf9cKPzvd86KgiidUXsAvps4OknSTfqDyE+JNIqcWSgfsM2CqzduaJ2m/JZGhcthzYsWmQoyQFb7
fsE/CBxeapsYNsig/+iBv+ysEKWrQxAjgA5L3sSjB1yLOAj1Vr4SopFzf/9xQp9By6mfutu5w8vq
XoJFvT/J1kmn3BPkXetFIfuq9GjDGlR2TKULyIkZRbA8YIX3h2T1USLsHvxEaGq4rl0gnqf1GWix
oXbUIZhnWaRlir8OiZA04/52fkayTcH6MNH8dHJt6iZ4LDG25lo93Ub7l+11rcKwGh6JNVqF+sIh
gGyOgEei8ye0kVYdnOasqtYIdfK8iuZJUomvvU6Ub8EB3dpV0d1WvANVMoQlyykIo65K7P2PxmaR
wrsb/zWq06Rz6p4xnNDyc0Ei2EhPAaI7B3ZWedu7MTEOzQFblX3TkDAdj79PKhO7O3BoGagFq4Up
uKQQ2EZMOyp1ax7ba/4o/X9K7CS+hBa3j+Kr31TYQ8YxGAqbJqG9l3+Kq7gllaEYz7x6TnXPIIXW
Y/TAm0JI0UAFJIuXqVvZGbYKpUL4es8NVYwJ1j55LNZgmsG2ddbtPhpzxyYlMmp0khUlGsJcurS8
JuRTZZ8ygTRW8SogvdQ5oTAQbdegM7tyV6e6E+MrN+0197PnrsDla11rhBZbkTCPdCR2UuR60hXF
uA/4Y1VerP9yB0+ECuATWhDJpFPerj1ZtcWzoWZUCcqeYCPJx1grads9MOEMCmP/aBvYZXnX/UUi
YwZ9OxxIvHGEl7wYvfAxVYTi/tWAgM2p7PHCOLrDDgjduDLWwYO9aCaPv63nF7GXYW/yTfzV0A2t
vKTONGQeE6DZiz/dZY1ugBcCjA+FdZHxb8cw7R32foq4uVS+AV4tD8iYNF+J1wMqa77ahv8xDGA7
RLTRZc3/s2lmJ+7yci/Uk84avgNF1V++3BFN9+Age3NI9Phsj+yfQDtI3CCtKPLfXQ5m8fCeX+b8
Z41Ai688zCSTu4479NTpsqoDSSgh8iKWH/MahRYM6ArPBxoXLbnWh6XbByP5YMwnohyZs95kFgWj
pQJJpura9MY8WdByqdFLeNTrvpDs0lZ+SgJovkYgWOUY/U2CPvy6eVzwHSeEbzcOqiFrCT60RHCK
E2u8fzjNGOu8/o5jNl82FP7XEBo8z700BxAlp5gKB7ZQRqg4fW9DfI+gAR2s/W9O7w9CoiIvo7ZP
hTgneGNcz8n4C1ns1E5I5sxR2DuvOQ3CoDQxoJHhq29isP3gSXvBJ2+Jb5CufdrJoQq5FISHpHOR
aKDBpi+zqDcIhcohxxB575sQhV6h+X03JNK80qAbFa+yw5WQjZQRhF0OGGOKPQ/LBd0J56Q1JcVO
/fe+rs4qvaYOH4yBoF5R2Rh6rEXnmApBA87yB8tog6T+fbuElyq2Kd32mf3wH1dfk1faMgGM3UhA
8LetbsrFF0M21ws4F4DZtrjUsXiE8gFgu8HrkyfEWKP4b66ITS4uLvZdZzqLR6Pay68rh56/k06f
liemMs1364ngMRS+7lC3nf8DnqxokHz1cjUNcsF4Ebi2trzMvKIbt38OGiQRu+WQJ9AlICqzS9CH
MN6pRhmr11RmRFs2wlQAg91NDTLcNwAheB7momTBFeOLmM/8zP3CZ3ldyLu9Jna+r/0jluxuOxWp
VmLun6I77MaOKoOO2N97KwmjqJ2tfd9MP7PvxAmwyshHNiz3uaAktKTwq5sc8Po5XlRj8G5iH1AC
0caNtfoqMEIcU0jHeeeKvNoq/iKkCG5ZZRD/4GmcQeeiIQP0fPwnWKoxcKUZddcpSQfl/OLBTjp6
W9I8iD439J/MwAAmJflk3Pi2BUe+pTlh72Fk7PG/SpWhJnQW5168J3xjn8lupHeMFMrB1TwEmT60
b+yMyHxLC/Dzo+dxcH1w2WQqUSfKAAuu5rg6+vQ1ByoUO7xbXQWEUj9sUxvOFRQf1UFsXyjkwI1f
mHzml4Zv9TDGGB8BLTcFdLQST7g2vpw8y3pOSsHF9YF+zx66tZKrraAJEZSCRABGD9lWXUYKiaY/
AVaHQ2zpSajI8Tl5q4xR3J2DuxC2rMEjFLaqUmLUkhOklT2tbTU3FsStnrh2MRt7QAAOv+bgV5jn
0SiX79QzBNVqr2BUGr+U2IxA5QCjXVtRGojiO5/RAabihHNb10dxFIK6q8s2lP5DaChRpz4MrDIm
uTwX2WpXDC5WWSvE5F8cOFBst05+at++XXVrzXAsk4oMM+qe/KYNQneNxvVN6PyxmYkYWlkAgdo6
kd3KcqqqKj0Veqma7+FuLmpvOxThfhaBA9tIf1ob6qDdSjZ6ZkB9M8GfJ7siRCgsy5CqfrEpgfF7
gCX/nEmaeMN4V7UsrfxXdnh/n+pNWLPnZp5Fta05XjD61evxb5u6cEnN7L6nVn6uYGGdp9XKo88I
m6cBsj7/1c/KPJEf++5jHgGkuUcvL6khm4H+OfZkDovRduVukjXrjdeHETO3FdlQbiUBsBl9Cd47
VS60sePVuYx8721gcvnBcEZQ+AYLXjQTMTV4n/0bBilhMprYi4OhVdB6zP0w5Kw8/e7dFZNgG+Zb
g7pLGjE776E50DoqJyFzCyk9XAzBjtys+IUFWEPRNzOZFypOnCWYqMca5IhSHUElYakbtJCNkweY
teDQPrTHpJi8fYs5NDGxEReG6ALM3YRhT77ukB03e0ZHU/ZYG6CAz9t+uv6ojcpl933q0sQ+vpaU
c7o76807TaQ7UosZmY0AnxRr++Zv8OayQ9pSS8bCRGeWnMWurjQFB9JDTRsQhJFMfaF89z/9YwN1
iHoCvQk0MOBLV4ubLGN42JIpou8JzSnXVRtAzEWNMeW6Ay2qUElIgkJAWL2gV8F4ineVRmFwvxff
sxeIrA7eJYnrsheZGaEtZDnH1+CsNOwfJ0y7wdDidH8912VAPeahcHrvQLZGCU/Kjni1/ejyzeL2
2OPJEE+cAZjmfMC9cE1BfTvZd92QJ8CHUj8UrWnIg41LwJNs7ISq19lk4eZFlGDpGe2Rp7Uzrt10
GMe2h/xO7wctlc9ziGFdK8zk+Mtq6mpWBtJAEeZhq0pPSqO7Xihigul2q0f45hZg+iKaQ8FUaqFY
CJT25NC8nxq0FbgdEIXoooY+Lkk+/1Bhh5mlGZpj8f2r+fDojwJMuZpW1mEwni3cxPXAy0JOyWEI
8SbxLpXecWjnZNJ9GeVqRa3HTlAR2/tNvJ4MtFdLLcc1qr8ROWcXPattQS1u/M75GFD5S8Tm7F6W
n171XT/Cg2whoEzaiam7uxGtD6wT7hEdl/xT2l60LJSCKc9AxPFtA4/IbY5xrTrJ3CDwdfDtjSST
RwvmauNBtK76VySEjNEoVVx4quiFPezMo0J7UiWYE6OZcgCpPYJFwNPYNa1nV/NJWG6BayF6SA90
AXYheM5+tBmpriqsGDcKYDlDJyutpYQCA4c1eBC+LKFR3F9LD1P0SAMjaYUlURkeDQTHyPcqIJKR
Wo1u+dRJT7n9+kylEUwPV9mZz9fozPrc8urE0xLzG+dJcBKv1TVuGYlRc7P1kyBcqbR26dqUFsiw
BWwWE2NPKs9pb1vI1rMfpx5zEhRrR2dCUjXFQcvtNirKapTkZri4NTYhjs800C2v8OXbzU432ZOm
Auf85BrZcoz6NQdk3zIl9iLMGj1PmH2QGzg+LQCu1k5Fmdi6KfQmQfL8yqAlXqQGtc0MOdVrsGri
uiL6msQMd2914qj9pOR4MuverO/8RA7EAMWpwgMthHCYNgouB7jwWrJzsffOApifzi+C+G48+hRc
+xFFExA3BfrpuXbbkukKjZZp7jZ0AUM2/YmiXJJvC4mEN203jsQsxFxlgrm0J2bphXDtc56gw6J4
fK3sDwMxv0gXAyuo1eZGG8jIr3R5WmiyFL3CK5hP5ZYK7wLorHS0vCFHUGWT5ZS/zr1eY/NZ8Q/l
W3/JNlx/qlsQRVdhCzX6+ICmoZdvgX63VOHjrFsxm/9Mh6IP8YEriG5OQxPf2jeJEZXEDogDqL+2
5dApEdV8GbM9qavUaFxvQtRnRUgZZPYke1fDN6XTDd/DlJ09DdQCOCDMhvdRmiGEDARgqKIeYuax
KwhxaQnxf6ouoZeunpWK8fPuRy3YOuhqxOWXuqItculsN+Q0HtVJPRmyZLYuzE98PueueU48Frbw
UPTadFOhPDzxGKq231gtCyUh1hvOWFf1kwBcx5yKNm2WLzQRz/kG4fw08gLg5MAlX9+/Ap1nxvFP
d06Kc/RLCYWyAbKMPLXsVIUKgeXclHxaYqCIJy5tXWzomizcL67MOvAWvqwM4lcZuEJ3MUDMNcCC
DeSmO9TRjhxr6vVQYXqTFtpngiqI56Wj2FtA/tLxpqgMQ2VmTudh3em3dVTP2C2yCivpBJtQeK4l
/8DPF2Pxcor3khg8+37/gWy1KAudY0t4k1wOPNV39KKhyOYdzXWcf0yER/2XHMs2CU5mGrzMYePO
WH/KYu/mdEBfxXxBYqVTWk4HP3ooJFoniAQIcfemy7g8tw7Rh1yndFRVcNG6Tk2O4CsDFkHhKEIw
8PySPy5cWIu95LzX/Ksme6u6jAwBXye5y4quvxskcsEgUfg2QCFwBAHYm00+yJSsMkkUpIAa44wm
9tMXY6Ili/HStqL3b4Sub6G3AxvAlvZAM10iLzyI2sxAMiUH4chtVtC+uUiySjmRKityww2QAa2V
da4/AQMeT2LlSbayEWk28SypdUDFRjp+4n8Y7t71pyx2mVzqkC9763BoUqheHuce8Gyd4K/BA2N4
uVD5vrxFj5OHo21whFnYqB8pJRxKXBAsGYbAAlUGVeI4mhVGoumOG1k/IodfBlpjAIfgglUdAS9C
pvATSraeeG7l5umoldOnlFTameX4mnEA8HTvSrHOPG8RQs2Bpw4z+y+hYHuRTQs5jSoTRENDckOE
ywuYM1eNdbtW1Sz+taScPCoQ32RQ64SpLjpKdSdZMqPJ6gKjwSVfEgIX6eC4SKKA7mIX4eZFRxSk
2U/BcmgeYUFf2mMGi96qpnZtUxaBftUl/rP2RGftlEGB+bTqpYtFxme7CksB2OkOCUGiBRrt7/bl
qrmebVa6zNC5Ot4F7j3kQr05Q+1Q73jBolJJbJuhMvqQeyidil4Iig8tkm1TfSI6YYmM2BekCufC
jXJehUsX+O9HBSWPGzAehhs1UW8GMtcRzt9i37HxXV90gSsK0y7A3uX5+TB6tbnREFQKTA2VZw/V
Qyxp8HjusgGpqbF4msHqahtu9xB6bcOvMsK2/AGIzv7CRcKKzkKUmvvjoJthv9KNgDVLloiWuVgQ
0dgdkBK00j/8B9GBke6OYkeWI2YDW6gRakWy1P7j/ig9RA48YomEsuaZiW5mhSPmWXZeKyBk+Xxz
iQLVsfqnIGtLj1AeFmssoWx5mPjOURRYB1GHKa1MOs7OIQWRlB/324KVYGFsm2sYmL+Rlw7s4cdH
Tpag+uWNH8TvjVBTfBwzLDVM3Bn43ZTtdYXYOrbBOMGxQjxx0I9Gqm/3T5ZsJiNbKA58bpnW4B+b
UrK7o9yuz5frAn/2CaFmTmhFpX3js2woOlfReXVK1HYhPuCTKLKzD04m7c0WYk84TgyP0ONpV5CM
vIFQpAF1jYcMiKkQVSw8yLCP09jFg6UWpnkFtv9Q7YEqol5mTtWnVtjemd9ET++dSY7bODUHexnA
Z5q6psEx9kOk7ncl2Mh0tBn8hW+Kz5iOpRA+pG+I4btqSr3//MfTWFSj/WI1CDoCSykhv9Q5wWqi
LcyyQI5sq8apDcOGJpi8oZeTq31awENAqcNzZijGSm8AIkYrVEwLu/NeuLOoE6nonH+uilvpDuyR
qTSRD27OrVFkgN2MqYn/bGUKmWvv6DQVXNhaD31NXu/pGNseQCofk9ognZaMLlWBO0Jipsw2NbYv
bxe12mpK5njEpy8H32JCDaaVIl/+RAV5iYbPMHaqyW4PHFiio7kTkqs61lPRRTH8+A6XvUD6R9g8
N/yCS+t/WtQeh4M+5k0bhPWfSn/H+G8/OcjohN0hB9fzSN0Sa0X4lNm+RIPgI81KzTXRyH9WRav9
2YILA6voZvRsmyctKTJwYywU6n2hpT1M7UIHdew5GYLRKu3qVa1ZhVN+S7f8JMRp2cZfknHexOIy
hzmMJ4LBhKvuPAi+A6ghULnTIFTgASQDiCxMSXJSsZEFOM12oTpBVYKP2s5Fg0jeyfpy6e9QLwrw
ddwNxg7MqaLEKgomUXo9FtYblPk8L/lOcBWPc0mK2GVs2wGOecBIrswQd8wHhUvHni377vLqC1UM
1PsDy2ZqsMiRvBwYIhLZXKvXB3iQ3hWSM/9ybA8Bmesddu5atNcgClEIMJPeOTTfu+DTHfzRcNW4
636xOiqC4vyQdwP+IcM+4vn6guyslKOSvG8xFfb3ldsZFjveAy/ptWG4Fqy18HoSjVtKSLQW2gDW
04/k4SfS70VsSUTUdQBcF7T4ZVu2Vng6O3PDdSeS664tWObksytQqgGK1nMdrVEM5rYpiVhZOljR
YdIGXfxMSUuTF8UPmV3UinXrXCZ0ZoX5jdHUyuYmxWknf4UGhXtSslmUc5X6xPEl2XHYy5sh3MkN
DXDoOFd33d/L+/veTJ5E8/WmktcO1wuP1qFkoDZLR58GNB98JdRNMhOn3yGDnna3FkL4MNqN4kB4
gKTWErpvzjyeF2+wAGTrv/FGeK3Uo5VTcXhH63djGCiJE+CbOX738vfkxn+kkg3xjLOVMrOrp7bH
xgF3r+Ny96nnNEMv3euU23Y4aZCxm9VW+jcalfvY8UdbqSvhFfgqiC8mN/oEMTd9rMRN0m4NnKIh
bj8/Lpyjs64gqnT6xdJ4lSYOpzyb2c2nDOCkwh/lbsIh5sE/Z5SB458ttdF2p9PbDP74S/3FZHaY
+mVJIwVHM77kG48xgPbG+yzoiVkHwC8RYHCiHoNsdX7vZrr5WDSO6CZDuNPNf8CSEOJrmOw5mSU+
a2sXYdXrbNtuwB6OieyMmAWTCQTlZ6eC5A2XJ/xK5n961c/g5phqWVyeThdmHzMhkei6aeJhQp3S
ZFgBo4rO4vMwVJCV00n9kxeeAPzciDylmAn+Erbl6XQCDLrvc16Pj0If2NLAGHnzF251m6MtFATp
ajex9PJibI3wPgECtjZ0MQp/Pdj668DTweI2Nnz7BZH8wxT/ofBI+torVVVhNJ0iCVfIvtjCEnyK
JrDgtjeuFHwPEX2cTvzb/AOC27Mo0beONgL8mP6NQT4sOlUWJVYuu5N4XwV/azQ++41mNQos2wzr
xkYGPE9z2a2Tv9O1qVsywMAgvDKenTiRW+2C2N9pontUGYFO+gvyi2tSMQsZQ/HtZ93rbuXEu5RR
89jbRcGAHk/p6abMALTtqrUi/AQO8Zu9r2G9ubEP5/3j2kdpXdOD/P01EIg61yrN05VUBhI8banA
k0T5i7Q3+EJRw2mSrGHQTiRjOdR4gd5Aa9j7eSxlFKhxlyl56WHnxrowatMpGQHNf12GekThy3p1
e4YveiFmopsbBJI9FSdZKvkqa9oSht6lGylPqnSfsPjIPGX9qbs2WGaNxs3q2LN1/3D1IMJN5HMB
TOlz7857Vrm7H1+tsmR7Qm0IczJLmc2nDYMnWcGMmNYU7ArMGx0/M7T2B1ndCO5gtC3eH/MJ78qY
4S24UT+tNsa3nVZlm06mFZPyGn7psUdGwkO4s8eQCy+RyGzQ4BtXFOS+ZPBHnA+5uSnk927G6zup
wzBdn6VG7Hm9v3Pflf0OKfhTZv1jbTaWVPpQO2GluOKl9tsZtEhsPEqmar4yFzH19bprSv+VJn+R
YQQNRHWHg/ir82pwHx6DQGGh6Sm9lAb7LwFLhoscwRFcLrA/VQYiw4cM3IV5epa8WF0ZXnTnA2OQ
xVyXqRMNZ6ybRVuc7PJxzQjN3+3RtoZkgVOXWvi/9W3Xo9DXzEuhj4a2/X7JBOttITrO2XPwSix0
JKziH/c6Bltkebevvq41TK0RD05QD9nVFEqNNRTKVPWEGeQrN97oBelMADEjoPbu9Tr5dHvBJzG1
aH2WHylGeO9czKmBgGHtg3oXIWtnat+DKZz1eMKRrLolA2vT7OqkptfMgfoN3nINLaVlpjEY/5RI
/TZPvIbVgXRdycCSXqd6HuorF/uB+ZlBAzJfaFjVI1q0W+8hYmmEx2dCf4xPEs3lIaY7viaOlw9Z
HwVPxtjjpxsOvvZGFCdIce6jDNLFSeRihY5UE+SKZwHRCDcm+/CvPUdJswZPeDWpfA3mMOp+gNMq
yINEYrGSz7W1Mi/6IigQ9SKjYCa+EcenACEwClNsK5DxrOJF6Fy50rDoOaGhMFr7q6obrJzQtDXE
Zh3PREvs4UqyMFeUebNlLR+3gKYMSaOWzHdz+eibY5Q+LbhTGeOg9YOLvNAtDbwzfatpVgGoLmJ7
dhuG7V+6wyMYt6xMvakTkyEPGA0yT4aN2332su7ssPgfc41QxHrsOBHJ3DQrcCSjJ+PMxMA0M9T3
Y0PfSH+aiAyvux1ugLQb6imQSJd/DIN0d8Xz4SGXpQKspevrMhl6de27ddG55hq8yIoraw2tDA9X
BmLI8ZFVC+ejSAfPQrw7x7PK2hXYU9qz/BXjQfm2LiGwsXTKUPDDa06b1OQBBrENLv9W8ZP8N+NO
u5hYxdHoWI/foxQJO+TGGXyL54rQUyauuK6CjDPqyRTW3t9z2vY6ROv6vQ0/TKMAZUmPPe70vTWu
aWNq4eZYhVYCMk3lRCIL5hh0UP18BVNRxmE8P+VkBZ4I6pJZRU82BjDJF50cAQmhiwWPi2dGFupG
SiElV6qya6vee4o3YGOKV7POQ8W1p9TGrpY3bEraj9zynoGBs2UnDTFvVz5A4HRX+c/IEh2fHvuU
6MzhTEkxy7lc7SHce6Sow+iz76MBEkCpxQdKXxmiyQaMYqbLHBRZfvl5qPYjszf54it86B1xT1q/
X5+no8R0kACAY3pYSQamZp/E4Jy/9c4rwSpmqlMp6g1wsjjAEeY3razasZUTyGv664TxxZCgEWzD
eRAD8AYTbXOPhUYZcqK/ouR7Ngx67nhHPxnW90PaiawPYtWm5RgraKiS4WR9n0COpXC7C0QBqSAL
RD4KY++1QSvyqFANPZCRLXmwFGtsFAAhNaDuoRTkfOBU8110Qwxs3vDG7onmj7eNo2w7t2y5Z3Wf
dCtNU0LF5Gy1QJnUMew02xfnHgQCEvIIsIGhyTG7cYeFlv9YnFMeobYqCuC8KyTY668Yiu+7xTb+
/YatDgq8kB9sTEHSwVCDtQ0lWjdTY4v5ze4i4wS1T/R3T9R8shdIRBieZvVpC7InGgzEvIXA+Mqh
KRFz2F7cn/7iIFYErjhZS3fl6rPQc0Yt233H2sPbuRyMniBXMk+YkU7LxGlkzE5KtXuth3ILzwV+
aQAMWEDsTFTuonnGbQlP6G330U5F1VxMsBzBx0M7fGmiEH7yBSQtAVP6q1pkvsgS0QGPbLc5K6PP
B6XC6l7bhzkljRQDxOA+cY3wOZg6BUaGySDyUEyYqdlkDFR9WffgU3ZHFv98xg4YwdWo8bcJZnQL
r6TTdxZBGtRQIENpj8AyaWvCE6DkbgHVqYnK9alPWIikCdMCFq8t3AMLzUknD8LkUXnfk2Jn0um2
qEHyHy9F9GNMdTeVxq5ICkiRLICXnjFBVaar87ES7odMK3CRXU1XSBc7rTnBEcNg9FiGKwVMV682
kxY7rkGpuO9gL+mhcNQ/tu/OTuCk8veK1JU2ETP3D8AU9+Q6NQKG8W+GJwTaTlnSqIsW2WOvAdp5
pdEeU+byJPCqFKGT1fcDDC0qHvNTte2pperaVxj1KfnArDcnZQejdD+vvX/w1pFLmON4fqvgBfQk
Jnl0vBeX6PKDQl7ZUrUNhWE1fCGEvPoll/N31s6330gYoFQFgn55DmuiAXi45jWpEyYL9wH84QXj
Yjo/1rJTkxsIrm2Drf87k6zlaN7LXj6RTzmLuUhQkJH42UBZHSHK2HrNDbZ77yuwawtNiSTzWxWE
y1CllD7s3FLgCL7c2JZYiurXov1pgZs7GYeFFm5p16EjJ/tvTrmO+EhOPFz8vTghedk/dvVslzaC
8wZI+LsObMSAIpyMBB4hhIX6uWaK9BfF3O8Fkkp1bV7ERua2PCVmjjWK5j7weQJ3zFMfG42E24AJ
zFuuJpdfl435QwOqK5aRNjKK1e3+HuRRVMP3PBzyUzyOmteMUAqEfFX6QHwC7KJBzZdnHw4K8a3A
Myqwloxi5Vf8P583tM37teSVa7o54dOOkM+n30wKmZGlDMsj6ht4zXDScWvy4AI4CA/94CiCVK+N
3W7pUAPjHAJMWr7OecrMHY19B2QppjHFSIDuZ7kDMz05T0YRrGz9c8uG4NmHiT5Pa+Z0XMjcABZR
ZM88Jf1oHuiIwcoszidRu4MxP07b8WY6ptivCXYWTEp1ZWXUPT6vGWXw9p4Q/TWpgtsPHP+A3lUw
hxhYAO7zXaSQoCpmghreE7E3zIZqmO/63H/JZbrlmrvkLtJvTygqSeRfZfDOcOxm5j1L5UnWYviE
5nkKfubnEFkOhE58Ro3F2J1e91Uu9CFmDZbtB1TJfZBhXmXhGcILitNlBCS30WwM3tMMX5Ivs9Nu
If7gt2wQXCj2Hph4DMTWnkFp6ZhNlx9SskLTYLy7PoXz2+3f4Ay0jXpaHlJPGG3M+YAZoQIkDVkh
VCk/uZHfOkFgAYcTvSmIW7DYOTvslow/geJyhq7WmvCrOx5dh8vXkRofWMOaaoYDfRuH+o8I2GKr
He4H8cd3fQhpu6dK/UDJLguXaH/IsQRf02poRNZBJ00nvCe+65yClnBhARmu8j8wM0dIvwT2mMJ5
ixQpcn/CkRjgolRSOHQPEIX5yryMOdArvbPHazcIlasSkqWEQ97MV/kUemtRwiKpGoxCrZGggYkC
cWJHPLSC9M5NYfQYVG7poSp9xWSepDKNlSUUljLCdhInXg+I4bzxh3SM35b7Jj/n53v+9u1TchdD
76HE0aLzQVDZY9ABU+J/zE29RAcKsQlkjF4MTMosftlf40dVF8dMAfUhQAPIuEug0QOOrarz+UnL
JkfTKYcvZCBzGEeoSAiNW+PrLMLIri5Qj+9M55OFXZx/D6DXssR+woQWTTYSwZij6Uc17Nx73gkS
ke9HwIfIY3XZU5xs4ctS2D27bqmUfX/nDoU/j8yZUnw2EviQgYYn3hrbgtRJtbUeYgwdlBLZXkiC
aqO2hY0ACDGz+4qow0G/hVq9JWO6yj3NQDtncPyOdotvayhTdgY6ThfgorMZomQ/ahPpprShhTbm
dcUEPNUiKEjEs1slEkX5GCqkM7ZR9jdEdRTXZprTk7VuCdlTXitxesCKna+ECSkvsiewVszrToqe
URSgHOBtvyGat6+KT2LAFERyTcycvnWo5a4oJHiqZUUxq/4MkLh4a4EUrg1E4/75qtoVqF85z8ml
I3Y6XZHZW+MWE5Kp+N75u4UdZdoTgQfrKs9uWc0CynBQ9DtPDfJCJoNhsiCjsAOfFUswN65ayt36
HM321lEkrCO8qIEkrE57dX5rejrWCsldnVI/lQ4Xt7bc3I6gR5lgC2VYQjXXQ6GAq6ulBbsyKSVt
Rn6WU4UjMgByCinXHviUaZTis0JbxqmR8kDoHgg/0zibUXDCJcEznLL3u3luKVE2nSzAAFlKmGTF
KqDGgpf2Bb5NkNbtHf84man7h0yRJJPf10hwYLYo65BD92nCzDfqDEu7rQy3w/CeZtuysPUD8txe
jrBg5xLMvIT4KWWBpFvl74WF6BNvAETs75REghs9eHXrRNqo3SWP9tOjzJJnbrs7JJ6qsLjUxB4B
raT5cj+nYjopVDW8dZ09I0c54hmXHLvaOlUj1izlm8TwWtxJ/fGvJc/fhUC9ER5Z78v1rx4rf20h
1kXp7AOGugUTli27K/55vacjaYlBvowynjOIFqtJ/dxwNiq8yhN71ccl8bHtz+ccIACynhvhWAxl
3TFSnHCxxsSxX/FQPpYtLDD0dv4W4f4m+Gnjc15rnjykNOPALC65zQRCCdfMAAGlAGS6BeGygRg2
Ca+rkl4uJeiABLBgm6Qz1EqM1+zSkqXtdzHwblYe8YStTPtpss4sm+nROpmP/XdkZ46/K9XnL4k2
Q5vTQtYaDRfvu1HHEhchsfXwfVWVe/VOAyfO1Me7W0SWgHQJdHcrcx5tqQX9STMkCGLtYb4J7qQv
Is0XfV/MG8rzHKuW546zoWZ/0lYTQk9AW3CVssnd3mjnioeJ0Z5Y01FDQ53yZJG1ywA83b3tb8kd
JHeG5fiGOS3XwkYaUczXnWZyDoWmbdN5Udv4nJhMKqFVRr+UBJl8mWAKsxEA7krHktbJNJyNHfqa
cXYoFzsCJ2hhK0MNiB9p4zX1iH9dHPJ+EU64qn/jbEjYSGsUAuNngI1iBqbaIW8U9aIReZXQ7iLh
kwQ9VKa7ujjC7hLte+3B8inh7qnZVjjUt53Y5GOvi4qPZk9S6E9hoUR5uqUAwuoddEGrUOR37Qkb
Put3WY9VxB6zWUxc/aNIMTM/OEaBQ0jf7ZELdAlRX2JCMifW7zjrZnwPakUsXuaLxgZ1YgtHHi/1
mhPv3FprAfr/zDucbJ/VNat0g6mGyPVPFPi2BMmXVme3+C2DoACmxyAxyCYaTfRsthQk/3JomUrV
5/m32qU0k/r09yjxgEmrJ2ZcVhyDSctptBxpp/PQOq8M2HlfD74wU2sZrnIyHc7CnRMluDMOYjrO
bucssWPkM++ul71FaXD7dFU3uHKqdgAyiRuw8/LjBjSbWQfxj+Y9K3/FFzxi2UATlBd99IZ09k06
Jf/hgtG8oPkBocA1Vqf8APDNu6ML2jFom2h6OFSP8xUECfOv7k2w/YhspTc8DHENsWMdq8dnOdrE
UEF2Gj6Rq8WUIcwc8748qZku891cWqPyrZ3RjYGQXQgibKPdgy0GzoejsvW0SIwm4ocbEUPMsTC/
oQUOJsq/HgGweO1RlwpceEpmBqSIYhhApfN2JzvMDISfV90m/M7CRZxdrqDKgsy2CgsY1QglLBNN
AhjzqjaOqRvl/qVvcn73XOLDAgAodze3O7j7oKhrz0A074Jb0YMqc0+yHVkvV50rNZfO0qehiAPL
pwtQNrmMQT2JiC0e9QzSlh2JAuOvmIrBUscEvea42ZatqmAQ0QaHN7/EKdsl1+dq3y9RVDhNMqx1
KRvq+XD34vZZPCMKEkqwM9KaB1/iWRpAjrKDJiGuGveVZy9R/4RXsvMGrHn1cq8ePhugdWsJWZUR
smaylbeAh2Zw6kQlQuruSPliUHXXzQplFdQYWGbLAkVNMaYMmvcAzktsGQRy9oQhLPTuPwN1rx+c
5njK7By9q8MxkgY2mcWC3UKDv8PcelNWtrmaaZRT85xZevD/dzmz1qroJHdYVCYCuTz6zhKP46RE
kq4FnvJ+YmMQdvTLtr+ipQamAtRlfsFnXtgQqONOPOEOWQqQIT8hrP+/+NaGf6l/m3edkakJlbiR
nJXtHc74OYIqT/5Lx6SkcxFF6SdwRevj0E39i0CdOx5YI645kaEQ4ZMC/nkwliwhCEqeyheAARzl
+4SilicHcLH+SbBVm+h8vWJ4W8sg/0TSubP4XmmdAxaA7IeUDdTA4i3SMXvPbQn1r1SfTNaQKeYE
fm+cVfLhHcN9PQ7WZsaw4H0bc23GMJB93uB5Rh5+IB3l5kXaG3E1cLm/hX1RTI0/FxXT1+X0Pjc8
DesImBYWPY+AGIL0piyvnh34AsupSMEvqUbwOtDTxd0SBLnRopJswSQgWYCY7WLT4u4h2m1aCWPq
eN/DqBgZjJZNCEa0HuR3oh/NpSWXyxgt+1DmevzRJmcafOEn6OtYslkY8UwvMoe3/pKuoLbejOdg
T7gIdxXO8WT+RjwCtVtJSLTXUfvp0c9TZRPmU//UnqpU2EosoTNWz1RyZb43jvBIzb/jR6PRB9uu
KByoQEWctI/U070PUnvgbnlE+VBjjYLiWDmjCEdu+mfd5g7mrYZqiEcPyPoiYE7ilftwtQ+h2gp4
KJYRWE46ka0M2cgPY2b4ku8/RxErLcum0mSN9nQGO/WfR/yLHZnn6h90nIfl8YhfEnwwi+sjcEBn
kzxDd/+JK98wHkzKbpbwpHcWO8sLq+AScjFq2CJ/2J7p4+nYSH6zTGvZxFbLAjv9iY1LDX5ZSbx5
JLAq/oJsKI2pSd4uuGyI2zB2jzV8hI+6XtdC3p1v1aXsKhQ+GIpwI8TJvpOYb+DmfTtDYT0iEJJN
d8LgK7hhF33Y/Uurw4carfkWnyIOmizNYpFwBkvcSFSFG0Dfk+IlpaS0UImGDYKfvoHSNC2bgjTk
lHmuqYiHtxj0Vqm8KeU8vEguTYyB2f83wvazk9mW4IiduktL57NAnjPWZExlHD6lv+p5/iq+8kqo
mXU1Rp8mFI3q9SfTpZx9Q2SCa11XOrt2yit/y28gmAb03sQUrsAhqxgqf+FuhcH3qpFJ7I9UN2Rn
9bhFr8EEQM4wkmIUOHg2DVtAlooUjjJWQ+22nRVM2ehSh5IRlVt1hsmkGyuAVdop9JvcyjtjekN/
SEvionFjYkPL4+Kp7yIaXMGUJP7S8wQgjQFFvYEUxcSpHRfMGR1EXAuGAjtAF+AuNkSOke/kCOva
u84R2Pu6+1mqpqTmG2AzkeUWD5pB9JmBtojK9dOEYdbi+/lY6VN6X1bzV8adXpWdU4el2bvMj8e9
v9tDjjH/IfMKgpMF2PyGs0nMbhnnALDQq4npOvOyXIrxmOaofvGPybDLFMa16yjHOmPwDq4fTNtE
pMBydBve5ryOd9PRr2pqgXQ373SUSsfFBfKBsX/vORMSk/UqHXKButIMwpUriUnY2cvSrJdT6j2e
Q1KcJRiJyfljsgWwTjI39rRP9uJht4pNqaRORcoqfDN8n5WKqu4q05HqeUyW1YALhgLIZB/4ArIT
1vnJq4lhdkgOgyhjlqAZqbraLBH3isXa/ssYpGNuzBmw+WUZ9sw4ksKU5dawKMdQXdefhrsS6BkP
NtUjrFmKEuMp/Fz7G7KGUzlHR7FYmD3Eii2LhCXZhp73NjwYYR5j1JCyBMStddDvyyhMoH8OhPPB
VuEmYpRJxeVZ+A5Bswl0cJRFdH7bJRseJxFA+xS+6ZGGLErfenwDYgUFxmXftnPdJCWTKuhEfN4l
cXmDkYsVsCAsPqjl+kQq6ROME7DGrVJEsbhFkMLhWyeASMznx1L8aQQCq1z+BodPmLompnk+M/Mv
X0k8B5DhU8080RANmsKmqn/XCBhY7l01SqZVnAfig+nK9phjDloW4Ojc/b57aRfwA/Cfbd4uIih4
29LxRhI02oB8HsSzPX1kGht9yADGNfGx3jbSr9L+MymX40g3sLZ1zDxyHXa2p1V6E33nso+ybb1M
SCVGAP2fLr33QukieLkEUuJj2kfwi671mlprapyM+K6bMRLLknb7KMFTr1n32GLhExCB0e9YOPys
K1b2Zmw72S514+br2oLqUrU0u4OYbDPIjKR0xsFOSgvLGwjqgPmvamLFaKIJthtF6RBk1Xyu5zLx
FfmyShVDe/Vw0RNyivjXoWV5H4jpZ4r64ONFBMsZLzVGsuEvHBEt2BXR/egxy+L64WtGMSkelLsB
EWxit9+GrQCp8AINESLC6tk9GSRzTqE306SKCX0rWJZL9GARBSDeZZxorzf5Me93HypO+fB3pIdk
fdQgpUTe6eIsaIZwdJuPaInYEti4W0+u/0ZGw5rlJdvxkCcssxf1fM5SQ+RPUh0IwUJrdCujS3Vr
fgZGcZT8CXB3oEQJtJhJ5JjZEJeNgWfgU6LIMH5eez4USICjtsrovPYOoUTPYnbDhUhDg/cK1Xi1
jFBK5o8DMg397Zmdi01zWyVbjsR7IS41ZhKS4lvLLcQZ0Nwfb2EKcIOEiPb9X/eaT3Ymy81uM0UD
vj8arOyugEotePz8S5ca+VOMCSyCr01xxQa4zUhx/niRmb96rwBEZB2wkGAmbmx+dSqVbm0nz2wH
+oiucHex1dFLry6WbecFuFHf2b4jWUWaKYlLzAtLOMUSGuhBtgl1VCxCNAIF3ghRVrXUVfa+F8X0
AXZqC8e86Kx0BSupRn4ifb9+SgTgQLcn/v78ubG4xZlVzXR7QdfgFWLuL9qNPG3rHrNPGbaUxVFs
sQJ6FkIsN7VJ1SBt2Enk/635MT63GexerlCCxzSeP5plK3nir60wd2Z3m3ELhSmq1OP40LpDjdY3
Cq+Q+Y4X3ACQpBlicflDfXcUtQ5PYL3n4cFanQWiqEecX6oyymfYOmb1FKRaYLlbSqhAePIwbk45
1gA0BGaBDIgheSKu5tsvyIQBv1im2M5VEd42ND2J4wMVaNYkIz0ueWJTWd9Z1UDOSAd+LxJcx1Al
bxi856w0N8j8qVWS39wl5T+RUvQefXv9aEgwWeZVgWP/Cg7JjltLM2sRnH8pIOwYtgt+7MaEdy6Q
td+QPsL2106QsUuSZM504RsWJc1Agc+1x5WbBv2xfZrgKVCTFR3DHeuClwcNSXuruBD8jh0LEstM
lT6K3TXLtcyVX52XHs9wfJtUliMZ89T13UBglEwRU5aLm/VdkmSSQhclxdouDtJSgZ9DGKpPZnfZ
cqb3TGADNlBtSSItxPsP6UsYdSwVhUt1+DXMf39miCzZAMRF9yZKLbGFqoYfMvpVpD9eMQcjwH/f
WkVCJO6vBkevvfv1N7F83DFRzYGD+5IEzHahfDWagSegjFxhwKJzVis634xjBQwN01FnS+yOzBud
M0B9H6EmvkdAlG3z6egbSIUlllcsSCcdiBx+WEV5Vl0pPJ45ILeilQGB8p1jTPtKR7AOrCSwAEP2
I3Ip1M2ZsbkW2AM1rmYDjkNFHLt55hkU1+dPPG8CWe2y/QHkdWqbiEl4mjfn7CWVTFTnxQIAnEkM
oi0EbgccJipLU1y9zmIS73RN+A8THjKnwvzF7/qYn9ZeBkWdryMHHIhG8FxovoSAkiVFZQp9mS6q
oW7Gveuodx+fbe/MREszUnJY8kag6IHFvAWfZDj6h3BozbSw+1obR3FY3+ZtlsjfjBOTWjkBvjIL
2dCiPBZp1MwzULvlp+eJerAt1uPhWb0C3TwHtLrbVceoGwj6W5MDXDALnmmR3uHcAqsR2gD2j9Xq
S0VOzx1sNWSmm/TvjmZXoNGBLoABdaqUPfpFkkO9e4CfWKedCEZdgQSD1/7DZP1Az0a2zkTK8Ozr
eI5MM7CoFX1K26JLdP2hWoYYPBL9oT+z3iC8D1gj/o4xkUcVXJs8ZdP7f8pTN+Yx6TOP+/leeyFB
OlUn2yLmTLHJilO/GNphhAm1Y0/1uSgPRPZzJdteCsa4WZcLSgH9Whc67WG9JRZ3yw2oi8JOoO0J
PKBVCGBqc1EnwVd7brLCtyoaUnOriy6u995Wqm1Ysyx8Js+vU8C8AylG9GZsCtqwVJTJHJc23Uxy
l8No2FN9Zbz+JNd1okp5Ws9u31XJpxWXQrdl5zJZNiUOl9vhycjbTz0ykGu38w2ngZrG9rxHcprZ
HLur5YehuYxgUrDtmutNF3UY+gHq6lOuzKnZ9pdsDmTtsMC50KBUw+qFwR+L+I77+s934DkHHHfZ
6r7lDz9ejuQTaHnUKltUC8CkHuyavJPS5k7VCgvaN7mJ3LRlPbsujednkZs8uqczjRTSk46hSXkI
M2vUc2e5n1yU+HHwekFH9ukjH5PLtm16CM8hNwcRVmFkD8cvNAILfvPtFR2/z0G9WhkXtiIN2BKS
J4RkYCI0JQtEVxLumvKTWXkiSdOpMVDUvQG/RqOEJVsivP595gmJGUdRFJR7YFpsqhnbNhQkl+xm
7Wctw5Uo85CnRFAMi0F+xnhpwoC+izCB6qCDaNJVDaS0aLDdbenY6DJ+qfDZvLrcrhSBQ5uaXB53
JSxQpFsQxJ5tWmLu6iUWXymFMh9UIpMZBpf01abtuRC4AtDfGWxWysnvYib9M9pPn0ZjeCTTrLXZ
MojscoRsfRDxHp2Ogt+PaceVno83KRHCggtxEkJIu50VP3grvRCbYJITJXDrnth5nTYEP6K98tqj
OcbNu66mVQkLhW/J6/V7Wrqv6Jotk8DrE352BhWjOKrYKkaMIoJ9xHyQnou3UcLcj2cLvUpfynUb
selPChJO5tMhAqxFpDelfjr8xKgXP1cFUDfnfCxsgBZerwzldhNPYe+UdFEfi8NE1qn/+mLaVJpu
xVHBG2x/ox+gHvWkq/sEni4EPp+XcJD4Bnw2Ov8js+PhebbemzcEFwhwKlmrjo+A3uFGYObOWWrJ
B1A4goQyFL1OkoCl4pq9J20QaKOWxkMw5sAb2iKHN/2nFrEDtTMsAnm0nj7tzal4VJ6S+GyOi6+S
V5ufvQmLoFd50gKMylGIrcrTlPsHlzksrPWhk+Z1xE38rjbqB0oSG+91Qh78Hcl1UZ6HRNAoycpF
NdrU2Hx1Ps5x9MqIgddtGZwMyMNnqNGVFR157oZMW3i3TvQn7oJkBiTEvo5FOJthoZWipVOg8bZ7
to3f5zOALIFMPDsQBXlKFkdSbUmYfWbPXPaBZTLrjzE2KiIW1zHRq7XZfsuktsIhYzSfQl9nFgT3
2xtKS0htZJz+08XbHwyZ4AKJExc5o/1sZOkVte8VZSgi6NK/nmuW5BLyySzLQJEMLbXs5Uq4RDqp
XySBIdSZfsQbuo/ex9/2uqzP4HoIXqH9ZDszVBwHu5pvlYm6SRflPB8g6XKtHcjAJ0ENK8Jihkm+
+eUYQakHhzd1+xCDNmGszOgcA57aAsn0gvckmYH9CLBFVKOV9ONbWvGUOjXhzF6AyzGAvjiZu/ty
7vLvVuECG1PgBiKy2vQ4V0nE1EVwPSRC0XK54/cgd8GPHeRYQJJKAW/KshIil/3Up4pN6F7F8Yxh
rA/fYbIW/wKmqpJeLcZOon6U56q7TbXA0WS6b0oAX7DWzQ8EfNfFN0/50Kz9Ui+0EMuSsytKcH/Q
jw+F9ChrOGSq8ps74vE5f29NoQrCyKaTrP5ZUrvXeWc2TU36gyC/wDH21vCezVNQn5xWSi6xmUWD
s8LzjcYqpwO76oXhH+33XQ5C9M7HOIl/haFvtduWR1Ki+5Usj7448FI0Cm9cC78zjnWTTMtkaJHb
oI5QjrqOr/VYQtc28Vfx7RvlBucOXc5orEhbM84pTEQviF2kHqa0acfpJ9TSZeODJvJXb2Mt/sM5
d1M3S2/xRZk6y35y7el9wAWD+qqmcpZBN6Y3oba8ZQU4TQ/hNsb4iXUsX2WShe9WdAuXdwaXkXjA
Ow4dDjf8lNpE90nmbmiZScqdBIGpUxIUfu7B2umVhXaJDQyyaKX2cx/tN9wQsj4fTKkrMon3QYzL
wRKrGD+QhKzk2X9c/bLZIF8MeIktKiOOA5bjZTJ51DEXTxI8aqZXyVRcRFY7UPteyRFhfTU8Lw25
SVTP3dPZDDtMpD603DZIUYr6aC4srpB+9WQg343o1FiKvThZZOkGoMypwoc7j98r92sroBAP6d4z
tDhCWHZIhWTJW99l/C2C9DIVaHaN1tRFX8i8O6DNEr6ljkD7CzUyyXKv8TtXxKzec4zMDMJpVveY
21rNK4S4e49pkr89GwOJkBsfEIBjTlHQegxTjjq1DhyHZX9oxjsBM1L3IjEURUfyOV17uL1ZLOHT
/JA4AlG/Q7+4+/S2e/QPlYix152avPcdb4bKqe/O6gY0cSnOQ6cCtS/iNkrJG2HHVYNy4CsbgQws
IfgpfMDCrHY+Oz+YuFmYQP0ddE7cpagvVvF7MLApPqMGhlemXGsY9CdMuYpuW9yCKvdWyE0gke/H
Ys+/dk32igXfJE7w9YNQsq/jlzgsdjK+dV4d7j8HgADkl+HpIzCyD0rOkZ6N49KmoPv66VXAQWjp
LZcF/a3NfmMFML5OzoiTvgG1u2apO06YvpGpGg6/JqAVsuKgZBzUf0jvUwCflgFbi/ieNKqcM1DX
+KY1T4egRBR3UJvBprx+Y791DzdUpO6+9vRF4BoFzgf+1/MTqYmt6/i80jEPccYW0hXyn7LADrSm
Na5ZS3CYHfEBKYEpFr9eWJE2CuW5UaJaMlU+gdpEsltNgOC2m3i6GK3z8RAMoIsX5FbUy2UZ4h0+
TUYZ3viKhPWMb7yoxJV41a50eQCqhKEGp6hGMfjH20YrPz/dJb+BuoGivLD6V8YRUqpc8gtLZfBk
bAu783VK19MByvuzrBDkVVT/cldLd6lYl7Su76O7wyB/s+WsMeCZA5cLSKQkN0CP7FqCUBsloTAY
YnshE+M+pCSZAF4yZ+Tte9IRnoBcHBjlT8CSgWj1uGDCcR7GPAQpstLNvOW2mV8dDZIPU//QhZa4
og2AO3vhzxdhLp3cBoaz3OV69aGzbHynk6VaiCGx5hadlMiV5meLrE4/yNzMcSPaJ167zhIvJIP2
cUl4e7Tf8XwjrEa0e2ds0Guc0ZiuXwRtI4+6Vt52NRlpVUIHdTotDRvPZWTU6fRNcKnWy/6scMv3
AUM+QjsSTz9qPK4h2d0WetOcY2soVC15YvnFb16G6fW1IJ1pNvo9MoqvPJS9cv6w8zqoLTO5S8mb
2FOB0xb20ChBorWVxx9Ke9QLSB6CbgnL5QEmTLIyb/BA7gNCK1drVnpXFkWToEQOBBbamubnkFiv
JEFXzY7bYBCBTjpLvbKuECsHb2YTMSCSOqP66nlcYG9pgskyVTHMDlO964v2OKIwRAkOvJd7Pu3C
4Y766YHDjNK9YeU8ETxRsadOnA2Z64CFSHbU/IzijNl4iRGwnqJzjCn51dtnjOR6k2gxtxAO1feM
C5lYFFm6zqB6ugY71xC/zPUaRZwavdz69sU/SMhSrk4+nLKbinrBqm6vwyebGPrIp0IHvTU7X/ZH
bmFGKBKwNsfvixrEqPrV/mqh5DTj6L8sVns9uO7sm+FjfseV6boUD6AMDwsa0itnEghhZh6naDfG
c/W3rQET0Zr66OE3HVLU+cFvDzqhnyiMhWMjvyJD0CxauxisOmwrc3gSQFh3HDPRRl2CaOKQq9VG
7VyBlnBfUl1vfQ3RVGj7eBCmoxI/pwjFS73Bzdds+R576HaafgTzYJ58guIoqB87GYbt0Tf3isJF
lEXWlE7CQKeDKXPZOvAQ1JDVBjy0dl27/GpTCsrBz9T40zfrU4MIzqzeoYtEPKYZUPePoUQkrlG9
ZWS7oNz5oOCZ8CVtDDuinDDTZ4726ysp8Zzm9DzCaH/8aMaASml/HS6St91V1QiIxL1Ri2P+v3A7
D1It3tLfaGenz1Oc75c3YYwY6LkywtqpgCULeD/OQ6QQQTMewYWu6qZrwn0niLZbGgCi5UICTZZ9
3NzMIXIrpntYTttYPXH7eEzZcmIFcoQN/gH3n8hIc7mkZ3sXjpgHsnKc/JZE/pGcNCB4QDyq09UU
aDna2k8qN4/3Jq5EatTXMjnTeAJCod2AR+/v0L5Htl4Qj3mgoegp+dvjA67DLIl2trV3fnSEQwMx
afwZXSSzziDEbeOztN7WZOFZ+s3UhHpSLdKfOXmwiu1H+E7rtCduo/onr7YVJAg5JZVLYRz1tDAv
Chr15VDflUedKvx1fwLS11A/GaFxY51g/r+NHm0/IVaJ3H1tE8XKrp/J0Xypd9CRZN66vanerwr6
1YWCO/kEC5LLzAMQPf5DRikiUPWPa1/fksAGVdBWJx9TbY9By61bLhIOzAyAlErRVnzGgDbnE0QK
QA7/sslOhsL7/SipnBvHVkxu/FITX4E64LZW4pq2i/uW4Ih9QX6S9VgmOIYe2yPbnTZ0+k9DQCng
E2JYANqVMNDZ78FhVtvsdBf8KW9LEd+JrmlgBjB8NLI4zf2YUWAKPsSJJjZVpGKx1Cf01fdIvOx0
3D5G/mIZAUOE4hSQD41Y/HbQxyfw/gTxhkN4u06lHWrb+T8fSZ7Q5fxMEGEJHxgh9jE/k6MWxkOJ
3GVn2wTFk8PCX9fWUQnBkNaqt2LZ7UQ+V1FYc01sDCNufQng5uNFmVVZL1XI9UqHiKwSPMyUu1Zf
qb4uECQUPubJq+ZCYhvWIU81NyVMJvORYhzH088K8ktyv2z2xjugHGm+mCgmfrWcAvxsk91HZRmA
t3sPn3MQ0x38LJA3CD1fB5XuqlFjAZFrdz+JwBpEiz+aSxSf3VWBoogViqqHYZwA19vkQkTlatNR
J/FwzerNjv8wPSM4WkwT/FpgrpiqosVkattaRbZHUOdYWMFqOP4RPeqNH0NoYact57A2MK1eM7kH
DPrnyfFOUS7BF9ioqjqQ8rXUMf6MXG0upHxdH96SlddlN3QPnWwGiPzKaNQshAnix+dkPQ5TS+yp
hNauydBnCA5wgYaBVA4Mqluk343/mmAAHyx3tyjMkm51t4YTruY+QgK54O/RAOHgm33CeZGYsR66
xDJ/+ac69jJVS34kVXf5PF+ub86W3rv8zNqxfV19veB+5F8AP67NZlkU4if/lJkqLyt1+aAkbBuT
ZUgbYlS3GdGFqnNtBwsQl7Ec5gydkZVdb9GEvQUpAncc9hD3pWZcy1DcyujwlKZAKvVBRWME0r9K
/5nGOGtKMkmwbNvR2/Oi+8x5t2+L/SVNXk5czHigOnxOYrMJ5umFyVtP7KZaKeW8GfnKmcBKhSr1
ombjhyB1ndCFKIzqGU4nfhiMG8TZSXWA7iSTDpojJWPfGQ+HqmeqSc5cieIGqRCtPrFlrqpJJPlq
0IPOIrpwq/UEYWerM7qw9JcU459FbM8Es78hW2rGu2AJG1WQPA+gIkWvUX/rh9UoiURGgxdWFnCV
BZKtKiy2fsKtZM/hi9KBRbp0vVwzf/XN4X0cz0uz0eWJMUxSPODoISM4NEHIpTuYPba53w1GCxvn
uHMmVEHL9kBuOnHkQ+07sQ1iJ0UWwmjpSK1tTKNlgWqNoZVt8+MUARgdoQxEZZK1HW98G1qe/yTo
/KJK4eJ18Rd+jOv6xuK/S+ytpoTu2dngWo76m78eaqR6FSiqCISJHsSDk9XxOHHvBv74uQdWaHDk
TDSh07TRcd0zgiE3UOyWaXdUAUvZrjAm9NJLJ75pGRE6Rcm61ziTOYHaa5o/OhObR41pXfWbgOXy
cp4vBFbhhPhPj/V2Kwb+4S8Nam/r9D9nUn2kVD/Bz5rz62vqbppC2F/MHRbiAAE5foS8rh+D1bMT
8aHyXo9OOPbqcZ7cI1G4988bNAHnF+DawBVPoc6pTtV5bhje6sqgh5zr777YfWHBv4J6t+UR9dmE
Z9Q1nG8yrpo2WI/qjMEEzBa09nHPnK97EWkOu9ztJgoMZrAMI7bun/TtMkW6TZcLbzNP85ZvuTEz
2b2gwxj4sL+d0UJAqUsM0SdUSZL4xFfSckllmg8MgZ5njb3p0BYqkqSiNVGuJOYv0PJ+6RyXCiJS
3MRQVfyEo9CphEC57lS26cjYDDdBWyS9JXR4jeMEW9nU4W6cgQs4cvZKaBFUeyrNc+U2Dv6KNY/A
FhFbS9QCXGO4zovzpQgVVt3+vYsizoEeZtNK1Tuk05UXirEoHp7z1H/SijjHPwR1tEn9MYPwwf1R
5SfRFtvCd4GZVrf8va+Jh12J5D6iVZvr2KpNynQ2AMYSeNVH1mSP2del93yT5gFhMQOokANN1rsw
I3kECj3XeKbs8ko7dMS3aKF2n4eCwen8rD2hlrO0pKhBsi/JIOYpmBzFimHhux6/ryffR+9sN+9N
aSJqmrG6eDRk/O9evE9hgXSQJrA3Hisqy5Fiawpth08mjCVBfPUHD+PAHrZW0iRELoSt06Zb/wRG
QWIKLIEaIEFp8xlM3a4SdSwJ0GSAGFJLLyqmaPUD9GfgtMUUe5FHMVW+ddZcj6FxLvHzqxgNxxhz
ApB3i23uy2NzGjVixMvPwGWg8c1v1tH9j/HQUqX8G5+GIbwDRA9NjuTHCh3hbhUaZs+ovpq8YpDW
3lvT97sNrSiPOuWgYOTKMIHTG7VEWmQrwd5aGaONyXvBI6SdBcMmNJZ59mIxbmxl7RlbcoV/EoYi
GbeTvrWUGGuRUB2tzbEtoTwBwuUIizPzunMZFGMGIFTTJt1aBHhP7ItYiP/xHuNp6vOowBTyxPXW
+nc1UQr1B3T/CBB33bswpiEvBrgbN8RLpcCNz2H75Ypk0U30jC647KhL8sWuY8V3aFg2jbFsGko0
stx/TUFVrbdqr3gaseO+aVhB83nKcMPCiRTsqbrjjnawTWjVaqD0MyBaIQzSfv9fEhzDJ6EFhfME
6cEXnOJkJLbjGNBvwVxGPktTnCKh9YksxB2VhYwwclltwXPz0j+p8mdyIhJMKAugMrpTSX+/9+32
FA0tmWasx9PTrQuFNuW2viOT05n9MJLeWU9ILhJhNwQkm8M1IlgcKEwhEOwFp8MonbqhlW3H+H6o
iEKe3bdLbMMRWQWBz4gXQmkSpqheB8jWpGRl/Hcmm/PscNqmxzh3B2b9XQTlUuFS+AMILezJL8yv
2Q7jIEIQGkrSZzhYJ9u6CvD29LfzILy1qw1JJIFDdtQdxgvi5hRb9Ip5tn2zfmuzH9l689Ouo3h+
JgjQNjhwXuswIW0kr8rNs8mZBPvTVUXQaFMltBMHvPi2HO1qG3NRjZufAIpCOyJRGuyorQ3ydkIG
wPhjeR3QsX9XRnfKndUQH9jlpFKEYQG9lTx5iYUU/qHiAqSGm4tkYeqfrUbTte61TQ0CwTkk7O8o
hBhOr0SnOolyruwaxIjFqY17jQFS4W2CDa2xYXEEavYhfsI6qzpUEE+go0soJ8QgQltQkySmtVVe
XYsqlN5pcoktF6pTz3W+hEXYnUO7v0ZuWZGNcofc39QPWQf6KrNpMZUh8n2INSMbVu5CFhYxcp18
NOLyAjPsCsRx4xEOZ/pcmzCprI8LmzurlRC+DEbCnjmGaFqZ62r3J5JXGuyfQ8xsit2vz9FrRq7G
PFJHWHDr2Ty/Y9RK5lKhK+AXeSH12CAJpcj0Vp7vYstReG3XVwNhUP7TTFX/OUXDCvv4ML1Hp9SI
mcyYH8WqCpZErkOnN+Cn6j75Wt28nFgdzHW6o5mxSKbOond8jZPiaEbM3eydBbISY3D09xpBSoSf
bFDuZsZihqcDD+VvpAVTA+kyh1P6MrGU2Qiykw1oaMkaK0WGaBxL8RVhTTWUnJh20M9dx3NfStYz
vWuifVTKjdeE8Uvoqk1nVRR8zBL0ZxJbYsCprjsFU+FYF76DvPoWi/zSVfv5LzOc+zZsgBloEYrX
oX2nHwcLBYqu2XZWzuGXp8vPufLcNYc3i/hbqtbu4sNuUtV7jCzq3tzAknMgnnOlGuzyfXMjysQ4
T37wSVDJASpgw7oSilKFAj09N0Mx4Dkdm0MOcs9IMpv2m1wywGws7N7nt1ihYh2bK7fuKMq86YRF
ptyBlYblA9lMo0kz0vY7mT06TSED18IQXCxpLseD85gHZCikpuLx7NVU9678mBPDBhZSX4+jMnAn
6ei5kPKkK+WTIUbxvnAqlXFp7/gXsHkHrXUAERtziGYnMPk8nrU393Gn9cPsLbvdS/1afJeE9Sv4
3TCB9LK68Nh/h6gvUQR4lY1gVRGg8sbUtC2/heylhRbJnSaMIuLpvfvzEmp6J+pf8dApbOtb6q1j
AjoaKUWOvub5810LK+KbL+CwRUAejw9wcs7o4E+c8d/sxmA1CDd+yodJ/AgpBbXID9W9+Neh5C75
Ar7nIY7GQz6m+sYhEIpM3CAV3v42zgvn1Us5HM+/mXFqz8az9NAgcgMQJ+9Q3V7rs+QeJ7nhD4HO
VcSTo5hMk6JvOwy6iN3iAK87IRUyA1HfipA/37IWOg7utaXtCXlbdEqgp0azriLafQnLv/QJQQoo
dwxRR0tCMn4IHdQMJMNhcfLutb6LjVzDRj/Syut1gNMrtLnbIBaHifDhSMnJ8pPLIP1T2DWTtDbZ
gWryEvRrIDaBcMk67zG3MrBcIDrZzmpikZqSo6G+3T43g57Y1TK4OVwewDS4SIjMyxBwUGXK/ydA
MWxdEyE4MNHRcbymIUz5IRWrfBoNLy8xI40T9UbqwwmXBsBSmKYOovrapNkgMzHa5HVi8JxytgV9
gfXt2ATPu/GnsyvhjaQ8orwyw4xdmUKKAbSTUIAsMAik7cNmx5I7c2yVGguzHcadlnkAJqaGja/v
4KN1YOj8qRrVdd3uWFEqp4K02E66Z4/d6QNo6iv0lCfWiiOJXdRWUQyAGUeB16Z/jc5PvqI6vTAr
a+2BQwVi8FCe/+ns2glelfzryKrEZcK2jPhBP5FQtIvzO+ct0eqY1h2co5wFgBaI+XBRHyf6R0I3
tEvTPbVL47dBM7ykJ6X+CZBgbWY93ppTZItYaLZY+w9hte6bEgBChtsZ1aGg8fn4/GIvhrVBGCE7
b9wrkwcFD7i9fVq9mwNRZ845kFcEkfx8RHYtnt83d95phmlzPtgItKjvXVViuE8vzFwkBJ+cYHM+
88BUQ3RY9Sn+M10ZMWbnNFAl6Y4K/XG18rAjuIp7xAvp/aVkIpJEmrLf/6TYCkuFyXBF5JIGqWBg
GndgCEEs5q1SVTVLtMOysnk7QCBgtBRzou9afrgkjfsXplyMYDPoAvUiA8ewVII/YznVI/A6VRTl
p4YkNEFbrbH5f0h5G/8+EUZScQH+Norm4qZGjDJT53awnK6Sp5l+du9V+RQpCvxRImZMqYtTVDaU
lFZSft2M01hze3k8/Hw3qfgXqqmBSwAIz0Yi8HbfHnwRScxe0jVnjZiZuBDEXv22JSGP/kqTEYAo
iV6Wved/sepBI57qLZvP11O8cRxmOsNbCJrwcn/q0G9sGT15a8TDz9GiuiaRJHKRNH4p/HEXYaQB
kj38J5lACFdv683M6qQdaF5SrNlaOb/YdID4g2NC0Cn5TzV3HN7P+jhMOp2Ifi6vZdQvGiOQq3Fh
e6Lkz3Uvn3IqEB9sl5g3pgCu72+QnnPaZQdMLDlg7CLYwzyuri4EoViReopBUgLRXCEYAW7sB6qx
+jrMBjBKkG3LXvlcSNXWe7oaTeq/SupJuWq4w1FcbEA/FbVjFXubtHGDwCq4NQwcy5cPKipKwl4w
yPal5yFK6McYRJgJMUIJJVuGvMxqt5owRJIySk6Bnfs7BFK71Ah+rS/P/hBoehjIq4iF0r20pb8Z
MtTje4KN8iGcJGExh3JAeUUn6DFlGBoaWR7U70j8VRhwdtHAScc+yTRTSAUkUd+sr2kdhys6Y0kS
+GssZU4EhOED9swRBvUsS4y2VwVG0TdJmh3XEoj4l0bdZ+S53Ika13ETWvxD1TAkXOGXDr0wb4E5
kEmtqwCzb25t0RRyGb9rtRMvmSeG9kQ9GHwQhkgLOXXSBlPUL3wgRcTf4YMmj0GskmgmkfyfN6kE
fcXQDu69jqrDGkXAXHc6JWFJOt853+djQAXFZpdi7RRh3l0DezqmiwJIQmhUX0VrZf9A+/8dUkH/
lreRmQhRAnYpgmRppC93Bz00QBp+SplqC1nLMOC/4kSvAqm9C74LqkQiW6eImB/YqhWHyUy7El+j
f2n/9SBDyOLICleFKrN50QQyytRMg7mSLDCnad0zOvcSsZqcnvzWM2X3DhuFS06xG9djZIPI9747
5vnqbYYA26yrFRCFPLopbVYFYGfsToFTCzsU6CQwjeEuflPOfCNtV1LKPPKN57fNcok7bqGWfaei
quMX1wyV6BR2/PLELmc9qmTTHqbYQZVAsdfPOhpu5jDAbluhFaXCOASPgeR0CW6XL7u6gRZ4wPj6
qUQAIcmMGYu1udMwnmrv9a4cPRWvsUux5gWqPxgxtnjwfBrjZVqCdXZw07DNoTitUcDLjEG5i/Db
Dnt4ZUuH4keAAn5QYF6G8woQfb/jNR2MosZi3t+e8L6Nfpty+BJvTpVEhWq9vUqYh1Uq5VcRMDe3
PbTSrcGcKmZX+Mm43LlMYC4eJKuniB/A3E+22BjrKnhIfWhn9rGazLfYmJ4eWCRPKWc4pQgPkqvX
oCH52v/fdrqMTEW3fiXr0Ljt4L4yjDXGbcfoVaSz165GRrsgKndP8x49l/gpuAohce0MyoQuNLYD
OhzJ/GzUVQOQp3hfbXZTpZfgQPqulexw2pi8Agj9OdsEzLnq7sobGH38i6pf7oNcbQwRRQOAs++v
Zr/0sSdSuisYExe9QvGqOFLh3jqfQLIuAEnRI6E5klwv+NnhSow2hzktjxBcB51HdH+006mimeDy
kP43SEIVHi+u5Fu6bG4bIn2mhV1AfrtcqSetdJpqZFbif5MGuSJL8gEVdxbdigoJy6jTFIufCFMm
d0vfz17lERnS1CKWbEP8IkfPwnaoN+z3XhlsdmIBBapYnl6dSepGDooz5e2Lc+cOoFIuFSqG520o
8LTJN7OtdI2uCxGG00RYHcyaXBqu/lsxhPYnSoj2U1q//i6onFMXDehm8i08x93z1Vdce1ns8HXS
Qnt/qlQrT3sSGnSh4wnLLWSnt2h9gkzmDB1qNnLRLED0PhqNikwqeb2aMKMxYsgjTHEFRd6T7ODH
QYI+zI6l9qdON1za7iTw+n4WCAoUDHeiYzrn7lfbhFUi4f0g+jOosRdhQk8VcS3JzCrhs0+sfFqi
Ty26lArn42VW33lpMGrtLMBV262wAhwNklIgtDyyhuTd8bSd6QsVsIWsPaTgydOc2TyqMtIiYTGS
s5web7rWAbiGLT4verxn8nfRbKsvPAdB1ev2bogDyBH5zCjw73PSep9C0xfdUxvmB9AKERawxkUE
gh2VzEqFhgwa1UpfLL4J8Qbfqrx2SNJD1BXWd3JBJUi7xtHghB0tDEVqw2MXy+1kRdYCgsddoKK4
FMkn/DwrIMP/G6107S0rP3JY7SsMAsRN8LgGhgunz7GfyHGUlD77pPY8CSkGnGkhAZvPFGoMfqEc
kcd9/ZRKrp3yjQSVUIbp2IxNMA96vBuCIZKjqcg2xxNhhWbg+hoV8kgQY2eN0VLnI/kwvyPDSrGN
4Je5M5TvuYH1UGLuc8PP84ZrNQVg9+EdfEVoJH67U/5dw5El1um6VGqYPGTAwbFkI+oqCDD4Pko7
IieuKwAI7Dsc9OLN/+QWlyWmGA0z65SOFDDiFask2gjS+W2fywP2deC0Wz/q+q/lcDMLbP+hI0z7
pBwgLWr98AsxgqYgb4BVql1ARdbAMK3WD/M+rLdOMEVE/cagC4ug3GSzSM+tvUSKzE/V2RV2UvMC
Hh45uDvg/Hi5/Flw3kwJhtDf4sVNU2V6udMrcVdNCut9CSbrEOI6kyRASvJ6o9ytI7cwJyyEalR/
z4SWSFjS2XJOGts+DTDU2uU3JCDf8fhE5al3eTy5gmMRuOZCo4ePv8REnwtWo7ywU+JheSqlai+b
pdBF3PELLTkQ+Oa5+VDDJute+XMdsszVLRS85SHcxl5qsLqbvb4lt2zbHh+yqDSHCnPGC8rpWchW
EVPH/kPk0IPXRWzUcqpFyMsCpqtsI8PHmw5DNOG6jIfsxoNrA9esyYm7XzuBzd9muSls5VbedjOJ
dxVxmw8gLQXUHgZmVFiidyhIbe+8rqAbazuoflAWj7CFkLenLpako+zEtVrPcHy+hX9spsxpaYcS
/ct+L2xaOSpdOH/0ad6Emma01V9Y+yql8e6vz7s+6d4EQO5ax5XaQ9ppjZrglpLIAOLMtGVZWQBg
yOteM1ZCqq80QD/WvQ0KM3Ag4fqDYo5UWD+Jiih+ysLwpRpsvpVemIEuekFXc96HN3L6RJA7x2WL
V9h0KAiMM8cO1/dEe6HPT6sRox1vAOKdfQzt4nt8A3QvR+98HsyymJTXFmNCx2GfprlbhkerAXi+
pdNmzWLzr3Uetq5gkcEU3yqw7fs2wwQ7XAwXWhTycorZJHPjKsbKVsRgZf1pXtOIL0cKj9ZQWGHj
APtmncZx5gPb/AqVYLHr+RcFq4YrkClISrgW7yvOehsfOEMrIw/jaqdt6a/gq2MruZPoi6akgkmj
kt9CZEapdLTLUyt/VZBZwehfJMVHMytcnxqKifKMYT8sw7smzz6FR8RWKU4GglyvpYIezK44gDVz
413907cCmAdPXpMxnhA7NRvugmggba3CZaPSOtXjmT4dAc5OPbU9Elo0jexS2b/7nOoI3QjMh4WF
K3wC29KM3vxZ5r6GHBpl8jWHwSjuk359EuUda2ifBCD7PAbYg4r65FIaENkvTgIz1aVE48P7EYxl
/pwBJDjQP8GqE8RXy6ARyb5642Q273Cg2n/TqBEiZOqVIPpyxwsoymfu1YLTD3JWqJBNvaoJvM80
yYy5jumMnTdtZ0x8MUfE8+y1VTFkIlRbizGFTw2a2sRgotKLkA1pasdMTTlaY4Saq7ixUtSPZYk6
hf5eY4tClZQP5g13lHCZp9f/DLYgGEG8cnDpCB6k+Ll2hvqDMEE7+O1eknAGspIWzToW8fVbcPjv
5fa4QMzLNMVeaFx0jQnNr13p4BiH4WsZdh6IrW19lBEZDiCBZ+vAKS/f0V/TZWMMoGV2MfBjRUUf
xEMOu6e/bo4QwtaAIsov6t7avXUzRq8VbvO3sAwCw9gWPCaw78QH1FDaYZU0F+3s1XrN8Hj7W9Qi
K33MFTr46lnI/lxBKleLYJ7Z6O30r83U3QFiZ+RCfHK8XP3db04F3jGSwXy+LnwdL8/PJNs5hL3m
3/YAKatXPb51UhhG9iJbbSGbX+wE548lJUI8yBFNfYNbr/oCdD1KlJ7Yn0IVdn+GzIM31HK+5Yox
FohncxbvGTpcjhT8Dm7KRb+OuB+gjfySb/V5Zosqm8ytLKk+jR4mFEufEU4eJwPwuYp4Egs+9rNE
F5082zM6j1tFWt3wqwLrqYgecgS2TySh6pZ0PasSolZ8ncZMKa/RaD+zg1dQWvhaaKRx0NeLcJ51
AaTPqaNwGo3x0l3QiqYWs9fr4SO8+waY6FurEtzSTZ5NzHQzmQdsEgA8Pj4ikriewnC0NPvMAeXu
hyeSrGklITYMrRJRGT9aV48Ah3uRfWgE7oVU445RyF31MhThaN+Aud/a+SFgPEWmSpCyA8unU7KY
z/DCUVtsmaM0/g97NNNmrWxHjnC0l/nab1UFXC1B5m8WM//SozBK/94Yebc+LhZLRwFn+eM4bYhQ
qzZ5UffUcR/4WzJILbovXYJOlKYwxwmKKXDSOHvrWAQhY3M1/VWHn0Q5MyFykYvLDf3HLkMwr6Ij
3lAqjZg43Id/eqKxu08S1gFq5G+RDft3ffD3HR5AebNr05h4+n8IUg7jTpWYqJu94e1Opd/KaGZI
7LkmtyQp9PkknCUrgQMPhAs3++0Hh79qL+s4wes0WXccXFU3dvJ68eda2Fhgjiw2MbWdCG4q5mJB
LXvDKk3XHUU95Yu/m5tG9crTUqdIDvv4CGXDPmzsDmfbNKSrZyo+2BsXCve9kP8ieuvfuvmFRww7
H3pXu2+NK5QUh1437rTTq+XxtZba9x2Em3v1s3VvDYBVcSlLcve6C9Y5QuH84uJe35MWl4rZEivC
3+7yMuf4zHqx3/FftURmdXiUWF2TSw7sEFYnf6dqw3WYQWZ0eo5VkJ3fPidiL6aB6MF1+/r9MgcY
tS+JvBMmOW65afwC4Gy2JqvUF+RrdY8TDevluJpntd4mnBzOqjw4dFLYNnD9tEpeGpaImdtPyfSw
X/9KzCzj5Au674ME0Y0y8DjJoSJ5Wk7OQCy5Yr92BPPmRuMV4ujel2BTKX4I1Ibh3Y3f9QKUkAu1
3IEt2zgkze4/p15OdfDg/EqL3ZtLM3kA6pMv1w/Y1o+DumNzQcjvBTzmDUeS0KRsL4QxSimbknCp
2PXGGXx4YTIp4VeWkgbV9kjsHNGUTMhrsQNMpvykI334KUpR6zvKlklby3sWXsWDrpSIUnU3st3J
SqTDGVSP3OpELmJWT3+nFeuswmiPZIdrYx2Gvy73pQeKO10LDlN3cBia4zbDO3mUV7uqVTH1IK8L
sOdvrr3bo8GcX6UMOK0haHprwB0EiMdNzmc/hs20DRu1OaIwsW77/NLbdKgU/rIKuFdDuU5Nkd+s
QP20YhXeNdD0HggaHjj2T2A0WcMISFbbFMNQKB7IPkF+D+iKFm/mxTuktiVtvB9MKpIiGCUFubqK
YKIc0FwKKHL1yBLyR1S5oUREPloyuFYhb7q6L6qgccmTL2AWGvM1Jk9g7+cudlcGNxpaTB3GMrpL
0rSJv0CV3RolGudjrjU0obE9z8Ajr/lDr0iet7f7h/xl1VL8N/axQkciJ4w3oCJxoFZAlzfsJ14w
FdFlDqURkIkbwZPtsJxmnZPbGLbldYZti15BJKO2aX0gIeplkb4m072pw0ZjQiBdq91WWdujKMEa
GR8PtrNLDXip2MSMgaHbhyDQOuAV2kP/Mp6EM3x1kspateVqsGRpTR29tU4OTl8UI5eLB1jMxQRY
X/aHiGr+hmnGZcXqtK6gNZsOgEndAJLyFaaAoLBX5jpV0A91E7we2S2LyTvT9DilZfa1ZQI+Jvxs
vhZa+OsltSnqFU4XYya4HMcw1tOVFPiB7NdhhG6g7wJmof22uAk03H6GQ7zNIZL5oBaTmDAncrIh
PrMTwiGyfVEESms/+qWLbyr0KvXPbY6BUU0yMk1flPDmRcdeeEaZskPMS9+7F4yVIeMpXZWlXsD3
rTLH3WQRbWCBCSwk3qiGrgyicbvlrex21lUOW4Kq7GOLTin/TYRjvIxWng8jTaJ5Tnfsa+k+bXP8
7WkkQd8g6d3gZzGfmlCQfgaMehkExE0fqHBkHw9hO5zg8dEi+h4YpcF+U4jxV2MQHX935ux20wKs
Ocmh5yEjRf0x1BTFRAqGkeA+MSNoqlIxnvBsPrtGcNsOuE+0B0Dhk13MtNOYzFEhHT2V7sDmJ+7f
ULbukJ3187R1rQPD6JB61sOthjWh13d2ijl4RnAgxsStOqoX5JC3o7KdAjH8EL+293c4VGljzI6F
ZeJopBvp3pxASYrPwDWEEvu0Nb8vrV5ODsd742sa6g3a9GFh3MLFerlMClVZfCU5Tz1bb3hjjaBI
dKOBzW2+kpbzKmwKOp5nJeNN/mnzVNSKMzCQPaiyaDvVh+aPLHqeqvMQ/kobjNu/2Tt5TYQPkhkF
ibOtxqymzhZ4z5hwrDvqbIKJVvhNs5u76kvd+OvVgl9nx/Iq1Y7o8AUmWwNLOHgQFR7sbQQQSAvQ
Br1oyw5CYUuUIWKccmWjG5bl0mibePPVFAkQfC3EbGt3gosXxABdnNs2heuwHwOhSzefrbsZZgUJ
K8aO2pXhlC6Q5o3hPFHpBMjK9Ez9w/+rt0/S39DZtpT5fMSLVRXneGVFThrpv7OeXZhZKFtr1+F+
UVFVepdBbLkme0YD78uxlDLtXqRO8RNhzRTnjpjV5Ogcrr6I8R0eWOGlUiXmjDvQU+RC0RbN2DpJ
mFXHY0IBdFegpyNb7FNGJR2gcM+lP5T2IB59t+N1sIDmh1q1hpdcHDY8PJ2J/oc8rCwShiusMqkB
ZkPu+uHTrhcp8Ixfk3PhfcGUYgt1ZzoqVAqJWBzq1a/qC/aoqziBLRgrB3/wBEB49+AGMbnz8qln
SQ4b4Yu+C/8BzOXj6WIY5VdPAplM+51XX5odGN3Vse5gQ2XlKw1yz4k7+lBdoXvJ0hdOnWa0SF3E
Lg9AqJ3tVtS/2+17hOFDTgPvWiqQPT45rbISSX13WdlixXo8NtNfOha2ix45+44ItzqfMi+Yi05O
4tcTCmOyhcKc5MBn+E97Ae3FGKVwwN2mNHBUPQSRPMTAUU1yxYKZno1lcRlt8lZuOnxYUqFtJb6g
VHNmQ74P88ye+K1WYyP217jPo3GLbTExBDbq9hpj0H7h1XA6oIP7CzALJoD+tmI2p4eNbCIa72/f
Mo6gIpD2J6/HDYWEy5Erippu5wvv9Xthw/9qx1/aUZYfwOe1lHR2XEGvPr08XV+7mU9U4DfT9BeK
mkOE2JvCFJmcJqA5JtBfHNZY3yATu2bc34rJajkG/DyG3k6qygC2Ol1NPVg5Yt1ouvWSP8UgLDto
QjHDM5ikLIJCzPUOcYXkEvxUwIeyAU1iIR++HD8kndKnTKTBF/0Cjqu0x5TJSvHgGY7jgWZ9LttH
YNNi1ZIQTawVOTCsngKrmJ3ZMcToYg8AqG/fYj0xUnzgfXQSroEGoisfhu78JWZW2qE/psjI7+wN
JmxAu5WY2UNRl7AGhc/lJX6NHAnt3Wcr8VQd3v42e+53gJLMdVJ+wKoejkPsxZXjgRH+Bf8SlP3c
yXB50DYTshqwHMMdIenpTSpIgQmSydNJ8IrlLPEGEND5/mWAC4d7OZs0zA3BVDAMY06vJhH8/ohi
A/Dfy1/HHIQGHwh+TmsF9ou5aCwfE3WzfScgXRNFxx44e6eOahuI9ZuQBCEQioafv16RjaHMr95W
W9OXdOvv8ZGKkwlYFohSboefiEynq1jJdluYUwEQoXuz17oqq4I8EbXD5LiXGPfHC4teAUglQsvs
m6gPKzHmo8fBBmHrIPa8/bzBE+d23dtncazGlcjc+avqRHe55NJop2X43xxTHvWd7cV+F4DtldXK
rIcbceAK68W4DN2SSQpVQ+GWYgOSut8IC8jpk2lb+kpGOcyL1QdNLPkYgy7dh2hzXHag9gWPGiLr
RYvoadCod4g6+abukF3R+57vBYS/mo8XHMf64ZbV3847Z2f3FP+L8NaQVAtns4AVQ0+YDS7Dd7Xm
lOgmL33paEohJ+ifRMEZN8oYkuLWJ85JbTtbpCt/MCXBhxlv8qVL2CyA1Y3ni1L+f5sqSaBE7iFr
xk9IM+KPEMMGk2zNngOmjqR5SvcgPltdI1cewVFatQf3PfWDroViz0cfg4XSGC1igRbcS9N6MkYX
RBTvJ7S6PDv+QaCsfG4FWhEg5jB5QDUFZQ2I1ItQzOw6+NQmY8ZvzyvBfvxrqeHFHALq4Eri9DDF
pu0etaCVW86fCH6tECbf0BCIH5Wy1a/ZROLWtZfm1A1NTVHm6kwiPt8Ynjrg7SjDLH3GCtq6tXgV
3NrbeYoj2svqnMKgI41+SUb2tTuhXm2pwpo1Jhrw0Gmin5OY3Qhd/jmt7d2pB7FkMUOOOwwQZFrj
1H/ZLU2VhDfleNDTYDayk4QwOq5O1kYRkp0/ej0mGTT34ZZYCHKzLoMx9zkueu+/G76NS2nkos4G
fuhn91zDuSfsr7+1mxkJqQtvFDUkIMYCHrQmewuZY22I0zXj079Ddw2bzrvTV/8cq32A4TVgM03S
TcvuS9LtfJQLMbom9UstX4xgiOYO8Wrrkcu9TnAxyQWnBCDgROnCOzlZeRGYImjFNX4rLhaJTQcR
zXXUKWGiJclPgMTWIc2iMkc/Gx0LSl7Y5nIdDBixUgzGKz0BFP639MFsEqD3ZJm0D7rkkn5J0zhk
KD8jaB7kRFMVnbN9xwGMLJ18tHHNBrKu0xUIYaEFdKsdOfA2clTNao0iZ26Y4n94ZZKJGKRKsoTy
kschrctmrvDjEZkYp7/No/IU7iUr8CGm3qBIZq7lqJP9t8atXEjkC3FoI+HH7fnXw+n3FBWMpp3F
uVb8E+vfVkWR+eia7O1IuNOgs/+OKdsy5J4VOmOIY0NtF6tYLmpO7HDe1nU2f1g9IQ/cLZE/Vp32
BC7huSd0xKlxui3c/6YL3ajlHx3GE4rLAnYFWwX/f3TUU6bwWpLxNx7N8JWiIDa7NTvsCE31WDnl
jI0AMtGjknEb1vV76IbdS2yvdglc8282DJY/jaCVvSuCp5vYe9LZIdmiqu+tjrJgPqZ0aWu+cboo
V42xbftC9cfqzJ7QqSbZIZZh1WXHUu6CA1bWI9op6g7QiHjc+cZmXHsf5y9vbnrfqDEEkp8plH4l
nECPsMndcIlqIP9Sr5b6dtTuyUm88BwEsRDYJ4DZH9hGiKaKNMORSx5KYSMr49AbTsF2Ikn4Df/N
bE5vlr37/LB3LlSjtHOVrdTqWUX/i1JF+9ivAwXc3OzjUroJszuwQFTqJuaaWIx4DkQa52OBu7ZL
dRv+nYU1U/o2SHRwpC46vVIAGDFKGPMytjS1XyOeS/zO9ZL7Uh/pnW55RYv7fxA3d+83lnucnxjz
IrWnU51ICbWQUywcQUygWA3xaN3+2fTRtzV/NQQ8DJWs3a0cTjr5jYPtMgubsul1+QbCR0EYVVJY
BfCGkPFuZaiqItSoQ6sbPTEpGPfCypYtVWtgAshPbi89eGylF0JHe7pwdBRqSqY4Bohmz/j2XoO+
GXunFFV4TwsaIHX5KEAOF/t2tqfVB9/zUJbzEJpxhXxODk6nk5JDoP2RnSzZ3WWgPvsy/nZ7Lv3X
C5gwPjsslXC0guxu/Ib5q/qvk3pWlEzifEEJcsDnGtEF2a3jIsw3DwXAcfWP45tWqP3AHxuv4fvi
WLfoQ/ctwB6lm8FIf5h16uv19isGa8hAMXxHVdSFQ3RIKMSU7kW5KCIx3z4bYO/6q+t0t32Cl2BG
XuA5R6qJQ/o4qUjjR0dd4DKzMTnFIniofs21XBLsXxBE+00rVcUW4d78Beb/JezvgEaVHHrm7De+
qXx9gqo6y22L/8EgLumscTPpkZKvmtAtFDmINdzOy0r2sTLK/m3nyaOVIaISOcnlbv1qc0R1B4SR
shQ5ENU2f8q1Yi/2TZvufiPGRZrHqVVmIKYpR8Vwww7EQQmlnH2TooPojckrGBxqadzpWf9ViNbR
leVHMAXu5vrG/l8sAB/rBKnF+o5wPNXUP7pA5xC7LWslHlATRCDCmQeNyCb/VozP5U7K83r8WGUo
EYir8MzAAs6WIgISaI15qgFsKWTAPx/qvKRZBNtkgTrw6Rf2RKJr2DRdJKizyL0NpZLba/MAI1lj
Z+GfoymBjixEx3QwEpwpI0NJR2xrgpD5SyowA3I95CDw/IqWRXgFopbxZvDhlm8BH4WEroeO1hvL
Pcf5ZRFW+WcZR0LdmfDw5JjFEPcuP//T5XF1gGj22PWUqgJrn53L8kHmTrQk34RQ25DZZC7bOQMU
2awCuWSH4qcobOtRDTEE/9Vx08CHUPnHwEdDa/jRVremIsTC6hXIUpcJfCqHfcUS0GlSFPi3ZipJ
8orw3ew/BCiCDguboNSWtlhrlllzK9QXfiQbpGuPvfxnVazzwp8lS2KpSEBaWbWBbeun0pxWM0L4
w0EpjGuU43YVY4PVEudein6BhTzIF5AiagijAtD3M3YKykYSvFzS6uVePvEkC2EsnIRYyaiD4JW2
Gts3JpPWjhSiq9R9bbLO/Oj4Ri5Ur42yeKq30N5WVVr1bujxBLaWyfeHLmH5E/4EOzLv09EkdP4T
IblJ1qtyGcIcJKeLnBdDiBsj8X6r8aZVr5Gd2aExYtzEsKCz06euxeWlY6G2hEDQq5s0ri/DLnYr
dFL72vUN0NSzP9rDJ8RJA25ZgUWnSgJqikqeFKc1egD6/kIYBKmIUSYzEk9K1fqn1BYcOXBYlsSC
3YDHy/i2vWiWSNSnb17F7sF/MnKPRKd3zegIWRDS6pQorDCJ8uzMfAR6tonUk8QTXFVR8+sLn+Wl
pi7Yk9RBvd8BflkFR8kvM5s8eNBL50sUOrshuroiDhkhwNsb6OxKL3bFRSa5ncy8KQOxnn0gcQze
hdgPnqnBf+2TUd7PkUSnLyD8Qh8/f7aUIOyj+8VzA+wtjLZ9vNVF2LcY8i9d3I7cT3X7/+4Fr1en
s/uLsMgljPAOR31HD0LU4LgxFiXN09O3hpYb7UlI7+2a5NzuQtK79Y0G2smh+wfJl77X+e1raQCt
CkMnB6ykXjVdM4ARiZk7+bmHYGE0wIjS/flIbvf+u9VQmRK+q2FJCTVxIajmeE1G8F0i9rcKnsFM
H/iNP55XlN7EMCiX0FhGCHDW21Ot7etXvXhwzveh19fOaXvG3fEpgIo6oWvizf78MDtT/8+LKOhq
AglKkMO/urOp8/j/GbjFEG9WxUzPX9iu58ktDFfJL8/c3+X/WcJ70O/R0F0J6ZJD83W8DtlZKVjm
YlNyRVU6yqkWQ7bCO9CWK/EvklKDTjPU0F0fRVHoN6GLsWnVtCb+FGEo8Oyj1GYigfpUkNJL6JT/
LuDBME4OuyacSnf0Fu4oNlqeIHe6WpoOIZH9kCVkKOpQ6DMJGPWKIm/iuJkamFJLxLHgWlTBooUV
tFH9mPsS6LQK4TpbM9zfQogw6UraTZ0hQFlvim91y9axRnJAmNa7l8vbqhaVpZsK2xvhMzG+Vy+P
De+8jBgGagtV4p4VNEke23ayG/T0rBYfGaUgr8V+PHQtp/Cled00Iy3Crah6O18RUlOS5snCmNV2
+xJ/BwROK643+8IN+L8w/Z+QP2ryLA3KEYVfhOazfdBRjlvZUzZUY1MCyq4fvSjmEXSPyY5bQzx0
I/RNoEqwr7dDj0m2AodppvBNEiGr8q5KTZrKhnUgoi8d1LKEni2lDDV6cw3oRLNVrNfZvAHQfyt9
UbdP0XrTnbWzmcdhnetAWUHkCzLmL2lB6zK55mPal5pRVRA4Z+6hKG9uaiNghd6eqYEl52Pye6tJ
GCJVJjkU4p+3DBvjgN71zNU7Jtn1rYG6aCkpYnCjwT/O5mDqxfYbxgLvDpz+d8u+Hqjky4lPGB8w
un9a4m+MfHxavQ/av8ZduhnDJNafixTu825jcDSbRdww/xHOulseI6xm6NzpeUN5fbq+jWjMDa2N
v2a6yZ5PzFikRHixXpx6foEPj3/Q7diggZIPNDfrS0cDGoq4Q3qcBdNu000+u+5wmsVPk+koIHqB
DaRu3WmdXc6FBE3XcVNumI/7cu2xUtSL7ZbpaksywzoI+MUdFmu3jKMzy7/W6HqV9tIocXHHQYGL
reb8DyR0vPEa1ZevpW+Ypzs2/g9Bcj69/uYjMcgef4tnEOypV2OdUNebmCd+f/3oJq1gnToGoXTx
EpgU15TH+OvM1LYh0keFsoZUHgoYTr48iVE23FYC8kZswiBUtagn9UOAWFssubgmnNsiZ8gTvemb
ayeos+xGmGTk9xuzqQFkDow6zSnT4xeRyFA2VerE0jNB3Oz62J7XlUs+BK07qH0TgPjiPtsWi8e8
v2YS08BD6YFX4VE7Zed36ay0Q1rkMILBlgYyhtfnnIFIHkx9ss9HWM7db24g4Hq89BSPFcYvqX16
HXGfcKztMhVAO8V8Kwiflu9ERE9gbcNNnEoQAtp6uxU6uIV0cQHle9vUHNcnVFRhnEEUWwPK1m8m
cbKeLGekG0XtvwFA3L+7tPbXXkUacW27gAkviWoJzQwvP5BmpHA1fjPoEJLX9pG0Mu1sHJol03MJ
4HRt1J7MiWBo2b6e03b48F2PcEZ7GzC+tcqhhUpCsU8BydhYLfQHi0MAofv4iUkQMxcWC/FsGxLj
bVdcK0ENN7NQU92xuWyNJBpTIt50yCr8FR5BT+E4Bcabm52vQILN5u57FnxljdI35QfsltI80A3T
wK7zzrGD/MLICmth9wYa2gxTYDn4SIXQsXiUgXdOWZwNE1O5W4nJHG0u56JXhSp4ZawSa0PpLKGM
gp4D6LfiYly7ZwgdgGX1cxyIxAUgZHkBf06VhcAl4OUb5Wnbz3vWDpjs6kQ3bA+rRLytXc86TYlB
+iCw9/5pvEi9MGMzrPmuGApNYzIOoratSIaYUvWP7Bb3eMyRQPqXz8GkxZLVYhXic6DSrUOCJTUj
94964ym/yBpoybAWS8XAw38PHMulZaxJXVGCXaKGBBB6QD1BC0I/gUib6jDi7gN2YAl+6zm3iByP
ueNNE1anAarOtKS2rE4O7QZZCmWwGGwP03F55/tc70GGZUEex9uQ6jA2q5VtKL2pdAZf6QB7VFsn
LugWYNN8COEb0gB2Oy8FakckZ4rHXJ2XbXbnQKgXOnr2id5U/ua+4G+e0nY3nEsoKiZVuStM032x
5EhHgM/RyxRoqq/DgkwtLVFOu4iK76wlN7IZcRxnHJuahOluqwAVVQxWEnL4TNp0AwDqlpm9alXD
ISvcyT4GxNLesDVz7izlCO9hCjtWR33b9ey9Hybsh09gL7HmadaQtRz7/9DglFkunYMY843Cf3ud
VaUD7GBmRV1iE4MPF4rLz3NS/bEWvjzGFsIBpF29ktuywfXUMe1TjiWkOXHZ5IFgwdBVWcE/LldM
poidpNf6aqz40IGSB6gDS2xF3KqUq4INJ7pz6X9PGpHAdNaj8+VhP+eRJa+umXqP1XuLYnScU8cd
Y8rZODJufOWPBj+PjOwNsWTxngcDxXZ5e/fVuSFwoRZrWqtafe3xOdj0iLn4JSGYBJ3DHlwLuyJx
WA59nnKGNPMuzbXgR1DH5t+hI2nr5oAx4h36ftOB7FNUgGgj1GhVctb3p5M7ezyiywJRP5xHvQjv
PLRF71dYEQa2ohjF31Ew2MFDW8A0IZwjE1Hxg9NUb3c4JnwVdDqqL1MwPhfU+YW7VxkILtxN4b6u
UdQXR4v1sRfLQVQE4hD7UIrrH4faK2siJkP0dG8+k+gCC9DWLMCE8k3hbcTxjutN11xv7XnYukIq
VqEQhF9qYzsrndVkLwfABOdq+t5rhY/pkRqjp18VMCbnMHMDnSVoGsY1RtG6IMZ6FMvvd4T4hF79
zD/rqivnQ6yP+vDJiusj7qtkaJ1++4rH6+fIZJXZrxSx54nGAmVIgdQMi9qSmxZQgv1fjwQFPkGP
xLJR9aB6yTBak50w5d0eL4zCHcUEkxATOc2a0iAZ9+ybNubQHs9NbsQDRsVwVo5sbfOuqCWKYCRR
SfJ/C3to6Kso6V16jNcFvO1VJaYNRMYzGqaz12834f5Qc/8did9ztT6o0VgDTktHy3wklHx1w8gc
uoq76YLwm56Ef09OZ32cUZX/O6BJ/mpAg5vS0XvQdj99hy6lJoWEsvZRsyghYzuRtMk5eCUVQajm
jUmwzTCHPcNR7kqmp7nxmbuXRdo6zeWc/1oga6D3OA73ATdWK75gKG8ZslcFSMrmyl4sqffq9cxC
NFFu56a+u369I6C/PYZlG6EeSpFqPu7GtzrmIXrHnwkZDSPRKfoAomXH7f0taM4zidddr96num6u
4U6jxmm4OdDlgAZV8xRx4eZVTVRNz8dklBoAR5F4yugMUaRjPu+W1V5XeysA15eocBXfcneKBqw+
klOIZjzJurceozClcrYiFWO919U975ZYT29nBf07odO8SJGQrq5CkvVolQgVbjxBcjl2uf7GDBVB
McSxyLKAQUWKIZIcKMluUSV50IEFUtC+BSANBhLct/rQX4yi5Y7l9ont3sLfgTZaSXu6HKkpHtHS
kt2wM5H377CS2GogfCTgnAsLrLTod9MQnzegcTKN9mugFEX1csEwd3rmYt5n4ao9IQ7z2ax/GBrS
jbGvS0naDo0Nqr986ek/aq7KYUERu/dGU+QQztm20jIREvRZFz5YZMlQ/XOXBUm66A0qh7ukCFUk
I/SlmW5jJe61GGZMHZ82bp2r31/mLOBm6pEG+8TtEMLJJJLxKHgou9TOj4lDRLew5ir0MlA9/pQx
+jWs/bQqS5VqcRl59AfBaMjD+fAWOgDEokT7VPZ0/gnOteWshdR1dJvUj3WPAWKe/NoB6ENlBnDK
GbwP6/XEmkJlyWsgM0JLsgQFfJhlugOmIE0vZTyHDrLYSpk5dnOoMHFaBEC6vSGRT+fIf0lSD/tu
vgKoxSFdWBPIYcaLCgYKMBLmjQLJzaDkRvTAucXs/JNfAEpKILGOolBhdAXRJvMHNA3Gmjv3SglC
6tmVDnIXzrmH4i4qVZwAV07CNJmEzp6oGNSy7yolROnUDtX/SsqXx4oz7JyeTGLzzquTlaZ9J65Y
szwj/5ZIrLkyVJ8bhVP+EOXPxLJ92sg+51jp6lYaZMMk/PN8BeXQwjF8+d9ylB9FU2/v5JXv5GAd
ulHUFKTOslcQLWd3hW+6PO76QMS6KGM+Md6lRvJOQ03DMxD1rcp5q4edGmtWAKqbSpCyCjv+KOKM
BdronZH0x+lRx8rfw430/e4oKIbTPtp6NYzQPY2mpJCoeVyEpPN2y890JTOF8jN5HNMFcKWPZX4H
vHJ2kojz+CuX6E17QThqJDAQzSxJ5raLib7/d9JjgbfKCvPkEnDoR9lWZy7QONbuiG6PEhC1cTfn
aKRwfHcg85xsgW3TKY2GLepesnXv5X11vGHCQy1Id/vc+i7XGC34pGbq8UL1D1NQIRMpVvqCCW8B
wb7sHAweU1E2BLh7pq4+BNx1qIIBFpcpn+niDb/yQpWych/hlsgDGNmiI5+/fHTRbtsjuzCdkZWd
yVdfa7b2d8MTH7jIVBovLM4SCWB2VUaqfLbIbYq0q5x1RpZKyJ/Y5j7+GAjGW32I/Swf3/hvAtlf
rCiAI8rYdq8ItgwZx5nTtbPvE93HBWBxSme3b2HLBde+g75Jz/vKahj9sQKJ82wsiTjMuLieA7Ao
WRQzWoHU4gAsZzjgIS/r0w8e01SW119E2zOOAH5xrF/Ldw0CGlkbUf1ATj9ECLe7QVAaTVYFaRfx
HsXlGa61r1w56Y94Vh9T8muEgeGg03ADcNpgihHKG0pxx/+PFZ69zSX+gVDlwVf2Gx83u+vpRbJW
CsNvxOKiD5NDvisMzpKnH/TCOnuaTYMtXCSshr4s+a+MPxNb/6MPGHb7w+foI5D4FeiSet99q9fK
L+P4Ux1J973DZEt1lwaMifNY/0yeCHWKaAgkyVeYazAHpZUvVynyr3lnXmVA2JIq/rN300fg4ARx
mMzeVYSbmTirqaFkuCXnX3DEcYn690rAOZiyj+3dZ4QlnHwqf4y6qh/w/6QbBkcXlFnt0Pvr6Cd7
Mp+g0tA8ueKDhtu1Bu/uWSS5PAey/Zg3UD88VLhrC/jSdcsNahDHBJBmY1oFGbkXwTqy7jinqzXr
+4QRivyWy0754VQ3CXvB5PD90fhqwnXjBW/D9lPyU2u1TjLZDrtN24/WeZPFWA9hEXYQzm7w1EDF
bLOclJsqmHkmOwHydlIWx2IRTPz/s6yfSI+gA68kMmTasWAOLOz01QKlFBJ+OPWxT4VHNyNtqUf0
K7QuMYBLLH25NlX3kmPjD9M+I+SFJ8rNV3gTBhjgOaNbiW+GC8mXsOxLEyikd64PtdaB1Llg4WGt
fXryjnLLZXtH+JZJr+G+NXXzv40LE6UQ/UE2iI7t/tTbVGx46Y10z1GewMPJDzeBj4hiDAkFOCg1
U9W5FnLXtUTlZTGxTTYAy+6i83O3k7Y0nK0wifTxuq8EAuSgPTTxXNRWilrw+X5BCc7Lj+iiTJrb
ifQNEyHvtz/BXkX3q+O7j/6klVfgOp7+kwygWRnkFBmYyulJIF+SfJUQWzpyPvmqfbgzviDTs2+q
KbNrx05jWayv5bzu//D89sdTQz9LlNoFQxuv+sGEK9aP+E+eTdl5hB+dmMSV0O3RGubkS1DgD7jJ
dyO+2mPg9SwnQ0/djFc57sUZ9n09FyFsO1RE/jUt+VlDhz87XaJYtxkRd8GukGWKuX/7mKKvlItS
tmO7g3Ph3U+xFs+B/AhXuZUHbwKyMXp07MByK1C6gzjEcdNKhOp+ExC6LYEm+q5F1iVdZPwX6JK+
Sg4M2Fsode4R0m5pvL4g5U8zjWvytihSDiW0TyBNNA9QFSnhLW8jQeLffJSMXicfxFWW17wF5zT6
spV+D9d/0ZloGbU6oSp97+y6Iocc6yEEHjsI6hC3WEApg15BQKqtoJNCZ85UtdLUachRgSICokup
jpf6GbX09Jxa149Iw2GPW0WJ+NDr3VJx5n5oVplDjLuJ4eXmggPg2n/P1PqagCwLDHM/QHmkwiAo
WjoEOXGwYHYNdh/nuhdCXu3O6cCBMV8xFdVtOgZOwVRZbTm8ummscjBBj3UMoG/Y0rkYWhMLEb92
LvpUt3jKd7wMeGEvZd2vtoowQCdeFHDK5Oq4l2z8GdW/YnvLsSA4/iR7hVk+Ssl6uCbMb3w1bRtk
pPosHq9wlFwDVgEg+xJnkxVr7DDL7E1b8ABY0+I4F6KmdEEgxjSBX1QHZSQPHbDbn045YGF9uVUR
oxyitmnqC8ZLTqZc14Vla7u+34V2w2lYufvIED75zO3WmPYAzEANNmzXjHoNPTsP76VeFREWuVut
KeOE9JCH/nAp2mMEEdTY6xT+a9DndlW4THtZh6Uka85DWfHtePcMuq8HOQwtIBYJJQ24ZIyYBVfP
1uLEXD7XIFXgVOiIZ/5g+tivBJfqWh5YRyQtAaXS8Qmh6D0MqmFG0sTA1Cjeqsj+pHCD+9sEbILu
5BV91wwwNzLoMpZ7G+Q1v4mHQE1wJOIwv7+kh39Fb6WevQH78jGr/YG/9YP+rG88MNFYCRdNleny
NPjEYJYOd9Imh3NtVqAGeM7DuTSzI7KR4/nuGYlcSs3STRc9W97v0lTfSJnTbo3joPX8K8oOonRq
Ya4YFNEiha7tuBhm/jxYPL5akNLyD0WfqZU5NOquE0XHBdE0afbSlPexNV8Om7BYwMa6RyQR2xWw
qBraZwRmvMYcOxW0JViJDPMztvZNqD4iSKjixhnHLavdz7xKSrrWLj85AhfYQxziY8rsy2NSerq1
ash2ni5p8vHfcxABiWw2u6uvMb89F0RJW1YhST+x8cq2/Scoe28k1Pn1XJoRi1ohKRds4Rw3VZAz
E5C71/7rHjgoM5ixZOxpYw9+oYDeuezJIHNU5yiIeCofaqiv5SkMkkYlAvItBZRv0uUoJ+Jk6COn
LA06VikCE1U+5dWsCIv1w5Qyh1FO1M4hSMC7yMqQVn3IkQfEkQduc/GYCeA7gsJV335dEqtFNxUw
j6cR9sObW0ovpkcSeOP7ohgdn8h36KYsQuPLDvVz92JdoUU52XNZ8TCozuAuG2ynyOP52ABIBc3p
iGNcvjLNhKXbot+ZfsTB3DlmJIKFb3SiPHJLm1tjI5mQPP/niPdv+jSZt+nyYxvGzNjmnECN/B4k
GcWFQNiPzkeSzc+nzWV8bzruM3DVOfcpcwfp/NfsfUzhoSANdLDVuo/ebz8rmaLb9KN3X82oc5Rm
zfZz7vsufFFnY+iLIpUFJJXsKCALEbCQbXDYC2IslPgxRX0qbmAf5jNMqNZyWI+g1pXTFsqGG4gC
rFIDGAwLcXCjdpykaPAwBfx2faK+XT6sOmGqTBKRt1i9Qky93jLD2HfLAOD4iXp36Yys6bdE/4Zb
nBhute3WtXM6yst13JVvJUTOmK3zyXRwoDRhgYybkpeoI+OUt3vzNzkj4pD3QsUFdZaSakH3bTYs
EDt9w1GQFodqkB8T8pk0+hpxu+S3QhroEETFsLcuwiRZtqdvWnG/PL1fuppgInJqLB+FvOUlSLa/
WH+HQ03y7Qb0aphB29YlcASSRD6estE/QiO8GE++ZGMSRdoShNDrivnIxf7xE2WLhhCadmi7o+CM
B5jpt04lPU0SubVcYU5nyLgoolgwjWMqUqIsz94DTBGoR/Ddxm2yn9nC+AEcKfLq0HuntrjJWn7C
L+SlHwjErCcdqqoXtvH5Y5THOcyejKIt6kpFfJNvF450jQXgpkBTILq30bN4oNXa7leMZO46B4yo
BGY7SpqMkEQLKZjQiBCYyP7fjqTT6MBk5MgTLXf5VST+PBzaLVR0H2PEIn+MpZNsTt5heojFLFbF
IOYrlI76IX7TzRe2OX6fyA94jBkHcChEYnYtrxhpCD4iq1vt3FpL+KUu1CL3Yn4JVslPHh7AMmGI
kMhN43k57y/L+MI1n6Jva/u0XzXKKWBr+YCCfYjSsKiHQhEbdH3uB5cIDF5D7SV6H0XHekCw0Nx0
aFbIiYT/CzQfOj/w8VZSCJDULPdNTOUSXfcQpVa52si3pukEHfFBg4E0fPrPTWqnmO3Ur2cY+wX9
Wh3O5hc/iSGdIA5tyxstIW0maTHhSJjKTD+83EWJcu2i5obBhaI0nxSp8/oFQ61xjQwaEWcjYjih
jHJTmzvGwHCmap29V2J1zbP+f4OCMBqD6CQp0kxtR7/wcLou9sZaQMfJYMb2vUaptshble5drF6B
yM60lzIBdfdnRUGDsJHVnCPUKLxMpuCcVeXSnKtytUlvAjmTq+KT6KQS2q5YKuJBFNTM/H5Vwe82
M8rhDX1adeZU+G6xKN8VDZIZKHA488x82pU7/HbRQdJe+gtfhrAa01F8IaeFfOeASRaw7UG/WVz6
SZLVdpDYg6/Jn2zdTy/tZn24CrF4Nj0ysep0fzLbfrk+V89SJ1a3OhrE8lGtW8CFy1aRwqepFole
8t6nvF/mwxN16/HG8iv12kLdNhGBJSmUns41o/hcvnXjG81LnMag1Hd40P1cjDPgVLKLVc4Oy/iA
+7VH1dz6IbdELErfInF7X5sy7qEpQicsnWJoYPqpL5R5yT5stAmqCHXFgQOVLdQXlLc1jcEayBwj
3MwYHgR6wl3hu065M5OXmSDYLNImwVLtl+1AkUgwsqcU8XkQhc0SK/cDdI/kSUBg27hUeLxk2XvJ
LI2w3tw4gfWtVR7HIgCVvEJf+jeTBfu18W84QPt1bSCk7siAtUBGtUZtK1Vn5K74vEdosgloZlAW
OfmLRB2u3kbmw4l1N1lnTtjigrgCEBRwrC+ZcdcPMslQEf8sYqx9mwS370Cu9DLQ2s+BaoiF2zCo
OnDxRMnE+T0R2pEX8Klfl1M3W/zYX/ZA7K9qoWO5tAlZijCz/dI65dQ3+RCPkHAsIyd8mteoEF4i
W7mp+gnN5UYH5PqDJM3znMdehBCwAcUzQ6bH0o5p4cJrjIyZjtf9/RBDasaXRxFyfFqRUaZIZkZQ
rSdj6Jw61kHfjNJ9agwxmfR+Udhqsu4UIFlQQHP1rn/+5XtANGJoKVyoKtCJEAnE+j7PDBGtJf27
8nESrMI2ZZ3TmREXjHeq00MGumo4CLUgUmPaVScOMPdJ1t6+pzH1qq7xWjdTjFf7/LckrOXr1Oi2
OfN8DVvSDDEiwZT4qsvgpInpQlLPSg2H1bV/FTXTDl76VnfXguflz0k//G3q17bxEKS/FpcQBovI
DqSW6dCUIA7jX3KBFHxBA/LRNBv1uxy18rJqRUZHbWvB7mUjcktbkfwRGA86TYTHWrQIuYFHK0ua
adJrXmMorA/5XIN+8g+7+JQPQ0Yo9zZtyCheco0IuASR1h7xo+gjGNEr5DrdYVadVHISDMrKMWZj
KR07BcR/KdSEvwZzSVXZShVuHGcjY7hoPZtOEPBa5Dq4UPItmNQiqfRLZ0EDMvvhwpMIhZN47itY
QP+vAFaG0a3uxe5GKu1qLXYF1BzNdgvSPpwXxWhIUHmPXOuOeGb6O5aLNl6WHXcyolEsjYrcqlzy
RBXkRiB6BcK6vxhQ4GrLCUTWZpxFUQqCscbS0SjeQW6aVbF7v5LNccTf30Qvpeluo/wSuQX7nrTN
Uju1e8iFSqebsOxYoHk3AJJc40SCJ/ikaru+JZxoIgJwmjzhUZRVWIdXl0RohO4kO/GgwTi0iuvf
J3a1rdr2qBdY3LcKhvKdw24CrWth+p4Y393KqS5uMHCH42Fkwzm7+R5vcoL4aW/8/PWx4/7mr7I2
PBNLlhmc8vCyMSzBCl/hK2K4aiEmKC3Eq6VgLSBDoNBiey04VRRVmqJoJTGZmXE1/KSGlWNLWgDh
Ek9FVrRg9VAp+vNRYbtjUx3G86wdJb/yybB7b2yrM8sy5cL4m/ynk4RwE3dt0dH8LRkLAs0Tx06x
kvef87atfYQuwFl6IuBckfMoaXUmfrgJ65QW+gBiwrqy7/L2QsSBIGjUFsa9VFdv9oJuRHh8H35U
J1yMliI12eJDCx0Vq7XQJWz+ota/lgeKAXArI4wJQn1KDLfdc1bqV3LdbAZcjnEbOktFEeITh+d2
rpMhWZ1AM8B3Wo+/L+D3lQzr2e7axIEIuBZfH955nB3i7dzFwPR/nKLg0Lvn3m+u/tu6zqMmeG9s
xfJdk9On8Vhj+4Bfck3n6vAQ5jLtspamHuwTL/lkt6yB7Q48pIS+zQRkFr+SzljcxLafyx3LMVML
7Dfegr9al1+37mPvCH0MVYqCaWQ/5CbGhCfxEqk0W4xjbUtlULHEXy+2vEfFgZ+O4YNQWwkUpTjg
3ltYmljb6HjL7g/i5m7JXxZNeWJS3ABS/ldg6eDWOhfhWlEeto3h16Q6bq2MzD0wrAJUZBaYPjPM
9ndb89gWYutCP2M038wL01qxZdG8nGO3ISntXR88e6S5A/Amkb2ltbRGcW2qdTPqAOmW+/LtiTt9
hmnwBaAxi1B9bUeZb3p1b0NzauHuO7y+ns4KFqxOkOzww10W0pzwBOpMYG5Kr1PjdJ2xd3dtBk6o
70h1YhAMndS+5zqqX2L+6zXgRx3Sd2y4US3Uj+eqz3aG9jYFZQ5lH1+WO8nRFc46JOU1NfgaKlSI
dOmkLcXIAdamRjh97Gv+/iTmrjduNn4jzbteuvwBlEFsMU7pjU82TldPSa9JB4r/Mn07wGbdgf8g
KEYxD2L8gqrYZLVsau4UGCOa6PVB8qof52ME1SjMDzsDwpuqIvh6U+Vs8vHbH/id8KF9+hSNWyQr
6WueeN9J2pvg8ct/HVGTppDfF8OZ6caMjzY4mdPyDwy07wUA7g4dq1KHrfUrjLwLdMLhtQ+LwVW9
ncBdJGV9PrGLxmO8BRAa7ZvV8NSaXZlNsEGv65dsAi7yyWBiU6Om/IOZ10Bow+W+9t8kMxS9FBdM
QLXDN8S6cHHE1NoucCYEx7FDDUzkbzVqmUF4GDzCECe2kpWkkaLo6/u5p3gcJ7EsKYZonrdfZhs3
JqLXPQDEVrrDsSxBWjiSt+pIPkQzJJD/77owHL9XpLInkblj8FUk+TCiaonpDRHKFOJFZAmpdW5n
MW5ZJtlUa5bHpRSVbLl0eTaQOE+ipqhd/qjYJ/Cdo9bGJcCGxe2+GXp50QNeMIXV+yHaiElscLjU
k1YDbnfHcyn1AD/r9vGinbFzQGbf36yi78AY8+qOokqfJyOUuzu/GNjaQ9P5lXvKctufc52Tib8f
G2LQfk1fX6u+DMare5GTLRbMCXTVP6S6g0KqEqns3ruYoSSRg+sBtp/HIw2W4WHhCJdipJeyWQQS
yY6RWKobER+8tojOUKb7H63NKQmDpwDqilqkSghKIctPmqW5QFg6AYL+8xf0FA5nZqBS8Y6/izBj
MDZUE+k4jXfzuY8I7XW+RXzkrBkKWtIivSsuGctHWEKORrKh7pb37VwV/r7zHPNgpDJRWitMKbf7
zLEk20F5/t4nobyQ+BKJLxodTDc/nkRt1OjwkoVGEolDSu3b/uZpeDkeUaWRsnDkOTO6C+jbOskp
USJu0nlAE/YMtL8n20WJELLNxGJwzwFiq7KkzYVAvFRaaF8TGmhRxyTllIfatufXoYZa35qLkSou
nR74gNWrIisfJR7SzJm2pVZ2D2pCXBFIO2X3maboLysDrqYto6yc9vr6ut7hwRQf7mgLihwnbd5Q
3Imz5roiso6yuFsEUmvOO6oo7oe5NLB2je+djhY+BBfYo8NHMByRCwDqiwCB1rrBQCqGvCYzeGsQ
66uH40Nc65uQiJE1ZI9buQ3nyTAFjv9wptDcKhp0CA0C4Qmzto5+hMpPu/+x9PUlOseaxBwrBvY7
y6k62zrGYCraITYLft37jTLum/g2V9a5PGx+Ro5Ll7T8RCosSAC5G1R8+3tE6X7CW98eDE9CCU8c
rlVcZ9yxhNZlGJstailwvK6Nm0E/2QC7TyVvPQZz+MAFaiwREmwgaplJFY5uSa9gaD/DA1I7mD2k
Sb4MYomvKFSWUidB2wVi/VXw/TamXiM4C7pCSEu8kkH6FpK3rJotLJ8lpp174Sj1dgQLi0VA5IBs
kmdceXrsl/OjU66dGS0IQyAp/YqHNW7D7CvAgT0M7+NNWhp6nyclMKjd20dSGs+mJw3UloB6OVnu
SQEzdNST/R+IV+JYe41AwrbafRi6IRVBYOc6ILEZFV0ipxMuT0Nnk5Ym5m+P4qTZFUxlAhXQil1c
Q9L3hleJqufCXbMTGR/dksZg2CM0wkx3szyUbRvo7UJ6N1Bv59B6VH1D4xVfnHQMIJ4Efif72e06
U9OWxe44sd9iGjaijxmY2trKs7lRhYK7F9BOjJqvVMfmUFqr+udGruUJIdLhK0P1INtLb9rrHfT8
6Sj5Gz5LpVOh1crkpGMyalaglImiQajXyLojn0MlzR+jyKo58uVgAyHTWfkne991R70igsCb2vWz
fDFe5V6UiQm+ChrekP2x0EDMuA+T6tYEBmkinCv/umL88Atpbjwjc/PGEnU8iWZDAv5eNDVFcfIR
6f8WM1d/oAqeuciEIgh3CLQpN0n+aWtPD2EI9bKOjTddgBMVtd/uwHRQ6ZQRg2tYywPIPtcTYfaT
xv4mVHl8KVqXDG/cRJTZU/rue1lg6VOdzUbM2TdS5jGCydIh3zTc7o8gcUZMzpU+ZxTl1Bb/8h+E
NkpMkl6BUVdmzANk9KlIpZzzSXDsoPFNZYzevJFYtfMjawM/AydO62i8OWURdFM50ZFKPAg7CLbw
ssX2LeL1RZHxo985nyIVPTfnMvYNN3nIxAHe6M6yvjx0mZKCIzm0YsBj21NCumUKnL2UQwMSLapM
yT257Zy1TtM57R6FmREEDrvgJlfx+HGpt8gTQ5jxHFTd27NKIOlfPMd73CMbSd/mMQjIIwKLrO0o
otjRQSBBZPI6X51X8oXo5vq/jmjq2RZr5FhhQnh6J7wvjAwB5uGKjXtdKg8D+pYlrgH05T53KwGI
m07M5Ts5VeLbOixGfxk4lUiMhDQD8e9IztgFWbloPAFyPfn35S7EVxZL6niG0HVB91QugVT2kwUy
NP8+ymCLNb8PLpD4gh5W5IMyhml3rZCNHDNmJ2HfgZ+nqz1j1ibPO0URgbWGzhwk2NpBVitkGFLU
JOI7xi2iQwVJsayi1sqLm+3BDRrb+QoNpiMvzd4eE7kVVcHwNUAiJqsbLSD6sqcXMfOEeLBxR4Cp
6Ag0WYioP8rVV+o0E5VG8T0Q1mw8TwI217BXyxa+BBmb37BhJTVgiTEsBqSFCvDKEUusQZzhhPqU
3p8tB76+ZqiNQDzJPSGBSUmTiAjTWXFkMZza0EHsNFb3uePZq118CJi87+vMsrk+8lRsgCb+1aai
drjJZlm6w2lCy3vq9CmwOX06CEqI3/FoAKhYvKuF7brvFEkGwqbDKHYUwV+qlCTebNzwfY1832/X
OconChHGOYEH3tHableuw7xQTFPDa3j3PaP8o/k0LaAlvdgHLKgak90eOIAUvnc3DFq+j8EdD+rH
j9NHUvbNytODhb0N0YBIMapsKz5q3MBMbvCRVBqIIKuiv6sUOWEEActXq03U51kS/WOSS8v7KJz8
y0BO7YoRvjWDopsPGhcjOBrE4KN+I1l6nAKv+gnH+1Oo0PpJ+V29w7Q6wxcI7Mn5XQem4gjDGqRa
X9W6uuVdPBa3UvZggkYOaYvdt5YttMCkin/boJpkCLdMTcDtvhTMoo1wCoDoYwEmT9jZq/uGTjAz
ElTK0hqCWHlGUJQPFUAPjYBV0qUcxeP2M7GXIgj4pDOZa0Fj9Gh7b0h0izsmrotwK+PVp7k1Wks5
Ym0LeK29FfNeI9R6b+Cc6EQitGljLFheY1ucqoLbBoqWbbj5RE5ZP6uBKkc7q1XOWv12W/Oop5vx
TZabjyiz5CLkdtBnoBaqmKnGprvHOTlSJRFOdh2ViaucZhG6Fq8BXdar4UqGge7Gke5AJs4qj2w+
TWtpsc16tOb93s33ORL1VJQrzy2a+VmEjSF+QD84wSxzEn0lxvTe1vPaoQRemBa1kr9fW1YS0Vck
QzvSAVdr1AAfwVjBjX4b1EiKs5zizfqc8Z1/PC/BFu6kBi3etqMhDsRsV0mR2Hw8+Wl+cV5OHDxV
wj4rn52Jz7iNKtMEaC2rDnmsHw12fGF1rcUJguqHf+Cyp6+Yrv8YcrKeAT3vJ1gGvFR6Xe5AnHAK
gVSuKodxtSw3ZHwLckG2OWKsXQmI51Pg14MWNAuvjjAWYH6TbKsVIAce3QASyxdOCQmdHS1cEq/7
RVrNB/anw0NawzKJM16nIsniWZgb7MKjs7/QsMWH3XbxpaIjI9wGXJcJKvp926HbAodyA1kZr/PO
Ck5RzdKHMLBH0v8IY/i4A6GZjMMOeip1UrIH8fqVTBZe6YJz5aANZORFP0bPxav52dr4Bak15IaV
2LBv0NNPekTQLwI811vg7Zg4ITDltRQueQkIAxUW5W1+7M6ejwqTgF7bYG6X7xt3UEHNTjj3Yglg
pD3BFejKdyZCRmu/wAu0VbytytJj3+EpHZETMsBcqa58p0TL0r2nbrarh5DPMK5qGs4UMjpZBbpH
d5O03XvrkCpgxoO8r4ZUpHbw7uwIGOLQc500iJ3K5dnAiPp9Z1YktwFa6vSl+YdnpvBIAvQ0KubH
kG5PwPpqYlnLaEt9KRfXMAfEIeojH/zWJ5Ffn1pnhAD87sGahCyCvg+MmDIU11M835VczDUiEFEn
ggzotVjOHvWde99f6O//62sYkbn8S7bs/+XDbIGtmTzOyVplkQcrSezjdnat09QBRFrucwKKgs0+
G8rbZ8306GMqQnICoFWYLdbMj4q3XbxNM9ETeooqCjLHriVODZz7qK1PwUeZ/1E5I/tj9ecyd1iN
ZP9w0UzuSURQMt7mPMjXVYpCpWq7ni92pcf1N9yjSRCS7jXNRWMMDZi8vW5pwHC1qcI09YpF9OKp
ou/3e+HML74kWdMAbeVfspTOhWTEOUeP5eSxZRd4eTcJhIIKMa39QRac38tyl5eXzjOBpt0AhzS8
7O0KbqUJbC0+imoJ8/3EA5GxBWFB1P6V2PEPk0G5DdNlKXUxXEJ50WbwY6v6BVUSWq23MsJkiw3W
sOPBNiBoMSPszVjYP5eiGsuSkJdSVTp1VocWooVXfz4X5DQBub+0gQPQj19wVKUNnKmQ22ThOUyY
/7EmeRlEZx+pbIeqJFOpTWlJfWywJRyWZT64BsK0meUqqFp4tcROlwGtPoV9wBFQxkGjawgVHifZ
ohdIrvjPMV2xKJmURZbW0GiWcLv7/KLY/AcCgaf8l1XBrflJTys0AsGWG6GxWbFrBw7MIoe5wvm2
5p6SLU00z0X3YHF/YQV61x6pefF2dopEihyZsVpoG59ncZDJK47x62XCNs8cwr0EVfsA5+9XlInY
Sw3bwpp21Be2IZnkXS5V3GjK7qpnMgi+BFAt8bY5a73klm4ZufSjOs1pkdVVJSUKvNJFGhTYFI5A
KPIUM/xBFw24cXhTOtvNd6hn/PvZoVXvtDNv+9hHFy2INY/6OHZ7hsJ6SFzVXT25WXOtGY0LCiTJ
b+WVJ/bIf9j3+hhg+5qiGuiiYeNvaGbYGMunfwOjJpep7t23OpylOlQzv+4rFI7yX8NEejhiL+Dj
p0K03hEFo22NjK1vgHn6W0DpyCOhJ5C1lciztv4gK2Te12fKs0OAKRazxPCSuhV6eGisOTqgpaGd
g8QEtRqbsAuakgzPNTUziCOIDMmhWJQ/3LGDLnqUVSML4Acu/PT4tPpG+e8QQPXxtzF96bpO/4gw
/pc8eD6fS7YQ/wh5pcnRjfCKrDjmH8dK3jRPwmJPGB5Yw9+tti0Qd7Pi6Ck6X73/LT0h6/PeL2uc
gN+4t16oS3yPWDJLsZBy/Y9Ve8g1uIpR2Vc5jEZVpmI8AAnOhmVBab81O2dDIIb9kTo8yXabjivd
Mh/CLVtScD3A4RRL0J69PhFlO9r31l/dsIbLXkQ/mXb+li/Tk9nOVcBJHRfFCJRksraYJCJn2Oy+
tKm+oDuAw52S2LXTsDWmD09/mVKKESmoKn5hmgsD6+k95mfNnYGGUe2z1imWVKY6+PmLaYITj1SL
AQD7Bvrlt5BGWGsHms3OmAfKqFvZ0AM+Q494DdSgH8/AZDWQbFSd/ZKRRCxbUeMDb3qIslQ1bUBr
0j3LnXT3XYsQ3AHggIF3eCoUaG9KjwWuvnYTebufvlWo/jnWOBUqhdGVSsYCfxngzmskcpKV5E/M
J1cyerlOmuL+KKcu0EeGDnZcM3sQrEuT4N+rQ5a6Mt4kdrgqHWe0hG4SVT17hlH+QxYJJGc2xdn+
/d5KWx0g+osJweTykzYfYDtW5KTh6pOieUOyVe+Pk5PEn9MgBNMFq4/6ZHMYYOkNFsgqOrbs0bKG
8qdAmBrJPIWT7h/XAkPLjEADoqnYlXWRGombJmp8hIR4Jy1Sg3K/81Ervu70hw9VqKvKlAB13A1h
QK3c7y6dRBoSSxJj8Cksb8c1zxAmkdx9WuU3CqMPgn2LdyrhNhFfNkM0k+05LyBwpV3mWh8fjLTz
ISyMkLQ394ryVUm1s+iqf9PI/kXr7wl4yn/q3YUwJzhpxt2IHC8i61OzDPSUX3YS2kR612/XGMZI
ZBFKBpOEj1J612zibBmj6oRR3GsSQBoXTBhW2KeH8rNJ8c0pFImHneVgDfWD+hsSSCd6GPQDEUh2
BNpkZOFEgSoj4azFlKMCqdRItqQUxsXEScTj0geQFi3fZJ+Fam+qk75Wc26AKHfqXMPwk7QbOOmY
Sn8crVcKyxuehUm2vpGOH7szsqocz2p+8B5LFTNTNzct7q4l9mRHng72NT/0Z3xoSQ35kJ8UOylP
DJNkwMFmI+OVjilHmqyVhoISnAO8TMnyVvg1hHlE7eVKvXIcj4mn/n0eJBBEUzahf5H4HAbli4hM
vmrqumczZdRNmt03fhGfeN/KoMiKWDew5N6GUwTF1ja8DHsi1KvoFFpvsjOjBUBT//HB8sXtMgvj
miez2QX4BnKoLTQztP5i9JybStPewJPwb7SvnGOseDVuNkbxCnpGnDoYZ6WNDLBp3n1mziMV2dsJ
Fc7n4q/DHym+Sqf2WqlgWnAcqBULo1oGVFGW4cM3LRFgdSuUgdDTEG4vvp0F+EIPjT/uOSNQe28a
hCIxJ7iwQ68GZ76grXz04Sd71MmT2nJ4OHjx/aPSG6bgwCaZ4pvasGDoQgpU1yes7jY/FRHQXjBM
ddVPJXg0saw/zfzwNhxw8dmCDi+D5Cg75HDKNjPKOXA9ziO2p0QDuk9DEjVZhbZiCdY+NXR4Q2C4
W0ftO/cyKvjmfueAnywh+kh+Z+SU5SdxeW2zeXxVREqtqTPprkjqfcK6f7/kvTLZ06/+kcPdvCOV
+CEltCdKs/UDDH+Wa6g090Tq6oYFTQj2TmRTOIjEeVBpKcmGlfygT75yIBRmQwfwrrl+TtqIaR67
0blrFZdlwSNldF0A3ArtLNj4df9U0YnZdBIvp6mvL/+bSfT3pHD+p9Xml08XOgCXwmocXgrvRDKG
zzv1+Q4jg/KaHvUVQpi+U+E6nbX/pbxjUzyE3K6MLKE9XFzGkOp/Gq2TsPtYxvYQx9HHUDFFiSlw
zuPlde5xfSzADJRQI2MGFZSt9DbI/cW4l+Tln2O+MbvPazRKdmRV+8xOX5TZhgjWejqPPdmRAu51
pwZs2kfF7fckuiXJ47rPDvkUC8L6E/cpKwESO+a4OA8ajUDZ78z793KlGj6gBOKE7IfY4GFantk5
r2FEWq+T4hN4ncdSw7GjMcTfQbRy/9itqW8zIYkF4GShyfvu8uuMQaOe+5f23j019SD2aHEXvI3P
MYeXUSXacM9FUfCwgsyTCcm/pmmkNJMT2MoeqJaXslwsaz2XEv0jkb01/8MeeiGsHOrqi7IAbENe
dmCqU+3VuoXqzzRhLFKdt52rH0/CfLrSw46i0Y998WqbmaRvSrLz5K0oklGGcgWnSUsaXPMMwVE1
r/nOlLORlzC2X5MMtDC9Q8mELKifjwlrIrsiuWB8DpPyc9DXXEcxnuNScfpZyGjKnNX6hxn0lpT1
f/NsvyfLMXcHsPVA/5i9n2xe9XREcGjGNN/xaauPQ3O4EO6k14ToKQcqHpMy0vhKGt1gFXT41Q3M
9E0tsd78envCFb5Ekt1gC994ygwFQyGL2INd88EMI+u+uQwO3dn1sn5ERSGN/mw6lPcO1Fq+Sp2N
Tl/2tXardUqQFuvWoMt8aeY13fKXCT/0Cbx8TL9we01viwYLIQaYiLVbk/OvtS2lEZ7RhkpuHCUd
uSGHxPAFEWBa62YFEIUmFBgeCjnV5Wn4hI40Qgky8oTcc/hNMlUVQX7OFSNPsOBzw/llPxERT8QD
WoCwzrsv/IViTPVwEmsi0lMthwWc1o+kaLXGvmQhFSn1RvSw/vIshaQKXLfhdgT5hYE7fFBhDjbs
wY3e/3V9l6bj0bru6WGaDJ/BKp+ApKaHTycxIwETsDe84Vqvpl1KLnJT/whyzqScpN4CvkZ2LyjV
jXRlJa162vb9oNg8vubMxT9eAHQLfHEVY3+bgMl0wvcHevxkeVExbb5p24PLemGIeSr/8x703sKc
mL1uqpcyow/dKDCwd6lHQmniijVWJHOoYXJwDlbv5HWhNXWHGktwUpGTW5jfQj9L6DlBp/6BGqT3
ZbjwbbqDn16aCPWfvQsoE16wbi8BgehwDQY4LPE/0HfYEAOZZzIQTjEl34AC80VCMnyb0bpvsnNm
pueod/jPBxGkyzrVek92/O2LndCA0+FSABAlya2tiboOrD7ZVqzUEx2FcbEjFN5k0Wa5qHtK8Igw
9LxgiVkOkRBkoz9aPFEGcK6+VL/RG0jro7v1m2BrMHR2AlaJBfLAQhNhORo/wxcwlPb/rSMfjKlG
UDXgwRy6rMvvf1P+c5kQYRAyj0oiqNPnEZXIvTO38htqIq8GLud/e4QQ5zISBf9RZCqNRTvxrgsg
+eY67zQix7st9Ss7gHaQy5XSen/TjwSFSfoYpsWRYlkOLMzwU9/7J2LQPIKtDTz59jBPPZnl5X5Q
m/RFzkMIH9aDQUqdeXF60TISEZLNrshUcWbXZxJnU/SgNr35mnVe7WfMQ6ebnuoe5dU4w7J3xSaY
obgRLMaVGT5UxCsVzKfUkCk4Cn3Aknbqk3GAnUXv3Jfqga7paE8k0TBrJzS79Oe9PdSDjpxlXDH3
HGiqKXRP8VrAeEj2DKJogKXNtbW/YyB4zXRPTgydJwNT/jK/wMqcqW6dytSumQxtijbHgmlxQN69
8TakiNTRX13bHv0nT+h/OXir/jhB39MUsrBwKERNs8t70eSAkV9wuK/uCFKQpGdxzhQvP/m6GSxn
wmhDSthFIkS4Zbw7bYISKr6BuOqnBXCU5Hj+bf4z9+bdhR6OLyl6o3FS7iyAgF5uNE9PfRduVoGT
bPEDm5IVMoy7KhA/qIw9pWYZcTeNzjE6Cc/yJYeAGiU40k/B2Do3W1jF6zdxfgIVUHh9xDHfs09F
tGYGMxM/inJuVUyA8Q7OSxsWJypynactFYsPfUc7xpF0BQM1lTSfw8ot+MCtDCWNOCwZUwySPAw1
vmmNw4l2WESQhPDO1H6dlzSEJKz24F8LTrlYfDFLO3msSixO72pDroiPJT+by/7Iz+/3fz+2FjIa
xWniU7wlI42m4hyV2NIMPOWhavkXO5s8kCEzIx2/h+1pgWNLxCU1JlPWDT9Z29QZL3x/H1pG0gPv
R6IebDqPETLUwjUN967wr/Butti3w3XrfsQBTJAI62SR4k61+deA9jNEF5KxzryAHym4ZAU2xLN1
fWwOZIrkQ0xfUYy3mOq/vDgQTAyjn8VqtIUtgyRMrI3eVx4voMYXRNXPe/PpPdg5UqAF0HDvr2uj
847FNHlRtnrhvJ8LcrcfIZGr4IiFhENsxsu1cPd3rsUsXdY3hCe85EIgfrOx1WBmJBQ+t6OJvw83
JHBZ9Aqyk0+QzKDGl481l5/DJXF49gpzp4X8rPiyTGvQw2+OX8T1gom3VxhaGcIdBbQZyLfy+y6W
NZu5B62h6rGCxomDwH05GdxH3i3JkjOZ0dRHiQ8VJZavkyCs2lhBYNRlkdf1JwHM1UyVV4yMUPXf
RhQWUjUlgLNfpJNFtz2Smq3zTNMBbVSAnQfJn5eHns6X+TJ/Nd7wqGcmdJZ4p6qrm4xpln/5e069
ay0a5luUNJIz3eYt5Sdkj8QS3DKxM0kP67p9XXjpqnOZO7f3zk7yphwIUyewpQKpbCGbP5IS3xn0
ZQy+P7xmuoPWDx+kC16rbemVv0+jacN2xla8PhtnWOMAwkUiU8ESkDBqqix/uhO7kNA96b5qzWql
yhwIhprZ8xBnrqZ5BsOaN/8gB6jpt8jj6WFPH/quSqAEkKCCgQ8grtPCmkBB09FYJeMIkejbf9Er
lhW4rjHyL5NwRFeVxEbNm3K876rPY0H/5JUMJepbVXbyf7JxhTSKlpprXCUJdQNR6z1B0EojbwaA
oMNMAWIwqBN4DfrhhS/3N7QBx+KQ00b2uOSR3X0l3JgXI+7FXuTy3w0c4CXGb94qZe/3GSRZo7iJ
43gBaNVlseJKxYgxQGLasRR4q1FWf/SEZCdv0thAkqzQP2o8+n3ZFCh3VAiq9SZ18Dav3XN+HLbE
z5KP4VCeVFGqhy1CzTyCGiiztYEDFVFHKKavDP29PV5vY7s8OrqErDlBT8vk/P88XSQUZ6M27vD3
hizAHoyGM7Fkj9bLdIqf6D/bQQ8ad23mWxcZaP1M9Fv+YCANSZiLtj1/RlpAvHU8WhEjUqiHzegi
aMMiStQXQt88h4X6uNcrBbSem5ao6lLNc0Zm97TZZmncRoGZeATLUwettE39HFEP+0PlHvBaPOmd
C0/UNITsSQ7fTmWmG06IUOFwWKrDHD68a6TTF/xft4elN6rFus5N2WK2YGwUwuReKs0AapsTUCnY
/yuO3EklXxZZh4M9YmS8TaiHGNK2Mu2HWe7WMR70q6fSdJIcjMMqY9PHpHfD/7jNDQEn1OiT0oXK
+UzxCzIqrQmPlDwjuqhp834GF3odJjlX9QB6lay1NHJHvAjUMhM94ry4k8OgF82+fbMLBqhcUVSX
LBJdgBhFjIWTZV1N3V1czaH7t3dtiOnIoJjJAhA5CPpiFvz5bXhqVimRoFHWtLcwkC7GMqG9GUs7
1LkkZPTko1o4G/YUYDrTLtLhls1MEAme2dV7WOBpkxI0FeB4u+/elrem9RJ5aO4rKgpP0clvO0bM
u1ZnCYaHjmebUnDGejKGWSyZsxHowrZwGmz/CbFjgIc2qPup51xxeieAWBD3rcMP9i6IH+DwKh+R
7GjprnLFQmKDZRShWXGHHCyjGGTlU2vbYD/UVtPZ4R9uLNGCoRh9cD2U+h6qYwTSP2eCpGIh2Guh
qKfP6xL22u0KeR3lQQeOwvch7YLJVJjQUt0XvvXOAqpPt0ONBoK+Z7JcABZdOtYVz96Oeo6VnD1L
buZR6lTi6exoyfKfe9hN2gEagDyloPcfVfKsvmImUyJxvetSKLYWWhfOkMYfJGZGUfp3INO2xhQu
Z2sAMm+rcj+upqs/ujH0EtEul9tVRCRRvvxtHB/JVo4ymG9eI6nJHiJlowku/5nxK7dzHWNwRYLN
yDQ1GFylzPkzIMdLvAfev8/TZi/TcDPNndsdCTpRtn7oHzJoWf0AJOLkLRURgsela/JQjaLiFbZg
g4A0CwZLejCbQt6sfEwLEBOJRs0ouliqs8Yx6dUnFxwyp0OTG7t9spEqTT8p3UFtngPVc7yCQ2/K
hlVro3geAcTgCumOJoEsybnMHpRauTlQbAO3XFujtzH3mAmWxOEVqBiJZK4iNkxSVMbiywifru87
p2/Y+lKAGSU5CyovnyN9bXfqlDTceZABxX40wJss/9zzjVxnjHwib6mzF2H+44vxD8HYAiKgB5CE
bHRbTE864JEMg6EPcq9yRwxAhoI5J1+rt2I2FXlm/uks4vXYLUlUoFcr629ns/CdsrtLj+DkT5VZ
V9Rl18unVAAUyksYrITGRYUREdmdZ3KqMY4gW00Foxvccsi2YdjLZvOEsiawUQC5wzzgmkUG4BdN
iYQRPsvDXOedQ1rdIan2UneCMxowLSWDt0/bq0az++ZuDfTKSZNNrWjVXS7Xwi/nPcFgul7zGn0K
YaGIy538RsuP4r3IuOG6Hi4ymeGjtwRfFG9sRB+y37x2tj9hlZnr92RTxBDJPE7XvbsjShu4HoqT
I25YQUnJDrQBh1b1CoXr8mJfh8ZmcDtuPZmxv8TaNOBbp9bNgBX3oILlFIuB2qpy/iE9dAYrVODw
+9gKf/GjI5hlxF/BEk1KtCzJhfTKUTlsjL8k9zxUylfbUmTWGZp9Cjp1kpfp1cE46bgpGuUZ2XWw
jV9KM5kWk8vvrEMLtN7P51zOJVYfoXYZUT4xQwhDu499mQLEn2nzPpDGBZap7DT79ZwM2BTkGE/X
ZpSQvCfJW/DLGrOQjK4DrZ1MMtx13qsVPFj3hA9ApK6hOaSnumj9cu+Ry5/riwkWPrgP63V5ElzP
RObXmGkO9TvwHGTRTaxPz6Tt9JZK1lZBrgfMuNnT6OPUUeDd0MhO84Fqv6HfF/6JbZXmXwr/Bq1b
SDOHc396uFNcrzOflU8+5LWf/rJqr/R0U8lrrXozBawfMj/02wAoQ8oTHN4aBOGNSlKvWJya3nCl
Fs4uzECRbZlYaGz/Wqll+oAi7uQoJZ0SLY3F4PEYlD/cF+qRhEZUG0TzmucW56MShrbhBLbo10+L
EPUkPZM/tr68g0eITk/64tEiK0L6p/GRk+43VVpiyh+uLVIwnG3Brrh78accuf28sU3WoVTokwib
7EK5klRa685ZUkWP//2juZvjXvoVi4rffDMNa/2CPHHtSjBiqz1MZI3hQm48yJi4qBWNKFTsf2wk
G7SGcidBHbkA0PYbKAKkPR8d5tCvYm27POtZDxd8IArfuOpkL4NnFTflg39jkryzEucC3xak6E79
N40SCFziN3O2Wwf6uQTP7ZfbRlctaGsO+hcWw2hHk3gTOkuKDHI5EdaT/XqaX2OI1LiK1foYXPs/
CqDCRaM1Kk62M94WxAch9nHPPIqjM0IOg8U1T60lGvtBQZOLi0QRn9saKl6CiBOfCOVN7yPatwuu
oclLqzSwcrXjv57UDDXjL8iAIdTIyLH2s1bLJ2gP2V4DasFILlo0UCQ/e15oK7NBeSuv/c+vKlup
02QmpHnH5Yn9fvUxoNhwH50giRvOcnD9FTkvMHc/hgyQDZMlX43YjxRk2JH8lGTKv4aLpUhsa/+u
fV5/iF5Ublv2z2ybSnipp63kgBYG++zt330y4jL90B22WyCV5AkLYixTnpGu/nehqNqXhv9VVq4u
lsA7uCHZXIeqQkeGYtKE4dCI9VR2tvI1ZWzphrfrhSAmf4JsM82dEAdrnfrBRAIjsFH1q2iTm13M
SH1VXIws2UVGqYdOhWgNvFSWl+Cg/55cUKSY5GBDlc+3R3aKeF4sQQ3ZPgXeM1ZzwnSH9vWPFEpo
J6cHBeVtWniqz4aOfjbsw/yGgIorkZGBu9T1qOBko3sTJGTS8HJnj6EYKAZwlcZyX40IkbGokYvZ
hq5jYw6Kl9J3ySBpysWdKZm3jzNsL7JdHi7QC5JpNEf7X/zpG94j3qm8OBjvf6AQXLVsaVBHXs9m
PmxopsWS+KJrfI5p2JTHItgxPFHsv71CnQv2LjnbleN+khzmpYiV2UUV9zb33aGNGDY8W5Dgokq5
+z559dG6BirCfnReB+9E8TtTGtXtZK4DOyTOgN1w7zGcHnPCYy7RibNjoLA0TF+6vie9sdObV2XW
cCWaZ2YeQE2zZBPf0QUdTz0kYuohVjMn8lIzzDjulc4GPYwot2nONZMPhhyNeUHip78VvS2VI73c
fpkY3h0DiLg6Y5WePFNHMX/8dCeiFDB3Jtgz3qYYR+b1WmVbqbdLmf3is6/Sy3/vLHxBvbe0ev5M
1wU6bGwccc+6Qt+V1wHJp7YMj6T5BoqT6pnSJIO5kg/oUmozvWfzSsiwVZVbFJX+TEQImnxlrd+6
5p+wCSRA9nSrh3H9A9WJeQB4h5SHmjTgFJHO27hau9vk0C9c5fXqCjVm5Sd9wr/Bdyuxo1/3g6IK
jvfoLNnr6h+0DLwCl8Um/bBszeyszcnzi2KviK3vdURUymBBiIC9UeAoWDkQvGsDZiTyCTPnCLp2
87NVP+Y1m8OTixHsyYPdwuWTWEJH5HEe9ZsXYgCSjnnLVSwJPxWczguVceiVkR4nBWGBx6oZMvAv
nr4A/8EPpFypMIOZ3LiRV5DiiLyW/QGliZ5EFl2JPMXi+SIMHtaVqVW2j+CirfNnbP2uNnWVh4nu
76rJBNgyZ+0p5+70JEuIXXYjHBwMA0HGBhiRV6K8PpJChdGmmik/A/dOY8dHW4/bApyEt3f+kW3l
AJ7GRRkiQnk0uoYdN5ubU3mKkjx1ViTW7ir/Es2XU9dQuhMJ79AA84+h106Z3ur7zM86D5eYfFgP
CooZg9ybrYyv8DQ8iFLoAv1UWgMJygHlq3k+pIWPbKbRk1BEFcpyRz8DGk7XATSpXs8SlLckwNVw
O5j24mNwuUp7H3HUfcsHHyLeW5mov6UaEgMKYerfab4iWOXQr3IzlYW2sWEepuZ5Tq7OiuHeSvtm
8nJCMKjo8bi0VCNKCsMw0PMVQmlds1qEEWZkqAPaumlkZfVDh+PdspVPuDK/rxMXEcZRBtBv1WmM
wJl9Fubtg9PdkVLvFmdzAnD7n9nl9hSGQP9gPsh87cS2iD7AJhgGN1wPsvQEpC633DTppUoMdYRB
NB52Ecc+zaVwEpLUY67HIwjXrMvVeKkFbxwl0DJ4YQEBFdvkuHX/ooopUdJKNnjZEt1p9aVROSUw
fLAhFSYfoJHokSmO6+mAXrnNn7yjUIOVyiOfm4WboZPjJdpWjrRrwhHBGGf2X6ptMxcaDDiPyihy
sr0+SrkFBg5yWk0lA+fbQy4x4JNwHqwHX1g7I7DGrUmq1SjORGke5ppzSPuddXLUQRknNm850qFV
kNBbTWjpTF3uaS/iVSef00PLLzLI0O2CiXYuDaJujWRk06uMaf4w9gppThISo4nA+1+fyYdgF/0s
7E6EDcivUpHL16PV4Wx5PmMl4s8VxZcB2+RCBoXfN6kVYy23E78ygu95jvgeUIXFutYMhZlC14QO
PIxd5nSPj9/p4STdmFMuC/UGX1CtaU9uNdaIN8bXDdNcQUcAER7LlSRWZVHkIdhMqr5i91KgTAuR
y7sYZnwY9ABXQMb5hJP3Sh56M5RwmHbelUyv7xPTiJUf4ZG2gQjJcToUmhH1BXIUXzPEwnlt9oQU
trlVeG5pylmsfzsNgOuGvOGnPp1F9YtsLAThd+ctZKcNYE+MUUotTey0uF8h/tnT81TIjI3hrHUt
WP0dFQlmawckYEkPC6BdJTlAdvUrngqZ5c1FPQIg8V6FJnpHeYmZFgH2Ea0fCdZzr9Sh2doZ8rwZ
A9t7denks4RmKVMCM8Ta6I3rfuDi07z+x3/wgJpONuafBKcfS9S5/Ue+A6dimP8SdRM+QpEv8tPb
qwDmA5UTn0XvH2LRDgvnyQ0mSNDLPc+jIRgh2RQO9KdwNWaBhFqNqtrPZqkq54HOczV2RG0RhDLY
oILAotyP+LXF9UplY8leUNFx4NsDzFcDv/ReU38wkBW7QJPEu6abkoxmehNd9tTIhc8xaQL2XNBx
x3wOx0o4ZWe362QNwCxjsLo1zLHbGAOuyvlZDg+WrFdK7XWAHHW2+m9rjDun0Amea/o6/Ht9L3Rp
bOXZNSfhecxGoM//U3Nuj8g94d6oBxsxrBcJ1Zbuoo1Wxx4x+ZZy+s2zo1OIQY8ZR6GmKervWayj
VKIL/WqUcbcw7EtfC0Qdv6YAflzIYSWIsLIkUJi5UwnIHm80p5fIlqjsCfTZEYbBNbv0dVWXOthc
tR33DSb6BtImPx4sPlefGvnEsgiv+OPnpVYIvfv8zn+Uy2tGr9sTBhFnNyEZTta9RCxl0Z/7RRAu
ohq5UgYxMlat+Th3UJh8omIXSaylTuM+LKdLgN6FiNaVvYl6K5mxW1CvM9bVTRHYZ1NR6xKvs7jn
+0SDFQytDM0eDGeAziGrJrg33exubyqS2rG8aJQ4TOZPqnn/vy6XvaRiSE3GoUcTCCpCpV9YFG9v
9RHzXsDphH/TNFh/C3/sCTL1SU/m9b8q1R9udU6fGY63MTt+PphI8gwOjx0mbrPn9DT8KO5FCt/F
WDFboZNQ2YdVfdToObK+KKoqqZlZR/ygct+osd12/DjdecHLdnu1MvAaGB5/DPeqtxDcZf0CN6RR
utKTdarVQ7OBVSxQRH/lWTu/WfQWe1FWk/ICaWVuBcffkQ7FJ/s2MNQZm3fnGcVLqglI0GXmjuXY
AeAkYQ5WanqFJh9rKpTIKCLrz1/CXlW2hgvoIw5XxkwOwjcd2c2ua4UllrU6+9iraUYYWehkUL0r
sLNbYz9Y5t48Hno0icWKwFKF5gJbz/ZXRGiC0TC8zxximXhxzFp2kjH4k7+8uQu1f7gL7RxtiTKd
m5paf50hF7KOsvPgfIpnX2QldosqH0CF2Hz772TJN+yAxpC18BTYvszM7zkF/GNSsr6um6CRE5mw
sWejv6W18/LXIFM408VUTkRW3rpuV3JhT0kO/PFn1Etq6A7RbZ9v47Hp33VucLiebbZ1V1ylGWJg
mASuBuStlkK8nnyhQPXdP3MYDYnW6d1iKAlrcWrv7fk3iH0EU0ytviYLbjoOJLUTHiPhvgF6C3HV
xiB72ham76E83SIR0+lZf4l+/MIxKBus4rrYw9ScPPjcgQeOHDJeWm54tVQ0SzFLpmj68y+N0dQD
rFzo54x5ima02pHmC43QbqEAJqDldqd3c8P/zhSrA7zrWLYI6jYx6xAY6/MwkmA9fRZRgkw+qzLh
R5j1QwHf/4+8qsvpHjSy/0Q7paYk/MfFDLjSuiQsEwqJWrtJw8Vj+PI48oDKe+yzig17+Ar1gvT0
iS5mcouRsk0srhy/Ii8MXAr6+D3I4m/Qq7H3XPaHERZqSjWi2zXsE20AdsthxAgbvHarPlgNG02W
SU2fDlS68WGHIx4vQXmOK4qUbspfR0yn40Bz43RZgkc4/9jlTfdxTIvEKJDVKmPtW3WrLXJWN4K1
jxIz1fG8EMKPfXoZzqp5uV5afskNKw53PorRnidRZU8shs5w5e5lj32as4T8ki3dgCpTDtoUE/6D
cL84zCHmOpyS6el7RCFV0l7Fc0fGzrFhyn45lHXhSDMmH2FsUVOoMDkoeyPxl9+cNHYE1iDFNjsL
62m9m5j0o8CSiA0IZcRJqI5wMftwoXdOZH59ZfbaQQmklRE2RIWIOZI1IrbS+xrUzOZhaLFcR2fH
1/G6eOBawox+i6X9ylrJg2mD918YOQZqYAv9rSaQfdftOxxOtxEudSu/XOZw0zeG07pZ27UjjSgq
ZHKaKKkBOceJjIE0+HJXNSi8edI2p9Zeiwh50X5Nh7Vz8mK+ADttQ3ywhmS0S/8njAughYJvy4i0
Bj1RZHBBCcKwvTqoHasWL49zWNqdAcmywK4FSKalkEv59S66PZHFs7FwZ6MNC/jx5+UFwcp0cGpb
kyj1n3026cwGIhQdpG/pZO519Tf4EDd7jfbCcpzIRPtAh/SBMTmrKOwS3YlEEaVlDbHwBJvkshcB
xMxLi8b2GSH1lX5yuLsTqdrkH7T6yFHM81QXgPn8hb6nznkmVhi1jNnwo1krNhe8rvffBaaSREyy
a4mpdDWTc11pUWbYtpcUxW+L66E90278XeunGW9iMkk9drwmzOYdsjdHs0q0ZnUX7mYRAMoPmnG0
ggI+6RT+n2Tgt8BUD4wSFfEtZk3tynRp+ewGjO+TWaRdEmJzbTCMYEoSPRkLeibQFVgxDEkU/j/W
qGk2DzPsIKVoebe4hpghflhx65lQ8Bag1AycvuWS28kqPK5NfUWDXaZXsjlpLMFwNlIoLs/Dx2XV
patidZtHSSFVuea7CipaVKb5Kz5/GbtXVQmqqo+v4bGWY67P4/CL8LUkIGzQRkFmwxUEyeHy/9Sa
VvkMh/4WJHPU8GWWgmnmPmD25tzD6CFH2k7Zr0133eXBJCosmYPb4GBpaWfAKx8FcherHOtqfJd2
p4aWU1dgNQGEQplmwcgld2efFv+g3tAOfx2PRiUv5niCAYDgWjN47dJW5PguMfWanEmrmANW9iRj
pM9TIOVpOUV8jBg6NLNeWu09O/Giu20jZdtOWNlDf8lvzntun/36Qm1WJjuxH8HCBMSOs7MkDp8J
lA+GKN/iGapoTWk66YfopHZGo5abnrkdiBK3LqSd1zb59oMYUaNanD0SoPzuvTapPBfXUwBdDpiK
QwRtJRKPsiq3zjyucvIACH6jwyUTITLwSH76e+AN/GPxCu7hc4CXVoELn+Yjd+n5579hq2YOvkqc
SuqwLGHZFoF2OnnSj7smolbaMlDwPKd20F/+Q7dmp0+0/xHv4ogOkYayqCCea7TuC3cnkCuHN0TU
1qPh5gHoG73VL2CGdxevxGkKhNwX6pfLRDWXTcROkVehJnlfby4SbXdwcRd3iZwD59D3ITfKYmEw
E2bRbzqFTvvVwjX3TQe3FBnKcitwCBfkLcBHbQVWCg1BxaeTt6RuCAyrRSugD8WDJ6HDn8/aBBdy
mEnpkz08GgprvN40/GDtgbLuWy6mQ74jw4X31SWHaJJ3xGzKz6hgdn5r4AJCsXniKdDQXwExtNhX
h8hD9/XzKeuG3HhLB9fVlicswdELxNbjiJvlBbEsgbc+UCCtufPax5gUUVBRgHH+1Yf+FbGOkOaN
K4BOEOoJt2tsCWvBeU6iC6dbfsTkg+bX4dmfiF6lpDLNp72O8p/Nd+ZGCK590ysvj+I+NPvOrFI+
JySoj7ZS5/Exeo/UBNzj2B7o8txHqtbpJo9s4Oer/FAzpPA5F0yyLxIv0bYpb32u1G6c026zmT93
3ej7y8c6ou2Xo6XxdyIWUM7o2bmVVo6n5D84bvzfyYfA9hUVVfIxg1l983QITX/TxiHXMfwQ6/je
BcP8vNA1KOdeRfvq3R1qtRLC80n2mnKxtf2h+r8lTLrK3k7kaFfFf+i7+CrSJ3rFxyKw9iZt8i/J
YdVN3j53h0+fCD+t7Tdd8Enw5trF9iZqplDvJ5ua59BaV3Y+YGRMib/GmTRJb9b1VeBKh+xp3uhh
Q/3n+b54+JCJuImqH+QrCZc44Aba8HE3xh+rRwjChVEfyepX12tVDgAQzHr4joRE/RrDEjEjSDT2
Kw7h32msakGeYGc5Y/wqnbcnz8IXe4aOush2G3BwJbzY1I92YVZj1HiBenk+mZ7+YHYpKuoanAiJ
BdOCCihw17MJkdIsr8APGeRwCYX8vLX1O3s0ww6D1JjbXZ1s/rdWoZ0GtI7JSyFZRtUrYRySe5Uv
54wQ+/QbBQoZO2cfXK8mO1+/OwvjOvtbWtFZuYyRbZMPKSAUwh8ZrmhNEFEYw+uSQbulBiQqUPc5
o2L7N2aMFEbcFYV+ekp5p8Lzl5SE+Qrd45fkTgVkDb1JX0p+4hn0H67vPu2kA8/viMyzZZawsUyK
UBY4UqxLpc1b9gUHqGjJgHWwEzMHR9OevSV/5jky7lVi1J4eyx2e9mDZ9wgKtU1Euh43ruwyhCIf
7OcebB36R+BDewKjmwS42GoSeI+uKlpa0xNUfHKmGr3bLPaiGIoa5WY4pbopeY9Ru7OgCyTFBWPt
z5Y1EYErzVu+46CnltgyXwe0rAy8pS1JXb/9wtC4QF8whDPRcGk2FMsTa1GsBAJEz07NIIfipeNo
udDPcoTxTB0dBO8zpK6naEWNy7mw3y9rzDHGuN2ChKrF7NuTCv3W2UPeOud0dCtFLpxDw4pgrEK7
94VeNL9hW3OFHYJFf+v0D9AoHUO1RCA0/81Y281QBY8f6wf1A2FyuH+2SO/MV+zlKfUzi9wTC90+
hvibmr5hRY6s40q4EkPyFfF7AK9VjW4z8b8+STgmZ146sVq84pdWT4g2mPRfRWv4tnJp4q4+qh8Q
MrIJHoybBGRjK9HDshlCILmX6Xf0N5dNhwnRowYBusRRg5FTjVEarUMfroUkNPR2Rc2MHBCDKKL7
Z6IQjqz5wXBaSnIvJ2/xTO7Ivpy1LxF2mk5u5Gr15fL3ctqiptPAWHwUtHxIU2eU15d1Cwx/YMza
e/3KbBYDIlyAHYRcdv4A/j5fa6SvhuDvCaxedEX5VogFcyZSgCyX877vGw6rA7kS/qEqLuaoE2iT
tcyRfTx85yDyOi1Wk+ptt5Z7jLd2qAQLG8sipCrG832BXK698WAJRjhUbp/0FJintC21UuabmEkz
22BMcQDdu5bxslBj7ta/vzfqJxzZ8Nnz9JogfMej/+/rH58gyUjMNCA1olLwUkD9ooRRAmixwprr
/BEFyf0QzqBQhQmKTSi18zTIsvjgd0u8FPsVrqxFfRoP+VYxntJVoRt1vnACf2K7StAQVl0J6HIB
w1sq0WSq6etjt2pev4aHblSDtdW7DObLbQCj4VmBkOjL+XNZb0/A6KcNMCw18o3ZBVtsIfSzUt6W
Y1Jk783InBnol/EqKb0aS+qd0C6Scdz79bVZOOg1a9DuzonAp67UCGo+W1C1INQuxqwaeKGQRC1u
4WM+Wd4DqmpegtwIui8ZKkhxR64jMFI1JbHqR/bHu5eZtLH5PTV+CdHD1vOeai920Px8BNGNkRnK
axfOGGQU4/Jb4LsP0x8aBHVNV/XBpI/MCqi01KkjC7YzlGwzTR+znN6I7FPgVhpmEp2kGxVgD776
6puzDcTDpejCia6H7Ew6G/loXqyBSWSdo1pBkRpOwjstsyEcsqz8hFHP3VAuCuKwVij6e6dSduZR
xRndA4Y8eQOiy9cftjxOWVp57yxiR6Z9e/s5VmOlAkjOUuCKcNEGpNcUnlcHioONvW3iUV6+jEfJ
P6Rn8Jh25mpc1x5Hw31MtoXepLx4wnkLobHY9Og0iJPj/Rti2xUKjwYay8vPw/+gjwPiBq/y+vM6
JPlevCyONpLTqh296s+z+9w5Q/c3oPvK0iILoUewouAIMlCz5OFrrrktf2zXhUuaN/DYIMKVX7Dp
A/RdELS/hvzUyDmdl34LtY37T2dbdDHOrCgjpnsEKTdJkYD9v9GxrbnT6urP6dVHOBM6kX2r65gn
3UkeohhIEscje1mEBkwvqvNFXK/7ZQWl1jidutq9GXHh+3s7eaYBd8mWcgzkaxF6g2mqkuP5tzfD
ekY4xg0iWW1JpkT34d1SZLmz/yMrwW3JY6TEiEweh2x/3OnUGapLKhhepO7kWT/RN+WXsYPxSkHJ
GYhd4Oc2ATtLxtTIwFeETS50U1m5Wp0ZxZSqg3EwIl4susDG3Da9cssyMU+vi4sqgncZH3b8V2Bv
1TePbRwA3iTQg0hJs7DDPV1xkEbpPfcPg7p+19hgmr80BXnWTSY7EuqyU2IneKJbL7KUP1lr4076
Zmz5ofTvF8UIhXRz+wcUwoti24grgD00Xg57e/MlHNG8LtICSOnAGlKBZsSXIQxF6z82/CkZ8ufZ
JD6vpA+/J6gsRG7W6s2j+Z5KQVLQuApZXhzvjzxG95Ort+8MHQE8FU0Y018rkR6XoHmXmqh0qbWS
bb3OpbcS3ifiJR2OvsqqjCTJEPR+gN3+EX8eLG0mdZgJKCqc2HqFkw7+ZgUsbacYyS9k81Jm57EY
Qicr7qOkNF1eFIh41K8nKquoUb+qxQ3rmSzgS9Ro+lvEvdVA7tjnbONDXzXdOIM29pdjKhkt+xtW
leD6ctwUlwoi2OCGyv88I4VbhAzfSv49JK9ZVHlF5lZF3mFzBoBon1dfzrXI+hHIQWqFpcYlcyP8
Y1Mj9GQDGfWjrvnm9iBaxnIkNPul4dOtrM9X65+BV6a3aUPnkksdE1Wm48+Xl7EMufhuD0Nnn84j
GUEM5Nm1zaQTthsGfDF2t3nJNPT006oOa///6qjknO2mWjSQhEGiBWBxCPObLgM6speN7rT0b+iO
8JaZbm2zlRFDa5dKdUJufYDsVzrzs7ZIFWGmVKiihGUtUuy1UpW4n3oSZJ23Ib9GnNvPC/Oewxg9
hpmBMB/9sZ2BkTmuj7WoBs11H39WRNx9yzZC0g6Cwt6xy06can5JgiBEHMUUPClX5tLW29HdFjQu
FWpmr8KVNZjhATw846IAZ/C8aWcHq67xwiyDLcgDL8qk+NVUjaHzXO68qNAUDiFqvdR2L1K3PBgZ
sPxgBAyMBUNSySjoeH0EAnI8wG+pP4gRnQ+VYMSx/ocRDWLc9hyWM/k4LqRAA6CfV8vpepycvIkq
OUXwnuptSsesk6WI+8Uls9On8GxLtlvjz1I70Rr9CRhvV6KuCU5wL8V3uA2IPxpjL+J7NdSLN6ls
2jjoc1SPYWtq11orH/uNSTYHNbap9nqwBepRS9Siz8ND6doXxw0A67tHeWTat+wNNC7dRzvKuWkN
1H6st1c0hGP4q5echjNJhrsIi7XWLYBXPjd7tAXcyxPJOGN0vmGJO/3p/ZvKQBIQ/BYX46KOl9VE
uRjIpFEa6Q0qXrVhO7mP7/TZqn2SxoSJOyg5ZxOpSUpNBzY1eii5fMW604AH4rFlvu0KXXLWxd3s
PugWfqt0bsYuMGhuqg8/WYtr6f04Im2XPgww7a8gL3LmwbWHsXTLwhdnIECMA/RU5cCHwWhe5Nml
u/zG0So+dQmOrHP0cjWatPXIu9fu1AAVrJxC7LDGoRL89vXcXsChfyWYPkHDhbb940Wp/Mz44RGj
ejbpPODziVyrrpu6i55nSQ1oMiyKjlWsnw89R/hfPQxU6PKMKFYZY2LOcqCBY/RtzSZhEipAjGL5
FLwGCatnUW5+laYuPcEPAGG796bp6FQE0+Fcwjg4TC1ajTXktoRTJRBberwJxIv9QB8k7sgzNT4J
NLFfybJHpknRpzmo3HKxgQpD5NPQOvrCT6sj6rKMtmJ5J1/S7RUZZNs38BDduDnyvxABb6RtFmsK
PeaWxdB7aG1BJFvGCx29rI/J58murD8Kga6CBnh594i2SpFoXf+gYpZx7K2LgKjHBCaXXoIvQCSX
qX0qG9ae+FbFTHnVwOXa5P1Lf3X+Bd1HughkvLycBwJWKbobcIbG4rCgrdKg/XGgoA3UuAYV7Cn9
rW0yn8cJ13/k19Ry/OAvemJeNZnIvdgrBbJwmyFLkYnpz2vjX4Fr5z/x7IoLmaeQzmkR4dVneUgB
jet7rEU5mvOKBHzR+2+ncBqjc6MQDtUcQXiBiAelZVIqVAb1zFmmiOPwiTdtDKv8gBx7cGutgRJe
pysfIRBdtJ8sCHi+W+oCSdoTspRiEj3L9DLYjSs9SBbbXK+BTjoUgXU6eUnqKkyC9v0wc192a9Ho
TRvseiEwste5ommhealfdd4ZryJaRAKHijR9F4mFEDI57zpf5Rvm+BsuPex6kLMJsvWcQH2YBl1z
UMNYyb/WVu6RJR4GLtMG0aKn3Xz1BgZNqUmz+G8q+A0MHaykOlpXcBvJ8RQVqB2EXmbJet9od3m1
h+l/nCjuxOzaggrfOvADaTil+SI+emLrVes4gQXTlqCwybpuYQZVBXKfXd2bzhPmXRR/dXP8Y7ak
JcVI98WthIligREpecMLOy8lj4B8LUdtrpvKwRQ5aekf2iZl4p/QAJJQvgs1Ifyse8LKleXI2D4R
4BmEz0VZ5om9hRLn9tYUfIl48PhPDZ+/EMwTBRuvHdSgIdomPOos8PA6dW9dq+vDC2lGAFqw4BXe
1PgDJelRC879oBGNb0wyWVfbWYAkwWjSPO0KA9t68VnTrcb7hGZMNWtRGj87kQjh18m8ILYQWPZc
OFadj0IqdzY7bDspjcEzeWedAyzRbVcIA5Pe7/Gzh2UXXHiCjFt1HvwvNG3fuDTX/SufjnMF7YnB
j7tZlzHQbIoTK0DpN1K0NcTKqD2y+jKE0BWjDLRzx00ajjvgo0BXuy5FhjbEfezVUPHk72O/PXG2
f4hGLIgGakYHGNd14PFqhkGyp/rHBIyP0EQYjfEOcZpgbjxnq7Mrq/7SAtHH8IXJzGkcO7bJnK7l
8nu0rcPb9utU04va8mK3BwEGFfRfxud7PYdjOO4WahiD0guECQ7tTYGoGsk2DdPXWse/mrPrOx/r
qNx2az5f35LmeX4rMwSFvO7/MvMI2w916n6SB9CDjp2hdRxw9cowTSDWZfK9E8VY0JaEV8J6TpGN
6+hB87PFOfPVQKT82jNheh7O23AzKkahBk9xaXoOYKNFEieWGSgoka+yVfX1FIlW4CzL9rCyWzjA
o0ngxPJNoVUIIYL6ApoGVLCq+KyWLp8Xf5QqQLuK+mJSPu51cUZmjfunDnzu3tI5TSG+k73iRXkx
qGcKoqQ7bI5D8ce1RGHJmXv64kNpQYE3Qy15/OLx51v3YFwAf2nulPNM6M/Wuqr0IqyR7JOkUcGd
7PxY+94OiYt/qgtcAZLPNo5jkZjyUXOxxLNQv5slri9IjlanD2HTjdS7A05ogUm/flY6Y6qzHdRF
fo7kMfe7zaz1vuYAKDuxwqbaEqtKJd1+PjnJffEqf5HfAHX53ZbJW3LqDOkTBl8VvQohWmXhXCV6
qB/FTxqRThBVatXyzCgGBJ7jS1unrNbxythwaMDcIq9Cc+kF8WlFE1t6dPQGYGWFR3263EIZqKIY
YqndK3de7M8prRj9BwKvotn3g3yDAL7yjcz2d0sdBGZ3pbApivjBYMzFWmAg3V3MTaz1miuW1DMm
yFu5PrjeMCyVStLyUG+z6WHNIwWOZVJKMJy4N0HQlaOf2fA4NTKqf4xCYJx2rtOOlGbgMpyOEnq/
/oB2W/1lhLoIxkqxybdAY+jC3LAVDXXKeT9rP3vyHdz+w7pPDt9uLTAAmxEP66YBzS+gWv+aZcyq
vPXLiKaO8eddjXxQukCsmxQ/yVjDtED+fVqYFg9gVfJMae5xAXky4bRb6tBBNKf5q34mpVUsjxOd
u+gHulFtzzvW7uPkjxx7cj/CXF98hpl1LIxQYsUznvTtO6proM1UFxv4q9dnMnbe/4huH4q+22dn
K0oQ9ICFh2X3BB41L3IL1inwtIzTLjngmnZBxdYs8KAm3MXiL2BBH8mh/3kG8DdO88QgYkw0lMYD
hIuJr2T0GvcvKAxWynlNzY8MgCsHqHioRMs0H1wHUBImhQ4rhaYZMv3I3psaVlTkcwubAlrXkkcl
iXG7tK73ZD8Sg2n1TiskaA4OXWTe7LooS3wjHIsmj4P4cZEXmVd+i8KCKdxto+gmrcI6PYlp7uDU
k7AxIPHSBwqE/tdoO4fH4hgPxiWnFZwcKxTTjeVFCe0c1du5Eezx/CJ2B7istDxP5aDg8rS9/tgS
fFzhy/IezRbKx2KNuO7x8n/vqc0zsbyJQ27+5HU/qJc/jEpV2WfpI8o/tPm/gRMmSbrDGDGkByN7
x+1EslOu4YUmUP8pA3xkPyzstgO+BZ/N2VGYojuBAFeWVsrtVsccPqG4m6xaYpMEtFmo3TltP5Gq
So3sAKWSnj5WQC1Tc7giPx8a5JOAZnFH9VQLg/UfoXEyFuXeOf/bjsuJ8WhXoBv9PlVzy9rCsDu9
/DtZUnP2kXNVwmx1Oe5aEb7sfiNSi7XLS8tF2utB+P6Ybi5jiktAyyAVtIcyq0osxQOplz9tHRBx
s9NhJjNAB6esLqEAhnrD+/qt2jMHd1A2M34zRtMR01jYtEyaifldnyY/B7PSVsoAkz3HXDE6Krqr
Wer8e32a9CLbH+fagXeq8cyYgwiOb7bChVJ04/W9EwASd+RsIPTBDcBBr/3jJA6XUPmZsSLkQVLc
ScUhMY3urENV8e312UV0Zcc8/dSZGdauJUxvM6fB3tiHnnzGLib//YwxLP2FdNIZZg4jP+zE9isb
YkYQpkS1SDFwceEie/x2oEyZkc4ndKPr4S15jBC8LWeWBHVCs32ieAS3wo1ziDl3BZ/YbW5qwcSS
7WcWwsDxVKTVVZk57no/nGodaBJiw7QItm3o5WuL5BLjeMuH7uribCpxMub8OYiK3+plE9hAwvzK
F5VZxDoMJwGW65W07uA/goWZH5mON82X+TD5r3FwSsh//4q92dz0BoILSM4IoRhTpNVZn0Z3Zhn9
e6165qwe9RJ60d5RX2wEqNo8F8MmqChlGFG//Ng/tLxatRWi2E5ZUte1Hiyw2Fmi/BTdgqooRrvN
d3/7/GdBQ60CTY7bZMOazi1fFHwkWdHByiwAB8dv8AIqf1rv/WF6EQ/j8U4g5qwhcsvBw85ON3cp
muTVJKDeA/NcjmqJU2e5ynFCwb+iuU3P8TLn5p2i1XRJL7qjYxZVE+qyDs1neda8r4bdcfuvTAhQ
W818mYF9xodjHq7u6u5cFIpVrS5DrexUIBT50ie6HkVXHDQAy0OHRLs5Ql0OOUjyI+JJMA5hvrhT
MAHvm62Lq6jSz1HOwGHWQWEa2w5jwUwEJlfROddfeRWKYUTqz5tW0hKeJl134OX22OYqFzxnBmyF
xs3gGCgwC7RYcRtSSH6O7R1eMzxvskzGn2sl5E3gegGqdGWCnyZywKg0yZ/ttz3wR9vpJaPp5Fad
gkak03fO6EUPhLioQao9UKQUDXUfCdB86dw0PExDgpEJ1bM+irUEhg5NfULR3IiwD3IfZocqOoSj
YaolRpQyxSDGiuqYFPFxxYFgpsVei2HSrAqIILv4+mfjHkLXxSxzj5fs7ijX5b47IixU/yZoQc0Q
SQqSKaaK4vxQ5gbAPkPvSgHtaOoktavnVur1ueChjznjMQ7C2Waz91HGoySBdD+oHWKa5m+Ipkxi
6qJCASXi+tGNmcst8NaNV81H41Yg/pQMi+CVEvXyoAqUHf8C+vD9Vav6SaAvbY7w+MCduVoBHo9y
VC/Z2yXuKnLYzvYGipkaRrmc9OOF7PZfXhlYu4f3M49RY2CwEnW7yHgCHojGxLGiB0f1a9cdQ0by
mcqU7hwWEymSQyZr73kqKKshXAbAjbyqP0amJ/6ANWtAy+w5jegD2S5uvHoF2qISjkiLI63lvyej
DO6MWu6JHk7RRFA0dIhxloR3iUMe1UASzRHoBjPZLAe2/hB8QlcXisf1I1vnqFXY3DXdAQeMscZ4
k1Z53K/c5ITJ+Nja7i1qqFKOr0zElXSyCQJdgK+kG0Oen5AtSF/kb3Pkq67u4cY6p921iopyTYHK
veG95Ho+p9dcpWe8ZJ6zTktlgezlAHp01+quGCPClO+FpCDJhaSH7H7aCXH76AYM+0ixW8p5u5IY
EiI8jRZaLnpbhmqDgChn/wAyxYHF1akmJB7gJhEVFJTLz3d3737x9bpZVfl7XDZB+HrivruvqOHa
bKx31yD9CBbD+z+xk/s+EESOFRqaTtFzmFtXwB/Z5xL4nFxknA9qnB8/4CaZQCBKkDPdU3kXuHs2
SwJovTTl24M9YkvhOKwSPf4yBJsryYkZhEml8kiLqS5sujHGClHg8RXBF0zHgUx1XrweFPUJJWBj
R56xIoyuzwpXVx0MD4xxpTaOnzE6b6s4xsMeW19QVzx2btwK/Z8Q+59Vxe5EWPw2C4V6F+Gv9tlS
MUilyQtizjMZOcNQTtgq8gbIaCd8Ba3go6L1K2Z2yYVIXaEFDlyvdhihMeYAZEzIJ1FNU+dKr2jA
441S7Jpe6jk9m7BX7dVIK4QTmj5D2ZALUyD+29sDpmZ+p/y3F+4E75splBnSnkAtBeb2yMX7hen8
NHF4GOUE2CjrJWcqGUQwFqqLkKu46DOXjwQej4roTRLEKhR1yZE8C1o7N3G6xO+FMASw7YqJjkNW
NL6D4d85x/ZZo/EzAwH6zshKv/cHqC+7kHLqNwMR7xvV5AoeGFuC/zCWracaYwXuZSnCCC4rHU4P
qWYz6EAyT0qZi7jBGdOo74XsbsjvFugz5zFFBxwmafBcbC4dM9jP7ZEpKX9Kk28TM+JD0hBULp2Q
jfJUllZ25aLYJL8+SgvRF6iQkW447rPRM8xg5QGe8+Jl59RIb4LnyS8EVnHbxYAV6v31YzutUnaT
TQXxBVHpG+xr9riL/k2vi1dhAMccBW9tY61o1Tf0QD9EbKSvvZvIW6LaMzsIauiBoqkXMZJ2lMh3
dsyZnMcN2Ndwgnk1WggrqM55v46a1L2tPxLJvzZvPrTIJKJJeqtsEndlG3oiqrpgpb1G3ycVKFxQ
KR1HDXtqSVMitcmr1lc7yP1IEWRvwFylgS44NYQptvnEIqLsz7PdU0Bc2t0pJ/KG0f01a6rfon5Q
HoGNJsLnC9zXGgmYMM/O4jybGjt6o1a1iQ8orOZRQ8WPK2xqNJItdJRQ4hXmjv8eKpy/E1Lk80xp
zv5K2Yd+5OoL7RcKDypd8Qf8hBTe4JxZQTHuL7oY5PcHnMLAiqQNdWKID9BCbt71bpqT6ojWERus
rGY8WZYl/5nkZq5jeiYhSNqt6mJJ3OPsH9Mk9vSFYv7LHQH6UeSOwq7wKQhUOgw8fzZek5deIVZ1
qfBUUBgSxwqKyjCs8ERMFFjuvztIGqXGMs96YdAxS/3ME6SFrgCltA5r4Jmc1rY8w6JxZ6LHGDLZ
1cMQvKDpLGHSPFj7zJ/Z8V0Y4pTR0uOwwrDOtIEmpz05VHMCnRdmBfnmJHcqhBqlPMLn7aVDT+Yc
n6kIdAJeoXbTs9I2g7KNYXze1WL1Ojl7Ob9TP5qyZg5bDI+ZBXcdJbxdjus+OJbbJXNKZzZKyk45
k8fMFv0eR68aqbCgGbj/BPABwa0Th+NODlXkvSxRCbcKkBr40R+FfizKb0YFtfCwDywcfnVORBtq
d+PMLz3CmdE3xWPoAbogo8ooRWPBsCi+jLbUzs+7TU5UiFK5gPvRIAnmh13BDWZCLtJ1tJcV6jjs
DeIQriZBPvwFKqTIOLVTsqQYcj+tiA0OVDH7yN1vAKToLIPQMs7PEMFtJKT380jN5Ttpf7yzPyZ1
T1pH18pK2CiOqaS/h+h8oBweMom0cqb9wPEPHl+Yk5feSw6I465nbxwxmQE/bX1DlabKNcAiWDCG
UYDmwbZRkyoZMgmKKTaVRUL92wygGnWHRAJQ+vE0p+2UEQqS9WDwiMXJvsT69CodStK2Ew0sD551
ZPrT89CIKHwmCgGAxY1dXGbJFHrKRZokOOXHbSRF4+8n9q2gSGjgYg7aqr1pRc90vQRm2a+7qB8p
DgD8RIHRJYM7N537yl7ph7axv/9e2Ye5rKHV0GwYWfgOHimWuo0LhfaoMgjFls152n9KYKRPLanW
exDPcThm4h7GHkpIkxYQMpliwWqo1WVdccwPCsODlWGl4x0zsICQDrI4Na+w7396xkzbLpGRGryQ
sYkYQVMAzJp8b510lmGFvCdvcphSLtgzhSTiBSArpHgph9cg0FQjHeLFLohfVBDiKLIZlckbz7+w
XxErAK17IKwZIf/jqODfHTvHHhkJ79wKiyc8sWsDKLx/80AcjE8VHBcvec8HpLRYzmGF1WP69nPp
+9+4vX5SHM48Pa/qXvLNVXHs0nciq4cgnC8MXrgZiNzjP7nluxNAGjWbsWXayNMhfHrlucXU7cES
y2i1ibiJ9eJfo2Gu8683SJmRGUfWGUJM3+53bdiUrRoFYjy9hIOCdIyh/r/c8E1T7EKLYCe2D1xs
f6TZJem2nw5pw6EiLXZuwNBEDQpSYmkEujqnh/x++avz/ieVgPTW7zP/2XH7T9NahvTY1r0hPUiO
JIJYXrqWXLvrOvO/lBnj2CKzXcjRcU1e5/qIyUuhuo2xx3SVXJsE6iVGfTOX8W96qIh3vcrW8Adu
iweO+e06FFwy/AL8H+LZQP3FboFzOjieI505VHQEbJrdLeTlEf98YryFsTOxXTWvP8sR34Kh/dxm
x68qeGscGygko5qBTdn+TKopzc/lwjSOWTggcv1T0FTSmf3YvziejHbHnFzpkEOrBF/az9p//cb/
ryYuNNBwBRHoawMFbZx/aDnfmW3OLJsjoIWB2FX3NBC07ozpkLEGRpMjNvzrbxqUFLAs7LoJIRJF
KD2UEVkvPgnnJB3t0DJIwjiK1sqBRq5UQeubL2U4rSlSzUmK6yoIYM4eSxSmZMZH0lFt5DQEHccP
vc66Jyk4b84e3ycMcCaEM8cQk9nqzZ+kUIt2azhhJbn5Th/HPrpE6aaNEkVgpKrFR6MjUgw6v31h
22regJF7Bo4zajymaImbbH2u8SSSufHi+1knK9TjF05Zu0XCJ32w6KSKoA8fqjGFBcjHR6IhoSiR
g4GTDE7gCLnHNkf/n9v+MLEOPG7rkpwus+s7iOwIerc7SPi1Lw68UI64UtWZUhNXIIKS0ploOVLE
Uzb2JpQ1XNHwz6IcL2dUSn6rrWfWWStBwxFBwOYmnillgDtVJxvQo0LCvfbLLtW9ANuKn942mayA
MSyTFu0lwjCRfbCRR6/GBuM6F+Sjct3jzKEYrKcMyob+0M8Mjp3ZDuIwRMm80ljMsB8+Zhupzkf7
G52xK/WFb3zzDD7Gy5gSiJLfYEgCojj+74Llhi3dbczUb4+etQ1BQROQ0aUHM02MqPVHDfTrx1Aq
h/E8bRNn02+1LcRorEfBj3DXaYno4207livJh/08QqdqH1fwM3MxlDt04woiez46z7yYj0P6JrRp
sQaK4oZ/g71to8XcDjavu7JqmIMAt65Lh9dpKgIBb6PHq6M/5boY92VPAZJZo0b6dsL+haEGMmUr
8mseNxN6NF3+CylZ7i3uepQAj1k10IClWXBx4TEhZ3kPK9e8nHvjHK0NPsN/VnFJSJhjy0UvRHc2
qvpjW4IgPD4HO/U05b+kDYQBBGjztWEtn7DLQE6mcfAQmLXzLB8y5GHqO+DO1OK761jKpK3GLI0t
5ba8zlhuaznm2V+0La0BpYI/3jtEADgX7pIfc9zvwa8PA74Is5oMCjPvA4fzc/LFU5bWkhYLhoa9
tUhD55EXom5aeuLpMp0GUkiAwDm835CFydngjUTQMFQiYAV1X/lBIJTjKkwNxRrDu7RQVriPQp1Q
RvDRYtxGjZNAL8aOS9V7Lf/KsoWHJEe5NHHZEaI1fArUOmbxQYXo/VZX5B9BN0/JyTaOeMU8XyUQ
2D81jSrLyI8HunN14kkKNVedF0tjftC+81MiKLvOsYihUOx4LbHaAWNhFFmokEAw/YAsf8esPgec
0eoX13aHv9wWM0Ur8Rb6gKKgCkS4SGWiZZcAut81xth2HYbw6JpGX4u0EeieuACf2CHqazHzH2LR
lRHp1VdukLaZ4mwkVxc9TZpHjV+T3jTRxGpU96t7tmuEdPgvMA3fwo/Q0HylJL/LPjR4RE/fUzSt
N4YGVRiKmwjSAEPSMxrbBH+bIYHCy0nBL5yrRVSmQii+cIPsj7m+NjKJ6CJUHE2zg8UdGYW4il9o
obml+Yd0oBVdiJDhNnBuJlk03VsK5NB6jzMPSnsjd8LarT60KeMyQGx7O+3QFjlf0sJn97rNs2FR
wHuTdw5G4TgAa7xSaPvYbd0j/v9YY7DYzY/ssFQUwEBjyA5pOcXH0Vl7sdS9h+8OT11Gn5trnG03
0rS0Z0tnEFa1n6QyHzzwfAx1PV+/JX7jkmQGqnPYs29QS+unspJggt5WgfttvUDaivowFNzFAB2d
ObPTKLeiP1JpbRRR1qejmGq7NISGO9uhXJelAVGfbb5nkA86KWczCN+Vyi8RDY7HjG3aV9RSjRLt
4I5497VVfsDHtD6gWu8NUO9QkW+0NamEdQKpuDZLbqt/UrijYM2IlSw3UnR9UkRmzstm/heT2/pX
gJqOyfw4SB5q1PUgrr5GV9CXcYciwsvx1TgAPoq1/pRZU1MLUvdCTJr2rtWOrzudGhkqVEQnQJ57
hEcSSvjxazzDzXHSGjgKglyNUI1K9mWuQwI1RkRQE1+qfWWtA8kcqODY6dt+CjJzLHHzw7Icl0pq
bWnWEUTQEYpGjZR1TYvPnhmXFlanuIvhXxB/LH+p2w4pWlj9aFc3Y+xtnY2O5EMay1RmFxoCEBOx
fQa1f9/90VFmIgBpDvxFEmynZGV09N9H6rYo7gz9fwR2y9mpwTvZOGaxii+ol+X098pAALJvx7ul
ZMk9nzka/5QrQb5jsn0UiqHD6kCX87zYCB8fTnjeO03MGTgLOOakBny6TuygIqHuHeiDin/r6Oco
/7zm3UxDQR3hHX9F8S6/9BVXa2B3UL5VhTHwQSP0i5NKNQ253ByD72yTXQ0QI50O4yomnDN/XTGP
fP+1GGazKlKXzvUdC3G726vq2grXpltCWOEFBk7bQTHps6bnC1piLM4VQtutNK0zoT+fWB8q1CEd
G1gjZXgpKvbtO5DyuHY38jHL8Xyog4Qj1V8fp8ciZkq8zh3wq7u8pn+RHAr+a8eRFxlH5X4x+hTY
Ec026RioxuHiHZx9LJwhNPUWTU1/Kf/HEjA5u9LuBpV9teOGWUAcpux1z80HiRAphbA4ozzJYX1t
WVFWVNqMFGcHFgJZ1W2sfcIcximE3IWfXQVl17U3zy2rk/XdYO0qQXbfmJLHjY9tbu7m0Ra7MhWh
SIBWgKhgISwntxIzmpmc6wJByLmtDzxA/HJyr6qgXGoB5lkSPTRQTq1MCE54TZb1LDQVrbkeNAJL
ut7uczedZnNQDP51AX5ruHHq/bkF/bEvViAh25sr+0l0b+b5CAQAK/SWPDgWSqADhOIYHccdCsXQ
7PHIFLcUPMV/2YcB6PVbq0EUsi7JFgdFv5Bww0DepEkznP4A7XnObPUudyj+v11eNkAHM3LE2GIo
CpUfm9v9rWJnOQBjd3Wr+HhDp6bQ9BujnDOlr1Ch0UMMgCv4LqLOcspucOwsNyYzvwpiLyglH5VH
vbT6xse62Mu3cIXtuopIvijf6i4p4PZCmaauCENtffHscaMKQeWJuqTzRIaM0ZSmGD9tPBCab5kw
H+Y6T+e62hHpm9tcRaMVMZlXHj/qaYp4OgSVdt3e2T5n+LDsQE64oHWhzsTpW5F2kPSxh9MwPFS3
oW8Rf+9xn/HbSybPN6aRxowXxc4KN1lxKsppCTiHDdvAiYaGFRe/J4YYsnXWv/zT83dgGDjsxnfE
Q17bjuTbRc+UwQUU12S15MiEncNdqF8obw7L3Ezu8DfVfmx0rFghOv0YteNj6jkVN0i6q1pVnQQc
lorhT7pHHOEBL7BRX2tMeiReW64xpXucle5cS93NfKgY/evmKgC7tqqL4zuqH84xqHkazv0g9M5p
PA/6l7V7QcGD91RAlEU/aDOvjrIwyFEpQWNd23gLzljEQ3WSKigmqk6wyPFDDddjWDLKyCY1Zci7
hsM+wqTO++oIGyzl/OhXsELPkKYNoiDHZOGszy4rFPKEqqpAezA73hUHlE8XRVii2EB996C5A+LJ
3Okti1EigSaTCCEZdknG34mK3Ibqc0d1ovrMHGdy8u31U40ub690flH7YBZzIZFr1EBzqoxhkiGs
WI0+oOHhMTJjbQucBdwIYexLTRPL+5DhUe3AnyEXpKFJJ5Lmu4Rj0YSAwU+UppXGLuz2FynLOO6P
50+YQgVyegU8FirKv4CDd7GkcdiBLNgWrD4wr0PvZ97V4h9vKXKI4Yi0B0hbl4jrqMqVxt2e61t+
pKSh1lP24kgBZqkOe+F2iHuCL8n78vuqe/3yle/7d7WHYXCOfy8Pe37Bc23BC5cd9r8uKAuepWYR
5uW4XrAJvZkkA5do5svyQrC0PxuVYg5PI8NJ/OclHaoT7w0FQUro8z5k24yFAiWhEB6uLWkdZeM/
KLwpwC2sqaiS0zYP/5l8l0ra0I7lna4pJPGZ4mey7aPU6mQ9G09rWUNLv+2lsiHK/T6A7qpIUU9Y
3GOI1hdZcBmdQzT7LYSSZv4x2E3eUrC651kachKLkbh81mIJHvhBhWcI3epRSzT5MyXRysAPCUvy
+DJ4jiXxz0t+OEJQDZbUHaxmwpVIErn/T3AaBhpIptiDoHp/fiSWVl/cpjlYN8kI4MP8P+7h/KIC
VcRS409eqnF2BeleaepRwhDeUTxDaiFhsB/GLMqBMOJWgwgAbP9WxQurEe9a1ghMMWigZzbX5FGO
LhucOIJZJnbpmcY6OutKwPjdYc6aXSjyohV6qMFY3/yHBFZBaXMg/DLOEe1YF2oh3AyyY6Hr43bP
RcqNuoh9QNG8OpfLSDmiy20NbkZe158WNwaW9Xm58eZ1itLSFvj+fizC87K5l+oHDu5fvLM+x1vk
auop5PmxO9DLMXuCKpPwuNrmqirT7xH102ZIU1iarUQ9khFaJ5NhJQAWnZg5v6vgt/WNdzzLdzXz
hgngfm0hLT2Muk+2amF2J+Khh9muYycZIGbDOeVTs6BnMfcQeYYtaUsbdQgdq9l7+X8/UHQWkimA
U4NyGDfCnow8CYSQThjNrAMQ8kgFb5uruGj/QyLbFLFuG0HMUtulDeikHt1MId+5I6UKXGycuO5T
xsHrBym5MZmvzT81u5gkly+CEJ3/vt+gPdTbtMt90n3q2q2G1LR7XGvq4fnb6Q15LgnUJFY2Bck2
SkIkGhtHxw/ko6D+3Hm55VllLi5w5L8VSrgvRcN/I5wF5f2beQpiCIgYlrx6t3cX7EF7ApKhrLx1
2yTKFGIhIlSb/ta5YoGQRwmhBpHCz2Z7uQGiLFBLsM+Fywx3+eRk9V/BB2kWsGt8itvNtuqrbMte
3TxI10QoqKkVnWREQOazJKukIO9aPsUXi6kN1iddWr2t605obBQM5lYOQ2egQbvuZZY2tcI2IlNP
qRV1JNdg8zZa0nLfo2IUarQowq0exz9rPyDautG3mC9cLIu7uCJCovlrCbqUPd+qKp9bBNI7IwuK
R391/2ULe7Jvej8cye890rQWlB+OewxjUeKhxAW57e/OtJ50d4bxyRdPJEDD1k26EwnmGD27+yVc
BfaW9CPBhEg1kkyP7T/QE0Ya3sxOv5GhxEatpOOj2RXJJKMpX4n9hX49mqlJhELKTmvq81Il0dWv
EGzcfprFCJ6mza5t8x1+xshTnu9X2/KcWQjSXKoMySL/p5Zyohb4T8NcoNZVkjjE5Ra6iW2HCvZM
ykvIjnXlCk2bTG0hZyk5QxA3/rl28PPgnYn6oo0hVpnzU6iXSkVEH4P4/7frGEXXKOK/CzzCNg3G
E5weKPU6wQ81QBSLvjDRoLisb/mKtSqtPV8W0k4SdT/we2+NWzJrjsZ0JH/c1M6mWGW/Xak1JzXT
lEWZ4FAZ4RU7f9Orhj6X5JtUwkKj5pXIvw2lmL2nvz/M1Ikx1C4symY2nbXYvl4G1J+ZW3whjYN1
ur60dVybHob01zm3zmxnAYhf+ljB1EDC3NjRnB6IxP20VBGQrB8gGHNwA0QewRUylFhn4NE6XzMH
iOaxrSaV77WwQ39VjW99rPz6Ow0y6nnu1qsMivYEJNdsQSj0OdAXA9gCV+6vlyGGXFHREKBFtTCD
xTZ5iIecEfAgg/sfVyX/ANuxPiApOVv+BIIRbmp1keBFvn4hb/FKgmnZmwlT/i2dWu8tHL8Yn71a
YTBsNG/dDZya+1M3SQ4tlX3sC+Xs3OyT8nPxXy6j4fb0RtLRXikOoNsWwL5D02R5an7gPnSrvyes
4fyyvvXcbNke82D0bjhuboKxcwF0KLoJdVjyXXPZtZ6+Yg2BsBupcbaUw0+EmIeZPTaPITsnPASy
v08pQA+KNlaXeZArgo8luqgeFnSIAkNjwfEfxkd2XEfzYCIOEHnmE02RpFWU9RTkkhh5WU7Z2Gub
Y4pd/9yxp/3EDBjjuziVAiMrmDeC7WQpNUYCbE1UDbXl3GfdpmQyj3yuu0SpuCwsFXHcHI/L+qjv
IughfT9MwDjlP2RV73ROhoE5hgBhwZ+voQ/dK2IqFKkpMUg0irL/AR5D3MtdkvwZ9Yw57cgSHzg2
LicG7hm9jLp8PNX8r9hkgNnTP1nEad4zVCIZnanTnMxX3uZCbkBuE2zCg7xRLTOxJq4lHLenxsZg
3IAmwrp8KzeSlg1HXEl9YH7oPxLN8/IwniKDo0iv77Hh+U5TFrLY16hAtWLOnihiCxRWtM1JmxYL
mQCvnh2g5hEsYO1HGjf182uNMhHC/b283Tx9wBf5AhIA3cD5jc1nBCTqHLrFWoqxJm9Hd3mknDU0
IJRgBJHsgHYKJek0rY/AP5vSL8ucKamQrgDNE15m8+8+rpNQi2DU/drlxl/FiKjshR0gE/LTysck
cVgtqiL826NoeAsr/ijh5TAg/5l9n6y6ghQ0qItIR0f4EObbXh/BnGF6IWcQLj4BZn17yP8xwy/j
XeFLvOm8dy2NofTIy+9Y3iM8Nuiac+vFx5inRI49uMTZLUy6PKIgfNOkPZDu0fP2F05TmKPMsSUe
CQooCbVXbl2nycqrC7REF8JDlq0f398dIJaTVZfROSsSSepo6d7132K6+r+j8eb6d8EVfN2MMsM2
YYP7r5qe5W0QBX+E3rane+r80NvNHq+A6tLxgYTVKgTYGW1Zq+d4Fx0sHJF1Aw+Co2O3VTyqvPQB
hxRlM4AMH0Xd8u+A1rWaapiWeARYXUmbqlKH2amkRteBOBRO8fGva3I87orFuuC0Yu35nOL5fRUv
MGe66nGPK2+DO6OOS9w3yXwVkk4V9hXxfjIpBQh54cseRlHXpBEUZW6ERFUBEXcG9xn4MibhP5FF
5j/nxS5XEUHsZhUrqPUpcDG+VADRmiYysZMX8e3283GbGs034nr99Qzr+QsVFDYo2FbaaZHQQ7FP
naA9l6ZO7Pz7s5u2+DfvFWBD9g3TERivOhzIbm9iG1hJxKkhbdnIeh9fYzc8cpW97zzo+oertJcr
EkbUSXaY6LXhFaJ11McaCuK1DjNssmSxKCDJdIYOFAUMPJ1cddiK0sucNXcITBCleIhvVJc1QKTX
ytUL+lT8vSWkCEWZBkdv6LL2zWki6GQUxyZ6X5OswPZjwv5eiirEIe+kphfh3+FnTJLTmfm/mowu
yNucOlu+o6qnB5CXGrQEWd/n90Wz0FlPeSgrcVEn6BYh3/IQ7JdFb+B4+kfimsvO96DEbWD0TFnC
ab070l576c/Ocn8R/0ilWr33EHg6jOyoLsLMLne5X4PFFqeps6FoseZI+X3IIlNT/xF1mVhfPlQH
55A++GJikhHFI++Aj84q6XrLzbauWonoC+ppUQUDO1gtzjWUT7gxfdUWvPI4yq+EWVncj7qd1nCM
9LyB16vQ6r2z1GrOAeTg3b75g+33oBQSrQYRBspMhvmisEemhsScd2lzVls3LP/Ndk326tNt5F8q
qIVWqDU7rGo4Y+FCtcdIeib5Xie1bKpE/2f31PocVt3av1FhPJnUyJCgVqMnjuC9dPDk7rKhjb5W
61wC6hAioEBZ0ETYz9TUSXTNkU1IqPrvBrkxDSk/Xp60WtHe8NiN9osdwjEwTdMZmkzRO1Qit2DR
dK4VUOvOGzEedfSuE+YEj9AywXZo8QQ+LKakzqxCcI8ejZ0rkvmByks8df5ohe7khOMGaXP4QAle
TZGXRTCCcU9WpFYZUfnDG9x5uiMZ/u8xvPU0i1rUzw+RGOmd5VP2xEOJDxNQBBMYfAA+fdrbyV6J
S+TMw4fiBZjjm6uERyQzPNunTDp/2X4Y4QnZK9lR37we1KUo9HZLwFT/yEGuRrYxWoVDF1gk+zLu
krvBN1s1DLt2SaNBMNbjaBnwBHtAgmJdY4YVnqB7OU6yNIbI1aWmlff/7JXw65245hlQlRwOeP+K
QQFlsFA7WWRYiWtddaX9D59fhEHHTNRYqcdl8/pZ/kEEHyTnmt+RYWBkqgvcdTbZA9JQuBvoJd/e
zmzCa56g4Uylbr4ovJWwGW9YW6JsGZiYzaCFouaX64uLHpdd57kzqgnAhCmeU03HhKfFW8OSkpBN
wDL7CpoPsn0//VHRf/L42kZdTAIDaLP6wrWtb2chWyJgwUNW742PrkyfkN7PnHzTBqzzjFDIpoRk
sP49OgWZrCvmHZQCWvkVSceU/ifO/kgLNfSi/oRjV6Ot541QnL9tSi7s/6t6KCaOu75/twts3W2q
O/TD6N/NAZwIcY/6VYCx3xvF63w3qHkCW9Qkrky/VQUgYrzWh9bKDRKFDVrY9LD6qrnQlJQheTKY
i2Gb/sDWu6VJoR+2X1aF9irB1JUZTW6SRfHVtUDfhyv5SxXW01re5dS+gB//rdAV/w+ahEjQLvrm
L/mfz+mmT80qKw6SGbjMx+d1DOS+1JoYCAot8iNiwYiH7xS7rpjDCi+sWf2UPZvKtim8IibP8Wu7
AhFilYvmjUc6cNiVGiTB3ZaP5dS7psTisn8peRoYkpsi3PnI5tOUB/0Wa55xxvZL/DaE8stYu/Gq
+cllmpUjzKlLAnggcwOLB349RsogM/BvFezBMbKpsttSvUILa0xEUZaB4E5B+7lUV47tBVtYklYx
1xRsMlu7E6KZ9UwcqUBUhhLToLu3jJXewTrmVx+klTBYAlTJvPma5FZJ0nFj39neI4cA1pbyDfsA
JTYR1dxnyzbtYFGbX/1y6Yx/amRfYIVlyq7H1rNcLaZ1ePH6rJ64De41Y48mKQGAnekGPbLxdzwc
mpgxssG3tQyaWqTiFVtf8P0dPhqcCa5QU0T+CIAsB7O2MJ94dtBaQGS/FwZe5SOjueKFtBq9gd2h
5wpo8EZsaSBnuO6nt9IN6CJoBq0Si27TSjQIG6Wq4Aa2OYHTdmdt/PJiBtujIysRURbid443bn0Q
O/1/LodbaxHSS79oLuwuap53GX3w38UdEEpmzsySJmYDhT/JIE698jjqoIfgsG6dZwhVNkjNK3oP
EeeF80yyEf2XKbZWWgRg+uJFRLY47/+cQYnGhOPsk18Q5g1ZuGrkB+Y/oInGTN1sYQa6rZI1jhK5
+j2rneECIEuBcG5aMSiONBFy7zVi02zPquXAnSMqNjcpZHKuOBe5apBO8Hf1h51MvToHgJeZji3R
u574NEVBVTmrCtkA3/YjIQr+7xPR5wh0Nm8OARLEaTBDYAHjW7xCUJi7SGx/ZPU7hZ7Gyqs/AYDK
QvzXHybhNE/9LrvJM/vDQCsQkK1f3qb4YnJD0NdwFvAAz9RErIxma+YJujFXeXgFPZ7OJYRK3N8E
YV20ZzRLisFKPW+k/w6ekEnqaY+0ZhvgHEWgXMDVMryLVlEw4rgVId64o8PLnn/uWQi2P/fmbewJ
x10GzWZwTJMgVEwuRcyAnIRfoSb8KUPydPsBrTNtr9nl9SpXsDAW6aZQorKEmretH5EWHuLa2AAa
ykUEGc12kQiPxGdh392AYE4oZtS0h7PBRcrPFQtCpNgVgiMMtC8F2KUlwBjmZBR35ALMCOcYL4jH
hS9O2QyjQ8Nu9/Yq0u+6PkSp7tlV1SfWp67GfTx1r019IX0ejYosH1H9X0PgRyShynoOt7cygFzu
1r7XfDjsXj2CBvDRPISXl/4eN/4wscCsrkzbNA3sLicbJgbCYJHOTrguG3nAkGck+NLmSKUfJ+ha
7625tahvPtC0RyS3fczPJ4SlFijMK+tb4B4Mm6+SvTk6Ph4EXaC0hd+rYnZa8VAf4mtKbAbPmb6d
AfJ0Jps527DV1+vi7fwhNuSwyiOcwcIaNJ9E/JQ4pnuJ1ltW4ZW+NFQOEHojT7QRPvvrKcIKmmUz
YxEdKzO/06XD7r+vzWVTteq1Vx/1h/j50d8MC70PkejFFOim4DOKq1prMuSolLguE9jNRuWq1hfv
yvAq+eCNcdmLukNKMO8ItAilD/HuLxNvj5Edrvp9Z9yFbXxOCu3aWXXussb+x9HO+7Vt12/vbDim
Yn5VgU+dveSYekHwZD+WqPf+xw4HpAJlSL7AXim3EOvx8cggviDCzHYNBOFDsaVu5U10fS9hCZf4
GV588OXs32mNt3Z7yeBVVzztmf+R/KfhqD7spcuFZBuzitZLvilPIcqbKMo4ivAmj8z4SF1rTFN1
PVf7GMqUF6gFlDNpE2r+2RXzaOg3jbdGrcWGSPnmStT3D2hCBXCrYVBokdC4/PlwZm67RcBvGT9c
hoFVxK2r9KGBsytC4v2xuFpa/5IWeNTF2DtVeGg34gGBmLQCyfakUY7ftwT7RAaMJ0r66xTknJZq
Db8JfWAnO6MdBcWYaGOnyfzrE/i+CS30FXb9UV0fzVIHgyEIeatS8WIhh0kvN3+0rmOGPGlJe5VR
Fvt/5CQ04YBpZTyZd4v1dsDYcXJh5hEi79aGT+ebPEsM9XOs6gikchn2jlOXAxF8x0K0cKiGu1io
aI5z76cIBMdkDZioTnkq+oaAoh6fyApFXGg0snjyu2esrEzl6VGCfqtixdQUGjnPoKv8ge4J5WY0
2OxsuPAgKelvUGqSJfpLppqFhsMaEoEgcTknBeA3HEsOTXjO09RzppgefYUt0cwKcUsLilhpojc1
WtjkIyQ+l1o4l2J76jJeTFvg98ekKJBILyJVUr4NbpNNuKGHKzsryFwZ93a+TTiA5x4nraqSuHr9
mXLOQUsfXnuJTcrEf8EXqLgHC16rqEg8PeL92fC//4k7YVcjWpPVtzkV3HobRpasHe/rUNyPNXA8
WR/thxajZrZCNTDXoX9p6iAbyvLoj+xuem8X50cmaVDCgFSALVr3FD70va109+Y/fUWB9+qRVJ3y
DU7cUMU99Zy/wyEz+Q30fwqhRCgtGKHcMpEQWBhhMMJJpKypN8Ia1qmCmUQSjLGyV2cnfGuykDYT
jifGddftWSz/LtAuBXARVU/gqMbJ8JnLJ6dd4J9kilxCLXrwUPDhH1iDv8wF7hM1t0ZvAKsdRU78
fkOAojXa3lSvSYTlbFqwgZSnqZjxMemqhhtxyjABqrY/uxoLK6nwQSWRJCp8Ep+Yb3Bb6mTKMxPW
W14HlW1z78axg0eGZcidKIaAwi3a6IGTX49+ZRByx8qNP1R/SKhY017DWLc+86mJ/EbJsHRqJnqJ
Pph9x9Y4Ssb4holiXMRzxG1Uy9ZImXpSA8NapFh6FYuP/yCqSFIcBgONqXlgjzG3Zpf0DRCj96+x
ZXwpOxECmYIGRGmJDo7c2rCEuXz5TA7uUMJtW7B93D6PgXfhBVtmzMEBIycOuKIcQCQ4mo7/gPpT
EEGN8TE/B6zIkIOk+faYlyjKZTs064MlRBm4Rpq7lhWJDgCqJcKnhcS1Se+vvlAzrUHBSjG9D8lN
WPFC18iEKlAA85OT1ZcxPHUKIFtWL5DUprugbFP8P+eE7ZW2EnQwKhnrc21MgrKS2VlESbkp8SFl
wdOotG/9biVB/qQk2YJ+UwYbvrrFl6LGcwQZw9qo/8c7j2kvEY1uqorJAyCo4g82Mi9uIXy/OVOH
fTOw9xGPUsawqHSAS5FOrSN+XatTfe7xWLbzbOavBVS9Tc+eyRY7zFsUaWkrlSPa/yvlNe0i2yMJ
7idO8DEzCtx9MGF4/riYitlq6bUL6Kh6cFtQotFCS7zeFXi/QpKtoS/mX3klrj5NAzZLq9f44UHF
uomlj6OdtWkDitcIbtUcocALwhY3uqxtvepH3hh5/Zwj9GK2BehHFr6VP4g07L9CdYO5lK3NqC7t
G8yK0k+gDMm4lRZm9eKsNiK5yI2OQTXcgDs8Wx1TXgORPyHKCRiAz4PYA0fYuGx7NQxzhIJlGbsf
4kgCL2caxpmFqNPGc8tWeeAKDjObMB+6ZM0ErT4J0vEfnd01ERZdrUFBdTccEIqIH/cN8BPuLrK6
A/OImxpBfM/D8tlluuz3ZsBt9aV9EPJf5skoypdL2R4pxryjnJfNGnjfYQWyqhVgw+NHkkQf5vSe
R5goZ45S8jrE48vn/1TbcIeJlZzk8FgqhTPP8LW7kksNsnmDOS+WjspCCUSPVFVsx2flTvr9VjkL
6C+IPUA5eqpvhu+A6xBZzFWxgpS2HokaMml9tBkIWMNQvCBKf+eqDhtJWU0ww6KR23bejNwp3AWu
4/TsLpShlF30AWmA81n+ApFtQ78FTFphr9o9mXRTtKczs9WQGHQF8HB0ouDIWO8kYNlrq+VTpZBJ
cNuKO4Y64Zqn37gC5zTaa682aXKXrNxqVBHhzZWa85IhqYB3Gcr8wYAymdKEAaF4RlE6igx4LBzp
3s5gBMEtSSyMXND2m8Om5ty5Stlgi8JHUr+JO1crGDLcz+EY+tRVACJaocMPJY2/vMABqnym+Slb
CCTvkL5FX0Dsbet9WQYSQ00e6sxOVApy2m8vacDDoo0WIWz/UwBz66i7EwD5MNDq2JKHPVLrjdQp
On56CtyD2LfV/TeAJ8t5uxcRCQB3ED4YwryncE1PdVRqPPirZb+BnDtdBfy1itl/SMrNcW35KACI
QAXqHOZFmEq9QV1uCF8EEVVJiC1HYTNA2Mt/5xB0HD+kJc6vZ3rYlbxKGiV3Cmv8mSeyw1ME98vy
mW6m1jRRIXAYmAJupU744iKTrIOf2DYOWI7M6Z0qOlyQX3bmERXPJ7eb+/ZObKSjvsRcbIPassnO
EtR7uU3Y2sFW31sfzz/hEvGapcDrHWnPJdY1i7Uak637GZ/QHMg09TY4L/kqhJUPqYBEqE4COZWt
uHqRhgCCKdYyyuopFoWe4ezjZQbS94hWR7dlvSbnK+A5bKkqJB1pf+ziWWBp/+I5NW5Ee9Huf20n
XTv6bUCpIUNcOydAIY9WGQix08ieNL5DfTrFw17tApnwP3tvLHDCzsz9Dzam4TyOxV8/zJhy7oUj
Z7Kk1gyvJVY64EWVgVaripNYVoZr/+wblUq5khZ7FuJ6vT9Fl3Kn04v2F5rQYApRMU9Fz3egfcX5
Ug7g5YSTKK7AiD5nIOGtXiK6+vv2sAWudL5cZqYSJJlYjF23JXi2WXSZNJ9DKpzCIb2egx+EtYfZ
ihWGyq7T4KDYCgf3CUccBKiJRlhqQ60U7LSbuN+jsqJBPSSsdmQ1l5Ks0NaRz5fwx8Kuo0ejgxut
os6cwZUnPqxmPWK3toGzDPYy7a40miHY/HsJu1s31uc+cvIKTbZ3jejBImaHb+v4K0GRf7NGFuRC
QXmy67mjiEXo2qct78d8MSnEF7DtQ0Bj2JBrWL6F4GrP+YAKfSM6ly1cC0teZR4Gr2yhf3sCq1sf
9VCzwYMsy5qfxR2stFl4V7kJi30k9JTH1MzB8gW+3G91LwHEnhH7aGU/e6sNH2JXMzEhMKbqQKtR
tEGzL5RDDzQpwQi9DXMfDwpx2V4XktCYmqMDMROnAjQzkXVER2LTHi6BU9ozLxX+C78BOW0AVeUD
/jR+rniGODzQrN2zRMItMCjdi0nGwk3TYKcZNKUv5+joHViBlUJaAgX9JqQhh9zSbkw1kx/Wlq8c
SWsXRZSKGYueB0d409E3kdqyh+oGyMz1qGcrwxFvo56MJ6ZT0kESsh1FaUpEZ8BIQC5MyFCsbG6o
zNSdK1P63oPLOg1RopD1mX/PNpyNFI36vhzrNZOpNtYIfYc26azM1zmFrT90AQ0+AY2BbHTaMzxK
SqGZ2nRV7RPUBLp2SnR7Y5EedRzRD/WymQMZ+st9nJZYSM6NLaIgzz9t5h49QMV5AOgkWOisoDH8
E5R8yPOyvX9c+B++yQjiJqni4cPkfpkcmJepNPEy/dtCqFeN46VzyHA3UMBDUMwLTgLbDwUFk/nF
O67HhZFshdpMbsvr7JaMiGeqaXnxBngKdwrG1zFrGV9ioDvpimgbqKQkSx8oT94LoLLSr9I/I2CJ
KjoTPGUYSznjDBoauLsnmQpFnWovNvQ5Y2stcMWVzhp3bnIuulCI/9qXQaju6a00PZCre0HYlhKX
3jcfZGPaK7KopnHleBr96adrg9RZWd36fMTvHh7+RoaSG6lcO1GB9/X1P41Ue3MM6FXnp7Jas/HG
/fRmE0KsRZ+ONhmoCuiNTLxT1iKrcBx2w8Ptsw43FDtpvNbn8u3pquKnO485cxC/5kIkDH+y5HZO
ly4vAIdytnxblqgeawelmyvVUjta1D0z9GwunFtZVRKDFF57doH8uLAkp2FW4UgF6NLiFDl5U/wC
hs4PtT2e09j0/J7Nrgs6L66KivcGCGlxqxwIRgUbYUHuoFYN0fsKUoTaXw8CLE60btIUUsgmaika
cr03J8mOR+8jZwx08fpJr2qpXQyxp29gUfY/p9n9UwXdrrGUIbocs2IoJ0vVwdKDb0DB9CzeSoyX
CJlfeYSrGFV1rI5ncMJQ4aXshdWUVmKTbMoNANPVKwTtam7tPmOlvH7AghMyvmsPXAm2vWkKIZFg
WXb7uBD09Tq1rw1duw0gJJ2jev4h9g/hwWjXe1uC8aSEvx2ViMhD2un6l8ZLS9vFFwefaH3R5P5I
BGz26p4eJd3OBy8QHz6zfM21n46dpnhqPpN4dSld6nUB8J4pOeDzg2SeiG918aXn8GVgj62s6U5b
S9LexnOfcVkwx2WDNswbS8vxztWfqXA6SjOsg8U4Y4OUmfsqP2eze98w68BfI9JdjaF74Nqizxc5
LQ6x52HxLHmGNgih+31pWofZTjx4FeRx9R6be71Ib60eDqeVP/DSFY5maQh3z820MMbeuLQyhVBr
b6oynnTA233Jhf5YaeHizNhmjvQgC188ey52VFHIl0TzhPcT0rplFljYX5629PHDhrONHFkKb9Pb
Wl6WCPnNeVIFlYj7XucDBlXr3hCyD4w30j6GI3csE2JimgFyrHp5q7GV9gPcHYHy+kwD7N+ia53/
bng9N5L85MWN5pJ+bxoXycbdrBPDQHFGsgTFCZK8VJwNNkyFLuYu1VO9RfZ/eJ3F7OdB5Scft+ON
LHuWqwUIcDH+RrUo2smtXY7BDilZn//XiO5YLvjs3VFdX6W7SYmEaAm2LW5sCWT3SJ8ZldktO0Dz
3Wvz2aNRSA5nXlzLZLKAVqceDRbKUIO5xccwPLPcFLoQZq9CF4RN8X8nV6WqduJ9NQt22nac9ppx
fBl6NnZxVlGCswuMfmYaUYSEKVaai0cHhtjyU2RbER84YVJwb7NreZ4T3XQJaP+m0Z+O3FYasCyw
+K8q+4m5j8A0SLuT7XzW+GNZszBwodjLN6BeL30dnNp4RVIhw1/ur7IQjva6NNYe1XKxlOvm5NTE
yO11ltE46/wCgTy/JYyy7Uc4Ba2P4/7wDhAYNOGuzqFcCsiPm/qI1J3EpUdc12++Hse6GmWCGyJY
T/y/jr9eoOLSYg7yeFB9sY771B8YgerMLeuTnd3mpzR3SeBrhkrSh9SlyLFMZpgpHBKXRadBwNBl
NR2g1ia5cChq/hqG0/aKcz/ACEfAfvxpYxzZmUxZful/rtVa3hYF0f2DByBuV2iknvoJVwQdEdDW
tCUarD5jqm3bKXylFJ3O9Bjv9mCBRFckXEjcoAP6vGQqgbikQ4+9pDZOp4JtGhXXStjOWtkY1qL6
I0BJk2pgG2CbGPEoEfnQMLLKbnXgsQNolJzfKu1CJ6yEOvBW/7k80WWW6sOnmkruoi+NKrzl0ZqP
ETdu06ETXRwLq/csYKEeF2vdTz8eyqiZ2jrtoQXIcjqbTLBLkWryxsRgiLDVSgHAwsvRosf5JDNm
uMZ9eQLuRmy7izDbRS/DaT7/pfCtl1wmfNeRss2gW0T7XPzDA9eGk6vpHBUa6XJ5lQSfkQn/a0rc
PbMBorWLoXQgYdnGvzinOb2A2CpHotYrRw1zSdpLTwR7UciZtJNzpO0rFkt8idFdxGQEsMMr1FAd
S2ZolHdHVvalcKz6my9uYooVlJxiPSNxldWkww26PhP/MDoi5bJxAYMH/0J/8+rK6HtZoeBDFexb
/YaTrZJmh6IsLmrCq1TEtyc5802g3VnsKXNqQaL5n+8AUiXuUi9w4URElCuKvIu+roefx7SCM7Gh
IyrJ4jyiB1/mSohKFaC0oovpsaMYzSe06XH0Ke/vr3IIyxbOv2TXkujprj5zSVS0j0y8JKrSDuiz
dQSmIk+dj8fw6g/dhVjV2C+e+/TeG6g7iMe0am5jayOf//LuoBEkwdYt2fzB5yJ88km1odEY4uUq
Cdu93EsoVEL8R0WftjmdxjFxkkyltzbRTHar/Al2tCyIAX/ZYIcAkeLguI3VDRVkxWxANNPwgW6l
eagIjcdc4VViFGSlJS7GLDEA4jzQGczfQwVO8pWvCtZ0RwPBP7KvYzy3NyIGuAuVI7xS9BW6xbLP
0JZ7Yq2/tudbLKUGiqNEdGAi7Q1HzkSZDP5nDxInEelXqTBrbH+nvnWRkjcabMImRl47IiAv1yAn
dKli/v/ttlhi037OUE2C24sz/EMCg7m6FxLJEMZCBupzWPxV4tSV7MP0zGI5/Z9PRabh7FWGwxyx
UpDJs9N1QEiDGR7Cjq1ulQ4QkETkSvlanAwU0QZEbNzvmQxsDtNfvH8NtP28K7nwXB4quWFyVOSF
2kIGYvJXGpsbiqbPX6CdDzm8Rt3oBrxSmlx4c+VD8cOVL6QasDfBfA9yGY2mN+lSCE1Q0wMT139j
mVyVSa2o0OEqir5Rd9TV5QDvBY54OJc7RTh9e8kZlQGASdeiFWeHxo3pxDs/9UauRohLDo4QOsF6
rHXj7HVJDAiibBG5Ef9cr4T+9Q1hr7WhcGiu0kneNMAnEsyrNxRf0ujcuO7tKgsjk8WUHXdgPavO
DA/z4/zYzRXIwI4JQgLYjoz0TbG4SEmhpR/mKtuJSd6CCn0mejczyzylxmiB2MZMQuTCWXZuU4qh
EB7VrX8zAAiW32HXbIAKysogQpa4PpSpQKODkxWHGYe7bxquH/LzyOUE8vtljZJhVpNTg3kXGYth
Ef6Jf6HPt1J5AR8/S08GUwGnNfCQ8YbPGFYAdsjZ9zgS3q0khs4m5lkqEBIQnRiM/kyr+wlIO4Pm
vzCT1r2qzCoPhQqMwKJSQ5Fh2X0zmm2FSGlPwugKiT4+K8wq3Y+oN9C3lcY8k8LbR1WCUg5z4yLU
szlltiw8brLiEevx1wv/VnRd1pxNPy1WAGYTX8/MF5WLHCcjqNee7Bi62XV0geUcpvUEFkYoUWL9
B9Y7oYlpmZGK6Ht9sZkOVpYzTzLUHWvbHt6ITbpZ5ZEySi6eVSN+5OcHRPYVonJa9eRzX0XxdeaJ
JjVkOOvDKdZXQ+I0GLeInWlkHgZc2vx+m4QAz6MXOwD89TTnJYvNW/i2molM1CiVlVCM4sx/YPk3
VaAXFsUBMSJcVdZx27HIOZdxxJkniF90qvVY+vb2DBRhOg3KPba6dfx1+eS5Srnza+sAs2BHT6PM
gveF9fppUmzkeF/lIs/MTtTw9VpgPw/aJoBGGEaAfWEexHATPN4326pb2aEBQvsiKlZ9zDSAxBzF
6nTuoBpeTXnVFpZ3xQZMWeIjouX9njszkQ1wNbwF2gpiojGDFzY+dK50h6U7Km20Vna3gjs16d+n
aW7Ro8PBAvZRWPMEqWwXJtH9JRPV7heAluMzqJu4jz8U81zN+YOaX7oXuVP6vwOOhlt2cSe58i9r
d3OHgJm/gFBVZzNd5UDeviMWdDy0olg/RTxL1GW37c8jsDAAWQa95MVGXEgwtYWb9aVUXEv7wTR/
20qimCNt5kLegiUTSBwraHGpPPWXvWlhhlnGnPD+i87Jv9CcLEVcfXW0O0dx0edC07l9Ag2OpgAS
pxkfmKcUdIpoYY+xMeGlKGlK87NCPj9LYUHirjvsATWGyNiRhAHyBvSvGshV4Xu3blO77Bo+9dtX
G1Y9Kiokl55aWnl65fqTIl7WoP7vvf+7FlCLgR26R1sFoJhZC55yCL7TAFAwNzO9QW60RoiobDtW
3OflO1wRu+0br+kgcarxylR+QepEaBG9fn9ijaefrIIIDFn6q0PZKWeSxXgAEzlIbeEhLZJfEmaq
EJnIQyO/UKhhucIi0d4j4bG3729r0r46dTUnjrHwIYpc3vPY2L9QK4dmIQpDw5AjpArg69EkFoNs
1nNeltYHX6vI01GFHHFVQzV+Oh/zovu0qpQKHPZ/MVTxhH4deJrzAb1/qR5XmY1oHa57u0G+Nr+H
O8hBXdDCUAa+lIcUKYfwP7Ed3zgCZEvGyuCmrsLa2kLcbWdQAhNsLtt4gK10IFCgiEI9oskXP8fd
4ze8SxrHGesJXlu/MuzL5hjvK9+EQ5Z6GeRjWzMfQfd2ZrSu0c+npfiDSIT5DJ6BRd56etQsxzOM
DOY9UDp5gFV9klkTqiSv9x7CZ8JVXmC3twae87MV26hN/vZIkshliq0S41f0/+HCWG3GmGAoU1bq
bZp9zHIb/oBdWBFW8xE2xsAglx9WtmPbyBJeFXf1k0So06MxGmM1yFb/KWKYpREFy0GIDUf+xMFt
cqgRwjFt8jfAT8ds4zc9w7JGccgaTwQsC327ABWBKVdUo7kHvpLMsmIJEzURuccC+mWWD/9pTqil
+FX+hsMY7KnmuPC1evbz+WcKXitGqL0w701Rm16FzAaR9c/34Cl7iWEikjgGt+O2ZdPc1eI3uOc4
u96sPrln5QTxIENBp32Ic8o2eYOxyYcMxbh2nau/cno1hntC7nMesJuT59D9vTcY0OuMValsLwku
bQEp46kRXBFXRRUFGOQFYb+aHAp2zDqOxQ8m/vQD1MZCPxBMmkjH5hwM4QUWLINKl4wkq5Ap/4/K
LCf71MW6S0BB6juuyFKuvyPD5pA5zcpTGTWQYY+ec+xnbunicd81wCfM+OijKZD6eZzxW3/486Zu
suJxdO5JJld/tGjTEVCSsUs+kbs51xsgbSKt2qKIXYAM+lGpla7uk2vrVqRKThX7ss6158F/SnY7
cwIoLOcrkOtuAHitt86IxGQVTtAPkkLypgDE9H8NHfO/UkoKbrR8lXUcf5TJ+WxssDSBr7ls2Fy5
9xELf7hK+rYHGb0a97VPAB3sPwi/882nvV2f3QaPYCgJy2EvCIwJto68jdq14DuWz6CBAcrc/l5C
Wf62MZRZ4iYpoQUIor8iwKrH2gNaAUpHpeHp0+5UUtUHldooA0dno/+vlG6xaCpaAK3g77dA34R0
CrVD877PxBeB6z+CPvSse/9nBrg9tze7bGSaTxhgRMInruRPBOhY/DyCbjZUwQBO1oPUy3KaPCyW
Wq/LyVpdfYLnRO7UxcQz0VL+iHV6vDbVrj3dE5Bq/N4gXyDogoU7j8ByMSwOMe/1nNRc+PQREdeG
VI2UExLXB5SVre/THb5Mrcx0ImUtLwQzKh+2Tvin5bWuhaUMURsrmD/DCZ6RWyiXmInmtmH7WFJK
4r0o04C1b27MRJS6VbDogItpSefp7C2uCIT6oDYLvHr3AoDF3vh1Tbt1IdJXJz3pLTx3lfX5zcwd
R540ZIkrCqQeaUjM5HKJfwLWvnJH25FAXL38zeauy3OTTO3R1lwHwbSmu7k7NOQJvjPJ2Tws2yXu
G1zw//s4FAuqJVVBUcmWb4YkrMWRf0mjRIeCZaSzpAjNKrHyhtaYTJCvZGzLHi36MH0+q3iBD+SD
Qg/LfTX9GPQ7IMwzuGmOK9SHTE7ozpaQ9EVz6It6NPdAzHPhdkgzps+QGSE9WDjKhg1uCTlyXzcx
jcBneiJ28LU5N9IEGDzCKCd6OY00xwLalRc96MdYlDWQbe1Pijg0MPngaObt2ozUSrnJk0dUve/T
0+ApbY22KSyw/2PZmlxU5SKS2j8Vw0FemEe3ykvBlyWYAvN3Q6Qa3XHYsFZXfCqF/NJpkPB62Kp9
/efk1kspIwRdtc+EcjRy8ktR9resTy7sSJVywy/JTv6+yeZk6HBq2GLOh8nw32irFxdNe/ZZLWMk
sdpIrvj+PdaEcXQs/RVE9Ndu3H74fZDymhYbw3OyIxxNCVzR2A6kxIeAlcEoNZj3VCShazuFNsma
njL+yyWPZb1t4gABs/GIBaktqeUR61Jbj1wkQKvfQT8UtTmcsO5iQYJQRTXen5+lBxSFceGghbYD
87kUzmDKK3qa9vhJh8sAW5nD0iVC6x6Wydr6vEISBTLtDdKlbET9Rc9OPL+xpt86EQvRkHM/zEZb
UoYtHeq+7rcgyBe/AEIzNRuUWc3iB6igEeWjIgn/M9QIiuYAauUQa0NczO8jowNZXq37x55vgSJZ
WkVqTjVvLro90jrjUpn5KvHSv0oZ5J6lqd35AuRPiJePcDSvCnZIMjBtr40O8TNZAEvYRj/l7Jxa
WGnk5E4pKtATwZTANsuscoeQrEvEDzcqmlyfjASKzpK1a611uJKr+jKKJ49/0Fi4P3Tkp/L8pgSs
XQndLRvGanMU2XDaJcW3xuNNCMfB2TtpXvgb5h+LE8nlcL/wCs2g+1QaYQj68UNLoFoLAv/4HG3U
OkxNNWGONmLYjlon4nTFLQJWZkYEnlZ+2wXp3z+O4YFYu7e3GJTK0SOX8GgkkzwOWIR3Rbxxfb/Q
INNGPBkm2jPvgxsStFhGWd7cIZyX/jgt/iE485ttMPgNIuyaoANNyGOOo3ugi3TXQSc1KM06A7CJ
8TZ8R9Y3mPerfOsIAV1LhiLqALN6/L1xcz95axpUyGL8n46MDi1OIJV1uDMPqymmQ5QKkHIUk3kC
GJ1g3TgBo6xHPGpd0qAysHAfVNNb2IpNailXj7OAuiA/KKck9/Sbw2La6/eEQ8vILqdjMwvpPAeE
IrG2qdDcJPbWkY05vkHqS7iMalIeF/IPd+l7oY44G3fhJKWRkLuRlV124i1LVs1UImux9iuS4hhV
ZvzruYe4mJRGZ6OTBhhhVZxGAnFfwRPp73id4Y89ZPi9isqbues1/PdTZ9G31jZFreupI6EA3fAj
5M+I9J4qcDtOkIwKfI2swxzXKhZSiMqKfHW1LclIASBw2QaOE2U2mvfjjK44lRB1rXe49HROR+V0
NDKuFt6Y+ElxSJPVqwBWfz1zzQqis9HL8hzdkj3sdS9UNYcskQlzJ4QhExR2iBsX0InKrhEgngaV
YrBOwOq5YecgiXJKgGPX/p8dJ2phPrr8t+mX0ZbThRq1QvOpCgp/SihiFIMdjHv1OyrzXDi8vutI
O4j+J1s2GuftZ0Z/BLkAumeXfX3OH+1qfavpLqRS09CEekhIY+VLvYLuMKBT5McOqlOs0zcii1B1
JgZXlVMgEKkNcLiYJcmSK1me3pdovObmmTPqQYpa+Ud5OLJLE8oOqQ0o/Px9pBq59OTWrgrj4Jz9
FkYTgY6JZbH3fwHwYwtvwomKFEhCV/Y506YOiDwV67ysf7L31Hz8sq5tkmdQejj0+7MTd2OTKJvn
0kqM8J84sXYWp3qUjFVBpj/aeQc+M7+1nlLXvLCWn2mmk+01qgx8UqS68k8Z4Ln3u7x0G8Cfv6dM
UmB0vwC+e0u+QfphJ+B/lRHU1jARQtgYgSaej/09tg4w4RG9HMwmY82HEnAsNnu0xuz8kwKFvds5
pjgz/BzW4sVe5VjUxXNSauqZvAuBPnX+O01QzKP6hQ3vLTkF4T2VBskIEQxLMo/kz1D7OJGaO/ld
ZbSVXZABMMLroywxF+1HSPTNcJu43iTy4ePEjyDioQQciFanOq0nhZWCiDQmdGVBd3KIq08jnb1M
vuWPuyKGPl03/LhX6QZIYvyLv1CMzTJFxRDik3e4bpyB+/eRyGk57YC5B4Uta65LI/Xo8RQjtdSa
mgK4Dx0dkgwEg41EL5YplVispGsGwrNAhe3Xq1fU7KzR8iSUBU1T2I+zzBYGEjHf6x8cnyeGJPUV
P9iuZQImrpf5GzpHKDwIuxajgUoP3X2FEHDYMg/5pR15WO3vn01cFYkRCQRbqiAAcLVcWHNo3G4s
eaSi/Va0182+sWT/JeaiES16tBfW7EFggFxSWTsCgUc3xh9otDS51hscVhiMGwGbUr6iU0D/cE1S
QSlTo8Mo//AsLzZtvqJyyISDKEzziUQaF7cnK4YvKiOsqAzXmdUznHXjaqZCHN06LL9o21A8JveM
uo2b+m21ZtDOHFkU+71QcbadO+zaL1gKN7Rimvke/L27roGMYstH9RDUI4xfK8HDvwOJGuoylbsK
fqy46aIgQZ8Jn/5V5wgmfP3QRcu2cZ1e1rQuTATsX7K2HMXvjU6qVkv/KdZHvx6vV1xtBob88IIf
/AjTxy60tcD2fmu+2idhCTyrYn59I62mMALqXjiwr3TtEIFj8XMnKijkCYKPTwZEus52pnk/o/ZS
EbFBmRKKIoikxLtuo7q/8p+F/KloQDIR/td3TJg+2nNG5spUlgV79fkqsA1d/LgpRPVxkv96LlTZ
xgszEIkI4We/FMSPXXVEDWb6dZ+JlzxD7u3s7rnH/K4gtF6Xd/lxpDLB2bVs9Gzmbx7HXvAjQ3ri
bnkC8jCemo/RIBer0fz+px3Yz05A02KEiiYAT/LM5Eh+DvqSn4KhdVcqBjfpyw0NkyQbVV5VgH76
lpzBSf7CDo6Z13/7N36pR8JC2X71DmMYvbz6CGXTXNI+3fu+cp0ijSUmB0E8gg14mNP7fDQy3QJk
0yiLKaReWRmfUNDEBuUP2qnjlxOe+qeHT/8OnpHMcxwZoTvgd/tFn8O4b2i4dZzyooEodq1ECxR8
UAJxfB8hzEGrVTyYn62P0w2JRVSoZ7fGcr9vNwKk4+U5jUWFzagD/IzkGyZduOQRjpkdj9QCVt+w
AeS6TuJbw7NlkKq69eSjYd7454wKx9xYvTktBkmr6hYzj7YcsLmmxIgX/2jcpL3tHXp2RVj0rJo4
8P/WV9ADM6mlscIche6V6A/oxoi0xGhrTEfdtmAnwN8igJIctdXUsgEPJvYKFP4/G7xDTrbNe0a2
o5+UbpUMtoGH0qr9OoiJENRRPaCpw5EdNLAPufd67v53FtzOG0ePQoa8kanVRAJRQAqbZPH7zcO/
2qsHRKZjcm730ep5B0ufj3CIWn40vFavvaotcn6LE3wvdPCBQCARo84Ovd70x6QyaiCiZlpSQtks
1uretbV5h30ktZR8/oObXsQ6DxupK3192dp/7RL3wb7C8Der+uAHK08LYAC/rN/n0bJtiwSjQHM7
Qdge9zXmYOW6VJDDyCXT9+4JkfdACTCzNYxyhj6n1wKEZiJtqfHbU+AzDU/Y9Z5fhCxZr7SFhZQL
YBVbz6/zqnk/iRvjHG2QiDSJNY7ApcZIZBiTcvCCOpOrGnVHfiU2YPM3QRYIy430/WwyCY68R9IA
+c3P3LNyAXIom10gbF1bRwqmUHzehfDYnid5JV+S7aMTOpsE+0ByuxX9wK/gYi12wL3eqbBi+dsJ
DiHeGV39nfVsqyvqWSxqK453d8skzLWrz0qA1GnyM5EzfqR+L1Itd1HXt75TBhkvf71cP+Bgecq2
dgpSXVkYtFu2k/UQu+0got2lpioTwDEjjImEOQdHQHQOcg/wm8Y8xSIK2mj/+hMAg1U1BEE8YNfh
JQ+pI2d+qfwSD59/+33ZUSpCGhhe/+7mRv0Kie5hLbyiB6ScgIL2MX/5RXTYB/Id8yJ4oSrs4a7Q
PCwBk6RzDT1uLpEsVUMHTDYAYKSIThDLOoKsrfrhilAFjgJ+lc7NCDfjjxSGX0D3pZIZvb4QIGom
ikDnVHy+l0v+liz1MG2D1fcyAhTcwpSvmg6vMcB1t0XsbRXc3txeFh1b7KkU+B5iZA8qHRjENfvz
6uTXVoYex76KqVKKz2p9H1n4LVRg7D3BjUiYW5eawt+OFv/2+OPUgFOvdzL3Iwt1YEMMJNaYur7s
KjtJw8Zm3Dsdb/7hpC73KX9VLrpBfFa4ZlI8NQLzliKzxR+k2sfdKkeyocJk8VYGqnAZA0py97Ui
zfkt/WaBDIaHJ5DHlbvzY43wn1S9zfRgS5Cg9KPxfe6gKwSznRrE9uY/5erECBZFWGaeHMNY8a/6
xRV6jZ4HXxY9Ju3TNvIDqlsLwP9XyCUiBIn/UlvcCtzDku7HJPSD8oNa1YLPY9umIUdVKUPKHQgp
oa8QX3mVqqHjJrz5WVW0KigYgEYfy/4CnPaqAmmEFtQj2DUoPlCUnTcsMFcN4lb0VvGVqRSeDHRI
8qVzFSWD6ikCcxZmNtVbn1dSg6OLUIHeZ5OGaxjsYjGrCiPIC1wNtvWlRRpXtT1QvUWMB9v+Uh+T
+7kWD6IJjYLuBulyp+sCxv9eKWIxiBjE4LZ0xBEhkA0tr1j26uhZ3Owx7VgtDivHEzOMLf+S/cAp
MxcCM/joq051SJ9Ymk/w/Tqo2raXnRPtLJZNb/u5Puoobfgg1zm1QttE86BpzDbAZsp4JmuorDj0
SZJbD4aK5PJJO+wA6uGPuFPND6x5COI1qv6SoRjVbK/DcnPYM6vr4VPou+gxi7TaZLSs1YEJyL3f
rzgHYX/rm59tulNIVkNmvJBR0mnjhDKf9PvssI7IhY9IStKywu/g5UVLCFQ394dQmvuKqP3AwD5P
YJWorcuzLkvABq89tBeUQseRnMHRZg27pe1N6+l5lAfKSu0jrysWfyM6TLGPZtVdJPezo+iejwFV
eIzt+YujOZOIx3i1u2peGEHC41FnQm6rSFsTkwvZYM0pmWOqYvnCH4BrGacjFkJUGGiB5dMt3uLm
u7tgb81WypIKJ7tAycRTEfhk6pudvakw7qW1GgRgl2ferxLEv3PbUOkv7w0Aw/+cFqrb/iHvq85V
MMhmo1CevQqQa8v2v251z9hCmKLUDGCxe9lPItg5NNOVaCw1K0P7o0mH2f20x73LNI5TTHmEXAPF
a5xOXSsykwaEgkGzriSS2jqIr6/q8XNEbiATY8R0bEaMD7kujlfvFivmCustuwA+chh6gBJTXdQj
WuJX2JBjhreeag2/+am8A4Sft7PHcAON7P2CDIv/5wm0J4dNBgM+70Q7mcaML1vNkvrKVcum28+V
10LQHPYem1VOo85ITU26Vp53qF1q8QjLaiHEevLtNC99nwA1my4a3pE7Gr84P7T2q6Om7hA50Sxy
5yKx1oheA1vHec+vnIhnd+7iIzr4F6f0oF3JaE4HvAI6aLFDQFE1X4pL4GVnFfy6JLsEEV5Fli9I
au2lHDkxi4Uned+NO0diyRhbZE2xOvlIbqoZ00YJePeXL5dnPI1c4XW2jjLxuEHQene58HSId22H
JDAJXOUd0lv2VVa+aSic8L0CusAtaFF9BQoK3ipRqPrkcjvpbAQ6aqHjChkT3vIeubPoL7tv4R+R
fXGj317LGWw1P7dZm0U0NDESaF3c4/26PhdA9salBjc2i/gviYg9zrHJEfaszutECQKqKI2JbnG0
v2h+NRni2Xg7pgpGXYDJ7efw51wKG83ADU5Udr2xUf91cpnTbARQM6UBI82bIdSuoHqPa9kswSzI
DxRS3sqTvzIL94rZCDJH0+e0j3NrEn2NjVKyUI0GMm3pIEx+4Z8HfLWTuyZLFsSR32K0J5PmyJlN
OqaFhYHZQ0ml9CPbK1VrAz3UXwCbustWGp1TlCdzs6Me58GcgHbeXjuDDuKcAw10+RKZHKl9A3/E
n6x1kKC7+Bk2FY5BjJxCV2d7PqaCV6xGc959f2bqc4L8UikSNg1WhU98CH2FfSreHK6T38IYlP0l
nGDdKK6P8fOQfrq5PSb9pFCuOoMyKf6vpuzrEpIz3ODdKXix9Dm+ZZP4sB9Qi9NzePCtLtqanUX4
QRCrX6loy8X8d8kzpdVrleHf4Yn12I35Yp8sq8IsSkJ0lX0Zp0WE2dLWITNwsWxu3QfatSSMNXN2
JGV7fgIor4ab0r9W2RyjPUf9X4FttTuwN5E0AwhvsUgQG0AUTnfcVxz49PL+bTBtPw5wjUGNvk6u
NUnQblPByp6MYBI+S9A5m+0uwGfvNfELc9j+7DQW/OfgHJX6iRQ+v0mZ/JeMcOomDXR/oT4WsqV3
9ur3+7l/TEm1Op226Dfyso0I7A6bgHd96m5fVxhKq/8+5DHEraXYDoV9WKYGMC4+gqgyK9rYTuno
SjGjArZAD8CD54mWf/xXFfj2dz1Otj0VlTg2Yg4VIEKAgAQydmKZ4EIWJ79x4UMG+AHCtQSsVX0a
v7n+8F7HnWfYaoEfYo1zrQebLypJ8TByLUZWougUcJRwkQhXpBbA/2xjOTNvmYGGDGAikl+2DbL2
cjH8s1ysP9gIszF9sNDeM0dRSHsiQdKPZzczPR2zZSNqxS5q6XX5ib/4jWb+X8fC6vExZXbwo/P7
vGXx2Gkm9cSaAjGovr3jHBYkxBUT/mlje8WAYYfiwXmi1balubThGyn8TJY49yENaKMj68XqX/aG
HsTqgtNtW7PViSnM53dRwmxlaq4tpaC7pYD4fxE+1m8LT2+ibvI0bPitboIOnzWNb3LA+PtF43R+
ZdIKHclesXWJkXHfwwFpchihpmZ2Pyci5MEuVBBN7c9JfOGKwFPwtE2AOhXEYAFgkh1AonrRiLk0
pGh35bOKPrM5igCxtxDhFP7De72qIWv+gjyj6ifqNZceZIlzgRX7q6AvNoZ4lwKuzIy4YxRBuM50
bJL0vjcGUnpJ/PYyMQ3PWACar1BnIezlDbE+u5bZ3rUxsi9H6hnTtHC1j/SOIVpNSYXx4+ffB3B3
iD+bcA4tCXLVoGsOrZfGTrQEZAlRjA5rTE6HQZG/8n185JZ3aWBdKDNK+4DgZmYJZ94sWpbVry3+
zchi56SxVUF0le6YG7jZtc5uDIDnGuLANQ9Hhl3AbfCgx29O2mop325LRlTNZVd5uUvs6z5bt8vq
XQvNfXfQ+GWV+EEv301BWUiQASxMxdGSZ+s5+lc6Sm3x/cFnDbERc7mlS0fPBwK2D7w7909ppS1u
sjeYrAJJuZL2/SBaWiUiR/1zgGX6d/aoCt6NbMOngyxAbnrK73mpVEXvP6ZrdJ9FdsTit1w0Z7WF
uqaWL5AZdBFxvwQXLxDhtdH5ZEMPgpYXcDDkgFj7sAwO60HdbpkvMhcW+00BYRSq4knAMsyHMBq6
n5TzY4FpVgV4SGbufTlKW5P+iUyuPyiRj4SewqzD0oDPlnqitMs8db+1U4ZdXN7ITTWTZHJO1Y4z
Vq48niE/RwklSkUwGDfjhJc6EFN7cYP+5Vuu8bGSJVpqN9QH2yjhjVOPC5MkF5YLIio7wUlXuDYM
2J3YjPUzWw9egDaEqDaboa62udcMIiLjR4YuTuinim0J7Wm93Czj+aE+qieuK9bdNrTz7a6jsDKi
gcaYAquu7DIHkahd9ugDuBDQLukCQDiyYh+QCiz4KRHg6/GiMk3oHAQlrv8uvisc7biNaASNlB2f
2pU+ucjzxJZlmTpVaYUm8owL6F4aG8tB6nsnGNv2ri2Suc9zqa+tkVASV6a470bMrVJZD9B/I04m
xytFLAaCxqoxo/KPyUqyG/sWQGwGPbnwuoLocyJEjHb2u35DBXB08VrSPkK+QxGAsAEdusvaKrdY
jWdCpKHhHxVbhXqXVWCW+IMDb87ujb7UmM9hGEHItsdtnFCT3+H25pD5YYOnX5rOVlOEqMb3rJ0D
aiJQEWVjYhJlHCYcavKD+EIQTzBRnusKl8Y8hg9u7ny+5NGkbgSvu0Ay5E4NQ29nLNQXcEi6kyJG
FmotE5Eri/RH9XbUgkKM5GbG6s2jT6DS61l8xnNARpuBd7tuBNFzCM8zBeNIlM7y9CiUqCxWYp6g
dNO/6LA+/pMYfYmqfaMCa0vieJ8wzmwc1cFhRLzylfq8hwhJaJPERoE+42kRD4Ze0nN+AEJCXJcD
hoyi+NCjcQLsEUgzMgv7o5rDYOWVuj+E4GgCmAM0d70teZb7yWBSjJjF7P8XHInVx1Rmhcd6IB1q
F7Cq8NY7KcJwzWmE9ad7ZBIcY4DjdcknBuKNQ6IP3QFuzPRBfv4ouPf9f34Zs7D/EV6yG/9wwKx/
IhETa7zgbVJn3NdJj3xX/ZxyjGHtxomTCyU32XfdtgM6KJPpKx4b/2J4IgJzGmYYB6066iT/fZNG
44+BuPSSb/kDzv180EnkS8eRsp/hpr60izf90cikO5/pbE/d134e7EcI5Le/ikzksFv0lR3zCRsy
IEVD+10gMM5eMznOcKrNpLYtQblSM7mIir4FKY1zEqzLtphO7piBR/CiAzCKXpdo0wAnZdpnONw6
v6I2OfXHrb47ScKxJWQPXthowxOOE4sZ+6GUqti4aWPCbQUQMOTMhIWKISZrUCkjZUIIKI8OGaAS
dj4m7z4UybMViyuj9WSYGpE00tsV2+zpZEkCpJEJv0L2F9qqKLhJaJZ3TpXRdwAPDxaUtLnDtwiu
nw7OVcfOxxu7zU1jxOCPBkGdwx+PUSb6rKIrL8dAIKibc7i/wcgSP4GM7dLzUgo11mD0L1VTDGd4
Kb2Bty6iowuUg0+Z3deV+ayFaHEN3hwPXGEeY4rcLerugbQeCfIFo/xwedm7zb1Pbq40oyKn4l4M
yZyvoBFGE2wgM3kV7+spRzTbJhx5+LvSYRcuKfXTCxxZYWM1DlcGj/MHAeb030tMFcHiid1tVAHK
Nrx3MOTRCzESTR1znzXk8sZ/qillAIzt5jn+RHQzlMypYSDhNG+sFOAbTB4VY103r0uSNKvoUeJ3
R3U+GDbf4kXkJvBTGj99i2bOcIpN5IWBJ+1mt8PoXMXmgzPYRMbYyydtX6fPoRLNoMXVpfOsACs7
26pWdg7SDY9JPNLNiJG2fcOaj2pDAN1CmOnqFn3tagCziiLUdR/ALQ5nUWUKH9xaAqyRxCCDu7VA
jvAPmg6dMs/VWcVAzkc1gUrx82q8RC8Jqqx7QGn3/MXw8DEW6KYszFdmbTMcCfjriYGncYfHHodL
H7f0MOocm9BXrAJ0ouRMmulQSxGk74GQAlxViGBdMscNO1iu6e46pP17mIZoGkSKnDLlQ9F7Joka
H8Yz090EApd9d5/Rzb5yjmYt3gUszInURrN6J2npsrNlTMPbLJEcMF7LpyX5qRP+SOllcwN8enBX
43T8VIvqoc1DeSkZ/OUqJyQzkL7tLRs+KjhYFA1siwAH5GjHcJG7m8nN+B8B80u3XrOnN1l7C38v
xeyTby9lcLbllfBv4vuUpAm/qQY7TRIPQovxyA1X7HNLXEaZiSxR/pjUBSKEWFC8V6cskLJktnx5
Cf2Gp2PLLx2kbxvFSX/hd6p1KjgcljYkuzGxms3ZpPsamuP4KJKQE8tLMeH+O3RF/5l7Lqecr0Qj
PehzNHueByq/jCT657nZXNZST8m2BBNNCNLzZ6boGzJBj5SIFBBOBmJCbK5QDsdy9M+HuY1L4jv/
Cx3UQSqHsMhhiSBl2g5mzEai7/Sa42jOfB+RXXtykBzgSQSJQ94W/GfoJXJLB0WY0gokvs76MnhK
T9uAgFfGrTxuApDkt30UE1D9M+vlNPqx7D9J8kywAZThYwweJTyGT64ULumbScYZETxxIyhPs0Kx
m5Y7XoU5m2Hyt83TecEkEzkdD3MGFYVAZPuLfexBB8WZouubjX1LT3MjF3v50CmvuGt+20YKUy61
2GU5XjznYOMhhZUgeX9ybXYt6hyDvgWQ2fYGBj4q7MqcgsZyR8NWN+sldPjyMKjepL+DTMEzff4S
xWISV2nEap2CPYs94LwMRU3E9hheZZw4QlzG9K8huok3P8hgFtRDLDskL0OYazt+VZAqXUfXEpGd
eGD5zxSszro5u3jcDcAixwZnb7yFuy0RCx+MSooLPrXwokGIx9dzbIGatdOeNijg442X2CRDtoBB
1CwY6dMBc1BfSZVwQQ0IbcCxAqHB3iTwcVLslv8h/CyT8yLlZHAmI7uHtJQzVQmp4Ntfq0gO15D/
MFjieBwNSGs62sy6WZcF1de6/utLrpGX+eJAh7ZNCX86EsA41aiLgWTlPcmDObibFgW++IoBp9wx
732tzu8hSYFvY+SZRB/kKbfgaWk2WZdVxmpEl0c7Y1wl+4Y0jcDtWq4nUc3jn/1jXEnA6MYfvmNg
Ao1PJawm5vXXi/Al5pLtZ2leRXBtNjajZ222WDeiy19emk8cVkWJj9Ae/LDnUUjRYiPd0Zoh2w7u
GjZc+PAlWt1xVqclETvRhWlu4aaCCxGPhuB1J9uXoTgTrsyV6lOSpSNmuyuKFtN1wsAbV39eY+FJ
tyWR1K20zx+E2Zdah5otRecP4eNBUI0hnPp7d4f95sn5vnWVi2ZKnEqzn5icQhWetFLI5K5hEBx0
6mssn6GLdLwt2/BmeqTcXb106qrquOU+t0bIoEZvYuA/rnt59PNyKwJ423pj4iMf67+dHv/r9Q8D
UW58OsrJODnZknkd04fAKP7ueJhqRir2InQze1sK3SCtTqe67Wp32T8JufVRfyGB6yhw7d1Z+Mr9
WMDsC9BkFh6KL/KokqaBzonxnM2Hsp4BaeGmBJcC8r8YOPZ173abD+N7CoPfMV8/1QzKz4N357CV
TZTMzv5nYiEDpgY2Oye9T1sXiOkiHtNTzy0NSThV8KGFPm/nsEIMsPA7bQreYTK/8VF76+sMaTXm
9nxpeKO4fiRQ5TWVc4bWN/INaSvIt7Cy8GhqquldeyUt3Ilo5/XfWv6v3asjVODbUBN6oYI7Ob4x
9SlksNu8sxEkNZntx1vEprRfXn0EVxDylnnQFms3KaFLzuTkBmvIXrSoq5Or0plcm4uS/KZeKAKB
VJH8O9umUQZ4l5onfmiM5d7i2UKbWzOYVN4cCmLUpzHpswo5uIYaFwFZJfpwzmhLKKfSaLCA3biP
/NmWljO2HWHu6PuKXZqAIQgY8IOEyoJsQFxCmxFZSF5qfbnwPi2F2BYXgrqPRct7pmnSm+S21CnQ
qZf2UDqvHoucEFhYdhsFgV/lXFlH5KTZ1OGkrP7nMnq9tGWT6hIUcgWGKgyESRfELLSF08Y0DY+R
xSDAYJYEUp+I8o4rFGLSuCxfnpctC1CQ6NTmMofp2gAWPrtIgvljjiLWHx72ci6LTPkEXJueFuA7
G+Nkgo5u7/2Q3RxWTjpRgBY+3nx+qL9fzkCUFVXxZgFZzNE/E80PtX6hhzZc6FWHN3ko/kdUT8sb
8lekUDTD21PfMTHv7zh4T6Z01xVdHb9pSf4lgIC7ZTJZc5UelJCUpblmDsruZFxLc/9bh/BXKBD+
/bTDIrVBaoUc5wmv9iOpDKOUiBvpNEG5dQ+4KDvTVwy6wVwrr3C5wxh89GwhXxcHlsGTLUkfPnTn
gtqqtZxi2vKoNzAQDo44TT8ADlJ5DllNOGnrU+NkV7dZAYPaPOF2xPHA/7cRIYv+2pYNCnNdXH8y
aMVbtzeaIg82WaUM/Vjq4a0qEVO8DFzO/2Da9jRIra1XpL+NdWEE3roV7gqHhLeypLNFd+xlO7b6
cixzGXI1mPgfd4fO/FRZ3gP2tk+b0m2H8IeA5AuC3WbxVv3aSiSSiLTItTM+xikuyUdXtXilIm1t
4ZJESzSq4EI9EVgUqxNSPWAEuEsUmS12RT2IERcw3s0occeiRpiDaZn2KnVoxfH6KqFz60ft0s+k
z4cFtWYkrUIaMRrbE+h+IRv9RkEaEBaWTkIFS80L8S0gF82oDaPDRb3FOzpn5If7TeMqU78Kt0fW
oJ7YAeq3mwPfgrsPuoN3A7OzRaJzCOIYKlyoOeKSL9MrnNM0ZAB0bCrjZ9ylzqf1Ne4e9f95DEiN
1ZloShBhAVlxVPALdKa6TZjrVphB7U5YTdQ9fCtejaQ5rXWxhjGJ4AFCFzxFJHLaZyHPiMHyvbsB
rkKfizjr3dQneX9c0gaAZCTbcFijEJzwTgDGUYi8e07v9cvAHskYYYAC9zqZfL4h9O2uBetDTwjv
TKjhsZBd7onUQ3OaZXUXgOfVMf4/COZHQYVs8exQaHIxGMoBHXcGFwi+sjmxb5GtkbaELrwMtAdu
Dj7MYiZ3o/+mkPQfJfc69KDKmRd8z2s4RrY7fBAEeeEiP6206DGsVKvYE5XEGDFvtsfMe9dFynww
bP9/drMcqWxJg8qXp+ePgPfZ7Ok+7LzZPfslun+uXdlS/ZZTUdX1fRMM6l1jgdYuL+kYK1iRgoDg
paSs8P0w1YMwRabHcKPeuI2XqlPZRl4kGymV5cnLPxZybNWW5FfMOSc+Ge+9xWFGRaD4m/xpqYxj
F5APDab4wUvxkOLy5VJIJ16pyZjKrgt+obO68mBQTNKpWaM3Mu5rVkh81oL4vki4/g2e+ywUj2n8
Qjuj69XYY8BkQn2nJI6ZNeVoqKoeyAlWSsVpep/OVXwPozP92EEJXYEiO5xJUVn0OQSa0ydtuKEk
ZKiHX5uyMywfixTwod7bm3Hu34n+/9g1jP9obfY4TXnf63+xSOiTR8hYlisCpSiG6+AH3pvYjUmy
wZf9b3KKzpP6MQyPwh83Gmx1wTTVTTRjZdwviSFYiTWX2v4L3TowrgdOI79NXDxWZAcK29ItklXM
Q2ZumcKPmdtGHMSQeZtVvW1JbDHXwqqVFuVshTq939PpmQvxb1RdctverK6g7vdAa/Ll92Df9u3t
U1Vdjb6TsW3IjaXizH4sJ4rBqPUXnE78H1vN1LWtNC+5wWK4epT0OmPokfTlNCok4d/xPobre9oK
/vMOTR2Lpcg83iqzPqLp0DX98w/Dh8YA6AZJxt4kRENLz2ge+Qje7bqTc0rtcUw5NZrAXvvb1dKc
HSlwvZV7aD4/dFYeTDyUFH9nQjoFN5MzTiOMttUwogCFJP3VcBsQli0EaLnl+ksVn/O87S2UjLdj
dMXW6ccaaL72hJEg4Cf7f4xDbQuwfQbfluvd+2E9oKDzvnRaTw+6cICzyGZFPhJqFjMWSSpvXJpt
ebRyq3SGccRQ6iHxMKcJumxl4B4rjXwJTXRRTQ73P6EVgSyD06t7r0oThUxvOlk7hCDsILwEQvWG
hkFtObA+CB0kdkJAb1vN0Tuvo5iWcT+WbEexzGwnaHg2cum8FDNn0t+Vlzni7tHgAGFymD6FNimL
9KqElG23VBIXjKrVeNhXkB3XN6hUmV5piDtiZfWSZCpbH8J1JETYNLEQj5mVCkE1uoxwejsVwfC2
wytweG5Cl0PvlqcGaIN2YwRSKyyKvbsbqbWaanZWLkZu3oN4PV2w5zj2b1Mbgexkz1CxATFmSg1j
zeoxCrqimZRj8YrNEAdTsxl30/ks4zYW1hX68CSugwvdD08Ry0uvnmtU8qmBRtd2MEqXqlqqLyoL
USuodH4mAfUTz4UqCcmKVaj0tUdHvp4grf5v3a8W++s1jdd1NbGVrtcB9odSJ0nfdq1MuztQEIZv
JBjEuuOvud/fCt4CI/S9hzyAyFWUpZcFFnEs9k9YwZILQfXg4Y37h5ugvjvSB2UbygcV9mYU2AVu
WEJo8x04CLtt1qkVZGmLVO/mQtcRyrjwEZ1NCIruI0rSPEX3nyA+7sZU5lP8+2z6nDsvKFSzTtd+
qi+6KcFGPAselCnGmftRbvOPuY4bmTumuzfsztwWQBDGnR31CYtN9+vyiZ65OrOdcWbxA3GXJRRe
BFP1+7qQCZ3+yRk4GVLaNSOEf/HITq17d6k6cOaQeNoyv2q9eEsOWkSEKBzGbjj++OEQUtMfFwta
kO7KtLWPT17AiGrlMLkIGzi2Em/eVnmNa4QzttbIBR8RG3kzgruIumYt7Qcxl6FnsjdSMoJ41Wp+
3YdgNAdIHUn2n2QSB/3b/VMXBDU6IVSeizKJoARY6Vkd8tUDKcxZvZJXlxoFZAJwNygtBW79ZMcF
2zjaKJmotWJMOUlrHjrUomLxIIL8XdRlH/b25RXjVqsPuhRX6NbVsg8bG5vw3rM2lsOZiQurgUH3
2ijQFFZdtCwNE2f4Zuz7aTWkvXSq5WjGfuWOJyEDEE8jJb/VNChgi16fhUz3FGtFWweTeS+X+dUH
jkNrDaXt+Y4OnaQsLsipRgpF9rwjD8zP66IzET3RqIIYtUOJcuGr+1xLq9nlLHVVVCM11REmqA5u
rkUwEgmn+ybck2U+fp0CdG3xen6HMQLxGEVY/DyddY20EZkg1lngwagVcTe6PqT9xLeYDHsRtz9V
QiXZNa4uGsnbbg3HU5Gy/dH09yoD0C1GXTuOxtwnj6xSkySrfdtjxW2ei7wV8ekRb1DhFHLrHciL
ReKYYvcaKU6Ifi7jQuh6ZuwGrHtfMsS6N3lzUZKfSczKeBMFQN9JzN5u73FPagzcc4bE5FBNHI8u
K3SKGNyKBpgbTesKueZCZp4LB2C2jEk2LRCm2G5kB5WNb/pjANC+dzX8a7TGHS8u8Rh0n0sIqRb+
wTBv7hrVCiuiSir0A5WwXCAlnoQAO2n3olShpzgp7H+BW+c1pLhGln1pUEbrfsbqcY4P6N5ni+tD
R6mOC2wJ0AFIV/nJpk/SOMwrXhtw7892gJy9tcjEuxsWepMsnR4sgFDI9kzaVAgnSmbzl0CnhAQd
oFu482S4Ps+hmZicdHy7O6FQHpMXOWMGei4huve9bk8ba2OInNsh5/QXscciPq7cz/mLtainT3Zj
2uzVDuXNWhS6WLtr/suNvlXoasOc1XT5BUQylTRsXc7PqnDLFcZrqrHxefiw1cOCwE+gQMql0Qc+
QM24AzbmC/n9jBbPCpdWNDu2pnOYwnaA1w0ReP6KdUYuLencAIRQ9l9w1MmfOTLY95jKd8lZEqcl
jjqXVfoo7TLDwf1DyEJ5EpxAhBTkbTlK+AS9j2Tm8NF4jn8/wzvv3ixoHIBcsyEMXC2OzurOttJy
ZQ3HrSeZcmWpGYLAhojVYvpKnhTVQ//wyXWcG/FmEDIRjMHUkeb0envOb9Epfr+Lk7tRs8Ohnusu
e1FncfY4kf0GF3N5gaYXvquY1QMsFAZ7MW3pbRL8MZLiCBmQGC8AAAX1IHmmfGzLNdCeotQixgJz
5RBvtnT7IQpfnVUFjxpFcxePnSPyjd2OeUD3pR4i+K1U3rUVtYDnyr8qoz+Tm3DE5D7z7chJPEbB
wy9+RD7k8PaqOLK73obAqxsfTT3VyO1ITspraoTgpl0kmwHXtZ/e3/iEExLhUsbyM9DkdVSDyx0N
4H3+XDrEij/EJgda9Bu4LS+N9mXB5GfCQguj8qwYvyF3Q8Veb7t65XYSbAd5vluZ/hkLLMWFxFe1
mGCM6QfISxVjn41iXErEmsZIyLlziffcy0/XPIJiWmrsN16wNsgsa2a6hE9CUDvVNK7FtMBri0Ds
rHHmyw/5+dEuZonxMaNrAiPYkgN+aOz9acXHirPudvhWY2BnQR4tt1Uxoo+yvugaubO/WJUUeRZm
51dO7r0Y1cQWYIWNQwWuLfT1YElUBwv2o3ZIzUZzPwOLtOmU3D3GuWoZEabmUS2bjqjBe/90qHD0
mPxiy9oPE+VOA93qvIbAoLxAQJun828qSHM3TSxvOLYCJTf2cnI3jL2sEAHvFNzBI7z3skszcu8G
g93KB+xCnJp76D03OL+BcD9o3LsX4pl60cL4p4skdU3reTK2pnBVk+wkbqju0BiXuwhm4Pt49Me0
s+nKtH1bEpuT82e4PPQSZEBUvs0FLbSnvs760/9IgiLtomVEgQvcCepJSC3RhEQ+cPtJy+D2yaqd
D9greq+02qbZbOsdysupSbv6WMw9NU5jqi+kVc/1nU2HrGWYaalpxgAVe3yqQmHRJtV1zgSMH7hP
Nt4kCT8qGO+PmPKfmhbHFn2isVCJeffF1d17t3DUSV+K0qJa6l6QwZXh84jjIsl2FaeMiQzoL0XO
Km627whmioCnNu0h2X+GhbZaqYxvLbZgCJYrrw+jEbabMqTWyij9YSVq/V7OqnD7R49OkX4ZEy8f
sZa1xZPUBOch7GBCeKqeEPOxx6HVQTbR9W9a3SQKjePuj84Z6GhmP6p3lqHb8P+aw6L+4ahveo/G
wmIYD7r+O+JrcaQ98gkFXmVATncfOs5aPyo6xCAoTFSdGaVnKvLi2HeYb2GbUAgmudBYlCbTwRjo
eTQJbuRGh2dmCpMAL4dCSqEQNdqhbJTYhuClIw0bb0ptjfsCtiJFgEAITJJSfs6Etm4OC2B/ZpCj
JReGHosTbE/76AvllzweB6zB9wpLvxN0NsVWZEeLjXQl0ejI4mp06ZC9svOZsUQ9XyF7LnHGfQ1g
l5M7NQnn0aYoHF88VJeWYjz83sZogCAE+i0cnHGChNpp9vEMYpyeX9P319hyRnsnaweF54VHiVsA
WE/DuRFjTpQj9EHT38sg6GCg54d9NkH5qqMrLnZzyLx+TaAeUCPJuSnd1iYjm84DirzBtv1pvVhb
TKyn2RgsE3dv0RmF7dOPTWUt6MVwAOdDBLxMhmT8rloCKPJyyFp8K+c4L9DTBSrVJLK74hUThwrl
HaRL69LJbL9ppvU1Mj21o2/SwifcvXOeT02XnBQqzrBXs3BDfOTcyHdldvFBbAQEUKfGMVUTG3bU
PySo+2ROXOkoCAIKiel4PS2zAX8+R5vlRUMZUQEmDXWz+SCN/YX4emBxZuXmjzp0Q6BIBSvnbZDP
9KsNOlKLfamwJ3CbvG3ugMunvIHPwPRTnxqLIJJ24n2yMOpDu1D8g9CLhiIB6uDcggqfwffzqtma
sv3i05kmNwfXp6CIV/9Q2fo8uGhiZcEhyjsjDDsZ60BMaH+Hny1q+TZEHFDzx34cEqmHMEK2HTPd
jV2mGuJjyTxREKHDAUnz8vQfQ0E5tqIzY+2ZL7XN/YpE4wAapyHvomxBjAScUchSZRFIhLDcI8CJ
ynNEOS7rJGlLyWvjvPQCLn+ArRvRXyJrnRXmQjwS9JVO7PPUTFYs5XwPU7p6K85wEWkchn07dSP3
2gx1tXGWQnzZR0Po+RGt27wDEXHs4BhCh1yH1BZ/+XlsByTsv0dJ9FZpUFg5nzXjdsEt7NiHcr0Y
RPIK/9zOu5CX+GhupqZQDihtOcOQOvsKnmdHz9Okx5Bc5yaPQu6xOy25a1tdJlRZEyeQYY+MOnV5
9n+NtA781mYpVR3VjwJtXeipmmAAqw9I3/Nf4imif8TXiGRtQhgvKbwylQ8cgjXPuMvQJ0wRFdeG
K75r0N5qJaMaIpvt5LE14D1WETsJu/vJ7bzApCkD8LDMmYI4cUMFNAyicVOlspQPxwt/jxXvy07u
PWzlOP2P7yMQwQUMhxptfX194fDQGZbb3yxX7pjkpi8OnntKFybDc5LoxylpsbZEyf7PyDWglTKI
jmOrwZaOQelIxJ7BnjiE/zvzC+zfj/07TKKPmLXw/F2ozQFW5/NYVUkvFBbmjXStprh1NO4jAvy1
QLRZEYUuUBymczKrKsRIJfUjfcaVOahjVDudONYTqQ9Y8BBiAByISOMq4ni2nQl/KtrPz4dXKH0x
u5Jks1W/VPur3rsBUWPV8O72mmIHlTaWsoAF11bdI0JQBe3wbEDOs0kVNU2qm26y0+tLC7t8qh0n
KWrQmtjNvhLjetMyHQPVdXxo2P6+i4E0TI7DF5UQjQ1gNh9gfQNZXntF2OadBCsk5LcW6A+Jbw/G
d27CcyOAt1CbZ5M14m5GlZKtTKk/WS97TQo+cCP0Gx5FR1Zs2wjPj2bRF4kl3vSBsicMOGZr59EC
9YowWeI7TO7GABqvEQTPro09CvWKiz6cnIIpnsghztlAWilIxAhXttRNN2Fkkh2jUwLDd88UNAQ4
OEABA0k3bHU3hW6zVjKvUsJWu4+OenHDlqaMH7Ad7oqm4PhvLNHiZdX/g5xnaOBGILNKsRn1eGPx
FlqZY3ZWFX8R7pUgnEb1qpnsyRDtoye0j2D+dYGftAWqZLaEeoRN+gd5zTGU0m1wb+4knUNesdYD
o3zpm0HyP2qnzUDiPFz6jOxnNx/GfCO8cIJFI9y6fnPnJKbJii02XDgCbIQx1x/qlugFhfTS0q3T
4R5gGzxZDzneUnlapoS8kUnC4kDurJCd4IAB43yJr78FZ+BC1IbP+FElW6RevI0GLulwICcP9o/5
kCxlWhmbOke3VOfvs3TrfH4zPoDVBgeoJyS7lB44g+AjqUQ8Nkh4D2NuD7M3kDWJhu78cQhLqGkQ
Dx0HC4PLBo6XxI8ShoS+aM3c73rZ8enWHjLlPWUsOlYrsCWzGprp2+YnNY4m/y9WO3xK+cbt1J0V
NF4Yc+SQaGIS2GPrUAVvRJaBO+4fMKh63JNVGWYoHG5pXu+E0wulFaZMTbX2j62QJF6VeYbT7HGu
Bp3LArAbNR7C+4zvyIMHIEodHvKH46nQP8CsjL3ybCMEneGxp5wv1phy8dCUoXzrLVChhel/AtRu
knAn5MCGQ0xTYNSmVT8itZT6amoiexCenKhRarh+kt6KlktqCt6U2hiI/9BLreHHrHzEtGgvm1lf
7gVXaEi48CWNV5H9K+0sRQSLCR22d2oe/JA+ZKLvhpMJLnSOxDViUJ9GUvDk2EpfVz+xUOTNYmyk
FH6llf3wIhku9elR9IYCvbVQgrCHikJBUNp+JVM2dHV8rDGcZci3vo5UH3h3QibWPsyuSgZzlQ30
Z6VEr9ddmXy2ef8OZP2hjuop63H6m4fCSOByQqSFv0dsdfINpJ+W2obFXHmxosUtFTVCQ0UYJU3G
1vy6PfqVZRVxvUBK0LJLnfn/X3ukDrLV5L9BYrZVf2lq6MCcFN1JtKfovaL6EzV+LyaFDFwsBeGk
d5Nu/Eu0FhGAQ5y5TCK35LZGVl2+yXuGb9l2Rj+1kvosdzBNwBXAAFlt5u3HhUamZilxxP+faT82
U3h05z5FCcPoXR05zew5IqWLNITWPMxZRc4yvFsE+mY0Ze48aT3Er0U7tSSTKmNx2eSZK3j1/Ih3
ugJJttiiZOXpxE3W/HfRlcCLwVIpVzOlbJMz9CrX8lQxEM6Nz0j3NblMAKdzQPEkmxgBwJMVeCPB
5uSps2JYOnli/kF9ThkwxEyp7nxVbgHavOdAMbZnW6/Wp6GRXx7ZvlFAJUAimyWdD9IhMEGboAcE
lb6xcOcRXEGFirpeEfL932cQ0FvRTEEfHV/19S/llrdquIpDh6UFDU0pguc4sdt0xye4S0zbD38D
Vbi8VgUpR6k7RFWQqAoNn4zfyoW4H2uSvQAw0khyfoN9aOumx2ifJYrZLG1QITlOz6HU2y8cKl42
/B6QnPSCUj7E3Vd77La8d9jMXWQ6D/Y317j4koZFuS1A8tWDJXQFJ8aJjThQ+qr2VEws4y/8DFjp
JSLbXAf2D6x2K4YKL32b73JCB1KN4JJOZ4c8UvfLH34TyiYkNI9lWfuyf0zC2kXV4Y72E8x0LsjX
dnb0Hj9nrIQup18gj4AyFQNUh9pnCLoSqbzyQ0NwfgrtYuSM9UBI0T1v9KaU44s+eOeBTNKXJfN4
utQVKzUZeUlqsCX9pW9E0Lh0GrBbYJOPCi1PJ4ph/o04Yv0Xkucw01b570GPM5aNQIuGPTGR7Wlc
Z2loETMyC23k5s6jh/QFrZJpfO7tv5v9yANIkIU58fX7RqpYakfFgd6bZOzFdejobvee+x1NuaOG
EJnpu0fJXIofQMsrXJEbGJhvrgYxpxzUa3SaHAAZXbyx/sAtk0yljVdpOp40zJvxKAsZsbe4JUtk
c0ieqlkJcQqn4skD2snhXwW7IVkZydkHMuDGjNbQswiEOlVlQXU+LdTuLGbrhRqgysbITDiryG5i
JiknVBZrMZdjjJrm5Zv35bkIrxhf87YmkZ4AsJVHCSnlaC8YR/NS6iTXqbcgtneeCzHWayiyE5Vi
YZp85EMcSPqSta7fHpZg/ms+4sARskuhB1mdHjP2zjXZN+TAQMHLhZCeBhA3HdpVQiBUVMoOhORa
FY3rj6p/6dfqUj+pENQPmPr6k8rTaSE0I3uqcCQ5DWPjgdkIJwqqn9R6B7JfrF+gAo+ROHyIoaBN
t9mAbPJx8IrSpLOgdnBmh3IcoeTIszidyph36HSG08pOhyDCfXgVTOv3hoOMoJCM4PxVewcu/Yit
viw/KECeGLAv5cPDx6lT017vvOcdykje8C4FQOFZeCOCbxqd7LJc+/IiyNRfMoMp+83K4vqKReoG
WZAEKdlzHiiZp8Ak5Sd1PM3IxrLxJjE4rXF1qNBRtq1bWdBHkBhXLkmbY1k84w9/OrBeuTCDydLU
NuzfKZOkX9WcpBxcxd/i/1iu2mQ4EAYVlRd8wu1B+KcqsGjk261ASWUl1xWvEIJQPFfojzJ97raE
b1bSELxS+V51yFTCaXiF/7E/Xk+Cp1YCzHj9kD5ibKaFzqqcWJ8siF7HhA/GpS8mCFuR/xNyGfWL
4RDS480NFOjia9MExI6XlqgxIIoHOfZtlzp1a58fQ4J0LR6SVwfzHfr0usWBFfZ2zYuy38qV8BzF
I7YpesaO0CqhjwOV8Pq/Zw2VtZCspv5erpKeMJgqsubaPIF8a1bbwX/TPSWfzoeFoRyc35ujHFu3
/nb3biP5JQZ+GJ6A0qMMwEufvnJpW4dUMtKZZZJdY8o4oWLSoJwIVDKLI+xI/q2RNLNB5mjWVGYk
QP8HLwsPouYAQ0PYovjWh85O1MsIWSeFgwdPrXs76mHGuG+4wtaD6IwlQb+b8lovXZf3faNU3Mp4
a3Xu6bquD8vVz61eAyjMNXtphKfLFLWg5vlmqxwBabQxnBxEypsL2s0zd0dflWK7XZ33VErKYW52
B98VX0EiYpJOGzxYMDCMqnHygy5OZWFpd5ls5GnP9VU4+VCB1m/HTl4OBLOsCEiI2FrpOEPFyNAS
Ce/siiw4rinvNXJkwXSXBLjapwOa4V9WcIHUyhlw/4k0juUYc+FXyGl+J18TN6eMKogyMPOKTwn8
oNubj8QwJSJNj4bAoJsoBjzMOrfmDXDK4sfeOfjCzOZVKfAClzMpbDVX/3VYjJJ5r7nZAEe6zYpP
+3+dGVt2jWnW9m/FWUnrxc3TbW9Y+6sA5lAUdJt+12I6L2Gk6VAx7cPsIWQz+8eIdXmw5VUvTKVI
LVF62IhpflHWsUYcZ+IHns2yfMnd67FxpR/KapPC2AF3EN8w4W1rgVmOteoksAXcGFqYte3tAzFP
v9f/42rsoLEYKR7WPlKgphQqM13J+ItA4uwHl2yTHKe631z2F5Xwfl4CMJ66pYhjhGdi3KLpyxRL
2qeSl/OBdiPe/ZHRltMZVceHUsbTaS2k9Kfxq8h8bWJZc6n9SdwVemWKBhd/hrI/WBC6RGoYKEsR
vpHdY0AjuHCNptOCCe/pFlkHYYiAtG29b2NxDBnOXIcS09TgK2aUaWfSoDv3qjPADR1vlQ4bhzPJ
BegHn90F7+bHm2/2IJNMOmL6/Q35CthHPpeUJ9UTM3yR25Ya7c3p90cLWCxCVewN+t6c29rGl87U
PAUfMc3bHNr4cxb/MKcCKTnvAG2Ti5ewaas/b53i8OKcNIlI5lmTne1QrZoJpmBlH+SxIMbm5c7Z
5x9aJwMP7E+jmiRfmBHSCRClod/OvdOUap2ma1ujp7apIuhfWyRf2d8TU1bX7ELFf2l2Fu4vYxp8
zMH17wJ0CFUivGCnwHqLhlhG0heqfy1gzmYkgnKhdCTkYtLfiIOpEQcr26WyG8UBGO4b29ETSlI2
zQvIk+zqBBafeZcAvjjkVm3ofH/E0s7vgOHZNPm7fozUtL8tFV2gzD1nk9+a6zNvYlKAN0Y2WhcS
qX/gKbGKLx0xL9MZxY13QM51AejU0MNxDSDHKLtprUX0AznBtLdZvNkfELZsl+DnszRiiNnKSYMA
M01jERsMc/fIe18FIROHteO3MZnRyeiml7g++QyRHWu1pfUsFAJydNw28RhGtYU6DSyewyDmi6+q
BZ8UPqWZDm9hdVAjonNL4Lg6zNPvKrCBJLsq3Ehq2GmheTW+amqJ8hkHw/Q1E2LKJigvATNkwsRd
sNQ6zB7H76SJo3V/DMh4zCj5gDPlDnMouVvi/wpdmk2JbnOJjDlVNls/KNRuMP/pMGWBr+hoc4Xm
LGn+nwSzm/854SCqjf1sWPfDKh7qZbY94nbs70zMWogqCWqdryx9j7/MhQX9c51YsEmxfa13DMRB
A73cCht36C07Es0f311n8fVygE0N/7B3HJtbZfOGvd/DE8KTdSiNqjuQw3YHmyirl5WQ6QxUVAEE
pmyGkbwfm3xHXdr6GyfQm/p9HJ+AHxqEMOWuRbkOf5E6KHHkeFfgcYRaCml5TwiXOpygj5K7NYfK
sBlQPts/X17tp93kvlFEorCPsY7ZKeP3BgJbY4H0hmMOYMizxk/TQg1aeYsCrl1NLDBx7AX57uW6
ruNer2wkYJj2d29U5afuUFbP0YqHcoWlykkB0dETvnxeNexqzHlT/RQkWNOQGf91oJJdt6wQFd6y
mvlIdpRwzwQU0HxvsLMiW25MFdSQ4YXTZf6ClwTRhHXvDdeoNBnPbzwzMoAHYc0nkUpljWH6xMrs
ExbelOjhJfNTLK+BYTQ0tGJaZyVYDy6ze7m4BBrspWxp51HX6GtyPY8PG8DLqrPIYDpk/+2FLzj2
z3Wm/t8BLhGvJFLPIhKfSQqlpA3Lqf8kGzb8zgWJlyzmyBBCnQnbnI0J+xgkaOoYg0bEKxgTJkMX
8WH9RKwQJoDgASa/HOjajF/75FJWogDgTZQA0I/rfDrdOQ/Uc/0DGoNXy9YeaVGE5PcuHR+WPqJy
mIY+43fJr+kKgqRbNEu6QEcVymnmWgZH3m4JOYZp5RkDGFhkpJ9nVRC/bmHSc6NduG0CquiNHS2O
VF6iAnz7IGcQ7S11SMvyyyYTU9tft9zYDD1T0nkuDINczwivZnraKUgtOZymEyhpimOadcsnMVH/
JUngse4VCIZDMnyuIFSrWyVGxsdv63gIMgxnvOTpZvkdOiP48SLxIqwNgKqjPzXK52QJeLt2/1Fy
ceFNX5DAjuvrvzi6Rj0zuCaUZ6BXu8n16BzIORgw7asUfhNa/TO0JAjD2BcnYYDITQwH7EiRw+Rd
fdfaHGAAN5QEJseODOtOApBdmkoWANHJvoIWZGUODh4zKCM4TekBU/mUOrm0RlrZokKC6nNUD+fH
hWJQ5+HvQR/138nWBDFTe8SneAdnFZ/+FgeK8LtbvLNdmkI2PzJY3ZELy2SPtqm8f2pNyu41oX88
E4uKd/zl1ugaUq6q6tg+R+dV2KneX3zMNgj0lR+eRkn/uZNOJlDCXPWXyv1vACeab9taueyDioFx
sffuOjNbw1hILlSEayAebJFdHQbunMNf5StL1XZcQROtOo87qS+KuPFLuHddBjbQrucwgk0sr9R1
E3kwqjKGXngIJIOaTq8QinLmpEniW9ZbKmJ/dQKklB1tXNj/M1mMDumcoIxgddXODvf87sc7Rhe5
6tUyAeFZW594V0IYM3Z9OikC6gdj3x3ZB47/t+mDYB9VF4E1M4kPTtdo3viNawrdotcok7J6qNsA
pPPuruHExhMHq65ZZlZHCAjixbiX8a1QF2DTtWVuWj8J6DD9HKZyM2NeJpkmNu3DYo8cTu4jufpB
Gxt579IqfcAqVR8LrDdHSwKa9y1hq/NnbECXijQuNw3fdlGA728Peip5w5HT4Cx05wJ9VBKlIexx
geOflQ5a2cFQ/xxKAmHqrSiSHfb6iEkBJDx0LePLqJeFQesJJiHtfy7KBq+pHYHiZPppoFSdhx7w
kAVWot+1CZWNzYVy1/9m364sZTc3Wxa4WlIfuxvgxpICfxFhLt0q4kRAwRlU0lgaZ7Qps9cIsduA
9poU66DBc6gJKvSi+87jTTWz0L9KpOuLCDzhZMt1gput5KsooQT5mmTxlzVetZ2m1lzXSrd9RRbp
rx9prYR9DyhLmrLx4+SUMaXOddkN0palKjB2cnE3ui3zfG/oq9DPrKgxLbcOHL8Fyka7oWxQ/f8j
mqw45q5ds7PyjEZyisqTKj9HE33eBBXealum9RI4DRN09Ja1iDjLwUe8TZCAB39JJT022YktNpWd
8OGBkNnSgZ4pGLx2iSrlKRSIQIpZ3r5MXee4WoHU0m1Ypu+1/5+Nr7Fni1+zGiL5bd6HUga+RT/5
2Wy+rRbxawnBVLSZVo1DAvA8aqerVV9ryu4EroI+PHTX40XYJlUttKy6AHbF9n94e7Ab6FKTP3cS
UjJBvePd5maRerbvj7u/0zQOc/FGxcGj2lyjmujm0UQ6f9e66CgAA8qoLxbzxkyzLHMbeTs+i8X3
OVHyLDeMmusTplOr8dpNQQBXJkWxadoYDqWhl8FIYtw9hAUNRQYQ8X0UKc+0ZGvPItkYaEh1h2UB
uoMpivUNRv7aypaMT5amZ+tOtlIJ9oJZiGhjJ6g2A5WrlDRXD12+dDIduuPci1I2jmXUzw/02EbE
bxdn0ah0J8jI5AOe0fH7DO5xlvDfnNRZyC6IUjGzH2XqxKIMsK7BqjoOWuIPehuYlIRJe/8XS46C
eTfe9XgtnHwh3gOnbjfmZYjrc9OV3CYPVOPjhWaTmyN+9gTXqYfThNQv9wDGEmTpjcTWBBGoM2ZZ
2FXvfoznLMk4ErC1n5ceBfA7xaYokfrx5MeO6rShlr0AtcrpdLOt5f9tVZFgpQPsFatvwRDPSEwA
54WeR79xZAuMoXI9JlVYnM4+Vo6B30tE+5/HlRKrnYzLvK7skM+FmQ9ZaSbriaSxWaq1MUaP0XnH
sSS1CvAxy7ToaIwOpfEeDy2P1pzAfQSWzB7tBf00fT+2wdh0cML4AZ89FeWh3T+5jGl8qtopFxGV
q8BLdBu5+UVi2yrgm64HJhVrf5z3WK2QmFAWCDYn1UNTloE+vm7qP9Zf+N6GqIn/eN8cPPjII8Ot
l9JN70c9yTRDLGSienlAvWtOVZP71Pk9ALafHuvX6oNR+OzhaK44373FJLeyuOE+FE5oxxpBeXio
pxorYlfhp5R2cL26DXWTwE4NozksgItFQKwcX5hXq5KTWiD1fZ7XD7BXy10oXmK1+C2ERNtzFwr1
DT2MuOwJk1HfXzy+Uj38JdRBDafGhP2l4G9WY+PzBtATJOU9AVvFejy6iam33sS70DM4XaRE2Q8z
BXfXJIYS6kPAR+m0wYXudkRlOCL76jD+sN94uKTkqciD/48Q2z4VfdulzMoXnTjlha3W7P3K2ouZ
SniSO49XGmIDw8N94rJd7Fp8dgcDUzdtK2t63ox0lJ8jKtCr8p78uBXH9f9UDcE1s8wIurrCJ2mf
EYPJd7kpikDMFtRixYzOVyOjyGJpF+0+gLZnKfQPojAmyH/C58khpCN0Ui4X97m9MtOyxyS71g7p
y6KrtdV8xAwlR2Vypce/hTckxOVsP5OevUrulGyDmaXYWsNyvLdiszjrA6j2GlMa9MHjNdvTvNfY
oxxSogHIAiE67fkVGQk8jg7BhPtS6BJY3ZbVuf66P9xJB56/SSvp+rM+4zyu8W3kIGOLwdHsmuZG
WdHaU8fqoeuYk6Out54gFi3aEn+zLzjjyLk/kFA/xGc6QtCYxYey/2RgmYyg/rPdiA12AzvCDc7f
R4zmNqaXphEmV9i8fnQu6gUsFkJEI1KbH7UtwmAbQZVeeZWW6qmOJmf1A2q2b155DKm4jYYeKSJ0
ZNn5OTV3x1pZ5ExmB0re7PbeozAtAvHJ3BrTahf6ikjWNVpyMpurjKHtxzgoI8racWSZKzEsWSGU
rBIormWFUpUrYr1VhllR4hKcB7XsYiTXbImvIeWBayUbE645d1R2BHfIOknht1OaXZlH2WdLv1Cj
OoGZrTEox2TltSNBpU6RZ+4tXgfPnwRmhScMCudQidKhnGjwtk8c0PoBVVzp/xGXIE0SoDO2rLLo
lCaqdUMGPT5PkNfFVzWOJvtdBl/1l14B0MA5vL36k9gd7ya+K2QzewREPLC3o9sgdcGpwXgT57Ki
yQOIgHByMefaw79Fv8j+SRk15R+cap1414il3QNcC6teoHKgwJhwCalrMYTwMfOMBJI/NSb7pENy
IVPBaT2THpp/qVf9LgC7JYq8dz7DoO7bLoiqgci0CbFT5jKu3vx6g45HlSfiLwNA6UrWdA/7fQP5
JujgwpahGeqPQsIqAZjPt/aOs1OpXiPtL3S6/1OaefBE29NQ5woos8a9yx/kU98oQqSaWNfdJWeR
4mXSzTHW8NECuVtqP93SuEohPncVTXJp0bvEBrX2zNey/RQUG3MVIVtBGvyVbMS0bWE2DFIT3Eph
wIU5I7P5WY3yxzLcZpFUNTjBJNKrL+UKRdgXlU5KRshB6FIq958fQAgN0ToBgr/jOWyTtdGWUPNG
fgUK2TC3M4l2RALCPtaiz3lwzFcufbZDarKXgTojzPZ+4oTQz2Vlg7orPNiexgu/26NkzP0KOALY
6OFeKup4/sBcjWE7iIjdO856FL04AL7y9+e0DczvAlNSjq2VxPkodNSrcxj2gsato+Z2TCs9VAdi
E9ncncYkwzAtcEkch52YqnIf6/wonJKDNdO/xbJ5allbzhq3g9S9mxQTCbV5rF1wSexW1hl2GsZw
rv2wJJD/Civ8pFiV5NB9Ez9ubUXn3CJuDOnptGOsbQ1AntvRlsLiB8opwIAv2Pbwi/YFFFGcqJaf
07y9xLMdZy78l5Idvj8KyX+lcEOnRSmBvZ78KpdpomfDRCZIyO9ENuJW4mi5d3dITVByQg/edjiu
cJ4wyZkMRy3aqXtfJpjzwchv/YvW9Tw1cVKKwZPIuY1JOy4vV31a6nehzjqn4URUGrXaNwpFttWq
MCV+ICii2SDji8Rzsn669LLr2HuunjZ0lMZsbXR+uH+ssh2RaCTyHydL4T3VNkG6AHqy49vBHyy8
bLxbhihLc0w5Cnowr9dwb/lZlXFsgV4E5AHx+hxP5A7qcUR1TY5ahKkHVlyRyxoOBgDPaBio8jEA
el9U5iuw3q49BpzIjVVQpvtVp1rUlA5TLDuZ2cDIojdfIf96U9ihiwWvy2JewCALKL8r87RYIz+U
S1sNeXu36QHr0xXSiY0FKbiHC3IP/X8xWmmLVGtMl5XMv3BcVLPbjE4hxUX2vTGbz3f5ui42h9bQ
74lexrn3cpt7/oga95PV7tr/ZzsVN4Nh0fspOuLFYIxD769PSD9PxmdNC9h38ewtRSw4D1xGjsYR
GPPRmt8qp/HuZZnWzGqRCC9CkXBD4jXKGGiJ7jsnaXvg1HXPFRYU0sWZNNOHESDnffM8+CoHYrmd
jspGDw//lTo2muhm6fi9A8XVmwqZt8unaKqk5ADfzCKPnYkaVx/QTkoZB5JZUD9f92oDau0fbkym
GgMrgyBpzbOOBfgyLmOqB64Wdz3MffyxE4jWr7I+ogFYXL4uwuojjfZhKbM0bb5i8+IG/QymJ2WA
Cvby5xklucC1zfSf4h3AhuQG25SWYtmQ3OVIzN/JqP3vu48aiNrTZ8GMDf3dHAXTKV/aOauFPkik
LC1s931q0/7KE1n9Ha6MofX/GBZepyxkFlAr/hlGRFJ1UDB8XGL/FlLwFqluMi1EWLyiRscL7Qb7
aEq5YXph+cdHrugteKznkry4aoacpkL1+mdyF9t6Q7+jNiU/Juc9MYJZ97uTWRgy5zTKsDJtQZ1T
5K/0LLrT1ccw8o3jFtMbad134SLsD75Ok5pcUaoej2pxU6JhfatJajuiDEppJ0E4Q58ggIFtY0i1
Z6fblFBawGQrEtKNn0kOlDYCcXlfMfidLUZuJzUbRypbzAxGXp2piuJPhl14r4uGTvzpBbLr/D6G
tjHnnDa2ZihZAiS15oHwC8IWkDefIFLqEzOqyWrXepoxX9sVXlrdbA22PuoNF4zREYTjHxZqJi5/
E9QS0tl7ui2CXuT/8KKMMSbc1aO8Ua8hj33dG49Jz1/M7+7rcWjr1Cb9hSO667bkE5eqEyN6bp9k
6eydEs5A7KHAGQv4UMjA+0tV3chp6WkaOZFo6ie6z5jkIsquVbNXIYz2G65HWoBCsLSX4OLWU0eM
f3J8b1YwcQHoHQfJuUaK52lqim4LXNx3xD3J4MKm0reUc0KSGMjAaZJtbTdOc8j5YkwFLx0gtIR4
CumTZ1gmiGOCBHyPqcpMTaUCrHS2aZm9DJKWpJtU+SSKOw09e2oA5FG6wELMXnAVuyIiK06Vly+b
J49vqbt+iBGmLFgCM86qHbmWkDe78O8RTi755I7/NCd6KSdDJHcughX5qrcn2cEwtc0UsT4MFQyy
ZUxMFAngW5DlxmjLD1hTHLbdgrBRePnYbn4zRr3VkqA6W2INHMqdImuStFS2ygT8AweIMfUaT3AQ
ajg6CPYx6tXtkuzmMcx9gP9h8QAd48Dl1hrw0eTyilgtUxA970+JTlwCQJe1WnucDeQOo3D7HiOO
NlJ8tXj2Zm007/f0hmFn4Ut0jHYvfM2QABExCAcYzSor+BFtvC5UDOOnalwrHfbHKknox0FjSpoG
0jIIO+T9lNQPFJpHqPlUjwb/a/K6l2j8FVEqZyKuDpP/zvpAmo/j8F3CusVhW0+oKhRTlypq8/JG
NvZybtVIdoXPkYoyS2GsMjdl3Elb1zWS/BzyQgi1sOnq6BYkT0NzzB31tbCiWPF688JGPbt1vmwA
sthjoC3sgypbud+Hn5HOGe+9IcaNFvUaW31Swr+5PeMeURvD2SnZCg1a7LqUfMqf76aN7DAb5DUj
z3YBzzclnegI1ZqG1YUv/qvzZnqhVRFNTYeFklPPPBlFu5MHAbGQhZOvvEgRVxwBwAPza6SSjZqH
xMzUVSA5ubtl1ph2ld0E+fguv5tAEGktX4cRbFbhcGq8zMSdpwBIAKNEMsYRfsZk6Ra0mp4KjYgE
8wzjXE4guh8HHgTOVaZdkJjI9OESX+Uata6ZEgMpujoBoy0UIGQEOINXQhNjmDACdyjk/oNNsfAW
A6QcuvTR+ARqZunvqD8wMZxlTdyeOgIoPC6ywS+F8/TfVpUhQ9cZxVQq30Fj+q/FEuuGmHz5HIUO
AYt0ICLBAmfKB+90xcG50uagKcn2tzp9ZQdwIIC95/Jt/331D2wSVD4EU70BX581j1KozQ6d2WYK
o3iYxZ8KP/ttRGb54DkI69ZRBCEHFjHBUpEHNDRbgmDEjd7e0PnRLTMiPAc0jG2sQKWZC4YablV8
BVzhoAb0boXVVdLx0GM5Aw9gqGFzTS3CX+dY2QJKVsiuiOChejj1aUq3eNHFtoDuXZ7j6wPSoo8X
V88DfOvtzExyCuPQbArrdfvMIU+0buj/OCoR73+xKLtw8PJPKQ4HYXgs5q/xUi4rTBiaAvZspzXc
N//XSLEtz+cFe9oa17DDMWx8U3YIqacbpT2CM1gIqeoVUBn5zjX4ccZLf98GNDsxN8UsKvYZauPs
ZgL5xZnjVgoLORBZc//5wwcL8GrX31qGGX6v1md0kHdvrBbs4yGVuDttMD83Bo8T2+2Xt8ARB+st
831NIiae9/SeDsT51XPWD0mVkp7e6VMRedYhZV1hQM6VZr3FlmRIkwWTi8TmSATGpOGEx6BsHzP0
Y0IniVEsmT0yjvliOzkAW0uxu2bIhD6DytgiMyg1AGKn+N3665f0O80pgCE24rRa3ZdZDl3b7RSC
HZ7JXmvE55ztEJHzfyPWxEph+gopeXRl+WkQITlXlZX37HC+TxNWAETQy5G5hnDJys7N4O+A3G0t
wTUXYNhrY03kSVuSzdTnTfuI324l/EfToK3EWh0YmZ0Q7Kgz89EaHo29LytC+5tJKm8YrEfpz97q
DXvA7wKEPj4aa7VizHFDHHpzm/m7P0U7WwiguRCIuArYRhvs7rDDNp9x9AjO8BSP130QDnsr2Lxv
pC2TZ5s6RnTQeVPpWnRfUtXZZjT2tKYl6x5dzY4wKrrfseykoY0GnOsMGlHtbaH/qSxBQEeOtYMA
YoNSCOGJDaXtzpfnaV/OgdBnFrEhTYk/Vqjjv0IewuMC2pQyaiCueiizWNs5MgVG26WGgnefLLgC
FRgRZv7Exz0zvZyKQglbsCz72ZwHauA46WtMPa0szFABAcoNuXBH/atDfCITH5eN1dUWjiDegFeR
FpD14LCTIKniRLzNiwKv5QGr6ky8tNwUJlQVJFb3YzrqVNBk4fovbZziMPcH7qEv3rywkeir+Whi
7hwpKR3Zn6R84xdveoipW2ibOHi6aWIdTOY+f8nExagpe8Xhvykvu38ZG2px1Rq0bLUJiI41DzpR
gGPPrjCD8hWeMDvaSGZWHjp+PdqMoWIsK5J3p3/J/YbPxvsY7V2Tn1Kqr4BMtRMZAD48PDii+z4+
MupWMfG0N6zaqwsCymadnJ+06daar96xYC/2LCHOzDx94Bae01mFHqxd382GKZ37aue6Bc4AmrU+
Hn/kHfPCY6Tr3v3YJotgaCmBVGEHzcCeuUfQjbAxKH1AJ0MPEyg/56uIQAgpJB32ZxsL9mzwgVNx
4vKGVhseM2rDLYIbSZHxFDFLFUcmqMtoyPgnZtrRRUQ8z+PfZfscoKDo0RNALdIrEvmeipSkkH6K
8wPAU3TIeb7CagLR4K/4GU68SUtsTy16zprC4Y7rQ9+h7P9u6e85V6DiLoD8ZgifB7u6BK+oa4Ff
3V2Hc6QQTWDWRYO8u0IPsAXzhO2oSdqMir0CKAh+XObNlQP0vR1ZIumzERSQhln1/tvFrwDkFHs8
OmuNy8DcmAQex+QbEIRzOyMFIZaP4rr/mQ8T5oMU9Dt2v78BtS9x5MOEF+sTagqjxQayhbZZ//ut
3hdrw57YMAXKU5aimLnWDIj5DJWjl+vV0pEt7BdLAeyV3GoHQGt404pjGgkhAxeULea8MBO7js/c
5j+LTdoXf4BXPJDyBrRF0QIj2sjpsQTYvoHn0j1A9LLvdBO0VjC3irc2zwK7ucAynFzI/NNBZBTD
X5mQAYaa1Q/P6gTJVMBysyzI+wy/m6sYNhEkCehUpbYBmGzpUH1unuejth4D1DMeXQsM9aIFpF+s
DFZoOB/VNZjUDAgOSHyghx6LTu3iaRzxiHFN0Cg2Dac9+nnYLyTW2FyNMp/209yTnsEoYBRyTW82
PdihNN/mXOcWZ/cYuRFht6YJSduEB5HslJutM+jnakU/ZPII3Bgq++C1/efRG+WzKC9RDRX+piDP
UWKy5h8O0nTtEoLgV7DquKbv5TfHByGq8YbQD7JHY+rmC1IKkLuUE2jNF9/pMI84/LL4zTDDl2VU
Bce8ZOY2cfTBneWICk/YSgobNVZGbvXZs7WfDexV0t3IPFQrtDRHTJdOu7/n8P8ab8qwuUzL7Roy
i+mjqusJ/vcHIz+IskU8zrkbGJjXKLkIAn1bYbPfUTbu0OrEndaia+N7lpu5xrMD59qLztg+xRYJ
tuQK/8V4Fai4UsmxaKOybgSfUO0xBE2dvwRuKsaOdtyQdoYE5RfRD4UNmniaIa3OeXtiyNg3QKh1
183iskS5Cz0u+ROVzC2rQwivC421mVBM70ozgETyhvon8ohwyabpM3bv0fHo0QIPSiB3H4gAmEVN
f/KamWSSagFDTMzDlnwr6gENglAYUDyUM/Ugub/KYw3/BosUTAnWHufKERcWv0RANkUVby+sq5/v
AfoiC/u7hsqUTrHUc5cbA2nHDVq3AdNm7lOQrI/VKB55iPE3cjJ7/tWgPbuhsYO7bAJOGtaveOOf
dzFiPHD/0TUbTvZ7b3+rrII7UUi6IykHKGJgsXY7GRFkbiuO461iUroRFdpZThXeUghf6aK0Ic1y
/mpZxAGQm/Z0xLnbSUU/wmxTsl8hyGrG9jMnGdlUCOgITfqd0omSWqe7C6BGlzNd6J92ejx7hwtZ
LxdU+ziBaXuGQEPDO7N7ZDdgzGXvHJUB+8X+U3n+D65HN4FdBiZpxubb/Q6eYY6Fnb5yga8MkSme
KFw0L+FMnf41N3A6VD6f6YJVKQqWYSi+HGUUDUfjspsKpy68/fqAnNNpJPdR0EnhtE3ux3aCJLQt
6qgezjXKUQfxCDF7j20NKUuIDwqYFKUxdMNYMRp3VuVd8PeKWsoR9ER+0ukLNGCCCQEOBRQ4Og5r
9VkARIc76YGxdXcIBh2zq1g/CoG1xauA9uZZidjcvj9yeIc8Nx42SMXl7juaeIiP3fwwenGkmy9S
C+wkE4RpiNmBgq8SjUdTnS75oCOU5swQ9tTPVH8lVPDCN0jV88bO9zGXG3ksxGz51d2vZWLyuYcK
9aHBZWLxVjhTYpxlea6FmhKsWPh5J0LXoG1mSnrTpmhHoW++mhfaznLaHDLxVdRI0t5QOtWo0rWw
AhxKanGV+arUAndgrk6w7wtmMjR9P/wTxp5ntaDn17lqvEnDqEmIH3CeUGBGOOjmMoZYN31kMP0b
Kn8CMKyMRZ7jgv/h0k4ODTw9BL+M5y9gjAAKbGklJ+bl+Zwoixy0VLsebC2kcLbaQbfx8twaFJQx
6T1zKn3hym7Gw5XpwKtXye962hkAdYGA2B7cELP1aNZg6n6B+AnQopJmGdt9k+U1fiJ+LS7/7wxu
lkm/Ilz0HESc+JmrL3qcn9eq2s5ATz+ZMVmV4bdXCm2FRgxZFjvewbO3+f9iOZ3O8o58U6MerFxJ
2rE+rHw9xSSCAdI/+LP3tGjI3KlNUXjXNSsSwYAg997UyYLt9r1Tw8BV09aEfjP9G1wXrhRz8Peu
J2mAINimNR3lCeDx3EdD21vbTKm+MYB53eAqlan+V1dAQGgiH0v8/RymjpAuj2cBYj85P8EJChkc
6YhFbVDS7KRE2cEN0R2g3oCT86qDFr3vivtcWij+vovvzkpRyidAdyXHijTB8ARKmrJ73EaTR8T6
SQ1lXGLuE5fAwAXaWn5YXTUuLaKE6OztWhmtknup2C3wHmzddC0cPYZCESsjirNdSaH38TWlaf1d
41innyAK2eKgdSAfE05JtT4qjwvXyL5RlaPpXsocotEl2rgnHCwPKXrV4ST8M+J+tUziEcRNptEO
/WejOlyXtVe+DXTXtW/7zygH/zrTMN47V9FXd5pNM3pMbuQWxCOw/yRomFgTjcdwGJ4rA2NCDd48
y1dEk1C8WD7UHOxcMol/cPUGHQvdd50xvgTV2F8KQ0XofvWJp7+Kqg8LuyCPT03KCzGDf2BF4/+s
RfBhqu/lJK7i5lLmf77x/lxSsa9H9h6A/whThXXg7kTIkXLeC3Fi+jc8TeIoDRCEYuOdziD5eVj4
UPaONYsIS5sl+FKj83cpaRqaCWcMP0Kb/20tRNfATXUuNMsa2/RD8yH4Vu+z3t0Si8L2+zwlg8Gs
r8/WHiao98lcQAnudpcmKtr5JTsZhDB+G1vBuPoeXixeOUcJ+u3kA4hJfpmRaQ/tCE8EtLRSaGBj
AGMnyDGpRazsZL32cDTcn82stxnxUgY3GQEkNML/r2ifkaCK3ngt2yMBez565Npp9YptRYDJTdgh
FPkhC/a9LBpDBZXxhpVBv3Ax75uQbUGenhrL92ytEHaOkDHDLlOq879k+fCoAUZIXNpU7Jf4V/qL
x4UjXbV8Wmst+Z+fxneoqDcKY+I3hDgd2xoNfcgtohDKBIkB0XiGXsnenebFLbzMWKWY7huHz/ed
dK/jcSom/zYoVkAEBfr9S/eJb0Y0pqn8Q9ErzlG6VJYcOfZC0XxMrREhhfDnU1ZHZnZG9YqyeYOa
eRGv54lkHCN+m4Lxgr4/rUQ24Ox+fBahQe2FvSgPuFcydtKmX+5DNP14QxsTHcQzEOBOzCfm8gMh
aJqQuqap+uJD90VmcrOVCgmb5GfWF6lldP1vOi07CZgaZphYaso1jXzAZm9FXTqpV/WhN4MsCsSg
aEBItrJ80ZUCdjgYd+3uh9GzEgz1Up+wEm9ISO7Kw62QAgqLf7J51xGRzj54Y4Smf5vE+2ZD0dGF
sWnP2KPCRkwlfOnO36wdTODgjeRDz1avTBDWD7/yVzXi5GqnIJpoKSC2uzB6HCTve7l+2DVC6Bth
PeS9L6k/hkrNa9FjsEHGWjztFvtAhWkZWKfM17qkTDNjCqChHtolvh0wudM6PORmTsYY7I3QgNDj
RF39xbFLdHHyxxPb3pPvQ9A83CM3j5qvZrne/Gzr8IzMCAhUnlNTWCM4+P6wCONoYvbh+znL9xrS
qBJdciECGsshfBqGlNcOFuaUbjiOoHC4CUnXOafuGkmCSDK8yZ+MUNYComDqJgRax+wqq+Ico4P1
OajbUN2YcMhMgcu+dQ8nRD5anNB+dXl+vs5/zyLBSs2Mk8TRI6sOTYxmtwPST9uL5acYTl8C/QJR
gCQRv8oSQbGuYNtDCC0siHk0M7nMokpuc+rSFsCVwXZFPU2Li6NXYqk68AXne4Vzgy9hnt4ctJ1T
nnpST3wIDhzn/GtC09xX0GvIMWtSNG/EO9Cue0N3mSCQPvLHIiqwTe6DT2xnmh2lAScNrxPpmz8p
sglDUYO2rKx5pFDA4wM0zZuqAdePZGboSfSMUNsZzrW+u1ZG40V5rFE39Lz61K8uDfhQ6UyLChmz
Fxvs2ra9I+nbl0fxwW5xK0dv3ypTNd0AfzwW4PFjNOwJEhVu9KZUx1Mn+PXmZN2l/dnEs3SUkx1K
ZRT44RBGH09EFRxe0OIJg5AtOH9mhSGcbCMnhmCTgXA266aUNNayMARuFU79rwkIw283sE94Obug
2JPpAVOZJE+ngldrwseUbqfGpxRxvOnrNljKcDZn7173r/sJtZw7yc1xr8K32AgJyOkuL+Bmmfza
d5HrmC76GM9HwCtYGmBp0Bi61PL+l8jIfVoWVQoH1MA5EnUxqpQKjw5+7k1mp/qAXcFyP4wb9+ul
Ds+BsolrHiuvDlp436Vv2S8G+yvMkB9daQK1gfU35ovKvkcPAhB5toqj/PlQG3dlfRZ29Px8jnQX
I8LLCLC8faGn0iMhyBMwWmQ6efgEZ8Wc0EMqJxSkRMPFuVOwbtVpFJdtEoFaFCW9E27xLpaoZNaK
rNN4D9+XyNHpn3zlLiGn595eI5v/EYgPfR2sWrhmmeOY4qPrTr0jFm6XB1CZaZ97trJYkxmA0ch7
sF5EEErkNhrIWtge+dqnspv4HHVzu8ayK/K26c9HHVTA0Y0RkJynCgyn7CD8VaIH7/Q6gqLj3H1q
tu79AF1vjS2URuo5BAScPBZElEVbslueAn+uZVDj4GGd9F/2YpJPgQ9MaBSRbaH8ZGqBUTAaqPtd
bZiW9OsYZB7b83f7/9KXmBpvFXrYMrFENMaDsQQKzYV1UfPCIZ4OXqxveoPRigx8crphz8xQEG0m
ZCXcHPOgH5uMAZDG/0h4oYenrnQd3wjyP+D9wxjg0rF3OyVqC49gC4dlE9NazHKruJxgGVC56Gfg
GKYEJ+nnxxxK6h8Ar1zAP9maBSFQY4Lt0OthpFZScoxxN0J9ot2evFpjCcSFOmWAG0NOiTaauFSu
woOnqznl9y/zZyoi8WeDIGr+As5FE5xNmRdM0kjr5a+rHtSgzDn2W5iDnLeybqav1muO/nrD18zI
Tsx/tnB63osKeo/7p2bHFwAnr1/twlPxDAblhB6DQgAdl4r9gb+niykfNSOu6USwxYlK4u6qtjcd
22sA5QfjL9yTI8UPZ7W7CThNqGfoUvNwEGWxOdmuHvAOT5L/vQCppZojDBdTrZvxMCII2ywagNK9
5ApcwpSt0O5siyU++8mu7hIhhJEwZYQ2tUzTyH8wwn5unkpdjPxXyGce2tjYeEnPpnIBTLh88aAt
1kFCtnTPPHHN3nbC8S4+N9P19HA06N/rd1cGpCOSGo5FcBcSTukLG4u8jPzY2YwlSznDJeTFSdAA
amTwwT+1dZBCG3xQ0BagERCYggtD2p0HDFf+K1pyHfJg+BVIL8h/avGVeVON4nKfHeYcH3Tn3/9p
GNgp9iR6GXN7/kZ7h+cTYZX5RLwI9zpeMd36HB/J2KZIgYl/92ij+5VmbBDxQpQ1+z86Lwmcn/aT
kamdBSAk5tCMXYW1OXGdKWd7GEg/7QiM7vJPJCXsMVI+k9otIREIKEXRvconeIWCoIqRr/glVxfZ
FBzNm5IW61WKI3g1Iidf5Q2sWjeaSyyDUFYRILDEYR7yosJSMmoffKjzaI3EGP7fq2C0HtWqFFIJ
mywiTFuB43uveUm/5wzagu/lLIn2JXyMBZLUhKAeeEAjJT7lePGlbQYGcqY+nYsSQbBFUZ/ae/VU
piJnnrXVkG1jsqKmDXgLCF0qrczM20sMB54w/2o5kF2Vk0NRDpJxbzeCLUv3I40i2ypyULi7ZfOC
7sVtWPPtkpteJ+SxP2RO7pL45KjNdJ9lAMQAVXzpVvQSH2hoCAz9gMGCswlMVgURDmUmSUjJ5mT1
Wmu6fxblXUOYGFzyLGbyG+HYXdSiHRz1NcptP4x4SK6f+gXzqpn/yLKwSqwpUWNLsRuIKDYimHxB
VIKmyTIb4rY251oYIKhEj8G1XA8tQDoJa5BEYHLcQrU+8Lqav1MEsloZOg7SAUx6M5NEmpngb7in
jKC6FTNn34THOwuj3vRq4K2jcMdp6Fmh5CFHcPK7FnCKq3GpTh9E1KjQhK1+oAvj2LcML4i+J6a+
/5DDmk+8hvFNukXL1y6PgaXPdPb4GTJbsSlqbDjmE2H210NTFbHaDcCjNB3+MTXqCn0F5yjywylg
KssjezqdWOsiaQjKwPCrC+2O1/iwPs4lDYFjFzlnDdWSX2gVIsVOOc9MntViqfG7DWVJpvK0rDbK
XwA//VED5gYBZeLnVEOsE+ckMs0IEu34ZlgCjVI9i0ovJbNORCBqY6y1olKoVAO380E73qmzEFjm
LsRfcpwgrw2ni8qEG+wyEWP+1lpCeTK0tUzvSRpVjP8MyJmPg9nNH7gk6Ksr5UqD7hnB+4VBibRH
j+GDIUlWxAg0P+zkAcZEhHvASqWacHiqVDRLjnv9zTWq70+tRoS9QcrIZq3Y2u8g7U+n5lGishA6
T+k4O2TO3ZsnOzI+lT2fYYwJmPeB1AXyqIHfJRH6gLoQfm5nPdQ0uZuN//jfmBcl4ld68fvFD6Oq
AmP6SoGmTqMrGe3vIy22JzkzSxdHKf/7wnPO89IvIIanZEy9wuPxhH8kGrX9hFgcM6C4oOZClZz6
++DGsg1tpyw/EDK/O0troosUw2JLbtxJ1M0M9ExsjY054px8cenXR9eidxRlnpLKrBMQHMCi2liz
vEQ/yI6mjkj4ewXNqp1+K8SALrUm+0ulIuwIKC/3rCysFZ4FuL0OBgFd2j1CSTcBmN1k5llpBu/0
fp+OQULyQXelr0eqW89bIqyXLraQYGsfVT3ZsF78DFuBmxR8/j/OD8W5RUg9kKqdsev0rdhhUpWf
DKist7bHHKf6YWZc+5Bs/wCwuAmxm0tKHZJ8xlWaUtKA/PLrgT2VB5CnAh59MyI1cjyaRQpfMUka
Yry8e2BC8vZ/I49NICKPaIQctqBi+oSRzN8nLc6V4/bHFqYailjpxtH8+hJLk9zsQXTPnkzRcqbl
MARUqLJ9YLmq+v4xCh5rQJD3bl29LurPZqMbu/HlCbXhLHlDb/DsjavhPZWu1jUWEDUnWl+zUOB2
VEikf+kaT/6AyRajDbx41lA3NCrYPLxKk243CF+bSjt9g2N83eaEhmTI4qZQ7LhfFF06FB8AmOl1
EieBZKNdwlo+HceQgERC0c9J2D6DsE0NulFgh7aQ61q0L3Nbr/4QqibsEYdyzoCJUM3v6SNlgzx6
G3DYTBuwavVuy6clv1Z/Ah6M9javMTuQxIH4EsdPwChvfO0RuuW7KyHBIw5Yvo6ro9mMbcSrqRF1
zsWi2Roxy1l9gFKnHsP0s6o7Lmpk5jAAeAQWil0AXuGU1+jYkHTvC7hZg0/cwDpQW7+fMoULOE2N
FXo5lO4oaIGiRLPDC2rfvUJVfnrw874ddefVvGysbDQnsb3un8RAPFIOl8aB6dy+HXa5JLUnrc4O
oKaTGSTleX52v6L0iWCQ47Zv26Z/shqqDuDvkxmslKIyTTqH6CoTv2a6++G9OhGIuChsdSbSlMn5
KPHhmt3oRd4nikg5bxyGUKn8l7TG5pgLjXtXBYBYbM7JdboJcPsz27vOHfh++YUPmn/jaPM/lAl/
DV2yQmdq72ho/FYgL0xZAJUDxrJn9yFSyNNUQnJo9Jpk0OhbOA5Q8irKLI0jMFhxMmASenMO1Gr6
ghMtMIL8ElQu/GHyj9styjppyCL3xIeD+0S7qPZLh09iTjaE1UfrkA1Zc9FdaMhaaCrBTMls+gEQ
L0Ae54cYEK8j9HsnLxqgdmn7irWJrDnCrZaIGQPaTd0pm5jjxNM+7ivLjYeeUsF1lOShLGF9fAly
IrZNakS9JQbMnGw+mTb5NxUIt2AwZXl2uzFGzgeXWIafOCyzzsv2VnXJNVp78eg8+PtuG4w3o/UO
pxWwV9Wg1ASkuAOFDuouQvownHs2kcTxZ95f1PTQ1A6r+bRsz72rPjzdvSrM9vsNyGEFYkSWh+ot
j5NUpnCLO22mdhVYJtuY2Xp+EVz4H6oQw1D2rrQ3hKRa2mWXNP8//D4HzV2zqRO+T0NbPcixvG7o
ZeHrM2aEE2zMZrlrzoqkvblwXSbGI80as0B5lpzAOwc4y14QBo5h/TUoLkftdR7J1ZfdcSik77Wk
wEUiRVhEoFze2tQSd8JJLXF4YZYi7MpcD8GlYQJDvB278PfW2FADbBlHiTuH20Db7iER5fIf/0PQ
scRkyOY9aqp46sB5Y3EVLuahaMo6cWuh6WSd3unBQwlnCUi+hXlqu/3D4qxoX2AT7GUAC++joTVy
1Ho0A0OBW5oXpS/ikJMbxbwMLFaIG7+BPq0tJTJjwFVk6Bfi8QlvSH7bW7cAPQtsseMnj4fR3Yd7
bF4YI9WEJrhK1t6VZUAO/HCZyR794x/YGt9kBp8Hl9SnX6ixcb1A6nlr9l/bZYUteNH7YvmHbZGg
XTcao2yn7gI/U4CDevs7Jps+oPBjTzNy4lPIVaEPE0xm1PGMEOu/J4D6FVr/DIS5GquvCHy6/99m
VP51s5XsKJBkeSGu1OwbXbf4GLQ1BSfIrLf6zZcAIQTh9fbJLMm0MGBTE6QkJ8Twy5zqrwHAjndm
4FYtoSNr/qg+z5Lgi22s/ZXMipaB1PwSu/sNxqJpMb4Sbv1Zoi4PiWpzM39ekkjF5mWcMszXvPCl
D6evy4oYIqJpSdzt0tHcrTVHxEdbUqZvJzT4GSs9nM8V+jU6VflbbgaNcck80jjvq9J5c0Ug9H8j
gAnGP/edBq8mecoumjjtCTY01dG4oag5pliW0bxF6XoUyYr9JVeAjwrq8s5PpHAbMRpOwLSZblI4
VTi9UHzul1qsEaV2B6aMLCO1cp7U99e/QoPsBkejgG0EHyox0jYFKIYDFYrBvNXYs8Z0G2/NACQK
1u+kyMF2KfaeDs7EMJwzWhkqQIL2WM583CKvSWUS2R7zboOGFBZRuX5RnlMqhVlHyAooCMd71wUe
44xl7D8qt2YhW3fX0ZyKNwIdM1cjWqzP4o4YLDoLEWsjlESiKl8Nki++TTt8u+EqY1q+UwZQWrxH
LyNy+ynio4MegbQnw9SG94LmI5/78CdWWwlD3XWJWBlK8hIvMdfhEzBMlt+hdNITgYwA6+G1djBG
mRtW/0KGmbDjeS4AC9ikm9uHPdFrsFci7vQhmRoXDag5cv6P8mEUK9yvbi4ePZF1mzuM8t4jO89v
04ZDzjtOLNoyUh4J3h03bkH0bYWIq7uInePyN8LUhOk/+WBGDdAfxfqnf66XYsWe450MW59ZhpWN
NvktPn1ciqmBBreexKoGBJauW6QecgjBuqclUbuqLt13L6sdxlI3aSx2Yx31v9icrcuYE2YvA4JA
Zs3ckIX7K9N5HuczlTrnc9j7bPUoeTgjMibiwwLw9ddh7+65CbfvFuB8kxGmAhzcZRcACVkIH1iT
DnBammMaw7dSkOXNOFZISBFq1oTJVA+OMfM7eym/P5BM+2L0w734EaOwOa7NYvUkgs65wy/D6xtr
IfHgZRqbm0671j0l8PntVk5XDcjUk6q18d6NxYYoUuZ6q3dlRxyj6QyWlUCfASD6A3+hdQvn37eG
zAZXCZVuurjf7nM9ttTKXWWmpxN3ytuvC5IFFVHItAxXSgA4GZG6q5nwvr5vnsCRxkKvaDn9ILoU
+cvwGJgGledO4RW6AHucdcpHdBXrw+chU2EKNx33GvwG5I1Z1aqO5gC3p8XkkgVz9f6ioX+OdVyB
Q1L4O/ssLDM+3VZa6c/X6O46bYsMCey54mw3lGKseYwX/wATW6Kli3pYeqaGo8QVoPnDHyJ0gkLB
b71nVcULSw2RtJaoSl11DBzIfKhRO5Pzc1vWy3kCnKxBxeucspjb3AgMz7fLNIkLomg7MM/obGVh
NOunKiF/KlnsOAOJa7VWhvRCiFYnAbE6OlnRva4ZxQiH+XZpP5DapUJjbAWD60W5jC6d6ppTeyka
FMJwgq9OY1v8TCdg9bh0Gglt5U3bhZc6QvzgCBpDW0/QA9EIi0NLTrdTp+4WbACUZy3ph5sp2ZpD
K8oWPce5tWXWjSF4erpovuDwFfA+/0koFsMnm6XTidf/IIXPXfhVdNpWHhpxNDFcJEGQYDoEtGDR
Wk3ClKb2VdYTOHv0cR46Jv/An6kFTI8SkDwsKSivcdZt1EC80ZNkbvqYkXjD9XT0f3sDCEdfGH+u
sy8TXs33iaKcU9xgAoOGvPRzvvUR1qRRbCTIx10Roa8v6FIHJdpMfN8Tr3HU9SsmSfSoiFHg1ZLI
qOeNrqd//OjRUv6opHxHfj7fEFDYRks2CSw7wrhjROeke8U16JOd7ZkR5J2jKCJWi7wK6hG5xo/w
p/ZduMTD2u4Jk8K+3i+zBdvvqoY5wLjI7mufXjvjbe+inll9m7s5s0i2EOU2keDhHwitSSug1WHj
lWXC7pp4yvUQiClsEDVLVEi/2bQ95Z77v9LnLJObgsuWtS5pIlyk8K+lI5keikzNTXwYHGedrlVJ
Rrfgy9W637N/B76PbpzEnsTl6CNGCUpmXTgIdjvkFVZjneSIYbDwN1NSyhNzqVyr7EzdIyQj20Ax
7eNkaKshcFOs18EDswUCPhJAqivz8LFVEE5ingT78peaXZkAOStdHqdPF7lLqwiyG091gq1aynPD
FNALJKRVRSKJF1WkzCm+IIwJ5Ig6cZP85rCPlMM6M4dnk3amhj81khJB9Q/kX0Jc13gvreqooJa0
bugFnc9Mm3vZZUfKm/UUqe0NT4cLghHsG5ZDYw10iOkH+PUIwfkeLTZ2KWiLpx6FUNbWwjeFXlx4
dzn3AmzxgSPOcdkPcWJGkybh24hClCVvOMzas7fZc+UCSA9Zj5mYTTDUFTGgIOGFW4Q+jhfKJsFG
2PZ3fu/hGIdeZvBkr9IKXNDiavANDwhFvMZ9pdwtz8VuGF5sl6NkkNicco8P2QynL0iQMA0gZrED
k6k3B+nWiAwgHyfnTX03ymCBs5uxLVorzmQLoQ0KV/4CPEXH5QgjH8m3lBxu96cgMIWRzf5Vgr+D
QTdhll/w7cTNW14eDhgVLH94s9HtBBPLTe67gAY4rdNw0C7oMwJgXSlF0oxulAVB02SuzWbCGIw4
EJT6A/tMiL1/sTcZv5S7hGAR8meLxoh66kRGBHBt15691I9Zh5VFk7Tcy79rVIiGPyIRWIM/ur4b
sX6OCFcj+HzLE57cfcGvMZi99U8dHBbhavhdNwEHzvu2cVrPbzDdVUY5fZ2SX8okDonxDWQP9fx7
6Agb1aGg6cfuSJ10hgHxkcGbstfasZ5t1ek72LuES1VWaZCM1hn0fBTndc7FViRVDaIlTGPjD3Lt
JnSEf91hWpQ3babI3UZSzlzCdOACS3u2Vz8/0imn9jyzM/joWh5Mtslw19qp2bzwFDUiistNBBKw
WPVVfS+0MQdI2R9PXw9OrNFSOiG1XVqJckFwpnE4HTBSZhLjlPJIoB/aufe1p1FQdZMkZiJO9/+4
woRbzU1Wo3CHDPtYBrMi2QYWY6XPbs2r7D9tgi+GgXq1OtOavMQ5UFx57Ytan0lGnkASElBsD+AJ
zRGmjsI2T9/k/oVciRg7X9m1+EcfDNSGW7eD3VW/VELpodseboTfbCHYhtOyJK7YXwO/LY8v+rX7
vJnVTtmAm/nxbpuwL/SmME6r0scviLmgjcBAz9jtIIeR8zTvCuAF1beX8me/w2LxlIlwFGc1V1Tm
YLYm1LWiIjF2P3NaA8ZRsIX01ZGmY8PdDAa7MGSXc95JbMhjj28/kDOZViy/82WwDAAH7R3DZUBj
Zrbl/FiSTAQ/8DnTT/sxP+FKEM8dGmkDMvqxkzTBTkGCk+BQhgoo31FHzmRmSIGx3GQIQy0w0l5V
1gEncuS6Bff2cPlskZYsKMLpLXgILsN/HBeEJEvTHK7Vu68s1Ds+9AXnT0cSglNEOUKf6cVVKngI
uC7QMr65JATanVu5KKh7cs+hCJLcP9iWRdnZFLPtvKAWlb9pqEzw1P9XOrpV6wtyTPAuR9oOMW+b
p5kmxKEdvjg3LVg7cjRlwMSXISmAywqfYwhWb/n7WI5JeNIghLJ3eWRCYZrElORZ5wRiS6eYwe+l
483mgjC2Iwgj1xh6eCb0m5d2xAzrV3TOrGenrC1S50X/KGaLahv3wFPlQaCi/ZFEOdzYhrbWoUDX
T3A3f4L6fTHwQ/ipMGKMCqWT3g1t/bjBp0SK6NvegNOLyrshptu7wEpgbd8cNH714k8MRzRQcark
/piOxBbg+9BnY+m142ojHubUtSoLMARkFUDsR+MwtEaj+50qgymPvMM1N1XFSBIcax+Clj7evKnf
wzJ6schxdEwBmsimfarp5AV5kcpmVo7u74fUeWeLozbrZqCzM389xLswR55UgGmjcNDz8JcQnhNF
v1lw+p8xf3Cz2iR3sdXE0/nF0PKPxptCQRA8ItMH/1wIKmkbqMwAaTnaW3pTVtDuLi74VB1jlM7Q
bgwzXz02Ji8pNZaGNlLIXT7bFHijt6GfHBN56xDpfxcdY6kPHy7TiyE5lwFzzSdn/+P8me2d4TQ7
e4vYlkScttz2gpsF2MMkSp0d67URF8Kre6AHMg/nzihLoaXQJidxq210RrlyrpilnFmn5Jn5bLQc
pFhuF/ZfrwumsZwxznWG23MAUouTUUu4OvOGEf+i81HebtFqyWJQ9bvvjVD5LAnZ3OFKIwt/ODap
TMbgiqeHNfn0T/YjzW4zYdpJVsjYEfxjRVoBfSuBKFjHJ4LrwHeNkt4qP35F7D2+/8coG2OVX7fw
7gH3HISHUjDl7TYXt4o2aryXI/8nwhfCdnI3rPHQ6xY+VH09aT1x0GudxddUrWoLH7X1dU1gP78E
Ae232o3kX6BGm5Y1u3jp4VZO8IMEFFH2TaBAHEFXkCFFix9iqQuuxvdvuMjmNZJTv/LPQO7lLCr7
pfGhwYXW/8fZN9wpP1bk5Tlvcz+vzrd3jgeelirdcSo8FLakdFNiEcQhzIsYTfgInEzooXfQbutS
VbIsXn7PDciGs3crh9nEYWJZU62Eznh2J+hyiZLmO6AOvR7BDI0CMt9QGgUy5THZvhdGaBPq8Jpe
y+4LM1isFz/lAx43VFizJeFIaTQKheAC3l7u3L1LQuxa5VuM3vQJ9WJXLZK+xLBuXnMCO4Q/nh4T
2zwbJz0OpROw+4pDCU2wWfMip2OS+urF0khDhMAEA8UNy2rt4tnosf7kWDff8jczbfYpqEmH7YFV
PVN5G5K+tBRCxKCCsMKPXB0TOY3/skxXpNR2VBawjsRvcUIDyljcAdc2Dk+gjrEwSFWCBU2VyStj
sDVqvc1F57Ms9AcW3noMzCLtg9r9Sng+AvKO9+aUA9ZlXrhZ7kZ2qGCHO3539qI5j+GMLb1UPzEq
QlBXFVWNSsVUo7ZWHWTAqsWQP6Yg6PZz1nMJVxiRT9GggJR1vft5iJCeXh7Edu5b0/f+FgsJBALi
qTR2ETuwho5nz7ILfEkcIp0TCBnpiA0gBVoR8RjXmmZI5Qn1WXuUiOoMuuwtkdM18v4spm3HVeMt
MTQhY5t9FquuoOiYKPPFGb5RvEew2cl8qrxjJfj7Xeve2vRGYO0Q+jkK1771c2OchZKwK4IMQ4ct
fXPobkmWZzLAgTbXorOcOGGIQU+TkNUbaXQDxztDwO/XppYNE5e7jmcoZO5lSalvXP9pYqdgLwEi
vwcEW5nZPdQ6txxzXqvb6HUH1I8rDo2+/lEhI0RMU3LElZbjVKQ50gwCP7nHB4MR8b1B+hiui6GS
Rg0N7n89oEQ1cYVzJi3ZV/FT1Ee5mk/KB8bHMNY2KnyEVG8PnMoVciiN0fmINdsQuYOnT+oU0zy7
qiL2ynAwup6JULXVjglNPnyNOmuH2CBCzeahkz+yjsoz2st3XYx+8rDU5A1AkgKpkJaHPvG+SOTc
gxQOP8nE5oDFJ6Q/8MhkuXR8W4/BlRIeHpk+XxRh77+F+SDRgQ3YaAOYDTc4NBIb5k56rS32lBMa
kJHXMwVYZ4Lqwk8hlZBvKW854t3Efe7ks+9sQsniMR900QoFL/35E9IQE6eHGVwcakEV8ff5GPaS
8rOwVveDwLSmyMZg1Te0PRjko1gUKHDX+q69qfbJB8hXmPEPjS2VTmMMx/S/4uBz9Y2axIsg1FKL
jzCjdAXW7Ekxq4FpI0P4beh15Dbfrjm0LXzA3Z/LeuVgd0ag84B+Cgm6GJJHx6LQ4FWRPYEfskUy
YCfCUEFG62wz4SxskKyJmp6DGzJIkZOoezECtd7MK1CzI6iX/YgkB+gvGpcW9uVMzvduNMRvXQY3
x3uB+r0gHPUNf1juvzZ2IOXv0aAgp97e7wqDX3hmYTYZCcgx7JxFL32AeB6G4N9lGmfPPX83iq4i
JkWDgSW6vY9fC87bpYLUR2cNTAYBuxuLWNy50d5GQnJFs/hMrsg2LH2gCCIzlXSIx8dZUtXCIbto
Bxy/kTYI63sNqhD2IdTSw7NEBBuUJpu4giLMDyAEQ/of7Zel3oHbCgdWlY35JFkaB27m9KBrcDl6
ioKU7B7LDLinmXIFeiSXUTURnVglBMofXtwo2Wen7Gqo7wC/NScP4uRV2f+YdsHEILMAdeRtSXgM
LapyHrSpT7myNdGVoEEHTMOFG7NyB/jI20WJhRrE53KnsGI0lNa1IgOrEr6mJzboyms4YMHvMIe/
Mosoh3MPSze2aP1c6gmbX8nTjehK490n6E1WOZwE0nunneRHj971e9ALwFM3BqnEihTLKjnW9UqQ
G83ZAgpJBGGYZ7vnhUYpTlfAWHn3dIBmViwUvcei3+sSdCkuzEUiZfULhRIvzx+APKt/QE37Y9Ir
ToVIomrdZCKofWnx/dBYlliCq+huK1Qha0mwAim1PjlupAZDCyqjJ/qVoXBgOfW2dXXAqNPApKDr
n4A24p4v5fiMi8wJwMYbw9GLdVYEpB/JReecSmvMH9jtGwRG9n/Io4q16xs126omP4KpGKYR6FMp
ueXw83rQbjbiSWaTlE2U9dlnnXshnedQwtQ8GW/eMfau/7Nr8coWr7YobsgMfhv2t59mDcM2cJk8
qWxtaDQmPBkdHttohrlWhpITjoaiQNxbIpmQ8Y8OjyJm7k/Pu6xIs2VW78xaPGIsQFbsLHdUvA/4
ZuUxXbD/aUhdbgz/4XgzARLJ01Trp6qZBVuBSv7S/wGgbcwz7u8foPOfxPH2YntNN6OWEGTCU3xW
71nZsd8d6WTQzuOwPNjRcqELuicYx0YIe6L2eHQYFUhLWnPH0MXLzi371Y9KhlCUKAhJ6rpk5rvD
NVt0zvzAF+b3AfmTgBLIHLv9SokRQknRBbTWTLbjWlEOBvGWD6ivNUpK+h/XloL7uwvHAr6/Mlyt
s4tO8K+sy08aRS8lrJ0Xgc2ekx0KleqeRbbyBc+2rIQ8+S6Z/i/6q4twsWb7FO5Su3/gDwnEa9jW
1vw7sB+5EoMvyEcEO9fXpA0maVDQefICOQdu4Wa29MY+4uf+cTPp5O8VMn4b/lxgQvi4m6754xFn
V3amC8jy6X5Df98vV+SUjTlalNBXOYMS9MSD4Gd1aIeXixDhiqbXipUWKrMVwQMBP6D3cSSwTB0s
SAtY7LeYX5tmf4hpWlJ06IGo556u/pl5vs92ImUXmpDLlnjOHfKR5DkdEwZHaOSCLiWuiiWyet++
YTRCdqOJvotTSIt/AxLFUNR3HErg2a4FCQ/jFBCmOIplQvu+kaqMlyrBYptQgHhSYMG+RRmzG0rA
ffkAgAHN/mHyiwPd7Qq/lPS3FOFKyP+3Z64yfaRYNzDW+4+/VGNPOSAllKLKqbi/5tR7jm8h3NRk
gPl8uf1+/D5IGNa0RngRySUCXFUsdWUseJfaymRhV7cDW/tT4syX1H2KcKyQiPEBFe3n8MVNTHXH
pgwETQpFEGeF3EtzvHU1tyvqOnHs5K/fDw+RUgRE/glHzkPRxR6k2ROKIK1911HA1nY3OI8QJbIL
8BLWnCiVZt55k2Mqixr3YuKxkOP2pLljLJn1DsPhf41hL+vO54Y5aCcT0IwCEIwtsB0go4ctl7O1
NaCmbjS/qdrbOgU94i4LE48rexidoMBsgfTzVD9bfFkgNMsVqbevz9l8GAtUSaE342Q+1Wfs95JQ
jamZ0doQ0/7b9N8a7lIOWkCE5HwXEiXfu/by3yBW/6AZThV4sIutTrKALwcp6tti4gVvCANnlogm
ef7UEtjEsX3xoNM7xqKd59GvAl7o8x60IpVgxuhaXqqESjXEg4RGDq9RqjyRxYbA9WSdY9QuZiZM
uTXIVWQuWzo0ARcLrvo4dtnuNKblNIBhZqfazaEo2kb/ShN9DK4gi9GsFlvCHiSmZ+1vsxkAfzmh
S/ATmbtnONtWlC9Mj/BvWbdbMKReSxySmOqLcbdSoShj4PunJGirhhdlia9G6n5LmfmWJfbTEN+f
j9rUilN02KxVuf/XZiUEeUIFY26zroSQDi4K7/ax/r2ommP6nMkxCS0dCBdqvaH6/jXO//TTXva5
DpP1zBcmQN6uFGamzKoxOI9G0WGiAko3b2Ndwxhf7aks6eJNqubOZZ9+IZBOzYz6jO5fUFExt2C3
vkOc3wwcVA6Vqme9l2oM+AutXX7VoUPtlA4HcqJmqlnBOHUCg80yzdyjxe/6vWFWzJT/hA3Rulx4
jeb0lTSzW2PoLuVF+DLSADepEswuT84nk8Kgjb6CM/HLsRDy9mHwpShluQCGj5bpHcCfucjuLZo9
x1+6ilHRj5ahKUbARuMGzdD5nOpSXwzIOCDWK9+SG237R0PmeJK21aV2Ct6ZE2JC7wpZQDcl7t4C
LqK4pF5dxf6SbIzHeivnMIzSPRfEgVZUJ3329PPKPni4asnWKHLAZzHQEpoVCYJzuO4iZj/ZDBvh
Qcoa8+Ul6oLfCw60/76hVqTzBX7kosHP2mG69e7sanqFv5o6dHYsbzroWnmgCuAIhgp6o0gwsaxf
+v8jOco+mprKyWYsFfEFhVp8XaRp9B3DzF0AYA6gtpiJnEqNzHJwrZLaNLT4T3jqZ9fL3emfFjFr
ckMSmxqXRvb3fGDEpFLR5bpFbu7Q+iysdoFy3LSEfHHZq5c5nI4506Ka7iM2VT/JVQm37GcGZh3T
hsMvj2KmzALsN32fqG5EyARQGgOzFXQYqkQttDxwa1jqHXhHCWcvO9AlafLvuEf82ccnYQB1EgGw
vTCPm+uDsYygSqeebv0AwTLvjbWy8Erz/giI6x062UkDF7i7wTc3JQRt/XXHFOzhTEUxjpiso1xi
ptX6jDM+whaTM/tiapCpoGknNPj433Z/K6N5W9TDbslkojRjLurw8/OdxBBWx3W1KDNBcTOFAWHe
Cm6zCYacX9IzkZG1J30+vCuMxnVE18pR2OFyPlSDVR+wtHdIIyyWV6KvyAPYV/fsEDGLcFkyVeRR
2098m60EUbpKGrx7ZAMSecGLs+8WakNfNQ5hPemop/UncBJ70JVu+9XpsA62Ofz8uIq50PipHD9f
S/ew6vRmHfZr67fMRCabikUR9FXONexGKlp0Zy6ozol0H34uuM0jsxr0Vr8XHdbzCQQX8JCG650Y
Lpehm/3LUz7PZIVj2b+k2xovpTHOrrslm8nlELJuRfqZhByURWYh75lAmtsXG5lWNOl2r0IHOSGO
Ud1cTHni70hBf8PCtHRE643kWzX80zthLf7yuC8k2FnJPtfx8VEtt4EDbEoi0sGsZ6Fu00hIxykj
sQcFD0zNmbaGmsnl8YPA3C5l44XSc5l7bUm84MxpchYrRz8MngYntO1c4at5hiERUV5Nii4ApYTW
1MFlvvPSmjKlqHhmz/O/7Ejym1egIxl/Wz9F3ejSYeXyTYQkvPcGx+YxqscDMkNuKBUaysQknqTT
N15gE5kBaEEbohwU5h3uPsyr173DlJfMoJ1RhDVlhbuAa4j9zWfKtz0ZE8cg6kgcRtlQDXeuJ3td
AqM9Tg/V3vCfA3nECDVWBSXIKCu6xYyUQu98sbxFlKczpMBW/FZWleoMrFx+SvIWV4w++bRqk3xy
DBC8C3XIorjTmcjEZFMHF1FPphYpRpAYR0zniexCS89Y8ESZCCikXRX9xpg7ltqfI2GjvUuEhKnI
bySiGkbghpiVMeYaeAmeMyLTSqZOe6tK5lzfjgCSDmoERepk1U8ZQCR9zvO6HtA4sWjU8eU6dwkg
PolnwI9aPcTSirHjxUrcN/zZomyC8qqaE0DNbBabmDHoGtoJxcZb/4d9l/9MyKBuyW7YOb5F7wWV
No+4CrK3qNUiGIQXJqBTE3IfibaSrdAKADvjP/qv1QJp2LixXwVS1a2tj67Q86eWyGocToxoG2aC
GGdqvSvZI9REiwEwCri/nKZaitTd7miIkusUTxSdfAeMqbOV3A+yeHKCLRDVNdiSTdcLmQeMxo2V
2LgckL6vfhHOOVLpV1oKV+fgIcmte1reViTMsw7XpWZnvWy9c/qeClMD+grKF8JwfhKvphv6Ws/v
ppiz5/0R9kuTwON+D/PZPGpUVGskThoEun3EtXNOBvA/8H4LDuVv9Q1BR4D9M55QXvzM0AXPzinw
34VHIFTWwraQGWe+be+hMlaT14zrGv/xRmA2je1O5QBm3n6anHEEgstQLFaS/Nuk4o/YSK1eZXK1
dDc7IoWIux3mDoM6i5oUqKpBgHqFxxC9Cw7vdxPRu6rowjU04YD0hoUkKIQCzchifUq7l0sScRNK
GOUyK8G2dXG4wwcYMEsCm3021Cni4vY161Uk3zq8TcJtz3sC3Wt7J95AY+pF0ThTJUSuKXalK5Rn
sYWIMtwettfI+XC8SKi4+eRlQT0wFjPt/G7JVwzTpZdz/PAWvrVbdjNOM3rOClUVwHyYDB3JTVUP
UV7P+RnZC5NUhwkWW+M7fImZLcE++21GhcpPUWDW8FxqKf7fQ8EAsjFs1b8QNVbzBUdN40Plbhd5
QMF2+osKAb1ByjfT42ZIFRMaC/u/hA4f0ipo/kPsIT1Jld6F7j1aMfSvPPc0H6QJoqy8EdG0O1X1
abgy4y0OZeDI0EJ1ltx3jbD5vnyvJ86c7ZSmTjYdITwqWBE1KW1p16JAejY9xvFTz3f82esdsaUF
zsRCYuGkf1qzEYJrOmyJfrPZbscCYyEpko8JOCnuAX6eUwUjueYniWd5EbVu04VsIJjOXmOl0VuY
TbD2qvkDtbvOVUuWwmLaN9++aGAQR5J6JjQxQPGZhQnsR2q3Obq3VK8quTLLRzBJPX0oKJ6YUh5w
/RAJ3HCQQDZLd2lnaFBpBP9wI1BuFckDkeI3OKv1hgRM7Jw6Im3PubGv3MRm/2NRuSbKhzekFhbr
D712UKcArta1yVJOavlGy/Oz/cTyb/NThD48ZlsaQTMoC/zH1anTv3inBnN8VO1xyeJN3jF1q0gY
8R8DBmsXLo3aIJSyiaNRewrcOrw4sroPi6duNZn2x4AA3U0rqzx3pzKdIZtawci2RLBi+Iaugam+
mDa5XF4MfoTd1nnIdBfxgQB0My0CQejbRnYwKql4Xx29CB14tO8q2qyUl1f6lA/cng0YMayXeUew
7rIba9gGzOkCe1uN8xA2NDNT3xkrinEUQ6hgY8JPMjog03r79xjvKkDgZUJN8KAl1hixzc+JjYkI
BbIfbIriU2cmzlsgtu1GE3DlBwybuk1uNf6lU4JEhRwwZ9YCPJ3Lyz8w1fE37n6ZoqYbYsLsTgLC
4C/fnsgDL6m/ZQExqiVHwjygutrfxKffwUnuIuYfKEOtR0dvekcXADU4JLvnPRKaJbVdZ7ZiBUYl
ALiGLYRY4/eq0xiC7KSYay98WU8hJ9RDcJH5ej/SshF5N334WEjnCcHpUyKapHNvB8JgVoUT3WU+
I9gq/JfyOMuTFQdxbdevckp3w+BDTCh+UZ6J0oTzKQ3Zmrics77/3IUNmE439/MSHZgIx+6t53WL
vXlzV+zMrkC1uL2tFFHModptLrY7p0EmeP5/w+xVmNxeIuor7/lMvbxVybkWz6opfUdsiuMEv6vM
gCS8G7oCcVblSlsIad/8Mcgmw/pS33cVijre2wx8gKWMuMjTnkWYdvdLtMKvzqrL1M/PEyEBrd5S
nC0TK1m7bwz6jFiJ2BFR9NaF/eOSKlhTtkeTwiwDdGcZ75oi1d3qVKOOsNnyYFf20LmdD4z4c9EY
0SBJf6Kzz89IvqYY50LGtPHQ/k7bIkQ/rHDrIU0WfzMHFQnH+HJhCljlKhxs7O93BITa74ohkvNN
YEA27pvqd/CSdFPJ7101XTEJWo8k/0c7oDqMOptEsZPg0PsSaZDSd0URwoWLN6hlUX0KLf38hLov
Po1Ud6GSpB85Ypd5eXN0n4rFmRg4P7oUpbC0yPxhwVWHKF8x9i0yWxhYxQIQmTZNWiNnh43J9VXc
sPkcfUG0X26VIEiSOnViOuIkmVeaUsjSJ3/6eYFh7mDRemWqnmU04qeAdihLTflY/csAY+pRRq3+
ECDoSx3lrPEHbgv6aN1SWtEBq0mlLFtUQzGrtIOe/jKazDuhO9wF7htDu9O34oX4Aok6hV09tzLB
XF3Z50FlTG7cXgXxz9IJAJvRpJG6+VdatVPpzb27lYnfIbvKWAQN9h5a7vQSqL9CVwoWD0Uu7Y5m
YtiEo8xYF5WgxI6vTF/TA/+4ifv26EXU9NV1vxxhc+N3LqWg3OL8aK2z4N8t2WdOtEebJx1rhlQZ
Q20PMaWa3sRChKFUAYhA1jhoT+y0DnukFarBHxHJfFaYbGlGp8Ygz96J3gSZO6jqPSz4nkwHv8E3
BIN53agH39ZL2vomqLHBfh6GjGjGTDP7Q+zhhzLoGFd1zBe1SFx7/hOidf99Q812ASQv3WgaVFHB
feYBT5Arqg1I4OrjjmhhKBkcNf7vnhCiqPaDwtVYeqGpfWDQelL/20HTf5Z+l9MtztYArTq9fvqJ
nCqov+wiDU0qKDxNwy4nycNiCzyGNtiKqmhJwcjzx4R7edqvFoGAC4P0WID+WxjTVsIxpqv3WFXc
tcvJRFkRsc/5BPZ3tXmUS1IxtZjuFa5QnG90/qmfCF97i4FA+ka5BKNOrvWRRe+P3/Xc3PD6PX+d
/WYRwOs8GgCQwOBxhQHLgvIMh8V6Lu5UswM/kkQz4pvgRYX/b/EFTjxoazT1lNJ6437T4FwnV4yC
mzEU4MZmko/ZqGvnBV7f1kCKE9zbrIlzYhiDvrkAxZYZIG76YEabwhqt4FHgfOjO60Akp0V9W5Et
apcyRO4VxcRNpARgcpUw6qLVqQMS5m+u7VOO9oYmB3qhYQCHbH5+l3iaAvqirH1j7ul+q+R+N+ub
ule2Keah94BYl7yZ/iK5OH8DmLBWZtT4PVY3Hss+7X8KTSU+x98f7CXUAkDN+tvKPK2rfViBK92x
WtumEOpdRK6FXfVPgvk2CzDFNrTheYGtIbC1MtBM7WqHUpkkmFecLllGolfM0c3oTj7qsgPyCnop
+J1E7FrvniPRsLO7P9/8Jc44qOgKmxAg3XiIdy2TnaJoBDElcwCn8CHerpJzIszRD6YkhkUaToQ6
japTHOyYDEBoMnyu8cgXvW1bGL7Yk62BbL1ik99cuW0DkuD8wKHiYH8hEhe5dH30gBMhjK0Fo2w6
PtDPXbUbzhXRtsYznkzfERfzu3K23qoULgz3YMjPCukbcOz596o3l4kmtGNvbji/jcQxO/EUSQ5T
jMl61uFXNwnba8Y0lKB3GLdtdx/ne8zZ05GPr7qLfEz08N3f2xcMCPm3bMnQdWwQTi5mWMQ1gURN
5wGK9BIqjbz2GO+cewcGUCXwwqSByvYggwlC6cv/VHlFQElz9gyT1njHcS5xjubVgaCy4RZyCrxg
LK9LPcBawFPF98jdGlcR6LuwMqPU2jvRAxnsKJQj/MgKEi4N0SZebdlT6iWRb79IasnipHaRGgZ3
gMT+6Rc7cpHkJLjGGHLGObx16EOOFL6v3rqsqja+u41HYgEqjBMKU6c58HdO2OnVYjNLQFL1WYpD
+acneP56JbzwmkJe/nqv0l/aNLmWWwpPbNjneOkkDgVyoT+W0TjWnMkjlrXddaS7A/E5sBf6be1h
oxecVjmbt7UvSSZ4BJAM1g6nARQTosh9k7rcWEuhSGJKcOmcz2ZFpfYYPiTW5KZZZmIP06Vy1j6Z
g9MvRlwIK4L4s7p6IfCBUkC7R+Ji2jGsDz14QM5rlgIk0vbTpYVrc1od8U9tnzLHitZxNqplMUqP
X9VTf2xAP0xP6Gs4+sgLdOk2yXqRpaoIAzPWlmXvLrVXxGGXHwLr+DOHqnYVLMHKx1rJe+Ty+tL0
cB58gG4bRPCZdFdXTKe5yXG1dOgub6M1SZ2hd46T3z1sAt6kKGMdnQMpW3NpbCXfTgNIXs390ZQ6
m5na3Nl4INMvNcrH6oxteWP6iOP74p0pAlgnQwI8aU2OrgFs8GijVOGLjn1r5DTyIyWJligQlgfs
efg/GL+xzOEgIkBsphQpcaZAlqnelYTHR0iJwulHD74mKn8Ho3O7QJYaBNcaCcZhgAfPSmkEIV/J
0QiGv4tqUjmezWwrvwT1ZjxZGHfinqzAEpUL9z9r7SXIw2x7aZaSURrMIYH8LhpTqlb6s63IiRlM
MsHrdzJuL8o6h8LqVsVYFTND22gXOJblswsZSm3JnEZPRHh2QCCTaonCYfdorecaNRJnuJRc27Hi
1bqVxO1II9tvkCRKuweJCkg8QlM9W6HVkGyo/xsgh8UQhX9blstshe2GKPcB7ot9GK3Y7Pk1fVLV
AAkc0cp5T3Fw7/8igty0pjKnBfvh5yKix0qNuEFJxFJWixYnZ4ljchDwsKc5x4uhwvPacg2fGcHa
4oJiWF5j7QBnFlLhKjy1G6RA5NRyPRvxiDdDLVW6J9z3j7TT/cam0LH0vZYZJz88T1QaNe4AAJo6
9P6MYJ+6iJiwIME6BvLPkx5yBWGeuoiyfYssDXWk1FJOOBlW4ItMyg2dNMdrxgopwcY/r4Kei4f1
FG8enSwybqt9nHeH+aouAldzlxvpl92RYu4WXzXKpqZn30da6gFYvmuhHfNuW2SrcW7GPamZMs5t
j4i4RtGmMbrb7eSwxNkd2vk6AfnbGyBok+TAQQ/9XeAGXrPZOpianuqXEUVjNhf8Me3xJONk+iqw
AIZOMROhMCHJQMVqgm9c0BBbIKnCQSrH3PNQlNKk4SLz5HQlkRbt0uSXZKYnAjstNO4pQoRZceWl
RB1s2W6Okytmros/tVCWKB2dPDP/U9dZ83G3sWS3jGqc5d1tztnnP3t8s67+UsTaZgUISSNwmBSP
LOocf4m22YXRW4NmH8I0s2Qd9r8F5P9Qj8fsLpIjg3VjvW5gtCQkaJD0koh2JJYdXwBwM4UKPC3a
6GyqLB3eHsGwqTTVIrnJ0DmSnNH9bWZiLB8frG5sbcmdWGKd13hPEuLHhm5zcYunwd6idAQgQF9O
eo3KTnWuolDKuAGe1HMUTG+5phs13mp9ApQWWAiKpYG/iXrfg9CaIugTTg907jJ3uQC9KgfXKkP7
v+BJYfS4g1OzetL9tZgE8ardh/5PsaFetnWtQrrmmFu4iM4oYUmZnYIhE/ee4y5c56UO7rhQWv3H
fmcBYrLSCBN8g2WodxJeaaadvCAoRuSN8X3aytL2+QA5jJRZxeP7e/3Tv1Jnxr4l2VSICHj3wjeB
UOGTuY//OdBXkEB+BIpVNrcjQrBH8LKTRkfH+7rQZBGYBT9gf8qsGl/glLUNIgPK+RDlnnimyqan
Ut/9tbuKt2SZvJs1rZp9JbpAIrT0Sgb9oJ8rQfVGeKL9iuSb2IBtyc9eWfCsZHOX1FqPumWfh+8P
zlZmoB72AZYyOnWgPlM+uANJkeuRsdt+ujW8vNnjaUJvw70ytDYQ30ZO9qZs2qEXmUxdS6zunocr
bdcKVlkgI01mmideyh6GQIr3nCInBEEV7p/G9USyqGIFm1mx1SZtec15qKyQT81oMr8KaLYSiB/o
KfJVV4l+frUaKsfP+qBpuAWmhaWcVxq6N2UCO2eg1ifVpPqKYbZA1OV6Z0KD2z6LrBOO04pOS2gE
dhY7q7JZNnCUV2DQqZcJ23BtbQPah+hu9FA0zuxcVs8nqnEVkw9feOwXs/Hn6YMowRMCHFOWIo1j
9UA2NQ9Hrcp6Kzf8JvKXBht6DjrBqz1ch/wyglV7umb7xk2d33pkykaXVYls3RY6mtxiEAmUyc19
YAFGX3E6+rkT/v+RNx6FKrntWgH6sI/t4F6FZJqerJT2lwruGhanO9E50Q1AoNKPcj4t6tXp74/d
3+5QmgjYWSPyMN0Nss+NWbDaCOEziyNYTmoxA3VbxEyUI/M435gUxwX0ICiZqzOiGGVKDHhVOH1X
sRc+o6cSm2Vj5xs+o9cf8IPBgFBGaT4PdwnF1OWh01ONxvlopnzCdPSudt/8gACug32V0vA5if1g
WlZ8JAy5q8h9sqeJfK1KRDeUgudOtPh8Q7IR9Gqgja2o0opLcT4Z9UqOAW206yy6yorHs7qWUouZ
l3fMWo8DC7OvAcpt086p6LZ5AdklKqtYHiyW6NUA2wezkl3Yu9SZ9hg/+Yvwu05tG9K2U6Iow+uu
uc4pfSQhK8XVncioKYFUXcr3OkyHD2gEeIFosUMHH6jj8Q3MsUNsTAdnwBu3A9A9N26lv+FyXlJP
ffGNdbxrERV4fLKNdPOmPKAiYPaTZ9QbZjKA4dF06nDaNxMA0OS8imCTbE+OkdWYCl0Y1gTquLX7
+Ivuz0oB22P/tjBoyooC2rox2NSl/Q++fp/DoPfaCkJl9njfLB67+v+hhYq0GDLcXWHSl64K4bHc
uziMaukfUeVNMvmeOfYTQHqU8skOo6+P6gc6aqUoFWcXb3u7niqfZL9Y9eX1VRYUOzPx2UTyy+Zc
2q/4TWtm1zhz4SkkV64UNe+EY6Lo2+dyLHBU6rDnLAYJcdTKfaTTJ/KygpTI+aFndPFji+F6EYUz
axBIWSMUWU0Zy66gEEx6CuxR7N4lUzriIKsDXcXnR/JkX+7jtdUZqU90PSTuIUy2TztjOI4trVi0
0qPgJoVuVIrmiETAoih1tpjPaS1e2VukvT4OUnrvUpWiU+FVP1/+zOS2gs2pQw6cvKVXz8b8ruiB
5xeB1SP0xuJEAfeTu6RMjD9so0K/TxMGkKaB6950toCVGQVFNMImWjdekJwudV9RxHhB9dj4VzqE
06m+3VuiJQzIsvF4D64cpqH3bm+K47iWhxiiwPG3iLJV5YSHxR/ifZeo5NR9TXT9ocvXgjJ+5/Gb
YpNGGaaC154FUPG7mb9swsRJx/8yvIZcLb4gcA2QY45t3ZXE3PURbojtOj7FFHhYntQZzBmRT72l
twtaD8iUFJQ+CrSe3qRZBN9gpjR1ao5J7ryQuTRnsITAZ+p0X3t7xp9STYWef9X/xkAakkWpc92g
Q/IOYNT3NHFnXGAeXXKV+hTUSc6yWQPm9BlzY3yojkgdFJj0vXZJ17ZF1UVsgT4ZIIUC25xDQZS4
zphxfgkVFP8Klg8Tw067NWItfOzym6vKOGi0QinSW+WPvCx4jTWuAUBbdKv+0Czn0MZdXSZOng5f
+cNQ5GfBKBt5Y3/LtqVxWkiIJqVld7FlnGQg2cjljjZTyzcUbCBWWZe/ShJ1DWGTLl34Tzb8gFYn
Pe7jgxbIawN3OKxpd7SNlNLbCfd7WJATVeWiZLffiv/hzctmZn0+t+jNEXeL5O29HaZMfzrAZ0q/
yFS5DdMQavmmxjmlGOIawyeb40LwTbsZyoiIgwlNBHba8L1IsX3PNTO1VQtK4oiLFYRy4fiEPIpO
Nl82M6joykMDAQ0i1utLIvqi6QmOSRe7k7fd4CMShg9Ugbah6HWSAnQEwAfjNqeZVmJ3fGOUTnsc
XUDATKlgyKaUpdFlHCNbhuOcIxCk6q7ug0CLm8x8Hs6OatYNsGQCvYR4C7cUVqO2dA93sPgOkq+Y
VK0CXAzr1yt+3my6rgrkN20YJxnkwlmFqhTQZMEpgQjORjGo6x6/X6nfT5WdK1m4wAf+Yq5S3Jc3
XMdRM1Edv/L44t4IOZxqEJMVfaimsOTFnU1ubufZEDXLZEiCZ1iCK3yi6iKHZg9+kE4xmRcYOHfw
KofzjjYvZfquDogoEXDpMm9nwjmCDbmyIuIB7Mlhcn6qro44g4zg6di78wtFooev6lmkNwBUEm7z
1wfGdj6aMJkqbu2r6+pWLWfb2Sf5jovgg/BVhxVcAXa+EPAolkfgbDCa7hyJcV30KNvsywWEW5rK
Nw3K3q1IYmXE/iWy1sONKhfmB+oRCOekbyey0Ju1/c9SjeQvxb1E9ERdtLyIi3UhHxKcS468dTyY
qAmyxIVdN8i8aNqckGmM34Xpfemua61ZiiPBy6VVd5SRvKCZoSfWI4eEAh+/6cCVsskVzETQH5Lb
b2j14ol398SmYDKEgq0tiTTbH8zXZWMQqrrGSg7nFrane3zmBmrdzFXPQ9aUlJrfkyFiJQFQ4Ku5
MQ5dopN92n9233b+PqwXL8zboxNxQKV0Fzexw0s2tbRIrT42xWxFeLVNu/etz0uSzFqzCvuqmkiJ
6ltnuisr4p+nTUORVJ5dfxSBdCxY+8jcjPuzzq6i5t+OKuiSqZfVgTOz62jM6wRTCQwm4mMj0XsN
4jbl+KHUfBmHUqmWQkd/rLxtGfXhfxIs1xrINefnMCYVD+wSjJoahqKhU3oS3D//jQYKb6Bn2nk3
6SMMNKUNjotivcOzrDjw7HBENw7wx5FeWqg4zPvKe3r7LkS4+9Cil6MAluTu/UJ7RuMHBpHy0lJv
L5t0IastVH2RruqWMiefJNnfkLh+d0+a+KHq0Ic4ybWdMbqZtR1nKKCUPoaScwr5b5feIzoGcV6J
MDRbiYUOl+JyHLYfvX4FfjhNAqa5BvQijjuix8OSJivv7BpgWgu6umxmYekRfflor7JB6nuIxRAa
GFZwHb4VXEwlPWaiOXCV0dBM8BTSexlfD7b+vts42LwKDjz6rKg4771DS9Sj+i+xs+5EfFp9aGdk
w7BglxFu5wzdBnkWl8tz45O0RFos/LFHvJRO2ahUrhEA9gR6XCmI4p6RD8KUVsHI3gMqwycJV1kM
HA5evm/sq1PN6RajTAy1xpNRmf8hFozXG3fEcbR6QpM3SmWhRm2AfjYzU0tOxF6hIUIzT8n27fZ1
/coCyyxGFQ7OPOQWfscfBPmMUigxzyp5v/l46VIXQM9znAfpa2medX2v5LConK3lATnn3wUO1sgJ
kmxu9Ntsig7dtj+KB7wzBn46v5YLuAi7e1jCqI2Q3NFwy1vD7dnCs4ixqT2Dk2zB+yrzBO9uMfsg
G1CJg3sPsNzZtVNYi+9iqOeK7a4wZGNeeuvb4/UQbTCuxsVocWga9iF7OUjpuEgAcFhkUvyWpCbW
p1axsXwBIO7Zmb5n8cR3+dFsDujlqsGfvtfmTwt+u+SfmTNrr61Nb4cczIAQi/W7B0AL3Mx+lQz2
no4i1D2OmpRAOQp4aR9w0IANAvMKG8VrJqze0VPTOf8twnlqtqf37kJpg7SKlDcq9Hu52oJFmSBp
yk41AmwV/ZQdGQY0Te4GN0zwxfLEschlb/qiKuf8iivAWMCLEjh1pvg1GMW34b+zr1OCHiEn/vbp
NIJbbN6gOqz8Atdx/ahf4aI6GYUzwSpHk+rQ8Fmb1+wWj+TUiRWWS4F7wfGa4fCrwhQ0ysjjtmCF
FfDxucBf/M3IsoQmlaihKKBCFwSuewU1jjQEC7KVOwWr+nS2Bu3ojLc9HKkAZOZTqLZMGBEhHn36
wL3lh2GOZF3Zj1rmHpu7ljwG0ufFCJhgAt86tsRALWoITGh+/VlZo/Tb/KqV/MAGIsFQt/Nytzg4
ugGo3hr02NO/SBuKeXhAHoJUtz+a16Gln8+cnano0xMNy8Vb9brV+Ug5j7gZos5k34F2v8WTi3oD
GZkA9WNdCH6zPWc1uXAKcEzHexlF8+wYQp+LEK9MIyuhdc4v1ODcNpCrH1CucccEKt9rYABFUFr1
kcUio0ItYjM1Gn6UYkRphhXlIuzw2QrVdikGgi/zoieRnOpvK2zbg+ahZS9DRqqpIbsmMdjCHw1W
Z2bpTWaSppmFJGkS5UtRbntSyL56NngPFkpudKTHMvv2aNtHRKHqdR92e/X4L36xjpviU3yOem4P
gji8kperSuUAWGSw8jL2ThDeZcIs634vb2BpOj8IsP0bAvb5JgRcFCTalkEqsmIsAn7OTucyzIhE
j3CAONXxaVW7/Rh2151qfzGTp6DoI27rk/CgOfxbcO0zQp53A/YRjrCRPrAKfL96RZYUt4eVu9XJ
Ey1x6KCbENeeuoGcwWfqEzhwzFl/hS4ZPo128lxilHAScamEKfVmGMIU0bVC1R+R9yEQcdMLQcp8
IPe28Up4UjKNj5/6bqWVC/gPONxKbcHU1osQK2lHZg3WjdFxVMDKt9I9HhppGwHPEgNHPDrSQSJ3
tzmymbDH4c7hEdZy6geYdickRSlpTqADv0WHajXY88eMH7zwNRprK9Fte2pfb6Xo7T9z2d0io7yG
hfW6w+q5rIoUxqfPv4IMfcn52kBMh21vTOvOfDlEBfW9bWcerMz9MVxAN+z9ynZWKg8fBGMbr2su
AukfpmsmgIPAiq4CprCyZboR73BkTgsajKmBKFXE4YqFrEGda2x5OV6Do9mU7t+GVAWtBqK+xQb1
kSZXrM9qR9GEl8QaDHDdK/qhk/cf78AE3mYS4dA1atmOjV4xkLQLRgNnGTh+u7c/poiJI7jcN+Dp
DRgkLbhsCWwtKlsc2n0BuDT4oqp3+BovLvmBdR5uFNMy5OvGTgsyMAOkU/Ay3tlhAqyezoRff6cR
Zl3bTgA84OXdNIFs3v86blndQo8vpgq4fQWHw0ecKOiUYRHGuRoTfBkthFT1JXONBmCWOk3JK+C3
wicuj6awE0jTDyNDsnIe9vi91m3aWVQQdql+aZ1eXjk+swbkvLphH+1jsK5YN8N+Sex9F0prECJ9
amJFp3Q5OMzq6lYQzpHTX7Ve8j4d1F/1yfmkmDw5ZpooWMBpNv25xoxz7ajzhJeFjBttYyLCnS/j
XJqOqfICw6y/m8S/81ZevmJuwouGxOO9wBEhHS9GUbwxV81CK5osAgRkw2OonwVzVcCybkhWa6Sa
Iny+6hXxW3PMNRTQ7T3177HGfbntfQy7Y78kGP2fOPGCFubbZKrvuqm1UEexcQ3SH8ptrrMWzrAa
9rRCPaROc9/Mq+u/pO/I8m3qN2cqHG3zR7zY6h38LgM/aF9SWtOZWDpYXBnbH7XK8+i80E3DhQTA
+0r1Ow0aEv3jPLHvhwzfN1kbjUTl8xiOJy2DPoMhshS54QsJVPnRlWWM/ef9JzieOODPyp7y++E5
pKA+6ID6KkLSJdxNqAlLu23OBaDw6S3r2CtU5TOoJ5RlMA0iHNCg40P2jhdEMR2nx+pRoiLMf5mi
sQkaWbh8XUKYNDGnlpvtgxPcB3zVQJYiJrGfjpfdHhATI73yVwpIyhIgK5rUxts8XQ9H8ZrfOPua
aMWYK/MiFALvF62+gXpw8sVIr4jWj39EEyetC9li4lVMnx19Rq0TQCaWlpK1xgfnuCYA1QHrF8fV
sPgmr01faGCjmPEydmrW8JW9cJWY+mYjCS76PZSRQK00kiFHr7HsE1+wbXSs0BmleMG/4oyXul82
vjosFjVRNDQo+5CApqC9047viQulf3AeoZw8ViwKBfY3HqdPyYePR+8AczC+J2dhrL007EMnI0NO
NWHwF3JtahNibbu443wUPl/86CvhejfZrMio61k/cXIAOkpk/0sg96bfnLqiV796e1RvrDIt5iOB
Q9+ZxJ25UyaOzy4sKXLToGh5+e7NYqDu5zaI3arACd75BZnHi/2WUps7B+n6FbHLq03E/LcqKFO3
Y8XWuXZBW0bRH4x/K4MuvBW5a9mKB3Ot4Cr5OpwhCUjZfDLp9oH54NnBC9GLMsh6ed/ISBiTE0Kc
bSPMtt8mi7bmfDfrX8SqRRlYnU9uINIfJAqWd77mN1RADOfuKz3KTDdQUt4LcHine5SZ+82n9StR
0zRhjNW3R0kC3OgRr7XUqPYMH+Rrpm/XQ2ZFeMSwJ9+9oHfYIskswlJ/njN7pzj+mC9QSKXUlUtx
bccIlXHC7N5DCsXEFhaoa+CppceAEOhIRB86ri1lHijIb6lTwCGsxIjtZ5axtChPf0jLDSWyQHwS
JRSyCmWVgbaWw2mDUG/P3gxBEQAMLlUV6TEbx+0MiK+ttm6vw+QC8glcKfA1eN7kWntXYYVsCMxk
L8zC/YAadLdHCpqnCmj1L587vNCtoQOiRXXinIMQS4KT6QA9vff7U2rlMN1p8rvriEef5Va4iv5I
+YUIqWh9zMS+GVFNG7I4dGBQHEgwwCfzTVK9Xxzje8IrmW1FnMwaFy7jEmU+7PvZ3muv7+ss0Rkg
t5rOKtiN23WIus6dDl08mGPRHznTIy2pTi2Ha9AXjGnD11aju7BMIxDp0731WH+nUzSx4oxBu+sT
ftVSa5shFIy8YOfsCQgFUL6MkZVnBTgsNKe9immGvM5udd1kWbN2ZYXA9Fg6VubWsPjoxStTeWlt
mZ6jnUFfDd9LeaUr/gdBUCCbGFyXuSRwbbR4mXN7TE3Dt7Ywf67WVZvVwaLfDxuYHZto3rFzU/Kr
/5lqrcCp6T7nNHnuc9hvX4jIQx/faoyYHAJ3yI2JV7ZUJrTaw00UoCAifXtsgjE82Zakeru1a/Vt
6wk1Jhb0iV8PZI6liJsC2qx+vEYmTz/O7zAEIKO1uaO/Lv1ZR0w6I0Kpc08POc8myBj7RPt6sEcG
0rCrsAWCODxAEXdQVroop82x7bfxRihItj1PPwaEpZqBKmfF3W8j729xo5Eh4XTzedWRxEDx+EzO
8X54mbxO5e5vn7qv1F7N844SFVBBBI0e0y1899kd+E3FT4EJC/IMMqELBvyNo+n0IAIjh5Vxvrm4
E9hsF34+AWguRlLL7O9OGtaKwZkjukEHgnPxKoV8P62EPgsDYnBfiWfe4XZMtkgOxftquRPDvqwF
Nq1iStBrSCPtlR6s+w49FfDKG8Zv747kEKcCbKaeCE322uwXjyV9m1N4lpNtg4bjTr8Ed/29GIaB
dX5bmrBu0YVWyb25s0FAt2QbfvouxieTnCjA4XZtMv0zeyduVAfHQDnaa57CXFUthiMS1PVLgrLV
ZOmpWw70b8PJggtUKKvjNFTDN+Evmz+gBqa2cz1zqzXVFQClh/grixlLP/nAVwhhZjQRmpfyBvG7
B3//AeUINCY6PCPWwMkjny65TsefzAEZfOtSTu2B0Q/sekZqA6TJspvVYqdnZ7Kzs5vs+31UYJgu
2MgJxd5j3trUvZJyR9pymKZV1PvIY19dkK6EI2QkkVQztJPuQeG0N4qlQYoqzLFY89spqkxA+uAZ
BIZGREnFHmfdpuHET5jiznaDHjSGjnN5Dw1kjoHp8v7lIUQEMlNzrxPQ9RnXD6YqKbSjEXcFE2Hf
KT7+KcdJgjCvFyiRKRDQrVpCuK6HMTxIdaL05mizXPJFOZgSL5z3lmmNODHGRAIBHW6UwQBQGmdu
jLCSqdtmjad8cFrMnh5laPPCPRJUG8DC+Ke/oWaiFaGreAEh/txZznXKpfUsWQvJx0UODMl6401v
rFiOXamIikdW9dUzZFm0SHuwcgvlXAu+8yffWjH29UAPwcuwneh+zbE4F8xrWDvhauzK6fQapJlw
t7zwUYEssNbx2c1mv/kEJMzB7GwOrlhjqfqYqtRZ33rjLBCLMZCP0ZqJ+TZ4BJZbAwgoSy9Q7bOp
Va55Pz5uRQubvMb/scLVCNslX2/4cdGXDdnGFDlx2Eop9vcNIDxgcz38wdTrdoUTgYvtmj1xflBt
/gHcV2gusQCWqMUPY5pvt0lkHHzo3h/l4kn2rCq0vqxSjrFNjlmRrEPV5eF4mzDME08v/EWi84qQ
O+j0v4SRtzGoQR0I7k8jT7aMNVh9dGayVG4leXacfgeZrwLxRNDVw/B2L2O1GGrAmpT1lP74QTnO
ZtW1pY0JMeqPq+F0c0dbb+N0es9xBRfvq8pg+Jc3dtdJRJpF0YDLVCsBs+okTQgi1EwPVyAWDrrg
Q5Ofmblp+Zk79Rdqm7xAx7n4unCCGmx0eQLqg26llCOYAs8iWlPRKWtkimoGww0p7MgJhAeq066S
niqpxXtsgrEbZW7fLTky7T5SF9/RQEZoHyI6KPZa8od95iST1M5snECpWVukg1P8toS/o/sgNE2U
I78x8nmTWFFGRkqKKKW4J1ewGUX4xycGEEXclNNX8FE9pnrByjGah0szq3NdZX1weXBFNUSVdKtH
uempGO7RF+1Bal2yMjkbpPYgTGGZzoqhyYXWU+vw76m2l5GISeDLwliNw6/l3OQDDFWX6N3A2l7w
r4A2GBZdwyZ9tDjsHmV8jPAYnQPj1hwHVzanc1G2d0j7ln96JP7dvmqLiSguUnOWeOG/CJnm0iHo
mgNNZ4IcvJzVoWl/BpMFPob2kNmY5OWbuTW9mf/qRDVJ8W85VbcoDLKdI7+x66KsAoZnkgm9FrYr
dGxrybcaep6LpDzQBQl5BMW+tORqavtlsr6l3/aseB3K0lAi6SwmVyBSZhld5MA4FNaZ41WLFPEL
C/wp3YJnYdCU1sH87Z2LGaRNPxkWoVVfGS3FcGi7zLdq4go+dWRuOkTz+ZIcngcxNRTjGQ6Qpp1M
yDepizqw5mzeTl5VpIcJ9L5trwJqmmmvfVLxCxf3uiItXav/2zHkb8JMTXxYJACJH9OYV1ZQ0JAi
UHHLRxrU8E0ImJoLzNlvIpqVStsfKMy8SLNqj9xhqOYHwloRTv5k5ny/KXtC0ZfPc5VMRM1jITkz
adllMRKkqOQduTeOcDHZN6AcyN8BWfc0E/BfNTOcXa1MEpMgyOXWGQ+Afl6FpnQwbqxXnB+S7VE3
TDxnH4/fPNQzKJ8bwpTVcJU0LZlcGyuPys7p2LjsuF7ZNFif+ZvZpCEKTrf5d2YayWipXFdGo0lm
X+mEO6f/9X5kX3pycfWp/06+iBMrMf+a0FMpks4UgzSAwKDejuEHHgetniGNLNob5zOe3GxkvsEX
oN63PxoXGls8pi1Cczx3YibPisZ3Nodyi1bldCPVatIiQ0I2GhbDBvdOPLNv/D2u6dea1GB8t+Ka
w0HNuOeGOL1EUJ/xw4EfhuDiXIuNKPnu1L/h5qR6kzc3yghtpYQuwg+CGSM4GzccJISVc1k3cupz
sikjXof3NcaZFyzs0mzOc7SWHR5rM2GDGQEjOayaM+ANXRmDEKf8HpCE/Oq0YaBtvuXF1sPPpvHJ
e0oqzWmW0d41mCZ21cM+thvyZ6k0xaPWrIKghy6wdELhJpP57ANi3SZTwHjVFmpwQfk7xXJrJsHJ
+2OJUgVJFbTyWEqz5oHi80acV4bXF8AUMZraaUOokHp8sNVKgdgrdGhogiEGEuHXi7TrEgTNKGte
azPtx+bbJzO4ZDEWtJ/ux8Qx7iVaaRgMz/e6d+WTxt243x+2XvR4hfx5hz/8wQNGRrQ5/5wEhJ+H
mdxWD/NsybdLNdlwr6QO7qJalKoXTZfrPibIlPQVBT3Wlqk8kdX+aanGvW6kmCJqj/gfGtOED2EC
RyBxT4pJUcAojuQnbB0VtC5b/iVHbiO62+q8nmjt99K+TBaCKN9bAY8Y3np88GhLHt4FmQBLDvnb
dzEEQsZ7YQs8Hu7d9jeZhFgp1D6QaTu26SdcImmjSf3I0mX4xvxGA20Q6DFtc2H+Rr/2cC1vNFDH
/2jmTRDoIOsfIb2Gm3/1t69oF2zctbLzjza6ATtxtPaipdntiICueQd6sxQLCnnDYE7XqXRNSI9T
7FEREL3k+rbEthupyQUbEN3zyYmWx5qK0DsB/Hztg8DrkZB1e+nKqE9ywB85CYLCS++wHAi0hx8v
AJYJ6hGoV0LVUHNaA+AjM0Ot2MmFs8Ut4Cm2IH+sd87XmV5fOiwbSQOGcp4SdPpl1kIhTWbn5/Tm
2bCEVygWe6uBo757Zia/SCQwYdXuSW9EKV8u4DJOmFa/aqSxA52q5byYUhyVnOkZF2xkUzR3pAhV
rSCFQMGDHggvSoWRRdJZwNFYLGOXRXQWvG+cuIGhCshJqL+EOvnL/+IclhY0EBq9u4LVv80o3nt+
OEqxnSN7ZJ0MS3NocCpryG2GPND/ODm5c7Xs+DwY8deX0vLwzNuEyhgogQqa+K5giFMIUc//CRz6
Pey+XUfkrLJZCeaqPoLYcBAm7zCPfji4DBdVIuT2Rui2Mdw9XVMOALvEVquHg7L2ROu9Pq48UMAS
8eQ39vur76dg5CfRBYpq89L23pmW1scJX1uJRsTGrjE9LCz0rXiJVqPHZi+WuVKZqnbk1LWQ8S2n
sxMGIsTMz/UHf0Ns1a/pyI/OL5rbzVI6k7iAfWfk2guDwASYlM2QLfpHvnEbq66T7O+wWJXyCcqQ
GKnEGI6xy/Qmp/XVNBeCvAaRRKWUe5IodBVD2PVaxtgxxFafFLrXhwDcfCwZy3yyh/hvl5SRQExN
2B+qc06ARDlU078wWXTU/3cE2/AKLJ/pHu8Mc7MgWExA+m7iCcmXWJo8flBn+fPljZTcibQmZhvY
KQS23xEZ4iildIevQqStRCgECcxhIUW4t5hkqtI1mJejMM0m0GQgMaNcHTOJOqPqOz6jwAzw18I6
+2jEUEHVFSqjNQzbDYa3sPCM5mKEdpIeFnJHONPtnG9jWl0WzNwoLHuBvQgDhdPCs0yjUQDcKGyN
s+xgBCBcVvhiNK9O5A+vIvwrGl8umeESGYEI7ffb/qrgnDvWyyVwbz/UmSJO5j5YgOgSE+K6B1oO
iabiiJNUrszJyzmqsz8CetxBdYvq+YRnF/deoUtpZW0vEnGCkDnoiDvA4vve9e+61e7ZEERvDKcW
2PVTNxL4zYyB6eeskzLkOQhShKLYAj36hwA/OEceFxtmkzrsJgtfRpGL0VfwrPi60bb7NuTTvEws
Ky6Sdrg/YO51RjIg8/SXCG4n3NBcTuMamSgpHxs1jWqHiRy2C0zaSMkwQMRQb6nIgWB/7unBJKcn
1JshOudDu0cfGkzazF66tiISa3421PbxgOOlxZR3cITFkexAH7VpvdfoI0g/+ziYPFf51ApENh1z
lsU/r4+x44bNSZ79NNSkXduoBzjjZvQZpTIfOPQ5e9/RmFiqJVN4a0QQlFQBdvnSEfPkQiTaxTOg
fNFX3PMEPKtLYoWJaTeGTxA4w+Sn+7p9qyIRFkAZVSW8hjjBkF8dhuKnWZMlgGwR/1hC0DzsXPim
nJA9PCAPGoJTIY8HBpAkIWdSx8xYQjxQ/eFws8bQvuSwQeiMJik6tM1tMgIYGWB1+21Rpxu/W7zh
5ef/dV4tciBwvPOIRbIOJLBWviro0VkWEONyQCE+HMKRTnsje8XzEOwqAQQzNzLru/X+nztt+JKg
eHCJ4J4awx465tqS2hnwCdhnlQ2EDOmV/21Xwk6SXVddU/2KXAYea0IIPInz+8l32oUcLPWn3tbK
S8588aRXosGpTygZzRW0hctWnrnOsk84Hx/otiBB7IeSZrY6jwYZZ4XOSoOMLnlXRIJWfEkjua/m
NkOYDWTXBRZ+xi/vVhp2IiY3fi2GjVI4j07RtRa7unrJEwtfd+TZmE4x0XYxc9dy9/I39u7uCcpX
mSxxmGU2TyvjlUdqc44OKHojC/4jtqIbdkeNGcPd4LTHCZNXbKDqTbWcLLvPVqnDBfDJZ5OdK9kX
/iPKAR3ygZ/fmYS8oxTG6dh6FQmpbJVVz474IN+leLtxY3V0M7d9oGxvIacYuscO2EJyxdtrCYaP
Mx9DzNSYuFiG+Ow/U73txcxr8/e/02Fa0Lp+DJxSel+aZa+g8sm0Koo14Bn7Jrpb6XsFAb7aq29y
3niMjHlOKWG+T8/B3AtvkUfaQGD0I+K7+gyXvGV2M8GuFpSs4ELEDCGXQTuXH62cyaS9IX1hkQQ7
KQgLcO3Y5JV82tc1z3oX2HFlYSISBlqCKlN6HJSvQY9kEaeceAl5SvxwusN7lJXMU5e0I51RTrNT
OTiRtMhNjT3dGJ/WWGN9T8LVsYZm4NII2B+OEc04iqmrMOgO0rG0ggN9ngUJo2YYDOUZEblzAFQE
WL12dTNnUwD864Dys6P2s6RzdcEFu/eewOdCQS4gD8vwx6K623aJZ9DmVRHhZlTftecizulfUOX4
k/2ehWoAskBIhrNilZE0/bpjhf7LQ1W9SUWwjvB7QBDlsuPYDo0md3qTWkKXEdfie06HsIS2Seyr
UHpLSor0GDX3mA7vsZksVVehQYv4UPpIUhyrJFc5VOJdmrVPQVi6wAVF5EF1GdKmTO+ynsdmaY0O
qebZtdy1MtaIxU+ce96SmKTTbh9ghYVbFUdYOOExf5ZVdhQPMyUi3nBLVK2XnWrOEyrVryZ3U4w1
YquYz45OV5U+QItZ5vBdPY2Rvq0qbkl7LhRNaX3w++lRp/TqcYyuTxY2UbcJI1I62uLxcfSosGp2
RYBdekcII9qbco0mJNB4QiiGVb0DLD815LzpdhdY3Zp2AULpDXduvb/W9ve/gBV81D2gp9fXcigh
y04rxysBprnpN6TnjiIs4hei6js5k7EhbJEea9jQ2d8sAJmvHwgOsgTyutVBUAPVkdUBzPoLHCQc
DdbGaL1xHgURn7oO/RAad3IKvapFwKCJdPioOBAZvxRDGIWy4ckwrm0zU1rYoh3QlCmZnIR64mue
ZwZBlpjlCN8VHMF+wHiryrlsaVDNVMPnmMQ2UuCIg2LLS+fJw3x9TwwjXW1+2aCvAuErRNsBbriO
Ql5NNf1sUpKpu257QferEn1Ae4UO4Bs3Lw2gZSAa32NSm3yEN4B1FCRKZzduuNLBxHoAky/iTNLc
AEm9cSS5S8fV3MpCudyVi7kalCMmQWHv2R4od+t1OI1NfFJP4a5O2QSG9Ym1ZqZtvitZnm0XQfPm
4tyu8aHdBheUVJSe8rtrDAigSj8PMwgBQLCd7a7qQbD+w5i+Fu/wD2AjaNBbyMDRvARuJ6hMJrr4
qDrMSUmIePg02NPajWXfvlZbynUne5EjBZY6J3CQ2y1PMAWZgcMiLx+T6ByY7plfcXbxYGpjRDYa
/HOq2S6kxx7qX1FgjcvYe281RBCds2pMWY16Z4YnJ6XlsBdiE75zcoCCXAeBeYTRflS9cS2h6bl/
O+i9cP6vW97iCcgnsWXMP3RTQfsRFxW93Oh5+EbfkldWnASR5iakdNjN7ZTa/9N4WmmAoznY64ei
I4ZLmWt96o7Stgt5EyxtZjpRF0qCwB/JWVynfz0zW0QNTQ8apsrgVfJLjFUHohWv9qIJxNewxMG1
rSFrlgq4V/qC2j14pLVglAKWkEm+i3dR6nCWNcj8ofDbV7yuWUsAYBDb/ttbroPy9PV3b/y57m+I
zx6tTTC6UkLvBV7MAOihHBpxU+Ij4aaNFMwBSBZrH3HmsReWr/QlJc/MrqK8/7EpOlatrHNk0HlH
m+zp54LF4/X2dyymrZWQ/HeRalNjdIPwPyTJFbXD7eSWUhFt70IHLjrW3cZofDkaLtJBKYqT7Abe
uIwkoma/Jh8/xQoTWpbq1xQU81+sXsH/h5doe1POv6B2/zQY8gVlxEy/UHAxO7yB5gPrQJE9Fzxl
jLf82iWFcco7B/JcLP81EJcOmFP76O12k9GkEkusH999fAr4ooVtFuU+5Jyg+Pk7MLphgLpj8a4Y
dzibNApHkCZAutn/ngonr9HCTWVFbx9NaUuur7LGatZkMbKqy434btlCHUSUP/VYN8AtzQFCip+R
UtPX69bGQOBKfHGu3ZVR9b5dnpMW8EKXGskDVCa5bhDqohasGxRAQX/KjmeNX6nblVckNtpefMKd
BEfLdrUXy3bW0SBYNdyA1p6Qo2uIICpJBI0QUpt+PSAge1U8AIUUTme4mOcDwSrReBPe+rDgFNE5
QcwBkE4T0wEdPGRhUhg4g73/JGMf5PmK5t52QtB6oPoJOir77g7jvITq+PYTBuhlz9IDqILgd4EP
yogJl0r6pDDqDLfHj32AmXUUe9wV0dY4A+Ve5IMEAi35qxTDoG229oI7eGZw0h5AcjYUYRHTSR4x
L3+ECbx8rOn1ZtFts1Ce2/ELdQz5a3GGN0PPNwt7uS7GnU0/uK6cTnApcN8XnbbSRzKgk3quOBBg
W0xsBgfVULYVtG0+pyI0QTVoTJ0EyOIDh9rpvxTr8V4zK0l5zPqBKLKsmIcqyy9ealhGu0JIIOI+
h0jCVB86HIzLZ4gMPkP5pJjccRSikW+nMrYJuUUNXfsm2AekWTZexOisU4HMICrbe2SiCZJyEzDo
etpM3rSuhpomodyGeCPTNyGdSeEc69FQgUdva3TtB/oqxv165bBj1vhkj2r3MBhKztuSnkxjM6pP
gJ1//E5Yg1x/NfMZAIHVEk4/pvd0ZnSPCfEpTxTeztQkruM8o4Gi3y894U2oXFdNEOYjaiLuxgwn
0eLXVi2eM6n1rYDj3fXqsE748x1zcEfb40aiS0ZOU/JOoT4tgS+S8u4DqJmI9pu92QismmwMR/q1
dpbqLTy3BYpJ6Vz0+/FyM0LYvb6jnZskkzzXGd9Ep9bMn1YfmRfKZw38w0RTUDdYmXuS7fgNGh86
s/mj6t/0HYcFG31fSXnyvTQhXAtSaBIBPRZcexEc1lsotngaiB3JrPC8UWspRTRJtq6SZz3xrL+V
6R8mCBJEAMW34Tg0PTDSDPqJyolex5bZbxiX0fsF2YfXokv4SUd0Zp4gtjchRJhQKJ1/huOJWxoL
rc8kBXAFGu1DF2LZWOAqoWeF/D5MZiTXLFk76hxyAE7bew1tslzfDYWBkyO5i8Wj2lQV69X2bWCn
z2KJSAh3ZqXPyb2ooRomHkhEfH46YahYu8f9fk7qi2I8cuZU2OOMCroM0eNnIth7Fg4TVuMBXYBw
qPNwBn5pP1WcdSsiKsgU7ry9DevJSL6LvcnI/CqjYVbLaP/5pXyjHXTELNqwBHLcbaDVYz0cWRb1
8+QcAqZtwnTiOS44lYaGl+uR4SM0NEvqfdI3vla60mS1qvgt4Oy6HmlH2ScNUl6ah/5e845Zdj+v
GYCw7T6EGtQ8CQBCDHIK4G8lzsZlVHzMTCNzw/f1oUFEtEB+WN6i2Jsg+HatjTu4Kp0td1/O28TN
g2fOOwrahCnoGFTPMoB59Wuzpususv0eNstgTzAhVGqR5mXKQeltY1a4Y06CC8ydvyuphwC9A+Ak
0n3paojKBQ3O6v1XiV/U+ppeHOmi2WKjg02eG6gM+RCT+50qqGi7ndINJtij/LbOVz2fe+OdiXwZ
dTYOXjAX/JmBLaDwFd7vrj7gadE2zlGYH5289hS7pHITyAt/BibsYNiK5Xc23XMd1eTHUAZqbW3Q
M4t0Y66z1HrA1q89P/CtrX2e3GWcATVIejHjj7bYKFeKzubVAuwpBgG2CK1Dku4wOAtKPVpcW6Tl
vb6S3Y4uo/PUdDL6LiGf4o5IvxEP0H4hQ1ROVn7nttecXqDCXyybRc9vodlXu0lWZxd6Dbd9uqC1
xcEBYWGYXkNiezyfwQXB/mgkIsJOv5XEUxj942nPDiV2x1HadMLOdQ2drVtIRTMKGtKwg3X5AYM7
CI+VZ9rpT0TrZIO5RD+v7y/oOu0Uo03+E9MvKbmgv7wNO1yqE5nF3TwZO2QoigL1nUoFU+W4idGn
kV1EnfJyka+xYTSrZyUMfj97CUvkXWsG2CzVP24g9oyrJUukzmK5kpm57Ivzi424Yh6mr/RvKQpe
a8rn0LRVhd01PcZ6JZ600E4rVsL2bQD48Rkf6WzqzmxbPHuolBATJKkIuNC2h/kN+GfgXc57aMJJ
DlnftkuYHSTzlR3LyFiWHGcFUuvQWGgemU2V9S5LJq1iLDMVVYCA4wBLyR5Xv2Xn6ruueKNisrej
OJRrAIpweeurzqCqASru6K2kP5WhPJnmCkCfhEZl2gsDJGOmvvYECnDRU+2WlX44xovAaCOmrkd3
h/zyxRIo4/fTk/coTgzwslb4o6Utt3nFTAJQYjQIae/YpkYOKYw1VRZ5fVWjbR/GUj+kh6uztxqs
73QGMTGEpMDZGO0IpZhNrq6x7py70t3RsUknmG6WvgeMUKfSTAITBNfrEu//dPDT0LNO796BBKcE
NgBj6azf1nWRJhxVBqTiL/C38ptVDCqp1VTmX0U+PyWbTQhY6X6b/G739Vr5UGin1cvUS/W/mQmZ
ZHEIBKapAeL1CgKheJ/nMkVfamxvR4sSy9G6R+hjBA9fmnbdp1UxahoJ3k7Q/3KCElwjwbpqa8Ww
kwce4Jguw4mLmUUy69AIrdRKdURKMUqJx+Lm5rD/f9B+JYUMWrLG76OOIEMmMwP5DSm83BPhG/Mx
eRY30IofdmC7cQb6FHxC1HR0WqJKM9HCIjs9YopsC6XUm8zrLJ5vLuT8bLjSN1VPTseZ8EQXIxdF
kTBNkOiWZCT1yktsUta17Zr6QqbJ0smfHYPttIv1c/mj40UWO7BIW6H32G+G/d1XArtPM02s1NEl
SDloE0+zq866/RaDSLT45wMnwxZY1E7jXBr8tiUiJd8RATwh1NphfySV5vzmzRLQ9UuBFHUI75eW
Wrpsmk9RROUBDcYJUbQkk9wyrt92s3ipkNuZiyOXiZyieX3/uW7EKJ4tH2NAK6DhS2Hqvk4hhaY5
91JCW4zWQjsLGQtQ/Ai5kn0yaT6gbioLiNN2XESJ0gar4TKIoi8vV4FedGsQzZf9DcN2sipuSsMT
Q/EE39TLlAT4rpAZjPetdZEqFsspT6JFQZj+O2vIqeB5eE2kqtAuFU+ldd5phG1Jcc9HAXcYT+nx
MMpd9ievL9ILS6y4BTn8UwX59B6RE4BCmyG9zzSBnIRMJdorK84rZ60E4hOVuJmqHAAAeIXUMODY
B9CcHtjum9du4MaTp+JuM3d9ro1QTy4RN9QFb7TWbN8JanXjaItxp5Ech9ql18JHSj5Z0lkgOjTY
iZib4p7kozTwDW9A+73tpWQEbzoebg6mF/B5CxiY+DHbQ9GgOOWQyp9nDArGjH+w+S+5dHSxvcbH
piRUVEuuS0YZFrdgsiD+QxiLS8zbeLyvsanZdhh24b84ft/M6lqDFLjMGA+dAO5rwMta5nMJ3kdP
p8QXyk3xxFeXh2NK9WNiGo4ZSv4uOT8nkbYMcSvW3bb+dSkpZEshvu+gK2zNKUd/lKdOEUL08vmw
Iq9LbK41vWxZGsETHk/7jFLXJvCJ3jda2LGJZGH8lviGwdw8U2DAjX0F/ag2RR2WCgN3lyk2NG4w
/rXZWO9JHjH8T2abMSNdiBH6kvDRgo/pSKE/LipTfVqOKj83DkqQa5D+cbr9CtafylKO4bxZ7j4e
to5nk8Znc5B+gUPHzdT3EcZ1gMklLgBDt2jcI5G3n7XocCnN3FWGMJhoIyaX7cYg0Hi0+3zDfE8E
mcRaI4ghYPeOGOrgv9AGXng1707x06flrzrOiDAWk6byBYoOc7mBym+oir6qhHla7x2NU86OZoDG
cJzliQiELj7O9uDOOoXyAsRO38HXtmKvMKs7BjQCl2WqgvuM+NydJ9c0XCfUl5/z6bLJ+772HiIm
6nbU3geSlsReaZTRGZpVCZb98oKvaQJlj5B7gofIryJ9t7uIBqa5tVgxbYZD/RMf6iHBwV9ktceM
i8t6cKcTOygg2ZiuQShDhlCG0Skmp1wOjjsWTATu76tHCIK1DWxf8GDG93t45sxv5j7a/Ihkju0s
AO17EIDmRO47CoAl68OSGcSQcwUbEWTjj+lIgD8BPtyE7pDfOSm9ZOgUw3yVb51a7ClmL+x1GlHQ
KFGZbC4gWXFaLPM2UbluEejzlrRbUCduEXVSgohdcVCusG5VAIbtSvl221xpaq11uJxkCUlKFx6j
/UgKpxB9fdx255eknvCFd+lLQentuTkwLDvgnjwfJETHfXLUckwBteM5LWS7JLw8WdB+3VgvsY77
lO6ZkvJ9eoE+Pl+FptwH/Z8o/VGHtoeJNYOAYRipX677LSfslZD4Qi8xeC4B7G1LrW//uLrsFSdX
Y2JjqQUr2vgGcFFRbWPA/sPlsxGbsHl+kpMvpcxIITIK0l3jncVTSYsNBxxD1aI7j7WgluFAqMEU
P0fFtc4g5MdpwiVFalFx5u7L8b7N7qaG9SqszDA/GRHKHLnmB/RGQ5V628m/hfe82crDZomokvEs
3iDXa8Vixl4Q9CpkFKCCsOZNaE2E1kDvVdxbur71xbAHdnUUEC00l/rl8KfsG+I/Z5IkqiwvKqkl
BaWjYyBJm8lAjazflJpzCy9usBODV3XSU9EahWZEZoFsZnLqJlsqBa9AxCHhLtoGjihEGeeElr+h
6lk2yp06juQoI8/NXJUFalKNBdL8FuuLE656iQMJxgyqgRZA5AqOuNMRhIiqELdWJ1EEzNiPaDe8
GZLT9QZmQ0693F3VrrExvw3op9dJoloSqU8WZhbqO/Rcjb2tc16fUf+QL4f9FrQvL0zey9NE0bAP
m/ZJnH8Tumf+5K1bbVe9J6Qobt8DtQ+U4X1Y+tR64YkdMlnMWTSkjorQMK63e/uCngWyQWK2Wot4
daV41je/fI5NWkJCD0caZ4jJ85ZQMLyyViwBCLgGkOn1Rlk2vYP+72xAWdfPWOq4AbRT0ibKBtFT
B65Eov9enMsr6+IuKLtb8Suy8YiIL2IFWVZXNkvMJ06sFeNGzjnfqwoCk3orEjqpTe9Tua+zGh8x
VrP4FjTRPTqgYIscAEtN9SAh6OyBuOWlGKSSj04N/WhJwf75WwGlk+tkLyVdDFRW06ihSr5FKhGj
/3Wj0aM+PShrWCIUr1QoMA6NVLZkn3qYOvGxS3XCcmtit8nObdgATEspkDQXFWbGg+xiM7+Eqv3R
eH9/bzY4Em2jwpa+bAU9m1NMhpMGPyN9h7ZPzU3qb3KFPZoqafCuRjsZixPeAQfHlWMj03SZ2kao
YqfzrRT2pjDQtSFH9tLim96RnmatSQ+Jv5uiYadmX5NmmMFp4vVtp2cSpnfG1IFPQ9Foo2rI7pY0
fFfLfeGNyGh5SyETR8HsKI+gqfamz+47w7aJ/ZfUZ3WYxiCsrgbHGrOy3mXnZNHM+SbfMLntkbQN
KC/PVejLIg2Ga9yZNRgDvtABIAdAj9lfthYuywazvKGzyGTZluT+1Tx15BXE7DC1qmETN05DcdWH
tnq+PD6trur9FmY7tYBC8l7tsPZbUjf4PNU3Kajh4whzKhPMA2W+bhT7etpSk1XpDof0oaDEwhe5
YQgJxjbUUWnzDWcvZyP/i1wjiijgphNRjahROdx2mva/972RuRAJM0tjWoM6bMAq0tqAwzP9EOZM
9BhTpVFjojeHdvxZfNFyV/TMWTOLoG+nkGboQt8e34vviqYlC9SYKiNJWJrHwJpNs12K7qsUTheP
SVcmiXTo4ytSnLd9zr9jeGWxXqmuBxVY75VXntg0JrOdAO9DmZJ/CUgmwhLCEIl7BvH4c029iFdG
lhVBNpI3GgLAFESEZgJA9vl+ucSL/uYXNx5PZkVBEjLEvf+0C7Yx3a9mciaHd9yjVX7Xa+iIVVc/
sclFr+Au3kBeq1Yv7pZ/O7hWNFShXSuMBxDIst6zenpNy1PfcpQfqijWgQuAfVQyi91AYFS9YPKJ
Trnch/4nHN3V6PabXB7a1NErG/drONsmaKdEYov+JVgkB4XKOfncddKevGWXA+9Ztgj8fWO7icGG
YGecyzWl6UKEyBnaMwSkoXuBStbooFeMxIgBXzO5cu94wyO3i6x4TFHIEnvo0yVLGNA5n+2wPCEv
LO8rEj6K5njh12/H/q3lxT9XL3hwkK1xC0Q6/UB4Y83Y9DDM9rt1Cqqa2G21r/vg1yzegAYij/Ih
0Um/JToskzPedxLrofBTVJwenmDhg4iaM+5Hy52cUu4QeJEhxDz3rXCul+VnaSSnwgYwg9/btbXT
Uxp0LzD/gR7b0AlGo6uw6QlSf8Ozmpzt+K8xSEGsKIf0P1QcLfoumKVR0t2Qj3UzCuvmZEyZeLX4
VuxVvESkVcOpXXw+hHW1ogb8RmB3RTAh1hqQ22ME0CMnOJD6toVReO4LTUgz1NHzoO27gdo+Xb+x
k3qMZx0nc2EfRolrI9Z1Lr5tJHuVTOz689FFpq/qmbKud009VGbAkEsE0e3+0IeNYBDX1W4XiwDU
hsoisj5rT3LhsxGhzr5RfUecWwv1dz4U5ACOXaTBsmQOLXQ0ZHYId+lNrWKvug1nu6fleegZeZim
WBnMg+bGri5p3/M0QcVaVh6/i/QxrD+K8PE3e8KfyrpM7Pfj8Ekb2XZtrfh/GKygQvHz6l5FeXy7
ybdk73My4EhGbKafv6z+GP/G/miF7EWWcDp3L4Uz87nzFjypPe9szZfMT2Dqxcw/B/BlYrLdI95H
wmcSLaNoSsVI9MELjeQKIeXnwXSwHdp039w9tsZIv68SAGfkIU5ib752a37qXe/TMucob5xd4/HA
+cnJGQ08HQgY/9PRPFl3Z9kahzcJ1veNxdfP97cgkOoLH5FmKsGo3vpSEfnNGsFxfvEZV5yXKCHu
ADpGlecgieQQt9NqVDpfs3YfKUETeA6Hl5/DTS5BZTKRHonD97H46Wn2cpfxlO4A+FoiTcEkgDV4
cq9ITi9x33G2/NC/TMQ/5hHjdRojMcI7jtBicHHJkT+E4T9oceSLC7UowCJUvhnuTAaFxvJ8m0xD
FdIkHr0VrOVaNOo2Ch4r49JSXJXB5r2AxczfIQ3CCYvVf23ny5NWBio7gML+hPaEh3hY8gET3POO
ZvGmugQ1O6F+kL4wIPJymR6zMiAnLTkeUbdJ0BMZZvdETjSj9BnxP3G0TqKI17c+t0jvH4K0eFlP
/R5TKjgs+BmVrjXimMM1OiuNVyVAF1OP5qrIWqLvAXCCyc3KXaGv0MvCVWkSNYDIDmWuhcTRvEGh
YtLOzM66DQqNIvpMIqDMsCZHh8dGgMzg4LX7osxxrFCOzbX9IOaLD8fIVXbOlPnt0gDgBseVDS34
IcA75KMqH7Q7tF3OdIANhp2GVm2hs2W+UccTMyWFFy5j7nyXP+kofy529L3w7koLDmsD92L4BtQ+
JhGOiu99DcJ0e35bj4FjDF1mjBk79On+qtn5NOY4GdePvlRJWOhycPqMgR6vhqG5w34mC2uHheRM
6R2Qf2A2rpyWKn9UBBOsLEfLXg24Rfui4Z1ZgrIrF5eNRtAIhDUN3JfXQjMofQKGAcLcBttmC+2B
0rI7mHC78zVyDJh+zpSXz7GfmDqVKk4jU0v4oxoYV11rAAYjy2kVW7upbNSHMaNNY+LkHd5RTCHb
ZQ+fsz4Q8UKlCqBNuwje805Yopj0ahVfi5SuOOYaGfLcoUk2bekx4fPNa5vu9VlqP7J4z1fF+KHh
4PWF+SsUIwW14FRe9WE9OIdr3S54ad3B8449i9nTFB8prJLUg9NieEliM0v2SqZ1gCNuv0zZGZU8
6TxP6vdooAeGlqa3Z5jo90uisCra7yu1rNDxazPO2k09OQlGsDdkEO0uzpDigIFjMoZ/LlNczDzo
Rbj3CKfXxZoOwW4vxiNdHJ25Vblw3eTjPkA3Uz4cA0q6qfjBZkcdyzHXZcOcWpP5yBq2JdGag8Xa
wvkyhKB1DQ4hieVFGFfS7tjIq++TLhG106pcQHn/n+Ro4udu2mxT1aakqP/YLxT8LtuY1D7tuWyt
HYFVaA7DzcYHqroMqeC3O9GpRU79nwhxqn9crc4/oy7C0ZyYUzEHdHqSlRtcsIb+qYcrTLW/o36t
lcXb2BA9/b48oB5tdCCHTtFEx4L6qV5Oc9l7BW7JeLtoN8U9AX3wUfy9PydO0pRVQBIoasIzzujr
U5hozXmzPYZI7Cbvs40jtTbJLoaFFM80IYo2m7bIzmoW6yYWTrtToiO/GB3eSAE4QsPoDrtQqCdp
mouUzJxlpu/gJOSATdYO02Q8YF3R72cmB9f7cjdw4OFWY82muqfoQCj3d06RxlCoegQqie/QHwt7
Rz4zyF3LqSbZDUS45Ed/BJLNkK3hMq/oVhoPdDexPd6/VIoKqotvy3HIuhyucwBWfbRWQ8J8PaQ8
VGs6Y3B+ws8FPp9EWIf5cLQv9opUIw+8zbDglditXXNh1MlX3aXcbct/l0xFLWi0f1s9iD98aR0t
UqxmiZDyo0ovEMXGbzHhUxmNAydUtoP5tRQxIbSyZ2lhvOrT0wQyv0bTpLP1Tu2at3nwtceqqkG5
K71uVsJZEkIxam1FgHfp86G+k+w1QCZpSi/Z/fXg/jjslGgE6ggDMUAiBB52DT7xdO61knldCkLe
s7vQzWFLCyBAqivvlZ43bTvzVmMpr5B9A2r27v6IVp8GLJidJtAcNYIuq6b+Lu2NHm0hQOXIqwNL
9s6Kvt9bK1SViG5dSCvvOOK7V2i0KnNWl9D0POFthKRtWNV3UqrlN6VufTFaLU3oFOyeiRxD8Cl8
FQA4yJcx1hfdx72d0EuKZ9KDuoY8Gi1G3vJ63s1bhvoNV5hLNkoYBNL+AMbJaU47EhhQxktWReR+
ctOH6EGc8dnUWwzuiA7qeaic5M2GdcNj03A24/y78q0NxbNkYuCg8bkTLFfEiQTkWiQoLGsHTrJx
LAyfRzinq+H6BYpYGxvVYESKIxeKUUf1R0cwoVTDpzvL1CzbdWum9aPiJJXo5PojdAGzgt6J3lNF
1tOA7hU6fNt+SsbI4gZHemdVi6dhTgB5GdFjxFoWdtvxdmXNU+RdFXdX+uVvarbCRTQhN/DFqHJa
BPjW340AWQHbXuzBFMP//eWwxWjDLjh7MaPH1/bah7c7lMpyTaM5Z2ZhX4AkDKp/jgblRCJxOIgr
s3mpVxti+acP81anc18OfGSVErg8lZYfdip+vaSKgUUt4wDTJxF/nLcQHL5Z3CuB7Y+Q/+JtEpIE
dH9eNi3rCn8/xKDt6C41y+SgFeDlZnTh5OFeNw/6RbG57qf/42JxJCIY2JA4VCBexw9QtnVexDwJ
PbAMI7jp7bRgUAUeN3uZ8Hx7135U/9P81DBssIVVSrPJV/hAu7Ty6FhV07FyL/M1ENLS7OWbG5Ln
7i6813RdVO9VE8SoOghQiaZtHut3X4YrDkNSZBevatDN7ZVts4xhW4mhlA9ZkL3kh/6fxxDZwTef
aF69cfsCx9zkUUq1iSx3X465zGTUSq/Ud6KoEHZOb8I5JabCcgWHQC1kyazijJlT6wQGqZ2hrOrB
X2hmk2lTjC3vgOjTBlLZErfguFDIt2dJBVCWpLo94F7dzG2JsulB1IZvglldRrB7kR1ITxFnL5Xe
94logBhPTmrLihtxBmhn5upb8Zl1Hdx1QOjuAURMJuDNXUFAuH8o2vSzvUSZFuyNDcI5pp52wgJR
XkvZ305iY7lFN4Q5HSUOVB5XfO4ttcbUoEFlimRNPc19IyGy4QNtF5JM69KbGv58f8Xz9lDMyZRO
l12Rrfmj81aj6BF4OUrBHwXVozP6J6YBEcLg+mGcOqNGCzvkrRpj7WlJB81VfeLpqykcLyhYvCJA
zTlWnTBeOPkCh6jAntM76ApIzZNtJvmt6cwdd/NaPEkWEpZQE4IIieZXvlUUgxitiLyNgaYzpJne
FFIX/M0iYfLRwG2eEcDQ5EVEbMEnXmt51dyRayM6dehkKbxZfw+OlVsV9ecqw2CWWF7yi4I9mo5T
a+g86/uvZmWeGem3xs4hXh5RvONoRKUsuJYdXWYrNy1VdUnYUyM6nCgbrVGfl9XrnlnvD2SuclCe
ERqbDxXuqwfp9Y89nZgZ+LqTp8h8LalNVItNCt0i0wZCCvBBBSzjYizNDT+4aEWxex3gKHK+fKIH
0iLEuf1vZ8fOYKOSxj+qZabmUCIlvvs1j7RIU84LQtJlD6YVm53FfVrLoWcNgD1lYyXFWl9rIqCM
Y8YwE7CcgS8QHosoDJdWUgg0syVjamzJrQGm8c5NIcYp9qaQQb6DzWZl05kQh3a+iE5XoIeQIJrw
bZzgIPwTLEk141/V5mqVNji08hZhDeUmTsXcHmG9EGJGI7fQBYl2LkDUtqeY+8jmH60u6NDAAc6F
CMxOERwJ1+ZcszFylzIQV+s6cN4XjnETG2WeHHyL4iXt/QQJ4JfhuRPdfbEVVlnUZ19H1Qpy6aaO
UopKYhRrq2X6mHi0jS1J+Mdo4kYgbCSyg4Fo/JbeLQrq1gwZfp7kYyzWznDGV5N4Bc5Tb5NbCdzK
MVgu8UPu3R+74vi5XcuUOG+Hy1aCk6bjpZSnxy4ITyqfl+vb1O4oaO7MY3gLIU4a8m++JaMJFjm2
dfaJGHUeQRBKFbfC9D1ZKQhsjH5CIX09wSR12N2Ulm9VBIVaaHg8TKGUfi1k6pga9X0QezJa9tmz
91UfqwdBa35RZJbxtnoa/n2/Ztbr7mDXZxuRDI3etxurehIyeQUiM9zIF2bWxQKDYLK5nQGssIv9
3RPVB4EFSGsfFNis8UQCrfqY8w9zeq6FjKBi8hlGGVp3HsspLu9riIvsz1X4XyXcx2RiJVhZEoFN
Xrymh7IZZomUlLRV2ndTG8/kCNhdvrUGH5e6x074qkSpUBTgi2dXLHqAqMblsLbbv/Z4bwYfOdHa
4Tx5Y8Nh0NkEX2Kj+7zeK4Q+fBa6wf1wt2ZPJkzvmPmVp9Wbn9cTMkqLsYP2mb29r5WRWurusATK
0h0CWu44r96PjIHugcILLA3CektIdyzdpzfqDvJtJ16+LYLRG9Me0ABP0bD7hDUzXgcEu1W5eu2s
YYPNXPP1pZkQ11pq0oZODw6URVbk/Itkx8Fz4eBO+JnnOet4lqiUFtixJyuJIX5JSQtEVo8GseEU
GuhORuD43Sij2v+x3JhGP/8rJ4vLn0/A2dvjoL+G/BxdeDXt6viI0kAIpQWgJekDeLac+iMuoQZg
PYFK0/TEecmCW1PpCACtYkBOgIGQQjLTHaiCeRjcRjt/CHK1sKQrguDwXiGPShOOBxBU70boutjB
oeO3j3CdNPrkCo1w9wSXYVhQQ7Kl3IMZV75CgNIAFXqcbO1eDX92pSqvG3hZNSuxqRSoI2Y1UKT4
x9jsHaqjLjoZcbnGtDaiNYC2i9+XI/l0I9zw2BNFLCALhwCcUZPn2IF89QlXdgVGXiSUZCyRhy7l
cJv7TyOmMGCaGp232/sFTuCQkd3E+5UQi1Dm58Tq7rqanEJHsiaiUuR0YLm8rI/vneYXYnId5xa/
nbrgZCqxZaIPZ6zonYha4WjnIFa/jR8DeaqFeNavKhi5TgOrR1MuyfrBBYpcWMZLw1zAuz8vaazM
XKHOA9IwJWK8EvKM2YndUVXtsl8kKt1Zny6xrQivkRjIKY9x6L7UTZDK3Nm0Kwj7TvxI1Djd7Fgr
ByiDIcqWvqBGnxxQDAvM6DLzdLEhKf7bEWdVxZGrSSvW7I3/cdPLYY4S+fEmPDrInd8mwuPzoBs7
HDmuZkrnZ/D0yf28Km5Hz4aJ9USEYVj/ntPsSmil+JJ2rzLgXCysSW+cfU2h2y28TAtqjxLdPS/d
O+Ko+h0dDEAvsOSZbtYjdyKLY4fwlYeVHWUPfNho630bUnVPW2fZep00vKTt5MS7jJMyFO4t0htX
GJA2Q5NgoRZ2LjnIHFtxQdFtcseGuKuMRRGoTkgjJPLQywyNHkOH2vBIBYiqPdol1Romesqfzicq
mzR3Wz72+vuicUxOj3V33aOMEf6ehTFleyHgzdx5M7g91Me6qvF0DropJOLe6kjGWqSgEwYQ5AnC
0cgTeFccVT5RlwmsTzY5ZRi9YLZNuh4i5XMr4R1eZGjl4kQOvFbee8x7tdUUjBD75I16D51LxcdU
I7PZgDmJDP1Ku3aQAcxfhKyaTGGutoP1oz8xNIjx0jK7OHwjrs7pQp8TO35BSsfSr5009n0ZlnDa
bt61LxqKPeOAtiT+WAr9RA61ffgpNTfVMMZlVU3W2VfSJ6pubDsTSby4Hk/k4sQz77hOK/qoyCuF
38repngE93o1XYWFZu6AcyGz6woCR5Iv9Hr8Gs4rqPJZh9T5bVAJx+oNU6Z5/OWJOHEeJniOzkfa
Q/2QrCGgKrLAy2IVL4l2fAiCkcPOJmLGNHrmjHO+p9s/CO9aJ8TcxXGdAWiajM2Yd1Lnj3uzowaK
RfLAjoJxbWtmKpGs9rHWI73fk7FGV1xvnBpo325HlZLYMB4FBCLTn7StVxc5tzRL5tf3mlzBLvqD
zr76q3Jwj08bHqm2bEelVhpp5KBuoivNgOFsKcMoQddIr+4VppCqvd2+yObKL7CkdRp/I7gSH9k7
hvhmnw7V0dJrwVi978DP8V5wMJikkvEmg8hit/h0Ml0VUGRZDm6L9gKMOGRMTwRQtzdVF9D06oU+
CZ4P72z6qxkM8O6toc6rSbe6CCLAfV2QzbB7pgltCfSNNeZ9yOm3roMgxNXAXU/x+r2hBsSzJu7p
UjxfILXaKYMmxzfNMUXC3HPjg3mFhBd30zHMdaNiBHFqm3jqqj80T9YHXJz8CRP2at+whYJHPpp3
pCOQ9pi4FQrjSa8xCxb0bgYzW/PQKn44sXZitJgM24HR83UlzEysvym9aLT50rnzsusPpZQWfTDp
tnclHnQ0GmaX+42kWaqGRPjkS9nG5utvmH8zImM5wzEq8uFW2xLf+DVz+RykJSdNnc3VQHX6u5wE
QvmKfeoCudesxsHG+xMRKxy+4PaXc3phIp/9S1RJYOAXjAqBFgeP8xlWwlveuFK2e6CWTI5HLkK1
thtIaY2lBZnsLdRXuGE1cgdlJy9BplzB0tA71emZICiUF6Za/xLu2uWrETaS/anbdXAktAwUTLtL
R5bt0xEqTZ4305UB7ea8BISh3y4toMH7bOakLebuxYxtwzQgMVTGA9kxv8O3gkqNclyh/HvAgCGu
mHZ3bLAZGRIYaRQjdFl/ZW+7gBpLZeU3QqKjbvqku+8EQQXFZHvuyNHPkoo9ZxJCR23PoyTr1qDw
EEJu35LkU+9SN6fHL3dCmAiDzSeP6opiBiAcXbjMzSvZ356n9CM4ax8+3geIoHn+HZaZg6nLnJRW
0vsBT73F35m5fEf6gNQJR+oRNLThyoy4e3KI9TzZFCo7D/CyXV57v8XMV3859chqJPFSTqqFSu2+
4beFZ77w/i8z9iNgwMg2kQEmfvYoiySw9Efq7j0adUOiIQF9qQL0Pqc06cSeHGJ1o7yxqM37l2XG
1mBYMNzxDXOhncHCmycMFelfnJodg4Jh/V8JMsgyfz9AGazJNK49sXQ1x9uJagoxmdx1DtV/dT/T
bNvMhR3Z2BcfPK8rgf+xFmcuk5M5/S0g2Ikp63vempuI8DCQWwanDgpurQhQfQ2GVgWR1mjU42L1
yFPzCJAuLrEFaRogH2ZTkSsBXPOL8AXBxfB35LVTESuQOj0v9pSrogKgF8Bx4fQZorMRNpOwKrU3
D9gPr9mullIkJlzOsXOaP8VkSQvmaE5uL/cKJWncR/jhy74AQwqjMY+oiEN29IrBKiM0/OFyEZ48
U1HJHzgt9OjWrqWiRECSIIJBTqn212stMTKFABMuz76tHwMUVdw5jlGTIx1dTIENH2vjJ3T2///0
JWAV10+rNFFwRYDYp21UVFw6VLCt4SWoVF+e+H4O8ldB5LBRJQbDmqsQEZTvtlZX7CBuW0TqRpji
1kYS2FwTFXmIuyXPtoJSso4S4Q04/AhxHGeZ+zAgzZPT6ZjCD1mgi/ZCHqL/h6/XanVMFEd7juwM
D7lO5qrCUDZllP2VldUa5B/P7KPdIbz0RH75YrhbNBcYACdU3jZySCP2OkQrByjxHL0iTyzJly8q
YAHyGfUTRScQZYVkbq1VwV4igGq/6pJvHKS0AOumzLt77GzyD+jIwEVy2GRh/nPJjmGtfgg/Y+qV
Uv8kzp5+aH3yZJ6NK7SDxhF15Q3cncn89h9Yjv8qOhBM0pj+WdTrXAxNBrl7/8bLMNKbGEn2yUBA
ov0brXxSJtn9zQdrnQ2dGfWrB0AoKXQ99ctP/QrPfl7NACP3g9HRGZdapq/9lOFE11KRkV6b/paP
gPhAOuXGtvWbOahzQt/O3d8DjdbRFl2QRGvu4Jl5JD0swBgTILVkMxIBEStLy9JgwS/8NwfIAU+9
fvdXtz3GPW5rNDvTlUWAhszPRO63B60uWxmKVS3Z4uLeNC4QrgpSPWr4kp0IJdTHsz3lSAIKVV2C
1JSEwGh64RZaf6FDSNS/61J7Aan0748nhP6PEH11LsjbSGn0A4eZJUNL2TpMV0U+6ULolqJgXb6L
MdaCNF7KJOa7xNyRp5izTAAhNqvvgxL3knn2LJiAHEc77i4FBcZZ1Ah79w3c6Q3qRo6UXzyAYwyq
nBqm0P85PHWrSCTD3Y6I6Jhj53bFIPEokYaW9gPN1AAaTBuBzkfOPYWV7U2baKUsU2vnVgmQNbkg
3JnsuRSS4WWAcbSi85iAhww+Vbvvls6Ce8H0tU+jg16Jx5gCc5L4c5NLM0OMZT/HPwO43lUFLZ1T
TzTQw1LeOLkJ0C9EermXdvyvJnEbzJ5v0CdhsgJnZmGEZ//1zA8rELnQN+ZTA7pssH5FY/npAo/g
/6t93jLe/JU6bt0Y9nCGUR81LFX1KuymQ/7arBAemvuExaQVCo2Qp5/WUsAwIY5VydY1/bmoRTnD
pR7KZOR6AzrepYeTSugTBqnoqadupL1tSUygS1fl4fxW61xa8z7r3sbDBgrFxvTPEQIjPfA6B7QS
N82rmAyUG5jbC5MSqRKHCsaCSGPzkXD0gI1DJuseYpHsLDMLSb0EjmcXDtOjvmIOzBGuf54nS7KW
rd73JbhFlcJjzUG+8MZ8YG5LyepJVPFeCqUCgdER/ylxGEYGgOWfV2EX1WZrn8DOFXAxaJbKlniS
xS8UuIQ5hNAG7uQjGUGX78IA23C8CsR9cH97QEBZikbP7UPmkfrd+emIGBjNGxGAvN0791HREMJk
Bm3PvrnffMVfwc5ajMrqyYBOPVLHrSE83VxftI8MiEvEX4dmjqIu7U4reIEEH0sd0i2xMovywxBg
44zANsMqjnkSkFpGWMOKW2IeES7kArsXFzDqzyrEfXkWsLLnri+bv4r1jModZMAxQ7atA4iYlILM
WYW9c6IAlOC/ZNPIF29fV+NFAv0vN9gk/z93qUKae6TYgkODjiDKCmOfgEQ3+B+h2OKjaCEy65Jq
t5JXz4heSSuHzijYJM6AaqY0/KWdr+auxgyzbwNHb2uLaVNFRzwJ+qggHmZSKpNNVI8PYrvd1Ke3
iCQqhMLdA3h+dxGuTv6BTtq8zVs61oqMDhvcqpalyUClMz31RWVCO56XSv+9jroIKIX2q4jbyJr/
zW3dQq/8fiTT+qwmOkdrz8nM+mdsrNMD6xgedQPScaXo3FSh4OtrH+ZGKR8QWPnD+WIUJwc8Kn0p
x3vtD0YdiQ410JSpuXQcRM+v0X10yfBCU/4bDsL0t9MiP7h2CaDMdRxE4pm2GvQvXgPw9touGkXy
yS2fsZFlpCC9aWXA4HAPO+eM5iWaFBub1Etvgmz6g6urel/Hz7DX7KmYGHjSZFz3hlKd7maLEvkH
vN+5tDuVLHZqohfWZtj+8UWynu3OhRWH256pzMx5f5HNkVZ42KrcX6aOOjH8pIACkSHW9dAYSg3h
KRzJFC7AiHzBkPZP6yqSL+fODuyNR7dAkF0uVpqS0WVHZK9X+8nimMy7ryv+D/NIzhTrQcN8sH5Q
tMHbXRL73N7eLrYHO+VB6yZYutuugCdDDMB6d4RE5pqh0WsqO0yCKdOjm3EqKXNbtTuVPcjM3NwN
y5Dqb27AtY/jj+lf9bP8fE97iAeY+45k4ESQwIH3vBnG5o9EFEw4JGLL1YldwuuZ3F9Jq9TeJSM7
AhJixU7pN1vYYkxo3h81dvlVYTGQDhhJ0v1vINArDIVsO3d+ws+Iu3A8XdTms7ABtIVm+LLVLNjo
qpELExtKRVu/Q85+iIrItlest49DzB0UpZzTr0xfKkxOC5o+FEHAchM9qrJdvWIcuCWwos5g3AjC
j2X6+RYRZJmHEU6mLvH3rL264odvnaF895U/F1r2Z10IO6aBckgfL71keoXzgKwJF58aAbkwIxRi
QslM0LUM2HxsEwKC1RbXyCSSAhtBX/C3rR2cYJTryMFUBFz0XTbDJcryY1osX2BxYRTCU6XdMVkz
jBeAbtNu+ezyq8M0DzMyzDlJMaV1BJKUVazUPnEnnbCtqZY4CkbSbDaVrgOzZni1PUJc7WjUgiCi
u9J4rM8O3plqLiIHi0CvunxkQN53+ClFIfkBNGr0EfCOr0MlEB7NnhdLnn2XwJ90Lm53x/qtyi8/
p5hjqmsRjj1roAWS3xgcjL/cwQcXb9/8zNAyXfhaVzKQQIGt/cnPdd9OiAK7zE94Uq/V70r3bTgh
ZT3Z3W5IbNLl2Ve8RMzalSFy1hHGnRzIfK4FmUz6NwdZs4DFFkf7eqKFzMMMAd+5lin/qbHQtO/I
gXahrlnmyvjfUGTxZn4WzM0PpunGKJm358bHr4o8IdlCAmHhPankB4vJdAHJdcBuZ/cpj7Rgxxxx
HdUy26ZmtPkmZ1aYEML7L1bvvc9yswNMUPLf/R1gkHZwqAk09hOggydcOcicGscGlAA/KKlxdi6d
l8jaFjVTftU/6WZGr9P+I0q4VdF/TgtfSRyr2zlFL0FFkf3DMtRHDFjfh+MljDfVDg+GEOS4UN82
Foubp8rfo2o548QibXHwpbrIAt07EwvGHyzOJLdz519oiW36uWXfHHSjxq1BdBdMR6rW0yrQsIUA
FSgqopFookCEI/qvZaZDlf9i0AVj+Vh3G6UzjZkJMb2UD+w7sF1B8bKWyleUnDj5+TSBjBu3HOWX
ywSRw0aIY6QGOks9tvhPY9FvbENx0T0RUMELe6hCYG9K6XDLdktS4VJ/QIjiylXTCyoKggqt4XeO
ZwPi4+BYusk/LqHCXTSrHtO0DullgIyV3Nj/S+m0LJa+ivHoY5eFBNBqfbTr1bs7iMfuC4dEuN9q
+7yjLPqnGn5i9zYaBbvqfJsGe7lXvJuQihR+LYS38wYNvQp5Q0UCpFW7q+PX13Dr+bD8+TbsJ/Mt
o4IjCvmkRkMGLaRwm/LHLnAZ76TmB1yzQRoYNPiarUsRqaIhjFUqAq4vzyyrfSlGdkVmxV7Um0Ik
V01/lFCkoNLAA3j59HTH9p/0ITXsjJv++boAplstaG90IC7zrQ1E+UfZXsZAl3NLrT4buD0eSo05
Hg6eEtsc3A1ceLkNIgCIiv7PzdOKEEP3vc++pWLACcRtaa8GnOpHGQ/GmfB6L5Gy36mRFDGhVqgd
LeDA9roKFUxjF/fxda+3Dc5S5a4TxyUOXI5IPb5ULIrNXQH2nMimA5kFSCpHxER72BPzI6nGWdMv
5YSVJNFR7pJQNEjg8bj+btH7baw6nQw5kPBmNgdlG3hH9haAjrZftSwBVM2/a9PELl0FNkk0DNN7
zE/tbjYcHu1e4QQ5kfPRYaf0ueYX4DAD8wqM7IObmYw51rzXcfoR+et65KW6z8wASzzZvDNf2aO1
Dw/IQNIsWoHlqy81tAQPbK/RDg3egFRodNUGaERHlrz+F2OvTGu3UlBVvJCQRoVVv3uZ4Syuj1Ka
ozpM7XeEBMA07ShY7usBV/LQJiH8S+CARp5B1Uq7Oe+OTjiWXoXNFhK/Fn89aX57X5o8/zwCAp0g
kcsXDwcifl98Iol3yb/p9piqgJtf2pfZVKwpuYrXOxVjVxmIQDohDoVkGbFvKo2eGfzZoHENkHpg
qN7sWSuQBd2Zc6kfaseGkac8OxGg/RaJH5Vl+K861Yi27Lz+YeoKlM8VlEVzXOv891sYZfjy56Ff
lfcgswUtZ/lrBSdYyQTcMp+LXXEIU6YkIoJa8JnpkCPiN3dZJdNuVRMaYXToX/scu790Nte+RWp8
Z+RL/BRyWPCZhbxCErSqaHn9Zdl/R1V5/NN5N9dfdAcmM1Nuj79QxhGllm3m9ltUcYAtJsaEnmcM
hk9e5FrVqdPw/OTY2ghoq1vQ++fpodHKziPj+/lEWEGMT/+Zg53Owe3Gbf7rF95L2NFcUG+RcttA
n966/V6NCHNGeztqgNV59vf+NYNCd5pBdZPqWWd6nOvB+xMYV9e28wDtT0SQt4fQD4di9ljBZluV
EJ7LhgD7EBu2iQPAcSAAlns/s17hMEUlD0htlXLFW/waAfW9g+ehJGa77lz3Pf3cUs/FdRSwWLEM
G5Ro6OJYxYhyIGlexmVtIYfnDIheNF6T9IjFGEeVA8AQwZeNH3XY0N3tnjwwhdEezkaBahqw5GaS
UVw6m0mYCHX9+qA9NQegFITP5NAgjeho+vw6GrQ9jupRd2mcfDAzrASRkda4KGIZXhGvFNxTSe8U
nLu7VplaVr3HSzpfVZnuPRqzcu2oDSeFcSU6RwDymrg3oQoGffvIEuucu/+SvypDvVEfNMNDql7X
eF5bn53zgQ26afvl8Y8hAzULouNYD4AzejBOenyEAeQtYR26ACyQa17n7DX7eeF9aalWjLrWkHW+
NCa9oPFch47IrWHuQ4oib00M5Q+r3l7KyeRDGePXVqmahGunFL2LVBldLI7YLrTwDrNPZlE5/lT6
UJCav2726CaMyGg5kB7HDg341faCx/Fj2pTQa6tuguv4sRjX7yfkSr0fzvLxLdpc/P6mC5TyVpHV
iLEZBEgN4ZUk+ej7pJHMJB2YLFbM7B5YFinw6lO7Ob5zgi0wwzF5yaMt2PImJgTysuMcUtusviDr
kuwjvLVVE2QmAH0VT7EcBpr3m7XPQE/k6ynSO/L1BfFdmND5rdg+YoiMUZg7P6BjqmX9z87jNL/d
kIwky7s9HjiiEIrfw5hSfOFdzC5gpJLWKno5MfBJf/OYewn/RjZ3lnt8toafojgedRqol6YN45/F
HIAtyBhyNXGeKGCDSYORbF6edcIw7W96aEOdDTHh7P7cec5/e5j7SzFwu9sSs3M0Pr94atvHoyVZ
qKf6wH+JkdQPyl6jqOBJrwuEXrddH1YJR6yCJ0pnCgSUb4kcKiCAFLPa05ZkingdSb/NKH15U6GS
rp9QVEPFmN9cRHaWcInUWvXP8BbqWqed9aFuDnQnfNrA0JnZQ+hp7moUW3X7Cw4k5p1XJBv3XXah
+Mo/ADvp2WTjmojugn9LB+5L/aUf9+mdwLMHFW8zTBm2Tg/Z+HjFJF0aYOmq2KKMfPHX8IRxVic9
bk5hdrsn9kzm2/f2ekkkn4CN/ByMHlnyD0puP7XWZzLKLQ6vYjEZ4rm/Np9e/NapZvpz2Bi8olmw
lsPu6qsAcQ/lri1s6FUI85rmBIBXwXidLtoYbDJKB2MgpDS63Q1oU5cTwQe454tw97m8Bc32QHHB
/f1x4o6XaIXUT/qNcQNyDLP27GEU5i3UzEfkDwAG5TVM7mqJ/ViRuYmmzVhnYt09ZGOaIH1C3kso
Ci3GYUyv5oxYzu5TRqHMuRYZN7R0iENFtaQEjbaDkocM51CKOV3YopNHC+wEL7KrTjl6ZsIYPLMN
QfVOujXWE3x5HnPrILtQzgoC8u5FBak7EsI8l9yE8On3tfFiotNcEqmXXX088JbpZ6ZzsDU8q7et
lSebIcQmn5J1mtti/U/Q23rUcbZUo15DHtm8OBknITsN9nlhbKxkijU3L412KIJzUfRdehZRAGyq
SADXW5Wf63bpPUn5QOycR3K1Bw0iO8fLhBp8RjMEMyFzs6wj++hQU5cgAixDBiQ0ITe2x68szmlG
Xc9p4k5QzjfKYeE37rSi17NIR/FHNI12+ucNuiFO2w5Q2irbV/351zpeWNuCYiTVbMob4d3U5MkJ
voWlFuRpuus9gM5PNEF1g3qR5vPUb07AdYJFwoncexJuKvVuioBpc9yz7ELw3h4c+LKmm+vmJ08h
vXwxuaCtsxjicRivkhVH1s8FUfzyjxSquJAf+50DQcCo03yoT3Mjhchy6g3OSpJiJLxxIDnebhuO
iJ2qRIRuOtuo+vAbKjSG4cQkIIvmGPQz5hFNN1cF89qhUdyg8RtU1tOryceQEjdyz2lFLwadnOcO
9LKY3nP25mbFMIvD6J7r97oUHtY4i3Zg1yigg6NTB3k3Bu38fvwemSytogLnEtbgwObVl+W4JTo8
Zu8HsM+VNpyZ5YdSB0WXyb5UM6sFRTl1fkxw9MSWVYvDohfDxl0PYtPaTDLNFeH33Nv4nugn0XaA
ZG8cUvLE8aDIPm3ZJZ8oAQXH408YjVwjGJnGieW8PGtvnqymlIG+lyF+IPYW6YgBAOnFYH4N/Zyh
OhcOEmY8Lh/USs0UOnEmbsswP+vIDIokqgvEehqPl5uR+BiMRoWRFxGgOY/5svGqQCDnobFHQ6PR
FbURjjtTxfz/3TT26D1UZbkUyd85aLWX2gtCBBHQAWC2LnNOMUdWS3eIoed8zpAKGg6zeLNCNaZA
oQHhD59MnVZaYGnLqyeLoXXDZSo+Ejw7hy1uIyvcp9gcWoQz5OP6rdVhYC1SdReIvIWnBGNpHdrn
NmUayo4djh7g5DIvHS1WBP7i875KGMCJfVZBJ/88DfPPnaaoMi1KP5SUz2SNC4xqOogJi/quIBxj
48DucUOGL2rVHtTco784X4Q4js9yYq2v3GB7US/uw9wGNbPlTejwZ+NfWtPhcd2fnbo5TwP8G9GA
k3bZrkz4pByWyK9mz26cMlPvnZE8iBJ5kvIDtC3o4h6j5FDkUurW/iVLl183DHBMoOV7CRSewDsI
aJaItBQnrskHG1eeLCMVAbDtL0WdWkMJqegcS7D/lgct1+6b58+Bm9U7La8Qr2RrsYZadMsRDZca
sQc2YA+rXdFo1HI/tskD00iPO7lfh/zv1zuqmcp/irJ0GICQgFhiKuAuHs32A7NeBacAIHxWsNR8
PScTpjkuCfKOUduE/ktrCVpOp2POTf7Sg04CVwCYqXUXF4ykr4kWygH7cWImjEJrEqGnIHzLr8+G
Qk4qgKbPeSVbqyHBt2/RQUt2y08X4Z5VQ6ahnjb6plDH//byx101IJ324Fro7bxkSEHlXX7X3ZP9
PKwEIMGl5cHVeaASCZAB3FBDSuFjftyFyYBQI2TqVa6o2FJi8mv75/bBL9y7TRTPLaz3jwTeIH+n
cqlItygetZLzWluOHa+N4jp3jE7gpcqBZL9rECXmXWyLWW6EgOfJxWKLcOMWLcQatCZ+OLtbsO5G
7ME315OU0ueH9otAr1jnR5b3WBgAFZYXyHRmxvXD6OWCefan5RpsRS1Q1T6yFujFexaBf+jy3F2E
J8H7adewNNNOJPUMno9vnfO4kqm0VIQt12eki7lFvi3dd9YJ5W7JkSazuxLkjt6gkYcarV9Ir+pX
M1rcUp9spR/nqbJJNuvZxtYd23wug6iMEa8FsY6PR1JZ5f8M9ZnTFSI4R6RxmyYxhNvXPaZBz9S7
n+S6bjPDtqj+jmbUxiYVJd83WblbAZBrolJSGZbzLt9jh9ghLOruCHaTeFDNZ4P4VkUjhxbBzeoW
plPBLo19l2npVd893tDYI8dto6lxW5sti8rfT0ww/r3yJoU/saPhPtCwc0Rlys2zGKg4nx8L1rh0
vxt1nNWkxxmcWuqWNG6QmWphF0f5qfKZI0MoLuOZlOsD4yfiVWkxG6YnGKjB9Dxc84SqhRRArE0w
9k4E6SGUNFHHrx4jHyKLJUTz+RY+G6ipaycsivOUPVVlJJpWjbtoeFxf5iPi+Sjh2vDPXvQGnpKl
ltHq7Hr5jAT/k4tJpnWgTk9M1FETDRxMVl14giEHroPuUi7u83Pckfii2kL0sm/g+jHj8sSWbwyj
dV/POP+7ttXxLINRqUXnMoyLi+zAITQAMjM1rZ4tehBn9EDdnYzSYEfrN/niDF9tB3Ja76MyLm4F
xF8zdDvGA0MNDU1B2JkxPs9yZrN8/E7Hv4HwtlzZdCJSU4ynjnuYndJ7/n8q/980CxY4Cpyax3UC
6lfFSoWD1bTQs9AXbajh2rFN76mjS5ySORBnX4h5gMZGBfCPoRsGwFQdRBRzEfy0j1k6faBg3mnn
SV5KIssHpwYEAhSKTMBYOJ6hJwcUjdyP0DxXD8XxLUI/y97XP5EBObRhWX82PVkqa0JTYhC2mB1N
G7e+3jriL97RbIsniEEud2Len7McPNLdXrXK+/6eKd8RMSiSXBvQfHcOIPZVI9vd+LowHQwQARdV
Y+QD7hiLy93ztIPKq9TE+4ln6VvUfT43ZBtNOoaauFtF64DE91MFnBD2ovRFKvMQzYBu3kvw1qQE
HIgr3KneAX6yW7Y9vfb43iFTzqUF+tl4aVGXveyIoGc7L02B1fSdqTg7ESe7yagTddFlkdT28wwm
xb27nV4a6GPUSieGEK2s5BvEjy76SyQi/Bf2Trm0kcPltfR/sDDbxEcC/eYWKJ896VnFQgCtwU6I
Aqzobq9mrbDBw238XF1dxGqWU5QviQddBKJmfGk0WPvjcGAvVq29Haf3Gkv5y4F4bJcYAXdvRkH+
uc3tSZItTWwyHSqvSXeF7xA1MK9sClX6mjz+nB6AHf8OjMZrb0a58tmw8rSG76btedZm4cUWG+6i
aVO9Quvb+u4HENadqNJ98afkGmSApIA4woOad0o/B2MCPap5IU030edt5Fnlj+NGjYJZ8akWSDjl
WNq+J0M0+pwUTSwkLrXn+sFgx3zbR6Qs1wLznks1YERbViicufz5qxGnJRzFj4fOrGRFEUEgKrPB
b/XilrsLuIeXi9ICYcN0Tjy2GH+KDkfVOWj15XyC2YVLmPkODMGaiF0NBVWFi7+GFs4WqVCq5MoC
Js4Vj5yriVJEYisA5PxVZJ8dRqMMwsvF19yxdo6OjVz+A7DcX4uv1KbtY+SBHHE+vCYXdyC9H193
nMkeUrif5cxI1dt0kxqUOiCYs0PZVl9zKKBW5bajV8zy8HLXtcfrHLqS6dfrx0iLbYJMNf1+pH2n
nlZPFdSbkNyTXlw5lgcKPUVG1zlShEKKsMLeI0R5+SvBjG1RvukPww325Ahk3oCwzmx7k/lWHsVz
J9KcCeDyHKIdAcyFinJEiuUy7sYvaRdt0i2LFtDP9s5QAwuZ1pCUAQWxzZFHttYUQ6vHGDL2Gb8m
V4EOKehfCvbXEMw1Yj9xCjPS82/NEkpx4hV+USPgw483cBBrGGLeQBMZtEI3IwkfRGn2hGrcoZql
yHC6jUzrYr1q8TeJ2I8o9LTbfZgIAZdt5x/s0md3HLAp9VykQgVbQnWg561VPihTovvqeQM51Rm9
lLecP9Y6SYeDPIeHKzdBoI1HRgQrHsu6gwood9CcOzLpLf65L29GcYW6ZlILfR6e2MMc4WpGOWGP
0gXGeyylfTkvg0TNOZ6VU1/4ZnyHRo5C2FIGNF3I112tJTYgdLLV2Ehci29gTLfTDwPCXr50PF6x
76czQqEgY2xKCNGZAjTxImD+LXwFQqNPSJr8aqAdHvQGpe1vhXxPu2/5rRjB6v+UjZcn9JilhamN
TqKjmdZzneiWdlSiSnsiHUwaVPByGvI7kjUP0o6/DHjprfz/5qPbibAu87wz+S9ccFDnd/Do+s80
Y+V/4av7I+RfjByCJI35QB+f/+iDBZwkRWqUHkyhZQpWJUgfQkIYSq1/qtisbYE5p5d1b7NR6sBy
JaLVlDXPFvTgy0EfMuM/tu3uy7fAX5xTVl/y57GcQAH4kV1FWp9R6jGa65umXhllz6TTZvAuLSwq
JQNRkL0unG+FvYvetwbPSMn26Z6uy3gxs9EM7V5wHSD2NvrJXTbpmJvA9UmcqZg4RZ7pGLUErd6W
RbmCFvkTZ9YK+8C0Pihav1YKeISa/QN8ImTrcuL7ZC6dHClDoT3tsRRsQ6IHqsBmeoEhJNsbk9Ew
TnjNukxZPOMMWti/5n9kzwXQQQZHJ8+JFd/SUAlfPPQu3pP5Vt8EKhko9Y+iRzxdn+T9kyt0E1IE
clpMatWrPaJxN/2Hey4xHZEZ2QnPrx2tAXrNMzhiLMfx56I7qJWdayGNkik1JnVeEWIIFB2N0C+1
soILo5mRstGBeLATuDIyy5oqWN/zEOgCxueJiUEY5HNh5gnRR50S4hSVcXfMxALbt4PxRei+gXSC
CmyDRRfD9kdDUplB7YpX0cBIv2+VlrQilCqDvT1TY0K3YTCHZSMbF3+xL2OMYUE+RRDrgKEPBN1H
bfZfDOG1AUPV4APbPfPfusbF6U+NBryhUM5trvAIsN3n8EArOYbsBfnZbXlvbq1MXTeNOe92KA7v
ynFVERrl9dLm3Da5lfi3kDSgf9fDJMKOiejnAy9HJkWBsYeFrOlA8jRjTzlFnbjbJDopmb3Yq7Un
haNJcHSjtq5n/klTftm7SMeFQhUchlEpptFGI63fnvd2VITQtAR6ZdsOJINdgwpQG3iuWxaFDklG
FkCW45vOG69ArkpsVTh+T1j76SkvstxwmC4svMyLAvAzUcnEeny6n+6XapnBQOToKdBWRpYpIKLr
YEUzSlfSY2ZOykmMnUX1GHM3h29/Dmn0BCGSjl1N4Bs+VKJyS6TwL/10Rsqrifb5WPqywJHESgu2
E3+/i50cMcVaZFV7c7wZuOPcbqibDnhjWtKv/6OSTTMBrcLebRb9lRiZn+X8HXfY5tw+iClAsiku
dC6MloiFJTFlDCoaatcIRCplArqLo0xUhLy96PIY2hn8TeQ01+ko+ZYPkmdzH1xAe43/x+tTFZmk
u6cTav76DcX7Ef8H1DRVB6liWBbkUfo3zRHRgtTcDNuXu/loMXW5NKn4gd9Dowc4xhC+Lhsgyluj
OTDS8hVBSY9xSiQ8ANqw2WNorjo//85d3J8f7ouXMz8foHWfKiz0BAAvSbRJ07jtHxJd7vs4/qt7
F++zwufRHv8ZEeayB7oAqvMyxNdrtU3sm1xQlmKmL76/BHifQ+AQCKGJBwWtNx0E2DSV9LGPU9AP
tpzAfdFQsknXVzMIIGQiOXcR/XljGY46vhE6TA+ncew2pYOGAWZrg+0MH4bn7/+1HInfkoVLvPvw
GPMNt9CZEnJBGLyc6nPpQKTfQWKY2jBgA5MbhkBbYhtqeKI4+VW01osYpWDvNyOhyHUjHmHBDSwf
X+/R8Awp9VjUsbDfFKHgQb8xU3c0Vt13/Ygu18jSheUnSzI7sui+pIpPbRtbfznYgupys/Ist+iT
abzjRmFlWQIyt+zsm4+ZEndFIyR8C/RczlrKCk7iwinRQ2KcJbJ+veEarPwmhoxTOtASLzTf0mYh
TAdImojiWCMSmHU5Ua9cDd9T7k+KpdhR5LwOAP4pt1JZSCY6QGU1BosGX+zs1852S5UVf5+WmdKJ
n5ikhCQJ39icPlVBGPy8t/XGxL5EmJFRQS2Hm6vCBBTPSeImqBemb88qkQcvHoPT0RnD/Pkl+op5
ckJiEASHiNfJV5Sp+h3p8m0GkkBinsHhVp/Wic/Q9Zk3yBzP2I5KhmxFdrBVuCh1yZTByBcX0IsM
+Vt/6+SeMjqqCwY8HgDw5UvPB2EepreF8IvFeZ+rcirdxibHB6xG+f2mux5/62PHbQfrbDIEwnKk
85A6teABAE+fEgo7BVNDuWGbqWrjzi0dhl+4mgihhbBHR0r2jbk5eC163gGFIzf+PE+4KRXxEdil
XpgEbQT09GJE5KFa1RMba+uS0MpmnAFHhOzmNTo7c3wxMG8I0wqWr1Z4IO0E0qBTQvUOLWmNb1ve
Yj+BIai5jzytuYoRCzExnISO8oAP7opBY0fI2sy1wFIXel2cpC1t2ZevoM1Ni7TOS/nlhYIXOZLE
eH9IDGhjylEe6o9a7hwTuY+yjDFxlMSTWLi5/3PPVrf5oGvkflu1ufVZnL7f1m6itFA8rXe0LATE
ksbsktG3ntax7GMkG1LZZ4MGfIUDOH8MX8pBb8+vSlkqnRh93C5j/ePRrk8Qts6Af5dALAj+myFB
CyIgZq+SyW2kH9OtOaPkkccJZ5XkgIGMWAOBjsjeRRvh6AJVLPjzeP9QG3me260uM42lHWvJ6ahN
2LFRU/VLJwO+PfLFtmvZ2DTF+S+v4V1AMzMbR8w3yviTVAcwm968yDrUy9Mja9GtkrnICvtT6gYx
tpUkkhFCAjukbIjk7ywVZluXOpPNVkzzkCUx+jSsZZTSFCkRHpzFYWfNrc7VxB3Pa4/FDzHD2HAj
SF3fP7shzofLT8yyfcaqcLYlnuZ+VNgPFRjQ40WnNGudjUQvdzB1mfxktyUKSN6gW0Ew3o6pdyPd
VagZof6CmjXzqk7RFnfGA6KuTMfeaJvY8FGpiEA1l1yOpjvtjV9LvajAU+fqDrZzsu8ntniSlRuh
7Fli/RGLiQv6OLOX7U1C6JXMBIMvGBlqDHULddDxeX/p3+Ux62ZLm2RO/RZZAPT9Sk2JX+aOcQtD
13A6ekhnoM2fpChJyr47eYg30EKUTcR+9rC5393P7ParzIUqFGb+aMqWOacSw2yDqpwDHPk5goZW
dKc4cQfWF9eqpI9jNM8GJQf5sXse5e6pM5drI5hHwllhNJSlEkHP20zTdiENS9juKe2taIDiHhCm
CIz0lPRi4xHRYLiXCmbx7u5RblQljmafUzfzaeUMlxdHy50UPeBs4hN/GLbYoGRTRWuTJlKe0qhc
GZUFeAMvUq5Qy4PAey7UKI8Xs8ksDUIUUvTkubwC/m6b2ErA6jCUXgL8ghM9+sdSZ7EAr9lRDYdh
GSmvRMIKLmEKsi7f4BknOk2qRUaOICT8d8UmC21YwrKSn3mHemN3vWzznamsvHZEALlWOG3zXo+/
J2ODVRiHTTDrqT+um57+zV9JNoYFU0SsdzOC99CV5B7TD9NpjJ7IGwuGQy2haJINfKh7W403Hzry
KeclMFM5t7RvB9CxE2TqFDcch1ZL19KNwhIqoekeHO4FzaLrAkAFyZzwWGXsfoFE0mjOAvFZFX4O
/x+XVjhNhKcJkMtXNepMyRDq5jR3d2C/dkA961DDmu8r3GG6qD4WCl5YIfii4rpO6H/KCGPecXdd
MBj8mbD1BujHAL2Xk7QgzpvlP0aQ7iHZev4Z5bZ49ePiHyYYGUeX+EVyNlvQw3o0IZkWo+YcUgRK
JMWRDJSHzyx8J5wjDiKkg1NgnbwF0gO387/LrBaBBBGZz7tD7MsR36yd/dLe5z7GGOuPbOO5+OX3
rl2Yx3r3Q9QHUi/CGZT/dr1YdzWZLowML1wZfLjh0dmGpZdhES7Z6oF/9ToPVuv8ya3fKghwOoWI
p7TZ7/00QX76WnLhyI/OL/hHpG2bEh8ePqxHPLlcVwnrQITZQ5/NjabiTKR6SznmbNx95iUbMB17
O2vYAgHoj0Xtn81IG4bmpoFfS/BB8KnlkhFq3diIjAVJpISFUx1mZe61aB2WcsjAl23yxkpzpqSU
5zcKfsMeljFgMBfzVy+gJWQhroj/xa281mT1UyMcetiueCwkFZLCJlsiQKs4Gmfkk30lvhjzRzsF
8zqtCBuOUe208s/7yZGWeSGUaCjbTPkqYH+mHaBAJglv9MhfE9Fw7Z2ZhpXf5p7YCMdBrzIqTJkW
GUQ9UkOCewQGRkJD4Fe2PxTH/2gjGr68VATdFcS161TMS+0+DXYSl3cKSzNAhWe4pQMyKL5iz//K
NRnwQ0q8lQxQy6JBvQfw/e9Mf4Jgt96qEk+KdDc/0nUwppJTdxtHP0cR2e5qhEgABoeJjiqNN2qG
jFuusXItIZ7qrbBhzBDheQEH+LdQoqCiirsWdnNlrYDcm3okF7uN31rN6KYx6ZIcUffE8QSnUsSn
cU4cgy58vOC1koznEa2x67bJxtvf2w44Tf/a+hWWfZWyrLoNmy2Pz4+emNxL4hU/7dh7iygXs0E2
ghzBN3m6Pjd8chj1MQvaezuUd7LuE96VFh67iGQdKqiEI4YaPibzZrzVfU3koVzEHxNLPnSjN2Lf
pObEAwePPU4gqXBS92rvKQbMxooj7svMoQE1r/itRgsVSvlWcJWMA2ui6Zj43WEvyLYQaCgmRTHo
+irDS2NPW/dhP2C9wb4sWDubL1I2XE/pmP4uD64S9eeDfSolzdfTkMTVNTuvgpFaFTeM0OQ5kw+g
njtFE4EXHPWbi47yP0yENMbTFgXJKgISpuaCweexbGTwJMnDKeB6cN24zxZiz8fYsX3JY86VdQAZ
Lo0jlwzmForW29xESFvfreke5654PCtomoR1H+6P9xunA0XJTBEazoCWUz/1GBZyULcj1nbFEeWo
g69fb/WF5puygp5xNFs/2VFiBs+7YlpgwRNJLBtrXL8vlfhIoahana6EgOxMNIy97GBnBVmqCOFf
AMcPWgO/rlF5U+J2A84fA+eww23cojvLo3o5uMfkArUuUfF3Rn9Hw8kl1TONqaPSMAXMR4EpgqTL
kD0Slp8fZi49IunFGj3PzAi5Rd+6ebObsDSCjGIlJ7aJTMcnW7Vjtx/warTA2amPHVFhLUDpS76N
CxsD4QYD4XKUL2KdH2QunIrbz+F8wOwZQ24VneYVKbUvW12RStiRcV6JoHUABD2T6wBsWj7iz0A6
OZVhi9Co0J/78D6QvpnccTnLYSFkADI0mdeQB2SPAQN4xbJLQuewgG3RSFRiLikkFihbA7tsqaxI
sgrFBtcZUJ5Jg9McrQFBrdxYzvCN1zpeBRzecjxoYl55ItFKoh0z0VC6ucpDyFxtemWIk+Y2rDwx
2vQTODEyayd97kcgxy/av9T2XDOuVtlP56PS2FaBEKVWL22qkkBUkE+A6920gyJSCJQ45auwvoMP
5cgNkg/7lGFaSttS7omVV0V4A1B2NANTttKdjruhuaLe8YHMHIcMF04nOOOr+ZWffQ0pZwfqTC98
1cw9fqLLYkiHz0EpDwn2vqKFMb5OMgjSo+38zs6Yc0iz+F1wCvBCimlqxg1/uQtluda+y+I7Pq6k
v9/1KtF2Iq+91eVG/93OzZue9o2wCxTu/kM1C0pZv/TPxtCfeNTa11Nsu5Aix0x2ZsEFZZE3pBCv
qHRPrkMeQh4u8uocSoxSpg0Y2lBcfe46jT4xPslKLsw5oR8a28HYh6DJPRMbj4aVExTET2rLDer8
TRbCg2n1t782t7HNI0MJB6r4PD/pz7KVdQWqyEucXkKJNwnnRVzTuS8qYgD4TRa3Hz+8EhINdzZf
ehEO2Z+77FOMu31/lxTYwV5+BkSanY8bN6tHFOjhsMWkNWYWwn0yOekUTg63Xn63Uj0JVvzpwJ8h
g/tCDseof+WuwzKf2jPUKnr+kk7hLqwprDmK5XsF8/Ri2Ao374zAj3q9J6WVxhx51ExRiVOyfm9q
ViuHMTPAfN5XVRyDal758aEBOfXWteeFqyVgxJGSQx8B1xrOjVjYRLPMk55iwUrZ9zHuyKcWy5lM
T90qL+Sa+ij/AFGj8r0M8YCzRdhWaEoY7VuHh6xH3QTQkMKsrOpQK6NTIDjnjjIR5zUYOBPI3mM4
EH6gCFpkx9VI9nGHEXU40+bBv8IAiOj71G9xj/zKOQjSmGeRD5979pgwB7GHd1AoF8dmAZLc3feh
w9C8XDovjPou2wsc/e+eos0WUPQYth6/xpHJJw6KiJBrckg3QgTBdXhT+581NLyH2B+xg4ujs7uI
h/S1a5iaNd5U5PwHbdxardGP9f0rXRtrJtvaOQdTyNMsuXAJGkqhHb6Ww4BFSNJUsFM5fi6E0CfW
W5BByWEelcNpmU7m/CdvnzvqLszgG4CaYu6C7MdY94pr0tBFWn/jUizraFtUx/NFG3apZqyQsVft
bcmES3PKNjLGL3ylszNtmfDCcW3zCQxz/+Eta8600XMHLdyneAXtdPXmgFTfY1MaAOYaNIltIqtl
AF3X2rC3nAD2XL4QEa8H70o6VhdNKeYri98Svl8ycoqCBw0gGKlLuxpCY2/U7jzYXT1lzgLrEZsD
/4EDljwkVpcuJRofoLqHS2u19evjFiGOJJKD8GuJDIKgJDok7jyxwo0lkBDRK9TW0CqHVgOWg4EA
0qGlljUMMUuZU3tRZXGuK2Y5qtSVBu+t6ARi/x+XlizAH3O0hW0yr3UNBgLDAH3OvqR0e+A7TEYo
bcJLxMlrUdzZZK664gOT1NUysuM4nsCox1ZbVWdpQDn6Nnudzk4pw5jE1eybbkqG1HsOQEK4NhHI
1HCT4RFSChBhE2GPWWQ6WfY42mruXEqxR+nA6AGteyZMxIv8XhWkhiiWh3wjs/10vgNjEiB2qsH5
Vkwb9lzKOxiNIvmEvON9WD+R9vlfh4mcZv+Q5+bKsAjE0dDiMhx0RQBLdBAKC+cZyDGRYnoDiLzk
OyIstpoNZDyNd3iIRDe6aP3QGsRo0o2NxIF3xW6hsvKvORgkcLpx+zQx+LXbGNqnGQSqEws1N7qs
q692bv4+4nKdwe/GMuP9L7Pl0mIYgRqF+K7sANaJE+7d3x/JE3AXwMjG6DvSffgoI+aiz0qmpuem
YNt7b+2UXs345CiryOJ+mszari/SZAn/oP/kudrN7Wui3VcobIfTY6kB4e65cPrTxpltQ8cxYIvh
tAzJndRLpgjxNCF83XCoDg/3bdbTY38xYsSaEJlM+IJv2W8Cd7MoOD5drxSATI/Al9fPbzbATnVN
rsH9TpyCRzY9Vfqhpfw2I7SP7MODJ7tz041qHES4O0GU1i3U0NXYL22j/X8TSsmVR6HkKwnAqInj
OVLVcYXHnWXfUopSnBcj/NJf6s1iVVmIWBGLKoRLKoPNIhIKcMi26BHaIk8JF/ZgMEDAEyuX5bKN
oNakRDxc/hKK8uhQVEs1YQOAkPO/M+1dOCrRhFc/Z9+OZGvXurmLyveXBEr4VOR2oqGP/kWAVyC7
KndUj3cFiv+htpl1meKxP+DGGKu7MtKUGIwIgtoQdW+AgS7Zl3pBDurvIzpk2fs7ZaKjgKLHmCtV
rIVGbJgXjt76v7sHm7zk5dN1Vapo2caNSZQ1hxaV/2FHXr6y5RiQLvRgqYu0O/ollKhkZ7tTwgCF
6MzQXKa8VpW4rNWUzwE+spWcJLfBB8HySlmCnu8sOZbwFtoUbyI2JTtQZyzbyFVOhMnLU62O/wxU
GyKOqkH4y107ei72rL0pIYrKun/4LdzEjGWZKRjd9WO0YCjLzjP4bDOaKydD2LW/tpsBogIWx8tO
lTVMHYJCBhMYdF3BO9v6AuPC/30Kj0+BW8AiqkcKxIkvHiXQzUtcOWV9LDcMUGAS9B1UDO05yEtu
2lFcpcGswCZyF/Co1/ydjBYPnz/GZkEGS0jQtD8QT5G98RuDiVBfIhGNATdMucnZ8EmgbxluLIKN
3eOzB42bgmWjLHfS0F5noxi7i0fGUTxFwWyR/f6Nf3od3yeTIc2MQEafvIinMf5JOsERlUluyMFR
867WlCnT34+FutJS5/brLXqEKaB5MEBU+whBFD7cWpqUIhGElW7adx4cGvFX3ctjsjF45mYdkJNJ
JbcbEVQZBEeNvsmWGqrWlkKKRwPJn9RhyqXSSkaIrKqvN26SslH+yFXHN7wwsLjJPkR1dVn1i4aA
2VeLnJD32VfgCEYhBxlSBX/QRsEJkGLuUscR7AMKvYdsp+Brogfsjop3nZMAmPYJJtiXEwOKeVwq
uLoaVCi3UDjmEx1XzR3D7kcjeXyLb4oyuZWvCb2VGyJFSLC3I+I2Ldr2EaGyQaYOGR2lOOh1oCTy
3RHDuXvn0NT83xIlDI3Y3ybVHLpxwKYozLizSRSMyUKIp6iRNmx32Zfbactr64IHn+U6tFrrnJa0
Gbit+LlZQuOlnc89WDh8otSH3C15B5vbGgU5FuLb4BUxWGy8cpdcn/xgvLgRQSvJmSxUamI1nS3f
G4EUnrAFaazSGux17fvYW/P73Rr3boqvR9e7N9TvXII93jgBzYqJw63xMJcbCRq+HBM2EqwOSJRy
1ip/8LgAUvnKzUCYAmOcmQ5UIa4Vn1JM6P3QJy5oLBJP1AZN3ZGz/KVNrgHIFVoE6nZQkP+6OgbJ
gAq/yh0i6Y/MTKmnsYntOQNY76Ksrmg5qoScgU9FnabpT1BnO+Lu3jR8myPckYW7mlnrRXIWbdt9
fBhR/cgWr/ke/UOhsPeHUzcASyU2gM11o7QSN3yp3ulaO+ifHKmpI9py2SoG9qj72ARbBW8qX5dZ
ndhNbYH+Qk/wRZnPEL4kKiUBGYF0uVPEqG+o5zLCbfBywkMHlo9WjnXKHPhh0u+jxQHIa5IJeQ/t
OWCBnRlFSykxZQ+YvTpneIPAb/bG132WgeMmUOQaUGgSczOZ9TQks9ZqDj5fmaQsa+lxqSMt21Km
OsV6oBpGdF7fZ11utbjKHTB0/3/QWhTIeNqhTNIES+iRhmx4glr8CtJikqgBKmaTQnbJMv8CDR+s
0Zgg6iphov2hZD4nLbbze7eLQvtuO7OdgFAW5Y8pZ0UcU7aEkDjD/DeTI/a1UMoTndHIue6xz8/M
1H3DZ9C+XqkZt8tXVewk8CGqueUM4P8y9XueMZVhObtAIetuJFA6hILg0ABmUnUYmfKnQfzirg9u
6IYgmUP4X8dOK72Rq5XDI/MOD7bTeBGajMm6W1U/oS/IRbJ2EnohQq/tokxtP8x3mfYR3ZFYY1Ty
KrWk0YK0hD2R7GfqyOpFo7jHqJQ0MeYlgD6Nupd77POBNjDFzc3nlp6+rHkNXb4lEiwydX8y6ajC
Pyqe+WMsVlf+ykg4Wx8JQ3Ym+LN0EbmnZMDUA6zTxOPhtRlTh4mGl9p6bHTSRA32W9ouJY2b78MI
jTS/zrDM5A6+lWtUyZ3LxtKW9JOrRuK3rv7Yhsi9cS45197uIA2UOhGIugg/aIFRVTpiC3tesyr5
QdYi5LZlKaV1gNFNOXk4LA+nfZTa8gDeGOJzcq3cIVok5LjtPbFjCWfLtTBflOaGeZMDtAnMAn8s
o1CcnQaEaAzyKHtvge5Wpkj0lYs/dPM+YsXYXJyG7AN8UQYWKiciZrO7VnVN+GDXQq51/2LrGhvT
uLBfnwcw300yqJTaV23AEQbG0V7fnQk1hFQwm3Rp9BrGCTqXfhtPph4GHeyTG58Y4rZr7j2az9tW
GevRmV0IoD/CLvJBB2fEAFWf0T1xbnaJYEwW6bVTTx1XKLjTliNnCo7EHbmX81MW54UzXn616XXm
nw/NWxvWtsDZP7geYtCO0OvJBOguadlGDffohJB0bDvDcl6zCHJao5w/Q+fX11K4o3gDU0NTd3xa
SgcakhalmPu2+l7UgHC3hjo6Kn5CvnImilJhwSwJ+71R7gzQK78dUmre0UsnD8WKVtiPKUV52PeE
UIrVdzpLJw+vbRRPVZMrtYhZikYoxc7UNM3k30wN808GbmWqQ1OkTMVkRxLkcuXSEM+LUtpD+jUx
rI7grJfkyIv0SJ9vn4CbKDDsfYrrJudM4AnJKkYzfozlP1dCHHUby6yHypKFoEXrj3cHHYBEEKKY
j4+CSdv+Xc2d09BHlCZeaPxF41hk1ClaS4s0xY8ZfVLm1aCLDnkxV1Q8A8DsoztJPg+bStpNCH8w
MYs427AKZcCINg9r2+/8wNocECwYmdLLG+fN4iSEg3ng6lRKvUXuX+Nda2mpgAUdt/U43Rh54jrf
Zo91RmDFoskmL3ENarw+TXEoz8PY1XjmlLcK+tSkyk78YnRRbKxdHZtn/AP2pdXy8itWyaIAgdBc
7JyezNic/ZMdm/RtYiceiXWSrDN1nmJXisVrKwtVM280pyPFkhkcPfkvUutXzrAAgc8UfvOJoGkv
CFkR1gTXMSuf5vVBB6AayGc01OG/qFUbLgL/dLi2oH2//twGw55hQCjT8XE6Ybni6P+T1FZVxQw8
7HWeGJE7xU6P8oBCpj54X4eCZ8cBnc88XeSvc/Tb2mO+vIhgOF0zMX1P5RLgn1z/xs5k+Kezp5p8
77IihOdj2QVFkyWoe4FfUKjBWR8dJlyPquXCi/YIVjxqywzIbYtOorcKa5BbwG+RnDJfwAOzRXs7
D6Ee2SL/dCzTVrImbELRP0YPPdB8Qp2wl5XN1GF1l6nuvhQhSz4QHaOeJIXYfpIoBJF1KVArS78K
lB8eeEjcLEdkckDKAFz7HNW/hb3gxtmeQg5LuhEl9CKJ5z5jU4nhdy250A8/oE0Hd+c1na2JNm5u
DcxuX/ygiBDkF4u5n0SbOX74KlQ/+bxe1ZZ77722psHHjUhuwJtAAycM3R2/OefIco7GUP7hHBLY
KuggyCYMQdjwLKTX9tIiBREq1sCJOPyYs2qkLAj+z1aivSF13ckdv78SnhC6BSdW32+iwdqzZsKy
TA6RitO3D1Lxq8g/kGbzqEC5BOke76Vh2jfLjRDfy9DYYNSX4mV57S+zrjQRH5AsuvAgOCTv2HPp
u8ecY4PQy26zapz5Q+LIVCaKOz+cNYmyAS4YTTVBQ/EMpEIRXLGu++6tqr06W60NvQKTcJDHCr/c
bLxkSI4A/fdBUGC6SyKHa5X41epRVC/PrIhrp5vYqthhNJRM10Lu/ANxj1SF8ROr5wdlu/fDDzCX
HpdRiCcByCuSiwJM9JHxuhq1XEQ8qqvtqa5POgE6iubY/aLhHUStOs5CYBa2OxEK3K2wpESmzHSb
9xP4icZmZ55DRFep76CoU0gzIhIJWOGio26aKKs7Cul4B2Fun776bOmOZNjRa0YtKb1OkCoAuUM/
XQwBqYHk7NiRqbXF1PgvG38fBXdRK0W+n/Lo5tUDig5CM4t8IOQHTNXWuiwDCCe733/iTwnlowVV
BSo/7dMqGgXHxpje6JrTKgtUuS5GD810aeZS+p5roshfjMuq67bdwbDN41+a86WrpQipEuSaae/r
4Mwm4c5Bau+c139OK608H+CRU2MHO7oTjKtOeFcurv4aLlNVbTTLNa9qQWBpnbX6n90kVJ0RxeOA
t8Q3461f6szLqrmR5bS1QbMQoDJ2J76VyhZ9Kp0+54PmmDU2pK5K9V/WNu8nNdcKRiYn1/MPrfpX
485Y5m0FeFHaPesUHjCM72/pdcb+KHhy5SDyyOCIoztoH/Xd3Hy2VUtM2ae+Df/VMWj5QJhd1QdS
OlbNWQH07SSy18ZiYzo/TAuE/3wnO1wwYeePYgTdCGhyD6nGG9mt3SdPlmYZH/lAH7TmX4JQhOpw
CZ7fxCFwYKvQ+dWQ43fkWmKS58IY0QOyZXB9CEtvHHarfVt4UntUfhUKarh5XwE6CV3mbUDJgNTQ
RiW3rzu+UDhFU4hOg1R/8/QjqeB29rQrmJv7Wj2Gly7cCrGIT+IZ+dKMJMtNdFUFaraLmehXSffQ
M01eS0fjW38g5paKQ4MHbpf2fg6INi5o16ocTriPgkr2JPHHilGESffuGkvrrcdXI1BQc8cRDkYg
YzNAG/QnK1OrKdTQHOu6ioj52+7p15LxucGUsJx9zG3mj0p2nrxijDs7wWKFsd1oBFmfnkth3zNk
vQqurUHUXlO2EImfXrcM3wQvVbxk8pNc3p9DoX58HNdon5v3YYH3GNF54vNRFKkQMIveWzabk8un
/V69dczVbL0CuMiBxobzu4mDUYIPb2DMx2rYiMXX3spE3JDNnJz6cEzTpN5aXgeqskbqCd6NsW59
gUAoUwZN9YJq3u3di92RMfF7kL4FMsBXFUe+ywN8yGwpYrNLS3TaFJyCodOmvBwaHsjja1MoCuvX
ikwENQh1/LeQ3BCBaJa0jP0tHW6Yt4A/zWPx/1IVxtUBltJh5f1ApBgkhtE1H2X0ePiCwXbRXo0s
anb1j7IKwm6blhvH6KD4FezJZ4tBW+vxEibJyyxuuGb1H5r90gZ+8ietQIA6iTOuJ5z3Qrri+P+t
4y4Ad1cidM+LChlx6vG4DhttaBoUgcNN02lS1zLyiBm6rhV6VkCQatXtTpLsOBZhUmNExp6dJrUe
d14HtxUdBTeAl+0Vc6WvjZdGiRjyO1apm77UnzH6FwrzQHiDW3EqznsNQmM51b3Ex1meXZafHybH
Mrb4a3OQPRJ/v9EJAcqUyEH/had7Cu/ngdRPOHoY5O20aCjIg7wxgRLlipcHzI6NDGzbVel2IBtn
JfBxdof2Rih2sANoNIIihRHimQXNxqZ8QfZtS5akCwPBvXrZS45Qhug4ialOti1/0vMjRmUNoA7s
JQTpPQYroXpxNqG5jWCIC9I8pfYIIwMzYHbZq8ZmOS+/u37tCkYrnHhKCNlggtFoB2agr9wfbY9t
lAVPSxqTn6AfytFFEUCiMAI52AnXTlyT1iEQTFgRzr0irP+SZ5Atilea2QBFlulrN7Op2/xP4cTs
C9aojGgGy5Gpk75cw8gaSnjc67GStvw+GSyzUSvEHcO5Z0YIa7jcqaI9TFuyrjfroOC+WmbgIaiI
uqQIFsqSzwinSQJ5GUs16sPcjmgeRH/koRrXpvL126mHt/KBN+v34tAvreTRHjo1/MVTk4yD0F4G
ikRFClCSV2A+OGjK9P9XRPnrl+RDG5ro/GUpafDpgqEKuGBpz4F7HgH9KJ4l6BccYzON9Lsp2sS1
58JiQyX7F269Ig63zbnlVd2q1WdcbyXLwbA0njcvVSJp8myVsiCkiL23ZQW6rTcZ5n16sfzCJd2n
11ZsGWNMA/OHdHcJB+m+TBAWnwXIP0Ae06cUh3SLAI5Ia9cwHxMn2JOv0XD5v2yr9P27CioVIOjQ
ZFNW6ShfhQsg+GEwz7BGHreuZaAKpzpo7CbvND3TY5KUMaMpfXV0Tc7LeLvn4Z24UMqroao935sn
UIQW45NnHc1h2PzJ0iXObwzvQbCIYAy+REAgc2rxQwP+DfMz7+MXcEJ9GwQmctHtUzrirPPWtAJB
hKilepwcrF1NVjzLqdWm5aVvl8Ho0DRQpFqy193a1N4W2c5o3N1lkP8ArwjbOC/JCLETSdqcI9S4
p/Nm+esra6gyyCTf1ltcg5YV6vxpO+CTwmYAvoJRJRdeaxJaVEpPuUxYFYg98Y+3j9I31Pp+XRxH
tGZ31Qg1C9u75khZuMo/Iu74NnNLaYOxay4khGhfCyHk6IjP633KfRTT6OzQq6Ws78CuXjb2+YfB
bq8CAHs7UhhKzEuxUrZCWqY61nCclw2PnsPKSzjECBr44qjN51A8ySRQv6zj4dMfj83YmyyWBlu4
tQvGUqH0K/lprhE82WSZxEpmKpWQYovzA4ZEyTAp83UbVqT9cyndty5zFobTJWrAwjg8NY7YYfDw
4OeZ74MfN1wLoPvYZAhd2d3ByT6VBbaqWjaQ77IMyr4RRH+99fJcCjN+0lpzoRje6MSygyTY/OqZ
v38cP2N0cLj8/bvqwf8ShcPIfAoXtCuCZTPOP1it1LhP8eZA8g/JsKGm/qbvOm2zSwV7xVutrjiN
73Ag74nswwnB7kytwFg+440MAtnJT5QXva50oWOv35UDQzNXvPvE5z0+wQoezKF9BA0B/4KzlUSS
+e+/Jmbb6vNqnq4PecE7hReX1ORpTZJrC+XyYyCL/XzELM0eTwcKemhr3cqJLq/WDAiHFdv1QsNx
zTNaSPsMVkeveMQhkN2gscYNKyPASYaWiMbJJrvwVyY1CH2J/TL2n99/nitTgmVBHCdWYzoEyKFi
bA2ti5BQ8lKm0Qdc06wXKdP+Ozn2WyywKbjdVmLAEJEKy9BP71h/YtRRE98S5XI8Jx4LNVcUnq5d
FGZ4Jb4/ykmVvsWkFOA1PURSd1WUkapHIDbUNP9XB3PA3jNCExC8BKJPy1nZNY2MYQYFzVK2+tem
dJFTgz2gcMP1seZ8X/RspmqhklHCT/6mttPvigSpOEOO6NQKdChdmqQ+D516qis06H75lseoS46h
L+kMJK825PyBqktdWW8jltE76lGK/ywM8uif08WSv4tkobvQV4+aruvj0IMZTlopPYkJLkGHH30M
L/Ygzutnt68E3xgFgUMh+3pDQe7dKbUMYHhA5QeMi7r5YuqXooVszXvgrBNvEIRnLme/6hvdSpxS
CoUP1ns4IaBlvoIyspJX/DCH/A3G6owAdQIeaocNfEMaCwhFGVBuAuXGKYvscfSnR+GBpzCNjwmB
ddLwWAYf+5GuKaaOxfLPU/30sSI8ExwXui1oYvu49b6q8QVkOmVSBn9w6cBtPrKYr9+vD3jWP1/5
0vBqGL8qLyxp0qywc9Xa/xuWGPKU3Ta/iQobE55UzeVvbIaglNPRv0rBzLrIlA95qXGDUCdYTIdW
mL4kjM+8wdLa671V0hnXHRDpzDQVjRjgGgX3sQN7DCObHyAxJ/TCOG2lJTm7nNG//hcDUXzZK00H
hYCb3n2PnF410vdhPTAOx3aKMw+KYw4T2hXogXRyMwtWDuJ2TVlHA3fj4mhaZBnsmgdCf+6lBt4J
6E/rvJcCwGAh58EVtarPaKupwRFL9nm0a834594e7snUgda5ZuNjMQYTWwgUeUpRvnx/Ad4k4zhO
dDfvAXOmUHd56r9RDPR3OatoI1WGPi7kQ1DkHm2NrAd8E6OHxvnCQ9Yr1sa1s1mxrTk6gG3i+W48
Xev+e0knSWD38ilBKX6HxpATX6Y57Ullxqr0FrDWYb3vFahM5QvphZW4IhvKK7nxEONoTDRXEHdK
6BHHIirV1WLstjnk+VzwksNueDwCQnMdLvEve6mo/BKcC/ipVbM4huxC8nOYqvQjJy2FlAq4Tcnj
9FgsdFfG/JzUmfcej6+ljxqpeegrswo3pbkodCOG9Mw3JEO4JnHclChI5BhIHiXYp9UWPWxg8yW3
wl9x3KGkJIgzlz/7aXRRoHptOzy5sW7BpZuufwM/ibL9bQufNT0emir2GuMp9Ar+bogS/kZXJNgZ
IhzGzlPTX7zENO4CzHCtj4wRqIxsWXUvQkTJ/uO0Zp10SAKTugE4tKVe//DsUi4ByfACWZKcbL35
h4MrD9WxBLcwbW61Qrsy4Op7EZgd8iXq4N//U1wJ+CEaogRRsBP7JzY/A/cBWHgG6eFFTBdbki9U
dvMKzgxvXAik+p3qojZ+zYa+xVrdGShadFsnJ4K0LIQUX8x6ebrwNb4hK+Sw7PVntrp7UVDTEtCP
2DfVlT4k1ksBOgeZnWGKbY6LJbtiHudIUgc15pNwdj98zpRSTlVmP2K+VofbHy/hqlZRFLUNszQt
vaXW+dhpvL4Btkvh9TB1nexNDoNtwNIwXYyFducxhTWMPbzFdcYH+aoQb50ZtpOb2gaclyj69/0n
709fIgITNlOH0i/AkQHMu5jp9mu3Hs0TW6llaQ2he2Kq3Ictw7qqc231OmW+CnJzj+dHJIZ+Nmek
q7BWvoioI93g/cpchU2sTLyIKqZyT9gLbMh0syy4MyAqZeXQfLDSUwPjZywVnWADolJt6Rmi0tNo
+80FrE/avmhrmNZFD9B40sR2cgmL17uUVQtQ9B+XPYFvLtQbM6JfxAOacIIFcwN8ir4bnQxDDS0C
/xrGBSJXxNl3sR7hvpcHZwofBdpMxKakuIbKpctBeIF7vsBB29exPRM0dmjljlIJ0AzJ6yZyCPXk
jZ0l3whqMBPyjPJqvSTyR/lqx8U0JeF71t+HeZGnpN9szcKJjP9QFCNKMs3hmDz4Y02NBYpzjU1S
5U9Urec57dBeJtEeM+tRlwz7ACf1pX+cMJ1G0ahl3h0TKg1xC0FjmHXP/KjnMjqAnoZH/itSiyxW
BzFq9dfM/W/GLRGjqI/pOGXcb9GJ3QeBPftu5Dkl1hCtSWF+T315VlyQoPboSRC4LW3TQU1WRDb1
Xk1MFxmOhBjAEUTZhrBiIeN8xPg+j1B9NIC/1O3uVnS+b3fUkg7Q9N0e9Lw9lQHGzUJ26JrMHiKb
eY0LyTuW49fNHV8PgV7vkZkVQJcGjzq1UFrhm9DWbPZNHvGWsJ3MOx0YypJtqXrJutq1MtknjWpm
H2B5jTwXtkSeu/GNQxla2mKJ0+zs0PdTVbeKqxFiVWJxKNyWFCRmsBLhEuweqgmnAQUTEg6I0QJt
OywyuxE0cmA6iJeA8evnaWpPh91mRiPeevN+yDSpNeFAXv2qAgHCDBiKNIx3mNd0xH0BJxybB9Ui
Zm6Wxp87tuHk5B51t6NVJZUksqdpgRT3zy4ieg+pcYwX7rsi52M7lJQP+w7l+6+TJrttkACythAQ
FOrdyjBF/q/LZNYSfucfMAW8hI9ZKM2vjl+U37Sbokr7wCTxEwIiNd487K4COAyXD/sfDJRJIHMv
isOY8tdn2HnmjZTzDwoN1igOYfzrO2YLQOEob79qwG6egOOWdjHAPwmxBQuYSA4k9v6iZVfCfl8n
/0hml6fmib8SqNi1azdDzHzyCYNkaykRppwFqHGoPYNTZqWd7iYbk6YBFxWjnYtUoFEq+hznCeBM
pqNZo7KBM4fvn18L+Y7rdvmmc/ou1gFwX6Boamy8Xk8N1ZUYEA0Zt6e7oDdFIVUmrIAiINvDlAQn
KAV1rf+vCw1gn5ju7sEmh+vGJ7l6dw4UrDrfe232XObje4n9b6i6bAibhFMzSzxLNS2SKWDRMEtb
myTkjnEooOJDh5/2zRU/E3vjr/TVc5iTlxBu0i1bx4wbmgm2AEgjoGU23+fNS3I9YG7CluEMiZEV
gKysnap1zVSGI2AXtPXMp/pc+hdZGVHMRSgVwhaFQ7PdOUeXp4qRjspb/i8h1aA9eJ7IZl2EZyXR
21b3NaIz4Emflo9rq0kqFORAon/XxGHjdFjFHHwTGBvfkmaH6D7t72yvMRi7fII9dKjaosKr4Z0n
Ks+gwm+WdzX7vXFjVdpQjpMBhOqGP9vP22KsMhAfiMRZ+fISnzqFHygB8hGUHjGyGTVd4Riuu9P8
UJevuBZASIyfS3Y8+gAelmIMmMwfoPXjFEcspGtuhWyOw0QWcIn1gjK2pk0tzgZDpHj9kYDic10x
Ti1OdfHjFH65yGgbx06uDiYSS9sJ17XZP4TMEJriS1p9CsBhK7ox7+FmO8/N7IOJQytM7L/37sUs
PBpx8rl4PIuvsPIYGBqmAo6bL2zIFAcXyGJusqKTABcxyx9N/xnTDicf8iTJlEn88V2Iy1kzhZD5
05hjlE2wHXmWrl0bfwQcbD3FIo4tknVvjNSTgNy3C01kF3ANhY1qopOJrKcFGiUwZYYx6p24B5Ls
RGpS3Fx0sCxymuhjB8TuRqZGkONA4uZyPS5M+601/VpknY9N8YVaUjBHxdKLHNKXGRKu+3JG+ARE
b2KipeYaUw+F8UkKOUvt4SCnZmItVIzKRvGzUaqHB+yqxNwflmtjs32Cv6by9fsG7zwlrfk1LO86
xhZ17qbGXjbBuU71VwIvHTuXjeDsjrhZ+LiFRNv/PED97HsC1dLQbX5bpuS6utQI25v6YtvWtoPF
HsLEpcm6XvELv1JZVv3p8VPZ811qj1kCyskOcRCE6NRYKUpWDp1h+uRrwC6GUzcNNzmBUokB+mCD
OYBAohP9JP/cZ8SyU8RxVd8WZUUr6vGxuKAdkvY2BO6fFUpT6ou97mQv14bHpHc4Xh0spkV/Xp9J
FTMBKWqywPpTtaNQ/jEBvaSoiYrhPf/jn+kDqGvPywrn47OQEDr0XrKDIkjk3xa9lZim03HrEq5U
+L82KmprBPzNEhYogRJcrzrEGS8YEhVUTy9fLKXqFMy118ldS4XE0EqjFk0KiD7jbg+T0dn1nFWf
k2hvIS4VUxPo4N9KQJsJmmqceJBM4bz/MTEQUFdFZOdL9OL4aHBTFhMIFGYvqrP/YFuR1Mfve+0+
vtRvc+v3TejCTb3CsL/vRP1PTyN48RvriE5VLlBI3x++P1T0QTzez4R2DuMDqjBCq7hcTHF7x0QR
r5EDs9+YPFfx7QXMkNKYAHDpbzpDKI4agVpgB7z2f4d0Aft7sfSOuz3CwoBaZ3Wz1nnG3OhEYF5y
jEkvAxGaWIWFeku+jOlM3e5pUhvshOW0t2y5E3mCY86UFmauadMriGhjzvlwcH2atUWPpyWm3nFv
E8Mw7r5RzoOQ7/4wA22Dr8jl6ZjjtqrcSLMOwBFHIKEumDUr2iuORCDvOwQQ0YTt6s8MbgFNUM3o
y45ccrm+s5OUWn2Ow7LfDtvxLPh5wJ6d4uSQcW7eFeHVaf2eK6oWvwgVm/6w+HS3XbkEv/CyPhef
XNPn4B/CPk2kSNgVJS0+2Evgk2uqQ3zCwsWA7uolbbOnUbQX+8uQ8617E/shCHV5QzPQAvZmJJiU
TtRpVUCdotUo3wL4qjlzJTTej8rwxZKgwjkD8EX9NPm/9SX8IasJNFFeUAakAxnZ6uvroDE05OKL
pbdeZVYScwu4ovXU485lk3kBI7uY88g650pkwUAjvztGi/xj60CZRQCatY6eiOZmKwFygtT11xII
lYT3OEQaZCg9VXTDvglEhL9Bzmm1rHz23BLgjuZRapIrjownnuPRsCT9Q5ASiRgsNdxp56NvclPO
pWViJV9bBUBsIxXhOsdHxkdOfVNiS1NaC/+5/CWDFaY1CsFL8lF0WLj2t71MJMtKCAxFxStkt6pA
Br/Cz3xgOb1Z3UIULbScZtMBMlC2D9s/P16IHRwKZIaxFO1NWUKYzrZ/LKpaMynQwOlWUWXpq0xD
7R588AQQ6j+q0okM944k2kGLgYmD2MukxlHWOxi3PKOoJH6SrgXWyVTTP00k5vi5S4RSJ/mOA8bW
BmHEEQnns8Gmft8KqebwtBOm/Zoxp4DZHA9bZqCBJiWKjJaadpAiFSbBIOILBGvKHoXKrJ0ygywr
AO7o0scJ4QrySTv0xRlDHcFWFKhnAZTrlQQiFynaOU5gz0wZAOVb1FL4NxsvrFSHp4ZCu950zWxw
WNDyV26HVQkKXROBX2krSaCtDsle1jAUYvknR3p+7yV6titFpsyzRJ6BDYBSrfmp3DAd5xXd4QGB
w1fsKAAhyS+8hg6lll3VfdWH4VV5eKNgCAxhX+UqJhxt2PuihiG/gW1T1UVxaNs8txo07lKSws6f
o7oH4v/PnsnKAhe4tix34WEjj/kshHLCA1ykvPwUt7ne/J5SSTshaWc9aV9E5X0Bjq9+etkCDJ0K
+qhc4OEn5ej/PQDN5MJAliXurl2cGyNY5YnMHQecKCYMIngY1Som7DJzr8qRqSA30gr8ZBrCNr52
CSEktd+pE/LiwgEzv3u9X0/8YTBbMfWHWSBUSyj/F1k/lLnKqVBHHJL8g+NVPMWytZGa1t4Eu6Lk
pqpBoKg1iJPYCnkLChqWP1W1Ogx7+ZEaboDdjDlBD3SvlF2XFRrQh6hVMuyIkM/vz/YLzqfgsQ+g
wiCz5rEt1kDG4nUrqTZ0sPwBgHjV6XIZqDxPeeophFCClW+zbqo5KJXBCHP8YKYTxCqpHmh9pj3o
h/9vzT8AC/2SEOoP+LIJ9PjKNvKC7ulSXDeh46y1UH8GRyCTU1xWfW+zFWyew/gIR2wDMvNCbEF0
WfUQj6Wuf0n9g959HMWwOLMpVKi5wq8ZSKmQ9u7N6arFznYAgsOU8YAoMc0EoL/gVi9F1o4W1lq9
yXuS4lZmtSd1qQPTT6SHtwqMw5CuwHt3+VpuC8YOqSVYhZVU13Kb/3bTsghwek9j1gzHCrx9Z+Fm
IFVcI/Nhcv36bnvxrprrYDXoChS3TkSXWPLAz94sO/yStZuFHHnXOp0hpc4qSZhxn6dACmk0jj25
03x0o5uHw+4PZEDTt7rjoXS8dF9dv2ZrpGrow1X75HnuFTu3O5BiSrO5Rc/gbock7g90+emBFSRc
yfxFC5cvw/vm4u7TZzarteb6KyVreZp7IPlI4fUSFMKG3y1w0r51JQ5BG+zUml1J6N1MWBXQdGzC
lv2GhXHYxa6TrWSj0Y8ifwIO4uNqrIrHDDBdW/PX5WWXbRIiexQd5gHyAG6I/W7HooelbDU7RaBZ
9WLohf+qvcKKNyIjpUwKsop0No8xK95hvn8Rb1+xCfz2OhV53E+gF5J1pzM4ukaKNoLYMYOp0QGq
ae6NMREK0UD0hYIeyvISCGuUwCNydp8mTAjc/qzkk1LwGKPzE2ZQB+S/El9le70klpWzcdZQHl2b
a5mG2PI4lIrwx3parzBs51opmR2lUxPI317mfioDeejKuqE7Z3GN3hbuctzEystV0fFagvV4p8FM
mH1eiNnh0tFnVZ7k01PVe7hN2wy5zTWVcvKKS5KfMePz6Qf8rBjjEqaxeJMjb+UseXV1XoEJn6Jt
SiCyFgujm23ea80tlucjCBlc2cKw8G6CP4Ndn3C9V/rqRXGJPcGy9dermFDQSRxGapryvfEc59gM
ERkk9pxvnhSWf3znyHkUkZtvpT2eUg52LCcdJouZBCGjclvSXtrWh1lQAPlo+IutMQmaSJ2tf4jX
zFJnpQkKlXUGNGvcHPpL1ozSRvZmbr5IwFC7GH46Oeqc9dpZ7uQkuhlckEIwGS2oEJ/tPf4wPuNT
jswwyDK1GID+3jGuiNg5IiM0M3ZjCNGoA9gTF5uM8RlSiLrHZ6gqFyTyUkiOcoPJ1Ojdudmv2uWF
RPwIQNLVAKqRjGQPQjda26i82N1bxVfmkzYinnzOUGQF3z1rm4Z6JTocXvJlGWB0p0k7WCiSG3OT
KLBNOxUWdEWvvfRcQt7D4qLponUOAerhNStMhXuxxpyUdlVGKERoivXQj7sg4X3CJ0IAgW9e7KfC
BCuzDjwArG94GarhJwdhEOAqYmG65I0MMi+J0J69MWEgCZ5yQY1Pxvxf3ZVswKxEDguV+N+hXiVR
MY9rHBy6IK2svirsDVtl1BFUPS63YZMXodiNUDLbsWXtC/eJiL/Wt3Wp/2ZL1QeAEb63qRjPezII
e07WFT+nbS8l+ClrYWlY9L8x3b+qa93/XMdNAJ/BM2XT4TVq6COfi3cEnvTgdd1+sFsz16HVR1f/
pBlxkG4QbpDO7zxpYCJm05j9pEoKFI8iRudOwWmKuurK3lHXVBB43GnNQoSduQnE8TVmKYAKwMoI
emMISTlrbkfTTIFMlqVQYmF37TTMEErNRQ18P/Zr8PFsHSdplCgDrVVLLINlfNkeTmLG1RzD/fYi
QrP7grE0LIk+5CF8uCWK3p+EVOCTra46Eg8O1e3ikHE0+JOWVAc/haxHjpXVO7zvrE44FH/9nR0L
ESiEIoji4EfB9Xn4CPDHDIrdK6NDu4zDqE30hsZmmMGivlh1VpIj6slRo1NBJ058r7wpWHDEENzR
AvNr5Sd+HAKk0jvGvI96/N2R2mhq73+C1Z9Ydcsho+ZKDGm2fUBtsEWB9Zwnv2uD54F7a92FOQ6B
px9hwwMMFl6ls2EiwKp0Sa4xPsRD7K6DINGQWPyZd1FGNCHSXX21fK7hCPlwx4P47yo3gsH/UCU4
dEbdtI+9gfR8XXYMETO2grj6AHUM/5Xo6pPdHEyf6gOZJx1pgdapxLCjWoTzAtHjTekbDR9wCDwn
zVu5vP2XH37HtJJxD5uY0rtlLet2/YOx6EaHtkmhWTyGbhnxNTjLTAAeVlXcoPdKwK/ldKECP/5r
x/+jAMIIf+Gx3/qO265kSHv8x+tZi+t7Jh6cwLundz0tTBEEYAfDoCo6gHQgL6w3c+RquFECKQqm
AyOrHrA19j3gk9CZqhd7/3Lm4P+Zwemwv7H4rHws1g5A/ffl8iW50aT8X5EDF3bOnxPvpaViC98v
t5iquPzXPMYk4q9fBvbwfmh+uL8tuq5hgULCszP60icR+IPeusfr8Iw9AKPiXjnxyYbxc2VsjY5/
a5uacML6+DYvBCBOdoLxnYUf01tseygNu8+BIxAWh6PBmHrq2n1i94nHBYgH21ECQa93je3Yug8I
352b9SbSc/ti8jN4kJuSEU0bCoqMV/N3JXft0ya8Il02HJOyJ//yBB0UUuZSjeDvpZtc5iQnhxpG
CG982tvHHZKk8FZyB6vf+vPK2BKgeLfrFccjlwh3bqViYB/a8bEbE3fR94s6Gpym1vHxgYHqsjse
fzO2nT9E6U2Y9pvO6nV7/qeKLgxIHA9Iu7ok6h9rg5eH2KLlly50w+J6ScBS7h/w1QC90gyprvcW
OSnyWZM8T0T3OoFrUnXYa+9n/HpVI8MvcdoZ7z2CPFEdF3XPuMqvyPaJdbeaztTPt2whmn1NCaat
+30n1wYvV4mt5z7dMpC1AID5LeEDmdJWCisb8CHOkqAzh7mivJst1DQFNlL1LqxLC7lKYWxR2fME
2aF2cfQFfvURRtsFJ0oaJxTaZP6Gd0Fk309bBD1CWsR4O2d/qTRUmpIdCrXcEViFQPP9S+Ncnkqz
o+QtJyCIpgk5HDRkHkS0ql0H5sXIkGpCIpibUYPTsldQCpClvdhomKiorO4BlTCQ/Hodu+x6NpBC
hTITm72QUYlm/X7JXuXAwPr5D6F+6ZSVkUVHf4RF2R7uZcEzSuPH8mQ9J0D9DFUhktYyxlzoBPti
cGypjusbYP0KontdJTvcOwMTqC5RjwaLMGXq7QPCVYjLvoK+sUCkyaiLSUwSjEA/t7b7Z0F2Cgd9
/SwNrls7KRRydGGgX5ke5tmk/POzg2ZvFxGUgFh+v8U+HRWe29sBYM1s4nURw8+E5JE8IxzFqgYh
Y4wKiZ8244/UMuKg7iGGnc2rNhRTcMAEQFaa5+mUERu7Ux4hB8dlCqSKlkiRvjRbo4pyhDUhKyub
6MJTkNrW6+XY8M2HJ7VdJZqHdUetheqMZzFiBGw+aagiNc24bzXihvmEEjvdTxiw8qs/NJBinfSF
Q+NQMOFDc9q0PEjLHV5bC7oLDk2GRgoqgQb23QeA93xx4/YmBTWtzf2WaoumuxpFA5oC2YprZl4i
8Bfhm92akKX8e8qf/TrEoGJcrIFC6hENG1gkqOroUDYevDyfBQKNLu9GYe5vurVMgvhkE/olbIWa
H8yHjTbG60KodTN+QPWSuEZzufq3ts/G767O+9wAd5qTD3YdvQwfLkNebHNSZzM8hjrcRTsuLLNh
74Y72E/oFrE+5bx2cerK20hHeniSQAyjZFH2fd6liOwg/osSQ5aWoq4nIwXNr1fgNpTjsywHYsPa
uYNzhlrmQ1w/WXOrcBg8xrFmRAyDBnY71gBzcN99Cz9slLg+VynwXAW6dhY0tYk6AdHzINEGzZqu
eUzjJTLWGzpmtQ++Ms40e3IsrgKIwnxPiRjlaDjNKFjhS2d067lCPHriuW4PtGCv5CSexBgutyxT
Zf3qNTT94BInF29BMkK/EAxQBj+VV8r318v1mezCtGuhVvi9goMGbPEbrozdpKq2AsPIdarMT4be
cokg5fwiwWtOKPny8aMnhCcBGu6gUIUu6SMEcjL1K8+KigaduVWv1Ni7eZ4K3ACOcCVpHkI2ln01
lYWd6IWYj6/vowq/Bn6ExBiNohchXFnPboM71T4ptmotCaupqMOXfXEUlzYg82jUigHqde5US+8y
/XvtfiHv7xMbpwO/8tWXawktzLeUgxIX54esZbaITubHoh6v97uC62LC2mXzqfrVZ15EzXkfvUGf
Ipv3sMP6WihEpITf99kiMj5UgHLA/QivHMl9RV2WM/4Rxpate1q64kYX13qKvF04a9wO6N9pI1/L
zXvs8hYZjJZPztzGt8b9VKE1dloXCiJtW8H62zkZY9ToCsoSeti2iYMOm89BiGTDFJFsYHFvMZad
Nqe6k9SJlGL3hfqmC7dMSPcQbYVXv7bHPSKWNb1uwtjmctMNzbLeavAP/LEL9mi7Xf6FpTGurjDb
bBJa/6cEw9WbgoJRW9F9vw7Qa27wS4QDxHZ9zNRAt0nQLgcOkmFXBUXVxvn0jsGwIOkcQ591suZw
6cgteXXjUjenBu/1fAQubk42uKgMexTFFs5OnBJUC4y2QYewQ0POBjbuEmkno08erV7wpM3HwcX6
3ixGZLiR4iI5pkS9t9U+xRScTg0XpvYIQPUjUp/3qeXXw2XTi2nZInBGyA6Dzi6ap1FuOWT4SqMY
h7JUjD4g4Zv3jDnyXQ7UfI+fe6xjwfL+QLsn329+td76zS093NxGHfHlT1TeXU5NHfncOqdf1FRk
apXUqm6e7ddIfaXnB7M7mvcmVDfi9Al8uF9kjbXOIMh+a/zBYaOfd91FBoxYuQfXySZwzBJcDpg8
l3WYxQzX3HfUYlzeFXSD5ZF9hAQVZBhazR/ZU5FFhzmRZhzBOXRMks4kb2tdoNLg4g+DjGC6wGB0
RRUZs24qHwfztq1ZUZZOL9DO6nPgQhMZMTVC+X/Pg3UeMIVjOeZHDJ9ZHV2DT9I2zr7/1USjE9X3
BN5cUTFs+mu9LczUBm8rDFkyYejGi29UUsgB76TXiZqstmsn3JutrPYksL2YJUWAn/bdt/m+1k6A
iyfNXa6MwkoTJv9GLehmN64avi/HINJMdLw9V4yeZC8MAa5oVC/MLWKS5Z76t+o3LA1BixITHAOU
k+lGU5XbzyYSQIOmy9mCLE3RxiACMXsTa4RWOQZi55GyikIDGc/IJ7RXTcfrqMBTyWEKOnPTuP8k
eKgJFSRKn3lJvr5MXCGuAEfeRp/cpTpDuJN0Vvy2LokQS/QkHkhFK3Vs1+6DXAo1ptHfRxrAyLnu
ApaL1vsbaefnBBal70PgDtBCeKzUY7+y5X0D+BDmumyRB35V7iD0kDXeG7KI2GGkjvNBSahvLpTi
R7vpT8Tq3yxJOV2xMz/5CSASFbHFKAutKODulMU21k23ryi7DDIVD6RjGHZR5t8QU0dOrUFtaUJ2
AC8sAqVI/hR+gHVeNNM9EGvNFBbhFfWmsofYDOs/9usH0+kRjXFGPyYA42s4UvGKIiJT+eC/K5XR
wZiMXWT1H60K/ppI3kdS100vm9zPp4g8zxqu2B1j19CQRC930bS5acvY0vOU1V+2gyZZG+C/tViz
COy8Yjdng2sPDw07D6PYwNcJmLdNeLslPXt+ZcTJcKc9iRKvSFtnboZM9xCTd6Mew8PIAFitKc6a
e7VtNPpvzDEEnv2W0S6xMroJ1J5hIMeViUJu4mkBISqawgsZXLYICEYHpDNr6EPZkESqkV1apdW0
HzJ8sSsDy1WruWFW9uF036DaqKayBNW6fLFR5oZaj6WFtVGXt8HQB+jtM0BPs6KS5Z8nn5RkqAcD
szSa1ayvCAHjqavF0vo35qfiAQsVc7OPLfgBz1gksRpWysdhdO5E3kzBEESLDBDnFqWaI684BJ9H
1qYFb2rtWGW8GI9YLUADDcrSTbxVYF/0VgWjxGAvB5JegG8GYvSXVzfteGz8ddCLJ0k58sNXiNwY
I6XEkz7A754T4kXsaqZTDr4bteCN1/jM0HOwUV7iY9sPTM2Ah8+XzuC9q1BjE3SfH4ZLndUiBRnn
gCJwX5Ydg4NwaCKwqkcX8k1WlQRm4Vuv2FYEq+4QUS9mkVtWMuUYHuep29onx3U6brqa/9lfAls1
u1Rdam349vO9s9xHe+A1GK1PPFvV1/N6E0cogkTcD4PeOWnKZA+xfxTBO+ovEX6SXANQqI2nmtko
1NgUHf3A+5vGEz4qZlGVqv4G4W5pQ8rE9AVCrMrGCmCj01buiRUIxehVeMkXVZLJEJC9qq8CR6Tp
pTnU+rK4tDoymINTvaofE+5kpZY/qYz5+fl9/rarCJBsq7itmHz2knZFBJXrJmOmX2RZqtnKYUXv
uQie15iZ3jZGc8d8axVY7mkyuBYITV0B9bRNA+PLowAwOBPuPxfyE5incaBXZYeXifTtO4wcfYtt
/6tFM5Yuowc9ozRJkzziXFaeX25UEmlBuXvPxmb/UwTnWM3n2iJVob6ZXcwOicCV20EAzriK+U1A
QYP9iSBNbM6z8Jga9qdgtKjgx689ACVKrTKTwraMJ5tfUUvXtaqMKRaKCNigHIXX4VBNK6JpVjgu
RsYo9/K9d0kEPVX9pgrsf0SvSQcH23PpmWuHSsIrGzvLMk5gPC/cKQsVQw0mqk6rUvgpNIwAWsNk
OBqZUdSm/413RjHVgsrTGvlprD//7FrT+n8FY4ukTBmBCDy4wqCC7rfYtFvmjceTFlYaYXa9TMwZ
WoouxErvFmBNlhai/BMgRovhAaKL6wPQ5eetP3lUjLzbBBwCrtvqhhzn4+GPfI7apL3u0rruA0AC
tEWJHky0qZNm1ZnNzE8NntCYAXFuD9ekE2ZmKMiP8zJKvR2Z+QjEMADWn9IumO7c3UhXipyn45wF
JfWFsD3aEHV2DsVXpdhXPDn7Ih0u5fvnSxAXp7E/LDqgTemMQQxGu1chaZXKoRIrm94Dshcwh0QH
R+8MhHifw2ic8dlGQMm96KcpYAm+GTYr+/F2OfzrX5uL2MXIxWcl0FrNNXvMITWKwq3FKKMi4GAn
Ii7murnAcN+rjdKaUOUdFiG0jEvN5YCu+32YpGCMaissnBwEhAj/E8rUtFx1n263xdK4vLOQIRMC
oiUT7zEIl5rSMOaZfWFoddY6vk5SC/bGlkWtpI78d9A40aFle9MYXb2aBXcneKoA5CASBboYzXFJ
/3hGVafkLXSSutApDq4aH/7hrn4aPzlM7IC5drfNevry2ibkLLaHhx8KE8szoan7JFcThp0UZoCQ
LKGYoVWUXPj5p0rzWxKKnz8WFeqrfEjI8+vo8X9wYqThnttAgEmTxGFRZNGYfRlfS7yvaNWxr4by
goU3suAg4iy0Zj//nICsmWFyXvw8WqEngiqj4TktS/wFmUsLnEJUYtYlxRpDLjQSOntCXwGAsvgO
p1sDsxiKPmZ+ssRh79sdZ0DTCu+k0cTOaq91YHy+DKH/2gHTYFNpsp5BVjmuMMHV1HQGy4yehQlQ
3j3OQ5PVPRQFon2i3SS5uUyROOu6eX0ex4u4o4ExkYG6CUjeGRo4Wemr/Cu70vThGklgoO4/l4aE
Ixe4GQKUbQUADmRdelALmKdGAlxCoxqbrIiDRkHMFMpgVPhHKiS5n5RWjIVnl7LMgBDUH53i6TZB
B54P32Ye4nHo8NdDNpIxAoiHGlgFleGCk3Q/SVrRfS5qDMc4jsfL4ipb97ED/46xicdml9YQy+zm
XoB6e8mDDEQY6RIZ4ZqswISlqzx5FSmRYmHjFXDXQ2ErmJ9GyNVbiEM3HuGBu6vA4kJRSqS/EfXz
OFLuZPiVhVQQcTd3xaUT/eIODae56YDRitpZ4rlIoV27wu/mp1J0ENAsbq5+1c6FCPf5KDkOtdPf
ILazD1nUYKoejCSzULtQhv9/Tb+SGmxUDejTj8gw2JrG+CUFTx7GY7g054Db+MCpO4oVuPKvSrxi
eGoD9Sh36Ji/PQDaoIcKc0xuDGEPNhQALTkWxzDhb6PzgbSFbNVCJ/NvWIpHWBb/xUlMRxak/oue
XjErf/QoJT+pmnHn0rkjtANK2CGq39WA69gjchUcBbfNI+6AJpqMj1kOdlHP1dTCxzjRkMAwswq0
OCt8XD3OJOT8qh7yWJQOZcS7vZPfAy46I1E+ptFMNdI7s0rADk8osyOvQG9YwjC5hSkPdlUfjbPR
AKPlrShqtV6KYo/jTq93KnAWMKEYmAiVZHluS1+I+OvPz+f3jtFImLzLvbZwjOE+DQZcJvTnY6rR
bc0atUA0ze+So1BRFSPJi5Oy1oi7Gn+M+dW8etDRQ+hgPjIWrudGGjCGrNB7RrccHn46mxSDyFDw
KtxI4+WtH/3w8TS7dKy3X1sipZTiqrO2TlbvwRHseKLvS5354lK+lBpLDnakz1vXPNhQkIsSrX6y
DEjYHON8kGtgM6lpLtlB9K737h02CsHdkN7Clb0ICUe6FBsNhvaGl8ebO5QBSSgXy0dWarduZW4r
GVMMT5c0Vs7lrk0/Cl7dgBiCsP0egQvicrG82SeprYDlyLa6zBNgFZTLinOpZF3RqbbPWZUcR1WM
Lne5geOXQk6cKK5PfsYSCgpjQ1oslunetJ1j5GrgUnsazWqjM+8H/EZVuFP727+CIU9uwSGexIbC
DT7KLCpnufq3rz40gghx1BxnzfYkCyACeaSLUAKrSEBpkZwDXl1H9rWDmbT+2YwC7TsSe5I0Xa7E
hACUi+scSCj7KYYjF3ek895EBuqfADKRp+mDlT/tQpCvZPnAXrPHz6RsK76hJUM19pg4qIwkjzt0
Pg8/hCAYh/uEWrr2NE9jgfYA+yR2Tg3QH772p4a7ZRRfyCzyF9Rf1S6jJSXcVo1d7QURCaU2vlnD
OGlweHT9CMods1BeK9bnc2BMrGRNDH41AIPnNA/dOWKe81Si5mIyBCQqbiOJowVaojZZQm2qCeCV
lLrPwkdszfsdbpArCV5bungZXwWlNFjKfjJIqyB3xgbWd/tPA9tvCLVbITnVkWK9aRGy8HUDLQNw
APJLIcVAcltgV4ZuPKZwyQK80dV/Ben+vgA6hQ9f8X3NoVlBC9OlckPUEMNPtBBQNfGhGV6/nmV2
xINaaWdv69MAYsh8Vcnh01kSi+cwxaMcZx2yxryRDSaKxFc432e5CFaHbDaHrGAkIuG0CoRljELl
yc1vPXsOOTahB/ucKSrqtH1pLd/iumT/ZytefN1CHiYP0Eii5fZO6oQM2kILh/LdWygMsFwawdIO
3k4X7tnC8iux1JOU2D7ySmSUU/6Rqof9FVi6zkuGOBCAsy3kBbjXjxPUBxX5Kh07ON2qwvm7qEkp
qV3+46M0P9AmSpReRaP22h6sRB/cQvkVKVyba3tup/lEdFL4cNZmKmBJJWvbDVIwtuwSNQAWLRKS
HcP7c8MEVPQeiEIrBBYTxTaMOyuZB4n+LI9NmMQqR5fSX386fMYJGzrQu8w/eW02OiE0SvqSM5bd
8Ow5uPCco7gbd/TuwTIMpo5EJtJlCc5iq2S1Q3MpwKCHZE553Lc6EkUnvXKPnDcsn6X296UuPo5r
NywrIVwHZMCqNiSHZeevXl/NM3U/IL98pRDB/h1VyHXGKGWp/z1SxAflogNpSfZmO5BsB+cYKvkA
0fxzEIKvEp64xGF+7wCkMy999IacwSL8SoTrxt3t3PyjygtNBNGWLoP37UOuhQFWsLtMsmzLobzT
fG7ks6SaPXyGFZI1jX3hs+zdmacRcr1S4BNxJ1If2lrs8gQJcdL7eNkHyBMfxXv8we6k2HRbzk6E
5Pg+7emughuM1HSR5q/tTdEa58C/79TfHR3j5pzR/FaJmNuC0UUX4F5tgnfB0EVqZVSi43Wb2AXH
KnUGiTWsKXSSWQ2huNB5gzsQDYD/vexe7ToLYcJV5IJf26ovUYJ8xLSBsV1GSkg83wYA9F2+Ih+s
dlxuKcmj3QXNikkywQGNiWZfBWN/w6KOBCCqR4ifVflq7UHg8ihTXoGd5bb6elwrJFoHzKiL7exN
twIf5r6SdjRV6UvpwikRzN+/r5KrDLxqQIq7yCTDB0g26K0mQ6nsveuyZTq/yrmVTNE1wFKO2JGJ
G29YEMb+Ya625gPVZtgeKFnNHrcW/EAmst+0/1Vu/InJk9WR/VHdRwpJ0wMCE3eGZiVSneHT2VtD
P7cy75hO8hJ5NKS4fyIuEHjcUMpmyoHiwF2tc4JEL/fjfi+4MuXTwgoQBFDnV3MdtlfasbkYZMg5
+Sc7jW62Rncm5StFdpKoHvYzdd7Vpz0cBWuIHvG3kT/PB54UNd/YQiA0VxHyEFNR7eEU/UCM5XLm
9ffI3qBV2lKv0vdARmpauE9Lgr39kqsXZI0x0hFXclfFFT8ug0bDAB3eFxglHKe/1n+Pf0EGACcG
f+SVUanSJL4cmba7EGaleydgj25kEj2ZH1nSC5p92ICiSbv6QoR/+DbPEofDnaOGYoB5INPzPDXK
NAwvEE0loIX84Ikzv9di4j67eXuRBWSR40uGd5wcV623rSKwaNGO1SDc75JXRQa8DfZB/ZAUP18U
c8slHv4oWB7ecuJsAGSSSjNBiZkFvrvCpgiFQNSaDEr/h4RaeNrzIktR0Eb4mUclTt4TCUQJipJU
C2TXnAuTookeTj10DVKqD0EWHnvdhTyGR7vIefxMZDztGD3V3vn6QwajbMmpK8pK1Yj0KNBC/Ik8
xLstSFULz8/PdGKR01g+Vug0d/HBwmenK6TbJHK/pqwwHkLxj9NcvOxP18uiukeRXrfXbse383Dh
xfTOBThOBBgonBpyHdH+txNOGfee/jcC6g11FOQ3W/CTIQQGpBWsI9niEXq47mjrQo2fcgTmMokx
ELs6NjfcefGte2yXJjWlx10a9DmwnjM6a6VcMpo+W8Nx0nvrfANiUPY7ivPdq1VoHd32ER370XIG
vNIZOeDEaiaLIZrtNFWmL0Ryyw6yCy1J4K8URNJ+yp+JsJ7pP4aXs0ZS4RW2Q1jIOP0CGAgM4clZ
AcvMiqUFdOH5VZF+mJ2ePEc4oeVNZaUR0UfjDBg6SwuKSypNEaNNTFvM52I1aBjNckEtU49dLjAo
BMtIJjPBdFdtg4AmfH/ZTUo5i/dLZfwzp8hkt3HVQJYsi6e6+8ppj7wvAA/x3IAUQz34GqVkywpG
WGt3aBG0pOaWrI+ySh0KBA6ZqxHg231mqKTZmu8bpCi+D33kXHk1X3QofN/CAazFqoHCrr+qDUet
Ajy8fGRBpb6WzCOh2YNmGX4o7ceGswC7blmAxNudwm3F72ei5Lp99OT57P0Y6GSNrsPqXoC/cCQr
W0gHBRghCypiZHLIfmoF6XRp6SUtGwt4pwty16Z1bklxUwHI+IdgRDGseW7NSif9tQU8j2C+HHd3
WvqVddSdkqpVY8cR1QKnKwjSzuGHOa7qiiel+1uujQqAU44Sy9EVLkEJAGl8It1Va5RSK/cQ+9GJ
YJrO8qzkXnlA1N6aCzudi1wbQ6Cm1fe345JZA9sM5rTL2HELBKoTD1w0F6oz4sSkkEpTKjJbXT98
D9BL9irImOMiIZNJofWx8Bq1rjzV1ZCweYSwhZqou0zNmoGh8R1siIOWf2ppasD3T+JYwxsgrsBs
0ZIpw58KMIUexne8yaW/ROLl+RI/hUDBpACnflRaQACP1S5WcQ56J7v0/emUhFDlkPYfaZDi420z
pPzGgY3VMAXMe/nNTGiCOQLpGEy+qNLHLc1PP7sc0y+BmqBfBybEEEOfmgmb80s4lUJd8gfVkupw
JcEQdxw/kvtip2eGwYq7ALVdVgov5DmsK4pJ25pHqwIN/SQ5PEexkUEqPZr8yZXSzc+9n8+3Y8CZ
uWuEo6q2YrSivWmjaGPKqqIwPL8A6KoiszbsiC2IGrSC0m+kQeTAEVnLDB7hRuuoWbe74RgRxxpv
5Wogf0oB4sSoIOI1qbBpkwkKV7JMsj5Jxpp1zRFVudfd/9fVXWFJ18GuW993ghNH4T07Aprd9Qnd
BhqrZLg1pPVsbzWr4o6mhfEVItCaZV7FOkWRWFg0ay3bUlSqlNmVEfhZCpiMoTtPJcDwduLSDvOz
0dKxVIRkOIbJg4t5Niw0JJntH4Ufrqha7euBYkCp4uOjpFG+tGTcE6K0In0+Jtr4afogmxDKD+V8
T6u13ucUfnx++j3qjP2kX6cpqNRND+U9TqJSr1lXkRrRCLrh9IKjhBIbv1yl2Dary3p3Vkpx1znx
LnjrbgH7+FmDVNglV9rojaBp+PLa8P1EKwZXINu0W9zaK9z2OUmcT3YfkZZMLMDTUCxXy/ZnhLYM
9nNv4mQ+fz+yWcjlfSPcjGkBAstVys+9/ou+lNniF+ijWsUzawedlWaNAa9AWHG2c9p9viznNZep
NthIt1NBQ4m3Sg1w0gGMvTZmGn3zajtUT6d4FoDfWWf/ICwYNrQA/18k+o8rvmfWFI3IcwM5MWhY
ppU+/l6D2+s7Kz93LWpGH0WT9lhwZxUWmW6jhBu6GiaRF3323MGOpN1sFLKCXQjWadDXkMRHJdac
sFvHFg2rvG/RfqTuWocaG9DYD/SajmJ5j1nS7LfNW6FLzOT0BvDXLZNzr1beRZpmF+3bQ49TjcKK
f3DtmpuftkNZgKBmo6Ts3JOQWojoX2P4lggTKWc/LhhF4vBcF/Xf4kSC4hdms0zaC7pxDMihAwGM
aqv8ETGlVEMcwiZKEntG3OKTAC2qN/TLcaab4M9FgLoyOPDduMHXRujHsHDEz9ZZTCRMH83cydKz
9zRo4prKt8aZ8NkL423XrERwaYH6nQHYXvcEhobPqx6Ul579vSObEYU6OdPLG1HaXNqGSTCaczCz
/Pv4jH5ktk+z/fxVQEUSS/EBRtdewCk8B2Pq8svphRh8EixrNQq30A2EsUt2zyQ/ULo4PZHsZyOy
lAgmhqPQzbWekZhN+m9uYlEh6FgZZLeMEVKy+bEvXn4fsZ0CcAiKQQVQPfXORIbLQ8Y77jzb7H88
iEXt84/XupXbnFdEv9x1tD7Hu69gcsW1u3gHGDz3H+6h6CD9KfZYLTZShwtxj3VzwGIg/BHTUlJ6
zXwbuUpjollnTe/TnLOw6+EBLWJ65ZE4VRfGVj4Z8nrzY6IXRmUFHB+c8NchL3MhI22Q+cjdBobx
fZjCWJy77NOKffnLjKG7KRatJfh2tb0brhHzDvjPU7fBdbrD1Q/V7VhywEyTeyMBPGgj5T8Scmtc
6cKqTYtYc1hiOn2EIRegBqFxu+VQY5yjRUnVgcnRnqbUJxUYItSEieB3k3DLi3EuIqavg5LCq2Eg
wpGcvsre0Ga6GXTReqT1czHdDnBNXAynnLhER8wQU9KRNkPad/zTafHl8clIHed8ppqRYel+NaSv
0h33gGvxIEpvqaH4d3qFRKLRWy887oPTCyndNJ1IgCY3eFjFWg01GTIcQ2QG9akgJbNJ+ikH+IH3
XWg8YmvGuzzjJa37a2c0hkny0t6iYujr4IgqQL/q1nW3oaaDA/Ni8NNry4y91M2kHuB8SdZq1SVp
yZ4970+F2t/OjfKiswcJgOzWkuDj6UIKeU7IZbltFj+fOTl1hjEm69+EJ/rzQvUAGjdOESSW3sJr
Sn/QFMpFzQfMvhqyetEF0T5NP66N3WDOCaSjI+Pt40h/KIlCbEbJix9b94VWPIXmw5UXhP1Jpdjt
x8a24BLCm5FKd+ouwC7wNOEiyQHh7SoQAs/c5VXKmktNI5Pd4FTZau1de53RVfQzzcam8tMzqqfc
0nmmPLl148mhbsY2eVS7/OmTfQbM4Oe87mfIKa89o+k1W6Cx+TuXSIgty+afbwzCGpG/ukiu/Q3K
Fxk3birlwvp0VMet4VWd0Y6hxWbr/9V9P+FFGZjTpUq2gUhSVlD7JcPdKEW7TlEx+1Uow7Wy5fUw
7nNWgOnGeonFJIkZHT6RBvrtlqCWQQ/YtxoHl0KHeO13c7viKWQ5SkqooNj+kD+dg5xZek/aoj76
BIJqFF+omo5U/t9mEZBaQgg3BA/59Ist/yYzdVROcQE0ggthvBkcSa/pdA+3P2zAacjE8kWgFLLw
KDQP7fDCCe+KivkEAlL6e3hlGQ4GkKV9Ns7vHZxYR6xbiMdo+Uryww+/JJ9A5NeJKhk5NHpgSWc0
D/FRnsW0LZ96Yr7lD82DWIpQezxA+iBWjox2J+kHHksoUjl/SAlMepBpxllequ8vPLJPAMSlYL8Y
90AnwkX/u6Q+ceEbXxM5aS+JR1CwVUA8pWB/XhLQbeZtSeaW2vJScl755FWKunPE5+wap/ThU1Jm
p8c5ZCa9H4BMiVZEIUZaChOEiOUN3CynNpfcLJznsYqLIRL9GIOB1Hxvia3yzl/f0dcpI7D+7eFU
rKkSxCBoxf3mGmBJXyJ1c1WQEF0hYx19hKr7aCuYbh1yNygt/iIkH8aO4S89oI3gk2sqISqjAuG8
CNrAu6xrcwOEGfCV5/7TEw1MK8agCxppiPojDtJwdAf1WyFkDvMBlCKfuAuE/wkUwEp5VTjHNEio
DQVB3lLnmBf8qXKEcqGH3RZSL64FS2erJtjiEcf2TVvv6U+crh3vD26WsBu5u2r9KLlGtVbz8tNp
Qujo8+SaMklW/y9VAODmrR2OgZzky0XIKKHrE2+Qn4A5K1DyMgyPde3LE8AkFLcwj+wodk27nRnZ
nIVRa27gBO4CCInSpmTQFszGqXEm/WdrlOlCM73a9pB2IgxfEIpSFzLGtqieuK1t5Qpw6zoViGi6
gAP9Qox3coOEJy+SgNrsNv0ZzFgeV3K0WHvmvbKaEr0W6eXKrTjmswEOtKwzll13+XCmUWcLYncc
9Dv8F7AjK0Ff6vSVvMVvpH8feHv5o+YOThIv/0+aS16jp/qIt3NBAMQnY0WzuR8lyrRqn/2zwqGR
vqvZSvPI2CKr6+now+YrWGBbNGUlvYFtmbxc4+dq11PmbFpwz66I69XQDkm/xXR13TF5APoDAdcc
ZK+P+DIGUdtzK3F4sIAQxpQgk5sJv2PDCYRQiUgG3vZ1bzckkZPfSCc9G6Mys1AQtJgGvhbRf/3C
a44Cim8N5NXxBcs6mbk8mZCiHVptxkm2F3pXSge0oAs2FnrvuwAMV35OMUUdDMBoZDBycow+5xaN
7Vi+ocjDop+wq1pUZc6Hg8U3D9UG66TNypog4t0Wa/eYCQG1557rO5Td/xAU10majpLj/ww9G9gx
kdY/6Tbht7C6gjn00o2uC5Etc2+q9bvtBDhGmW6NiIksm5S3ILrc0vT5q48o5oufSwE3Mxiv0BgB
g05fv7jPFc0Wm9nYibWpNkg7vQroNbSyKyezVFJ15PdXQrHK5JzUlnZluD9IsFW1QhhCe2hDC7LG
px6rf+NTEo+Ee9nvWudiohOc3mer/GcJaCOJvwrvQgY5qWp+NglhgKigEljd0S/gJ01l+H3kGXCZ
oe1D01zZ7/miAECTtUNiMSQRXBW2bc+2qGSF9cRGy8+Sa47TbOsCeqgJrRKOiiak5B2J7bAWvZEK
Iyz842p3CCwFIcXjnmb/9PPci7c4za88Iu4uXk9W8q1nD1QJjBgxAzZ1mKrLJuzixf+VzVCtWNGl
As2hvH3Ou2w1uY4TIiLnxgx10aQWMW39Z58nD2jF5PDKxwYQJuAiBpY0woDL7bgFY04bIrFFzoAW
Mof1Z02Izab5A00TBt/SqAUHaNta7RDDXOGhy/PM5eZTAOHNaE5In3agner4ZlrairAJdxu40e2T
4wuvfXDA+MNlcPmjy6fI1HYxOhM/HFO6uHUPYyMS8J7nZrm6N/XQG78Qje6VqrBccdV48b6CkmaR
oOePKETN52nZQuEGZUBooDhm8m1M35a+hxsx4X3/ibzdUPeMJPOjVDSWGAIPd9a+aPK7KrHQqMwP
R8THBqMxg86p94RL830XL4dwgdrTvMY0GOiEfWwii5PHCfL4FT347UwToFo+eomdS5662aMy7dU0
c6VQKy/qJ+KtrbpJvehq2tF7xMVjJZOPSUpdQ9rlYxmNFpEt9hxFbusMQBLFAFEKgk8jmApJscZY
Mf4NzCzOnMV8LwsjnPTReCNjEDgS1erZrvLyvDycOGBLEVL5tM2KClZD3Qp2rgRk1t/BMxSL+uCG
1JF9t8+EmFQsgo3KP3mQtDkVLXkGGqy/qodrPeRiMxZGgfOGVf9QNyOEHpny6jUH4baG+qjEJvgk
sNP1gYqQfdZ7ElSIA6t4JoX8UQlyT6etd7TBWmlneFsHV+XgdRQaecFXWqvIa7ORyiiLyA5bnWkQ
ndbk042vTx03Nqe0g6n65fn/KJWVI6cxAo0Zf5f/A7+c4l8dJphOaRPyOnfTzEPn65ESyll6GMAO
j4eU6MTwTwutRSJOt+FCyIjKz7c8wrM8jj+dUr4vCHz9kfDMyMVrSi1HyfHHRHa9BJDLkoIvMKt3
K9Decqw2m2p9jDgqyAvB+Pxbg+bcMeedvCHx7c7tEylpjOH/rqgAwIsnLoZKaRSYmljOv0AyoAYB
YG/48uOUFLpeVoop6KrtLKFIy8SkDRcssOthUNYAIQ5iUjTGw1qyHAe816qtHAQOKEtWNbJNx2eD
N1j4cmH+LBv+uyuAV+UUPyYbZWBYynNPX8ZzLD11p84jMJpu/dJdmWMkuIYP0dzU4v9/+TQv/uO+
lC9GfmxIOCVHS+ah1xsRaKpjl4bPoa1DDZoYLdzKvqueK5Vm8J5GT+b3AeLeoVvoaMFVuxYlOvSJ
H5wTpguuumJyaqHx3mpiMxCvRrPPguhuDjceyDieqDR5cgzKzJUM5NdcENz8s6/P7ZdgX92MQv31
7tTob2B8Md7sIMYgCYFlmECgcN0R49c9QtSHfi9qjkrW6jY/M+pdMTplua9LSHJYjODrJ3D9ogBO
bfl/VQnX04c+pzJN7yeoiJUfFVQUEF/nYI1Q+cWkCU9l/fpfBXxoX2So5tURBkYB+TC4ozI2H5A8
9vV5F4Ey9p81bvj1SYmu6gSpPr4Z3TC8sKqVhmHJqhjKlffM0rUBEUR9FbDRoHkapMhLcIAmWbiC
eFWJnR+Y7bB/gEpwRkrjlnh1DkxtUWrKSthLUXQksEKgnPz+z7OXee0XlxBlOo5lLFcx2swvIqOO
gOo0uIdY9AWgn5kAqreH6KVjMCtze4T1hDEt8QU0/eyz8SvSxmghK9PuJ7VDf0/NrC/lsDtFmuo8
uugUJ5RmewSInEp0KGsO9+Snzot/AWGn6c9rMk9vCyEpuXWWWH6heSLT/tKnG4LcB8FBpBh3AJWe
j8n+xxpD/IL/ukcIISvCNI+nx1xw6jTC6sbj9G3UCl+ybQha6pwMJBNdV/lZKe9jG2EmHLU8VEqz
3uM3+Z8+Suh9mj+eGsevpOlf/g5Hx9zCbzhZw9VPwYbtL8CPIdh5jJsNy5BmVPy15DS6VKBcQW/j
DIxQjYEyhuCQQzljE7GuVYv0AIXctrCC/diQs3ZTUBtsBsz/TOyT6hSycJbnYLIlg1dHJz1FnyQ+
CbQF51F5BSa/FKd3lk3LPDUL0rmMYpNc0hAWUzzQGSPk27FD52ZPl79XNyMfwDjvPE6tg/QvbuG8
g9jIPHMwd1bZ6ZmFgJ6ahbBSUWrZuwn2jCOigShOzerDRNAXeVydQqaF6dCIi5zIIJzfHXupEfoG
tMFi5iL+3XSel2bNe9gZSek7MhSvxsvx9RXOfCp6DJn9ubv8ddU14z8+dSBBoQVoO9MRXc1xncm8
7pvCS8E3SBA0+HeVuXgQcAEnaj+GYjppuyROGJNj+DZ3wIpjxq5+ApSNl6LVTv8AGSvJ5arZbUBH
+RGmIUTeMrjhsYLBBwEdrg/a62VI1PaeO7BAqwer48Kfg2z01b0N8WGySjfdiM4LHZ54koTjTxD0
3LPuj8MLeEtx3JeYjnKdePVrAVyp/12blEwOlTc06Ota/gy5q+Dhb0Eq8jzJw44j5E+FrcWQxIqy
txrKFNGxCsiPMw9PMad8jtRz2eG9/MGyXJjU5/Pqbab1HyySui7GKpyfgHh3pDtnSO3Mbv03hEqO
ZCRY/jPsoc4KGx1vRU4w2GTi8OOcDEysqulqy2j0rSlnPM38lHkJxa8vYX3tpHboA1YK15yZ55Zg
rBbBL+GFql4I6iTf9cSd6RGy+XcikO4MQHqs/KVW9y4F3/RT7kYpOgeHbN2y9HdNTnkvCoN3QRiU
yko2hBUL4Kfbvd3YVXPBovnkeUkUWo0n2LdYumqZf4PnNtrw01tnGE78xXQ8YjQ0ud8btpJue/LH
eKpp5Kk5UV+q/UyuqtWCu8KBx4jTQFz8Dt7SOtuR0bwU0bV4vKVBGoLLLfQgrsDxDLwsHBiuuahx
gXPhO5nCcXSFNwNrY3XlYm1tck03MLeRonM2Vxy7d7M5cSEvblrZRLOm+iM/FftTRPAHAJEgm1wN
H5xmMVziyXfcn5t1YpmBMGTNJR2pvwKVxgX2TvXulUXahjYQjZGX6l35PSDe6aRkHK/buZf9OPqe
2khHjGolIULSgKU87iBNxN+OWeTghzRZWm199eju/jndR/66wQ+s2QuTg2brQqtL5Gz/KXewkbef
LSTExfTYaIxES/yJOWDgOPVEg6qMPrGjV2UJh3+KYk8m56aAERLbMB4j32nU8ylYYVaI17b3JGjU
0wkkqkgP6ZDdkC2gkauEwwEqlNMchWxMId9M3p+My6FylS5e/nBJaxga009xe7kNl7P3uwKNfgON
abcsMrdXA3yn38yCg/rxzbHu6lG5NM1j5N79B//BosQ4/OS9TjQ9jmMpnZJJadc1mq37CEqivVeA
1pfDh/GO9vWD0xnZd791gGE4OYpCmqGy7VLOrD+of8HaGNMnRiHz9QPsB8au3vFOcjopksHTHWe+
AA/1IZx2T/TgmJ4zBCfttixD+s4bmp6wYTAbBCgjkbqH97kJHRtQemogsT5m5/1lKRcsL0tf86fa
TuRRtiovXB0cO9hvUOPeAPEo3g1hGr10FEzcuFsO6SETNTy7oUnyusgBi9pcXvgXgUDL1IpMS6S2
jZM6rYCykdQl68uV2WcVPL0l1vZ+KvCkqHzPLr014/Is+s/SEo6e8Ebqf3yCfFhsHd3pcPBIsrE+
bFkQOuN/CZCbmb0DaMzuLWvIWqS1yjWFn9fkbNaloPAcNBuiX6wTnWWgpXVpWm5b3/NgoiRvQSiM
1+VaG4tjFFuGq9JAEGl5fVwZXAGa2AFrS6XFdfWR+jlAxItP0zKO10SQJiCWOFXH3EKabd2OABZY
tnzHIcb9/EDh+iMlqoaBJZhFbpz8EXCWB01MkVzkQohzE7JWRKMYtcn3bJc2VCga/H6K+A4mLf79
891wW+sURopMOkU9L+zgjvzqSAjDxW7J6JmUfjbGz6ikgTd5G5uTS/c2h4CmoWvfeqLrxYXavyKA
+83zAi4BCihe0OCYKZ3vprPF4bXvFm6CjoMFVSUN5dC/GPDqBsFwBCfG/iZL2CEXgA0FN5M+U+g3
edtPp+/sycEx45jctP21sQg+a62vir/LpRGVN6rc8wAn/jV9hrnyclRjk6RuyLdT6uRE1jgQWged
N233JgZQ64gLKutYWC8cvQzcax+hctpputOHuyLkg2jqlPVrsQpRvVi9h1PWrFN5uhRpooU/v9yP
hkb18LGLJs3abZ2cltO1YOx/nb3M7JOXpqyAAei5E6UatXsTLZwbSh336W1PZRjQqMTkbv6PEIdf
vA1EOR6d0QeLIkRIx/wi32Zspnb1rc19dsvXcZNjhBVguhjr6GjMKiQggF2Ot0yR5+zDQv8mxncl
kytjSs0BdhcXK2XbELW634OnIl5XDJ3S2+iN9fi+WRZy1RLVq+q+DIk+ZRytiJ0qUwmYPo2i+cMl
CgjXEka/NS4QmT4ia6xf9Wefnb7bBWSxLmswlhhF3Tc4c/3UD70bNiAd6nV6aX3F2q+vo3R3fMuC
x5qHJAhdRsVSEEJK70XAl/Vb7QDb/J/HG0I2S5a4sGUhDujjcskcrjMk5kmaK9ucYa7QEZElAJQp
jic/2ueQi7+KMxJ1BwGZouzR8F6fQiOpsAWfMdyzckGPOu2tTmWS0aIyM1c9HAebmkThZEG3Ph+x
oDHErK3FBtibChk8+WHSFEh6I9iHAGt020WlNhaJWmEP+MEYpJIMZWw780qsBvFc4mDOSfiNIMb6
+rhs85TE+IPuRxHTzD2Bv5Ya27MJmIPMM9P3wELhkazK0I2NgOKhMktHA28dhJEhKbL5r7fCmldQ
yRnb+IkG3kOyfPfXL23t690V86RkZmD1dhOAJC8Ag0jEpN3YWLhHH3C7s6ObaRlhWdLST9bBjVat
OqGW2fuh3EI1sdD6aE9iro3n7d4kfMB6q9HRA/q4gXx0UdPqP6jE43YQWRFSVZKREs0hBffmIO2Y
br/hf0EcvdARLqXJZEf918nU9cE7Wh/EqdTapQ1TTa3bcCf6Gq3qCNG0SnFnJMjlZAGqhkXuMfdk
PgWRA550XMZCoDKfmY0IIE3V66qfi621lMVZ2P31iIvO/BsMuL97swMYXQa9yNNd5DdL5ofr1Iw0
ChxBTO6KKn1uHtftnm/Nf4DMKLZ7ynBinWTibbdQ/flRfS5WWp12jo/gBfzfTOWPkQwjI9atPoTC
C94EMExBG/pQTNJLZ4JkdiRmX9ugccmg8Bn/zq1M/cNOiLRtH6Ib7rCc2aAvDz0Bmz9/ENFsPAvt
NFg2k/xo8aUwmKDxyydS/ggXTYPTUG4oTiQnrao80UDX8sLQu6wD8N0DuZmLimE+ttx8RXWATEJk
6ZeJdjY4+XHYGWA5ISlzt9tXlelDmDu5aczqUAh1v7eK5XW7PSozUQu4zyIuuMnhCcTDrk7nhITg
GHqckbzsvzw1e5TEP/cFqOFiPXOvdDoNa6QcF4Eva9WQ3aXhQUAAPyu6YORFLC72BrhUZjFnAtsW
JNtKVgxiNhRxGjFDN2Xb17glec1OHDtbejcwicbJ1t3puZucCk8FMkQhi5ksJK76qHRVm+xDWI3I
XEgtLV0Cz00ZJ+ix4chJ6crU7xYXghZ8OUU2SAYH27m6Jv3H6SbdlKRm/ZTRQ8dlBSgTBwsO41vB
yKHhOLXwu9aTP4JSNaG4v6eqnKy8pGZHTmTep+dm3SimJJEx4890iVxTktqfyoveSeYbr9K/fbOC
eYrOLvSXHRR8zQIKpJj/0apUMpgNoV3LNbuOMWA3xmuNbK6y6yZBzZpwfFH/U5yk5WSuoPMoISLc
4u4gI5BUqYnSAqnH0kAYw1+6mTgmQXwLPfHBoL+/VTLsZkicqLTkwCdmWBTMqWT5ncq2Itd3zw+m
l1hCHeSzWmLyOqZFwI942USzsag3idahlFqyR8xzOzuaGumm31tnyxq8P147cAd/bRUtXUMA9nLo
DGA1HtMtgc3jLOvACRlI92puK90SSAgs878GnWQzeETtaxduzhz8CMENWpQNrz9c4j6PdeN9WXPA
FaITfqeaXRCCt3nzJ6SGj4sUNCfZL6Cgww1TPuVQ49SfFDUpD0wnTm1xbmJvTqLMQbTumFbgHzCe
+wxvqTiMQD/2uwbIquMeeJjedMMnyh6tM70GBVpILuf2pfmtjefjB3MTgTca457eJrxO72CjIqPL
u30JPt+QN2u7q9AZ2Y2k61u3LHCiapHNzNJPPcDhiqbiZlc/fmfx321WLkBIzEaFnvKhDiBYvp8E
sQtCoDkkcs4AjjHFOZv8CpTyH94hpeqcCC/ixvw40CErCjUcaCB3W0itfCn5oyKB4Z9SJ5worpwn
x5SwNsZLNfDjQBW52JaMHAgQpIMr6xjbsCbtQKDCC8eda/lu6GAD2OnWYmefr7HOzyc+bJ8a//a4
GvDWbTxSktov63w3CLhnJxuNyoq9ipGreB4bmP1vuXr79xGNlUCtViXTo+Tij+BQ6lI3JNxPIQ/y
lMJJOmIFXGrOCw0BcFMPRWql9PuYT0NimnMnvsf2niS40dL6zgGZQlX3rhbNdwQFKcyQGXL0AGql
sUiFHR4JDs/Pi/q1vgJ8iFcKZoEkARNL1BVez79aGX5JBEVqBzlRdbbymSyDKTb7pxt0glqtJRl4
KDAtdLF7nqPkk5CckZ5aHBc+szwU4+hUFkm4H5sH4Zs0fnyyphPRja7XEDxuyySzKW/3XUY0yrAq
ZhsrXRBEZEI+fCrfI7l7COkp1/Begfs6a8zD39I2PTCNImz56YxnfsUGlu2UHTA15egY1g1jR2Rx
cqcV5A1VH9fuIJBUXjQ5Rygew4mwebXds7gWVa0ZVNzcROJels5B4o/nZsR8vpCU20V1uxeWyqvD
hc6N8zZhK2jmOT4zCpTESX4tiG9BVufZkvb2i4lx9C0Cyp8BYiR++mNsMnl5lfzfTK7d5GBCGm1s
EA0IySkmRWt87/dYw/rGXu7bbp6enYJWIWTHWuvzINboOU1u0rt4UwKEm6vCLyM3umdW4U8Tm4Sl
PKJtmDd7wvC8/scP5hinCfx43/6mcZfTVdc18QQEcRvzM9qCei8lKg99YdQGddCi8HhIy01qVUy3
VSTWzncGMx6OaDrhCNvyrUpr6GKCBwNmdC9sN2mIVhPJo0SCeR8oosqwVuY39QabG6gy6iNH8lF+
RSvJycc4Jt3Bq0w3uh9WyX8yVuHD33ikKW/zSzW+p8Xm9sluTnrS3zwd7ReN/yUX1rdlxhjHDpeH
csvpueU4QrD6utPxGSmIohaM/qTXBu/2/29JNQyyEXp11UigBj7RzBTeBUQH+7C8+zVPyjSe3RIB
4TVR5ECpJ2/2IogbprqkivJqWbDaP0CPCY7yZxfh/1vDQj46tFS3xwWhjgBjw6lZFOAqYMoqcw2e
Mf4lNPGFAIZhZbNysvM/pB5XI79QU+TT7E6HhI5OnEbMmT4Fg0Kc00AiOBD4jxmYsCRwoFBG685i
vwwzpSyicRW2e9WBKWHLIjna2d1CMIUaB7kmlMLXr9UT4mbLDO4C3k9rSpgWY0GFXBS/ZHDi/Xcr
OJQgnIOR86SIyTSIdKBs+r6Tbgx/2EDuPYrCvoFDrRzlfuPmMM4onBmQbO41zzIuabjSlCl3obvw
D0Dpl7kpHqTdorWZu8zsjBqj1J66SsmjiXilUXJNL9jYxocJOjB09/TmLF2UlL0LhzVBaBghaklb
NqOXORujQQMUqg/o1lt7P4IIUASJ9PGmqozCsfbs3en20kEcivokZpgry+P0+g9WtDYqsGN6ffcY
nrOe7bq/8pVFUgHnkmsLvxVgkjCh1B1G4k/Kb+XOkqQOUedC859GOlPTbUu0bdooAlqsUvZVjih8
2UxvsvedgjAOS8y+XpcgnbggwFWKLVV9c+ALcFTwLTHeoONpVAxVgbJVHYsyrWwlxZTBGKBwn5IJ
+Mdta6Av2HAXXLwpMkgj5AqayNAxQbi2u1C/ioKICQHNi3RJV4FYO/hh3ZPEotRsw7wz39fwNCm8
cyv4ol3N7WAf/XnQveB5NF3Gcx1ypeELiEj4ZNqUQ+hODnSHf6MHl4DAXxY35E3aTwfpbTDIMNS3
yfy+URkRM/RUF8FZbuU+kkah7f3by3I7zRvXbzFGEMONQkjUXC4ztLh2stPZmddih2Lp1GyEOwrJ
kkPon4LavyA6TvRzu6ghzsHYVAZ5JQlBk6BXpbzx7tcoOA+BM9HJ8y/i+DQWQXdFPSpUsDgyax1J
GmVm6M52vwUJyfZHdi5706ZAIeBu1yBl8+eIfUmcHsbyZ3JSEZEsPZBJ9uNF6v7M9fXazgsCA3fy
bpavq0KsZZNU7ZqbrhqlBnPE+UeOJFbRgHS9XviMzbAMihbpZtvMAwvgL92k8anAhynavBPriNm7
V2JVzBSXA4Zpoxd43v1o+Pl3UHu8I+vozpOThfJF2/nhKLAHI3xBBJIXEM6qnhxPuonITeLPdPok
irR+hnRh/u+gNcVGAU2nrkbwBgRIhVrrUDMng1xb75CVh7651pUNVOcMGMCBjMtrA2NfvVl/fj7D
masJGzxBD7qyr+KeE7Sz86sVy0F7GqNX6nQuNqCOEa01aTNdpmdk25Blvei3lAcWlNvaYGfIphNG
Q6Z8wQXE3Kpee8po6jJGZSTY4qeYfOby+PCvG5VCx7nFOVTSbcwIwrnS6L/3xbR3NUCwnVT17oaZ
PYw9CKmgdrdeIEbI5vRF5Z4pVV+noOmqRkFymjmJEFdL9ci31FYmgUFnKd4wpegC1bh2Kr5wUxCL
bnmIvh9HSHrWwcboNe05l6Im2zYOq7qoNqLMYk078yLiGQODby3XPl/ViOybqK2TYB+RzEoyX/1Q
9tIG21S66g+RBhOpIQbite7tJ1P5ANUkNCnesR915+J3C5i02LpYVM4FkSY/tfES+OT+dSEPGYf0
U7sxplj+8kAhES8FSTgdMwqnnB8cOA7dJmpMrwYmU8obli95KnH65wTUcs/mg3fFLp6mrr495Ak9
EcEx3TwMzdPedys/tZXoTguveo/Z9LpRtC2NT+3DOZrIkSRI8c10udI7GyVJfUmjR9lGsAk0RD4M
BRNm2MQvCxBLfoK0+Daj+yjT+sUo2N4952rOph6clGMUl/tWOEpOpiAzElkJOkOeSzuZlb6HpqrE
+jvThNqEBXVqZZxUpDaIAbUv2vrLevd/Sdpzdfvgc44eFrO8lDzDNJaW7Wd8/lB8/tDcztf0hXHH
8YkWkLwd173BZH9E/zKir/iAKn6t8vGrblAKmbuwGhE9mDHJ/5/jLrA3msuu0LfP3eBaHD0MlyyN
c8K36C5OX6S6HtWsgthNAtfaYdoMk4g+NnxDfJhvPWcQMYdOCc1zjdLRdWDIDYjaP/FIw9re2XSu
WYvyayK36hOS4UqD9VgOlZxw2gAiNHlp2MqfgGKEByyjgry7/L9HQtLisoeY+291W6T/XzjRMJnT
37JdIRc40t3zkMDHyruYIjY5CZ4h5hptZmIcr21Kb//poiMxV8UZQXA/N74EM4hpk3wBEQEsL/CZ
80lnZT9x/1aMQq4vbaZkavGJnc8j01FXOhtgyQDAjc6ECTLWu1M37TmlWlpsa/3lePvCtF5IpXtQ
taNd+RM9M3IxgJ8fh1BT+nSEdiX2Szw3sBOs9IaiBQ5OcqeTY9xC/iJqS5oh1okIh76iC9LlhIAc
IPAWpIlktEoHwX1CB3hCYjTUheMJIxBnwlUGqrkKeo9SdBBehum8UaiwYLmAMfiIKnMKJ5d+YQOW
aU8NlclSBHERIKigo1wt4F5wcejzunsOCex/fNNKxgxe1nSFeWHNbEjMs/j18sSHiwAcjp6xJz0Z
WVtrCSNWGPWJ1UHOCl2548SEaLZsQdxZzc6rCsf4nctXGQwzKd/nLcwfKaUwQ75OsIE4SejFYeSb
pLnU+E9wPsuks/LKFUGAe/T6ptj05NdLx1JRJE8XoEmvWZKqHdoEZ7l5wjPmWaTlSH9bGjhFQlyz
aymf/eHAq4iwbDUAh4wZ5Uh+9hwDZWCE3kho88w94qkTYxSkPA4bBttDysb620JbhgmlJ4fy5mgO
TrKep/j+Gwo/7gLbAdCYyXezsKaaHzygm5254AFGdXim4sH3vyqldi67ABoNlg2N/CSGSV5zIHp6
bef2RN8pc9x8xPdIX3rkvQOACti6KyvUeqQNzxam+A03LXqf8gVWhzq7TCJODuh2Tz7Cucws+zNU
m3pi3u0IfkHbbCxiiSvEP/25k32E792wgRtHQVu9GG/NKg6x+lmZM+TB9IW4/fPDYPNHpzup8SQc
FVGnsFPsD8rH+aPAhW7g3wsGZFEUp4dD+VQerTAnGtroJUFfGSqAk2hgAYoaboKVVhyTeVIlSLDY
VH0gbLD1bbevkxtGrbTCG4P+BmB3hq0d6dwCx0hAWCeEFxTQWSTQ3ZM+kxgMRZGP5S04aSrw2I4E
mDdtMSWS8sYl0dH10ASBj25rbmFw9ct4ZHe9zzNN0ei7lXreMmJk1q+PJCuspkt5OBTfwIh/cTOw
4DptqOvefmklpYNCRdJfDJqGVKj8tcvC/uqsHbPOQRv57QVm+LjWMg/CPoXOS5xEBaOKHEDHsLdd
yRUeYmWc11RELdUPQFcJ7GHWOf+vL5VdIJj5pD/MD0y2DXG2+Ozy/a/I65am9SjpYBBjrNh2bbAa
J3RUr/pB8u1nUzvvDm1mQgY7NXGkgvtukmW5GHDjw5aw2TP4WZ0aRKDqiYgzxfiQyks1K9snhgma
KQbn7tNRHyzRzwcne9PnTzB47KtUzmELr6mwhRQo2ufXHRGcrmEOfsEhWDoL8AtP9zaiyWsK2xEa
TnyC4QG6kc2+YuXPJhx2XF0D9khz2U1WreMks5CSDeXhKOsB26HLQRifmmKv3QBwPCEFowGS4ikK
Xle1rRxvNN3r6aRuO1u/BPTgCm45ajLEwV+LJC1EoNivP+txfkKgKPv8u09U7kOQYnp4D7zynl3P
gc4N4OXcvRBQrmGK4zme0W2cKcePvrUkACwzEuTQrcxg/jZio6zJ6Rrtw+LQvrsU97jQneVsdnU1
95hVhGgPX4bAW1QjMNpMTbSohM+bDcz1JLvrKTvVIytaBiZwPzDKbyi26akkgmRbngECZXiPEKpy
Mc7z+LbVO4ckUka/0v4yBHDA9Gc/AKQh/G6WKCyiL8Vl5J0ZG4OUp6/l/hDpMimMDOizFTGoQMpH
nf0Yo/3ZKZiNXDTaUh0eLjm9u3KY0B3mS3OUizvH08cN7mNOf4kkqvKaDDo2zcBOsdibZ0UC5/DM
cSjREGZU/129YuAcgYHFrNrQupTk5+l9wkJhTKQrkFg8cEIXSftxWojTZJUw1oZj10H7i4wxi/wu
P4WZxgXe/s0EGN67YQvA+mYTu86T2wRXdDWzPtsSeyt/rzh0ENn1Mg8Fuik4mhO3R3u8ZHYUrovQ
vlOi+Ds6XVAM9SNCdw0IkMmrlC0jB6BJvIwG5va8I9fJxKb2Fnv7F+luVNkUlgwm/88P/uk24GkV
PLwJXrP5N/+bo9TkPX1U+xw/L41hM1VmgrwzL9AdV47v12RnIT3wXJdGHpivT/2IvFaB6Ee0VQDz
zhTg4e2kvDuDN2pQEY0CyDJcB/iKsC+j2MH9uQ+kgA30Exmx3K9C7AXupWe8udKyTbRrJxXKOrO0
5qecQuu/B0GVzf/ptODwEZ47iyJWl5pXsSBPGcQ/ev+NiBJiAVdt+pD+PN+xq32hj3Okl5VwSDiC
6V2BvtUUUOWYTzhCGW6GgTluUc6Kpo5RrJL5glheqlsLD5il+nyPd9/Hi1JPZCHPuZWaE9PxIWXN
rOzudhsTEi+jqZkXjcFoFjJgNFH/9ps1+9jDPZ7WFqk7UfqMlOxZ7pQSgdDDR+jw22kTvThVMBoO
7UyZRlD4zanSFFOjX09m2arjidK4cs5TwylvDngvYntjbpPC07wWEeKE3KVAG1M26rTh+9b/YCyu
NuC1eMXzbONcUAk7ZQceiNQD7reUowvyXwv1bCOOmVm99jcf2O9JDxS2VZIaqbzLaUAvV1fCH8hZ
yG/X6zMoUHQF3OmJtF2cLTsAFFgSIYJXFrjth2v6OehfdNSvZycVpCE9kRtAnees2wBI0SFjZgY4
8KDUdjtm0NFTvqWS5D/6ROLwmztatuOfyJ7rA6hMkbzgfejIDdynE5L6PA3CqTgdPZ406KYhJH8e
NDh9TYWX1ss+Jdq1Q9BCaddztNKUuYL0vj78GqSQWqBKPXyv/T9nyv/b6vF7s7GTchpRXZ4MjX8x
mNfuJ8/AeMXywP24J8FiftZ7kGidSPcEKWgXiMLOqfO771i4Hi+w1XNCnRbuMRgX9BJBir2CUdP6
FrY4Zeouu8igWrS+6cTJJhrfDgNPNgmIKYWvhn+CrncZKkcl0SDTFFoWiGRcVLTpq5VoJDsBV9jX
LLCerrE7Omh+9a57sGXTCAXPUTyg/a0/ny23tzyCt06jdQkY43lkZNLBhSY5RB4zo9lF9m7oQaYU
WAX7KwpACwPNAdqqTWeCCpmnCwc0Y/lHOKkkE2krlG2twbWS2XmMRACc52DWr2pkrbIID3PF0RQj
8/2bEqlBK8AZt0GnfO7oRB+NJ/kwWtoDoewBlMfV3BGIZiwvl+Prw3r/YnbtDNoKlOM5oUvbuH6X
OMMzhzoes9EzLD5Je6/8oJgDnpriNYZpYQ7EBNUhZ39ftj3ClESffsiS6XqNAnGVehLVDSkTUASI
mur3e1PgXl/vvoC9vmzP7sLa9hn3imA0PsOdwVN/+ZVGVyR7jMuF99XZmQY/ucKjehUwp0r2t9fD
H4X5US5Z0EcpkR1UZvyPUxTQJkV8ExI20m7zT0G5tUriQW5tDFkzAeL/dU/GIdpvZp7QNgVEQG2c
A3hM7EMYoCjKVSw7rnKNzWW4HPdpTWq885WzRhfdise0N4A0O4DqiMQVdMHp43yJfCinbrg4lHtR
LuDPKUzHTSmJkoDgjvRX+moeTPJdGIIVNQjqBH1+8ifnhzJoJxsJbuFG6SLmcAb5io9FGNdvE5y5
TXVRqcvaeIXP4czoiyY9WNamdxORfQ50Bc30aE/OYci6P9Jp8YwCQE9/KCANpjdRapqEFSmOpmvN
T9UWo8lchKqxtHzFk0BEXDeYjJp147MNTH///tkxp3iGPUQKOsMtpNQ63LceuSjg/v25svY1pVHe
dZ798C7DRWrrT6m0bkTrFv+9rUZryBYlynrJ3S4FfWxIe5n3h7/xTZ67lETq+z9gpp6SGyVGo7Gt
I/Vs4T4i2KgzSt1uiPhZ1BQ15oKcnXZoZn0XplcfDOKuSGuj/MMua3E4cvkd5cIxqBmsiIYIPtV5
LVacovL0l821BQECMzuFqYkhaKYKOMFBQrFyKiuvwly4vJFiBFHLdK8JCwQEUBbkMGdmBL863+cB
7Vg9xFHTdXzQbXigMBlPZoivFF0uBqlXIiUpF15dnycGl5jIMC9ZsbPVtzYjvEWk2rBPBiEQLbxd
r4SudcHY0TSNLNKDPdpYti/mlN/u2zlmNdDvA1bcNyttrh/gQInerv/H7LeXr8FMO1fnHGv3Geq8
ONNajYQ2o8Ho9wai/w8nPtLmlM9fDDEW/PVcBLocZuJkHT3hJ0T4pfWeXNsjMm0KJu7yBtB968m9
Bou2Pwv4UNzWv02JWUYjYN1EQvuYOA/GeYymqt0xxl8/wZz7JD0ow5AOGKNptMJJwm3yXziEz4Qa
LQZmkg1touL9zK8KlVFuWU5xMSst2CiVpdrlsSJ6U2PWNeaLGBbqUdXQt1ndPn4BGeNAAQ9u6QPT
AYRCAeRU3zBcnle3duOxbEon7uLxOZLqF4ZXZShNsC6rMSxOaxRPQJBCg4QByg7M+3hzsPFjMvYd
/MS3srUbH2rkjYSRqf/XfEGzg/ml3u3U54GumRgcThk2O57bNAxmemFdKRgiKQ5oFpndJYuu8MNy
V9GaxmskNRDpd/ZXWa2sti016g/jw9xRtENcg08phQBIMBq/A8DOQ6LH0JeponcD0vjiE9TFc02P
mgopG4L/Uw6FQoWMGkhNLuXVUqVrS39bIY+G9o9WTcsOk3yzP9tIq/EAaIIk5hEkshsT6khZtm4z
KnqGuYbWDQHc1kawvwYLPygdPGC59eZPUk+nXpenA/kKMf7nrItJdiukt/8KjroMHZyWZPyynxNK
htbsqIgBdmNM8EbMRXUwbkrXn8UxyoQ+lLLV4viCwzM90X7AaJT+Rt7oz66dJFqfovq3TtqRKqMb
uNHpkgOw96iiLqCC1mcOXyCI8IQSyB4axkt0DSN9HWqOMlxOAGxEGc4vm1oecKal7bW4wYlKM2Q6
6qqo5BsEL4WNrjV/59oolWas0G8eKNqyllBR4eeN0xl+QbKBvmaIKrfECekbztInRIMrGeV90+9d
aMhYej/6kY5JPzFYrgRU2YXPkhQfTTpQ++un0/00f8j4wKAyYxA+pWraUFzQx+fMJeYIXVNYPqxi
uI3nndpbScb8eIdhO1zILSIs1Ggjwl2UzewOWO2SDbJvsv00SLKz0jKXjrhKWVSNPklt4s6rVV4K
24Rnm7qqjzbn6IDzPtI3SXvM8sln5coCrMG04Y6WL3X1vLfm8N2zGVyF5nkfecvDH1lXC+gV41x4
M9KPJAPShH7VP4wu1ip/B21Zf+TcUFxhxoo0AMG7M2OsSXe22o5K/6fiHhfomqbjxnODgZ/MdCIn
XVE0/Gd04MkbVLswKdlztGZXaH/uJrvEV6JyUDGo0Ljdsm/NRV7/qAFjgW1TIspXHt+P5OaHguPl
wYoWJxluasGnm6KQdSt/fE6Akxz/qU8anft/gUWm8hgE86p+I1JjHvTLrVXIgU1orXnHOwdQgPid
4+drYLniaQ/fozAwsEpLMVBr0ZZD5pScQpHcE1dlC9tQaiJrh9sLdoEX3geRaoyeCBXMlpDVC7/R
tJsSjIK4HVq0Q4AMvjW7xQaP5CzFSQtARE+LMWR5kSkIgPvw+lDAw4eWJ+VwY3Ha0wwPoWPaeIaP
iLEdCr8txXLKk+M48O3ffxRF8qHGFzOXHV6KhMSQTm45bm+E3JtKl+KLm8lXgqAMLxkXPokeMUWM
k2J4fBk/LP61Vvszfhr82F15GlPJ+QjYZk0PX2NowYgKJSRrhdTxvsphNgkI9vgNw7you9gbnkgC
+WJoAOpvdKzPoVRBTO9FYPi6iO+vbgOFbyrpNXUYk/KNaor9FHFm4uTfPwJk3WlgchWiTsh3WF8n
P8v2M4W4nGVaX/2Xi+W6gM39nvp19DE4aqUmmltVSMM+tnQT+Z0xXVk6/5UlidafJXnwQWMEdtZi
lLaNLDAPXCGi2vKRttHbe3/W6nbW7UfSRlWAQT4ENXotXXEJu+x+ulXVwxceeBayUnL5BuydX9AS
gDTY3enut9dVXmc/W972j2YJMZO/I4YOJYy45RJPdgzSDq7wBJ0xRtyjfzXCVV4bE6jpsJMdcQri
yFyIX+bno/btj2siUXdwPJxZ9Kj5co8f7OXOgfWWCuywoBY4t8+Tc5VOCBuNTHhY6TfMcb9gZ3mI
Z7vxZGtt6bVfMaVD1EAWTIPyjt+o/D5G99tsCxv+R2l2OBT1tYjGHL1eRZ8xnpAS7y6T7dZqpECJ
kMUrAG84oue525Bbh55JCAkiyx/NE6kDg//9aQDlrwiFjEAbNG8GwzacaYJeCvNWlaymUpftx24z
6MWu5H5LFf54tZyqsAnnQkMNaAzuuIA+4uzGSODrOwxKyRyWRqRDuB5pBqbcY65LkLWa5BS5VyjD
9PHhb2SJc7qJ7Lgj2HCdglLBwFVyefN8mZa4yFWp8srrxVeJVBxSF4L9HK7x9G9vuh0VanMT2/yd
wectysm+SFm/K65u9UYuXaj1X6c13K4lyK4ChpyygVw0TvJ1Li+dHIhSY0fF0wtw+NRvk2R7dfa+
UHHtbR6hE+jaern3KD+xT4CZ/t1E95VZiz6rauotc238jyTpHMhugd+DBIsatk0M1mHQFrSV4kJ4
PKj2Po20nGCM5EIW2DVv7mVTQ0iaMzAo8vLqmRZXpc/+Qxb1Cda40Txws7eNyUJO1QDj7F23HPfy
GKGESKGmlcbKGj6NdM/Ttsc1aL29NCU9wjw4+Ob70HHXyXqJ5cTyZLSV3OE7Z3w3JB75PrXODnX/
PmmLcc9+Z4jhYRJyzTo5wmjuzEsZ+poYjTsrk3csdlzI5ViCwSQO+3j7B2OUg5/2V7bgLzx5UawS
ge0eqGE3/0vBNd29y1Rl0mp7VXwRqGKSkj+3odKg4BqWzpX2smKjgKxenzZX3A+ryqWhjdv0NQK0
HldXKKjMXdGie74frpUZl8t+r1JVOnUTaNGbzGTRtdjIhoCp2bJx9ft5ndnUwyun4XNfjmbvzBKT
n4Jp3+wIjahR7bDLkWG377jH4DN4Hc8kUtYpMA0MCHx1VxFJ5UdgAT+rbWujs1FccrxE/FM4dF5C
io4D5Mx5esBkjMasj5RKgQsIeLRCPqL1BFEOsELWFj8r94FV78Jls23TfmYhNUiUcWQsOWJmafZA
HepoHqcaaXYzFT95AUssoZrUPk0vs2264gCTyzQ/s4TCHh7kW3+i80BJC4jj+6FaCXqBw7p1CFoB
qjB9trPHgPcSn5Fr1xiYc5oiYOon3R/KlkUNXpRdyzWGVkP145vkqjrf+TXIoi5uK3+Qy6k3KGqF
EXLPDhNHpxHdfmjJLGaPTwminkMhztZqE6WXzdS1tNylklyPKOHHOlAnBntIT80EAxKNxc2AAian
p7Jazew3O/kVIJl4FdfPNwia4vteJXZF/8H1qCkqxb2SKJHb2wLO+8+IaKc3G1hKbK/JmhR7r7ac
jSufN4TfgfIMm2Eow8E7+V7JoNvA8VvqHj0UjaZCJtliVi7gOiph8a9Ex4sYpWdo9XIkmlae+J94
7n8exEA9JzbukQOIk/cOufCD+xCF6XWpF4GRGJ1qo9KLISEmk02meA6ICy2/9Ks1JTKz+pusZhv3
FJMnY79ldGVAEH3ke64knlFuC/42RD0Pu6drwdkBVMh1XWT5/DFv+8XavYTdqbK5NNym8tZZ6vR5
hyXDF0kzkR4twj1kZSNA4yVaOEJXO65ITawNc8IGt6JVZHd05B/hTmSmzPGSfw+cnh2wYPgFhL62
MWNLq2tKX0EKN59KCnNljS4erDRqJIOcqDvQw1WH3PoBo7xiWbkxwdsyKgJd7eBW58w1jPDZ3Hc7
kFfaeUCCFEapjgIhCrxPyKof2dYosbdEQa8/9OoSgPc6XH/NRhWckQ7SGBTTn9NOMzCsf0QOCAQa
IE3N9fF/ErgqFsYhHorg4e1oSTsDIDS+xLzP66XMNb77ojz52Kh4jiJ+AMuQAU37g5qj/eEOJ3B4
RqB1ysh/6kl7RlV+W4zTe7osKF1Lj+6l/vAyiktbD8jEmGPjXlwxXQjQ+JyCjT5RaUc1+bpw28HC
lhwioAUovVWxayGxD5pkRQVsqF3TF4un+/t9I9+2iqYL05dS58wHrWevUWn9xoL2tyW70HUl4BTE
kWxjffsHqB7dtChQVUi+4WWNCR+bOiIWRLPRNT2Vqr/Vm1/h8x66TRY6Kz4Uc66SYb0DhK6sTPIf
fk7Z/ICfJ3K7iuQInhjUdHUQ6b3TMOvo1Rqx+PnE7Ot1jqGhkgOKwQKrA6+MhJAWuvAM2jIXn3qQ
48WGVAWptyLn3zM74btbw6pD0D/LaOYATZ2eS0fwpUKX7PltfEZcEKHBUXQzn9gzKIpdFPcEZN1p
n3qlaXQ5ACfNRn8i5GDP/BS4nicOWj2W8Sims5Et4hsvEGcR4ZshJ4uGOIl9tv3Kh7eDGQ71RrI7
O202cCq7HmaG6tCPkhfRBbhQrCx5oKi1DMCx/YeVT5aVIAGwF3h9rgCkDqJ3Qktd51v9UppZN0fS
alo3oUEmpXpi+7VoRh836HbeXH6N14RMPigNAcqtIqxKL7XwvNVHBHJvxzD78XH1wEVfN3YE9rk6
flxhsKP703mMsFTt3gnNunuHREmU4wzHxbhdM5oWClbVxWAYJnGkt0emB5c1Iqm6KecoXjnU202d
sPgBi2bji7+WfVAp75Furaxp1VEyX2/ImfcKqO6qw+oQu9QVrnAthCvBbapSve+InctzM7lfNgBd
2E61worg6RcvNnwTSN0fmuK7oWI79IrYhX4nRINj0QC4XP69Q7dYSAJElVwuCtZosidQghv+SHTB
Kr3ECjc9cvWPIID9frbCMQIxQbycz9cRVQSCM6HHR5VMj9zeDoalyPj/YKfsgKvAv9mKTnYQc/li
eZydNXeM8U70E/vCAkUOaFhEBDmZ0Sz+mc5xvQ+8JbbC1FSjPY0dw6LlHhSdxrFLHCXZf4ctkqF7
eLHmTWQCZb///4pJV50IhZmZpZiGu21GFO+gW1Na+WjkprmkQym10PvJz4iZFJRdejEsghKRGOIu
cwxElbbcLhBtr4JIIRuj35CWhJiKsy/+HB9UwAWyn7MQk4B4MDzwoiz2PvYC0yBB7NNJrQtnAR0B
K22CB0h1sizikck0h6kNTeNhPvRvn3pHvN4Tu+dVFhU3PcCHgM/uK+ED4Hh2T86tRBCwUZy8QfSs
SNKObqeMJzALl6dpe6JGXbN07sYiCM0HfG+S5VVHKtp3xLN0D1dk0A0zR4MNVvLAwaFJd/Gjgn+d
oLmvsRkFQkgfwLUwtgTqv57GUU+4xTzoUo0BvI0F1atONC9saHHko1xb+kg7VmRe33XbdpA7lTbg
u3M0EEhnKsYSqGLStw2IWHfzb2JUZxSj/6CkO1xLhweQHvnEWBMIsdnWkUXRlANub/Ig8XmTTR3D
Id5zPYBl5L/pWZnW+AmG1IAbNaCy2q0jYgw+RLs7l5W9d+p4zFGCxp3wltDggr6gN4kEiE3bG1gc
h0JtFaA42KCvUIvm0vbZQgcImbuDNZLKyA6j1HdHCUkcYCRGpaT0OHznkDTOVSqiVtHNzw2QlUtC
skXbshXY5timv/zWsAE+IVE/2zKvFJ+M+J2wuZO6+sJhgCaWwwHfR15EmKO0IngBTjTUcQKRmFLd
6Sp2inVY7/fl9zGcpIYu8ucGr4vWmkspoVrpIEbBlGyjVidAIBh6+9GjcKVH55p8yk7IDLCP/gGa
YhWZostxuxlbvEyeCIaZzpPsQb5XJJjJcwBbTz8PfFFSHXowWtcC2gNJiDA8YwPq09e9JueS46IP
MqAuhbgfqbAMoQYlq4011/b47JwLnYCY9zOmB7a3eF7coj5E6ABDoG6OqANAy1NkxZHYJCwVqpPB
xHI6tbgHaMlRt8ixQc2Yg0DsZ3azkr8Tz0j5j9jqFsrGvbICazZU+M7Lbuc0jfaGlEIjn68xWHo/
poZp+GUjlzcr2xF8XA/aMZ87mAUVeJDFtanrWbxaoO9Yz6fhLl8INjF0dzENWfHjrzdU8VHg9QFC
9Gb9IBOrLHCx5pAbbCpHgdE2fcbNsgQQJEJQh6Wi9lpWnUKqcqs4a6besi54cbH7/NoZoxi8nuLF
djPrKg0gM/SRMgCu2eeO8YL66EZAxytNGEcb0f3CwJbYY852SCE1+qekiM0Mm/ETk/Kcvmg2LXlX
wkd/vsbEC2ywNqhil69814EZZQ2C9DjnaVbnllS7SwNVw12SZaRFpbkHjuIWWWXWIf3BxcvcnSKX
JG8ghl88IfWEfLMYk+dsC3d6ou6n0QHHawkZGfspcQeIKHGBJgN2t+2xdSydW8YHHC5IWjtW/xu8
rJc1gDncPtM6HIltB7bbiCBIlOxNi/ZEmbgJZk/Dhny2aej3OAPfBEBOl2EIc7855e5OebjVGICO
RqDzVrH+qvdl1gR6gcRxZ1gjlBAFEKpnaijzQrVVAUqLpOxFOQ2HDjFIFeH1miUDYzeO4/yWT6ny
hZZi4zgt5N5Qmxc0KB6BX6ydPG1gbR51eY4cngEVSY9yrttX1bBef2+O8RugFZQWklX06wONkbQk
AeMtlBIFkiXvO8RZJ5DJFNpwIwTeou1gp2Nntg+QKmUGYqUqYxAJcyzOaP3r+JF5WWi0/hTVWPEQ
Ci5VCx3lHNtY06gIDMN1V5H+e06OoiWGh2nocOSlrYQXNek2mcfoZ6+my+Pqeu0yyIUbTwagJuw7
SyKASFH2q37LeomVrKAi0o/mm6aoJHT8MwY8VDH7R4brEFWm3Df3GHdRiumnys7O5jOcnqRADzAi
UmwLeVoszedr6UA/aJ5p7XS6WEn98g9VceLUEv+gHjns3tZka82EFd/nX4v/EU1L87+RElXkH9iq
7/i8EaaCuC7C98VJWxxTqCbe5qgeyUpjmIJ6hV8Oh94T36mlCJ/paxG86bBriqWY/W6SUvRWXiOe
e0PAIPWsu4oZ1VKhziVndGpSs+24OJe85afyGUS9obMbtwtERRk1mubLTUSJLxxl0UH8CuM1FE/1
zAWsVq02ZCVVxY17U4fqyZOeQMnoAzGRn6U6WFbkcvGwwzmWpjjy96gufeAe5R6Iw+/heFm1rc38
7KCiOjzmIramtdS3k4/f3uf7KgemBDEh8rWJHN8l/PfEakOlxMRno1MTlYLYoKYMRTiguD73dLcA
B3V5UcJRncz/r3NjRF31UYZscsUoW44aPXJ+VV82Tqtm9wHtsmHkOnWXiiAdEqjP17pCie6PkjsC
HC3u2m/Y2QcAwrAVmI5HSN4SjcHyOD+KPAOm3J2BXkaYjVY/Fe3rDDbglvPLnqktPEfQpTrcBA9+
0+nc8HPy228Lag2pEfgNRIHCxdDTbBeauYcPH47f4Zg/H9XIeUcASucVS+fmJXOO+sJ/flz7BNm0
G7zIjn9ZHbQSostak3L3ClR+oL/97Y4//Xw96z+dnHANtqaT7W/hYT3+rN2FSmMJ4oaKs7juirFI
jpK6IbTfRfmeFAm2g2lfJSqGIMV/BH+VPNQceVH91fY+YR49tlWCB7gowL1xYCZAT4ienkj1YHOm
ja8x7QZR4uD7eaeHKZrq13UFFHxneF1FIBq3WVjAXwSjkQDhnkoMfJ9uAgo4yTm7071WOxqmTJSa
/vB+OBGJtOvWWvjYZHEdVGXomsZJ5uTAQRHU2+wlJ5wy3BjS3Ri8YxbXtwSVfBKVBQ7mZ9xcrH/+
XWV/7lnBRnFclW2eX7q15b78xiiFlPYw22ojwgVjPfeuN24Ayz5XU84rvc7OlHcbdNhsrTHRXhII
tSgOPQI1M+vgySzvJgEhYU6LvzqC3oxLyP4osXrBBM4a+kELhhi6U5emJYw5PwoTbDxTx55J2NUD
wwS3V6fFylKPy3IODLgEdqFtJJEA5h8VfkzxB6+QjcUBcDbHxL8tYOWEW5oMFrdb8hYne2PaIb5E
7BX8vLpNBEH5LuqncH1RjbM8lmABqoDwlswRJojYSAmsRT8OdYxg7DmYYSwUkPoNsUojjCW8cIzK
8tOjQPw948P4O1IMN6ijAHMvfuQ4HLaETguE9zBpRSrnNMZTat+gh5rCTnGkvRDb2u9eUqBsyexD
sjLQLkfG5QAXEOXfHXanDEGzgerdheEmXQ/tZhh2XbzvYOz0zVY4K2dBTNdGegE+ziWC0COGEA2c
gzZkjA+7nW6zVY6kzxkJF9cqqOSe8T0oMRSLt8BwSf2bD2xjx/nANGqphU2m5r6KjMgD+WO9YB5W
Qwljjszl2esk3YDHUh++K/t8GUiTuBIJxZ2ktzIspZ4hq4/cfsrspkZFGJEHUyd8YeFdXAa38sTR
n2xXVwaTSpP7jNVqu0ZlTm46t84rlW9wg/t8dzSOfBFuF8YHQ7nQVJJPhVLhg1QhY0TVO8gAuzGb
JPHh2mTva/41Iys1vdw1xgKr7Hlhy6N1X7eAm6eQtbrLku+xbY6p3pHyk2UoXCIB59BActHEuN6z
ZYdxsvnL69ZOMUOdibizZti+2fo5qGjpqseE7zAgTj0BZ1TRod53tb8s7ko2Ceovg2hBpkUgwiWl
zJ/Sxs+UwyNFqIid/sFNMz2OdKtX44DJVPnhbQN88gi7uJ1h2BF29p9XxQZFUib9RoGGk64ZmtQP
lPNUwpOEC6zD7y/cT2VT4/TYKkiMZPyA0mpZxtYlWD/b+ySu8/JgDjlvz3Yw8PDimQlt0ttZ1Rae
8KKCeGQylZzvEL3e4Ebd0ZpCmhlNgTpyLlKkSfrmyuQYGD6uwITreNeDLnXKlO7K155co0Hq7zqP
ixE565ZzvteNBBZwIFJN3nu/+Nt6kxgqMO6wMLTaBifUnhZTqYebjwbKQATDWAlzPwKHDgFm1x26
rM0EymEU4TMl5NiF+0Tcvw0nINMfmQcp5rnUYr9RMTxJ7RCI2hUbUH9Gk2FLG5Sg/1FiycrNbCx3
a9XT9Wj3dupazD3y1FhxicyefTBq5uR2i5UXiUcH5fI9mubzB8vutX4DH+47bhusoJnzEra8pBf0
JIQwEwjC+2TMQzqsSJl/gqtuGNBBSpE06qPhGcL+x7yCXi9IVzI96syVcMWmZLk18SmOJlSyMtdl
cjl02G6VFFEox14pxgwPILjFkQ6/ZA/n1ZueSXMPBs5Q5Aov2L3nxqP0a+8xh4EcTy5JsasUr+83
cBAOkBzi9m8Ct6fkwZQbnI59svRR+RrjgRXhGgOpq+SR2Afv5Z8SQNO/KfjLaTPLOAbaup/rDJT4
/B+pD1qTiSfMaTziSiA2esrISqfzK5tj8xCtgPBDGVSphdiGVFcn0z9YQQOj/qxne8zXqdHi1iVK
AU5zbMz+fP2dpPGn6OQyskw3AZDaYyLQpp9RH3fZ0kytuNfPbr1BHxOIfzvtnQ9CAb2dMLA4sIsB
RCfv9b7aOQ08RuaRxFEmIlrbkAlapyt4BrhrUsNL30gQaYNdIzl58QtmCbRq+j+F9WYK85+Oisat
Ku1mL6PklrV/vSgNa6Z0bea4jzXnkqBxVApKIZQ30RZhUxsgv+qiwGX3TG0PZpeg/V4ZSoOkhRHe
gfbOslxd8NbD6Xj4Yyv8HKqpGW1U7KbMxWhS+GQsboIwUUTP9bJvBmDt8QBitgIsPF87ohVfWEyI
lA1k5LkJs6g1qlGieOEzLlL/+Rszcebk3veUxvVUl7c95pcDaiGoxs6tVhnr0uE9vo3v/witR/jF
K8S64NL3l2omDYkfv8X/Rafg2K+3iBZuRuEGoS+Yq5Im2o9NtkmqVpy5ANBH33CG+wOrNg4ULXkO
3s10AlvgeGwL2T+cscWvEOnPYkUS8dnTX7ZO2ACrsMfqAc/tXU7mIl1XO/fBCH/xbA8trsWvllbn
lqXCspXPkZdNwfhegLtadGSEthy8hpUNGEkaxGXVdWPCHsxzVrYEcAd2uV/cJa74rW8OwAJ+vL6j
xNsFDl+TuwSmK/AuGZMXM9S83eT71P2E6EruSvtVz1J5+p3YwjuJq8/o4uDCgkeiZDFFmqMOwdfj
bKqyfSHQpgUqhj8eU0Qn5dOVPQzQs3VQkQt7Q+RnnJBlFPE22L0npDCRrfjDW9rXXtwXZ0qCnYY9
X6MV0ifaO4p9yb/JTwJkr3FZllXO6c6WfZKUH2X4gtsQaQbVkmIxVkk8ZHb/mjau4bMewXjDov9S
dJJw85I7Y56QaPQ5vMHJBhCD26OAymqHIantRUE3ObzDF1+kKk2xd3P4o+bWratmxjw+nS4toDVS
+ziMK6/NIErBDNIO4kgvWPeShcNlASn29/GSr90wV1A5+R1HBpn/ENEHoeIdb25dVC0iT8F2rtkz
Nu87S36pyCPMQsHNi7e+BI9EAAEQvel5YSR0AzJid4WkPQFzS/0JJ9SeVYlg/CQ719p0BXFkwei0
ViTwVvilduacN+0LHkZGXp0BK2LV5FU0X/L7Cb/yE9nejF8HRY+2U8/WDaPKSw0T1Ne1KIIDP1dN
5EDRPL3BnY/MGnULA7EYZpL1eVimQMgsH6FMoCVtySjQ00kMD2UybxcOskomT3HO71jyTUTT4UBT
AdrF8lvh2SZ3FvPH2uZa/LuyBD0SnaIdA9BksNh8eyhlI/H9Ka+lP4BkWXGUIg8wZJLxeF6LBpSQ
JNDyrbNUB5V/R5++kmx/CMIgOtP4HTZHYyBfPzRuaxboML7NiIJKX+PFJOaiAoM8vSxbgsBVd7eq
kMEdlNfSdeiBDkDx1kODRCz5+f6qlp8tleak7+J9//WoDOEZj0si6vf+sg8gkPY4frptUL6IsNx5
QQtNZFfh2AZWl04z6SLyZIoF0M/c78T3RTbtAMWk/v4Cwwl8A8rN9xrJ2pQ65LKpngkds0lI9QUu
OrZIVLjyAtaQrEWjs7BZtAy6t9CkohK1fu3QfDc2N58pCLEit/n9mzPv4vX8NZJU9aPQvimxI93e
83al4gCXL5dG6rjuPThLSNZl7fL43CeWSajCCkuLQAivzlxYRqZeTRBMEAtkOwMw1n9PsKOM5t3E
toLotL94IQIgNvXQuu/p2ujMO2Xc5IyX4FMdzzEAnjePfUcL4g5f7r5hrlVZAd2+VhSfTDQ7Chfu
hO4avxYgBo3uDEpEXTaDDfDsmiD9AeSGcuiBCWuRw9J9oIoifCFoUOxOPJltipH/vs7JfG/AlPLt
4eEzmvnGXvyFEwTZT70DVtkWqSUq9kOX3AmlJv7TOjS7/ukAxXxAsIJ18JIxV/tFPQ8WR/calnK0
FecJfu13XkYmGNs46iIIJp2Wg8o0wSN9GQdCfGG69RW4kr10BheT02L5184h0ttcOtXQ2/P3J1th
+dXK+oJSJ1yKIVB1qu2ytm7hIMwq7d6XFX072cGwqFItqGvbSula4d3vaANiQkkZxruCnU90IiWs
jjR57xcJBTviZa3NhQ6afSQIXk0IKccQG7WAt0G8NNVQIl+yAPhN5+6L1Vq5HsNR3YSZYCT6EXTB
TCTalQQHwxHxKPAha/a7GH2l0WPGsyEncob/FZHtIzEx5djd/x44ZkFz1bj0gq5wie8WdPujk+hH
4N4bN7cVBSDDA4EB7DlPiRRzNuyGH7X5E6ONEC77uyHJsoFenIppnewaafhuZ2PJ3YBQYgUcZJOK
anWWyrTwprfadC4kxkUx5n/6f8ZmIfCDtmRRSrv/Ggj56WIm0l1hDratJlFDhgiugeNMzuukhj2k
f0QEu1hBGxZOanoprwwWEBZXXpYeQe7muqLmizkamOnSPHx/mQ0BWpwK/5ep4yfzDjuxtRIn5wMl
+rme028PS5MtJR8N6l4227XVrh7nxFr4dpunV3j9FHY7NPj5zk/gOB8QmOlReIfotZ0c8JNjFAOO
ATGIWIR1iDTpOxkNivO/c6q3OGqPZ7L0OCeRWbrLDMIY1xdcPCEqnlOtg9OllxKhtMD+9j5Gn+W1
X8BW8AzgdPmOwuB9TDA+9/lqhX1a0JNjoYewYr7j0OenTRS2AuurhjKHzWWbyKxZOl9rUUqknCUb
9rJJLnUj859XZc78R39mfykHAIYVc2LcA8gWk44Zd8o3ASTK3fencR2ykDq6fiH0+cqFXbq204Jx
KxkytMXJ9og3SYj6ZUa80B0dXqjVBcY/alitDQZfY2O7OvyiulpxKfmMWkj04NiNH4E+KRmRelcp
sQSRsxOTfUvMj5AplAhW3E46dEB/T8FkMa4o+WdyEdS5kxpmuqxPQq0PuvZf6o4NU4lqAEd2Ldh6
rPB68fAF6OYyExWdusbk6vSYB5cxOcSUasAHV6nZOReP+7ho+AaZDeVfkbV44HjDYqQDQINuzvJX
wH2V5zKoxZxxVVmMoSBUcKEVk87Qy4185jxjCgitFIjztqVTnMHffWRbQaZlsLeONWEwv9zRXIcK
v/hkNCkh9PHhwUA9ClDbzAO+aRi7zLuuQ4oJukiMbGaUafgREnrKI/5ajK2P3OBr7dklntg1lsVx
IP4iymsCSYg2DYGlEBOrAEOcFKvJ0F37ZQDBOLRJ3AmAG4NQ1iS71lczbgvmMjigH8OgIqrv4xpa
kEwCd75UQGNAUN0s7lZOATscwK/7xaaXj4PjCqBjn7rCDZZRILKVxRDhY+tGWEcr83dT7lDMD9Wc
9aeJQwRQpXgGrt1ROIQ96Unc+iKwtU91zYqzqH2T4mtCR9VLuBBnd3bs+YPc2HPMWbF9eVrD+C6Y
6kpzXiFtWeUeYcelJt5to0q5OwmiogeMucGLoCfX57W83ltJwPo+9QWRW7IzKMKItM67/Jh8LF5b
F+oc8MBJmS/7Zlq3lsam42GUvgkG/ZXIdvJPT3lDgb/EPhawEfzHTTFYjp8dO/7CidntPPhne6r/
IciRcaUVa7zu8Rp2StgGl9vL9nduNmEb2uxsGtKWtKtIJJ6ISkNAgds1KpVBUP5I2Y7ZGJTFYClu
XOedyrXsvDDjSxIMNy80JDEaTjiEz3O0wLStdP4IPP+RjQblHDQNMFrtRoW6DPZ+SHi5zzM6Uw89
NCmdQ97ALgZIXmP9fbWJk69guzFCDjfR64OUipVQpXlrg5YEuby4EmABGHAItc03FlAp85Eh/TMp
5C9wn//SNh35XeFvLp6N+5vE6kVw5GBeJrJkXPeAXqyXfNWQ6U8mkN/VpqiIopBEe9SISoEEBa2z
SWxnJvq7P5rynf2q6kt1tnZFh+pmA+OmCPfb+BTxDE00Kcdho0AVlDpuf2AjM8JSLM53Fh1kAV8q
6E23pZisbfr389ngp/LRzmsWOaksNjdyy/hb+hanafeypF+6um2fKJ5yLdzayVAc9BqyonF1gGM2
3IdsgAD4gT8bOc3Gw4I7sd6zQ9Jl2hRoYvF1fmuWMrohZFLGorzMsm3SpGz9jUPhTS155ttj3C4t
gYl8qCmdTDgpdcVTFtBkw0y+tlFPvTCTGtsOwmGW2P8Tk7JkrB2okSI5KhKWLn8YlAvnIjILkpS5
MGxxG2UUWIQw4UEKmp00ZG97AqKHd1NF4PPVgxRx+Nr/tEJEFE946Yp4XWTwoz6k+MEMjbmND5jc
pVcguDKfzvgFvn/X2aEMTlP3zIvAmMgMM4PpK8e8TIcSywEChus3t+KbXedgloDtjos2ypqI73oq
XKOmhi7ts5RjdYemUzl9Oi2QfvjEV5owp5Zn1qtV+t3vSXzBrXvMkkluPE7AxGBCjY8yA3yG4DsD
DnoReHmfdllEKVh4muv0aKmFPRhSKb2NyFiLgIhyZ41z/Tm1vG8bzy7enWfsMAFp/1Mahmwvsd0N
E+9ahvf8f3xkXP2VHqJkzWbrxcgQnCUmJxkJtq9r131JO5M4uYr3jAMRhCW4D4P6J7R0QBeQLCqS
hjqMegTJN98qWt68IBt5HirptxnniJi0eWnDEOY7gqVgoneQPFAvzCeUyDHJSn9tSDC75tZvcPE8
GgwoTzBKYm0CJlANEqKf5y2ZRRm7AyPd1tVeksZ4MA9CC7NpQtkosgVyIiJfY7a1AnSHRLYy4idq
qpw/hWO2j+6oy6vKc9G8lNjwA1z3dLQRGWZ+IISPSVu4SukkTugX72fhljLqviDhn1G3jrD+FJTZ
/X3HnfKSfWDU/nvK55laUIjLe4E0Om/mTO58tdEDTCNPQGv4Yt1lTtTV6o9mkDVYlsX5rXzAg5Wy
7BA1lTLSMIx2a0FimsJ4+XP0hRWCYQBXM/yjX7iFfKt42WrFlSt8RIdsPpZZEodlJslO40sdaa+E
7wTkVGBWHEu+qTtAfVgKQZBaAINyHZqlC65i4OkrSCI3G3HXSiWngkshJO5C+69yPXXZgL3UZc8Q
COJlpDA8L1bsC9/QJsS9WuT8cExcwRIcOhzsp8ZMRKjQVhoeJ7ZTcqDM0KuHE1dhj0aTbZQdOYqf
MMiHgQ2DmbPnsnXJAs9SGSu8+7qitRQDhtYjme1yLVHrWtwN7U5ZYMBNUaHv/3I+kwrJHJbLVrRh
StWy4ybRpu3ONxSgd6LsCmQl1HNtUScD4m8KK+qom5XA4vVxdDQTDEp3uXPRb79Rr20U+kGhwVqe
OE+gxOKsrPc12vJ0ZQNhY6gpEu1qCwFzLje4IRkgvUmzZuCMHhRa9q3Bvex2Y9VvJWoS+l+sjNGc
pnl4Ve2h8uss+7oMN7+0eMVLmvHMIhQQSQGTGz6iWKQCNE2LLb1ltC3Hjlq+Cclw2faQqV9hIvOC
AOxXlJKwh8onZE6VGUF9MWY0LPjIWx67ChoHjKTd/uROllrSHhJye4aItQrTtx8E6BpNLLjmYlYs
BTqVO5z4RUyX5X5hVdKHgMjMofl6O7ZGuV1V6gP/UXVlZYC2lxepr2kQqIz6NTxT+75OeTX3H/Lq
RvcIJgr1h1dgQfMtZ9gJELH76obutEt1Xh4KlENrxAiGXfVaj49zwvW8TGuBFvWRA1PNZolkEKRk
Trd5hdla/5g0XccWNrfgjLri1a1KIoOnUmNmptC3N6zLHjJcZPwX8ufjyVVqaN7g3/SY0YtuxjXQ
zHPxPci4HHhgaDBEI+37+5znBRmFo1+YPeHki6+YeJWPLzpEzX6541/3e+ONtNwx9Eyd0JQBL+gs
N+0mDbEYIo4cBKJiA+mM7gBvyhM0/pOIzjJfT/ILvigVFsvaRWDeVhcUTKXI2uCYvYmM9ryyKgMp
++FE73jGATplfMIMh2fIOvzAM05X1D2rjFunwK/M1kdmHyuV3w+dFTgQ7wbRXOKCiK/TKSz3vlcA
Q/C+hU7N+IfJSuNgQDu/NXMn4dolLkiBjNPVIePKSxKW9gcAiWqHzSmdc0u0gxi0L2bsAJ3cvGuq
EZTIF7LCKtbPjN/8hf88OuOYoO6oipfhZGIOBIAua9tq6dO1x1Xfn3uU/17Fp1U9uqTluKY8v5eb
Yi958v6JFOcy9hzPwQirFo0upI9S5ur5FyexdXk9g+kulbcOccWkF+Oe5COOEnu2uC9y8vVyPxIp
4y9FfQPzf/vI3zVBqh8SHbb39rKFsziBSg0EU/J2UWxWiFLF+0ILkA+NE28UlVObQcA9M6UBTmXm
0p0eJN2mD8N6Z/TiKc6rYUoDNsBSAujmk4dTTjvFMa1VN1+/sYUZsA8O5G+D47Vv2A5IVExJ4oQG
3yJEn5lu8C3wTKefxxSgY9zpLVxViGfSXhGLYz8HSjj90/edSXoHMjf0rwCN85OVD6STSR+81S21
nxT56wsAwPfQe4mhnl8Qg1m6qDNT7J3uUL/+PnqZHITlWBUwe6Bk3HXU8uBZLjQy58dpfJEZJ8kS
JQk1vGdz5gfz9VG0qthjyqv4qxHZlvwFD+iJWDqHr/e3a2IdfZczjzZKCA2dXHjwEOFN2KKOwPJ9
GGX66epmzd5XWk8CvPzA02OwbDRAz0FGMYCU2Fh4CzzupudgNm2pU7/BQxaTSVR/+iOVQv7MbR9j
oEVsxkSwCSEY0DywjF0KAPCWBTzuw0WKV68Cz0L2KRoi3ZNfHDZk7iRBVROMEPG4tudcOIGGjUni
CHlGHq0cy1qT0Wt0GTKqB4vfLXKsEMl5YjPbW0XsSMQLPypf3enBKqEyaZ6MlKIbGA5jrZmtxsdw
N2EimEDZuxenOT4SCHbPnKSYhkC9UXNF49DmDABPo26hLbrY5RruUgxipRRfabSlUvtFlyM8FIgZ
9hTnnLpIvfHkCpDxTydY37r3RxEo6ob7hjQUsh0RvwMC/Gr/ilJO8rPJlhzRA384/9D6f0zprr4Q
BFj2qZP61XmX1SvFQaXEJzoT66BJLHGtwiEiHwidNVa0I5NoJYFJKpEc8fZFrdeg9qVsQQMI0lWd
I7IdOxzqKHlCyrYG9+appiyKmWcCxMc94dkAsJb7cNMkQSXdHxccA20aRcGSb3D3BKokP1hN83QQ
7oe6RD//ALqBMmki/1D6VmOirOSKVKO3CY8AxX8DATKjbUy28TN6aU37pITvrya9bvPuAu6ZmBQq
HNsHHIxRDSoL6S4llV8TPGqtaBCmfP6WV1c+yxjp8+bL9Hs/StE3lFFdDCZ8RlLgiZpw+xd+DnXZ
2ZFQPavgKBtmZtpvnLqL9Enp+gSFhWUO+iF8/1X83jlz/q0h1mF/ggBC68hm7dTXygKDHzFcoM3E
abw1RtVvRywv7QM0t0U3T1+efMORSkuTbN9EZG/FU5wJCK1OiQ3+beWC3zBOTvhA4U8yBpo1iQD9
uFjuCT22oDME3GhnRNstAZQ4du9I6AXHmlEBLQKvG1vNIv3xpHK2xooETTTZqb6/rxa26GEmAhdu
fwK5K6kZGDzl+EF8vBmyYIwvaEvTk4/Rr7rjG//KfjkCC0wORuzG/XgnX+/V7rVSDVrfycegWDJ1
h1Y4vXYFbnqRPy7u17RRCXuVAlo+bFFbBoCNK4yNipd6Tm25RhibJc4gh10H+nWGTkPfAZvOreFi
QIMNHxQ6TlPNmV1w+IENClNS5RIGXLrq4/+pdxHGXzIFIT7l8eLlAmTFAID0hQSxr3WwaWa8m4Rs
48aCM3PfgU7ciaARwQIkTCbpeAU4HGZkGXrLG8hUeh694ANRioxv9dgk67yADt/pw/9KXMZd4Xby
9pxgv1ct+dcCSGuXGT5YGbNDf4IdxZPLqPJ87hwxz0dXmT8mCj3ZIOId4i+yeCgdKSjhc7nWEDtQ
Y6OHfofhVgp6LGZ92rDap+gDX+HeHyl6QxGRVab7oORIQMlDNN1NeYAnUBD40xWh2DCfPqn+Kr1j
e1XPdEjo68a7NslrBscWbrlrSFPS08lJBdvVhsdSsHKTwUq71m9dNK9pwJq9OrHxfqIOKe/oCyJM
jrYZ6XPpBjONK4aKrui1y9DwYpykrpRZdY2eWebrccm7yq8NxuKQYM5R7N7v2+MbCLQ3iqsa1tE0
Dn5cjbWcua+Wkg7CErHDHsIfK6XPc/TeKcG8j32ozgvHO5Yw4DrS8CyEQQ3TOZOE0Z3bhznWtJ68
VxxbQ/0SAGoTp0Kw42jrVFhaaCm9k40+ANmqc80sQowMmLDaQZKabtJO+LVFpigzn0luBGlUXPxn
Bg4Vm2w9EA76tyxM/PVnV6mEF4FrFlTuClsf1W5Zn0Kd8QdGkkjXTmcSOsLqoLgywbtATkWT7+un
oKHYeOQkyc9WzqjRJSH49q4NgRbHhSFy3iPna38iwbrVZm45h47Ao1o0ZdwEj0BmivQbQZ2p1R3U
PGByhKAwgb3J8HmtOxfzKLrJUnfNynDQpRrJstA8L9achYBfZ50xeZfwgYjD/k95+metYRu81qoe
SztLxU2IYWg802d2yme4HXlUxhtgAzKuLItpv9puzm6yeg58Yk+FnxR6be2XhewPRz5CjT5IqdCN
FFBkxKlvr3kEDC2RNm/HM35SEOT490cUxElUROsq3JO+oQeustPmciRGunZZJi6A++zFjU6g6WEn
oRN+yrbzy7o1Vh/0D8vdPZuiGOmi00fxVvKfzMXNdx8V5dvX7l1TsQKDrfjVphvMRxnygYpPqs3r
FXIwk0AIOVkxYAglm3/c0CZtJ71R4aBIag+uZf9CQr9sJYEB9Dz54YLOp+N2ZBWpX0RXneHml4/l
UX2qH4p1RTbyMbHTSrf7bdxlYHmPfaNo6XcDPgVtrBpVaP7jKNuV1eV5LXUOZr39NDJ2M2mzM8WR
FwoO4uc0/v1dfhID5hBemeZiEo3uRF7hN/9D8hr3ER1xbg9wKzmEO9r7G3uC77AhDvNtSA6ZJ4sS
t2Sma3HB/zvBtXUwscxAmXs3Mvsdix7MkJfChEFqHjRmFM6MUe3VoUIy8n8qKqDO2kDeTaIEuvTf
lAGc0ZKWqAvsJSTNHihtaHtj/4KJEZJhhWS2ciB2LC6kBFARppNDSwBcJUeszZQ+qeGpb+fGeNef
mtQ4fOVaDXNwRlxsI7ByKOilLD1KCOeThW+CPwsvJrfoA009YqK01DJQT2dMlfZtE71+0md7zZgt
vW9dB0VeWyRxF2XinQpiZzF7EQOjWDT6zQqSTedUyC/ceyOs6uKQubftI2aukq8HTEcmJKEhqRsf
x5q4z/aRYKcY7Va1C27fx2NE34iGAsoT8hDDXvY1hSU8HV+/ghdmEJghixFN9rPOWj86QSLIrJap
qxGe+HTt46EZaZ4Y0mOEvbQ5wDP1kWyEQI1gFmGGkIj6KQVYP6ZkJIqB9159iOfgu8y9jpK8KRjd
YQ1tDIKFUmhDX1cVqNcUSN2xul2kDHY2EwtpRHlrD1T7Gkfp5coZI9Od0sMa+izb98Vgec0yHAjY
po/qH/EmIGPW7KwAP2kStn12IRkseo0nyBT8P5R9bILinSxjgRqwSkPOHQv8682fPlSAiA8+Ghhd
bDoLVscTA8nDyZJ43NgLsn4gmdoIjGcoKDIrUGdsYAqdfY4RFw/FdnDR1BzkaS9e77Rd0l7brf0V
xVU9+gGfkljS2wOBSZUJD5RvWRWzj4B1TOLqH7B2vuehFmcfc+Gtvr9sI45RdEgVHDgfjmTssmsf
paySRtro0K57eXtlxpKTaXEUMGOl8MIH77EnQMD+y5z57O5tsQ2kQlJRMkJEiZ5o8IcGYd+3XsoY
/i6wOHhYbTYn7qaEtdKN/7hNwRqAX6EST3hjdtqEzjeCBT4Lo6jhakcOS0tiMLSFjWJWXt9uIPKF
GoHmjSpSZRn7Cbfiu5JKBEdC3f5lzso08DspX6jrNmqCaAQVj0/T6w5uvVSh6PcSA7CrQjOik83w
3jI1WcKVuLqTa/9kQvJSsd4suKil+Gk7M4o7NapD9I7nUw4sw+yNlQwa67eVASPHnFwgCfWO9sDX
zZEP2IuCfB9SmUJ5D9e/5knearCef08GId1P4M6fOuehGBKsFjaa04xZWMEFsdZ2RxYG/MBJmO/U
D9AuflmRT6UjwjIIFsg4mHDPs919qsVZf63vZm9DgMhG/HcLFuwGAtKnYxRthPVHR4cW/AfPH/d/
DLZzkU3+0yRapXIjiyiX0L/PB7FKzeQB5kqgy7E3S5K0IEeau2o12RK7UMBxaKjWwzBoGub7HcxC
UkO8jW0WBHauahAelP9JzT3uks/h7NhNwj9RrjrQ5QXYPg8kKClKJ9HYlanX9/AvDn0PWwaBVoQS
jNw6jCntJQiefqIsq0a+kB0tthytPfk9f2+tWOvEeTSS6R+ZUEB+frqvjQO0hnk+G6K5qcVS+Y9A
hwo8r9eZInjYVnY9u/fLFAIHfE989h+8lCj595XoBtEVQ/Ktblc6yx0cCoDzJD53T/fL9VJ7ybYL
SjMOiX8ldTs4M1hHKf+njXapube+wtdaNoE8fI93Dh4rHZ7Hy+TRy1ij3EG55YAAp1AfMVSdu9/x
0ntEoOUF9HbdipeXyIRo8JLQztyGK1qhXmNvfjD2jSRtTnf6EqjuMeP1GFbKBvc/m8oUqazybqRK
+ziaiphMzV6Jo0H1d6CJJJ+0uht3KIxhjplocJGi45Ov+GdAS0ie3CzRxzpmlJ2P7lWLg4f1nVXo
GlyiageTbfZiGTC5lU6ZZhoHVyw/xIJbG5TD8VXM/+rfAInEkOxQEUaxPFAKZLW82TyX1okgtuBT
INbEIYUvIT+dwtXJODz8OgxoCx8e580Y5mqxHsQfCK2Wt+jN8r03+xEUa6IiRrZr5/DwovF0POhM
QMuixD/NR29pzhCzpikctuQqF/Nw4zRlaoq8tUMYQq1ccfhTl8Z15Yw/4VjQElIx7omolM9ZOrGV
+2ckEhQeMjeMtpmUFoOZ6k40EcnIgbPzAQJS/kjISqsGTKF3XSYUolZMvBw8UM/MZU8kw0dPwm+8
gj6yDHCoAm9wiYEOrZ29OeINTqeUkYQOkndqZzIlm9L3Bijc/nNIjkrDFE6gFxKpgaFJfuKnMRj2
xgu6tXEtKXc2hj35GnV2rSD5jzSmh0S70J4FpiSE0JssgymdNJUFFyEgCFjg72/zL+5ChlS/ESQP
ZhNu3DowhC5V7twB06j1z3o2c4XJZWUe4JsQOi6RZ/9yH14DdFL6TlcNBfXB+weDbQDoMHZ5iDz3
cvdM/CLXuheOVbASlJ3eHEe5XLybqRjDsImGHJosrVbiV1ousTXqNJ2n86J8bFuJVggv+/dv6Sq8
QqJkRKVPyU107/DiLcTb/8bBXlqA1bka0qqB31DejiUXelDSqL12VLcSvqdwGVx9iEIuuERYHydn
jrqyFyDPMOTA0WPr3Zt4E2V5WYAYSw2OxUcbTOZmVXFyreyjJWzPYSe/DIUizYE/PtLWLSr3n04L
QiLEbCLl9hancQYDDC0OldabLKpNdxVIUno/GgQR98Awzemb3z1px1Wsf6OE96lszJU7m3rMpSd2
D11ahBeMhkhDqsWvGyTWEDT6iu5xxITu7GbcN9VcTRc6mxYgQTbruQ5oFwhsffXEpCtd/SEXrexJ
jrsucwZXDBK6OfLtNrXuhYDhOUvpogPFZb/jl8OpaKqwPHc9PgQ+MAfPJ43pJKHiyZa8SWN1PolM
UiLR7XQP5Zrd//SXCdoLdgx0ogD0TL+rq+ye/AyfDSZ0mcCXnZ2ryEylKOgc/e5URmz6X3v/lnT0
+UzV7Gy81D7x+WLTI/5RucBGiblxMjy+iTKUE/iucvefJ9gRmQmeqHahphlOF4vk2XuGKlnAdWA4
EgMvMaFIT41H/Szws4E7SQx5Dj3IA+BLyw7rxLA/g1r3B96A+Bg83jgJ84XuIFvDh0KKJP0ac390
yoHtWCNtCElFxbottlJGatUtyz4ZHz+F7A6kwAPYVw0NaMmYgHrKnnQCVXTN7UC2jDXkCIFzK2+o
wFzN/dVqMwH17+2jUTudXqnXcJbw5Xj7nrVD/JLJJxewh8jLlNn0npGgPoIOofdhXh7dZTZh5zjl
Xu3LC5PkDzxDg/4XZJrXZ+U2z7SNb2u9vTwWw6Xazdhqqi7ZMZg08RNhJn4DaAUMf5jS7JB+ZQIR
LdgbAhISwRW+Z7ed0cnkSWMAs0xuoB19v84DEoWUoS+7dvirpK5MUTAlRvB0NR3iXAl1XMZFwAnQ
i9bqTzt+WLftTrsy4aBYgy8SLi+VH6ALC3zBAUVPKMe+UbZZHvgKOATQwCjzDHVNCGBGI8hA5EzZ
DhVWE41sniQ4DxtZMS4QjP65x1WaHK/T1wKYXz0ZxvkxEBGYVKGsgcoC5jUaBT96tsCqLcUrY5EM
WvxtuxuTYFHRfck1HU0s11t6vcT1sLjoY0PldZEj2/FlOwiZYpuv6OoMrbq5j6iJ9o7Qh0PcNW59
3CkrK7y2KiV+ruBnnBf4CUgt5iDGUqx0ZNjFH58H9v7A+xLPJMhltoL/L9TV73i3B9osMhvxBOZE
y6lrCT7napLcIDE6MnvaTXgTzLfgELnLj+YdC/4yGwVR2J4Kp42sABEOG8m37UUtPSBi3EvIiiXq
mll3NDsUvDj466spPFKxvNT/CG1LWaiqYsYyJDos1IZVcn9Lezw686BdFbxh7Ec8r/GtVK+wjKg/
JlBxQIHI4J5W1tb+KyQLvVYJPJmuSFecQJBfZEpxFHWc1C0tGEMX9w3YJi2yevnb262TcAn+hS38
p0p0lYwGYl9fDRn8kcY+AwOcuvXKrJlb0l7BiqffDr/NRBk8wGkdeP2PXgLLSw77IFnX8X183I/D
J1uIyVCcqeGJiR8NY/W8ryDaXEgCm3+5rDI1RHYtaboj1Zub/2nrKoGHoLYNtP0MwUBoOXS2CoSu
Wes/+28xGpVqFSCu1bWTnVjd70nUkhJ5INo3FF54TGZ2HPVg2dYqxV2zvISyyFNrJY0p3caMBze7
80CRiNCmRlthSYhoDK6H9ScQInytkUcVqVgxSudKQnN7hzCvCPBa8ISlJ6sUoRzMt3ZsRxp0qGje
f0bJl2utgauc4RTQXg6HaVkrf2GgUVQ6ASVicfG+4W1VzVlIKcOwvVjXbUcO6O90pLP2sog4FViP
VQIkG458XfuCAF6ZLidsewtlfhr32oxOufsjepGB3Cp+sW54Lk7Xb+c9RmR0zMU1IzPUw1tEOPsR
OjWudi9BFZiKjK2aYDS5sl5dtLg9I9Js8r5s2lowxC/QTceGJgNmc5ajShLB9WNd9mduZUoWmn4U
YJ4md+pfdgnL7UEJikJbyBtXhrxkNtGfAu8hQkIx+HsT13DHceHWWW3y4sc2P6R7ZBnEPEbtAjjB
rNYR9OajfK3KiZEJ4Rr2H6fivc5s/D9H7u5+dIFd9Urj7kicHKqzG46hRyEV+aDuqNAn4BZg2Wb8
WbODbOaeysGOeFkn/avBifMHYa96fhI8CiyUD5ZHu3YONLhcA4qK/F6MNQ9E9THsZUG2jWCCOZ6D
8CBFm+3wbydNil6vMVty9X9hkxg9zqIbmf7GM1vrUR7fD1KyiprxizE+KYvW2UDR3ZduogYOysw+
ayQtdEnJ56cbiF8Nv/xxym7cxEOBx1S5YRDZ4rSpJBsSpLN6c6bOmPL3hThTYtU9SBu9oAi2EOSv
VAJL24KED+KgBgM3LGw/QMroQmHR3sXb6fyEETImdgjqPPRi+M5nh5vytdWGjtxBsgswFkdshVIA
1jRmofWsUjP3xCydjpcY+mMKSPLfXcCUneKR3kerIIvJ5anzaL1fBOaPdloiU+kepUKQKdIIW7tQ
KkNKhzFE9mS44W/7cZpYMJKac15rINeDrN185vqccy8tDMq3/Fk5qB/PyDhCEBeA5+nO+iPqSkLJ
9T1jJWLRRr6BavjM0OGgGreFspYICjjkkLlwy6p6fCYEXap7uQgMFQT3dllDE24pJYPtOlxv3Ias
+dGJoevIWaiIpPKoZR8ewshKGD/LxBAzVz0yC65+cPnYnt1f9bsm8flhXER9n90lTs3TlAiK59gm
8RS2tK5ENrPC6yB186zOaKs4txn8Do+PKXk/XjX9rb32WFNU+Hkk44TipVgIWkzRz/KRPSLZqe3G
ovW6twVEZPoeVZxIvXqH9+y3pFTFoM6AokmrGsOTKX1ZmJ2iFZK8hN+CIfmMLZYlePzaiUx5SagT
D7n7EmzJsdlkRTJvrLe5RZQiSo1QBMtjHYy89kVPJAYFWV0Qx3H5Oxu72xFVyo/N4AClg1F1hCHc
OiTK2r5CTrKRj6nR856gCJCezSdD8EkxJ+u/wbEz8hH0UFcW3kJbGexHw3EhqlV3PFP3zu9IEylz
mhRj+xqTeROOmFfJhI42AqbftoG6Ua9kfTCm+UvlU81eMNxMue2BGXWtqR1ugJUjsxtUVI2iDcc4
cqXp2Cwq2uMp6m/rDbXxWiC+3h0lpF30dlkQ0WFUqh2H9CxDM7/1ewh1SMn/nP74UONGpOOy8s+l
FdPCb5rN1y5KfxSifPeLyZMxccYjZZAromCrczkFYnwKksLSLAiNIXYbKJc7jaSMBm4lQeoSgwuI
JA2mjdGI4SZuN/OMlD6D/Qxse0j9AQ5bmfCB3HOq/z2rwMml7bPNiTTrmJ0V5SQrtx8+5x/7nN9e
8L3un9qktiT4HQr8kO6pmZr6761xcs5ye7mEYbjXHEbzh4cGmCHs0k/PC23V8HOYcNhFT4FRZbkI
vaCZP4u/JTt7zMOIE7XgoERjxHbcA2U+YjmDzWve5POylEl1xmrXcdZuXj9gBPuK0ywhLwB9MkYX
gwg/ofy/mYEYzXiUqD0ZIyi+LqSUHleh+2pfrziYVjM2ViFQYX0AYHuWa9/nTp61tVcXUWyCXAXc
i+1eUk4RphNFlm3MC7DTQeSe587sxQne1/jhpMC0dhZMZy32jgDTVoUR55ZGJcHv5c6PX0XiWPA/
O6zf9Y5EmJt9CCEKYfAH8+Tcbzyby6+UjSMOEOhSldW6RZ6zhUiYjSzJkkFJYY7s6iw2C2VZE6Kw
KLz6eU5QvoHqmBQyFBCDI/ih7aeQdVEmvV75uxVTBdF3nH2bdS7j3nTUPAFqPD7beg47dvpm3+sy
gYRfXORONJ4OB+5zDpPSO4rkF9btk/s3EkFvsrEIib/+ngK2KRcxprPmmmTsQk+KPKE+e37xacmD
FIaM0iMStUQQpg02U8yamdIC55Vht8WWOMbf5wOLvEPvGJsDEDWTzXoDbfBccSmchtr4HTCkNAZw
VN/Xep5n1FmUqb1Ac7HzmjycE927csicpWt/YddRk61y1EG18rwZMd+RqVairzMRlkvNESIXEG1G
a6rcHwNhGVmMOdb70rX5ocbhThmqR42NQzVZPZuk+4Tr1oSsZOSTN27DOorDBNigis9HUkIsle37
MmdCSpb2bdrMO15N/JF21trUGHb6PfU1oc863p0/A/+/VekUz1D5kUteCsTWrGDs2AxA/Twksech
LDH7pZmNsPfXa3DPLCtz8h21GDiQviWdbNhVmwu45Qgv0GCD0PUhZVoj+AxXTnXH0zajKQjimZJh
p4js8oBkf/FGWehptGvkIqf3vfwmh4TYqPD1oO88TTn1VOttgCohcGfiCi3eR4l0ky90SO9R6lXm
gvo1gOMUhCvalz3J6sanVdiYEjRGz232oE4AQVTRi6lYB5FDTiyBNug9anLy1MT+QFu6Krre99vR
M7gtzmp5movQIIN4LfbZio75O2nFNvdS+V2Asj4vP+KOWxVi1OfDWCBLKjtfm/PVk/QDLqis5z5i
yKiSUY3gfsKmYAqui0OTdaypsEbl9QeQbHYa/+TFxpiyeNDSVHoIuALu0xfKGZf/7xPbD95qymuz
Omm5sR7JYFxjiSfPw0/43MO1yzoM5FHCxmS4QEsCYuf5m3TuAJQamyPgLcrMqzxfSTV6/tNC6NNH
q8a6mS4f/E3MzRoCpb3aB1ZqD0oseUwImjZrvrFOvMzWkfUSw+QZ+fFOLtuGZATA9ZkBJkwK/gJq
tTJaXqleGjqAujaEqvsY/NtpBFvq8nV15Jm+wdNrN5Lym14FGJfQedc+xr8vY1saYHSIzR1XXeM2
ujw4VBkjJAJMR2hOVpIrSbUFNq8QGU5fxeSummvZoVTEjws9Xvc8R6sUAIjozXT2nSDHHETDHn/L
w0oDgvExuRE4YNIVALsOhmMhDMW5ohIRSdids1Hp12gCJ7TmztIM8lH6qUuQp6TY4FmQ9xls/vTn
EPphpkdsknwVnA0uXJly4k73dt5Q6mcg+8qbf0t5oiazR36ggnujK1LzJpWYcWeFizICu+a3cQCt
aARV/2vhqMjBbxkpBYykppcWBAFQPR3GSUnNme8Akqiv1vN7SkQCuJGmAq/1XzHhQ75r1vrU0ksH
ZhglrKUVrabA5gRluETDGbtqDLoG5QNHbzRvohTgNKQ5fVA22xZzetAOoTMFJ/5hAKdC9JjFGUgP
O7/GNI1Ea1PExe6HNiACgNJhl4nSCSegIq8QTP5afPORKzlEKW5F5V0CYsrBl0GOGwiwW3dbh2Tk
CvBvvkZ470c3T11y0etoghW8NvceJTTcSjRZPJIh2QEth2WEY69dOilvczPzPxtPM1f64io0QFyA
pSQIpyfFAct8PUezJfJjIQbVaQtDnDmR1WM27AWBKSYZe/nmAkhD1SnqRFcjTqCpceK+Clo2mkwj
NNpggenwtngk1QnUKqYclWYhua8dbi+0HvUb1NumCJiDsH9hwoNQybI6Yw5YlwJ8q1dIMKOU4Bjl
8FQ7nBkFbYtbzlR+i7EYuQVPFSgNgC+0unabRzRPt+TB0fHiThDGTUEJMIcWV1Fn1j7UzYe0ew5v
vkxr7Ilg7SitmEGlQGHwH4cZ4Q2SLr9GHnWCTyOP/TkKOT9laCC2M0s0xrMGqg2Z/K/G9k6dHVqc
pdCg4Il/xgD+r0UysBqR+6xmmRMAxyU+BF1odWfWdO+lF0ALX12KPjR4QIHBQXPRsmy6F+3wyNle
oNSe7Cco+k85vNFqm8A/TPwLXF7fkRwHRB6DMww504qDV7AdKUxYBUrD5mu/914SrFXSPEId3ZdD
GPvX0eK6zosCHpmBo+aCAyvPBES9pxZkIUwB1eXvhFy/xwVziG/OaZgCcXUrsF5yFyaAlJhmHs+l
GiB8JX3stijAxN1j3Y0pDPgPpoBX2aidtxhEr8KhHS8XirgUAJCfSQPxtIeTIOKjRU9kHK/apBgG
ksx9OspIrPofsDycjLZbe5byD7np93hsz1tKyvd6kCuPFw7+RCbYWlSV4mJLzZWa/v61WA4If8XW
i+RyLaimAz2Fks/m/lZXgsrFNQlrCvoKqWsw+H8NUVPUQJmyrl4POB3KxZEq7PKiCexpmZX2akxJ
xA9Y+kxtaFqNCDXfsz/kfEa/TrIBEetAaQLbWazio+erdRne0wQ0FFGbLl8YbwIF3jVZfFBet82B
7Qt1BYJ2VGr0ErdLVGHq7TtG5ChCqqutTB6HiiViqmQPy3uGgk9Wo5y3KBAKd3kwp7dIUk4R+pXV
FrU9DojMwtLeqtiXow08PiNdR35mZzm61lOHqT7BngGmAntkMOiRD7fQkBllCtNVSfxfjOM05syt
Wi+E5W5vlbfY5PSQwYgHWf5E+oRDna3ZT1F1bS69vyTBidPouFuOLVk8telXk/jpVara1Z2APAdQ
58MouSq9n/3I9e4Pa97o98oWNZ0JMZ+LtiAZYm1RD5UIM7fN0osmWGIF3TUb+gMK0ri/fmind25z
GASXnzCfQCqfM23ku+oG8DPRHhSxtB0A1mmABInocCV//YkWWeslDeFX59yVdBj/a06ObEnd/mC9
syYiPP6vXo4U2N6wQbC14VXCUw5fdSKJIOk1ww5Idp2jtLq1RVbJLcOej7O/Xr5+Coi6oW0B18Rd
TYLJPbwZ/WVm9JC6ZBqyAlZg6ClER2nOJzcj2FFhBd54Ymbg3Lrwgb5oehFQPm1ctAZ0ZPz/Snc2
H/+JXt+afXy1MQBEfWgWZ9vx68cBMAFlsN/vKSuiLqOLu6JrAtFed/yxI1X5eBV7XvEi46TuDO4C
0PfNpVNVF4zrEk5kW6WXb/OiHj4X7l5i9FO8Oiowd4ScM38X4IoqM4oxh08iW4Mjit07me9WV/ho
rn1s6tJ2PqJRypvDx5yXJkIzJMsi9c0+VcibH2bvkMfNfO7KCcwMEFGq0ePY7dkVofhll6Q0w1CB
6HfsdRxTt0HC32p4+8F0sqb21W2CDRer6wZdZxMcLbYBx1wmyE3at3ZYYBSYmrMzf0Ajj27oAwdO
h42OIMo5A8k0L1g2cCRd3sUAq7XO27nHfF2XkUtjZar++IorRVc+F/5NaYVg3TTcmMqh+e3VQbHl
L8d0FkbNQVZRduhxvUVYI+xvpTCGkR/Y/oPFLEfNl8PT9CzlnZ0ihRNHFw2Rmn3IbxWrU0ix5HB6
Ji1m/7mRjXm0pEjDikAjOzsobVUPSheUvvHRFTpMKTx9RoCdLjdJ3FG0CCQAoH/f6D+U/YTxjgRJ
6Z90AR9p3MZiKpbKpoP2RJBNcBxq44SH1ibQucL9RUZqc684S1hyqzmbUuttscWZ7YNH0iVNADO/
B8BOVVhAwLpws6kIhzX7HIxNobegzgyn9H1Ho/x/pAyIHK/k+eyhQsRQfUz/zP6GDvndfIe+EmCZ
lHapV8oL9yvfBn/yAuZXZmagobE2fGPEcxtPRnRG2Knrvh6BT493vWTjO6QjWZ+ZXzl5jemEY8EW
mZzqbi7Av1ObKwdgIGNDy4hEBrzK3GLWa9LcknoYMLyNdA7jCCB2J1BzltNIy/swDIF7VsDz5fOf
7McpitndZGOpsTMHGe+BHk1IlSruF7BVUyClqQswgLz5kpnqwNjvYpKmAonQbF01NqXN1iQpWIwt
a6EcT5XJAL6tvoIDg6hf6bTatrxWPHG7QVAN+4VwSo2G/2z5h9pPebHB9H9hhbMCKfol+FLC1EzT
AiwOABd4YJNVu6kBScqCGiCwDZvLWrmEwOrEHNFBx8HNLnokEzPndFZ8Qdrcgk/Cz1QbUzwjusHV
bPDvZCkpYXL0Ke1zI9LoFh76PD9W9spQQAt2IAMUPzZHc/SfF9Nt1Ko9GdJrMygBotqvwo7zJRdY
Tmznpkw6UnFaPtDhCYY++ms0dylPZhuFNyJmIl/4dVgtLAoAoHJhax4hhv0Esmb7kX66YCnuqcHo
Jw+OkTbdEuL4/tRoiAGHv0qd5K0YPvE3sqTRnyIL/OBjNLeUov/7sP36IcOFhu5CZLoyvKpdQva9
lHsHEdgise1zfg7ISLKxcKxU5mSfaGd/+QSZkX2Fq+qr5cz9T3LOeN6knLMkgtyKQB8uoAyeg5hF
4qaqIUf77MWb/KlBGCIGjCKTLi/Uc9SANdeavIqcBsxbazM3y1b6BaZZcbxjbHpUqhdNf1YZmypb
ZJZdQrNsVDwJ02IiLFrUXDoSWVgJQOHKq/2b/zVPyyG6/XDFhYxTtLPT0sGLDdmfjAYUKWUZuLys
1WbKTYpMAAheANqtXdS/ct7x9BjAplqksQX+xgD9fWK350QF6+x4gEoqMq6S3zEJyOcT03qxEZV5
8p7W/AncegFlJL2pm6UlBzQp+UaxHK83kp8lOp6mJuF9UR+uw873tUD915HUBmAkEdRiOSRV7gWe
BhIGlhfGKjjH1IvK40kURcpArYynqWR5KwAhXzkayMIruFxogo1Mo4JtvMzXXv7FKaVd0p38JevA
k+xJgK6m/xu0/24XtAW2V0o4cbq1biSZzF+xsGKkwMTWVi6FJTWRky2AWWI3eOWDPrTmYwZYEIcu
hsG5g9csK+j6we3cQrZi2iyOAQKxgES6VgKDR0IC/Y5iZMJagEyz76NmP0IeM1RNNNb0k6HzcpnF
0q5yZ57fUboDEuceppB0g/gj0D0Xa6Waot8odR26JuaN9tupXmmQB05FudOoY9RaAAYUy8JhOZ2E
wSmcMWMwzDAHAk+JElF4A1iBLrF0OlDm0eSAwha2+hIezTykZbObZ6g4NwLi7esHlMuBeiSlGCzZ
XOEqdIqP9ufDaFui/a8k3EMO5/qBXY8RO68j8RQ57spFvrYidp9Yu+mCRxJ2NjtqkbAYyCwe8l9J
5gjnVkqou4+GNujt23D2B9ER02+d10iiW4J3gal/lTJvLKySbekEe4SmZN0OxgS3GsbDwhmBQNp5
Ws+qBRTVhuokhfTWeTKpnguwWqIeHEjZt8OFLdH4DgiN58pf9PUHqCL33uShCWl4XwC2fBq0xYJ9
MetgsuNzvM9/efvSSRjy9hFGxH8wTp2SXXFdu1ByuWqSRYTOLZPsh7wCFdApfDLxcIJ803RePzbi
AO0yZAN43ujYVwl9sUCviPhvx/KV7Qs+IdrQl+IEcvvvx1W6KPPKA+T740ppVN1KuqPqSxt4i8Q6
VWLjPMFlXav8/y1QZj7NxbsJWSeRKJ344+ARpTE4SW+EaRot97zi8Oj0h3asiFwRBu1wYq1ORVUK
RVD9ffOsGctkOdRgX5d1loPlCj486X4qlQ8jwwmBxOacI1uBZQFtduCZ2NtqunN6M0JIK9UgihAW
aTulWr2wTRe+LF8gmQHfwpreLwYWMuLdDaVIkMycrWeAH+2dVWLc7NFSwaZvRAxxm1LE2Js+0i2j
enRuqI+uXc5zxqObnwe0ywWHlGxFZyQoPYu7wBvdLFvgg3+OO6AXogIC3NFE9QUKY1yt11K+55lU
QgEGMQV7REuzfTYnenBjWD+YuU7mRpoYDpI97oawkYXYt6yxSB03Rk8QylE8b2ZSS9MbTy/yHk26
sD9xu4A2WabZQrC3r/lGD+ldJZj76Z4mnlQtp5YiXRUbrlwwd8SL6dIdi/JknePvAFOBYHT2SXtf
yzsA5drh/lIXVWDsMgl7Gut2e2W45TH3FZatKpONU7JJwFe5BkcGCudSdKs/onfn/S60CjEf/yes
dmed1AYPArjtGE6SUZdUWpKdROJv4exm8D081rSJfD9luRFT3TPKo/5IFIKazV4ce2Y1reFY8elj
IqKsNPnswa9oYf0pKfaf83rc9b5vpUXvBeK9tcBv0j3L4SKw+Qb5WfUU7TGdEE9xM1+kFBb4lpVO
zF+faZie0fh2e6mRSgYfTDygo1Q76y+vVzzOgOTnFrl7HZYTklk5eR/KcMYQo/NwxvMV0Ld9kfq6
5T9gIf/VPdwGNiMWC2QnjKjr2Z5wb6eDqoq8+YbHsPN4oFbZa2vs9iI7uHtskRc+rm5cEzNohpqS
A5KupKYoE7lmkbNnLQ4lxE2ZSA8rdHOb258oP5gVglmaDNBBy55uCTN+3mOt5JZLSMuimG4rXQDB
/mHcK703N+/R7HR4+T3Sm4qw4Ruk4qKnVRFTlvhmNgbsBzeo55igSQMzRYuiQ5i5hvo3vbfKOBCL
+YmP+qc3CAgEuDTci1f5OzQ0zy89LJl2iACwFOi6ub8I5P2ZnUxYtmsLf6uOVBKrnUeM0+YcLZmO
Z5PHJ/pggG8+tDpp7ooeFksMgun6SMl+SzSTeP7ehhAB6AYBAR5dxHxIYJvF5gZV/cG6Su42DVVU
8Mv8E8LRxTNWtCY+D7wGvBFoxzA0sLLfdRjYFGHES9oFrbTxGCYsCdRoXJAGr4uoY/7vbD558D38
FujEcdHt+ZtvRU2zyetsQDlj0MSWIKI9/ujor/4om++5D7CJFB3oRVfoO3IXowHSabSEDDDz4bHv
2AK+Iv6UF5UvNPj3gBCm7fxFbQY5hz9zZIfdq8+VNadixuPoGcuKLgLgHlNOXOt7a39QyJHSJJs6
EH75DpF+aThteEAvGvXFdqyroX+TD+QawSSdzkXVLoVsQ+jtNM7KtsLRf99OWG6nSxxw0e53RU+W
eeW52RIlcjHOnQttS+mtJp/U7uVUcFkshyOO3kd4lCn8d4jJnf0LgKT3sxbQPadgf5MsfeorsTHn
PEyBgOMgVgIj1vMbHKJ3VEB4I1OLSDs/EEG7RYQVo0AS8JbmMowWwkc8bc5qHrgtAsUCbjGbsyo8
vQsZhi/PSunEIPf/yeSThoRWzHRGi/J/GF8w6fljKAy8bZyHcmB6KS6VDZPZ/y9yZuEDqXwbUzAK
JlWgZ2KHFtu8ovlopN1q0LB0Cq3026x++HW1UqMxUhA0Zw7LJ71ksOUafAKCGKeGx7DLGrI+Qnlx
JEp01Xd/E/6c6WMz3Frw7YUA6xIyAmjuolCZoDuiLZ+aPS2BW+lXpz23Rn9wgCVt+9govq+Y+EJo
pm3z08U1JFnXyorVM8PoiSqEymqS6TjioT2c6DOFJSJP+TodPPV1ypJaUxP85AVCRbAn+jTQyMaY
2FpZh/4F9fTCrpCXYY5AWkfDgXK7in9ShKbUpMHwQ3TBfnyLyjNhFXHDP8j/8wBGXUZB1eYJ2a5X
gsReBFiKRW15wdzB6RJhSOcIr7VcavDPEzkplCXGGjNuZew0lk9dO4GcZwwcscGuSbOEpGKIkTVN
o9uvztm4dzs1nirhqgdEIz/Wn5FHWWjdwwhq4LDYVbseH8AoDt5ifbAEvoLAyi+oaDyBbz205Lru
hgClXKvZcPQqB5jbdEyTdqQzpaqBMrfy0wB245kLD9VARAn0BG/SJoZQMpLMRW8CbEsunVkh1dYj
PgyhFIL6hmnrRFe3hoLhGU69ZuPkVqR4Lx50gKFPoCt0/TSWD4XGJr1CaQnUGAPJn003NId5RXh1
d5lvN22ilCRIyUFhc5ZC7kyaRfZI6LyEJx/2WEgW50RMNHnHPiE93O6UJFvvvQ3dxNLrc8X4xx60
idZ+oD2+kb4ZKRh5dAMN/4x2JCHpSOB2VlmHK04jdfWbMhyC05IZFeBLziJLpDNX+DtlvF9BFPGu
KDKXB01g5k20MPQWmmEjDy4W/dd8H34/flrgaiPJBaW7kXYgDSLfJP9wLLzMsW7F3IBFzZBL4auJ
khii7+lZ8NTg4gkmXLYha3sqG439nHyxMa3JlbnKmHu+Qd4SwOHnA5dlFvz2zzk6/vEvvp64gd7u
xP0Y7Zu+FdP/q81rX+zcdu/x/Z1v616NDFMfmX1IvLU/gtXy6+wgA7mTkVV6WihiJTuqUgWxuEmE
Z+yG/F7N1No8xG0KeQQqs3zYaQVKNOTvk3HMnibErgURBHVrNR3OKZ5OQCH3LyMLRx5CbxnFE87f
IX7Ab6J8SgX6omUGem2NAUUqedWfnVm8zi+jp9jS2+hSWaOG1vms0weLxD1lFGE4/fCK3VSKUkPC
Akmuh9fx4drDwPqH6fi/LFUkY6zXhnP8JQvcZ7MSBmTzqIJJVnMV/u3w2ykOq8SNaBxDFuM2J2VK
Hs97Dg423sigL/o5ZDDFuHJ0ie6sp2W+tDOKvid/oUtK8yTg7XPCIvurkhnOoda3UVaDeZm7f1KJ
MfrNRkksCC2oLvfZ3RZbauFWrtvMnz1eRvOIHkAYamX+kK22MJQpqac0cGS644PBLClyUijvrBN1
ZO8ogW/5pGYV3rYSeEVfFSIS9ld2r5cdkL54OqEs3Xo0rRXYWQJzVKiVQaaFeFoZ86hkHOe4PLY7
soH2QL460JR4b89vTyVEU6q7p5ZQhc4cMzkKH663Vttg9/e1gPUXA8OaAS6scwq10wAy9PHv72q/
op6NpLZmj5tF/KRuPBYdIW3nmaEgxNa41HueOXZWpD4jW5wwTSUW5+Phwy5zU37LsJZo2z3rZh6n
QwYtOKAEX79IU09vqosbgHe6RecemacL7RrDCFFh20gAz6PomIqYFDjAwfNcniY+x/UKZ4M5Z8aL
Wq8X+Rj4HD1pMcWBPooWFx+t/HT8FOzBpNoe6VRu+XHcOQhmJydP1o0ojTO6D8OvqMqx6538j5Pv
D5COHAX//WiVca/0aHPbDzXBGx5dbTYs/Ar13oZzX3w6870+rEJtcOdV54E7A/haoAbL4NsrE4Tx
TLV0e7LJYG7ltXHwfLl3bAqBy7Bs/l6lm6lkpanNQngFPpxAC6EFxYSN+IXs+ncA225ZW8qlCzki
BneqfAMWL7KnLXVOA1qKJwcbF+VJXgUtyZpNh5DSvGvt1bDz6mrl4zrLFLqdeP/jh6aEqoj3WeSo
ByVQpf1IuRhcDEpvqTzThjVTiIK8KGadPfHWdZmpd1aw2Ck4uqP+83F/rwqu3rT6rBzKC86UFFJs
Zl3h0cfcZNbvwAS2Go79SJee51jCND+fs6818aKH5ottncrAv6JwZx37qPwIyhdMmkDF/mHQetX3
viNcOMfg11TbPJzodlsuRsYsmD096Chr1Ueyj70eff1qC6g9QAgHFaPAt+dhU8Em3SrjRTQjAALn
loMM8bfAI34WyAzLFwUXsq/lFuFvTh0ku4iiiit7V5bEGr7P3lSeV6M4ss3t/auJFjJoYlQ1rMSr
1WjaxW9NPOzjcQmIdd3ZDfgBsj+WKMXtxsdnT/ZsVplwvwmWg2kE3WjTOp7GWV2xQT4et/oqrp5F
sQiXpH7hm1ud6r4qF0d0RsOKztyU4JoPrg9NOVesDDf0DwAb3GajBKiWKbyIfyS2F5dL8wSveaHI
Bpa3T2PwMapgIehg3+9oeHylJ/K4GR77wdoVvgKPElOoNfi4JasIvQDJ0ws5UGOJ9tWL83IFIYkX
eieBOK38/a+3I63GiR/Uynn+onjSv5mxx9+bIZNRHwPA2o+Q5OhyaDUxS61pmqD21kjvnQVGmtHT
EoOx3ohU3hFyXLerJR4cox2IbU8ip95KgV9zDfsc3Ea3GqolOF/q0PKtp8ZqRV7RQ+CdvQwKwJDJ
IJjq7dIZp5dnr0fWKRoEDqoYHFX6nnakjSqRILR+lPESUbtZfJDcU8KtvbjSIy5crmTBBNfTwBEB
qigGxB4oksgOpxhZZf0rHktK8gmxos7hzQe/5yyfusjhq2QBPlHLIpYmBa1S3LA27RLEaA0q6PWU
Mcg33K03e3gySPJH3QqSnGY1Gvw7V38m7V5NtuRM4tLK2jJ0ZuE/ZvKl1HNKcKhTCJ5glwg+pSxw
pklLHR0PAEo1EhgLi3bWB3QZLcsh2xKOHeoke29Zagv371d3JmqfyB4Z74laJBSJ73uNwznxkQnC
tzJCuo32Q2nkYUBQP5fcL1eJuB61XKpfCNfwRMPuRFPDvUWGaHfqxaS8G6ZH+aOaJQCBc4BElv4a
Dwg6i+gJq9QFD0cgia9N8eaX4njtB3u/F3AVx6035gWQIAolc3diyPqViRCVO6h816IY0jPVXXiA
Hco/BTZMOaJNAnbQefcmsAmIN7PhpvLSzHgd7JCWPONNrgzPSGe+CPFxBQsCoBwdflSbVqol1lGk
tEPB5S2xSljnwgRkKsftEk3iGjV9Xf7Z4Lgdta3MugGvIYCUzP2UKzUa0YXxB61qpE2gAi/YOJeT
T5slxECJgAlSmTQH3yY3YU4C8R/znE+UCumafUZ8ovCFW+67k+PG2BhIBKEK9LBe2hJAfLA7w89D
fqjjvGuvwuBX2iD1HwKst2xuunSrRcCOezYZIvvR3Cwe4r4WOkYM8mlO0Lv6/CwlDqvelABOCZV4
xCrcR4W98/hFWsPFKlC+KAfJaRMHyx8YYgPM7zbvUtidztsysDCHdoM6ViZUK04q24K6PUJNYlwS
0PAaxtOjPXWvTLF9EMGOOaKnwHqpfLWx4/c2GKM8y6OweXWmMEjggft9I2VxBZL6FKQdNiQEyfCG
5DoBmmcuphgvtHwrIyTpoE+zfW+faw74djt7rtqd4VvA3z9INNVvI7ITLx9pAu/K5HUXrn4A7TPw
Uq2ZBT/m3nVZUfha+PUx8txUL7m2IDbL5a3LU8qcWCKM0m4qdU1wS/itLmUT3XwyhyUDhmiVQn0j
qyV1+886X1hNy3irtpK1RjaTFpd13dMV3ErBk3rfZ83vqIJ+x/x3uJn2k3wiDRP8LUsOMyduquBp
8jra/ZmPhoJRMPyk3a2enpoS78FM8oQXd9Db5JOPxe3aTJPEWILmlNVirSrvWvtyn5d7Y+Vh5pmM
9hg56BGVwhVLo64KHpadu4rtELNsqRZpHvn5ugLOb0N1nM0H3K5MJYJxozme7VWjXxUXBL5AiW9A
UWLSM84ayBy0IM1eX10ERQyqgGfh7hqVHN6oNy2GUCmVaSrq3mHK6UjTZE4wr5MPhNCZ/uoXBCX3
Yh4kmlJgnRxhVCnqRPV5hLToTwp0xrehDUfB6kaKPw4LwJPG4a2+uriRbYhizM3ZkbOVJ6Duv8fb
LCiKIb7NlZK/bhxYifBEK7bxThLq3mD+YAt0+s9mUBc9cVYFTCWZxwRvXxD+5sbfFYIWoaFKvJob
MQjJsi8Gx3H+Coz5FUJnwJZ2hJIIkqRMt5HwGGHYMjyLJibxEaiAttTlQLzj2L65aFw3/zdCuj6p
Qv39wXtUzAw20klriM2JoeGavlnbYaXdLv/tnOiEX3f4+a3qa8MDiwligOcoLWMNJMBR9cZ6XJto
CTga7Gxdvpign7Fqfi4MQ3Q2zojNwdL47gt2gJ4GGdy0anab/fNDyNNIvxoWK01ahTbwqN+UBEqM
vEIZoBNc+oUSUcmBAbQx6bOalIaj13sQyI5s6St6oDvM2AnN+MRpk2AAPslQtJeyEosLKJM75N3S
J8V11+KVaast4pyS80RiJ5MJQvZER72tl3k6oFQj4Yj55dwn/jQYIXSJEUuDmeeYQfxFx5AMkgLs
QUmwS8GG8BVkLEeEknfZOzeRgIiywB42xXHTSUiIzOnYfny7cMRcNc6hiwvKrJoY6Sg7aqP1dBoE
wVCCXUtXwksG/GgbNp5ykfcJ+av7oZ512N1RkihJ++EACRO5LXOmSoTvAesZ6nT12JIe8Gj/ssgL
XsF6iQl1jug/i4rZ7TErqv3mhtkmN2PpB6fIEAaO5wczr26GekgW0qbZvdefcazChd0eLdLo4OVF
WMsXQ9IV/zrOWGuWp/ctsLpx088bRAlDgBTVTDTtBOIXj5jd4K6XT5qSXQnSetRzs+l/cIDpLDeD
HMxnJ6XiKNCzF8wX27003CaxZ4V2MkFT54VLEJ99jxO4obDj9QTL/4+X7rDQMzvSqRw10D9paBkd
c4i3Wmjb9sAT67Ig+MhIsFx91v9KRUtDl4SMKjFRhHq8+JoDOXLhWvmyAR9t6txk3wk+ShfQ15tK
OGgygHxpzVQhc08Smo48uvMMlREuadxI+VK+cR32TlNE1v7JYZWR869aesAzGhn8HxESmKpWqExs
i70EPy7GhTU9t4uU0wyUG8AA7IuFwce3pR1K5Yi5CSamTRwmRAh0QcbXVzgLFTI5+euvHd9ip1y4
SbJ7nuDH/N6PObWQNLhdNlwIPiMjeXW1t2qBlT+ap/3VGtsevEy4ivGCDJtfDdLqrDbmZmHTbUmE
UKptar1VGhUgdyVFSGMlXRmnsLKyDscqBJ6TVHgxBWaEe0cwRfIcAJJ1+2HgHE05uhCWAxOU3TRq
uU6Mst5yBUCLcs3VezWTa9rg19oK1ama1nP/D2dLEr8XLik3EQbcalRTtsJYUNxLjMOGUQ+4JRyR
mo7HWa3xDb1FgKPjD+Q0K/eUAC+HchNdIHfY0YwAafy8v0zwWfSgL8coMShs5hjFx2dfNtjrfJ5U
i6xguGafIJPXm6rCM/rgcBFGvef5SmYKjfBoKuZImuzc8sYSunGN7AK23MMAIoB7neoXQff6RYuI
qqtFlQn4WySvKwsyhTD/ptWFG61CBeL0CDq0164o1guAkGut7uAz3dU/7eZuB/IhrkPpIcDm/8aJ
DwvMPpC71g3J/ufPjyvQ5eETS0uG1AqRpQdb9DJQAahUwcttXItBabwdf1KYKGg7Uf5kmRG72s9E
aCThM+uyi4912+MuAP+5MgHHe9LUyNWPUlclmZsUhvFdTLhaowSk86ghEx8aKsVqr4XvYeMxxSem
/Rsg2nUk9W/wjlgnb3okNU9S0VIdmw1RqEITFsvUWoOzhdnKSFCGYeEH3iXJJqO5izGgPGvdCEwZ
WrNaxyPR/rfRAPoSfMw/btqjhchxCVtuqkPdYgSaxNaXy3KCEgRTyJ9yVMd6qit5ZaX5DHeKIkKX
3F5EPi3yb08pQxs74zvBPT9vi8aVoWOEYszzht9yjC4InNRWbXdsVa582Uk3vJuFSdF4p37CwgZN
38DoFvbyGSzON132m+PhTlp50Z9cwPyZbrrS3NqIZlqbzpAbSET1nWBVlgAEL5ucJBDb++ZveDBs
CDRw5JoqoZxKJxif65KeLAfbZEHsFMllDMslIWEOIANyEpKmYWT3IUxbN2R8osEZ+09aX/qQ+Vrq
wc8lE406D9Lt1csyW+DM/I0lmTYfz9ny0N5zxsGneBFSzwi2HwyqSRI23j1MCQrRL59appmd12Do
rhKQfDSUUYZng1JMldlkZri3vpqtIJ+lNhtVSAxC/DwcRZlxbfjKdbhrBI5CrIqRPJF6UMZ2it4k
24ZPdhP0Rl/PhAhvYvzyyadK0rHW8cZlTv+qporJ5AYBZF2vBIKDxWuqVI+Ub8XrXeprZUUxf55f
XBWfD/y7Bjwsn4DufhchBXrmCbj5MtAdvC2dVC6ZT+5xoxK9EwV0yVye+MDXcsLu4G7kRFTmDmJ/
r13yxX3fdYRVPcUsrv5/UBz0urNaArtn0QHLOPiDJrIka9OukqaKNq/dONJh/5/zz91757zfwzuG
nXf1t1QXG7VzBrRdb9vfPLtycbbkYRBC3WvtcEzDd5i6HlgPu0gahCCnxODrzEPtDyyFBxi9js2b
uQOL+Pki4+LOekphCcIAT9VCgk1G4CqKvP7FDcSUoOmJMmvuRZI2kIB/mhRSXnmVaxjUIgpj+vgm
KANIu3bwI2dkVkO/TOCkkuIGwDm7QCASocV694lV4BpBCChOH9yQS9th6miV21cOPBBNIeZgsdhV
OIfxvgQc/RvZ78nt+wXEtbVKKF4dY5keWn5hqpCFTImUiRdkESaPVRrfgTX3ys5FOiiclvte1r3H
iUXDR5tBJBWnenTWLFvp+OdNLKO7HP7y86Ch8U4YIBmY41Ef2rh9QnbUtB82b1qNmS0hWsLOKMtk
xMxcX4mZvNUadN6rTp9ajOzKzz7troG0jDWMjkIXg7hVNr4Ph1DBfPonNIkX9HdEb706CiCEkArF
0C8PsQDj6vQQoOYZSO8bSzIn08WaUGdPPjGy3dnAdRgeOp86NBpAhYBZktQXT7yRe8RP6jOnutRP
dElMYK2Vm938z1RvS4Sc38Us+QsA+1NFgNsg0kk1QkJGR5qyzyP+6H2meOQPgiQuEK2h0HLCwa0i
Fs1YgzkxKRFLGQ+pwBHKOGCioyTNPs4DKPIx3IhOx8KI/H16rRsuzQBUcJV8mWnEBmD1huawLIOl
k7WeEromxULLK4KTyCey0ZGYIp/Ac0aZSXf/a+zbQl9FMfZvLWVqrBAKXnIjGl7fzZTxyLYNeyLq
oY1TY+tSrOEaIcj3u227mlSsCMrfzIDIidhrAXzA3RKlU+JvaPvkb4npkfTcEmJvpdyS0dPB5UaH
LH5m+uOS9MF96JGDahBbUPVTuA5bdJq3+jgotUshF7THm7il/WuGAZlyWmN9suVlm2ValZrFbt/S
ePxqF+Aq0L165vEhc1bTtNc4asU7Nsx9aGdYZyYI0F3SPdXbIkGnUdHr4ORacFRm/nADPAHqbXfE
TSflvpw1d0s4EB7BiXgelyTbKCciJzULy0hIGggUsJcDKNxDuCWbfzxqSY6i/MLFb2w0VwlBm7bL
RJZ5UesZQcperTJc2fCGVcXxl42PGFWnfeC91+jS50Q21xrFfN4oAjexSqzVVKn1zbr4FQusvn3h
p6i01ye1qvQYcBO27NhPe8mvmzhnHKsfmVcv+PsMZw1Z1TqLta9jYhy5mQ8odcklaC2djlPcOjKs
DDvAQufskr567zzYlH1b7CmAk5DjostJXxO3E+kgfOn7cmU+zpLBD0ZgQIsbouVwC6ddgXnTVEN5
Wp4UNyO8WOYHm/sj+oS69GcrSiSLCNPCXeMyolM3TrpGslJ+wbs3uyUf8IYrA+v0sq5iwLCcRmxd
B9Sv2vzB0Q2l6xRcbEZzmFuL891CeBDIITGV1TEUYe/xwYng1lh6jt6OKAaA1jU6bSVTvPzj5i62
b6T0Ik2+xmHslB5OhXazXkHeyFeiMfZuYxIDdgSQc65gpDkfQSNfeMg9X4CW9KZlTHX0YpbH5U/Y
tXD5mB7aC1h1dpWYLbyI4M70xMT79ChdLUJ1Qezvd5i9X8Aha2U26j/lGddc99Q8GyzcTuSJuP25
sFPzJktVLxDXKcY01Q/5p7zijhN96yk87Rhrso153w1WfHeZOoxDWOmYdc7trd/HWb6srWozXrXx
niVIYD698DeRaHSTAs4ueh/bdrHPO8b+PIL0DuPmVX0l1ENusI/3ktY+nnoeA0MiL6uxcgRCCh1C
V1RerxS1ntuEvsDNy7L6wYRF/kMch0Zm0ljLwhaO23AsiP7wAyI3xyzJ8hSNnS/b+l7ZFKdXx5t2
pwdyLFhQQSF9g28uLUMmnWHudijupxmRyWGzxtfNf7JyiK3Mrhw9pgCgC98RNeGLxH4QNbxsXRrD
eV5NtuVFEh3fhi6EMy3z/bE+Od7+OGegz0LVDwWe2GskXcgK+vi6JOSfQXLzWPqOVCihG9PqQWOE
uthpNxqKWHrJxBmJgNbWV6q5BHD2aentrhZKCuLkJ2jsuqfU9MCNRKBb1ZMCACEqlu6/bgOgccw2
tzIaRQW58b++njUn+0s1JdK0Z6xe4xABKfbM3iBk1+kWndbTh3amhu2GgzeDgZrlY9mT0Y+zPRR5
aESHkyr2Sa85Thlrww1j9DBnTvY8JOsW07q8dXN2QGpJxe8e1z8Px9IvLMXUjlR96UH3CHLGhbib
vHqTE8HoID6Al1yE56LOIc05vHl9LmRPS0iDcdkEwsAkIbdPy4/+ktbvDoCnq63IXa7wFBNsGC/O
pAVu7sHTpSbwecZQ19y2DF3qq6N40tJdO2UdBJ/FdQmgxc2+2NhiedZjOS2bHyVl9gTWInDo+Mpj
DY+/RT7g02MILj7insMUBkydtPLz+cFHqtg6lX0o4OYpGFbjCadLtWqDbOfS+rz/ErHklFjSoHDm
duk01+YrwWlxthPUFH+p0xJyaRptNF1xuUPi3n0lqVI+qMxIio6sfx4bWychASna2wwUrBGp9YV5
TrvkfpwzpXH8Ta8LeSiDeeuRAy/8crQRNxz3CosoN6GHnAWd8SRzOHXTNGypkzJaPUxk16ThZL6v
DoQgGEitnu/dWRf0oNNGB/iNF43tSred7maOOYZeaEPm+xIHmMQfriwDaXZ88m8le43cd5ahHtba
rxfk/Wq0Ns10sxRr3ZhUgCQF9E8gZHG3ZIdCsLp+jH51eOzu4ot4iG4aU4JRHncsMsY0RsYCExP1
0ksn/a/wisZE+usV/unSOSe0fLOBcKjl8SyzTzg6u2QqPOkOBk0AuE34mNWfn86+UuAI2LXqy96N
Jt6YQ5QT9WhKQ678kkPncqVfEmm/W4/9GKZwKZ0IyldK8Xc8uyXY5fQJxDp8fD0uN/r1/VTVfz+y
rWR4L5kgNTAFizrb7h6KEnaczRENhRi9ued9D/3PvBPtzpIE/zsflbPvMwzXlbUBnGZrR5AezvMu
G+AiHEC+yELfohlhdxpFwrcabC6pv4IWhy3jS2qMmcejVALDGlKWZaYyMtplZd/ixX7oDVqDNtzz
h/mpfSLl8k2gIZoY5vmhVXwvPoJUwr3Tps5AqVEgXcWI0HQ49MWOlbAkaGJ5Sb0Xg/JjTsb8V9gV
pipB/15xr7q34rfpYA7//0DxK1Mlba1MIzWPe3ECRnuo0GrgoApEfkJk7p1HE1Tq20Tn5372+XPx
f7pxTYgWmTAT6DPh4dOGtE9kX4elsPmXMhXAbdS2KnvDMa1lyd9I71fiOKad4AnoHqwjCRptaw0h
vuaJsP8VMOZ9UlmYgxxPS4NrR1lWc/i3XX1oHzQv6htD4JiR4jtyGv0hGLSREqTgBWACPlBp2a/m
Rp0gQGoc9h9neRhdkRAGsW5QuCXnXpSOMnxd+RAAhlPGifhdSpnDRRn+uLjKtv8BKWfoolwZiIJo
nD81IAQaVSbEpEBLrsJj9I9jla19npQn3plsvBKdjdea5eVefhsq59P7zQNkbmS1zam+Gha2nEVK
Oy9Ib9gWkzt/HZNw4GPMzEyt4R6IYWL25cdgHYaWi9D3c2c+BpCl0J2Kc5ZKw+jnqsQ6Hoq/B5tg
RBvdOgUbLLmin0x/gXxklpFSHnM7R1cgyOgwp+gk8BuYlk6EaUsqNfHar2Xug/pNqs8TFzObUPPp
bpithgyddGVTFdKVeJgjIBDtsyD6hwuMIjd9pstCukKXDspkpwBH8lNxlMB5DLytgrEWuvxtdYjr
kav2VIHffXr0qsKwh4JJe7hOk5/GTWhoINZU367gu+DSREzBEEXS6aLugGJrurENlCiRNfDh94Uy
lHem/aBY+Rcc0JiG+lhYwqeisczV2g0BjjqA9gKnYtpzrKUlnUr6wxJYA+2ovvz32aE97cndSStD
Fekr+ZyL9CTVtFgaxJnhPG+8S2nC+1oumBVpByWI2Rtarcn0Ubj5niFt+KqCPHVsmEHT0gZzCoGQ
5q9fFtMirItZf98Qx8c6VhaPm2RJD8Tra6au+is4Iv2iziKiygXyqoMilLllWFMENHlsw8eSX9BH
KYFeuBUBhb7vDCQv610wIPKVJq4ZHY91OMCEHU9W6Q7/v0Ee7KwBv+G/oHIio4h2mmQivadCk35x
Xq83KrOLGEoBY9cZWSL66rv/voVagt9IW1JvIBv7WFQFl7HFtwtwx6Ta/yWqms04Z8/e+QBhvXoa
0NqBvVgeXV9W19yRZY1q2SkTlxDKU5fGnJar2Qn+5wc5+hKc69Hs5LLd0poP3hlwqUueOq578mf/
+d8Bs2DKZczVjnJ9hrgG0PPJVkBLp/F3cpemJJKDIY7LTyDhs1M4mIZupdbNNSEpcvcXJ3Kj0hFB
yDx/+njujzekLvLyaiX2k81++A953D6CTVMaWvpku9u4BupVThissC+S8AkZdlKr9vLf/WLu8y1A
xQo1r6W10+ZptSC5McjVk2hMoeBLUKzFItibrLA6K5sw29lfKlUgJ7SuHSZa71aMieSTdrsPcPvP
FBPBPRkZ3GWNpHGb+E2IiNg5K+KK1Xu+xVYhqMZth6wFD+s9HOZJ1mkrOicYxtF1JeYXhGp39I4a
O1hh2B0IV36ybZZ/CIvLiTHcWkODWUWYuExSETevHrOnI6V8qlGa/o084tM2hTNmSKY48mNzbzuw
iiob9YBVEtTTuUERPS1/YsTpEr4B5RUtd3aa6bQNAcuvr0HyHfbkAiKVPxSOvhJkO8JMMg+a+WTY
3cWjs0oxPmGxox9Mo+Jb+HXtF50NlRCGrKggCAmInRkNizJOIwlClPD1QSOlABQUKKxPLuQtXQgn
cxnFluOxdtCCmmVc3gV+j2yJCytGRQLp86z4obPoNA7G/RSfncuHgzBuAto8xF3wBNfQTOqjlr9j
2FpumfaL1jxEhpxqpMuXiadDO1xNYz9VBuCwz3dMUMA7+potSAAIsXOA2Xl3z9F1lDEljWPFsbIR
uhv0Y1faUw7vDaanz99Lh/F3XWqfK9Lyv7fziJeCc9WUPM/8IpOoUBtAmHrYFWcEXsRrsPi93avC
azSTw2puX0a7/D4UO0jKKtEgUbV1lcGLwIyWsyb9knYLa3xeRZ50J4CD7Y1p78cU5xvC8ZeS5q/k
uzi/DISrA80vw2zH/pT/7Ez3OqJfJkjeqkhBx/uOR/9SWODyMR3/fzhAp3QcgC6xbCYuKhNVVYpW
UXVNyJcyRyg9n/3p7C/2EL9DCMzekp0jcmO1QOvOuTMiOVqd9a+gUY4tF4WOmUBxj8eng9TizQ9h
k0nTDBxpAoWAT5A/ZKhSHRLPoQ/SS0PZbRsiXphj/THhNUOblp+z/0Spbkr7abM+R/JlBe0tw0X5
KIf/LZS3GmvTy80mLvmgdqJOZc1cCTWkRh7qlt0Z+IJ9upqMB87kp2POFbgaBIAN/dPZ+IYGE1xU
Yyazyz48be2HQelnemI1dQlZFfoZe+xP1QT5t4DwcO1azRNAwyVSwFq1VaGsj0nJXY518jqHkHsJ
0aFnsVEozLStomHMvOjOLEkLQr8odDALrTGX+5iS4EMbgUmf2KN337NC0s/5ML6g6oUgn/Rk4gr3
yYwh5RZ/Jxq8DCcETJhrz8sk8YOMnzIcLY0rK1PL6SVjgCBC/jdnOujbyw1XoWKr8ilaABfgGzi0
4Rt791VtgqA2J+2wEE14ZIIJSVKraAbAU9h1h6KlsLyG8qJdEi1ev5CHAAnOJdNs2M1EU8DstW5X
AQjTjncgroojAUMHZzfwWu9Q15dhamZ33897jEUpqF0X4zWNsp4yEUNYKKl/aovK/DVnCAQLORB5
JMG5MtKbATv5GZpxVO7LDz/ymFvia8PgV6vZpVXxiTpX4IkaDyW1BZxUMbSfn4IerEpvr6a+VG99
VMBfHEQRLONqnBETBHJQnDmCbbMTMq1zu928VjDi3TboYb257WU7pYP1+mf8Mj/3vHkIRdG4k6v8
Q6snbJHsqWyDeCHj2BXLvjEPRl0FfwJsmcvYDiZvDCe7kqditk6djo89gANjGJZzywR6Ku05UPuS
vyB2vp8I+tkeQEmQLvn0vrQaP/A6edLWCNAHhq3li8oNlBRZighhGLWMz0Yl4yPxxsUPNlsBO1Ri
gbDpm7RogvsQ1103i/2cIaAUmW+RxhWNoXqt4wdG/Bc6ONmLrCq8yLlbGHhU0/VsExAVLBrZORB7
pOrprxtyjBV1Y7nw8unSICFkhkSa+ajdx7W/gS6+0izo+M0KFBtbAID5jj/e/rHXlk50Qq1JW2yr
LlgcYxmrGW1FwNmVqCX8tMTOAgws8MBNkygv7FaxWNeuMrsn55/SJ9TtuMjW8RbsZ78qfrDmG5+6
HvFOCT3f0ayKttA1/iStbOYcB8TnQ9p5TP2pppYyN/mGAv66r9c9LQfg7J0ZqhFYD/wDivTyhShb
CMmC2Q1ZagZMKQXLt2OKp0D37oSTSYPbMCgbvNDkOLIIZf45+tW2dccSV0O0wrJ94HqV61+TewrE
f4+uN7JzqZw3T8kJDNyqIUHkBz6y+N4hhU6NwXBcAN6cTh378l2+9c+auKWVoFsQt68ZXJMr3mj8
xgTnH4Fg2+ov6RJZij36EcrF6jQsBE/qBzmTy7JwqxpB+gRwx+kzWS2T/LEbY4Mz4KWiaSSJ+hwA
b4djbgiQ9aJadedNuvp57pIRthjP29+1+5PDf/XeWx3iBk396YKCQOk4CMX3XtCyBUpTJNgl7qt7
irvxciPoRR1OTs4pIVcGAPB7ehR8ZSj9FTf47h3co+oMpqWONY/VZUlSABchuUOfyxZW/W0iEDzL
XAxCJSNLJn3I5jnzKL6mUZME7IioDChYMoOfWER3nGC2XuOQJIRRp4LudtHBL/foQ26yfDE0Q9z9
R9zKw1U6YJ6M9cD/XwXRIp0wbmTDGsTjKcbUBUJ3f1WawT5qd4Oduu7HLcyimwThKOagVi3vnwLc
X96JlkWwItdVGBIklq9zC+6t+fFwI46S4t3Xm7H6mbrych5zpycDTKdJL8274ikWaA4x/OCh1joG
txLjYmxF8eyECgWX+8r/I+PwvV7g194FciQNggn2jEZqZlP41E7PbwEA4vCygl1ckJuqo5eZaEMx
sBhP8zZrKW06lJSnnDDvOocX42XtU1Y/ZiCml+5xDAmjQr2irQbMjKg98NjvIPttLWLaBwpaHCeR
Fsqm8hTGK4JfGzrr9Ku4v3uKCoCUT1JBusiag5G587EPUXx1hLZUW4Vihv5LkrH2Iso0UgUu00t9
YDTgcsTpj9Jp+mj8Gtp1VLyHKaiddXI4sIOVGo54iY+A4gup3SWca6Nuzd4E7Ajk3gVtqb68YoDk
9Wrbvbg6pBOpGwiZgtcsW3YXbkh6Y5l50dCxvuXcMZKGH/3uFuYMC55t7k31+/AGjJez+s2jVGQM
jPxPyPB4e4o0w/j7/3RZFxSoDaRAEYuK0GBGBHGUw9JhVS4JxWbRfp0wfA8yBx4FoKjpKbCJkPpA
Y0GWpxYLLH5fc21MCCU+ueuruR5tIdldcDx0jsE0oR8Oh9fg44i/jch/tzqkSajUfLPjX4yd8qr0
JkeHQe+V6gwdj5GfKRQ6Uqh33CPWCTAf4s8+mnc8uJvX1yUeXkzVtLCTpna/rZCJ4/8vdurGcGs7
qRIfQFTfAWju0HpWvIhMh3mEKH4bVcpJurLGKIYGunE61Ns2NVITCJYgLuYy9X4LksZ2Igjhp5wd
i/LdhW3zn1E5ANm/wbaJU3mUE1SazTJh/nXBWQIr14/hS99rBi+Brze1v7frtLOdrrzAMm+Ou4Ml
yxyL56xZUt49XJKlWsGCdzhELvwPVB2Mct9aIKi7RgLgTSvaRmUiavocBCqbvXutI19lYYNfYUM3
dH3En490hAlkOQ2KM4D5wrAg9p9Ckwf1zbhiAlE0mvlpc3XCiLOoGlU6PbCgx5stc295u4qfqmo6
AfmXnWt56dg9adf+Ok2x2zpnwbZ2nCNW1/K7ZxyJdUvVU1tbs9GniozFNIVb9EaAz37h08Q+9lnO
2zek3wcAbwCifcR//YdsTcKI30BUTgV6VMWu9QBYfWFAE4O5iKWwQsjs8Yq19gyf3Ah35WD5KHog
lxBIZmd2lwXKsafMRa/VPujB90QXahjlgZJZtmLzunn5e5fqExCOQtr1U22twvA2qQg4aMofVy9Q
vsdVbBz9zU7V3tn0Nc3zXlPHeb+rWLl8HFwKvfnUuFwWp87diT6930WhYqRD3KQxOjDM9x+D4hFG
BfodezPbGtjY9DRdMtrTCYZOPhXvdLSUOh1a/TatRuUPhLVPEFyMFmT/OmYwP30FZxoBSs28eSPb
5YtHAPAxT/7c9unCQKZ8qtGvC9uWYR7XFBXx8GR79bZXhbTFWjOXLxOqDZtgH1g7WbN5yUBwSeTR
OZKpOmuWIhwBzFwcrue/98Lgo9pllfVIkH6EKsRABNP2kl/uvoa/Ta+gKo7bBgGUzDh68U+jxnmY
6xtjfMO/F13TxnPy5HRAuNuMNARU2xgZaGCObmXS5lOe0MfYzxEHAazR9ZnNtExFhpOhfMEpVnw5
cvqtT2fI9jkuZFg4u7otJ75lZhxclCUxHfzTOYFT7gsJMPiFiso1OS1j+YDpcrWe9HUZgW1nXH4D
AIqCCTAqwgcr2IUF7qAbjW+GJjriYz5nxzFVh117qixuP84v0bs4zaX3XWutyZgVwh5Z8WI6ZnjD
DtErOCOmZUGMm8t0N3HjHAQopDKWiO8aec1YzaklieF6lZ6JfOcTvTai91JJISpj5pVEr9xyI/6d
GXYZESez7j3yr2bSGY6iPup5hTjlX+YnEkHQOxT77LROu2fZ92jU5Trvfw+GE/t31hGfoZe2X103
yRGzEQdVS+lQbJhUi9noAc5FmCF3Qfz1mdqgjzGBUuQvw17aHiGPAZqG0EckwhHUw6/UxuXYT9B8
e50MALrjNhV6rfpJrZ9TIYQx4y/YS/BwbNDrB6j9VZiFArO+A64fnnjQM9y3OJtJekuxZshCdRWE
pJgp3UituuqXbTnBUoypFPP3r6k++mVIUS0udYntmq6819ciZbRrx6bIm3A7sBqgdPjPYq5Cxh6/
U7xwEROcHdCq+Fklr4O8PvP1V6ivRHRki3U6bTW+WCVXSM/VeERrqlbPJ02j54p5f9XOt0bx2VeN
6FgVFB0vwB2CTHzEHu0uU7YXszaybzG2ecMchw+0E87nK4GS00eKVC+4L2JJgGawvcdPEZv3KCvm
sPCxOsikYM3E3LMIQ3fosq0xsn2uOwVfDkpEzFwUR5YEQ1Kkysn5TP94leA4099dmgmJJ30JOaaf
uAdYdSIdIb1TjwF+Urzt833QlqEFHw6x/Y94i4nf82t/VEvLr7bR5SQUVK6jwivj1erUeST7eGzs
PAGZhKMGo0V7SCixGsm8ThzNc0bzYAVoxiB/FA9aAolR2Z7t+VQHxFwtIqpn+Ar2dmKozIEg0ARb
krSaDY8N+NqusVWQtFjsJlyrLI00vIrP1E19vNrk+1jod89n3Dpa8nE/zF2ifszRIFJSp7BSp5e6
X9mMH8cZMxGnII3ddTTWkWPMWT0u7zWtUziANVEjx6MqgH10X/UJorVZRymr+gyMesbfCO6XhbeW
ac1xctrNTivnuZ3JoHszAE/4uWQZLqiDkfClGYTSwoTpefP58npG/YgQS/dlWOP3IQuFvaFLOain
ThdVu5EhlQrL2kNMDmErC7POfaeGNO3ifJZuF1CGjsEzPJ8xyoJRi0ueLPvFSz9op+UPqxcIH+nH
w8c7EBb3gpEqApCFiZGkBjL19//DEKyUe/1k5L09pmboXdc0HRCgNxdQEr4U+kJWTKPr3GA11dsb
VJFGVIsVw0PrgIeZsUWJzhX5pwjJrpWnO8ho6jIBd7r12dUEkUCEOgiWIGhiAPfSxiIUqMlrpwTj
+ap/Zq4IQq46KNhH8NLWxYV1AWz4L6JvlHWTEID+SIUKNmApoyyN73yNI8J6LRoNqmmN28BDpsGR
Nqg8ncm8cML1B+XP/Q6StbYWwsKYCY29LfAmZkIJR4cvYU5JEOJJZ98Pj0W50m3pmaQOC2nI//0I
NkKQteSLksYMgS9AYRSCE65n95QU+3+j1JJLOHImo1NXVEzGvHWy+og8RCYmjnDFcuN9QE8UxMCa
mY1SLWnCV4iFAHTz3CWCsFu6ydJydqAVYtyq8pKJ8iydAAB2DXDp9lNhQuIPewyKDaEu+KhcMa7X
xlLWdSFNiefOznSEdTlVyROAjC5cnpzKH7Ihtv/i5+A8RE0WCOloAF0eKGRpszL3ncwJyVj3lnQE
Ct9+qL5Sir4WUjm4s3fuTccR+sSqEcrJKyk7+vf0FlGMC5+/X7rv+67hAh6/fpy/fnSZ24WiCEpa
ByHbwBm2wFbi4pG9HLC50NAl7CXsxkslEDGxvCdJnbSzc1g5Ks+BRdw/9sfbrjHcjaUcUrzoBNVF
E4gqV9F/qLGHkm4jOYs/NpiaYhytbuedlxJWQp8U6QGDwrFPbH72IJdR0u36wbgwRGU0TmEMxRZu
QVJxyagjUUYKSYsLleaxjMLeOS7PtUMNxK25hh3IECUtOqciLO6gRfB+y9ACDl9eBbFzsgrfKtOs
6hlwY5lgeR20RRWDs/FbeXNbrX9Ilu4eyYaby0N27ZblFe6boKQiULvlKR91gwul+IIA5CHvz8JZ
dbLjs2Ic49RrNIUVXgPsrxDV5aKggfCBTyv7go00aneDHYGZ1V5YS1/wHXeh7D5F82SuQB5uaSVZ
XSm3XRLnaehqnV3pPJw7MiVJEo39eadbqU8f2zQaLgSeQO0DBmTKLIUDK/sCMUCzk5MJ9Fl0tF2p
86vejjEzwem9/p7BGvlA+iKpmBvSDzMIp0Oi9e+zjMBc//DMNksUSkALC/05snBqVgDSk5/XCpQe
BgDJZV0++EhvS3D6JKzGtLcxzR/UORk9CVdgL27tm6qJXLf5ub6iBvyWbc+UNPz0WC3cMmMqsN7u
jUiVtg7n5QfxQRcvF9mNEMZTUfV4rflk12fNJkuU0fRzCJpUXd4Gk1/me36l44VrXvlKk7tvnGkE
GbGI7xuq/ySgzRErKJaHRFU66tUX2JY5SwIaTIswyvB9whi0V7fKgrtR0k0UuN8DBqB+Ayh8Xaqc
JQcMo2w9ozgl3oiriOhO6mayzB4CKoy0+2SvctOl1dx0DBoGBackrHb4Z/Y3SV4U1Ex/XXJ+UT8O
fp6iqy816NHHMoTeRc859qcTkNXIHJS2kQtlUKopgafSmzTvnoRPbZ2/iaOxEQqB/N06/de6Ttdp
RL9aFCk7c8dm2rGkwIcOqt0y7VVcX5382IamQU4bVe1l1KA7XEDSrL6K0Ip8TN0rg5ylk/vZuITK
y67d52VOXKZJAcD+3AsIFpLngoTnX/t7bWddSEiIn2HlIb8N2t13EInAKYRZy4Crw30Y7JGUF/up
MvqxaLfYOO3wIqHeN9D55UV1Boj46s/+zDoZHh2ypuZeytPxNzCvVDMJVDF1NnXqBei32jCvu6eC
sjh8MZLyPTRHogCNMrAuw2CnTIvpWa0EkCFlQCSqmXtuv191KCVmhfB+cG0nQsZbeymflb7/4KE9
0DG/CRHbQawV7SAjRc9cqU9pXTxcGs+iBnOjQfBOyyrAKbGan1kFXWRJgORrFTPolISfx4Z82QFm
t4K09SqNy3Q+ZrHOABedz9dHld3GN5TnEbSl8uPLjpF/okDwvmlTgjuA+RyWgCpj/SeQ55F25RIb
HUstbzjHQHEnWJMo3pquzosNoOEl43Kg2AgF94uz+XTJL1kISBIhdUDjEr/2SXmjNE5ME6ndHPZp
xDiSG4wWQ/M8OD0B+ji8ySLF+jEUIc5ZavUAHK6SNHQzJnwU8+TtLuw+mGCAqq7SBkuDcVYG4ge3
ZivDUiJBPPkErzaawnHF48AxQVGKFUIAraMkUrULhO9dOlFxKQaMCJkz9PgEA6DH4H5PujV3fdIu
ErrqMAa1dqCDgQN5tkCGOXgYtv4EQIBQ/XiV71KaMXTItTYhAJ4jvP1kkeZXlqeyF6J78sDUu4z6
HOFA8xRVw/O/u4dhAaZBmaWzCjYZRKncOYWvnYPmKU/E/IjUqkMs6DO42/g1DhbUJSIrRq1xlX7z
0U5e/1lhgB6iQVFdivIa7ufVRXOi9O7OO2u3OaauTVGsq1V+U+bKwfnEu73gyzO+56u8u1fwYMKG
dGKvNfXWUJCnXoLT6lBHKZdup/+VyNAigHzMeHGu+ODWENYJRPqMwW1+PsEBbznJN3uDDGnpc/p5
bueewvuWSLsaxEb8ZXQU41ssm5BNiOeVinTjMO2rQDs1TR+PSBdS6bP1boEJaZd1IyNyZXwf6EJl
GUT1dDRl12gl396m50GQii7tei0bGOvc9orvQ0an0AJkq4aFV0bKYb6jsA/cebZDdUaLD2OqW8kw
XzPLNV2tRwGDEVoik6b7Z9vfqWMtJHmCCRbWAAKoyiUY1GKq2qcn+EURXzJLz/yb9jfgfEWCq0WE
vRHgIl/rLUp76cgrZxurI5kSdzDNmaHaPtlk99iQB588vdxgcRD/fTWfE7wzoeriUQrHRM/aD5o+
4huai0GY/2vEG5gIoqZUsdIzSLHFlxYvTnv2TY96EIgoJ7vDyGPIlNIq87VT3+BU63wogIs/Dbev
G/1hFflGvtE2DfdMHXmC0PFOF51qZfjxmeljMuBaU1EOIGcOSvKVmgeBIYMDimCqvmbazoIgA2v6
wK0lYKfu1m+VYNJbO2H4Bo1JdvqcYzR0k2oBG1KpvHqBY9Z3Yf1h/uwT84pHU7Z2y3YkRmKTlc/n
gjgEhUsE01WVoYe/Z5R8r1kwHHpZbDR/mDk0vN8kfgpzSlyLULHyT2PiIimjKsbovkRpTfvFvGId
VSYVEhkURp6GqliPvRAozT880wZ/ZVjmmUVvdEEGWxtbnQgrbUKayKdXdduWY1TBZZv/hqDP6Y9H
0dHZdIu21qQqQXdZL7O8hj4oJHtjFVl4+pXFTzJlaO6jyxslVI8jyVqk29CUzsKHrnjgKucpa0Nw
cgYZw4PNkw2hIB1kYaQP9QDnS1/zDrdoBiTxg73LFjt+hTL4tuqqEv9VGr2iWRySmuunLGBjhUYA
HWR2KQiHmqk8DrR7DNIDwpxJcZFE2rqBRpPkKpUaDB1UDG45EO+dIORZNTY2tR+FhVmJZH+jAEkU
PHbugMRjrxrK2OOJEGskyfnMmQ/bAE6n+huQDociVnercf9rdzGvq6qZyvtAlk80gCYREOYmTr2t
KftdARbEPpt3CyneufxvMcQMyhohtAw7mmgEdqGVM0bm95vzdmDyZd5ZIymXXhbQItVGPTKOcw3m
9iU8SF+6iR1SUih+RKudZUtgIiC9A4Xfj6jjzbGGUZQP3mHUm5dqFc/0CacxmqgUMKkuVM4kAZCX
y5uK9zngC/xkzm+pmTMIJ840i212lwKLcJj3JVtZEqFETL24FKSZj7/rgeaD+4oVleC8J6i2N/5c
QYifkTorieUe3NlRLKtnAR75ASGipXurh5y4xnXK83dg7HBXNeoMOvUup5KtBjpwdS6MTH1K5Bxe
tAFBrKOb52WS4IBm84DehnU6NRJYqYjb2Q2+vkccRGOmFfMTQL6NxecJFSZMfj7Edl3nD7JlyJCe
0/sz/Cxt/HVSnbDSwy7fE838L0jr4zWzxIdFyXROdMw7qUzyAdCRjb/AiXmuon++ZOoZZjYs/rTe
wyo5lRvdb51FEoj/a8WZoODePM0WDSeVUZ5pKdKHDtFkIPyNxxyj4YaEHPmISnZMUq6E8rt/szMm
znZ9embjKg04IF9nNcvtmxcnuf3oCJ1KUy2zKXlh8bnmYdOubofCcJRy6M0nz02M7Kt2UjJS56aK
COkrqJeeQYjHS35JCkLPmgZ8EFka4SU9xH9sTaSWbdxKOahOd8bWUF0YsYgAEtlUNJ0aMXXyVqTL
H3y7pH0yBELspz5ALYeCLgulWZh87n8Vgz9D+cyG4Ji11M7N9ZPsleYEbNYjjLAflhAGDfe3d6Lo
XdRDHbnk+BHRd2D0HADx5oBtbPs5C1B17cHPFSDEe2hvLkA4eMFUCCKt5izjPa7IfNPViFr/9T/I
L6Zj8eJkyYRrrjV71UxScUoZW2MLT2Du/JghxoFeRS1hspSAtrwRjQ9k7RFydUeMWMCmBhhjNV0d
crGs29i8/1a83grPs+zWbfiAAdyQ2L9DbknF35IFP8IGjeZxpZUkM+JBUXlyW9mOrZ+ztHjwqT0Z
/15wfr0xUMi8j4DpDDE/TSAnJRty7M8VwihwKFThAK0c8MTzaPUAe9JRNpWjwtSklPD+SqT6v9Am
dCy5TzgczeJUpEOTUdJuDrbC2cXFd9Xk2pXdWP0K3KKvZnTvooVm63eZSeZBz5qAuaUL3Vbd8Teo
jpf29BtVEsy5AI7x7XzWg0DTkxr+Gga1s9QGHce6GnCw/Nac+d2AhSEFf54v/qlQ5W0CIS/MMyne
jWd09keZ3oh2yUk01ZrUKDDnnJZSMzCatFnckSjYqhaCHIa2VJJeUP+f1wHlfGMzsHNXbr5S0Nte
+yIPh0EKuc6rkASBvdXYeNApPZc8jlhfwlB7SPCpMDj82HwOF2qo1m2WWiGSJUDuxQ4oH0FEB+bk
8D8RgDlmPvtyPCJZBZ2d1hYovJ+1a99Xb2sH6/5yX1ikRMfz8Olq/1EAVS61e9AR//QlU9YJDDiV
fjRC9gDkkPhXJpFCMZh08hlr699rn0DhU0T7RfYDwbp0Ta7kmevnnVflFzvsTiFkP5rw/NhaYrg0
lIxhPPcyMiQKVuFsBG6rbmI13tcj7QwAyV9xGI5VZhbnB3Ra0mavKNiHB1eOUrop1jQGaDDEdhD7
BWMcsF5X77qet+2s8bWdBaHvJhweIdd2Z8cNFdYe1wu0bzxrK6S4Ok0i/e3athlwiSl7oKQp8/xE
bangWdDpIXTC4ZALaFmEiaiPaJNAtUg9IooN7xxDPdWYTuZuG2JqsdqB4zi/RnVYjCg3w4HIQ2/J
i7iLaKiSNrQI1/vyx7FFnlB/aLqOey9aSF875FD12U0vbvrbKoYGfmNAqj2eqAxyMpFGSfkpRJ0R
uwRw7M29cWMenuxNADx79KbLPSyXVAMeUuV5sPQ7koPmKdimN9uEU8MYw5KlHsdnRjLbi/vbLbYC
2PmLnw5WbdNN/3TwgERFRmTmr0Uhd5MhX1PKJ6VyFv0gk99ezKOQea6J5hdiPJj218MzRa4sRyw7
XPQL0dbVx3lqIH3uwt0C3gJFhHk8Ip2HrEgPKNv9fksNdVoYjl1yB0KNvknOeckTRIxs19PudRjL
s5e4jnWhPfmcNxkYlwMSKdQ7xiVZHQGIjHVD7xIB1r4uzF/IiKUAYjZF7tCDxvYqdhvrzF5T2vJi
JV8Aje6XeWPFEWrBBXzKK7BTBAc7e2kVmdOOKIJYbYWm18xfqX/6oTHybBJhLaPX4m/t7/qXdrr9
vgEULCisZ93Bcpf3s3DY3RUiZR9SpD2AJyr6lD5f+pJYBPFGJyBL7SBjo81UttJAXi4k+g09TTkb
q7tCNUyb3jgkHB/fVyRZPYhUu5WIymO0YYiZdKNR1+EOkcAYhUG3XNGha3RmgFnzc58Zs8Qo/gKS
g/g3/IifdO1Q2VqqakHwU+U+xG9p4CxmJ5ltbsr0twr1bhTDV7MCRw7cA6KtFzRZ+LUEb+5WaR32
PrE1UC6rudvQ+ryMF43WbJmFptHZoL6+9JTMpgyps97VriiYn/Dc5f1LfiYDU5s1FDsL0M8x2/2+
r4j3ItgYk8KnxNVtHvPwJ436IaapR4+/VucrphYo+2Z7ZfhUJn9+/LXpKsSC2R2IMlofbKz7Uite
yq3pyoj7srqKDwlE8Dv37TVJuYBIeSkBVtiDtAgypiIuVBUoKik4cJcba+4r81zkKxl96Lj3WZgB
GX9EopfLZCuC60mMPpEe8UFkBl6qJAy4eqLOUWNQbrQyOZSb9VX8OIVk3TM0BU0kFT2OQmIMyyxW
al8ZM12u9aRvNRjjpw4tp54ynpZdt+qBr6Y/TnD8WJ2iaf8rsmzuFjj+Jp6yB5uzS4HJwJcBNhCB
l4/o/Gx2HajmHO8luGvlIjw4c/Va23jkPoxMHT4t0Pa3fDcIBlQsSWqzTWOzYT0dPBFOlItD8+c8
JJnjjZOB0vt/F3YJZxbuYSmRY/JdOytbYUmh9/KQxxAHuIGUAmxjzp66XaOhOAwk//HlVI91x40O
rX0BKjuRFHXKqQnG8GpJFLZxnbSOOKLjLdIii8Re54uinLsDMckBKdPnhRj4mbuE7KFpLA+x6Qm8
GZqHVKpbIk1LEldMX28AMMFIg5uFBOixT8n/kkEqRdxXTNH+n1KRtcT6YFMBDnzAjVIBjilSJrvQ
g+JvXvb4ZeUC4lmGPJaXaZnou//CUKo0QXEzl7PxNEu9/SFWR7K73WevYZC8uTFUFmgaRP6tGxz0
hHLrPZUDpxYUt6mNWeRGKhtxHDqiZ8MVMKLz4PXWDh/SGMNZ7g4FtWT9rXA7UYWIcfVI2R58KlCI
b54LRJZwy98tD8jpOX0Yyb+ZyXUmJ8ntK/c1plxIA6Xfd41tpVmEnzbqhcI/b4ci+xCXzgkyyCgk
5IjGjqzZrKEqdubZcLFNu+7+/0ZVhbp9E118owy9JOsx1ZKK03M/hXn7JXD5liHpdWcJ5xc/m2mu
JHUBo0oSE2Ye0M0wyHfRnwbiHP/nZUjHqO3wcS5rW96ImyX0aTFgL5YkBrySmOD1l8jEgzgVoLsU
rX2ELac503u0W/Hy3QAnhd/83Zvf1TR+y4cAIq3q2B2txu8zGdzR1TjQrDWu4bzSTvtHzuN+gI7d
mXOA6Ggh2LiPol2HzftbJGYisgTiVAw9qnm03G8JgPixn524f/LzkzrpqHvYQL7dAm3AD8rjObLt
B8BzuBL17osymfGsqTXw2t0XvTB446+5GVkU7NqsNFkee0El36yd4C49vdZ1V+I2HDPNjX6gqbfL
ploDgX5U/pAGxlDit6wzDXHHIIulXucdiyalgPJhUWYBs0ATTq8JzeiFxo66fnJOdpHzMA31eISR
ahDans8WjK2gp4UHUgvlxU+LeO7oUwBvhCqxdnyWCnzgT1j9MLXGBh90E2AF97FFBlGlGVIgdCat
ePn2ueSFej3vv+lZv2f8fRoECrw1nrr4i6KeoKQSiPXJp1WQRcBUOy7T8VeaUVlmWOVR0zIAvVXx
y3DzM3Rjtk75PUGfWRqB/Hc1N10igLPvSHGVenfEl/N8qxo8RmRFqxJUNt7gVKuVImQjCSR7tkgD
EIaAmU52dlkBz6VkgqT/rAJ7VQTLX4YrSZ/Gm83zqWTv33s0Qz+z7IMajd8+wr5JOLqsBzRftdlC
iBjMXEysJNIh0W05IEal2YbQXpMcseSjcAZi2Lc56bvyjGP0J2Z3vlTOyGl7zWyln2tLeoexswoT
7/FWIqE3eNstZXlJkp9/9GBtKWvDDN9rFC9HiKqJYyFKQezHtwD+3xqgCLbfCfSUZ11dVADbxT+e
iJoPAlGPoWZZhecSUyympQVWEcDhJSwFpEl60J2APnHIxkxpKZaIjLWS1VuNxNZOrN++IiZtmYKd
PoKXMyZaP3cgqXYjABzhHIxRWpaVlCSFCnCgv/LvmbfFbkdwcupF8ELsevcpuHaIZytfnt66Pcg+
zMCQzCHFvkYy4WVUTL6Wdy14nWHLY3ela1qlGOLPccNYDKiiygVV4doE4mRIq5EilaCRK5VAx7th
3rV+tQ9Z47vjbMokgBgZu63AAOu1Ysm2AHXmatIIbc6q+silczNl3WOAuUGc+lvCTefuqCvy89ge
Z54USWqRZkRiqNtLq2ZL2w951tes8jsGfwER4nEAQsp5vgKID1sLqtaG9pRFN/5X3OS4KMhRmn6e
A8gkg7KYJVAOzvQyRE4l7AvA7UjbXLIOZW5Mh4LZ622/DTYOT03fMdoYWoFQaIkK4pRjbNlku3+k
OGUc2fYT4ZjM999CXk8NZqOpKRZgfsywQR9FwkLFaOGkzBuM9PZf1a01CCvlJGUQunRssIA2YR0a
P7byrGZJlOU+GanDsJvNW4r0jBRAVvDs2tTsIFZaYZL6EOQErhdrhsFXuDpSeAXDdovunVNKL5rh
sr8E8/BpiGKDBqFT37mdYnjKUAcERjPzDI1wVkkjI37Ye94lbhEEGQxuAsImFz9Ft5ubY7LYZCjs
0DDO27fvURYWwtWDu+dnm8upkAijRi9kh7mpliK5lyttQ7GZGrdhZD8UprJ7yucoZw5uekFNiwJy
m2CU/snFLJC/YeksuZ2qgiuhvIr5QOkUs0cqPAlf6NgsqxppHJOzi+vp7PqsEmNt7kbD9cMX4HYu
lhxJEdJPQvj8OKKdK8xBI/0AmAOXzw097OUX766oTNgQHgEbHijMpLISKSpnr+YBzepwF0FUZuLm
uDoe/ne8poHddkeVAybe1aByWeCpoAIVRQHUYUBZEcnFfeB/ubZC8nqm0eb2J63sTpRGgw8QOfuX
u/iPl7DIUQAuDsCwVOBxSpieeUbYbUgwUV9oAqPa7H5hnltjLi7mB0ZmIjZLeJpMMEy4wQcyw2Pk
m7MeYAmNyHrxtIxSmBEKtpRbcMRiRA7OY1bsrRF9+CRlyHcaYLc1mgPJJ5lX8e33qziLumKLNKiX
fk62ztuFlvmewyz8LJCjPAHyFHaxi4pJDBd5wO9cVUeonNSL5N2qX3oMyMmEyoH1em5HMYgPhgv/
9xPpBy03VwmRDoZVKTvFOgXl7xwnKKDCi6jI560h2Na5ZqVoNADtH1cJC3IxpaaPNm+2VzVUjd8O
28FMIBwL8SIRTrmUzCXreVioDEISJf+/WaS/y111X0JGC0WZYmZ8b7Ai8gJ1I3O51Os3fX3UuNBO
FJVYELl/Zr0wGw37U12vwy2Mgqrzn9ryOV3zYvaegb+Zuo58TtZpTDXPReFpBJiwNYBXOHVjJdO3
R+Ksyz5v7eQl9gTvkp2iJBTfn5u9OMOmkFsjNTyGJad7OKdUQtkAu4+UYQdM4+fyKoFnaFFh4cuP
ds5RPI4EPtPAgLFwG/fIEYVqafzXxVyY3KuNE5g4vO7xWxw66ajwueJtXG9zes8kbYU1Z2AYGpSJ
wX1qK3VsssvbsHqOHnCp369zw8mZddZ7Mp8Sv6m8XH3CFarSkZBJzArP4isarcljqbsudYRIxmFx
Hr96pgv3bnmgYOFaXsgT12ExW16zlzq8ic0sNjYeyo4RIxL3Z3HZUzlnJxeAi8XJBxIMG2lf4b/x
1SGnoUVUjpOoTOOEV/PCSUFpmAdtu7yw4hWcHWeaGrz++8z/JiGYsurNEi6vcMXhy9PEfvb3qO9a
zyRTaokkOPlTl0+HXTYsvY3ANYLf3c7BoxJZFjHKaQri8NDmbkEU1D76UdqVXxcCxqnsbIERwL24
t8wvvDm83m5KuyzUIz7AveW/QdgDECwxe/a2CGlUa8EcHr4XOiO+iUYGeXEOGYkYoN/mQGWihmpS
xGUli+JV5PXF1XrDT6ub6Y588B3z3juLQC9STVRomguV1yYJU8AVzz1Q6RZay2gVALFX/F6CeFrY
6RoreSdIkjcFMmkY7IaFhMTmBk7r6U1u/xnjGBufq+sAVSghfpqpmGTO37qR5s8U+yZmj+BPjNEC
S+0CAmvEgVPsiqnJIiiI96ukR2j0pvziJEmZj159dTbilSphM40KkgQAB42gs2skUEy4xDJ+Z6/T
IV99vUoVhr1w/lquMysCwQN33X7pQSckknNS3L9sF5lB0wf3UFIjZ/OcNaw+zZR6//cfKYwKQeNk
UT7eOfgYPM0qwIuNLm9QdKvMI58KFO6x+dF14EEwI1rXhNET/SODsjDcaokDn80inssuojE3HEZY
8OVvfWvZ2yPlZHB7kSndQWlqqqrh40IN8H657Qgz5sAnhf5GB3JTjYr3P+Ywysn8OpOZ2MN9yvpr
7VX4/huv43i6Rigv6pWqX1X2Z5XeKS1VVU4DtC6OsvmtDAEvjkc0IkamUTuOBTLX0hceBHQ2smKH
bD6dz13KxwiIge45Gog2JFtWI9KuErhD47uX53t+mJrbDu1+HMrj4MvWp0w6OAA6OQQrYrvXD6P+
sEN5h+eKWVvS9apjDpJRrMQMzobhjJeAWPYfNjfHmOhcJ4XP0X5ahUYvzMEvkXlPaF/FoLDfBOBM
LQE8pzv3teEpLRR/rp6m/h0oBZggvwXKrkBplvrGqqm1+jJy1dTDr87fdgsFy7AVl9UPCw7tRRXv
z0GWIQ3r2yzUM1owv5PGwGJe04a6LDSoLWZCs9Ih9O6PKOICr8yufQ+UaL6ZKGG7u412cCMWRMiP
ehG6IIWr7bSSOgPVEY3DsKc7VDAxTw98kFvx4Hh96QD6NZVWc4MY+GY3nlcfcw5vnOw4fMe0Q6hy
7/Lj4QXpuK7W6EVXVx0HFpAG4mKz5LI9hhBTipYIZ7dP3C2RvA7twehK1lWlRVdmJ3CeZDD/9wwG
A8iyfRqqcpt0EoT0obiGXDowz81cKNi5lxTwboecU409KS+BY5NP9GFcMaR2Pa2jpR+5y/QU/g6Q
tBY94mK+TmSsqaHIHCp5X06R1vJdK/a92+2ZbpOsQJ9AUzNHMS6w9gVUZsSqo9NUhlT2T+WfXU8m
Z4UzjIif4ahFiulX+pWbDtlNDRlMeeoaz1aTsujmI2WwpR/lLL4qlp/qXpwv+s387pcp0YXXRVU6
e1GmmVFxWmXvGf3CBbyglU9t3DWgcfnptnL25tX98UaH832nmj47x8BD17KypuZ1+u0nCHE35ZW+
/ejFIMmXX23/+64qFYv+tYDaIk950hA7Xk1GbX2eM8LH/AvulM6xKZ3+JH103QHwSbfM6/2c3QiT
BsCopuqEaH0kUZNdKJK6Ip+zUlpSi9uR/mguhUqHFO+3nuqjg+jfnqw5Nssr1IT3GzHNjmC4ub6r
MKFm+wkfPoNf+ffTwlfXoHMcMiBLHpRxkEsv4VXG0bMEmQM0LD9wtYq9JxNCgU7AMcza7YLEttgx
UWB7dEljbxiYSvlocJNUTs1DW7Y3mDLwOMpMKqwarMEOQ4dY2UBValGEG/rshh4SqeA9qpudNYF5
6lqGMsPR4vjPGJEJJL+46sOrU3O1LJm1+0+RKB2Syg4V7Bp1WYg8kE8UEEbpdV+odKD272ckk0MI
cIoMA+NBAdq6ehi6lV12mPoJYA6P6taiWd6/dLEmAkQ1otDwXYdlFQP7MWoG/HSI/S76Zq+Aky37
m0GFP/WymSwf9SfELprbagjuR5haZbdjzD5Yhd60sZwJIrHG/ibIHi/tA9tO1Gx1nQT63Li2I0XD
ZIe6UH7mhbqAWXqW8T/Jy+WkMXvzAd/hH/7tnNIrEbPmezsE6BCIT63IGDcIkJVhP89eQWYLl0x2
6dRhwY6bb2Ep/+NprcUkjDS6fskpzD1+FT1+QuEOCbsl5URyb9LjFy/VVS/QGrWZEqoSXBVXwfWT
w17wMhPb5JeI6BGyEVKCCYWXlvxIjsuvnwIaNzvnGI2kQNlpHqXEQsGxNm8YG9IavXjMJIliPrBE
OcP5jKLwovfp8j6/LQz53SQSv+/3MA5SFU/MqLQJOxtC6DsnJUNCab0IBuuGZp7ecvMiflrlKdbY
AibIwaybvmqf2UvmKdyOpnBdVG428bn34Got3rDsdu23eZ6gd9P689jl3sMbQe7T6ayFFqiC44Sk
oTJu7zaPRpIgitdNEG06zMHX2gp1bvnjWBne9n40Stz/NKZ/GEybO1TXvkke/r9jiWTboHXFl+8l
Mf7wNzTgT8GtEWm/EuFvOtgJ9g5V+ywif86UP2gga7vM0YseO0py0SOYdCtsLrCcU7LzIAyDe+DQ
Mdo1NRjf9m98eKOvWqXenAIsydv+eTRHpetdMFyI6ePciH+XQvAIsOn1bNNWv5y6Bwk/lJR74iSh
lXQZ6Z5N7zpqr7oQrUYC2uCkLabYGO0/tjNV3RQoUnqGVXBdkXNmcILfzHCFeedkVlj6NJxyjzep
WXmg8df57B1ZQKSq5Lrx55neIczWjJBjKNWtDUeNBg2J0N1QfmsfLpJRDH/eYdMsTsN1mgDfeCGK
Xrg8yotlw1/2Gmzei1jUby0a3IjRUOrOVmMRVJROjIbHM5JW/yCFUJpSLbJBB9TIJiXWatz7mefF
/jIlaAiDfTvjzD4Ebl/gQa9GfCWpVncsO0EzlyriIxrAWyZ6M9FPXTIynyxiHEYxJeH+89xAjP8U
7eYblCms+98ivudJEuVELpgdt9Cz0hxxELufXk28Q7ZLWUUW6c21hjDBTTs3g+u0vfllWlSC5sBB
lzgtkP/HsVYH144wt3k/Nl7iMuQIROSZmjiLtxHrnJV3jL6U8/On2UY7hfgtwlMVAc7d32zc68ZR
3wV8MAwUq8YWFxliHjlqq6zEoK4HlwOaIiLWU/pQGw/uJZfnFo+w3xPM0rDc32sXYK88/uokak2Q
Cot+YPCZj1wjXld4IlBySbVPv7ju1Z8twXDxUrCW3I66JwnJHI7wqmHQllBFcAKA9lFeN2G4Vw5j
CavHSEX71aN6+IVuwJ+9RWIaaVPzoHjZWYBs4RhPbfYCG9RJrJplmVQMuFCOGML/8PAk09kg1BRo
tFXwoY/YP6l6oIPu62lUC7SvkQT0Gyd2oAS2c8Z/wjovBAzZ3Nzg0bq3WRv38C//EkSuswQsN3gK
Pnea80T1rMC8UmEqZ3bZYuhN8wkWHxbyS1XZFT1scqcpHhcgmG/FHG6SLqlGxl0hVQQx5kbsGkAp
sA6CfY5L22QQRuNfiqD2oDTZdeki3n9PckNBFM/1YAh6IvhVGERGTPNOBz+n+cdosVRp9fs6cQsm
6SEpioRHTx28RX3r2BObxbHaVr5u1CyrG9Ky6nPC3EAw9xxfsJjGFDXOYp/YyZ4ztv/UhxFBoBZ4
Vrp5P2oeNWltJcKGoZNzdPlSOdT5Hrn87mIfUSVh0mitFVTnKEUSnuvYRjgWBobrpJ4xW0cFaayD
rtMy005PP+bInFKjAUESR/YodMq3LqM8o3hezeAYRQRZLiHIcXSIy7wMzMAbiY8ah4Uvc/1nVLkh
pFmbaWawj8UEFTUyylvXgpSoq3I/0cuxuZ0YYplUICtdBOAFUra+Yz6L+C8S9nDEKTlfoedoy4Mk
LR4UF+2Pa9kdh1o1KPtSrwlhYbC/FJZJLQRtm1m3HUkXjHkwZPQ2RAa8vv9BttxIWeAUq1dZQmUM
ElDVaxw1tNJAelhIFsN2ZcG29kMA5UDnWv3/s86VZRyDyVWrQ+6Wpq0k3XHMs/midlTjFUaeGXSB
JyCM30oiZqYn6SAgvtB68T8PAHfa/WXj83G5Y3EZjPaxqQNT68WZJOixwybniNP3qf2uYYlL8+RY
oFXbQugEYM0ifHXeVE3s1c2op+nRJHvLbnDHZo43I8Z08TrELRogjNulHbu8nxyJyP7Ums3XwqyP
whF2Ceq59NnxeGRmqE8waTebGM4j7T0M4cSsPu1RW8rP3+deDQyA1KbJJI1d6Aqkgrl03w5DBAoj
GlALVL4g0C5wFOdpG7j+MuIapWjiexosAGYH+Brs/eRmE8jOH2nYJwl1mR+/E5IT34m285cJZtLZ
xYu3ToqApjEdPKs99zyf1aI2YnsfOFDfOL0M8bvna4OqpwNUBVgmN7HVXqyVEV8punqYGzc2MHmK
VtoayhjXFLkFpt1PMzIS2Gj4bacoIxfM/ynYnRi/oYaG/nJr3LImvG4Vos9yffPRCjPVhMVYEGf8
ARIm3BZPMEu8hbVrUxfP3clXZSlrTQCPTLZCz9V48IX7/qUBKMc5tZ82D5BMp9BLKgN6gplnuFkZ
AzLeYNeGL5ualVjkMnpbB9Sy3Z1rP//xDd+2J+xLFSRWHNwPkcOmou4buhoZiZIrjGGN/X5k3pBc
uZ2EBHpHBRs0+BJI33BaNHc8ouKPn4N9mwGMC4VjUKK1MlvrLvNtfdzB/UjWyzFW5U9lMGcbvDlO
Db4bRbwjOHSuk8NJ1MtwdrHCd4nsvjdvWuzOLaappx0LHLUm2vPnBsJ6vdFKIo2czE7vpPPRg/Nt
VkWkIxUhRkA4Ji8yhFZUMvtTwp7+zv0WsK1qOUE686oP+lZG3kIdqJVVOccsqZ/bGzIaLMBIJHxu
38uOASM01MsqHeIZQzpBJlGNpaY1wqwFMW56DVd4e46S8RqMXRtMRQvEndGy2JngPVyyUn+U/pNt
ko9zOg2S93Aj0hMtlCGyoNIExUlKVkXXKP91k5BxOXvwZBAW2cMkyetuxJiUh16rTusjmb6T4zUK
BYgT6/UpLusZdQLMq1oZDJqbztAxsdw97fkAZUPl9JJTQ8C5CXF2JIohNB7cL7p0fGNRPsp98wIy
JLHZ8V1sPR9wlOg0eKQXvd+m4AvgnVfkx0xNsOBUMKcrgn8A8p3l7RQ+Im5sw/dE8f8I04H3qYn5
aCrkqIVyjPP0zqMpFY+93pf4w24qrdXBXTV1UNwLFbrQKOu2aL0RK+MCVf/Ey2T31101ArEoFORE
xLaGfZUjTNmaUuVOrS/97xgPR5WPx/gTedmsYAQh6pbApWaKJEZDtAa3R84vSAk3CDvxr40fmGot
TdqSGzVgm7qZFHHhEc98TJ1N4w2WbQTpTDr/ICF3jT4AQHzEJ9Y5rBGMzJMvtTP9o4SavmEMM/u3
ixrwz7pq0QcFXCrSPlE48KtOEe3yioh3ZSRzgB6HF2Hb769EuItUHQ1IjDNX38yWLhwRoix5uf53
lwcR7eKwG0FlGF0yUEAC7HDOfoygDAAcSuf0ivMbNhmeTEn97pBYnBECI7ZuUric3E9xGEhGwYST
AnmfxeBFZTGihHgRw7f6ixsfWIB2LQXADZHj9rnxZ8qUBaxzgRYoPhnjFy7irDzWHyaTDx476tOq
OJqsw0/TmkWFRmwZ+xrQWGyUxmC6xGk+Axrms94Lnsi6r5BbBk898xFTY+P1las7/eyBMKbSWEBn
htuP2giabuPWbIeSKBak26lYkLTlj7KMtk9RoAZ2s/EbepClB4O1RrxU3Yr5DP4zDYzsU5MS/rlk
KMp8hg9V8297XDEaCXycvkOuE9qzzmE0gSjryOM2aEeJveuGdTjgTmoOoUPC1qcWSxkW7BMnW31j
nZOwvy2mKCx6zBei9sMdCwFPnf9oFgX7cMNCVAz7LN1Lvn+Kb5HT+vC+uCJvl2m6lOD+WYsfypej
bJprvNeZclQn1JQkj5v+rS88JNaCN6Tc0ZpPPXmDxM9FqK1k4S0zf+cE6y0n6IM4eSeGmGdFGEQ3
dvNv5sdUgpwmfmKsLDgmPp23SktLSGo1mQg428RPN4hTILhC/cLFEC17xMZ0hjqdeeREgaNH21iG
j8LiYqg68/hi5/biqTfT/BU5GZM0MQ+qzIcJKr6ZnpuU0Wn/6NKZ/lM3/sj+3klVVkzKXA2ziNGP
6Wj53epOJSxHjwFGiNMACy0ncfwnF5JOcFfa9ZmHpyf+n0zWuVgOWr5YfSdAWEifsPpFXQftfCFo
dInfzRlqG/Y79mQ6XrPZphPvs20B/A0WYqm40kY/66YudNbevCFFygllqqNup3oahcpuLkEeeFKE
UypwA2e0LKQBuB1YRk72Rrijz5QflFKGwV7GA52vHtcsUsDQSibYShKq6Ud6gDdGYUDq1pKqC0t7
9BGXKG4bpOVTPIl/BTn6FNX3uSFZ6ElFuPAyKVo7cyonZ5e/0L6WDf90qkPNFtUa2L7WoOX5Txi5
aIxDjDD4NKnydCtajRYJj7GvsyftHtNkUqqC7ZXKKci0cB0+h8KwItbmgZmdRWod3udRsaG3ajG5
CGzuCPVBLVOGifqHQlA/zHDpdwCSFUDQrTTYcmDZcNnddtwY0z/dr5sq34Lgexze5epl36UOZHni
fK+SejS6cRDLYYor6S//ZEaBb4rLBTAsF+WMefibPC2U9bkcBEvAImlpSYoiSQPzMbLQnx5Z3PX+
U9U0lMOiQ419TwBS5232hwFoao+Lecw1fzwCc1kdhAToLYcYyYeugnUiiuUcLpXiABdO34/F/nc+
B2tyle0HznbS2spCuOmQZY3g2d8f8WyogUzcj6msVxWD156OJUAyGwFuHgutJ4hoq/0jWy/ugNgG
nxFznHWZPgzP0X/ZBa+dzyDN3DlD1gMJKnRcSaxyi3ddXUm6DqIr4vjMYA3OfnYh52xTnxIk6wKB
mwr2lNb8DBIF4vgUQJ2OzdnCQXNu/7aB6iCn55L8tjztyMNzWc7SgW0ByN2R3tdJc2VbDxYIBnGN
a/MHjeppbFkFWgvg4DWbyz7y/oXH3I5UWVIa+vZ/bEeB1Z9tUzWH4r6tWRqR9oylzYWdcc9g7JzF
cwZKjOgwWSHFhReEphKYqC+H4GzJqe2eQt7Drq8RVN2MEd6XG6mr7sQYgn5RNN5CluJs7Gsm5vup
9S5+bltFL1kYA7BWrBcchybug8bnASXEiPKmbhtSX4JnJK1j/lL/Wx7vDPlLfroD0w6YpQu3glO4
SlJWsirdaykAJMQFqySNetqCr77Cq2NVaiG+N13fl/C+sWrdCQYeF6fznsNB/eqW6W3SAw9FvOeT
el8RWDPUgHAtnUSHhSrvrHfT9XzArLuZJAvW66VHx056qdg0crbf3lBrSGYSVJjTVHNd6M3k9A7+
tGGa32d7vnLhUG5qg2iSeeYVwLilv898hCZVt4pisiaMdxEF1nF/pYr1g+zp+uxvvwy5BYrx8Bnu
WizttM99uBoX4v5UrKFRjNyIk7mOExGTaLTWFX+Htbevd6oRfRZc17vFcpYOKVi9Hz+38sRzZF5F
gDoAOmNIuLrVWFZIILDhxGqVjT3jluRJmRSmq5y/O1Q5WcbyJBmtGP8gPvG3NCm+t6teLkeYiOyy
fVjZgElgEXNfSCE2ds4PR5uL9oy+uWLUnzriXcPaT7YyMHlLZsyJ/qhlX5dLgC4ABVpW2ZhypCHw
bRfNzl2uuvCyXJTTwVbo/4UIRCw/uLjo6BWFEPAUImETPgCg8lXi0+aQ6oMxxGr2g03UGCjfJ8oR
QNwODTHndVtnlBqe/W/TzJ/KA2uFRkaqM/tQChTvH8mGnGkoxqA0MOMMZ88NXoSEePUqWmZTxhil
4UQaG8qGJQx+CtJuVI1qOLmNJRuAET7eF96XK6+jz/ytA2OygYzRKUYCqHTInw6O54Bebw8/uL8Q
Q1Qv3kX+qdhupyFHHsq9d9l4iI3zWESPExGckEbRF5MnA/xWhp/+CpXrp+W0unPb7932Nqko1dxE
zqFJ6uRS/1pi3OIfc1eMqKDtn4RvjfmPynu2pCyFRoYXRy8toV+Wk3SI78wcvTgU2EiL4cxz6RKV
eCgKc69c4+CJxr4IsRvKDToDcGZ2XOwhnOAW/96ZyGw2C2yXEhF61QJ/ACxbvGw0jW9NcYawlDKb
N1PmFGwH42AlW9kugwn1U3SkSqrB+chuBasTTLpwsN2Xgihr9nf5TX2s9AAHCzQzLRo7Aqga2PCX
qN5zDuCIHSE9M0RegJMhPcQMXPF46E4HVX7Z8NNN28UdSEjlQABB/RE+apmAyjfZ+pv6s+u3ss6x
WwtWbKXX76/eC6M7K3MR1Zj/kMJod55ZOYz6LFcmwL+I/jYhLVvg/vzUJ8rd0fJ9tFB8iwRuN0ZJ
JLydAHHqXEjFKd3e01cQWbl3BmFAXVp2hlNDguVGU29ebknuFbqBNKDN1HmfchCn6LacEEGwTZAr
dEL9J9pdfSFYq/HF07EJaO4ffsy8//c+eVuH2NZbAP+eg0X/K0iW3gP2DqFXtTOmmcuF1xdiDuzr
nPdSAYwU/eFfJnYqhFCNqE8OvDKHJLRfpdNDuoX5maN2lkku84Z8r0dQjdq3t73FdRBhfOBnQDH7
olY/ebKG4px02QJtmcO/TiA9VQh9weerIz5fbUpmGO+0Bqi5V9LDE0ORnmmQ8lZPdjh9x/7SxLM0
4H4vsvmlRuyiTQ6Q5spUPr1g7K9FFKI/fsA8SQ/2SuSrkXj0hvaMbn/SvAo7i0+2DB4KMQJFqEhZ
WUMP+ZwGLWh7kv4VkpH2J+VeYYtLCbzwDB57NH54mL/Tcyiv/HCniQyozRiWf1SxzviszEnJv9hr
MalPX4rPFeD1D/W5gjb+xCvQcu953u47SuczGdqGhE8z3oZVL6g3G3slbXhDQZHMshY1n0hNCqto
q9gPbUs2ohXwwCAkStzBP02u0strD3A7me/bLvdneDwNw2ZugpoFihBvXBelGhKX/I8Ibo/bELGo
CJA7Zw8FprhrGbygMVzrSMrANNzxAqRbXAUxzJI7f+19AZ0aCRwOgheQ10hYh3Sl8loEIcX/nFgc
DMfCSEILmROCkxTH8o2HjtP04J105zwuMYoF+5crWSqA5EXe+TEOukIpfDxEbXSUSOfVUEsZnaJL
8e4OkqKR1R3yrtt518gZWG95D4ReCub6U+OO/ynqNYLJFCh4f4oGqN32hjLdPHIbHp/jz+91d3uc
IrwrmMj1JSOrMAtn7yaOFe8Gag1Iu3Gnaz3sT19PDZ5qhEjINzm5PDccp6RiChda2KEsRlUSqERm
LmxzXEEZ7GxorSAWw7jj41KmJqZ0X9783BnbIRXax8L7lGaQ3xrfE7xpGyWmClgNCRcVrmrW2Nck
2Cd1zljhs7Mk5Ipsq0EP2e5uhy710bmZnxEDFsAjm26l94cOHPzlLDkqddfXoJ/+LNMPPCWBVevd
+CCudyTx0KwqotHjgQuYe6hud43KftLs4gw6YGfYC7WuIonLSRtaORljzq6Wm3bGC6gXyOwXcyNQ
x7brPKyuoAiFJcz/fwEAge9/9yDUpaB6zXn/cYDadb7nvhvuANWqxHdLrQDZiqFwsvG2AaPa6toH
OX5YT5JIkV9fRg0RnwOtvipq7Y82vebp6xsNealdWBEy76zQUKg7WqGpk2AJiFUbxwTv9yPX0qCh
mBQ8+2EO4JcbWEFSztYxPxx7MSkXZXPRYaT0ymy8YyLNk+rStyzyygerfEh1ptmJGXLrkM5BCTLc
hWWHpywliZkZXptcDBUA6vZ+fiGqFzCBEvkA1+ZZ+SIdDGUyaa0skEODeaFgOnuIzrwv8dnvtfyZ
82AbXFsgxEQ7iw152syqfJunsw/x1imgf5yJx0y0BNVQVeWITS3/ZAox2YRAGOpt2fO1OX+I40x8
bxnoMVMTnAXryBRdwFaYcQ0bvUe/E8gAuqNO3JhdYFsxhUpsUxES5CXE+9/fB9NMOv7z29o+2fu7
gNGPhPy5pqTfugzOtX5is4rRTIZ2E9dRYOyBxAAunC3pHqw1S0Wy/Ew+0mpZG5j2mr9IbDPLDJO7
lywky2MYfaLNsrSC7Ryc6BTGvE4eHiKo/N1pJAzyPzNfKpUXt573xjnc3DCp6I4jKAipN7/PdB0/
h4koGT8y193KgB7zRjkttsQJxaGvdzbLUi2tyHDXwsD8SjFW4WFPz/i/tnqlWBqwj3uE2bz/gg/5
mTQWXK2rIzVdq3wbBhH2FgcTU4z6qhNla+TOWSiS6Mz1c2ebUzcfUq78uw39/1aLL0x1idATKm/7
xX8Pp6hpeupW2ee3REmbXtT4/I/mvZx6WQ66iflYg7MkbeLUX/LGJ8w9+7rNHomjUtyKoqpifNzr
bYhXi1nC/MrWAtA7pI0rALJjO95hSuruCqPyKJSxfJXxJH79OYHJxm1jfqijehDorpEK1QUvMKtc
VvQ8StucPgxSvUcc0LfuixlB05dfc8l8ANT03QX6NuoL/RtERi1kXO6L+j71r1FgYGUTdEcFLHII
2bYX40BAAsJIlw2VpAbnjOb99fripkYM+2xD7i7Rj38xT3EBqwl51NQKUuY1EjAMjutiH8xXGMXy
JQg8HKx19OkpO6s8FzOoSFoUP599U65EgN+exoX9FZCTskwaSVsAHLjIs1Ic5K6yZy2ks0zC+/Xa
IwQAOmFQKyqqjk8x+plaRcBB5kkPRXtiM1U5EM93u8BnCFD55Gc7fFHi0C/stkDm0PF3S6s+MVnJ
uQPNQ1AlcqJB6FQRbvRONZWnsVqTV180HTjnWzR5YJ6GXFt0tj8clKkYRFwhGusgNMehuH5PkwUp
8SNquMLcvc7V9ztcShTuo/fvyOMCQmM4fQ2Vuku/7Am9wtfqN6abMFaWTYiNuUAW/7m++JcInvLE
KmZQBp1i0U9i6P30AxyQXjbt9f+VwEMnYr4cDAPJa6Bz5aF84Whggi/+TcenPOLP3OUN5K1hp+2a
0sccRzR4ISAOgpUrSZCa9pXzgpr5fb/LiAEW5xx/69XNEvMc+DxQIx0794Dd3vSt9Ihq60NCXmC+
WrJa749feiggplQ5m0Ra7PW7B9t3m0V8Vr4ffsnPgx5IY8w3hhg1fHohkTuXASQlqMK/njtnFPD2
SC1olonMGBWRF9xJDgg5QTu16Xn+++fhpDi9dO+2w7Cehrsaqw1exiDbsZeB8Bqb/nbxAqVyEXq5
h996VRYS72jbTRHBAbeZYq3y75Q2XqDKaEw3n+guJPRGHJ14zNMF8touVDlmpf7nnnS2eTH21+do
7ZoVQRxKGtLrzO+ZsO2EXvGjiCWL8LcRTu9BQprF1brkG8Pgn8hE2aOZmHwqoQGXD+81G1mJ9CXD
vsXr+KASsOv9gx8fjjhE5kqKw9kvgzfA0QU6DnIiC7c1MOEZ4MuhUMCixK+De+H1LdFOqrnoExDh
nqg78HO0GdGQo6jvOHFH/ZD19u5N14qn9t3ihjuSAdGNX9hKGG9jtWWBIsl4fUCHiubh8BWnP7b6
c0ISEO0NwKJwkLYlGNiQUX7BURvikt3GHnny3MxQwWIwO/4E44xHi2DBJK7byzVs0AtRDYYkZLf0
lxJiVeYU/Ne/ClkSAzwZBgwFBv3pxq57JYfHhds5kfRV6KEIu4kNPmaWJ/HuxYF1T6t6Ob7vE4mc
Efu1YkEqEAqkbIwwEXq0EtV48u5ZFobZnZdtZ4cTLZA0br8l+P/vxo9MIzaQM25xOHZyV6qaO7dR
p4eYVjCmXM+aJVit9eGc2zSszSbVBVk6+rzjwGdpQAArUBm7NJAqw8ilpyGe4bHHJgM/PuIQAolZ
TukqaxghJmVp0OerHxRbxWXoeqU/AcHRj9h4lfZEG99IOfyoxHDwmWgGFnepezCUzzc7I1tsu6BF
M47FnyEY/ObnbS/b7qfbrs+yiJ4RiF5mvhTv477kbrCF0NSgehX+DD8j2V6P5Od0jOkLvL5jkYpE
QGVm1n/UvRALzWz/OxsgGNA/voEtTnrZ06qo9sb2vLvhGJBk1VzD8/Bez09A7dTdc4MUgVl1mdRC
cTNir8vqsgcUK3A9nDBTIJyvchjIHDV4818CfMI3TwMHALx0eXEyKXEsOEyaLlllPA/oAypFG/W1
u49HkktDXxyBy9xxYnZTCp2+AFZxreBnxWpef6dIRVXv50i49LxEhQZasxl5fK+fqTFmHoh3K8Zj
5v/dCbwvKQT50041nQuD/qPcQLBXp9fD1jZ+tX2nJG86YIOtNB6/2twaulG+KAq0GRzTH+QDTS6p
IlAsIMb5Xiaw7ySVniJRZjnFVazR6tZi4YQB6+sWtT8TfhibJzfY5vmWrpxxBe5pNYXKQ/jkaM9e
ygv/efvRbdk2AfWpPmeg+VI8H7A1h2mZNyfij6R7cRvN46RM6WtdTpbhINeXIqzTX72/yjoUQaWG
sc+UiVSjxqVtjq+rRsoBXIxn1q/tZFRIG0ytW0NlmfNoEL/EbFYmOwmbHIxgouJIBRFOvMb9Du8d
dNiCayLOv3/5WxIsSgHS6d/APN/aHf3Ipli1CaRvAOvuwKttGO1zCy2d7zd13wsanIVjPBm5citK
0DxDtUu4NbQvvXTDRlNipYjX/eZO9VmG+wSBEgYQLzQJDV84XYpeJKgNkOwuEx0FYXQAlY1iSLe5
+K9QC+90yBWvvIqslEn3nsqlcDVPQXmHf+56h7UJXz1vveYrqOcZDM+BptR4DC91nRBE8h3T3So7
XRsE1ZEJEavcPDbCistzfi09Z9gOKwJPHiGJ522XWm4KKkSTEnL1B8UhoeHVysf3bE6Feqi94/25
26XO4H7vpm3w1Zc0E6zFmOppYnAWsYnGU5AE4COwDELV9DMNl1rrsb6b2lBKkBGhqyrWBVvU8Nx+
iw9MlH/sIkwaF4yZQhpJFXd6vj3rSQk/u9QSTYEmqSbv47JZ8hr51bVHRolvQcTlrglFVsLYUsBP
sit/Mp6z4vPE8rPtGJc/2Ry2VpaiW9TK9rs0VmzdgQVokyad5w/yo9xfcMU/F67VkQvE0oHYxSZe
Aiw516tQFDAF810C8j0eEa3SF/WiisMJkouiro4CBgvl/U31KVnvVYhMQr92BETgm8Bpl/sKD4zt
h4L56Np391lQVPDsWYPK1Ee2GgkNG1V2gv+hPpV9E197MhW74gl11YoHmzH81gjWTZlQS3soKfDg
AmlVXhS2+3WPRrqVFy7b1eFv/7RJCOuwlWS6wt7wzEwxoY4ChWOA8Er0kWaTFDmn0a/kxQJxcOcF
vH1NH8/9tshSxRU+eqWgMSjXcosXAY6Bg/FUed8S/Xe4PbVYvsoAkmBP14m2dmp2YSpoFcKQiPub
cG3LcOVzTRvgn70Y4yyujqRsLiGNYlkBs8akcWViqvn6KKoI+Q+Fqqn8seg9vs5if1doIkt3z17k
K0lIHf30WK4Dv2PHReJFCAXKVUtofoGSoU5b4I1B1X/IR9NL4eTA/ZVmuW4gqhxNF10MDneYtQ/a
+mwU6Y0OhEC3E/mS6Cau13epdMCtMAuVJ/rQvW0tvZjXnjWgsy6HS+Nx6qxbQWIUYk0uF9OL11vQ
EgXnaZ+ZiYHgXKEAxac+m2Egfr14k7o+uzBAufisilSy6tLLuFuGrCrVMT+Nlph4PhUwMBu9J2FR
NiIBtd9SYxDvxg36jcqiWNwhQ8XZbU5gpgqVvn9qs17M7yFzgzS4GJH7+gMVWmUXQqciMFangQGD
DCHU7jnPzHaneAgazbmP2olc8imh2W30Uh7CQmy8f+OlOMDL3oD0l0Wty89cDxlJtwPzD7VIUWMN
hJdL+Bq6srzN9I0YjIQCZaenBuCx2xAHVHG0RmEFx48DLfucmddHAvqC7Qq7Gs7/YeSpdqax8rAB
x3/SRLj6ox726+QbwgkA3OiEyOcWk28Q3ZlZVBzIXzlLNcNO4vApu9eIrqboOqy7eTuTi597dHyS
3Z16kqMp4ladEdA1vsBGYARBbhp1ZKHSd0C89/kYbnqrQf+BC+V7e086/yBV24yQzm1ZBRDhdcy+
rqyitKvRg8IXLYb6PGQhnfLLzAqaNo1vBdXAZmKw7puKgcdTHdUre/t/BqUGJV6hDSIHljrZoScq
h3aUVUPHLhuP0pp94uFLipQCe2Y21//ek3WJeuRDLj0CbvFmub0zQ3bDY+MwIt8hDJopuZLIYhQt
6HvJ2OxzVJEfBpRVmhyfcUee/7FnsrzMP0M12boCS9oFZZTbO71OMs/qfKAMdcG5rbmILs1XzT8K
nD5duv80K4Jhv/NWeLb/mWc2K2iR4WciN0V9IZg4c0FYCxpeJ25X5WelhXHHrNXMU7qlnMnSn5eG
KdiMb8Od3KlO9vOKhnRH9WMTyjbn8MSMxwgbw4KYtr6TSOpVzmczzgtBEPEm1MJBOrF6nEoAdXT+
9ivNJCdKofkIByLWVoZG8iAhNRG1v8KMiOZVLYgdUQh52LSXsNeaZqpC2UA9v2p1OlRxDr+oKMEe
7iRDaPJzqGjBePX5Y2m1SrQAD5F1NsTdUolLm/eXAAMe+D6nyldCHumfCPzlHS9CmtGGHqslqO7w
o0GiouX9F60WFmACDvpJZ9X8ebLSiEGX0ehCe6g4SJJt/Cv+xvHWwdsxwqlAPJ4SgS9QaQTEFGZm
sel35akhxuzh9bVgoFb5RN9itv7XIw0fiFtAN95+hZsOGJipUBecY3PlSp4RhzSNa7V4DFQYu6Gu
UiMQZUmwh6kDnsMrkOUQoQweZVdn/u19u7y0+69gblojv+2Dr+Jjhz0qd86Q+mhqV0SrLp5jUkQH
DBmWmwumZzN/Sm7CviRe1vEu7fiRlVo6oQmer7sAm9ihzuyPgtbgzo6PttvrdrXB0vX7utuEYf3Z
0CkPnphdUYm+1M1G8PrPhGLiJ8UzTrCp5E90WWCORTOEgBb/aQyQExDlztHJP3uNo/AfzGJs9SCa
y6+ksSDYamMZJWDe0Bt8T8Fwo943kdZQcDWB10WYji1GW/mlhsvCbpTaWzYYIwND0p0+DYiiY3z1
N8wyHCoOwdK8BAYBP2JbcjBO3NjDFthMgOOmzbJ9eyRumfcTFQItrIKqFzeGJmNCsfRYFunCywNA
HTcWVce5XJd2PX7z9JOweCnj3ual5jVTpDos0ZRZUCY4W3GDHs142VAjaxMCsBIMiAThc1J/YxOT
ZWYcdYCNoyrmgAxO0lpQM1moHhJ4gl0ZkO5vLVI4lH2653lKF4ysq901+/nBCOz9P0IyEuDBfoRk
NYpbd5+XkZwY8iewOsaJWwI7I6yaqraxfoq+uvVNbtDK6Y3HW7pWgI2whByVef+GvtPFDq4r6Uqa
owFLWC4070mtNajy/FbZ7a0QZmFDlqp9m9/jH74m1yTqYIV65MBUdvgjzjipS/icAa1dLyIq+HDL
WR8U9k3rvoxuesCEvIPIL6JvOqMEjm+7kXve/djlZBTSYzkqcnGUM2UnhuSZJ/yNM40xL/0qtBxq
1YKHTHTVrL/MfQaf9KpxEM9ZKhT48UJUW6oiWz/GbNt5xZwJUzFluZbc/AGME20/1hlZQg55M0/M
niMtZcZyCmy9cg5jPU/fHg6/YcVS4bXU/2cTdX9yzVbHLUQGZQ0/vZgg6pt4XpWHVio6v2qrwUbn
tHhRNwB50herhTEmAH3L/hPwyjFZYop6AkQiq3GNe120XFefwb5akcuadLylFRy8SDMIREezm4Bl
fEhWSwTULWXjWieav5jGBK5ClcmRHT7F0gjIFiXt5Qm9V9kn6q3PlPdAbfsM2r4S5Ob19ru3r3Dk
aOIFVPBI/V/tC2tmyJJt9ZxDCWC8ijfpoLNwcNnQ9xIBK36AUs1vO63Jb9nneQJX3+awyAis9Jj5
uUG+9C0ne+rpB8RG1mrPvemDdUwpr+nIHF+83NPxv3dv9XODk/MOqhsBKJ3mxlt+2FTP2b5Tro16
ozCRoofxsDPqgagvlwy2W6VEo0YWeUsB1BEg1EfQx4axH6MwjGIngRy8Y3Cnh/LthT9rXLkh9BuI
8j2uWDNSaI3tBALEua8C0RR8fiSlWIaf8xSRamTGEXjN5hM/8PKEufMEQobPRtYk9gMh0Ak2k0Wq
yBqXD8RXhyU/HalyX6RjkuOSYRLw12aoklfgSiitl/hvEIhP7RtPNdrXscxKvYNW2mUKwl8nrTfQ
85SX8DqTraHWy+JST1zxo8zwWf/Y3tBUAd7nAghCYybwRsIuj1q1zp+p13XmaJH541QTUdArAdbP
Lxqv8+pFJCQ9s/+L++1fTM5/V4X4jTVf9wRLprRO6MTWGijePygTZ9eImaSd+j0WQoDlG4yn1FwS
FHWDaTWNwzw3eWXRZKoSHOfLk5OHMBQVJ172S+7huO/P6B8rpkNhWZbEAXXRb99rUSwvQatxSXtn
cKCWJ6SfwANZdAESTZgWq5D4ir+Fc7XbJL7/Xgk0Hpp8Vpt/xeqTL+ip+Js4qr/l8NIHUQDDJRjp
BhUEr6SjMzV2PUfit+kQ/igTA8NmWPxRprh3/aAlDs9YGNlOIhBhhcFExxyXrjR3A0wKzik/slWi
9sHHUikFklg4dcq4vskKIs5sikz7YoVDMeoifzU9jcRr5nbC2TZTWQ8gCzPbzZtwl5uvWENEJSmU
nT08x+iORcUEVYhp8yMGzwh+aXjktjNwZZknASgPuGO9G1ypOAVbWlzy44C/BZCDfSx+6xfp5L0M
a7WFKq+R3vIz5IWXqluBHsoZ4BUci5d1fTYetWBzQnEDH+lPEJG0Ds67BiVlYBGV1HgxSQVUWURe
mOs/h3CifiI+8MxrW5hphRUTG1WM0TXeJxWWe9Z/4edBsrvcvex9QBVQcQ1UkkjStf5kJ013Als/
5WaadmfTPFbsQvnTgzyjWan9mnrpoHScnMRvboSIKgTGxgbPB9o3NthBAwLwhpybR9XiTr0q1MKF
8WGjR8mDvcx0Y6fOTbhdx12D4tdCvsiMzeb0p5kBIxKAScj47HQoB5UzJ+Bv96n/HPSClg9HI5mg
nE2Yq7w1gSSZUOCtlgphDWhr5qTSzsTm2dxvbHIgWWeNxdk73LUdMo5SUuB7de7uhz8wFN/NXnJh
iCF4sNYM1TIyaNs0LKE9WR1jRPPBDf2PqkQp3BnQqBnnWF6rSp5JscHaMoP3nQfac4Kqj167xVqu
SZzwxiPuFLxVNq6pnyuJWLxWGP9IfsiR8p397dhscOgCFflXvGcsq5S9SLogmCkam08xExCU5HlH
WCpazcVzwVz0Sy5D22JRcWQwH0nlj6qK0zPjATWDDS2CZ8LKgTSWja0zqdVJdscfqVl0cn7DJl+o
2VCVvfJPHG3fPaTDTV8xnv8v48Hgv9VOZqksWhLOeH4PvyW22Q/cIla3i4aCg6h0PIe5PSVeUnRT
5d7gPk4DhoWR+km0dJONvSl8oRS63V9tmm6fuYpNeaPBdZVC14gfdDb9FZjJ7w4qIel+GIJ63f3N
bjwcjGuUa4MwCBcCrwZXG7rXpnrsEuZ57e9BBPgfVC3GD5nJe11fh+ei5KmVvtdYL01LUZJw4JBo
dZWcVfe2iY/z2rjyfROvG6i8jagU8NKYe9LCY6yLrbZWaqLDYP+cWRaPVtpvaTltYQIpagqh7FAE
Nq2oYCGr0xysIQMUZrTaCrVRHjMGhiVCvrokj7zYHkx1awQmLcHAydz0ltx147EKRhUdwtFtFJfP
o4Vj+DXGRMs51/vYL+rUJhioZ8U0xQxzR4CZt+ggFzW3tnXzt+WJAdRGFwRLx4kzLHLEcce+pp8P
nBM3eGlKisd3nR6aJu+0ICmhsxoU45M/pZYq7E+e24AwD+PPx4M8+ZpSButBVcOo6uOd7QXUDt4E
Si13Bt3ZFdy0qRNcfntFK0CV6qishGivpujz6JEqlDpKv9cyWlKsPozL9LRa1nhNy1N7gKRbEy2t
1sjMMFo02VPq/+hD1pYIe97otd5z8a3mkaTGZEvxYk4fJxhqp3eiC2G4Vli0CrNfSVRwEWA8L6fD
4I+C3C6U76Bg6k5PQ5EzztHXt+Wb3KzEfa9FpSbt20epf29Fv+CFQz9ip/2JuMTdxQcW5+uDTomx
bRkbUDdAqGvMHa1aFTi0c0/hE1GOThofdQDdFxFEo/+phpvPxKpRr5IgBU87kr0vCYPNAzvyB8j4
YsCM6b9Qb6nx/RTEr1Jq38tGRKgzezcaNn8FMoUxUoobJJHW0dyCA//5/6rqaMNYh7HxCpYphYvG
A+lMY44M+AeWzK2kGEOnJ484xSYdVdBcNLj3cmYaFp7yqMHT++ol925qC1E5rKMpWz0SKd25Q4wx
Bd/iRM2m86tqaTm4iwm+pYf2NHZ7/8LTuevTP8EVg+dFlPcm2mryepUav+cWCPgVvfvEEzdRb9Mw
WuiLMXWNXVSRHCyePen54VoxFLxilQ8MtzMzp/YoZF+WEgd7vFQ/5k7P+9dt61p/SS0MLPdQDeA/
YGFGvpEj1Ne1s3m8c18DAELvB/48v1zZgdhVc7aOwUVAWBODyzFhXOh84IBTQAYGCll35bf9MDMU
NrG59C77i8LO+UMHBGKW53nL5J98YDPKTfo8TZUX1i98Tl6UBvT3rTU3yv1vfpqQ/MmUP9Lv05zH
NVRrDiaGO+/FXmJ9nPgsksGp9qWFZEp9uaZFXtY5QukTemre+1m7s6dk3L/5pS/WQwqU61oFi9oC
BlYmFBfni9rCGfcELTk53I+n8K1slWOMeuooMbar0LepBbk0SKV04S5DmpoN8EOUNMh8IeZw2I/G
Fldo/soBudz+S0bY0CLOvrJA/bajK40h3GlN1eS/famnHfFBivVnGRhOpwaXlKGw9vetIF9qElKd
f8ar1vTli70HlY871c3s153IUTtUTUMxI8ZTpaE/z2i/POTtxEpHGMRbyrGXdjSl/xkO/JN4Tzoe
sjT3z7Q2nvRDw62tPqaBQurpeDaGQC1b/ZiT0S9wCaE18NCGGUP2O3ZsppqklboFis0pwixk3xu5
Q9/LZ4URBh7XO1Ya24JCcfxAVinagslxws1vyGot2bJZv+MXJq2y8IjDd00XQQMS0rpJuqb00wDR
FzNb1hW95tmo73ym80C7WqFeOoC1k+xX7tpLcxE6ocd8YgRbu2AUJqNsLpUeLpkZZrYO9thXf4//
hrRx3S7sr5yQwtaZBp9xDNy297EPQvbGeketNu6pgNh8+P+UGxWI/be/blrAvJ68+Nto499OjKAY
f9ossCWQvoejDvp29wTYTlwWFE1tkGZddr3qVSAqMyk8Sb8dZBhTYIZPGsXPcAgWlOJ9kQTcUrlq
wWNbpawslM0Qp0/nhHH2u/mXTzwEoL+rn0/R4vztcDl69FeoYuvU8bEWFKL5II5MU6BYGu0U1ieW
bwJwxeCXJUax9n3aA2l6xNW8jyW0DO7svQXiemc/Op249yRG8IJ0718naw2xM5EovSpwV5cliQOh
n2icLYU0lygHbpEJQcNfoPgpdVkTz9FPcnRLQgnDzo6VTk7HhAbDRadPA9rQrsGozWLJTBerPYDi
SngNoavgSwGSr2bl8YW6gaMWsmRp5XMzNOEQVIxxF6tPc7ry/7jQ2Y9G+bnNUfHLw2VEEOaR8Qgb
M7wAwQLo1EJEGeSSp+TJgCR7TlXAvZcE9zEgkNQ67qg8aTqlk1Bkt/2uvhjYfjosfFjNz8n1sX4T
txIB67bp/t/NS97A4FT9dKQlxT6WdtM8qKPDSbtSulbQwBy1Z4QnI9JoL7NL4jqsiTRQArxMnCUG
WhGlC/vZj1W1o4p7ENMjp2ssE87o6lGeUykKLFhrL/nsli27Be3NAvZpjoYrMF2x4yUOstAeDeax
IDTBT4F0ENqZnvmVlXzr+VG3JY/SFlmQaR3bBm3aU/SvonYB8VUkYsAYJFdZRBsB+oDRnO1vTelI
MfNyr3scjyqWU49jEdS9/HyChtUrBXhOA0N3gUlP/VtpNVzLVlzqIDe9/Yg2TuDlIyaOnYEtyTNL
4HtFAOWGCuv6TFSrB9FyTcwMsWvzWTLB0E+Akv68JfIbcENviOT/BZicN3bwnMdh1zqlXMM4e2YO
4cqwkASwM1z0lGLUDpmJt8yQDSLC8bWnmyIKkZkUNY5r/1wSmjvDKS0lYlPy2UqnYL8fX6Kvs6zG
m2yaEVgmn2d4zx+Kb1ZOI6EBM0JUhEPrKnhAL+pWINlarcNm6FQRBoYe4axyO9zvbnHc+YJPN4dA
C0BQAROaCOwrZIFvsRV7Bgarf5U/ZqljvH/IoE2YReKCjMkUwgKRazgsmHoLEwnlvPqAY2xO7Zck
IHFxhc0eKgtfch6Phd4ARgeDorp0N0TXZDSJ2H9o7Gph9fc6Pl7TaLcw21PUF0080uul/b9fIIlO
NFfWz5+ei4o4kXPp5cYmWyJrrtrpnPhk3nyrnMT3hE5QEsiGYlIYHOuX1d4u5B/pPX25vDeKG6fv
8ARAyC91KpXHkuS6FSG88wRwfhsGcgsL76fvNZBYMxglm9H7KX/JbdeZr3021N4x2E38Fxmz2QkW
spk9/IxcQuxW8HqY4sJ+pP/+jRcD6S1/hL4P0pTShZB78MOP77oA36K1Nb3cPeFReobx2/X7ZxSb
szgU2KA6qzOaCbMM/Uj1rJqPeGnZsCkDt/MBtLbDY5nAu7Ws/3B1H2G8A9e8QQaKlNvs/N6C52An
iBAfleT5Eqeq2hbotqMl9Q9Mh/9HGWo9/JFgkDFOBJ1oyIPcAKJJ7qQ20e/6Y6WWDHQ1UrgZqdM4
DPaRxM9VY+a1SZm2KO6euTWwZ+8qEoG9waPj/MguzudlbFux+9RgnWVuKLGQWNV++m0IVtyGYLFq
UYPs5ahh7PBEedoLwoC6Um/jNV56x2D7RicWDsJ+Zqib5z4UOqKeWO5cpmLCjd4deBcrtsQBZbE+
StVe5rAdtki0WT43X/XpRwmelXyVnQDQ4v7dmBrmFSn5gx+xSjzkZt/y/uaFJI4YrcVGhhsAylUJ
p8DhR/HzQvInmIQA/LzL+gbzvopO/WpcaSuFbohIeTNtMAJSHF5qSAbzd9OOmmTYuiHsd1u36rZw
b3odNfS3lUviJ7Rpn8hD69C3cTBVoz679inb2KLAKgxf21gYLYjlwY5kaoe+vuGxuhorTN2qTH9z
AeEGcGHUGMci20ZBAmvAkHy0/5cFJme3qB+8z8l+9UUntELR4FZVuiM8EB0iKJ4G/Cx99OaJI734
tUKb7cyBPVXwCPrLuWnFJz0M9Xt/7/PzPy54sliwLTz7lYuF0u7ZOBLroPLJFi030PCHJuM30YQt
gu2StGBbHtcNx7S3kG/w2Ns5+l84h4/p8FDGwEHzNiMCR73IIFWWA3hGjkVwAG9iUh5PDqz1uLVz
54tV5U6racqWMWXnLmoITmmSaAQ548Zou1aGqDlY3PjrDaVWx/iD4Cw4xcyrH5w1xKJevRhkT08z
i6UT1BwCdjpG5nUBt/5dkGOJ4QJi6fFSv5ann0cJBWEMqDb0wpaF4+9BUSNuXqPqWQnlpzROvG37
PEKoPvBqOvk725PXWgiKHnM9z8ALA+HWtDcytAkknpBHtW2RZ+11XwGNYL8z+GjX6FdiIcAz99uO
yYwdeKceS8ZL61gs4os8syFXbEa0O4vI1fOhy1odfXs3T4OU8qVC1QcL5iEagrGURUiKfn7gs12T
fXck/LjfLzwazMjMg1wLH05KqcnojN5G3yX2XiLyHgJvLWYi/nGJoPRKs/J4qJEK+9CP53uiF5q6
H/JgpyRf3CS5CN6tdtTftVn6Q2NkEQWx3Ujxc6ZHzvvb884wD2fMf2d0Q5xrJMFrNob29blUpK5p
z92bRYJA9GlQh3e80OOACS4odgPupxpUVTt+XOUd+x9cXGmrTOhvsQZiroEBaFXIEA5IhxEEPc1g
949ah7VAsRrKErK+4NiEI2lKyOLwSN5reH+M22IVsuUjaYHZSZnTw1JrQ30Vj3xi4Ej7lSajsjJh
fVD2YscBzyON/T30KMfT1EHaE0Z+JwD94N9Cq6Sy+oh3kXxWFKIJxLFfGlV9JAeld9cl+T9Enro+
rkVxTa/ndmH/tkIj9wu0x8BrzQh0e3G0k8l16BH1lTUzzU1FxwkYcWNhpchhUZNLC2+5+9lRH92F
q6tBr3dGJ30Jlydb3p1IRlSzTscv20r5TwLFBhTvhBmqJg302SS9auYsJu2i1uz5/eHiRU4As36z
HccEKMny5slwesRMjTcxYipb213rjWnKcw5E27fTNyhSkOTFcoCXQTAOKEyysWTv2h8vqlrTxxGq
HChvH7C8HBesEfHi23tqp4Us7/LcTNvcULMqYMrwMCKCHB6PRFQQ10Ys+uT0ujmlSLTeIniayfwk
tJzCJ2rg2XJZon/MB1h4v2ziSEq/NDXot8HKZesYkTFV5Z5Z+OFPSCKPUQ8yDHXEQNBoCp3WjOv/
gqLTJzcYezVRs+nRlE+qkdgHIK+ymd2aH/O8tvPzl7Jfbl03CNFNSc2KiDaMIq0Fa5MK8KQoSNBU
NBCStKxTXOrMtc7h6I5JeaSSXZogPuPJe9cTXA6U549ZM6Se1iIJyzRSm0AIR1S78YSfRtgCWENF
dAxf6vMgQ7rNVr9qUW+k2TxEGEFlOA7TUqer+5dwzjGQBr9iFO5x/jlC0uCaa97r4nvZpbOeblvN
krkejYaCshlHzFLf6gKoab9XDcosgxP+bpMFwaJ3pDuErJsauXOXWyaqSFH5LOWPE0ccbYBLzTh4
Brll9Gymrz84EnkBeYIzWTt/7Ah3xuLoi0AefJk6ATfickb3f4RVK8vwJt3XAi25ZprpTBYEAbCq
aRK4dZ5f74GoHd2Eoy47GKFPGeld16yJRv8QvdN9YGGDiC9V5sGcElmjHI1QjEwHQqjDEIpus9bx
MM9Rkw2jnsZDGeJKJFVU73CndssjmJzuumxwtdRdr+EqKvUFEj8TUEnbvomg5BME9SzpVKVmDGhG
ghRrLhJvORtJBX3pXdmI34FkAUoIwMHeiuJvFKjiIIZP0w66ceuyCZiYfHoVB78cM5gSdRM0Np0K
10Grdo974jO+L6/uEYL4wnhC5c7E5hLtXDwkf5D/2MiG85YghU68hNm2RO77BleLfaxzOAdMywWN
gpusn1BqHfiHw9IKx2btpYbXW34Obwjc7GXUjHgi+fmHehe6g2xMctzBcG244SD7YmSSHrq9NarD
dUrtP4v7tGa5Q2pZkjoq2ziIrxI/2udjmuMJaf7bPYQcxisEV07mEpXMWFEmwbAUd6jQ0NeM6rI9
o5UDPQmvdXjIS1TP8V1XMbONmj1/sewLW5hvUxVn738maElkWdsGbQsWc6yTP49c9pKDfttWc2w3
93HGo4qqvzR4k9iEqbhh/6xrW9aLowkfgxUky4GuBeGtCq/n48Vv42sgLTHt+zYh5yL+TH6tK3Jc
/6tGcbFjA2S4Ifc+jbJ6jeLN0C77kFFUkxrWdG0Js410NJgudJlAlyDxdzWFmwQmcVpr/Z0Ir1is
ARgAEqN4rLCy1KVlO/nsOk+sjoMysK4O0NQe+Uh5MBXxITb6W1Z8FmIScwD80LdQQpAdP+/ulHa1
F7W/2AMgQJsYnXJlqSdfOBOBCYDmTCsOPXZhzLpQJUZKeTWgJTkdTbzDMGrq5X59Gs46n3tHmHiQ
1c8JCflVCHdWsjKL5D/g/GRNlrIn5hERucQ9xGJ6AkeXPs3S/EiMzQ/2mX1yBfflvvHSz5sKtzDX
SPvGdQWQMhEDsZC2d4x9F2slRzHNjebF3JGFpHTYif1K79otFg/9pE1+ZF0+jKvUdi3aqeOmuxCI
V7AGDnuaQrF9Uqcjx6/CCtMGWQB2kd8VUA0pR2Crpknb32i6KrRpmcxG8nm9867Fd3YJO8ADJMGM
7i8p6FiKb1Ls8s/nbWfN5P+ZPfH1K+gWmbEqiqv7906vivk/tykcFVB3dl9p6yXhI/C4fDcq812O
tMMxGCIVygEApD/FzJkGKLuno9eZJyG9fDyMu5u2V4TrJydnpB7rP5vOaVL7dkdHGXZTzRO3Spuo
EY+nAPtbxxjQbwbpdN2rnjgxvKRunpwViMzYj8F5bNb+tQm5w0g40UE3hrTtZ1iROUiW2x25Ymow
hdb+0Zi2bQSI6F62w5rjP0jODARehq0rY29X7WlqIY9Mvhpk9UdIlU4Qoxxvo8qOMqHpr2QiNrvy
J7+D1CLtQaz76EyXhjorzPGhLjpH4QZ6maJkHvtoDsPH2s+Qy1EICWTy0ZptWyNj8p54ActvdVcI
ZECg/2zVnkqHWGHwC2bJKS3tZeNX+yD/JyXHOF0meheOGOz7U6HiG1tLCGv38PZgF+FQvEyW7+P7
e8EK/onfHptjRdyON8wbczgwOqsz1/PZEF9jIouddYVXABf2vD8AGvCLvEsTVEM8HSRHJQLbtMRJ
57kDEF91/IMIvTEHjjdPxK94XeTFkEWgVgS8GhvUDaYwzR+sJEtE1uD7J1WkPh4QoehVD9Boa+Zs
2RUfekbozCzYTh2PxKQ4yJtR+dsq1gqmulPS8/v6Nfh9WnNDoqRmS+rW0/lTEAj+FweynnwDX3z0
/89lJiDOfCk2koxWIQJ67KOt2N2iq1TFAZYLe6FvNJ+g8A2Akes7lT6CIUkJjE+DPf3RMevf+aJB
l5ADpFN++c76K+1UWDxYKBlnO9mbLnpZg9APZIIykkOLzXpOC04s+QkDZqSYCJhWP/XX7zvho0I+
cEfKqkl8zekfyD2SvOYSUMpfl/1wieMqJsS6D4T0Rrxgn7eZ19H39u7HipoHE3P2d3jNmRv4SXMk
SuIEIKB2AX2YGb3zoj9/y+bdTv+cAXwpZpFLAMAYoCwJ5BmqiI3lfoRTUJRbBJnKlrhvXsiW2Yhd
2pQ5mAgED564Ks369eJk4+i1aBgD+ezboLDYnftRkb15FBVT271PqYldGu+Ooqkcuqrnt9gLAxIj
8N6i6VuT806qaQSEiI6rQPdD+cJVTi9LMmoreT7/k++nG2wPMpoyYqBX7fkeTHTS5aLKBVckdLHw
SSVOmPADZd+jlQUhTtpsignsbBwoGRBNSEz4ca7a75qaopJFaMXbkHgn1CQmrFj4P2vupx6hKqvW
FZUbRyNGRAeIypbEX73Lhner30oPxty+HX4k94VNSZODgaCAsWi+oRzV3R7TVQdhTy9IbyvnwNl2
GsfG8uVfEsvAoY+tyfgKlxJcgJ8iMrrCCY9JaJfHzllwb949Qm3j6QRnivwAVUO+YKES5j3RFLyf
cdJEY6ZsusUZewlpCBEH5dgSBFXwRfmi4sRhEUk/IMBn6Q0lAalVopFJ6o++RKpnpZWsQ+4KzcWS
vBvG4/kica0rEodpK3rP3sCg2kgESZXPGHk/NsyQYoksP2i0tznCzVx16Tq6AL5f7FqTMERI0H2L
CfT+gSKSJ1gP4jxtd6IFqUFt4OhU7zLegCW/jJO0Gri7tOqNSCwyqoHZvjjo2MuiQ8lxxnK/rOTx
9PTnCj1SM/m1+Aryl2Zv1jvbYh2XyCso/3AcPosZ94tRgTLUeYY56Z2R67EU1vjYPxd8tLRoIUBm
DttibqdR7gYBI/mhXC+sRJGGKYhGlkXXqvTpZ2dYyDrmqy88VCJV3UGT+XxeuZWeM23J1V02/6Er
TI/HUjlRgb57rZyosXeEgJ6sj/L50XOs6xIwH8MsTRTdVsw9rRraxjyuODxjg5kE7U2xZCM6OKuj
DIK5HU3AnInWo/s14VPjm8hG+uPwgCpCe2c9EZi/ZrDi0p1X5lKOcTRp+5fI5VOqxlo7+8ozlm5+
kbrxZklQVonTKAMXc58o3iFPA+l0TTwOfUsodeDwkdGQU0chdTxdmfsB3+LPVgmTqefbDezVIGLU
ve5cuLeH3wrnRzz704Y1+eKIdkWsi2ofzpaSDVLSTJi6nUYpZLvetHpIHCFl5uN5+9LjKnCb/RHe
ejFUOgRhZpjlXxqW/MS0UkpddoHo7liysRJ1FXVAjDYNe7OreueIU0tPFx3vrGr/oxIbPnLJCiur
XMm/OqqqEm5clreAKc7H4cLTSoujnLYxYqSOK9r48YLfDw0nkf9YfmODXIlOTntQGHSZ51R9psGV
Y9Gy07Co3Kul8KqbaajPu3ngviByITc3AVtZKjviWX/BkaV9NvvKpR1tthPkPFSIfEjBzh8WbbhY
syM0rz5UQpBa1womIQajDyvZOWP6zWSeL1MYPa3R671SlJYQ/pSZO7hKMfvuL7VDnHAVs5/gdFqh
I/JtdMq9znnqv7XWix21+fAnkON6I5zLec+JdJBcVKNjAzlI8W2bLXOztSOCg0acTsUE5eGU/3/E
AhaDb39KyrPmneo073lNuDXVNhoo2ori/8xQSo+ocVMnvm5iyYcgn2LwMHcudZnhE75rm1GJDN31
wncjzm9PYSBmnWlCFEWjEIQHt6eXwFzLz7UN2e5p6wRgz+Asv5vEfpoD+91zP5qZLsGmf4zW22Ez
TfGPNxS0mjRFRKwtGDbQy6eYg/oOwJZKgzlF3oTJ6F4OeKQDE4pO95/30+u679daBZn0kBfx6z69
giUn0SMKts8GC8TJ8heuKZdy6bOeAbfqyskUrglVTMJQ/4Rws5wtI68P3cEx7U8kcPxj7U27QzQj
w8MaxmXJ85IhPQkXLzIKRbgQwzazPGxpzGsLhqAr9aNSZiP8tyHUutUaxJ/k7DgO7sPWDaeliLU1
X4HexmHDMWn7X0epFeHGHJD3oQYJPF3X9Itz/efTOZmU92MAuqWHWzkG0Efg6XT0lkrzz5+YeNvF
qpA38QO2o8kI6h3HWcp5Vd6sb5ubhgXmA/QqyWnlSsRtrBpxcfvFnMJznvXGX16HL4QMwJun9eAk
30xzJnKSoZ5mN+lAsN8KXqsY/C9FUmlDi+ygIFQKFoyncLRgvN4qeSv7WaX177ze5XPt0qJxKoaN
gGfLdyyQ86+1ZJpgFo6b6NfhxeutkcgjcH7jZ0FXygxIcC30AeslFSle4hzOwtRxFropiTaHXZPP
dmuCeegs0r9zRCgWySMD+uLz0Fn1KRDYAbALHHjq9IP8qhNNK/TLcVTi2ZsmIyunR2kSXJHnUuhV
SmRYoyzCpmakpNceUCASaXArMF4pfmVBzYLG32F+PD3WJ8X41V682meoXc9mcQsHGsX9uI/FF+AU
+xvERB0daGlZEOty+CkKofArw5nbM3nt+MrXPzW8wj4A5sxAUSjWxjqj49O/Qk57vcgNhPUAUckS
cytK0OMr46DgIDKirJtIJ/sEC/LXzCcBqQ5/LSEs5WyG3gMTXPzKPCuNAXf2IRfkfCodR2D039AM
OtLUmYoWwzR0ryWcXq1bkrjqLXW5PC9R8JznCF0j5WrZ8THILCBlTFXZ9RXp7jNXdAtAGF1V/rro
rU6HO6E6r+joR2a+sBuxCw/OK6+xTbPbCiZfv934wzJNqqedr7HmvRA9W992rUMcwIo5LPrBQfJY
56xfCKnBM6fv+/wHDWehUzkocA2VB0BSqxkYTf5ccJPFCBedIe5XgiPkPICCx2iDPSU2gdIsc6GF
7FcGX3TJEmCwg9qLpMgaoICoGcwocA5rFXnPROqWRl30lCuvqDMUjpOYsvt50vkpFIo024MwbzxI
5KNybeoKA9780iAi7uJ/yDDY46y2C3OllO4vqq/qJJDtb915VB8/GCsRwW35gUKCqnOtX6PLhlfq
S/KDrHP+fV0WGtAf93V6XmWpn/v/toOu3whkFJ985KQAwHs4l/KgjhPLs+88bJ3DyGL7LCX2Utya
a24TIrIkFbKlsgWUlnseK8zBl+Pt0eqJ6WDeZwzmFNJK5lvVm4zs0RksTgFXk6YYlixMtCv0q5yZ
RdkM3NyGFPLLBAZ4H+bPUm/B3QcfoVgk28h7QFpM/kApToP7Lcj4aQFk7/JqOLbgujNKud8b0oYH
x0Gdq7dYg1xQTu9peUP7h2lvh1HvHmwBg32dPcbyGc23lYFnago37owCCBzKi5NXX0kELAQvsWMw
TI1yg6bM9lTS2JYEdX2uqOPJCt/+JSsEzd1sPrPsrS8sP8bVRsFwi/YnuJbj9n2ZhTC/S2u60D9g
btOKaB89Obdk8Ar93qWknVzZV20qUri+URE5ovxj39aHZX5U+la00AUFKOMxQHB7CsbjpLslkpV6
Pa5kcIypa/RWJTQOfmNkO+stDmkXNyGKkfvNXeLx7LcPoNWXJbmaPa1ruXzUfIKZTDcfHwEFpKtS
Ojydo/Gu4bw84uQFcZ0B+GSfynoKC5F8ABstB/u/hoG4f/8XwO2LiJiGOuMeuvSbqYvcgcd8lGNe
Jv3oJGPbPB9es+cge3tcmisE1DqwCb/8NFuO+5ZB2yP5/kmUK3w9djmFdWRDWwILuhsVolqqVHZ+
gz0JeRmoaEFB4QljCWyVGXCjc8J6hWWJCULf31HKiqFbNlUHZDCxQu/Z9ojmbehmi6FSeDB55svo
QahVptVpCU1GX0+Aqg3Bk6M7B0AvYpA0e7SGONEqHfZMesZVSGfTbR8RmbLshqzvgTGC+CnXDKsi
CR2NcNwascWYnVxU0MMvW9LsnLX1pAeBAFmP+yiGFp4yDHZaPc2Xp8dyitXteMRWlM47VvGx5Pp1
tHEYkaXe2WuVXc/Ut4INA7hvoA/mOsNqMOXg3mpkCuvTxeXWHfNJmk0gPwd7PG1k4MCmO0lQMT3q
lOE/GDqGFaKyWEc8duiKh3V6Dj8Mhrk8+tinOpSDtDHp0QXNmreIATFFdN8JY9LfkNYwg2wFbwUU
P9SefLXvQGQtlyTPHSnU8n/kQ5TBtChmsjXFJ04J7jZ9SF4e2NgRx8gGc3hv5Sa7RJQ+9tmxB/Zt
tZaLIWjzjBAQ2G1Mf6Ja5hS0L3FPO8+k+k8gMlM1egqOHjHOjvQ6zWhNN9w2j4+skRZN64pxqvoZ
DyGCIByV4QFPmj64ULg1IAiZ0fTwQ53hf2waHhttSFQBV6t7hf5SznFHD7BsO9XtToV1DjL4Adnw
FGRBroRx42q7Ym8lKEzvYFAbyswrdTEP7ck6py9OIIUw6GlZgzE2cCDWU0W22WlS6xSHzRvz5Dxm
egLnBvnpR5EH7qf2MFz14wZVoe9q9wW+fLiOmK6vS2q1Jxy5V+D+9MqnMMr0frcZJ1XQuqyY4sR7
TarIeJ1SOJ48+c21e+Nm3MFWS3pc0eoDCzw2f4nB7Ae4WflbM6yK4EUEVsxLMZVx1FIaVDqtjosT
o8GFI75TgNqdLK5Z318KOKiXHWJwT1zKwlH6rNj0vsZL958MP6JKYnTmRZ0IvcH0SE+096DF9sV8
L/4QVVZqpASwG2gOF0hrVw//7nJ9jOgMYD70IftlR0TteM14RJvJerb/5qyegqnL1dTAOUgpvS8X
vPusg3bz2lo8iW+HUrqD9DY5r3aAdXAXiI1b5XxIMEG6Kyor0WWaMLY56MHu/p9OzcjzcZRAk+B6
m0OwNzfKqxTZxm8b42TeNDOeZ/r1Sfnqi9BYF7T8bzeT2QRZkZadlZRcruL/EH0t/2uR6d6C5oIO
qK7PHU0gxlcSU+l9HKw1qIB2p+0XQ+ECHbz+UCmHi99YVn5N8O6F4OF80KzubO2coLXO8p6qt1X3
6twqCpDUskklFW0zNE9QVkunLMbCFKrezVh6CRiCIvf7Qg9VLFQ4xVOI5HLUuC84XTxnic+VIzTH
owBInDH5npxXAfLZbz2C7zHbkZrAt47xWkRiYFpMm/aDOQtzn7wqLSOoCaWKakFaQcLqPACHDszX
HdsL6SJRYn1dwpUc7sfPS06DZa30KHRO3FFu5cr2SM3+nMyiYCwB82F+A8HQ+gi7onfqo8D4eyuw
0Xzp/NbDdvXM38DvE3ArJBV7dJI1NmVh4TY6hgnUO7WiPLtzQzx/ehFzBUZgqNLQ3hS4mHwAxu1C
mZSqJI2p7smxKpvaKLZTV8ehVvIA9i/2bUdXCl2PFC0ZOT6yiv1LLAAEbs4yHYiNP5Dc5NLt+jMr
H4mpqF0I1QkiKGrIO1myCZ9PwjBXIpV3BEQIrGbn9FblBGQc6rkMmEnvVk8W8c2haAR0CZVDB57Y
mMJZuBa46taLqOs0yI5TjrUqxXJ65wRQ9WnVnXbJjcYtrTLKmDC8ItagQYKCeXCv6Bpt0NQlr7pW
51QJ4yQPImw9rd1RtZ7FBiAU7YlOR3eAi6wODO8O9jDjH1ktaklIjmgrtfrtGmjZRrcsQl738WYd
W1YV95l2ZYq/iWuA0Xu5xtu/0+cLU9qFJc8Tn+sC90c/0uwP8ntVx6jJp2OCbTqYFRSAF8VmEkep
ZF6cnuMTLb0cpZhoeeM4Jf/E1u3+aVps8YM88iVia87LLMBbKUyCz8S/p1BsB6K+3a/keQfT/sal
26LmNCihK+7Mz02sxRswKkpUM6PCvP9ShgYF1Ws0HPZU2+Q0OHUEr3BL1P5Zw6a1pdtZNPOr2IVD
RA4eA9rjj2Hkbu9x2vfXDV6nf3z38YCwDeG3kcEWhPEmJZsTAIp9rLRAKyZkD+ltQuzxuYkcUJdN
nPgL7MCrZba3NElEV0HCtaa5p0KIkexYGstvJSRlVTf6/wW9ci5srtbeLUvXlNNMPmHgq48YJ3EW
GI+fxHUT4X1fkV3gX6lRJnJNNBXshnYy9IIXuXP9xt4f01ikuuGLs2gckkMvAaWKWKQon4+ucYO3
51pHmZ5DgXZZwq8/ChwZfMinTREM5t88WcDuOxOsae8ObwGffSorWk9tFCdlqaFIUVHJJsEbPau9
ub7u8T7jemIuFvQdKHyyEgCUb9FcKC94KkqfTP+9grQl7q7jvLqwnyqaX53rPFUzfRZu5hiWQZ72
sgFLaKHqFfSxiRg5oi+V112itXLJFTZUYSjv86tiyteVba0sdB6KslMrwZIt3/t4vXnXvxn3x8jX
s6fROyD6pmkOKXtEXhAxGEA9HPG4+/jWsNyh7IY7mzsD2ie1AFQ1BXRkDVJ9pWHLlPx0AdtiBkAx
wv3yHSIeeGdBwViakRMFPFGjfC7oFy/Jyt5JsbbVcEgWTXQfIrTxYGWttMriNTStvv6tOICKftPZ
4S3LK0ytxx0ZqvrKuefku3q+3+UbS/nNHHgJjB+ear45Cwnxw4jVB15CI6B8Y9XOQgX+Z/dbzF8D
XHkkHMZuuXYk3vVP0fx39AxN94Zphh8UN9JR/hyPrIimbOSzn9nBu8EB1slsYbCANILc9IURsi86
rkFbVnaWnzUdTGwvZPVPSn4vHkhrSELWf2YWt/iUG7tzh94M9J6NrYtfsblwxz05o0umhn2vVOy7
giC4sC4sf9Ds4v8/yvVR4Dlzrdb7BnWsIyqSz3SVoE2J+DncjUlOTJdks+swOxV1Acps4/tuYbUB
5X+83piQHikkvsIXXpejXGuiFQVdCHPLXubz9QBxpngN8LFBEhetVm3tejepOaRg23nuJtD04EpN
LMa+Vxzk4NPxXtU1TGCwAvtj9K8dAsmrlRrqvkatvJHQRIgRkTV20L6gdXM0k0vbRXObaOIn7AJm
2tl8ouwBQ5cX5vuANMqXOEvUKERc2bkqfAGlR4ogG6Ry3ftlZD1SokKRzalRWqSXR2i5jnPZJaI0
Bg4vQrMaAvz2UM/B6ZrJVLdB8ZSB5GaIZT9MrOaaSI2TlobYp7G4kCYiCmI3+Q/3juA9Wpxtd6p3
c3WT9f26KZrDmdftqQmz5e+5CuKjrXId//bHtCCg4fOn9oDp0/6pK35/S07KcXSdCeW84X0iprYh
Osg6EaXubbxS3ggotc+snYD1+zIhhbwnJmb94O9aaQRH5BWpbbB0Cgent1mb8AnbYqBuFaZ/oA3Y
M8BZ1Jdbeuy2sjuswPHafWmVaFTA0o+ou+mL1DRzvHGZERoXT2rT4KcZ3j1Jr6/71ovrtTjqr2rJ
P5ajqrGuYQM7SGTRR+Exz5v0if595nJRRILL2tRrOK+31nx40YcmfDxcP5Uc6g43gamtH34QP6ZF
lXPT/c3YzwMRFgp8WpT2x35A2COrzF/eXhLVyAoTPZveUODXYCY+ZCnkRQ+LxhTwcsSQAVC8r7lj
dGILlr5SQoiFyHakLsxMUMkLqKq2hvWL1Ue9gt6F2wQWWLNrcuInZGjeuYVUZxofPJYnX5OrUSQb
4eXqKIxaFv9pNOlGKi0Z2fMjSSjh4bxSKxRG8/A2v1XLB3LVDw0oySa8joeZeijbU0c7GuTK0P2F
D6bq7/NU/Am0Mgyo0GjbzKinHj6VvMoGMu1k3k9xwCVJMCtqr5GUqdQigzEyzvn5Wmmevj2cDM7g
n7BOtL175qA5HnDnlCY7zYKL5WMB+uMTc3nhsBW9/f8TXykxL+bJ6FOSi7oL4lqJAI4c/GnDtMNI
M7WyoXqctm7W3CJiO/MZ3rjsneqwQ1vYnl0xlhza7UyuIXGudip17cM4MTA4ujk6z52QkHcE1z12
YwISfvTx4aKNcNTJPBq58xmv6LJfGduiYrvNS6faIWVCohqrFa+FC9DrvVhzAF6DAmYgSbe3xX0K
ijdJVYXmUJVuED7XT3iurqj//wAG/aZD2/TJGD2A+X3GPtpW8xSx683w9QZNsu9LoTR4wLTGewGv
UzLiHIzKwfrbL9ZMbvRChKirbdeADzFpifYMlAkTfetDhVKiydhnbblYBmEV5x2utHgAADV/86UY
mZ+36N0hMGSyVlJbCfPLl+hh3AYhprZofXhUkNgVvnvRd9GfSTTcssGmJ43XxynZv75BsfU+gMak
hC3ARkf9LRBCwUmG6ybvLZZCUV3bAGKMdhZ9pah1AK+I4VBhlOLAljzSHt5frxo04y0Oti7R50q9
dmhQO/XoZZeJ0kcyq22Vx5TXHtVoNwidZwz1aSTzkS3SfzZmXTLkBZhJsvKoG4u7nlgXxITU/RJB
mhc+7iUiei5qLgBehA7pd5JPCJ4f0798rElJIyIWcUgBH2D13OLgO8ELRQqaRsI1OTC1eebffxK+
W5d3TojzOxvTwpPWgH3h6cxhXW3DM/fD89IbnHOMz/cJ0/seNVPFeeC58YinLNcoGz9OqdOy/W/d
WS2lTl3C89hGSb0/Qzqwo0lLLiKfwmqHRGTIhxLjXjOp7ibcAemjGR5tZVL1gg11bH7Qr+KtcrHL
GqYWuonV2LlgUFgKsDYZw7x3W380wI4rL5vZqO/pBt3oye8vsaZHk0j4wrSkLv1A3/1n9ogGfNIT
5g7eNuyj/iA5Lqk3Gw4lU/0S6ZFvoHE1NpUynAtv7lpVt2ckkEycRgxTFPXWjT6PoM25uth+cHZ7
HxM+1VrfBu93McCjyV41SRZP+q/idpYQRLeZQumLXlWRS7o8IMtrxRv4WVFqJXKbffds1BWD5A/I
aoB0l/ZYWLQDtfDIb4SzJbRDNFqBl5+JLeE5PEi1f2jwKNu0/8d+YQsfaacTXt54N8Z8HJU0BvpX
qzbYvUjedB309gWp3Dmd+XrAHE0YoZgeaKJTgGmboCA/p7AaiwZzKNpPG5IZ55RQY/Xl3afFC3mo
u6CPM9pzhDA+M6KZWXlTaelgpHeK9ZWj3XvWSsRU2janIFFPyrQzcUaek0rwHD2P3jPeiHEcr8Oi
52TlEbgHRu4cqGl8H1pkR6yM0yuhMj7akCs3qBxj6207Spl3XGJgaA7U5HvTnHs2u/hmlQTNsxhM
KdDvrwKbm8NEfPOPC4er4pt4wo0Bkh5H3qiodt/4GlV7S81HFHZkf5187oQ8OvprSc2QvlFQ9ueU
S4BJIHG+9oXy2suNFUBzGMpTyqb++y3Iq1EOOv/Mi3gtPYRr/FLC/lJEussHo5l+L8SkBs5qYpHj
Zg4ys27iopB7tmSymyOpm9I2/VC2LVQr7LWsWwTcN/WmanElFglUAiJmNZacU++XovwiVbXQolM6
BzGh0tADyPaYQyZKm9PGSlJGwAHmSTcI++yiUTpBzWrjMqSaIk6wSVGA9YySybS3uxVPvRnjr7Wo
6DV2guMAIDnkjIWZ7hzMfiZXrhxQMbyG1pHkp4A2c3U+aLvsGbJfDHELtrlHywgv35R3XAoGqxd+
hWuRObP8reci5vwGtEKZ1LDGo0jUxUj8ua11Vvr5xFUsvuCc4QaLhkCXMuwNL1FYkH8nrFXBu2qi
0087PeddGnX8FL1oNoYus4ci762sLrSVRoL+6sOb9M6nwBt8eWmMO4HFnb3CQ1A9RwLs1j1nN1hy
gG8jOrXz93f0u5SxKvL+cAcPbVHLBXDPc0n4c52AqJ9SwdVVvqYHWwOS4ihGcBoYQPAPG5EaaNS5
vqPvXIkRDaLjqT8HP3QU4bbTYHQDIYP4vY8u3p2zxtHWSvUH0tlz1cDR1fRNbu2Ns4sPD8vnsFHV
Jm2HxcRepTGe9cijit8Kex2RnOPPf+tlS/60RXYwFXI2waNgDbRro55aCt1P6byl5a4Jmu3OrwWR
q70PnrUO7nt5AkcN6kls8xrt1Jcs/Hfp7wkd4uNwcFu2+UKh6Mk4V0AhcV8eC54NKaZxe4+2QRfy
FTmKwyNjurQNmfGmIdOFusBXd+EDSaVvOXVt7A920AiuvWvbUXTAFgrXwD2Ve7pI+IgVyBI5P2Vu
TdkWkwXpuZhwQfcHwDmO/IusG4D6KhM0gH+OWM3AC2XazfeJ89oX2N6DunToUHiYcjQltaGgpfEO
MdPpPilSonLz9oggxi8BYnhj+053BB4cRYbs2eYj3wBvq1FDwv17ngdZoA59bWX8Sny0032SAUhb
ZvJLeItexJDXKbZl9L6+a7JXdBAjJQphoA0mPM2XGF4OXyJ7VqZ1iNrPg5Yc705rgZsAY65QVWI0
eX/4CgPotX0n7c+8cl8FjwXrggb4yjKWEvSCbOV89rvi4uMCFTbj81H2/EEGk9yw3e28Dib22XtY
wH2iZa2Dz0NeihUxbEqpOH4GSrOHtkezeSgACvFbn1PnfufrDyDJrMcpPOq++P2MtKoib6Iz9oF9
I4GgB3d65pq+XNW6mx+2t4wxysBHKXBVs4jW5qCXdDyYDb+RUjGU3ZNaHVV/h2kkCmpdOM1NodVd
dYbQimQIxS6k6+o/YI2OX46tEpzieIy2FG24J8iE2YHyo/C2IiMQQCbGwnsfABf2F2VGurXjgVAN
EJxuDAwDy9Cj3j4b2w1aVAD5YnJdXV4jIFmsDVg5Dje1IoX3lw0dVul+F9ZD+z9TrcWsBCmYHToN
mfhqXzL+Sxe6tb4u21ZIQOExXoix+kgQW2rnaMAL2hGGNWlNGpRvA3rYF0z93h+Q2SbiXiVg9Ll8
b9Y6RI+83Uf5FlPykkb1sLic7H8kV+UjKpqOCzeB7ogHiRcdzzqzuuSJecy+HtZx685NT4tWSF3F
TpzIBv8pKJryEzQWIMczjqhFxo1k/zBsqGU/y8ixhqDw/3QKoev1MNgOyeY1byxkDpPYDe0pl6mN
FW8vBSdoepBB0Batwm41+dJrw4W0Eao6LBVaeazUwfl+NVLLDTLpxhwjoNKQbaKCQ3jpticpYYKJ
Jq2fjC+f+WfOUPi3OMZFso+cxQvosvJ1kmSJDW3w6i9UBzJ6fHIyVMp0smjcf7wAIqK2Nu/Xsfhg
H+QVPVaOviIn63o78fZ7H810y41G3EryEaOZ/x8xmp5TGcoNwoCv1UdoJNNrqGzi9J9BrfdNpkuB
5+1VP7Bfd4ynA/T5aSW/oFkje1a/E3KSqAajqris52Iq3xhsxpgXGcfU9QhQH31KfqBdrrLD626s
JO0iv912TNXL061cc36dwcAjpu6npmYn5PxfT7fQURlLVZrWJpoBjQNWdtHFjvHuM+mlVpI/5S9X
Z/woTFJ/g18ul5dYb7KGfR0T06Vumf57lFlhwIEj1KsCvUbGhIdBtgsdM53XL9AgE7oY6ztCOluf
WkeeWgB+yokpDjuBRz4uhStzQ2XdM3gdhqHHKo1/JXnJPk8YCzFyVTsvgE8T8ovCn058X+fabzTr
Lxdqs0YVrGFzEFkS2IQc43M61iyt77PqQ6p9NaUiieHTm25c8Na5Do314weZSLxcLRoyX4c/v1os
T4v2bM7/JFtv7mlwcsxPTkCfC5E1a2shmsRWI7Pzm8trWJou6Wbyh9Cr/TGIFm3DvqUmyD3I/dXe
W5yyHFvghF2tXDZkxrKEcTKf3Ro9c1WsPxtg89dDrMVu0rcSeHhw/F04p5LxDejm5d3SSYd0Ssev
sGonP/55e/1DsH/HMWuZr0wfRc3yH8piAFBNbadtytUWd21S8SfSoOx7xq5OKRbp+SVIS9AmyNGf
tXsr9AMLkVfs0Xck+UuQcdZTnXHGo9v+a2Wh9Oym8uKDbsS4OWRhNWlSvw5LVJyg7w4WIJXHq9LI
POZ6wXFkvoGmcRxpq1GlYmBpBe1Eumi/Ng6yYwdTfH1zXB2LUOMFmCSXSZkRcnt0lHTVBvVako85
+PVSa0/J03kVaUJDH+j4Tqp31FDn8ir0sh8Cphybyn3OfGBxv7sXfJyK8AMfUWB3j5/CvLbKuIB+
xKgXROrGhQgwSnUTKMFFwfUrUWseLfYdNq9hQwFeo/iu+8gY8LmKi+/Po7/NzGWgHw/kwtbftrxA
YFQ8yGhMrgcN+gPb0bXMnogrWqqnSD6SYSR508QlJNNISZHN5Melesd5TM+LsqWt+H6+5fZEIFCi
aDGMcIhrcG1INn6+zsU2ePZYpW9sBWfVfLT8MikNZ+vVjfEc8uZfFmy/psIftNtbp77lA+iQEyuO
kdZfrNEgYO2OxfJD8fNOlisRV2AV6Jx9cYzGrOq5a27Zveh4nG3xc+wAV8G+XWpNr9RR+J0eDC9H
QrXNOqVPa+Mwgo0gPZiTYkdREZyFgE+/qyIsy/gW+CEV7KYmEAvb/CTIUDwwG6RYF0noOqQg/kOT
2M8cQ5U+o1tjWn61ZRZ3SYOfgrz9c+BFE1Ohnd5jvNuDhkbFG8f03fxjz5XIhySFhMJoyIiV5wVc
5NYwLNqjio+EDMxQdgvSluYGoOMO0Ew9kboZdK12eY94tGl7Pw4Ib/QQS+EtbDi/8Za/m26ZpRtP
k+lBACebE3K2/uXV8nnmFmoYh53bCL1kXQBCzZ4D6irxc6gtLS5pKqf+q3KJAmUXtJfjkjSvLHAj
Dq6NqFP/ZtKLDNEMfHs0Ak4S7ywIDGu6+kx8lKMLggQ9vPJxXoAd6ta97p+gI2DAMn2xnyPuhDyU
WhlGo81eLt42RTiuTHKnojgpaFc5hl1LcbbTTt1jGs4Dk3sWmYNVpOOa+t0FV+Ueuq1Ay6k8Vpk2
uP1hBVGlwPPW/DvCkihReh1lkV6f+7KFFpRPfIzFji4rs2NOzuryqFHAFtr/eCrW2jM4CXclg3z8
pH6rrm5qtB6IrHlFLM1XUsx60TTLwkfqaBdd6sa814OBqjU6NxebJktu1La9pEPfeww7YEj2lNru
HAbe72J7pfe/XaADQlel+FOjpGQExR5I8+7cxJCHrwNMrLX0A5tJpgZ809uK0SvBk3QQvcMlkUW4
Uge+Yfh7LW3mE0okOaRIQ/WiH3CkrX3j91cKPlLbM3A9aXEq/YQikUOa8+Pid/fU/EOFXQD7tXgR
tWpIOOvoiEvOCiA963dEaUn2ogP3Y+sGs1It1WkIjv0VpeF/P2PDUbJR/g92sIzyX6YPebvgEkAw
FzKthu7PV3h3dLvjWs39iPBWcvG9wPerDCnwAz3Wn2oXyT12180/NaYR4Ue3Cju0RsB5dYtmTuIH
aJqe4fTEX6tYMDG9rxk/jmWjAhI0Vkv8hsr6l9UHbOqZUeP6x3W4sHywdR56JGF9/1bw4lfrpxqS
xMt9R0JdVKI8XGRUwWNH6SLX97cesuhEqwmn8wR/k6UGpiYbbGcOmw9Z2cxM+HZPpkcJ3jDCGPKy
HQaymSsu5fWzIiWVIC3+iUxrgeSOjZRPPptvwhPHWKcR0H7wMbySnmXxGSxyy55SgzlJ7mT3wYxm
QbJTJ196DPjDL7hkZMU7/qeoQ9Fz8p7ixx3bekGXMkVfefOovAH/fTpiGVT69Dgrpk0Vis+WJg6o
ExApnrY3DUt+RBbA/yoz1Zi1rIJyIxyo64VI7b1H+vUj3Q9yJ+LZsN9urEup4WSR1HpCe4YVVlen
MjoURl+/PQNhUjMgD6OArApfYcu8U+RVd3RJ8w2NLYGw2XObiXckvZEgutt4EN0AsGkffZ1VXVax
6YJk3pxA8sWErWAKyT0XG47lP2G7c5UOsWz9Jwsc0EsUVgGL8iXaDyE3jnpACZFGVqGS9O9FT3Tl
C5Z5cH1Sbbjx3I1P3RAJkzvhzwt8RwsVJb3hwj0rtlW7eRdSoN5UlQ5dfrgz0mOBvDhsKYzfWqjV
oNnUe4hDXeri4gFXRu03qeeGWjhOKORLsBTtwkEMgoGJUfwc/vvT5njx44GpujLuzK5pf2xtYsi7
bV3nHU3HkiwEWGqpBy/WeAWMV5HNQUFXJEtuwCKfxVpHQ6CMCfbRESMtXhDhzB9BktMJUeIrJPcI
FVUQbIAUfLZuJmF5gWrN6dx5aqQ9lWa+vXMJEiFQAz4ISAxMAO2CBK92p9OMkBmK1D1ySOy1GnCh
bQO/LwffMnno1nnB2Iz0Ku598AFCh6fzP04s+E5yj/AaQpOSOfUdx+wQx7+MSAVTUqoMdmUFN6FW
9mYKcCwpNaRYPspLfpZMC3wYZ51Kqua6wRDt5Cufo5wITJ2QqpS+bU84zQfjwGvmHpziqSh3zSt4
9qpBLR/oZhu6T584WdT1umwRaRgOs0pKNDp2pblPYreSaw0U9l/DCOeGPLG5GNSP6ZdMB2kgclkv
jIOdggLRmaE0ueFnUWG61sLkGD/jV4B/8zkfk7QI3Gqdv6+50nmKRumW4fgCz/g50HTBM7JWtbNP
0yyiXI+AHZYMB7idGRc2pI0/doaMh4W3gmstjaGfyJFwKdvvVhM9LToRj866SRFV2bbnrpyP8Yq1
0UMSCNcrn0qT8VZCmD9Pp2TtLGv6M+UkViaeCjLWBua+XA2fS3vEKsD+UmrqmH6HFacvyi6UNF0K
xLKVewQXzliCPc52j/EIDnH9aIZlz6xmczP4iIyI2+btJ0MUQvGHBxjqFqC495QIHMOCDenN/Iel
Ewv22zswEZxXnIaFuGWxtIenvomJ3RGlDJ8Z6g55bl4VDKZEVXBKr+7VTupo/cuJTGeCVkDWCp/p
7DABADP4uzPEEI4j95tAIKIKAMllHXbyca78mDnPEIbzKxpKx/iXUW9BfA+swax1uik6tR4lSxEU
g+KuxPSlgsJks8K+lyizstcbRJKwLUX6BtNqaSJjmQaymqRNi0O9Emju+bIfpdJPgDmyfho8vbpW
M1p5zsJnvumz6BpabOJByJf/QDgGfOyJ2pgvQsJkKnVJDdfGvLx/t7m/ckhoTV7ZSHbjAHBTRYi8
zDCjo/sRYuo7s1xYZ7M/gQCvH7ocW7kU/wGljaOiRiZ0lR/CiHmUQPRqewdHN0YyhtB9OBrqjaaE
vEqGaDChzKhywtiPHq5CpSRze6F2pan4VbMEkNsHmvWOerWYtFznYBrvsm1vyjnqmtf/hsd0GWy8
Hhq8eFkUfB0qXJuIbqBOtBtpvBv5aXbeNDyEkUsZQWLnazGhnjl+1litcN5oaeRN5EHIyTIWQPsl
KMgwgTwN7jhqs4UNt4UAZcsC7ws7y637ACejJcaneG5c9p/c0mrHnH9OmeV5lQL+ylynECjZh2nq
I61xq7B/uXeanABBdVk3zbm5U0qIKesl1m61r9dbtG3WVTx4Mn4c6TQV1L7HKIGeEM7cIt+TbMV+
XlaSCYB3nN9DSQlDfmPis6xgqEowVN/ISG6oNlM7R/2TlXvya4ytPMs51xwzmnQijyc8rDEsHxIX
G7AR5mNatyG5bVH3qc0pVSlpRMkOBaeYdKJX0ERxIFyKQm8VtqSMvyAB5Ew8ieFYyIGuWqOEbL57
U3QMTmP1STPRbQCb0l1xOrOWp/aBo/MCMWgiMoG1fNKm8l87sEI7UGyv5YQCAWY4bAQb9TyPNdku
GFx88A7K2cEknLPt/CH9YADY0DZyq0xkMfSd03l95S/8aiQQfTuH+uGW/E7ayduF4V6mdL2aMi61
OekYt7eqOnWcLKVgLwBCHB3SvZJb9C5Dj7adXa6qsCLmKdv9sVomXFfVq4e0dsXs1z8ah886KfoX
2LCWDfV9N+SOldMiwzTWo0J7kGUh8mnkrF/qONKPLDvBcYOxWwMwfgQxOUAHwFhGIMfYRh9b3loQ
w0rG0ADG5ayEWg1mJFiOw7aRplb0ECAvpbsxdGAtX2RlUuOa74ysoRLPnh+pNrXPCelELJdLnmmy
ld86nUKfetuu/dGNTYf53nD3xbGDQsEnzDz8Rb6VA9jasIpy3Btn7x8zfzWnmmrNtJ9UdGH/X2p0
xj/adT/7J9dmb28s5xPuWGLBgK5pyMhgFr0E4vBFIce6xMJPL2wuJVHFCP8wV2V+5TGxQtAbzZds
doiiaSg00CPWA5Cp/M1/vRJSqmDCv3aIKK1j7++m2E1TRv4Wv0+YfB5RAcAYXlFMOvrfKAVUHG9W
ny71vhUomm9BUiQnY9xTIa8c4AhnXZ1lEUZWYBpZUdMRnhQzlRIC0QWjNpkj+BOBWXDkX3OOShU0
xXZk5tCzNeGa9h9N/T8vvD5eEP/GhjU4FFi2Thjg8LLtyFNqaznETnFp/A5hnEADz1OO7xImCIyl
6gdBgJGoZ7+DDvKcUnBRP5SpYIFPYiRbIMx7YbPp93+m2PEhuPfho9dpQPTJdgD6YqIfRm64esFd
u6+FFRysBT+u8OZlESQUMtr6ouEsAaOzwFUNNz2mjwUF1/c5kq7ZA31kj1nvZPOBBF4yREmWvTI+
p1nakL6KxuCaBIiqPcrQ3Qe7PRJ8+3kUVRUEx6cxjfIpEF1s3jAYnHMB+5Tuf4Ng5/2jCPpnSBW+
tvTT8NgpZ7VbWB8V4W33UymtK/u08AP/EW2IpWH/q3t/tqMCvZStjwgVi6EPHRBRiEb4VGsKftWA
7FhtN+8ieLZPJZHwl88hBJahzCjh9iMBJBQONyWvW7vDP+5HaDltaNWwwpcwOakKnd+tLmXiTV7L
1gXhLxmNjGOzZvNMVrj3eLhrgJHmBmwqAFh6hqxJwDn/Ri7uIRadgs82eHoLFTkYy81hKZLRDNGU
E44TRpNBmTeYNNfDgfIEyV4TSU53EpCnPLAP9x8jNuQgcGga8J54z/fCOlrn/6vJ/IDTAxv6Evru
SiBkOGA5Vl7OCvXFnmsxY5AEZDMdP9uIVR+Qf7cDUJZOlpbTySm81mC5yTGl0qLlxEAYPl5bIFD5
/cPM2vBIr529l8OzftrXRLRliHPOPFeTf5nAzBx4gSF8TlH/sZSVZSLxOojeChREUlTZFiwMi1nJ
xx5s2sinPS+zR2dqiK/TsGg5hWTy0EdUcdkBgo7n8SN8RNdFNHVM9dY5aAMSQnN36i44GRi9OsoS
Tphb4SF+Aof+Q+oNbfuvmJ8/XOUakza+OgCxM5i8nu7AU/+WpHZhhwGnhSqCFANuET6WyNxLWidb
aZav4yi/VL5EAQB8GDfrbeeP6mpu0Em3dPb2a2IwMirWRZfG6ryypJ4DWCQeR/gOqXDwfcnEgdN5
D/Rnb24SiBSDYVGiCGYVNd3I1KYxy2nP0kgCph8tRH5V+SLB16lr4XbmG2GhRTXpMemw0xlcIX+6
bQNfdLIuWeh0gT1FQV5bqGFB6Vg5vPdlN2h+QcHKnrJIinAqLqZyPD+puKuOWYQROyDJkpiAib6U
Mg/wUo5mQF88VUijLddpCrXX6qHs4/T9Dtdce1ZnomdEgilpXfYtvKYamPWWqJzXBlpuxAysSruK
yNNOnnOl5cEub1BJSY9AYosdhztK2vt3cC9pOsV5u9rHfVLyAIBmU/U5DaB+/OBgqeyobRNq1GlP
mevn4TB9PYd56Nr6bDjIumH1C/qTsKwyXsmXsDAPImcLbylFanle04vkYw7P9e41D3IAIJuoKfF1
ev1f7PqCZXuHGB8PrRMHXIwMZxxZWxpng4ebTA4BJhee3ZAuceQl/l4k0/5bb66hjk5ltxNdWXou
QSYJC3TRnEUffhIX2rvufYbX+s/N45lbDIl/9tbiKe2MoOpDstaTN0wTWzpvSF5IKtDBdn/Obaw4
7r85cAIoc2GsrNHegT/TZFlHCJGK+3KuEqOHNIikyzFSLVAbT7E/JQqB2QruzhM+Xbk3Vd8hB+px
2bi1rWn2ismmXHCxVKCk+J1G96HLbPw8QDdP72R7yffy984PK9861mWuDH+RQq55hEmshwvJva0s
dkpJGzb1eTCkI01/6NsNSxzGFWcb9EDc0gcQ7NcRX2w4bhrjIhkoG2HkcCoEaxK5+zSO2LKnRdNv
yCC8727Fu8iBG9ThHb6ElP/IgiWmLi6ZqXQvZoiYT/KeEz5YcDlsflPuNJtsTjXArJqowtEC7ZB9
vXcjqUNyCreVv27sRyPbbXdi18XYvW3WHzZ+LkFbqQ1Hky+bZ7zlQVwm/s6WwEvwuQ3lkGTW4iWv
E/LGyOGDlZS8MMOtzfOw0OW89SV+Qs2oQAY6Vk68C6rk+fQMb+dvtX6Tfi10aE890p0KDljf5vDs
8ebjT5ykVEn38N/jU1qQNMn05VX7iNpQyKlWsFK1v5CI0/VzWfu5AWMbhIooUorb2IGwjDZRuQrp
rPQJQKuRUU9jUtVJpAxKN8DevvtLU65fu+cE7J7/8cJ4UM6cOtorlDcUrAFe/0kiA4vMY/KUzXaG
IwGjmHiKUqCx3VVy38XfPn8jq+a0A3bNrs0RANkBw95Rs9tR+SotLU8tKOQysZG1qF+4MYaovwsZ
+1FyL6B3kvNQ1bSHJDusiMLVcqIluLkZJkBQYvzs75mLCgs506P4S9leY5QWZ5OmZbuJN0ki4779
nWz9OaYdN+CnyAAMV7QC/WjaMB8JUnCDw/kXxtLRTYkzbYWdsh8wPtt9SSJzJt0eteEb1JdkIY6o
n6K2pJp6rmh2XTA+IhD+b8DF0KfhJATUT6aEBJOuHZlVMZiOzN/LYit2XIhI3KDx+K5664xlzR02
gYBypnQKJDqOjS7Pjd/PWIR5l00/TuPVAl5qIkEi/ZDqHzzY3sg8JAyf4XnExzKL8TsseCq/3c3Q
ZOlmO5UQFiRX3zirIDzKl9bPgXct0FXe6k/tMTBSEy2xQmoHXCKnYLep0PVwzUiu+7LFzebz2Us+
w4S216kywBITtfmldvuFXESXZD+lndtTM65MSKNA8pt72VvlSL0rzNJ8SCqTgJw4O6MG0RtZAZMN
a5SSHCtqQjs778FULOL8jQL52LMB+2V3nU++sN1T7M4JX1SV2g3oBGAfC4eck7iHT3f3avHbl1WD
mpdSt4FA6Yyy+/a2oFKvZfd3wK307Enf/O9Y+4AMa6bpZJ+aZ1MSUNJyFDTEkmH4VtUMgIr8k2XB
uZ4y54Q1A9h96Yh1bKyiX9NCmRhAEy23sMcHyrEAjxwVcoyykuFca661cZn7c3nNkSRiLHLEYMqj
FqbatpJ/HytqfLaNGabdhLZ4UCTRAN6df9mbuwjLFJQhYM0+ehAm9xyz31kZ8YIu0Ps+HjA5VqpP
4cunEfkL7ZnGQcjcSHVXnR8qaSdaWJs39qal1vUa/anpKeh5wkeM8tzb3sjQKGhnsfOu3Be0p+B3
dEFvolRZw2EfQWvtYerkcBljfDsKTqxRW2QRY+AH3SxWQEypZl2nxmBpPtON44cBEitern2UYEJH
F4ZbN/AKVylm/Igp1x1AQ5rnvhNs9xdGGNDVubYcmGus+FDvxFBGG+ke0wFrAEbFZCBPDsX33YXz
ohC82qk/Q2zwZsqIbvcT4B4abiFNWpYTfbcfnn3j/sBnIHN7inM6ZyXHF1gP+cZKoFUM9aYnJjNa
gIYrK5HC5Yj42NM8nNBATdlWjsp4UBH7B9sAl0mqepqgzS8ZLiYAyf5z0X8hNAcpxsRNhKx78XJv
mgi2LooQAoX8O0/weS7Bh2HrkDq/ASaq1pepyLhQtO7r00mJdph1/MpxwDEI+xNETkyFUntxz1Kc
7dGvbwYFPoPCBhNgyqBpLghJmT7uIYsbMjNYm86+XO8hDh4/Klku4EHBN9I+fGgRugELNhILmDpg
mN8p9wOIU907+Mr9zW5jmvAtFDYAzpLx3kP29v3PBspRX7T/BmiNNlxxDvvEoef8Toc9vSE5sPBz
BEe6yY1ItqwRqryo85hKdS+qQ4uDaxjo80LTTHouEIPcJVZmsQhlUs6v+KyrnDjJY9fB1VP1eQ9e
j8LGFh0NRbJJ1lSLEhTau/cL3WHJ41e3TGEmanC73Fkss1TqDaVONwX0jOEP+2vr6aaQL86pDHw8
Tf/RH4nHhTauqjRPzHWenYAmwoxn4HhB5CKjk+wY7qkyc0og8jyC5+lljR8OyUsyBLMSeE+e+ShB
Sgj840uZDVHmzkgUfnKftiGrnjfpP82WXU5b6+WouJDe/wOrpUFvr8xCxHPW3JsOvkojd5Fr6ijp
21Rvagh5e5knMzngdnH9OAR1bvKIYq0sEprjIuNAxfB1ev1DFRR1CKrfW29BYhU2aDbCeC9FZH7A
jGe3Iw4CP32dFbyD7Sxteg4oAzS1yK4O5puJQ4bAoXmRiqE+xXtdgZTrH0c3c8CJLMwYZ10HRWDZ
VFagrUxri9jMVxX4NKFsh2Aa+4OdAMxTNQuuSOXgeSwCBy91zTJNU6GwGpCunwb4P2UTH3w4nS61
fGRozowwkkarT7B6yfpPojz4WswiD9hbIEnYqNvQXovp69dUSD1K9BY347Y3hl24t06HcyXV5O47
Sg8VdwSi1tDN7Xa1lQJnmlMjrr3AQ90wJ1ZW75dpx0JyGdiyObsWvwJEZ0tBdF2Ucxo3+HkbYmx3
Jx6iEwolp76dAb54eXwBKIPCvg+kIMzNNw2jON/zQlMlAOfWs0IOkD8aWRV5YJz/b5X6dfdvI1Gc
l4pyUhgvZ8JDL+/ZJ+7+2L1nBcEuLBsOwmLKRhV/BQ+kBgrfH90XiCVQfKnaWY2SQLp1zXDwsd6N
rQ+SMAlBJzw3bjL+Tr660D0CdQO9YCiPS+rWDeAVX+Dgf7F4wgqhJcUGc07Es9H3s7KtaXVbgyQr
+kaRQunfsamsQMoyJfJgkgqKPMtht+YRcXALz9yMwiBjP2yoUAtqDataOk116Sa3UaTNFAwVsjzh
rFPjqPy1w5ttZ7rtHo1ALouRbFEhBuNq3HecAm2fYrpf6AtGLZjhCpJP8D4w9mWgY7RTN8M5z0MF
P0VpdgCGYByHE9jKH9GMBT+Dbc/yQk0PY9si5/wQMYJDNohfVmZB9jEpLmRRbnek+ZqzpZUlMEGJ
CJOylUJn14t3AYIVZ31rVH11anEBxsdnRApGMjnf4WaEog63eIXBxJC0/hRX0Yks3824ORXAaoW7
Hahe/9el27WqEMI90ptu5+XdbsniQsBR7ffplscEBEN0pf+Gj7Uueuj5h+bqZCgCFp/WucU3M8lt
ivoxiwZ82V3Hcy/IzdY8nYiAiyOzajm/GRCF4bGVV4gDeFtTDWhy22OgmK0Gnh+bRQZTibpCa+uR
Cm4+V6ZOvGsyazZiqZnPdk+PX7K/if3E1kBMlseYYWZfTNfvXS5ZgSIYOD5+nAkVpMDnOXZcAHqV
uonubSwy6/inBnWdVT6Kt0uEDtA7OeL4bZuqyiuYSHB/u5MXqymk1WdxobAyHC1YViWSRIxuL9k9
/RZZ/BAOtjyWzCJPQ5LrNgVoxmJyyW26t+JArleTZNL5hD2WcSJ1d9RVqWTbo5CMVHPe0fV+ryYW
9ZBmNT5HSCqvYhp41oTZuM/y+sPn25r6Ll9pM29NHeZWneZ4xchGQL6Fcv7fly7uVHgd2OQ1Exx3
wcUi8fesvQRhKZwYCxLDDjcuW/TWPaL1y+3UoE/GZ518MqRioBC0m5JicuDEYOGhVhISEDMp7jCm
nUD0wPgi2Fh5OdHbKHREhLZ3XDnOy1qQGReaBGwhZ7WANxS8kn/f0kXDlbLhcKxaGYQcgnuecxrP
1B0mEud0EJOTuJ1L5bOUvbODzOA5aqueAUjTWlvIEYBTqTIqEvh9pzNWijvj4lHNUni7l+mqxoLZ
+3zuwf7b2jrOlP9hUylndkwEuV17z+0Gqe0WBPvo7JKd30mmxFyNnIQcY3GIyqIrwSRUEi5I6Ewy
GajX9dhfLygD/XOrPWciZh/dgtRT6TIxNh5V1sDDk/yCfbhhZgh/PEbUovAnBzkv4wwAA6V7K//o
wC0FRUmfimI5WUC7b7zjneCJNp59bvlKAvE1CCopxEe6ZhZdNo9maDLRahSal4SksLF3w90A5Zmr
YhDLyxcywpYWXh3FkRq4wcDvZVaLSkGXM4lKQyqVVgKOIhdy57MY02QbQx8LylJ64g46NWkslmzF
hcL5/5Isc1qNbSu8YjZYJUtmcfuuXQODficdon8B5H1XabHgEP0DgGfYMEdKOTkgGBEkn0Tzd/7U
Pj3OnDni8h/qHc61n40R5iqbb2NZkNmjvfv9ljamyhVTONJQAbG/me3T3S9xXjSyanmxzGM+LoFL
CAOT5a1rd9f8kpr66gX93j8SLuKGc2P0WunmilKGB0tafpwG8sqbivy9S+MODLgstbSAaXrB73aw
k8yWbjnKC/+zeJYfaWzPz8s3ieGXAR/WsfVmGI20ZS3jy/x9HZZMI2okiYg4iN4Imidkb/v5PCYH
uhBb0AY4JUJhgTOQB3UBZpd75V1mZZ08Kc8O7Z07T6ggj9/bAjtWZIedHraOMw15DFAvzn8wcfas
Cc4oGG+fY0vETHqhXt1/Ge0F0/L/kYGzJQWjHE0T3qWtR0Qv/WdXOFJxip6BnO7npcsZ3Uza+t1T
Au8TL66FW4UH9lKUWgdfLVWKBJpDkC49yF0nsCnfYlp7KwK4iXs5h64znzaSa+o8HHM1e/gQRdvM
axkMp2WZPT/GOkBDm08hC93XI882d7tussHedYOsi4fL4cRPR1Sdj5yQ32lxpHkqGqfRYzcX8YOb
f+FOYQuAlpclRpoxGrB5Pp5cBqCsYzVOqaATbfNvf1eOXhputqdPSymxoUA6UduwNUb8Z27eK+FY
/8ZOTQWMtGmVtciFJep7bcXeZ6qrxu7NmahT0g3Pyfbu1HkcS78I2NH6jwtwUyof9HTOBPPIEZS/
p1mIOLQyXUHTO2vOhw7yu4GQRfDbpKzFY9eZkh2ZEXHINFJnNaBprdVYuZEE0X5mm2UIQLeWwcLF
KwNytcFeJ16eDEOHtR2ILR4Qh/khNUZk/WAcWqyfmu1cyQG1+dF1U8uhup9gz14ikZxArjmQRMbX
a8nM+qB9OwXK7FzwgXKPHxxz8Vkp+7Dzo0Dulr001L+FO9gvA41E7sOvm7fvyLeDsTnf7qa5UsqE
9dKgy/Z8Xa3UquWv+rYmch2vZyBalx8siTN1kvHZtE80yW568cT3rgwMTVWD466rsJ4ho7B3Ppir
74zdEWomBwLMiKIMFTEBRSBYXtGkjEPJ4paIaqDq7i+AQa+ksJP+E64pHdkVozwlAA21kK1G2OmJ
0134dwQVmgps8red+UP4TOGm3CWkDbVqbQ9ANxOsLmhrgZ6gKsJ9ENtL7lhnFVoD3t3E1TetCboo
yckO/WG+FvlyOrzPn2qBHdYgBlzHUKTFGyttfqU7ruHaf/+D779iMtB0fpocc1vdmm/l/EtRcZwX
wUPKZUSc0Iyn/l7HZf3t9jdgBReDnZc0xAJ/Zruopw07Y6kpp7q0r4823n3XC9USkQUUuBDHbjdo
6CsYmKcrt2UF0z3boCUlJkJxJBhoPsRZK+xax467qsk2pGxCHGPkHeNspqBj36YIvrC/Do9hnE89
N4tcVev6xMtuWDBIxoRZ9gTV1uc0Xq5Lw0F6jMnbk7g7kbRwsU4YNOWv/Co2SuURBdOCmjQ4Zehj
g+eX576kgXqJQzmJiPEggaD+T3rjHreGTBT3K1+WCR4zqBn3ROtScKg/3R42Y9d2knoegX59M7C+
p0dWoci2zWwDvjxQRi0RfSlBrClqxoW44bX/KxR4B9rFekmD1mYRNyLWd3NHxNnqza1LLkmrKOSf
gVCYtoUjUzCl9eKTnuE5L3AVJBaArgWcBNQnQnu5jI/XUlQKGbYQyDpkL+9Dw+Q/V0pNoi/5zQzK
Lo3ELgG5qKrw9Cb97hE3EYQZ+TczcGsyT2jW8yYauv3PcfBIjD+YCeiUx+glqv4+qgsRUZrKdeu0
HzrTI1eGRPv14m2NHqMY4JbxEiZUlZ6gtbGhN1yK098wJH8qoolYO3HOqfsAGH7rt/398IQ45CLd
wxpNdpaF9DVwNs98DVKqONuWBFYiAblUshAmT/xRaD11kxKNU+bGFBqRlbvR1P29hYQgBwUDdagk
L/uyDWQQd24X6mxgwi94t7lPx+hA4drLPrVt8VLu41+043apFWeoDl14+1DajPNRIe5KJhCx5ct9
XfH2uQFxl7Q9clOZFYknuNQ41EpwA6OYIjpY4gv6vWUCxRMjC6o/8/bDD9JL9xSbqq92G5i/qFQa
BRDNuvsed39Ve/I6uuvJ9V5mVpXPuV8jPEPGOxRLEnfR8gKQPnnpGwrcYDf9icb9+ClpIE7sp0KD
YPwrG6TdPmbwmDDnlrjmoKJqn7K2kFqiOYy7Z9R5BPtl7i72Y1RzqSYgLOucur8dY7vG1L+gB8jE
FbtCbVqRIhj5WhApAiXnTQn2JP3DNZAM4uR2XNZuV9pYkvP6jmyKpun6PWvawC0ez3b6Lwpsoqyg
OCS5IZjvk409gcSElsj2ScFaMht7GkpdN8jHHyTZlVHxliF1Vb78jCn83IoiWOD9OmPUp6s27rUr
4dSIswIfBBfUnWjbVshDPfUBrvpbcslc8TYmixJ3LJVH+QeRRGJfIhe8qgEE8U34FGc4x8W37d+U
kUvIN1ElXjhore5teIZJ+X980VnYXf1G4qBJrE3QZ+SlDRr7nIj6Yaht77VA+hjPVxhxb1iXDKfW
m7D/jEhzsr1skzaMvusyrN4PP4mmfX8J0wwbMlj8YA8DoImM5bLh4gxmbPwVXFAThoTiBqCMqZkr
eazxheMssXZeGGiaEweqSlnWbl4gYB6QEbUo3eO7IuzBtZGD78F8uJxfGQblt78g0u+f0+aKj15L
IvIj1e3HHx3h1ITHOpjvmhxgHRDkNpbUb/FwuRcex8/Zxf+56gmuUmIbJh9azp3ETwOvqApVV8Dw
VOdDdGy3PDDmrO+s05p+J/qeY9SSKtT+uEdm3YEe21WHbiRx0FZlpBHFDDDkASlwH4D4Hc3D/KdL
fdtJ//ejWYQrkpHAeuxSBDedgurLW0xZgHFGgqORweZRghp+zh6xopcBGmwJxnikRIPnSG70AI5Q
X72RxQpqDKfSLTPnrgMYnXT/sqlI22Tt7xxUmn0+aDf3PBqV3YI3BPNp6d/0ck3Dm+GB/ePc6aVY
UjVd/GlzNAh+q5BocrDhcajh2Ko3a4m3QBJNRSyQx0K6kDchfK5xPWdtYsmV4ZGvGTYQuhGC0O8U
qW3IJduzYbv/JZ5Mgqh786HeX03GYGNN76t2jEjGYDMt3A/I2rZTow0I6qZ0zciKAkycARGQhDUX
x2tuBw4bDRfRP6EE/bVkfW1z4TqsYYC1seZegmsn6mA91kG3YvrQlaZlBuOgPGUi6MHvQopcafUM
86B7/J+TTR1SZeEMzqgy8iCJisd/MOm1ICbvn+zKYT+Pla2/TfSSOLSw29zcPB5BFxmawGIOxgRu
phOCAHCEqoypID1I1qCh5Sd9N8ek6lrah8Z+/9Y5KlirXs2gUiq0TiASoW6b2AQH53PMwdgKXlnf
NZwfLkYhfxR7ELhTZWyi533MWrW6ubQWimg7WNnDg3J9GHnNGINZmmo4hw6tnDHFLT8jamaJvScK
1BSaqF9w3gNYX0OWNSPKMiuaIvzf5/jr2tMW23u0c/XL6suT+7RPT1R+cmwCMKoodyi8kxaopECw
EUQO2fxy/mifq1gosmBzj1AWsaJXvRir6HTOBjgaVRj7AOmsNhxSOM6PPrR2x5dO+tLg0QYnJ6ig
PiubXn4O+EuI/syeYfrdApjcppHnBTqUkEYCHT9TcmrWPywHwGBghtmE+4rZDcWoT3GzXBiMLXoB
DNCNll0sF1kWEGMwwyp999RA2301iC20QLRmhdZpqaNRrfXV3ofsXcRFxWwpf8KLHt5nTlyijNRL
UaCsTmyob5aMFivbfjrxDuUf/ILhBB0jl7kj0WFq7eeCPwXgEiTtahiH6pHjdV8Jn6vvoD1TeVBw
ZhwcXTFkwDA4/F60XFSSkWwipsdaZUjbDKmHxBZEYEP9T1+aBuzIhX+ePOkQkhGnYABwIz06wY2A
qRak/5xjIFxkFnn02PtQ56wTbVSJscPjpCJWC2SGGdCclNOl7H29GmnsSCj7rbcbhQ8wX96OCCRp
YkFsJUY/a9HWPUIrJS6CvOUpq0hi6rliH/CbrK/U7lqy5tQSrqLM5wN3SCQS0ul1rqpPymlJJgsi
s2nojv63w9IV9FKX9GT2DGS4fwh0GvOvvodmJhV8dXLHu9NLq1Ke4kCAe7jsVerIgAsQQvdEzz7F
GLRHhh3L6ZQC0SRvnpbqVCce+CV8ZlQTUCuF11xVcc+0twS6rLH9IWdSASbB/+KK5sT8Jsb3bEyN
RjsSWectBhQuxSKmeZAjMkE4pBqJieghzceLfCSb50kMzwOPil78AnNwSV3zI9zLAdHROURFpfyC
2soSmFtXAN0m6/D6QbHo9nORUQVEZc+yJXLY6mF/nvgmoMHmHaALdFOMmB7ichuhAM7hYPoYnl3/
6uxc77SGQ46Ux4jJWcvrNtTjRAyDC34lfGwFK+PFnWZP1ec1ab0+bYA+J0jdGSsjJ901JQID51Tv
+u8+AkXhvziwFyIBCuOwnXfYRW6BT3jgSw7vmCKrDq90CVYfCgLbB8Y0JWMZmhYGwPcX087nIHyg
I4c06LPN9ZZxstAS1di1p9HiYHh+mrg0y+K2RPhPbdJiHPe2IZnJK/YE5cdl/sZx9mBXIZUDTP8/
hmXBsADYq0V00LgkPZNo8R9jwmPyuKVYFXSR8mzida/jY3rgQUC2+F6odAy4aZ3O4zY9y+yeDX/U
hud5ON5g8MuTk8XCbVd3A+8h0EtUbY4zQMSaOSLumlL0lyrDGPoTNJNEAsRaOF0WGPxioNZLtOXX
M0PZsk9CgaXr5HdPE3XtK2KVe0+KiGGMblADws+kZG21BnZY5PEp09bmqusEBCAoUbdDAzEZmv0e
uJ1npe6p/8SKz5m4EfqHJflqm/m7iUzBk9ctrDtaPDrUfbExlUSAhmxCY7z1ftoy1VayMbwDHfKH
aL0GbbYocvRDlNUjJz6UhBVbTp4Hvw/idP3Ztj1CDdDtx5yJiDxaVTQA4Oro3cJhj8bt8xkPW+mf
0U5suPaftPSURqg+feBmPZlOJ/qySBtJjhqVkAPYQ3v5gC3HasSgEa/EOO8sl+lLinHAjO7OsvvF
70ik0HbasYJTvpHhuckfqpznagrh0JZslWaOA36B5Dw5sb7XWDn+SAkyyvpqezoL6YWOtPIV24su
nJC0tU+MVhpnHhWu465A4IeSzv82YOrWg/T/677FWgay0+xupzWfeVrF+CXx27IzpRvYMBeJDyfW
Ug2a6eGB/z7CcW3uKXn1+KYgD7zj+dptQMjuuTVR2eZUqwpJFaxHBB6k9wL6btEW6+8FqQ64WioV
4XyU1vaK5uBtmp2+QO0JzK2tha1oq9ky7JOcoKWSEpDKaLrEeL+cS5COdFQ4M2zTPy4UyfMvh3yI
AaxMbmE1yz4Y2dZiempGpbgHaFn6GQymD3CHgj1SlacMNEiU/zjvGy8HaiEhcMHecreV/5Bc0lpc
HJi+ql8LnyXVmFFypqjJIdHosBTG1FEiMEuod1UKSs2upxzxPmhdAMybWQfbCdusNoBd3nAnerEp
jk4AEoZEP3vCtjVGQlbPu/nH/meziM/unG9vukR/QjKSUCBc72z4BVAT5MLMEXaJ4ZWilKHWF1PY
nMtLznuDv8ImzEoaadUoWhdJxy+vZS1YqyAYscUyMER8/eVBIONKLEujs8iablL43xmOCyGRZya0
CsVIuDffYwTO0accKJAN5ndnWE7cegq44ftOP47m94hSxyNs76YVctOr7nXkrh0Z2A1POh1Kd9R5
YqW4ecTHA5NMkhe1b1cmLGA4edVM/iAIp4qteoN9mO0TT9Z0BvQiNUV5rtpDAIQMlFpcXkmta76u
nVxw32M1VD/fWOJXittALxjSyWMhxf5TtHg596l0nxe+Ss2jLEmFSB33tuXXcMNVfGPN2wNjs9Dh
VKDvlsESoF0rvPySm9l/NMbr/gdPZCVtHbVijrPQT/KagrkVc6kafG34c3byyzfRT4lE5IhbVPXl
2UnJFqt5oF7rrZ4c9cWwePfI6MHAfJ153m4tW+BjTMka+ESQdjSQigyUxbQMfTZTO99it+tZ1VdP
R4BcYLZq9RkaWIBLw5pkplId2VHHtk3ZEpS3VEOke2KAw5wk7IbnVicZSdQj45z5DJ+DEyiLwCaz
lNuIhZbJ1ReWMuFJfaDvOnNsII+oduX7TiIE45Rt94gj7KWkX6+nJBSUU8bJGxvDQ9Xq7h1629FA
HRtMol8zFHEiHP2BClzCJKNNbseM5gUlPXRMTPxjHrZZ0YFlRmMqzPNV2eIhpBhYHaBUatPDoQe9
Q+5T6rFXWAlHh1DXcmhApIa354dYS8mkF95g175XcnaGUkx/BMRmbAob9LM81FHDz5CNgPUZhAG/
XAB/cZp0fG/Pds8Y6StsknYh9SuZkbS2NLa/+E/5f1qzAKJ39fmYyIVl/C9yOOWDj5sSqAGtsGAs
G7V4Xac77iwYRaiGCZvnN9aIN7FFcsG3HEp5WRne3THBlDn0YpXL2r3Hxzg8LwSg//eJZxSlIpGi
qSz61RsbdbsDqokjdtiNU6eJhvh/LJeAoCqVzNaLNGIhABzLaBbvWTHEaXmY1DxkBrDx/LbgSHb1
DwqkAdZ0Z0BBuvteZ8t2g+uZ1hGGfkT9KLOdPchqKEzTwVuQYN4kYmLUzRxyKjTGzWPmnem3Z69/
SxKoAt94t6onVn0jVR8GIAM7hGEJ+H2xuJElwSbzGcBnRD0HczSuiHVNpKlvWy2wKHzg+mn4uHsN
aBAgwmky0zEDLs7xWlAXNz+/MHwXQVvSI3N+iTyNefJX1s4lhDgdiGiFcamwWZIvFg3OnGhQYLMV
4ImB5CGkO3vp8Q2+5hAZcc+Nf13aYySrnXpY68z+GXI0NZXS1RpzPdesN91SGL9TfEeUcHbxi6Ku
qpmsYVqYgUVskBfnARw+Yqk5JixOeHdDTnZ009bAAPBYab8xAXIj3xETAXEtHpHapTNI527ON8uN
oPgicVfsUsETJmrt0xmRBbBuCvSyEWlO61gVACaOWUrKEnIm39Yvn34NClFHMRwCJ4PgrMkoQnmO
1gidZb29AMlzC2SE6xTEe5O5NW0QZszfHHsWGeb3f8bS7wqTcNBF6fLjNaMimOQCjrfe1MfHQuJi
Z9ae1e16coSPTXhxV3tQAoWp89Dq8PiwB4CZsOpJGt9Z2pBV8Dsc6aW8XA7ty+ofrerrHXt47YG4
+52yDgN+R8R8m/MZiVRvjT3iVNhrwjVBhwJqM4vsNI7B0XXKkDZqPU2VNsdhjB+k7OQRKJN3CPYH
gjuE4DBTvyZabUG/YByRdHXJbLEDBZjwq+7FsNuCFxNz6IKOPgnLE37Igan4glvWrWe7K5P+k1R2
7UA3/DnAcCIgmHxjMaSygI93lKXzoKE8oGhg1S+7/QnRFpDE6gt5q1gdPflXeTMUbPe9VzjXDpb9
j8uq0v17VoOWNZgzla+eO54LyuuRatv0T3juoi3DT3LweO7w7T3LkA4p8gwWLrI6LYcqltKMrTBX
bRybBZqzzZKeMV1jgf9OK+5ro4Z5z+QNbbVCK8HurCDEYUKMo2ekjuHR/qEPPCQg51g0e7P/Cx+g
h/u8jvQcN2MhSlPjB5r5pFVpT+rqXtkMOn9qE+ebZlJKngZU9gMD8tVNbwg48ERG8Cofi0rmtObm
mV88BO1F6OY2/sTLK/Yar6yjXokrncUo6W89GEqZtkabQxQzSgJgYFjdm7MkC9ElNZqGsIXIYfnt
3yLOOI9cABgmQU3CDlSh2Bac5o0tREW39RxKPVelZoLvIgvFePJsF70sByuJsZm9QBzUzUBlDNBL
RhhsSYkefj5aNc7cbLW8gYGo0D4r2h5EeK6UQfIoQ2juzYFP7pSTWgVR6mnplVgNxmUsOjU4q8AU
h2avHuHTC/XYvD7crTgeifOZfvPm2TTXuW101pJPnlxFDxhDMsJTyKOXJfuUGy743JdmTcvZz4UJ
Axi2izljPWPyClsmP4bG52pNDlH5yK9XjRNQGdvgSlh39sZaXpvGUL99aMy69ZdUYHhtx64qCYB+
9Ga+UvRhPMnytert+02GQNqfjcRLQqtF6f6wrrHxqrF4IQEKlULyJbd7uZxeBRduIQLn4qCVR8oL
u+Lw0fM1GYxuSKOCk0QHr9SqY7Qw8gUhUYCENMVBuHaz/ZmQyVFIO4O34hOBOmyJCzvP1AHFv091
uUnx65Jtdsb5Q0aMFjiXb9Pc829t9goTE5auQ0oGjV9xuZ6lTJYfAyAtsDAXfMJmOR4yD7zaR9Ss
zIEZsJU4Q74oglOvXE8XBEwwyPPX2OQNTNkB0QjAnDsmP/4OzVnfWZXhNK6apya2ShWTD0yKveV8
pA9oD4Nn4BgWVlqfRgkqbzAGFd6dVxarR623uVyw5cYVmj9DqcDDKEN+R2rSttbhr4rkkZnNO+GN
nXXX8utSRGJTu6zoZSmCD7CDDh36VEROjz5qh8rGvVEF9iKbhqh5M4OZZhHQGpT2jW4icQhJzIdb
G1lJ/gYxf39ynLXQWx1UFvs1K2HqbuLd/jLxgyEJkQUYRKeE2P9Oh6mNdybnv3pxbRcdWOxbQNTc
V2fwYCf5Pwm8Laiy1P59ntV2CIgQOw2s9HJt108SGcu+duRbtOI4uJOzPWegZHMBdSUSmBvQUfo9
M2594X+TKjblLvsl1vCxt8pZgouhZ3vrTqDViRrLYfXeqHN+zk+L546zdbjC22H4v5gods8Xy0YL
6LA9c75GVCd+A8JZgVFmcG76HcwN+Ve1vVjiLLoVif2GT0hl8vDZ/pWIRHNRdyptqkoWkEgThzcM
NC3JhhDSKc479x6SxFmAUL3icVU7/YUrvEBgcwPbYXh0as2rTqnEWj9g/XKYuGqQEPswHodGChnl
4s/ZeuAdns4kuTUSr9k3uYgdAh5nAapPkAeQ2M6NpTzs0EvKXn6iapU0zPVMkq4x/PJ6/wjhy3f7
+Ctlj5J9P3hImPysdwBCqFIWI9Nh4jZEqPU3rmoybjAtJLAGpZAJVgxdY10TR6ot1AW7MNPFyqpS
2VZhbyL0CQ1F8t0b12zD4oppqyTLQN39Bq99Hx/SNlYvLCeo8xsdEuVsjpOWGgaMu18/VLDALzdT
pKF4zjOwShxtQnOpeNJXT0hcEI2zK2G3qe0UIXVyONSXN6+H1QQODYD46ur24oX0tgny3gCKT9Ld
atqdQxBC+lPP4rkSMNmKEUChbD+zRKqE4jaAxLpYiDBsYhIwEFX34eFddrEovz1xJaoDOCBNsjxK
QQkDSeHmOvWfBR7yXEVUFvU5Ah5DLvkYwdh7+6ifGDIWWeEw1tOfwJchKHvbXf/KdVRv2heicQXl
AsYEYD4K5woFnUqIEyp6YtokeCqvu2gsE60LQC2WfOsDKLOEofHGE5SSBU3d4Fpi2da9Q7KCkHmq
ruASzQncDXWDTRQfgPPypUYpXYgJYWwZsbdszU93Gozn0+FuSESZRTChGcB1WLn6MUVFDofGfgUK
ipkqJmRigwBUmQmM/pVuImmTxmkIp8sGOA9KllsmQbZMbgp0kS+9sgV87e/CJRzOV5Vp9DvCP0AB
kfFn+Psoih6icKOAeG/r5JuztceoXF6cpKLE4Z+l8HzfeSpzIiBWcM+PtcTGpbZ+g448j9h5oNLj
I0O6ZqWfHsaAQQfJhA01rpOSvEX2Cr1IGa4Yjm2X++Tq1wfa+bIGVJ21byP02Ea7yhjFmYzM+OnR
NzDlbZEg3GwnixY//+FvWcAdpH0EBZhhL4O0a0dAtmdkh1UWCCfo+uCHrfqpJfSAkoSZuvB0GdVR
5M1SHZmhwb68ivgA0vl7Nww+0sIGlgUgidUiHtY5Rb+BSImyWxqjGdixSq0+RaHqYhwHXwWFOFIp
OPOmmBiOnZwhN2o2D3+AE9FOphgGFtTUt7hZ/8aQllEVDrEbFjs2eMvpRue69K+08eHihz3EIvga
W5zqG7dcQ14Oe1tbMpqCQsEEztgFAhj31WCikBd3uXzSG802hXSD7cSOWXTsbxDEaaOeGU8gwH3I
NYyRyJ0jv2F9ozswU+xGcrlLrSR9yx2GoK7fQprZSFaoW2SeWCFqSblW63OtsLHo8bAycsY0iZjI
1gCkxRAIfoiEyPBE7ppJcOz+V28Vv7dnyk0Xt8VYoURch0g5QvcleRbrh8NhdP06Ddw/WAg1AdCH
rtxUmOjazzGLwowhYPix09D9Ho5eJw/jFFNr6otrulS0gHuIRSln0Atj09vJ0aseuEXzQK2vrgno
RCF7hEaKRqz/ZyhAbBju0l6MoFwE8tO0s/fXBXEMH8jw/m/inFC9xJV5hfF2fYIsmDdnKyWB6m+Z
YMaZajMX1JvYRcdfSys+3JFUq5tdSuJvG+Ly76NSSgpnLETe8IPI5pF8icrUCL0WoGMg+KAVIiSq
mZa1IhI08sNrVzgCMw9ioupgS/QFkn0v8jH6XqHU7KyBXqTVnbkVtZzqPAafXnQFV4ldEZIVYjc7
/Jdu+9qhoS+qysDef1xhT4Mjbtb1N0o60H1Nnr3k36tNRFQJPOygaJwCgkTNkmmgbFVtfCC4G+/f
XJF9NAz/gRbav1GJChYYu04zlm81/QwER9NPxv/rixQVifjO7Sg697t9A+mVOBNgPqC5/ImpFCRH
+OAy3ZAKGuHcf/qJVoP3OnX4e5ml1QFA1BhP0oqQ3X4Z554uLMpn4tfJWyZlRGAJ7b+kGx04mgK3
jcSIm7E0vSo2xJbpL55v/tQrNEi//LPeKFkJQDAKo4lLDHgIsJDBeYfPVi2WtVNVyMJR/qmpb9CE
05vGGpesla/QRqSjmPAlTxkK5WemF/D4AvEKeXaJxu9PefzqSvhYgj53igeww0gOHFGo9mcvwwR9
uUneovPDEGIZEV+6kVQ18IIhX9qa874vY97MKxziFnyak0mvoOXOQB4onNek/D8pHI8pAEpsHJ5F
7ElYfeT0tTvRaRXRB/ZAq4aXc/BgeyIrSfPtA5nMYapLMS5VH/jqCttEPtuYkY6j5c/jL6kPq6gP
3EaP/USThB+9I9scijn4vKnMLTuarLa975UWS/erXAlpDmwPRrD7sNPcrkv99OWPLN+dLs5YKwcF
0p5FgPudqHQmbnmVs9K1bHFs/heodqw3rUfOt9UGjn6LCI2iRb2lyWa7KcdSpRQCwOjkttx9mDOQ
5sMy4ixyQuLvIkYtr+bejY8u7+jfhMZtF1dmD6kMhmvUlfan8Bvmz5mJPtWI72JOBTTxheH1v/pe
pu4xYic0L5hrkZDYKnf58vUCvNlO+BQTqZGLS6L+aWbNbzi2FZ7xBT98iV4Kmde9gFbIK6sPaG8A
8yusvvm9x6taOyaGNft410y1D0oe/TpQoNq7KRI8pq4t5QYc+vRzV2TnA1u8yv15BL9HQdYCNe0J
uCQ88675ENYA5bWtNjvAoaTAVxiPg5GMkDD0GZbnf/xiXLh83bI1A1TzvaGPmKDLOjfMJtzhKG4b
dFi7O/NsMsvqPywus2/HHh/iX/N3YDBKQ71405fMdkbz5AtVOAIfIQEAZJpG1vdWGyFMdVMk0rD7
yp0KsIWIx1r6oviWHvC1yKMdbKgAIQY+SgNDSnoslaYRBAO6aI31k70ydsfaJ/Zv2Ij7DUPc2WGr
xv2pibYcNAiDoSGH48Y7RyY4QFadIWBzRYQ5tyH1AAXFuspJOBXGLLBRrPtrvT/OiPniFw4kd/Vk
O31kOoGyDVEeurtpnZWTJGK74cjQ6cN885tCvkyrjbEKr88Iu1Vb610MDrfsWvH4fONEPCA5fgnx
aJHYEpex4ycKO6q1gbIv2+9hrkJFY6R/thnVIg+Uc+ewIJURGCcK1u3oI6cw0AbnvhUNEjbaHjJd
xe+xKdNvMpuqgEkOzSI4be88FFEBW1IUDBOEdiYaiR8xpvY/tCG0VO6NSjWAqGCiHRunoR/VplDv
rvYYiB4KwMXX8O9iYadyj0yOlEodUn8orQjEyN9dZLSWpyiVRnHH5n3XU59EMs8pcqCLWLHHhfHx
PrH/5hINwJ2Dd719MYCh1cr68gN+vW4YxPcwNxGhv03CjC4jUSYY2ocOHLhwoR9hl2NiGglz6V17
uoaF0b84eL6enDDWXEXn6paBybVKr3BN0i4fkyBA8lCgD+z4/55+JqxUEXEqt5l7IDUms40EFMec
EBUlXWpWHeb/2cr6uecg0/NB/0zbqx8dWDgSvqlpIEpANJF5sTFSAbmsTIyNmkgqvB4eqw2Q83h2
CZePTsm9KkuV7LKyb19AG0MsNc4/+TkIXtxMtftmHjpySOZwDsT//oMbeBtaZiwSxU62Yr28ON+t
tD23PF5LgkB701Meola6Rf2bK2mdBICYslznZADpxXycSD7IVW3Q27Hs/K6aLF3O4yYn+pIri0Oj
KKGAGbqGhJ4z+JrTnbAC5ZvyP2CXPktR8BvvSD2VFBiyKp7oDr6Otk83JJOLISCFXpyuAmj1iiwK
w5IhG+PZWLaO1pUyn5aaU3+afZo87ry6IePZzeKCYI9i6MbTZQFH49JKXWs9ewnyJn8ed9xUY/1T
G8LEnfE1oD4Ubv0FKA5VZqK56kMCfLeYw8ubvMrMvnD5T5rlrNtiw0vJ822J1IQaca4m32GHstYR
76H5GLK9bYJzbIX4ZEiuZmNEAXs2psc6Njv4klgYMr85weuZUHEOCXfYJSvoFU/Obyf8dYoozza9
WBPn1ZhsjclAE71ETlY5IIy8UIqBPJ2QhUMv5eSpKQAB0uvR96JhxjzvXP9f1dLj6yegDc+bSVJD
kakP2xMF92bAg2MLcKD6maG117i21yrsu9qukYdiTpkHKz7vqUpzsvYKDOWOp0ifL2Ae4gSPiQNv
wPPlFDo4o3u06wizOn/Bx4cRBKoju31KDV5W0IB63VVmtYw1X+yj7ZvsVANXTiWW7MyFEjY/hFOP
Gs5xLLEAvFVZvpmdwHBuSBaO9Ky8jpv1MtqiMhIX78RZeHsyuchzJ31qCEbd2ledEHu1earFhqcJ
z+dyiu2961qi3vqbDxqvlLko0s2xXPLW6T8AhMTE7uAVxwCwtIOowDlvvhfcgwDyMdauPh2IYuqn
ZTPn5v59uzLHY4YuBSeiHtyW1LvezkNFrlSPePseR3neUseTx63QaxCBot3SbGjdQG4HZlNNr4bz
DrvE8xW5BZd8kzJtEjt8UY7HgDYIE9iP1KJHpgjF5oQnYC2qtUZPUafEUBKkPSIuQjU8bKv1HXZq
fbQsgXRP6tVv8pCDnJ55MRRGnLA/jAN3YSLvoLPgxe5J9SkfmwuXhNviPAXsZnESk5kSgSguN/Ap
LJPQWTt9cHVd5adfQDtJW8YkVp4fMrFIMa8m3QllzpPANIX9UTr0Ds149JpkG+rgD2cgrci79dfB
21sewJgf4FB9iMdWzT91nvU3k3OPyh43OV+uHr8yh5CpQSgBbctrRLfY7wW0FFoinB/GV9tmogM2
n9LTFXL7yQE4SO6vDEt1KK41RfheD0zhnDRI4dXc7eJmf8+d09Q7/GRASVpT0D5qly5h0R28CwD9
BMkr0rQOwC1fIk6w1LPYc6W1rJudRpNe2vPZqEgMN47a7vmJs1u8SeqC/B0Hf841cM0BSn+yQnM2
mKvJEF5Q4ndIzRxGe+8TudRQhyruiCe2j5aI46pb55a8WniSMDCKJwFUNLj2qQr5Eo0Gyx6fm8CB
QUOA+PwMHfK2zlocfaiyqoDmhaopxcqtuGWJoxIOHnCJ1F7vfKB5AglmF364f7AmGn6MajckKRtd
UTRLBIc2LT6cychuEChx06m8bUyj2yh4zB6Moe/GSWWL0wyZkC0Mu6pFT2pJyGvYA2ubXY7omS/K
1CTWcdr6+dhWnKfj/K1XOfwx331pJqaAL4gUlSuhu+6dUKmZPlNe1kDwF0XwONexiz9OtSmWNgqg
Ks1RjuwCe6i6StPmAVXwA9SJZQiWTXFhhqIyosUW4tnakfEHovaEqQbFZJFu3VKipYTPE4/kKFx4
OCMsd7yN42IfAXyJtBr3zd1inn9E6EGosEzDCjbsYPojqmupbOvS1+d9B6fXj2kyDusjn+q7ev8c
v+LEk2+x8RlYIg/Ukq4XUuHjvNVByOwPxKDG5jPZQNNCerC+/Fh5IPjNj0Lk3n4B5VlHVNoBasgJ
jQ5xdIezme0/LvgRb/cl3Px8w02ngqq2u2X6up+XYF3qvRwoxvqbMo7SWSxyrWvRTnnM95QpZOyw
ZJgoOoAJPU9XlG3g1KkAkj1kbP933wDkyh5AF4vvMagxeqsD/Hf2ko3pitrpy589QcmUqQu0eu16
Q6aiK7Y4lj0dwUWKVxqDknBTvvj+FrRT4uyLiOuEnSG4zRC9teuhGlpJcR/AB2spQf4kv/0Jgz1F
lDrW9lGb42MhSk2wsDK/Icpsxh2IHWVCDevdQVsaT/B2H61+9XxdDnzi96T/QPNVt5TMAvv0BQuD
JjigW/YZtXQbUFpX1ORgg1ww1OgWn1h4e7vKtWwBjXLMeHW5MuHZh4t9qitCyoCIDo/fJUboyCmp
i6wMwnd+7y7LZf51YrxMRI+u7dnbWfMOfZpKgUxQk7zx35/IDv/Hy56hw9VUyYJ31GajcV6dsvyZ
H42Fg+TBY9d9sWt4Ad3cCgQtUmhx6f+6QPxR6W+gtqkUlh8oSY7ZLTED3awIHv0w9J1aGZ3b5XCD
J9JPIDnKHT7mhoLJSOkm2jjssPkyae6tdBpAp9uxXXWKGDwNn1M6fKDpaJ11EwZj2ttKvGObPNTg
GLz1u4jJwaNJZvpLAsTlpZFQypYl1pZ/Ctyexofcm6oUi2zWPz/Jz3b9VsZsnV8tvHlbl0cfncWi
LKdB+yOsSVnpRwZ5a2A+q3iTEUVLbV3KKZjIsE7V6frzhC62/+TklxyNro5SHmHWqIA+yB38dRP2
7lzO39hDYUMloz3JXFFZqqO09yQYtk2ygg1QqZ4bWbYg5VQyrjS+3OyVTFyWuzUnu7PiJbools7n
E4OxjPpKjVGoUfpSStyaix7fRLQRgHJcwHaArigTbCGAhF4+x2Jd1+PBCEQ43tVJSNESEAf7UGsb
QycITb+qS/3SV3osnbOIMrz3uyU9CW2aXrMlokQE6v6Z8mvCg5vGfw4S6sZtIQe8Plq+Lisg6gPK
YpmvpTI+bPj7vHp43xXXgPiiVimDh0j1MAnvi7zCi6JJItZlNbtvKTQ7iiamIjn7q2zWPIWlYv5Q
0mgCxMOTwT/rx6HyG28hbnZ6D670F0RwTtrzFMHl8wxjGTtkYoY6Olt9epnXbqx27FzwlK/k7y+L
YoZNokuUhKOoSKNxp+16YwJ3noi4TJ3K8HOhVKuu4Hub9h7OG2ReWFKR/K5XGOpyoZXCaiAr+aFG
DJTIjLbclkt9Wqo2DZZOTre7qDd+9gnbMe/+UfytC+IMXnco4OrXUtAJhp37m0sINXQpWTvnGkZd
/XgQn3EAopUje6yhbMR8BHA49A/GYAjrMf2cWHH6VnRz+9mtbuatriih72XEWZKyMIlRIhYL/OIN
2zR+74VDDnWudUOcpRRdGyLWtnnllSj5tvTccr4xTF5TVqN1iae42vQDNjIj03JkCz4DRpRxStrd
P7CLiNr6RXJooNAX4TmA3/8TNMPcHoj+cnLTXGKekCEnDe3rsUMpK1P/AGK97dUuauPREZSglj3W
Oca8D4idxVNjiM2n6v6EKapFrv54iaQtFySTraIQItHJMyg8Z1hdW6x0n7t0xAzoxmBqxag4oFIC
WK0XEiaB5DHBfSWU/aIDkvadtbBBSZdyu24t8h+7njJTMh5TECHUh4jyCVHK+myyd7ok8lfQ/pG1
R8hQZ91BGYTRnQp597H2T7RsKY9F15Mpom7jpm1lv32QjRuBsmOVgoAfzC7c07JqaiHlo1dCtOyh
b4tkFu2NLNtmQ0uEUx+qHd5Em5WF1Dt9QBP3kw0jthFhv4GOsDI+m3ctjJ1n/plCOmXImDybifBy
nGPGkKPWqdizYTKUrS7Y3TwNPftpCB1GxcvoPCILsEAZuY4Slk1Fp9bYaCAw/uzBSBKpX9P72WZn
N7BGiqXcQdth6E+WC+AUXXCOWL4Py/Xgg1FzLxEZAt58wVvGBrHkMjmyh9IANO+RvhpyrhjpxDRQ
k2//hU+Q4NV+YP0ZAfMw8mOjonKnqp3rNBLPJbPBJsGx4MncIN7OrEuHqwCA4V8OqUUnMPYAE9v0
PfGFg82VEa7WvclfAzT1h11xLyiadlx/Rl44HoSBkUxRDpHcJW5/d2FBy6w/V9yjcgfwbtZoeKBB
FR6gD/dz4VTko+5kYuC9Sf1A24ERxHaBh/jRFsnd1TkHcv2tKDnMlyPuUMYNDUgDL9loY8dR2JH7
6z28Lux3qr/475iI5HQdnY90St5WLcWWGnnJwGZO95mmseEuvQfGQtvX79ZgUcC2YSlP7J7VSNBl
36l1hDlpn8XDQKgD8SlWUAZylkYzKDciIFaBfcHDcYBUJHt+RVjCZcDMbOJU05H/8/fVd3KUglg4
XnoE2OtHbI5NvKK5dKApMzIGMe/rXmYvVIX99psIPAud3bCtILrrZ7ENaBVSyFS3DZ1wxrGLar9k
KAb2Q0ySKlJ6bE12jzPx6p2x4OiNy4wmoJoK/7lLd6F8qs6rS9heTtKoAxA042XR9lDH9gUUWw/L
JsDC9ZamS5lI4F7tBbgXnx/4LIGGISb23N1ii8obh7gl7e90fs1Qs+La7awRUt+3+qNwKsCgHmLc
0zAOSgBSyPx7jBnyuUyHWfwyH+jOEnCJYoOHGIwc6Gg+hAg0s/p15tSIfu+DbmX7JS7OQRmDDY6W
rtNRUjyLMzEdBCzB02u1R8rPGvqYakDkazlrPic3ztg2yxKF1LNLEpMvIWalkEhutEvyQGAgmZbv
xHx4/GCBklLhiOaYvSGbGUX/A/CLGFsfdiZ/MLO4xSCKdr1/qtyQmgV7i8lavH2s1JkEBjdnHzu0
SAjL45TAuo0aEV6zdZdGVKUSDpMo4wg9CDhC0huwbFSVMuVeJxOvfxJ4ZUYcZ59g4zcJaxOGuv6G
yXgtN1LluHcZj+cPAO1Aoccr8f/UkzvrKXlNvmhElZH5ku1XOENPpXDoe5l5/VUPA347uYCmXX8T
kpK2k2jI72t9sY2BT/2ClmCyVYFP8inpEeKUth6LuUB6z3L05UtqXghPy3eSXUE6qs41W6nKSX95
R5gIR/B9qIPxPw1BLSchp7pK/2xEAIwJsh2pWbS5qK/3/yKNPaGlh7hYd1uAAgkzI6tdPd/egDRK
Oa61+/82fBgiCiqUWcvL8mxSihvv+WxbmxDHuuDQ/p20oHXXUHyLa1PgJif8yYvB47aIlVQQNdn6
7W6iRvsRVWFu/c2KLv+xzvVGh+nv/+jRSAVaNLkw0X7c7AQq5cW7Gqr68p8YDnel6MDaGzw7xw2r
YEh0SaVrOGWrS0D4zEn3djx7jWMu2VTwKONNMy0ROr3307dSUfM+pvbQk1TIskZzi6rfLuuY0clJ
NK0aCjugYQhfqsil6WbSK5XHFtDV0eWZ3mHfkjuvaF1mArF9JaqiKTm3tX08O/i06FZQErNMyCow
MdFx461Oqw2PqMp7f5yX1+DycFSWg2hvJ4DtyqV0ZccPW1BX9WJ426T3B8Gr5vZgeyToDYNOZhDq
w9l6wbIWg4JJMHU26122WWSmp8J8df+KkdwNehBTlGEwkmH/S35EKH7CciNe4lLd7y7jTxDRUUU2
U6WGQqOnBIhWlarAY2K+tv3YyW3h3KW+R7qWiHhxc/qjkBPq89n6P0do/YylwY8f8q6FfJLqESO5
0+azcJ3lJBRNR2eWxaTawBHWCQ+eQ6Htga5rWKYHWfyGzzKiE6CCLId7h1WtU9tPDpmFBa2+hmNp
RoR/Hon64E1zy4NpOBkVnzNV4uaW/GvpS7BPX+v/GFoe88XtGTV6/oUPkf/2OlUbBi4fNaXqf7q9
ZR2IZ+zWWFcMXCMekAjIhxLhjvpy9ReRrJ/1u1D/JvmnJ4/m7oyaMsGhMRq9p5tWIwLgTIFRzAiX
SYjEuYHlmJ7rhXLIvLO0Y47Iff5MCqIZt1tPcILwGWlxt8H5HeTUKhmKBIGqV5bqH3Jw5nLVTaHM
5b0dGZBsJ+o90t0vhJZX+rkDJa04SNzlXNJmigWSqaoL0d2gELorl00XFbCsTwXLTu6ek1DUHYWN
ddGQMTY9HhaQj6dNLJ5hUklHft03lHt3A+hEIdydK1aHXldMXPa6G7hblr3KGdttaBgwr0YJExCE
dvALF1WWt2Fdemk8dzEHU5MjRa0/31EDJLmnHrslZ7wAmV4PRjV2L9C0ZGV3dK9en0oo0aFa+0aS
88r3p2L8ehgmJs6SDHf2seF9CFagGVNzwcXPiyD54G2DlMLhAl016AIUiNWTvCWcEDC82bRQ+8u/
qnSMIspR8d9hzntIKsLFzenyc+VoMzOY8DZU6EmBUNZQj0bd80TcnOyXzfgbfTy4aOeqDSt6faMX
nAcXKEoUgtZSuOcuZmGUzWNUYGPY29SWtOPExGYKOHd2yh7yt4KjZd18Svh8de3vXPoZB2gCoba9
LE9LLoyX/J/JBxAlVYhMzFJrkKEraat6I3Dt3tMhOh9AbpnhoGjTT8Nz2H3N2EgPPg7IsDQdyig2
yUMRrnUHAqO0Btsv19XOLB+aY4cQgsM0dFcIzjCnrQnz6Ps+3Wmplvk73J7vyHfaNH7ixUTs+iwW
0o6jDfkwxF08xytIdKXUF1gyIeQw3PrZOo65RaI9t+Z4Y7Yzckb4gl9zkmlH6jyb1sZZdDqe2pvO
7xCD7dDq+0IzuGrnDSXcifHib8YyfGQlnN++O+XJZ8aGWP9KOjsiNDCyIRUzuDSx9h3RtGi1/xDw
op4R2o7Ld15hwzLKw2nF36qhNL4/RsUpeS6CAKmGJdIPlrDkdkZff/3+e0ZyjYlWKvvBc6z3ptkT
zfEUCN4GsKrZ2Jtcg+Hp2hZC/1JLoFo+u6NqsgFgta9FiclPhw5JaXT6QqJVKADTvLNiUIJ1gE6O
hudjUq96IEIWu1wqw8Xd2FZ87lWWP6dCHgHfq+VrQZx8QkHD7FnrEuwSXLAH6jC2ZYJlzDolvEu7
FnR1UI7CkRJgafPdmiZi83CgdpgzMyn4juxvOEvPcszN9gU0k4aFk4+Ap6XsFq1PLvREc3Rr7MI6
8vtffMMUanCvtEgo0y3Z/m+ajbAwJoNECg9kBQ9fhw73LnuWsQ30Tz0ZfNOug7EUHtzQPuaALKgR
rfbO+eQD5xo/Ht0hEcZiJOdKxfrSbV0faH9Oyx6W5ayfCYqsJYy+Eh/YxKeRQ5PZ5YigJTB+LvcP
qCU8bTatj1pBRYhp1NLwJavNPyvpRA69F2rEFDxi2iyTYTqf88tAm4vPGoLuxDiNhwyiGPVrkqmF
yiX10Loj3dP9FIKR+/jbHUD0IP/xSqXFKbGg3Kq5UJvPjSSmxaC8++kslEQPdbiL8Api8anBxvQt
EfQuLQ8eNEP8TSyA4cPUgl3TDtxGBlOxPQbF8W9g97WfKtWhEx1MJUnGKX4kjuonb2entJ8+RuRu
4qavngtdM508H5UjijzAjWOzd13+TCxo/buPLtvOFoGjqGAnNB+49qDGz1hnmBkOsO+iHjC0/2uf
vHtISDvERMcLhIfd4SPcMEkC/RRGxYZv6oR8+37cmGhZGYc2/IuBS06BqUGKSoZ38LHwAE4VAnhm
doyLpK1KiDx3I1U/qNO1hh4G8Ra345Eed8e0bNUsOMYOdq7L5tsJJJ06srEvhlbwnaP8AcB+tOOl
RnZM4V73/8nZB6SrldW8HSDf04XJcyPy8PUNUib5rN4m2myQS+KM1PT9tDioa0404nMW8/YQhpg0
8uYPqdBaPzdQHYViRBYmx7MzbAWnl9OKiuLwyTZHmstO72JzznrwWduARJfU7P9n/LhPy9MNFm9y
wj8aHsinYbvfSxnk9T6zVfZLa1I03cf6cNUMKZFOcXmbsURq0nUzKdl009DqcpDnDCGlCVxBTopf
dDf/D64+bnM4Y+8T7x35T1CLWcGJdkMs6uZvLMLnzxsV8olx3SNSj/mgI77SozrPzjPyXnBFjoG2
k0FU7QhqsvSNAfzlgwh7Vv7abrubr9958EqsqAS2lXCCsSoe2F766gymdJLZtVDrsoWeRl8LPA3e
Qbc9Abtw+BYbWxYWbfp9aBrwGxHHS8uOPttFzcnH1cqBCpEqJxduU8Oke7TlLV91PT3nnVKU6xmP
6AwvUe9HrEcAfIGcUoQhmTigHit1o5cQjTffW2SkF1mkaovzdv8vYP+GVLHoOTguD37JdY12ZOxy
1dCSfz5YyLWP6GDp7Ogj8VTl9q3WRja1VJunIsz0m0n6ZDxmRZUFThcKfVtigmKiXYtfWFwXcX7x
50aVKrh3iSXC7N5P7Hb9S9nZYXoydKybF9met+Li9RJDKsVQr3M6XHDC1ZzceTMTW2tKFgq/G08N
/q/6Lp9CvUyUm9cfh6VZHrac1H7Wi5ld3b2q2ZT44PgG2Do8zo3WkSpUB7paz3Q7hU0zkD7tB08n
EWnSxlE6e5HHOQMQXh7fyNFCb4BcNboj/N4+o1m6MFbTZG6v1gtOr+R2Rx11MUHZRhFgt4nkybZl
Hwc5aVoXPUxE+Phm5ljZ/AFraNo6YKfagzgh3RuO/miPR6Ugn0+ZDEYbnFLgtqtn/+ZwsF4QvEPq
3BGOOT+GVW7CzrfGRMGHpko9c3OO1RddjvVfQ3uk1Vs2FGy8ypMP7uDy6PQb7xaHC2luJ/HDJ05p
yZdzVxDD79Vl02STvJpyIQPHx/VvidSFQBnsqdhDCGU6WF4QHz5C7ywFVZF0tCFPxbIqqS9UJ9QG
u4ixq09U1wML1sJHT1HKyNRKTvszsXumZdgVgpi2h85oxgrg+ywMTwoni5Hty+Zw+iBa7XdsiPbH
dzF/r/tU9Gju6RaCiJP8uR/9PRToUA8dEXMt0vsppM9od/Zp413Kxfd0/n+FoYBKpJQOrcA5XSLE
Igmkj1lpRWk45Mt1GRTTR95fjwRQYCcLFtN9fmFA3d0JNFQbCLEO1wUB0Xm8hG0vUHQ85dpIU8mm
WQCIrdJAzQkLtdCmY+ZAUIOD/ELi3zMkcs5xUJRzJ4jSndY2SFB/ct1ecMc+S4EEeB7XPT3+Tsll
yyj+G52SMuky14fLM7WBzZzOizHFmB7XfEX1UOIVQJJY5Ob2sC6he1NiZ63b/+BEef3IWP9RUgsJ
r5y0+gl+ilTUCPVdUcyEanxnhje2tuse41NBIg3yWHD48Z/seTcsV4ACXlSsp49zF2Vn/9yMpdLt
3DOC1iYRI/PMzdsCSU417H+NAHFRj4yBzd7Flt/W+RxpRutKRIEoxu+0NO5fZq/XNAbSiHaRXOr0
vc5dcxyQ9eRnTjZJNDb/Yl7d10+w/xPwEgLNfn5zJwbJ4G4UtRtikagWs4SJVUN7HkoviPkZsG+p
aAu4FJfo+MZJbaqGbAu2ciY0dR3s2svxI/jvIJpT5Wb0js1mtc2V36mU5ayxhqOy1/u3/9M2JCE0
DrZvGdofqbk+/pIkv3sH0ODtzvNzLdxrfHIdbHSPALI7TvHLW926pTiSE+46rGJ8gxczVjbSB7Jm
YpkvTrFKTPPLpe2cnT6URb+sF4Sqi+Svk73dQR9V8nEHNuzJHmNU435oh3a8oEEZSc8l+dJWUHFk
Ze0Lx78EtAx3xNS0bGg469E8+V3O336KCQvppf65Q+TT3CDmK2tC4RX4lH6jIPO4VbRqkXN4V1BG
4D+hRhUWaX2Y2JPQ8JdBJX8PxY5pVi28Xuk6Su5DOF9bWax27ys4p5N3zEKpkicRu/UBPgu/+Wni
0RKZBU+XjNECORbB9Uoyhy86hvHnScVJ/kBeTY1LEipBSOaoIVWv2L9qedNAICgQA3MP3WopFbhL
ZnDx1YkBaR8MWVPKituEeJrJCSROZrqTL/zO+ufixfIewyUhBrbiDDCalZa0Ae8O+lrYPIVOoPL2
j2kMBjKMR5jPY55byXi9RA00t/xKZfp62CNpNKVB188U9S/mWaBdLBOy7Hhcknqyb7xKlzP9B2y6
wPNkprFdIzn8TRf3Mf0+Hge7h5Xp5Z5cySCEjhEb7IR5oR5uUD61sJ6qg0q3rNMRsT8Gx2fdMZkx
hxMmyCNC+T6LvdmkbTpwfW191EJDT6+8/3C5LmYPEq4sybu+bcmO6woi9Q82fYAYIFJDj0MFnaW5
3GuIvXiNb20R9DpiZgYoeUwLTPuq4lklaA41sXrUy1DKp2onUv8tYwdD8MjZA3feg1nM1MVBSbeN
owuKSNShcjyxxe7YwljdEHMAlDGi9DT/AEdR3cPUWezFIlin6qFUVgUtZsm9X4ZHS+59CIbVN1VG
uGKbT94x4BkOLl8TxNiP/W4Lv9Td06wAMsaZCkLHivkUX102rAw8r41czRYmUNe/pco2vtELR+dT
KqyImS56JIsl70nM8GW/fzO5hYv5kpVht3j1JuF8+2tkGVoDeUdepnVGpYMBK09bpo/kHQaO94IV
bC+x1rHW+EUZ6wTxSvWVlb+qbdVvv2IWSYasWe2/2NZEv5JYHo78x3QxBiytcQYj1vW6vmf7wcsS
HeaHxEUYVEZLEwRbu0Sq0shOKRRXpgPAAbsY6i9kiS9GZJpTN63FjeKrOQmEisMzCYLzRNH33m7L
sAi3zVQoPgNC71U2Hna65Y3VPCmnw7a2vbCDi5zaqoDyvjTIR+zbM8WGi+V70pwOxsJuDsxBYer9
EFdgjk5iBBbUVuFIs4Lul5rlX2L+RwDy9i8sRQF8yyEZsEa+p3Q4t2XsAklnVC3PuaownDyQFxQN
GAXQU8p7Iqhwh3uX0AscHY7juWZsMbzuxGa4dzdJczwXxJB3jVNfr8M2fNc0L18pwJWggsy4f0PN
JF7VCAQ2U0XUQD+XopZdz9Zze0pGOg9Ux5o7RujfcnWGt86ydIhwEk8VgM5W/yzPd/vgksaL7q+J
fF1sl1iK1gcoxhA2RQpKo2g2v9Pm+kuTVXPf8CXjXIwGSg/disXVFFPuPudBIZ7o6OZHOGoytKgJ
MmEZBPd56I1awDYT1M5POs2SLjLPvRr3d5DkW8aMlPNHY17ox4qxtRswPILgbJOGMmO9u2vRJWmd
rklO+CFRLlrU7Gf7W4STBsYz/BqN08++yAdWdV4c6z2gLT4daep6ts35qSwyD+575nTuZFqCOYxs
oEN0ERKbwOMcSN//d8nrU4RITVshFOqRLB9UILuk0omwvSywl6EORwxLhJW2EfI8j/NuVoyih6RW
qVynv7vUcozZzQ1R8eofaCVtKagYYSOG7Oe22RROr1wW2PdyjY6UI87YIczFk9pZjGygRDrYzFKA
W339adj0T7eUVH1XXvharAoo0juFe4KUxaWvid3pOUz4e0jo7zqScQPFa9KYCH3SMe/gdDRxvPRV
tpjHtZ/9uBsib7wik6pxTuylBFhzLGXiYFUcRsR3sgaHf0LPD+ptOZ0GphcQuKJ2YFbou1Bhq4vx
1Wj7RwYU/vKLOyvvLccAJMdLlUxXCnkq2XcaCAiYgIEIPZzpLl9yh8SyqpSZItiO/Bp8EEp2yn3t
Z+ugzmkHhgQrBV0pv57fU2PWN1ErGnlvBjEWUwCY5GmpHIFEgy2psxy9nAIRyism67fEr7+DS68Y
uUVyRVG92ZVsSNjYeAQsfddoeDdS1MIOxUphuAstBgX5jSXUEDhv6Gh2M+3EKJerxgYJctx/5Hh/
o7+hYpGaotFh3V24kPDyuHtdwvq0kjovAFxAWQImFz/Imee7AGjtHlBjCF0IleG6QloCff1YIhp8
blTkB38Ea8uX1LB3wydmfbtQG3QZqNTdLPd42XPETN7N9w2d8vlkekuCrN7MaLhqbVhn+iv8l66p
kNhrD16XEFA+bvG55M9Mdd7GzRi9hgd6BCkGlAsHQrM7aiiLLoyGQFO7zoHVoSFkDLLQV1aVZ5s3
VM4bGCTxjcecNi14FrajoHMOhhbrdIcDLjBXxwLixls5hrZoWXA7M+bZg4ngxMeOP4h0/Fhebfp5
xgpTEzjJmtGNKbmZsez0DudhRClboFbhwUqMhvEHtN/FNIegj0Hl87YkAjm2EJaDq3Xg2FDokVNZ
DNry5uW3/uqur/m7mTz/YKpmrgb2uZTJk0NSHVwyHo6/OBaDFZFNWCLyf7KUrmGVr5E96X8v/nSu
sQJu0n6IU8aS6cssDv5QSq2X/9lhmFJWVF+N8xMY2hfmFIKBpPyV2uTAG/cFx3p/3T7etq6Py5K5
HPxf/IEQMBiJ6XjXlFZRUNT5jBDAAYanl0OmcIXT+gpr13HQVSwKrp2vkkYIA07cEY8LzLRXCbO7
yUK4H/gyvMQl47Ic0qKWVItLcpTjiuL842BS4JAP1gEQx5b++rfQw95fPEojazTFefRkuZypL0Rj
TWJTH+/TkoFjo7Tb3k9+ojWzadb5p04BZn3V+dPM7C2+0gXp6HnylbSXSYXNz9icSl3tFBGOmUZg
ZApaPGA8/1/P3YSywylkYmXVEbjN8mrABZE9tReAdGLjcQEiu6sbSpiM1neCMj1FW7IH5hur3MJr
9yuXBV88PzDT+cT4wvLkZIqoo5C9XxNgjnoLRmGn9u5A8CGlk4ZWEHPm6cm1v1ldOkG2xnU7vdzA
hQvyLaV3r0Z94uI6Tr2QDzE1rkyE6Toru+x31/eB3fS4s7AQ0garAlQOT+3197V017bQ56qdfhHz
Zyjs5v8gqI9usDU+/wjP3GLAq6ds14wpPEUmTKE0DGEBnEl69rqJNVFijF2FhG6/+NbEpYi5Vmc1
CpEcfd8oZL8Hd3keqIHVhiH5v0ZDvjOs38Qm3oyqR5mDi1h8P9Klcd4LuhuWaFYOoEh+ouWh97ID
8gR8/0nhL3UiZf0ZbG9IaGC5g7KZXkiZqr10+KdR/Tdb+ipfizvMotHl//G0Rha3WC3OLgjMAbC1
aPIFqz7v/023Th65/WYNdMFgP5h5AfRUAi8e6rmnt2t/kJZByFJrlBO/zQLzXjo140uc2IQrJ+4z
CmIvakOPfq1TVWThBCUhCPYm0a/AxvRxiTkkM2K3ghpVQVetpiMRg3VVd53NGGPoatZs2CTmAlH3
nCih05PC2oG4GGCBFlhzyV7egF9dCx+tmoTywaFgQyCpnLNCBEwGTvE3YsF8238hRguM0XSWpKqF
0E16fWhvbhIJAE+t0CO1d24UpWRliFn5yocFjNWLvfdqi5Lp/Prt48dnw1vVUTWusU1HUjKKPGQu
G56ZIs9Fls+opn/yR13vaczybPMEbOMxh+10M2mZXMfMiycqk+AW9p4jwB1kvzHVo/smb+9hTndJ
FWmvjSyQJteM0NKMoPju4/M7d9j+58oF+m1vQeEtxkI3IcX4BK3UZ8xNYX47uIPFoID0QnWHkY9U
CYidlL+5TqGcQ9cuhflSSSki7dVhudth9kYYBzYOk0wB2guJ25CsutNc1KKFzRB+c13N1LEFUkAw
Cwer8QbDUlgRjc4QbAKdrGcsywZ9+YGKJX3hgMpCXQUUBN1Z60z22tDy5l2AaGEtnq0R419wIV1/
pzo1e6A7soMIZASakwIwxBXimIiPfnAjlIzZXZWgWMKT+GOUYbH4azk+tcX5R6TcuB2lS6bnbvuo
Hzb0l+bSn9CU+5I589J8m/8ZdXORFduyKgzWzwkZwfRpFj4SBv+TnPPjvqnyErajtMlgVpQrJG8f
axtNGf1SHeTkd9SbMiGaHKmC9ZOUZhqCBjrtw3HF296Y4ht+jeAK6fxKAs0NPRK0NUCW4463udrR
0amhZODEW6u4zVtJ7tUJHidgoa/P3p9del3TXlfapufJTYIARQPgByCjmGKh8+JAhb4yBQtXHOh9
QRXcNioDNhD4Xp6SUgKj2IW5OCtyEzYaVdWfTYTzH5nIEuilDiBEKGrnrcQrWhW3XNVBAAfENy39
v8ZJTk0WwZF+H8upl3TypqUBMgrdAjQPJtv9HfR738glya3jUNIZIK1fzMeX/vMPBa7eyNAHc4Hw
o2y5+z+5KfvIlt4g7Q3RLhltObOTyBe0xt75im364u5APUsBJ3o4V+CS/v2sZeisxRHeAP/ogHYu
mCebyepMGJ0gUhKhLtO4b0UFviiawPskfMqBBTpWUGkbsSFqZ/qH3sxjWep5GucNt3HGI8FWQGVs
US3ucfHv9UNPJzS8KC7llI3VGvmRXZcoi8K3gA6imuaQoabpDZslzx9Az12ajEedJfKb9LM4fQAJ
gaDbEW6CY71n3+wfrrmSVTPseTqTC51sv4O/bZ2ic/2Kr2D5egR4Q3OGzhugnQy8TbNOcITsFKyG
U9GXkXuh5qhnSw0iwRPLJhTdL3wcvIPkZxQH2lVVdzCuWqh0UHQho6FbKMZAadadOE7BRfb+REDU
rPqlsUpRNXd3mF3ByuIo6z4+QFZRHxFkwP2PM36rXlB7s+2BgPuSl1CV6OBgHphznSlyxhGDedgQ
LLsDH7jcKY/9H6KfMXxVOAbVRe1SPTNAei3BNDQAC3vRu5G5BAHv11rhJpKUdMPZrBDR+VcUvBLa
nY5jfDDIeKZ9GlPo03kc+XB6tDc3FvegBNVCh41pAFOHzgO/FruPGiObtqrqL/4EAVtaRfEK1afO
Tp3n/AYh/2xvPOsYaMNyMYhghGR0KOrwsvK7kxPuGQHl1IHcpRz03cOE9K8kI70s/BfF5vW9zC78
fghQOEEMehmOF8ugBr3seHKnCU4vuegI2f/oY8HBhuAQ0+6SSIg5oB7kKKrvHf+xEbq9MWE7nS6p
i9uUPAR5PBBtwK0F5oqqQkWX2N8WdGXAHlsVFSuMhy/m7Wftfe+EPc2n3EnLkpfE7ytoHfxaJ2QZ
oKOrwrG1ElkAmaTJNvU1cHUzLTMQTF2fvpVFFddyvziNFrbFW4UUdVEceSmcT+lbdY+IA4SzlMN3
uLZrEkbTiSzFg/Ru0Zwuc/kaoJEDd+gIvc67AN1D21vp0DcXPNM0EQuViRVQ//6iEPIs0F2amj1x
K/RiIhxADdHwBQqbGMLcmnNfF/iw5kwvk+fl97FZ4kYbwuhuEYKi0QLUl/9o/zCfJDVBsSIXVO+y
JqWMh3UmiZH9pWhYx+0eQHCborN+ORaUKingtnggGxaLnO9wFEESR9xyKVNDOAwDofbdZhK7KKJ6
+LdhACVONCkU1bZypy7mvOJKfDVawKvYRPgLCMG99npbEbbDIIAPkYifkedPy1DV8d494U95DGw+
3inpJTWB8uNcaPQJrZT2ezimzKNPqdboobuT3gTk80GWnl3ap59IEb9+WSWaxbIEPpeGEH9ihz8G
/ul5xqjyLnlMECE1fx2yqbiYbcbgANNgwkIFNSOBTVj2EcNO9yGw+hE7Duc+QyOolRlcgi0a5ST5
2++T+b7nkYQZdmRJ/Fnk5KQ3SrMLLMV1Y9jCrH1cxnvFLDdFplCQD0MivM+mUp2fkU7yFQ9alhNh
qMRYRVWCYiqlQbWVaPfB+YnyMxd4s9cVwJgLiOYh/TjA8by12DjvjC3E9e961qyPKC1RdPU3DYPZ
vRZj/ojMnXOUnZ8i2iYwaT+ZVTMxr86Gst1/M7SDAHFgi1ntQuLokzJnYmy0qkP4yVnn7m4l2a99
jY9F9z0LZl0g9XmLwa9wUV6vtHoJW/yX8xgjiQcWLerdZX5Ga5+Jeryn5IiOCUDdT+zPZCqjapYm
Y5f7O04y6ws3ow2ihSSiCvLhzgzGV9kOA2t+KMZxKlkianaUrXmtcdaHxtTD4rCgM3XwUoq8Qrem
RycoAFqMursN0VZOyEAsqj0enxQKFcGVswib50LpJRuG4YIjjxbhY3cDt+TV4y4ZfPLBwbOXr+GO
IoYuwAXpaKU4OvZDA16OaYlX8x2pMMOtoycqczbWS7JeTfjLsvS+7GqAABHbcc/fZ8TKmF9ET3L0
+BgDNGtUef3LpGA3Z70y2za16J8soF0RKzska1J0rxnWq4wtncuSQk/aU4WpXDV8+Qm+Ss8n1sre
Loq3L2mGYHvbHyas1pQlWwtAhCJ3dSEvQ54iCa2JK2FyTH19uc8fqCiUJE11P2PGCCrQ6C9QC/nF
aqatgEjJed4bOxkzAwsPTBNENrn4BPdgsX9RLxdssRIKUoKxY9RjR53Vdz9TZsvIwNuZTy3LMcKR
wLfF1OqPEO7bqJGBEyUBj7F3ZhNNJFiEbbRzg/XatpAvPqPi3lgLU+QVh2EJ3ugkcHluO1R2yeZZ
avdKKKv6FelRVbaeRMjWSp7LFiyN9W4/k+ENnQ6sebyS/V4dlOx5kvEhwm3rRh+7eSPAJM3ULyUP
9SHrUa9dhvMvdGap+1VnRfVQgZuVKzZBestIAOk1FUMPzI5l05YkutqWDQ06DVmhpnXMbPkOCzQI
VHkzDoVse4mxkoRJUOXbjXE4ZojNXdyORkjfIoAipoQUPAkLhXsXTv3uPh+BP+qGLnXlSfP2wZLA
EmqbErPMnfj2rNG0F6shWfBXirkgxF7cXGvNCNvmv4qFSWgAWATxqn8l34GA6vMgCAPe+osT+Du1
rgPx5NzoOgu+H/9+uM+MH70kfjo59C7WEdXZiX8ec4Rb0JcvQDHXX7JzuoA5PYmkWVn4JuTGzHfv
DEmbKUwzVVrvOaidLJRDjwOfjXCcS6gEiXWuoNX0xJgdwrLjsPWhMXfmXVKkzjaoGoZepp99rdGb
O9s/7SXk9XWo2jmPGZ20ok5j9ospRUY/RQLBGfc1FCgIEU7l0nXtiQIkD74qIB0XburcB8KhpYJg
C5ChjWODYlsNtGGyscwjTkIY3fjj2rWIAjqTnnBh2cbMeQjE3gCnh2ICQD96VDwBuoaXqiQZsuBD
goW+YD4TTbZ4f3zzAMjnNPeQEOZYknnid0sODDoJnbssoUAvtX1g4vgK9fIzdHX7BVRh3CLke6iy
BSzkCgbbcFvd26IQnurypziBRy0EPdyj+lyNTCWZQYX7hCTA4p4LA8eGXMHYJNYCJYJzr/hPmX0H
0ZeAoOABumwjW80FevFkEsb9GsU/gqWxnIJ4duuIKrK+4NhnC9JXUHY7Jh2u8jZV3jC6sbkQgcIU
kfLFu0tAvBBPJD60/9WAYUtlFiJ+UhLKj+dgPhiwWVA6oWVSbjOLdnEOggWPfVOJ8UoqwssAglJo
Q8JoErY6e/BIoCSuAo/wGyu0miVuAV9hwNLvYuj3Qe7e7qhaHGavEuGfhT7h1RBYJs971lKWFjhV
uOSCJqGYPSQPfY8t5Avpawut0u0pBjwRPMFkR6VhFOQkXPkrLDH/KtE2x29aDieIj2+1rYOsre4Y
v/i4Z4t+BQoMqJHxr5WDRPVbkcKAqqRVZRW4eX14vQ31b9Fn628FNeq0fhsvcLO9EBNCqqEvOXHR
qBR1/4L9uOHVvHUBxlIgoqVwzvcgNY06leY+KNloxahvU7VzQIhMlWKfuq7xtyBz4IbSaPm62hx3
rqJuAdGTvzBL/JTHE+qCCFAaHJReQ82Er146/K2myenGa0UeF8BnOOcg0tAjslSJVhboL6wrI0it
gcqSRxyvyml0upIvjk7xxoM82J22RWZthxEuvI/AUg89OZPwOMnvYK7r03RGHhyhsUHN/y/96sT6
57EboPFldIxiVi+8MMLube/pZ5G9TNNXdhndHm7CysvfTsK7PHm8dG3ahkXMBBL/zcUuZoC7ebR6
X6Xy/M2AWUeeHt98Koh4/kM7uUcODWr4ePzu3zCT8yrWaPsmIwqZjM3RuwY/RzpesBFStEReUpCo
s8NqzQ/MLbUu8WbSvlVNpgq/oWhgV006yepgiQBzs4/zQj1rHy855zkzMOYRihrageY9q4GehvNP
aeHUHzgWCZTn/v+4RiH0belddBmvrC9J/Xo6EMz760k4/TVJ81uDCTlV/lhua2jqLV3mKyQTIjcD
iyHwYR9BXaAYbqjAns6fwRGJw9jl0GdzgEzT2mSXj+D5uathlIuMkHNTiBUipNTrnQLrkG/euBe+
Ox/iFhXfi0i/hB0gk7w9xZmAFMpi1NCdwhYSuyd0spauFxI6xx8mlJC1KJNT2BZbC2uN6ZBDV/OL
NKzSMmpL1KV7dxDuHLW6cYvG9Pn/+vTBS60PoetQ49GTTrkz2svbU/8ZsmXH38ucR12Om0YTdYaK
SwFhxskWdlardwWA5p8fT5lrOWcNE+S9vWqlAf/StO+E7asNf6N08RC9S9iDDosyEvMHmHpaXJMq
RYg8VBw+5scsmwydZap2C7tsmzhhwuCvKuYPB/L2pSsAfzOVo9Jdgsco7z4y8uO5EsaAfuXRFdlV
c4Vz5o875MJ4y7YfDU2xWgvMwW1X6g/uFS8M7rXBGfXEwjTcHLIKW31Yw4T+MQVXRNk8LCvY/vQ9
kinFnrY1w+GAXjUJnk26eg/+CGx8aqTRKqZGhc/JqeX+3W1y59eaXN8NOSDZrqgmFfw5GaB/4vyv
tVompFaG6VytCW1AAJo03473AwA7Tf9BAVcBA0/8VyKYFinPZF0hVktplZrbQNZb1ed7Aga1hZw4
odjWMOm29d/vfwad+c5glK+0ns/DTdcApoRFrNiDPoR2XHJTBBwPpf9qt+DFgWGNucBB3V4sZuvy
ywrmtHUKOeSAmf/wtNS1qPGgzCsHXxdd9oblrRUorSpVCJsn0ypr2nHcjC7AdImqGNkswpr84Bhe
8zba0UcGCOslG0fvogfv4Sn7XPI7IMbgf7389hmito+S4vu6scT97XNYDhcYCuEJafcyWYQqsrFP
v5CnfpCRpNao7Uzzp3zNOUx2yIi2uHcikCjJID77qoRebz4cApKR0xIiAWaIWgF75Hk+pYi1n7bJ
EQgYLa0aP3iz0lMYTSDN0k90a2a0dw9LqxJxHqc2Jf0n0tTZJ1I2fmSxake832LKjDo4WLZL+1O2
V+fg6Ej2nKFvyl27MC6Z4uMSS7lQdj2o2mbXBVxM2HUGFIbmYD8LmR7Wb1T2ukjupNslU9oQ40nj
fEdj11Xun0jiVF9ejkkUISiRt53Qh05pyjp6MxV3EY5q5n6sL3lgTgxaB6tfS4Ye0pBwvAkWUb8/
30jdeRCCM654bfRmox8LgHtfZ+Y89D9t60FMWy3N2N0XtlPgditWjJ6Ufl4JyprCEweHHnHZednN
uBtNx3LWNsZn2ixdFJhQFYU61Mpm/Y4xYsXZKVTeasPrs9lgBS/hVH7ZiVlhiqAqmkJwiJUU9JF1
3wWALgYIoJLkTJTH07kLmnGwQ4rCvopJw1peTlrbO5Qv9bzMBuFuEpM6mYd+lnPLClLo5lb6ATqi
qw0DGOBKWHrvr7+kCRnc8FkOYLsebGKFb8zhCLnjBWk0xVyHu0Mt0P++D5zG3NC1t6Skblbn7j0E
h9RNQRhLFKzoPa78v+imJaswUb/uLcUsiWcyl0iPqk4/sFP5gC5lo1dq5LJYm4hbZgGNNhwA1+1f
z12Tw5RY5DBmQP3lzaCxa8oT75ClW9tye+gQ/hgEFV+WF/+2C2dd/P5T5T5NYgZ+vo3OyKS5rvFv
M/oXuqimvdJkjglItGHDS1Q2m16wCGd3cc+9V27p0dbLIjQMPRD/zXpNyj9V3mKj0q9JANPoFazN
yqiO9sm28Is/tzaGEhhDBgPG83YnAgxIVOzrgjpqVPbkS5K1LwEmZHTbHpd7CjB9Pyaqse4ablek
S74Rsfhz9hDbz1SzFIeBzX0V4BNnyCnTtb0XLMs+Tl6NniRxWrg7bab09qvnLvi7rfUgl4wVrTYM
PmCotUvcfQF2M1kcel7Bjur8ivOv3tkJ3O0lmsTIUtbie5RcOwLsawUYuiaY/tGyR5icsqCagXCb
vork9XnbHoFI8W6o1QpmZ7RNNG+7k3L9VFiJc4WTaldDF7ulStRfG552o1PRXzNX7s4MHio43iVw
ZAcn1fZ+quPLvpdqs6AOe4R7KRCV/lz44C8878ZSaB+vhH0UbYpXHvtIw0v1MdiGEG65DK54ESDm
2+6EmrSStqUVMvA18d1mZHWaSPzIwwX6TJR6i5Fb98DJlylj0CrJmZaOplj1TxDT+IIhGSaSAnt5
kg2Qw47RTemtUbNyY26wN+EW1zTQ6Kek52DDfqss1i3TBYI4FW/9ggpT0i/2KRjt+Jfl6owPD37b
B8uCS/3eA0rPrf4W1ACFkceS0DUGXR5oEJ4/TgPVRfBZNwrEylNdDi1Pi67MpM78OnXHQYK31xR8
4l0Iat2bCY7y/j8D27pz8LqXk30ewgfwALOPPFyWWnlDTqM7kTHz7EHEcJzE0uJbikab9sBLJHTX
LpUw8E+4tInogknfc/LyOo3iypEaziI5gwhF1LQvASyoTnKaJxSUs8aTww1Qg+K4ZqpE6hKP//+D
J957RHwq3PT+45d2Rm32fB/9qtA7q1b3f3juRZpz6xqwVzLD2yoy2ewz74Sv0ylj91v5SzTxeucK
GX3bgAe5piN8Zt4yr9SycnmLLVVQCoIFg7GUp2LmCPb5O2mNg45fZoTEXi4mJyuIOL6D1Az0YVtU
dfMLKuawuMSDdTv2Wh543G1aQInROFLf01gTAo0a+C7+BwPOlZTER5SnNiTqK/bC4PfGHAtTGWnB
pqjXT8A9nvV8YiwRcq3XxFDhJT7+UoNTDx7uskYP6kUMWQrahjkBc25i5L/4QWOpQMZqT9jpBMLp
S9yQBzSgKmKrRzwu1lqDzgGbujlWAgXxz65ufX/k1f/Js7ibOSvSZjHqBcxR8f4YUCE9I/Zh2GaH
kkcIL3BxKfQmIQRkw61s7zZSss+f0uIUlTeSvP+uPwbFG4R4BIm32Ri8UuvES2exeRsuDBeOlpeO
beRp0A6YPWeFUrAht8iOHe6c4WfAlI3RojWl69Glu1RI2aojEpGAMebydEypNFWrxxosJVprcspU
2HA8BR5RAP3dLKRvWL+uU9GckeIdTXWGv+aNGqZ6Fxwcjy9+cD8Gcxz5gdSGQRTIduNLRIqmXXug
QMXtjPDOrASb4j7k/wU/tgOKKGDLBsJ0LgvuclKXcqpf66rWmtdSfALz93gHL5/Q5Gecel4v8nUh
16Veq854c7KaaMChNtoOEj21OlG1Bg38QLuHPXiMO/FA//u8y6GN4ijXRD6PDXWdBy0cHkKBq+Ml
QNdEOeovsXNS1F/GOHXriAQEEF1Pjq8xTeP5i6GUubdIKZ0If4/XElgW/CsVhcfVBl6UTEEeXR4U
rKwcYZsH4Ge7186wXSL72dzZjxG17I2WEV7mm9hJgwT07UGVF6jRvWGAVFsBxsLlK2rmxOqb471q
t9sV+td+py4ckMVUoM1oc+Cwyss/qMo9IYLaK7RquI/s1VvuM5QyQ1jzSn6fxJMF+yUmxTvqBVas
my/Qi5aygE2iJIny3CuqpFfYBjLwIebPZ/jKenPw8w4/mr1Al90KQHjrOV3bl1ORBNxnU3ZmkicQ
AeKvyjDcB4HhMLtWw2DgmTSNMP4uV2DvAWXnEXFN1+NguzXntKkAAVoQ+6l8Ispp89ePQ1YkANJC
xN15JH15GDc7zbF6QzfJ8EAvCI0NJ2IA8VF7y8xLocjfy6kPMaxXuyZjWasQb3oVn+clJwcPsebv
k14JGNoAcotqKNLUHjDcHe570TGmUfeiLEsodTyFsvI1nu0VICTXyzd0vl4/qnPLVT29O0nLPgmR
CQRHLQ5S9TJUkm36QpxL2ZN98SBI+NqydLh2tbPUfVrJ2Nut5vqn/jE8VYASQjizeI7/O7tsLMbq
CkNmYw3pk9nZgixbirKitYBcDqyf+6LX3ZpGOIvJgezJJh8LOVPT5F5UEoJ2Y1rtN8ChdTwg7X5t
qZSaKRZYUZrSLGPpT5dvhpHOFk56Sz5/pjCeunxqQ56pPNMleKQMyPbXKuv0JXMLdNiyp1X1EKoc
nwSpGGwii8XnzX6PBO1crlWIez85JXGGfYsgA1QxlEsacuzNfkZ2XaXHKUej1bRpbcnCm4F5E+IH
kiGfU+H/vKsrekJcVAVxjggs0n5CvhAigiJewlylm5swERLs70xMdGImhKr9m1zuNy6Sxseq0LSq
ctAHffvBNDuqKUnTZyZus3JZmwAh+JGzasgT7kyKieKasSaV5bGMeeSXQ5yz7+BP3bI6KS3Mp+kA
xa7wSUB0C2TwuFJfClO+h2RM0bDiLi91PVabmeEffk5PYUsWepQd2E6S1pE+ZWYpCrwzdhbaDn0F
qCKQjw6i1QoA4wL473bCDdJ9RjephJUWxkVRSpjt/Wa5uNJa0F4d45m8Qj8hu0V1MWvlqcF0IQfI
C7BPsvBQ+5nsm4S5n14rK4KGo8JgRSXDzpMxAU/6zsEuVyEUhf0MtY7PyxTPooThOpYP01RQ8HDr
9LfOdKm8yU07mtxx9vS8PJk9JJjlIYmDQKV/t8DjLC/Q5whUUwbXsTQ6QqJA4HYj6AKH3Tb6gf0y
4o/uWImN+Pcolmo0SJckxh0tUY4Son1CkOWIxxkTs30ghjeGQslkYP44W1U6qvbl1Hifue9FwDvo
tQ8WI8a07fa+/GG2aIMglnXMrdPO97PyssXs/Xt9/VKMaQBzGXcABLuX2vZdQ3/x3kLmqcmFZa8n
OIUIj67fSP+IMVVdEI5WGNEvWKYlHFxII3/tEzp4K39aeEnuxWnFKNSqVpxXH0hohKfXXEBTv0Zs
wHyog/Wg+eoy3SlR1nTpV4m6o/1E8nr1knAV2fQk0DSSaW9RjfFDVwqvVT1F8zTWP1DGelIKuu2e
Z/pEOiJwS3oH5Rp5IxwPNSrry7ZuI5yto1N74F/lrygRK6kqvhiMgCxrtsRl1qpeulfOF6jrspDz
8146us+q70blW3QWNvfSWZInevsbzmn8/qtpvLSRcBiUM6YiHzpPWkowvPoR74mHe6WBElBB4gsG
Z31TMSEiTFQirxBmDUa9XccleRn2HENfp3p+kAgQLs3x7q9rwUGHXNZw3CcsZkLQYRlZhpOsZgPi
/R/dQXZK0723hK98t6wP/R6EDhtFPkq2GWNRDpd7VRtRye7PymnwjXFnc/nsSGccUS+2/CoPB3gN
GgILUhqoS/aYSbCHkHRUniRnRCOfvQklGHOV0S0hKcnFUClpCGcSXlPbfpBYTN0USCcXuINcQOAR
EUMwNWoBJZv2XvrUyiQSd43MyGaw9A3EfNSl/inLXuAbZOVoWagWoaEJ9pdQcvHsvMg1KlclId+V
xtgqjbhRNrBBiEzNmaGGuYIxkPpWP91qY1GCS1yuW+Rwxoa0WE7jBMgu+kMSn5JoMfAynDKwkliq
kUzFWQqp/WmUXLx+Za09YwsXQOJD8mKxmTw5oHusMh9j/suGer7yYgr1v4nvHvoEvx5lbefGgHi6
ixT7FMJExAEDxLMc7H1YMlZ9sr5feCr1PZrASj57ss5KNC0neJKOV5t9qS4Muq9/uQxSr6JlZXWt
bV3s3sKNHb4HGLcygwOYCJGuxViIg0+vNYkeA3eTsc1vrr0DZNo4w2a5YiAXuJUXnVQjycuDUXik
42wHD+Io7ln68tviiErR3vw2JrVXHOxM5XgO44FPjBo13ENWjOT5GmMiG/fyUHHMuRZ9/7GedPjV
rvvazjrx+5KHmet7GNZKkujcbTWrdgSFmVcFlve1U3hbzdOViyj/+NIWJId5Ctx+WuFHWxIboQjj
P9UYHRrGKjjjZyMFZBZoBYA2Yv4AZH9KI/lLnf8MVShuzubhouY+AzcVkXwFBI0GUTPV3y47XGpV
Ok1QVYUzDa5syorkuCNPs5E7eCzK6YIViRSuO29CvBhKTgP8Nvj2FCRQMcrB8shPHY55RlO114Ag
IEdtugYJgtqT1XL9pIbT6+p2KBCBc9b00h+mnZZ0pUkbxQqA3Gh+hV6sI8XPkUpieiwoyOT0yIxv
JYHZQfrfD3fQ6MoNUF5UADuZ/M6Hj2b22PMO1uBeRm6H8ruTyoa5R4K3P2KvWcuvSU/IPt/JBPQ8
J510+fziUnXrsbEdjiWOmqaWoO7XMkpk5+DPo3FOymAOz5Q3GrjB7skJzvmCnKDwafxy2JT3KHhV
0Qb4pK3yRQxZv8tHMZ+2HoUzoKWhKkrGQ9pOMd+kaBZ8lvQqHN+Db8XK4tWwflIZPE2y1PyvqpXJ
z7Kw0z8EbQk2jDZ/pD4nq9kKjGJ7c1qc3wupNcGCxoB5sIqiCb4/iGQD6VJbHM3gwk6u+cC5671n
wgQpiTTAuqMVkJWjvyiS/W+vK8QsnExigGnmaV3jKYna610ayKwVdRrFEZMR0dtdFrbxHGkEsBiL
xvo5W30I8LkmW+V2Yrnei+ll1PuFZLhiIFaZ+lg7VEU/fPOSYL/3w1vaNrwJJXJ7OyP4NBRgf3lK
6VT0AFsCaz1/Ip9MGuNlyEO4AFwaGKKZPO1BAFgw46YXj4+Zw5dBQwinBSndbxKMhSJ+eYuY6X/h
mOslu3PlBbOLYO7Tzg24aupRCFCRaGBhSsx5k8M99wBrLQXZVDVYYMMYZerO9D75xmfAkYC5h9u9
4a8bAaQWcdW9JOr2Xlf8TKoC9shncRp9Kd5dsYx+XMMY50953Jqv72wudEOwsysxzrODWDEiTI2H
jpwXUFL3BNpRseKSgZNbQkP87j6jDtkTDSk85R+OE7mUKUP9TkiRUMkkQ9qc3SUAPfgrBjN+ycaZ
izkbOqCRbm7cwdqDtT1R3Z4CNkIYWNsnKHrtFrwrF0Bf54PNyhyt/NC+6FZpak2gmFwMKIeOcenG
EJM01upW1hYQJSb/Q4WSNiZYPagiwcaBYjZCw9mKfpjMAHM9AubsND9o2OKoTCJ85VkfxEdLDExg
OMmfmV2QigFgXcgXs9swX0C8S0RVGke7v2lbU+m7RvN3E9qP1wVE45rWYhg7NRdKctzZlbuQFSmy
S/nCBUdev+MSFmS1fVbkSe8jb0xWULmrM+ZWkx23ZvgP84zmXj8wVYV0JhImSCFJH4h5XusTz/EE
kfNR9fqoLXUhSrxZ6fBwfkQegkMbqpXYJFdh8DwQjed0Xp23n8FxiRN5d0FVeX9rrCmI4BD249F3
OM/8KYjLYITC2X+u7MKDTk+bcXem/1xxQeZC7xDIQyi4SSomQXeAyC/aFK4lhK/uBj9P4uL8BZtz
Y9eyPfhhg5N5oajE+q43d1gYwQd7M1+KUmG8lk52i3N5pztqgRMeLL2+9aqMDT+7Wv9c2fvG3wfA
hrt8vzJTcafWHW2aa7/jRtbm7pp5w/1LeCbXC+D7wW3eg/bOeDkKkBvy+4x3sDvqqwzs2rXqes1Q
IKxI4Q2XALymzsxQ07dFEyMD3f/fodNnLnayKlduxhCKgPW/S1wRy0cVXnYfZ8Chtetmjj3U2SIC
VKRKWTi1O5/6J0i7ppM4mgrtjL8bOnbotgLRkWbGymn1GkVw89BYLWtlvr+5OUBG1etMPW/sYBc0
/8zkp3Cb/ZjO0VHORTwFeSUoXq/NhDHY1qQXPj+KwD4idUXIzs+CyP97IIeA8Z0EbQqEcdHyl3Xs
RGBv45KXQ+SLjYNuXLZB74YyYMBnkoY0bc3IfXEtitqinVvWPLVzTBfzXEqeNQfI3RU8PumNt/ID
1Y8SucrxFa9mNB34nmvS2SqNXoCmqURyjmefMEzTJTb+NlBh3GTn9gMtXoJGVK4mGFSzqfKaGshb
h/f7dkf4l8hshVsSGAbMIk+lfBwxwhQi2e7ygOLgGnnAc/ZtO7F+smIeJwYEnms/t9NRrLCcTFwS
PbPAHUpN9IQM47hXmklUGN8qMABuRp0zrW+O1wUomyysnlky2ZKzoKsHlCvH5VlLdi9lX4OrKWH4
nScEZ2XI79zwlO0hY475tQbdoZ5pdIWN6SfSyPLQ++5xtik2yro08c6y8ey8eoyMCq7UDfPtYc08
bT0oRy+7dUhYHRftNtWfLcdVvqQ6QOxP5e0ur67D5DlCknXcEE2mJm2SPl4CxwEBvk0qdrwyqNPz
YYgGqq060eir7Prx/dwvfo9kYqWLJIn4tpvgn0l8BGsg9QlisRfLq98e+5ve/eBGbmoYcRknOHv0
N4ZqQzNUroFLOnCXGSKHEuhJz68kU3l+Avs4lK2uRUdHRvjHnfIiJmOqCk/mSqXmnH5wgPocnxFd
Zi8S9o9qWSMns1MyVEOs2OHGf6XBMIbnYbHDZmamtbahjAi+X/6tQKK+phYxiypzTJ4EvILBVFWn
tTPXG7OXgSaJXjjV4BDfggE0IXlJNKOXmHkam1imwWPEHl231lRC5IeNE0PwrUE/jV+DM+d8U+zP
9ubmG2NQ/Z8icOg1ePfojee2x2B/GTxYUaOxeKlGhJdm88WIM/svm36byqDGA/wm12LDRdtXw0j6
9w3Cz90xqrlQb53z9aTXdUe79fPtCIUBs5NNh6MSGOniGLJBDuCzomUFWWnyWUp2sGLfKa0YwNuk
9Lt2azS+RpOQXhcuikUnDo6SpEu10kfmqvI/qn7A9wNqPSN3tJ/vs2O5v41TXvO+pVJqWesQIbav
FyCjDpy8mGP2C3ee1zwY+UKRbzHfAXmtR54ynzxNKosMrInsruus44bjbvpusxJHCw/VjQ57+JTm
JXQrLxqD7XsGQV0l8DAcH7lKyKqjHWWxGb9FTJ8wiYDJSgYpwtbUrIYrSXQUcw1Rt++ZAd5iX3X+
4LjXmVQGIrYObbzD/8RGPvl/upYvfqKaH7p/pSSD3oAM7MCb5fVxxDf8TH4Vo45PF8AHjs0vP67r
J3DKqvK8IQrU3ZCsRtpzNlCU+TUm0bmC3kTYnxo/ZeuOQvV3PAD0wpMmHlrAHL/qZi7glpFJl0+f
GiQ/kHT5nXDGESHupDth01kJ/sft53HrCwjnRSPvaRcRgOXZ1JUt8xJS6TZ/SAuQpkvbC8Im5NOA
DaNYryV4ihElRQVo+zKPRYEKoLdgqxyOq8KrbZP1tPAfVuOTcszgIFr3dszSxvIyejsxLIZD/xXX
gexOpGDYR2BsrROMKdejHceLkLH5QYvBBAF7IU1KId1RpFjhETEutcRt1JMArJ2k+v1YVrNmBLk9
CaENlqmOjfD7GVfRy7U8GV3aud/rKj3qnLwc3L3skWL80byNxLIB5T1/211HllJiLb0XdX3Ytw+Y
2VipqzPoLgnuC8wgzx7b3+Jv22sAzXHWwgkFF3ziui3st9t+Rlt6vvCYnjaAwSPJIu4P0fcx9Nn7
hbfMaQdIkqlL/nJcQOiQ9+11lN3eUbEN4AaqZi23nXUxqyvnNd3O1csQvQcUgOwNXPrmrbux41Xe
NrDqLDwdsOPgC0PtCjKtgcfV6YCdXyIwquJE6GXLijXm5kOVcamhT9dnH8kUR2u52Fl1J50tY3e/
Vt7zVssPaDikZF98tIoMJZxG2KgYel7GwskDboo+HLrgFItqysFajk5n7ShRjYJvNtDubfZZz5+D
dENeXf4scD8iHwWGAUV2DkV3tEz+lXm2MdFXmUn7PL1bgRZGJKXKwEqM+nyudl+6g+N47fTgd6oD
k3rdBBUwqQ4p+irrW8ffVStOk5gTkmwLzTGVi/imagjGdfU8MbYjGPap1ukz2/NOJY5uWDMnnarS
iyHZmXRQWTvukXY67enrQulnaHis5K6GXC6GgRXFvxDu0VxdglQFEfVu9Xm88X+yFf9329cpmizZ
MkFBvaqTL/azIDUtcCMYKtKUzNN8q5hXrEeAfukG1FZjVd/ceWo3a9aZNHoiDYIOv11tC3HOxSSu
blDNWK/2O4rQEhttgrbJC46WE5X40ygYnd5DnS3rT9j2tat5CZsc1JRD3fhNZNczXgbPh2/E9H9c
ybnQ86jmbkzy5Pq+My2tjXS0XlNCxmvsr4QrSrIS1TUewmKWUkSdN/3fDiUEa0nXN4Y+Piw9/R4f
x3oZ9Ct78d7TEUziG9zF8SkCsEKQAoIrcLYJpmys3khxdcMY8kncHaXjA/hACH5aUCh7H9HZLTDP
+AcBlIcQkA2tMN5EeCChxbJUzC+VtbvZgGXz9rpCoA/bEY4xOwXuww88khu1tnmiis5WtIa3f6vF
66vbIIHJntme113QANSjjYQx68o5YpX7lVHMx9nvxE3ndWvf9IpQY/TzRKs9Zha/VbuXHAmz5qWm
Z0NNO8NMDGIFQKzqSZaUy48aob9ILiWQ5am7sQ29t1RG4eASB6a/UqELLIKCE/S2zMs70BKYFBaf
dp7LCASnoM4FjLIRHF1s8V4tD/8X8X1+7cmiNbKiMCSO0nMmogxka343OM/6AXFJ3rFs4qb36Got
MsGiVJhZmm9jwcCt/N3yBYb0JyIvVD10qhKyhX6QCS7f7ooG/o1ti+ARi6KJ+7RNBQgThswMGgM6
gGu/GCG4XQYxU/YiLPx7NdciQ5F23D3eXTYjEPPS9ThgrEl4et4OsXvU5HIOOopnJl3vg4UG6hqr
Gyn84oWSxjc7v73eHv9DtAmGl+ikyotMniB7DTRuw69nBxSbX4aAWdVDGN/nt2Wv0TtSVfwSoXIW
qZmsd4pyvRCKsswEckt9XM6EmZoygEQFnP0Qd/pZFmXoKPv/9n6X0iHlPDsu8fWHsmglAJyoj2Wf
CsmW/ZkGB7bUo+YK0qMDUuSGmPUSUfXrED+mHXE7dvYUv30g5qdG/IPEQi7pZPhiefmEE6GbybP7
ggclFcqMff4gLMLvXfA0rBaGekLvlcVhzgI5R7mCXq41zfyG298jfORCJ1G0Ewe7VkeJvTm7vz0u
JiDjl3xNg6GFOlPq3iggFdEGrT7jW2B5WUzUAZeBCIc/GOno2BrI7JzaSbMzta5G8ZHDSmuzG5AT
Trk6al1rZet/4I4rq6hcAqNmqM4JOqXh/Qg7mOlrkbStxyU734MSr8+D0qKNc5yeQSUrbyKz9WBm
K4RSJWBW7Urj98Zksov7CNYaW0+U+r5qN6SBOjzFmhZ50b7OPg4c9YAll1K8KmbgrclApcD8eDX9
G7Lo3X4u86NooZVWBHX2NqfVYq7wbIJfRi2S0iW/Cp1h4ruGvl5DWJiFxy9JarC03//ScMJWOiWH
FKIPZhQS2Dbu2RwMkm+vleJfaotx5KCU8+T5vNZN1+p8pMnbyOAc2wB+EkDW/TweF8jogjPe29W4
r7vjGuOFrjDk5ltTY3Rgqi5UsULbYG0d7/Kx3h4Cvxf7s7F3+h5jTAUHtqo3CVdjoqJGM+UwmGT8
j+otyjzk2wN5RcE/D/fkuzhJ9lmxoNrkgJxE8XcwnUPyPg5pLIKSxbIMbXCvTbo6fezMaF8AYrQ0
oenLuAgR8WyOc9z2l4e+2xwYm1pL2q/qy2iP70HYNwHNgfe26Qw33P3PGa69yHYhCN7tswF3VD06
ZRJImAB0PNlphdJOeT9Mv4WeAy/YaeQU98pLJA+eGQEVFSxbWAn5znG2MDlaJBhR51oGcq8sNpM6
qx+Ucwin/DVIqMLMjcGDpRVWs1RepRB+0VL5UA6OGVr3V8u8pyzxDmxdrUXdGBv/cwb+LpcZ6UaJ
y0AoVVCNtVPqSm0Lx+C44EBhw/VCy+8Ii20i5J31kkdb9KM/WtbfHiRY6d2q2jXIKuUyCVBYLZSp
PPxFXz2xcYWQYj2FGdFkPNLbhuGnlBO/BroEs83LgdABTJJqhfyqcSNzqCbgUnpvr9DPmWSo1N6I
6pg/qQorFQQGTf5lJSgt2mBLpfCsNrbcvPa+j5KB3YYYF9CsTkx6Cbq9eBziObL123zNk3ZuP3Xg
Kyaveq2W0PxghyAyY/rXwncS8QZcQ134o+2pcIJFxlY87227uvx1MnBqdZqLVtgp+NPcBwqr7nLa
+ksD1ioLq6cjxDms++UYy8ISpYVzGD+SlBMRQsXtthyhcC8E7xmjkKlXYcMHLopdyQ83h2Fe6UbR
3A34wQ4L0hFWaBfLG2UfmudG1/hn4ByN72EcAsp1i99qaPiL+bqPXQ5rV4XYlAH3A9SGpbBbfb8P
rEx8+oZVbvsC8IqiwEG3WsiHxhrYb6L2M1b9yuZJ15V1n8HhvCJzl/BAN3pKTkyP6Mp+w/pwTOS6
99JG8pF05rEUT7hWhtXsSfwF3kpYlSfl5pWEvu34khr162st7vVrtYpwu0S6XPlsuK8o32jwKKwN
GMBoMypoijortjQkcTUBEwXv/5Z4UHWduEXony0whdPbGriX/TXHCJ3bv4embKN5CzloY0engteZ
Or/9EH1q+sWnWB2rjzLdtWwPbYH1aeuVqetnIR8p6gizC+TwzbiOsd5BhFYBWP17MY15HP8ozbcT
uFgffJA1JemR7+D0+EKQD7ePGQ8QbW/g7w2Ad11u95t+csxgS2Y/XORQlEjJg2GIDOG7wWkzmmOX
wyRET4+OeKyVzpeM04AAcEhJC5K6xMl5co0xoMmNoVg7Y6Suc/55MTA68UCmiy0ZicIjgIQnDG4W
f4jkrN53i96OsBY0hD8EyusCOQplyP5UM2pNKGXJ+8ZI6PgtqijIPTPSuqWKgbOAGtiWHR+PJ30Y
ZRIXVoyMXsR7j94kOU3iV7YlX0eIPaUNlt6enHbpBRyGg7axR0BZOWTk7h+VmMfM2uVBbPHbD6PL
JyOkDqj0BTjY+l5/HidahERlYJLNoxAoJTF51G2L1x+rz1YT4agMpP9xB1LDY45pGO3o4lC/YDBJ
0GXE9BJoAaX1WPSJGqA6LdM7D++5yEnhEcLgzFbHL+tctd22FPbQnZQCWQC0m/AryCkx9Qt5oNkg
oAz+pgy2exdESu9JMr8hOpl2Ccllw68L08iuJUHEcsdBddNcCXrupdgemtSbxQrU/JL8Ec5hqXYL
txsYOgA6fRP/8XdQqPj3Ypcw8RxTH4n6nuWXZf5YVLuT/btAIFrbOTFOjuUBso39drps9bWHaYVQ
oRZIsRrik0fB+wQ9s8HOSYUdJrYhFH5CdgnTRRFeD1/TsLMcl/5bd+nwYESaIoaf7ecKj8VcLB3q
jYAJ/b/A9szPgycCa+NRufBZydfmHQ5eO0z+WYN7/ovorHD8HsGVqefHVTfeoN24HZMTRtOalTxA
XwxYqtEB0u96m1qLjnjJIZdpOuF+fbMmHGN/K6piCWPMhA0wY+1K6j3IxoDtCI5kbgl41dwQdWeg
7NIjuBB7eofA2DVFYhmDGI2edrKZIkCkKklm9iImZG1IQyVE59w/arC9U7YlAGEiuoYiwsr0/jkd
NLC7xlj+E0X878adM6OXCTD5azK5rbLVetizCeY2l17vZpzy1kkFzWRbg3155iskxrfVMJMk89Wd
QzmLm1AgR/kCB830CKyoCb5xmcLg0dLuNoaW5fB/lzPzP53Q9sTfdqxvUebaK0QmRh7EGgBfy3cD
u7ugGqYEB53AEBZ5KuL7cC5bnOCDrUO0fhJjQhcWlXm4S8oO/fDFMRUTOKOZDSmlXoNW0WFMtGGA
k9yyLKFyFC3VPyqqDZryDmou39K1yZ6Xbgqixrs2QA40q5yq5tUdmdFx3MMzc50yIYDhrZK9smxl
lGt1jdZORHV/jiI4E9TKEWs12YTOQGFmu5Vr+EPQiiI8yYJFSAwxirbb+g7VpQGqiU9szmQ7ZNBj
AFSwRDn92rDU6GqDlrZa4t6NXK2irBtvhNX6HtCJG3TPsRuxNoPJllETmedpK8v4tWScJogKr/rO
kTpur4iY51EcI9qdI3kAHKJSCh7DoAGBbqLu7vu5cC3+7N29goMtAnJA1FNbZcsiGd+cltCAk4Wo
eyDBJxdKWyCmWcP+UA41SbGL9qyIci1G/Efr5DXUtrcu2Zr9P2VqkdN1cJlcAkC8UVPNNeWh7WrU
nzQZwrWRea++lzanZ2B6Y38tXz5cJYQRIUxqi3X4GRdAZ+GlxhgMqAEuwlbwlnfA5T1rcdLmpFf4
9jwU3yD2Np9eZXUGWVFe4J+rK9tBZSyP668+gOTrHe16RhWDQE5PTcrc8rBPSO0B1fChzJhcWRqP
vgnchc9Kh0Xk2KfcHRe0AQGmo8EYej1/aT9jnDqMT9q9g5AYbuKUICrbLb17d94u58P3p2YkROw6
BC7o5M4dxjVJifG2xnHYHGe/rRzcFD5Z3uN/OvQxto7LLF95BNzAqZqFzf2OYb53fmuyLgNNiODW
Dop98aSPL5stblTKA5fsR/BufGLm5feyY5lTpLQ8yE46cnqPUJl6lkgGxwqjW9EP1XmuUEUqD+GW
8Dfox60cgxwdzHBtZx3JWjgckYc4sfsjSJF1qQ87Eg8BFGV+lJ/DhDgpfduebCeLmQoY1iRljLeN
7B49xwqTa/7K94m3YCWOLXPFnXpziYENMfR0PYa0/nO+zXHcpOV/wIH4dhecE21cWwwtMApRxF4l
9NHm4kxPSYzbDxNFKileQOO4jxIx3VdalWxxtts5hgpCzcUsnhsz8h/OZdziUNNsNXTtcJ3h3zLf
zIvbyyWn6XH4wT6SMir+faqYm2fxgyXk1QqNiy8LSqm8aXDxpQXsGVBp7cDx7UJ0IrFxsiymstLT
IOPZtzjueksWEsiCGsIhvoxBkNYzF4H9LqPEji8K0XA445VY2wOFgAyBa4IvKFWStV8q3YkOgA22
HYr2qNcqg6sCCE+TgHv6AAk7R4Fn9J+LzyH8Tf5fXasNlyO9U8Dcru+mTQxDZsMrO+/U2TLpNRSk
0ZTxqgV1RHHgZMTu/obovh/+djbV7TZy+ULxlOW0EYgZA5uj0yembDkdggE8GdwSYjxRBYK2qeR7
ywZlWkGmd//MZsxfjmPVN3c8jvE7FAIxJ8YRVPh3pnsKerphVMMEs+Epb2exP5Bhl3heOO2to15z
fqTd0Yd2jPb8gVIBv343EaWzGbbZJ/2J1DKtJaMCTHt3M4tgjZT5aGlGTFdiRwm9iIKRB3TuMIpe
3WiR1wviCzKlEGDsOs59LK9faDUzAyR3fKkGiGTnUblT3kXWxckWdUVuHlO+nrZhaWVrTGdUO2de
sPFQkwyW7BkKbgir4kO3XGMqxaKwcF+cB0fPG0+Rc2CotuWEGzBBQLXy2f8bZ3Ae2IfLlR/HJXvj
+UoEopozXgYaJV6Rc04YR42owTY1sKU8qFI/InxjnyneDKQDJ4b2hrGtB76K6sq7rt+BTdHA25vd
e2OlIv8NXhqdHOw8vPi6/mMYRErlbWYYnTmS/Df55edpmIbFE3VMmto0dQhSkGvlr5S5Vg263ziU
juGa/zu6INL2JjJAp2PNf8L1cJIiNX+0ceyr+Kl/89RVvj1bgzDT2WhtEbKdkWB34SmGhdxM62L2
io7eJsgXysFUwL0C9KuDgE7lVPs2S8689EXF7luTjVOUibuxJA7FnWSYc7yE7dT5mnHwf02QpcrA
+D6yNRHF6uB9kydCBh3JJSu0Ls65MZo9sR6of81qPMat/gq1Z7vBW9wEEl0l8K1dpGpeJmHs8IHX
RcFzjqQMNP4AO/MWzd5tuTapaL1/TkhRGLOEtIPWhoLUKHvXPvJBFjHySALE/z4hJHsn0jeLtcl+
Mfae5GanPP/Yk9mepwEu3uwWrwY5SFzPlAe6Sq00sG2KEYls+pG2cjPTy90LABWeJAx7mlXZ29CZ
OMrO+S1UUxqPTmzR9u8fL87qUt+lXp7U2x9pO6hAcWq02koZ7OVNIKtDcZp4LCrh5rD0ovVZX80l
cAYIvFFtEQLGAb24UsgeBA6FJv+LoCnwJ8Z1iAk2mjHphAakRyfNV+McT3cD3j/GIjoEu3r1quGt
W6/sJRufknsxE4WO/lQnrmxC5aEA0PTWObbyq4Mbbi7pwzsXDZNutZUb+g1HyF3auO87EHGhic4Y
EztvGygC3d9bbNiO2RvaA2Wz5lRuYOXLsKlEoBIA82x/Ldrt54hn7vXsKHSBjKSrWvTiPK4myCwr
VagBqY3a2bUXZIpdK7WrVT2tqDxevKikH3rRBLSYp7QtNG7Q3UcCU6xZxmgDriv13fTgvghu2A/q
l13AjtSSX0+EVmZirf580GG2/Szrc3KjrMfUyY37AqGMHz54A9Wkgfk8WIQbp3XsyO6dJqviBQzX
b1J9sKKe/pa8m0KRl1wCQ6k09CW34sdKndQjeXvSgHuV0+5Fdkpha6TJCmauZ8PX9nyzmMdxqhGl
NGyfgBqxhXEe73HCDqgryhGgGExsi72ucBvh/PlZS40UtjY0ow/KtHbKLmX0EPuaIFP3VMsnDVsk
x648GS0dtAdnXWyt5XcH6cKzS2TdGTm9JU01g7cRYZBGfO7bkHBDPFctYgdjXAPHaJyH1KfGZyKa
FXqQxcXFwCDkQVt4IDsWkGtnLMtY+UqdT0Uczd+512EBPqTyuIYBns938PvBPU/EnaowNygvDyLp
qAfhJej2XQIGZtNy/mVmELxizryLCHXbZvfxUGscb/PMMF4KjEVeBMIFAHNIEfzFs/DoVE9a+/jt
jzLvOnKuRwvE6KPm7Xd2XO7Qym9vDuBPVpcaqW1F4Yfs4S+V6cmoF1E1vijYrwPliRirb7LKpWav
IwM3uwKIHO7IkVN6/A+v8La3XyL0qqCXhoGwLF0/Ultr9HH1FEae6CeucGJO/Ndmv/EtFQpZlCo6
rYj0uJS5ahGK2/mCXUt4+unp4rudNft2bbHhkHatcc45j82iL4a2OzSfoNaSsaGn0bA4TV1fWFoE
DOY7K1vlowlpIUNepdtOb/4vzS14ipyKVEpFrCchdPaeOn0knzVD9KBNxiWRtX49lPRHZ2iEh7YS
maPcdsZhcZcYZX+9Eod2IPtMGVDRRTXSiGReHKtPrTa7Uq5UuFp+olW68namY6BZUpmGElnc6WLa
G7EWI3ktjOR3X8fOymfhSnSQc6+C+kOh9Ir2WoFpyibgJUboGonTYnsDsXftjj7U8ZRkvpXlL1VG
5OjlWuYdeapWs1WcCfu6HFcTleoI16aFv8e+TCtZrK734zUOi8fV1n4EkM6Pk7dJMlz228L4eDA6
G+rIPqyL53Mbys/o17eS5Kz3rhFVTkB/EZBYs2dfwC/y01yYd5ejgwzo53yIdr9axd28LliaGQjS
TsfjWwoMaa0r6maX2adDytOv0B85hkomMp4layjWssWjziY/QQatJxlcDcb2ASYzU09wRBkkOT5U
/Hp14jpNWrjuozeR7jqoFiY+8hsxQBxBz+nsEZu905sjqlF9ke3UvHkWsiX1rM7I7qD3+chZhmB4
Y59RIONhfiVTo08eDwsumbUwYKtqdgdTPA7gZZSliQcFoR+Sak0gjoOuwKVIRPUhOSY5Edndj+p6
KpvbW3XaVwIDcLvF/01Jz4ND2rB5jwXTLNgNNUBb5Z36KViAG0z0TMp3Qhu0uUdDSMm70wFgk/a8
GixMEy1TzyPAodHO6MJXjBjJUwK9nU1By3ePgIyyutQro3mx5rwluSSkS4vJgsY6FwU4jJU4cjTF
9jXYSxBzkyZkGlRSn7iFp7Szab4LW6qCUyu84V2wLo8X48hYf0ltYzxoOHegS6AoSuKVxQlFE9CZ
ls0nFs13aSzjf2QyeruegKDGSkJStoCmf84JkvyQLuzC+pU8Uay8PNEvXdKiEsOLwwXg7BeXIa9D
wfIAwzUn+9HIgsK6Qf2gCqNdgOD25opvzHCAK+RydJTy5peRmT0h+dMVWgJWC/n91LwtngoLSnk1
rKSQELH767E+LQWxzjUspWd72XxJJ661XiA1Rr+lYTtAEKzXTyqH7wpC4/51VfJwIz6qUYbG6hYz
/qSYkaF1SapsTw/wtH5eIZ0+yhf/gJr/nfJGgQX6oI5o4ajiGYsydVwGoEQPheFOyNkeNCDvUTsE
VTo+5edntg8knlUJu6f7Sh9SbMGwiPcF2jqxa7slDp9rlPggbH8UkLuOgMLzn+cjeRmjTXDVWDgo
/KdvtzRLBems4ZcL9ByWV5tB9j62+mb9VYl0yzApTNSbeIFu0xgNB4vx3Fi9mUTWkLliU6ThT+cc
EOcwx/Y4j8Wvqp9z0fI3F+colXF/QoioOIo6tWT6ZZiVv6PMVJFiXSXdwb37hhFzy/GUbFaaOX58
YwUcZc5EHCQHLWafd4VO4xIXR5zPwXaUZu+clYdZqh5YJvGNbLwlFF0KFAaPjoDNv6L0jBo5v+rj
O5CElxI8vaJYA+pn6e0JiyCTpniKM1Sopa3f35k3j2UUd4tOYKjdPUYDkuqjwgQ6VCbCmoAc1OTM
U7lB9nWM4tQ7vYqfav4iU2kcxy4txl4QoLRWTIjXusg+wustxQC8haANAnY8gjav13+aKpriFj8Y
mFkgrtXu/VQxjBTfDy8AQN+a3YroD1wQANV/4zDS1AkLRCdFCCSEaOehQVwKD6U9DjegNBucYDOa
MkhB5UqegRsa+zyMDbXdUmzgWFenfg3wyEHiLp7H7iaXR3+SeIGf8Y3YCEhee5p30EBdM1D1Rn6P
s5M+cWHeGp6xIilaOij8VUz1Ux6r7khW6gIM3ZrCCjTKuyLlOw3zGq3BQlSSPwD3WsIV4q5RZkeq
a1C3A7PgkpFnauWuA1qvaFoeDnv7kqLarNHsf/MU0u+ewWN/iOUrzyVXl5TukBX+F6Jp6aNkVQsc
mWrxM95YmY0nelaapASSz0eZ4E9uFlmJTqno5Jjp7Zd4Rofj/097/QiQjDSpleeM+wGhYXDod9Qe
109wIKDf0vERDH4uscGoQ4ii3UWP9wCjB8CTUYwAQhZ7y9uEfvO6sbIkp9dwH2hwi8TOQWnj9z0H
fkw2c0XfUpNRAwF0Id7AoY6+4KW5XxqaW0K87sG7aOfDl8hlpQLFwUE3nUa3e+upAzyfUIUC/g3B
ySnq2EXJJmFGINBfTp0iMfoT4Y4YdmatPNxF67vi0PgAvp2qwYNATDsNc+A8EF4c4JnCTQLgp9iT
Ik4vkcqCdIzFNtROCTGlbfiGmZo9G8AbWn3sYEj6rruvyn9ZRGi2SAbCTIGV7mu4azCdOETVOjNJ
vB9JqvRErxve0iDmdqJbmZ/N0ofue3h41BQ2OUyDISl5Jr1H3CuDVU2XzUwFyV6AitR1wx39y6Ol
Fsrhl4ugDSTYu4YKDfdRXhtg4e+1UNtdbvqikbvIDc07wXZfxVuM0b6BXh7iQPOjhT4yFjWj3MGY
doN7vX7Tmje6gdRmz6dBQEWrKVrHoT4LbJxX3nDctpA9A39yGgLzQ950oFO+1w5MhOUAMDmntMbP
Ex20xZ7vY7dLM2sDjKpwBZbmLERao6OtAQ5DTGop1UI/xpqOpkcCEa1io/QPssiBYrKAL5GllqNQ
FOPTphJsQjGdykdA9qbWV7pdGDvGpc6QHemrcb9jdQEIS9GOoXXIINlkla0ABn5t7gTqATDh0hLl
cn2Xn31yLVOTl9Ijk81i3dZ9+vVVJd/vEalz2UrAxm6xAMEs6wNEtoyuqSihv8JoZUyuLWA9op5/
0nKKujseEGV0Nvs3EfuYkC0yhmdXgm942cIIij4//qrwn7DStDuMN8ZHCUqVyR54VmYZJ94QYOXs
8TSatr7+YYBM/kR5RUxfXR45RZdi2AhWiUXDMPqy5bpo0v/fSN8rfsrSezO2vsBGMMgJwIJDBK83
iAH7BClNpkcaC/4TvS88eM6YJTDvvSSRiCmiUt35Gkz4wZbZMzCqajgcBlIA7POBy3jKf6mawmHt
ViBOLY/ZonJnQpA9ZNHAmkT0pgU1eUbOdY/yagLa0JmpDwiEP3f4Gc2YGXxJk2WWwyXmQ3tw4+ER
aTj1b5J6UdujAmmVmKXBVD2dk4ywaqK9KdPhGB94/DbxsKBm7zbwxVU/7LdkexmXuxBdd8GMLUe6
u9ubya9DN9N10LsWhQcmQ+uGnWJphrqf0sqgnBCbbDnxBtut1BqXzP792yweMFAqZpnO4cDUz6I2
GgsG1Lax5mTteTXebtzBvj9e4eKmnXaKV7atyC2FMgrrRmiPiQvIFA1O16Hc2ia0jleoQlB9vcgv
Lb33PIpEYGYVliZZNuPhAzhEfccnsuU+XpjoCDssXevgaycL4GSRA7sXjuPrMcxRhmhTF3H9kL3Y
WAcEQMI1Qj00nxeNrmDWyBlP/E4gyCHBjRS3wD5pEWvc1kncwZoj23O4pd0B++Xgbq/5lFMe/irL
r7/bIopzJK/6MBnIpwBFdDP9RYzycZRfztGHp9RYIQbyxosPX/44Gb/OsDTx7uLANNkIc4FWtILt
AKO0q1MUwQESQYvWQsFEZanQfxE5+LabmSnAxdKKOSA5vV0kcez0Kdyi7zDtJGxx4+Kgz8dM5V77
qZ4nWiUCR2NsB2lphwDZCWMpFxu0T/hbEidDS+EO6T5M3BMH4hO1OSOrN3V54TE6o0fn5cQjyrON
KDcPCmul2qHZJkAuzpOgP2xkUsXiZokzDi0uEI8eiXdPQbvYtWRwOOm6fEoUJiWk2MxUqfJd3nMO
kHQn3JEcknwYB3IXLBHzqxOhVdjgrjS2Hngj2JI6aRBLQgowmwnuoxeCLIJ+y+SNMsYIs5k4m2Vs
+MHAxn1F3RyxGGnawx/N0i8+BUxQCRYofeM0bvmNiQdokjxCgvAuZ9lzql/xLUjylp+I3mumzTdv
RcoR/3gjl17/FqzVFyoeneo5IkSyBmZGguuzJTzs4T9MQpsvfvmdTh0tyNkHI2EEBkV//8DtZDT3
axd+vxxszw7GoBw3ZR25s1e3pI0UMO+uCyJ3kQASXx7uBxfyY5iM48a8Mx8dZvTr3lSzcnVfx2Si
WX7Nwk6qpjgPQ4/xGVNZGhLqK9YaODLjhrUfTU0SkULQnL/4S2lorsb4PvqsTll3UYAvDunQrITk
lXC6zmDjTCBhvKChlcAZBxQv6MxOmM8JN4Sa3Qjthpn14gWOdQHc3lD8LoccdMbwKsz58oIjP9ib
DLa7EshXYwIbErBHLpd2ize9BCEWGZEtAKl5EOljoKaVtoSDS0sw9uqzuVO5IrnEQZ+PlLDrzGaI
HLEpYTwTN3kLIHGsMzsDbfWEaYTyB70FEF02iEsfWJOwdHli/EFXBfQNq1fdgS9Tcd94uMUlQcHr
f+qmnQW0weXu0LJBj84TGk8E74eemrx4Yuczhhi64QzD2+dlP1oeZBjBNNYg2xclu2mb8IeNlenA
OT6oLSsEY4LjbUYVqgfjxKChrA6zGGW54NOTRqgn74AzSp062dNWpnaOC2jYL+OP9qUemeey441L
r5iO0dBwRRUF5shi0m/wtBCH/D/8fcH38X4aZGAMC8BLOmLU6RmZK4IFSNwmI0cxXTZw/x3F0gjW
IYZNGdzTVYViv/rs2B6zbOiTYziojJCde0ZcMXCvllhQCmgqs8bS0O9IFgdW6V9j7pWSrpcWxrmf
6p1EQ/Zcd/gI2NScwxk0H9YOzIz+Rd+82snYEAG9z/zK2QDRmLABVGVgetRsq3hMEPOjdx+oxMHc
6wjUMA0NIRf0JiUOi75HFW+BTnRat33aB6Y0An+a3rT5L6aPUmdXzQtGMTWc+9/6O02u0c8gDK1z
R1a5WPPaDDYL/1n1BmM+co3o/UGFJ8pKc5i3rESl++49kjvj90jHhOfMKOFaiNaxkRTG3g+rvtjG
RWQhgpsId+AMcQnFPA/hg/u8wDhJSZEeFfFpvHTOjek3/Zs+mOLTB0uGxaMj64TtFCseZeifUiBk
XS5p09j9xh6jnVtImFoHOIuTbwF0YYPwgQj5GUX2iXUtu1D6Vr36FdcLhU+NQJLzNao9Fzly3wZp
3exyBLqLkorMFq2oCAlLVEeIIVwyv8ZHfn52SVRYnEdPhTg/O8DmFVD3aIO01HYCAIYsSqrZmNPy
Mlmd7ovB/oHYs+T9s4ms5aUVsgKex7jg5+TFt7qI/wBziLzHwrlRbcWg4b5asiJMVj+ZXnBJwecj
sI/WxHnGJ7aAMQbQjwu1juk0colDb8r40x2qu2FFP2gZZ3/wk1IV3IKEqyW7CHxCyiwZv83L4yvQ
gXvugklvMZFX5Ir/XfnBRBbq0kRxof3dO+ZAe3ldcZLE6+2nzf2+2oGhvIvLm+JULAWNCe1gepyd
xlJWhpuKw3IjiGE4aDS2U7xABS7GCH+c43D6rwBAJaebeK/E/QzskSkDE3BC6zqLQcK/FNKQNrj4
9iassMZBUao01zYkRoTg/5S1wa8X46wXp55D8fo8WIyvwXWc8TzSpI/Kk89scqlswtVaMce3me1Q
Wd6zXN3vNo7oOY7X2NvRE1bf2v3VpW/QmZOdyfttvLbl2DFpE6iGE5nXZjEBl6PzFd8QlFxw/6I8
Y36WI5KgfGODUwiGrEAGpFdZktisWQUnTvn9RjdI6R3XydKmnTjmqMw/djxJxg5wspUtkyxfgju6
NesI0g0nNf55K01tUy65YgSAHxL2uvP/DJK/1LuyR0jl9/MYTBTjHX90pEGidvL5Kgc6an+je93N
LPqgzESlbPhW/59NR3O8M2m8dahVNwK8fDuYl2/3YmHfhimEYkBkwuvOIYXCxrcW1odoNSBOP3jN
OY9cAUuhSOGAasS5tcbu+AbRsymPNjjJVw+eZqIr3V1ob+g6raqQ7P05nvNqv98raqdun1dJKvOf
PALkArw6y5zM5Xw5kqlX57jV/XDJruXn1R5utKhVGlVPFMSRYV79iDyxHMjz29o0yzdpkLN4sCsi
m2Uk3e/VuWVQBugdZ+YP635Ensn+/zJjAOAB6Avc1Di9a7rKMlSjH7jxj46xDwXeQ2BbpX3ED4Y4
46H3lOmQIwEDgWp4VHTnW13hnixOsdu0/VCT1ShTmFxV+ESJmYpZ1Dfj396Mq05yC0iSZTepWrLw
8cZoNlVB/FYnheN0TE1kEA5MCu2vNa2TIIMKc+YsUffD9UMyJbbKfSU0QVKJKEVlCBHSC70zG4/6
/Q2AiViF63ftc1LLz7tclyVaWsdbITMtwjnNnh8Wydiku8m36nQwQnYd2LTEWLQ9f3Yzk+gW1Hlc
JRE7A7mBELIQHFttHVao4b5jTqHREyXccGBvfd6jEifNE8F5V33iH06GrRZ8Jv3iQWyhUy2OdWwJ
W85H6Mt95RKotrzrOgJAwsnFDkUqLOZKd1m0VCoDolDarMU09eYGkOxiQi+9DFR+6YsMwlHcvgjm
DSfV9jWtJsZnF9m9Kpzf6twim2QnQYlcAZOvI4mo/Yiv6XOR8gkEzjlvJ2UtN7wX+drLCAqkj2Vx
JVXrRxGIsG4LdyjCSxCjXyRlA8VbH3/5b8nJJ/EMC49rJS492M2/mxRtwSVXlnvofBg7Gu+meMXM
uxJzdeldM8Klbx/Tm61LapFPkxohfKF4jL634OQZ/LkN767oeR1jM7Ksr+eZpZhZJYnRsN6ztRRZ
mZ6i45GKsfcuz1A0c4IPS5ANvgEzgNhD2J9JBeZuzBadNGfacTU4ZXhyrfzkzWrNP9qdyYDAaRHx
BBVsHmDjW7a/5pIqChktGSS2j/8vDRWaUqrznwUI17fbOkEO0WEMEaIt0lHWxi+l2JvIH1LY8n5x
1kiTUcy7Bmp/3a2K5glkL2UlRXL1ZLD+X7LYw+JvyvefVbSHCZzQs8+6JHTv2ku11WhNa1qBb15f
vmnvhkWMcJwchgkcXcb8gNj/L6cZpkYTPP8VJzow80OXR4d1dws+rztVqe+53VxP0aldY/a3rMnG
1cTn0idMZty3eRxZ0CS/5CFx3G+mZypXeOtaRM7q8vl962xElmUPIh01qK+IAlCcSzrVMaDjNacb
yhpNdsTNvW0Pp1aSJqygemstqzpO0PLTPe6Vt9YX6bEdl+414Tk3+Hwaqd4E0sUpmYKuRsbwdIGk
YGoF6dWSC+egoBjgnr4s5mA5PF35u1J3pmL3esX7loUPKcVuoCXOpmPxlbhR44pWtZ3FbzdWmBUH
nOCHRSzGolKeAh0OW4ro2lZMNcKDjCx2D6Z3F4zYQqKd7IckyzgSiNedbN2OwI0udgB25yME8q0J
T71GToe0rNySc9Wo7D/HI04J8c6745x8MbQ2MeTroGJX/dWhEDLBBSff7AW/eM2ZA1gPSFnjwbm5
WMPhh5PmIk2WdPLrEmfzM51kusafSiw49LJ1z27xFt2/y0srFm19oA8TcAGGhVYmnt9PdfmqrR6u
rCo1padOTgt+/W9EZsxJcKSS25wuocF/gMjwVJeTR4vqK5PaQFX83PYxb59hhNq13jxSCjf6xaNo
a0IFuvZ7oOm+PqCohoNYG/1z7BOpfay9319cd86i3SoF/Z3OVEn+5oe6N4mbnYn8hu1soQFdYq8z
4Gf4tc6HSxHC7gmfBGgEAQ4TTqOFKPLtRsUhkRbQxj8SAZ4zW4Qv7muc5FK95RSn53PTLZqwLy1q
NHC+m826NZD8hKry/F+w6Frd2QJx1I79WaK5CcHIf+ZHugeRu0QgmB5W1BxhNTxQUJvgOMn5wZDu
WIUywSbTWuycL9STdBBE97+Sf2S6f+RrSPvEUEla2ulnUEiLduCVSbWaa1GnvwPmn8/m85BPpJ0K
owSLogyLfYpNIk4tfJgwRvOSqyeLPljib49fZRbURcJ353LE/9tApeWKtaA+sD4nWXAmLf40Ia+b
KdDEp3vQRVT8ml0HClfbC8JK5yJKvETCnHOmY4oWL/+zzlLZkj0cVPJ8TUFZx/F5JXbF6z4gn5Fm
d9RisGKDX9VInz9/IC9kL8MJbxMVLqx3R3CMWFOMvwI6QxBQ+f6LJJyzfN4cRYeemMM8BaDLTr3v
0/GMrqVnivA/W5cI8tyX2V6W6/W9NsiGRzzAdXLdJkJEnWgqt8H1WR18HDlIXCohVM+s+VDPXJDS
smibPRnS4GeJFFxXy8Up6w2UWOpaycw/ChDrilRTX0KCkAKhwVUReiw30AoCaI3daG8OQPW8/EPG
zc2ZGz2UpFcxUuxyId2zGGbpmbOlqHvKulj7U4d6o0NuUUGNi4OAJNWdMDu+zLYNbk2L9Njcbtl4
kQ6xpc9hEDlwCG1ghtVP2y+lCEpF6lBbe8t2A6iI+xP1QlnyWYQszGr+9+fcBegk5fAQtFnS5lc3
VO/v+zfFitBcRd08q8rN88mZgvKWH2kT0dskKzlfMPOeVloQDnmNqu7dWaFOW03GISDW3pk1WdNo
OeNbHKyTm6YhvFSkKBa1/Zl4u1krxQ/wv6RaZBE4rAu816tDRB+VgyP0nW9juC0EhO3L7KukwQj7
BhWNg8a+JH3/k8SgyFC3pauTL5NTRXixeYn8g5cx+DqqfykRAHdKtAcGcGSfXy4CfKcPL3a1uYhX
0NEm04TjKnzCfJ4jX3F794ck4DHwYAtfeD66dMVEucPdJX0HTC3qOBlxleTEqugKYeMAt/xEtMOP
DvUbYHMXQ1YHSexGqCLM4LIBGnEE+I84VmKl9czJW487PV4TEcD7Ve1TXvT+hXThPPm0YXfMjjC3
QI5zS9DHEy5eZau7Rya8tMk95+nf/FBwuEd5KBhL/FRO8H5O/Xi8SO16347yVIN9XmM/32BpEMw3
hRHvxKUyBKWxAidntYR7kIxeIZFo4VJbxh9cOb/3C3+jD3Mg966rRrvzwQ3TwhwDGIhYIrVPf0cA
ru1HzQjb4xnzMapatPXEYrKQK8YE4VZKu03PLMo3/Qb5MQXfUWzSv3FknuRHqTk7qkM17rCYo+R+
kzmwNd6ejqnaQgCJJBjhecbM41rhzdcfN4mhXZ34hJfNu+wpwBMdBanAvEZHMKsHOZxdXyJIIgsM
H4T7kxJiN1JXCtr2BxNtvdhPmS8Cz1WgIxv2OLKkSaK41ClXXI0OqE7o1NvYYhZSrbMrNtlOg3HD
cEsz9PPkN4bMAUF8kOK7wbvQgVwxcqtfZfvg0lRZImoIlX/TUuQeEut1HUWn2BPb95Aakacd8n30
bHxSTvDXvhOmYpRxIjUErzU9G7ygTkP2ikgh+90ufwPPrnZZA5GRN3nlYu5JTI/jrgbDZ8suCj/l
r3yHt3q5J8sFs/J6eUmFw1TdX/DSpWKq12qAcrkOe7gig5VmJSvFlQ1lTGDnB84AgJ9YuHgwLcoq
KApKxKnmSARfFyirzKVqJtBAzdPWOgkPUgFertkV9zm2+VcH3VPX/OOps8INJSel26AL7R77SNwl
K6OpJCq6A2NPhugG629orWYiSvm+MgMWtvAWjGxrDTIUfoecyAUHXfPdq/74HidWEJlPFHqHQx/z
nuE10IWxLsinPRZ9+UDH6/MtxUBNt7i0MFHlfCDX1qd8Kou/eK8fEtU7618ti9PSNZRmHw9CPPU1
IIRN7TAkqQ6vE2CVf9YzqYyAM0e935TDCLkz1DZXxZHfEDb6rPTDt00wTmNY0POv4bOC2Wu8/+S7
VtKOpuQHePpmfoCEql/0CUwGKvzgR+b78v9wpwLdpa2Nqj4BVidpd93o9FyTW2IcWR4f/U127/8u
6AzZU0Nn3gyyy15tT34sC+baFCtakscukqcJ/Nr8wfsQJGHQ/QHqcs1a1cwhaXSYMSD0pp+us3AS
GyESTCv9mAH5SnfwH7JsRIrNyd59p4M2URVpZS35dtNqv3gNVaK8NDHU1DIs9OBqjeGaw16+9MX2
kPQqVwLHh/lILY1iyK6VLo/YFB2Kp3B6q/xwJjhZVeo/3zNy0ZFGVDEqqwlkM2gbRoMVKFJutaU0
OgGM/HQFqGTnhog3IxCfSoSWxU2s7mUS9CuQEVbJTrf8ahZw0jEUffQEL2XRhmzU0poJfcrTAJ3b
UOlW2rohIQCnWDsIGLn4lEb2GH7xM7VGBYizNIZPZ4MoLSV9GHB9jrANErEj4MJVJcv45Xc0/SKh
n+ZbnIbiLwppEPLjf7L2uqawTUK4VwJdxAEsYU+CLS3yjdRinhnhn8qY3bA2RUewY3WX82FUCaSa
pwPcujY13LPyDyB1lKsui067doZIZJQfnyEI6l/BOFBpxgapE3pcZXkjWuguJhQtINZeaZoh39I3
ZIvVCDP9UEzqxvl/00HII5/spxBYa8ss+8jTzH2EP4LBuzH2I+Oq33ihQRO6snNcQIRe+s/NSjhy
jqKrSDi835J+RNuReaIgPk9jVSf8PulM+dnAgaO8M9lxUc6byh04yrPw83dXrbdjidqSoBoxFAI8
sj1c6soMxG/2iW5BSiSDQmzJ19ksf80XP3e2eWel6nYlMCJjZYUS/q5nDswOP1X1e/32Wfnj69hu
ZUA659z/T4MoJgLlATiwO+49icGUAUem/xACFSKMbBJ6jzAJantCfat5Ij7NLq0CiLsxeo6wstVc
Qx7iLw/1L0pFbgJ7hrMt0k/i5UshW628gMqsnFPPXG0YZZO+hIqd06GKWNmhptgIfzZwDKYcuOaa
/gV9j21dn6XfvRtPc8joqUz8/FhAF3Q+kacZjxgYienrcwEOUztldUf/hrLlAPQa+GmbJQTTJS6g
9nJEZ/tBjTnmHggzztWWVoxg86ljQqgk9ouutylZj2f5KlTZl1Tb86U47Y9ltKLS+VUgNqUEnD2e
YpFhiNMgHZ6UXwRlBtfvQsLRzMgUuA5p2wU0quf+yM+OCb8gILLPG2tJpPzj3k3O4yJiTaJFhpoH
R8JSj1Y/hCWrR7Q00r3szJPYNCdpx/3gTr5i57AaYuBs1nTrUfcvkZz2Yt5YWVyrGIr7q+n8blHH
fzDeCQwj5HWOda6PPp1QZ+cPQoOsz81JuHuzuyvu2u7t3UDQKYxtWOGWD/k7D6vMNWq1dDngu+es
Ao3WMMch/POZKsbo0bOvl/Toa3X0qxmDhJHrM+jQKCTttQyQLb4qRzGVPWjW2wACwxUCxDOIOzix
xzNrc+jgMowTo1b4ah7doM//86aN0QEYOvBkD8cuPKXXkL78fTW3MqG/yuKEPnLaCDP6CU8eaO9n
L4wtGOcW+6KTHmN7C7IoQyV1pvA3Bdb4g+YcIcPZNeLCzVnqgTtkZ519NHJv8KaNhzmQVe6cPmKS
dqmEcFwMkUe/yRShjcmLpwEnqHXXJ7OsRi1nx8gP8Ma5m6kRSC3itaXehdX9qTD4/eAp0ZcezG81
txYg+mrhcYgBYXvucLKGXA4hsC+HekV/5A0RZlqJ/D1vYoNmior6qiaH+4o1mMYRZVSV0ZaQ0XhI
DvRLz3FPJMMxB/JjOY4OdudTYJE5jN60iIwsRrj7QkcxPbofljz58g0Q9rPmaYAgufmoBbXWNwH3
z3CHSNJ+RYKXrpSK1nEwggDzUNtXmxNecctFZAhkG36VK+SLHuOAnrUto/x+F0fRR+ueVEvAML7L
GzaFdCy1DbUxO1Mj1c0b0sa32R18AqYAiR6Cym3PzPFAjLc5koFTN5l2CXcsre3eY/Zc4fSCqLqr
IWgO0wKwt7ZEkgw7042s3ZCbHh3V3DPRPjT6WZZQOyC1+YNr5HtpUtTUcUMVp5js14CAV9MTiLt6
ChIRoGrzftwOjwgg+vCrqSf+Un6XfeXCEPevAHKqk6022A9jjKqQPxFMwGVVsbFgkXBtra/GCUDS
wKyP82N2BquScHACSdOrvZqGSjPFYZTBrcZraADfq3+XmR9fSwXoAoZTUFfVYOzfgcExsTFjJqt1
J6M7bubL3NPLM6cCaZL+8RMrOVRV4ko1XN4Ez18KIAk+aCJQvTs31uIQ0W+yBjNyE7WNGpn58FZN
rC4kmbwyemJorGkdsR2z45yZFJJkcXbjHCkwck/VHcB4vweFaCYv51o7fg3usHv+JE2PJzrYt/my
0rfPeUQjB1TQ+Ui4rL3t8OkhFU6aVmpW/wwJK4JD3T70KuWl7t8yTRHDEt4M/TRwS3mXuehRK8cr
8j3QnL6Yfw50F4tqhz4YkEQc+ezV5+DRm6LDBDoVqB0fjoKY2NoL53uNApYhYGspuk9/0VawFVHJ
d1jrN+gwwUmsojeOW8Hx2apmeOgwhfYgfMR0DhXt41nWV4rZnL0/K7SKe3TcqkKAP6nWqtJfzoaM
hC1mOC5XQOTeydmEH39j71iFCTRLsi4aftAZPeulc/NuPVp6hI9PrMFaeEWrmC3Ojm9WC62ZIP/m
QOx6GvD7/67+x+Sd5hxllwGYo3A5+8Sx9yumwTvennkghRBc+ojbvRCl13H2DXOb5Qt/h2vwLyni
XDp+qjkkOhTlLaENmTDGoM6/86x/MdofHKToZdM/Hpusn+lByUdgHCueHlh9v2oiCewYO3vfiVXK
XM6zv4a/ML5cUZNYp1DjxvbbKGSk78l+SYY9rKpQuwTYBM+cgLAm+sFPL5OnCjhsb+L680Y82aRU
S1rZiGfy3Rjf0PWuenkHd1dwIpu5CesigHNpp0nXQS7ft8JPeS/LBCfksKKptz9Ta2SeXRwQRh7P
s0eSHAHGSL+wChGb48N4VFzaehMIiJs1X8MC0JTt+YI5dGI8cIAiiKvMoAGoMhHuhcG6pPnwL6g5
dTRJPDF5dTnqu1gvityXCz1JtuYRJxcaOpuuXIeOpbhtQJjUN6YL4weNJ+uYnOvqN7P2Zy/k3WRy
uqjMFoRWpsqUhn/LvCmbtRWjlelqmbXxb5CwXTbkgAml+QSvw/JU6BDlK0YFXHTt8ZY/pcyZm4gR
DoMdml8mDooSMYxonUGIEmlF3r7OiLqmQgXEUR3pq4okcneZe7tSudLOoJ/xIblKhndOUrH5Bi8u
XsPCR0hQ9brkjlRJMw6ACEqx1t832+QYQY/pFsDe7AJG4uy/ohoSwe1XWsL96jweRcghbS13TW+L
z0/njhP6jJLskzTRAn/puJvQYtKsShKUyVUwSaHiHpZ+XUbFBT4r0V28rvha/92IEDSqfpyqmrHD
l7yZMrw+ngFjVYvT6VJ1IRLpO3athEp29xdMLgfZU/jJa8Rzha79BBqtjpJ7oe5nCOg/B0glssSZ
pRdKcucPl2MMWwTTYuH9UnqUDMh5V2OmpnH6t36N4x0eorAENQOoZOynYIwssXoFy2C9DW9gOWBe
CCJzhUUYb/9chb1j2qc215COPfDzDcImIs9KVR1A2f5e1pagJcRHfZFhLIkdj6vsBdUcjcC8fSEK
PYEEZjnbbBIGc63r1BeVQjWpQLT5W5vLykpVp4LL2/EsM5iIzSkSQCRs9vWD5gqfVsMQbsFdKjbo
Sg/SR/UBwTcp6kP/dffrRZmDsT1RYbpGBIB4MaUA0n8S/PCcpmKEGcwkeqvR00rLbvpPGVY/aJfI
R1vmBBZzzDbzUcQNDZy5Am2AXTtvxtnEr8P3k6AvF6ilJJy6ns+MV3NFCKD6DdQF3ncjM47E0LXg
4SDGUji2X1GFPEJWIC+xTUtsdtFEHfigpDjrfa/oyhNGE7XDeFQVbxuwlB0ip/X5ET1cfmvzqQxb
IcakgPxkLdkT71Z6Rxw0I2ji7K48pLfRl11IxW8erUyQMMZd9GrpsSCcz01IxinyovF5Vhrk1pWC
eWqiLvfYz4EBHse64MBqujeXH1ri7tIZ6EdcHqgVz99ocO5esbDilyTnbeR3prwCmrxRkojPHaV1
kp50XjUH/QZ5Ov5Rx6E9c7gHzxfBtuDNju3pCZJCN4t9L9PBAtAlaJyOn1ztASB9a+9iAQCEL/L/
8q4biDDIehDBSkvzA5znJcCHi9evgZhQbda8qGgvjXe2AbV5cBthUQ7vNpDhsBI/mWWpCLxd2LO7
nkfIi1w+/DTp02Ik661XAztaSMq0DagFlAo0B6V8+l0tL6Rw1lpys3LbDsrdYKxlsCSsXJyTbqCj
i8qV+NTNOwWtOmKYFG4L6tCSduYc6340riu/LhVw1+2yTcJ8XIP3C3z4jq5onDb8jFfvzFkD5Xso
XvTATUHj/ObDGic2OJATrlNiqgqYxYMzP1020Iv47CHQF523abeFeAL6hDk+ddLcU7y7A5tE9Yxf
tKx48iHaVoWdFapfX5nYvHlgKxFTY9WXSjfMD0pctxYAaXBZDL3H7FR4xpZB8cY6dzslj3bN0HsS
AlTf1wInujeYbBRkZm0rp5YPAoVCZmgOirlmNpE/ZHL93bp2k7htJhsmO9fDfJZrbhzufb3IooIx
bGpRA9OiIujBNc/ZQuYzZTuj1SlRErU81dvVi513mWOg/n/J+X32nmpOTkNK1c/x3UMxEMNXTZl8
RJSAXje8JlMJ/AR8jPlKq0/j3UpU079a+iou2hpGZubUWKkYqCW9Qun+8trnfzzkzvbU89rQ09ij
L5mNh34TVrmxVUY1pV+6r6S3DUSFW3GvI/NPOCVnDgC8Xn/0hGpKnG7MbM667LYNSJJXLnjfbYAw
1hJ4Quxls6/8pSVLoLHMinHExYVymTb7WFjUiIEalxnGXnzCjO8/3KQHs3RNqOyyF2R8bi7iJ3QC
gglzM0VmtQ9iLD04T/R3BtA9HFOTs15fIFTIL4aj5XHFBVoI6lAUdttzuBHhbW3D5fhR2u6S8DQu
uE1Uhp12HpzyvIbFWj1NHLpYDIfEiuVBAm4Xw0EzulAmH7VmjlB1w46HRJq7T/pgYAeX3sLT/ODt
GzRmpgp2/7YZo4nkeEVvvCIybpM187Erqgp6QUXo6XnpNnTWsGTwuOLgHr92dK2N+zBcwGzoWiac
juy03Vxe63b3NMYu0m+Lkpn+0ziuOgJFHfOMF3tGAkKgSiX3B7lwIwsuFPa2LP4Y1/bkv9oGxqWG
D4yS+5L621hMVf81xyCewYDWziKFA73HNB4Vx62wlGVuTyBXEuSi+VXNfYDbAvLcYkddGCyvXI/b
1ra4Hjz+twrQuhYQkSsKQMTZttrAHzfLL9Y/GV6gscYrcYR5L8HxaufVfRslxY8CJaquy+udWDPr
JSux+64F9E+/+VTGbCX3xPlxm2Ph52/xEQMb+dHHy0ErDWM8hsDtmQybL2/k00ToOiKufCMQOPPj
ys3FUm4x3R28izSzJy5tx3ZwK2Wq2jsimV+0CPrN2QdmyUX6Q/66jSgoCrl68QSsZHNtcUZKGN7W
9s2wuh4Cl/MYJxUZbzhgd3LHQkt7BRy6WgWrKRmZLLmn8lYrwKWpp+tQ/qTklmZEk5u1ZGfb+Khf
pQm77OzUN4f2QeHWIKzMQ+PRAEgWbPYj/vGY9z9nWoxE39oRDmKg29vnb6LKKQMK/MyEbRVujTuW
xHZxaeTtgijFg2rIcslUqlf3RInGEhiphutpL7n+lWASDNo+kLb48ZrBWijFSMg2jtAZWMijhGtX
3UOsxUxIJ2HPlmOdLvUk9asVoqcfL2pAcpDEE4T9/88I0SnZ76jPSrI6E4mCsMRLWn0IPPo3wcA8
7TTSrJm7xGTeNNIQdlTEGsbLafF4fxpt1mjZ/bYGhed7Q+JUmSM6gK2lY9Juy2qCCGcakZm+pN1i
p588WWh+o8wmaWAoq3XoUYW/IRkrZ4bvL0TRm2kf0Mn3dMigjCwNG+is5ehynBcImcj/uv2KXon1
0mI9+Z+IB2rBMz+tPp3cPSlQEEkWF1wT8dOmfK4gYgbqY1JVDqMerSSQg4Hfyat1991aRB/7a/KH
pPU4WDyJtKYc+iUntaTJkQO8HTlFHrQhYdBcPjST/3mmj+KhAwdsMiz1/Gu3+F6x/Sbahe84S4kz
lwzLRwkQSkdgvZJ5u2QL6/XHbYEHV/oXcP5XN9RCZ7lNWYQzJojbQOwwLBV06guX4bdNEWx0y7Q/
lPQa4fcBLo8pWdCMNQ/z9tpIRpKm0u+Cv8c7RkK+V+sVlqm+/V/E6WgtS/9gxm/1PDfBpzLEYLlb
X7pAwwfSKxifddhWsvXsvEi4N1v0J3R6U6YIfEuoIwt88BfbWukdIepr0sTK0YGTfJpJjaA1CddX
fQ+jyIV2aDBqAVzREpO+LJyjb68hzw3wtODVe1M75EYpo5xtWUlaCdery80J6sOaJis/8A4FmoWd
ZagFBKd7CBJW3NEiLxQWB/6Kj2l07ZMrRkdlgnWUtJWGxdq5sjfGknfl4pQMshRDvMjN5EUEBh9r
QQagVEBcHE7QAlhGj3Ct+xb0wL3pq/qFqAqOhub9KU9hBudS1ghIQOuXbTrDn+iW3oovXQXj/5P2
6IDGdsuX2fNmXTtZqPCLCXUsF9b9XjbUOvWbLmWdf57Z0/tdxTn+a6fK150tW6KLr4WqWMXwdUJU
63EDEqBJRAkJBn+BkNoraOb3cUe8Kc4l5da5RyDP1V7tKXtjPy3sppZlMrTbyZ0AoaCXt5NOTIX+
VBaPRNlxnmXvNkMmHTDH59TUuwWoFykxSBhz02jVFtGqNwHCAgH5lrehxrQnQDGOCc6Eu5u8hfCn
P4P1hOaHzZjZ6OTQCM4woZ2BYLkQjZW+ATCOXsdoY/A994AcMWRBn8wh70DP6arACdwsKSx9b6ne
UbnyQTyZW2cJQGNHDYqSC8KzZx22GJGU19WUV/4VeCYwXmAz87VFwH6NcJbMmRgplnBoraCItLih
AzKiQOGiVasm7tqFzeb3RFttfj6Cio9Z5Bmv6fviYvBT1NC2r9D0Z4aP+Had/U9IbPNllr9vN52Z
FhyoLHNM6ClGQfa4m7QsoHXJf7QuQVqw+qYkn4i7RU2Nx4EghLQGtv6n6P4GerrJoZzzvS0ZpNc1
I+4OpYuMJ/PTt8DSA0CJPmYECm5v4PLfe5/QhcZHiMM+w4trMgWiTsdK7lGrbrayjQoymx3PmuVa
eRXM68VWPtxaz3uJCZmMFWRZdJIxErg9JPgXSQpy3Hb1H4tOSVJtcSgmmyBgufV/GUTxBYbpWha4
LB6jS4s/EyafJV5E+urBYW45VN57S5kBrO+3tjbDXgCBaTfDgG1ARV2/3TsCNDOyEkdUysG0sthO
DP1gkrXfy4/eclhT/81kF6uLSVDZbqRfQ0/ASdxYIDUUuNAxo2zA2qlQftcpDY6D+/nM7cn4pBCu
1sSobLiLNotXk1wTj55QMOjtCIUV36eI1B2JveQmGeEsZxeE0CX1u6JLKukgUqKTfT+4OLsUMwfH
IC4hlNKSuns3xPhathqj4jp4hDiibgyUPsT9nKq3AsKS9uiRBLZCcsy3UAIL4XpmVHwdBHfZwiGx
36M39AMybYEgQOe3JsG4lZ7HP6Y8eDdyhJUmxuHWK7vFag9ohIt5B45Sgyd1/il0m2RG1/2Ohop+
hH1i+4y7/UnihV3m9EN7lV1SwJZeQl61j1oqt+NreO7izjBc83GD+T7pAmjprqDKCW/Mtp5/NsA0
1dwlEt4+B7snIdSUG3/HuSFDrv92DEuabjEEt5cv3RCEM61C9vfa392fq9ES9Kif3hHtuC/hiQ5T
Od8Pc+xSVyqp+HIq8Jay1SdvmW+q5012627vf0sgMW/SMeBoorHyVSBqtxL6Mi4M0ddFJngkrnf5
byP6hQJnptA3MqoOQFTfx55LJyQGi5lPItxXPJjG+HOem5jsj53kr0hsU9hZbYrXBDRz4332YoaW
Dyts5kjdn/OlbzEFwuTBCk3MEljDnfVBG4u9KaI+1n5tVCoHN5x1Z2XFQDJMGflFl5QkmVICskI8
i/TFB4hz9AR3/jqvGPCyrtXZ+spRLjEUMbySPrn/IhfJekyktITxueQV8B9pdYbaEAYgkV3DT7Hf
02mUZ5VlJ7dWpTefRmAxCr/aNfekjUAbwB+R9bSvdFMhm23LUcSxQ2RiJpwMpCgPJGN77+7k6E4R
te91MbylkNrrobDibigWKgquvqke/S7xBGtGoCuHm7JdoRnF0LW1wk1QJ8lOtv1m+x3MLJURmcms
v9JDd5j8cty+m+mGeymPdcJZU8IohrjKImNpQPszxH9s+bYZAewLH8sXJaxMeW/DO7Z7JIXKusUD
rcEMtoXlOWCsEVn1XX6DTfYcdNIDwfP1RUZ9c/in3R5OLgr8zCYuBw94evIZlvam43boVUhTkzJB
9/14qWWSmDau85+ZtAqL5joHPfsT7rRs/N5XUcAW4/SnG+PvlM+lTciXx7ON6kuWy3xz9ujs4XKW
GAfnZTYuDzA93y6u1hnLLUfZCURzHL9xXB0ED5fMw7jLWO7IlUSb1FH41CYpG8GAT4j9xLnk9Ec2
WAGZ3nMJCCprGO/K8AU4/6qQfgNNjo2O4ePzT2OWu9Kv45bm3kL8YG0oOqlgO0yw+Mb2hDiX1Dj+
/bHXIqfQq7LuUFa2U9IPI6isoQ34buMl1TX6ss3j4Eg1LO9FK8JyDD8eWGULLHWgEy4rBbApz1qP
liRSnbZizHByXSkzmGFjdgGNDl6avXzZAVOooqamml4AZxJovlb2bwR7KX6Vn2C/LJp1Bbi6xiDu
FO56FDh//VNtnmGvTIWMWSJZ97dilvXopSVEoqJRKgl+QL1zBYlyFo1kHdUzy2xHdMF+m5gMBjFO
NP9jYZx6kT5FJ+y8DX18Zzf7Xng+C7xKZawbFbSxhuWjWjcarnMnDULdD0lj2PpHWzryFaNDwAv0
fsLIhr2Is2NZ7y1ag4TJnc0cJ+7iJ4lQIcDG0wEuedqhAvNeCgaw2SHga4fTk4MR4Uwu2HpsNRSW
mU6VDGq6na4Ci1N5+IRLbdAAE1A+ZsZ5+6W0EYVcfz1WL+BS37zMwDWzRO5oiyJFg0fTpPxmwLTt
vJmXng9juTHk/pxqFm4GTQ7oF9eD+axjlY6/3sFf+qJqei3sk+1S1WXi7/+39HMwHYSIhrIJf01e
ENNI4tg8ss7V0RQn7DMsfucW3N3AeHT8Uyz0JGEH3jMjT8nOD/kLqvQYAEH7hEyp8sOTZjXpUN+d
uh84Xy9/1nhOXE8r6Fm75QRYNtk+4tU3ViN8m8D+ZApdLS4E+UxoWcwc8uAFZC0wYPtjEV+7EhtQ
2i9ECZD27W1h43cqaVIBL2jAxgXiUOK/ZiYj7ZhGCszv8I2Qv+MZkJMogVbnZrOvnZRSEewN8vcd
5v991jTMtx8+9smVbNBxoGpU1oXR9C27xQc5kdX0Xdt9qrYR93rBiVWF5/GIIYTwfibid0qAxXOk
TUY98noz3cGLCpHpFJcGMF7BqWRK9dlGIZbmnggzbRkqyNFubl1N1vaUg/922JPbn5PcJP8+gpDU
WsjuhYBDEzjiVewbyoQqWA3gkQvsPNw9L/2B53A1+DGN426j7eXQv5XDMmhcr8oPv5DdhQNYbT5j
SU4PA3Hia3an5ZS4JZq08SXl7BiFVqxi8emmKEAjHitkVN7Mtav3I/j1+7yYR2unCk1o9dcKmxkp
fLd3TyfEg87kXClx+wvWrpxxwOvhhvbv7UuTxDSqgwK4o/I2yfBs4NBR4d4OWiiCd09XTbNT+jiT
qf3zAhIXHF9iobstk4DiHCpbdQ0u9PZzO3dsnIP6EtdL4o+CN7xoVU6ozc8XcV7G/mxuu/Fdf63L
MCP94trFfyTsvW4/z9Nk1wI/XEDQiwm+4tCcSYKaVts3qAVxFoJIHJqKbNueAvvyfuupClpfWbZF
0Zf8DoABQV4ZQflNVsToHfr+dbpzJZWW0GRQeg4lwwMpz50oLtPVruyeTZDDz83cNsjCN1Ol4Ss1
2lD9F7+aaAX8+Dom0aABog+iSWLiYywQ5ERqrAIiWmw4+IuAmVyk+eWa6ZFRBGPRY71htBRJnyyG
7WDVvNBGPtZhAbGS3bLlSx5zwOxZN6gfK60/UFSaLuyOXaK5XWpBwDQtC9qNHX9l1MNZTyI0W+7G
YkRr1NfwYSi1svAOzBbbyFqOJ6cvB1Pv+41jWjBotGJZvt+9o0P3XSlatlvCOl+VyA6dnqd1S8pb
ltu5N9Qh4grMBSOtKdf6Qy6Wapwzs7HNDWShvVtoiFkDne+46Kh9oSvlztgCBeC7zvxFmBS4S73g
A+2vdKcWAyVr3YP5oQb8V3O/W0jVGiWAD+Wy0o0GS6U55cN+xzoypNV+3lJ6S8DLEwhK75MWZDgt
nHx+08lA+D+tneEJFHahqPx5rZ6AL9zCKEbDsQm4SvCk0yuuQeGsBYcdqgSWlTPKfMyXTPH6uHIT
xRR82h12YYhGZkFcAWNM2F3eAufux68Imkvm0PTn0S7Dollzgznfx6vKp61gGUD8D6/WYbe/ROVW
/eVfjIhzKp1SFMOcjiz8LXLsamClTYkqlxdCnYYB+CYCTfMxIdlkTRpzewABmWcCBM3rHocCVJuZ
6rUL6jpHChO4ywNoOVuvbcBgYTTNC9CYOgvNCR9kS5dlKdj1guyYJRtB3Qge+Y6gRAbxVt5MS3fI
ufAjFVbVjcCcX3RuWjgt4OnMo8Hpe2jQn05JGSDxJc1Sdzj638iehlrtF53qDDlZHlr4zBe1Y7aP
PvusFgbTjGRfzkKQ1hsLaDLVdzWKalAdfIViyhWlaMkHaCyVYWPPtJHHVzc1ntggL4iUdsBOJP4g
MT6MRB973DeInyG1hIouKvIJK6l1mIM2FQqhP0Bc9Ks47CIwk/9EXuD9F6e0lZaslvLvEHhAmnXc
HDzx5HIVe60S+smCLoA/dxK3gmYz30CVVZIZFWzwqA2/u1xuKJlKoUkId/DfxQcRDpXzNj9BBx1G
XcnRjQycg70QHUC7/SZ/aoOdxxsYfJ7aCWDFB4G6AL4GdZ6+NPCPbv5sH+Wk3A9feXFk086Vvhpl
1RloLZKfzqJmrMUg8zbyCygIpq5YAYSeSyzu7p4xHGKySwaFT8QDTA3nnBBVNejogHtBZIRgee6f
I0VEAKHO6oECiDy3hjiUInZBuVoUNryrqFr/q+A30HwoayQ4Ok3OKnyj3vyqqUNM9B11id+GlJcW
sk/eBS692OnK+flUy1z7dZoIEX+/GgkaP4V8phFpTovQoNTTyW2ucTPfNwse3/R6ediXQi9Qgvy3
8wiQwoq2Eo402cW+eZflzkb3yEQGLOWGUfRDisJ6ZJ2HtceTvM51ybtidHBd3x3U7TWNPU6lrZny
Dcn4/ithqIivStMJlzGryOs2x2lLo8zZuQrH2AXst3gM7WrXOGPHdG2s8T1tP/ZLeRlNEvHe1akl
M7NcoLQRAIVNSng8WdgHvFLCXbM5PFdN9MDVa+KS9PHtl90a1L3QQahVRTje5oINgx/UeRhYsuCv
oEpThtYiucMIgPa6L0ZAG6X/O2sf6G+x7QaY9rLqxJOD4pgp3hlZfCnTZpwa9Sdrf5i4Yu3ty6Jh
ZDlIbFBYwa8ncFzJWLHszD+W/vLJtBTABwiyZcM8CY2QIuLk6t1CBMBbjAgtIozWFg0djYBKSywh
pj85S/t9Ld1+lLLzd/HzvMFfpdEumjs13f993ybRIasad4OihtctmZeBoxlYpZMoby5PEuuiAWE2
56q9r0663BFljTwIF8jR9zglb/5TNr6m3VAaWE2+N5G2XtI8PUDfznESlzn0ZWaPh++Yst3KoDHG
AJh63a73lyljiuoF1zpuROJjQToaH2W003psTzcFyi7WXIDTUQNnr0jverkXDYviLreT7yPoAMko
jugF/7mg+q6XDGiutE5xV6HBXwjU+YDyLNMca6AFTslBoPT1vTSMHe7+YfuovnLgI12qRQyQQkbe
DW+wk54QwAiESQmyZCEn+G88P2cxFoK4+DY0EFYsP4Q+f83BDBEXN9XacuNEOLoGJUTPWUG+dyxP
9kV4NnGj6R1n8p+rLVLNrGEsA//9U+Zg2LADMkBiwnDIJp54OVvH+EVINQtiPZjTytRaANCYj/Uk
ohgRNHMFUE179GT5M3gjHmliSgBt06YWiC5CMVRaZpNMSM/XUwc0FTvuBI+k08g/Kxdt/XBEV1Y1
Fm70Uw4pk7s/RuK1bavc2CF+wNaAadBIBkSXiFkGeFcZjGOfuAOxWiZymw6gxNUvOuJFDUAvxhLj
mf+VHCWXzLBm2QRoA2j2RMExLCvR4ytR76Egmfsh8unQifw/PIaGekGKmGBBcgQWbeD2DWxw8a/9
S1pfqkqDljRKl4pAX9JCUXno/LyCztYQ9MwlV20vftqNn0ZTIWksQcgW8e6csQxHeuJj8XmHkX04
DbwnxeIZtKMsOMe/ghSO0SZRYpY268PKF8yl/u2rSR+3RN6a9yfJiiRcmgdM2y8gH5iQ2zpST4IJ
1mg+B4KzQUgYPmGPibj9lmCJRFT6VKUcbq8VZ0AfjW4XE+wKjxmlfcN6znoD9p1q8xUj3d6QpuK3
255RZ5vfQGR+jlz2Yx4GvqKK1eGYea41DnTkHRQuIRnQyFx7LiLfZOp55Wfg1faZk9lCXwWYvXzg
PL7IKoE4tHJ/VXlJaG02vMCi9x7oER7ptz5c+K6LsySv7SL+JCLMb2zNHgrZyFyLlxa7m1oeod+E
P1H/VeZkAJqIgYvzaYQE2F1OF4F6nnwipYOCmYPwCdlEdFzs5jzj1evn3D13d5TX7jrHQSB4Uj8q
72bbyWkME/MGffqGMhKQLy8wVKQgnDDEqMHL23gYpBn8LkN/gYFfFEcqvXsbTvn1rlqsmodxAKls
1REVoKpPSv1IAh9qYQdTj9WWeX0j+JDg2qmoL1rDLn1ZrgWk8iODkQMInZCftV+8PU88VUJbdTkm
Yz8tpQxUBhUlOfWsShs3hbAACY0HsPtjcJ6e8WxF07rN1Hg1EFfjcRPjf7+2Xiy7x33NrzPL4wKm
hl1pgORQETXVQt/QPFZQi63L0hXPJMvdMtM0mCdR/TOO52cvVJv+SemNjaKJpc6pculK3aaC/fik
sy3webFgzn8OJvkwbu9TEcpQg6qXYDe66oIHIjKjj+eCPJdtCg+v06BHmKFalniUzNTELK2JRJGF
xjwP2dxT+w4sDbRWyaOmAY+VgDASiFfc46PWV/PeGl2z+X/yirbzqMJ3CL25NRMRwnkPDGJ4uAv9
2frJXUZFAQMqQLeKkH1MOC2ezlUqejUVxBP2ZNZ5pQ/oCnBTMZ2PFmB+YRO7gcXvmZZYNrt7Spro
Jmo4BHWgBAwyWme/IDmuNOB5Ii/EOeegLGZRla2yqgyrR1TJeKUkNT7e7jcBWrI+2hQqcHkoyDuV
+HH5Yddc7cz5IAgon3IpSVycEu80tSau4Gqeak1yEk+ThtDXqAxgT/7JDiL9MWXuK6x6vUa8pIuM
AbMdPQTyvW0IMtD3omPRGN03lciWHESvSvAIwBxdiHmeaKk62vnnHDq7jQgRPjs/+n73LQSyrMjP
7IzNy/5zM9RhYBPKFJtKbX2YCD2P5DOVIEOiBQtspUka70LUnZCbd7YDFFt3u7sQZSkcPCvf1nI4
JnMSxxALSBpQjEnXBERQ5bUZwCb9s2snz/rCtCY0V2F0efec2e9JF5pw/BU9XKdovBbKZGxWqWmT
CwsTADuskFKry4KBL6B6lAFbfnfzLMWgZaoTLwGJ/YsIBBr3a0v8QtLdG8chgdmmL4U1WP/MCetF
kSpragb9O3Na+6I+iKMVVn3n10yvDxdTXZalQ35V+cDdlc4pHXL2JfVVahHOZ8xfNDRuRKdFOkO8
zCWO5twga1BUg1hff8IlSpk4pjUUp4PhjdgF2KMpInD5KmoLQBuB/hWBbZ4ovvM75AV7Kl/H6sye
Viuiikeg4ZRmWyqR6k9w+75R5av1lWwgEIdzs0TFaO4wot4OzwCflf1zPTu2m+++olsPXPqcCBBm
HYOKIt53sInO+DuqwhR+ISi/8DIHhw1BTEURE8ILVNk5jcsFqY8Qp9TtYeBZ3XXK/7gpLe2PGYyT
mSJCy9Q3BJw5CMLnlbuSlhySyD6g8KWpXSkcr1tw8L3iedT+Pr7mxB5enAj9qvlzl4kW7HnjIIxq
CRkPaEj3sDVwTl1uM+t7xmC6JcUDiZGyMBASCx/Fp+kPUeuGRY8Fwu1F/RCN1kzMxwj46c06g+jR
1kzdHtZoBucTFG6ryhlCJxJv8BfHS9GFWHwIaCbkeE8EoINPWqtfq8JHTSxpRdQ44CGWPzSmuo+k
clw6kbjCwqTY7DHfLaexeDgkyY6u4eeyNh2I+5E8OIJEbGe2RGvsvMmi2wpPor5bsQa/l4o58yFl
zl454D52llwIRyGAd80D9mmvNZsjjmSYHbYHHwkjMWizf5xavLKOCUA5+hN7JmtiXoJJtVWWt6WN
8G1iAXQ/OPKbqtIxV2yTexb++fK5sNp7al8wnlpOoms4chivFyVQFOYS5qfRNEU5rd1eqqL2uDjb
W1GwHKJ6SVwfJ4ladVLH0qULXGnUdfkLwQmVxfqAJlYc5dcnCtZUceMnENFYW77s9Ia4ccY1Ejlq
2USzEUsy7AjxzRAjzRXVZckCUH4DoBmySW5aY9SDrbjd3fUK6JSW+5CPz5aeflwWydgJwRLIuI1I
a57FKEZdhF4cJympS9DJo1k5mEuP8YifoaAj1VDB6ed0MXJbk4dUswF65zsXHbb8ef1kQ+IOW0g9
Bpf/jmqSAXk+w4g5qgj2IQ0HbU0d8Q+w/G4tIE/bz7pV+RFplJRfjLgbsGu5L+8qlGcks/g37slu
Z94qAJE3VkhQ6Mf6kLfUIbeHrLK0wZ8CVLNNASaJx+1xe8VQbBSswJy4u+NIQCJjF1ZKkOX8uGHm
53G0vQJYRpJA4v8gQAKIFNxcJ7RvEPoh2bHLRrTa90C5Y7XvrB4ZTDaz8HlrS0waEYRdnwulwaLK
Y91bxg47HHpptMtVj3XwyY9ckoD+MRQTaGf0VN3BnLC99TvP2jw7fd0g4g/OSOrJPXY3ztk41mzi
QsFF4JGvjL27Hg+fPjEvb+E5hqTmvPpyhVKSTbo6/CN+z/aN1A5krnHFHMGlFcR2bbsBrA7XrjG+
QKNWwXiLUrFLFh47DgYtMHOrme5yDgb1QOVNTxUqhObdMWlaiu+hBGibFPimcqt0MVANkAQOpuP4
G/w3RBBmDC7gIixU3xBDBkILr1S4VHM/ieWxhQTAfaajCTTIXzfjW4ziqYQ5n9e4AqdZJ7bVat/M
ao57aoxxgAPWCSLC0ebr+CtitJYG7ZVrWHEKdnDJRnNsHj96aZkBCC2VemezZPHYhlKv726qogSd
5r9rflTUzDc1mhea5A49uXda9bC38jRve59Bf2BIt5nJiIXNGcg1h6OyfSOOfF2YCR67hJnFAeCZ
LzyX5zumS0NDVu4vlVNWkBC/wTT9rN5cGx4jq4MMzRovcK5xpAYm2DEz8slijJj0/xtjExwtFdQR
unbSzC3zoUDeF5tilCF+dF+5Fa9d7l2KuDI9yvOjDSOdQ0s98F8F3AQmT1VWmfaf7gFfixg/7stj
7f4min4OwSrjXrHZTk5zHs60yIWDBBZj7QWDLjJk9Bx52lZQ6TCM5d5ayX7tJpyURzjC7axIKcP0
l/yLYwvfS5HgUHlp6FR2sDFqNTlcyHOrfCI0Nrr90bGuYiV/UgZllT8zfwEI9ploQkyVhroNkZWX
muERdmPW0ibVfbZDw2P9hJ6FfJW5DUiQOPEtPU4S7KIeXxFIkSj8zbf52gioLV5hSbklxbDoRDTd
PBDtqFHP/73jRcY2ptVY5U0/OAUaV0q2daQIRzOkIRQyt83b4/9Oq9jSf85+mT1phSH1z3QCtcMU
vH0IJ7ruPbeGtriMdMc4X5d2Db98xLdPhRO67I0Is50VpgSlhVgtcfV0wUb0bpibLGV9xD9KGx8m
viYq4GoHrVfcfKCiYejduWMK2E8tdohtPknFhdDCKA/fqebOX7+ciYgRDqKSw+t2GNbn/qvC9gbk
frsTku0kGNc/fpJgX0MeV8t8wa+xJqmWKobP9MUFf+fGjnTY/rotp/kYrKnA4v2L4LHmGEylbdzd
f7Cc7y9+alrgnb0HE++lhS+nAM1ZqSdx5QgN1aY6cNxn4YoVf2jvMm3ggIr8m7i5aFlInQlG453v
d1G/CmGTs44XQ2uU2a76YQYTaKUt8qAHARZ62iAde79aMVm0yiJ9Bp+0UZqhhiUDsH9NkG6lXjlh
B4/y5vvSY67x5Ymz+vrR09ntiHxVeiTqLixSiuMaSWD7zUWcazLYktro8VA//fsAh3SFykDlk2lX
njUeT/FW1LZhpTtWU+Q8dc9kaq2DbyY/lEfr/BRQST4t0apyOFGxHqWraEKfGz3wPbiBjzORBkLv
LF8qJA79fzzXvqgU1kxnWMi1PAhxSa/WEV/yZ7uahz7uoB4Fj5nzOssylZOZkVSUREqM6+2QFhCI
LqM1mLO3Z5+gqMNrAYavQLQ3FitftSYGKiqIGKrNvwSAkn0rrzgEOmHntbUR11E4v8g5P+ocsneo
2NIUtFqcGjt1COiN4DfCtCOt2Qy5PRNT1GB1085UiwFHa4WNWCGIzTwaUhvruKJW5tGFPaDb1J2F
TgwsgERP3+Rw8mrEU69E4XPjHdZ94U01Nkbov0AtoZf+x2VD4Crlu3JlhSMUppYHj9nkTaPoAO05
BC9LEB/TOpmMQstFIaNyokMn47at70vbNhPcHJ11AXXU76Lp0okIKOa1Me26dgNdEP3bQL8p2yt4
X+OJ+Hmqe66bK6+1Kpzjf39oAwoiGLwAKMvwFWCty5VppFbDpzN/jQVp7SDh8b2YyWMfczvRL8Ld
0CWEfjEWZqePwL4uzmlwYjyOyOAbK9i/0hQOe8iOdmxLv+WlL8cjBC+A4zOVXTxvKn7eRC6gZkUg
d62uSMl6RHuFIdEszlgd0HIiB6lsBb0VV4fA/kVESbqKSz0MTK2cksikt0zpXwvO2hJYIAsdD3Wl
TloHU4JU9caogUUwdTUAEZH0COa9wgTaeU3f8k7ZQ+gbMB1hCgFRrDZd3bmm7HNiCjxQSXFMHcj0
hcAsG/YhkrqZ1iYvJANQIyPb9VMIfEHOaIxjhv6GJtdR2xzHPb3snpDCtmV1Rcq+0t5PQiEV+oWT
7VIvgYQU5kA1ZJUQ15ReqJEE5UzDjBtY/zS0taFw9VZRxbXLSSOwj0J0Os5/MJst93He7HlNn3ZJ
9LRd82Ufh5csKvA4RzoG60RyftzNUQqr3ww/qULFhGk4Of2gNevlA0jb6hilVGO6eKZJ+xzcombD
NACxmoH2yUD29uKArP/Z3t3ZU440bDGOqGuCOvIF39X3layTsZDDkrFLI2HJUsLo2yjALOzifJDK
fVPfT5O+3EqoDdznbcy92AZ/nD4AlOraL27qHb7o2WPxFdeyebVUxrJZWKFZYpNT9sfUNW65RPE7
Q4vHRFKqwG0X7MTJmvPGsaLLH+Jm4NEb6uHSvaf89dWGj7aCJWppz4NqLNaiTP67fqWDz+6SXNPa
cBYGoU7qSTBe0FaIpKprwx7L03dhctWiQ3Ko8ItP0NoEm77mb9GWmJXHsoKN12gIvG8Bw4VEo3OW
/j4Ktoc5deC3pVJQ1p6T9fzW+HFOd1OB2ExEeaWv54/JcAoaIwbI2yTjlqWH7jXbfG1I122URe7/
RUoVmqo/b+10gRDd9LsljSnIHDEzz3KupQl+xuvwkDqALMvN++0TxyY3QqtkRoSqU08gm+VtVL5O
cBGU/bztvlBUNral3Fjdj0t7EgTFV2NHHtLDxzkEJLScGeGiBroQh6FT/umgQayiQ/7j7lOLd1UX
+R2UyJX7ahVHI8BHwcl0qDrDwtWnAt2NXaKfhXLSmwTxF0xxDveQvUrAIB6bFiOkfXOllaRRKCNR
Pkw2hpdi/yyE3DH2Bi8apobkCyavr3kp7T0yr0Tw8bMj5oXv/XncKNpNnIfCsRiJzdkFRYO2o1dP
Ue+vqWet4FgJFdQqYa7NM+Xo5MyYBmQLXehIiqWE+AJn4kkxbt/TXtaDmynCo0OfoVSG6sAG+xnI
JKRAkZ053klp7tplj9buHbjcw+RCsaG6/J6Aog1gRREKin1KNnuixsSjN29hByHmRZjpaNuZl6dr
UGFEec1nMvxExf2RFrir0YvnHhmNcVodqDgBxChJs3b0MjO28nH8Bd+89VceylUQaJGcurv6l258
Eo6xB+28Dm/7Io1/euQg5sQaK5EF9xUumexvkitmNRxLem7TbfjIf3QHp7kT2/2TGCp7kTm9JXJ9
jpKy+7zsTknWy/+xeNbMToVr5lE4fAvih7KpHiXVmFiG21bC0EJQ4v2UJ2XHY7qKzAF5bERe+QjU
FyxAP+LKfA/B1lRm+/F+5Es7mvPtL4rDdFSWrdkU698RfXHGHz40T4YBoQnv5kEKB2YYwPJ+B2b8
RWFZYUDzDYMjGvLt5aZlWKcbEyM8U9pCp25IMCI1noudjBjNgu4G+gD/iW8EXgp0JJ+XCyZJDHwe
DRWGU/GlbJkU7wP0lbNDDgdFu4R4xOkIRKOqd3YKEXHSUw84jtX22FDScEBWXP+1aYqhBJtc+m7/
fkaVC1YRGduz97egvVt2liu7CJTn02fyZLlZE1e3JfGBBj+vfMU1HKqyAiIMoym0UJ9kXa0WN31W
yxlC0e75tJpD9g7eA6L5M+DBKkNQGrDg8EE6gU/YcROnK4wUcMdVYSGgKBB5PHPR56GioJ1bVZw1
IabqxYJnS2XyrvLo2PNWelui0LJ/i9GPNRitWfURMSX5/i5P3KHh/XM1OKcoiTCui3r3CEy/I5V2
zGmP+ovoRCbcnwL6DlDIk4f5DJH8/tE1GJL3F/edhU144dkSdIkdenWEw2shUs+09EtQjxne/aw4
4ofqcBghBTcI8fOlXlkGWVkFDZGhQYr0VUQNaz4X+aGtS8jN2XggDBsUfk8QN2kia54R2z9FCYz1
vI4yrlOqKbeiRZOwJDLcmjBIGqI1h5/xnwVu0VUSeYLJuLNvzFsnLhVbvqVc9dWUbBkjtSz+zcQ5
86KwEnb4dj5di4rhmrXdF3sp71WY2+pH199/dwEV2UonCjWTtl+FC26HAADSgvYfOqzqQSWuyj7F
NGn0W7ISBtV5TFxaaTPdbBWckp0XZeH1KkocYjm0cUaO90tlX+x3L6hbQXYMfLWNP7Cz0sETtopy
5Lq3V5nYcmv1l9nAAC8El34tBLqKKZNyc7DuMJo+XiA0JhRG90Ek09Pzpk2jARKIgPUU94kzQMbB
EbDzZWyGBwD2p5Xni2raYnZPHK1p2oLmM65NvE5xiJE7yDeHlTIVFwH47CAo5zIlVzf1OdKeH6+R
wQB75UfBuijwTZnTvlHJ8qV48799MbAnPC1YXNkqvyd3aAaxvOxWS/WVAWS9cwpQRtSW6Dn7iORo
emR/Dimsw9CLXB2AcMQCOtOpjuj1KBbhNQcGdzZC1QsaVdOo/amdIzitDI+wGnlJSBKpopcyT+jq
Eqs60VNAloIZCcYLKuDEaLkncahgwYhhcnADQvo3AGepo+4Pjk4tZpWtnbhGXYK2BBzIx+WAB5N1
yzqK5UYWB7TIxBUk1a3py303OyQlEX/gqrN9/K+gBi1lKnFeoraSJ/cPAbV/VEUZnGwiUXPphuuH
zm9XoRKs6/KPhkEhpco6EGxflGhub0+iMEwl46f80fqE4vmVAk/qivnbjQWF5vk1ntY4KBU4kZhQ
O8ZwWLMLLXq4AS4wpMOXUOl7Mbx39VjiBk7MWBBuSA/VKS/XpGZEHq0wSfPyjhk48JSHqi27qUdz
oa2TfDLtjkn8ItpkF/vBrK75WDvaAJU+GI0RO5s1CRky4L2SN6uwseoPskLQ1bl+Y2CQ+QbzQf8M
nt4ug8h9kwgGpPEYyEs8+2AKvhjamwOmOYjlI3MduAOZ1zmEvTm8kkFO1wu81GK1aXKOI2lprYbn
9RcUIxt2wwzNsc2LmnLGkURZO3V4RtmM1Y3Nmf2jXG01N04DZDIjzZWx/tMaZwqoQ/XMCEjv8Axz
99mCp2FnJ4caC0Pz14Uier8Bn/Uum36QR99jqrUQ+Hg4E3DSrZRuoSq26ejxL/H11A5lj9kUg0We
ZeESiKn5OWAddJUcrkLILzqwrv/1kC65awHYcHrWDQ5twVPL8O36epOQgyrwYRQTATjyEczmNlX9
qVBDSi8hcPbD0DRUgoUAhBeEwJvVQlVjzXCobpOXzt8TmdV81gtglP5AaRuzrKNYw7ryTFqD9nYF
smH1BahFicvrz+P0fL3fVeYyCaJGPyi9bx3YUsiDoDroH+E40bc6yuho6hvVWEW8XzDkkEWjnd5I
RJl2zeEZzxOXeurQ3+2a4Nr5G9A1yqWHMmF68aTqdAD/4OfiI4PZJdqmgsGaGoKhUVtBDTkfyS8S
iV8RlM0aGBEkfopbDBMGKM7dD+TkdCDZHkyvD9/DKtFTezARNF7PEp4/Bfhrn4ObEvTznvqLf/Ye
AnO9qxSEu+M72wTHBkgB/QRqMZ3dYuNpN1m0hZo70SFi1fWQDOjQWw/6EQ0hvUI+I7tAEU2b4e5/
y3MOON0/WQMK5cGwoQO4LeOe/E0SeoAk9hyDowrBy4ce5ibZ6CfFAUtEkESHn70dhcekCL3pO/AP
F3Xj0J15alSXuwIB1RAcMpGDy4ctoWIhxNQt2CatHNyRwYWhw6VbOlTGv3U5LAXEKzuD8yPGkz4b
RLpwnvT7MJwWfrnM1hbFdZ/GhxuhyYhF0rfh6KepssQ0/toDiC/MLL5RRlU6M85nEw2FAWAGpodP
DbbuYfLEmzzhZYZhvFNiNeAls3Bng4R5t5iPLr/03eHjjoDNfo0xhMyP7ALIfSQuUqUgN36GfqQt
/6/JV01nIMWItbxoU6covzld9Kgqi4A0UntRWLYzjpRgzDzJOmEWirF64pFNHo9V/vIHKMspwUIB
p7Y9mNhpnQ4F0ZnpISzS2RRg0yWuPnYxgsf6FcBpX0x3aBlkLIhgVOEYjt8ZWOXICTTfbLqFHlZG
FGulbAQaMQpmT/tfHMWh+kwmZy0E6e536nygpAwTOWmVoF6o5GRvbZONjwYXRj3+X59s3ykIqnIt
bzJRw5TOQmOp5gDQTfeL4xym96CZO5AWRYwlZZWM6uoLpv8OmSEThppMOp2dwfYxDO0ffjzT+m0d
NDEKliOaNI+vQw6ZwueeM3DrlCxxmAe+PVpxAmxWmfVtotuEuiHaLUIkB47fx6lwmKsVQgILizT1
z9Wz+UX4ol16z4snRd8k2znCnRKH1Pt4n47WmoqJjYBKLFU+mJFCrmEOb5u1XOWOB9gOLbw1mRXy
t3M5sUUt2Dy7c+GKVlP1JBaodb1/LkfbD34w7leLLzAJWO77S52iocxZ7+LDnF8OK0kKzlBqXlOb
8Oj1MLNOrDRWRdNRjEnUbzxuuf+F8FWtG4PzzfEPvpf/FqGF5wAIO30uwnb77UG8oA7l64k0lE0n
dYNDeLLjcWPnWogvxgHQegFotAQShFKfcm/WtXbts6Lkg/NGwes7nM++BiYfHHjwHGorhSl/UwTk
lKOHAeB5I9PI4ubvF71u+vGuH+AUob1AB+X7WnyGKAOHmm/vkP1AfCqgoLP8tWv7K2tDkfdL+RwZ
6Qwwmkmsvb7RhjHTBfpNeW/XewVM3qKL1W4sKIgcVysxXhv+JLuCCszULj4zhJxQSi5jT+Y+rjP/
EDodM/PTl9VynyaVyQBg9Q8rHujXHfZqSPX0uTeCKqemzCvUXIWVPeGdxUjw/f03dUCSOG8bnocK
cdqm+XFqAsmC+BER1b1bS0RYfZLV6OgSLFNIAyXk0h6cm2Z9d5JcFZCAzF5V8fe2Mm5pA8eeOsoc
kCyLPihlx79H9/z7A0D2I+KJ/9z3PX0RcqQKU5VJplSR81zW+Vhly6bz/htMVxzEmn2aHA2epPJJ
yWsI0OjVhBrtnpnviynU2Z0bWML2GZ4UFzMUwDBCSQuz4aEcP4owZKcQHHKNsGGObY/2zpLHI17a
rdijuny+nYA/5HQK4eYZcfxUUY9h4LZ8GifQtS/T+fw2Y6IdY5MTMnCUXrcREw/ZJ3Dbzq80b2DU
MtmBblGbhlLs4Mzr7nl1zV+IxRWyYYlFhN5HT1SDqNxdDYlVSiixFTtPNKEgVSnjntIRxA8mhK/c
RUVhV9mXx2JuMRDy1BTwAIZih9Ntk+Mp6oCvwtUAwUC1jbvWu6CtjLz7+yiOf7x1QWIGp7YFOXxf
jRSDez/DyqjKFVEynzoocU9/sXLwHegnYmHkLMmeQuYuQihot24gwuN9DQLTyOiF9WEneQ6DdRQw
gvr8b260BTTfk7CK0VsU4uXCdi/P6Ka05CTPQ2zBHSMZZ+cUsmEWLx5jE5XJFI4My2BBh9jfy4J8
uTQfuBWsj0+HF5sjrxmAVDR3XaSjn8G5X1kZgxE8okQwLG0GejXR5FHNzIMHr+76klZM1PbCuICA
ezjEjAZlwVIDVGJ6YnCgTDCKC44gBEQ3qqqnyuEZEL0sFWbSiEgXwP6l/n+qkeTJVbL84+pSmTW1
Zx+c1tgQpCM2kU4uWzJWh4p6SjjniSe+8xtEvAwvw/xXpLKAz+L4dvQKyt7+X+F6hKcJIyx8y/4s
WjCcKof2vreWfIha5p+uB1eI07l/GtGFRmly4cFtaujgURkq6UACBJgR+otO6Tx0I/Cc646cMdmp
J/qT/jR+QLaMzehMVbyDxGRAjuUMWSu7VldkK6hlxSzfEjHVYD8zQ69cbYpW/CRz/ijfI2tIr4jn
/aFTj1tOxaJ6kBEGbejgIJp6wv2YNbFRCx+JV3Rg7M5VYRd9SYTQYw27W9b03UaPfEjcqerFvdKR
O2IeXX+0jj+LkcxbvD+XHprO+6J8sRM0/jEp/i3ZgcGgQnGFsWv/eeTxZGV67ny2DcWCJBWJZ+om
R4g2QnNXMJeCkToLq/LY2Psex0ed9G6t/BsHGrS04RWvvXKow3imdCo49IejxkCk6jqvQbqlh1Ag
P4JDsQQRHTZvlwQJ1mdGb/9umxYQClAOK5AR57l2Wi4mWhc9jksWi9QxCr7wd20SAPebKN7A4czt
Hvb1pf8Wu9ksVAzRCdb1zS7NHDHaXR0QgbrZnYItmOhofMplrS7odWQf7yjurruCyZxXUtXh4h3H
pAsOgft1y6xTKxwWYD8IVF024nZWcMX2FgqofZ9VsHmMcHpAlhglZjdZyMxUKAwhNrnO+B9oKG1+
Xv46OkdHcsPslMCNxufkNY1os8bv73JbZs/OoSmo2WiF8nIT0Jn0tdHltsuS/Qcl62KSilBGMj+A
ARE67p329mnO/825v3Y6nEki4q7vMEWppw95g/ZqvmhMF585IbTU43LjF2j0dc+0rhCGNqQsGUw5
HidL6YXSksLS+bZtWniL3zHbRYARoOta+RRrQzMtsGBPN6c4P0TNHQnCF4H01NeLibcUHrSD26Nx
EpEjN1A73c6QEiZPB+hkYt8EZb4h4dYDcj68I5amETSu88W+dMTxKiR3jVfT1xa3+PAFZcq2q722
I9bg9rYZC42JaBI8yRxtV8OhVhAha5j3VxS2lD9HjPtoMlcf+je9bMrbgyDy6pEUyj8dyhIu1Qon
9xyvvSrhPQveovCGPxXkaNS7kJOZtDyO+o+o/lGQ/eDd+EVOUPZYphwKvPvyw/OmoOtRbKrhBpYv
3QVUKH6MhLdUHkL1mblp/LirVhdLHN7FdLoxnus+J/smsFUNm/4LL27uZHMndThhcycAdF9EBSEz
4GoKrlOCTlK+Yekilw7+TEMadsKaaMeijwlCpJuWRZ3saQFnZALvkIgOQFjvg3JEbKj2Vl8fSZPO
hNCuqSK6hf6fb/LX/BhSP+HDqm4cMI3tMfZMxuMZ3PK4NPuJsfyEa1n0GR43k4myQ1wJhc59rlw4
XVnstCiaaEA8U3pWUnf6jJmX7bmXhLSIw32hi0fPqtkUQeB7Pi4UzwCA+geHFZTssWumtpxY60NY
CZ362HF6zhhdsuVkPaYdWjdU5Y0S1R/GE6LUiBqkHEuKbR2Pgq4Lnxjka7Sk9hhajmuNncs0zWEd
BUPlclYFKDhZdvGrjfZc/A/XtmiQRVezl56ZkDy3oEI9GiDiXcp0IG9V/EDhzZ+B+YYGd219LkgA
iFeUDBBIFzN3zeP3PIlRGZ+R6LOpqRJ5CeFrL5oiVdc51CEcjHIFpJpY88iXochGFWA/owutR+lH
jMyy407koUdAi9NVf9UlWlIckNp1CZpiV9c1NrJUtXTgrsSgJxTBFB6EiJ3p4UbrprCYaLysuwLP
ay/UDBpjhoWZz4YsE+PVEOIoqi7GJTxGvpWdn5zeUk/mPSq9SlRxe7ASuev6yy3o/2G/wCyO2sI9
5Z1hY406W1c3EK81vP0C5u/8ucBp/7Q82iK2gLl+R+vahdmW8GhOOuZqG04tqLfmyYGU1FnaConm
9vySKqKjkJOUyuukkrJfIUsXgb+9GDGNiy9ugduvg/nJpQryWXEyI0GrvCc6E9p569BG+iB2vEfY
6MIcJWCUV/x3GzXqN3TE00xO/74MEjGN7y8yt18w9gPzHtT0aWUkdVoDzVFxSL1Wh4hev/4/1who
7egLebDAg/WDtj3NBmFNEd5YgPNPd3tpIy0GI6NfaVKMgkxFGwSw5vYRtmh7EP5vy6GBURu/Gd8x
l1YmGnTkgq87oJmDZbDLO5jHhh0jFRSvWvnChuu6TaWl8Yyq5wG5BVApNm3eIBPMqGBUBEJNtD0S
qXjhfxF4cfFEhQ4VnaLq0gSTyAN65ja88Lgy9G0BDtkdlRgk5fncaxz1Q60S2aDDCeirhGxf8d4u
0uAzKXVvvzQnUSoY+BPNU/JQ9GCMUKLQrlOhj8BTx5Kpr6HwsAQ6m0Fh1o9hPkMa9FFlSg3fVvg5
mOvHDd9ruT+UDrrvKXNPC18XM+RJCuTSgzzdOEIzmt3bE+1P0cjtPgbKG530LST09L67fM5wJEBL
72tZEOBmuXHKRYjg1NsSIakhC8GsxnpNaVML+oMTGQ933/r64BvF8TrTTY/7DjHolPVS7OZEayZt
TL+RzdnyP5gvOYMULe9g34bD2SfnfP+bTpx3uqCdpdNQTKeYKTAx2CJ6qUcD+T/3C7jue9AFJ/Vy
Jnn3APY790SvIEpW+CEdlfMH6SliiaEj9uACx3d4ttiELmGl6fCkTuinRQxVju+L8aaZ6sj9CmFj
8jYbzG7VCIILC7ZzG5AmSnBZumRPGjUcn0HqQKw9sgqhWT0Fx8P9edqf+qciFiIR5uB2S9SwSxBB
hnAaMI4OBJsHoGMEPUeWFLHcfU2T2/lDM91CWr2CeXkoW3uo9BX3NjRSIE26cn0hL9jKFZWvWI7y
g4Rdo/SsYRsDYw6ikuaA/4MiZSWK39EfgsdtdR97dvWfdawKk/xgvKjE9OUcKLOGXJSdgnLa4R1R
NTYQIWi7Q+iUxIFDP+yhW7GFia8KviXLbn0GJX2R0EAfCdbHb8E07QMVeFbIR8q2Tx+vSgfsv3cX
14ckXO/06tGxpS3kwpt1hqoCXPLFsrrohYC6oKsVs3BiU0d6KC7qUNLx102RAaTyCOUL4A9FpfAT
v/1xJy/di146O5gMA1PMSTH8BwKGIpd68C01Hh4IO0gri3fAVjyvNRiSbcFijbT4bvirzOHAyPIU
vTFqU97zRZtbZkRfC244odyQD/nxq/7SNHJduFmZ6JisCEkAYu874sJ3XZ4kk9gUcbi7hXgNiNEM
xMg9KhFpehbivUHmI7MVJTtvGgTMFm2TO4CFmqq6u/FQNEAXi9Q/xbAUUWI5oR/PWJEiwGaWdKiT
0qvmMzpzRrxnvaGJ0kLw9vBseqx4hAYlEIWihHhs0ImJaL4VQXFxp/ikiioZ7gCaQPuR/GFGdWWL
5m6rMijO2jAidUhxnwORB4W2FeaIrZA2JKvqNCSlkBNn5QeoeWYUc+f/8WlBI+r35OUClBqFyxN9
YZTQ6Scl7qac2yUbDK7eTqmW1aTAjwtQXdCT4UUtupusxJzxYPqTn9uKgb7Hgi5omCTUkrGYKqJr
c21YK/cleZQo3dZWJKV7aYPofrfLZIzulKfMEiIEpTX2VPrCvBa3F1doLOEmtSZq6NXu2yJZ2h44
qXKvOXuGGTn4zcGbMgsxMEa3tzXE1g7Zw6fNhLfsIPKU8mue+lEa3Tyts5D1zxx8vHgBnVo6fD+J
49AUWKbnNbRCHqtkmCsSneb7Z6g5yp8SN4TKc9mh3g6bN6mwjdnm25P1T48bktHiUbSnUPQ5X8Cd
F0jRsxV1gcNM6TyTa9O1feVVOot0ks2hbg8oTm1uvcnhqWcpbR2mSx/u1qdZ8SKjw4fMpfYz1FVI
w9P3le2oZfB27S8T9RPOuJRdQxLSeTJ69NqCOdyfYkmBKO1dwo8icdWUlOmZOAOaqQ5s0dyvoeFg
zbTDZGRcytuVEw6AvuhBrSuhLGRzTy/mhCdTi5SXgsmq8iBUL1A2G7O6+9jGLU5VIAWCcXWmIcdQ
D+G97Z+3Yeuq1Bhdhzjkd+q6Jdg6Y3Fd180D4WAndeo8aMrXYKe+aGHhwH3n7+E9fadHPfVZDNgR
DKzcTvY/AaKmZ/mqNpd/MdjUFJEnWzRjW7S72QggWtldbA+OnwRnVyScV+VPumK/ApfSBwUgKZr1
BQkcmam5ysSBiOFs6yHtuR7oSLV/mluUGIIGWHZxNNlUR6pA+acdmsrWGr3aMBItmrqfw+HgNRCI
xnl5+AEvD7MAvpgUUzCLHMsx6UO1z/m9dfSSIZDkME9uQlUq2cUdLOSG1HGjrf9XZU6BO334zg6w
Hlfr/h46wxjhq3kp017eQXdHVz/bMW9c9dhXV/18MyuUXcQcjHPnm9MBI+nMGg6pJVKLHZvnxIvP
8bcLO8FFUeHqOowBvDNdAk99TTgOn40BmTLk+J0G6q2AlIDdfsIyunrBrETUblMfnyEjtLs7fpxv
1eJ0XmXrEouTV7M7+gyAetvVWPOEly86TxQ/FDZEEncGG/bS8/D7Xc+0JPXp7nPlrSW8vJ9W3pim
WPFmtzvf+93V21obOQV5tjyX4DZilvuTHhrIuAii0tMPpKHQSkHAk1fx/e07s45+dctpppK3MzDm
1NItyZAYQu5DALh3Wupc3huxCiCgRo9gExK2y1wloOLLswKxEBk/A99OWFdtnKaBOTfySTJrV0jV
mdMqMB4RlWgKWOyEUdrtF/4rep7npa0wNFKjBL16iUDvln/OvjlL1H7N7xLmDE4pue64zdNosRbN
pZEQCJ0bHmCibdbxMIrFpJTy55uDJWxfYpAXOIBaDz8JmNlgRQ1wNmg9NVrkYCuQFrCY5Lote35Q
qIS6jLuZqR1+g+meN96SxQEpN+6ZCJ67fC10DU2niKDKxsl107H5P7v6nlRW7ehFfNOEKB0gjdBy
FphckSBnB6bbSmt8PXzt4bIGbSL80BGOVdHv7DqPIVw8xteGnKYLL6RldEg1SXYA7ypptslP9Xem
bw0ZT3VhO112st6UA6xXYMKBCwLoo/cyDLGU/SEzIOTn5lXEqReMFVeqJR9s3hU7cjDFqx+cX3D5
Y0RdpVY2QgK+2kgSQ9ISycEU1LxDwG3sj9Km/S/+A/6o5aGdQFECyXW4+L82u5DajAzeKkuzrwQa
8Prm/dhQKqckfKwmAHGkS+Eh4LeYVfJ6r2QssC4ZzTslzO0Z/Bhov40Y9s3Kd60ajOUNL6AJxoFI
f+oCUffmWGsDFsQ3kIBcAskhoGjpl0vqs/zO7Sb7W8XBDIlBJlIFPENctk7vlxFtwVpf/DrIZ5oj
JQwDuF0SbORjciiqC/Tbs5KA/+i/XqONaxzU5+MFtP+1VYsvnyhJQD3em7bYnIs85DHkdIhOKEyg
2N23jgnFzSZqZFeQ7d2YLc+pdWHrcon7w+0YOj0lWPpFdSDR3a3Zwk8zrj1J+1SSkfvZ26kKJEba
3/ROcNnODk42P0vdSWBNEhzA3S/JyloXhtbY0ihdmEf4sIpoZOoCTLYyjEc74Ss03dO/wyLn+56y
A5xMn8bY4roR3ZAs7PbykwTB2J8NztIiQI9+S0ckI4awsjajzqEDRtN58YnSP5NIs/D7BCuCZxnV
8zCkZSDXTGK0BB6wlfyfFD/g0IUotr82c4K4SJa3XKbMPAOzMJAJrQYwH+bcqSB6G1P5BclGyPAi
IBCVcXymhkViP8mh3z0aDMpeHlgkIpQjA8X4g/qjhOPMwz2sn2FwN27CqfemCHjQfe6GejS5Rfbv
1eAqDLqqBa2ovs/cAiG3gTtGlvYo41g9efOhkUurkUk9zQa/0iZSDLRS5bP+0LRLc26+Ap/JqDE0
xK1IAyG+lKrfBAHl5rKQ6eEDkQIHGzIQjB2epGB54msl0Jp4Mjeq/iMiMPxOrPmb1fcBccYS1rdJ
+t5cv/adXaNChGeKUpklwYXKxPH9i5FRvpYGCN5ZSpGncGXMHJ3KbOkNqFQ6g8H/cSL0f7nr4y6Z
8zdeM4taraXAAQvKq0XNB2dWx1EJyHku49vpjEx551lA/ONynIWFe9OjI9Xm9Og02mjXViK3yTIU
suywYkEI4ZZphsXs/8+pVwFH9Ts6aBo/+gkJWtCgPgwrzITtC5TRGVSly34rQCwY+LfopVHQOczw
XTgx1PbI8dv0JH72A5sr34mxsyJjIA0awFTpqWw6/v63+rucyUjulmPmpIvVKAb8dHi/LFR09ZV1
1dI453cCFcJu9jXTspzXnm882nAYrI9tWru5Sv59jUjHb53D8UwSYtGF35vJ59/eoq74r7UwYjhX
CTwN18EmUq5r2MUkGVluU6sEjPTEJCZnuQ7zZwcuNaVXnMh6+Z0cyUS7Xe2NHR5pKW4g5m0H7gLH
9H0lESwDmALTKkp1rSm3WskTuatl0x61jZLEMbvQxHKpdUserQQ9TE8LTitZU0uPLSDiDpIzmcGP
rlGSNhJxDEHy51I6TLe2dDcViP8lVxNS6ED5kpHs9CLXxshVsoECnZTo0VWZ3rFC9iNeCh5RaALx
mTaRiObWrAQNqbdwztvG50mHfs1y+ix/qfC7bGo+UJcoVCOOxvr4Zh2YL45G3UWtK7uEN/g64YJL
TyW3z0K8HE30gLEKrAWsu40AD48IbF1w3Dav0qVhZri3T/Grv5lyjwimX2cFYcJJt5q4TGLduuID
BP1QL1XAJ6qG+pY26Dba9gJryKH5r5XD3nWeGca3DHeY0D5zme0GZ46yOpCHjwy5PtJv6sy4cEPs
m3Epq42wNPP/DEpgagOTGcxEu7JhHSXwpVN2sNMzi5DWi7S0Q+x8oQe0QZbUd/LMXuEktFOccOfz
qjfi1ORQnNoRZNKdx2TDwTod1piO6FX6eX6o2zPMapb55Pb2jkB/oG4Cq94O3IqTO/dCJ8W4uFhA
0xtE650g/1k4uGm5Xi0V82FkczVNNTu6yAticbfXPAfvzjg8DMBXCIi7lCEYq2jVspEZZCG2snif
At7NxpBEOFOTUDTuj7rtKbjrDkYESFsO9OS2fD8AxsetxdAX2FjS2WF+/bu/cjXbVTA/CUekveGP
pP3lLUBDJz3teqHJrwT0D7krQTBqNJfzq7gnsHHwYXcYXKM36FO5Wct442ECQ7NzUnH0/z9TVrfS
mvpiFyA9VWurZNyjroIAR97Ecbqhf/I++BFDFte3LErhkZ17Yqwpzwa+chWGSKoU+8FKaKVS54ln
WO8FLq539/LJGGvrfA7apyXiBakxK6Obl5XG9C/dfAV8AVE4e0TZDdZHMiakPQwmUPmIC/Y41Aa/
yYr6+ukQC8h2pieDlBPAdJrZCnF2v+b9zfw2ul7NIY9qSixKXQX2rxsvbC7TAHnrogUBVaWuJlmN
hPa9gpP8cijT4Bxq+18QYwxhJQyJNCBVCBWNNqEV6wk2EJd2jf+4o+tM0rbQinvxZIcr3oLN6kB+
dD+QhK6vXvlWWeA3c92p0DkW7LAY5JRC+AWojmk/BIBmz+HOvXCci1OfzZQ/IwhOOLZyOfcZGtpw
azAYT1/yoyocIAzu/hG8J1AO7yXl530B0mSFeBVwAnSFtqzHNqIHreMkZ241jG+XKW+rWoAKDK0C
tLvqbDKOswLKGx1/Uh3dPVY0hPhm+jbkoc/wHfna0OsouSZ0CJ8ybu6qcg+PAeGGuO/yPUqgydlW
92XbJN6h/drNJOqJEegZpfY6D/JygRGjUSSfq1L+zEwkAjLSd74WqrXIEUFwEAxsh9rCf4xiOaSD
MVFdBjezRB5/CZBz5UtrwOHgUDom2cfvGnh3v4XpS4vXBDFm7YSGwreAjpVjDYGmiS98ZjK1e9r/
vLf81mortn2jEJxq70CcfdoYmgVCHR98pKHXfFKUAmJ+eSdJG/dH2CfkFzZ1ZLOUdojyEpZ87SUQ
5du23hEPAojj3bJ54WwxtI4BrNP/+OL/1agGpTKRqZankfzWHVVfq4PAqv3iwaYQu9oHfz/WtuAv
nFC/vxRBECBINbPrQITVZ7w9GNVJNo7PHFpDMF9uD42uT50Gv+uSU7OLabvUm8QeIVfPHpXeRSb1
iGOZFojcC+NfkM87+mtKzOJ8uwsm4qqOYdXiJKIxREq0taraObIS1b0dw3Mi5W5DDulUmiu/1XuJ
cfrVd17GJqkUn6eTaJ8m/cmjglD2OTIxiRF/0988bU1ZVhdVHX/MxyCx1uHotepHkI+oi0J3M8uq
yydv+rM4GzA4B4rdmOH1uHYp2YsMjqr63axiV2aKbvTfPmc16kheGuMBL5yQo4ELJYoasEN5wQS9
i5WbK/wm1vrUHSt3gSPWz2IYU9pYMRp4bP2Ry2YEvUn+SGlvYFJStU5Q61+4lmOBoyI4H11SPe4i
Ksp+oTFnVT+XxjO6UzF29DyxAr9/Xtf/e9w2rfDyUb0Exxnb0b9feBTuBwheEWT+/L8eLsT28hdA
dYG/xUbmht+bcKg6WiCmWECOm/zH26GAzOljyKbFkE4OVuVUgxYbdX23qjLZilsAubg1W/klf5tP
gbWLwqHKeE2dAoP3mS7yLlct+JVwRvqYRJe+/BBqhsDYwU8MV7AuUXYe8MILTL7hKPtSFxTgjcwp
jJnRe81f9luZwKQDbrOCwbWnsX+3DXN+wEEqG0G0Y0v8rVq7HDY9L/edcE3uhSRAuRIP1svycK1/
stRcK092uGtalFLLRkYL+CVCxtqlousXwN88yFWWCjf2KKnV0ZSCofQs3TM+8NZq1WbRp0ffTv1O
sjAUBMeCmPdmPpKnVkpCxV67aHX79qYPQ3/GJXJCmgjgvVOP72Xkp17w8h6vNq1IarvbLoLiuuR8
NUH59x96Vc+gnwo53tTB7o2OOuPbeYeAr6apROa8/JKejyK31tyzfvTsiIt6seWfROwsDB4mK6Is
ayNoJkc2o85ZTEO2tArwnaPH/OnCOMBixwcj5yW+GPV8ikECx3wXUjP49cgwdZq0ntfkPT+KORGp
96av3orF67MSUtnhGpwTgjd1F5yTIZHdfGYfD0veUVLtxEUSb3fyZKn84s2eIvxc/qpStyHiofwU
xlv1tK2sxmKcWMI/zylIR3N6HClljt1iM2+0kgNRbtHnXOd5mG16MZqZOwvzYDGPnGYl/lbvqM7v
gCvZGdCBo9O96PE/RoCyUQkze9PaAxL5q2KALOFdrS37np35DqtnjPag47N+keTYGwYBXTBFehal
OdEm5NJ45qmHD+WllnICXgynoGeDT3umftoDDIyjyM3Ru9gmCY55zzXstF1BbmlL5OOsMWgzHf+q
VBFN3Yap27ohK+lalfe6RjVhuxEeaRebVj+CZ/HJzEtUBjDKi8bqW/UcgbphrLRDNONttCD3zvZ9
PWn2NsQ47ME79g/rRRFqzqXkKMBUfCWg5DiI7F50r0tqME5kXamk5xfwEA7T79WU1x/VEI3r/eHL
nbpOJORu/SDugmRu1D7hjIdV/71KgUGC7x7Is27GMDfNuq4sQk1cBAZjEDtJYo6oas8ZXx/jN15M
ulvAcJy4YgUpUFMuZM42ufsY+fXzo/wPOlhYVoo9E2rQ/04DykxHOEjILOEFqhNWD1qzy8azPFt4
YrKnTy2bhFFcStSt/MBEWhI6lg5XSG8JhqdJhmX5rB7IKWxKG8pb02TzwK8i0wkxcos0EOKlE/tI
13xekRcA9AwYW9bynQpAC8Yh7S9ZYKzCRg2VhH+S5WwUDt2pwkble+YNO4ZvH/GvsGWK+WuKMWN6
WaLlqtAONo0YR7XwJ2znQynzshkyj108xT9u1uakLP2alm9ntP+XpHZsrSOaqcUgAjB490uWWqbs
ZD7umSh0PF/7cSrdwvXu+H8qUxPbDUXGT09xvmmeDle/dnv6oMkhgMYRuvW5Id4IGxoJ5VJldXHa
2vNEmrV+nN0UhknI2AcXXbOcJQylHUUpboaYFe/QdR/lu0ggFpeNEfMDrIISQLVd45JanGX3AWxe
/2/bJwp/RnuwflgGh6XLVR6ly++JtBnSM5RtMStjHUo/8fEb/CSD6bclZkB6+bQm1NrgQxpjIlq2
O0hi8aCkPPK3mKUxpaOZnohnKMz+Gb987fs0iZyEnVPaeftI0CbtAiWrkUZqDN4zlgFhl0MNWQzc
F75KJGp9/dew7onsYirv8MwOil5Dh+bFhkSxW47GI9xio6BCijo/yN/SXnXTbzXHe7DW7g55cyFj
cwc87jT71xlyAGxwewzH2+AsWfRG/xJVGBA9gk1BgHnrHl+Q7NtG3XcfmpdQT8xvHWKOlwXzuu4O
XIyRiUCX5Z09C/DEzPqVtGWhWKupgic3sEmfFcE5EprsgOLIpcAPjdGiBaVGUYTJyfeQS5rl3st6
YtRq2IZPnAgBsLQWft3+msqzhedtasqw0g0hoMnwdmfVwqsX9Nu7qV4+bjPvNDlsnjCvu26/WRPl
U1pk5966DhhN2AtmTFlY8QfJIwlOGfnOd6UH2aVzUwTq2qss36sxCG6ipUihVlogPIVbKHNWQ7qc
/6ymFclVw1MXraWkedBrasRiXd/GvUl6UqTIEK/+WuHl/njMXcjz5i1gT+Yzmj+hqoaeF6UoyLOh
+wUWSxWYM56zcLQezzhoytiXWIEUTfbpdniOyFkCF9zGoEeQYtBiN3knxn+Db80sqSEJDCUKAbJH
8yAaIf6bJtQginuXXOYM3P4kJGeev0uW1FHuggd8zfEikOj4Jat/vKXw4eW0CbSii6ZtEEXGcxXJ
SzRBMarI0dgwx7GDolz6s96wHus7cZxoksQxRdp+fE/3EVu5hIu9seSp+EWEZw731vXHnCl6QSXI
eLh8R24lBHHd+nBvhUnTiFs4EkojWr3ZSTKc2Y4Z9gnjt4feVtE/aI/TKatfC71Qhv+9D0DiKWv3
H1oH5/8l9hjLpgTjTc3l5KYGspXTbqrWvLjGno7iloyypTNGaC9sxe0PYY4HTBoqgLuiWDbACt/f
vil6vtKGSgDLEtiuwgsdCvnAEikR6v4ppyr6CfrEBaUd5Qpo+1d/mwXR232tRviYke3iZ6E/ad5I
yZCyEX/wMBen0aTUOWZ+q+a6eo6xBiznuYIeHYxZAJLjxsOwuhlCDcwrIFObov9h3un1/ghasFTj
EdoeWNDR4jqnl8yTcEuh7yOvF9W7tA+MkWK+r4bZ/7KtCkX+MOHlg33olP+pRivQVvd3nQtXaBGK
9SkzkSKLn7LemUrIfGyTRbUmL2QTfTQnocyS50cFpkkK8v0EnkAid20QjbO17KldWSwSLX7H5zca
Vpvixt4obyy9V7Bt+ZbdbN6ZuFDXhYFFYNdPAjVXNmeMxmGWM3xisGMB2kLRy0Fy1VnbRzq9w+eE
uyfsm1s9UJswYw9U1rWMj55juiDXFsGxSCUIwfNvzLdKaEuHDmxEtz+jlvaX63PsllLZiX8pex6Z
zxeW7llJ/h1ANZTE3sgiFnHl+OcXGXSW38Vsae8iDcbe66llYUNtuMfUa6FRSpd1vkIJ/B5DH3+L
bQQztYH6xLWppY+2eJgrsKOnui5kFpftfM2fq7HZBcdJMTO2PwdJckZwSsQA0N7/kthlbieiWHV5
1OPKYsjb4tI1jSvIYNVnYR6ok99B1j5KalERhmmcW72Rv+ayrhS+xGfrJcHyQqzANR/I136setfc
ff8LrgIMrQ0e+6LatqJKyfjw9+tdHby2FAsAX+BLmTbT3I7gUBbYR56G32qHpUE9gWATqNczJKOU
SlsTRm6iO1ZY6ud2l6va3oOpCA8o7NVjyIaWMa4WR3v1idnuzllqn1AoKbOTPnQemgm8185NUo91
MYxvuXkXFlh6HBAGnxxBd6Ksnvq0VUmQeIpKxS5hewn5IKdtmruS2LuEdDlKSBfBHH3U8g2dd421
nE8AjQyAoDFVlm2ZtEgueExIdPPefxXFEs0c0uAa3UeTtq18BIAz6eawaX7+DoBzj5xB39Lj7RAw
8cL9ULoVkZWcHqn6DS1pZuNKiQ1nsdyBmOJHVAv/+ZKhg/W9zJLLlAxbkJK/QQ954gRJysJcWNtG
BOkH5P5UT1IPcubEXHmMXpPJ4AyQ/SvL9wurzN/Vc/5AD2RUmxcPXaljb40bu/J94vVktnVe3Y4E
yaOrAnvk7KgBcc51d0aVnI/we0ARWcZbsTu8GokzFGXg3uCMgCZPZIvc2m0VYZwL1Z06+vialsz+
GZUk/SLSdF29YEXXFQuUx4U1i2zbli71/FhRHGvVczsCMI+1nMFKq5wWmEuT1xHVXv62VsihvIwh
g5xOG6Yn2LvbbNK2l7DqlsOnC27raeiMI99hRGFMjt4+ossuvtFAUC8KYs4eA46TEZl4aaJWWqVv
J1lc84MP7LVJSW/5nyaL8Wg/GFpiyeHoXLKlWiMtk3fP2ev02sXYymZ/fDZR2U/DDnXidzi/i4ln
PP1iXBUeylLBLZv4WlGoEq9041PSsSelwFXO6yqnMF6L3/q2/l8ZAndLZPhc+Wc0UzjsrT3Xu7OE
70oBwab+1+MhXs9ubCjUC9Jcyh04XLdQ8iTQyh1Be9MeAKzV61YMyNr8dgh3pOZrMuLWroYufhVn
yCR6x8p0fSB6YSM/13OSY/NOOAE0AFnh6lGNaMdJCSOCzokwGfRQ8ABr8WCAOhZAIzgmiH0YyHuD
lBVK95EiNAoYyNS/1qj8Oq4x3JH1my0ShgbLUhMBKu1mIO6Ypv8Mx7V7Dc1mPrCKTb7WIx6SNK3h
5hlFqE2QZRllFqYFj5FokwF58YQnUb7NTpU7DilJxb3/BeaJyuCaRA9pHV/RDXN9yK7XR/St7YUj
OQbJyAGfUOo4ex49ZNDETMUD7N4fak5tPGNTPv5V3Yur7Iv7nZAND6pQFW8Ojg9XVmw27iH2vYPU
y5r2LQ6plFidnUYXvYwgqbtho64F7+KORV/tAKT9vLBqFX8yXHOWyWzp9skW3c3iyVdv0PLYXvHb
ALAD0dgdLiszOhSlHuFcn/ixcHsx5Aa8iGj77U5zBmY35vexTT71IMXBEEJxW/S+dSGMzXAhd3Lu
Vbz0eIhw9+NlbpbXxsiBArjL1UKl0/UGWSVP9KPGMRLo3NCRO1rB3tgYD/B1W4gTZHmeeVqBFLmz
CAN1cUC5B/SSjWTQFbqZF5487Vm+jO92mvAqX0seUWJMXI8ZuhvJgtEF62DOl/ZYgwi/sYDCH5OI
C30uuuYVU6lUNhB84MoJQnrzOZPpBas+uU7zC9SGYaCZbVzTOUNClcuAqHvi8Vdq+G2n9P1NOAjq
DtDmZO9N61WPnEAgm5LRFd8FWbTrodJUEOTInomwzV8ozZre5c81GfR4NBM6WPJV39PgBOGnUtik
FnJcj9Mbh3UC2UZmPwNo05zlgGhhHYRPFKnP6eYLfI89yxbuytVyPK/DqzlMgRtnVd3xwoGJr7Qa
GQcajpyC5+lpW5DJdhQAWPId9m87dnISSftm7w+RlHkRpQXrtRBVWirXeivEDnSTi1oVHce00LJh
MRY3C1yQsZ7ovpyI9NYTucMkhTZlVNRR2ZL3p3NTlAxPzHH+UJHm2IamrdkB7Et6COrRTHB7Zoso
joudWvRJKJK9xjiT2X92ZlkDM4Ri1VDQH+4Sl7fSEW9iZZLc1kRF1hjTGnnNfaR3EwnJhlu7vfY6
IR4YaiLFxdnt1JcSTH4n25vHe9YlPCEWdEdf64lhFuCrqcysyLssEeC5I5nDQXkrhSnJPM1tG/Vb
gWVe/yiidE4eb9SliU547mt4byzLu4KRc2aRRg1LAhNK0qi1L4h5rSKXC1EoBM4TXPn6S2VEKddx
hqkurSW9RpG/XYxRMAJsyt4CTt3Zo5L3Y8AJPsCybkd3HQAusCPH9GbgrpD4qaalxYG2P1Az8N3U
TgAt6amR3ASd7Np8P4s3TkHfq6L4JanhyABh13djDwQ4zLk1hPpPe1IsIp4aQ0RifGqn8Xz7e7IR
WiDiyIBzN2OS/ijBXjups7j0bSzFn+0G/3dlSAawk4A/DQV6F2JQCLRANgjpdzdI5mXfOMddVtSx
Xjg3eifKXS3QeedYv+E26tq8Fh/xcYUXKVtJNOFeEueyT5/vZ4zoOmhXrKBXmFFldSTK9/9E/EUD
uivw6mG35TZ1C3PdY2EKJuFdJe8cRbaxQKnTuBtvVhON4leMNpHPTWO4Bhb8h9lujcBfXHJNRFGc
gHdrnDAQ0WzOW4OD2igJYE3TL+ZHxZjf/emp9LHUXN1SQ0lma/pkmPIMwYsWi0RLjsL/9xioRTvZ
bIqyxH+/ph4Mwd6zXvSOKXw5ovrm/Tmh9C4rhWTSW+JCvF05r+BOsD8jPvcRXOx9Agw1XF/XTqL5
hxGs44aTZh4JpYbK9mHtC24cklbPcTylo5ApUjxJU8ARnOviFXOR9H3hKWKsVYzcG4JM3CjJMHyO
CFYH2hNslJSDcEPEEkLscXsRLP7YiUufyhkAKwdouApsgci/Y1Tk19hfS3hlm2uxQfmEqXkn51Y6
rytNv5qzgJGFierchfz009Ab2hpJzTx8FKQxZQSHRjLGTkdiBYe4HWiX2VrBzkd7L0pOQGbta4x1
6JKdSH78L/7bpYLE1yAlvxG7lYgknnq+ip7YhLycsKQ5A5Xc86/kkP+r6agZxRDATjZURPvpbLsR
swMysLdtrEwLVR0PH1YWoTbyyIVCMtV8wb5cDaHGmHmKjoBOLKLhtSDuyviSOalnlB/HH6wL7+vz
9x3kwUH6QhcJLtK3P9lLi/6KnbZ3AL+O3iKq5QixKtsTDh1mwmh3OgqHMd2MVDtRoJqd5pKf7gfU
GgISDHDWwtz/NCGvZaenlkKASftV7NooRK2Q68WqUo21K2J/VzGvChhgs8xS7hSkeZe7bHmJUcDb
1gvCg1S5AbrIgvKBGHH7y2yrNExgQt+98G4c5lJgSEyWgg/1Ov7s7CXosOVD9xsBuPb7Qe3WDqC7
k6SMJA+uLf+HF6s4AKjhrVHIKbZekSstoaJKUfmMKL/NpvQrV9zYjmuBRNUxgeBm5jdnuMt2SyPX
RremyLMX/K1Fy1gpgsIyicQ4+lksw5EnuHcXYxn3FnCQJzAddy1U3JRYRzFhijX2NKPxzAFOuiIv
UnNN1uLfaGoWKGWojtEi22asiyx/d6Z9wa2/CwrM67F2fSb78Q0wt7LaZ0Ahq8Z3KhzW1g7uHBO1
TnoNGQ0HFrpbfAk8gejh9TZk5tBTzzL2RJ3jxas3UluupbKTLcLJVP9ldlhygSm6Xzu10nB5nyD2
eJZKccmR1oxzpJA0k01sAfpm11V+dxtwchFA/rqThW0unq+IW4e3Ujyjjy1/475AYG/TU7yMwyoA
/Sz3JA/FdfVGkuwOitJ6yVsX3l3yYq6IG6Q5gkcN2B8bZ7BNcxEWxuXR39XHS8zAEJDnqbkQy9cx
sCLpMGZczAtVICV19BmDgaK0BEHrTVkYJxkwNM7KFm1ugzwlL0JsDGPpCHDcSEy0M4WXdi5RSwrV
pBkRhf8wWomjVtXDMqM0J1VxSZAT0wV050ZyLoCCqVZMq5Zdn2mMfkN3gNwIWE7bHgXzb2uSx1j/
bcLP68DZKXylqpCBrsv7Tgni2n8OZ4VDhKj57gL6oFXPYX14tfE3+vg4lCfMC/TYAD8yYN+5mqYx
8tfifnvRfnRL3wkWAUp/ZO/OtWRxHO+Ux6My6iANZFY+CpY7jodGjQZd+eGfMnCOcawK4TEFJwdY
4+dm80wJKbb8s1y9Nua8XrZR4v4Jf5LriFe8/qj6JSCMFA9MkWr5SaSZ/0Rol/NBzr3YVm6UJb9T
AInB2WKMXRfKn6IZR0rapAS8kgTlPtUi55vVhM7xyT2hMMCcYypCg8kaQGs2A048RlVPJrhDxqZe
tDgRvkpUZCnJLX2zqGWr37jMkvElbeoI3/9CVgUb7tBOxvElhkx1X4jDJZyLIi26tvl2qOrsCu+y
GBtJz/N9Zp5t2CJ3+sFqf+k2TrBzG2n9cKaWmkEat4WTSK7TLeiQPRN7sRS5XqIOAsbTpXTAFgqU
YNm6uz5ZoLjYpXeajS7JC57BD3jzoNr9syQy9E38VlEOrBHyb1wezBUN/eW+8t40bxtKf2YjzuXx
ub//vULvla0jgtqLQPbVFSO3ISt1SVWAc2ucIoWE9Ug/oSWYFslTIQqeFWqyZihxgpg2BvnjxUG2
eUDZv4IgTI2nG/q2sjtL3Vc3avZ7vb1J64WcetKSJkv7glDNyCeux2K9f80EFAAmbIsaZISu5i4N
VSXggbKto0WZnrb4jI+FJ3yob5Nk1hckTFKMq+55+eojTx8nSfROJaT+zHq4ynxTci3+7jBkrvlI
KMlKH/mcehEhqHSUnQ5cn+fA6IrLT2LZK7OKi4YM7CV9GgtEt8K4d3gKwF3ssTfcuMZx1ggtIpNz
Ynxm8dUKMLTYfc9uj0/Y5QXBMhH6nM6omEf7c/WRrk50T1vxuO48Alzopo5k0BGOfGzzHXwIkpRk
FWXRJ3TDkqEP648U//zzeQYMeIkN1oLWeqPGGMfss3PqrlRqscuG4xrIgrCjOnHkwmKq15BljXzB
wO5vA6NxezKcImkrxrBv1IAthSlCTrNmPZF4QZ2KwjeNmI9WO/exSDRSSOtqjvKXGLU0l3Yscwze
TyGQuFydczBJTTIPmhmiUjnZbfavQ2axmoBHfIDlfm4U/Hx/j5LtHHPl6rWnJTLV3165liAjWESh
P+bBAPdYi0/GKk2gOutAjLei/PdsL7OwBdxJgWQaVuo5byJvwe42CuAPNgC8x3+lDi042ifCl0qE
SFvygpZ+t3wvdxqxiV5HyfQzVyfNsyzIXFY8D2+YXyfxrK3JEMFtu/WHyasvLedrlmvrxTPUhq6i
evWqEzsEziulEnPKRvvXKvycqQkFnJZQRaNs2wXgkw5nR7he9F+H42uGq+DD6eS7aJiGW5L/VfQt
711f5B5UMmkCyiT9sUDxsCAVBEMKwLnvGd0VyomtRExiuPeGVXXvEzO6mVw6TuJZkfsn6k1ipEsO
aeh2r7bUSXnqK8X6yxC+x2uJ7Fbvmdo8tFHDJcKwRtPneNpM0qNd1JGjqMkZtBOSYeS5xwro1TEv
rOqXNB9mTwXfAsnOplP+zdHpwUIieLn2/w/jsBBg9WLXkwpTdFoe8a65ocNALqAN3/1g3EqwSE3S
QqWjnyx89KbLFsoJUGnaYhLf4K/He6tWuNDuLbg/TJRKu5bT+PfMi88/PaKJAEs6ZyFbbyZRI1N/
lA3fRBnJlcN/cQsNncasgL2vXG5Eb/3VklF7yDi5ff6sHAEBOw1jn8/GZRtZtzacD+1oElYumSEL
DpoxdKqaRK8Bc5MloOJ5A3DS41loD0Qs7PoaIujdqBpFG2yHNybHXXrrz7D9/adBfYEjGNQJNHzV
djOXTbxNYYC/7zw3mMh91O4O5kSXausDHjydClwnR2y+Oq/UKGqYyF5wPdwe7JG2SRCdW2+0/wnX
nsatb9tACzHvAOXrzlX9YtwUlGreGzVBwZCKfr3M4TWcd01mT0wCbujGPXO/7eFG7bLHKhCGZMHJ
2rSA4odLACz/odqAfQP6M9API0ZD5TkVep+I8/yftXESFjMyD7brMBaAnpf86HcaORjGcizRacJH
YDetgkvk9RgcbWY6xjdp6sFRRRYX7+oPFWHRzMiofge8KVzE8uPIBA6j0nDJ3FSDBFMch2Y0LsV+
ssiSDwd1Y7Qi9dg5ybuoujiRh2EgI6TKHYgz6BzuN5F4huDXjjhmtEaDIWAaajUqVupnkKYvPV/S
+nqIy88W05nDceG9y1gLjaECUVGLb2m2qG7ZjjnuNwEpmBJuEgVw27tnhORm/0fgGBJyL3uHra2H
ukrEbwJzcYztFbZMurPOXOctESWwlh/XLVX2q8AKCskC9Ib9N26PsM4lcInn7GRagHwG97nMepgM
Vbs59lfUr7hwNMXDkS9I43VR0WD7nFaoPVVODy20J8EAbiUm0GaqmX33qNMEzXSorkKRKLNqnU8J
HPtk4XC6Q9hoWMAqj/kTKHoGGFkEdRDzu3ssAGCQmNSShG+FhepNizTko16xEEqdW4pbAdsXcGWa
KpTIIc0hnAHbsZEqCE9/6yiKlCuaX4bgyUUQPo/AzbLEhjLREVKumJiMXaAv6gMHpHdd7fZmGPaM
F8QfAEPjIHhoLXITiSq8L2zorER/mL5Jl5L9eeZlnKoZbYhm86j9jyY9gCHDs4+UYrAoredPSIyb
QWgFIszJa9dFTsPZ+j5uBNLmAZZ9JFXczcLzCfyqNcLy+q6IWAq2R3EDmhw1Ppr9IBTvAnP0ATv0
Pt202HVnuRJ/Tp+ph1BV7xH4eoHVO6Aokh5ydbYvfdSlUsoS40QVEII6U/oWjz4OWLsn62jaFijw
v//21+Vgol/SE53WqmGtz3uEMBGNS5L+RXhqTJbVGGQl6kEGlD9OrRli+z5WnpkW6NuCb3Pm0VTk
3tJYKhE9CloJ5ZEmdlsXjwryyCDSw7LENjGjUZrg4tS2fWBWofQKp7xP9kucTCl0mJoctpVjbtrG
IKdT7ZgTUw4kAEdOZ3L/iWkvMQr8PdGQpnf+W1JkE2+FrRPjH5HOsOuRmdOBQW8FrEaV8QxmTT9X
ULBG2GL/5h3NzZMMDDuKwxxcQxqbztqXGQn8h55H/oBOmPPgtks+cnyjaMsCkxojR+tv4aDd8fEo
4An5jMHeWwN7GGYlQbqKwls4gy5yCzVhuUvKsdHPz3YG0XQobIoglyzKWgswtihjs4/OG23oovez
cX68NC2ywzn4r/Yx5AOSxVs0vjWSktgOC03NrtmOgfawA3AM6PGvNpgsNk5BOVxrY2xqf/rv/ijm
pv24wHSoxDuHBtavD88N9jMaosbZt93j/4na9Vdxpj0LajFBrGf1EtoQXqCB7jmrBQIepuPC7dWw
iL4j69XG1eraEIZGHp9xOudiFVZGnP4E4EGuqDPP4RGrxYYGxrK9U3nF4XanHYVD2czsofnSdKi/
tU95FJ+VHiI5pCWkKs6abrSwnJ6aWhrl81B0wkoPkr2maMg1tN4nqxns4Uq2hOdE8HbOBzuPqThG
y8lFfgcrXRRQtXMQEEY4vp8v7o9z4SNix+7vWzC041AJkGcFF2cAgRxPd0+/CAwLDyEHcEqxxssp
YMwcPKmkg0KC5Qoa8TFmBp6KBapopUKD5ERo05keg8CUQP4PG9iGQhLTiWWVhFR/MPfsXSn05f7J
+h91tYQRTpbsqXZmPuj8CdyWQ1AkLs090+hB3tePWU7RFIQyvefFHVrJSdII8liOoC6dm3F1iUDu
N/Xug+/hbKvopPmS2LUGPTf/QMOs8T8r61q1GGPr+FTUQgxTXk2az6ZgBvRNea22h4VP0xxzAlhK
zIV3bPl9s9ObOXKNhdFsKMrTjKGMYLDbLXzAbBhC1KcRuuW36Ca80IU6jvQyhUYsbpZ9iskMS6f6
d6Pu5WnuEkTwJEGUc4uKQTdTTtZOHaoV20erisW1L3caaCXwY62MURjzc4nrgTrsMCZ9Go6AZDlM
xzqcj3gwgOhSqUB+kLnELzSk132sNdQwwBbJwCXygXLA3J8wLng2SrnbcRyXjCx4Z7h24zZz7kmN
MQDWz7DPRK9GefLGRzEuRkaMUybBQ6lf0Hf0DBVTYPf//KWtiFqYQVNkLv5p1xYEqOrJiFqLbKVg
aQprWvO80qKyXc0sVYHnQU9prb9XpN8cCQh7K42I4aj4ld+44L77vkCccfcAfkV1Wq11x0b+wQZI
KiF5BtyPVmV4lvQPGppCX1efqs5pNowMZ3FPHWMFWE/76vfpY9FHbqHA3sciHZEBqAh6BnydS9Bh
Sp5F4w8WrwhV6SSfmsh3P9oCOLs6l/udjwxzvG0R8iFgakdvOHJ3zLXRWfToIT5tukkPscGATmU6
WLo2HGuvKox3Ew5zC1Y2NXf0x4KAPrc2L1NseVsFuEx1/MLVSPDekVekzgNdewqvmTjXc1ljra57
ws6PFVZr3hX+39Yttz8LUJEynq1AszAR2MjV4Yf9+InmhB0++n3Amuj8RG8JNyxNkgKdBsKM2ugC
TpRfep9rdbKYjkE7H3NiN1YhHQG/qJVc3BSYs+gHLAbFdwZOcPY5+xYWQtQIWQ9acJb9iFcsFR9E
x5lcWe+4K0GuPaOAwqTInrofBvE9XLvmajV0Xt5Dip9SoxS+rxoADJhjusQC6+8/efa3uSjbZTW+
fkta7MJoDt8bvfrtmw0XxH5sEg+A53jpUq8IZWxkiWUE+aclbWZUhYLE+5/Q2pKrsgqvGLB6ESzw
vmnSU7cD0kgS/C/3zUGvkyjCtkhzUtsp4Fef3x61bMAZTg4laCadWGaph2+HlHfVbN8zINlMUFwE
AkPoXP9bBW7EjpP0Q421LdqAkfIm17FAm/eBRpkv6tVuDz844ZBpl3dwkNyHmx0zMX4Bgl3TLq8b
gR15hljq1Wj1ms9gDEXPUD4bnxRLGq8rMW5MrtUIVx4ZMGW9k6ynVwM1F76Vw9KPSB1Pyp156nDD
UW8Sh/+SzX8YWUGR8tUJ/zCpGwZDjFF5MaBaCPK5crOq21bYnpF+xZjmQmrRfGmzyCIK4z8sNuS9
ZGdZVisYqMY616xGwqO+KznlC+RpuIIHR0IRH7AF4P6uUNHDx6BSXiXplJehcm4XX82ltwhBP+PK
std29DrmJaNZqpw9vnrN8xz5uk35ecy5vqz+0+LUJGz8PkyM3bYY8ddUUKhcG6S6FazW+coq6D6J
tTMx7AXpCkoYynfq5L1tPhPp1srus6QiVP5VXzsgAwzPs7b3KNLTWkayCRL9ao1Uq+dUCJoLTOPj
1585Y38hTaxc8NwukrC+Zyu84RkjyhBbI6GuEfextb3fW3umRpbblAZyt5mroObRhHXrno9/xkTT
lfWtd31YJ71BHnKxJebqObQ+I8HaPZdV/cBZB0iR++Lg/DWClwqd41X+/EGrUHDCxk/4Q3rjfKwz
3ZT9Ds9yhlMEzrpoXEvHNQzoO+xIp6dLSRHQcmzVpxQLqmDMAnRWL7LJbPWc18fA4ZuBpJY2qady
sCEFxgm8O/WZloiPZ9feBq/tJIIEVkG/bsZvE94GlRl8ObEjqwjbFuMfdwNQroGn38mE+imbx5pl
+Y+oJtpUouxypnucez7ssgfQK4q1TjqxxeG+ovk3OW5KSS4tScNch2EvNqB7tkq03d8U6i2nI6f4
pt8wjkrQQjGcKpIAZnhlfFR3ToWJ2P9+2BYMcKS4VfWW8jDrXr/WYpJ4IMuD+xJntqxou5lwmN5X
JnAlqEepfRQR9ovgbReV0pq5fPMXDsged5RsXoMGhbdagyDNnSfEVBbTdpigoTqH7J22T5LINjSj
0r6AL2ak/+MadSXCEiR4yyiiM5IDx5sJSTFSXn8mYQgwT2RqAfKu1zJxY4TjFJkOfXekjabuWA9q
CrpY0kChy1c+p8R1WsiET32OT9fkDUoINCCZasNpHNjJRCHii/F4P2vTqfw4vVW+x+2YWnl53Mw1
fm1PLsQXiX8Qh6MeoswlhLe+KGoeczT0i8AcfWsSFhsNuyanBXNURy9s+vqSd0jiGo/DGYqzfrLp
TQVE4EKYv0FfGS57wLZHAhD5u2Mu8ZOnN6lpqqeA3ZuJVnmxurUx+mJV4T6rTy8fhj92RwDFLdZ+
mrLdBmmOIJ5gwY3jW7ci3ltlHs21M8YUPntzdx3B+nrxkTGPCn3s3eSQ7J7qKJnpZTo1w6USWgHn
Sz/Tjkz7gBU4HFu+m2BcvNhhnxIsE4S2zbmppbWuw49XP4ZRTWd5lCwEo1wRfY1dCMl1xwAkOhfI
+MHEjzswirltBa1NVImua+9+VjIgAM5q410+eJ/bK1hmFaiRqgrAMW1/7gCAYXkG9+HJdx8FDraz
/zgyqv57vckcgx6NDnjmxq26EVpLCNyjbY6JcdPm1tVffXJfopWwzulw9wfx+0/9TEfhe7T35St7
sXl45VVkZnJMIFvb3QSq1ndJ6fUaDa2yrgj1hHTSBvxkClGTOJn87HI2kclAV4huJq/sIl8IDnVq
69YDayaGOB4bRHOhNBjYwlYWtcpuJbMgbc37rpi/MjWtenYYkruUT5L9yZSjN2IoMl0+qMgPISUa
tOdzVZFa5LCawgqG9tB9KKJuZoEuSKSieQsbgxcZNX414VAwGvKqViHfsSP8vgowGXwrrSCum61W
UdVwEL+URBgAhZ4mn0gwclXmJuHzZrL8lPueisAPwEg8ppfExlR5/b5d5TujAEVQqN+3a/+oW/Ag
Xl9XjqYg8oN5xq1U9nvi9xlBG96MQ9VPC4MzF6nfwQ0rCsM7BciACps2hBdToLM9UpdR6QN8NxJI
5rAmVHoTb66oKhxAAogUmyI3m51ZiYylgayTUovvgPdIV1uGXQJ3lfJq1DFBr+SwDA8gdd66lH+Q
Dr56FRQ5fbixSIxhUIqfxVmzaBjyxGhVvsWzfL891XBashJAGQ2hVID6NT2aei1rLTcbWiprS0Yd
TYBwg/9dDDu/8IilUy1er3cmUVxFO5r9BPFNl0v++IF97+V54FcDTwknbq0jz7ADinfq6t2p2DrU
bdTu3WN7sMBP7g2eeaF3LSMAT1B6hGl85RZnvvjFr7SJSHGyBWH3L+HKjW1jurgCRS8uiLk2zad3
EwLmPwk8734atdmbuMuSLw4njp4rQRHvg/QqvPe3FVpzTykSdWgPb8yAgAteWWNorbivqrB3Qi8D
VpliPw1oh7suEPd3QaG5vBByNPsRmmYGJQKFBBcncVyPGISctrii+G0cExMIxt0Ti3Cb42RucnY5
snYJhDi8mDrjqTpVltTIreKKiF+s7iCCKrxmYjk7cLQNxvw8/S5ZpqPIwhv42j4+19caezb7pSOz
s35hE3sJe7nwjnMisq8xzVOUxH0tlJcW1RA+/IV+8d4l/JD7PBVR1KYh4uEOQltn1S1AM5DaL2Ps
2vYs/NZNe6GfksR6hMqyhhBMxvM1UVsYRE/Q2dsqdqTJHIq2WzbTYc7HbWjF6NRFnuLfzFu8tzFO
kGTPOYQG7TVI7KtxsYZGkGqZNLUQvjndseuHkJxXrd7gtiVEIFtfT7IvunxN65pwt+Y+moQv1xJb
lxpfIAodmcLwyDcKR3lxOk6aBACrdrKN9DggcyEg8CE4k25q0gkCHKAcH24d8AoNlziSz+ivguT3
DEILaaSfz2XOoLRQjcwPeogwTh776XSoanp3Ak3qaZQTZkMdsTO761E5RG9WMdlHS+E38nkhIH6V
dvsK9hKjLMCte2E0xcFqKBjS/gPsX0upwy61M3P4uTeLWjkjrs1o5wbsmq0SJ6/QPh90Llp/Z3ae
6gYrXxKNeUjKen3vekySDzYJPbTlwFhBv5sL4C5iKILJV4Ddjk7V44RFwL8XUcTSI8BUKaQbppgb
xeXjEVhQrjcoUHwBhG+ojLS3N37oK4ITe1zTeD/UVay7BbtZ+CnwyTlRQjK7kP88LX3uk5WJJ2dV
HWCrR9dCxbYX5UC6TjZq2Wi+SjvNRhplpw6BqVcwzTnaMxJm5W1iLqVo/nhq/He0adcloC9nQLFo
dQ5hHmpaEgJDbw5cKDIZoVv1htg1HLgzlw+OTP47DQzuhUk0TENBjvW+gGcc7UGNoOKIaTu4fphe
0faH4T+Y2dwQMGKDYckyvDD6rMrtweKAsi9dVTgIJJs40cjqajCdVvRPn7wtjwnj0mLya0qyP/DZ
cvzScUgWKlv7CFSH7cQUsqQcpBX5yyyqJTirO5rSyUB/xFteTKymUgSELwGvVQvWDrHv95u3WlSf
dtIDEVY3xzgQWDtw24odwblRwPPt2R6CA0/lom6qFqA/4hAkUcD+qQ6DN36EtiDHKOWBs+EzXlcr
Mvl97Xn35XlU2XEZPgY9DiACdTc0tTdT4L0hW0fQk3BO14fehISpIGzjNWoMNEwOHanMkaxTndJG
89/UZxCzMiBCoXgSI8At2C2ZfTqvbVjBU3smHDWVoroyfMkjbA3RrV4IPfaNfOYcOhccRtq+v2BJ
JzX659DUSEURJzLEl+o4sXf5J7DjspWfqL8ISyXitKkN1Izj935eNKFhzDz7dleOz8bQ0WJZRkzE
5Uo3bpflstC44QHi5JoCYUd875Q7axehmeLXRXYf1SktENcX/f1u+vi1ui2pGb7ExBJjY7vPQfFH
UvmRGHpvUmRj4r0DY3qR3tR3AZky5oQKofjbRKe+DBRCkNFs6uClXp8rgpzkAyx1ZXaAtgBIeQNq
29GqSoPEoFacJ6maAEGNrdZNt3yf9Ez+Yoj/T7GA3hHZFpKdDQDPSfUfEGipIiIiCosqwcubgkor
iY42lty7DUKjEOBesFTyWCS3VZpP5F7mE/G0BdEyc6GXJq2M3Bh5rQHGVGO7mG1dhLwZRkU6rzSM
zjgIovz05xWwCdcGW5ooXEACTFv19Th7ReK4kacDABTELY/VSfOPQED1xLawun74f3QPXDLCbeJn
cZoMWB41z3o13mZilNI2F4PQTQ4GOY+sAUMEmhUlikDiNrYbco5QcKNm9MVbIRhAbJBI7Gtf/vRO
y+cSuuuAfuakBRfhKfEeC90QZzama7xmjA2S8atymeZ+UGi5nWLGKggWFdcezsC1AF1etYAO305n
UbM90VpUAyTPYYd3fqRrfQouLu4mU28gZZ1TuPSNU4Rw6tDwWkUV9fuu26ZK1E6zCBD7cnUC5UqB
TQFww0o3lbIMKRqbc0n+a3stOu+fyQq8ZSiltla1sFqfuhLvtUPFlqeZWuGHdi7XiEVlSQJksXoM
uHDH0kcRMsZZY88AuH4HZixGFUK8esmo7R0Z/VO8mNwfv3bHQehTGI8kK1aPtoSUqF9DxlTFdbQ/
KYYo6NmK6wsepVNx3QE35593VZQfTPafJ4lLx7EmPfOkGj16os6sHnnIAWQ+ppUYn5Aq4ZBwJGkk
diDejkjoWW2/9eutZAGEi7vbEZxS99M8dodv+Jklv6GLsV/p65WcOAUQxedz9VyrYmJbfoz0mUuJ
ae2Tj+tf/zBWWx/nTlHUCgt0F6iChX/oRVQLGCgU16eiMIjZASA0297Vw3h/p6zsAdb9VXxrjifk
xIGxVDzbn25tnR0qvp42b4VeJYx9qg2qZCeTflsJbzI9IYJSwgLV2czCW44uFPOQ9Mk10Ytjk4Rk
0dr5y5jBUhM4fDx1D7ih7nAxdi0RQGjFSBOL+w0yOok5yUxuWomz0TBZIucb/2QsMU+vcymReM7w
TO+/P5UMcFN/hkzCz3YplrY3QM6w+MY0TSk1Vyn0DXAp09ct5ZHb+P/vvm/9TeACNAarheCzxuBJ
fBP8pUUqGwu6Sv6k7a/EvZBnDbtx5GmE0PlngadDvml6TfHBZYDTDp6ZL11hKB6CC391jDEnCLZp
OE45Rz4IqqI3uMxrhZ30EhFZ24A6KMCWTXi9jmgvXoH6vX6o+RF67dS0nOpTSyj1XJicdDA/P0lG
zUolY6zZ+RQQdADFUj5T+H1XYHNiSsLpmozYkU4d3OiGsHnapLpZpb4g66AZ3VAA/pvnNQHP4CEY
Z54T2/z5VM51D6uB/4eLQPJnLTMsCju6tfS2+XOz+FL6Rkf+8jRK7t9OIYh8XAor+dPJcftJClan
wDmCA8UuT3HuNTM4hJAUPBHlnSkLxQYHwri7geBDetr44AvXqSNXqV7aDKUMQp8xoWDQTHve0k7W
kaaS0pHuZ421jKykPVmT8X+49ypaGzYfSkKp09eFu4lVaXA/rbXnvJI/IAQUDIhlwsfh9Mml4Xnb
RZGuhL/YYqruUhwp/TDA4Y2Vy9TH3+cwXpLeSG23GRZqMW5F6i/sdqVA7rC1yy2v541vudh9ijY4
4llTgBlgMafx4t9cKO9ftYN/ccB14HApnFb+X9XcYnuaSWmGV7r02PO59jqWWlBGRgGkTlLw9xnk
+csTCiLE7qGtJp6Z7fZa5iAIj+jcndfbz7bYDmvsa/pLjoPOLeMs7/3UWdFg+OhOL4d1B6zzCdX6
IhbYlgOk7yosRzJlfu4b2hzY0ZpYYW0B4esxukRhNelKNLJfB8jwKNMcb5EC9CwLnr+BeiGJD8O7
wTw5x76y3ymaj7kB5RUTfltZ1WDxC5fK3rdUWduVIaLNzOkBwBnxM8x8Y07l91uNMEJ7gu9CU3/8
af4rcAJRd9939jc9ECSw5SPCye4c8cLBgMdZo4byeEtvX01pS6/PCsFbm/bbYLPIfZyF3mvvcYWF
I7hB8WzjxyZXcavXAB+GFxF8Fa/BRjVKEH/y2JyPxc1XofJwyKL0/b/tUvVihQd+65X93xT3Psvl
YnJx9ICFgZo0O2TcOcQrlZt/tv1z+JjKGVW5r+Jgo1jn8QJHd4BAI+pnCjk+XPfcywv+jEP0ejIB
+UbgpkFt3aGbxU5VTSAuPjucEessu/mvqwP30isFEaSvLLh8pqkRH5y4zH+dgNab1Kn1ojJ1bVtC
sNZEeJPQuu8zSMXdM2EPlj+rFS/IKFQw1Hhux6qCOMFn8A3WRGO92xzU3nlgxRdCXT73sbVpeNmq
LKXvYW0UPHEfwhAex/UhlLlWt2cGjGxpbhd431WO0xGi+7nUhPQ6uEZFkjIZPvGqva2QGyCiu7Aw
noXVSgXZ8hSMIfDeBE1TMFdnnXrYDwoNNMb6uXz1DJsZZaOeiUdonIEvFJeIThMXFxdfgX5X+inz
AaURkVlaCypoobxw6f2u51L7JKQXb1UaNLNeiWKX/KjSWYW1BlbxiW7HF1Iuy4rz4g2bjkSTbOSf
SKNUC8N89oA3IKf5eaXlcQQv0V72mBjNtM9Bv0Ae4QTG1KDorLBe5M29aLTawCLqIVwLqHBsyr8N
EEk5tFiB80hIcboNce/2o2oG+LzNRT28UYgsIj2GBM9sa2rT7M5SiI8Nu+hxQdoq3wgxATuspsAJ
rtIPFbT/yy/hbzInuqHnXc/b0fhbKzC4tglUIR8A9jxU1C+I1kCTHpyKCxNUWkckqn1ldtNo+rUC
O7G29rtzlOYYN9plk9TckIMTJxN9nzwCqH4tyyKYF6/pWGtYse3/0+uNSBuAETVsbVTNFdDCHMQ9
zOt4kbL4xBj8xbOWrAXqMsMd4vKmxCOxAOs+tLGR8IEVlyhqv9oDdEbbhYFFMLG7ifmJyLI+GVMJ
KbU1s4oTZ6Ik+Dny2Mglk7I+CZL32Y/2y4pxXjm7qFAngSE2G+OQXfNINxmV6CxWehzSUjPPYDZL
9OP4SXRGs4oc2H6DHMCHxPKJvWkoE5upWNIH6g5EE0yQBswixumyHF1dwrmAT37j+H3npEyioO4y
pd5FRprbaRgi9A3ZMRbH7hSafOz2XcqK92NzEdu8iF1e838YanHLxumuYkaTGjs/8nEJnE94H3Cw
hQQuKvGY5lnL1wB6x2iuI3KGBuiHTglc37bxveKJdzwKE7U5D5PLux06yNlX6prIBiuTY8RTq/Ld
qLLXyT8/PxYlSA9+IOPNWZUi5tcmxw5V8VQqHxsVJ7ER0sdE7Z0t0MZVtG81xjxx0XU7LOz/0gAY
ml8eABIvWCns1QDV/pBl0EdAKcZZZlbBPbRybuMoVQxQyqZPo7b8+6XRCG0/0xz1SqXMWZp2Ta97
vcmfANp6kcXdE8QwEDB1yF9zk4/IJchV93TUEr3Wz6nJXLERx+Dl69O4b6pw4kBfAwnEKd01EAf9
Jy6Uf9p7U8bwCujusT6eEsgE59g+rUOFqgxzWZI3a+54cVnBeDuB7Ub+WhJNLWWtErG/87tAFruM
9ZNywQFRovCBLWxUNY5ktDWULeQ7ocjhcCWFhHS5Wd+K1n3v+NmPDlSvL3wHaAxF1eAxxUbuHQCF
XBRgtOGMpFTXU8oUB0UolcAJT1IBF7KMTIBhnNo3zoGUr5cLEycYN7LKODjFt4I+N9EWo5+A1Q5v
EgbsGfvk4/Mm+O0DORPsLlbKAya9nQLAYhIEb1RaLgHmUogbu/0jmd7cTuDUree7ZLMI4rEohUXo
ja8sRX1/cwtrW3lu2Gxul4kLxOsouxE5fSkX4ZM0joHI/qptiWT2exvXtw1oFfRwqkamExXeN2ZK
KuFI7657pC9HHyGI2rqa5RMTdAydUYs1E2u3aXofuxrNYRPaUsfOEYJTtOkGqgYnzKET6EQCNsTY
xRUlDoZbCkY3tJEoD2fpLEWbZLcuC7YmaZEDyIJlGN+Nh2AnYpu/I0VeWh/rYLfeO37tROe1FyB3
Gjc6GH0MTVTzS25cnBi3HZff1lijHqnPNhlMlMl+zpZ/vViq17JfWLX0kOFmAHRJCe2ZxDaTHdPE
Y4kYnjOayBKXvaOcF3rY+Qtwuh9xm4XEKMMkpmOSUunW8AwH/9SQfVyUdZCqYmGwMEtrq0Kiolw8
M1eETYBahtV5iIag9DCulSAo+1Ab36zBOIMmPWGNqWSTLJLv/9MqyEJSOlqNvd/J6K5qa3sCtxJP
b+R8IK2M7ojs9WhV9ttAq1yjMtoekQVxO4ILGSFAWgV5+Nbb5VgHeOvYWvA5nsP5BNfz9gRQ18r4
9Fs2gMYdWlCoPCSb+2OvDtMJUbddKmBvz8jJdgZhvBjdi5G5Bl8F3CgvF2aFQ0zPPWPOzGLV1X3k
JQ9oLzK2UQXP/m8FT/tLx38W5jLbKbkkscCvAErBp4Fofo9KFk3xskOr8/jLZPlDNVx7FZApXAv9
uj7vWjj35K9Xpvr3Tfyi00ExgkyejdeACdyatqnV6QKnJctv3EXx1Co7m1M/LA4ecHWBrNFH2aKJ
78Nc+cdOQnkkXxLRSTuZOdxFHHLzKFyBkl0PcEb+kFgXpENesVax8ajxJn7dtZoLp0CxW44Tx63S
cNbPRrUBZwtstEAusLf69U+bKSOX4UB0+byRRjFujQyiEbxTWWdBKMsLVGTyO9ul6crNnw8tLqD7
bF/eS6DPN5S8J+uIjxfWP85MCZbPKldPSiOMaooHLt55FrqVx46/6FyBxcF/2L39Tzk2vWdRYQeN
Rjgy8u3K7T/UjTtSm9NQTS9qNHFUmSXqe8YzK/O5ucrzfKNCPSpgCgJ22Y94sTuYZ+n/JLnuub5a
iJ1SCaRPKLptNYu73tWXwSh2L6oMnICp2vejWWCJLlb+neph2+BurLD43lNvLlTjPpvFsIGisn7Q
MPVSoO86Kd96MxqHVuC9O7/znsdKwhYz3UmfheLlnQeHxuwDhNpCEbJSwy2KkFBIP67J33KxEGRQ
gXULiIoNjIb7XXB0Y8ineYfjWYfNYrs50ivvcqp1571IAmQyie6airC8SVJgfYYrEbrBDTdM/F4Q
VrWNShkH3QrKpDVebkB8BUOFs0J5MNG5s7Z2Tp8RWBO1UDAcnh1b0H4nN4D6Xz/vV27xSCz2ug0Q
ip0AG/Gws+JNQET4w+RK9qsjD/ljUlUcbyP5CKbTlzaTTM7w9MoTF8gBPgIfnNGY+hRTWmXk1G1m
/a13er+5hwt1ISJVqj72mLX1/U1RyxoX7YtqgTWUwJtNP2nocmCvIeVfCj6Cvyg/bWIMNm4no0uC
fY+0dYcsXecchya05vu8DOVAy50vREGNOM/Jd2L2jp+pWO3i+8bJ7IdS/ptlKNRrKAz6wJHiAGmv
9BddGQTKJ3dSpD0sDT/baHe6a7FujzBeI62P/hpCkduBDmnx+FAL/KsjRDMbR6i8I5Uqsiz7+fQu
sr0b7o6hFaXijwyJfpiA1nyBvrrM5mZkGOXDqCmyV+rnziT/qUTcarYFytHlaTztH0irjwW4Zi6b
JbCZUMj0pZEZe9au5ey0UzQ4yUxTkNek/1xS11ypRlL2omMKmNgM9EJTSxnLsYiL2m4/E8eMS3+9
rQgsFVg+mJVDkPZ1c88ga/F5NrUzcGdgVudc2HFC8igajatcgf4NFiG0OrJTAN7kj7q3q4Ti4r1S
2qlO/FljprX0OPl0hZPRFENyCPfgVJABwtyAUr+0zSUu6uJrZccyzBiEwfdkZg83ZGLL6A58TxnW
9lgoBx7E6ezTLpHVZeIJ6o7MGg/ZkaCYeh5Xdmx1SRlW+GF9cRMnrtO50V+fcWSkxP8LsJxBbYlt
xQ8GFHrELm+NBxyNAbgGf7TXZhol4PbJT9WMJpNnrfeidSvmhAS0XMoUVm4lSn+vRJ3k0MZOwIm+
OnpoAf/6u3Zo+xOwJ1BXQX2zY5wfz5jKvQEO6bLAZMCRGj6dqANXPfnUYB99lKKjJpyKq4Wwc9Sj
6zEjmt1u2s/dHHftaWI8aeJ7diAod9nOkroyb8ANHZACmHQe1t5xk0sRZMLc0FTwocSCcCcZFfk7
Qyj1W9sSD3Meq6WJu/9v1Uz7JR8SkD3j/rn8If1qJVIE53EWkHoH3Eql2htX8VMy1fWouyK8xD2k
JvSnRDeHYS4Wa6RMs0MDJj/5i2HN3zppBHXDG1+qulLB7LxayORnRFwKjrTErghZTYa4M1J8ieEe
kcDz4nO0fx/R+5Iyp6PdlZ17nxT5kco+5I+1Gf0d+8d8vr5qJ6IC7jk2PzAfOS2rvmRnO4MmQgvr
AuBL/24+eIuvLs/NWZ74jAtmM+Fz7jjW1BEVkQTT2JPZdi1wqdT1Q/sV2qRuTnqvtE6lNdqC/KqN
tgGDrdckWV6NTHcTauMyIGA1WuZq/m5+064XmZYqAUsIyFuibC569EcaczzDEIDbo/F2/9F554np
tom32yDnVWFdgYh+dIXH16yN+WurGA90WSUA52AKDYJ8w/LGJKe2r0BXwaMGaFsR2/Hp5Jc1GG+k
Jooq3Vr60rVb84fNq9ZanZeeqvuo4cAvKnHW9IhtBKUFobYghbCZU00VsYZ8mGLJ8sWiA3tRcLtY
gnLc71NFVjOyMDbw6HMP1c4TKdwoJslg3NOt3fXY9ZZ9mY1/OeOy8qV0n0OQmAqnCURh/seQ5bjE
Ra48jpjIArzxl831haVnQObbfkyZfjNNHozt26cpHCBIdFtPJi3zTYJXLQZx5Izris5A1mSlaJsa
O3A59sLz9FkMuDQ8NyZk/oD5YAx7/G3Tn+4vz6p9H56rYkV+VNiByokeVJyw4VPGkMMtLu7+zRIj
rlVd5jlKwfmBoUsGQ0t3/QsqDOu1afasbJH4sHlIxSVyygSp1GmA1KH4yC8vte1Zn9woDgahyoWA
V2jVx3zTbGh9QMMeEpTzOullxCFgcrOTj/9yOi2GkcoVcZbVj0HRfTfrwuN7MifT1BeNj505QDnq
XFt8S8PoB2zAoojAe7CYysMQpHBggoCKRzfH/uW7BrfThDAM2XwijoWGSe7NtdokZa3xSVlv77IR
a/OHcHcbGV6L55A053mQ/QhxyYBv52JOKEohCQQN+rOi1tYjtNE0tHdNcocGMKcLc5ia/2Im91Jv
ggA9tEXzeGqtZmI/3sjnC0Y0NdATDsnocB4QV9Gr5Md0jwhl0FZZ3f5Uu9lq3WK5z/fRaAVYnL2E
cH3hA5rfLJa1AnBDK4CK98DTVWYw7GOtL8E50YTZdwREh5eTGv8m7T6sQROFuI8JlwGUDZ/6SZIi
9jJjnQThWJ8FqFfwqZIH4nd7cApkxnHRdpuLcbHhMHYCKdLxAZhF6QggLcBLynieEru+8fKpqsAA
fakzhBex3rfPQla+081YVLOrO5lmOlQaCBh2XPDqCHFrqia7+mkvX+I3kndb9A6bpDCAZ09Q26+G
ZhBAMY1gVmu6zO493kZJq0fJ0KE/G921oarJJz6SEOX8nJzRcN7YlsWU8EILWqvtgPHnPJ1OMcby
CJfmdD0UqceeD0RBQQGvLWKv7WaNYcsdctrPiXF2CYU571zhf3FBjvHokctgjmjPYWG2eBAjDW1o
Zd5NiojUJOJPB9nF19yMdqmdbPu6lHH/J5DkQn2xWHjHniKu0lmPUWBbmL2vo9Z79iSokkTOYgXg
2ttrV9umQSjQfIMri9vyNTgIuscyg/2IAVk4vvrDtnWGSyAfU9odDcQAj0uVKe4pnwZ0SwjGwgVy
zLA5CK6ZFMBrURvn5Yypz/CCewv3mNCzSMv1tNJHRpFlXPmYWIOVE0SA48SrnnidROdhsXloH2H4
gIjtDfQJMlbPxib2rNMhWJPN8m2Ju5NvAyHse5qHzHg8GIJBacXejsznLw0C2ctfG4QJv6G5e3pa
iNBqqwQBwB6zJPH9/u4lf3JQq6Vh194TyCnud3R9/+YwWnFLHBwo6W2KtDAWFB6Vyg9OxzUTK5Cg
M9QVluIBbT2rqnsTHjLjqrBPObUGsWTOqzp+566MxuWwgaFpYpZUwuRAu42dg5YF0ZwkpjwU0BJM
bEYTzdl/cwxgsGK4hXC3OWlZYPGTigZxi5Xh2t1rYB/2qk2nV7fWuYlytCe5kfbcpiGnIDXq77dD
MtjrLnvvwDVcIW929JSkx1InJVQP6qIXYCKb7Xq4VgkcLw5DUcgmJDCLJQJoDEBm/QGnBbNRZVQs
uR3AGFl93G7xvysgbTsaOjSKjfIiT7g2fyba00ngwRaS7WboRtemvtOwvLy1sSEZfncD4btI0M95
rhYFS1KcsTqxmEhbwx6PAAqUSo/rVB1xh1yX7kzgmJeIfzQ1s7BS73P1HktKSYsnnqHDMqzYDux0
Kb0nmSfLDnEbWMClwUXaEmOtZD0OjQWFN4JK5rTnIj/ej8etP81YxOM/9/m/9JnD48771lBfjppS
xVrFPbcLa5HTH85P2nPAm2jlqz1I0hY3r9ZMWvn6j3wszbaVe2o5T9CMnEAwkIYUwsoDQ6hmPbTQ
Fx7b7QssJ4bCuHJ6mUmr11mhYcRuMVii57Y9CowT1lPV15e0fRzYf8aGUqgQPS1mwp9Pn0SJsTEz
tjPocSaniC4POMQibk0NCDh0CjSooAqxHblnf0ASLCDiTnlvcvvzEnjZGn+/A7D+wRvRN1IGFcuS
u3bL5i6M5Zl0GiRskgvG2z5Lmqyk5lB2AaThBAPCCqOsIDsk2cm/xhoMCq54xirCeIr73iGuBVum
DlC1p9/sSK/bQolGl3mQqhjdBTzpTx4y6DElrg9n0awyWdK90ermucPdwKvGkTNHEcp1UtvxyvfF
yYWwwRsi6KMk5qT/h5VshGbKiCi1LZjOEw1ReufSERlKyBV72s7ntTJntD5MohgIGgyzJWGQTM/2
BaIUdLPmlTKeYY/FQq733c5L8bP4Jt2wV6DBiwUWFSgTekpVUcUVk4owLQ/zY4DJ4nEZHpPllME0
vMZdABRv27gO6bVhWpHNE9OPD9jQlA1IEJzA1QoIw4cxsTITp/8l7PCV8rLkortqhlbD7D6qNhbm
qoZ2JeM16HR1VNnMxpH74/SjmtKAho+7xKpff3ZypFq+wt+6yAolknC7BZCcXtZjxPCKeh9IGOKS
hNMyYskRxdSDPB9xf7X4xT8Lps2iWzyWkoseZ8OUIrRiayswaRYZeZED7vFxpBk0gi4tDysV15nR
uHvVwyYhq8YmXfGisv3g8G4DWhOAdF8giGs7d6dYau0h+M6GitrARS/LpDtx68EyAsikNUMp4jK3
4fyjqmpsepknwmGVGUO+yJ1Dm6kRa9zxoeu5arkTHLYxdPXGARwRgO1G+sq/JmwrKQTpqkFrU3HO
xfs8v+xoa8os6LWJTY57ElXHDzlXp6leAwSbAKTs7vdwSOweHzGPBtQDrw0MzQEpz8i29trtEvXG
Ou48mA4TDqK8/VWvLS0VLDfvDetyz3VbyERctaZdhQWOzJ08ZikHbJf+gE2cr4DVkpl6g+vNwAEd
yJNw+sv7G7QuMQ9Ky42BR+BtG5/vO34GUaWwcsvY1nhcp76PIL2SAblsaWnl+AGYE3fRzbsZMgvF
pTE093DlZyhIZyNz4tESizp7lXT1zKqfXi1HvK8AK+D4MtS0wE+TiuAo2Qu9ntrznmoPFEEHMv+Z
Iit5JG7l1miRycuBBniXvnE6UQ/vaGReecRrvTaBna8aYp2wPIUHvFlLgZ9RUHvqu2ueC1fE7wa9
WKiBoOft61H3EQQFDwSk4fWmJ5MQjt6XTRj2f/pobjb5BA4uhsoPjjfvBj4GZW7rBBCvE1S4ILRW
qZiPz8dFed8Kp9SxPfJuqriw8ANT5/DuvBMBYRkF4MZSrS5R5uGkAlGRcEXlqC/XyEoaUKgykTCR
0cQn+UuT3f0Vq5OqWWN2Qly+RoLjwAFXZ/cX7JThLx1lEjsMLEJJInWA2/A1X6XncacZS5hNLI+F
eOcZHNg51o+25sP0vxXh8uonDFhmsd/P/pn6jQVrdCwS5VEoCnJIdn15mt4GXyFkzkHGIcqoHdsq
tnoA5I4P8yVC8rG7ZkXulB4z15z6MkH8hbBnQorJKs1oZ0bImmxe7LCtGnWYgmImF/dYg7wZpKLv
5aEH75ymZ5Q3fkSKhY0gHrB+GI1GIQO1o6RoVpLPzPI23hLSggijrTVcrlai0Ce6u7R9AkeT8Su2
MNUZCtGa7InLF86n5UebgB22Vo70E+7sCpnPCmy92REtZ/zbAYLGWKbu+BS1Ma8hT2x2QOxfLo9Y
eDplHkqItUWM5HF4gwVhUaQU8A0PNqnu/2R0HUjukGaYHQ5IyShXgoCgVO3xdB3XlK6wpXdeqdSr
Uz85NMl5sJU2uVczi9W652FXI9rLZzpsieE5w9+DBy8dybwvDLLd97htbhMUNWBYVoke8vBlNVvm
okW0RV+KB6VbLYmnji9AOGL6Xvg4exwqp6zwkC+JsfBPOszkbDbtFsKxuZIX8Bhy8gko6qasHd9k
v8MBOM26XAITB5meDD4WO9M7MMYc59ygPC8IfC+uZaHs9HcUIKWdYjFrfFkjEsDaZ+cO1buW0kiC
Ww6QpBizL0HnS0mvu+Z4USFfe38bN1vwfJz98jhOVSe1ZTpuNPjv+GWGC90n8BF+QMBjI4ruY/d4
wTavYXSbOic+LqXgSQ4xe1mpmVAYUF6AIfA64AckhgYI7khpiO1nWHxHrE2c/3Ose9ZCGspuv3Rn
Oe1KYksD58IRx1IAqYi35zCGZK6GP/mb2Eo9KqivCS3GOETZXdVrZllXpreT5MorAgq6lCBlgdAE
f9jwYToAacrYhJOFTjfrCCVlSR9hdUPeuUcXbU5/pj3W2yTqilj/Dvv4elYZ8oUvSh8BOOeBpajU
0Vcadv/n4NlC5sSklaBMNslK4nPuQ2w53jgL3uuEbZiu6jCUjuK2Y1FxfRTUvITnV4KKhz71gV/J
6rzdpA3CYYSMcH24yjDbNLG16w/o6S1DlTDLIAs8uMq7ikILoS+IWXQ4KTlOZPl1r08aD0cf++QA
LfIA6YullHmvQUJa2v82sSkRLZ1lvDMRrOhwibCsjIN4hLBiSscj1OmnopONyLKX5B8qH8akBy0t
v+/QPU5yVqcM6QqLEhwQ5IPuLkE3i/qMFxgby6dZVqoj3uwebbOkfplPFKMatZLx+cBy3M0IjyC1
hkWdSjIqC0ltgad353QltZmKdnvBhK8irDNlqbLza+rFsW4W7stMDec2PissMSDB4GWl1fVEzL6J
zTa/7K9yDJGsUwGRpXF01uS3s/QsL6RXlxbhztEOmVGCEt6Hb+EKkiJUsRjpDrzbyizaq77oK6Km
KT3PJclhWAX3oWpF5dhjn7fseqMEqaevlRN5ZKpnfObABikigzhqX1NyXlh9lfZhWJI5UZ4NVEBl
G0e6OPqtD1UgjnRarbQH2Q9Ywj5c+CoyxEFSpDclZH4L/9+rj7WU7rYh/WnAnzQzGwEosSgHI/Tv
SlZ1V6TgiPRZ276+24a8LZKmQFsfxHb27bZS5dJRKgnvby5BBqzbQvxRoThKPP6Pfblc4E1cuGYx
huftEeKtMhj51ffXWp4ZANftcZubkvj9Eq0HGbo12YMK49iY4BpautNyplyvTjT+J7XwUZC+Eo4m
5wZWOzqNXiWg3mTrrMms20efZOL3ZnrzQqlTfEdWbYTACN7Q6tvtDwvqpojElpNaMdAkMysFFCAy
l1taJD1zhc35EIcvfAT1rgODNvBWmrK3DeHpVWIuw6ZMCw9pQ+g2YklKZCuVrd92eSqmHcT9kUCV
IvEouSFNsGX20wGCWTmpqq1rf82gBKtNO3IdV7TwlWWxysZKYY+PIHHEBIH3r/jXsRLsPDWFg137
4qo3HNHj+eVvxwchW83Rbej5pHOY93823DXJpZXirspNLhwP0KsTnKISWNb3wqnWSi06/euCbAN7
rHjOdyaPdtZFab+LN6aRfpcFW05Ls4RZYLp/TuDX5qMgLDvEzLjcpzJGCW2mPBse1dw3IPlL59NM
8XKEKkSkidB0KuZdfqc7jDiLf54itMSukZr1oFFCpc8zPyz62xK2ih4c7gq1uPBJXqowJrZUUOcO
AJG8518RlvRDAqC2w0BTCTdqiNnE1t7Fj1/jo5tPC7gk9XKivb+BFggPmkzTPvG6ib7DtXD/mwor
n/H50HBxfj+LfwY8RG1gBjLlmRl1UpQhn8LTi/xiuy5czCmcAm9wCMtTVdPxvTq0dpjd9zSpBz91
+GfWtrvpJjIqCHImDXcyAoRicDMCR6ggNpoRkXYQVRxSZ0GCcNMS5CnGkCo9YkO4BB+Pd/TApQ15
uvJnzoJDIzgZVpBiduk/NNTi9W2sJOq/4SWg9cjwbrJYuwGJSWNn+fQkNL8SYOOdy32iw2ZkOeWI
9kqxZstQz7E4/shD4m/pGdDrtclt57d98y5UOYN/5XGsXMfU+EA06QwdkbVZmqTEa22wu9gqQmxQ
Qr9j+QvkQcsOvOWBXuYhaNhwkkUSvaFdqXIkdj2mBZHBxhwtwjVtb/304w1O3PZm+LjOf35Rvftf
+aNWac9pU7W5bu7otikc/JvJgyIbi86rXq3JsZSznp6e4HeUYlE81Jpdpkd6S0F+P2g8wQpmA/lC
ki05UtHGlOGQF317R1ycjd09Jmg3q3dEq0YbVoxd9p1bMdjre81YgxHuVSVTaN2gBwpVEheaPF7v
eGQn8yg3HGiZzk8hp2cMmKvLQIdF4lbr4XvRG0Fw0C3nA4MI7WroLEPfXdJLIdHyCci9NukCyguC
qkv3HBQ0Q0CJhQ8TNoVeyLnHOQUcrT5WJghhqdov72lZ3HPDiHHJikrvjMpQ7WFTX8sKMBRooG3j
isDexhtrR86R70WO+45AhRyq/FY4RCp/Diin4iK4ed2tiTO7xsv1yGZ0vqiWhusDYfyFbvOvrpH5
6wiJIr5sevQQNIUAJ2BydAHRzO7xxOM18rGCty/fPlg3RWGtO8nTD0Dzoe6/Po/osjk62uq/00N7
aO83j+WJB23G/8lv8UuiKg6h/Kfvzucr0JdhmdX+iNpVzx5NCWOb4PuUKv+rkVMgN6dMdaRRiDv9
zQyO9eEExeXxirzC/TXQamsbZKgMlGfP8AmIKHCtSrx8H3Yka/KtYyp6jgyQOtqdC8Q/nr9gGmAM
aKsDrsR2eASqF4aUrx6cFcROo4uknXp7hDApnmfo1CkJq6N7b0BoIsa5y35ANNHFeY4BNVD9yDZP
P7UjaMp1QhGxCDWzGWa7bPSbWNWJqS/XModM2KnmFCDfW6B1eP9kjuQhkEVFdYCoSh8O4o7N7JRi
vAjQN+DhTIV/W2agO8jHVVbf0Oh8LrAu3CxYLR3ftREQQsS6EbytyjK99tWoiab8nMskIInM6ILh
akLZU+jxcv8k/mWV0SK+62J99siZBn1bIVYZ4QUDNzkvLsdW8u9nUICe+BPTICiJiA3nmkUV4Pnm
MoLyZoiSHkCeWxXaFbLLPvDCTQ95SJHRH8pji56Lfy022cFJka5mY2Oah6PoQ5QzjD48xO1Aq7BQ
rgcGfhadsmD8titxchj7lt8eyYmTstlntmTkUqWUi11DmwUFgnj/5py7N2muafAGfXajjN6snERE
FrE66ExYGKAw+qlN0uylb3uKWMKoMU8kWN5zh/qnw1i7lK62KN6hwgi8RX28mfvltgVaJW6g6TZv
bg26M7CzQvS/OORLaziA1Fh1RaXCjk/1V46EYRFCgBi1zmm0HfPRk33Gtkw/wV7mnPnON+XNPhjw
9NFFswDmYcWqmAL010i8+s44/h/tJL/X+yLiMK4n8nhM0HRw+mxzvLvsicss2aaeaBQ0WDjjPdD9
bSbGQCOn4s9eSOspd4QkexKk6mw/j7WcLOq+XctSid1lxDM0hpzASJ+KJtAur89qkfxAaM3FyG0v
u1lzgRz0vLpMQL/j/HDQhSF31DcFURzmCbivRjjJZeoFeYL+rt0s2Dph7Gmz8cAUl4dTHVBHhbhk
euE76uFHiCnkMBFyMKhKDWXtEcUQoG+wCKc9CATMCSORfDSvjd4Z3787Xi+k5MlBlC2TEyHxnhFp
eNZhNosAWf+w0+QXbjPrDsPyRxB+AGCJhdbi0gqnhNcsAYW5TNJjAB1DGZ6cOTnkP/B1l9PRXJwP
VOn8Kjl4ky7s70+a+l5okGQKJP2Bd/vtAlveLW+Y0qfMx7D0rfTKMZAzEq/3gd79kXXyyH1nfCtU
e5t1hQxCadHqgwJ6eieAVozLhR835VkVVCUF78alCEPE9gKf7qnB/RmsGVk6xdzwQTFs9/YCpS8s
9ohdGRz/Kt9xMiNgeWOiDMoS6ZSdrs4yRDaACaf2RZuDL8s5g8ATXHMjTmJsxViBIq6R5TuwVtig
6Vm4QosMKlltB1it7jiLsLHS1dBMDCDSbsFjztqXMEadE+bcEFB6N5TA/Y0kyGMfrQCht4bICis7
qtDP3mfRIM6qG9hOwdKjq1GPVT/rDVTFzbwa3K+5rxcKG7f1gZG7UzzT8T0nY24TlgNeUTWHsL58
fcrgA2vSatAIwg4ruQAG1N7xWf7lVcGMUnBQ0qH348OBXaJWyVl8l9T+1DVYyBs/O6tuxFadKyT/
gURsb8r/EI2u7cpMsbvd0TEW4lwj0eWux7ONCaAoWGumi0PBdSIPZK7vdWYCd8ggY53JtI61whf6
8JQgutz0bbYFxA5K6d0rw0AKVXeSY71XirCIquZ2hHd3YwNCMK6U80LQbUxQBBM+7+duebAQDnYO
bQ/99p7d34vJDeasZoYr4Q5yGiegZzat9mR28mS1+DBbzHR4u6R6BfsFlUcEOld7imT1ISvDaP+x
j38LCwuACh3Zi013mjQDuEHlsbtEHys0akqYL5ZAiZkqWXK1jZvrjSTACl69k4hPRWblwWXzqDLY
dazgy4oZkPHU44VQlPhUQ/ULeSbA4ajD9T5EtOxY5Xb/EyflXb7nQDLt0jEaVBWTf2z9EUz17SBR
qE4F2rHEs7psTfm10Ta1aMdpZUTdZleZY4tOHLJqXMXdJZFvxJ4GoFlOGIuIJEwMODej+MJtqVWE
dGsbmsedNrDH9tJRHWb7lklKMc0W8DVSTqhLVGcan+Kcjm5XMoAYaUWMUtzgQnI1uPfElOs2koej
EMfCzGo0zb73/FRj1hvTSviS81XPoOOIhT6Cp8i+AJxe0V/SkDDSmBdEaidOlIWhwK8Z8M7GvAEe
vnNGavgB9kg4u4SObVCHboacGg+LNxuGMGUFINrd0Cttz2i/OEQ8WHUKlp/4k38r3iETP7KQtAzg
c8P9sf2mdTLz9ISpHNAWRlk1ZWMVRmgAjew/KmAS647B3+gf3clr/vNA7NER8kMTRMvfjMxmf0Do
GwP+DcQzTMyf63u2em0ygHKXhLR4C5RaerjC1/oJftmHokvoE6EZWLWyKBuFTh9YRIwo1SjR0vDj
pxCnaoH1VQfpnC15VzUqailoV93cQlasVcB0ejMZ87m0tZlcVMHR0r/PIlKYzXCOU9l0dk98S9mS
YDhEomukDsIyCjykmtzVwjV6n2KatxyLpqbhXGy0COqaYMk5M5J95aGzTUEy3dwWESn3ySwCPXFx
PbCV33utjasgL0f1UA2t57CdlNza5xi+dogO/iUarQCFSON0nxmn9qOPgv+RxG9JTxnRAql3ylNb
4CkBVIRKl6MREwJDLrerXOIPWket16ofN5s+7E3s20xvc0XAE648eYz2XhS13mtZSB1bdNN3Li3P
Vdg+sw5BNF2FXTBX8/JUuxOlSx4JEvVbigBuQsGL/de/Qrp9XBPEv/FbP3YfCVtpv4Wy9b/gRIQ5
l871Ypxnm0hkzwWd/++v2rl39UVrc3x7YaFd32MT9HjKQam3qJw1p3AZ9QpSiDpaZAK4Seo1Q31/
8HhcJGh+PR8iyVWTyiB/HcTW9Vf3OCsHnBvzxX1ZlYP+4j9X8GSgc8zMs84nE4Z3tutlTAwyos9v
nfXAklqv2r2yTU/Pk+Re01CzMPFKd/3K/i01pJnavpurBZlDeLGgxpKSSZBslEn4PTdqnghcU5mk
cMdc2xLFTkJRjFgy93dpVv7o7WkrROKrfwm5xJ/13IZCSZJpK6ehWSk+hunaHttIym8UDvs9PEAA
MVrYkekh+Xpo3cs9fxees8IQ9+fHYudivos5Rlapfs+SlNR4dUujekhoH/edILg5SThrUnONwE3S
1hbZj2DPtQFrO7E4Ncl5YzyxrRWAbWu8L/gLVc3giUlKo5z3dVYWHuhYgMymQ8rABv+OUabynJqs
zlLrJBsguJESgtJRGn3/QLg0Y5miYpFZ06n6X1/TIIlE6KLJiez0mOnRQWEwPTOvfZhCkS9MjmiF
XFJ/PLD7zLN2hA5CqmfFfVB6BsCol0pjRUsgk+GxGZkXLri5AmO60S47QbufvEl4dUxwhTGxD440
+y3q36xJOndyobsqgL4cXIP0GTFn0AowHO16XZ2WarcN9BzlybjOTdYObucyyF2Zn4ZGZgBrbD3e
M9s18YWAsxHtU7jnYo79vQIgWO9eQt9q04xpMDXL3OFNNHIqx2KXdtFwYYazFkFk5GQI/HvYQOSf
yLpmT8nStyNX21l9RB2VpS3CzAieTs6CxDPiPvsED6oBzdLzm2yg1cq/ufTz54+WWjxRjbOPpaRW
/rNjQlP9Co8GdDyX1W/dyHvO7hzs9t+joqU+vyTa692QU4Itl+iDWCcSDuxpZK3C9wARLKla1JgS
K1Zdf23LEkB+eQ5cfJMjnSlGn737ydIQ9eh0ibH896mFFxCfHHyRNuL9szjMUkostiMIHJAvPIW+
uzNbjSau2ZO2BpglRdqsJ4TmBonh6fSQcr5h5BZfDHFN/NjU/PWLU74P9CzeMeaFzSRrKu0hjnXE
g0+mhM30EYmabXKBkg3IBciK+R5A0JDp/7TgdBcWxgP6+PXlJSjk1vmB19gkI18pSnyZkM+XxfEz
hs0Ikba7pfH9aTT8+elf/h6F+9DLOuRCDRQDvHrPRHbu5wsqGgODK/nkQsA4kU/cm/W5Hd568QgT
ikC4QYv4tlbgFiIPRMJ7trII6E9R7r0pp4acOgdcUzWaa6Ys9O9+obHC3QEImgQ/maoSptePgUF5
tw24RujJIQ6bMmGx9jh+kXkJolLKQEyTdVfOZ5+eqjgZGFJrVOgjLpjOYk3iVf5o5SibtLHfBqnq
GWy4kH8sZsGuutFaDAHyx2eqIURQQtxIWDIdc1/jUbOCfNFRb5zG/a9x1L24pJuy9okLbmzWKmyI
bMDY0CI4FXlQ43RIxigYg7C/pO4t9jcwnD8Rg9biK1DIZTGDH7kHCYbC0w9CeTl6XlX+dQq6YPz6
BlFmLW0juZYVKhtBajI1fh6fDzgCVxCiI8Sj2fNzo512lAqekcoLA60NlNVFt1RYTRHYtIlrge06
/3/47dh6Yca2GfCPdA29vmi0voJp1PhWPMVrU4H6Ox0RNC1j39YLN81drJxnCsTRf/+uqY4V0vax
e4+oZ+z3fGg6uC9NKmVmZcM+Ldn4fMGyD1BueiWXPFsz97MR2J21aiVR2Inm3cmaaBMfCQT3T/yA
xnBpwnU6JKQidIoaZLwUWGx4PbTV+VstAj1FNA8FFRJdPmLrm7MfAAGyrPVJYKnMYNI0H8MY3lOy
bFv847rfg6QCtatJY8uAEzQH9++Reo1necuLWhgwlAO5vsT2Am7iZiSPZBDl3rQxU3pQpg74wcA/
asisxFS23z9TekdkYw3/dQhxmiXLZwlZiHb7ZMNegOf7iEFSdYh+EXdjW/b+SC2xLF+qdaIP+94U
YBn2xCZxYnTf9XWzfzTCAGlmmuGPewQGBDs7ySb5gGf1b5S7ANJ5m5/gngh1iPxI23EwSbzpsfKm
PKsGKkjPwLYF4R5N43E0gWqbngZBXqUhKyZfJGhqwUlLfx2szlpBjpoJdAQEDvwV1sD6CF3rZU7c
XCdvwazk/NZwniADDCREu0E21n8McRJ4luCdHzxSBka5AdCIclguV4qQxuBtAFobSSQ51zOvYgMF
xwmfjSKC88sn3MmcMo5EY17RROj/esvzqKaE5Yw4KDF1XEaOIk0tKvtQHERAU48uciCwFEKlaiGW
EvUjFIiZw4TbJkK0Kk6ajI/wmA1/id4XFenhlf3MD0WMb+nJSFfQIwN5oxLnFz89YkILBW13E0vS
UkRON7oAwsyLyJkQSTJAB8TpLB1uKCinGT6kNRNnY8vWThldd6USE/035f+x2Wxc0Ed9Gl38EmqU
fIzLGMIlQafRVTM0+UzhAglt+QVtwcn5hVEy9O/m5vwqzjj7Sd0/R1mdaOjIR/xaV0dhIDUK8Zkm
T34OxjzZDdQuUP2jgxDR7ZQ0CzDYD47P4Hr2hTWGVoIewsAEwx8dEA7HE9GDETOtfrg7dJ6zoY7p
oRBWbh2ojXRqebJwTCE7uJoESvQ4FfCUZH6Smi3kuQGd3v4Kf75BPS1L5GPpmJ0Wt0HIR5ybko2D
gw2XghxySyIsc5bBYkislCUlKb98wL6BStdJNVNkAgYQ0OzrVWuKA8IBxVJ2S5AbW5ypyWmHMFf1
93SwBIhCsR6Ds2+0gywCDPNnWiNVC+zGF24Ih6r3iDceEXU9JeIf5j0RB3biS7Y1xKg1CneRBWkG
V4gJCoTTI2ITTCHbNhqBZ3pz2Tfd+j6mjc9dsUPzIyRZBmR/nkfvTCJCaOtE/lL6yOK+f+vAaB8N
wTjKhW5gE48JSqrDT65lmobyFqOmn52DWMKD0I0UXidOjQ5LHqiAoQVmoyxpKkmXhD44hjfrOp2d
lkBzqy1TDXycw5hqM1euiJdcavP8eLEoA+iIE61Gf/k7F5fhr+40BaB5r0H0GzEkvUzFUpg28wKC
VGn1Evx2JOTOrsrzWkQG1NbpH+uMLT//berYQk0NRMyGQkcRWjCMU7ntj7jR0WjEv+2v1IqlOFnj
APsFckXFyedrswaQ+TOsf2wqRWPDCktAJNxoVpvHcSR9rAhSbwkv0aRHx34lnNnHc4KNtYmSkRwW
glISJnr1bjnJslXiqWmxL4U6lsn++PgrROwiPnf/iuBMmkPdB4rRrhNMG1y2YKol0Uo1sSy0ife+
9iIs1Wa85/w+1v9OyzW3t2Vyl+jLk98FOffpQXFRiWHTnf8TXRSJ4IpHlJPzirDZk4hepNsnie6J
1u4oK93WdXJQBHrubfHdsrOJCmX1DZUw4gNrzJvKGmqUZjE3XfIsS+DU0w9X4ZvZYWyZurXL+ozi
s9SmNNL7EkRUe13+L81m0DRVYUC3/2ZxUmKHNwYdmAzwmwGYDiDQJmxGo10XVOSBduo+5Bgz2siw
l7zen0iq7Vqnexe0loqGyIwsFdKdPoN3Dzu2U55gztPLMBQ03uyWW7bF8Egj4Hparuji8Faa2ImO
CxmeJHuE49Lmd7c7iWtAptEftreafdESuzJ6XM1zKX9Ggg/nJhkgL+FjK/4G7pf0lWuRqCqFbADo
k5ZDUFFQ9hDU1YQz5A/IomQDbpGTrzW9K5hUK1nAvsnu2cJiwLP9OWQQdngLWf0+h+5R43GDtSjW
haXuPQwuslPjXEJUDIcI/gagt6XjbugNF5N8348WCsUuodiBzgRTVaGSZmdeoRkTV+T3xkRe5JuK
9CYqRDzHAgkvIqLnPde7Ab61kCl6U0pRSSOpKvNLMy9SgjeyoRW79kdYZEvsYQ0/NCcAcbHFJ5Lw
453BSQFh6Nrxk5j6yhLD+JDAboCn0D/v6TUvrFkV3VmSUN1Erfg5Hvlk54SUud8VqRXfe97nP5ok
JNmdqON9UBlv2KIRgPuKIjX82xnNecbB+72SVHxU1O8dHmrfTJKxeSu/Bo85sbUS2W3zSLyDHhVV
7tkd3IJSbKO/1CgaAr9pnnDztd0dGVPKvQDobLO/0k5ZJaoIB0TEMGiXG8PSnB8l1lTscX6hhuoL
NFoMfp6907h0PQJUXIWCJEJjlR1HBu/t8ggiX+C0q37bXxJlfkiTEttjr+HKBJW1cL0x/CnoVaR0
2cYxFsaR5VqpXoVzfHG+tthTIsJXSGNK1JlVeFZb7g3hEdCJsK0Dul/u1xf2ElvGHXnIA9Vaw29G
W7k7BBOhIfp26r0mDyMzUobvBgKCf2/MsYZY2d5pJOH2chE4zujNgZ5y0T0+sR5D7bB5zxzoUf8k
tjxMUulEnpV/YGtqMZHCj5Ag/Uuye725S8O2OxUhBdA9fGdonhR35nmoyc9QyGH8TYNQzZUWXl/t
ox3/H9db/YNHpFR+bLt6wq+6h6EYBwfRgMfQG7dpEy3xqVw2GJtUK00N/7xeZQZBxoIyEvF1qzBK
K16qEIN2AgWc3nrxwP0io4ZN5ayvRFayrK5p7CCO9/XrYhFVGsqfICM9N0guAodxmrWe5WdWnz17
RjtRaECSezF80YsbMtLKVXr+W+M6QgA+8Y6fYhBytmnhM69hfwwhkOtqunTcgiLje5VbjHG8EGij
9rNTlyOmdfXzfbXhOJXT+vmQtDFsbWXX0wHgZeMsaUmMizz075htSvWz1Dt9AQ7ZXGz93oSkQDNr
sIFY+EhZASaH4zFrIcjDaaOJC/2wH0PAW8cBaLOPqkdvFd1o5lzmLOQKxvWAdWZMlrU+epWQJCJg
5RnyxvtcWhiNCEKmshJRlE4B/hkYyGw0+Ct0Yh2t4GLnQ/aaeo2jnal9Jd97l+ArNttelJeyyKUC
l5Z05zqlpR6edSGBQoLKEXy5qkqROmliPMh5jxtn65HAZbNSXwr5jTN21SB6Xg4o1bjWE9B/JTj/
EYTCA4sAiWiWrLW+1LSesds1MfJctiJfhVZNpdub9HJNGB4LwZW+j4v+YWGxL0K9BMGS/mUo/qzP
0mehNCieW3drmTmVgUQVVPXBUXbdJ+wFxLrVoOSNcoieuVXbEEmUmbiIdD/gPdWyhk6HOQxc4Oi6
eabaOTkiaM6YpQzBcWNXcv4RRjAWxLZXVCWdgsqhLcPS9KE0xMS9ETj4UZvyM/xvWqNuquoaePab
76hLj2CnLlCoQDwpUdY1kXt4l6LIa1rOYgE6plBvqZYV6wwHVQqKx/CvAGUyAOAVCAzIpZh8aXtX
TxdtOw7lesZhoYbi3lYSTCb7eq7S0WupQ51sGUEvr+Kt3h1vyJMgWOfgXqhyVaNFfWwzn03PRUQp
AqkZ7CIrYIQ7RMRJmJQ1FWF4dfVy2GCadYZ7QcKqXj4fqTigi9A3+sneiDhGG7KvQCVgmw2eXA4T
emrEXXez/sR08ChbP1ImOQeiA9C5vc+BdiwGIewlfccmTpSS4dp0Lx1jS37wCZBDNqXqQqeM/vlJ
oHVvvWTjHjLI6k5JS8eg9lBxUrKOdGKxwpoPss1W3fWEEel7O2P7dqhnqC3yuHNT6rr1Ttn5pOuz
cGwG5lQA27BtaPlwHdqoRmm++3dDBtp3X5xxJ70fKKyjjF5X50tXwRjlzeAJt0eUwBhHCRU9bxRu
QCFZ5MoQIknzOzfeslHr6l97GAncTY7WqtO/9wX8KD5wenqgh/LRky4ZdInmY3UoPZ6DG0OUHSZa
jNhxPukbejxsZfexNNdJJhcW+0VejEPvC6o2oCxiyAJXRqqsQXTEsn7NrqLvWqknBflNoK9oFE5P
/nWukfb/g2bktmIJ33PiNcdq0AOZub/6virROKzVKPH7Q79TpVm5J+u68MXOQtdDn+ERWb9JmJxB
5YzLBVVLY7hRtPy/BfluHQ4Bm7R5lVi0/kc5AoDoTHx/lU5fOGu9Y9ZCcmtc9HWBr6c88hOYdkV4
w4RYyC5Uiq8LacmU3txU9Rqi/wAI3kVAF/7e80lRvU0/+p4qw5olKKMWx5Rcs/qULZmQttM/9UD9
wZ0pAAktK0EQU27siCrevwWrpzc3czRvMvETnBKD6IYAi2KnKVxMMnWGD8GqeM4otufcCMNAR6lD
XshifvGsm6n66WBDZnVREzMqeFal7gQMeHSK0xZmXn/GTo/cLYKLjwG+2w8nYb7J2EM54fg0aWqk
VXd54uRb9dKJPnCZCMTnjXV+6vBFfXdE5CtOB1K3GXNAP6/+3UkU/TM8MKXtJ3dfrWG2CIybLgw8
2SP5pwxxTsj12KHawU564GdECdKY8LphQbvFu9woR0NsZ/ceMe6ea13A8qMOYbvEEmYanWC9WN80
/0rYl0X6CxJpq9zemNKk2BBYzUSwuM494f3Frz+kuh/GocZV2eCqVpvoRAZRKzSBZnTm4DRt6jB7
lfA4U+4B9jliEpAQKd6HtNO96ECXEWhzwIOuSljB9QfrI62+UFTTHuMXpEYTPrS2CrFEE8PV+KQr
FLj+pCUKqiY4dv4E+vyT1vFdMfGQLdrobN1sK8JhVYqPh1SQF+wYIB1uaLYzJTV9dQkSQxhWtz8N
bmaeOGmNz2HiN+z9ho8Zt0wzjQTWOxwjlhWmzT1bbxbc0Gyqlekb+KDcF/bHOtJ+g18igvBW+jPE
+HE65MF2Q44fleqknwAQdEuGBTqGey+dVwm9fjINYytkUMp+WBj1ZNqTstDkX4oN8HHP4WDWA17X
Bfd1UeVnLvevYiTAVTTxvcy1DjSv5FikX33Tzk7+/hw06SDR6ctzspWd7df7FfRIWYCANsyUS4bU
2n3sKJycom5KgvPYzYjxP9P8Ux9eTEeF6MU9Y5gWdijZFenVobOZdaTHrSt5ZE5fgl7t9TqkFe2p
Vayr77a3cN6E5tTHRojM6upHk51MNboEBctXJo/PM7Dtaitx+xvU9lXYdWvo/jGgkn1Ju7bu696z
QS/Wi/1a+y72LJAJfdoXtbju28rHDikHlDggsQvQJUiFkNmxeCrDHcEOwdY8yT0CxulmXvkJ06iR
gTNzqsaHEv6cu7NxASHtYRMh/1jnKxk1Q8cuNHxwt3txvEkE4wdo/6j4Crg3E1o2mBHXKVcHgHNG
pqTpeFpEZGc0V79wWkWeK7WOq1uP0EViR9BdXh1Uhw/JEnS5PZxalUT9ne2dqeFhAqChFTDsjWpp
K5x36JCBVoR33wOVgStnxC01v1EUgFYKXFEdYrnj7m2JvGiwIZFy2DMlHDpYTVzsFIwwUg+jdr9x
3hwk0iYe2PyDskbS95SSmwTCXHo4nHUK9juUYCy0vH2iRo8huFwuguIXO0F2DcIWtP5kquU98Kgr
vuyhvl3KCyq9MMJwT2FkIeZuayZ+2NJQ391mCkYAAbWUnl7ooShGWQ+auA0Kv70gn3/yaNaM+D8R
FWImbxa6yd5GaVXJmmzACZJgTdPb31BWULDjtHyfzadIf6HsPhCosR5+Zud5OqlND12/5TzTvbTW
mypYCfYYMSmetlOft6O7ZMCo4KTKt7myM52jOJyIXcWjoxvKYFMdEwXO/cEagEInjC4CPLmZT5QK
HsiKcGTp2tG8Mv4EXlUbqQ3lt8+K7DIK33WHwArtghsLrvu0szULT9iYKJqZNH2chGmjedWfu9Jx
1OOTiK1unDB9Gj3VfUWAaPwuoz1sXRc2krFIOd7GDlHHEOnamvixBj9aTeDwQLBEiSt4HY5xCJ+K
2aCLgQGqy99pVifYVA2EH+0UEi8nQONQY2gG+SH6OcBVUh+Txbudi1z5Lx1axa7tr5jYyZDy3wWa
0iaYW//vsonSADZcCQd83M0/Ozup0Oqxg9gnDlm53HYOMGghPq/Cz14cHFOFRE+rVF6xPkgc182q
+exWIKHZhlsmkHHooc1STyRrx1I+yswZ4b3IFM8Zrbmwr8pLbmEkKD72OUk0cha6C8QICwxqDywd
TPHdk5+ZiDMhwA4ge3kGg/LeTfAWkol0jTvQqI/MyOucnWXs0KUGTrzdBT43bmXxNR5zXnnzmXyp
V/5SwQjKQr+yb7VV2O2vOh8Q/qbDjwxiB2S6InM/fHM3fPPI5u49xRI2fdTTYy6SwgNc7i7ji37a
P3kBtkRE7BfN3EylCgxzZQjHRJHuwPM5BoKkgSWlKa6JM5ub3NdUnArZijwwvdM69r4L3e021twZ
NnXUjbsO7GGwXMMljunhvf+agqv5NUK3waoUK2yWfGMQs51aWsIqNHyo6EomdaswNBCYPF3dU6Oz
chQezsSfur4Xvtcc8Bm/175F2dOQWfsGVDSyohVpkAYqVORw3Vb0Ry0II48L3gsQuWKMzO+51FWY
Tpd5Esgx75z/fRlFff7pNPZMYqj55ddw5x9eO6kIoDOfCalVlVP4nDtSmfSVc25fUCyJQuOpWFpA
G8NdCZAYqTNRhHf1v6PWZgSafWIa5qxRVoUK2pVJ4fsA0RcvihJhWz6PXp5CA8Z4VUtl1o0Hfm94
SjkpDuy2UkIdinRxQbOhDF7AiiRGTOaFfAXlKFyXKKrRFL/lJcFFQxOGixWOLuPfJaXbczdn0V0B
fz+dcgscc3eqSBzNEZEgxMO1nqjv/8f2xYH4UyDCdLUggqwJ12GkEFZ33uIh1Gt//VOWSAOJKbx8
vSwosTwH1GOp6o9GJMUJUI2TvLS3EL1bWFGUJeNPHgQ2cY3GtsTyF3wHYQY8ISWrnmZ8D8ukS0ut
xXS7FE7Ybjk3intnuaQ6DBJW/RsWIlcSieza8+57g1l9FPO3k54tvY3N1alPeTrYD3VNF3ehQSkF
hUmhfYjhuIdPHLCMalWv6FZtou7vSaO6t7FvSOan/hyHn1ghus7bCEJpvw/Gt4Ua5m0hNarnR72h
ZLzP/1uq6i7hGpgZBh97ETnQMRiaYY0h0gyn6PhUC89O3Hrh10bwVxgaWllOEfMYpHSjwgwnTXee
lFXgY2/Ldgf5UcA/YlWTFpFE4tLiqEA8rt+OxWbRdtSq5rs7Bs/mHeiLnSpQnj8Hk/2yJjUFWEFq
M2h6WFEQNkH2Yh41oV3aTj/lNdwNnl31GxXhwmZhGtagi+vLui1XmJf+k/Iam8T4ZMsEpfUQAwAO
5CVl1OguuQA2FC129IHUWjoJayFCf6JQJDXIALkWUxip/wAJpwOsl3le48XuAXCMOzLBBbKwxRlk
3uzV1C997wtSMCkZ5Xu8UZEibsRfThJyrYQ6DxrK5ynfZCLBFllzkNa+xyZrlsiqdsMp4CmPEHse
w3SRwB4v55SnhRxLEnkxNt4SxxE7QWS1NLZ/jj287IJ/gRn/SyaDmh8teFzCoBQpdMQlA3mbHEaI
N2d9v3hU2B/flkCSA/7b2I4bPmIuppE0MAUYt/+7Cp7xJ7172mrXwWSLsiSUlhzqEp/r+C/lCygD
EgQPNZv6fHdjKTwvyljwMMsbjyU1I8dhOJcPloa72AKCQAMn6wLxKfoBighVSsYdj1fNizO/YRZr
GLr+cFJOnPcXtZkXvJp31pcUEhHyy9pFME9Hm3wSomlPHQYodCsEWoY2ZkXEqKaxFtLuZSvjGpj4
eqJKJxqY/PITgYbrDG5LiNt32f26XuQujs5pvxN7g8YcJL25iVGPv9UMXYR4tV+KxP4Tx3fesjwd
tWPZkDdzaDFIoNyvouG5BFt+CbvFJBfaKiA9Rz3VjNyAF/BAx55KTivHh4Az1cYWPFzQiHfWOe8r
RspW7HoEbnXdNa241AV3PPPZM1LiL2z+n5TSjccI7DFM6rAxsPLcYuN1saWZWFIsksa84J6QKlru
G19FERi3MAZt9fc3Dq/isgiLY3Q1pFqVpxEML+5gNj5/YSeEJnJF6zmG/Yosz6fx5SRXxkqDx9Tt
fKTJx+K2wqaT4rOcbxHYMFYnNdx4kMC+FtddI5Vjf9pz1ev26TNTYUpG09waHALTpxw2ahAM+WUA
5H+nM8S3yiLDKTs9yUvoOmYBU6dBLKfwQnerDYNcXlfG+MZoWH2Ddq4g+i3/qyrSkAlGLeq/TDHu
gnBzh0VIrYrRpkUwghakU6GpJ8YP+o/1a2rmrnROla4SqiMayhH9p/zHQ+MhBPdXR9/CNEFACsm3
ylu6Ga4Hlfi+e+SWxk0frqqtnmKgeOn2iRMHfD40yUr/nm+7Evq1V+qNTFvXcX7yWgZTAKrjIMqB
PHgPGxz5wZMWnWvmvVRDMsXZD9ddOr0lw2BmqPZGw3zP6pq/xLvsbKG/wDSYB0daHRNcFT3JSuqd
+1CwgWOzfWwlC+ip4sI7TaJZQK1D18K6BbZqsbC1E/20FRRrB6vrvmCkGXFKeSQZ6hNSmt1dNNjT
4Co4oEXkvyyNIDm2T8Z0vHOh3NIUaCneF0z9ZO2hZ46rmm9HdmyrSQ0bfJ8CnQyzUwditx2Tq2K9
LK/h/MW9ag+uuwAbrZO8PcliLQkhDth4l8qRH1xML378LJDQx1d2kh8NWOcdfcf3vQbdiV55Lv2y
ahvPlgGN/OvRijTGQ/2L/6u89XiiVE7x8AB9cEoFIewtdZHsp76Z5H01X55lzxxl3rG4JvuoSFh0
XDEoshTrSN6bak50JqoqQUOiCOMqOQ2JMFRopvCLqtVeDcEMmpBtBpXnYRAP7CXkhqihpbsKP4uV
0ZdvEWmQo4/WjmAULN6KUITao2ZeZpBpDvk9I9lghakfN48v4cwLsoSdjc+HtiqNrePxlu8xZ+oK
QPrwvXB5aQLZz91IwZmYwTKSBhV6eN/deuxFwW1vXNPC5VC20X3hG/MBWxKRVtfAFn25C+RZhIuZ
bHqJfoC+wechhZh/OojYdhGN4X05miFeGZzu4X45pvaiFy65HUB6uCrjL+bUqnb5Zy/zvtIp5tKd
tf+84YSCuEJZn0wsXeS1cqi88B8QQpcSxBz8BwVf7j97FmVXc2xHnz4+hCOS304fRnLJBUlfbcx1
x6LE2WXwoLPQcjn5Ra+kjGdZClW45snskHCP7XUOrtkTH8K+rYTWw7AhA77Wm1j0SVNrgnKsCc1m
CAHuN4ObqPtl56FmU1tFScyy94nQBo2FBykaTUsWstuoapaTByTuiRPY3qNamlge2KNgeqt4MtuL
UdYaTvXWHblUnvxNWa/jva+IhD8yndG4QSiCHSlN8LPQWb6zOEg+Jw2OXa3DFv8AFX3Gx6rCTRyq
z4RiWYVKm1acRAwdS2CfL83lC+hRHEgkp6+nVuCFo7hZ3ZC+hF4radS1fsnLoC0qWirvmvZrpr03
J/M00+SqVzTsHY1e5PmL3TlXNs/WZiCSs1qSVcA4AHyg2kSULD5KjaA4TUUD3JL7u2Qqgt5xCUvS
8/mZ42Tozm/ufz2AC+TfoyZmGvPGk25w8KpbLa/ChLFOwTnWhh1BFiFJCLecJse8sHCPwfkLD2A+
UbWWM//a4JTwavLrWUCylqLj1uQhnAaT4X+8GpioLyV3hkPOV8tD96/CNocPIbQe1S3LizaD/oKs
GDEltF+LTyGzoqi4ZjGugDWP9HYSpiWp35n5YidEZAT61MgLX5Laj0znHIJwRBGME+HPkVkB401T
r7TJzqteYd6U93f0R8+BuAZ3xceawpHMFIjUAKRQS6aMRqls5iCSEeKwfpq+SuSYxyjYKKdMaG5n
eEM+GHi6tXiI3uvOTuNAZCUM8JFxsgaCPwduKfIgj1SmYk3V+l4R86ANxKxoO42qP/jR3vkOZx+6
6KNKv0v0kkKiCbJTQukzOuHaMny6LMJKR6q9jPAfbg5qIRbuUp5XhH72NgHLAxO4RC6ZIjYoDbua
7A9Ne/1kBWSk4YQ3ZWo4XczZdCRbmytfkKF4qtDY3zv+QsjtUXXi+3Ao/j70E+6TGNPHHL5sQnfD
5aOgNxjasQxkei/glBNPQhwOrLaenxJicMgHPN38HmEEDQWVG+ELi1ge/7SlxIObv9pEsQCKpw02
MMUMB/BSzYC8JnrD9xuN8p/vEkvYVrk1Xhx1P4QEemq8cItnTcGdY1QYQfkoHAEkNo4TPL5GSzwn
/XW4UojU75hcL4AhSbMF3mOsNaFiul0IxtQY/2qCs+iecnvyGtAUV/vmUobBEEEQDzBO4fozySyJ
1Ouk5/sHglzd94AoG8Ueg4xIR5JQr79hkMMinEoLJt9UnnTQCfI83bduKiVGSoX/12OLKU0jPLxq
ZXBwtxQTqLTzRIw3K0PuDYjH5qqK3JrLMdIyxow94e/PzBBadPLztJP8JiYPjJqVJjhlYjN5137I
aOELebkfuzBFvN3Y7wQeNEop+xMoL2ZGEUfRWZQu2LNzWbsFsBkXx2OnBwcWT7xCaQLVKHTMzWDC
DiDZCsaAo/LdUSp1jnQyCLhNaTCSAV+ErCWpczFH36KVjbavGiiZzj4v8PZSjdYIEhPAZqI/Hco1
Bmxo6FmQNHWRXviYDQhwfRQJjUAEeOTYf7MglJp/WNq5XN+wsHb4EHdx06lEgCI+1VLDrRTpHXy+
+vjXUgdG1W/u2S0pGcIa+qb1wlmoicu4V87KCXGkYYsIKDDZu3QRKvsCfgU2uzDFqek0WEPR/yJK
/5i9o98dKvKyHBJu2y9lP9wILEQrYY/g2QVCpeDBHouM/IwN8tCUYRrvO4pIQbbDtGyo5JucIMsa
CIgKNoSnwixsFXCIXCGw4fxTjsxTvpsi7hj1gGlUOSo98efA34g2V1dE+avluCAfh1DLMY8yZKSO
CkGYCzSV6SRAGXjELacWdljAfF7YGH0dN+Qte/RoOMwCIsI9k96TBqid6KFyT90I7Vnz2c8RH4LX
25nOWhCOzIDLCDUDO3INHErC1Dn31DJRMIQN19X5j5ayz4YMPa2dbLUeL548Q//qJ/Uwap2XBEgn
cE81zXVWfYnN5ftrjtN1lwV2hqFFg5gRUbdR+OW+vRFxy2hMdwYNAj2P65ft3n4Hy7Gede5uiDAH
sKBQiLckcK3YOM72Cj50ml9GvXIxvMf1R+cKk4XOJoHfwm6tVYU+uONWkPBg9P2f0tEoX36QX9X0
ubyFvN/ZpbOm0LMQ4ToVJsGkadqEoepQ4PPQAtUcxB9mPM4KTnq0uHc8T8w7foUygpGkc2oILA5q
DkBGc3DxlgrRye5yrR7X0ytSl1AO9ljFjTFhCBdNiYcc/2wUsKg+Mpss1kfAfC5PKOtBMvQNlAdy
16CBLNh1g0+ZbYSa7g2es0cfN8nGD3Zpf2WLcMwf+JUvOojq9blC4oke/p/sTE/RaS8saNnP91CV
7qZ3sWNCrz10blonXYDljpNonVDjd306+GVwPLzd6ul65DXWR+NChB/pdfcehOVBiXSx8SDsKmNm
K2yhtMVPleKnZoW3QzK4VIhtgldTZVYEQjTol/cB51I6sWAH5RtyrboTwQlMLhxVFuFBkEDvs/5A
mo5CN4v4hbieK6x5VxQWT3VFQbgMRcRawsPNVNV9xrU1GgcEIK+gMkEb9s5dWN0ETcke95O/VEWk
PhVdtyR4y4g84ewux9WlS8a3neKDd3BS/hXxcQZxwwdwbGdnncNVsH6C541ylAs2MbLxp8iqfOAD
dbsnPeuwIQpYykMjGOMb+TXgPZk8PQSjvY3OYQu64WNGuOp0ujkrDXKRpWLchKwBH9bEpnFp88b7
CtXa+yPYDSJbibPNiN50uLkT0XLglVOF2IOOLjpoP+xH8lhL4TMtNGPlYPPz3zJA/ZyA3MahH9og
WeHJg3oqz8kVAulNK6FOM62LHLHplHKFXIlsENqQocepYGSqRt21OTHGVLU1AeqMHcKvOMd3HMCI
wtE0i8AV0VCjuUR/BhIhGSTsdfaKJijnVoPmZFB+3undQcyWct8w/XLOChD7izTrPcKawLmyyQHa
eJ2niJr/YQBx30Br6rnZeBa7CvQeQA6Vd1SJGeVT8X5f3slkgI3XMIErIcZweLkJHmTWICCdU4p/
eWY5rPzWOJd2x3Wj9QmOyoOQoDS2JDG9iBmtzv1MZshvbZvEUddZd2nQZ30/DNzSeGAVJ+z/0eMD
EqBzWC66sjYzovoItX95866eDKYkeM+90AmElQr+1K3kVO2sE5QM+q60VmhM2m4Uhq3LF8hiNw8i
7fPOK+U15EK3Ztn/EcKOu5OclBULsGKmzelq0r7JYlepLSDK9FvE5lR5y9kJqDk9jvKUHErvNsmB
qahE0dLjqgOMq9Ql35rvzmgB57A3WTon1og6fILIrKstiKRK9Y30Tij0PkOb1CMSCClwES2Rfut3
GrH+sa5J9921dVlxJP2jJ64H7ULGjtoPHTG5PxhmsAafgp339LPkwq0roDAwt41T5bui4wogbu91
U1LKVwMWFhIyk5xkPQH5kH4E3ZjG5ILDZp4koqJwxC1CluZAVXh0gHoVJwA5YQIvMncHM2ZLNab3
7zj7M6LwxV9yHbD79kR8ZoSnOp6am6cj5sI//mzzgTcTBBY1e7gqjCNe8NxYtA5i+yL67f8s3vGH
Jk/F3diF0LzYo5BWGU7TxmAOAzOzQ8PMYfRI6wZKqe3KPFyLHCVP/1QZlCBL+BhfatUg7jr+0mr/
Xk4F8QF9meyp1cy1aYh+zY7MJ0d7r8SGGl8XRuro5TVfhLVQEvideKTPz9+6GQ4y1wQS4dJG+fW5
mMtfC6RpIIYnfl1CGbagctviRAaiyisNRKZbjbp/faYZa8+IVIhH977+yIHqe7mMtPIGz5yLOgM8
RNRs0ljHSyekKg17Mwgkw36RJF6Wx0kURzvT8ephEcnQNyuZyFv76dJezjJ9H55xpFeO2T0n3wng
Ro90uevqj6452QiRD7Yg18HHzhOdOoqZzcmTYTASwuoyPO7HTYJohB1o7z7jxKcC4HgPI5mjoYuE
TBoq6QYyf6kR+QyGnkBeM7cI6l/Ad6N9QseAf6ovU+kBRfzJfUj5OLFbCjNH0EYCilm+eZ5IHhw5
RWl++k88lMLDLABbQk+n9w40+PnAeWZNOX+WKB/zY0f4lURNpDf1JFeBtHas7HLuFWxnp4iO/x1r
ArZT/D0HA6vpl/555JM1nOSbv+elCgN53rrU2lQ3VHDas3WYKKD1gsazllCcoRi8vQAE2WER66WT
YR6S6MITLdnwucI8jbWqtqcSGGOc4/uxqf0DkizpJx2ILqPaFVL6Nqowm+uXv8Ox5y6CZ/9BIufw
mtI35c5Iq8b3BOjJU2FsvYQL0NkHtoBKVEEs/vRICuicHxDke+IbOBlKQZXZXtZg1R/pwZaw8Wl3
iHYq0Da/dTAIxnRzx+fA87t2Ryu9Tx1al4WZPrVA7sDWiAN1ysWm7N83pJ553f+ZkdsT490FgC4Y
826OEXFVXtVAIvI+eb3KSxFdfvIceXt0p7K2ApP37XDt19eczf1P5fFRY/QWXEBwAh4iQoG2nQdJ
QgB4fvVbYEqP10ZOUlryFq+H3Ye4n9vNRIyhyPc/vPfpt1cmvNUFGZZJsE3M2qC4Vf9fkzoiZom+
cFfmVfu3QxKOUXFbcrJwak9preWPx3KMSsILLmDb2WJfHrQtB0XCFev40ji39LqQ33k2+TwSoFtL
d3v2PQLNDZK0Zq4dJqDcYFr8CQfCJ/JmHw8dSzII3t2lQBSaL6YyW9H7p4vIloAXOMszHIoIv0fQ
w+jO8/iVJPg1xNdUjnk1mSNgVc4T7C5gqw+UMMgtfFj8i9aJGcil4TN8rdzfEJWKqV39kQd0LMVa
L69ZjZyyApjrQeTvLlg/deFK115M7r0GmW1LKWbcSA0Im9Q/fI7xSKbWxA7Tb1NuTh13le3a7rdX
7fJDTJEqjbEKnDUkIXQFPpq55ZMBnz7Yhcs1jQ2x2FffIYy+hiuYPix4AXUcyWVbi7H0Dvb4e1/G
xB6QC8MM+0XAJO8Rp2PlZyNBVE0QnaCZ3R0Fi9sTLOhkBw6VEBQU8cy8VvNuTl+lRSo32d1CVOuZ
z1O4foS1cHK3tKhmKdbGL/PUu7VW6xcQCtl9E8zZyYwOpQc8FVrdEl+y+dNbSqxs2beK8jch/Scd
CwhR6bjxaWVoJQKtKFO5FYLilglD7Dboqn6Ivlv4otnQzouSj1K04QbOerM2P0AwUVsahB1K/MkM
UPSaCABKM5RlG0W08brbqGhVpn2pwq4lCLrN5vfiUVyRZZinNjekjt7ic76k2tXB/x+ariOPL2BL
Huvx5GIUDqmMLFdyF+3l9WNy5FbLl/L2lQR5A2cUcU3FoOOFiYj8IQNkdC+mjedD0BHMXZn9obIh
nTdI0yNm62FH3f8X2N4uruqSK3JT8cMfsnVj6Kv+zOFM2gM8ptwNpq2LoUQHvyyJqpC9gQjHK3fy
VKPSm7C4kHr6bY17qncSbkXIUl8W2JxlyccLMS9mIcEEgcAGTIg1Tvn4WKMsGj9Uie6+iYJSI5F7
3Nfywb7Cz7S7I5An0/mRaGWXhu2qiMbO97pnBK61ahXODb5oVNJN4ejrEkSOpwDTcPQVl58JW9CA
c++BvqOjnXK1eqtyuIpOVSr4C/Ja/lC3LXuUuNKSLuz7XMsuRNfcq0CqNjiDLQtV5sheMO9LJJvI
70UnziQaqB37soB2FdrgxhvH6UmujBZobGKPEmQJQZOkewz5lR9vshy+yBb58fxLxL2vIAsoWU7D
83FDyzcQHBXNcjoWnE16NyOF8Iii9yz+S9kUdq3IN/0BeTlkRJoJ2alaMdY4KsAxuJReJ1iWtSD8
m+iQTPyphAlVk+DxWK1eLFgG3eWshMbeSsowvrK1oQNceelnjqAdGrw7IIPhftBDzkC01/9pRbzl
+9hICUijDzw1mq3REpyUtq9B6K4u+Ny0liVigJSs/DKvVFpxiLFeOzM/KG2+oqf73FKuIoWwpqLC
jIxcUdqu9SXs6nJUfL0BsKAKl89dIxWPwNHxlrCIO1QlxADvOL8J5KxrBqozKBMFJRDWQMYzvAAF
QsVV/vR30ABAqCyiubiRtxtsNJo+2HxsQ2w0tvTmGGf9StZB6nlW0BEiIkaWC3ywyW6taY9EQeYX
azxuqaGffL/R5jgJck3xhvLc1iqjOlfAlQVzd62xnBrhoazrKkWxaKouKmgDhznztamwtsxf0ccw
W9qcgMo6M5m0u5nC3O4rBVF30F+ThadX2tHywLrAOKZLWUET/mYFQmChVEXhkqNXrjNjWbOoK99Y
JN1PNhfIs8iIlP/OJYedY+n0eFw39JbVx96MKFy03OBl74MMbYJ9EqhDytt2jTn7ms3v++9S8X+5
YRKDcaxL/0B8wc2qMHDOSuQJt75tFjjDZfWXznfOULzGtJXA2TJg85GGWusHBmCAe2w5yNOSdsrf
P2XsVGsEllqwQufE/XzgoARpgIcopPH86lpzGff50VUiCnRqGJoGQD7R9Bp7i2C+L0gKe6Hrq+CG
RYhAcUasiCkSqYxK5weviqWsf+7jM7RRXyFgZ/jRALe1Uinne7HqP6Cdrb2B6lxvlMmCjoMLvdvt
yIzl+5VPzOCqbrTmCNV6YPbtV6UwHYzPxiXaJvUK7gzXxLo5WaJ8UJeR6zz3q1mfrBPwkaqqBTGu
MY8P3a2mPYH5IPamHo0o60KY+O5CvylhRizQq/Eetcyk8oW158aVpkdR1c9byGWMwD4qRgQNsHKI
7cPK9rcILSitelbAukVi4EhsXp2GeTskQyh5rI5bYNSuZbCPKnDRkl6qGnQkn4OWShzfE4BhF97E
EvlfqEnvmUAEkHe8cb3Vguq32wMP9jy53+9qMFdp6I55C9imeZD4DIGyjEqdGpis+TDUqOrdjK7p
DxsoaHR1zJwBNWESUkl032fOEUwvRg9cczXFlQ1Lg5l0mPVY3qEoxYZFXzUBEUcD/Qq+bEn9x65x
lkf02qRzKrRVXA1lVqEXthW4z2wiLSYkvnrRD+y2pEBg9lEqZUbF8T2gB5wnzWK+lz1WMyGNsq2C
/pmlhhV67pU5jwvAIDqTz+4do2KN/W9/f5muHg6lDvjEOP49iZ5QV6FLIUVe1SaflGbt6tSIesEc
xrQbVzJL6B3jbyoo/hdBRUYuHYqSXQCYsBBjK24pvha9h4M4XqPDpWlIXasDktxBwFlNUvAGlxhV
ECrZ6Sf/JnhgmwgQrCPfwPb63odlQ6lFZea9BY5t/JspNxJB+iy1Nyj3rigqaSfRJ1LtayLeRoNs
HPz2OrrKodBMb2ucbNkUdItlYb7j2RfQNYAVrnwDGWSya5YtNv7iyAKvXfbGnuy4cUpVyBn1sYOU
ZPpT51apzSYKaLwqixM+KbmObjloMYZN/ssQErzP982GXJae1GGHeL3nvhSR5ZHjJjRO+1ueQuRK
GlSgb1SdYOnb8XvOFQI7+YbiiNoG2sJ5Y8Elttb2OTfyvqyf40/PJc6Dqig2i1WcWpIpcJZSATRN
sE6TQRMlr9AYEZxA2Y2pyJLTAKaqUS4zAgIri3cezjuNmx/eL04qH/XIbx5e+XUEM22xkARqbFn7
mxQHx0z1E5FEF+5vMSvMuGe8W2riaQkfFrvC7raVDvSkLJLi2L8hmRlXquSF70OG8RnnqHdOwcjj
24xWuVz4gatd86TMiiJ0BmUjqIZqmo1IRDChL5NZ1rXYeljwXNg2WiZswd8rzWGOSOq1QL/+XLv0
Gpox8JUJCwbh1Zi/ar9GEGANHQ35f4Omtv4qy7VPnEkak6yXXlc5l4ofK3rmzjYVtGbyWqD+vDvj
fNJy7jlcDwdJqDDUKqPlOLoImIXwFUPkszyX3MwWY4l01Wj5+8PIsybreJ2L/+IsfyLOJMNV//Ru
BMhS/JmBzP5bTLZwhyqwM1z8y2EHTVSaRvHPKq/c3by0ai+g5RQeD0or7csUAtkO2DYNK9BcRXWE
9sJp1Rzi9uChzYVZgUSK7gtgvMK8ypBFJslqr2aw9FG3bPDYIEYpd76G/x3x2i8aO2RAhAse3cMi
/DNlqbqkezQdzFDICxTTEx15lxrRiMOZVous2N2WYjfDM+Mz36Nsmif9u6Q2RO22xs5LcXUFQBnV
BfWZsDRvyzbhBw2pav/tcb6uRxEYiRvK6Gmrej95HSRo7zY31zzqkAyqMBf2hgx6NfaGN56RzPGD
CxuD9+2314jGajq4G8OJGRO2hItco8ZpDa6sTSuFnX0ayoNF2HM5+yAVNuJ5GQiRWRR2ltZm0+si
zFruud1m/BXf8Uu2BRcQule3QOhPr21bL3W7tmBJyaclzRdiGYSlqvSM+6H3JPg5JbWPc8h3uQQT
6rD2lYPGm3ndASA5ZZLPsh9h9DozhE6NBaql+HeUTWIeJxXg0/Y6XeCa/dTWi2RBgH/5GDhqSx09
k/LdgYZ00Bg1JpwCwHVhVHVEDW/u02Rh6lwCxSMui4wUzUM2EmUSadMRG2KrXl33c5uOaNT2toqW
RHA4bUjHnhXFB7OGDLqP5k2LYtmkI6K5lzqzxuh5IAMAp7VnlXpcb6Xa43D3R38IH6tL9iPQSMzA
C3yqHYeq/LIlR9abZE4vIG7oUpqPgwNaAb046tF6HR9+26NVpIW5WifePRAskGXLYWRx53OOzI4D
aGwvwvWuv5M5squZa4MBnWNbwfkppf2gW2dTaQpHCiJ3wJw/Uk8qBe8R9q5FqVltqaM3Ty57kNMY
QkcEP3bpWIwCxZo/yk50Pcn4ATrwi0ExkgukzmO4hGqX90S9kWd6oYd31a4WENwqDbB2pbLAIYu4
r0wDgR1kfSSY57eKObiwR5So9d5YTar09RVx2fGC4xEzxo45kAmVsfJb+f2+xEvFfuZ7qtpyNIMx
7wrGM8TlgMAT6rFN7gxVzcJ27czKkOsBbjBUAY1VShlzvUyLqWAkWRc/+MouxxhHxl6guKi9uZW8
mZYMdYHTuclFDgW+q1b52oh2PfXijFpNdcKgpa3QnBt9FGL2p/mzi2pHH4E8NDdVtpa/PJMgPVdT
+XrCQJw1Gj1OGFm6P30m6/WMrCGuR9ChxXuc3QN4xRIYWmsYXitvOClkwIE/sAvuV0E6A099wCRg
PPHfj4i4OHhUdVJi5FywxonART8c/Cy8VOUrLFIvvt6v0KoL+7c8JwFdrIjrETgU4jWEdmXvggzX
AR9p/oEeA0q+ceBfoZ+5BWMuogBVHO4CatIPIJdN6sFcDG7FmaAuaWqB3jRuEwe3AaNyriDFSIyW
j570pUFAFLuvnNBB1vzU5xJMj6lClgzZMTMLofFm6sshqVgp1ouZsyANfcUzLsS6G5FlDrVjq+db
T4ZgNTmprygreOI88QXQW65buaG//4FY4hk++ObW/RFD/ZrvQbVm/6qfLwVjb9KudnUV5RiX1d7U
f+UktryD2qvqTqZZYguXlTpm40bQX0ZIDIvV1UN3bkG7/6q/wqQ0bqonksljcWzcGfy3dhRYNSLZ
GdLodya58Nhey0L8AM2+AW4f12NFBla0N4/Squ0jCbXOZt8JYHCoWY3YXw62JnpLYTkmaL4yuU9v
9kNVN9mV0tpUihZ6HLubAmhL6hnuoAfApXtbxc1V9ygN3iXdYTJ+vrEBkgnBcQXfFNHOcorwnGzt
fC2C0KTR/lYMeWU0iMQ0PiharlQy4gOI9ChUnGJQBB++n8L+RzalI3+qdMtqIHNRamnqSj2V77xJ
z8aI4AMhoyC33Exijiq4nnrnSRfP56rwJndkHt8AAw3nS2YvcD61dzwEie/hvZ5w2z/cg+NteaDr
H+inlqajvQpQXLVikqjvpX4pJdKXHoBVIwGlZnM47oHhB7PG3cI+62S+zY7+uMZb8lg2iI90rNrz
hLeVyMeyOLoQ7JvsuO6A1aS1hjXnyq+7QVugafveuhw9Itk0wKmKLMyIZoEarUawYTwhTyPICW5Y
xUlz0ESlxnstbQdtGCM0e8P/OgPEHzFA8bLq6u0VhH2i/0WBTXheIqkzTNrYkEo534kRdI4jK+4o
69UyhWa01IFuitYmxejcyaALdwTj1WdQhOddJP9fNl/83awW34Cep15LhU1KUoiCF0VVamHQl+Cq
JlY/m0GPB9KWgQ1JGBCZcxO/Z0qfxygcSR0k2VpqkFz+gwVMjjOj6imoios5KAIe0sBarIPzWKjC
0oh7/IlX/vrysFpQfpxkQI8IbaKuZa59Eko7/rf3WeF855UwCx5cwwFK2bFkeV7vY86wGedNxPNy
APwY7a3tECBVvF5c9etZaLG7DMo8NnFZ0GxTuZBqdb8fH8kVtcqKRenhTM1axMSTa2SsnxSMuldD
kO8R/74nwszurFmmZ4vylj0h/fo+UnZ5s55AKHyaW3kWMoiF5I/s0JCNBmmjSI+ZySemc+RL9qLV
HFkFcH06DXnH3OSWJAxlu5qQm1Ftq6tY+mNaFQJZDVPyg2cnZYvFXUUI7oGKZSnEiiUAZLfAJOEk
8scuO5M16h8IFyg2FNQF/5lDlH5sC/RkxJAJoFOZzsGstGGP/9ujsxAd5LrEbpI7NKmEXc1vczSO
Vm5jRqX0Gd+nhuGNUsmNwlwuomLQqkTDOiLzLjIfnGZTI+dVfdDZD6qMZFYT4HyrcNajR3yRgN1j
DAaYvFhplXbxJYFeN5EBv62wUDedlw6AT/k49LTQ6vzBBA1VLpna+0DTkPmB9mMiwzN4bBAuq66h
jFHttoXBhTv3kjbDNEkw/uQ67hjOK33MiOj+ScB7yqPkfH5+I4qhaV5hZAZHx7XmkXW2SmOwlOyh
9PjVtFEMy0R9KxRzPkniMwCbzMGBX4d05zgnbN5EX4g3cXQ6++7gC/eN+iWnLqT7lBkQ6jBIlRSt
WbE8KymsJw+iZId5d+jt4XaK2O2lyhs/54/JUcshUgzCPJEUjTzMPdz7q1aqb0vXPOdMLqiZd0lH
PhDqdX+R0Hp+TagH+4cEoy2tHLrBw/rDytpwiGevlURN+jLvDI2Mp2z34pRDBdzdQIIYdXnu/H0W
y3d9k25tlLWVc7/KQoPIi0J3N4/cSjOx071PXKtxQ47Ks0M4x8/jIJQ/bGcH8resaIt56EZN8zeu
Mh/rukwtnC8eDUjGbQ6begsDTvQJcSBa1dCBGgapctrZaPV8dG44c1zFxzBiL/6D2DYa6q3rPGRu
NBRv7228UXpWGTTqQAjJE0ds3IqsbtPIOIJ+1ANtkjcGhr9/XmQwFrfyqTKGGORtVhZNUU71Iyj2
Xy9M34GR/X9vQe44u2xtBlRLOJekSa404gHsRnclvMuW3ty19luSK3rLMDZuZ7jmgVT+tIwAB2If
D6VTkJ+AidS7VfyQTBfFQrOooKklKIwvJ3sypilZJWmyWNs2M5sCbAA5QuCgVbs1MJsMlGRPv0Dv
v5zFTMhgA2EV78uU1H3QsB+aDBeajBohAo0W60pfmslYCuQUvc/0wKCx+XWpsrktcjBrKhKcmN4p
dUcickZXUe6HDQSU5bTTVeUNuxSd2zt+x5t1gM4IEzGckBSM3WCY/qoa9tt4hJ7udIQJYPLLsis0
RH5PBj0hW73+ewq4zPV3neHJO8k0otrdKX97b3AOlv+a53PYFvleTlb8LM/paEF0v0GArHYZJ5b3
uTYBJOohJVG6bhbrTV42NQJ5yy3vFeoUb8tK40ZiE5fB21RGD3PWkKh8seF0x70lJ+oJQTASHB3S
yQbRNZ8IVm3b27HssXKD58Sdq/yQoGZMZ4Wh3N/lhAdPLf/tBUPnJep4y98eWD5AyzfqA0SIBX/8
LUn4R2Y+pPo8v7Eo95xSE1s/KYpqFXXrex1Svb8xva01jOlydeA4ZrVIQMqn0Dmy3mOxcc/uPrRO
VpUXuoanQLh0Vvbr4SwKhwwBaAs/QHN+jx15DLN5O7uHMWI7C7wvO8SH01jhoQXTrdBMFo3E6Xuy
3/NpD+PArwlKVJpkwt7AXGpNarf4sUNOv5Nyhz8lY1l1b9PwHaxFQxWAIa4GLVqWiVkDI8Cjtzeu
S0x2u5mfzEkkKm33MzU/mfY8+Iwo2jsuIXovFq/ib9NhFyx8cRAnKXLVl/+35b5ZBs6OsqhwhbFp
NGmln8AHoD5hRN5ze2hoGeIpQ7O+NbLjsjlfbivY0GBR3xtgAdfAO5zt8dXmq8rs3AIaIios4H7r
iKw11Cn34DzAnY6Y2qFA4am83skuq1rd7c/Fzgzfq9mo8HiPxUCIcJc99ColNCIpHqeNTHqSDESu
B6s9MJd1FRKP+X0metULEXQKsnSgcLyyk2RfAewiTkMbdoTFPFDod54Ohn22Z0U2ztjcqUYNldcn
aBWymCoJI1LlCrMyhhCf2CCV3gct9j9xMW2mDwerXDvfz9kJSrEU9YYtz30xvtOKsA7qiZthIs/+
YNa+NYjvoWLxHTCUWEniQ/FLNuqKkByN8ROPLKDDV1VP6ejvfqnId9Bw2vQZwU+4DW8mncelHT7N
OtvTFFs+PzcA/h3+rVtpM1m5TAFDvyLZMsAN/XJL8dG40dJTsWZ7P2CRw4CAKsSQh9vFXRKmUA13
iFB4m7WvQPIMTDHMl01HGGHPgDAgBZ5RYFDg/2vCGMl8kJtu+VRHDohReh9TRGY3RXcqIqc+cEjn
qfRUIChS+D8QFmouyWwuEoYsNkiwv3UE8TYu5bpS6+aFqzgg8obaC/OkkjCCVOlzQbeLng4wNnPf
DRlkC6xfWP84eAtZFPUWRHHs4i1iWn/GcEbj+oPCX+aGakA4JrWWx3jH/gXfTMFyTv65ueiSbYVv
5lSVh7Q9HowzEuyiPU28WmtB5PRerTGMB87XKd9nHP+DM6AovFDS31DjYUDqSDyziaENGTqMSRRV
czi9HuTmAJPKLuO3KSBWPW47e5x9aS6LKTAXTKtKZG3eNjEL2PkWFkMLOSJHRAAb7yOpcksrXbVt
X+YNfL4zbOer0O8aIyXFlNInYBxogLbiLDlwBAdcMV7lSbjb7v+M+OFf6B+tM7s4ahLnqhGcGJxr
KitlOomr5nO2ARUg2aGuxy+f6cUiVAHCnoRBdBx8ZdTxzSwXkvQjNtimO1nP7RfhWqWZoqepHjX4
X9BgUwkxhhyq+TB7looW8gjookxVrK0FT0B+WKS/3UIG/0EQ6AAh71XkSfcsd1FEaUFrsAXy9WSk
JBBypUAtSGEwsNblMmSFaDHlV7S9MEQqyioQk41e2JP1HE2KGPPYkiTJrYs+v/3IruD7cV+zoHmu
c0nzO8exq1ClVCQqtyhT7ctr2remLmLPbSLAVHVH9yUJaIOrOnlLi/in5U4HjW00TqJV192X6dgv
cvU28wMM7uDAszLMMAA0KQ6/I7PQFT4Dp7rnIJr+WZaP2tuKk4t2Fyda5pddFVbqvbwct1WaBsDf
o/K6ta02+aGIOO+yX/iA7ua15DupTr9Iodasjz9UGvNaS6jLNMFLrv844LKvE0IFuzG88cjy5YIh
pHqX0FipW6hyFtidLBFcauZV9doyRfUEoPCZ1ioh4sNYxfheY/FhIr5YtBWPyGT2DU3S6Ux9CX7P
PiOJeI/PyKPkmR6xwIIGHQuqwIN8YKsgt/ZgIzKvJR9SFxqFI9gMLqqzly+5PhGfKUKoRq2ddPQr
nvTnpPerSCA9ksD6EgCzrnOj2RrMG0Jsk6ZB0B6w/pMHJQTwO37DEaMQkgjvV0MnSXOH9OArnIoc
/Z0JaDhrTKcBX1S3GIHwqxC2xxi8CBxdXFC+7VUGFK/fo+B1lq7s0oXIGbxV088dE6oZXeu+drvE
C/OpV6fpz+dxcRv/EY9DXHb6Ttw3j7diJx3/KuoEPjzz35+8FvloLMXca95pdNNtxBuLZO8AkPzc
RGNvmywMQZ0vFC0U7wYyQycIxpneeFtXhVBxYAzXojnnyLIn8dQZ4yqjeJp007dmSq3q9GBLLM4I
79YBCmhO16rUBj0XhbOifoc31Vms7kKT+Jd6fyWn58O+NK7k/O/3N9q5f+KDXOFJcp9Sw/WYG2nM
mcklZiAy1WxafPR5jsyp8lc6XDb3P12mV37f+4Wij38hN2KQ5ykIk4wV8dkJr8Ki62kTIQf0/2FU
KCGtgGDrn1asaiy7U+WG6I0wvgYftMxELBiDph7FlwuI35Z+3DBm5IPoWG/WVKSPbuXuL3Gxy9Dr
4AQVrdF8DBNp1v5269/hbi5Wfq275dCVrih8GH20eHuTnfxwg1dVzWiL2H0TQEM5f9DtcHnXNw4A
2RIq8l36YoLwrXC+BJMM0eCkkuSIbmjdru26JCRVieCaNv6Q/b6G2nBWcVnerbF7g/VkH1hgu+YQ
zUBSmcxTrV/ckqVcNYEmJydTFioJepe+azim3IAMC23DJapxZBw8Qq9IQPoNYSLT6ZT7qbye2pct
yYlCuW46ICAFsbu/lNeHpLT25EZrVNUGTNi2EXG8vDB+rjvBJLTjWQd8IonK/SvCVKhRLTsyC2HO
9Xn2286Q1EDR2KRSBlX9pzz7BsxUFsLg0EB/qWK4htyV8HTe+AImU/rHBX9Ku3rfvHYlvVx4lkSw
5AHsOQ3zOIeIPxk3YdR3Pkmt49es7cBt4OCcJWX1t3GfHCzoFRMNfDttdIPXe172XTyucvRHlWq9
DFxagdk0sh/+rL1o8tzYtbNh8Qni0dnLRa8PFQr+g+K8EvVJg8+t/oKX96hW8Bh8TdHaQRoVi4+S
/QofhTo4hDOADBhDF7a1ek+DwlrxPLfAz0V9ZcVNm5Dz5DI07WCbrlXjN7Tuxzwsaw1HBkLJ69dZ
gOn1WIqTWit5ueojDhJ4IQejJrXP47ODOxgkGPshD9wsXR5X6n/vN6ygENZjvTrAOL9nzhs+qYKs
BW7sDxJwbACfY/isVSu3XebDRHrt7w+yGwg2omk3IDuk9nHfk6moY7JlieU4H9iHzu4L+v8t5QdW
DzCedyZCfY3DujEPV+m4FQkZjB9myJrZz8p0mj/uV1w1Sid7KIkad90GEnldHS5DqAK5UT41sYwb
Srw8S1wfpFLn5+87zaayrYgUQlzll3uStk6twT5cKifdFxR7wLpXaFhb0hXsTSQJD2bBwbXjJhz7
BZslgSPX1Jfv0ZTpY30EXgZkQKCWaD7cf9k+XKXeegudo5GK98JiCO/+LKEIaicXmh1SpndMsiUP
reYlNL0cvC6riQOM+UEKZnxyVK2CqbddghsXAbCN/zaiHkdSWNbguM4ajimPHNeWztXCYcJnJDcU
waSYgOdOJDiMzyZ1yaNjKEi7SiNSNhaTzfiCC800V6L6GFWnQ+8iNFFdEuHdxMAFFQ+jmjU7Udu9
e4GsHY8hkP8Lhtyi+/3PjpqGLzp1yLE0AR8r7aQ/wE7ZJ9cHpcAnWn8XNbP61Yxhka9fDiF465JM
wWQsmx2AnaWOJNjpSI3rmJO6pPP9Bnwo1czvzaKOkBKwcDPhqZuXE3ZXWH4/BDF/he/Ow1eM+Akp
k8KHHxO0NWNC7LueY2y3sHyULfyPrN3THSlanC4kGgtZeY/CoP0UbWOcjGDeqNRmlKLGxsSd96QF
u5LYy27RmMOewP0q0a4klbVYXCDe83npnW4xv3t7p93FyGJ6/JFwj4OGaHyeGaIkUEhs9KWcviA6
BSB4RYC9GA6rq721JTRAq0BTMQB0FdBgTZvA4Co+S5+71eyL8/GhY2ch4lQq2O3wRcg3MMgfS122
vfczo3ejNvVPCuJ0uPTJoBl/AUTCx73dBGcqaVM9nBWbmuWWTOWr3b/47znRm+svSiXb35M7Ipfq
6u5NoxYvQf9k3zi6QKI4QXYLV/PcSLEo+EXqLbuIajiINBv2r5vY9/MCmJ5DbnNMkegj4C+i+iWw
bkuCJfKILK8x5oBdI1B00Jvlp4HGC15pCMD/YTkM4l5eaS3DO4CgYVQyZiu2Cv9qHPj/kG3b9g9/
rbhLvDM+mppSA/Od12a2/TUCq6JZCwc7Q/y5Qm3xHhNk339pU/HianY1NfanJgeW1ZrgPUSw9aql
c4AvJiQiOxYds4HdnOY97wR3jyWICG0A2QsseHddRruQUlLzzovuEaNADZceu9n6RUObqSQslzKx
cPUOTulmwADcEMvGrSCGKxRTPgRpkKFgftrjtLY9WX+JQTEF/STuAJe0atyFf+7Czta9PSxKMWKm
mjdr50Oq4hIDsjKuAvAwQr7NXV2EfdBDc+exZW1JknG+HDkaNECwwatRwpZdQ9MCFEtvipzJZUS3
y3H2954EBtHoSbgt0SzV2hm75Tx+lSKI0zYeS7s3jHsAUOIlCuDuLS1McQQSFJvsoj4oX1pnJwaW
JWETyT0V8FoXfahPE0feCu18HMYQuOxZLcl3LpKW2MDIqvxzsWeHfV8izyF3YxIURP2IKqGnDuIZ
9fAv0p97OLHOz3KENvrjumn3ndVMFmC6+fzgAlpm23lg6ettmkG2cqLJEYvo79D2wVr1TdNQVJJJ
zswt5BAOwg/Bmxwp2rcW9/PzFevSjRrdlactCvqW/GG6JCsp+7VWKhJkrFTZ/7sWWO2dtSjXZiZG
nC3AB8E7InyZNzoB6Z6Nn/KXyoEa+M0pwHbDE2hQgek/GAwFi7J/FN6X8foJGctLR2jutBIwykps
o7E3DQ3j1jJCEzlKPmtQXDMfVVVUx8RO59gJsrr6RJgb23Oob0AUXIFhz/UlMoHMRG98mE4uG3ll
7qE1Trlxs9CcX8TCQb19iOrGTPyfCH5JFJ8RKojYoe77mzkG/3OQoM9kcUJ6cRdpgdb3Y2qHYMEs
CZ0uAS3uiNpiQ0IO5oh+ADuJuiDJLoXFCxZweB+AqMV9nTCzdDCsuJ4hJN1uJ7RYR5mEBAL2Nc8r
UyW8LpxZ4Rl4bLoXcKwTqu4OkY0Qbig7UqidDXQAwI243aHn2IrK+JzSS3C6Gyj7xk0qZuFx/hVR
50AY7QnGnYwXYLXBApxtbakyfYkFTPvStrYUyg36wW3d5rPF2YjkDb7fnQnKMqqTGmyktyhEolJh
APs5czRfaI5jIgjZHYuMdaWr4JHLfl21Bmd3a70ThYzogrKb/MEYy21elyrQ274jl5yzPO+Uz2w4
VJ0pMTTMCu7NJKCi+kLV/IS4LEuArUQ5nuQbpK++JMvvWn+3hk9ginCwfBR2ggJYlryOuRyXpwdn
aoAEl57NKeDA02sQZ4EMRKZ9Yp/NrtViWNHJ6CgCJpvNllRYuh7Yp1M1a5Jr9yKYEjC7i3z+E7ym
Z87kS4FXFNTMjYbVoAKMHh2WS3vOBbDzuzydIrMAmVOQRakXu1ur9lMngUQMvskneadjMu5IcWmV
uZ0GdUy7VWxJy4/Of/Gu8uCot2Cv5YO73sUl4gz2HQ8SUAzpc8xHNQfXLBuXyCTGHAb2Apo5SSoh
x7fsEXM2+ssEa97Lx2lHS7eX1mAt3PTaAQuFRYSYBXW4aS77jiz53OtvXjjhf/fRO5JQfiYsnvv2
U4q6YZGRF0RfVrUZ0P0Fhcx238CUd+5lX1Ob5aXbC7pXga7PsI21pzxYv5FBm92jTxKulW8IPPXx
2Mr1Nqdq4LrzksqOKliI7OiFnytuorZd43XY8Mz6X2hFca1dA4OL0d2z3De7WpyRLt8ADhznx472
U3PMDqHTUvDFuF3gmmrrCIOkAo7N6WgjSgoWobD7G1hrzscxlR6E0u2qiNqt98V4VBNDlAu2YtfF
mPKKEUoOIRjw/6D1+ERprmfqgQPxKa2oK2SAKqrqinkDXCpf7tslSHcaNmNNaC6L9WcmKyG56FXX
vxT7sdnmex4beUzIGlsrKvy2A4YX+RlVvH4fvwEQpI5GuDP/ZRKbD1s6DXI6HDSy7XgpWkLddFpq
BIveL1GVj3ttXHALgZ/TXBBZ8JZmiCuc8UMXzwcfzbChqSzyuuuJ9jj8KyeOFS3ye/5ndMZLbfb8
nqeFovShx1Dot9tTa5b/or1eLpx7Lwmuf3/QMS94TGDb7tGPnX4lpHOkTXZ/+FceU0r3uu++1Cp3
Y3YfQaiSjTHL6iKd0ISDVOhf8ZeU+KuRYz1IPV9S2gvky1ZcCqyFHqqYEo1W6esfCozd1CqExHC/
rTi4hlGL9cia+sVDsLbs+ebUIWplCrd3GOSGqBNuwa+nhKLziK0Nh6qFpPkch6E00Z4B5lyhjJx+
l/iK5VzxrxozVI6UKt4O8mwuhzvhBf9aei1TVLGZvOYIdwwJS5zxmy1IvKF0HUPv+Lfc1KIY0dMw
17KuCvbJg/ViqkDPJiYU5Okqf2cE7r8UVrYsdSPVbbiroUAR5p08Q3t0mma2oVCIQelQMPuVOUpi
4kCbJvMDyAZo4hYbHzZ/KC7uEyiSIjpvL4pMLN3JU5QaejrrmM/bqhg36t/ioNLdXlt15X5lmRbw
59ORd0pEXmn2j5WvFCffVwRGnfNM1le9LtNjBEFLBJ5iznSz7+J7wHc5PGWQdi0hBra8AxXKXvjx
evZFE3LMzMCoiL25AglC50VjHn7JGh/Ncd7khfanvYPO7yjPUnrLSMT8hO4m/mFM2Tuj6iKNlnXh
ZpHh17pemxwMj2djYYhXJQ9T+47hcZ9f1xt5xVc6T7wdF08ghVrO3QFwMXRFICDIPo8EgsoreMp0
UbltrL7xaj0PfexGvRzxQz8z5Lq7RLxJOGXSp8tHa/7Bh+FhKa/DXhrU1zPhwGlYQpMKfi9849Nn
0bWLCPlY1WoFCfvNF2KPkhcCsgS+J4pw77Y3F1fkT6+VpIu6xg97o2JwySgZSne5rX82+wMcAEBq
C1miIpieQhyOgAQ+Gv9mpLG1CKTqoAYw0sgW6HqE9UfkOtqcGYwZ5GJR3/hKrMo3iz1UAA3jRwQr
kxlj3Aq75W1PWqg1rA46wsP/zQJmMODcygtl+gapeofYw4lvL3lyrC8Z8HDUcjxGKCZpMTOBc/D9
W4pBlPeH6f2B2mudMWVwFCw9PPC59t6KR5LY9tOJoQYnKUf3n1U575S7U6uYPR7j1tlxvDbLzfCT
rkCt48grEjQg0iCUQge/i3kNGexpElZSgJThj1A3aAvqf2WC8d71wEHdtXwmAyyeRmTMGmO3Es8t
JK9a4HrBORGgqL8nCCVdvZ+5jG6Sb0feJHNlGt7UqTI1pyGeKftgF/OiePXtdESeRxyvS/7YJmjp
KUCBb8nwIkMxeJGlPEOfvrITQX6qL4xt8P7ah87M8P7WthyCuOBAGoLb8rAGBXjC8jCnSs+E6nOe
l6ewMohDnnwUFPQmdUQKUxcx/wGjMkgtD7HeoKSBebATr6CXTNjhD6Q705IiBLlc2h4bWhMvjVrU
qEEv9pjnUp6g62j5pHEaj9N/Hx+h6E4nx0upTjDARHrqRevn7nmOISWvfdKLEYEHAJ+AEvy/fxZd
4G0PIrWuOHVUi9U12xssEIhFXUPkaxy3yq0VZ5hyw9zcut4jLDTq4PGIoNlcdc7mfw0niXfN2eYu
84Tr56rJfS6Ef/n/dRf82A/3APEyAxCapicu9bnc8yzfHKW7Z7zzOIFL78G0UNhr2sHOqBdWrYwv
KHh6Xe1VVCIgX8rsbABHg14j4Zh8hCydzz/5Y6Q3mn6OLwSEXQ2EYclPZKEzTQkr947HXyYdrSrx
cJG/bVsJExW8VnlCC48RXCRANO+HNFDSXaB5Kz5cogV83NV2IRZdaGOi98wmqoQDU4B2h3vWr96/
g56Td+VU6mCj43DhCW72K0u0XyJG5q0LJ7SdPKOum/D54LluPdpFkTTP9v1q4p1rEgJ6oImyvvB2
iIg9oHe68+7y6impe+0yKfMclPESGGDHUsJ8hWdzSxpheDQibfch5IPviowrJ78QeEgQ8UoW5XnU
0yOlxdrbbokrrTSfDScVvMjIJ5l0YeKKgHOwbrnmZcvwd1PJ48ZImXfYcA2Y3VGku1kidqb9tox9
y3Doje5s2wv+nmI/Yla4NS1eH+nMCNiVFfWkEU8JEt4qSMX03fEpzP6Z5y00FmUIuvy8/ynN/8ul
wK/QzgwEJb6A3Bx8GNmn7F9obEvXPFw1G74F3HixoL9qT+1MqYt0QawHA4d3VdO705YnqqTTMA4Z
DUGwj8uw3SKgAeiQetpZYWfkiZZ8L3vM6QHuFagQRgzoGbZSbdqOEJiR9b/WmpuVaZy9F/v89rmd
5eCx+5QOUvye4oP3CmbLgzqlKF0X/G504ahEaAGAQzBp+1INtYzqooqyZbl6pYqrVhmPZQX6tRxL
XUV5Mx6MiyIwGEhwq7paqgyayPixyTvOYReWAQzITVFO4+apdQg1YDHrvojT7Mv3d1WvF4YN7JnS
Vmv8cdmMeoH79UrH7OYLW67ag13C9A/3WW/mMU4sQ/tdnR9niW37HQXJETFF6CiPGU5OF5BWMTKb
1RG6bl2kIO4Mwb8pIQOYYJ0oYmTVCf931bCvweWfcJYaanV7WYcFLB6jJMvg5qjS+4FiRD1gu4Cu
3tqmexP4hKjgBBbMnmc53kNckNflYqVVM+pY8GKMfzDOfLYr5KwuQ0KD4GIVSP4/9kkVhWcVgmfg
REVOXPOKCHCsIOH8MVIwkKbLNryNnHot1D/spPRQXIUtXDXwIn561SqdHFgaS6sYtS4qHBJ2j5lV
jBs7BzX9+FB4LwmB0+t/3/y7sTGpIkzsjZEJleDDYinsMkS5n6/FVVpTxD3Ad6YX2nzOubZhMGwq
06ydZEkt8r9gRvyTrJV1qFev3Z8Gk6bjKLflxZk31MFNUj4HWkMk+LcNsk7eqzWox7dPMfkCaviN
vCB8aWvr3vNNsFGf97oVJWA/86L8alFde0syUdeOm0CVHpOBvXtlM8L0N5w8WoJrnNTmjWxtq/GK
nN61HW3kcunjecFulT3hJONvyE04OKPXUWfttSU9uhVibHJIGAu3Qb2a2Qj/bOBLFqo4H/EjHqyB
A8fvEgGOTG0pfDZ4uHWcNJLOwBLv0KLS3NL1ZyLhpY6Ec/4rVdlgCDdj7VYDlWcv0iTK4rC4gJr9
crEmF/Erp5ZY+Xgf9tWVPWGFpZEO4MgAMwkrqgbMzZWmGgyTE0W/ESYrYMuQLVUaYkoO7nnVA8S0
TL+ItJ69tZPdGAmeyu84iq+lioOTbJZMx1q40n/tZ9Tj6LZ3vfh7mod3N/C2mLHOetAgHtF/7fHR
VU5FA61lsWXCvYzCSx5LlZRSbQ89VxptJP2eOnNNajoswDWSoygzmJ1VZRdQj6my2nLFOHA+p5cj
2uq/A7baUqpDwhMSxbnB3QY9W8x1MNgpeSKV6V0NxVAadUcCpe4v1fd8XYuThHnBdormqF1PTXfx
JL3eSlsU3ZLCtMgqPlY/C6DnDjlKww6gWy7O18GedQ7mhBqlPcdvMutGKS/qoiggfVfDCl1PYuMY
ejBhj8102qmGBOLln9zfESufllfV7V4rSbvEL0Y4amZR1++mrJaou8OqmuYnQjgHUoExzhSbiJJf
nGqpngNTKK51em36Ixi/7ABiiyFpVfUaWEQHfT5UBdiLMxp+9GDNuqmwm3Q1STBndOqDJV1VkGo3
i0kcCIxk50hn5slOTooUtvIL49A3lkxHIZpWg5c9Me1MZXSZmqGM9to8cSAuy9efP17fQLCVO8xN
ei68LkrcZMSP8ziR0JoYGWuUUhGcxM3ccKSRt53CY8W3YhINP4QB1kqs1jeGS2jmqDFpW87CWVnf
lvomclkcGwQf0bfabXYYjlAxuLkwTqVcHeklGxN7xdsCbdOL7O5lUPtVjNuQTv56O3r1i/28+ffB
r1cO+0ekyv06/N8bNOyWxSg6iQfpwkv6sgQ/X9JFrHYsacJt07KYNlFueK32YKSuQXAuOXBFt79n
jKRt5Jf9hurtLj0t8i/xgoisVk/UMJ2kXQe+3FsfNGMxyoOc44j4MEDd7pSVxyGfXmmRpF1k91OX
nbGREwQI6adlLVu2T0qhXLsDQiF5m/ugOMSlFfAe5oiHAOJ7OZgDz9FQR4/B5HGSwzRBe1g+0yWj
kWkuB3XGPRAcuGXE0EWgBjMREVMGR/RDAg7B7YYD+FX4cI/TJHp7Y824OWcAm7zFTf/b3WyccfNI
/4Y97zcwsAo6UeP9VRFU+aY5bO/u7Rri8iQ3FAZwQB9IIjrDS6U0D4CErFcyIV5AFdhSHrYrwp8t
22kCBrtReSbmBfvILy5uoWqjpAyVc4ehi8A3qodrgow3QXSTR3aumAM41Dcd63YW+WcqqSTvFvQf
1yEe/+cGZiWjjz0Qy4mCuKIjvuy0GCcyqplWCPgSeFYOvAHkT2+cyFY6hewlyG6pMdtcInSepc1h
N2PYDSdHwkoQQ/vfRzv2fi/+qgIj+kY7l4Cxa4iR0vXbCpBI7K7mXyoozZ/BBzKK+5qnpjXePRu5
ekPmtsxyArFgo4arzZOqr0kOx4PVrcAM68uHSFcUlDexwan7OGUU+52GcWuXwlE8BZmOTTpQS4fa
sAhpV61nvVqkIX+tIJ+VVC+wV/jtSWUgk9MxcCYiiQys3S3H2h0XyO8MoOSwINLn/khylHiF4uix
b8OWpqcWzNHvBjTTAK0p7/YAE8Qdnn1Oe+e3QKfX1FtfGef9tU70/9Q55TlZFMggo9IGp4iZ/NLs
MZ2M8H46QextWmNTR8qiSLLGpRjS03dAdrV/1y67pGoZH4ouzrGY09ZXlCKSQhglgzAFDUUzF9S6
EywMw6DR65KzSdrE/WMKziOrB2VPeWo0cbMNXToLbVZN/UEnznM4DON4FBmvd8v26c9CjIZGxphY
8wXA7mEVRPHJU9U035lBx470lpfsXKIW5pE5Nlm8LvUBWdhbbFwv7MSqx6VbTZG9JWUguFJ+gnza
OgkXdEN61z7U5comEVAW3GXGwD/8ePMIwr1soNKDPRQlkMx7HA/TP0JVwEDTI229z6u8kYnT+92U
N8a/LE0iHVAR0F7LmIxZyFuDjHTRJ+eR1J9TaHTPSF67xNoNybDM3lrqXlCyAeSuerHM+CGdOJAX
6wox08AnkmQq/ST2g8SrH5Vjo/eP4AJnDE01gCW0djG2FeBzjr1KRtJjt4kFhT25R9PKAQ7uROQB
mnSKbYbs0vtjGxFF9LIcntrDFROvpwwNB+5AOnClujn0LMEfsjWCBnkVoPhwcOQQJHRT2RtnIdYW
HcC45+79ohkLYF4kFZrOhycsXpAZwFBA1OvHzpMs9ef1PIFIF0JlC+NJtNpZZ+UTPMwSry0WbWhn
oFW1fRukb82wLH6dy5SFGsfTA8GOAGgui/SWDYd+fUNNuxP2y7iFhJ+3A/9Aw7QVB2XeyRSEMFGa
9V3Gyw0toEXZIb3+ESIKGQmJM5jmZRW0GoFCxrdXV6iEDnwtaIZdQGeCAP2L4ew40X3YkALAz4We
OPZTv25G8sNPz4sugmzXQ7KRqbtlrEhIEKQBgFiwGhaQn5T2u9Q11s9k4vWIE8lmNFmDLNAVYEXl
OdHLwofG2KNrLkKBdJT37Ai9H0pFsLXP3IOhbYhHJ8aZy9PGDg8zbZgFfTPg64aGU/HYmvsQtJKP
z0O+AZRlMSpnBdqJ+SgRiUpz07pEef4pL1OmxBF9Vqx2IGqKWu2yUQPAEMT47FGf5oaoRMYZ2koK
t9bZk/nbFkuSqwG4xz51Pvs4IMP2taHigyHFrIJN99TfUvuA7nLYmGm7wzFhCtvIfhzQ4VhgnTRH
zvD4FecTAzCxvGMCYbmM6YTLEAQ6xA+Um6XXzOIZhhLm00Ga1opTj7L6mmjo4PhcRxsp5kLe2aI9
lB0YpkgWm4IDlmTBMIUW6Cq3tF023Pe0g1k1xcFdUTVFmo8kacT6vNSjfZmY+cIyCKV+1PS3Vs+7
W0CpQVa52czCs3SD0j+Rb8F9ZpticJaCo23Hmg6A6Z4xoaL90F//x5ljGPueEqlMChBhWJBbXyKS
M9P5nrSF5IFnS7+SNfu5UPyZU8FbmHbRKE1CXUglUepvk3IPIYu7yG+4dusqAvm96AsjXE/CkthP
km6L/7orUf1L9gJw9tb4ITVd5gMBDF/NS+M2TSHqjMQ9HJTZWDOqlBtSTOjRSKvATpOzv4yYPvyc
5DyqeF8k+uhys5Ilab9YPCaB2V3LI9qkujIH5DscEoupTLqaAJrUCsbfOS6kfbRyMjhevzsYaR2D
RNuk4E3ZQLxluhJOISvA+2XFhgGxA5hkmdmNExxEjrPzoWRwWB07bvW2cVIpr5cL74JR2QbG3Pfl
yub9m3cELLZVHBr/6Gr2+8Di7cFsEXcdRqBE+Yb7W0HEEtqF1wZsJCSGLj+c1GGQSX/M8Hvd2ms0
aXj1SGoSGKgthQHTeS9Iba6EFNkSTpL7yPWBTAADu/J+aVf5Z4Tq3Ry60sI2owAIdwr04T0C4hm+
q9okqp3LpgYLq5a1C6ZJu+BmvhbPCW7D9OnMsxuC4/OSvLfaS9SRD8K4KLSu8FeXM/Z18TJkMfyp
1toTYka1Bp3LZ2MVKEMwHF1LPUMGFRKzdQAdCT11AoshxsCJSf0ZZ08Had2+r0sWDXYZP5Br9+PW
a48NTZw3HizZ8hjG9VIgtH9Eda43L7MjIVTGSOvEllbS2/02s4wd2zMLv+sSdKq0NknhZDXQ7xt8
SkDjsel4wnpkoaS40yNODK2y/SK8n04c0g5zvxsVfh6e+zPVuE1KaY517lS9n8oeshv6QDSiLpfd
/EZFsPuDLFE++ZD3E8vIPK0V9JHqdP14zU2Mso+w2F7AU0Ob4ialKJsz/K1Ybrs55G3Fxdt0dvB4
FP4kpyVS6Gp4JNEi+3n56YOa72x0aYUtq0LEcS2zpfna5h6c7hlNBgsqeDdX9H67Ji5WkdboP/lE
6DQlrumktppy3kyzuHsg0D3tNdY/hVDWU/QhfgC1vylmvKy88S7MypsZD4BC82cZIz8IZhBKR8zW
ljx53z06bj2eWDCHgQpnjwkVVKVbSiUhthsUHbHsz/avX4U7tsmpioNQlsRWQ+Sgawh72fklVh2Q
O6YcdG4xlyRABqD9M8X2jQEN2hjiyh/USeUuea5WmdXIXjDoT+ysqq5rMnbIeEhphI81SDEQMtgL
DJwMmMdBQw+roPkNy8DVvMD7T2MWLTNYo73ubhS+m7P4suMShfhJa0KYl2Gt+c8tX2C/Nm5sEl8X
3YRJUER//OT+1N3+KjzQGowB5YhSp1wbgmtSpWobPjRGSQ+ChU4Wulv9zaIq4cyR0pl9cn/t9fU/
umdElDEMjokfA1N73CH/0IOL4yGOqBr94PlaCeNIP206xAF3vzu3MnQw7pJmSKCSMlzrFPKXzBP1
uqQ7PDz+1lX/tFRsE686AoOQN3v9opnObkoEKckwg8j8E+2dkLDwofbW7zeLjKnn2vH7BrBnx0yi
RgvwCp2BGRgC9z1czO+TkvzYSDrkM2CturMonI3iOjr5QMYQye2hb2VzdjtnOiVRyfKDCY7dLyw8
gQkwgNCRct9qp4uFeJUxXgc/bdxiYZiWxbxipNeJVTS1p1HXGd90LVCDqmKINPeKvpZc6mBpHdKx
pLwEdkaBRlv7d+Biu8KGuuI+4zWbzXiIeEYbr5oihH7ngnIyety42gAcTr67aA2dpmiDp6vIj2sC
PTHlyz20aTAUb6SgttghZ5bFBCeuLkNgiitlrctMv+cZg9prDgTIIyBR3NaPHX+C32BZPid53aci
1KyMpPXphuR2jmOGS/49nyWs6bZ2qlKc3wuLiPKgXnrczsNAtPwbSYGeBv3tUwEwIXMBF+FmL1iJ
U/ryq9lJ3MDyzzpNUyR2cosWzmgY2g4zFHH32k4oqhWNRGcnluRZ7hEDqE6I0dUK387BXb1TCuR1
XURfKxLJJbp1kAR2emV9TqlXIoguelzehsp+ZpmLOADlXj17FvVwhAmI4Di5QiM0c4jEZO+wpmL8
jr3eqh3sZvcAIiTb2kOMQybqFJsat9QS7JQ6vo0vj+AooujpdJi/3koGNUGWoK5sS+55VrFH18Tr
tXXM7VtZXnd3M1LTV1+QWu0Dyf7joYo2L3pIUGVWf0dpIdIlY3go+np0DOkFptSKSDEQlpIYRDUc
tJHllZSkeHHDDqp9xhkHthvCWcufsxO6Nftc8RXS7z2tFt2d8n8NZithMmQj84/RDK3D8Oi6bP56
mm4fN5CuZHKXEnMAMBvRdssGYPGgd1KeNj4VyrRmj3Xe/GI28T68WaLlLWWdGrl2P9yqhbeL+svu
9hl0fDasfwSq14UIPyaOGnKWLC6kbnPAmNV4C8+oqZvARIt9bNJue4nHgIu3LF2HAJOI5PQxJ4wM
fm/uDL5EfJ+li7X/nfuz1CkUvOCTK3QOZkkXfoQfSPBbsRC0mLoQwQtfkLtkcLc2m0jrUBbptTsJ
xPXE/qG9twGlGVCBwXoraF32qKDQqkRgCwxxePpX/Gh8WghVmVWOagljZQVYlmXWPWpbmLr3qsh5
D7YQa01e8M3TFOHVDCVMMbKsRfZHpoLGDV8eQ9isqg6NL2DtksYtBblVGr+C17LjClIiPYO5mi/P
cqFpTLy3KPxS5zMFLNcATK3RD5/k4RqkHsqc9t+0j0/5R7BYh5i9NwYUA9QBzmEtFXK71sJVcSOr
2tghkV78zjtB7KN3PZ1NL5rxOOmi4HUPro0bJtS1CsWIXsetG/tDxD0fqCWeNkwfvXVobPR8MvjN
BF/Iznn3gUGvTgJ9/1sG38oGUd/n6AefRekx2LLFeo0ibs1BGIGDR+Vc3Dv6T8tqREXxp2aF76kQ
lDM8APc1K/cDy0ZZhR9/+jmibaGN6bqVlCmTIViBeLDDnqiSkbX6k7TOJ8c1Ix0fpFPEW21ZCk3x
hFjIMHFx4zNDtE2veUUrMjyAPNFR1P9QDAep/oY0obCHeTHxdGi5OSpP6J/8fCumw4+KSubK0uth
y3JwANGgZBJm33qbbDWuHQHZs4gjvhEFPCsDgJ1XjR0P+f9cRTX8zyw1Oic06K+xebnXhX4dfBCn
svoICcsAay2ctZDOX3r/kvC8vLID2g2z6965LjYE/E9q3STjsGDjEPFId/XJ7SKO/tp4+Aigd6jD
onQv6wwMQx8JPEBBgZ0aoj0pEs0DtcHR9EVOM31VOhR1qCky8I3+4JtzPzR4L9JGnV3H/aYXT9xz
eeu2OkkHhTxqtnpY7l4JPpKaEhP4/yO4IS1alRz4l8PE+RGId7WSx9ASgtTpp9ocwxxAXOGDxljF
bBiiD/4XTnTbIzL2oN1AhdeDAjLCYIZJi0L1sVsFWI5DrYBZAw7XrtpxUhXPuprMe9/CW9JwA0No
a5swJ6reObb1DFWWkDkz708+eggbS6cf+8uL7R0jTbdPwd0jgdqG23O7nUkz2hN4gE2xAsMFuDOQ
+xWWzc8rptsjYg+BKW25n74qICwevv/65uYLH8Sd8K5dEEAtzqLPVBhf+Itml5Q3fGA0tUMsQ1br
Q10j7mQzb1W2/safJDaq1EIaTv/vdTO7bGB9stl/burJ1uwYLih8c42NW1oZAtoCVLpc7zHzqtGw
FU4NorYpNMhyFga7clIoL9oH8TjJqMT2xSah8RePElbdwnl5NyKQ7N4vxNU1K2nyzf3IKxvuQLRy
aTzGMdSv2saV59QWC9RBUWjxl8qj0V7ENDZW90cRzvfk5th0P5BaCmWJY6Kw5zQkxBMPiE9gJMmz
k51TsQGhUWgRNTC1QFYCrDZ3cyXgR+Wse68OT++US1NgoyFGnK7vFPx3vl1DcU0BC82v/Sp4LqrG
toTrTAR/NMJ/Flzy8959+4XgiYEKFNvXzZn//vl80SZ9Dhw8FD4c96R0VyRxjpWZrl6AQKMvnciP
moTSHK84U/lf7kMY7cW2V3Y0Ubi3nyAnH21LLd6XVZTVh/rgQy02NO1JAwSkyzAkVRk097ubfrOI
pekKJcOcuFSj3DSQsmSGvWesjok2Ggzxqa58xm2i1J9Pqg9+5M0tXeHEhPycImBp4SV95im5Br4u
0UpL+wZTbAYWqXonWb9ZZ3VF7sEgBjLnt3SmFRI5Q/6c5Ogs5zzydHiwxHYVKjBJFo7B/iix145k
cjJcTwlPs5WcPUxga5T3El1PhpE4H5zTlehOJVHFNzDlUbQUw3yA2aOs4AaykBn5ep361Po8cdK+
9DsgyzWPNqRzcShcl+UkxI4XXqSR0qLYH1W23Xf6T4wL/n8P1CS7I32UH1zzG1QqaYAie/wq3MmA
lXqT/Mt9FstOf88t5l518xjncG/Ne2NcYZjfNR+EwYgHRiJY3JIypd8ZJvxVniftE05HzrWzexxi
hLpuYVNLY28Xurgrv32yDoo2NkCcSz8N8ae63rbAp9u7J/Rwt624PQjMqoW2LwdNKfkc6n9G7Xji
/jdSdOcrSJodWeB4ElgBvtrlf2RnVVXn2jlWOBbCHtS6oTMbajqh9jbbYZQ47C7eUu9JQXVAhY11
y56PIyhcBRzJBTPUHfcpcDiaZ8cFfcNVGpct1M56GVKIObl3PQlw6bWYLJJkksfEVk23FqZpf3bQ
zaNxChjQlf6n48AxgxWETJRMGYGujUVvCBxdJAVOwxW2psgoKLtyNo+zzlzdfZn8St4GF7SMGaxA
x+5l8fJTrYzSTqjEMMPSrl+1twnoApUboDleNThE8R04ziN8oVjByI/lCGUCnaW7DKhx7islQb7y
AOMTkm5QiX2Bf3e4cu8u6wqkftv2tX8d7AkpO3ZJM+74BaFXZp+6HzCpEXaRaSSyWfQkWh/Pvy0S
ibdiKsWXZdjpx/36VKFpCNfnWyNBQTKKw6bmauYAY0cnbvclXzfpmE4p8wXxSD2Qt2FsEmNZ0DQe
3gEbUwYk6A5IUPv89HDMIBz583uiv5EjKi2pPcL5qoeD7aHtzXEtOnUzSDTorVi42Xm8YT7Ecrsi
okI0flqg/+Ng79neznK46ZtTrqOkKhXIjkz4bmeGH49QSAC7E+rqJhKK2RRDqHBTTE7iBqlj7EsE
uT+dAZ2dWem0TRNv6zOiFaRyrrmBBl1kQcqCpoeTOofjHu8In2iugyvDDey6BHXvv6gwTCTWnkkA
aLG8Z6gobXcIwQgL8vTS3S3TxdNRJKWGeA3ej08caaRCtYnpBPyIYtVS2Z4XauP8qJbC0+13Md6L
Dqr0JYhzYgh/Hsew0xlhnjcBJJGeJMILIGHC9hu6iUMClGWWAGoGnoaoaJQ2jVmjQZRCets/7iZo
Igl3Z4I8D2HgrhDv5C1icedY7utbR5bXuXodlQuYdgH2jmFjEBNuHi4jGwK/tkQSlb68yTcA0WWK
WdKeW9h0yQ+iCsuI8t4gNEGcgyJUC8yopzVOSiC94TiNs81dRLD33N+TEdx0ysRKqSUlHzvCgbJv
smG7/vGFOKmnRgKo6UXmDpBbEHtnHQQl1dzwVgv46Uu9HO/b9sdwRfgRPrr7CInGLXWEabmXqIc2
rm2HEC2NqQcc0VbqSrqTHgOgLWQIx2/2OGLEco7obPinI4KRfiRu3EiL2mOhQKGbm7eFNQvJ12dO
w3jOYatolxcfJEjGuwsRbjT2Z3nictWxmmb0M+N9z4yldmMsFfogc9BUCjGZF+sky7nx8kpWQznc
A0eN7wH3l9BoX+dgTn1ZsHJV8gDWTXg8d6zJQpFce708EtDIFkjwNItGiv+PxoVR6VjhvVIypp5m
KrAyQFNPVYz1PQLXUQYkOCRJt1x4yGZsqZ2saxaA06DTY3MDHLIQWis5aVaSkuBwTGEk1c03WuVm
g4Mf/aDyEzgdMMFxZZH4b2fTX0hYgevk7wyiBUcQwu0VjH2dus3c8E5yqwgWi5Ky6DsPEwBvvrR/
hJgIZ3x/K1W/1DjS87VQsxZg7ADwyHYcyQ2ORmNRFg7bZ9Z/TXsQz1R+TQyf4dy6QOdwLYvYv0Yd
muo/5NSg+sQfR0rhHC0GMzUiABBE0SbDdn5lsqrqwer9nDSr9xcw9oQDYL4TbobwwNkRbGIp6xlS
zbY6ZA8LH8BVPGLZSUgOqV/CQxt2glxtMjEt36wL5BnX87C4IU9UXz8qZfqd2GoBoyZlJ1IwPEL1
Rmn0vX1/7YBLtmOULFQt8nceYverNwgW5TdyTqETueeiq3mY4F6ZdZaLf/Az0ZHcMnNHv0xT6HtD
2BMspH5RlFnlidCU/1toIb4PRkx+KdfiWsW/na13v3U9T0UNXcf3xvz8B6ZUbh09vs/5wjsYmGAN
Mk5agFp2AoN0ffUAas6eWnYHZasrCfPtj7jz1dsv7m9KRvL9n629RjK0sLzJA0L5rGYcGfEoFB5V
NowO+DTxI0oprUFwPzP8t42BQtztljoIjDxE6bF28qbFK9H1uSJUg7i1+uiuYvZfnIoaWQazYbK7
ovMMz7Rwp6mSDmeg3FwgaCeQGEuDXyfAAFdipP0o4OVdwsQ2UNHbJGHCh7U/nix0Pbi51Kjno+Ix
T3iAh/r6wUaOd9ynR7fOqYVEzXQNUiysVfLe+TAGOJkyg6Uump/4LcH4rKlHwCGUEAcTYOP0xGXG
6js4Qa20rFPjkqZqgzPhy75rfRvhJpzx/GRH1RYrhHGf1vqwW3Y+oX/3jVAKfH2eGHo+3rXkiaIQ
TJ/IB3q1Im/6IN3Bg63BPx0v8nOGyQJGOd8eogiT/MMLMwXpnyIlg/zy5ZQB1rcR2ey5/PN25bCM
SRvHwDtMmfjtNrW2HH3h/QBVvcRHCQ4JPxHisF7yNw1gDGIQO17crv41JSseU0//v1TxwlJfmCyr
FzfeL+cNHWqV6KdxeBZycfhVR9OqQRj30en9ljpkhB88Eesm9dwQ+BZM0Fn4UYHQPcCy1DAZBmOM
oH3e7lwtYosCGWmHXNq87DUCrg2fWYS7YTid2nNPA+5g8DtrPgUYccopWof9HS6yYf/a3IQu3fSl
L2S1wyyIjHkrG4qJ9MrSfxGvguXpaVGnsSYPrdOsIICW2o0HNgtlrfVjiY+2VmVrjALMl87/7/8x
GtGkHx0TISbNnYX7NqEci0sahLjwZpDDIgOYc6HsQeujgselwCXgT5zX0Q0NYMyCutis88pKEf5B
K/1XeZ0dJNG7a8H31C42WrZ7x3rm/FGfqDuz3fSigTI1Ubfcpen5/hycUSH7700JZQ8JAk4onHA7
+Ue//765dPigcGnz1gJO+0ZLiEVxyjFpeP8go9Wh9ECwd7Jzh4GoMjSBViZq0IzL3OdfUaonjdcI
RKBDgkA9Nbtzof44Klvj7KbVEiJwN6ErJoBqcAdPrLrz5e0r8soGZQyJ5+sdZchLapPk8qJ0oIDU
3+QTq4DjNpncXgImGbZcHpPR2yg+Ofj4KMMDB5NA1/NqIOcfyNXUApplzGhrQSITj48HrdB31+JB
jNoUFG7W8kQHWusbLNA0eUYYrgXqdESfC1KLlmwOuQUihu2t8TFVzbV3YGPfHIE9zRB+H2nGncK4
C8nir0e6r2dO+YmhjLlt7GoWPp3T6i4X7d1WBy8dDE5TgTAdsSESNm/l9Zhk7nNM5GvDTw7aRNZF
+ObZd/IRgTMuWAvYT36cQs3fj/EFovrQ3jfqz5SEOvOEUDKWdIEgW93+XVm3L/ahiPmO1f++g8SB
zYGWHIkpp//V2LoEKlBcJF9+gwHIqvKDCG2FuG+wsOQGN+ItirSLVwWEni9tFWUQi3Ls8M8+e4RT
WRro1pL7HH9ny7AXYOmUUMN8dPapQv61VWfif7rnj7IOSN66/oTUbEXjePHh/ZOttcUIzar8soXy
R2SUFmO8k0QbAcJ0+7evgXdHB2kogdvGAr0kkzSDI1UuRJVZqUbBBngcAzr/66k0XZ8rn/Pb5TjD
qrrJTJz5tCby3QIymJrST1m1pfuNmybJ49GRiwTMn+93mXPUsZx6rSzRlqCS5Lxp5qzEl9IyioQH
h/KvKNwH3KN+OW0hKbCuEWSkwyXkUov8H35GVQ5f0EROyIhcUSzjg71h+c8NBdaUZF227aGW7l1S
sNfiCYv9x+IPKdQx5QN13Qacd2g9vA8lRBXBVYR6hLgk+BDrDTa9vQgcxI4hGSBtjbdXAH4wzuKA
sb9beRhs6ngaZOSeADJV5ve3N3XWBqjxShjJHvHZ8FROsCnJUM1dClsmqVNQM7PTUs1ALk53G1gL
Uivluw64xBdJEv07MB3CRRG3vZ2NqZoP/Bj8Sz1UOqSLASfB6IRrpKCj/HQ1huiTunJQLIQlh6ND
AWBpfORGVB5KwsETfr/BKVHHBV9Ia4rIScp9+GzQdTJHaGvHJsvcq0yLV3jfjiVZJ6HSH9b1x2Cb
sj6tdpmFzQBaGfgvmwzcU/wP6Kjt6E6MAnZmaoEG7eveWOhTzGr4jYO6us3VCjvVjK5wqw1GRHng
3Fa3PW9YnEAxtVH0BAtYaF1t3MIJeVCYdju9caLSM9XJs5nyvw8TeB61yRCOUJCks8s0xNb0/3oq
H3pmGv9BTe6GI+bE+R3bVVxe9FLmB/80wxC9wmiYzDyMevIyw9wlS1sD8H3H84apTrLB1vMTJ0cL
tx0QFa/jv4p8btyUKENU3MY+Oj8EnYEnkn32aOYSyGmM12FKOShMyHbVB1a14RrqueJsl0clHBMu
bjTiKwoQP5/xMDuWeCT+0Dwj4Zz+VCaXDMxz/IOned28FMfYHRsAvzu7DKcw9ZE3TAJCibEpV2Ym
hboe0qs9sMqNGw/bo9ggIKmZnwEjMvM64KtxGe51O+qyRtHLDfaDW4wB1LB9RWxs+E1R5mTOqgTw
hwiluOgtrDWVUF65WEqS6gqHQ1+FAXqtqsnYxAql7yQVVdlsOgpyEuB0n38xsLfc12VcDiwXKjMU
QgQfCaMAyVG8G9d4LhacPLs4gw5GibB/VBuir3aldE/LRqGBBdYo5CjGma7bTyhmfBbu8V/VAYcj
79yidiq/8uAtJbxP23Xp0+aDyxuef1s3u7sDyyz0uOM4BfUONiA5WzNMWKYWEhZx32vMC6ssNscL
cpc9a8dYInBHryFTGDEBjBXVlH5t8wTWh2JQASNcNVCwjw9VxE5SduQbqZwFO3xl7di6UtH/j9Iy
24JpzjET+uVXzFll+SMSSS7UopWhHlPLO9giDYndJpsmdmDAXU4RxqGHnGyjzE0gW5iwsgMam6SX
8npokoW5HP7bl5M/muXUpVC89ZZBy7SRuTmLmJ0BIZMClF/fnbFgY7e965gcIdnng6f+ZsJqZ5KI
AFp2PxlBSyfVAjb9F6ikuJtY9hnrT32obthUNwdyJiWdalZWWa6uQyGeo5pBF5HuFZmXBBaHIaj6
qDLyyPzxiYHA3On/Kt0h3cpknl4G9+FQ7hklpQ+wew6yp27/crwlHPwAc7d6IJ6rlEvnp2CzGvFC
X2pRrCvyg7OHcTtzKKRtelWARkD3AvnGU7D4zDWy21w7MVsSs5r9JSasHk/23NbsZKA1W8AKstRG
q2E3t9wDKD4dHj/y1ASFTyp+17RNBrCC3s3uU4cB0Mhy8OJOy+m3T7AwK39wB44BcEPBqBDDgbM2
JFsmSzGiIDhYxIwelOhY+or97YwiKE4qQ6IEXbBliPnZTgYebX9GPPHwbLmCwM+ZcldmxbOZ1m+M
docPK7+aZdduoX+a6A9Ckf1CycGdCxfXvC9evjyGJCFOmcPOwH1GHWl7Nt03j3wegmnPMGXSWZ0B
8KqyAkUn28mw3Ok63Rc+K+fK+M4MQP3EVNcnhLwxpmXGmtrRuuYF6Q3jQqK6WFb2sjBAc5lPFqam
6VRG3CZCHz5k3Kgf44xwiBw8ezL+IPBBGvdKkoVhrpk61TQI2R9WAjruk79ltyc0VyWQ40sxATy0
WAmJBQBlBZ3bMRYidMGKieAaI80T6aShuJZ0paro2q/O/Bvg0Lmvl6fLROBWS/cYrYHhnCk2Awn5
hayXnPKChgfbJ6zBc56+5O9uyh3mUH1AQuSbY0Yp/VRQX96P1eiSxO3W5pUOgGs7jv061i80ULuf
7t4zcy115xw8bAEH1eMIdXiVYrP4CFHOwXB/8tTCXVZKAAeEBfNWK+tqN7tIleGmB1OhQ23Bs/mk
ys66hCCyhVIQmidIFcOIbJBe0x85bLQo9J/9FepWL4RM1V4KTzVgEyESuntVkaS5Wsq1zaPgXPbQ
l9oBSi2BA8mc4/ACCKVOQEpA5TPa9iraU9lQpMEizcIPN02J1/AXZWPRHWW3lJcIrlx4bDrnwmPp
3Au/6T3Uk6m07F6ibvGzEXImo6gAFY688hjyPr8ZWUraNn9Ims/elcLUd4O6ZNPFyqEhvtbcifiV
RXO3zg9ZSWbl01LiktIKTmBPns07wvW2qDVzERyV1kIr7nsFYTPIWU4pEOvQhVHMtia/58/6QZSV
1Be5KAX4f7fZQ/c+li4l15ZRbvWBlXx31+MQKnYrQWbqI/D3oV4Q7FBH8L44dXujvbDRf252MKbo
2ONmyuIEJX92QY87NFtkdCVfnfmCe4TQanmobJRwcj/RGpcJsjOsdXe/l6+Pb7aPBC3KdtjBSIkO
XXkoIvoV4Nr/GoJoLhezL5tASh6SejSlKtYkmMGRiUKeyx8Ke45eT9GDjyuOYLL2SbmbihgTsnoE
5oH9k3vyiREa+aKgr8lcYsQOcdtPgSIibF3+GUsCgyhLUEWrpTqgBK91XlQt59MgQh8bssWtVN48
+ROmgKcxE5PIBScuyETXnYWAFHRk9zY8/g0RooASexqAZUdOaIHrghuXfMT1T7cJ48gTV9cBMhpM
jd6VDrj/ItvqLbX34ptRE5fiRBfsixrCYJ1339qKi+JSjId3NU3uDIrM1NKY+NXY5k7wtl7xh01A
bNHdPO0Osfjd5XjE/JvkOoH0gBUNZcgKnQaoxuZ8a9mnTD6htsSWY/EWDOSserQzsNNpO202DRd0
PjHEhbaePr+xCFB55t6ZC8/EVaV5DuMJbl60TbJlZMVMQ1hlKSzRNxiUDniX4H9ubEdrKcD9B9F1
q0FWrNHyu18OT413mLfYeWAHd+H+wclt5ndc7vtLi+tFw9WPvrNxe79n4+RPVBzSr2AMwdHW9BRF
PrfnPCGjNN5+sCVI/B7IsudE47Z3UgofZcy+dyswiCZqavn2jKRIsEwAflzWCrwbRzd2SpcsqaTK
AR5U/W6YPPHUtzVwLz444FdxEw7gTcP/LG4YNkuFuVi81pFLgvgmKtioNBvnL4QPjkBzpWtMiDLL
MCMH+Mmcn/dtzIdW7xLROn4oi2UEDKjBBj63XK5xoP4VxyDiGQK2kSOxIf1W/DAu/3uSgExq9kmc
6wvhyUqjT9BQR54l3ofrakhtopyQnaanTs5UZ42VngL02RZUUAAVLRvlzLdk6YijmQMAHmzUVBlJ
CpAjDjlvPyy/1WD7HqzaFz+klqpUjQ+Jod9xl9gDtcGpZYKQxIKdKWpI3JxNigPUYH9YJfC4I+I/
UMwVKTwg6kt5dVMnAwi/6hmNPOCpZ5ldtSa2SXL+8qlCUR0HKj+cNft064PcHuJ6FCQpc7i42pKk
y0sQtgA6/DkEDltoMga/wvXB+bNCU052sKUMcnsG/f+it9TaN2Mcy1ShvyVdoxAxvr+UYbfqx9bm
KYIL8ayZMDflQrxR0pEnv6ePKzIno7mb5ivSJq11StTqew9iHQjRN3b9uAJ+ZUHqQl/yuBsdBKNw
SqFGLjqwvB/LoylxxtNyLRTmaCIB7+dBpj0VZfDQmGX8yKIFpEp36bgpam022QS/91Au3al4cl95
HSjdLC3dfwuRoLBlDaLBtb9M11QcU+VJLDrCa2nXa5IX3u0nqXKCxP7Jr62nyy0cU0jqIMJD2Twl
gUen76nOq9re0UOOnny2YeK1xHSHh0pSMpRAb5jAWBwHOAKv0Zw6/nkLcdI9Oh12qpWJs1RrqObj
BC6AweQqZtd3cyz/d04RK5ZgQFqadr0hREAxBtPOxH0eHwNBg+c5bBQCvYqDv/b68HqKLfZBGSFh
DossOpGCXPweEAI6X0ZxN359sjHk4fXY3DRYEBCvJJaBpaGIP5vwZ9fq3xEFZCGQ/gQ8HR/OBS+V
3/bUCv8ynHSn8a3A2U4tqc6rsDNQ6aVV+Fxkt63qmgycVFO395P3odI/EsDf8IpUGxDfhNZXWQVx
JPOIA6BLtKniA0c0S6iuEU6hV24uS5YWFMTWx5CrAm13izXlyTGMY2ZaoZOdkDDKB52+WCvw3KT8
DqBRF9BtNY8pmFmcVKaudPAgCurTd7uTtGivB6/HX407f/7T4w3u5zCAFWCZc3YrCQVn/4JqgU+R
di6+O9WvBk9IQQZS3w+GfQToxjGIXvHbT8zlVRMgcg5q1EYAHfv2tjV1jr/rAVfoLilhGi3gtSTb
22OZW7kOO0XeSoZl+sA+7CfkkoChYIozHjdOsa8oUMn+nATtbZywqPbfYDcelO/qUBfQyESUpOr2
NQjfCZPJOezInANdUT+Z/InXHcRSPtOyS5K08H91Ggoyc4Wk03cac/FUgbVt77jJVL6//8FZ3mGu
BnMDCRp2BZKUCe4nAgq655uALB2ut4qx8RYLgERGFQQXlcRfMsSrlkHNQmlqP5UTPVm7X4hkh15e
8G4iwisuIXgMe+YG5Yhyh7n5n0SgwrfA0Q6Xpk+DqAzIiaddNe/+/rayvkWEh5xXgpEfGtYjNKzW
YzAQt3yhOQOb83DqsY7U96jcc7t2zN88Zi+t2SRWe1a8fPUtS+zIL6FkOYX5fuunVxt5BQXsMTig
Cl2snPs5vBfWjmmSfJkF4wYhMX7O1e4+blURci/s2YpTqBHHrrAjyDn7BmR93coTS6hSawpD/skG
WEDdTHsoOFbwGsXsAoqdRfl3ceECWw54XmR299rjRuVHOJOOU0GYfX6lZzIVsJKVQBfABIRw9wix
LjgkcB90z2CkOLf0DCcGsDz28ebTWuWfi5hyAV0QOnw14hV8aSrWwrpM8ITv8KnO5PQmQhKzzxb2
xqp7ws+e8Z6++24TubCRaqJrOsWahOdkTWXWqkSEzcA9vdO06FzJjM9ocMg2ixGFgmfORmWnJX6u
Vz/qt4RAvCZg+3Wixj54a6GIovNr8O8ZDvortP1i8tzzgH58LTxnK+hTfEOhDoGtOIsCfrUEfllO
SHNS5Z/YLqYJX9AlS2GdeJCKl+J8Vzc89wHNYsHmJr3UmSMuPshTE4vvkZYsg8zyjVHf9EeMb7br
drkjaQ5zgaZQkidGlMoC0cYJHa73neBBS8alIVTz60d6Jrgk0DHExOFyBpUbktQVaG2X1ZYsW7Ma
QUk54aeKR2ILJ+AOfM45AWTzdVzIWE9tqLYJpGx61Ug6oa0f3VPT0hP/mN5IQp530GlYc9u405tY
jkMQGzfePLbN3ic5cdGDbMWMlwPDOCiQb4S/SBRQfz93pEWgWJ7s8DK4warLyIB/YoJeiuDtbsOy
YD8x50eIfAOBEWRFlvZrom8IvjgClmcE5JY2pFCkN1lC7qHa67ZzV+1PXP4HZontZqthevnHIlNh
U1y99vcLTHZYLsOlGlFUjGKI85oE6vtPwXm18ADJhOLPGsym3zGELDLqvR6Y9RlO3VLbjmSY8P4i
L4i/Kqr0j1JwFl6I9NHdrNJGsXEgXJoHuZr8HvmqfudWpSPvSdnA9ISRb9bl6ZVBP01FM7jN/sOX
yROI6T1QFtDpZBT8xRZvleGxj8FqEtgQ216bedmB3OxBrzpkBJRjlHbK8HqSvUKZuLUpnr7YjMiQ
w6NbVTKZSQuv4mZqQPOYIV8MelGyXZHqaC9WCxou5L0KtNTPL7dMvEsITMiv5fMoF2/GjxmW9bD3
c+1UJ4cN+3bkFMQmc8C4H7uJFRDDddQgxgCSX30LRi1CBBBAF1WA4aw1F2A+A7QH6KrTHOhhR0ZE
KZwnU3ahDIf0yp/+9NolhfQhg+1eXd4Tbbjx2JnGr8Y1gpSMc8M2gKXiR61SkEoSO+e1PlBNmiIF
B5gPIuYQRi16zWx6lY8bloOeFZrwUgSbrK0zx1nw33Q7v5X5paZzGEVlvnyWB11m4M8NNePZnIh3
A8ldPCu2rhha6xYUlS25wygxKDl+rtkFTHerst46UqleeCcK7OU3beSDM32u8gRVvYJ/dz4JoD6E
9jhtH7RWWdAfECw7Y09W8P+5ZAtgPcyrABSonzEKHIRwe24EnLX0Yt9mppL7n0jhL3rSOCjLI/z+
hSsof2oM/M+XZjjWavSwmBve61O5zZ3PkcqlJcGJ/iMr/5EtVOiAxfuCs/feZyx162pi4Hk05eje
cKaHzyZAowDl1Qzqm6Sf3hEZXrL5PQwbRlapMvD5eYqZaV02D7iSx1QFno8cKv7gI0gauj/JKHie
0r6+Qk6VvbJds9qUCB1d77dI69Ir3iNPLpgpiE9CNnS32j2WUf1fdEVwrjE9IaF6cK++zH1A0+EN
eXya3FPCf3rBtmTB3LbU4IjfhSNxDHiqhnCB9cmn+N7BqYj7urziFbVXQplFxY0ZD9OdSDRvYuHv
O5LsxXIz5YhtRRv802vPj+7LcyYzm8meubJdS1nJdXpRiOuQUND29Ldsv9w+Ea/SMY5S3FOWPcSa
9zJbceQ7Yjaalb9q3VrfhPAzafbM2vkWP1yh8FyNHxPiCN+FUPsAEl5j5KgxJijpQm1lCdxXGKKv
CO31HRJ5S3U87/+dBVqJlsVngzDxxCDOpXu9gqbj7y7CzpzZUBmO0fg+eNqKG34APDOzJ7VlfNnr
CnQIuNXVZfylht1IGGayjm0KcRBXCnyCvrYLWOzMSsNvulaORtEURWInkZEGr8+EtaeYFIfgnoGO
1+eTTl8RDXG35w8jvHcZKyD1FRXbvoy+yCiu9ErvcKtcac4NCXAeHfFyFpLg3gBLJaS3dWjLVZjS
1n0vmvO/hpFjoQqtfNWtpuUYH/pLeUb/04JRDBkiMMWrtKj7/6uRM5gdNmY6+XLaw4/TPTxkF44o
XjZ8zBfpKHLphLdkF9kDuB5ydblG4s65lCvJZ9jVLaHQo7qWQVYEeAsDVH5uzVglpiY8p8n+ShEt
Fcf4URV4rfBMO5iFQLcA/Rq6QnxyJnF+LSNMDKVGoj1oLrFTiPy8WcgExmDj1+K63U9YTm1yOBbS
0SOxnEKIITqEOOyBaeatX7WU5nvGYIjx3FCXQNLNBJeJ+AXUVYAvzXsYAfH+3kjOgH+Gznhwix5J
5ayINDrQqDupf9orEfs+2iw+Wj9GRr3VbqUY5iA3+hY8WtLu6jBns1Hkazw9PxMwuEcjqqSDwyL5
SoOAncKdyGufJ51IFtJ77MPP3lyJbwLpfeTnz7pvaZJsZ4JkAxQ1SeHyB5of+XNB5189NJVQv/Ra
mCu+fVZYFl8Gan1T7lsGiEoqbVV0mFtyB6Lwasft34cVKIZf02J2uQD/6I35M9DSL0XewOOWHZF1
FMg7rpnPb5yGYYmpkV9Dg6DsSZg4NsLQBfAbW+YyjRcO8kTJdAFqNvAXpAyzgAov+jUtNAsmXD4I
1xgRIJQbzt/56X+Qq/PAtrOi1u483zblhmquKGVh9DjsoPPLsWEXx1ogMCbYgISfLBBLf/9xvSMN
y7XCBFl+TaJJUEe0YvYbp4+GvbVFcm/91llUohtZilIzCG/PrwhATrITeaRLw7fsUYYrFX1dJM4I
J0UMqK6izNojF1BarHk/zGcHtA2goYPcLMGu0OJNs9GyH+rhA5ZFRGdS5kY5bel8KAmnu45WrXCz
qfnnUwF77pxODl6znVUQX2EVfVkVWUgZ7WD3o1Stnq2shqjoWfEcEoZQN2C8rRMx77hDsO20Bq2w
ulrn1NYWM5lE86Qy5hQivw4z1WetC4SAQ4LIq63ck009zh2fRgYbF4izxeVB+pCwZ+zyi1lPwA1I
47mK3Ron5uGQ9wjcFIJCp6sHC+imYvi+SDX9MFsVMZDcu5w1iVrpdoZYVwGi1gAcKYPI3Pc25Hj7
Ujj4Si27SCfvh78KAHdVJ9NwZjWq1kw5eMgEcqkG6ZdY2fziKYU/0oZqW1Ys8arv9CQ3Q1J8wAXm
aOXfVvQQ0E+tFYvyj/bbrddfrPGZb0/qKXRNYqDWGkjsvDTZUxKRLw4DghUQd1xNhFqzREO7L/jH
su+jUGO8Zp8NMbXjnGFAMpIVU1SX8XWR6+DFXwrE7Qf6mNKNlvaD12aIIhwoIg5cPNsHJ/h//BdR
FP9cM9rswSEGRox9ykfsmwDAlOTK1QLRe6E2II7dIvfKDzUoAA9wOjmrbM7iYgo2xpUYOqWjv26g
w3RP1MbHm/jUyx+2jPZzYSLXklx3S/pgj/O4tvANUvvSW65VDGmocrGg657my5IG/F229KqwiWRa
L8241JHEQ7KOH8lklSE2wohLShzGRWENBisBStav+6p+0G4/7fGxRt80y2ReBWFl39IDW/yML8Zw
KCy001yK42WoE4Kz/w62ciWVeLSC3jMV2y/1UilmOOTsEWpHz8yId48LOTZCmK9lPlYdzqQI+7sT
xbuBQYwBoHRCzKkELCtEwN3BH4eFH5E6TfAa3YHrGHqup5E6U00ZkUoGGFoDH4RV2rXl2OmqM9uU
S1Q8ohrFNrlLEa+XUtm7jYju31yFcUD0FxtxxjHUY9DZSKeqfR8eMiScE9sS2T3RE9RbTLb302e/
ZtHI210l7tMAJ+JH8eLzN+lQJuSXMJT+cNXn5f+Kc2IxM4vXSUp6bEXpC6ZzvY0XwYpKxbAaMRnO
eQUYoROfBt6FxvmYmWMGWC88dfBpAsTrjWtMLyK26BhcoOuZjrKKaT5TmiiHfDQXk2xKmxUET6SJ
KrLbhlIVZG4iMW7cklQDBYZNtUoc21aaqkjk0TV4Kstch7nv5DcRaW2M8a1GxKzzOeem0w52Atyv
ZjjE+kfFkariIEjgG9tBjyaxFfe3gntWWqogstC+Zg6RACYj0OgSgKtELIH1c5O8NIt2J55Iy1En
jHRLH1GThE3vuUNEt7iNdrgaHTr467DogF8Fa7cPl/kHMPC+W7jEHxgJ61P+YrRgKxgaKlRce1GH
Kybn03883LNkZkerHr4Xf9gnUQxWplCGiI3wwt9BQsEbCdbB+KLVvS38QIlPHvjSVZFIKfQ5SnmB
M6F026il8oHGrOplRSVGpiDHVksrbH94BaP3dmbf8/S9QbBbJBar7XPFfz1mY4kPhT5mfdD/Nwls
wlXhoK7/S89kDx/h58nyGKvGtK3027fEBMlum0kUNbqE80qw4RTSVdS3M9hA1ojrdv77034Oepzg
WKwS5JeLvZiIqM+5shHJFn1gONBxb8ajTlBUI12pT9I1gwkEE8fWSt1zOonRgCPJXjcrQpSSO1QI
Znh/mol97nN+Njz9Ci7ZJQfy2N5Pb1Gg0otizZmzxHb6wZCU6jVO9I6mMzcXpFVzKe86J5WIFQ83
Gil34f7BEDG3snblV6uX08qvHPZcTB6VHdSnCIHR0jLCQBvskUjZN/Gf/DLkW/w6uPyUsKr11qu4
Aq9Sn4OlM2aj91uaSMyo1A2pnlS23vNxiVBbs6Z2B63VfUqeUYIROi/Od1kby43gGHm2qJvkO/Ii
PScOBQ2m1QMgfyIJZFEI/g0y8BqL7pYfjKheeMVNTAsPARlPqtn9gaSWNi1kZlt4pFO0+8Roaz/h
TT7tU5Yx1HH9m9VpNfKvptaFeYNqPxlg94E5HMHg1KtHpqpEAcjcDu1+5WGNBf0pVfLR6raXImEW
YEjGV3DukjkiP5+1foCHKLby0isDe+FoSiXFwEui+orrCl2s0lh/v+yVEqmKbzqerTUdUT6bwK1m
Rx+iLoxrWe5g8aGExGkBo86do59IqN4cOZFmTIUFrXQ1nKI1CTtVrakDI9vsYe1tFXqeLUNjJ8Ts
hixlx3W3CGcXuL7JVU2aaAQwgwwws4n5naiqu5b3HHcG4fjty8LOTu2fYyeYY/qkYQIGBaAuMgGe
QdD2tFlkVOErpaaIdfexsydme19rg/ac0eUwusiJSDv+C5JceHan60W7VgcBNQ3QCH2OpaSvVucm
2/cZZP2P8P/ZiI8FIs+wciJxpZOvjCuQreg5Vk0hv4D7aImYaxau4DvYyTMYAk+/RlbrT/Yzh7OZ
mK4B4kJJR5dHDPyvC6yADcKYc4NlISY3zC0upPq3Vm58CPKob+cQsT42Mp4GtkKZQC0C1LTX8Gww
7kitWIgPIV9e757B1fKoXFN5NrUI+YiQ6izvRXBrFkh9Xvsxbyk7YZauUKj40PJ+0IYCxBeinEfR
pzpAOEdYnIQH7wgEIV4DFS56cLo5Kcb/qy2HTerru0T+30mAj8QAt2ytj52N1UvQ98mVzH2dPUQk
kFaNkO7WaKtueWPMN14HNWz7wvJbqlKNsVuBNEfr4ecnuAI8oaUpsrQY9tYM+zxEhx+H82PRLFT3
ONc89FdbRZgQgvFXJ13U/WzYdh/tZz8BfIR4afzyAQTcnSZVTV1U8mMUA13NqZb8zHiFX7jPrZVi
g5vxles7nFiLtDjTxnDWO4vd6+CM1dww5RI7xe2zbdkGPwCbLJKwkBObtfI8fEhGxIHDia+TUiPH
bmbnVbLn2kI8WNXP/FaoZe+Tk/6omw/6z6wOOBo4c5S8pFzg9zOXqOw2ETn0jx+FsmXwrpABBxHC
ChAQwkQVBcFlDOmTn2OCq17zKnbahrl8sZoltAsK+me3PrgRvCW7VmcIX0q0Nxh/kw/AdBVbND/9
q7/YT7TwT0iWuF4BEbbrNu+mZWEhJLwI8AAAKfqdUZQ1ytohLcuraIi3C6/7jbNT8ynpRe4oLkrU
eQ6JKDSCBIE+B1alkWjWviKq8jpjN+JGE9ls9TXAdP7C+gGtFU4Ti97yJme3Q1o4ks7kMO1qrJ2q
9UsMGsq+Z4llsythMDON1Cp695/BzOPTp89H/NsRvDfZJKf7jlvP5/3pCkBe/kVyWZIofGdefTHq
49DW7X+/d8K/pHGqi5O6oEtB7VvfG01RC1/mgoy3Qc0NBcIw+ubfjYdfJwMQbUJRo7TjbBD9bnKr
3bW+Uijw1vW6lmPaTM7rUBkXVnI8+7E4drzE+ng4AZWzlYbJnj/Bbh3Pmvjw1a/h8FIKtw2F3w91
9mb/HYjxbR4psL+1JGfSdm7/cjpmJ5PMc3pMVEZC3F2ZzHpdlJ1lkCwpWnRS48EAoXxeW4GoB6Pf
Ethqske/hGVmq+Q0FNfKmVVu5Y4Epw4/AwhKLPMiDFdUw5UoMnpJrVbB6aC2KTEGqE6qUYiwrGhO
cK5eWqhW3Kxnrw7UUOcbGY3HxYAX38dNgF8sOJwZ4zkWU3LOdeAjmzjvDeJzJVsXdQ+RzmC7KdmX
UD/8riLsOWoE70DUG0K5SrcJETlqvLDCdyMnaUf5vGa0CKUXtuC9tisvcGHdjhr5Vy1wg3nTvhsd
R5U/3OjlTt2AFGuUrbc9we/kVVLw8TDnGGfFf6JSTkf/wWBwEYd8P8L2KpjHWKiT4rU1h+BrlLjV
6VpFCs1rdnrd4oYAXhvp4eyzumOFId7NHy0vZX8SNVvOzDc9n0bVaLCtOcK0B3Srp2I539qbBtqB
jeueqPbGLeXxkVFS3hjiFu85AcWDdZngWv3D+znyZFICK9KlArhQnXVYjdTDYS8r9FbqhM5X8LR7
GgWSy1ir36zIur0fTVphMIVebAADXT/I8oZqhtZnAvsTWdDkxOey23HtRRl2faNz6rvrtukweWvI
C2yVvngOjWkUOHdd6/UX1M3xJSaqlPNoBa9/oekK5Fl0v+gt8wfK8ImLU2VwexxA0F3v1E7ASykr
gTCKmAQzSpkWMXNyxHK3t+tFnsiHepwzmtBvgXeOf2MypAyHBnArWcYd5juQ49WgcfjddpmeXS2U
l83ewpOTRNsDwQEL3IvfTSM7FlNDw22PCGj3WvuKNUDnw5GpCMn5RYHgSX0RI2r47+hb+5bHOSC+
gXz4NWDRWqnyAWFaBAmjv1DYdLmfcbkkJOK1vrqawwPqvUkaOkA0k9dUXqLQBAXLBz8EicIzu3KK
VoY5tBMSyf9wx3+/fend1pfOI1zwjdrR8nzNbIhDpt9je5Kq5XTr23OqfYG8wr9QFu9oWIO/h2DP
Gi5RCAiJOX19GkhBJnZe4Gj/ff4rthYTbpwjs7hANa+CP/7iww2VjFWKkltXVh47k1VawnKGw6tA
iswzPLVNxupTnZP6Pqypk7Iu6c7iS/x+EbcGsvQ7Lz+SRF8QtVi7EuR3zU2pKmUh4T2UeY7TxyCr
GTp6Ytis2rEo6gsxHh9CrGImGcAKwtAZSIlnZ7PoKoFi9v67oTSWDXNv3Cek8nAYr2IBAgBOgFNm
8rfR3mG1YgQRm6JPutLyuxXYiRe0Odr1SvIubvfwjnQ1VACj7LnVB8X+6iyJNChV80gCCt+B2i08
SwaTfjbUnTybbOc0ND629Ex41nyvMM+ovwBy3ZBE5dlrt0tjdn2WS36VvflbWzOJ9s5+W9DsvCD/
zr81CUaZTPZvPcbGgI/djguswZZjItbzelw62tsRnlrp8jGQ5/wASWkh29AcK21wi9yTD4d0ixiJ
K7gBMX6xfmLY0hLaykcJUnG4RJN62Np9O+JCm4ntEKncdY0E1Upl3PMio+c59WjGVZgWZJ+maxoj
SvtZYg3QW9vfWlVyDnrH6xbD4+pHBXPtEBWie/Ey2ZYmczDTNO7JIn+fmEDTTnfDmSm7CoFdnW1+
T5+0VHkQu6UPlAo4pnHUxdjzjCG9DRiaZrkwON+iqm+5Enoi7fXXWSiTrIPKGJ+FLoshOFXUGQoh
TD597reXXj5XEcnxDVC5xGvRaIRnqjZp5zFdKsfM2N+sSpZ97aiD/CMbPNMqeK83ExXalsszEb5H
Mm0Kl2pBHGuSoScTts4U+pr26hRoJ5zf6cELiDUSX877UQdLIYqoodxn+XTvWo4FZTsfHgpkA465
/I0DeOs2b4EfMGtZb4cieGLRnXJQDpbGzkdygmCelnwxZwTbfMnqT35qNnS6VfbFgkXVWsPUQFy2
usAsHNy6fM906rEIebCvX9sD8YysIk7v/oiNbBOQSllypdqMj2KXocp6itvBm0rc4qwPFluDxB7o
wFk3T3fOEhEPWBExCV9YRIfJoAc8Sll3v8D3So8X0h3+Iuz2VCQfNjWE3yfDiCJKc8ii72QHRNZZ
Qbw3a6wmp1Q/Ry/G1x9242g0YQk/6w1Mc88ZJQyWeFp9J4Xv3c9rKhe6QDl56YLAz317L6qF6NJr
uV7BLj1VIOqHgM+jPSpgBtTl6C+fFp0xqsfmVE3G1GYZWw3SHn3negeRS35gO9hYL5ox/i+dyrXN
fev42GGYJ/8rgxoP8KUR1KlWmSltQWUgJHb3Z/NKz8Z9PDmql7BEOqdyyb+ZrVjNsT+PJw7ekDVW
5VmkVoJJXsxMk9q8ekkfv+wwyjmT1KgdmG6bP6eOGt3s7VRN26x2RmjJ1m2h5jQ7y1D6aIqdmlRI
bWuLg0e/R+CYfYj1nNzbilhiOTOvXwj05KQCvgcaE04VeVuvQ5kVyiDwTDMKFGzz1kNEugf8AgTi
4K2sbKWgteI9fDo4QYLZLo26ewVhhCEve7IMRmgqNoRwQV4+yAyEDSniC26PiSI18W2lyObtLivp
iQM3bThvSEnHYkpUJ0DZwRjcD9uGNLdvZeg/Q0fPRFIOwRfJAI2yXcaZzGMNSdB3r2GLnvRNOU68
Tqot9C1AoZtbaH/GZmaI6mQS/7i2R/9m9952CGruHgBVEXAJFYASxzt8v5GDRdVND8lld9rmYkMB
ZtDVA5UyqandmBzciT+dsSZN1Tjp1U/+1ULJtH/aUKxamaSZBRhQv0PTNUQHzZVyxNLOlrYgffs0
CShtgyp5M9X99aRR/cVOEu3YZ9SGeTVzkZUDjj/MFA0JkWRSUonyzZD45OCE5Oo4bRApqIb9J8Ms
+BegCj4tR58M46mA57YBM+H0N7klNTrPZAKeuwZd7QKZMzi3e1OHSvFInbW5PlPSCxsWm0UmoZ1J
fSSmMMD+lx3Gq/u4Qao9dPFtP9UvRmudN+iq0+Qk8bauv3YmxsF6/phBcbUddhq2aUgPoKYI2zo6
NQzq8EBZMBsypewHTzWfWlC8Wpth79LwzKNTRkckWxlMtOJX2fxyRSOn+Dc71ZK9mDEPdLGLS/o2
Xfjg4kYoELYLZh34N5Sa9fI1yZM8tEvuPaTPNIYna2YqAOEIHsV7AKEM/HQoFJzUhRkiHmG9FZEe
X4QJIJyrOH24DM0L18YxJXdE3NjOlbWdiNP2Hjla2GdU7ymMqyU8hKpsq9O69xvUfmT5V/xa1W+r
FhOMjqzwLdzWQ9FWJZeuBTgChcEZf5+t1slZX4wdEyjGtZSkZH/fPO03MC3XmE7acCVudN0/wHbB
Fuj2SB6fK4OF22x4/qiuO3sy16QaquKXrxi2sILeKDFQBi61z8YUlpam4piCTe8E+0CCbjuiifHW
MJ8l00E+fCD7bGArNP6mXZlhGG/z2zxsAcpRnr32VCFTTzsL1wMJ2RmP+lda/lGPgY74rKOd9WHR
1mUXx9qZmRhp6Tb2Q70fZYkRiAH3DYnDS78PYSOqrz3NtZGUwmfAN/K4+OGalOvgUtnzUtc1Qxnn
tuV7yPAQSAL68tEcyjTTsSRw0nriI3GQNyAgLN7oe6MA7bPAvE/5vmVw7/f3qN2iPRYK2bRBH+Cd
fZO+biaOd7OZyk+DTgouqAWx2rmfMU4z7ativAMhTDiFvQE2lELlsGSeA5DdihBK+PstNildtqhs
8G+wXu08Cga2Uj0fTdZIZiby9znnNtxLOWtApyPFgMHq/6f1m4szKZe7Rqp36MqJpdlmvX807/vq
OEq0WiNXElT9WB+NqKtKNEpU/MuQ6ohf+SqpM3GudAtePTzTx87+/LNHDm785qTUAU3K+uWj3qI/
vFJTcfKvRzb3gt65ncYvWRW+es1TaQaDPmddiuQuKXQKYSLeBNCTZ1FIjITPPtQeO1HaSF9yIpn/
xNTs8FU3FHrJpWfZvyz7L/Ci4uhtFgzHT07xJx1Z+VgIBq//Euzp3f76zzqjq8E+KRI4bGOkf7MQ
nh6SVRgXrwq3AEn+QkfgOsKRDTBEpGFAjR5OB1IA8ZVV5OR6RB0OnqbWqmHbcJrKcoRfBGclXfvv
OTqE+v/i1lui05YHEkeLRQz8i7KQWOj018HKk4hEjSbIE/2fcYAhyd2UzwOhDzfvAXQriAZSOfMC
I12WEhUvTaHvwKa2vJsincdvUUZ43hNRIrZnCRql1XRWAGFgL5HU1cxHijAfr0S7jDl0xqu69qpK
nOMojvj+BQVBXaCKaJJ5qIT12GcmhZAGA5YZ7INMJ5JkhNUtOEssnsnz/ZyQcap+d+97elDBSnTh
8Es8v3BVVMKOK3Vp99xX426lIH/tpGfRQ7dZk2FrL5FakZvHNn0y434IvoDyqGrTE2ox/yDS3tFB
qF1/+Qo5E1o49F8UIeBw/0C4LmqhD7ur6H35xYxXZatGm+yXKsqvX2boSp68a+Z/FEblrO3YSuYq
gfboe6YHRS2qAMrNhqfppqkG+4/Nv1SrCshFttwEEVH7NmX5M+/W/+IPCkNf2jer74OAQqiyWR2A
1jHClkkKOQDU8sjUAPQh3qQXZ5X2NLn/0ucUVmzupF7wS1zNRGLrmHY7HPwAtHUwSC1x41V0VhPJ
a/uyewz4swKb3Ka4ZxYaUH8VUNwHt+9Ug9zL5NWHwQU5RVaZ9YmXyz21R/owlQHu9OINEu0al6rD
SvM/cnOCwfb69QWwRWrLb1XGwjqmTg7GULBsfIZ4YF84m2Urp5ZjPYhxVLBZNryGzBfTbb3CSMPJ
or0kGA86rfhOu0pw7JTi4cH2Kd/JDhzVTFko5JWP4dEQFGmFl2liJsXqZyQgTonDb7Vaf8Gn1tlK
1mkiti1DWWHEM3I4k7Ygl97lkoKol/Q5lb0Dn+S9ahNZafe0O/bukAdKcMDoyxPklulHWn6KTDMd
KUW7/o9UGhpua/LEF4hlx83NT/PbFC+nBhMT39vKh8rxDFLES5RYDuQh5rdEdoyBiCmAUCxjeQxL
XAq8aoXodZgRW2/P3Ox0H87kN59q4zlMxK1M3zNM89w2BXWFYOmDv78LbXA4OqnLzRB2I9OXhsCS
Wf8p4ymrqjwQlesxIlsUo4kdk2DuAruAYkdUDfdVp1w7fRZXC1qTgLMKCOK78YGW4PgOerTp/ams
TcX26r/1qCAHMzd2HfuCkUunLeeY7gVbJWhOD+HuLtkz3V+jdFsfvieJC3JSr8zHmSS3rniXoV65
N38OiPmA5ve+XgOrYHBbg/gCTPZi9F0nDOLGJHahLNMku2sFdPVukZn0ouAn0iFELIn3ZoOeRJ9M
UkI9WSZeaUNhjx1KtxjupGLNtfMgY2+zrFPUGEinmnJasG+mXpG23/pOSxHa+FUbZyvrslw+897w
xBthOlG/xKXfq7Fb2W2032rO9Y68JZtLmMtXdqJ0FCDGwIurRng1yVnGc/d/zxasAaBvlN5kKz/6
PuTdOURoNgGczMxDctGKv371tEkR6ld3ZLaXemsu9mRgunCviMmtPkDVsgBi3A+ikuD7dni0/a3r
m7jS0EUsBUipfp35Vx2l2SwF/asgN+USyH3M55nBBFf+rCdDF/nYqLUJ+sv2QJYItRr7Z/nlXYyQ
x28sldo3SiKNJLZue9CzoPO3FDELWYUiX+HAnb5KgBvKKul36GMl8Hwup0Ql1+18etWPb1E4xmLm
SfhA4hxAoey7ee/4ddD4RT1ziY5YDNhY3M8ifYczYNQJn2XsJsvMowrhb18UwQs3mOmTK7s72nI2
uCy03iBJX+yGWFK7ecEfp9VnQdbPY+Nq6SSn4GjH4pWbRKnZo24kVZ0grGhT9LzD1HxniGhCEycK
4UifeYp9Z4cdU3C4Sy2Zw0AcblvsL+ibzMtUaJjyi/+U5t4o4NlvkX39HJmtUSbo2k+QmhPt1FkS
7Lx792+h0rFSwCCF+YfHOgfGIrkXGLyvw095qaJOXVNnt+vaIgH2yHno6aR5wVH5DPdkYfIy3Q8f
jWAFZxdUOVPLNWXdW0JUNsxJ0+QQbj0YQ3KtnPioa6fFM4yHyG+Vi5hN+0a7PiGO/FA26Acwzrpq
WOJyB7THo1SmZ/viGE2ExNwGFsOQ5jNzDAo+0wIypxwlhmSjXK21NMeoERetBo+txSSXwY5t9fk0
G/SBQSnAl4LpMmahQuagnMKwrTWFGFyV+/GV8+h4flXGKXW2kD0WrICHPAmmwqk05Hy7PjP2cdNB
IZSPkKEZWSW4EsVMIwF2vPs35qlVDUXx8Cs3wz0vGw933EMSzAkltlnZ13xasymbN12WuWpmdx5f
L4SPhQYChWFm44AN+suN2mun+D96A9Rlc0BwRcF8yTjfsDUtd44/hKampZOCmd/uWAN9Rcsub8ig
WTyiy7OujRFg8E4nh+7q4iraHe4LNLecpJt1VejZqZe+Erf+SaILwxXfmrVeR4b3Hsku/8WG8Y5I
DihiMlnbIThnobaKYQWV1jtLwKEWW0kpFU52tO1o6LxBsL7xygLh6gochDjVvPtVQz6r5OyavWaY
7iqfka+2miZgGBF4yxfdEvuea0guu4iOqsYU2GBlffFWjANqKeGeH8Uy1PRRPg8Il7RfvxIZQWxx
SlBdt77mEC7L/kYnIkJ8pOrIORc2N5MCIWY/FDc8YSgywdGoQKsETKNpovs6ZzXSxIA7MY3Tfu3u
jd1ZQtkYtRuj1agKjyB8m+U3uD0TaIm49VSmqiR9GeWLf4vLEw3gQorey8WduPCdp/Gk5a8ZaA3L
ApQTC9aDHCMc3Uu3BHWXckuk1DTDrMQa+CSqpSV9uOMC1iiGAFgOHFLjB1RjpBD5jXP4yHWtmLiR
LeLpB8ZmX97ONjyII48Msd1o8Ejyn/izR6TQgv86uP/eFRqTrgf1xHT7XK4shLZsaXm0VUrXAm+N
UmvoXQmK/daPHhp0Yj/kmSNWGfZDuKcIRp/G6CmT4FH5agVvCdZf06M37O8w8cSybN2B3y5HZu5C
qjsDyNiy7eonArnrG1gp3e/sMoaovvqJLrr4IeKS91FTu4UNf9LOUWMozgIRMTR2QLDhafYy97JS
UAuvkoQd7XIuij5cZz616UflZyoSMOXgDwKu6TY0kPMFTZlJqAwaxl//95F5elW3uD0lXTR/dFpZ
y2z7dE7PLc3iVGR1zoaCtBEJz6/9oKqxYa29A/kBGnlhBPZl9s1myHgUkLX14S2K03TyBQofvDjX
aV95D+pMtO4owpuxOMh/xCpy+izJfP8dYqDz/o3n5yfFVWs/oQ5SNuW3BDOkVjqfUd4o3Dvvoaes
bJAsbtovTNPl9eQffn1sISypi45xjoUFGb+miT+MBBBWG48iih18VfoJJhNXXNcM180vOG+Qf2f/
VxHKCDIK7TnbPwO2PQQcH8jk6jnR826LostYlj0kEZUk4kilpkDEmiREZHT33/8QzzCozjSyMXvc
mnKwTVwAn7YxcqgbBT08uZ+tYfSONYmH6onpFJTN1rOUt/ddiYBHH492QH1a9JcXMdZsK7rDQ38R
Y07tJTv1cHK+V84R/nY4HnM8UHwEpRG28YXBfTy++Oku823z5e3oLlsQfKniz9Nd0s0qfnkwaOun
IfzwvqEswvw+xgIQMJIBx23/8CNRlyFLztXpe5m7Qmmqp0rKqC1aVIv8m7+tV6ykw9Pwbhi1IEQa
LaiTmZyGGALDi2n44M6MfkyA44jA5BzDaDEWzEaMCNuiY30nzr6X2iO/d2R278UD2cxNnHujfprs
mf6gujaH9WkqaZ2kWjK4IyUChgxEdCoIfhjybznvEZZyAL234qVuJZ2UzZO/XxdBaR2AcIYWRDqh
Idssw+zi51uNsacb7qTY6pZJ9Xfw6Ou5R3uEkRyMFuhKZ49EhA2bsOJ1qTG5xkCzFccNlZA/BjAJ
uFSMdsBfRnco40CMvQ7hxnhVka3K1KX3TaCDzL1akaoCP2PAMt9Jdn8EOleWLlA038vqSq/S7iHr
od+W2/UZEynG1QjBwTGN6//NZckXIRQtdUW0p9CiOj9OB1H8fmCQ9Q16D82vnuVw0n7K22xmI2Z0
TVu6S3wdpWoFaXF2qTSgEaEUWOhiEoqfCZqG9jgUMxMs1xEa8G2/r7nC5xhQlHLOFr46U2B5pKqN
RqP7EV67hUMoAMv4ctn6Dy52Q6G25MBUlfwTSZZhQnBLQ6GQGXkzKzODsqVSiOhA7/GhvwKuTbDY
5YPCHlZSegb0fFyzprwPq2WLgS6e02S7zjRRmJ4c5ENTLBn7ldNKStqdCvXNkI+0On5MXlHSnT1g
mF0hzUntQzNuXSqgP78eJ4DzBkN/+T/8HwE/59SmC3OQjkW3mEhyTJNTtdpJz5bKlGxaLpJ5+Lkj
jGs3xd8hs/0GEN0HAw5ygXrVp1F8JLDiBdRrUIUTM7MG2WSHak/8YDhF7ERoLcgYwlXVNAuhEZR3
Lu7NeVGplkHRctQ80clVefvwKzjJHLVSAARudgZIIS/9XW2DUCJF43Pz4WhSOcwJOdLfllDjuYuG
AIil6VoDXcgYI8h6YVzavNcPSZFUmRlbrpFy0hRtFURCxtnqjO+CbBclVeRr13wOQsSK8YONd239
HhUjLhbvT3LeXUOat972M+oNZxD9zZ/Cid4uwJRbRWlwuhPh3X2q5+sbAT8fVYfc59PnZMHRMzpz
ZdVWV3mUlt91fJxeCX+b+1MTVfyme/u4nGUSWtJKcnI654WWk04zFeqS0kszZswSOqm9i2zZEdtZ
yRTe/6l0KZCNv3KIUZje4FouCo6MEjOWr7wfYAXZ2V9eEoMkZZsX5m66wYixXjh8YxPnS48lA48C
Hbra84XfelctxhjVfne8njgdxf7nkeSr+1cJzqKF+ZFw938TWF5ckw3vw3hHa6Z9A1K6Pz2c36Cl
DxFgfcS8HUOYIwo4RNxDQRi2O/M21zVi6Lxtlacs4YHKNu2Od+lNo1Fp5CxGjP7mRQDVEpV73dUm
4x1j8P0FeDQ2wqoxpsnQFAgS0SEq4GSTpjqrG9tbarQxTw+XYTVlsp2uCMZ7v1o5jtvYxk7x3WhS
0gJ4brNvpyKfM2Xz1IeB/OYO1yDVqvCIXHHdGzXsfCxkNAKxvQVFecZMF5fBr+nVp8n5sbvYR2Hx
u6DCDWNZRUYzmTOgdSas6aGlcZnt8vioK/24l70kyR53vYG/HCNvb4f1r4IGAQWuap5ABTsABiEm
pj4elqzjTcnvweV+Wz1vp7ImDv/EYpgcV+TTNfkXBSQ6yzhc94nqYNhSJeuAif4rlJ9b2flgEZUH
gbY6v+wLn8aGda76DJrsp0WboJajKRX+c+GGlHX1xMBh+3AAhPzVnq1FenI7cHrAOenjskWb0m7F
L2gtbHSkXBNdAS1G8HPBpMa1D/l/gx57gb6wXSY/1TExCL+gaN4YP7Sbx80KvwYhdcWiHdN+3h+H
bUr1bxcYl7A8HPEbfNgZ+k7j0Pn+931W8/xWVc8n/f6qSlopYjK3yawmIZnoUOK1QCaAweUcGNwQ
HPVCBnF7KFAFxdlsEB1zuFD/oxWbKTBk9Ssg5c9EugWXx25gM02g8jjTV9PvErX6mcZa+AQ3f85R
irr6KjJ0sKcgdGn2nbHxgW4xTovx39uV2YnAZSnZtKjiELGYZB8XrAtS+63aacxzg7Xwwjx0R56i
XxtumjdbtXI1u/6Orj26gdu856yo4Cw6z1pKTK50J+Fj1OR6Ph99eNYlVfv6SpBCVo+XnioBXAsi
mIqXbQAHi9zA+7T4lamxhWt0gTM+h3EXdrwcnA9K39OBi9QZsufex+oPBq1Z4P/RVmKM1zB6akaH
gwKi1Dy2jaro6XK+3LX/sgxi7IdrgS7wAL6aF4c1oE+Wt5NzS0QE5cK7r8j1OBv31ZwbSqOx7q1G
JI4CA5XyM8F86BYqw3tbB3BH0lMyqSYZXEFsxFdqLG8nStEnq12B1PmpQvYjHqXiZ9OCOLQoBq24
N70aDrvfbzaNAro0t5o0mYhCE1aID3FHHrOlmIifXKkrBM7F8Jey8EPlOqQfcPANp0R2gRMwAp92
8q4WgKf0ybHZtQ6+bmQMgsFysf2CL+wFER9gmpu8LKXOZuZz0d87SbvP00eXrkT9pIabt9Y931k3
9skyoTP42tmauatk9JvH9D++q2J2aYRPqhdZZ1qLww/7++mvEcqP5/Ixi45EXGXzEHGm3L9cSrst
uwPVRpMcGlna9Ii4OsiQyzQUhRrwtRH0RpsSpSLEXiWFbernh8tb2/Be1Kc9/RwIPczloRtZqG1A
hU+iE6N8hPmpEfZfdgeY/5O4iYSlixyw0G4P0BFKIIzxDkDovVWk0czBxdiF58nim2rDnX/Ohsie
ZuKp0oJ58fOGVB3g2LgfSAe/kP2JKGz5UIMMhqzUIge/ehGMN+g4iV+PXN95bZCxHxp+zldRS28D
7tAAOU3FOKaaSw2UM3MqLeYQ4TvHGxZXGNOqKsF9K9ISPY6V6nVQzpJaXFXJXif+N+G2h2gZJcxY
pjCoUgmM+x49jCvfEYnkrGGijOc377+KEYpBOut1grz3nrfXMfnFsNRxWJJFGvnNv+smODBGulc5
qZMi7pJY3eMUQhfRnAUVNmydsPBaKFBySFTEKr4HW6WO6veKGyqO1qJV2uy+Sf8kW5fMxICA7qcP
rYCf1GnKv3iHWUOXNaKdZCpX+Em2C8zvjhmX7VbRt2S1Q0iedheJPx4BC768r86uPDhDakjXnbe3
IP+ml6vGaAC2DgQDVkU/cqthSHFk+1a/1aMjQQWD3ipqztMuycxB2mR75XZ2nSZsn8gQ910fh/Tx
aMMsfBSFQVqduHCOmW6f14+YDyQJi41wvxm/0A4nSq7PlfrCAGjJfTrSIVgBOyfnLBNgzPYo49rY
9Lv9UZ2wnsijsflHribnjgelDdxw8tc1P70qvrEh4mWJTal/aT8ZAkJE3AyWFNtcjezWi7ucH8JS
pbPurALKn5eVnDy+mwk5cMdGkrGcKKMw1kVC3Qj+/Bq8lfIvsdtKGY9CN4dyKvz2l3lLzJ1M7caE
0CElgjwruHXMYjHsU1jz20F80yjK6SO5s5pOYrAvHBysKVD3EifzQYTnk2yguYyRg7DMqTauZQvs
H4T+xHe8zmzD/OpKq9RqFlBPOQQOlGZ73M7A2tfn82YspWoYTJTeDuX5S+qODQ/CElc8MDsOYKjO
D7SMrHPxibYJjAB/8a5gHv+x7fu5D693Bf7paNHsjeXUhyoX4CmJ2AyS9nyc3bTLmGvoMu6At7O+
ceh8Kxi+80fApPe/Gv+yTEIC5N8PZ55WtQpg9+GC/r7fbteCzutLhA9gmQXCcnhFB12/ULdb/r7O
EEy3CSQyVMWtMN+NUEgpU48+1EXQnCTTESkUAK4La4ffQzZulWmjQWp+lYqAtuaEoLxorwlgVnH0
Ltp+ZsisrbjIevEz6CLIU932xAL/9xFgojrl0b9goU/x1LQba8Xg++bw2nMixRuEJ3D1vKgtzo2B
KK98NHAQaCScZNHDYfp40qXOSS6sdHFSsRO6ienqtgOW8CcCR8BMfenA9MngFIxxXyLl0dKLijUm
Dn3vfcpfhLUOzI5+9usUVPfa8MZ757O+PHe9tkP0RMkk4O6rWxQeuCfgWy8eK6t1o/mvkZkALyjT
y2apbV8ujdTZ1uGzuPfS439tk/XuBdPJEdHLUFo+9f9Y/ic1+3OudlSmfMV95xtQR0+YlrcxGoBf
6HjmiPe/giP1Tqg9bccaM3EfmaU3fJlNgP5BW76R02GE51EhVsx/HfzDIyliupZiMaXWL2TcD5Rs
Y4PsONQf+b6BWnOTfWK9ugon3Ce89lgjo0ciuMLJeAHt/NlqnickwO5JwFBqFfJ1m+xcfaofsnBA
205i4REx7zsO5wOgRI/63p8cfqshTvIS24OaJ9ANNaBv1S5V7aO6ytXT2gcxtTJHkNh8ygY1as5l
X6PbrTWvmz9aUhaC/7gZYWAKRXkw1t1y4lxWIPmfvZXb5jZSadxt5Eq1Ecn8orsBG6jq6VT7qFLg
Of8/GxcTVg8d3i4AVLGZn+VhSEEpLCMwzMI/XWUHetBx/9U7lwz7/M1+m5AghNnyK3FmlCc9FKnx
X2/2TGZRVgdChpDGcxpUF76JPmCAApnp5IGcw4pq/YbTTgKOcXGLbhjfoe8L7Fhr5DYhP3LcY0w4
ZjvjSr2Y+7kb16fzVv/OleSOZGJsflTKa7fbjjEuav9LImm2numUP2V2kdZg6pkwdadhmNhIg5tj
nLFol5T0wEPkoEqVmEe984n0Qe3raLPN3prqPvl+nWW55JRZpdC7hL/dFEfW1Rd6CTBfL8Czv3TV
ZxKk6m2dhNK2GwtWQBn8ZFdJ6U87/978oq7A/lOSCFBqvmx4YE5LTzWJ1CJtEDt6AdK2BgXlY5ic
QShmq6djY8qiZCc0SRJOb+5D4L0l+58nlCD9wexc4mHi55wydvzsjJbDdbNmpn6IopYwldLVfxv/
G2BqoPCWiCJbzQHOxffuaeYCwq/E8uVIeqFV80K/C5DnPsid2KlfqOp+0UtC+uhGkqCkVzt6u7Ht
q1eQxFF4Mwy39YKW9tdSiR1vUgng3/d0+LEh31Zs44lHHyAFmbIGNe0dpY8q5uMcpemQtNRUwHmn
+T/Ub6gz/encbs2LI42+jWLJS3aJppZEi9F6wvXRHWs8kJx3COU9NDj3MzLHmO4L2croO6oejAeF
6ApZO1/DIOtn/eM39uSBW5d9HKMJmyIfXa70fheu39VaBmkGHTmaExPB9WEiIJtV9tGHn6YnfF48
PIZ0XpA505AwL+4A4vAmktaMsTJpwA1+C8r+mWMjwqtdzJkQ14/27IuJ80zaoqXdK+kgKI5UY/lk
bxyoxZvz9zUPC8l5NcOBfdmSQ//lTI/bBKNwwXqip36aHxmyzGCWXeZPoSrUVvD/jDVolegHuHWA
CxDlYXLvpvI39SIvnNLT/1+dfWbnO6EEgknUlJp4sh15w8QOvToeFjoqvvc0QgGU8fgM0tVyIsbD
ttVyzVLys+syV205EB2hnEbwk9WaqqJLKHE8rPSmHfVTWxGUXP5BfugmkNn7qme501XCwCzXDFF9
azSDCNAth3K8lLNbM/m+YP270Ei3VLh3/xcu/UH04ZUzV9MGgtUVLfGpfV+O2zO51dDwDc5ivMw7
UiAjTCedWFqp++59fplTQtKoYqlmw9BgYKPJBxHI4QRPmCMnN4TnJeYCEpjLMPZGSBz3Zv/fd4EX
Ob8plda81oS+22MgjGJUO7MMclyZeQWLLpByDJgPbBcQuANuaw92Pwlzeb5drHKYfc7oYjEqdtPG
D/hyFXsKfhZIH2IfUbnKWFAI3oXBNtgvhh6wAY5FUtNSUMceyg4tK1+tG/k4sP4Egq80pOATRf3D
a3pcwkmpGafd33Phhugh0o9LrGZYTVi4Bs/OG/N5iZq04LhW6bo6Qor9BWwoVHvG9d2w1/jJMNhr
h/elbIZ0CdDbICgvJW44ULS8AS/JfbRVDpanw95CqnnAKbT19cdRcZUfUq2mhyqZUhYSf815nEW3
B6FYqFa/jrH0UmUSGVH0ySLyG4FmMSJWmRxrlcJtqLQOq0sNFqWXlNVNP8ugfZC7WgcSD7fk3iES
PfXIl4pc8Zy3D5IJ0f2SycAV2F36BxXigVoI27idUzn/n4Om36vwH7FcGeNmeKHAFBk+cE4ROP69
6hmrriFm8fzC8Bi3Ngb0dJodbMuZh7mIKSsvRc77EvsLzPGSUgTnqG3n5fKPd4KbDz4QNjgMWr1/
9asA7eOYesoOcK4esubF3aw8QU1b4mWYEOk5fgIa1/gyzMmKvzTBaLmn3seEz6bQcqETjA7cH9uk
U6/HjSKg/hH4yY9l/PW1oN9kcvXzbLpX+nV7v6Ur/riwWPes73G13yMdykHnTnOgc4icwRToW4gf
JYqo6ZkNC75Mf8jafv7CFv0XHKlYgzHsoVnqSU0Fk2xMlwZBSSCZxBSQj30H0WZQvIAPfOfD9BNO
OF5XvBcrVDBnVBnXH3XcZK6ugp2siwzmXD9zoK+UcsD3ZefPyFC765mMyWshWme7BnLEW8amDh0W
u3MnNaVpS9+imLxLWuEwfCWlnP/c4QOtpivPDufEXe0p8h+dKVK8fV6lSeZ5aBLwylEQmpkATp3J
ku8CPae1miyqhJuv0r90C6TGEyeFqnOxfnjLIxqIdF8976NqPegjOfj7qGLTIKSLUiIE1F4hrmF6
JXwo3sEILaLEO42NYkgdaQJatTjpQaukqwso4vNCdVn+Ah0SD2Cn6sVNIR6hCEFlG7VtUg2iK5GE
qiF0NNAM7QUd/JuEg7rZ0871ZoAZHs9BfV1+Noa+0rCU8+jz39SDWvSVy1JqETAXNJFldWEwuoUJ
2Qsu0pO3iH4yH/eYYwQHNPZ6PZq10No/RWCI8zRZ9ViaT6Ywl4Y3bX6+PJ6sSgp7KxYIPB8VXHQg
Y1Djx2p1U6b23fP0KQJMLRxjp+hyI3rFguteucp4yKBvREJwY0/hhjjJyULJ+scd4GJ/e1zhh/vf
CL8KpMtIQid6qwqrHmiR39zt4jYNrjzOcvTnMVVkZWVqanfc1cyHTiTmq70tlA7uosaW+PVEg4fz
FcQpN5pHpsZzNCIbJ/XaCgivMXS8XfgadS2oOxRWiiWMZj7TTzmP93jiffUJa6H3qIIff3xKZW7i
MrSL0kUEfJnRDTX/XYnfVpVs2VJCCdKMX31NchHuTkEXCigOlPDKZXDTuI3PPBPbVTsZlQgOo0s/
bLdl6lMfodKbL2AtQO6f3Nl1qxb0RlpiP0pVs71ISOa2FC2EC2GUVCSrJVwpx4Djs1AlKJluMYBF
xUJg/PRG5AeynNVpLx8tOEKmJ9zBrTplVwbECSRauA88sB3hknfu7uWgD5nWfpEiO0tx1Y+WhpB+
lsSvz+YZHTjUJpDtkp7sftswLYv09dhx7/OvSJrxotgcg9m0THFgTv8XBNqa5gWuSV5E13orJhdd
2Gb5U2NHHZLAYfcygtrYtt1/I19tGqPNvxoukLsWvEaRo/PvCQfofcAh2CjdWZn2Zhqmn9eE8/Xr
T85AfFlZWVPrMp+eTeaK7aYuniv8JjfVWdihKPRfMynm79nA+u7dw96ptn+TPLLoqEabJskGLiTI
KWsv1z0dVexv0X50fYC602FBqde4h69oQwpCpw/N5XT6AK4VZJIOBCLMent+W3ndnV+soM1bH9D7
zqcBikDPfoGOzoaP7KE8QYyklIGMJifSpEv1jkW80dSmWnuF9q7xUx2+BIJbzivAxBulKGcegbBg
1t+/dO93t7r6fK9PwhppxfROtB4/5Rnzm0Ge1IFc+KRbHH5oDigHppCpc+zfscdq1AqfTHElQcSt
u8GYMk/PKyVn4KBZUE4Ov866760QazqXODcC49rOTmSyTKOUOJG7UYZ0LfqEc5Q0SDyRNb9E9REt
juO6ADwLh9MC/xjU923whnxqUL7spOsCtjyre88qeOTpA+evUHN5B9EpLgrsTZcQ3lOCaXVXhg+f
BaYg3BALZrSRM87oxH6SnF9fZ588NzrLNfF1X1MuIjXhc5LWTadzCYJuMgBOeWtgT9cz5lw5Qtgq
EgzQAG8csfcJMO2VCn+MJ5BqTjk3ufKtTNbhPMLAZgrMlukE+tOQfavyUgNmXi09l90gJY3icZHg
1EaMusMkHcaqvmR4R4gjmFsPJfQ8i4qIU33unHCk3NgpIjqDhjKxwEGNmmGVLZ4cxT+4iVo22Xlv
NomwmbPhPeSDdAtv7l9HMyzNW50dKA8LulhChj0hHMvRZHuMWzhGoXb9RLOMdYXSkA4XazM7NKoW
jWE1Kg4KZwQmnZu5Hi9cao73Smi1M3C/yNahTZq0/h2gF2WwgMOL4CkO7ngYmy953CFCGwa9HdNF
ifwlWiee8edBxYxeSrIXbg2mygvLLzHO+Spp1hz3F/WG9pOvNTfLlSDAzz4oS+nOTn4JHk89OfM0
o7oW4KWjnh+oOutZrH1FdLsBEHO40rled11jospnuyJvA3mfuqRYIsHIIk2reyg1phVkzsBHSpls
YNy7JvLvHfSxJrWbHo1LglOxdtVgjTcWpgq73R5mmDheOdqZa1Ui9hnmAmCbAiyMoefCrmPBfB2H
yezcn17YnFiDHya9jGBjmEFVxNHpUt77GMYv58ZK8UjJ2+Ezsx2vt0eTSkF4Aym8PdisT7ZAoft7
EfwdJLmAteGnLSyInx0uweMRt79cD4OxY7A/t5h9jSpH79nSucKA2q7UlnPLWIhGsYbONRp7cAG0
Jn97pfIc5ycFZFuDRAuUCq84NR8+y0GoBxXb5+d/nq1f6f8dKvVkgaEjKFnpa50CnX8kNmuOhU6P
PMrSxdQ/oLL1KhP+H1DiqHJJ9QoFUVLEInbTVUPM6QlLZDajbzaJoMWuOMDEoKSAryjv1sJAW+1x
FbzsFX3DkTswsf7g864PHXfy/oHKgEm9re0FGXMRhzGop0TESUAND90f2cXydc0spW4SCTVxhSsV
Cy66SLMr/n0VkVfPihVfP3OxVH7AilPRKaZvhlTYzzrSgUyZXnjTcrVrkAcFLarBRAGYf6CC3VTI
IXFqoXrwpo1jk0ABUcrnFi6Gbof5WNx0FrqW1H/SmKFPvOGbpYb7WbYWirAm/PmHX2q1YMUCF7+7
qJK2huoFB92yZtTmn0WHkOjP8lwj7T6qoYL9U5FNV6PZcBTppT5X/n5tIOcXG+F0GiiDNm7rkPDA
Zd4q/MUYEgigoDlnDpYtjhZ6wD4T4OcuXmZCcMH6OGS6NiMPqt0JEXhkK4PZrs1gDKHm+28+MOi0
qhBlYtNppoF8dEkUp+u0PmlM2loezJlzC6kLWEl3TntDVMKpyNdxwUQB3SLSDSL6aruljA3mfANh
mAkdfcLXt97dXDYhhLs6oW/MRAdo/led1LrM6bEMq6HwkgacdHy7PsPkUeYj+zbnSqhhKzW9lbF1
y8Za2qwxyDWjTExN/1parFX5XNcegDdmUOSrMFwMuAlzIYI/dJncx6bSWiozxcVBC7AgzXV83Wvv
hZdXFV0QaWi+YHuQxO/D4RXziESaPKkEsgmrABt5101aqfEyh2TrORx5fW/9eF1HnMbtvnG/4Ahb
bVvz+3XOL8NfJ+WSuGccBXK5bdSQj7ULa4FKIglm6WETbj5qezIX1kKANFLRC0F0uTKFxOA9ZkAX
WI7QUOf6uh0Zi/V7wDiJpxqj9KkzfEa/fT50bXpeMLdFejHncJyjvCoQXgNXZFPAuHXC/3PqfsrW
6hxmRT3OtDFPD4WWo478U+SNAutF2whduinCyuLqHA7HszUc2kNpONEqNloaZxrjKfMvxxTmVPTO
NPljYbJA/z7a9vw4Hl1F/kYstrdTiwsR45j61EZs/3o2By4UhA7y5Ku4x5kJrZTkeJohXSMcjQ7s
+7Jb0EQnHIBkohE+0r9Gtpxn1pfOWcEU49UW5DXduAJGNdJQiyTgUZjFbNnVFC+vyS8sSWDjSho4
Q4LhMFxBe3xUd4SF+6PdvWT2TorkdNS9Gau9sR84eXXv4/7MVRNdla39P5f7gP0kKapMbWHAWbOk
4/BKSbHPERNCsqGKS0ch6PsRDxkehsiVn+2EwMwynY3gTR7tbGYOQJ9AtCOgGgHDgbRd508ocoS3
wEQ/CEFW3Gn+0+ZV5JPgL8tmeEYKkFDjQ6rq+YgA+PZrrnXMcPxJP3QJwuaUbq36OHhE0pN52CHa
6ZW3MfX7qfCIToGc6zJHxlI0q1+4fDfRbY1ofXUgsQDnYKF4aqDuOGjbgGVbj8V+Mm4ZmREj64UO
c81uuEVYrTJ4pvkxMJZM1YHoHhuNGQWqVokIVpXimvKyfsSVDOI6OXlmbISI+86HW91SIZf/sULl
g6NUUAtwIdyL8mVlxrWGw6YfnRaS+X8NBCjaaC6V/BA54aJUGWe+sQl6yPTFmxCKFzHhildT5E+B
cxMIc2bE1PsRdnGGS1s5dyr5z0w27LOe/yKAR4qGddrrb5NuMxJNro0nHHCGoyMsi0OHSNnfaoCC
kjr+/0X8f7yZJme7nXb+629UrcTOUohTFA42Bsif681aic+3+FdxfxbEmZbf2bXJtKKt/hVnm9tj
3+y+6qVdf1jlO0fpMlH4DUuzmRhhFdEruCZxWuJ14xwmEdeu/CI5inADew8WxRFuCoR2GEDlJ3qT
rP0rlUXw6gph/m0wieg1gcKBTfAUtHheJI85Sgtura2TRqdjMwfGNg/IMc934YHRusUkTyW/TpfY
aOq236K6hxG0UKusQRa3oQwG/5jBg02+cqhiUZyHIhsn5vJjTJ27YER74ZNF9Xudu+Oz+d44odJq
BwS/NlG40MH9ja1pFocVPiHmgWvFk8qcSkY/t6kMFUo5qjVSa++Zhj+eB86SnXvYxtF1c4QeF17L
0Go/ID46uWFyNsVE1Y/DyGgxRP/YVS1RJWeInbTP7AK+hcb04/K6ZHYHE8SRK6/gal3hiG9VzV5z
xe5mLKMKOW80dqSOg4qFQIz+ONVzGqQTIHP4Uh64dRJzKyLajDdt5WkeQoxd1/pa0SuxO6i0Uarz
kl+tsgfvU7kShrpj+mqbOdIjKLAjzbzk3Eepl9o0s0wbR/J1Ot+MZ4HAxXBUVbDwW6l5933ichx0
44vDSrGf/U7nV8GaMpDPHgitA8Hma5ZqSfaEYTbz+q7hWQ7azfuUCnunTljhZbl2cu/ygURPa8MO
RwFOeOpzGFHPmnRwASiqCWfkGBGU2iHdB3j2Ef+BAl25La6KeMYW8x6QIBZc8vWL6wb2tTLrYMQh
LSmuwNF7T8TbgV6xibYKqiCneIeRNhuUCaQcoqCLt/kiBCIh4T4kby/frR9D/LQ95CeS9FLvJGUR
Sofz61aXvWIo9YVze8p1pqdmrISfgbdwoZFcqL0aM92Nt2cwz/W9XJhtBB2HSATE2HKckGhu9PJw
46cma7QskBKuGXABqFu0jz/2Z7hCyMNu7k7wAM2dpkYhZgqvUtSlzhD9GgKXi46ecyqStgTZwbDN
GMwY1NcAml4evukm8WTyVZ3gweK1EiG2sGnpP79Z2tdPYmU2zH9QnlZ5QI65gqxX7PCtAKsVGpo6
ZNEgfwPNyxj3QIoOjwvHFNAmvDx6ki+L9yMoNUhtY6cPB+AqOkV1t9FuH0uUc6+KOx3hx/2mKZqS
5TbuGH09r4Wvl8REXPRPoDluMEcsZ6aVtrOifkgB0UFeonCWY2hA3ONZ91TxFYEcyOt6s8HtS6wj
KGdUe9RT77hbOg2kla82lf9XaLlZCuh2I1Se3fkgOqBaU2ilQI+EiiMYh12qk7kG/YeP3QDLGLKo
YpEZqDJCo7LSfAD23H+PxD19O9NNXabckyRL8StlOh9F8RiiA1QF1okFb3yZzD3aqRkgf/8lVvwf
sJYO4gDX/LM/Z4JqVDLnCJZHr3O0bmG+QZkCuDXZBcvgOykbVNWNKPXmz3EYqZDelLYDw7uELMle
a0xvWW9qhivB9ZvXB57vaZkS7yIk3TkuLz1hVVzVA+Ns2jJPHmh+Ntgjk7ud0v1X5W+5So4+HPoo
430IXos4pcCu/q2fYQAW9oHnUc/hHEiQwwmls51Mv7c+rVjN+9f8FaaGkQpSjMFDl4g0Vsq1W5rg
7GHZLQkkyTPoHBFlAa8rGuyo1BsQu72I1i9UWUfWqYCcny4BGlDZaAUG5qMOw7sVU32YbWHzWghP
egfc4NqcLyaXwUmKY9u/xPO0zQ0qrrOluup0/q6ncTBP+5BCmWkWeo7g07Ddd6X/r1kkonPSW+JA
VRgbSkMDNUSTNyJrHLShL7MsIHJsjXaqqylCty7XPr5wmZ2GWJZRih9fk//k0BaA5vuyvmJQys87
HuhTN2YlS3Gtj9SRHAhEkN6zshZ+WXqUCeDcE7v5YS1FQNnwSUnDW4mIjie0uosKfteudEMftuMx
91RDUTGlZ5t8kn6/XaEMlHeCdXKIwwTA5iP8n++pvttRJ9LIpYe36PbVliH6EmaWSwRqFiu2ZtYl
qDWFPiKaymErgFtbpZi1uUNedf0zoK75rVWYn1GgJYQMZ4kGJ9iFh5ZiX4YoZUrzLwS8BAsozr3R
tnUSIBO0gBA+3s8XmoF1MUrMqpXVbyMD+ySYqsROyktjiaSR51rdKgbnSXaNDnr9hX5mzDzhnrac
dqFyq8GKGVSp/IhXGuP3T7cmZoB36S7L8wtqzt/hp+B4Nq0FByh4w44C/RMepHObScOboUrsmRVu
NeaxUUWR3aI2Jw4Hd40mhOh5+M2XCB+cgf64Sp4Gh2pkUd6DKeMUsQkAqi5XPVxVQltRE8tX/rqh
uu37LKZF58hSXBJLhPg54d9X220m2vxaeOAWpGtC4FloeqDXM5Rear68OIqDS6q2EystY/phzz4u
t/Y23pinsh30ETzy0Hm/3gFjqf4KQXV5LxP7W07q3rxRhHrg+G1zOLt2rO97mmBi2tQzYHFZqMEn
tnMocSCHu+bXZW95y4xfYxYaIou++SjX/bqtYafDgMlgRszyMQDsjoojG2xPXmarbIkvpLdxg6qd
1wc49Cw6Sp1BtKXGZkwXpXT0c1Mm3dc+vWdtaWcfS3MSpI2YymuBdHl4lA17cNhW5RUS66ySWzwV
EtLzmMkELAuv77zJUYtzUl5P7WHYIpwJisMR03OkZwo/k4+/UlRNaXGieaeIgDPTp1hHqFz4c07M
6Hw8x08b4En1EuhfHVSf6gfgfLSenSId1qsIbdjLk8iGTOGGaLBCbzY3K7yaNvl09e5e8uLOPD1B
wUHgKUN/LaNoSReN7GKaiJbhivaEnHyntqGcTqmxbLOZXEiH9Uz3/wmla3KGFEqRtX0Pu5o6GTDU
H3/kaaLV+6T100l2QjIcrkjDz+TYRHCxEIW/bx/nyH++ROvNLfKr991iOaJ3Pn667f/HvkBOOtgA
4Cz3l0tHccGy2K2P5FclBJes655mmX2cngbJLaTyj7FGJJdxYpX5f4R+knK+JDPYFJw8BIXqRdcT
RY251RGpZRb0e+AWZ34MjI2jPeBez875DHR7JCK0lCG5U7l3UdVCW7Uvd3cIDU3an0kcVrHfrJOM
pH+t1ufXxRURDn+CGr+p5AUAE/2BRJTXGnY73QysG4i4gcXbeDo+s0BPzL3WRHJpCpQDmueQFBjd
QH1GwZS63RdZDK3UwcPh90tW1Xi1wqDZj9u/P6JzRyOxN3em6/qtKWLPXZ/a3svetNfyjZWYhfgL
f2073K8jMyebtAgsWskR7VLhE3HQfAMEr/C+so2eK8rblDVDyjug3k4gK8O687I68lqjohfZvyLR
VQazPasnIp2k4zo2ZEzD5ZiAEOSRN7vllkqqpk2hv4G5oZDYUR2uJfrg+A6kfZNjuC24+eqgt/rZ
9KDsffBnkZpqmColFg5FZmYuVaeNjWlbDfMSn/wasufa/vYaecxAcIg1S1WXMiZSE/988OcebQCF
N5dWjSiwugDIv7KQywPkFzHgVs9+gjOL5JYzf9svpsH8no1nUucTwN+6YO/7vD1i66mSmR4OBl98
HtCpx+mM2ySA5/NGCV093HExLGbE5MGpPoS8Pu1JeoZQkw4omplQrAT1yM0JJuqhvqlW/A2zJGfc
FeXs/PZAx05t5zKN2+bWS8Xg/PtYUzb0FqGP7Zh1Zvq/aTaRHJ+NHi9XRwG8dTJn84qgSwUeaNzQ
YeXTEKNeNiydHROFlzSXEC0ZgCCpzBlIPXBbdTPBbJDtybIb+M9ijBMGA4GOhfH8TdtczrHrLnQv
QfPjRriw2wx5O95jc5Yj1KT5KsNSr0bZrwkgqw3csoqrMsCkUInl1d61HUJ0X5pka0Qt8vxIEMrk
1Tk71Rtg1/+FutFAXKiCOVdHYVCaV0ySLLhAZ2pbpGg3ylLkgX2ugtWLtWiG1heyZGNPM/oMylEr
cBLhUWvTzv8/3V8/pVPUZ8K5ST5gX9HEibhlUMhQDc1nlCdBNqVuqKg+oGTnocBP44eHI8P4wlnd
METNHLDnHWYwHhmgTFOUFD/a/bAhUFX7WvZU5AcMwTQCh5qswq1Shq6y29vipH2rNSBLj+5Ulu9I
7ikDHJ6AIRyvplbWXrNcZbBX0SiOwdq7C3rKdyuUABzANkTYwVpOSa9zCBfzGHFu768FCvYyTTyD
0hcQLqtKpFD0CnbjGKgx3SDkfGMcjrGEXwtuaHt6c1LKPaYV4kMaDvl1EDfsPDlf/64WQkzPvCDv
mDksPzUu5BjJO66VvnejKgowLd2Xb8/kN8OxPxpNJfoc+VXorIMu0lZKbPhoncUy+SPEVBLW3PRj
liNFvtBg9/NP2ibFKULAcfKRsMthuxgCljb3QDWendzbQ+kopaECxLtGNQbutXv9b8Yfg8Xl4SBl
7OziUGT1jiN8cpuxHPA9FSSQCgUwJRDCS/Zk+sWKySXInBMGP+4EJYiPOXPxTYuCxGAcbsKwFILY
8e4LB3oYvp14OcaG6EGe17wejHy5nzBGexVgRViZrj7bTj/TmavUEWnvyTu188TflIhYEkR0PhiJ
0w6xJwOHHe8tFN22oI+R4kyB2qDTk4c40Kojxm4feB58KqunFvgq0quIePxMkzu5MlSlEr9HJYq4
WSALpuEQ9KOBMqQf6eWl+pyxZ/BdncIHAOPCA/YIcjQPS+pqP4uZCMD+0IBxy2YoqPzMC80iwGKl
eDrypWAIX9NTwzE1A07xJElIJo+osevlL/oY/MWVpwEu+EUKt2xVhYiTfkEVgbWU5oVMOCv3ngfN
lVIlJofTx0kNRB/guNBZrTG3X1f7U6bY1AuLf0KLkKhOJtr9IB72NDmVSJjcVwWMTOO+gLEGkOfB
gEiXHoUTEXdGo4xshZmzVUsVDv3a6YXAzzYqlPavptJD5s5BSZhU2ZsPAAM3pQnlxTOnPuEd8f0m
UfNOhpbue/4yfvqdHCWfxTLS5VTnzBpvLtz+S9t/3L4627wabkDUQ8QS8KXB4KY2YqGJkX4iNUQz
iN0C9DG6JMUxWL8jT6oLzFFOyaAGJuZhbujPZtn32gO+ou19w+CL1fmQpolC65gp9TIvDmOO+HhX
MhLXEDJw2Ds7P/UboF8iL2FqPT/Cu4lEtfK48N1vePjIQmn1gGWrpw+VnHcooW+vWf5hz8v7/q1B
sMHHf9wKi+c3E+fyC4WJSPGBDUYt/ZWbwSpg3/C2t1I+v7ObmRJXyNuYn75DwyZhePyHlKM9cDzf
zjzFTvUHwAz9TJLsLTxv4pX6n/PEEPj3WbEQskyuuzVmSjv7w+wFkZHqaeW92qy15IK2YWfw/aaS
rcQoIS4la1dDVmcPTCa4G9/oaoN/ychLfmulYz8EF1FbGL15z3oRwFf32Gt6j8K8g4vtmFxDCkHV
nt1I5sUbvNzRIpo9NLLvGpvknj30BG1FNI54Zt6F2s2HkE60xqFhouAdX1kUCN7x8JchcTzV7RCf
CiVxSFmGOXxZzxKn0ZOol1dswptYJxz41302qAIm6XbbtJfeHVRrS/UUa5ZU1pjpSnvXeLAfsCV+
WgAr6/VOVmQrzdSr1UsE2UHu5kiJoFTNC/mkkNFZif93v5Ee7dhkYJC0orBTkpQGABP//Y55unh9
800SOImgwM4zHrhJFd7vODxqYApDTX+rVwU7xo/p+s66vF5v+TEjYE5o9nbBmBSudG92r/czcJYR
GUo8PzHemYhK9rDR8e+oPOTu1EQZrgQ8g833d3O2VYwdMotKI6du13PCei66/cqLRksG+R5Q6/tM
rcOTSDhZ9nMQbfxTn6jh0HoYjsx1ib7PiIij7a8FYktgMTdfPbA8jqzoiOHWpTzH7UQO+IvKaYDV
d2XdBOSNGC7pVG3q5dyXtqFgQSuTvvYht9YB8TGmk4jT2nE4BnRARefhEjZyUgqk2s9YOVph41sF
8+4RNbK7bxD59lzfnxOUrDbl0NKyrIlpdsKEGXw5jUThdHQRSIP8Gzsxsc4Y22msrN/UkGcyIT78
Qp5ml3eHmfdFn2CRpvyf6B/Keol3ZLezPSijD7XK1m9J+5OrWU2FgqZeTN4F2H2wAEAPjbhjgsmu
tgItcw2o+jpCuHt77KS03/MDzqRovWDiYw8RYnILYD9RGxVvCs/4u/T/c6WcZogvtLqB2ZoOgtC+
2Rf156+TDlx0vR5by006CdRMmH+SQ6pQSHZkAFlo8b5fCyXPpBuV/uvwUnLp8D9u1jHWovROv1s7
ffi58Y4ZkM4orWeonKuvQQnj7i565ggFPn0SBr5PC+euT7QHkC2Dk2JQb/82Arshrcaqo5kfTBEi
b5pVu7qNUM1TQeAIArdyFQigX4rmJLzxQEjKg4lXkmoXi3LRu6lHdAxVn2g+bG7JgW2bfPgbK+NF
vC3QpmGaEhFx1fPFmo/GjUkzVnIkVtJb/kwt1ksS37az1OUM2+wBvmMKrXWYCUxcIhauD7QJVIeF
wMzZ71FoKGjRG6hfoUmkPPk3VTlI2BtWqpUr/JaG64au/6xqTOxNRyqifo3NbQ6lSsFZ3ubaucNd
080Ksc/es3FNHsAWcmsxsQfcxki90Qt20Esfa3VIO56XUVwMaolLYja//zU+yAX1jrdzPA9067sG
f3tsyCYr2UU3bvSBWVwhe3Yz8YWlFXj2dMB4ITOS9XqsIze4zdUVgqA7TIaBgJbCSatTyABCifqM
3Fi+V0MfLi0WLQvfVGlUwN9xdFs8/JE/3U/OOMKdgjpRAv4FVMwmlIkCgK83pGeQuGvhGin0A+lx
0P7Y3IIBwlDshvFRP3LYUJBoEhBrTd4qipLHI3G7CjvYfsAii49gE+yz+tB42WTHq2bKIWVtwU6g
7wWVIUoxHjn8YA5d8KNbtPvQkJKk7Kz6KMqQdr6BU1C1A/qqveIBQeXLf1k6gfnfTnYAMKrAuOU/
S7gx+aMArjbzvUbrnMO5wLqlYA+v1Sji3YISikRGk5A2wUQz32fKhREQbZ7KUWjczriPBv7RbAFA
s6JzNJ3b/L4sOQsSW+5f5VY/jzDJ+r44cx84mKXXfFjMG/zrqZXQduHXmFQOpYsZ+RzsdlPTt6ol
KwAOdUYfDcJIkY6QmywKLUTK0VqIMNQ4qCXQOqCiOLI5d98r4IcMdKbSn0tp6RkihRUhkpsnv9Lf
hAGD5f+rckJnpPz9xZaddt6MmPYUrs38m3dG4OWLIZyQYIMJxOCfiv1okyoc+UBZXqTCvHa9/aEh
YfSH9wJD3GZN59TWs9j2Ez+s+e2TOdpcL1Wg/Qw839bCyZ4PS5/2QMuS3gYjpVES6hgkLgwJFtpI
oYnCDGubXCXPkqE68IHy0zGjIAw/jRyxtE+WnLJ2tvX+KRVHGn+KlSYdMuwNiEjLqMBe0VeLcJOx
icYtgvDzQPRcYIU+OdfP2jOnYYFpnEChBV6+eb+P3b1TOCkdeIKXrPgwWG3bT3UUFddKmEIyaomU
2Qh1dTk+ssaICWmLdo8BwLcnG6VDbo2TaOMpRQl93jL51wR2zRQDBZORzMdaPbiJWt6y6PD0GU9i
r0kkP7d2rTNS2CJsUfYW3qBinvQDLPk/911rZD/sfBDuKNlIfmMBnJ7v9KPD1DI6UMtsMnCdZpzg
4Ud7rr1b7bk2tZ76ibELFQHkUZOC/PmWgMe0Pe4spm09d6PwYBGaLXy3Zw11afDGbOb2SvJcH3Q7
sSPjPNoDjaLwJqBnaRCfes4xMrknT4BlY2Nuxg6Je38t5cFN+aOAELy4eedsf5C6lZwOnivZ/5yc
4QBY9CVCukDvrNvw5MgoL+6oyTImBuTMTiC6oF7haUwjJ4iY/roUrOYlFfp9vT6kpOGDHV0lBgI+
Ib0WbcZgMwkfud/IWXVszmWVSr04o4dVYQyCqr18rX6xKGHOHr4e5vL5JIIquTrZK0bWVnj8kPye
aDbj+/h7Va0CXjdhQWZj/JSu79ISq0hKlpMfmgS7OHmMD2Z8At4dWkrYnjId49mstROh3zE9rfCi
PQOvluylN1lEaX7ihXunZmTsFGKFtfef0uOBVIeqzGV2rOe0yKSlATg2ZjvVRYlbvW59Hskk8jic
vnC0CfiQLg1kloDl5MKm0vY7+JRyj+6JasQj3akqUc4g3Mk7OecwKBmdep9cNWddEQi/It1+HpoD
NWdwnNAEnG3s1sCQxccVPNttWXkEFMDVthFSdrf1uplnmAfJUst0jnkx9aehazUD465KGK8fKumb
0y0747JCVi4TQknRnXLAz+Vq2MYJ5z8ISvl9GA9XA+EmZ/Wb1eEkI3/ROoICsbqBJXsZmWQ2LqvS
vs3/fmaZPwxFun79X4yEz96GVbki5uDg0HYsKdZkoZRNwQfeTBeat5aXjXk+Hb59NJe+ne0Zj1e+
HhyUI8rco6bLWj/Wi0oPXB7ebwZ0Xowig43JZwaodxU4ts0c87DOh3U4TdxBNKtNkd5lE4vJgA18
97hhL87IAGRYc4n8oCA7sxlXR4sRL+HnIL8NG3zFlL2U5UsstkTDqowcF2/RUfxiIbpNFq/mMTH8
O0VJ5QDm29UPf3A967czA1PxUWfixdnnlFNigXn2PFrohZmjEaDz188sYLlVqeLRN4OzskfDSP5R
FXCFOPP5oyQVbmup1vlLo/PGC6fBZx5UlUiKZGMLZhIORRkTcf2wgaPBhF/BayiC8tvmPiMu8wbe
xIQhyVp9MF21BYNIL0BkV0FOOdqfl4F48CdimOLac1nDqw8HDqF6/PjqkQmQcpSQF5MneN/RBLby
JbyZ+odILdhy3TgxOMIQi2wXKnRBQ09bldayi+tm1JDgL59cfwXtba4wQ+U2maa46ShSmRrNZX3J
g/37inFI5gCgJlf54J6bw71F+cZo69qvH/ospoGnD8YLtBoxQoBZu1vBVwXTvORR3txo6BiF+F47
hMdnIYB0Rk33+K9M3xdedmo323hVAWV2mhqFXCORjfbT3qEX6RaYb0oRDyCeuqak3sqQJOwfMtSC
2w2/qpPEmUjcOTZu6QQvyoU2OiWWOQTvN98gWwVH18kn9wyZKF50de2bxtwaCFr3HZIsbmm113zX
MXXcZKvRtNsFCUREhEhQYsk0AfBh3A+TIl+D2y4WcAnSQYFB8wBPevacMwzw4Bi4ZXMiIx07c/4u
o3BDk+ImcpRAdjrnfaXiq3YLQf6171C/z0Tt+gp0Cf9SoIykByncBTWpo2LDEsZv3IcJwT+yE1Y/
Lkd4zvWW/8Yf9e/ltCplbE8w575y0j7LyXVv+GrJLtsX5Y7O1mdYflC7gQ6JGHTzsQ7lidjyWV6e
35rDSpJOUptOXqcCmTSaHTlh+YGXeh5u76dvOC9elW6+Y/ExyEUL+u/3zBeEev/dbS72n1H20X8q
hmgCBKjX5+kL+yGuZpgR7225rMBfAA53zN+KrKmvBDEf/hIN7uYTx9vzZYn3lzHYccU13SXSDlEm
WKO7rAsMVp0xieEEt3UlepX/w1alvGwGgOrUP2/e66NWLC+3qHgQKJ+quELqNhRSsTSCj3fESUBY
2ZBUGI3JCeIDYf0WQ8pcAcTw5OtE/vbdIzJIaSp9V+/17wuH4iXBM4oFYPyB0yte4gHDD/d73P++
X5wKlgkgxHToMmWNSSjhU5OFgeAZ2tQNbgJUiKLe52nHCVRms70MkbYMIZ8WAH1VrfAkqa54bvNA
oOJIS3pucKHzVbGTREcZ+HLPoDIa0kwnZCnj9+evFA2spT+/GL+Xp8qLGrlrkw4KIDMHFWIjSI42
9Av5Lm9ljzySYGn2270plEmwrqhnVgYI5opv8PEYDJ0jAC6eI2bbjC9YnxKz13/lsGFwbagDPJJj
uv2hQTwBlCex/vjEpCvyxudXseamnou41ezNL7pCuW9x1Yhg/p6O8XhHaqqMdLuhg09D7WP86iPC
Poy4kEKaiaAFSCzazJWQJioBs56eFwPt3hMhxASRt52W+bCU0ro+bi+RqH6pe4rfDVEXLVDGYPsB
Tt83C2JBPfmK1rHsD6KItHcH9shDknQrly14fYz2IyRfGOYC1TvvdGMeoSXNhcTCl+TmHqJjQfFe
Giy1h4JC/x9ucgMKSxR9o/Mz2L4bK7+HDoZszEqCRj6jtQczIs8nw40aMDp4MfX+WzsC0vMKU0Sy
qBctkDpCwI4jNiABtDc4Ytl7O+uHgP/qbjbUeBKlJIzFJ5BbqPYVc7N8aOQ0iFxNWM5VwoNmoqBD
qY9STxatiY3MFV1RavYhwA7E636SvQC//DycDEuTgtT4e2TXiAHqW+ppdAQNb8xsOb8XLHpvY3JA
+Xyypc18rDEEDM2G88SuKORs4Lcst5Zo1G422L7t3IRXUglMbwlYjjDSJnWT6qZM6FcysKOdQ8sz
H3XQ5ir9icyokGkCH5LLFQG+vu0j3Yvfdw2w8koiOCYhf0lVWOXLnsrwzSKnBchzNrgL6jqzCbQJ
D+KDR8ToDKq+1S7OuN732ejAMA8WQq5tYZhxX3esZTpiRNe1CmfNxYXsFtKmZ05sQ6+a9DjI5u7D
VJrOe5pldlEkrPucDmooySy01k1JIjd2UtYL32C+2IB0isxOK0RLd5zlPQyYkfumez771jVTi7Wb
ShiBJVNs5ayrmHIcM4dk3neZ0LWw+Mjit8rU+Ocdzo5C/oJD9AOpiFjJd3yInpe6jy58c3wNxm1N
EU3NvPLX5VWr4t8/THPn7+yXovB9CsYycu3+YGNpgUfR5RJISza5eDLxsY5CrD6ANdYGQ4VcWBHa
rTQ1G1ij+oHqGGVJ4C17Pv661srvkor3bfR7bbMB3b4pOcZpKfPFdLXh2Ab/FAcVsnIHnyn0Vlgm
Sd/rEy3/DOjYT6m0t/1JRIWZM+4fnhsC69PCh9JSOUPWXL4Jfb84w2nxNPIOcyKY0Kjr9cVEl8Sm
YA3q7o/vM7akZte5yU/jPuh3UV7yIGYCiVINLbi1O2NtpB4ZuvBegbswZ9RFO7ATNHkjjB+YTs7z
zJN8+OhSQa7rPto5P9qa7/9wZQWTGQN/LJwHNhIOIv0HJPf+6yfBm9wN6i7F9sqpuvJyFfu1t1rb
wU3JHCL8hdWAr2TKxutZYvqu5lg9pNzmETfuDGS5REWNbZGQe+1R8Gse0016T4Dz855w22KzL+Q3
I6ARifuGIG134odU9WajtJB0zGJec1PFkHBr6QgsYRKVFqCm0OIsZRfYLDQdstLDLvOhvoa2i99/
FUKyhGVRqD3pzZYI4YxA1ZmV5ySSDBErHOnpxPfHKO4RvL7RsH4s6PbPcLnZ8o+seSA+OmWY+0tT
Osik267LXGDpbieAH/2znStnT2Wi6g1fmppBOBn2Ck41kQWy+wRUO2bVEdO74aPj9UUpK+fYZXnC
5g2bPlW3oGWwutUHP35b1DlXIKJFhgRnVf1SFzB+SSB7oXJBM8uHaeuSie9SNNzOHHhpPR1pm4PO
oVVvu1fphohjYvkwVXWAwsSC5Bdag1VdBa7ssxh/namzK10HZ9jli6AhXWJuORaa3GR6p2eTb/5W
/WndsNII+ETrG+WA+u+K0vC9JjT8xfYTqN/iMIrpcwCgeVScHYPvYBhmn+gsXamyGBb5yngaVk0E
WbJvDVt95fGUUn5uTN82wYyzHZGk53GgMsM/Eu4fMpYHdveVnUnJT/Yx3ljEOeaC94hVVwdlLS8c
Z1jT7B/7WMhJpob5QAMIgWDN+6T+bIPzHjc9HtGQE5OXQBBFwQuL6ghObw9qOS9f7Yv6Gn6g6bMd
BEGYfrkQJfpXssHrXn63ieXKzMh31p6/PnC4D5cJGxleYzaE27tVqr2WO+vjGXO7yoWogtJNVHOj
Io/tR7danH4wG++8tBdbES6vbqEehG+WbnIwEGSdTi0yza44Fax7pgORU+oMA2TKWlbRRbwBgk0A
wOJotb+NC25YNbg/xnIGelDOK08CDbnmS7ygH/SpMmy7lVqt+7nQJN1fLdaHgg4UZnxDSygVejaf
6jodnWsvhJzAaCsPoczCUwj61j2l52VmoSEgrZHKbo2HSdtD8bkWKT8/ScYXlNvf7AIRQxvVWx+L
DEeuccE9PwEG2xkou78tD60mkV/yPtnUlRsoZRjGL0h4MLeZlDePl7e9nd5qcb6rSvyknBO6Sr8x
kXTvGGMe3GPPxurO8p8B1doFJ1YdZ/9+xt93zIbkEqZLr2tec8QZm4lfYTUjS5zUoTbV7C53MARL
6A5Jthy0QKy4nCQqg+bWAMrz2ssFpNhNXnbU3uegjAUglEQgBum69pAbm7rzPe/qduvop5oJ6eD6
5lF91MyBFlV1ncAYgvP6b8OCnioN0ucUQa9qHH6/T8R5D/GCF8+ddW2Doo8T/iOPt3iknUQpwuZL
upQcbQMrqEcXG7J0SAhGydW0k+TbHWj6sRBERelwp7BFW1Shj0nThMUbdFak5RgYwG97tSXU1Qip
kxjdXJVKo3R5uSL2CiXCTIh1+N3ZNKP1xJBkMuw3h76AQhaMJWjsBAFAcC++fSWPNa60rnwP9zJK
khX74s1n5UafFDeS3CAp1al76UY1Q+LH+3O1QJn4FvOhm8gKxGV7JJ/j5tFhcXiEKAiiCi41Nh8n
i5cf5jJt66gx4bE1kEhk9IfkVaDk/dxBcZPL5B0R0H1qGdPqaffvNqm7ipKskG/wxaDefhrITVcI
6hFlK8Zr4IHlM/+OBkgZT/HjHFpNg3sqPBiL9icPRDJzeXvestnvZ5XtR+Iwm5cyQy+SbAhHlBaP
63Id3KgDH+tlrC9c4c15b0ajAULkbYzo2TUIzQleM50eOtre/XLtwgp1XUpx7TZQkGy5t7no7ScM
lAAX6hoCEus6TYBsFxQjqG3yqCEx4SlSWdC5fx8RZRzsfSWmqebgI07HJsaMyVGiCPI0ZVXlyRIE
swGuc/cxgKDWwPl8KbVUf4E/H9L9t0Tfx8IAX/HvN/6Yv90vlqPwnUp4ZBnUZhaS0ZglM8pyKEFk
kIOJD1epR4fVBtqVHsZ30nwxHNDyzChFodq66+xcF/Cchezc8aZrg7qK3QP0g2BNSl1oKxzTdn6o
sretWVKerGc5QloAEmUjzu7dY+tzaUIm+7CY8AkrM8AsuK5qb7XmMBKjMoekNaw5uOAqmBbUd4KL
Cpuy5a7w004Hd5fLRDhdntiEdJY+Yy3xrbrgVt+UB3ulkjmi3nHtbsTker9FHFAbIC8xOUp8x3sO
2n4qJAL2Fs9ZPdpywcGBnREelr7y3hRg7bNdb9b565M8/b9A+wzuO/SFSOSW4p2x66ns4HIvAMdJ
9zrE/ZC7bQ9hiwgTAncaF1MncUG2G9lbXNIxb+vvcl7Iv07oqcRCD0xUjDFpNQW/nzIsMYR8goAx
aCYtPqgj5XeXRXb7QGL6L+MfDaiHGozEuAkw+78T4G89/DIz7ClT2MyvSVQfK+IXvzQDUZXA3uSQ
/8BFV0kChv/wJ96rH6bMrOjmVIkMtBXCqFvmeYkffDsCZw6alxpzn/qW13bEFM03glSI510tf+WA
ZXQSKa2jDUpe+HX5rXkzhLvXQMaxMpxnuZn0syk5UmhFLKJsGYbCKntG31Nz6scUSlAFtM8Fi53v
vc8RqIjG/tE7tqE+jrVv9Zt0a1NQ56QDfDYGvHOMdV5HT4TWlw5MplDeEz9XEQ9yOSUKzd0V+H65
i8Wb11v5gaoZ3OSYTxT3MW5f9To5+wIdE2n7kf/MwnekBTbYZMQlvXCB8Er9duyfMTNDdlL1DB4k
Mp4waUBEkIXAZqS0TUsAk1KlDZ/OMKFEUDbE7rT+Qiys3oFBPvPimt+HtODiAS1bxANRBrxp4FCx
6W3yFwE2/GLyH//WSDoNWFmnwGIOi4mX6smrMCGHFDmMqnc+rsPGse6xaEbM6yXXDKQkvpsn3NcO
BneIEPbeUWPjuw+8N9onO2janxGkle0aWRV3rqJO+KqIw/PXKgIKK/GT46AUuOCHv8xfHcmxmLbC
X6WUXima5kjwV7DX6W0AshpeZfsgerHRS1H5B240edsZse9P0RNGgd5QPkqi3+OCu79Am2zL4GG3
ryuaLtENVmLRIQSNWpHk5YLhGEYX39kfDSGpr2pwWYEG6Q9yAl5m8bFjM/1I5jfieYoxbRNOw/MM
YcjfgJdCoFr91emOjlsvU2gEzWGjHHO+OUIvQXo1NXAC3yWmJ1NIDDEPYOk73lbA3OEtvvX2aqS6
hespHTvbsIGdiNcamG4VzsXsKRDwogN9bh8MAftYg1cUPoR5KUq8efFCmdH/MYkp3nKH07vboQ1V
fNL2oy1p/En/r37GxiFTxEid58TONgGoXnVxCluWa9mdv4KMoaqytorIh/zQDqlrIvulX3hmWNtu
2Tr39lQG8/oBm3eUCUb+lHwJBH9gGkgBjk3S4PmJvBiDLIZkpRKZ0H6s4pX8GOtLhv1XAl2ApxNR
yC4mtaTjcx/VKZ2rJqFvhcZToOita9FhhOqKX6JYgYjkm8pjO+5rJOb8lqwO5nRv4LfFQqdzPKEj
arXz4wuWVow/TeC3+7Mp70oZ3MxFunn3DP3CtfQ6bJx79mGFIkbkHzz/5lzNxYFLAKGdRl/38N7N
cRAs+KOhdySV4d1b8Pe1I+h7QVTDRQ6tjf8TElJKF0Ptg+sLF+OicAjaTQCstN6+s0FQOhHwaT+1
z9hkXruWZrH/23Tqdh3so1nyjtNg0Xq2nJBcO1yMuCAMa1fpsxttTqzTZzKlSjYKvQjEhL5hoQdS
wcmwakGd04eSZZrLa8hJDfEyCgZtEsZBr9qoYWrMpl6hX2MJ87OCm0g6tX0tTugIAuRW5c423na7
PCs/jXJaonyGFaPC171fiD3PYkl+6SxBx/xXSXogcSSRDZPTQSBT2BP4tGaY3K67dEg4MzxEuAFj
LGHG46PQIlJdlxadjBx6LG46qdNAOEYDvSoLXgSAMO3dh/juOTL3PooCHBQ+nyfpBpP2BprTTWkS
Q39vjBcF1QO4iQlZ7cEytIIl8f+CZoylApz6x5RDWb+zQOMiGVY+Ta9YwELrLX/xTyEcl9WOkPT7
I5che+6qMdAsK7WasCDdOvwzaBJWpkpg5iEAs6QEL1+fzL2dNkfjZrelJKzIm9SRvDQnoVncFl9m
2x5GmKg8HXZhDPQzZ/x5QPuGSkx1dfg9eBFYNSugSnOH1UAct7ZaqeQmuKSslW5N34EgggImXz6z
oCAVGCmnom2Gb4QlECgZd0pd0DTovDsy2IwgH6RkkF+h4lEum/Az3NgMlvcMAAnsV3ItpYVdxMsN
phg1qU/ZnjgMh5b1ZbxbGZ95x0W3PlWRceU1prGV5EakeMaisiJAj/xxuxAPwn6w6Jw8pB/t+dEE
Hs5NM9/KOUyChdsVOomLF7/MDGubpoQXvMuwmnS4hItEZvf7qkah1neXY//roDjW91Di5c7rxNUZ
2C6GJ6bLzkpWcZSdUIZK9DuI7KwZiJH1R2jzPEMjvhnTbS9CymwrHVHeF70EZSg7Yeytjv+3Lf+a
uP33F8F43oVecqyOVfSI5WmOMM0piTOb9+iD+DguEu0nte6y/3sKkxUzb8nxUcAlZMg5cLNexT6L
jynIQSuphSEcCyhUSve6jYDw16s6CAZdw1dqhose97PQDU7Ug3mH2n7fp6snt4hHB//LajiI5qG1
XUrTG9c6auymKmBEDvU9BVQyxcVT/mzWxTnno2eQk9zQLe3+UneNYSP6QZogz2D5yXg4lKhcZ36/
8Ys/fjHZh4KuyCQyjVtiY5l8D7347+/5K2zyfkOIRa9cb8okhk8u78G5YYN8SSxUZMhHDtg2cFx/
c11DykQpil1UFc6UY/GOpZT7ECQaVhKD4gNyNwrAMVbhCnoBNHJ2GBvbjzt5J/tOIokyki4Nsi57
/hVy4eRtqf/tXK/KToUCe5mf2wXNrXYJE9uzuCXP4Fu0cBf5WkXWwjjL+6NAOtAMDSJ8LAHMgCbR
Rn+bqKHXiVavE0iezNq91A7p8CKd4rnALNkpT4gjqXeo0NbelbKgPJQjvOOIAB1vaJE61nergZFd
gZlhO61UcHBmwPBgqxpdUrbb3c9Oh4fvQ6ldYmu31V96bgHj49KNzW9g2ifdNVFT76lBHp7oEbCq
FZrM57DGKan4DydhjEgl8IWMUuR9HAisoR7T82a8gJmCrnrTm9jMGFAXCmNwylKmkHk0nVGtIEG4
uJytfD9CgENHYTHi4cRZnClP1m0tw5Syuw/fF4V9IrnImk7d4eMI+Aqn8vGxISWIlo3Oixmn69wQ
L9X2X/0E6xCo9+U7myKtdklCh3GXTP88s+QUOlDeXyXgpCSXk2mewsqz4qhnocHRHL8DsILppXHq
2P3Ndk3mGLdr4xuHTnob6wvcwWqoDJlNpLEsztWBp1IuxWV/+F4u8TUqrllD4AFzdhCyWLqyqfwm
E0MKG/ThLHPiHYt1BtvnbQDE/jyp4KcvPl9UEuMFjLdTS4rk+q8lUH0Zq6H7GiZcp4qa4vAabX7M
8aze1Nh7UjVB3SyvJ72X7uA/bF5YghJvNWqihYNl29AxYBlQYOcr594XHpaOG0DpJ8cq/nb0FKq7
FNQlk8kb3C2UkVytEvUQVPvatAnHXOYLgUwsYSiAiZ9ZyxWvf5e1r87GMCnzaZ9+FdK+sRNzc4Fi
Igiju0LSdHwKl9VL9+zenH4XRoTahmH92vaVVFbFWOs01QvE0cE08sAqY58/1PL9C988o0zgEJvR
kd3yMekh/BFUShuU0NDEPCYJeD3G/nQ9tbeJJa5WQjbktVzlueg1JkISgbYrQZ2fqmxWWzHf2QHD
akwJs4drLcU/kAocd7vJ06CTALzRM4LGNGae3OP56zwcO04zASmp6xQ0GdNesZ3EKAgf0dBc3tNe
+CzCdOoZEGDtgRSaLnrdcn5UCWXCAXsnP9mXy78T37W42/R5luIbbZTUDyHvBrE7MccgdBI5Drde
w72ulv+884nQ6dQ+gJ+TodNl6dy6Tnr9fpjhCdrWBsLmKS71ZLcvdPNooiTSTt3lVzlRHGHPNewP
nRfsQEGfZGie0ILP7RjgBMvYz2omtNG/MGVgNaAacBuGuwjCHq5yzVRNPgmuiHeesU4mlM612XG+
N5CPAz02+5X2OnUdUrUJK/YDNHyPtnmgL2B+r+7ODZ69FKorNETk7ApMhIpO+szKYO9nrLq5Kuqb
DesNjS1hpe9y57nxPXrza9TiN0gMZfc0dQJcNEiJ6K9bcksCYsvbUSsI8bkfdkdTEUdCmS3YLTkC
60BsQRk7pIIWG45MiDL7YLxzStjxyQquTso3132NyuG9yDIAqWd2AuQqNvzQPSdYSHo67PIxYOr1
1onuWSRnJO8++0Z/KqNeH93k6B+xdKimQo3YBoDbfuIaGYtGsTClPne64L2ceG7V2AodS8TADTS5
VQWBuWPTtExz+0Spo00PcsYVlFvZOoFMAHEN4gnZEuxfB/0mGdw80OHatgCg4BGT9jxukafk2qOB
y9QYkIr4TLy2+iBPlC4F0I78YVsb0hJty7clA6GUA2yhD9zhO2tXyROzqmaXpyODQWxG6i9vdJbw
Nz0HHOmW5qbvYc6KuTQdIGiIm5VLTavR9R6PJBzL4fCQ6z2ZiaEmK2mjq58LuC+YxuYXXzG5FdtJ
UUM2XenSkLWgcJIu2RGLo9jqaI/M1cYdflKs1VcRkfeuqKuFchJPV8l6oVs6N7K6IpCmdt7pif4J
SbSHN4tHkKM3J0VhWXrsIKJ6v4G16n2dhIVMI++lPqUWUKUpelnnx4dF2l8f3CH7alSVm5RYPPfG
kdvr4BLyym9byG/rxlbBGewdWF0yUT+iShdlR5hn0qwrGJRLYABjjAN7LsnRAadJC+j/YQItQTgs
FPe6d2gYuRC+nhEU32k5qCYP2MTTXL9Gj3dId7ptsiyyfauLIVm8++893DKIAhqkbgNiJDYrqY9Z
rusoYl0kFRE8CuSrbXgWVFjIt7XTpjN1/hLBPsu6ONDOr7FOFOGl4JH8V4cbykDs3r/XMO3mksJi
YO91B8RMOzwKYW/19vPFx/aE0Jaw5hxjzLxBxyEs8IsDOaW0oRvgWAcT0KuRFfEbc6WAIuxFt6VA
Qm3C92Les4n/N29dQXCZTmhUDh91wTRPj7zLoCjgEYS2GkUPCmy5c8ke+yA6aZ3EKUlifC7O8YeA
FAHmGKxn7ge+uDeYw4XKJSpUoKx8hXEKkLRbS0xMtTXztMAVKS/i8pANtoCkThJcfgzHo+1ezcQm
2zLnT7m0LXtWxt37RPbmk07oGSJAMBB60qc3+hZUtny9TVrIxBIcsFUXJgz7iFhkrw1EBBaB5hQo
gVPWWbohEhFtu1PCawwKQeNUmkyizwmXFfO9zQPVu4AcE4jxZSsPA6sSorJE7uQDFskHFFw8xLVi
OMhB6KC7IdwiSLpRHP1zBvkVg4boiHjGsE7/qSmT9OUGfjD0jD0OW8/i41o0z5/SS1Xw0VdKHdkK
8pZ+99HSqRqd6KdcYfeY2dROY85lLi+wxkPy3yVDC/kU/fFomfC7Lr/ayRI48rb7BAtuIcROLqfV
Y/UgsmRw9uyCVp5OpnhZJ7eO+vhxNX+GF1HA2uY6Gx25BqGiDjpjLJzZZrthChKxe6VTMDE3mmIp
ctmEMJYIHxnLokgNekpln5swDPxURu90185YOSpX1qe1LZZ/h19dgo6nIi964qr5bnU8qw0JsMpS
P6n6fwdJkQnJmVVCVgmZ3QOR1radYyIV0XN4ciM+QUSt4sHACFuCrPrsVGkbkrAc9pv8GoEUSx2P
9B6/NluHL5gkhOOSpWGpauxzdhP3tnq218xHp2ZDA4hYs/CG/4YdSza4xLpJs0VZF9rVnYPJrRhW
uIvFKS2RjN+INWmrbyCvpNyB/qh+i1g146ran8xQc8comiA0hvx15HFPPdzxoafTnkmXldaOfDTR
aclwiH9H+ZZN+xvXHPpaDPnZzLmvwbtxZyPzn2MVP8TuTyFTt4W0RjHDdBuN+9kIRQ/oISIPUZjl
ze3Cae32cgEii6v/BSdyd6yAEOmB4CvxkBNu1EsHfRH2u0P12Q6FfNhGOFUvZ5iGio/lNp/vmwLY
z/jMwXlX2khgVNFd8oD+yQ2HGxb0O5TC04TTmVI936wifTpXuKiSOk7Jo11ghzQRb6qTXPwzqEXz
i8srbBcqfFpPVHUMsoaboye/AvM+LzMFHV0tJB/V5g7Xy2aDjpvRLcOVQeDSYascupgTqhBAjyRx
PQO05sDwOOh9Ddp2dShFUZLkc6YA1690/F0AN+4/eIa/W7iFOdMfyB7kdE8utinvIqOGBQZZLt86
xgktn5sYe01G1LXhUVqHeg4+X6EX9Ph80yOh/620g95Q9uQv/fzaSTB0Fjr7pORO8StMbXbpeIbO
kH3dGeFUMtzdUdHSKd/dEsRv/EAcb5f7CYNUfsSOjUUUxQxcaYQEkFMtFHfHmhpzgHh3C5QkjOv2
+VH/PCpx07FplNyrS4kqPSIIwHZ8g1aSUODI2E2I4OTrSGZwLJUsqQKshPMJwN3NCCvMWG2iaXrg
h7vjJc3rLNycgJO5iSQ3oKEm54B7EJTZta6aOrA/p3ZNygT7zZDRhg03Y1eAji6JjAD+DDFfdVro
wipS1IpcamgdB1uzMFwi3ojrZPNjWP3knQouv4w/nXhCxE9tAx1D7yboo8+fjc1SnXBLavazNupV
/y6LnUAPNhqtWTEpv3B3gMRf0xLQxI0i5xlOZe2HPufuAq8ISXNBNUQ0QeXpldHK/nbGgoRAt1nY
Z+2Vveks0ghanPyXk3+TBPdjnQ059yQqqb49AbUBw6LRUKR4Ag//Y7kU2KfRLBSXZjum943Epmhy
m9aD2t6yTdRdZQP3KPPWIgNpwMhyb/WEk8f8crFwYAjw7JdAgzXFxGgyUwmcUjhcPJYwtxRNYamC
LWqCBGruQdUeMA2nvKLvxGsUQZDcvCzS+UKV0k8M5zBn2+eQYBRHPDwo6WygW3SXXJWncQeuWBe+
+FWuHNiXpyBIVN87jSznKja5QjV/dtmX4oiGjRhlcjZU4kG8OpGZzV0e3MGK3kt4oHUC28csZGAA
lovxjFWbZL5RZEyv9Aibx5elF2SnFBjUbLqlu6suEuce2VWefQqSP/pkL9l/BJcnhmjSpsQSiHZS
ShZYtqi+3dOx6UiHzd8+xUjjGjnIXHL9qCg0jPKl5J6AGA6oJsoIIgD5lksRUI14pc3uYNQPGkxq
kiRRd5Koh6djqBfq2ixTevUicJ8MIk8jmsOI51RMKy2dvBAWF27JWuULxOUaBQnKJ7+uuZ3sYQ3p
OTP/tuPFDGveQdOk+WcrZDyJhraVi/Tyo03ZqpuLNbobLrNwvtnwC4Rhp4GofyrCeqY7x43atFGy
F9kihX6kuVQ8sFw5CsxfXImLoj/07MLFCJE3CFeMbaYxctjcCVII9nOj9lUHVM1TzhARjTOEh0h4
yu16/PxfbX7VaQEbj+VSmwp6BBA7S+/HN3I9pStjNcPx9HlIsgMAhtBcPVU+h+PlVJ+flejLseAh
EXiGsh77J+PuP+ANGyXrbHjCxAJVe0k/siKfmuMCF5K1vur1dHVK8a9KsOn4CtpiO2GyBHUrWZrr
CRKNXfUG+2RS/L0GTauttDOzVNBlg3Hy+zW3Ibu0eyD866yK78lUp5uvbMjw4YQVNq5FSeYLg3/L
asc1hsup/mIZw+RMHgg8XLn9xLMblxC3rPLrgugVHcxVr0dlWOs6SxzpErWypNmNUWdLUO1I+AF4
x0q7FRkDvNiqdVvaSRiaeOUoc4wGE85lJMEGnp6VHLtieK7nDCPIjvsH6e0YpuleoNrhYtElsyE0
z/mJAlbJ/u4F/ucj4P4MSQ/yn3Q7t/4PiCAMmFqIIw49SoyGx1dwprq6oaHYA45cPeULPWb3HOaI
Gy+Z2Yp7/2zXRVDANzPv+zTrECbAL240bXHBqXr7/uRjC6gjA08l1RtGDJjHMijM0C4DwmHlanRv
SiWvudUm5ixWJSROmlKTckkcAXFdedyUpq1ehhertDv8UGVoigN+Er04wIRPfMOdjSroR7+5NcXN
3RDT86cPTkpayFASM0rkeqOi8KXKEWZlj2IfiE+Hhq7tyhdi4IXo5ZN66LeyXBqFX5zAnwroQUXN
8P/uOWwzQEjWRGvha9njCtrEH9RR6NBKO9BUQkqdDPoOblJVhdiMmgmzXAbwIC6bSLSi0IVLy/P8
OqEhj0vSnArEg/qGuhlaKyBVwYqeMQyd/sQvLy08PLjrLQmjRW4cxs7t01RL6jEoS2eeeJ+vKs3L
wKz+Ix4kcaAAEdNMfaGxU5/cN8ylU5nmUzAtfyhDhvnYJadu5/Gg35mbaJYTqSPtVVxQHrgqUvhh
Y0Xa1cZBdR8l4sYKYjrVB6LpCV6zIFWAPI0SfdsX3rtLlxi9yHR+1iUIzd3sl9RqEx5XT8gjAgqz
mR8Z/O1K73gCXw9zDrCj0J0Byv1u9xk/FC3QvIjuFfkuwJWE7WA9GOUb2R/ZDz7xy7CM8SZ02ydw
Bu4Qq2MD4p7+y5ee6zcbVy5oC2BrZz0zu5gsg3m1LYY5rze1K3POfLop0OLiLsSO0iloxP30Sw+t
KMI8lfL3ETseeb55dITb3jRKwvEtWxRpCLHZ0+M4rzsMRdW+CEOpo+33zCb6BKgRt3sFML6FQzDt
J6bZ6V5YMOax0CQuCv545cZ752Rt3dbP43JvFZta5PDbAzOvE7uZNRWOCKK4voIKkp0W+19ke08s
1asaQ5MgGRym9viYcnfAFzqKXicL/M/vGf8oHyx5LXjuQ+kGlHkUjlS8CmQZGVHkLl9sllnSrKPj
EBV8JwMsVb0ftylF1zF8qe/JSr5fojXNMh+nUuelXLN6sia2ruXhtrCL/YivrmJIBpO8jyZx+xeY
hNQdwN/TwuOtoYSwUtB492oLFd/S8745JzDNtq6qapFVTb0mYAE+Dv6W8HY7qkWn4mq4xUHtPvBn
GPkV4feyhQxhtOWIWUgCnZGNVQcbQmakX2W3QuplkGeKmtff9LjqwezrYy+Qu+QipGsiYiudWoLH
09bI9yGl9eWE2Ki05U08SFyXhwlbUvveqdSzOlKtgNFN142Vzz0sJDmkZj3B26upQllZYucLDX+M
kl1bctFQMdnAHro/LT9pXZ1E4rTjDVnW1IWTVkhc6rkhXdEwOdKCc5MWuks/0VJC1rvL4UvTbWgA
VqbA6VmQUPPINnz0ab0oQbVJIy07khzdVY04WaU9taVHvRWLGpSDvOw4Q/TYXaOHplOTxULLMmfW
5qRAN8phAkIJviz/tq1zo0c835TZlYvxqh7ZFyAO9Q3QQfsgQ1nHR5281dqjUxUBXM2hMLVjbjlW
SjbpgRtXi+8S1GVOeUW7kjKZpYZCMtTW7/M79Yh7huvxGoqshCleLu6tDMBEeKTJUPePKau714az
HYSeF20iJvsbogc9s95yu5X1FA1NGWu056vlY2aHCMmVx8g96nB0Sysz1bGEZ1GBa5FpzIZCDPXr
4Q+Y5NDH15enTgmkJ5OVmVTN9s7wUsQTrBewKb+c/lClYHeCosy/LPRkY/FIadq/7UrmBWqE7sop
iFeG7W+Msqz1by39W4Tx4LxRqUwm49IyOrew4mlAMK6pNaP+bgfwirmaL0eMpgJIqn4eES+GHq2O
V6eviiykSsqhyKTQzhvCzPcESwcBoBtX+uo3l3Ou3XtlvE3z1SnwuF983CVpKQrX8GCVI0q5Obw1
XOa/RQEWUwIX2IE6rAI0SDYup5WCOHgLuS6crPt3ZfQ1vRl6RMg77Sz211jMGIqy25C6wPuxez6e
lhTR7l+mjOmdbnEUJ/bV5g2dxmopE10YLbDK0gHRaw3EQmJY3QI0EFN8hSxmDDBVFPy14wbvEQg0
NfYZbeuWbnxgpQ6us5EhBeeJ6dwx0hx9lZnxTOwo7cVLJdHKGECNNvOHHFtkIgzWCNpwEQoclhpY
wGSBkAMJy617PmZvmJKzvgVeA6sXScdU5EZMc6V16jmwONxA1b7BbOIhG5zuMLyCuG8AK1Xcb2Uy
hU+d5Mcanhqi+nLARbA6YZ4EpM8hGvB0yXKIi2pSdhqmk0U2wHe801ZUH9eQ2ZlaXbrsNn4hZaRb
eQHNVYnSSeC8eOJhKbS+DD/hKMq5kqxeyJZo4ZebzQr1qo0sdj5c11XPd7IfJtpimNSBAoH4a7Ps
MXjMYWA01gdR/DZxJguaSC7rFKhSXUvHCzUkL9uulLxZCATrSJDgAuAbj+yEfGLvawrrFSP8kmYX
holUglrXjo/SxHNvGwyBb+oez4zyVXLYyyKle/Vv5786xi4Zb7OKqxuEFuenu2EnHVVmGDBrnUZ/
jcWfGx18lU/uZiTzWLUdTQBpFyDo1NsPSLGlYO5zYv8Hk4jpD05NPs1rReeNnpvtSYfI0H1EgdyN
smnBsxPwD8z+yaPAGkLkXpImXfsLR1LDJm08pTQmi4ltjjtGyZ8ZnLsLSZxJIP3kE6rjOTZ4Se+q
8LQ3untBPVloJjeRvPcljWi20+wbQTPpIvYO59WD4Logwvj1YHVCdlwznArbW+89UW3CZK7rIKUq
7fu05UlrXvwVBZBzcgCkiU1Y2qDgEYS2FgBm+QaVwcFWITwP72qrLVsLG+d0b3Ts00k1DNCBRib7
2ymZUMly337pqz8ILn4VtqRxa9yeWJrK4o0t0NyvbQq1LxG6/6glkkDZWlQzXVWMhMGJiRpj46n3
59V5vpmq6dSNbTU3pCscNDTmDWhCpRPULDlAY8yLxGoTLOMOo1qZeUvfX7NWX0CcVYH4tyerjR6/
Tv9qhtTVgLMtFpLJx1U38NogYfRWQHdk79V58P/sYfdes0zqCB/tThadj3FDmkV2+T7lie/k6qMb
M3zn+fRp9XG+KmgExA0VJBLDWw/SzBqaigJkUoVuDvD1YKnK0aKEjZKfeqKe0VK+rbLwNVGpkhOA
6qSfrUGDw+u7+AiFWmzAvsiwEiuMb361jbx1Qc5Mk7fXSLj1zovBV+SCPBJGy2qdUE/6nOB8AQQF
8aRwuA1hB0dNSZ+TB3LBJm4k9uWD8uLtrrOdoQsruiiINay1R930cdN6hSGbBHIu8eoV4/FkhCjD
0d2WCTa3nsDFSYObvOo7SrgpmndYZnbsvKdKzXML8oce23wsGsBFUVhGKsQRjIA0a8GtnXHJOK2c
quZOfeIPklQFGqm7aRrK3pbi/vKll++DZU8dIOnDXRDrizscgJ6SxDeW/h0g4sh5RcnxBY3LKljL
Yb5ivnYMoGWC4VV1BJDZW0v6tyjrms4TfChTpDI3oFAoSwQBE6cehEAOIhi3MmEKvqtk9lM3cqWW
PKVlSpSkJ7tYnYz3pWTZbPDps5bBLRTVj9VXm4WTE07OwbAAuneeJguwnf688b6ui4kBWe906LsT
m62CFqhgOQlXAVa/BMBvPMNJ6PmhDYJSXnIIpAOVLSoVsw+x+/38O41HbDrhwF8278QLgLbP5huv
a0l4lwRU4c03WLd8If5xaaIjDxCf5IQJ7ZKUXkHOYrD5Dve/UYcKSCaPRzuBtjP1VEjO4eJykAO/
Jp9B8cQ1ifO+IrgQGqgCXixVA/4BWkNOa9mcjRTNda3jRDyw6VQFNkssgKsjp57n3GuysT3IQLIU
je19kalabQBDMl32IgDgUYQPK4UO6WuCcCa3zWL59Dd592ex3rfiMYZKVZQVeMM+PYLKMO5tDLmh
vzFkSkGqOCyzfhzstMfl0Adxtb38tKoNROGnrnfVefTx0cf/T/2O4bhB+1f4eOlUilR3t+4bfuUW
f2kpTgs+bwYeKh3Zq8F3yh8QSONvizwfXbmwIi6GdbdwTQQp2Y/xQZacb6WVSdGe0VUq81LSk4Ws
3s73ld/Bemh3QUEMh381SvaWcA0W+hBi9da+/C0Mokno3H8LETYui01huxt0uGzGb84H7rQM6vkO
Zzcndo8MuSLjWfUWiH5/+het4mXpyser7WJvXO8fgK1AbgCXGWa3XJdsf//ulMVDPC/M4WrnsxwN
JwdjXpV2Qb9vkoUxP/RYgiMqeQiVGP4AeoMjGolobAA8bVJldvA1jeV93VE4rHysvUQ8nnnVDmCP
EeIwfdslRtrWuI7ZYgY13Ky1mZwY8eRFo8dqqGwilpnYDjx0S9MbYV5/pe7wN3BIkPAVWFwYL9VT
gb6mKDXY43KIPHe3VVcyJIvr+3XeUWfbFcaeLrH7EyZOxb2S4gVYh6e0yYDdP708lWMjjVFl1XDx
m3egCUUIV26fMSwYaDZz33S25SxBIzniPrJkIoyNRxoI5jnFWuzqXywn72yQ1ECzkqZ5A6jsEKIl
f7ecEmZ8ugm9Sly3gIduP6EgeJVLNeX9cdsg5R//TtBlqC86d0m7pkkjzx7aIK//KGqXdJHfyAGZ
C/ynhmdqytfpPfjAkTb9jpd0lFJMe3m66f+yW36KrLC6s/ktH7y6uRNSKFV6uBfizqQNSGLD8Wl/
W0jgDGCsvtR9qN0KfykfAeeKHkBg0UHZ6P/LuvQkF4CLqwPpNMayFqpRzy2Ex5lABEPka9dW2yen
NJpSRpFQux5FbPkroZ9W0aehxTZtQ70b1vTcRAfjp3PrrZFtr8qNyY4UHXl7mxeaqVxMY9t+a22O
FxnaBwjMgtBEQOnMroDliYCIZ6dsmGNHvws6zFwPj9gSWm2uFq/u92hctS2ReS39l1uX5lzAjJ27
/g2YiTM3IXeM01PJb99XodT6kb8LYQqXoIx9FwbwlNa4m0xRKN5KYFEcFGGZTUvJxLPIqr3pVQ1R
kjQxbFsN8ukQ9eMA+eFho0vojVqByrb1/qefZeQ+VTH9xlXrqx0b2cgH7PKzg2GW/mRDiDKydUwm
wlKmXGmbukMFY2WoZj6TMf0oFi0LrpAPPYnzpTYp3e9SjxDhlgIDY/fAuvGyyky7A2b/thFv5Bat
PoNCnkbd9k9C0jx2IeC73PqcvqyM9fIiNhRa6Sa7WQDIvTEwXvxXOjO8s7QGQH6jk8Hh9ihXSeWp
F2eiqO9AU3CbjUD5SBAmSAwnrNdu4zKCtqdSQgwYQc+1vjDiB57trgzCk4Mv+KmglUYiKZ61RMLW
UltV1tH3FuPgsBtrdYLXm0LXDAANbnad3tYX2jBIG6Jg/F4lwMqSABRtk3F5m4rxLYTW1foOqF2k
LzyhEyIuWdqlM27KMjQIUftOBISivzl06l8k0dFphYT1UTT3fL3BvaVFqnlFGHDnCoBqfxTpuntj
XrrMZP8mNZL1DCBMl2qsPZL38VTRqkqx0S2B+I6eKoLD/Ztf5tDPoIxCufhy4oXXDamdv5txZY/t
MzDcmyh9BUn8PWu3gHSU+PYjJF2/a3BC556VzNIJ2Iyn9QqydZ8YJVgU6yxLRXYRZLGpMGt+o5hV
S2vpK/CovvD7e6cSz6IPttqZ1soGY/yTl2ncn4eyOd8GFIH1kADcdjp1QbjBtSE6P7oqNl7R2/my
r8zstzyLEo1StPvnKCtqNoG5m77W0xXquRdgOdHJwIQxZVU7m1xsiEBnqgbSBiQ3Vy3RK0wysXAu
PpxLTCNjy7n2Z9jPG++VXvng+sbPOMMiI+Do1csOOXauhSPKRcvUvLVHoUtFiul3OQe+O0WPwioe
/bPpXRM+YygNIhvsOBmV1gwobzvzgcKcsxo/9ZR+S9CZEksqB0nv0dbaSG3tGukfuU+pqq8se3nT
Q8HfKxo6UpPxFVca/WdiI+KjJe31qJw51jOUzJTn3suWjpJh/Ssk5U337RC27e+oMa3C0lL28ak8
Dob9t/F5oyrI8nb0SyGCwvY0FDNBDETbFa0smK1KWX9Be/akn5GLOqnAvDeIpQVKfeeHOC0VM8vD
iCRI6oVfnz8MZMN7klW6AsGKnlXVVIHy2TzMTSzQ3TZbRtwaPYs0nEuHr/K/deDrffUN93SlQvlR
f3bduYeS+tmwQJmAPC0z6V2nr9qb1jtmM821M+44jJoEpu+E5MruqDfSdA2tOn/JVpkgnxUMQmK3
GjF/wT4EH4N0Uuo8G6Zjzwjh8Jkg7/hjYcgM8p0uKrczuHRm9iKJGho/JQqrMSoLMAwel7JRL0dz
fYux4frsxUd8ahXtFy1Q2zUFxIWJ+L5GyETOTKHjLt25wvd9YbMk3TnjIDLZXmNOEU1BbZml8irt
IIXeJliWU1Roy6ZdEuNbDOmb/J03rPJ4y1dzJI5EuDq9J06SDfejMZc2DKqU8o5vad/ufZqP6FCL
Xagjceq8KHxkZrqCJ+J/B8u3Tloh8k5OjNfHFZMg7E63klcgW/eDx+bMXEdUQ908sVh/7x+3+h/J
GmKo+tdKMHTJgH3ana5hIATexol5uiIz2z5Ud2uYcbYSiyxj48Sbh5mxXV4l1VCQzEESL1+1TF2P
16uChn4jhnKlHbTzDLLo7tFxKpyEG7+OXunMGdrA8AsVIBpnmBRqqUmjnI/Sn67wN6668RTGayqC
eFvOwG3JzRuhB2zWbvAFHwJZmDBQ4T/zk6wG/qByN44lLNfeHr9Qj7ne6S+LAqQP1FGc+Yecj075
rBO3iUuAIbc0xhiNKKIqlsQo+cciygVAP1ET6C3XK3HtyjHebT4/IiaeKIfgVxc6yfkfWTwRiEvj
FA0SWpKpl2o8u5tjx2tiQ/bWo6CySOIZfO1TU7Ffrqo44vYdWmgr0TNK2RPQPGXGWxJWgLfkaai7
DRaJhWNDLajq+r0NhnFF4jG33F8pFZ9/iOFazOv8w1h0myiSV1JVBGcE2Lg+ulJrjqx6A5re8LGU
HuPY0zuQnDaZfKE4PiZnmIb3P4cMprSiWX/m2eU1cY43KOub7vEgoC1zLlPPgrPvMl2nC7+pXFM1
xdiKqebf4p0jzvUNyA1KqfAaFG1RW34Ja/AwNyRS5yisfJQn77DHG2FnwrRqpn2fZcFR/j9o3J2E
9MNPk88ja5v4uuidCsLiWuINBRni+ReOFGqqNVjMd+PZDIEdpRuzXM6NtWHipdRcl98jbAKLTzo9
i/yuHA5uQMLyO317Oa7uUn/IbHI9ApDfM2A9x6DRRmhinH2boHVp3gVERVm30pIM/6h7laBndx8g
JaxENmk4dHPYchXM834wFqcOgOHzfg5mA8twcFqsRCZumdf0U92vnSuwZyVx9njIMuw+ejr+WOqb
paTBz3wRSUhyovdBzsUYkmtCEPJ/oFcXZ39Vuu2h78ZmzhpH1DxOQQTnJK7ITyYxMA4+kj76TuMe
eerkkcGvnb5PD3g9IkyjWugVcn29stNE1c470iL2BTBNoL+feTcBqBkJJQ9PI1eaHob/JdbdPnTC
TU7IVqGnTJzPV1ce9pVSzTwCNYSLQtVGB0Y31RMZ/ff/2E+5FIyd4LZTLEvFvvfkxQrokygKjOY1
ePMU3C8OyqEx6CogHGhjhZKZ65tyWKuCb5WQiWnxQV9EaTcRWVy/ItaOCa5RU0oUzBLPFMxpvEkt
d7quYhOjNueWhNF5CElQKvFqJ5DWzneHNc2ZgkG6zakf+925udPqbuzx1i8N8lpoKb3yU97yql/k
3Rxuj8aawbZXDONLs3KrtDIDeXcyAgrOkB97aHZqmFzy1xcOBn4QVc5Qb5senFjz+L19DKm1XHHj
FWlP6jkUoVYAXeKP53kg7A72HIupyCh9BhSOFSWgXDPz1IAT5LCH9hLfGq3j5NXGDd6e/A9TadGt
CS2yUtjtQ3CZ4vuzHJyCfEjk+6rBIAzAFHfvZnLHXeMcmjIr197/3qh63SgeklvY2P7PW6+j7nUZ
mtbegEu+iZWyyv5G8CzfBPUyozM4jfMKWD9Xmd7ZvADre1GI/XUHoaEAbA7KdpytdnMXhR7wpQnW
UOd26wJv7CFyfEc7eu0Z8PZ/2XrtV/lrPN/mZ85B9CJSxMjEx5nfJ33gsH3qQdSHkQW1A65P6lfL
0fb1K5T6lJ8VOzrk+bgoIA3S7zZLyqzgt9kKjVMnce/+mZi2bTjIXD5u305AYjg0Jgf6nhwWezpT
Z40wpLtwy2WFsndptTlJtwWVlADnlCU3CIqaanz+2/xa2/LQRDkaeuN+iUsqWXg8nLHZap46K2xs
q0QAl8f8pHX6cFWQCbVPb1IW6rJRXlWifKy/4gAxrq/xMOxVhHW0zJyYGmd8ct2QAZ+zrvnBJUNd
P9fZE/Mn+0mi8C4CHmlhGE+648aBGSE/OSNlVzTT7gFCI8Mj3UB8leGj4PPAuC/ANXAryksp15fF
Gt5D+CEZZIqfIFdCMDvbAPjc/bQqKs8eOjr+qVpjjic/jkVjmy//eD3HyajHyFr7zHCGkJUmxjtk
/N5qtChKZbJ6aQeWe2Yrp2BRBKqkogOI+B6iKYtZDaMPtr3STquKMoQOhV9eaoF8E6HvOosl1Y2U
jweC4rhzkmNexstIde2PNboo5fzbSZSBT3iLyyiMpaA42+OMNrdyUDPENua58o08bpnlxyIhkB7Y
zDsHvqTRDS2JzXVwDDMu24h0l10SqK17M93g08QNIksDeNzBI89wMnEEXm3uaHjZy/i3XoPn7t1M
CUAjJAVfJm30gCf9cBaZDCgYTZOEKdz4Zpb2oyu1RBJsWAjfyqCJy+ZNTcByiZ4ru63J+aATJvHD
V9tNMTlDmzRSwIfDmg2xFZn4USQbDQi/sBGgff/CRTYQ/ufu6B+C5qRIFbnl9plTPWB43DOrDvjX
szmp3bgifhBowsjMmBVfTq3fpkTykS43F6SWnMejOjQG0iQFVJH+gx1pV6oHm6ZohEswdMD/G25L
NSoHc92uUPJE05lN7kCXjAs01jo//z1GMXqi8UkAC9v+JRtUfCEVptznBYA9SzSJRt6K9JyCe8gF
5e8pWbEqkh7xBC/gzVS8Zl+AGucFUbdsyAxjxs0mYoOZaxxL3IWSNjbwbzMJyVNxldZwoUCC/46z
gO5wMJUXP5fA2uFfOc6GXzLVbqd8xVil65MZ+16PBzgLh8pV7Tf2E6RkbQ2/7FIJyOTkvqrtspEo
/flxrI9VKDGptC3OUmF8/mxpiyYwTAt6BGSCFCa8WBANUtkno65fTHzg0BjSudU0lA+unn1mctgV
HPd6Yf1xZeFpS3VKCkB2zN0mxnP/59M0tq/FLjO28Is6iPbwc8R7Z3RcXfSnHCdsMbHRL/zi1ErN
QPmw26VssHaNORqeZWwVcPs1h7jC3EUrFdaNpZ/kb/PKVRid2ok89lZ3b/yiuL4PpTXk3Nx2H1US
df8XnFUiqMTdXsehyx9UiB6r5tkopYlptNF5PLdJse6tv2Xy7EkoEXSsPH8eG6/5Gt68Yj7ZYPDj
EZGIlDbwbW8UpJTBzwMlzovv4SVwE9VDDgxlaucCPIdmPWFOwv9Fch/w6V9i/I5gr+KoAoie7ESF
TT1srPt9R+1m+jCRURko8pTVD82A46r7oDEEFB7wYtXomOjFF9fiINIDZvWHUUVxGcUY2L0dDRmd
yKRMDMNNmMoBXILe2Hfd4cF8+u8VE5zX8ykCWmR8oM6e8VTJ5sMPTBaPxKcZbjQ5KA7v8iespp5C
fDYQ+QNN4xWY0kDhNYCYYD8mGrnv6U4fflJIL+asSP+vl6/9ba7DQzH9O2cekpsb0rmGUUyTvRql
swx2GdVQtB3zzTVXcH91Ltk/Lrad7uoxCD2oD7BNSn3wUeUPeWtvzgYFPpeTG0w9Hn6Rna7hi9Ft
lntpli3OSquIGm05TxS116w6va8oX2U+4eLnh1X2V7OLk4Y1EKY57UFVbQhft3G2NS67O8r3w5k9
Jmn+GdeqkVDO6Epui2GZH6JTmyfwUpBuOP1lQfjnGk7fE1BARU2T74ZcXRrFgnpD7LrF+uGcZFBk
d1km2nSpuNxvk0fXzd8n03C7peMsydt/kwV/sCO9U0eQp50Kpj1SsumMy2IvXB6zeVS0CL4iKEMJ
tjlg6HEV7xUJk7Nrj6h3Qhu7c1akdSoZsZP/yhM6JWBjGzOt771QyjXQyRe587Lb6gNTzDbXvKPz
CmVt+lnMFGT85cMzq9tv2Vn9v1NdqCrbA1kboXqAm5GSXMupOhg3VBzJyr+Nr9xwCPn7dhSMJYYn
xTGuIu7jIkdCAolh2PVhJHd60hNMrpAsNVEp3aj99IAVNJMmvJ/OAJAAHzM0cTEJqyBghNNiH+OM
LWcDGrzjuGqRk/Ut4DXt9TGjl3NVua/U74SCzFHINEWb8tqOdAaEi6vsPZtQWqBuBxb5CKAEI1BH
PaRrbob7EVRZhT0z5Z1oCKk9+Q4IghnkQ9FBmTflkhTX6WbdNAAfE5en+uujCKkmkkS5jP4ZUxpd
lI9whWwloAB+g1+GJXcQEkyjysRavPKWbQMAtNOe+sQDgG22qphvR1gMHuGqY6L/RG80Q9cHmsSg
Yb8JvHio2rwF3NLaLe1odfYyPJgBEZ3yPYhOrDB9JMswPXqt7+HXQUkbGSBs256mggcgIiIFlNES
tUoLOn6XH/LD8YKpxbOdNB5S3FWcqRGyozb5dHrTx9PQg8ev3FaoXoUmUlmpdtU9Gw4hLUlix3uX
bsclwoeuIi3+pYfWBsg1DUcINLMAz7dtpF6Y4dQrFuqzjfzck2njBI2JGR5vXmI5nioTjkLv6rbJ
Ql/os1W59ZPLvjINM+SkyLOpH76pBWewzIlRfBVGoAD1vm6SfVMFFgCU7sQluW/TG/9FOK5wR8u+
23XWw2X3JCupJtwqVDI2mgjN8VxtWa+uZ/lwCYXtAfJMFlIqfjR+JS4jc+AC0ODYVjxt22ao38+S
23Zscx3Lh7BExQAa5HJRfh6syP8fQGNsqcoXSM623uxRAwcKOOmkRz5hN1kR2taHDEBxbVNXS/3u
oaVoVXuYzzGSQv+h5eLdvYEDbHvMBGsrauwKxo0qDZkebMBuZv6Fc/QDyZfyDJqqxxzURca/hf1X
wE1GKPVjigEWwGwUfgoNEn/s+IG+QY5XXbM4rrfhYh2ZPxj1lf0mJDKkWWWMkowViDMjz6nLalGZ
8UfJNmu1L8rwTTIsKX/sjkKZh3lGB3naiNydLtbmhkIccgIWk1cx54LCdsm9RsqK9yBnm/c555uP
DSYN53N46xlerbwLg9A2+Db4jGaDaXShu+lzzY84UPnieOfWrLp+CSYCjFhFVxPWqu337Ff/ahba
27Z145oWw65evIHBrckJIKIHhy5jDD6668v2s6CeEIJAaTxBAiLZzjCb7kV2nV88U8FK54hkvu0U
BCN47u343uX68M06FxsUiQqK0mgH6/BI9ujvJHLoW2WplsBUj4H7gQ+0D+cMY3jKLp4SbsFb8ocb
oGUxHEr12lBmSkVEbb5RIewajrB4nUnSMZP0JqWk7PhbI8x7xhCg7yK/Fl6MBhGGNwOiV2JLO1ZW
cjVjGVswDMBH0fd8D6IPN3CINOCTOs13msxSo/5rku+GBqDZtjTFmeFGqyALCBkYcQ8vzJfEnYgz
FwF5/CcLp4CRB0x1m2shEyIhTLYoQsITr/6aGVYMJO3U9VVyJDDr94FIyg4FMYOo12415F0gSwSv
aOzOYAGvDKXGD+8Z5jdqkY6bk+++lMc8m0FXVlzeyM5f4Y0PzAYcltNhePkPVr6xT5uz+dpj28Ti
2Rf29NjG7KqDTQhlSXyqiEzlDR2l/yaOzEUL7V939CQRyeac6W7YM0XDndHu5ch6xDxjALclBM/L
3/RPTH0MG5jP2r4meZZI+6w+7SZygrWpzsnmY5O3eJO2eCF6Ao+Dz/mDjMB/BcirTrQqoR7STFTX
sa4yaoF/K3v7vtvW61JKF0gc2togioUisGMVqYYWehfAMxMpwUTi0pDIahSpZub458DAuH3Ya9VH
gcRD2ri0Kk1oLroGvJZsEkN11E4MHwvME1lyyleZQXLjZ7IqPXahTTLOnN6wvQeVsrU4usH5yibm
GW+vIqACqKUhwXMGNXeBCw3s0fgIV3nrRf2OQvYOHJuLcvy/7gXpc1n/V/ND5MpO8umB41CzjCt0
U/qW+FK8f9cL82Jh1Xft16B8UBOeI7RZy5FBjU/BbklGx9CEHPJzIFdUvAmwp0kuKcIU/o52btug
Bfq5AmysY3M7m6Dg19Eu0+Due3f1Tb68TADdJKoacAQwevv8xFu+736QVWBqzc5rt/080zxpLkSz
wd8QoWyxtawjhtS1a3Ward/mxnDFWMCiKaDMMwRG9U6oFKcpTNfXmMr4oLtREXY0TEeDoj7YqaHq
Z55L5nBfRqav97I7/6O8pjnyb4D+S++4wDrGgnIdPDyVCrkZf3oHGQ1d+PvvyDr0bC7dpr6QAJVJ
Hz3IW3taVyfpvmDa9WcprNtEZoCslv49wYaG3VMcIzosFwTlTUZojbS0g0BwPVSrORwiA8TRVgRC
ra0KYgDgdHn7rlbmSHFaH3tJJLkdY6TtMGHkII4Vu4xXyGqzQ069E+95X5W9WT9S0Be7vZJD4Qwr
aI2zLiF6MAFW2uIeMOGpUs6gYWx0+9TjOiwhI7SIhrJFBtlKMNUvCO360/fugPTf+m+Qc1qul9eb
NW7a7ojoah5paKERTPfUohd86XSXvrh1PLapg8O/RLV3u2x+r9V22GLUi/QqnkjUUfNxv6a1clWn
KLUCtF0mj1306bSzTZZQDgzaAhxuWvz+Ww2fMxaH1bHA+1S+4sFkdIKivj5XLqm3oNqWPRfxJ3um
RQW8VK4sOrigy9cViAOzoO0pA2WZiVrUX+LzBNNuKiCWEpMtrqIKuJ4k5T5K9ng26+3qz2GgH9fe
xx9oVzpsAqah9ulQmuTZdE4dZ1kotQBAq7neF3RzZTU84vt4KT0X7jcX6pDHhjIV34mFJiMS+n6O
cit7Dau/NikWIsQRFpIzm1cQJSyG551fBUw/6XDesQq/M6UtslFE+eamygbyryOHV871vwQcwV7N
J20v/HLhy6b9D4lfPABqjEirg9VmTLRBXC5qvh3vM3v9lsa63IsgqwPeXJlJePla6kSd3nWOdqq4
sKhkES/EXiT/wKWUdezAmz19Wi1rmgHLfob9swJrohDV/gbEcw==

`protect end_protected

