------------------------------------------------------------------------
----
---- This file has been generated the 2019/05/06 - 15:19:36.
---- This file can be used with modelsim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 3.2.2.0.
---- DRM VERSION 3.2.2.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect key_block
R/bbMphqCRqeZGgPcYJEgCasXIyTMrwEAmPzLDoE90K1tZCTxDGApsrVVXR/Hm3Ud8CQlARBkvuj
DYy9rxritG+auyaIYssuIIg7cg1dBAZLs6cjCCV77uXSXnrkuCmbIzvK6jGGsGXybi7JRFhaJqrX
W7HrQ2/VDMFoBamkVYI=

`protect encoding=(enctype="base64", line_length=76, bytes=827760)
`protect data_method="aes128-cbc"
`protect data_block
DSti9A7bEoZjd8is4CpJNbSRo7OkamG9W7hRMvDocs5tQupzj+zX/exa5yawFgh0Vj4RHq8r15UF
v7GJz1IGnXSBT7FF3Mb7yfNNxRUeDIwh3hXzS+eJUfzv0+zwH5kRwQmB0ClLUhCLjKM9cM+CMCH2
2FN4PDepS+hLXxgDOIMBr1JRZFM9HP/ErvrGQTHSZp/RIQukuHExQMkhNmE6SnFVyCShp6s/Q0s3
kimnoooS5KXPq56RG5e0EA+5YTEvWdPb4FMxMsxkv/AkuU2OZ93pEzbc1/B2Akkji4QijaPr25Qf
xRpnYTtL3XrxUOc0zFXocrEDzWoWOXSQQqHkWp9hEBUEegYbRQ+AKZg+uqL0Fq68vV7U8PbvrlbI
41+frI9AaYnHva80x909aApqY95iXszFwTLgqMLdg2dRHhwZgfO8Zcpu0r6r/HSeOnG3SRmwdHgq
lTo6FDzNUUe2razdwlJAe+Fgg7TMwpoVEU4Lomk0IItlhVSR2/j+cGP5MfINsamehFC0CGvVWI4y
Z/FlW40VDZR7oTDag2pVgjyg3T8JanZ0KRwPcOMyVaixHvv+EnWTFAB7uq+rzGMn0XirmId1KDmj
01WvAJW9pqySUBE8cmZd7zn3SIgOhHdquvAQRRsgtfdVgnH5MlTTXUe8EspbLm7hd26P7o6ulTgF
TOVxA2lHYKR1FcmtSV7mpzfx5TEpe4GOs+iOvxwf5olVLl2dYxr0sOgEa+GzMY+XOpjQnWPxZs5w
9ZBDqozqAWv02OgSVh8QGSOfJVkoigoGX4t6VKEoT0mxUf2aYHDe073vTzcNC3CnrHpaVhg0Qyy3
qBQFolFMX2McJTQBwg8IetBVBWOYIH5kxuZv7bWYxMDMa1lRQJVfMH8wsG3Eh6CJygm/ADN9A4zA
ROmG72lMTk/n9QWu7+YeLnkczlLwnk6p7q9VOZJ4fO41s+NHOOUUeciqKQwas2LTX086YhyO+wF3
WBstUC1qBIOghr+XQqyJdtY1fj+qLQb9T9TgvzVjZMwFK3MXC5uEL6uMQh6YTcxzqWdUWXYRbWsM
KbX8JjGgLE5lrI+1IBy8gDvP2dSDYrb02TCprs6ubFjgvqq9S+kBB+Yy8CMEDpq9aEqjRq9pftvT
nbKwPvXtqnnAQG5G1moNYOPjEueRpMQy9Cc6LAknECz6gO1fa3Dpjdn8IOoDsEMwQzvAgq2IBEeS
V3P3bcymADlm9EidEiBZuZiTbG+IujuPcP6jw9QVJq97MXRebpOu/XyO6kIXl0dcUpX5cxshwLzX
NwhUWu0uwFEhfq5HC1j3coghBgZWclkvfs1jJoCftonAfdjqkX7B4d+akWfIyC8/Jx+z7Cy1+eYT
TSLu2cNaG0kUSBvxzltt6Qi9CXWIbpooSr2JVItfNtYMzy6b476uANw4szZB/CagReZBLeC9ohTf
lE4Xmpalc/yzzb4+lm37yw9+gbSdlcBRnmoE5iTq+dKoOYm0MATCQzsE9zSVbM9lRo/mGPHa/HI2
IBqy4ErEv3pFuPgyixVm6wpqEBUUAI/Pl5NYhOIDhh9xOwGK770ok/HqB+PzC82OiegVBP9N8Zzt
8FGfrWqgSNkVfmq//WBp+uFOQyc33KKcA28vPUD1XcAGOc77ryz60DfAIERQsrZUGH8lRPgEH2/+
mIyp1XM03pMpniF0h8UlFpFwf3OdjwwiwZxnKIX1Dj+0Lo0vWUc5PJ4rGF7FNNotnGfDnaajw8HV
9hrFKsZSDx31JplxFdS0RsmhLJobulvmCioO/8x5bVVWoCcDC17EDx+HJ4Rx9Hk7GafpgMxrYth/
lTJkztp0oAuDPLboOnGBatjEPzk1q7XLfkcVOR35qO5qD/7RUNm0m8OcIGcaEgiFrxrCQ0XZ1X8y
3LeIXxTIgB63K3rtOkweN3dQZL/Qj7qs6RrhNJniZc8x7cEeKmkLOGS4j3q6Eu/7SPPnnznjNdDK
fodXslJ0usab2Uxc9vqaiHcYgp3/XMKHnBMsCyo3mtEYBnR70a2eEl8QDH77byLluvr7yHm1oKui
NjDX7yvK3ebHSbwsDMHgBsi18LGW8Ft8KW5aWAjQDhFjrSx9E+N+dGVy8UtUl86cPCw1UCDuXA1o
xeCF0zhD73zRQbwG8Mmfevp6z5TcNnKWPPYgqMUmUQATN/ANN9qLRkAArOmyaxmlPV1O6TEYDnbq
APk5mMr+qpsNpQX5vWxLcmceyjncM+2DBvvzyoX6S11HRxyneATW1S5Yu/TesPs9RWGSBKyywfQP
3iDlOIC570Sb8pGASomxvhF3lSrla7AJEd/KIn5JmJwvL5Nb/zX8RKcY3Kz6reyx2gwymk3NOapz
+YjqdlCPkA0ufzzOKZiPc4zKphKKSnJda+/HjGE4NEAs0c+uHCoP/GXTrwLXppnYL4lhyhAE1uhI
x/Vsdd4IRun7AkC0R4x8brlZunn+MkaWPIC2TpUOhYuL+1kJSHHuSSUV63WL0pQ6QADCO0kpJRCg
Q0Ek9AkHbX2tKp9jrvQHUvBNVULl6xaIj9eqH3foV3SL/0xMexbPpCeEdV3evJFAPk5moLD9AFum
zG60MxRoi+p03erCb4kq17mgnvU15RSioslTYZpZ+Vh/iCUiSsGKd9KNg9waI/DHct29l+A/kVdN
CByeSp1gUcZRVBSkibwixe3ehLnJu653do2DtEH6L8Sz9KvA/O4tCDPeTwv3k7Q2Xx5o2EU60k1U
SobdTaOa3cyTp0MBSU7X/65zKjwulSPzFWY9744nYd0Fju2MlZ9ypTpRvKNfCG3vUzB0Fos/DtxC
2foKlnKe4WDYOck8CfareJ/qU4zsWUntaHz1atV7pj9/sjB3HCF2lM611i6ZBnboXwDB8SWx81nT
Gx9W2HI7wfIZ0AFT5qcw3s2QnsILcYcDnuiWfetdQei+jrgkZNmBFnenntCvxT30zRKR2ouRcSSK
sVmGQP/lncPKnx56sWeaGNjPk76peKCEhBDoG8VOHIuLu2u7AzstTsNRBvHiiIC7q7McJECzbIc5
9CsQ9lEtnbmUXwfRb2++1ToYwiv4xzYlxntCxj89b0DKd1mDUooLEiKjhUOqD3iQgbP/aMvsdin0
mjNBjAGPP7mrtxGMMgjn8KccrNv61neVqs28Iy4a6l6rcWvATDSryUMrsHsG5iA5oITKhMYhI0Jy
y5jTI5TuSHKf9ICv6EoLdqSsFrju5bIzb21fOb+7NwaEKZfqINeKuU1D+AB5qCu+DwYm0pafmEf1
7QMjhfzqYhYFaUxwmv/xD58m7g73DKkiQtpIkj7iDOA9d1/uWc5ukS01mE8d6fh731Yq7n6yofsn
n3HWdtUg4owrKX9ItyyDx0uSfOCGCJyD6CyM8absWlxJzrT2rYt5pwOBw5fh2Hl50nfch+CMbzVr
MwuAzCecGuBuwCQl3sXdfMJyugEJdfE6uh0LA8fEI5jeFpyV91hugYna9tFCZdFPAKdhFchlR90n
tXDj1hvWq5fEWY8moblyNh+hSqUPvenXezfluJtdXE78hwZpVJy7pCkul1hDI4fX0Tz076IZxVT8
i3pkvPSfFYYplZHycf9J+v+hr22i2VWCy01Rv28aoZvBHMTN2CGWHUvLGa8Yy2VM8YWOpiMRQjTo
hF0cWx5jzkIdbKxJ0BQrfTCi/1WaN/0rEGxbM/VuLALE96DsMLh5RRohaZk+SSu6TzTGGJxzOczb
u0jXf2bEr2ggqvozUJrCqmTnR+Y0UFUr+kJ3Shx4D1J1Sqss8XP34T/Vgg4xzvbyKjbfMLqZfDtA
AkYCmcQCV36kFJYqG7V8N3JbjV76QXAonqe/d5ZVoiUlFMlREUuvk2QwvehPKeHKXC3hzahBHZx9
u0tX3utAEKqdk9s8kq04MqG2p8xra4vmclfxAKVx3UU8RDmR+6OiNfWhXM5kLp1aiPmcTyyMDVWL
PeY/8pygf0bwNpjnNUu0441FZfbC9c0fPm+A//bUUZcHlwCDO8OMgoa7qZwVNOHbisQyJ/J3dxEw
NOdrtWgA9C2sOqNSiH2tKxm1F0fqizQMpxRrsgIChxb17tPkKyDV4yZChK9c/bHOSK6Z4J4C0BTf
4dBbYZldQX35RuYYC3axU94/EX4Lp/Ic3bBwsMjNVrzXU5tMjsD7AUU6+41upWYbzddTd/YrrjbX
XkE3Hh/mea4RI/6eJCI14gGqGknHghq2NY1W8Hgmi46hZwgrFaAjHMiR16QL1isWxvMDb5BORCVC
OxnQ3+OfBw3WErNAwbM1eT40NBBL92HGjF47shqel9R8UC4lByA3/xEsaycyczvvN+i2vy9jQB+o
9owVEymOL27CFlp2jXr7tHJcWjTVdGD5swPt23kzpYtMmkCJTPlv5vgjh1L442F0A8JoDwtNuDb+
DnkTk7a22Gq1mS/xJJ2leXunyJM4OAGwUwepDdK6moFKx9toZ03A/gglFhhickmvNNQP8wRgFv9a
jghKfBts6C/28JSlVS39kzt+9deRy9wsP6hUtUyt9QFe9RTDiu9FrhHAfoiTGY2KZ7Hpc3FCr2rR
puJ1aWI4hP4lNXmygbRv7IOVQLT35+mmTB9+AIxxx9CrodYybQzocbeK1ADI1Nlc14znosY0rb5I
u7ohnzHuifdDlEv89ercf7lWvn1HtIkZoV4+zCrA9Vrvo2SEZVt37ig3TuN6kMTkBkF4vCuLXBMj
3ztwwZbvTjKT7FXgXxI85yfMqO9XuyH2GJIR/6g231GB1uyvlm6sO2J3dM/RMURFkFKkJixuJtOz
ezXg/uVvjc+ccUCQo6Wnfc5FkDYtazRoTipHcS3jcWJ+fqrmHPiPZVK3DB4FoWtB6W5FykPz4Lm7
ckq/o9+FYlktCNnFbhUiVOTlRRu6n6/R3SG3m6R/xX5qU3hZ9rZnwR9OXk9YNy5zGpNBfNo2+bwB
pPP25pvgkfDLEB8Uh37iaEEI4faDVIWibmdSsFG1vBiLfXyitvZgkIBKvmKzi9wTLiL4mB+qy+pq
ekCrVuZ/0gE0X/zw7BKaJ9cg60MHzGVNbK09Mi8IWZjXykHDzFvewMraeXdQe6IIaWOfGPsVvIhQ
9FDAOBMlT5ZeXh9DG5zqggVCzm6OKUcDM0rEe3togudaT3nJ6ShKqyLFzwHK3b7F0FA8tkjoY9k0
WAZOGtPkkrabbjgZrWKk2HEXrk7PL9TugHo4PeywY8XdK29xiXQXwoRtWyO1Iuxdi1RPvDl9c2ZC
SV6H/fn+MDAv5CCHUV4LvLXpSrbTM173lsqvhZkUur4XymjwCe8SrnVhjhQ0LiW0pVmIdkJcLXEg
OL+TBzN2RLsDpkrBq242I8dwqvlfiIqLnIjI9JNpFxqS2EkX9zPiYDTRDoNElWObHMgnrGclXgtL
Hk0XPHoQmBNKKfftaNCmYzh4jPdnkj/Orj+YrLlLpZuRhL3hYFtjFcr3W2/u9F/hzY0bMVpJx621
e2t/KNMk+fduolesz/uSqVfpVGUXe1SZMa+gST8h8RDTzrt0vmQOVqe2MMU4DNLCGYEWkkb9qwUe
4KBkLIUKkubIGexyJFMc6L6CJqi2guoLWRfD9GrEmwJ0gY9vpBExNhEcDT+O7BruHtWYbGx71dV8
G2NnwIgo5lnJN/HWlBTSMQsd2XJ/SEw2G6X2Yqi7ptZnLdhNQrYOrjAW0SzyqcF1QE+lne11/LBU
ihiUHnM9i/uhAUh5BtNitE1nPNI+nJRKA2rBKT5I3iZCXiRE4QYWbCcNv53Pj+9sZ6NTqg8P8/mY
wAJgVazDyigax/W1t7F8Sto+O/E3XnO6ZNV0pQF0lMDOq3JLMEsvwx7kiQ8/E3QgVORYypuSP2VH
s/G1Yvc8IqIjpoBSQF2S96VnjR6T3Q2ok5r1OaydrL83wswUoEwYV3WAj5dyB1g8rLREmsP4dKbI
xHTzH0JinBUIsBGPkZ8q+mMf30K4f23dKX66oqWTWKul4TN7Xvp/UrV8FWmKFCtmanEfsUyANzpI
0h+iCNPy2K/0gMOKEfwOAVYckv3G0JGvFzVDEi4rJ1iKn6P+N6o0DJ6WFZ5r6iwP4cqsJ4kZyOF3
78Bl2TDq59odKcA2VtbQZ55jUwvSSvKmCvLaYj7raj+LoZdaHutk67mrJZuPSG1uwHBcCV8IcIwO
EP6QSwFz8OoQNpiMnqOyhDCj/VZKQj0o8qWGR94UOso66g3vQOEp3B7aS3EfGyPg3HMjYV3lqZDP
+08hkwwUnCad2rjldcIYO0Ts1UnPMJzgCbgccVYrf97eglEUt0Q9DaOeXqDOwNAXGDJTSSdeGAeX
FWbu1U5SUwpmIs4JF3R2GmbydHbcekkvbA3wKMlTpPnt1uWunq8dVgmqHLTWy7CK/wWA337FszqG
+eW68n1D1P0mHPskIrfIxXRk86sJTs3Dph7sq9367snuZaEUOtTU9gXPj+F2pmorfdKSnPz1clsd
SDyBAK6W19Usu+hapsWIlpog2Q75XEdHwEFtPMtJoP0x6I2/TyPnSj2Sk54oKgmiV4YxouunXeq7
r31qWjjNMCmKeQkIeB6qxuMTwhKPc+l/Xm6DOswkG0hJOMitaSR3T1JAcq+7rXwh4DmRLa7/g9QN
LZzdewd/9aFSGRzGlx/YOUyLH8awYFTXn8/IYF+5PM1s+3Ihi9YXO0MrDqZ9960vsQtR/PfaIm9e
yWBDVvYxHhtG1b7CIY4i3Y2lKHjX4rN2Jqc7SFWKZ3b5zsgJ+GiD9cVwOgXz2dI/Q9Zl8oscGBBq
BIu7g+m/nhjUCEbe+qizUG6I++CR7wKuGmaYXIf7AF9sblLbuIJf/jR/7HVYqTz2ZDDLWkv29QOQ
tx+PgN+v2VwGp6BT8DnjS30OwF9q3LLKsw4VSyTvzhymTB+NhzMJBmqC8G0I1n6lAAoRxLZWNGXu
MGKrXNWyUapNTTg5uNquglyYKvkOlyeVrxTXC/+VAbtjsM2qO1d+II7DdNC+JA55VhI4/DHzhQFD
tsxOeEvKKgUb56Ch4N2N7hsvZXN9u7tpbvsncykacyGDLMVeabN65kQZ6rKBVtz1gXW5yg83nH1L
ttWFVdveVawTAQ2NcEq5oVbVDQOvbWIcIxyU10mn4iUkDlQFCLTlDKzWxjcAObFTVKg9Xr+++DSU
x+qDwCNXm0j8t/wtJxrTTw98TuZt2fFlBYh3RoMd2T4vIvy5hX6Dtdmg/1ZWTH7R5z4XIXm41kbH
HR+mJsAbmIK8Z5K5cdn6eNSU7Ysp9pEe/FOS3vOr+5h6p2Iqo0XWJKPJksVJphiDeeh4zOD11MNf
WlGCkSeFqUfYJVlAtaH/t+LWVi7QxQjZ56f7uRE8fwdxxRzwGM+cryyuCgVJp7PU59umeUcubVWB
p8/UrCvpazfk3TNwMOiN7SpY0JQUkfEE/50Uz3fxD8Wp51QRPk+AiPZUnEiUZKUfK9wYx2jgNB7O
shRwhP8qNL3K94sIoNPF9A2emKB1Cte8dKv2Bu8a8Usw2wsT2/CSbNzqo4PoudCIc6PK1NHFDh0p
9BNZ7jVsrttm12oO78OlnJ2V8kvJV0is65R+TM3uUCdr6n7k/LLgaVSeT8ZAVjGLc53V/O5F67uL
x9Txly8CsRiH5Y7gfTLWM2nkXf2LjZScWKuWlKVhmkqR8dRCstyZ3ina+9X2MdSwNnqsMnz72lxn
gvQUVk3E92Hd+9UfbUSDfwRF/Qj1rjDqDdcp3ZDuWyhEa0ngdkZyvaFTOYmgny6IT2E1f+pkEpb6
R1ZX4//sOaQPZHY90x1AXjFVeXyequWvlNgwODU/P/RUseWndOwQKrq5bvQwQHwj8gX35v9DtlB3
J26ePM5sfXTECwo5yFTTH1X0ob+JWyX5YcxbAPt0W4xSJpqWBmKSpC1iy8reNGH17URAt4tz3CH/
EF0O0CUamomqgwqqexz0oz5qbQIchMK/oLiINZAIm4PGU6bJt1jgl3FYqTL2RfBHw/r73ZMNZ5iQ
+sFzipg308hCp3/Pmm54FkgllBc8YqLJfCa5QR14B+I9fRRLxZUVylxFgutwDLHgiPqmib5J82zI
Uq5c7QSLaIryKIODcNhIxvb1Cg1vKzkMw1jxUt8GsDVmR8J1Uukpa+nGbp5cYJPqaM8PFY0tbaC/
qV077Dsl36Rv6/Fc0U8BssulHcKW5Lf9NKomCkjYJRco72Spj2YtqdTWHbv2mn66uKk4P4BZTGpB
TGKyY0LioJS/Q4br5KVw+Az6pWiTQcDSImHMUUtyW/CN/WtbW4l8gj6aLL60dBRTWoVsCTylmpO8
aitDx/STbQUQ+HCmngGYsEkR2MRUtUxpbmRhMo0obqU18sh36fCKIRLShquaqpPWw8E9kA4n0NFR
ktdnUafTIFBjxuL10uOTBVQE5pLAEWyN1ydCaYNp0lkBQuZGYZu4xoGxqDt8QuLY8Qc1/45LbhmS
2xC43yfiB4Uvml6/IwnidnUk9jcaoarX/aewSb8BrykOsvLOywkKlHBwLRSW8X25EwPNrCqR13df
WygJyLpxMRP3lXyCahfQXpGCfvP2er9RHgsWodlqPsDQRGCSDfQBhlpReIN248uYgqiEjijEHHXQ
Fbt6dEF8D2qUbCSxiulscOmHmxeYKKMV08x6vHbj/KDASNOsgR6TfAHlSnRf54Yw4XHhR/qnUCwl
N5O7fRm6iq7DioymPDzHdkvF53EJNl00oZn+1OjRwMRf+mu0Bp3E6Vbs+PyhB5PlB4cP2yylIOsI
mmvZIqk8TBM0BHDKgshIIQ759EbYeZpsY2xu+49OL+JBVo/MP5oXRFUWKIhQ4InaM7JXt8qd9vj8
E9jkvEMXZyhSjZE4g5IoLPJWne4M9e6wYCRXUWj4/ROUBNm8Uj2z7Kt0wQ5fNU+1krgcy2+OOFVP
9hLMuNJKG5hw7YkKwHMHqI4cyBBJSmVV+KeGKOTdgTrODSER8NLEy04+tVQQ4S61fSiy8q93jQJz
MHvciDj7k8vNCcQQ1HoqulfHQVBnnciq97KJ52jKsJ+A1k6lZ3O0JtRxk6AoXmRsnU+P0hOEfwxc
cZOgvk8nYt/HMj90RxdsbV452Cw5pUKXCgfUdO8JQLmred+FoMomyaJ6YUZXxgG4JrJTblM7RuQl
HzjUeynjK9oA5JmRD/g83MnD1sEbxdeTnRo7qXoLTHG18p5vYDhmi+F+RoZkznEWTtbTu5z4piX6
suLeks78bZmdF0/f+jrZ54n9UAmkoteHwCCjPoSDaaqA7XrsBJxRIlzlUeGlt+K+9tlN87/dYzpY
U2QJpVa8EBPhEb/BS/ELZxdD1rx0K6WjxVTC3Qz2ftzf5qxIpZr4WK1ggRhkNtAyr/VN/UdMl2/1
E4JM2e+pFE3INE2diO3/+/qk5PYcyYkTBygSo86lsny/4uER2r4d1GTUZuUHnu1V8maxDzUhj8sO
fKYqnIjG1rNvDzRBE+gD69McPufTzDQ5GXtcPOrlBe/u6tEOqgb/VANxJFxLATOF1uw0RN0oMcOJ
MLHXp2VVzROriQ0OT/S+9CLJnU4xdRtQ1P3FOfLwNebpnDIRlV37h5zynTRellA4MNkaVfdjkLT/
vEfjGwnXbLCi1n1rKFzGwRyWmSLyVW+bGFxCoDUek4Lg1d6K7obTjnxKrEDKmu6n4W8tTxpF7kgi
cxG5fGs7//HQG2Ziby1vX3umwE0mRn5Kx4vnFj6vfcL6UM3dPc3Lh8BtkbX1q8YOvGUZ4Pp55Ju6
uW9W+4L71WUuz9Y+iWQf2tz8CG+HYs/CwhZxGFobh9g6eh0i4mB/U+xwC2fCQmPoYCaBZeGyT2hy
/CUQGMdIkk5r2Qp1bd9+XCwq6dhxYWJ78eKKR4Xii34TZuIEKYCad9FZjBwogadMgh0V+FrepIaG
53MZTqEriqI/cWT2z0IPHyMhbY2w3Vue3uC6x3LIEuXhHirTGpfwN9uAQq8QYfjbu5th6e7DR3fg
AHtJpgz+RbqVGvgg85Y9ZUGyYPSnxr3JjEGyr/f+Zf7YKnDD2OOqd7ms7mNZ41z7rstjxRjdasUS
rKfJtZqhIaolqVAx4W3fadzYjCvTrPVZssS167+avTxy1/+K0papXBqYbb9uvQD8xOITh81zFozA
X4htYkIZPp+raye0GGuYA1gLNddO3M+eLjIeHFeF6oXNSyI/vIEZ8IBKkPCtd9tM9uFuUEtrwoAO
71XTxgpqbM4NcMRoph5iZuWPVqMLvpViSM+eY2ckrhLTJfeP1yAcfCTdlfZlsSUaDr/D7csg5k0s
LrQ2gbNaaAZFZ8vQBlqJ1GD8+196XuEHrBBCt4gOZJ4vs3mCO3tHeJ2QH0SWb+S715aRWNOT9TVr
admsoXfB6WTSeUw+WyqXbSCjNgddhEu3Do4QtYh+xTAw1wd2rrAzTIIhdvjGZjlf65/wdhipjaAB
xmwF+bCt9bWp+DRLfQCQCrn7RBtj1nZPbOpktjgPeVjjlFdNcTtNxGB7506LXeB8swoajL7ss3p9
XLpZbq3TrGSZIvOhHg8/0DDMk0lO2ySjYfui5xJuS26K4eponRYev47GcNNvoJv+SmsI19ueWjOZ
3JbiTkeyU8AX5q3sIcM00OsIqdkda75S1TackFMge3vadUfpt2HuxMjK9Nb5oEGxGK0+to7sxY/p
P51XNEIo12qPMHcaj/PDlQA6HOX++kXMpGCXh7Zm44jeKlrm7FlYdA91HPWoGtAAVNFNyjU3DzRk
gEoy0FHNq24PSvh1xEjJadyj8+WkvUrSou70Fu9Pz/xHzICyROXP4rPX5qqcl1xIq/7eHR7zxTk1
UNHd5nCNx9LahLanb13kAtU5gQeyzsJE38oYb0YrXyMeBshL2h7wSZb8NaN32hYBpuQaQzcdXAl2
g6gykuXSXsoN0U/GSVwzBuwziaE2eYQlaEcZqlFdxEY0orjEwflDtIHDjFzSy/wE6R+P4/uSMmB0
KmHCc/0VkNwNRrkGWhnNkvUQY6Ylw1WkT79c1l9pZQnIgsT3EQbHJNrXu4hWcljR6AXhAuCifDS2
P1GIe/+EprsNi1C9vuDVZDoDwLoVS4uwih89vRetD1FBzNkuSrqqmbRohgvmb/Go2kLLFjlZH+tO
OcprqGo4WAc1xPEz/9nUKKI2CoZLP+LbvoVA+TfcPGveD7TI4KPy2nVxUju/iPjtoYKcUn5Wih+4
BSqWKhOoHs4araXAnou4QwWLFeRUr4NU1humTD3KXzMHol5LLYCuImiEbTnBL3zLRuGktqBNQ5ki
sfOGLbAPAaVEJmE0uf4wnopZiktKaH1ZXTjRTYxJdgsXPiIYyW1FqA73b2Z4iSyrBO7i4rD/N53g
mofd7tfh1NdYQlt47RCeyvmxpcdD1NW8seUATgNQ/3vLwPV2FolL8UuLavNm+RuzINd5Q+AtHfdi
dpESu+l0mrO2lKf+zk2UTV7Ts+HPyecIi2QPeqf28dlRpb6XhM9ZaqUxEqf+JwLL61MNAIciyv3+
LEz2lDGe+sCdrh4eb2un5J8djdso8zm0Do+pNncehd8WNJ/zCDUjvI+zkQWjDOIpYVuMaOuD3Hm0
hRoTpTs/jlUj704BCK405dnQTEwPVuxY7RbNBt0ceFeIykeeqw/a/n11MixwddanLAaznS0az/DN
Sh2jOasKe/72KQ+OTXXvKgrnEm1Ie0fDVkg/9Ddp60dOSO5EnjDHebPubsiP9ccErdK0bWGDdhXG
/y5QYCVE3D6TzP2AFjtLyCdWymkpETisVmL/Y+9057HWRl82nD7BNFGcLLQk2rRBhWiLYQ0aihPP
wbLJZY3oRqbE2eHy9EwaEM09R5zB4uB5MjtSphoqISK3p3KeArHirZIvobW6jouR1TRpRyWZNXt1
Bt//k/tssn6PDuNt7cUgmJaGKOcvSBEIBFWkD05OmKzhDSQ82WoDyAFmvmq/aOlCvhjwBXTFTAgW
AMVhUSkRwNgFW3EU+693Z678CE3PJpk1ZzgNiJMX4p0snilgUyxxMXTSA36u0PpzZ2p5RzMSPxza
XyYhcTHJn+x9uQURcKsILjUAMZZGQODkMaoedDht9NfP4nEqBFFcTQXEqF51kZzqrnFUJZ4xeyvU
3jEdrrAHJeWLZFZio7N49SdxSVntMofHlwwByq2y5XGA4nJSWUEaSgWiUcvRojQYXLrzpxNBTtZu
M6iqWPYErDZXC5DBthAQFQCLJgzoEbOW7UkMeDjgFU6fRm52Gr2SF0/TdBELiDZJkvwuzW8473xh
JcN6FXbq8cu0XYyxAI1uaBVfpI3JtVHiclv2Q80mhlBLzqn1/MxEl82SALbU8nrwOlqShYh7zgW/
1ltrC1/r+opjDJ8G2TE6TPWqHglIgBu9N1b0XrJi/yuoR9E+RcgPBM7IFxwCE5Egr0rg/fZp5CsB
LWCQSp5pD+meai+nEnbeVHysomefWs2my2XMValu+yqQVS0jlN81grzGEO5rVNFXRRSTUY6RJVue
jt1jpNvjug5ktxjrZjFHRMakTFirxj1Hd9dhvX739/gJi/8kPeBjwWm+2G6kbypRQ1ohdNR8Qz2G
iEIvuzlOE4oKx7tiJ3ihpGToB5+D94Tf8jOS03UrOZ3XBhLXRFEZSjLmPjkvgwz1PztpZEeV/Yp1
x9d7r7IRKRKWE2uCEED/kxqBgt+fhBREqYctlKc5e0HUNnVl+aVaoXzId/Nw2NLxxSe4qk5pMLgv
b+zV9hlFfbFJgNgn5YUBaicl1nxayWdylcFrFtQNEozL/GcvX+/o1jVXDvfRP8ODHA4TKsNW0T9I
iZNBip20BEXXrAUP90dgtuKlyRPzWT67GhZ2WwFinmG98SIdJwDDg41ZDkovxwU2nIVZrrM6WyqA
cYSVVibXrs9gOZtBGjr72uLoKVxW5xeT8Rm3p4IaqngiaHmgW1KgnqiWKvLnqKa6KI4516Tt8U5b
8EFKD2UPJIi0gSw4l9HESIL1s3fCJVfrAwLllTKV9ZDupYbgRK/MrSQ/5PJ18rjjl+kWyoRIQb8d
6ato9zxRNqML5k2LuRYussaPoYRPPGw8DwqOQF/5AY09NR9xKxb7rEqkesDQ5Y3wd1Dw1/fglIf/
wnJztdncIDe3lFWtGXNgFRTs/lbkJCWe6vIVQoiW8NM7exhw2hFWfNYgJ0OGxY8kbwYYNNNOjhJs
eaYEkJJfPXL9hldx0XpH8plkn/SW4/ZfhF0/hh+bj7gkJ2BBhPcY1EDCtfGpsQHYPqE0+ogs7o+0
90shRA4c3u0GfNmSnMWo/TA8j3hf0IsrAs/qDYXr04IteI+HSFrnm9yoXfrV2TJiiqmDjBWcZFIU
Xy3v+eb8l6KPjW6nSTduNl9dsIwh0hwxLVYB01RANfiGCyXA6pZ92HogrOXNHBJnB3fg6HWwwXLL
WF8hlQYGxK8iNt4ons5Ttt9IRBN+18MHCCqcB4sbEXkrg3x5G0/CDcrINYQk8hCe9P3c8UfAKhXi
aJjEc/zfX0g5fRY+nBrRWbbNwBRdHPBXG+ZU9ABr5SZrMd6SDVWU3ZG9KwYg48D+nebrZLvCgUWw
DU7KrLRljSYpHCcrrsrhuA/RiHqb8//gpRW86HJanQrsJrjHcZY3/vMDRUs+Fgta5HNjL4DN344P
/hcaTsdJPndi0V/Z9bGbFJANIZWFuvJoq9Td87ts7UnzCDm5UXZRT8Tk7AtINBB0vZSkFoGKUujS
lrPFZ3zcNy8bIdsUJGz44hLtR0Ovz16Z6aey03HaeMrOCj47Vx/t/DyJqdN5p3DRq6DqF8G2S/MF
3AMzO0acU/o151w96jne6R6b8/9KSlenLD1SfG2+PNmqQ1DS1hILlfa+xcBm+0fmMlc/GSOpZO/F
S1GDGCUsFkcPCdp69gnjvMhi656fZuPOBqMBlbQSwWTLxG7sFNFQq1+w2SIP/pRXnFoLVm3wjRxX
XlpuliZHfIO1Z20rXGeVgOBGECUhPEtE5uYInMkFZFDXiED86SKS5GlqoO/23VAPHc8JKW15GZ2B
qCTVFi3dd5gJ72OP7fKLKC51TUUZh0JKK74BlWQITO5b5rYHMrNMJONg809RDHy+lXcPKWtZhQTw
c1cCTXKwyPKzUoSCzfawpj7dZmfeH0bJFXPRXjb5DPI87TT2SX/ecsKj0wH/YGezkGl70zcR7yrt
znSi/R/qkXA0SqrHQlXV4tXoo46lhhYsJMct6AakYoK5uz0NLja+lboACr4wec2KaRYrmnqzuAdU
YOewCB7zX7QfdzTiPOfw13CmvjpOtZS8SU/M43AUz2eCUWV86QwcWQNavGDUrbHMWynU/GJjhyDu
vszD+2jmYvABuW5yjPB0sMy2fmLu4ryTmoHJJSuTHcOHqfD8/tpVwnZirwHMuu1lwI6SOPBa7aoG
WQs2yseLqpL4T/k09k0zLGCMf8RpMudBIrJctl6Dxztouh9RFuG/EdvtINa2agIB0QTvAcnfIiZM
sQAJubCYoOZutF32w95eD/J0UxRi0aEPXMqUpMhgrZ9+Wpr4kZsSPzIiEZKdPFxVm16x9q/dYcVf
s2UN1cV9i190uqdhXJFy4qBrj89w9ZMdJQSlcqmynrUFwLXcfLciAZi0WMr+P6GNVZD5MdSS6fFJ
TMDf9hxXq+ol9/vqog5wUKq19XWulj/AOkKqnaEPErCHmam7rJ5EbuoS6QgVvoGkMz1VCs1oxNN+
AsciehZ2Demq3U1JiM3ptw7eWsY7zr7Gn5aZZ3Qb25c6p8veF774rpCe1/xjLzJJewu49wUIwNmB
UxcbUtjdNMWeJrYUpS2dHSfiz4fB1yHtUN47/lNB2rwGFO/TWSiP9FViDVApHizgD5W2gGUV8mRd
t/gMPPMW8UUnGNGlG1cVChKiSAQx5IOZbZ1XS1JDua7Kmo15LasmlxYCvGI2Rr6Fzml7qRV5MPDj
W8XoCIOzq1UKIe2VfdwQiCHSZclTETrK1JHQBdcjYOGmMF5ZB/NUWKnSdzG6aJOvonm1dR/GVrzd
L6DH0+hzM1wsyLYN8Ey1UUySBNfnVSfFQxmW5QdcZ26fdK0ejBjZfn60L4VZHOV2f6kS7Mluc0pk
T4QF5o7qjJLv8Wnb+erFws/hNjoEUyEyU55V/GXSi9T/eDRGa0KLIio1wq3CICQ+su+wbfiFr6kS
s8RipLOmKUTGFArpp5V5FuDBOs/UP/pWilNMopSASqziaxjrwgLTrgSp60E3mZfJgP5/gGH2e6mk
QwixQ78uPL4gwYUzMq6kbv2TCMho2cMb02ZOyEElamCn0/bLcj5fBRqleC06zRM0oylJImXQ6SZr
v8XkMMNghSKPKGd9qMoGXwDay4ErNqD9otjXXAFculwwkF3pVkXC0fqz9pRmE592n90NcpUslSBi
VxeBuV0dVv2aFj0TVi+oqbObDm7f3tzG0V4YzzfP6yxZVrkyTkcHoyM4vXV3dp/XmmuaOxLj1lfH
Gngo6FDZrmNY5qUprSb3h83IEeRsHibnUUA/Jl86Li7/Wn8pNS9cAatNcPlSQvYrYoyfgPZHYgeM
Z4AWwHAFZr2TtLD97JviwAredOaDCUJb6BA25VdO0NbiEqLjHXTvV+6YW2TZpsJ4lHZxz/oqrmJt
HP+A3RIq2iT7oPP30v3gbRcvamRf5cc/HHOb4/jgQFhdp3Rv+k6MIQxqoMdoFVdWg92oEEKQ20mu
aWkh0F8OghJpI3WBNvwxBoqcqaNQAt6oKSZXVz1as9mp3PySQpqnJTQIEtPQkveesZb4+q8BitLm
5guk9aDnOgduXoxLMZ1mK0ginueATtCuWL6jszh3sLG+KLYJX6JhIrf4ywGkQ/7xvTz9MTna5Wge
PchZcqfJmzcrNHU3pz4ezYUmvKsdvf6GGFDTzq6e5ZENJwCnaUIMWrNgHeJ/UTMb2E76JIXlZ9b3
+x6k4wIqlhBs4cqCsGdKY0W5opST8uGeF0B8Il/NskiB9dtCbgMagBWy2nIMv+oiURotgVqxM1+s
0DlE2YSYhOesk/EqERH3vBEhzR7zDLtyxG4oqfRwm6i6PH8otZIgUzB6X7u5QlJA/0KUl0IAy/U3
VInRAEVDbL8p7KiAAcD3sHEb+RRhrKJ15kXZJrb1QH2Pm8hNN7UGj1P9g7aXsVQnxmLyQtV8iNpm
RHMU6kluZ+VMZKjNbnCdiewDehVTvzrWKOORCGkdt9jWJPbAqThY5fKCrp8MI3SwkV11IGKT/QZ/
BYY2SphoP3LeT2f/aGYbO2uXKLQauKiYKQeJxGUSb0E/8wgYllQC39TeyMUgkJnyl55SlenixF6d
OxDkbpkfZlqbbNsFltMsnSq1XQHcX/Okv5rE+AheK2gCngxb21L9yFB9JA3fHbM89mueg+TWYf9/
k17eq0J7gGtmP20HwOncQkRTAHB3e3E8fk1RUP24FqgVQ72SjTImH8sYM6hQZN5CKhywSIOl5lx0
cuajvy8UxZ5+8916c34uus8/LCfqSyMS0bbJDli4ebK22hBfNifaLNdzA02uv+pz2L1IeHIHa88I
Wpy0kQNfElqUHNjmrcitnksMf8Q/ldUtRoQftN+wERyif5lg2pZwAC07baq4pUPogACy5Wz/W/zL
ngmKdlyaWIX6dRT/n/qKPpyZ5DRzJfPSe/pGYiPi2HZrgEgdKD/nLViUfHQEqZ65/eghD6YJl/M4
W1LQJ6uydAz722zfy28sJ0Ap0ZWNNfwmFiGS5AcJZYtucgZQwJlyfob7JtsgvqHuUj7stIqZfOXv
vWp16mvFg+8SLWgI0AOh73m9BkyDfQOjBTKK+JTRcwO/tuP8C9YWNsQjiDK/yJqqVTl/7X8igZg8
N5igqzn3FtWbu+5qWGqibDR5wy3j+m8mtz99lhs7okZwJN38PLaoS74CXwhdX2hHqT6OtFzP2tdJ
80wL6xjx8innKFhuqt2TnG0Y7LZ33+Rbca8IBvPOIb67UL83yRgplxG7vyaVwT+SEONrX6hQlOCw
qIkwW8Ck25EHRg78nHT+3Kd2ompkNF5xexfBYgf76UpwXydcbLigA2R2wBtV7stgbPRGFSyxdhDA
kRR+t6jkDLZk82/MFNmEvKi8VwI8/bl+0rDcIvmLWDj6SQujhRGbG8agptbAt+DS8bKmln/ZcVbN
rVmiMnybv6+7U6/wwrWErs/9omBG9sOKEzMLoyoJ9J7R+sbVj2KKLtCkSBqiGKdpTW0TrbSkgHw6
zX480s2NNygPwXd3ldnFTOg2Z9MfUl3qQi0TJYz1wZcItTnD/kw+LA9d3XabaEvULzKOT+EdN186
k1Wq3Kq729NQ1I1VyNeniOKOUyDGF1OhY2KjB1plzUULB7/8xlNAORTUBN/L9/Eob6VIn/OxVTno
7Ut5CBV62O1SLGu5cxT4jEY85oCjV1wWWSa0/pjwy9ED86wSxG9kpw1NwDdoK5hKsrAbNfsBgDPk
WFhSNvAfRqUs89k1gfirw2fWm9PmR30mS68o5z7Iq3zDsHl/LeVHF7Z0uL47MGJKzrFVLmTfqCRf
Jak/wUJRXdkGiYeOuTqckqzg49srwhDKoA5rYKtep6d5Nv+A/VITMH7V6MAsMY/uDMjuhxEfjX7/
8bKfM4ROjuNirozHW4Ia5dbm4ifH3L3dvETxKHS3fIIJ5kAur4wSM5N7Eq3BVw2fUOfOZQEkt71r
R1IQYiYdjmi8PXrwtkT+yP6uQJzdjbj1J7ATZpNQQb/TFpwrDihFJVjh7IaSnKj7s0CMzHgnEK8S
R8tVn6wRbyh5s+OKEWsuMj3LYYt65F4M+fIRtJUWQ8xIJquhDOf3ZsqabNn5nv99GVRYMNUYEQ/2
vg8Nfuz8MtBkFctS6/yog/gkfoQa/qSixAiGQqy49IQDYP4hHDXLG9r7F7IednEXOvHYRMOJTyG6
g80CdQe3mIaGs43Al57HeaBHKyrqJrR/9ddTYTvYdD/Hl6kdRnxj9IIEbgRtdt7isml6r72A8ITp
rDHCA1VyPeJVBCA+dQT3f4VB5YZxiNHUp4+Gah1KO1EBJ2c5/6xVhT6kJiwjwHDuGmTMONX0mXOM
FXXsiWIyb7QI7ZADgOKMNYwoVlmTg9hGpQQ/Y7cVZFofNAXj2OIlBeqGFMQfMayobzE/6Rqr4yDo
NFzZvQfd0zwmyX5TuXUXGBpoJUHUAADaXQoq6cedeuvBO3DSdozKoEj7i+jYi+qM08GC3lZWflvS
3bYxjMry8z5uiyuW0VQnYmemzFJzZ75VVEn22ZvYa5zGOSYb1YaCu0ZGOeq1pzbi91C5dpgbmqZZ
UuQJCzX2g5wJcaS5pUgldlZPN9XwdmSt+iLzXbBI3yJioAuFoIqVVYyehy6i81/iMmxW3pu7rd9M
zjXX7JHAQnZ16nu9Js5dQkMc7u4aeyvJqeqcIvAXPTHNO1XU7QCguKlHkpE7tVQSNoncVazXJ72e
SODh0gU6Bs3Qt86oxYxGNDbXPDSJuSaRZyJ8my2RY97TygERzvIgUihC1+Ptuf5GimE0axwCttGT
vVWHfKucbnn0lZFdCncYWGTU341Bg3b9qi6n0UeJ5wSoKGRwr2bJfra8f0KmBzH1B6N781xl1Zz4
Lysc2XA0g+lgZ5v+am/E4dRdLGBYrqSDp/fOZBLUsGKDO5hkM8FRN03jeNqbxdPtCqcOnIHxCvFB
280h6met8PbZ/i4iV4IoU8SSsmsrVXvVDe2ZSWXlP0u3uWM+y5HA4soU6QdTqcrEqzutBiPDag0a
L46NWwWEAl2TmAMAmDqtXRD8wP43dLVoIy15Tbr4GXXn8BNRTALLt8gfnzM+ve0msPYYqda/cXPR
ipVUhsnoN2Uh/dfdzL+pO0cvAM+GUPZY1A5G0BAkTsz6XtuL/+IRNfedZCyBnnUNI/1hJnP58bJk
AyqhQtdw/a9oPV4dHD8Vcxbp6skXSgZ3mhtpr54huQKXLNa4iUNuERJHZBALjN+b7bpHyYCIAFfA
XER5svkBCjRtBcCctkZIGpfNT6DVKvG6ftW46scmmKxLhSxOPm56818iuzMFjKJ/CfwVGcYRJg8a
cTf1aLSBlDF+ZHU4hM6ykcr35e7SnLF51bJWzEgtw7b14knW/OjK7kiZX0vghi3GnGZJVBJqWeid
4hx9+eoWjK/7nWn9vFccNSmImj0j+G3gO3P5DDXmMUKsykfdhyyQVsSBZDxMm/aKJi9EhmbTxt+L
SWO7aYS4/oCm0h+1vfN3eIUycMLd3+qXLj9IHC0cUngddSsN/iPuktwPC5j3qBrYfrrSM7HyKAub
Bn8+SkyRt3ygNKrgaxfvumVQmH9P5rhXmCyunupr4eEOAwVxVaoMP/+1lsmAU0H4lcRRHaIqTeN/
FVvnrb1GEwdRztgbYhwWoTF0FeguN9c0EmYVr9M43IFmHepIYs8lU/4qYCxW2i2qqMzvvVozmlbT
ed/HDbn3PRZmLJxSDFh5A9tkWlHQEutwWFNKApufxDAN8ErKXBf4RV1Rql1KZayU6J/lWQyj3aPk
cgCK24RMF13QroYZKbzegzN9MjGmsZTrEc5wsrHYZeeygcjSPU3Q/9pGPLnpWlLkeoIbDKgR7oiH
PcIXrWGB/oaa2jSF82oTn49f4BrfPLzPuBz3Lfc03bKujxejE4kweNRoRAxXlyFkfWMHXnZ5537L
eAgIWY5rb1h6SY5DJteNZjqhWCSDLDvWBWS9eeLXBX6a3S76WwPSbUZyUtQg91zpDiNe5Qtshukj
4iITLf2s71N5oYtwn+8Mx8w/s28eY0sofj2fmswW/dbJQYmQcYhD0V48uij6IvxnsdjwADD4RQp0
+aFj+MycGujZF2rc58ln5+/mLKR/aptU++ecagyXQaM1hqZlbaX8U2A6vrnMv9YnNr+7tFZ+HKVL
YmQdSOk3LorPcfc4YXOUhSCYZu9ZUzSujmUBF48LRoJMAlHeoRGUBoE8FEs74Zkf9O9GNSmNqdbV
q73iNmQLklA4BlPMdsn4PaAOFj3umgvA6Iubb4jqQJTHIk9e1XV+iysx6fI0yinu28RQKxPBKoVB
yWChZu3DBILLu4v9UuYSHyo1vz0h0ew7b9D3Iq3IJLz/dG6H89+UEm9sayWr8wtUz3m173Iau54e
5nwIqGNfYAXjpjnnT0uIZ2QbvRyjS0ZNecJ4jmKaE+cTrDpvEc3Rak+qa/CcGA5c1eb1UQM0MvL4
pzhBXJxF3hY+UKaFFdzuPyrT1WbBvqEgTay8EXvvMmPLGsdbEKxwfFYfk44I9H39ab3bXIFfFWkC
/vuxRyfm+KVmYuh48LWlfNFCYnpowOynghcKhAVhlRhLi3nD4lSNdnXah9uLDoUQXqaKzCImXMlL
gmC4GhviDLMOEVE36AWCSaBGt0jfJqqlTTUqRVHmUuh6QBu7CS0JTVFHvyg/UlosKUQejuOVu+Gv
oJSZGDS2ErHMf0m1m6eDT31gK14vhzoW1NO3aV9fpXFn7GUi5mQRk/gi9sesInfqIvBuhqv+ekWr
6vetmXTUk6okxy/5GiJ7S+rVk1DGcdG50UV/NuRHXKS9kOaH0DYPsIbdb1ew1/3XEWbMxkgUPw4I
Ye5btsc0sDLQL5hAOTOppTc779FQj+mwEp4WVOXKVH5Hw5BoMC5eV6hBgRTxgnKq1bVKePSNeAkY
e4NWGIXBk4xnd7ZYGlFZbObdLEarR5xaQa8oKd7C/8903ZQ3DzFdL3BMopx88EpZdXwokpZ5b6F4
lo7W0xZmq0HCPzNh4dBGxEC6bRbsRYctYjE4cl/cqggE5s7tEVx1zTqT5YRPUf+jVwyjlhSRc/Oe
+eRQmHdawTm7kYvy3OfIGZB6f7QPSR3cX1YpHwGpGAGttxRwzpEwMWF1uWMlrBf2erCyvCLwlaxW
7p48Qep5GhsRiQor/9G78951+cFkOvbXL3rMgLM563JEzZqRlrrFu3SmORHJXPGQw7wx/iFOUYmQ
kd9Lpeovb6bM6ayf6PNS9y70+MGTmX2/F5oiuAwTUFU+ZqKaZzNldPFQwt+XPAYT5ubMv2QD+Etp
rkWVPBYk/PPqhIj8+PePT3Hd4VBqhytZeJtweCpTCjo+TT/opLXori7wwo/sDU3fS9g4x+IBYLuN
GKUFzoW1MEPpcxxkiLgxVqUP4qeq1Xkhw2uM9DeFtQCma+qIho2CTkx/7PPfz12B41lz9mFzetmr
N2MSel1B2U/t6+9GR56zH4aw/FldaFrUP3Moh6UTll0UGa2gbtudTkm4a0GeuRObvPkDS0Wom0l3
Ainw68MsUYRMPEqGOBLROZ+f0DZFrxP1chbLNIdBHGLoIO52bHkXjKzTHeXEH3xeNCp2LyqAQ1eI
a3pIKh3xrKfsD7OqvmHLxQDlMzv9IohJkAxPg8FGCd5ctOtxK4Fk88vrEEEIWXby+sGpFBQRZNND
FnIFM1O4ae4U91m3GiWJ9T6BRC27GK4ad+Y7HWEA2v+3qdgxzGr9HUXRZOGXJ2wV8GrXgIPuAjC9
zDCsebDrEGJkU0Yag0Pjuah/ykTulPxsq+ve1x8ljbB4D+v8HQZcwgNz9v+UNl4TUtD6rmu++Ja5
D8PX/7R4h1Urv8v5qSax7LxpBj/z1oay9VY0pLq8I01di694hrP6z7Qucn/WKS1u01O0VWurIg68
j9Cq1Q0sHV+M/yX5omcDmnEDWiQduAQRExSKMlahecnpZ9yX4emao9wKMubpOgtj3xS8M41KIG0X
dixtjfEvXHCvGKkdiVSWmoUWBQiZxpvqerOXX1KNP5SgW3vwpMSyzX1WL5L6CX8+Pmw/QQLxVRZO
IbM05tR1xIQ9FLge4Byxie7y/U4BhoGCFWxM19fErQ5sjCQYFg4JZiYh38Xz1Ma+CdJOgBsk/6ts
Ov7lh0zATO+la5gGDqAC4rKKq0oVJ9Yl2Nd7QrkfljWzjBOn5fjkh+mt/BdZ4jWZTm8HFT4GK9ew
bODIsg3BOUSlUrmlBr21qALc/6ymWISq9UjfEvRmaXHNkQxoj8DUcR1i9gZvEifahVidk34Ue73U
jkqoHPdhBGEdZOByP8NU06OOe1G6b6b9xArTUnagMYD9V45jshxRilpAi1ECGTRoKqG+AujF84bf
Lwm2JMKg1F6o5aUGSkJxaH4ZEE2znErAlfXCbx/CXAVYzqcdTIvDsq9ZUKCG3sqJVdVg+oLLDgU+
9LSOEN1n7TAOvX2hZ1efRuLGtRJzXgowixFWvyiHj+nJxT4JgidlLLjD8t7SlZ4leUpwCHTiWsA0
yLNe9biVHc40aLFhmUK13Mr2DliDToArxK+JhGUZfWUMSJdNFqSFmoVLunyy2Zo0b9rj6YtueZCc
44VZubqnP5YTK+I/zbwljNUM+t6ZLmvcnXm6F/35k1wyvqb5uTsS1fand5b/FOY3N0uUAW2uqJjm
egAcSltGVTWHF+SGmf4tIC05ik0Hm4w8/d2SfP008C8R1krzRorDrLtmg3wZWvjb5cByyDqjkrgn
iEoBC0u0MpQ51z4JsrAizbEMp7gw6cHDheZREjao8dWYG0dkYD+WWGNfv/r0wNYucrfAWh5PxGir
J/DWmGqKWTt9lfv7NCmsEacKUgsLeoAf4l14Zdiq0c6HNUIJfi6Dka0TwGlQAVO9POuaIjkZ+tLA
E4AdtIlE0RYddzQe/9k4KS9rWbxnLiJkIA9iC7BrZYD9rqzVUmDJnebODrXAf4g302tFkxVyWZJO
6y9ipEZ8fST/m8J7Ah8I4U/OijMOwhvc/r4l3F4dbHHQd6/xXkY8dxYekRRwKsUSgLxqutotIiaE
C2Gi1pJ7qdZIaQ7Usqd1e8zOqQdLKwg4ExRU31sO1WOt2zHPtPI0HEZmJ+h7tH6/NvsdR6YcBab5
sc0gbBog5LeSgfyKkyWc6M4B69baj/UnW+W17UBy9Mr10EJ422aKO74RBAGTdIX1msfFwJIFepSh
Fb35BMlzVOtgyeCCfqDHxG0GRmxxvZD0QopmwtfId+wztxWfl22RQry64bJBwmlusN6wa4suacLZ
E+G+MGZiGUzsTe6/Xov9qywbrYoePl+JoxKukeE8Gx1n7c7+87d4OVW9d/qe3FgOjw8S6gAEZA0g
9j7VlRrS4bGzRGd883aFGA7Yavo1Kjih6oV7AbYFJbTyMar4ry+5UDYZZcZ9k15JXpUxrnDH+nHP
7IXwPxxoPKiIHexCHpr2mZU8QHicrp38m0h7GcMYsyYnj0BzUjEIXgx/shnlaxoK9YEbXYWIGeDM
jlxrhNt7XtFPL9Q9WVQd2ZZB+0+14s58/Hejmj6p8n9wrpd6WBToYrNGchMUkP0g5G+Ef5kNVaF1
G9DifMHE9nxbU0P1CGbC8PWNEvW0uLrtIlpRmUt+6M8f+W8Rdf8Fmb4cb1WoeF3ALOUs944Em9lb
n8uU5hK6N8ss2/zgZgPP0LPJbIMBDVBnqHIdupHeURrNmjSx4iEWMsXULo29SwXO+g+cW06gdNxb
oppnZ97qu9lMG8JiCxycWEgyPUudjT3Gq2TaIyLlLCaS/5NgzWzTkyZgXvCqw5dPMDm44ANgaSNM
aoWBxvEaK9XRRGi7gGvPJqfRPwMc2OcClwJnKf5zx3j1pAkLi3hGFUWTl2VBQqIpl5R/nSB7Pf4D
4gPY5Q0CBnxRS3CjY9iz9ep/0+W9tZXrsUeo3HrnWs/MQilGRhmdHcNEwcWl2gAop7hwP2vnRXl2
5eTlNBmyEtD1CkttJoomOjD8djnMA0tSmUiL6aTFcxY0tpq/1rPzVtl/B/WdTRSIgYfq2V5SqlFj
BlX4dw0TmZZfJFNHigjl3yQPSovqKqXvVs5P1bq8IsWJF8oIyKAsFU6Pbu5UpMNEOEtXFpIUpDlg
CFT5cFvSRlqIrt5qM69ga54tsHaPl8lmRPD9Qxba+RlL3D+Bt3ILrys8ZefDRPWEzD518AseJf+k
pF/xedhZs1oRs7JsmUl6vzsJlu8zV9RDp3R5cGw81qBRZ4ZD9k0sTQNvqNFq5v5s2z7nwE8TO+tF
zQws5+5bImjvJvnrv0/lb9Hj6nK+7Dd7CIDO1pYcZTMCPJQDEY3Cr5nKvXPyn+1eQwhaw4UIhlF3
j6MPWSccFPr5GETVdPYQusX4t7ocrIuhJ0iFrqZDMbciMg1PzutGVDTYpsdfQLpY+J3GB+NgF06h
caHPo8gd4u8kQUldnYn273e1aO+7L3Kj8x6eg7VWDqaxPu3ktVhYHnMIQiD6ACSPKOQTokI77dl3
u980QB/sz3GBwxq8+Rsb0X2JOmi3YrXeQxlp8kM5bksw2ZSkTLtG0G+p+cBjsCCljD9JZEJVBEfR
IloRQmIeA7pD9AG6h5uvoxNOavKJN46B3CjABnyKWVKi/FgOYcTysqnZh+640huHTy3f+sr/lGc3
aE1lMjPITXyC/PWN2k85FQrZ1dm7OA73+dzr+BAQ5fgx9EDJl/Hgt1S+2RQ3+nGIW7egZ/mgx8Lx
TxzPlgp1T2TbDglkm1bdVoVLALb3ryy0gdltyzJHe2s7ZsM8eSfrz31wfLQ2uIy0imHQ4lgfLyoE
rurBdIvYE0OpGGFQadamIX6xD9EmRrFgSS98VbgSJnpzL1THJNa6j+IxAJReXifJqafrRFsSKyi+
mw5pDUW1VytKe1sYjqT7HIIuOYKS9OFofWnrb99Ho39g9lE4SD4Kj4GBlin1M2au0FjYNHYcw+Jf
SPATLt5QewqYMouU4J4IBzmiTXXThFr4chrFPGL9rTW0UM8HFT1J5xQTE17B7BdVYQvlDXofxZEh
lBpyeNfSjO5HS+A2DmEdJNvF0lYXsoEyH9nKRobbllQgERNZGUYc+aBlzg2/Lkh+ThI6lTwbZaum
+1R/5jPc3ryn20tUhiVjSFRQIhvxVb0rkBovb0gxv9fUfOrLLyi8xyA+oAmjpzwzeRLJo1EKF04O
XyA6blV0tV8nYAjx/w3UY+fSWMFKA1+T9y63QCryLnDyJYkrXtGFUnje8T/HhXp8XZD56vzs+oc7
zU52o34ReYvaCKW/SZaNdQsuE9BbZV9MwCS2ZCl58YsAqToJK/vw3+R+/AN2/pD31YJTi83uWx9h
YAYYZR5YZpU8V1H/MkG2Kh+3G3RK0qorHajtXnCQow183G4VkfEraSUhU9YdU1xbYc5Z217OaHO9
K+7Eq4/5cMwdnMVNwE2f32aUUWXbMQWN7Ab2B1vhSZ6R2xiB7mTvXJ5rKDHOlHMgLL8hVSXKTbCI
7u8lcQfa3rb89WT45Wnd3xahPi1uSY9xrAIhyn+GUKPMjZo9X7oVKjGUpPMLIwfU2+wmO7U8goK+
pnni2+9UesgJCsSdtJiPy3UbwFioyFbkn/U5AvcuTEnjihK9XOoBpToVbjcDljMYO/mhvDMe84Z+
6w9H2g303KEYpTYzi1HqbCCYYnhpvn9STYiVGOGFrTmaEMFQfFLNN/g9OnSzVkxc2h/Kj8CjZAOo
ixyk7CsPCFugTIHcFN8wkje2euDRapd2FpqCjXYQV1WmVj4UGvzbgeGyCu5IMtgbh5hYUBNw37e8
tXA6Afo4dVzD6vRu59UAFXoodN/vLoOGTb1DSe82cuLHgBrhthjNLPvoLnZ69ezjaqM7NvNs+V0d
OWcfD/iGBhNRzPrgtrTVZdCGtyJZJxYS+toR92Z5KgaHIjuReylYNhQ7UQgXFKzu9NaRWIzS4YAM
iAyVFjCPejnFcJa3BXv56ktlN30+GA9dcrjQTjdO0wXUu/Tb5c8PTmTzI/EROuz9X6q5nv0HFeyh
wNCHTcDKCwm71Yu2PAZMkgV17hsuNBHthykzRqo1Fj5dKBFrCtyxQ6vAsgGWsVnjtCoggonK2j09
GrPxlaV9EMzp8sFavu1jS4DxIaNm0d3cTsBGLkcXW+P8bVZIKStFtQUV5kqq1AxNJeLY14k6Ef+3
H2P5qGf+vedKF/IXgcwOPHNnprg1yHpSS9yV3+DItPPj8rPtYZr5oNG8WilJeG+09mUxq/0ZEACz
4IQteFizJxsDcpW9OS3fW0M5BJGHuw+TvBgzsiNy49U50KRIwm6j1bOtSDE8BrU5OcwAPaV21d6D
fPRGPCEL+9YyJc4CJdR2yYB+QOqHQoT/Y/1AUGHhfiP+vqc/VAO+2hmP6DGTfRJJOPwrdyLOfEt2
9DVWtHTGEFN/LKUHlKjohXz/LcomtDaz/tHR/pwedxm9Ozzk0UVrK7UuHv9p6BOesR6/6B4PgRxq
Uj8qcJkTYPRXZ4AW4j3qvs5WqmZL+38sQs+NFTfeH8EOcMbRl2WbwV4KlU53IV2pHO9tepYhcSNF
/iIhE/SRFITxJkbg5gffTdFQ/1tUNZGSPW56L0t38BlNrF4v0euQ0IxeIynHuAudzx7/2mfAskgx
OFFvXzcbxN7QvU3WZiqOFqWgz2Wqx83dUfNhU1/jR8r+kbiCayvszfCdpOqX51e+HZWEdYU8TLvk
hW1BwBcQbjZdoXIjl85U8wcXei9xFF1dH2aYcoSb5GRYt+l9fANDOFdEqQyjxgHRJY+Ko56yv8Wn
Eol5zAHlfRx8lMCZovNxemDgftLsqt5cYg+tdLeFW5E5SmW7QUj6DBNg3ki7yqwzGBOJxg9NC7dF
bJp68lpd5TfLAIX0ra2Vhzws1304ePFmMj/4sSnnF8l2kwQEFnId07HO41+WiqcLnBWQhLfNpIRY
qOJwECrkqsr1Qtz1l0rO1hHQcq1VEqA4ruWyciTQY3tCPPq1w7KyrLr16Mz1egV2JGI9ZaklseDi
sDN7lpe8a6EZHWAVYqkmugSNqxXX5BUEEbAcnYFd63WYNoaGp0wvA/UxclBfadfB7auOttduLP3l
GxM/ocAQ6hVeElsz0rHfJb/VHSvbBtnNiU7WJVMyP2ziHTaQCA9qub11aMX7EMi9Ql98Mbs0EUAh
QZRkiUhj2J84DJHlYG65e8lKKmFgBTYHiQa+HLIAFhykKx/SVAsGgXUSsm2CiW983k1z9ibrev0c
SSOuxmZgcj9Y0oEp1SyDowuYoR32ZjyAI+S2zJJ4OI29JJxIK0ONACMa/oJ47xRRpAROomSkujB2
qx2Sh2s3BIbx89opbCqYJ5WG3ZC07c22zvPyxLluI6Nx85OLBXEMlklqeDfmtB6fMXZmRoyTQEEL
4xtVtjmBwNv7Anvjrxx7Psnpn0hlYFwi6e29suVNSoVkYtozI93+Y7p0T0ayGIsJahqeMVIr9Unm
f5d9XKSGBOBkqvroyV1x6icvrZ17bnCFxH9UiUEBv1D4nYO4/e2qfZJHyKuFQYLLDcwCw1kOGBnT
eA3gczicgXw6ClOIL+D/F7Opn2tEFIKUQYrOCxNk8v1D87ixg2USwYvCzLscmqi8ESyV/Kft/JFA
T890jc/+eyWYIF57uqgVMlTwMKK8qbto015gjQzeLW7coyo0ndIqpPkw9WY8/7Ri5hgBMziP6AFq
v7osoy3uUH+ZaqsZwQEY9SGyBiG7UX7meBJQh7mKJpkjyl90zqHTAKb+cUFdDC6U9dXU7be0btqi
EX65mOG0xaBi7AfchsAgJh2ZF8o1L8bxfiUGn98m4Z21tphxzRTWME6Ur9CLoEilLWdRgfrpfBRb
qqWpnNoMZe+zvHvKARL1nOEW4Rk/Uoyth9G8lABzE0WaX6Yf0Wbwa+4IBdl+jOl8vQQ6uPx35u5O
jxxSoEs7zC/dnauf17/8Ovg/HNLF9hJquF+heMpcfPeIDD8CJ/FGGxm2YsMN5p3X3dPplXwDBhUA
L/Z52GmlhVNBPzKWyc3X5EWES/Hd86JkIlTZm2eTBcyxFy1S0ywMRM4+9ULq/g2G+bnSRSojNO4p
NjqyA9zpiCvGuXaUIV55yZv54+RKEBvTVlV30dEd4zjTGaFJ8cGYswMIK+ziLynYsrk5LMHMKix4
pO9bktxSuAsQJ1yBG3mgXN1WiB9qXYrk8Od/flQ17D26Ce3PWtmN+QJ7By/U+y1eyRqEZMX47TyX
XNs01hJp/L9SnYI3aPxSs3kcwJK2b6MVw8GqNO5B6uVNigJ1HeVCVPcVwAYcyz1YVjHrQQiqMyNG
76lCIIwsT6uJrh+N7eIchFNNJUNQxVB6/gLp3VM8Z8HnSOqAH8jL7giv2ZKp8I/sS6nyunxtXxdY
rDDp/9imnOfVmDNM+nY2VTtmklotokUIzYSSGSFi2133s3qRfj1hUqgyZ5K6MDZG/MGTh4jy92U5
qNcDFvEPUmVJ4vEAomlgcg2qutd42YGvKU+IyFo+OyCmHFKQbDuZyWTeYLnFSIjsMX3t5WLvnasD
as7bB43OozJV46cd8rTDXpEbnudR9bso6ARPT/gRVZ1SLU0VYlY3F0eURqREaZk8zsS78xIToUxU
pG+VOOTAwSKAQclzojRbebcisTLat9xCe+09uuTi2/BXJsNNpoTWFsW+o/DMCUqdfff6PB3odAMx
WvXhSphMLM7vn9qY8hFD8Q5FX4OWh/ezqRqzXOOrnnT3Ooth56n9jGweT/oEXNq+BJOz3+fQvDha
eyD36B9dmM1DxAE2g6n6zxv+2Z/lR9JmAohNc9WfmuL6yNbTa60xD112jNO+Q0KiPKAv43KaKWsb
mxCSN2SlIswJxY1ZGbNfnmiEU3eYHGnVthOdnIPdzwRBIPwnp2KRmjlqZ2o+fnMytrusPz76DtDt
omsoa20BXb2/H0xvTkYAAXYErUXBgbkO8elRNLBmvHUYGL3BRd9lrQeYoUAlOF/OZNuknRcJZIgv
U1C/6ICNXYjqPt/qQ+K1AcJdCHReGBaauafVGg/NwT70GnjW6Ii5ZAHUB8+Sjwng2SmJ5NhgQsul
e0v96Hi1ELcEql1/a9/VvO39V0kHTLbBJTq79YhuogI3nTn8T2IJYLjAmUfu2ftwuZnLMJuwdw7n
CKBcbAtk3E3bfYIakegSTcjP8TzAuqQ6SsRq9VU+0sYPQTDh0QtMnKE4jqmkKUpGqdYQOSxSQ1yO
4IhqQvwVIH2hM2pK+900gmscSbcG5RyZuLhgppf/OIIuyiBLdUkoojOjarrNktJW+UnKoJXteVAn
4slO5OwoUaT7EWDK/wn/BVsv9B6bhbDSBuD7Fmjnevr63D9QOKTKG1mSgqmOLbMdfjc3POiFLjJM
zkMT2qgKfGbIpx3seKqCAB1Uj3u3ymsa9TpFqVnhzRdyLFyMq416FayZmgbincgL0/PXm2xQh+cD
MBQIOaNspvZCICccoG/XybVAJjKgJdhA6sMb0sqwpkbXg7R5NMcdLWZpMjnztWcyJ+8wO59QZEHH
FtLSH4Pw2dyYwpWFVBli9V9OMFJOynnWsu2z3o4dzAZD8p101VtRywl0uKM2FUT3NciLZTUZG+i/
jzaQL0zCOkWM9bMaczvsTAf9w3ZHCWXskdEpQqYdHhLraXqmVXMruDW4FZugw4DYE6bCmhdOkDN6
AvBhNGZ4LikUncA9d/dmbka7eiRUEz1aldUmAX2aJWlXCsCvvR59V3tXjxrKMIcGi99lnhrW+E7Q
IiXjLinsUdarW1kYIgllwmg5h07h2oI3+f+0o1PrRYV6vUL4pAOqMHRtKf6H7k6kQr4nVnjcDCHA
jOfxopMTTVq8imh4G93xiFbFseFv4qukmlyxLzmPy+uNaV7pj+JS+WyxwKL20Lsk7z64wzR0Azp2
uv1zSIqWct+/ct15CnRJWy3SR52oYvHxn96+RBsz+PeNhRDS7YtGLwVvQqejR42wsGijyNZCjUnn
+iKto72ZuINeihi3b6AussCfOk1PBowlqcXaewUYHbRipNrQAGFZ0xG1JKS7pR+KEPER0Itx20IN
egrXsG9Uo7W1JOfdhyOcch13eV4/0SHPISHsqDN12RmIWqWtDpBOQjkcCiDRM2+mRnR1D0zLS1Lc
t8CYGdb1L7okx7bqNcvIC5AJM1uJQb4ihMTKhwbVJVfH9mbIb68mWsdj4RLJfuOSIEN+fvAB5wAI
lodib1//1P9GoS1tMs3rtfQeCbbt+6uo7YhN4/lL71Q0BV8uNu+3JkNSegZoKR1tLDSfS92XIw18
XMSnn4mA9rcXLfHdYbFXj7HUhxR/oSxaEQm1R4IZYRRPNqPqThpdzzpjzDGT/U5FzYxh1UG274sb
X9DYFMQBKx6xl1U3c8j/KTW3Pw1rqoLElt/NTPvDn9g5epGCAJiXJzaTebKULy/G6A5rAgC7+zjb
U108FYNXaa6NgGBtDHQC9zPkOF87ZIdGX+H2CCVH92US+3p+5EPpurbrkS8bc04C304zJ4/tIRyB
ktCfpDOcmYzA2xYo2oMQ2gep4MzCASc2+MU8yhm3a2Jsx79HxODh/2+i1QSiXkqNfYj46LfyX3Pd
I7OsqUh/X6QgMEWdsgc2T+eJ3abFy127IkfpaWwu29SCn9T9GD8OU2Qvi8HkHf+SSePgNqc9/59s
JTHvftVlh9+Ow5CYZ3IuLB+5OQXCIEoc/bxrrzpBvKucYdn/0eubkTLInlGOcKahl3mnu/8E/3zt
tqJxsRP0xbxmDhz1aUT/SNEVOM5RxTs6xrLnz9zfOfbWD+JmhI6nIsZKNpAIjkEWR0bDijfa+RcC
03IvAB3Y6oAK+4QlNCt69UyCUEE/L8UfQELsAAxu7bD/mdeLTITbApYB8WRCcuiZb9UHnEAyv0hA
gGJq0aLRyvd82vihuBA7seMTHIG0MQP9B04lr0CGkEeSksOTMcylG/JvVVlRRyA5akUG2KhTYwMp
OxkubBFufol0Hl42Fu1eaIDL66YMOdszr14YeYrbs25U51D3YHr/JRL81QUzSySQT2jWL+8Tk3CP
+HULWht45LnTqErMa9VbBWBYAmXanezVAWIf5SVXmg9bs2oLwIDRif9k2Uh5MmmEojdDEw2XaWPK
wH0bjjVEcauZw8m+P8VX1IZScQfiZEg5M++5etaOh7q+ad0nrZzAIjDXEuaxEJVAhrzqYfD4fn4o
ShN1ZUUuQ4EowvVJf3aCjZkDYPSPpTNmMoo+ReBktO4hUZ2Ov+G/yXH/YIVeIDIN1B2DSVNM8gjV
Ko7FYeIpO4va7VHE8BLoIuSb+qZE/oueTp8PHzIA8KKmbJnI+/7DpnTAKlv/YXYXizmcXfDQBS49
iInApwJoQzIKPL9L5QHtpAU3h5bDke4Z8erZJEKMy++pRiq9h2HgEHGjPRxHY2d5g45lhZ9zmOuU
ZcCyDVaCsRyOjy/CAoHMA3w4ipgMaVxxCBK9azdg9BnxIL04zbpdgawwtVmvFXn+uHY8WqTf2Ica
eNdSTzcuf3xUbwM0BBuLXdHvGcwkWGt3l/CMj3MFkmi7TGyyPqDyPVVj17bP9SF5HVcahofFKNU8
3hTtExb6JrkqkRi5LDYUG0tym7zJFhAq+6eVn/tmrn4y0NTekHxX9q+KGBNuGWATS8APMbtDDTgQ
qqHA382gSOAtrDpqvhoTEIYgh8qAORSiW0/wwRw5IZvjPKHG8GUEdi0Xuhzti0lCXNBx7r08u6+O
KLKY5KP0O3nZe7/LYcWy1YNb0dMHlaeM5Gjib3/ehSXxL7nIfy6N2/V84FobxvDK2NFbfSsJXuoK
np6XnMeQNdBtrygcUTybFkDicT9tIjMQbgZ26HBMU8EFankqG4kQ4LrUbGjr7w/0fS2V6b6vlCU7
tnZKhaz0IaEzihnMhERa6RUjCSqhXwFLEJRu+Qgz2JdW5SJDXOQu0peFmKtcbExTDBPnWqVIGSXD
0vNzXtubOXUemNk3slPYbuDklXymWbp15ih+cINl+f2YOhcKw4M2mBuhgqvivKIZDWEbMqRkGI0N
OWYJy1A7r/7wKIvYJsDW2Z81ylMdRe934cBfxLdMwUUD+qGtmw1lNeADWVw3L+H0Qkd6PKClqyKt
SgG2JDGs4ku6lT5sxIQp2mLayXlFejGzZ1/Pnsrp9STjKvDkk+iIAsojp1U+fX9djcrYUO7Gq+7W
SUoboe14Rxw5wAsxNEqLvU8Q2HLsSq4zIUURgGVxuM/VPfD/d7gjgEnNUBaz0S3Sp8IbwxOOzC6b
3BgfAYEv56MgOkBeDzZklr6kr8NCRAow8luHoxSx6uzEKDvwSkDzO3/3Q3lVMBVntsAil/GQDbZE
liw6JQ2a5trGDLso0L8lUkPJotgWk500eNAsXRPAXxsBH3cZopoIdJ1d6P91q6zdAQ26CyXM1hNA
IuPZWsAsbCkPDBvbRjwqHybb8FBzBUmTQhul3zteNuojQgQUYSRiUg5f3dAKQLJNADbghJELK41q
of6aPk86TtNT3v320o+JfXvkEeGUsBQQpbhuVJDwStg6Sx9g2LUd3dySXbaItYZoiLvIC6bCW8n/
E+QUf7XnbuTOzfF7kq9AYin+7Lk33C6WgDuIcpy7pVpClkgThM7ecI41lXmtcExJiFCrHe4iBhKj
/gI8ZXS0/cAMwVeRsfjYPWhj60HFo9ykyFzJEj0w7OAamZp/7UUNHa9bVeZW+QLkJXcIdq/3lobo
GmsutBQO9H79OH/oRsVa9T3KZEIf3bho9rlNwC7ig/Am/wY43ggECGY2HaMVMXMpNSvp7rGicAjV
WCCHu2it/+BPRTbNSn/sDqHbm7H29LAYduIxKfLY5rWjlAAfSC9VuqQP1N5eGj+UxIjdIomz+Brg
DRBK9Lr5B+ADbyyoM9QuKYFyIc64RmXs2iBRJOxUcCt+qQfkkLZ/ffIFOyokobaNgeKTjjANdvFI
OLxKVojpUoUDMTldrvgqh8QEOr3ZUqzKcwaNZ/DXOJsXOSyGQV3IRdP2p0zFoVfaBcp4JcZtgiuT
fzgEFONJbbS4nxDeF4fIVVqDZoeZEyrfIUocv9sUd2Svd23zGvNGEqt5wCSOVuH9xPiCCTi6X3/2
cmIUzaJnWr+E3ORM94IWP+pElleyHjZ2xVLGyjWSPs84QXGAAn3zWSKEt5aefjLFgmVgEKpKovj8
aXprQSay/h5Kau6VOcixgv7Ohjv7Y1LHsum+TVkl3MOY0fjmZeftirfUUa5ivpRn0mOMHYpFP8tZ
WA/V3u89ZoTMudvcXbC4/m1+V1bsrEmbMKIwtNYpIyrrOUnnAF2GeieMxO6v9+SLHM6ajBBGKFhS
JAO8DSSHCtSXJyNQ7zSV1PuQyNNohhFMGBxzHzF9naKyNhM1MoMo6ZetlUFKE2PsaqodbXk+Ke/j
anlaMrIHbyq9blyPUBzKnBN1CazlhtS9fU183FFNufHdyJ1KAhG+9X+cNjxn1tyIHvPLCgJiVdU9
fDKoUezlqM1ndIlDy8XdWhV9Jf1MyWoLPX3ye5nfoxYJYY6dHlTgW+9wusOmOrSjJ9dHYq66Q/C0
jGMKvScoe22MfoFvt6HnLHnV/N7wW0brpIJmgykseztVKeb7EG28Cdz0xV7KmOUJx0dlf2AeVc2i
/djaTOcR/2Hx+a+9x8Mv6O6jeYs7hCd638s7swwdBdYWWL0xRRjs1aILrW8+XugJo/E5fea0g98K
rq/MKDk//ojAsiVFRJ8RcCJ1p41gProucSivCtaWaB+UsfOuGaQaZ9O6E2VcTv6ak8e8pzw/BCG3
v8tsvHdCwGUO19ZmJg3JilOM0l6DNehhDELkE+E8VqlDyuOqrEIuhOvNp+y/WSgqyWe69Vuj3Nmy
XcyvTbjGae+Sl3VN17040KS4tKFVfsrfikJvvW0wJrJCn35871xsiIy4Aw3gvsi72HttgeWOBCpW
qPDZbzpL6WfZxeDThw6bB+p9nQaZWeuclzNb64NgeE8dtxWTf9eJsGuRf1ucaEcVkzEpewanYDVs
RP4bgLNWUdLLAiQzGYEprdzLeXPaAHWnQxOVfDpROZ7DfE7buba0H2D51neqz+zvMfdUIhjrVTiL
sAiRO12LWlCecNRyx5fPImNz6rv3WT+jLE/vsDGpPdLAO63Pn//bubdjB+lZ5D803PSV8WWVR8Is
BHWEqvl6D9Ib3Eo0UwGdovPnvFgLUs5DBmiQ8HlmqzpvsbLi/fro+VbPAsMkGuqLFNnCZ7yevnZ6
MmBWUQW/oVCr7R59mh5j5nHZTcI9ycl0E9/cvLt/WH3xRmHRuJMM4uNC8i9lsB1JIP6nfkJjCtoQ
adEWtiFC9V/rZGlv2d3f3gXoNlhUQYOZ4nv8FwUESMpXW1EIaySjgQk6oK8k3YWfmyrbzWgHGy+L
QHUNnz+gWk/B/4JxjvaP7i5jxliSFl0JmeDxtYDklSGUwBnHajpXanzkU3c1oB911SFXk9GvDZ8d
rw9RzFxKC4zPtypYLM99lsluZ0YesejaMbGS/ApIW7URshdcyWeWTpkPqMIRfctGGBMdJVP84YUF
YwhhP3vgPu/Dxp+lOFvdxSxI+gSuyikpy1vxzQOopdpYFgwGw/4TMXnYDNKARUymVm0qSs26RXuP
aYdIiC+h4MMkPQWbpAuwcXFsWYGb2DZGFrFPiKF5Z2a8MU3gc4Z7NXNkTMESQMpy0RnCY6hFOge7
ac82QeF/mYOY/DZ4KOY5TbPcyM97PuvOYyjb+f3iEkxTptVcfKSqGUvf/NkfHmq6vpjHainoR7/I
xXKzEczzMcSvYqqvY9+4U4avopfamzJaCdzc1NIb2HiMC+vx/mgwHUgqE7oj0TjGYIvgjOBB1CPY
7LsaLMNt9DK+1eHz5QufMTT7+Mk0fPW1CxWajPO8nNHv2qADNAkDedG1K6wQhLHqkR06sbbNqm70
Dtg/RYde16W+iYbKt+cA3k3k1oFZC1KIqSP4pn1n9yQKPeYr0LSJFJutqdAGgC02ChmgWdMfdq5w
yPoRekBLlUSNK9v95QlvDa5tCbqYEeCfiQt7X87lytMZRB0JH0Sna2w3MBjUTYFDwnvJssJ1qSHV
xxaA0pF0tR3r3IbT7HB+tFkUhAKoQ76exjy3YHCAG7vlmSQxZ43Wtk1mmSPnFZG+XWDZBn8DyFFX
Abc54jRNkhOYICHl7LnOJmMzUueem1eGUZccYLuARGdgVC7Hk5+40I0xB2DoNv8kMwnAIw2vXxvI
+6Pg+pbgF3LZOaV/P7xdcMueqMouzkyquSsjELcxq6tRlLC6ajJc/tW8N5l+KycSyQQLhcrrYB1H
LUtqrK4yH1vfTVUUqbqF0M0H7khQiAL9VGB0COXn+A597cFHjZJoJYlIr8Gogq7Q0E2RG1nDE+aP
4Y9iA10Bmv+gtPwNDb4/f95ryD/Pr/w5OXqkpt9G6sJctbnG/a/SHbOHjgjNXeulqr9+MI/cHGwR
1Be62GBYXXi7i/ThYMtqeqSkFJi/3tLKQbI7bp9bNY5WHifOa4CXjyPL2bpTQk5nG1WBozqk4kH+
XUxsNKAmmi2A/L6pVkpNGNavzcAjkvSXV+6w8KabuTzstEi30w/3vvRPtaGUanTmisYCNh+sJHyW
gIbcK+DWL9JmqNXhOCVgv0NwoUvDKUJRsp6HEJIcvKUe5dBY4Kf92FbEhoB1U0/e/Xv2UQ1/6EMI
wub/agQPXQbnawUzNAyq9u8UH6Svkurv1U3lgXNnrYZWSvRAXw0AZm42NS/+F+Jmy2cH7IjoEgQJ
e/6L7nj69oVeXVpiri08N0M3VjkSI14Kp/PQaK+r3gpxf89UWqTerif/15MFQVizDHtGTkXuf/mq
nrXdWDBup4Og74flhcjdGy8QNL39YCLy0maPvVgaWVmya9DW0HaUoq11EoMBcJPXaFil05fFpPLq
2W4xZyRkhrbgE+h7yVg5HwtzGU/t3FsUSFegfpdNIXZ0A1gDEh+XsSjf0LN4iBxdtZsEKqbhYDg3
aVm5umQ8tu5u1CrUGoDAVuAHhjLTpa9XzUEQ/QyjAY5n48u/fFCDi8lOXpIknCr0kvh/5k7mXyxE
D8V42KKQBPqDNlTohYbmWWtAU9pleHFALvGWceVMSESdj0GNTe6yuzGLpADJ/aAu1hK/rVzz0qCd
GNsV0Rw9NyLA0k3iEeKAR3a6haivMAeBQm6rMtzh7RUougKDApxcICQoaWFlSwjAmvZ3iJll+qZP
SdrjXiBNTwbaL7govS9Nux2onbE0dWUF+pMZ6J2vM4LbOaYdWNvvC5Bq4Q1MtxM2Y/nq5H49o95I
Ok9es0vQU7rJUTVWA1kPGoyIV3Y8zSwD8Knv7xn/1YQfTXyaW09XhHr3PSs+EezjFjBWcHSWaAIP
Q7KNgxnSeebI3tQXqyn3IujFxuVjD1yBhGaGKYDeiFeoWKPc+i2M73OXIIw5lH405i/uBp6psZqE
fNuNED+VVUhXwMZZfl80Rm3zByT4MnMOZfFpBoRxXNMIPdBOhS/lZ5q4WpqChEXhqdIXl5yks0mX
FRvKCm+MaDZEHYcxUZSP0FWq1VCf80cypHcan8Q287ykDG1qqdg6R8vk3dAis09JbPNTc8BXfMrS
v4cG5b+4fFFg8TFq+ySNEro1Hcx83E4mFmICEnAgg+s+W0kOTmzUcZY3LIQjGwYxCzozC7lficis
NYnkjTiNh61SRcJf3HZr4pgdvD2kLCvZyl6y2ov0L/Ga1kWs/8SPRS2/woGXxqtV2UDhUG3Nfeuc
CqdY90+mTuch252R5em6hUnCvEbZSTauuT4b4w8NJCQW7N/eS34uOPf6fObiDoz+cmIhpHL1NaVz
7MmaMAV5QXGXaaPHyt0quGWEDR0cIhleqB+jjZiiWTxp4rBzkB0IC4fszmu/9x3GCcFqixEFDIjD
TjixS4Hs47DbSIe1/hHMoGtVpZXV4zyPkxZ801ax0JLVWe5V2i6shlgTf47WTr8x20QZFIy/lG9u
AImK5s5xiMw1seHjo7TIpEL4xKm1D15ZS4p3g0HX7+USROfRluod3PFGZCCXuX3UEQqtWud6bQbX
2gAGkszF1XKkiR/8SizZ4nZl9l4/7G/cl6Gb3JTq9ZLMghmIOoulZPhn4I0Bks0Zo7g2Tf1tv8TI
hS3GxBw8uQUC4EVCMydDIVGrpg4Oq/X3vEYdvdMSDk0SybIt6WOszpjZr9U5ZTmjPnhwW2IyCZnk
aBSvXfZD1pDTyLp49jdZZcAP7YA5HpfasjWmkGt0TZXsQhHdZwCQuXeogb7tkDqgR+DWrSZmqKhH
yFGi/F/OQlGcPG7bfl7t86viMRQvaRyjXGxVs/tMNG8DR8RpVpk/7DBgLR/W8pM+lEIoYS4TjnSR
L/hsB+brraqXJHlWjS0INoghbcP0eZIYCfGroOyohK3yEbbkjtYDGjRsuiGoVG/Z08Qdyk519mWW
EBcHSxF4stXMQ27iVX8xvrcijiu5Vw1T32ckGaGQzvOyPNNw6HPKadpUeWeP1KHE0lkEwwwc4Bjy
sTyd3SoEhaZLCGoBss/35VU7RaSzUDJO9j0bPw2NmdFBS+SCGNQ/eNqA6lKha3aGzRn6vSbebF3N
j0GJMMVKfMMyuFkKhRQMWbRiBTbyunrDPMjnpOekdnwubieQal3ybOia3hoAk/ukCCwU2TrphCBZ
hUUGBiLQaPT1JqFWzc6Sgf6HLP4TR9J9AGrpQfhYOLqQCH47Z5E/5phfauxHfyPK2kz05OFUbdTa
usVlOfh/funLuqe7/xGiL0APxCMBq49ykthtF001//DiAKQWZNLV6OyZ801v91pat8X+AmNYsBfx
IZruDqWYQkhb9O0rXG8SuwR2jSiOUNcFhofRTSpbOLUAF8FeJAnjFfTCkiLsT68sCI7DVtg9LDhW
7RzrVLdS1JgxXzIpsc213kDEX0O7orUGnqXNbfSHVHmK7470kcw3RrDDPXuiAY8F8fgqvScTabjb
ll4w+2I5yi2JUsU/3b5SEFUZFO0uv/gEpdCq8y3Vv0EJWaeqoAna0TU3SkbBLSOtbFjXzWrU5CgR
lXBgfnaadVLzT4NVKrBkTwjy9WX31XCt1S439k7Tk294EncBSy0dCXBRfcM4EQHqk4hdoBkw61BQ
y0P6IbfojCsd/9S0jTOqHhafCcgJxB/xvbSJlgz0EDjuMhm8snycdI0KfzdD/YSS1ES7ZPFDxq5D
EUuih0vrQq7IrZc5AuOz+dqpUjpZc9x4rwVjV8vYyVkaL7HmmnphpfFLVy/Pl9h8+5EN6go5QxRF
dkqZE3YFrZdBPeDKcoD4IeHn1TFxHHUznFn+0M2BC+OzKqB17cKg7nyXsBpLyl8qeEU1ErbXB63+
XBSqKfFEdEFa3sLDv2/FcAcrT5MbUi3BOEwf8rCHoYxSx0BBY0iRj9yNhM1po4snLDANrk4MQFaE
6ZB1SMiC2r/RH6PSpyIGGw2L/JcJHXoR4TtKPP/TD2gZRljCWmuMOwLepX/FoJbIMp8mAjBDHpPx
ukEVhdL4EsVYXacUu8JZrslETtTlLqD6rjPjr/Pb414XsRA4U2tgy9oX0RYgXx8c1wZIGOtwsWwW
/xff4UI07aQ4QpLM7PZ/YV449nKhEHGAtEo6TL1OWgJXVePUH3yx4m4LjA1HXsEsKKurRx+Fl49v
yJkPR7SG1tn9EN55ZWUBXQ1vcP97JcENP+e5Vtn+Jw4iNsg26v+dime9J/K/Bh5FlhebouviIp+c
hOBrbNUtak7XgO8tvrJXjlMnEXarkzSyMFwsvYncma7AQ1l+BOiO5eTrUfCyOTYO2PQNgWnFsSsg
87WMuR6YgLqGXG0HEoOvkVXCJz4GnazgswmimrnN11H3B22lo6wFLZKB5IH1n3hkN84V6XbWe3HA
AVBzyADxg6zbvXx1hrvYjS9jUZ7Sq+t43DuC5+Y1qZO21eaSTsvpPRrfsVjZPeCzK3Epqj4yZOra
YWD8SBG//Cc9lC2NevrXgCrbT93jseAVSbljHbrE0bh1Ycprqs5ureJQgEOvBsPdwvAHSOH6qi1L
orslE3nDzapMBCqqMjhptMBbB/Y+JWsl2ZuYO1tOba86J6Uchja6xmbUZCuWD1GfaWyYz/cAim5T
gvtqh1c6HIbes27S06ufmy0jUIzWjkUxMNQBGq1D7ycx78QXV0lfuVDJ+/HkL9ljYUxlPxj9p+3p
w7NHoZ6iy1Ae8fG3n6HgCnoyXA7yfIUZT9fxw4+Y243g3db/Gt7C4B6mZw5Kcfz4HkcgBxpKEYrj
KUMbWwZqvTayLtbP3Ok4rQfk+v2gtACGIMEUULvdAIupe4a8sVtloJa2yzertV/vQQLFrfX7tlFV
436q6USI3kBS0JS5jPghMVUSTF25sbrA4hJqBLfIOkpfxGMyBBgmcGCB/I3ITLi2gLDrDq3/6Qgq
0KOT6iLNkmlMyYd2SEEsLfBEXDAI2j3XHFrADnBlF9mA0zuQT0EM/5P2bYVJBdxlRARbhaeCFYcL
uiX8IGwvUiQhyZih5JOXtRpaiPp1bdSs9xqDxKjdoWotcj/MpkAZV5PZv8B681wfXk6FwdRK/MMv
eA/jo3spPmhlqAnsNodN/EUU345sKxs5NUuAwXQzZFxNcoPj1B1wUTUSU9oYfwyUV33YYjI9Wcya
y0JrfiIvGFfXrz3BTrOswftrEZgZ3cHgPuIb2cBlrAL5WNPnqQEpvIZAnJOEVI/k+t7XvaMdlR+J
P569jYESAfKGn1t5vQ4UG7LuoRpjBPtqVVQDAGhwrKaZeZkuMNXvRI8gbqPC4umy77KYAxTBIEJS
8yXyim6vqUkvRGwUVRnRBQS0bBt3mYK305ZmKz+Oy21xtYLW3EN1p8JTSI9zRz7kmNR7bFAglAid
6jVtmItJjDIf4XQRqfPF84cqNTZbl78u2W2riWvdvMCGDD28rU/uC6sqtA2T6LShQX/sdKzgbbRx
OHYdYjmjuESsccqOkuN4YING8kNZxgayuzNa8g/08uTac9jM3j29I2m1sbLsU7iaSNd7Khi6K7i2
2EcJerSu1XO3g4ytYT/oZJdL7Q0ShssegDjf/ALlFxBTvluOmL0qeC8vK3A270XcApJRMdVhOk5O
iNl5qUjZ1MZENHmNkhZHZBcHj4y+9ZVG3Znxs/XqvhsuANUP76a9K7uohQuNd/6Lzan4+wogFWr2
2+Ov7TOPRh/pF0chNUumIdChLymWhm+NKQjSn0N8WkoWatf4jDRal73CWjtkk5ji3S/0eYG0vWmT
FH99QtOZidFjk4vMkfpNNjeh7+Ep4hJa2iU8eFTIWfO1WxbYWD0d31YvdeYWIxegJhLQZZtjAjm9
8m1n6Zg9a6ZG73WPeXVjc9ckCrs1VLHKWMDZNEpBmA0OnXdRG3NivCRs3EaM1AQp6rNauzyTR2x3
vtU/ernDruAOawEjY0Y1yb9yNPawa0pIKACtG1A345VbVsJw3/TxnZZEuFpWY3jxNBZJaePItWFb
619CuP5qRfhaAbCdw9gEPLVJYr1hYTgs3y29HOeO9GjdQmnNQSjKiKZslzCmxHbnnyDqg8lM1dEZ
c1v4ML622sdFAIy/bklh19eqKh5fl+fhCd5tsc3F2s5aw4TgDa7udxaGeWSwbO32flDRjppJLyQ9
mVLlhVf+7PWYPYFSVVVDoBmMSq2H6XbrPHTJv/mdBMq/y5ZrF6ldU08CSV6mSu3q3PC/V6Eqkndm
TsfahzpnIosGKTqNwHdp1oCRZE6gZVNiDv3drSbQZCN5l5bJ9qU9vT289MO57jYxmqALcrffe9YT
cP/RKWO0YhJ0cLV5eOiN9Nq3486h5MLk+kk2zMpncuhLLfGi7xt1u5WOiThp5WfqmQ/+I8AxgO3T
Y+xAghBtggjH7RTrFL8SNBw+Ohm0yYrQSDBDlRjMSNkv4fajYpCQy5qp6TQGxzZxHH8OE3/lK9mc
h8yjBVuqKIV7jPUdndp2Bjeiha4gFVxX49PgR6nptWy6VSUyDUkvkswEThKrwK6Ip6sNDoG7b5mh
iMbTqasrjHE+LBycyGde9GMpJlY67BYBoCfP0BE0t6shsOdLYKQpmY18wOZyTHFD5Dfidb+3yp5a
vBjEbMg2VjFRRbXTBirUV1ma/kbDVF/0ciqB32XFqufsW+6q0zh+PxIkUN0kvXhYGMwBrYB2onX7
RJLzZZWwxM1FKMbclOg+1AGVoS+JQCo92xbiIxEj9P4A2n3rQfjQMgtrPI/2tc0T0aYGtJQngBNG
PEkH4RNZJpLaHdIY1lIRg6offoqplPZrHf2MyKQE9cq4IShdRwGMTaqFmIyh/zuxKXii1Ruh5+mw
8XhI2KaalsxA4fSaRDCBMZ4rAlbDwAxntmFCRw9HxFAhT50789KZphbwhKNh+NDpgeKf6dbtLVu9
sYwCGpyExPREKVQNnZWw/uglqHAIbdI43GlQcSadi+uFBV5yv9zt8xwEhSEk+TWW6Lac+Y4IotqX
qM9TUfW0AFj9qha+56lPFur3dAIe8ruRlgzQJ+H8xwMOknYkRsGfhPrAKbrTMXhuunY2jVFcCp3y
PFaC3iJ2Gi1W8cynFyjhsVBHYynhYI+1tjTU5hkO9G7Rpwq4njYbA9qIECc3TBI1+waGMzv6rHBB
zaljnR8uQO1+9LtuOWlZQeJ9JpY5bcZnhSe56lWpRRDfHPf8XbImmvKyTuMK0uypxYc31f76SIXr
mWVUMdlQYs4mv/4USGePNbNE9kA7npoGm8S3Uc37cMSlK+a0D0bKCb2xmeM+QZviGjsX3oIPQKXu
rze19vT4bx96CznMrtUax681K5U8n4BU9cjkVpMQtM3uqHwbZvCwnmXb1lCexxZ+Nzs7/+AXUZiJ
1o5uQkIi89CdTCg7ZEQOifg1aHUCsD7OFIYN5NfokH014RGIdYR74n4woe8WB42hpcSP8aIUcdiO
3OyUlxEfa9qpL91LDYMw5Cicie0y/U4yp0XLSCXPtxMMU5fKKi57wvpwTXMsmzXylWfW/+3SFF8p
s++4CX8hKn7K+o0a4rhoYJTcMY/AoBTa4Y5sirVSQDqhEKVWOXBqW+4SCnnHhPVyJsE4t0UcRSvw
T7UhMh6dmWF/fvpG+nmg5m3pMH8Q9+Yr/FrzL+Zt4B4zia3dxBxw7tyDdSwoBNTEd3tiW28KltNp
BtopzidaO/8xzzLIgColO6efLfAi7Hio/z1XYSmShFfHMzGZ6hFgACSDZx+EdyEN1r1W+JOA9cVH
ZSeZQDitQaYWrbC6+U6DI0+HCREBgk/pBfJyRrE6CFwINyHJih9xoZuUY7rwqc5hHghIcuK1Yv8f
Sw94mmUpkIRRWUCKMRvSJ30qm8TfMAfw11T1cbFReqCPC1IUWh1xDbV8V9KoZFPlJHnTxe5UdkcJ
pqGqvbBKGzUXrvsu/dzn+vWZ7pfeFBCiDM3KMTy/XComtsfE9rLIWdRIv0VEoeZp7UAhg9itinf/
q7Y56KN61I7Sg5WSs5bxOpyJ3RmBkLFNR/5cB5fq7jriFtsJriNvCoMK7w+WsGa9XT7kQ+8TtrL1
xrsDJAbZDTNRrtZLH7PAc9Nx1Gp0VzEeOBYgy/8fdzJj0ZMawFbJc6mIjKME3fgkvwMHQiQRFNOy
lbHI25QbtaQtFraT0/s7ZF1YPHvlMSAQKv/RaygS0eYIyBx+/khhyE0OVTzLpa58ETWdQDHlbS2o
N8ShmI5koKPlPzrT8XDyh411BJkOZwFcp/i+P2iKtiRfGTvZdazwkcZ8c7hv+Yxn4L/53Prq1Ys1
pJeHO4DHWs2aRkCJGKIqx8c31iAQqSCl7HjqnZhciayqcO6NYXxf6Q6JhecH1w2WMBt+2XzQegzo
BqPPEZ8XvE67QgxfY9jbMiB8WuzrH0LCV9ee7xRUiTUI0xDvnMmL5SfcoH7fSedUDFCnKiVVZAtH
va+PjR48B4vmlGoBPoHj1sRmodWKO6ALHvkzsPS75EC+Ch4WTsWOGy7z7EgtkLHbZHjkW5cj+aXw
daL6zlaIwSSi2Cm9DzQea9zRAQqi/ze+eaXBqGwyvfeuMcuJHbk3aLEChJLEuvXjoeYnPQEjJ/3+
OcbrnKFJJoU0cUv1qh/eTq9Rsh8Ynfnr47Vo96uCGyxE6lmLoWASANohqc6acAk59lzQlaY7OGB6
9aC/h+BYmAa1ftMcO0uf1H6mxoNxWwFRAMHJWSJRD+glZMSdmm/unWiuV7ii42qDwjUi60dfHEMn
9QSeSNSYDXY6QpGOBWBRmHivS76Z/qt+3jtRqBZ0YTKWBa4yy57ute0WJnNzH3i2GVbjWIwY4DRo
hEo+rBoQA+DhZTmWPR+HXPH78SbeCj2U+Bq1CS+qEYc73XVydaHBy4CZvOznCm1+D8FlVL3eAFQO
hIrrravVKxIjGV7UviUlzVK1M7fl0lDQ5TUH6fRQQJXS7pYXh/ha95TUPoQxy3mOWF1l1wEEJ0a/
VnRmGX60zqG/cwNmR0ONj6UyiE9DEV7BuUIPm89hxFvLX/ZzOkkbtOv4uZ6n553jtdHyL5sVSSuG
iOxjEaM1kjWutSJMbw8Tqwgf8a/xJvGiD/LYJ6cRYzVDZR7VuMrzmSUAUhAl8/tjMdaf0MFWkMyi
dm8G3CeYOMf15rihX4ftjaxyhG/IwYKxISYnt2Lz3u8o4huz0UAa0+Socg5vOQ/nczW7S9HiLciA
rCSx0Njunx0X4VCL1KGi9dwRuVzQQZ88YhUc5CsW7jKuj6hqrkmsBR5r5d1FaBc06weg5xBzq/2A
8feM7bpOKJKez2mf9hIfwkBGtURO1br3yY5kBb3i7Tw+z6fJsbJuMFnTgQ7U8qVjEJjhfMP4eL4r
gxza5kdAdRfg9tfiWCV2hXZzYBzdI6GdwYkTWz6EWeeHJDVl+nkYAb7K3w8ZTIz2bSuPb8QIyiHS
SCzQuYdp5OLLv2vZzNdXDNP1UAtkOTjB8nOQYVWHiTL+GiyNbXf3RPrFKmrbjZTPCTAYKYVfB2DY
T5TrCQMN4VKyJe3A7hJmSl4XlVCQMLgCZMg9vqNtsEaxHWyI7vnUoBY/S2554d/gNqyMmWSwu433
8U4B4JYklZHejYRAVfBnktccG4wHzAH03XuqLPeGV0xKk9F0FACH3lrFsm6scVnpWXDNC8fQQazx
EtIYyEN2CSKDQcy7/5SebFVZUrZg6+robRsVv018jReICxEktU3rCJWIv0Ku6O8LP13GUBT2xBIs
rrhuukvfJiJ1ed5TvNgTicPr2zrhDgV+PBMLbwVuJzPdrc4ayNKpBo0WtqeWfiKlew1+nL65kF9U
APElWslZgkpBBAYI4upjWFGhcjPvWDx8cl1jUC4idgRCCUhl9tYRqP3PiuqwBTfWTXQLFpwD3+aY
gszD+am5OkbWysAZKywwnROF+b8r4toH6A6l0/n2T7Y51wggJuGvqH3nwIydwUOMMYFOiRDchAxU
8dhe8xVzXOAegGBwzDb+rygd6FZrAmeNZ3n+yL7Y2V6mWLo2OPBUl2/Y5Djp1AxcRKEWODwi93qZ
rw7XzZos+okHea77QwM4C7UZsR+awPY//EMK2Qmf5fjsld65mW1TXIlQoxd9X0CzaHlda3J2NpGL
mbRqTQ0sxkc76gWwJkvbwxjWov930MeEx5Q2s059Y8s2fbb80Y+7oMjKkccBY5lXaHt7Ogxyi3ts
XjNBqd+mjGCgXZMXcTDvs/VUB6Hwja2AdPq3kz8LOxmQoXE1cMK5gUHp9EIoI5PIee8gwrqNQFUt
80XrFLELvOmvRirFrxIJD6lM04hlgsS3598jvDJVP4P/zXv8pSw4F61t+W49JIz1WVLQH4nnavas
j80moXKfk/Z0f5B8Lb0ALF2jnrsUdSZ0q1wnaqWjBPY+N/jdTEaWSASyeTAOlTShgNAbFhVDJQPh
ZZcf2ThkP5jsj55EI29AEyzTQDarTVywMtpfPsgQKUwHCN4CkXSyyI03oFy6NOgLpTlWrO0qfDpT
2GA/0RmnaSoenc8517Y9cF7/FXBH1XLn//SGVdjgp3zWt06AEu0yA05I49qs3iSPqvZA8h0Scpcc
LW9KvP/YCttiQKT3B1vYCxgq4xSNrBUxklX33/ZxhL1ukUJ5O1Iqjws8qZAYvfuyxVAOmsuQLQKm
B+f1mPo4tDPYvQQKY2y+7632Wbm0OZYLxrXpKMxJ4yplbDZZ8CFeCkAZOFuatf8VC2UkPXMN9JPF
zmmCCmiYfQRpSwhwbRTP/dtrTMHqrEl3MjU/pcZoBfLJsv90tapWAwubUrqpuWC9arSk7YcfkFBH
ITbIM4pjLA0mIBZrYSx0lvrvcIbgdz4EfXEpExlTgFw0MX9E0k/xF9b2Vh3lCkyD15cvahD0/Yhe
KWiELYeEBIZsGHNCT4TH2K94DLzhD2cIZYjtAhM9yn0Pbk5k2NVhDCYi/oP9+kHtJ5QqIq6JE4U+
vHyNMZs22IYonmfL+tX3MUX2ipL+Kx1PC58Ut1DfKyL0bALu/1NsydYKCR1WYykOZ1eJGynjOSCO
bMlGoD/LtsbG2EFq/AOepb8GwbxPqy0OfJTOQFoEXtywtYepRJF4LiSV04NMT63LMvyFQ6RKkubS
5mBKJ4byX5+yaDFjLZX4aR9Gpx9zpIElkQpVOHhsXDdtAhzsFsAr3x3IBoc6ae6YvXX04ROdO2CE
NBDnG45YM3DR8rrVsGW54Nz79zTs72Ojdv9hh80xFqzg4z6DjbIHrK3itx2vvuJyrtY0WhSpvwuy
3T583ZXyEiD6QV2fMbOLn/VYE0mp76pBXHE+JchKUnxG8Lm/Cfw9yDeN8m5/dUALhdUE14ApFpIN
2quFMklJgo+GkYGAlw2/yd/eK5lzokfTpScSFEMHCTo6RcPkwHqwomvkjPa/3rhfkh+/WLSSon4Q
EpL1uyz25DHIlc68oFmWVKGwX4mdysUyd2Gsuoi6dnT45yL9gVrDGRdt1Y+m3S7+6XUa/c/nnqEq
MUoQTt0if+NPNekZiwZtXrNVWr4tHfMGqFBLb3i0uGgsCKITVzS54Qi0G/y8n/uM3boPV/GxVS+p
1sRgn0NlHaqrNlZnoao7Oie+SV730tCagqj5fMwxZoX73U0zB5WPEVH0m5xWxPz+3yNuRU1EnncR
xRBSmtdEyQNyEEG+nN8tyvVIAyIYk0ePg2go0ccc5g2bCSoeqQ5yjBTphl6Xc2x1Mn8qqPSM40QA
zydegAJlAb+DGzDqQF2TimIQmA9yP5Mo0fnXawkhfMUfSqEAgpyUuU9cjMg+w1lFIxUx/kqcrNlL
y43iRsilO3OZJ0VyyWACJxeBIEgMoG9tEAU4lDxHhZj377J3/zUyMy62E8ghPjJSUov10UISO5JU
mZs0aaTRxWoaUUelDL1Fttku2jP6wj2I9y+D4QpN8P3cTjZWS023PFOeRXda1SaAa/9idVMZAx6c
wonT/IpsP/DcuAWVFZCaKBq9j6HnCthnyVw+F06LAqJIgE75ZbwrMNbm9JoYB5/BUlPZsWgwhBuU
wsBkubDXWYGliVxZSKHriNTNQNSPjPVMzqRVl20azsNLFBqHREi6eoyXUBf6o78IvHTWnbWx3HuK
WNggo2CNKF5/NH7LhFpFo6ANtSQPK4sMABWbwESKmxIMy/cNENC98TIuzv5WcrNb8IuxwTGC964d
/TACdHucLCUsmMJPSF7Ij8GBO3oWvyFXuCa0VAGv9nqQ52omhI/kfsx8td3c4YqmbGxGrBDbyW/J
uJwPzBfQxzIs0ZRRv+p0Tu8rSU6f+wSrBCVDS/4yXii0Zeclsmo7Py2Sw5ix6pQWOzBRvtSURNeF
hGHZznjGdQWT2oS5TW06Dt5j1dsTBj8KxFFpAuht5fryQ0yFgL7d35CMf25qxpxxW2Iw4ETP5rEk
c966JFieSEHakFlg0wNkVK4UMpev4TTEf8Hf3oB6nXMQTu17+eS51xCI9bL1WedjdxEtmjYXeE+0
FYOs79DVOeXG5FnJCbvkP+5G7LlHo0fffzxUDOfQUiEmNuEovWiCh0w+/AtzcbumtlZ7KC8r1bDZ
zI6d0kEPNsyegP03QdYpGJqeiYkxZdsiVSAfgZko1z6lyO2sVz52nhw2gioCraK8cjgrpUOyGeZu
AIu4zzmqjq6f2WlOnpuhslzqCOtmNmFlzaTvuTs3r+1otfA7U3LZXsQcpg5/KMafU9ZWd7Tvf4eX
W8n+WQOuFkzqXum67b0Wcbdnkal+/BelMZvvXbqPVP/9d4NaYA9bflCilhls5C9Iquq1aXXSSuxJ
pptjgK8J2sYbCC2i8T4o8c2GipNtVcEYCXbcbl1hHXQetNRl2mkTlprfaOck6rloPSErJsIo/wHL
drGhxvJvpuzzE/XOnv7LWWeIXCzh8gbFpY3qEdNeAYUzW7TWD7klZJz2qTmvq0IfoJkRkIIM+kOg
AAN1mBMzCWmwS/AznLMkp4BERFKLnIKOra4nZ1J/WqWRzREUFk/6Bx/S4v5s7cERpZKE14xCCf8/
QBtdR4V7zgCdDQeCVCPPXZfDkO+67rcq0B2Ey/0T0elC9u+S8AduLFOCF1MSaVNHbXhV7TT2iUHa
ZxYAmDnB85RYWPFdDmNoTXCYmWmwQTOcrpBmyLN96lX/nAdlwWsI6ZYq35N7qvn2vP85IqPbG/Zg
dX/d4Xe8iIGP+GdrXWWi7oaZ6x3LeERsFniL/e5uw52CWYFRBa8jR4jFzRK/u9HYfjFEymUYWQLI
5llItmakWM6086itWR+RNrieET7YoHXJwHC+u10PXXv81n/THV9EiS4zZpCw+s6Z+jQK7F2/Ft58
RPrxj5/EB941IsQvjLyz7v+5J2hJhs9Ff+Lb/l33HoEaentXAy+fBdoCbhB4F945oG0zrl4RyYw+
/SJEDFon3ZysYxODZ89ibNbNJeHc2CYvTMuEuVyJCCDap+Bt6Wp/DG8RspnHXD80sLywB7KGnIXi
nwBbacvw0teFA2CKD2aJ4RdbCHF9Kfd4qjCXxfiZkmEi63qXlBsegBm6z1aju16ZMajiWXpr5Xb5
dYKkSgsyZosY+casDivC9go8qc6mm01T4xl4w4wliQDFdsO+Y3fnjoCAF3rT/IVcXj+KLUSvqE4S
mea7pygpvW+io7V5KjgEQ+QAWx3bOYiyaoNvXr4b7kMvtIMXjW9cP2/R1YUG8cf42cildVm5Rs4l
Kkt0EJ9M1bYWqc89IuWv+1F7jdv1U4K9CAzIn8qzUrLtZty/XQf2dVoDQhXmeJswvF4zVV8PLhWI
PG+CTQkggOlQdIooJWaSLJq4fjB9QQmwUh6JSy4qduK3QAI/TySo3ZRupHIbuhu2Z5Dg8FdjQxwK
Y4xP72tiMVzBM8htkaekJbv1R/Syf7QXTdyajxWhio1zZq9zZOsznygg0Y8WZnyuNohk/BV3WSdi
Kr1gHxz9l+Z40+4FVG0D8tYolIuV+3Fiap/8aHjtzrer640cQlB7Uc5Hg7Ya0xlnhJaStasHzIUS
+3auGvFkkO1VuGvdVQtXs1Dxd5JKIp2LOKUjF8aqsM21luJb/T2SOnQwZkEzYAwJ8HzEuvKkyhjv
N8jTzxW6Qef12GA2AO+5tFZt/Ak5/ODr8Z2b5+oA44aI9ARLzZDCop5BVzGYZ0Vs9lgvpQN3FG4S
clNYltIJyinRfU1xxU+/tIcp2H0Fc9t/BQDnXiw3EwZI/+pGF5oRhC5gXYcDlSS4PWjD5aLk3VnB
qcu07kcb9nuH3sHn60Wb4BtFvLRwqsjb7QCP6TVPuHIqi1xJSLNU5n/+zeIEB8WZESfMqO2lof4S
hEDhMJhDZobKgJIMhin/Br3ZdDpQ2jQXFyA2+2GmZ2ExfFTXAqPUoM3jYkYhfXwWaN0dadT73zLV
U1FfGAq/8bkd9rqshOTmve9GGdw/qtMCYM2aQ+THuOxNIbukrG+i1ipSjZTh71zSPmF+5K4Jlvci
F+yvTzIivBSHjq1v+izqv5yOefavnl53XkIlEtIuuhMYfSIG4jdiqbQKSKSJfqKFkLme/BCYO2fv
AJ9cpnZjGvLaHGkaT2tp93yHkHV1ULPyov0IVL1OE5OEkGPC+UH8KirFEF/FLluljZX35G6IBgAd
GjbkrjDl7JeEhr23tgeRpRKc1CLOkZngN6no6/fLphLf9UZucNOqCQH+rkxEugQDvSkWmZdGeuEf
qksHZ29Q02pgx9H+YOYzN6DMbRLsyWGN7bn8iYqsSxPSKJaVhSFm/057CoOE9tdj0yHhZFlHGZs7
RnUwugMnIuZr2HRFjYpSZI/ALyaMQyWd1sUcLVSTtwv54Qm2El8OKvZeDr3aa2GxHXh0iCw8wcxQ
lLwu+uaA1Aoy7wgWLr57KzG/fZVnJhAK5EvD+6eauNKSwnD2mrLRrgBRVrDFfCnnRs7Iaffns+pC
eEW9nMTIP7QcZ7YkifNOXoZ9dyXQGhIGkZaDNFi7FFKOA8JPsj3v8BkUQZCrZCC4mKlsSA8i3dyT
FWTlV+53R3jeiqcusOGTrpAovdq1AIy2UOC86L5Iv/6CT1ieAB5LhEYQVQglS5yNqSBgbScY1jz/
Ow+RZ/kcUG7Iip0GcAxJEWdNQG1azqSnLtmqyYdTGzpOrOur3squvMiXPFUrT4xS9AL61tTFwSWD
yl5F04/cwoqdsFuGIsd66DdXcvbP1VemsnxRJH1Zl/fbg0Z4Oc/M1V6dTbivzKB6ZBmqextwdVox
RxnzBUdktmO2eCEf/Z8mxTx0rEoUh/AYHDkzSWxpFEPONo9bXJvwQP2uOvZnZ9IB7VxCtqWWHsSM
sDSeemg6pxKREQZdApI1MdiMvwgbbmzH7nIxRVQJ3EnlyO/7F9yy2rFmoc9zuCWrakDJvNckGneH
YiQHWfnNwmQhqHoZxrdxGH0zAU65bum9KW4DzL+KcDOazB1xO4UmH1RkiLnHIBsUR/nVPvxt76OU
GwFyYAKjkK0hFjdFgY8tYruEoQNuqWH1jzgwVJ/kGF4goHh3bgwNZ5vIVR58UiYWqT6wqFBraHNA
LojK6W0SEiNbhZ4+hSRI+SqZZEd2uDuvN9VuO0BW7Tv6jDx8QWab43Ictr4THJRtvBUpY+jLRztB
FMCk6m+0wHM4MlS7lqC7WDvio9rJvF2Na1ApsIzeLt+B/Ryx49wK+8L4GSagnPA+EuV+XpOIUJ44
ePh1ilehHaTFtqHTJLJBtdDJXL5z0BYB5HcJjnKwyOLzmlIce72ne9Rr5UWzIXaNdTsnC00+jlUG
PuNftKA1CWgY4IDyMqqFE8WYliIgxD6v6XBCm40DnxCFklCigrPxSYM3gnLGLL5ldf/ILEuy8sf1
XoZr5vu7bepkdXuAuWNjx4SfY9aEajjNdL7T7x8h4oZD9tQQ1MI102qqEP0OT1rHIsR9IGJnXgWk
JHPpjJh9Mh4IAqtqBgc1adPTnogXdnjnLKDvkKWsmgMFawgRJwdFQC3E5Xj/E19noekXCYRk1NRs
rIr/iiqExgK5lo4hDEoCIDhSkN/HTFyKrtbdkLiZoIy83eqfz3Okt0jmAxm/5MZzaYBwhJG4aqzZ
ugT9W9+krcWNvUXips5YnhpHp/gt/O8zBFYRgusAuKCh7EZ+kg7vnO9EdQkrCg5zWkZ56zZfNRlB
+K76Rj+bMGSBOMv5r+Deo8qlGEFjk/2jQrydhjHzmXWjaTfK1OANXy0xFnsjENy1YOENi8o9jzAy
CmWw6rersIlnzd5KFGTUIUbE18YWv0pkZPizLHTicnsARCfcpMP68pqvFidN15ckAExRhMbEZbZw
AbIFIoDhGkkt3mZBodvzcVRbHjygHgGBTLvbVAZIcNdG8VSeg4TcoUXEpIF+/OS3DS6YvMgdSoQP
MihX9iAPnJajn3BxrdafliIglRfVT1DQ+ZNI9FQF7E3BQhY+CKS3AMHXgMnMo/i2Upuyuadgzgqg
ulVzmzsZgQ4yHgtpHOvzxa1dUblPyhuTVnd5hiAL+rLHeytGAAmMf3kffDpgt66UpAHGysED3Tlw
qPjsh8xNNEZrM3VZcGVNSuyijSwMJ4ONeTmIqZGTvcBVMIVAbWR9vrisMbRh+j6FgxsnKEKo9QBD
LzafWAZe6nzQqyLgfc2e8nz9neTAfk00x0T1oVw9/+p838JnUGRaFxMW6HEckUJ5A6XlWKBkLlv6
GfPxz9eU7d7ESnH1x4ebgadih+WQfnfYld9mRcnBP0GW+7FzVp437gKSCKJW3PV6DkFwW9Sv2Yol
mFBKUg0xQoluSix/AW1Lmk8SbKQqLADoFHtUzTMIUTZMcKVtcr9vOjSYEadAWpciqYBdlXdR8h6T
eSFJPdAj8epgx+axEOTQzOCqcRZIVaUKlNecjXHmITid8qXd2cs3mBc+kk87HGgI8P+OREbhGQMg
Qfk9gSG+2EROn/IAIqQGKh+qf9LdqFVZbXCUlZ5h4Ghv9gak/CgEreHvVtiQRQYtpgAILM8AhcZG
OkD9Q3eMUa1xv+2l9NfQg1c039nieEiREhSNy8/WM2YDm/BUizUKhkHTjjrEvK66XI+SSPdYwJaa
t/UXZa8Kcb4Xf4q/t1w7ziklKLH6ByaSnmtjHtt5H4tqB/tzkYDGab21c1AV2+QpOxLgRRSARfLe
EEhIqIzs054iteGOw6qr0d81hn1S0vR/oBdycKIkCpye+pVMIoiOxMPGZsjYXqn5iNyzPLlD75XG
3NRSZj8T2j7UIVBZwwNTTZU0plmqd3m939J7RaNCgHOUfeL6joFVMD3IMeZJTfuc4P0ALLjWO3fJ
68C31ySLfZZc9wniM0EHYe3juH1PFd9FuTv9O2BHEdxujhrS12RWj0C5JjzOTMuyevzf6SmomNK4
DcQgh3N++rn/U472qp+6xtjz9zcp5Jvdrp4QyE8QBYVlRHRNufMd5HmEVje/gXlN9cATyKu++YPE
1FsatDXagV3FwwljUTrLY1ABpGBSUPfUqjpASFI8XN9q7xN1JiGjT8fCZIubGkgyxLzYZOM9dfeZ
UTg1jCvRdwNz5YY0pE1CBlQc9IHZK6RZcyP+UU1EKKXp+EmLiuuQeEgE2qwN29w2eFnfNSoTNKxV
48r9XdX74q4gJwLiZWNXr8g9ioSA6vBVpmYj6XbGb8PXEervDirew5RYt6ONFPyfUrzAdMrOyWME
O7weN3hl5l6zrPPUxj8G946hgJsb7cjKh2yW3/z3YsglSkE8cHgY0+Jb5oOz0uZ5BrMu6+ZI/Eaq
peUvSg4+uPSidFmqqpUhDwXypldqy65BegEUy4yxTiZMOfQ3K5z4Ue/BvbBwaWPh6fzQxdbgROrk
qMNmkoX+nJrNXeI4gHbwmWsNVc6YZWCStDUgyPYu1GuEgagdu4nui5+a3cSAmL9H6PPg4VM7bMuq
TMcBynp/BkDpBCa4JTanh8bGnVmswe1AStjUjNI4z7fptG1Pio/cIeUOhz8607PoY2o2sRVdukKX
TlIAHnIMQGcH0cJ6IM2GUfxI96EFZ2/24i2cMeHygyqIu6J2U562hWo6l0GLAdQGhbK7AiGRmT4d
zuZ4DApUNl3pGdgIP1g+C+9b9JAKx49ms8UaGDwv+2QfSQEm9EM1ebEDv6eFqE5P2sOhbPUkJnS8
khBsjXSb+F9BBgaJKvwThAkJn8aDo8QI8kBIoUMpsi5BEv9K4/VX2b6QvRs2qqljOdv4TCECAh77
DigEvP1U7jpdo753HVNGOTtWMcyLkZLMGAi1sNHcvdVZHBfVMEk9okT6QNQOI+RJfd0zwrOPKU1Z
iQULFG4VUwjHSG2/dfJDzEZ34XTxPVMkLX8j+CyGNSEBWaQ/8DFu2xYM2/iYq0XFGj4mP7cFjmQP
k6jyW76VgmMXluExdZteahiIzL9tV/nd5+wlnB3/Y2q0UcOuJ519cwazvgJQPRTNx1h3FpqQ67l3
Q6B/MMWllx9jeZ1NlVqzb62fRU3/kcyZc4C3Jyhi+Kuz+WVvsYDpOBxqpI3fjCaz+D7SWHWmP17V
u7PnxlmfCXD1gFfjGhl6v9KCR9Ax2o90vfpqxEu1Xt/LEwmzCrdP0b1nNw6vhuqw4idE8rX4fxSa
f5N7MU19jo4BluRmOfvqmwCPeiBFAeU2JEthNSOAy468AlJ79dt5n3nyNBp4bGLzEOw4W27qzMQs
6zq1so49LR8G5naE3tEUPah6FIVY4AI7ivqwIoYr2Z3q+AiZbSNfbmxIY3QG136qFweEGjUXIXZD
aH8YyGzrrhTMev9tP40WF47b7KHbwbQF7l6lfPF0lDxHtldpKS+0YjX/6HB6gAaopguddiAIDkqY
gc+qSLnWLSDrplpBZ8taFgPFxFAsG1MU/9TFS9ffScFCbHER7ouO7b2xMEco0F2GMDW4LE5w8e26
u8qychYzvus5fvXAyjkly4xAH81j/+e5gzeO3TiR4rrvyr/Vs6bG/AraFHriLSLl1ZNaj1DC3WZt
0fDxtg8QJW4rcI7pUxYMluRcNrWR0EKW5LVHyVAaAkUvAMbuRsX39nEJdJpdx0dplbl7KGaTsGaF
sIkKR8rIEZZYVEBXOPrW+WNaiSutb0Z3yEswWe2mPsbHB3zdpB431kq/mpFZG/Q9yvu3XYqlpxDh
3wai8lkwGIGvYXtWaX5DqpVpNH84gGV18XO9ehRJZBwKkBJEYrRJidQ/N0pXfQznGLtzw9HawhHx
lQv97nRXoA61anH0QInUbatIzJ1/4nB+YpBESPnexpMNg+4BDOFuh+sI4bmGXyQQhz/ugibX3UQp
DddLK2e+vrv0sYyAz5TaPkW6RQ3DLwKW2/Dsj6MsVI/jKnp0wWkfQ42Ey9XKzUwaoPP73n4MloU+
OLFLSPGAflrpUw+J5KWFozQJnnriJawny0YpwDrZZk1aE4UoR0yGkMJkHn8HvDeujHJGC03Lson2
uemgt6D/lTckmFtDOcuFupqQbPDZKmDus/e6LuIlCRjolBsq1JtQPL787AAwiY6ZNkQtkNV6+J5W
9/evUnR+fe6Cet519wYSgFfkoH83rBiiiPQHxbyWc85zI+GGYmqKCWAqEsYvuZmmYu65T5C2se+i
8xiGVoL7+1M1KFRo6dFmu+bi8k6iScg7cz7Vnzn2fOHqoKpCF0Wyav6rWE3F8fwRcsAQk+r9mko+
1QZELZ/alv9zmUXMjKVRhnRMb33KkZfaOaAimq9QeLAuggmqj0Uk9sIZ09cvO7fcXtsb3MH+Z86e
0YE/6PYwqK+xfCl2c4sUH1v2bkYsxqa/22P6eFGusxIYGMV3wzj0FcLZ4fMAXG10u0Ml0BOAbMF3
L1Dwadna5SZ3o8mVUGO8VuiqVJ3X2WJqlcaevP+pLI86TXJzHlW4/adYIh5i8rFzFSBgiXtDBcgj
zWOECcZIzUqHxJEPFLF2Bloo1sCiJ2kgxCUNsHMgnmRKiXt1GawNM1/XBlg3SKNSdk+9Iga7f6mU
cGlxw31E6z0QnHmOPnpO+2eOvhpgwTewgZRQ1PLRGGSq18zInTtldiwZWQlRRGmPOzB2a/CzH+f+
Aju503jzsMDVHPRLPQ4V1zH2Cb83I1fCu4UVINViu1swMrc0MXxBzEs5hqXnQfClOYVmHdShb1HF
1kocnF9waFgL92CoQ5EctT5tiYZVzyNv6JrvgmxG8c5DVACpyj41TwqlmMF7ir8TyJ0XRiXoe8VI
NDaUxgM2x8xLP+bzHK25spgpf3j1fcqI4asSyianciJXFSawExR/t5HvE7rZMQ8KG9GhF76B0ET4
0QJSu6JIWEMjzY/RkciRG+Y1F0sSWREtplnemARUeQdLArw5BSik9/95ejdvGlXbZQOu2YGBgSLL
SYc7DSfnNzya3JpoGgKyWw6JCjJc+vWv+UXf9Bdu+xCL+65UHHYkm4j8HtDHDWrA3QIr4Y/zBQzz
GbKCDuXfSupOvr4aDJBShdcC8+rc8Q+OpwzWI1DbrpLRNSdUqdHJYkiWLicBQwWU/mOxpZgbNIWG
ZUtUR91q/VXLypZBUIfNuUKD8RPybzHNDU0yBf4ncNmX1O6DHNtPBrRCXvZdd/sNJFjI0lvZR6RK
etaMrlcCaRewtRMae/xFceTBbR7LpqG7+mgx+QvKlKYmkHUgCZI2g4LFUJSM7Sq3rmQJQZTGZXnp
QoR0ziancx7LmRWFOPfyPim3ZsorvdUDBUJIH1gBxb5Q0iL0jsvy49z/5CZFlSPiwDSRCVUoPFb5
3vlWTdylpnpfW4q4JjR34R6yuQbhs+TUOeoSbYuWaJHR3jpg5Ol7UPWMenT0CeYrI20oRpk0lmhI
FIf2ZxNU18tnraXpJhjWg6IZztxewqCpinJkKne4rVeXHe1QCShDQ4SJI7Vdy/0ixf/gPB5h3BMM
ZNPeZwOiVfSjlNSYTL1O5AoSCQVyos6BlV3YeGame3MYdaFb/Ah07fxI7Cl1vzuY1H/U98UCNkdm
P7RnqLxv1ae6CQcPqH1Qjb6V8F8dFaTN2fBMkHCBmbwFWxg45x3WmTalIwWcb0j/8HqYTqSb+cOe
71VypoqjS5jXZc+70ATLc/BXVaUqWSWx+5zegXpCFPf25CeJQPZPUFKdzDdD2CJ/WZvr44qlfyHZ
Wajn4jdBVQL7P5irIVhaE2wLm4kiKMAMN68WxswYKNiNKzdJObi+112+N2xb/cpiCuJCmEE3lA/B
KooKa2die8RpPlDofs8QRcNNuGUeELPXKKvzZbKA4E0mm2mpU8O3ls8GmVTlAchcq0K43J0KRLa4
yWSkvIzkiVbQR59Kn+AZKYZZkFwClVYQKG0UDYZCi+vd3TKhr4Zievr2FzrOHt8qBfz2Q3foX997
4nAs0WmdmXpqpjrE3dek2DBpH1wEyVhieVaOXNcQ433xheZEU0w1i5cp4bSBl3BW0SuRqMEyvNLp
5+Np5sN7wQJLD4+6ejDaubFaOmST390mqN6SuiV/fbTZBXlEhKs0y+scm9hqKJezeMXyptBlznX0
4a/AEj8GqoC3+HLPRhfGctuYXwBZ5rjIx/ZFheoNSLEqyVui0b5bFgEYmFmHM3Lzy4LrqFfwuasY
bp51Q2Z1E3g3cyWzeJpB8DRd7tY+yWTZt6tefOtr12dhnhan0CXzwEohNYzmpoVpnLJ4oL6XYQK9
WqIejCAPqF08RzVNXciucTtormz9z3OB/nrFXANmfa9Ys4JlWBCsGN+59J8dyAR31IaQj4N4AXdy
4NBQuUCBp9KIBNNkMULmTyhdUECBzBz41l7bGt54q+eJ5vFm0sbyvtuD/fnTGYVEJyd4F1sdm4v9
MJflg8KtnTVE0NMcBD8G+hXHhhpoiD+IP23HbHCeirfJS7JACW9pAgHYJnNhyD41nCSTWgBVzx4N
HrhhKkmuRdL1cA761wHfHAG7SdlxDKRFFdLc/jKAwqgQknKUi66ibMJOJFT5eiL3FMcSDmeszXLd
l6s2vDfO0qph6AfVoLlzoO8PwyKx0fsn28TUDi39eJ74JKmrcqZOyblH2jMO0Pu9R168H+ZmdZtD
upU5RdREsT+RG8wdDwkw0KIi2AW4PJlSE0uJd45CZlg2Wh4zqxLVs+bw7Ka+dJhh10HtNez4i6Qu
XxZAcPI8weWpuXu5Sn8J3G7gLCT4aby+r15tbGx1AjgPE0lkH8+2uBrwO8DEqPNgHbKNXzZYzmQY
WtKWcZpkT7Jxan2W16qasWTZeYFu/UWHq4X6a1fR9QCXaxVnRSqlULvQ5Yrj9rT/cnYwKFXNlIid
ecRnsD58Q1YlsP+k5QqPPDzrwOo85onAI2CajEkEwelj8Sk6fEZwlNuOtGlornW36MqQ6dL4FzeL
8Muxn8poxx2gdlaerZSs+ljp9k1a9f/aWLygEfV1Isa2i3qtmQqoOctpHBCQmL6oa4+P3bXtZUhg
/PE+28VdBNXdyEQFX458Qr3ZHdFv/AMl8eUuoMjkOlwDwWRw+w5UnPBeWwc6X9yHI3q2n3EHAspC
pK4yRmZrCGYtZVMxu8FctncNFb+cpKJE3DbuCa0LHMk97fq/Ihso3JY0MLIBjK8HSK6E8lMM6xcv
XgS5MzDFudn2oOtygQA4nHa2x0DWgnvvGscemnqNs5Hg9j1BCUxxn8gDJWJaCM9Rqcp9yJp+J4R4
caNRg08QeFRk8WhYLugqUbK/Ppx719bF83O/cnpWT9tX0m2/4NZh1ynqaQE078AczzWXH9ysy2cf
W+PEq185LFcXSY8NYgnbshqNuNvGJ4NSHUpgrRuTsVaOvWq7RByj2MOYdoaUyV8PXj5mFxuEqToS
ZM45ShBt2qwO8zXQdGicfLqXGbkOWQfS3aw/PtwVkYwjwNdgjVvYUMcJyk8ew2lRRSmUk6+j/Vnq
SR0w03UeO2BOtae0vqn8G9fop1hAdzdGF/iU7dbHzcR4nZ1lvQYXLmR1Uq8EZGRsZlVo0tS6zb37
ZYPgGsisxRWQTFySbV754wTFgzmBH1NVwwK763Me0uWF39z7LWUpwVktxmCHWqqUTki08T93UsNe
8oCj4YOwlDpUJWR1QC81abF1s0K5NESnd1l8jSpSZqpcyYOXAFHI9qrrtaxNGTXybSnyHNlc7tuN
DG1isnOJmqV2TxyyrlFi0SOyFU1gY3rgSdNNBU/wxxb1jfQOavzROWh5iPnbn8JBqG8czWJvEj+z
DDdolzV0JjE+zc43gZxF6VWsMQz8E5B4WzA8ixB9QHOFVgUhKcMzENRXp6hnf6YinI8cYLJKPqMj
sEr1yG0hK6mfwSqfppMDQ9DoCF2pXjPp96yU4p3KWRD7RprGIFigouDgvXLVWLk/0YgRyBYIv+DF
ZEVxhSgtHdADgjioOLm/bMPCvx3ksB+kKb6KoXu4gGuHmp9zPNQ3xOJRaY7pMVN8EDd5PhJvSFps
83LY/lKLVN8sOgmhMDpho2vs62sYI8hrSrPe7yfbWHUaAEFmT1ukJdh65Xykko1/tsIDAVP48k82
70G3cOag3EH+Z69oDTAOCLlq172XKmOEH4mnTT//6sKg/vFiVIiTP75eqmQFosW1d5NcnwH55Ddb
OnG2dJVBcZp/kp5Sw2LJ3MhVJ3MhBEFhGnoGIaIQUyfYerBhwc1ffDnOv8fULAuO4+FZxj7FW6od
/Bd6i6sfZNZWrHFiVkDflkSi4r+55IvpbIl2Cw9G1vNyJN61MEtPcNLGIdI/GYZN7k1wSmXzdI4H
WS/h8auhRf8lJ5e0pL2UDmGutHgRqnF/YzFzXU511F9Og4IwNk6ps1hW6DTKgkV9fOHcBpvDjw/w
SJ/CXR+0Z+C03Us3zf9BR3OXuGEeShL8ELe/lMZoWk2oyb5ek1kK6Y37cCXo55qQDbVsN1SUVlvo
Y7KMiD4hlN8png4XijWr1HlmHUsaWJrYpUb/f4WO/BGRRjDyovLLqlyYOF/WrRr0o10ORWWME6jM
mcuYlU7HmrlJbXm16k7nDg1iM0b2T2+BJPnCPD1PZSX4hn0h9VmjZDp5kt1HBV0usNsYfwEp/6tD
255T1oN+/8a332bAN8alLj7lWQToqlrExF0iT9Bjaiu+8Ji3SLqvBnYMVC53L4l8vfmkrSrxfy6h
wtJguv9UjkYnY7KwwxLCZjhtI0n8CCQnISln1JBDwo+ndgNlzNhoTa9yZpgjcJ7YuOUd/53BJtmV
MIawP6BdDE5ARXhdZ7BSLCuVqonfRNlO5QRJjzlBat7iH7sjfAipKKm59UDWydo7IBLbcCRrOUlw
UYxSR0cvI5jUH5qNVnza+BYI+ILQTEt18HwKsczMamy+bS9Q25MCYSvEkanOmJtQGzuziF7kqrYq
EBX0k6g6U41wqi7yGy2wCZkBep+CBVFQbQk/G2gAZ66c/LhPLme1fhe4/ZADdgqrka6c9un+/qV6
MGCYhgCl2eKFNqnLqdH26SrTECzggUIG4d2dJz3kj9SX0tuDtf9/ArriALslDUJ9pPBs+EX5v0WX
VSRe0QBWRqbEorLH9gnsS7RYx0vofJ1F4t+A/b57sopGHzqET7jAqOwaHCjE7tqwb7KqQnxiZeo8
jf6Yhf2wLIINoquJGl2Lo6PSkEj88KA+S6YaCCKLeYQwczc941E2s2Ev1rbFLWW7gJVz0zYA29OE
kFZXA5e8fgGGmLHvtmxuQ3hOXrjeXSitGIInHl9mRAtZhT8iKJzgi770F+VniR5UIEbFMTc/2bSy
Y1q5wUd7NuShDdAyBuGVQq5NS3WAAr0rG6pSjvvu5Ez3rIWeiNgVcvrOhVbBptHQLenRc01EMPGy
a0AQGlb4UQK0C1o4l2gWuUziVKmSTosc3sNToTugNbNJze/eOuMa/7z+NVdgkSMgMjUj6qvhII2H
vm1kf1OnzrXrGGBIaJqOR0xpEmfDgrrmQZb8dOPHKfdSySU5YHjGtAATBUMm/o02yRN29828q8g+
fNCzJ7FoXhmSn0N6RUUlrT7Nijc8H8FSLMkPqqeza0g9PIiUFmI8CbDfbkMo68v/ceCwoPoo3RBM
oCON4po22zQ/KMFU717JoxJYviShSZS0R9KNKeGEwNaGKuP6ZMGRRJRZCt0vylJCwPQXUBjZ9f2o
w+5Nb13zaf2WqSlSWAVFk/Z5Qz5aKChis1Ls9pUYvuKgb/FuojcmCYA/of8h/i5BHpmY6rB5TFPu
ZxE5mb/bCwTDNuckAUhOvNx+ntVJTJLBtjz4pW7SGb7hRa5Yynz0yCouhnRLlC4Fj8K1+JC6pnTm
hxWjNdJ/mEjPGRBBgmqVhsEkldWQLYholK2jiEoUIjCKAeXwfTSFMNnQaNfQsm+fUiya1r5g4VeN
+/Or1JScCp42uauO9tEuX4264OtZ+f8allx51Hp7CseZ4sRLmQf9sq+OSl9121zh1Jd9P/iJl5lC
j1hL1sQotEb+53fPTbQYaXorjsGsSnH+10alKzR4YDbAy7gADm8tlFqxDHwwLW5qaIk/S3LovKr5
vmbRJ6kXfWPcCYY7wJo9YpMDKZRW2t0Wo0mZHeh9V8RJWuzWu1e/to5gPQjA56OtsIN/5KgbgSPh
hBD1kK9zW01iseug+roX3C2pWV0YeKWAov0udBovQxr+v8JMtxL7s2got9lK32RU+ELFpPuSS4FV
BxYWn1omY3r4gqe/KzDhvWoLg+ehQFVGQ6cIqfueiKqwLMG9M65pN04EDCYQggii09GSYIO6ZAdV
hUx+LM9h+1gdQtz64c461d6L4FJfvuDmOWaECJWELbkVS6VneHc7Mjwyl8azxveJDhcQVPSb/Gle
OeerC+NTJ/KhYY3CKdGwfLO9iO6UVJOuwHll9Un/V/lAlAzDDiJjr3rWOquqr+83xyNTOZMGbrCB
DdE+7aIN0Ude9jo2cHYPlzZqpojtbIsdVSm+m+nIA/p8cFVdMoQ1951B4SQQyVueRWv8MDRfpJNr
TckJemy09hQ0u/6VrAY6cev+sKwNJpUs6iQhZpdBE+HagmTGfpTFpwhBys13QoS6tCElCTVqVj0C
nAjJ9APouX6p/5RHWsooXmzPm2KowaCHKCbVfB6a3UCUlyqPs2DCDqJrQ6yHTWposcNJm9r79U38
0/dYCSqVrjAtaVHJWf2dvCNU8xo2ye3yetJo7GX5DdJvHunqHJD6HeOijQetYIAdFMRxoOEMaLpy
/VgMRSVASnH9m4HNCJMOJadSFJixEVnLzCAOWZHg02N+ALq8l+Tcgg0hXtBvHMkS2ib2WowjcFqZ
m50KjDJ94auBaSoyMr2E6N+slpOsRT1e1Zt9S6gtQHMH+PE35Psk8Jv7MeuD0wADWdZIkiCTdGUC
7W3Xbx1kLkZqyBy/YCysGtS7T+y3HlP2TV/aXl57HxK36X4lojIBKGPKUUDzlcGpJRvsb8Ttqo82
04JIRAVUpaaW5X+aUev1twQVoKnx8fWeQ/uM2E/p8k52C6N8GqCekwjNyI9WMrokmNX1I90oKE1z
Ajz4gYqUgzzIa6+Q84rn2/4sHokpH7FOXhdJyXXxK/ltviWkc1BIQfI+bzPY+kOK8pFJKq3brN7d
VGI7jz0GUN7eULSNHv15yRvH5PWZusqHTU2B8j7Z5YLOPotUhx0kkZfA8hN/bUgLqmceKHJiBjEO
wZonyrmDnS9xmSC1anGjL/KMrj+TscUpbdNxq51ls1TmwsDG8worBNHWhccCi9kNhd7bnJ7YFXm2
Xk3goFHOnCjFetwWFa7ksGGOgp0iPseJWDhhlI2/rY+xGcp9SV/fAJgDSvhIXBILrwuH5Gd+2VML
STBN5jMNg8O+VP0tkUPmPF7lTrMsMqTHDGBgFOEgPr23/y+VX6jADqiZRIMh819Jm2gHy0lMOu4/
HXzzG1MAXEm6ZV0Zx4f2Anx+iydv/gt2/qygI1p9qfG8+1uFJ72KUYshRE9DNNBS6ahkXnJByxeD
h6D0VgCfM3ERafACO+dYwFPRMi1qg6/kEHM4mhLFvCgSzX6EbyVAl3E9TF29BNpe2iJzOVjsKcgK
E/ONBlxolhmgSuQNGmXPiuqXAzQM/E1hJX9M2zrlk3rjiZBiZdVZM+sx28CCnCowYKJy1CBUSrk7
h0/Dqgx9e0lAFH0g1trdzR5IROGVj17bT26p4rBZcdR24fx7fMdUnx0UM/2MooKauD15KSg5Uto9
E0u9k3xH7xOr+hjVu5aWiWxW/+wrR9rs6ktIvLx1QqOSwbQ0UF/VVyJ7kNiOaN0DdX02Fei6/rbd
stotD8/Hv8sSh/Due+Xmbhdd3U0x65nDmz6YJLbqO1sQWmda9FdIGV8kxJR3BlwnqFdx1D65rmFl
tBix3C3d5MMfKDDsb7AjUNMGPey78jPKVyek9TgsUpqOsDJunSaeZcU0RYcSCbYTWRWCr+c5Asd0
SqRfziaLNlZru6cJd88Ik/FRY9AxDTfL0ch6dFVpWx/l+Uo0ybEEZsG5+dJ4E2SFYQhzZXwuEr6F
QOstfmkDlmjwpfpEn3Nb/Kd9htZmCbyKUvybBPPaO5RZhGuZrsumxnyPICKC9AvsVMlGORAE1oJE
6OuUH8Sm0vBw9mcOVpi+WQhPLpN/eEqqkzutjrYacQX43hQDDt20RUaxuMs7qfgHJs2/67e5yOC9
TI5pdS4jTD18a3o2a4V3dfQ/q5hGWxYRwty5voSxFARcX+j6gOt0KZdpdGPJr4AGSrPIGMlyYAyQ
LrV1DC/x4CDlH8RPMSW6qRahd+lIB13YZtPtTJN7oTL/6Qzy+NX3EXsS76Fxsrxyd+X1o/EkGWXl
CU9q4UID0NkIGV9uST6bkggvFIJhMvm9wW40noSyNAlbwAgUKNLqZ2tiY+6/f8qWo7nKcp3MlCqG
55KR2zvMeptfRwqrfKbvvXE6E7th7ZymqcKFSn6C1ksBgF5pOAuY1r36ekENt4w6eLbJk/kxpMtr
2JMQCS8aSQTVK0rRzuIdRloEArYcCOeVtEPP4q6NVbg4u5WgRRBUqeE+SJBS89o/A0ugdsE+sk+o
c4mL10HId1/nB0VprJJSWNNfTwoXyZF73jTqLGcrZ5FGxiiI+lxMAn4ETWcxYfNE5DnE5CfC6Erp
lp1MOwMGFlvl/GxIY9KCyz60OqZuepDSTwq23eo7p3Mlbj9L4O/2k407rM0jjBgSj9TCImsrZitV
gGffjL20PyskSRiq0pXn1GJt7eByY/u9mywwiEFt0skLbhbfU1F4lEPenRZRxMTR2R3Quq3R2gQU
rPOq0JxWEGVhwMUawmD+e5/6MnYlaO6pSWr3Qff9gFl6glw5B8HCvNSw3aX4LhhH7E6SvoaqdAq9
qWKLl25tYrFVbuK8yvX4WaANfE2+F7PM4wyjRFJhEWlt/b5Rw1aGPQ6x0omANG3NixcZVPTNp1el
Yh4hlmLxVPw+DRdaiYVUBhWhpCujZydEGHvMtJe7jjZis6ReB50jl78rBLeM3hZ48VYrl5qrmfZL
qPcnx3XtcTC6tnjwwMVvM1i04mUQOnJUgQnmwbmwnCu9xnd4i/utRT8AX3C8P2vhOzehNqgHe4xc
HzkjUl/Yu06UPq56jvJqAH6SZYkfQkNFfrQgfDBfCIwYisqMbrN3N9MT80erOCbzMsK3nECQFECB
i0x1dk8L7yesHQSjtQhUuZcyBNZ/kdUylOjqtB9KwwvrY4SzGPaCUmS7mPkiLBWW5C/kS8rMpUzh
CjCg5hAgaoaNlwWcoJ2lp5UQ7RZmf9jKCexO0q1FEHgzqzZwH5EHayrdtoyB/olJo2nXJwFxLpPJ
wGJLiJ6yu9Z1qyHE2HXKMsd4DkhsX1qxF8sTAPHX129L7k2tBS07tpfHCWprXvXvmrOak82GXubA
iVkvP5wsBdcBiXzMshUOKKCoFpbGFFyPmqxF2Jo0YnFmyTRqN4Mw87rdwYyuldyquMb+1lAturGU
kZK1EMl+Qzdlnfw1cYwB0m0TF+ipsEdJa6livuvhvwLay11M0B8PGlHTJCoXzJXQEVHXcQkC5KLx
9rGFumLxHTaEzf0jzSMSCf/10U+kMRzeTNxnyOg52H5ddlRijmN61Lu+Oaj6dAb7KbXU9mVjPH4g
TXYwZ2fI9YqB/90tHLDIOwEVGolLMFFSWTv9LyQCAobahMUuwh6+j6Vuzx09hmweTTunqjxhjF3U
LJiVTBV6lYvGCUK34LJhTGVro2p27Pf3Y5wIvKmTLRVMKHnqNi/MOe/dleQpGZ5Zu8pMTrKC4t1S
r/c8cDm0jZ2tDJHapNiEpfngnTZL5TCZlDLZo6k5ZrcSOlJEvgjUEYP/r69V77z480S1Ssuj0z7l
qEueAVvkh6b92yNMOGk6Tv68BJwvSUA+PC0HQ6iBAehTk6yJkrBlhpNtCZSk+OJKd2XMGRIMajEm
kd3LZ6ayXuL5kB3Cne9rTCyw6F0juc2oMwUO+JQGoMNMelhq69rZkO3+8yzlGptjNfuNr9nxML+Q
dt2cM0vx2oDydDQXPVumEDbopE/Yh3+OgxhGk9M/IK0lkv/Sd+Rtijzsi7DHsAwSQYCx4HKQ2OVP
7nhPuV8suBQUA7wXYLtKyD9O0Nxr+GjJYgTwX0lrvxBXohoHjjT4jE6h1tGuEz0FcE7RO8gCoYD/
eY7fvS9l7a2wbyIl/rI5hEUY0rJran0FQO4xhgC2+bSL/UxNprzs79acbpnBD+IojfalOBVrmrOB
FFriOogSQE3b4aEXU3Il2JQ4XHNQy1DP6Yzdp6kW6y86tpmZh8LT5Fg4DrlSHrvvWaSdaCTCQStu
u3uxSVoZELDXPI9YfUuBFNEdowA1pvSEiWhEpufCzC25Rk4wz7Xjo92BdYi8nWm7d1l9WU+ZkRyR
foYIFt12fv/KLfr6bs7zqt2M/B7/cSjFWOqa6OJ5fq5CCV3NnEYi/OjZUkc7HbAi5r2vzHZtXC8q
oU+Z93ky90xtzwod1c3T/RLiC5fLxrhXTIch1DAl9XHofNKlUTMVgxjFFxXfW1quRtAxL4AljwJx
U85fw/bP1kFpqzpsa2CCu12tS8uu5WGgniZUUX40PBIibJybpfQr3Pf6zRSGWyLM7EkfSm5aFIpl
srWhFEX3XHz+hQhcr9aFTxj+wdO5HZrZg2PJFoUPHjMLrFmYonEAyQkMDfmltG8/dKJNF1XboNAn
8svK2BTtaB/fMjM20sQhw0VGnUZRrxg4WJT0if+Wa6fk/xpleoGgKapKnFbrmu9u1xnwHrOUYvQP
oXysUUs0AsgMHPEqFCTxnpXyXRf/+wjZrtTzSSxdeZS+eza3CviL4mRwMqFKnRL4JAQ+5Uv+JAfh
MN5aFojEViP85YXXjiOQ1O0CMpgbJnRZyhvewTq13QDdZUfe8wZxBDuWYkBjzYcDnW6XucwqMRBc
SXlxs161eXlxWjxbb4ACpo+b6eLuqPW5VNjl530U/zEuHAN5/EchVz0aj7qFZR8Re5tiA8T2UBiM
Nt5WQ2AgHRKv6B6vNL7d8SDYl3nhz7QigTDAxdWLV5lQFFXF3X+H/tbdjKXUkr/JUelEVWnE5BXy
7ZrQ8pzICRsQLceSC9WDtY9RmW/N6g3vTq1lejmMJ4xqlchp76L90uVRX6+GzhtkzD3NRj+hcR4C
d1ONHMaYD82+vugTwrcNeie08YL98d3pq9D1+Ub2T+/JnzJfvOasYps0wYXI8gTbEUab/BnprSuk
kSQUsITB/f8qiAc19iCJM/QKC5hEQ8wSQhtq8HSGNy0PgIoKEwC+nicG6l90YTgbVaKE6Oqd6fv/
1g2dLJqvO24Zy9XafwlvnyAlAo9DziYfGOJo+uVquyn5u1bD/NCaVL0e9WfU5Xxb9WsarvEuKqXn
dS2PsZtMuYwj8xt4pfV0Ql4StiKmc4e+X6WAOvMTQg0/nsp68/T8GwRU/Qcx39upG7S56RdISSvI
8BgjXIq9hrX+12FvX4cy2W9S1rcMObGoOrLPP8ymu0wDvCN4U7JvfM8jlK7Zi84vk7pkAKM5GGd9
3eXdHc4pPkEhGmOD987SqaWUztUNAKkdOutl6q6pbQD/N5AMDV9PhhsfhBUXWtf76sNG0HePRsLE
z4T9UHoA6CPM70zi8gxDN/zUPvU9BsSyK48C7d3W3ANzDcC8aZfLK0F52PYKE8mhBKo8pRvHz/Bs
6086ilFpSRxF53hUw+sybn3Bd535MeglW4oSX35/vi21dVkDr5Yka8oTcTmBPcI0wqsHUveFtSAB
DH6HzPlJwVIJ4lN5SOBZPPB032AomIkZYg2Xw9SBG91isjSKLxzRTRSqaFFk+4i+6DaQNKPLe56F
76iCtWL4EVXMDVL4mcopDpq+65a0yFFSFvD8KKSBLQg/xAcrrrYVPdYSbedTA3thOXYgDvzFN/eI
3VopQ5mxqVlw/FZhXazKTlBMDpPa/AIhCPiNeznIY/26ErtswM6SehDWtgycfXW7td1SK+FLumkx
1Oe46jQ5/Rs9+C+nCN4BdnJUqbiuvm1kTfp/Euvc5YH4UbUHTQHhedhZoXHmFPU+bg9PMN0QKAKc
0E1LYXWCRO/4fGzuspcffPH9hwHexjHRSOUowVPu1oBKYDohxGbnaM3L/2F5WyOjD1ZSV0qUSmTL
MLNntSgvj7oP1+wzAK+yrNPTNwhtzRmJpDCy7roZBwVvpVk2QoJmR1Hy7QBPKFJLRyRhdFZN+FoQ
TcaGRZHIM21Eow0GeA1fszzrCUTtTqXj7DWHenvfRtG7H0koxNyVJd8DrI2HgbWRtcs2AAFaMQNx
wVXFDUhCXfuG4CtzMeoHwAFfkOOerdlH4FVXpe4GRJmnli+st5qCJW6sucDzOcEMUZJxr6VK45w2
u9UgcQbtKAzcFvNQKtVawdW10tQzLZaBvfBRVTTPBHXm8mc6odkoK01K3UNH/BlncVRtUfUgH2+u
ABReL2KVyPfYZXcnQfGn5pMA3j2By80tBd7eCBUy9NImWbzoVZww7QsfgZN/NJz+QwTjdYLSnHmD
U9bXMzsZNfyf5tlN7VBt77/2t45HhjKbZzqKVyWlVRhDKE8aA+JysRqAaqhBCg84xEHRaBC8kYKS
G7w8idbqwEIMpIvaUmrhABH2K5IAMpMQ9u+CRlaVuyJVNthAiM66d7+u3euzwk8ilDtN0aZt/Yn7
hheSnbZPsALghsw5t6AHWwIaN/6BGsTsG1ggtdaeakLupxCjAqIhG4IJZa5Pu/l8nsvBvCfvS1+m
1UcuzqYJ5UKm2dv7zifxwuld4JRhOMx2n/ixe8IXiGAFRk0xYWtYaMdQllHukw8zF13Hfn/VSu57
a2d7B8RWnHj9BvTyuE9990neYyRfzpUbW0grYQ6TWQwqf5JmbS8c9VWACH3jH3+pTJt+Ndio4l+N
yGX2Byte1ZJmbO4I8Lz/MckoPidsBr+e5O3nMd2jydAdB/Ta5JmbEmTlPTJK7OKLGf/GwAwwck04
+4YRb4aMf2FpHOnHaa0O7iL58aStTxKezHSw1FaFAvnv8Sm0pXxoNiA3nAYRga0YrvOjv//z6eBk
ZF+myNyohX4OiDUMJK3QNhxckjVCE3GADBC6OUejowox0a4XrP37ExTKhikipwEW8rbpMt+0pwQQ
vvxkbTmJwY35j6QpZHGevsKNRw7dcxOVsgmC2rr/J9j4l2XIHgG/1Efg3eojq1FfidQF2HtKpnBb
Nwfu4xuPPgx+ZARprWv9V1NTOTRWCZj7UEXL2SlioA0Vvjrv/gy/ozSoHOQ4Fn05COoizGwfT3pc
iGuP9RNrFHb6Si+yTYDYFa6YFI55a8VAAS27aa/D0Z8NZMbwBkc/nd26cAFSfjDz4BZOoGb1LS5D
olB7ppHAWu05MgAVLUtXVlNbvV89LfomZHyg+UDO9omHGmr+SkJCwmA1I6ns1bOMJ7arzZrIk1jk
L245adAJMXCPakBQUonJhTD2m53yffIymGVfyiHRK7SkrJNn8wahaw4ZKNrSlw6vUqv8MQ2SlODf
MqXSeCYgci5lp6UIasO7artHW7/luD2hZpWK34gH4FTgT7mBBf/YCrexadIoKWlCDP4n/+8W8n7q
TVEsOJsZkCzgitTmDc5LMpMKPkTrWitlqDS8VZPC4Lx1v6zEYLivbNGxBO/HuKPs2WYLQTuw/PA2
6J/uLW96txSLa3k0OhLA0syU+cADLv4rByOKZcErYmXVVRSfo8Bt+/XxPTSsDOcFNFNEzTsOqat9
og5fnH7bC/d3LB7tFm2me/OKvtDgMKC43wLvFVnRoQe47qgrYZ1UO+CkNtNHZKsr2QLFzqgrJfZx
vWeXoRaESyvoIiWzzp3xz+4v/sGfVNo3oiKohJk+12KmMYRm+KpgD6JNYSfmKPex9FryU26yz/kZ
G0zC+W4G8mdvyAsoWxEvRXc0ozxW8UmbflFbCHDSpPKSoOAcrf0MJ0KXE8YTiYSZnlDTl6CJ4njs
u4V1sDmEqGpzFgZDToL3xM34Y7sKXflc7ckE11xNC50aEAVk/qOkITCVtM8LOGwfXz0zVWKMAX9r
Dq6U8BNH5+4pwsyqXMqfMWGjHLkv9A4cMxoBXYgHM8YBCn1YEWuAEWHOMcAgpH0EScxLhB3uWdWq
Z0yJ3NRGg5X8hvM9gXT3Jrndmj6UXKwOOMwFMtOXbv6li3V1FIhs/sHUPfLubnHCiBuat3KZiSmK
D9kPJdwK1aZYtBuyRoiV7Z9PkJs7uzQv/14WBx1evNGQ2AIddev1HFAWKuOxwyMe9RmkXM5ZuTua
8Sd9yO1PoHoVPBwBKzWZfoT2lfA4V6ApjJ0Qk2JGg58KlSwttbIbmEU+EXOcxeZkVparndjwBrVU
tLAX80vY/8OFO0Ed4tKQO4cfZZASyPgbvpoyOrVSd4F/jLiJSB80rLIVmJ6Wj1iZq0wC0aG+CWSg
44CiQ0ZmRQ+Dw/wkDdn0F8T/6L72YB504jETJAfdkrxJa45ySzU+NQ69H2+6k3ExyeWRbmvFNPDi
K4PlvYqBc+oG28qEz7sd6TGUd5w4fuIiAvUh+F0PW/gSYt1CCWUXta+6Tk+wnDd9dJY6tYwvXIj5
oC/wwUc91yM7vTVMrzroY32nUSymhjYG8Qtj6gr7A/hDs/qSz9s/xnOgibnOtvaxXLsCfIjYrgRB
2WmDYC8vG6nHq71K3TbiTXyITRxno+mLkyGAFBB0+/RPLJLBao510wAN6mhInVFxxxhm9MwVYQvS
zIFSh6BJk+DtM8tWM0S9KxlvEKkixMF9UcabQhmooVaFG1CzfQWG0UmPfa6aelHxM3LqGUlo1wX5
uGpTSgk2dg7zPhZbQCR+MvLhOQHc3e1v8kW4+0xj4SkKsTOfEm5ZScGlBPsMM8NnCmwMuRC7Late
3sOEdWKAh61pVQoHeSsCh53gLz6gWkl4wbGmusJ6oROcuCFkeK67lgg4t5yQlMJ4onvWBx3Ti/zq
oFYP0LHmCWPRclLZ9kCwIGYDMU+LcyZCB2L3OP2e4KtC+3djKQhOuCFOWg9eYWGbaYlu8HgGeU9X
0cc0p93mRALobNwjm87YWnz1Or9xkksflBaDzTkaNL6O/ayg9mJihx0OQyvc+mNNievZJ73dqHXK
/DaYStcvtovs9bsitFQGgFAkZcQkOv/uDA2+WUir+JCXldPQOze2/myiqxQndkd+pTs7QUIdnmkl
/JkEHMbY7PFfzcgzo1fgDL83Q+d9SA588h0+Pw9Qe0cwnwL2eTRyLMrQ1pQt+aLcL3HXwI33+R8U
NRBKCWYLsEpuFUO8qSShRzxdWrvT07CGtDpqq2Xy8G66ZbiqlOEqYtcV9PcUojL7HsnlHJILJ7mH
gi9ZPl7R7oG652HTmwm4jvXqbSxq5xuOTrKHgLtr4RLoJMTH63PIUA3e318FPbvB2wxl7r6TBSd1
Gb3pyxrRg8DfEPm7lw19pZ3GMTU+9KA9DW3mUQDeQRePZp/ZF5SgON4Y5dOTKotrHMmnEnQCLKj3
gqfRcaeHJk2EXhYF901Ti3Anba5FiGNdWXe0Tnoi7nM64DjDYL0As4UaklNR6GcCiUQyd0nnj8uI
ySx1GKTvZl1NgQH+mf+99M4LjgBnZiI+4bLfNYEYs79kdvlpUPpwu+MCU58b3Hq0w6/AdWVFBW2u
UMycBapD+srHbfSTDM48jVg6knVFEYciVnhJh8h1BQbLF9jfHx1nPQXd/TRS1LXuPAqsiewClgxb
SJjBrYFll694XWTCkCo8Q/RqXRqe7XZsznSRCrJ327u4I5E0ee0OfHDYVXxiQRl7/d9H5Ar4Js3R
ThqvNpaosQ+RZorw4NC475/P7a58C+URaZPJkiBSgvCuw3q8rCHrtO2SEKN010a5GLDsJqyluf+D
8bfHcoIl8B32FoHT7peJx12FXdd/dnt37/QIIaf+q6NX9tF3egYurr45MdNwb18gUsuRIFtU6qpU
2nqGIt38UVQEO9KHBxvKHeMOrx5RKtigA++ipfbjwrVv87iptQajjvbSRGF4ur1N4SNw20AJfZt+
lDZEIvSMieqxjM233dN//KdLgjRaR9n/ici11THiwzoqyIYPKdqPShFo0+PHqUvawEoXtIwC4F3d
jpPeLaRaqRn8JPJu9HbPMRJrlER0RImVuso/4wlXMM4/48sSXnwF17rJhJxS6XMwr8Jf71oOj2y/
t1O210h4K9f9rNa0GkTBQHf/uOzhNKdr/LZrsaoJgtsQsiA3xzDO0csQkUB8xFiHRDI/HfZN+h7Z
sgEpU1cayD7tbETS0IZAVcmz5LBjTQ4HPoslnDmxOBEMHDcMlxW9nueO0PyHZMffSGK195wyqUtT
NX6qkLDkPc2UXBnMTO0AeUFi5I522DxG+aeVrnbglMpAl2PAbri7Ke7Eyjf14KHCViSC8ivVq/hO
ZhElu2v8wEHnx1IyyCsDCt5eJYN8GcMsi2cyHDNfztPahDIJm28n1ticlV50oJTjxgxLIfAqfrd/
p1G8tousYqQumNzatm4T6qHySUkNGP6i4+GClq0MzTIH0bsdawszgPlHfAZ16G3pgC8xXr+ymEOI
mhpRN+29llfvJ2NIxjJrVq36TvNUq5Y7ukXtooFB2Ch+PWwjsNDCZAbwmnJUp9n+TF3BoI6xBQqH
pW77RMhYw3gnrAZiWIVFOS74+p6SV9P0Bg69hZCOPLhpTBNWCFkN8KrfuxPH/7cIEXOmpKte2CtF
hgsVy5FIxZK6PaaPh290lM6pw57fAbVKUTlzP8+sBLkYc+2Jnt7Sf7iGvrxUfUt/uK1/WkgXpyeh
+W80eC9NArSLxIKc7GrL8GXXDlZXbm2UWbV/5Pl+LjsRlvf5EhVnRRO8uRWfXpP53XqXxgliw1mP
n3joOQ6d9E7r9nf5fF2Z8Uz5TV7mTZ/yWwqQ2y46nVnfQWef5Ou7QJUjwt6OBJ/CtDpa9mrfs2jy
adWa1JcjIU2i+LdHnJbVGvkI6ju1vJnjOPe3duIFacph3qyEOyx4/XfCkGnWlzc3VxiYds2ADMEf
Cv1ER5H0rQqvdDf4e6e48wJD5+rMJ5tuYAMtjVB9LoV8bBhdJ3rR98toaHSiX6RNnCs5QURsTEwW
h+qkFTzDmMOYXiEHUO8KgDo8LJQEp2/kc2jCqaq/n5GJ54j6KEiURiu1qw0eKyQQ5WsrZMpurosS
KhNsFyI7TbEZ4oMMbRpXxjZ4Dtkwfx8fprJqPvvKie8nnWjPYTYSJ1ZxeSKHJbMMUtVQ/4Fe02ph
7eDps0fbvrYT/vVnOUXhwbfdzpsnjcSq86QSZWWfL5z6wDflsbTds7TRBwXqHkaMH2Wr1z9fmsIb
3EK6D8lmkolYPrQaUlpzckO6Z+rY+1R7REm+ri3OxX86ac88X4yaVDfDHPoHUdp48l6EHtAp6bvh
s1AbY6rqp2HqavV+smag5kIBK/2SkRT4tosrvCxPsFtO7qoVVOFb8enDFk6zhHT4sDQinrg+SC5K
LetAeeDQGTLNb9irPgVGwNqdfJNI47ECRkySFRzN5rq3N89XEdhVI3x9ZwRkyfX/z/i8eHMybYqx
WjiXpYkxb2WI5H5NTwGoMeva30dObxJb/iUR8Mc/ipBPGNPmWNBxjbl9ckX1mxceBfUx8eLiBtg4
EiyWEGTXGw+eyaGEYbKT06LxnpSKZqHArDH6Pk0c0bReESfnyIASKbeOzwLPehJCMhgh2C162U7a
sL/G1AmBeKzWWJI8seKyIE1CWOsOqm+koaWVwfYKD1UbMnzdfa/+hnRXxAHPq8jrlYWmeSXquqT7
0oue8Uw3NwumcpZDDH6hLkcp57u3c4CiFIc9UKECWMLZa/QPvgoPpEx0vj94gUZ74tuxEB9MbP4O
KGh52rUatTcf7mtLN5hcthWfHV29fBQ+W8cbs+8VMf7gi4+fO6E8xcUFmuLSqe6D+pHoLg2GP2A6
H+WX9ehFJwOwJTuPMPTM9KN188/f8HGYW8TuvbUJJhlJ817fGA5m3jfFriWd18gGJcB9jkk5jom2
BO0PAMkyPlbY0z8Aydy9nO3hne8Wlyx8GWv4JvhkTsuwskygIj2g8Jb331FO4u/HoqM9kef66YZv
13GElaSyoGocH+Oj4SpIwD+eC7Mqi5+ZbAUEbBF0SyOkQCv4TEF2bC7K9LXjhGYRBnJdr6c0KYSi
S528WTpv2LhwiyLpCtFBZeqCMGpUXkZnh1voH38OM2d+hXcFiDjmAgaTMFoX1kaKxdwXbxfOxS2I
bemcCY7FQLgKPjhwpRdT2gGJkwttAiU9/oGOzQsJEV1LZM6VkkONm5jL/0o1xuQBqasDUzhZlw4T
5xI45DcgL3xCOx1XfP6KGA+RT1UHvWF+y840NaoWZDbWwTOriRESRzFmZBMiEZg5iU3J+0VB/Cor
F88uqOZYreQumHMK6v2Ua8s15IlB0S+xkVwFWECi8ydsWxdiVjl8sF+vxX2cCTXzZ1dlM0oW/Hrf
sjWC48OwygoYk/wjK9gt0o1tYwkLvDWx7SAE3hWHXYe7BgunXXnvRCcPw+2HRCK9cbwWUiM5DgO2
srxjK+3YUMlIGl2KCHo7gU4GPBzyVeTbBrugUIxkSdwKjDUbUe+TkM3uYikvWEGGrorxod45HrJk
/3EmocDJ7MjxQvEAYfY3N/dNtJfZT91TqQiH+GNW0SyuvP7AOs0AF+DOcZxSnrmUEEE+togiEuZI
occ0QjgMuZk+wCTy3ARFe0WLbW2YXK6JgWvfsErGXy4pfI2SHVp2+27hbMdng9fhUgCqd52GGTM4
T9wwgj3gK3krW4Y8xpIDNmMUugfgbtYABqLK5wPw9NPdHhdzez15QfvXBBihuphWQ7+UGkSI+jUK
+w9HLKd0crZ9/JtZkZTXzr1zR9Fk8JgV38PPQvlL/MQvQCbAu8iYNTwo78zeCGKJJ/krUCWdySRi
OoPDzOOw4LUKKaNYMW5AIqU4Dpdn6OZOOZk15NxoxPIp4fh47uj36Oxp1KUCMGkjizuW1OfatYIv
XPmRHcp8AOGIk2U2QjX6DfhnyI/0oruZ8E37OLSFtACk5zlzW0lxKf1vX8k69g04YJemdN/OeEDy
r9GCNaAgZdxkJ56u3W7xTtXkmk4YqZ4sXgnt/BMczaT9gK/g9J2y6a/lrA49J4KM7EdbOq9tZlPY
PNVABK7u8VoJYj7tF//nPvpovG8vikaUno3AbLbjSRplWzKOoq/EbtOamjr0H4brIm5bcqMAhns/
PbZfCKD9J3brNzRX6pbu1tBLVooVJ0y82U7ODFdGNe6XO93zVQRyBKX3TyfJi1HbWxvweecvyYhq
5xzsy44BaYVrBbE6pwbSLAwImD3enQZDyHlaKYeBUngN9SJ84xCaGNuAKvTuqWfuQ0UdV9TzKx26
JPkcGRQq1oclUvl9i5EHfER6OWTVdeikR9HKMuPLvZP5vOQnInx2GNjiaixR4QlvzSWI1ZkQw/Jx
5KmiWI9uT486sIzI1hvmkyobc0+CGS+G71YlPaI3q59MfMxirjwj+S3DcM5dKqgKsMDIzCxuzotJ
FMkC5TziCeKetaepcX6wplpIWKED166V187i8cRCyRYDFDG3ha73+3SqApPhWXcn3RucvTgvstWE
NGxy64+rHWLiO/lr9CJB6KqK17EHWglgpIRLH+2oVYs7XPw8v+TBsUF+vxiSEocIMF5DbsDBbo7J
oSf3R04yUk11OpnLUuhFlrqJVcRl85TkFTeThjRGw7dksQNUssZ8en0ucE52f/86jV+C8Uwoh8EZ
+PUXJ+yuvsfEM+vIypLdJfER9+kdgfSK2K9uApaIK9mJGqXseL4Qx/enifgALj7nPaVAdfKFuHau
XeNC8AYywarPGKFwj0BodqWfTbf5P8Yy38CWgiefpfTJQN4ruXKKmsKZ8I/PSpQmqAvTcT8SOdQF
FHg7w7gF7Ka6s+5g+dvNw4CPhdWRuO/ZCCKVPtOUSmErmaMcd3Vv/acq7vQ7bh8wMJRjRWenZIP0
Q8VZXG23a0Mf6cqg6Je6BiPmC2V3NMEzYy51ALoQVd1dbLnnI6Lpqcu9j6q0DlFrazXOtdW9gegD
dkCEfraOhF3AA22OoXR0RPqmi3+hT5qE6Cqq317+7y3iyEmDlwxuTr9JlbLl1rxwxlu35jHQgCZD
fXmW6Rmuc65HYPUcUiGDzd5WRykWEw5sBv7C4l6WSY4qYGX4e+CWb/XGKAuNfGsqWRuADDOeW1TZ
daCYVM2wLzc/df5lu9csw77aCsc3Bm/3j8rCA4F4HJStDwRidF6zQcntuVYTR3pBVn/dEtxdB+uu
RIdtQNaAfnpWav53cmjaoaMEx71Xlce/tNh/1bE6cGU4Jwfdq9v0j2ebxz5H9V0acQlvdjs0Us2T
eioV33JA2mCJPg66BZYi4uvh6Ual6dbzji3QxsMA4d2WqFRZvdzxmBHXCuiQfwG7c3aND4zoNJiT
SRTPGv1YQx3zEyJIjliMpxflTGX6EAb6DaVy35On8FygnU4OSabFVghqH+lkf1shp/XPjO78Yak/
j+KvwoMVkVcHY04VnUO1BOnzk+43nEjzD/vr6p+2POoVFJhk8Smk9PI1Hny/hBbRSfw60op3kpS7
Bq7SHeoGVgo+F9R982GcQOEQvsxy95k7wrnf3EEJnkxkBDxe/URzD8AzM4JfG6fT4FP8aTx+J8d+
XseZhjdq6jw3gJUQgqpfRyyUPKXtp/mfLzgOdOq7t7abILnCN5WmFyDLrtE6gVGTrPoiE1cm90Zs
DH+gW2JkzwlSPaHfcVujcfBHEx+Mi8QVGOJ40gRN5bgIeu8hBuys3CF4DDIZuL4kap29FE1Yfz/6
Jy+kA44/jiyUsn1NRNZrEsyb8vaX/wVr/cef89D2RMXjuy+zMDrVmgJaVBzxmsfgU/9DpNyf86uu
yRdtT8NrUO7To82A7V2aBvzSWY8BWoJT+TuJgJ6j55Vf+ONKf4nIfOdANnKopbvlkndvRmDo03ik
AzjdH2NbFxpj9x+wNPeyYf4whrm0hOSjB37p1+H7vOFbWQDaiKGgYKu1+5wuKVPc3k0FSqITPxxN
lAtY50I9SoMSyLjvJ7yteHIZhapeqBJ0/iYTzraH50EOzqUuatS4iPfuyzd99osIxpRwD++C8qND
uXJUxHbZjbeQ2CdO+O7GKn0dNvjRu+pBlWyG6mJnIWX7+CaSiWzdbNb+2QOvsLURDShoJwdji6AS
9BiVO7czPF1vGD65kRTwJjUjHA6+Zu5SGEQNiihIMuU4cc5I3Y5KvSKs9MjIIzghVQHIhrqI1a+O
naxPChiZ/nNB4pB8LBt2jAqIB3Q8tpWQdIRly6dstldIS9n4TF2clMURMuzqyfVAoipAf8vw3Bgq
sRLeY9QozhDN/1IV3F2rRm8joQeDjq4c9YClZEqvJ+ATsobHO/lZZBS5wOIXQRTo/qzAqRG2hk5A
Acm+JhNMPM7P9jl+2cXzvNa3ao8Xrzaj/BbTWzBf+o0MO8QLmzLsSFCsvmWyEV9DjVW3lvbLtjV7
b7pwqlWRFtebrxljnVe0PJLrc5rdaUYKAxByoagGhtoyy1E+tpH0CMiQNOow+nu6ijct5VKSNhre
q3A0RDEKdh5Sc2eUUl7u6W4C5fLPeV7Ml4AzdnEnDHTxf6tjhM1JU+i/Lq8MIaY5uoGZ+2rbmipy
TaQ0QWOZM2ozbpdCZq2TXSCByd7zq6BIDCXNG3l1YalZcEnq/50Q1LyvWY523BmHfzm0yNmpn6Nu
sJf3RChsO8USkXh2StgtRb2Jm3RRf20S9dWOjh9WMc903mcO52ooT8IDExodwGTuED4M0YbRnzfN
ojOklZVKEJBC6ZVeZG2f5o1LID+cXjbzbjKtp3mlvlXima2shRQ7+8gxjqCwU/Hjls14XEE1NewM
8o3t4kjSfYXvlBqGXuVlPm+tsOavVCagFk9WiQauAzF4EsdbMDHNURf41I1GqTVUDhGgGfSAxwU9
Ws5llLm7GK67PgBinWmvJgNXgyBjYl4XFJ166w1cq6LTLC1KwLN+bpJbt4UVl73Ku6zZZdTjgicg
NhfO2eVg+v2o4Fj2XfzP24pvXConRKY/K1vImGKd/LhMUd4Bga0IhOyqjIZwgyRRXMORV8Q7nDa1
BwlbzI9umJlnUGODWafn0t30E2zqEOhs85w++SDzsDr7SeM3U4m9hY2umjjSDXH+SmGMlyyW6H7W
Hwy50iMYjuQqeifSyptF3MpO27qaOP+xudFAiacl/whuMCMkHpA9KOs+MGajh0yvIiBWCXaPlASZ
L/wJlLEiga4Ulc6d07DM7R7DOP1lej/xsiyflom2yXkNvAwEMOCsoqjjwpQY6Zjs6xXUkErueKNQ
e81cLMaIcDHCbmLyJAhtU5s8R331rTfHHANSKRglpPaTl4EtyFqp7D53PDK9cDKTOvmjLMOJfZa1
deSWsacBmoSYpgVpd8U/mRv2wkySS3gHSVeM+jEKal6O+F6F1CprWEodtX/MJkiRsSeEJDbGqzrs
YmsOHyKeRxbgss+/nUz6YOK1eaXL2WHcwpE4SE326Rr0twO1RC+62eQ3SiVz8fNYIuy9O/v3DR8x
7ZMODpBQ7McqgSq8hQbK2ajrnAUeNpRNsvAI1VC9qE9KUPZbQpJNzcu1fx+ZWdtgrkJr6dNXyD9I
fA5GLVykF18fVMldOeImWvaMwwelKEddyrnNpYfbstoebu3+0uPEJhUnbFUqXgXSuXHaDhdb1pki
hZRu71frZh2Htylgw862lqJmaMErziOQU+ORaTt/t57QCtYwOXbLit6I5JX45S+lOXTkXOkZ9Tm4
/34gflUFKSkze09e9BKoxHEIur22iK9bZWCK1617V/BzZE4y97qCE993wZ9/jGqpzvhvKyleNkpl
Ew/VnOqRaY+G6ZyixM0btaoWfUsbNZEhOtLMBuW/LJFJsYFRvoHxnNVUQAqcFKsIjkQQqei0Fjyp
ZWS5x8VGlyG1h8SI+X8kn0V382dHzJZSjq2/Gx+Ljyu8BvgJlweGh9suKWWyKySQE4Uq1RCqlqcg
YHt361MOCqZQYe3OxywIayw2elZImtrfj9pvQjt1a0aQncH4t+jaVfEqS5mVla9Lq7JCU5z+JM8M
KpEdZ5WL/2BRXWyeTlNg53Z20g7vkESWZNqLYJrnenwfRPO9n5dE6TbLs02QvUZ2sKesICC93I7S
t+hPKna0ivLNt5OX9fEIBkfuO05c2QswRXf1THMDpaVLDfU61F+5YoEazKFHCbjjAJZatDYAdVnE
3k95oskxyGOkAJVvuszafGfUvS/anastpL9mkkn84azYPwy15IDdoUdpYv13B5MloxTKXjhRU6Be
uCAd0O244qkLaHF/byunfKgXV8VyhUx8m463w9t7qDPU55Qq8ocRwBH9FA8yx6omWLDNoPOgcWA+
7jWO4e4YvbaJkMq/i1RuOLjG6PH3VVK6QCgPieXdaCmX/pJXbAiPsAPqJMZ6kvdKVwcuX3PT2gM6
x9K29HXrPQq6N0XqwfKRo6a/+CaUlEneBlW/sYSs5bNmsmpLF+XNNwn90yYylPSUzfo8jDIyQXdK
HbHIkWu6i2poHE+rqewmLX/xBmp4cXIhRmJ8cbdi6Iu4gVKDF4PT63DO3mVE1Stmk3gel+qsSuI2
xSuBCHEmYm4rcKAcEYpE3pBw4HRa3e7PzQ5+G2/whbECU5vu3QYl8wGdDASJRiJxFOHswCXhYhcC
U2DIYbikgiz5ilC+LIyJc+kFUrENdGWF7UrMkjAVbLPv9QBxS5/OuLCFyG2idFtIBxPSB1ofO98D
cB2kwV1jMfgj1Nw/NFyUGhF1I4fOJ52eDnCe7fNwog0erBtkq4UNcFLdtIlHNmSm8gJk9nWE+S9B
Cha5FLXAPbzGoFXmE+Qhe6SsT5gisf1vpQ2LvqBJzh8ZrgpWA1x5wj62wk2LZk0tP0TrJybMAbpr
Liy+7yp8AW/aTNof7eBaTGmRTTqUZF9OJIbsC3fmZcsbonlYJd6dDVctuMsJCdpTUfidIy2DClpP
qZ0JmkshdwRPtbpPFx4ZCZTc8MFGUjt9D0H4rTbOIb6+kH7Qdw48trT6W4C0vcCC2pnfw2OLsCXO
usFaNA3MQpgAYVDyGVqCoOgnhby/y9FD4pHwYi4s/4W8RU4E3YIHoQVKwdhN4VEHjY6SBcy6gzKO
NF55bqrLLnhM56UujTpbnuXgRJZDfEWaIPCKaxE3bokrcmKAUyTGWUYyLf2OLvGC8FxS8/j0+FmW
VkgCDWW7zHFe3hCgXsrah+ZCkjCHKhzNOIiDmcKiQWNoG9bugh5IvhLilsqNZgMGFXPSBkQrzVJZ
ped2cNXON90D63PQd2bJJ9SlVyylwr4chO7AoR3Jbp2fBeR/QAAqo+7Ca36S2WC1TC4SykCzjRZW
63Ne2T/wvkBX2FiNU2qxixjH3k4rXhw43OOmqrLX8SZi3WIUEMx2ba85NCmqxkWkUpPCAQYyVOwZ
lnAI+R+3p3JFo6r2qUDXW1ukC0t7foxcXMKxSoBRYk9yvWTaEXMnHSxi8hFZ5rRSZfMX29xQtcIs
jwcC6U+VKQkbOURThQ6ZySKQyuuGvXfc/pacLxG7Ygj66GP46li28xrmqCRsLWguGC+nLpHuOTvw
HX0XuIXbYgqOaoayMdm04fvGCTjxz2vyzmPlDOUz2cc0oW0we24IszDBTYhIAkVe+Meo10rmAX86
2yaMPAnAYioNA4gpwB1L3lGrZI/BGMnX4BUrUcidJa2VTFt1RUxjcUJLbW1tOSTaMOAjqJYaMoTp
GyeswrLsEr9e+ICTDqF66fv6T1C60AKJ98sS2uOj6tfbtI09Rwu5LCTe22gZ1cWDrFO9tgHh96zv
laaswlfWXS3gaEGvRvRd8CzQIDXVMtpzXLUnSxWEb26wVmPjDoHIENChfLazB5mLs9SG/k2j2JUw
G6OjPVxlWvIclhbFWkRBaMWpvXGMmBsdz0C7hKKIyeUCf2nhyFEwz8SfU7VEUWMmYiMSvLMCSknP
ndU+hzyY7AHHtb8gTbFX6GpqfqT9xadQho8TOsB3D7aRfwZUlAxqmvOU/fAzXEU26vKZbbPuNTzx
+2P2tpmD0cOj4VphJJ19k1grPYq2TLpHYuFB6cbcZBugg30jS+BBZ1fl7AMEy7Rbf8f0PazdEwz3
62vJqpuLBs9avk6DvVZS00fhoj6uQGtHDwNqfEi4WyhMBKlMT7CyWNuCHNj0x6M8JjSTy9hAgd4E
BPCqNEKSaghHe+XhlBd6zv/ssiPFT+YsjVWLLSXiewJ8fiDDktxTNlyg5x569EDwVONAmtKfvKco
RKfAvcLzZrCLiuzqvaSJKrkhD9bODDPVK0BAvjcvFxVqDec5ZaMiRFvyU787vrDN1ot5OXUsTrUG
q0BIngdBv3cqk5LJS+iptBNBmyZi47dP7nvVOmgpni9RXjYcBzMVVArHhKqa0dHcWwvXGolt89bo
zeTHMTdOzT0MdBKEIZKne0Tj3Myu0yDYc28SQoHDDSgrsDOewqZkqzaTBTyobiGysZbkQygxLK8c
QuvawWxiAuJyJArhlZXP0bBLl+t5SGN02rW6Vf7+yKtKmLbWLM4YjfG2LnB+ffZv1TcqIDo/dTDP
N7LcSkOlqhxXmtDstJ9wqtPK5vIgPB4EUP6JGux3aNiYhzL7B35CZdKIZzMzKBn5v1rjabhpk/19
VmricJgkSYtxOFMYX5fCK7menS32krAO8l2dDBES9uDIg7saPy9t6GJkIYr3RDAa8FCRUH82K+3t
Ruf0D2n268EXv6033gffhOJnisB+5Sem6RhGa+yOnwwHG2Y5AjSWGqV6wZf0iLkSHjolVKHYq7dC
g2hYSIiGyQhArLdb18cZ2ksamPjJNu6duOhg3Sw8Jn5cxwc1qOjROeOQn3MTGxnow8zOjrtT0YzV
CSrx8aHhHRdCGARCFlVLqY1V07U9Y8Qu5HHGaJVi7IIWa2SS8iqjOO0WDLVt3VauMbpxDYGTLpHN
sf93MTwW8ssKM49LkYuEC7Lt8RP+YiDse0i5XradGXtTR0sJPQu/PhaCufFBw9xAFnRb/aFTxOtn
bvZ/a+Ogc3lzMF5xWSSGOpxqfOgotLAzg1WYeu7emMPWI4qDx9wXer7S1d4JLdJsU14Ady3qXsXL
I8vG7HCMow6UljC3Snir7Tv6qgD2voe49luUpPvG8wJAsmBzndjDxfSOEoTC8Sx9bnqNtNS04RO7
etGRUYMNbDaFYEb32DFxxZV1smXpgx+2zfEIENl1nFp40MBSpqhO74fTS1hZDayZs+f6NyOWZw4D
sZLwz5mgFlpq6xOsWJkHfFsDg8t9C1sMAEiyOokZp5Ta8LavoExY1Ga3ppULkeT2m4obeJyWxPj0
gG63KFxKz9HomLJKKgxM325GRsdWTlSPK4/s0mekVatA0mf1R8aO/5jonnv5K9aZAkOKGOyfhlhD
GBtm3TDS4vxfAiA0Ilap/jpu44eDjK510lPCISdES/TSyiY199KEyq776kHPp1tD20h0WiHzKNzy
oujaVmngHHWq9jWAgLNs7Ob+2KUR6QaxVPkfdB/DLgINr9O4l90KU+ywg26fsvvOAk1B45GaKSIa
vkWK4KweADbQIictAFrSvvjbTZH0mOIGDPL3L8tyNMItDTnXQqLlMsiFUwk+mQt/KOSf03ekG/Bz
enTR14+/xx1hHzE7dUvIC15Q6Um8K0PQ8A76SK4CqHiVGZs53OKVfZVxYqC+YnlmaDSAKrnCrejK
SGMa4IlU+GPSOsuwt39M2BhQpKIY6Exi+7QC9vwsY3QNKM97NoorCrI7m+rWJGX0Nx5PGd9+oSWr
Xq8aY/SQ8mdi+J0+hfSVAPq03Gj3VWNyURFtCej47FGuONkBkXfitwjXwQ5q05+/2fNjTXFyA9y7
oVYF2nERZFgbDF8GLZ9t5Gupy9f+fevsdaMVqlZtS6OLczykJxYykT2vr5oKV900l4zrX7zGM+sx
9/QyrLRL6DvnxxwxYEIvMp78You27EW8XMM5hUGphEMWB+iVmTyLfTbXq4Uj+9SQHCj6aoLhklww
Ymfs5cEYlb3yqb0k1OFxvm0BsyaJGAccKwdQGDJq8fWxClemU714C8fDS9L+WdUM53TzOAUJPlmW
AYH/dBIdfmejf+VwRRuy8RvJjAKVzy2d11QZ1CHJ2/oK8ZJTbi+uBx0i1+3R39RCuaxBcj+lg9RX
xVB3Y89MDczaFh1wJRqthzjAlqogLxNylXYGDtci7O/Pz1XCMvmM9JN+VnGP+juLjrAqccqAc4bF
1UzCH/6nll8j94BT/PBumAFkqY6ihYJv6xGz/MWeUhLTh21OYE0WFFt/TfmYwF8FNqDYty8AwYQP
q1c7pWzI1ULzYAhD+418cy8oEszl5CeCCYU8hsYqIgPjoiQPbgfXGSqkfNtWxBxxWUiAgAbjoZUt
HzZK2AB7+TuWUnRWbkAI+2hsgRHYbbd8FqwAMLR/s4kkmr2h75pClSz0y5MlZtKesJrJrxe/JwJG
AeCILMUb048ACC9XQHdGJD9XWR6WWyon+87Xr7P8Maad6N8b7DEsGAk9irWIQ72PMQN3Kpy/c5Ea
9nz7ALd3zHq/6V97GcNJPMOUn7IgBz6/gAQbSe3pHZ/qDNVVq8Asm3E+uJTLMAs3NkNTbvMzrfc3
kXOB7Irmiw9DHQrOAomjNwJRVPOsC2Lo7IOC6GwyFSnoaBjxIOM8uqC5A5ZwMoXOLgpQ7h2ShKzr
zohWkzoqIcLQrl6DQCQK1+Lb5VLRjTr2Y40I7IYUtHcKihX4txUhcLlVFUaWlvqCIDtbD0wx2iki
ni2Ep6o/cu46Ogd7NGEK+DxA8M/+srpL8qr7cxVD9IfaENWmpugFhlCEBZvEGkbRbm/pgCEheVb9
4PADn8ITWSTej1OHkp/oBvBkIDAvTI/sufOZZzamdJzxOXf8HQ2TrRVqWLTaj3iJAY4BCfJH8OlI
cWtx2INoXzRA+Q+sOkAhqncWuvt+bHiM7/6UW76PZ6zqo8sUdL7dW1G70tJXnYCEl2z4H8RQiYjo
fLMf0UCjjucQzJ/QRk2mXvOy1gNkZQZ2TLoS6lwaa0qMLy294Nn9B5LINq4guEoOeZSccvu45qyU
9SMpx97Go2U4gn338gsx/McgsybPuBHjFYQuSk3PlYq9Xg5hWUYt09FpZoRKT1Yi5AdtG7btORSC
SWzVJgjcRo3Urx/XQvmfsXE0A6EP5dC1RZ1yDz5udgW1LAhMg6I32XOQdy8h0sfD7NXGp7S4gWLr
gGjLAeZsvaeTLqy6xouRteB/vkwUDS8LGj9a5cTtaGBxvXrnTlFUxfyHfTNpowYfi/mnBKAZnxwT
d8dXyAsnVWji0sa+36W7Y/D7TjLe3g1S8VZ/WO+kfMbWWLcULB6Bj+BIH0w9VuDApNcW6vMLa8PV
+JpRwzBSieuvlaqIi0TY+T49xpLca/o5qq3wK0hjZ7uxMawoqQ5wEUNn6fkR982/1Rd1VneDANeR
zks+Knm25AKEcI8Mx0H/P/GQlrFZfcMdzm6DWKAW9/IncgfxTKQZSLbdlHb4gBTpS1I1uz1njERb
O4TuzuKikL3qBwVd5wYdn2HoTfUv/1yjgI8q/vLtnkSLlQPDOE//Cd1yglUsAwOIfIB7OxVFOhej
qD0MUrvN8aA5b2JbMazuzLd7nmsWzhn58V3hHmPcAJ/YSZfn72jexfE3t0bnj8D0NtbSNBvShizT
j2D3HARXXhBqT0D/PMMVyzZ7RY0CHtaFQ/bv8Yb80+jaY8cqFF/d0K/rsA2OZnp+r7CEtzKOrafK
BQ/MLsXHBJJMkVMzUUkMYXCBBrP+C66wF+bi1wrU+yQR+28hmiA/HP89grf9ovOG2+BHN5cjMnIf
JWb/hJ1OHOuN6Am/xmiO+Rp3cgXUHAuCQPNOwtkXtrkQDxTc6TMWOMbUwgvUb5wXnuu18/wfSSIl
1NraZAkhbFbB1jcOegLkKLs8wyVcTSzU5yrokPTaNwVE5hk6sywtGER3qKz6bhbq50kwW4+ZSl3q
DOAkZZjt1zH2doRq3VGL6FY2vtypE2nIBw3EJupAgG2NiBxxztgJycUhcdODIGdlvt5XS3sBZ9Lx
pcVALM+QJsTTLvhNR4ZYqe/qaoML6fuOcrs+Yb5g6yIf7b3lg3b+DkPahveYZEpl/eLthcZwdfUy
ibgHtAU+bN+8lld26CxW0Mt2wcyndiQI4Ys8S68xJV/FshPjSOe8Luro9pkkM9USH1leuEIsYfNR
bx+QHYFWWRy+uDuYF6EEBhyxCghTsRUonRG451tU/OS+PaVh26dHuNhFn9fS7tfvNkVacXqoWdOc
fye3PKmAG3trwlr1O3bC58TjzGnQKUcuVqD3LeSprs/B6RUX1gGnc87kz7VTSsEvD2ZsE8zKwzqB
qBebLw6EJ8TYPfIAqC6pt7c84ODBSjg09RsyopF+gJ0hC5qFIF0HcD5cTa1i66QGtRaNME/Tw/K0
Wn/0wqVhrJC56p81xsP3cZdUg24CspMGN/JVLsoKjUeMc9SjvjXxBMwFRQYKtlcPxOqPiPBcoQYD
aYX2uahkpxyQOLRZOGa/6KMJ+VksjeBho1d7cUjR7omnSA/4mTvCIQdCzJu0xP9PgEKWMxJ3+fFd
bY8nbgeRslNzbRW2rJo7+XWbvLXHXOyXwTemdSJJXQ7pv3TB6lTTZOaUszT3VslOALVlxoTCrW59
cAw4KvEtvTrZFtxwcBOXYTVC7rSp4XEcG9SQNBDrIe2YBRXAkweeq8b+VIppXDZqrKHPll+jWX+B
0iYY/QE/ILC4EvXdAGAX2KOQL/BHCXvekVygtHB7KwKozy5dFGHik2Q6KIYbuMLfLAGQbbKmEEzX
fZLGBwCkjEc4j22CWnlkUB60uWNsrYf95ogtKLDvh9OU6wAyXfzBXGtAKcscd4PiedUDM2EpzCm+
WsJuK2z432CiLk/5HbgsYSNLlb5xjv40yxXsKAdRr9a9JCCiD6MIAFTWNJpGb3YEveq5vAr7un85
40MekuOM9t4ILH7x/W1n76f35Wy4QiAxPZ1UkuXBdrTU/6ArdoozziadWikLWrQmZvDEnUINdmyO
caeLmmdJ6mvKuy5SOQ6wJbWqGhS5h57e/C6Q+/eLRv50HXBh03UaPd8wg6jU6OoCct75DDlacOjb
aE8lnKr9w0NaCflMuMMPbwtXswiXhglXqQDaRB6ubuxLSaLbGOeH3Pd83AtfV6qBkWo3izND7nRR
gppF/6vporEETO/LI0wxe1ViZ/+991WWTPUUPDvPy2OySUmfZygQoxiVlNwf6GRVMjgBG4TC4L9J
C9jJfBmhdMlJ5N1+HGKilRpBlJArOwcpkpcW71CPDI+YDsALl5X7oc58iGnw1+Qq2KTjBCj3MVej
8RoHzDsHykYa6BEuKGmaxkNA8rfLo3jn21YCVCwxnu7QlbXtFkUL5jketyowTkhKNWOE3u3QGvxL
kQIm6PAmbjV+Z9ZKeGMIrM6LK/Y4qFmV8vHw4etBhLVsFeyPwV2T7rkj1AY7ltuf5xuYReC3Kk31
SfwmVRb74b+HYXw4ALeDYYN70BMb5c8hgWnm4Alpjyg6l8M5dBvUM2XPjmGFMMlq2KsXaSSfqFuW
ZHrAPXi8ncIDmhthy081jkBTmXmliZVwOosHhNe7jxEtNcRgrZqJRA524UVeRIc2fH5L+TLjOKg0
2kwLUXIZha3Ip7m+Bm+qNiaj4DpBMIvdC1kmKkUYB1siQ7frZykWwJU70RYrGQfOdF4dN/pgNU+d
rVXodTQup21vsmE1TOzYRPU/3SZZmBtGuxfMgopWcf1TeJ2CJsXWvuauKfpDZKcueHy0bWLsMLKn
xxAjTro3P3he2QrPV9krnBonYSG6wB6FjUa1JO0IVfkN1fZZZzoawycpGl8oyBqdXYyIYpjaVgvT
EiJz8X2c/TP+TjuHYeP+PtLmdSkprWclKiz7Y2US7aSnk7uyoee6FQLfrVWQedZVhgycSOvslD+3
2Lkkl1tYXjVGoMUbLdkyWoC/+I/M/4zx+t6ewoJvY0h/POV4vhNy4F9hYuE15Ui0qXHH+Jh3tn5a
WZdGU6KNfrszjr/BZ1kCYjk77xPNhKPprcFbFZywne259LcbltVDZZgN00K0TpfOZRFY+P49XFXg
+lap9Hdxx5ixM37Nwg7wPW8gZ7PKOhQDFpYWYo8WgInONynBqy+W7m34CIkUE9KwRFtBDHn/ohKZ
5G1cxhZsaOoKTCKiZT/Secs8ndJBnCMoKmb9tQDjsPlmvbjs+5nfK9utgUqTmHmos256mF+FlmPq
YFzCL4iLx3hXKplzmfDdQBwVLCepyOX6aUJ9CWQ4JWkktcalCCKaGtKbi8fgq12MjPS0mfNF3zs8
6ednh5GaszFB6Xf8sy8GAeN149VN0EYjQtIJjvaRsdLSPW8oI2WOzIW6zfEMGBzE4L/QeCNU+71q
08xTGVE2daqk/QKc/EywycE21pqMAb82P0rcWqm2HBW/bEqEUnoRImk2oaz5Vio6nIVr3BlOVM+j
ltMoXPesjECXI5Emq/pd+roD1Yh8lnK5VwXZ2Rv3z1NvOW/3gJtcmy+YsgLH3V75FdciOe07m81s
II4EbK0OriYfF4qtr917Tn1cMwNEUWrVWkMxk3HcsGlsgSjwbuKv7hn4CII/fcq3Zat1N5lR6SHR
mWuPuJ9pHYXOqEf9KHvLDmLBBM1+U1x+xa9EGYKsFb/PROdGIgzM9ziFgmjBkFbPJdlmlgOFdZrE
SXsMpWoL2k7gMOI5XVhnkRZ2uOUToiojZqO8H6jPO6okWtQi6lVyuiSS0RctIsDTOZ0eEEO0NXa5
70TFExcES1XT4zeyS/Egxc8sefdwpiy7Oi3QCkthgOLY/utcn1XwtDZpxh9s3ckwgs7r4d048tUi
Es5J0nMAiNX5o/3qj/WVbkaEmC0JIvY8Jm+d8fmWmX7giI74S2lWf79cqauD9mqIGqxCt7cm87vk
bB/wP5ySUgKAlb4/etYqSbCbrO3jzbFeBFTzTBicFE3dh2wiSJ0PzZhdpesYyPNS+Yae/LTGnuI8
7U19kVA809Qo5Vo96VDRQj9WvcsqoUUmK91DCDj+soon6ZGy85j8EjlsDmFFSxtGEKBL61sGWi1z
9gdZUK2aC0bK/3BW5VDyVm0uxK0+VPPwArUV28DyxkHCbYDNhN3euD3vpSPAugXZoQeCSok3S+uG
advMFMwhwKBV4byRoGaiW43FZusM+5hzT8u8HvHOTUW2fTjM7Chug9xd6jNBTpngG5YwXCj9m0gW
YSY9TMe1sBD8AZN28c+dcn88XPfDl1J0H5WocGPlz+PGLxAIaNlBh+vdN85STexW+RIoIXXE8uTN
KwCK/bdRWkmvfvxCopWFuW0N9D1NcOUbE0tTczWGwWswCO+Sf9TMXVEN+ns7RRAzuTp0lExSKUS2
WOIraW6eNJAmzFu4Sd7eFo3qrIS8wkI3cFbM3bcssEyDqmt3ADQMbEoILh553VEbclOFXb5rAyI7
qaW+v//E/BWHDfApQg4ROXbg8TvVTLocv8yXfN5icoeUPUu6Dn8IV08efjHMzKC+EVDbYG5Wl6dO
WuxNTn/rWEuoy9+T1xcvLquB6MLfv7jnwW5Jnqrk7GWNkWVqw0FdBxJdu1SSiJnc/qdVi1jsx7lE
cxour7dd3m8SrL+umPpf12re0O4txvqlUg0f7cC/qTzjstkKVV2LuFr2woKIqUHz9vSZW5KqtHz/
iuH8Ble8wM/Hbocx9+ybaCY/kQ6kkdIcdCnaLopLpXRuOV0U+0NlVWGm2rpkwtonk5BAGpFIsvc8
b4B6+CqU25Mj7Yv09cIV7Zu5qJJ1Px2URL8pfcvFEVOPSuwYi/Nsz5C1xrwHx41NjhvTivnCOFcX
+PPFpelylPsC0Djku2o/Dhf9O1XsGOAbRg95BmI7cHqAHMcvNbIV6Sb5h/HwmJU5sCbHJ+W2bW6h
VswQmDJBxz57Cm/WmeA2Z7l3DQi8e5qivkjw90n4hqMvSKF0Ek0IxW9lH+dHAqnpfZoFJ5FSlZcf
Z6vvU0kRKHTobNO1N/sGn/UYwR4afa4bt6He6vJFev8WTqUsgJYKqhwG64kY40wSzUDc0RMZl/9w
dEkTZBciqsqAqs+0rcD2ONCL9FD0wHzVT5PFI3pIYXiCAE89PySUoPM9kzjeAwg26UT5nSQqUYNG
Ck+ZmCmpqBzPm8c3kUdE+Ty9ywS24sRXyZjv6VmG9E+kTAXDlwUgcwrcD1tW66a1woNMuB7srZV2
Jx21q6GxWlQEsP7M4yPuObUwlLu/yVN3OICPmFclykd2kLw9tp60XFewxyejlv3t4s90sXF5Opa5
fa4qRHBTstC7rhdK0SzfwHyUIoLxeoUS8zFOf7ZSiHgJyF4bsoqmws3CvMdPdDf6/yep/vBq4BtP
Bf9c268I8+ahV8ZpEaEMU6Pb3jpKh4t7qNrXqUNDXwoKswNEeq3JpdkiEfbqmqnty4Kei6JLsttj
UncoNR0TJ2D4e+471Np6pUpjIqqbjUlgGJFBatmftt0nO+TePowPCRZkT6ZKbztMFqavKzHGJb4S
fLB2QFX1ESbb2L/gV0mlypmjUTBGpDM1rDWhRrttQNkKRLhyg91PHD45FcjZQRn7cLFY6ioRCphN
GR8ww1CbgXsp0kXx3tBgt8HnIwb3HdeUw+48MGHq7nImqS21Ycv0ydsDqzjN/5bmMO045+36v4hg
zIoBduJKfB3xG5WQj9fP3yX9HMxQKzvwe9lX9OSmsEhHGrS13OG+82KDqxnIqU+jQ9LeP0nEzh+9
WTbSAkCdDzS/FiQtxT0HZ+/6cQp+OIYtBcwm63YdvRI0EspP4e4ZpGWLRTeVUGQfJD4mEOFV0voa
UAMU5lnTjinhBIeJzfpGDQGaBfzJDL47u9ZHZOKNTz10BgkUneMwrUwGI3RmghQTDmb4c8MU6tsE
ugfSAXBrMGUsWmITmiDlEOvauIwEqdN1uOUtWzVxlyuo8o9HyZf4pDknf8XWQvz5ykOpC73L7YoI
2V110MyvLgJSm/FitSQP3MLIE5ApfHXwVVA33HNcsaiTVexdbRrVWvIJWuf4ELlsGrg0DuiXHoUI
eZGOkTVFrUbl3rLk96ziu75V4Qh1FNKJ/uf5cHt/TML3+fjp9o1EsXHk00jiCrJBwlJ3QW5744Dq
okuice/fDYD7xt6kXc8Jnhg50g+3nC4i890T6Zxf7jmhh5SInmlWoONgq0ajDpJxSxITDabJ8bvk
PWqlWu3huPoPFpI3V+YysK+JGjj43DH2yw3rJE7ISna7HdLtndUHIFtV0s47XyGKYpNph8uiOE9I
UezU/47lPIBMchbkmRX480SehQjsTJzPG7tuz2jTFW+KgkGy0mR0wINwqcI6zE+0viUVxzdZ9axh
iq2sTC4Pa3ZJzPiq88h5fHo85AKUT9dYKgrGZjtNhd2lSASg0GIJnCi/p5x3xY0c6vIWFi/imSZD
ErfoWlrj0+jYBDEpwmk8XVOpzft3uyv2yd8uLWzxyk8IPt/Mw9A8Sz0mA89EExE0aSJan3FaDIcZ
Q/Jyf72T5/PI2KB2rXQuNjieLR7kifJWL1k9kOx16icvTcR/96RMWeiMil37UMc44LysfQ1GxpKh
N1cBrRG/C1BvCnIGFrn4v5KL5WDJ0wGzjIBBhgeOZYx6W2oVxuOx8xYV63IJ0sMApI/2pHXwWXlJ
QHk8YP1w5/gFkdnPrUJyiF7uyz0dd93cGtFwd/67vIX47wuxcO5pCmP6C5ZRKM5aaiqSX+g5tFMJ
dQ/dDtIzOHeoAw+L3L8IpAjHGwz0/Du6sNYfTvSsLWYNx8navNbo1vwUoHdCRwLReD5Tdmz3+RhW
a7eYUJLqnilvQnccaBf04bKxnNUb/o5DsV31MdIT2VIq9+Z10lYV94KLiEB9RrbYF0LTfWFhiFps
KapKidV5NMMrtBHctxa8qCOBU7AdtctDv/hLhOy9q+CtprBKSRvPDLY7NETsvgRDBOZdmLOMz/nG
SVtOjn7SzcwZ2w5jmSCKahP6zhVMyoyQHxnDsuo9dVI9OZQsn+7ajP09oI6wMC6J5DviUdxrUIy+
fCf4+5/cvJnwbYkLnwg130ghZwboIURFgjoDD2V5orhFJegWBeZ0E5cM02jWP6t3FOTRQ9K6uBkb
b8Zx3xUWNEZjb8V2zZ0pe8dGPa6J3XuoZpI+YboFl/U9R/VeO5R96ugVc6758j6XMHz+XzWbfmqI
R/QyuphNZ5x1Vlg7f5aE3nxEBVbqFzHRsKqPEedFX+EKu6yNw8dSM6pRLS5HSMlQa2ktmv0+hOkU
WzMdG+faWwiHbxZVG7qXy+LjD1/LZ+RqHJ3XKMV98CI6S45eCYbWvLr1d8NA8BYMRuxuXJ3FgGkt
o9xvJYzFwvs4oJX3i4u8tRe62mnDzt++hAH7OoC4i7NAYjDQwxrNhXqG4b6pKdZPYOmsXR/aNodW
Hxe9R93ilm0hchcaCTUiPJoAIyveBSZXOUyBFruufj2EMrnoG8U6+zzc4vzgCz+bh+m4xZLk0ptd
EOMj81ckZyGQm8Gwi6fl0cXxaXYgjncO++8uI9eejPz0KLvUtdl08kbhi4H9HWXIkV/vFGkRA6S4
FsOlcRDIDfa07bRiApP0Lr6T+kWq/2GdeBVyzmjutwzDD7WJPZiqsPUVxv93HrwLdovDXW70fXqb
2AE88sajrcFBZYKJkivfN5gAZ21SOoNA+hQEYc71xCCIBXqlL8KwPTXbGBy3+wEB+78bHIYixVHt
ze4/oW+mNifNfJMIbylZieAlDIdiFltkUg2IB1CuM6tSby/BZ8rWeyxM4qqW8ofvtK9xe4N2QErl
wggkssxFdEG4SDLoa3SMSRKOZhf6emJsEWj0NUPnGMnN9/AzR2/o9O3Lbal2WLaoUZ488g7fgOVl
xjQxyatyBr6zk66vOyH2XxhneKGKTiHjjaw6m5s5jhWKeQbwiqpBARiHu2NmN+JAQMuAOvbHkfwe
xdsPeek/2kORoMUseKDfWsWnh8hkmm29rGKQqLQQZ3YcJ8U+QZOdYR7pPH/Hc7/2095gzoMNpBTM
Nt01LEB/RfRuj6J9LLWIrv1B8Fp3WHI4OyT/DcK0kAeTjmSv6t6vZazdAlxr1Eag2R4TzZ/VfYOI
2x9E9HkHkJFYpGUtFkynU06XZkno/UI/K6HSYrrUjfOkSfQScTcR+pnc8kqT3FWVgQ8sWmA8cQEz
il4Pu9U4EjE8YRmWZy6/k1IbV0ZpKXJgyP6F1tPg5FVKoyj1QUg5rBaNp7VPECFu8/WnbU+ftPP7
XMADbOWdX+CZm7cr7P1QXv+xYipRN5vKoB+8wUhGeO/l2vUCmyDHnGi/rGdXoXTtXOjyZCIsNMVs
u+feI7l3SYaywwip/v58GqAyWrptKxDVfOkLuI4GEtyNeskUhmeCV6TchsRIkyp0GhsqiHrOMC/f
XrrBceLbrVzAeiw+8jUUOW+TzZI7ci6pxWnlvOZSFA++ryyE/GbfIDyw+1ClZxpZ9TxEZUd2Vzry
C6Oxc8tM6U0ubHqJPk+JrAuzMI4b0kTUpccBMRSRRHsoT/WGy0RJlAXsRSqXcr3bH9DNzKix4vcO
79R0ZKGQf7QGxihm3fT7wXeCcs5pW4J1V6m1wi3morXnIoDE6GOWLOtGQjgsZTT0hI8hoaehW3m2
zMJWDuGTJlDdP3RR0v0IlrNqe726Cr2F1aPIbUisuqJj7XwotYvGiRjqKUqnAa7Z5N8CR1WEduZR
6tcWaUPJxvnX7Zpd35Sb4DB6b/A0dKiS/q4NvC/C54RaFOYielCNAjerEQV290S2jWcEXvdXDoWd
tkSUxwhaeoRvuVhsjCSzlqnrWkixyQa5dZQleuGHH1Wjd8lY+xpnY1n5/ACT0BeUrP+qC32TWpT0
6lz+7lX23e37TPo0+2kZ0jXdKtLhxSxfCOlEQumjz+w76n1tHpH2bBHLh07lS98OhwszQI6zAc01
3GqHw7Zpq4HbOHFMBRZW8ft+Vy+UyEPJCe0KdZMG7Q3tTTQlkkOwPm3qlEY7PKC1SmRGDXxWHDug
Q9Bzdgo49EZvAtV2h1Cw/B03sXSfD9+YBEl2/UPqmwyMmDc22rjOBLgMBGkCM55Lg4OEMH67Kp4X
/TuET8q6S+8BU28T9Hwf0Twl/oTxAjtpZVG2GmW0p3Hzd8GVvL28XAMiO0v55cGUtsXsh1AsLr95
7KcbRPY3ok7e3IJKrNvCAVC4taNqHKwoF6Kl5OWbm60I99uIYBhxi00wun+bX5lcIP/mSokwcs1L
/OQr2sja7MQltmcWr5dFH8LyZ+xoztQ+iowcL+hsMW1fy0QhRAveeJRExbnTCTAPCKsk/hz+O3QF
wTF0Ug6MPXv/20WVDzy6MB6SCcCIHozqGUzv40dZ4bE3wBV0Yuqrwu4t0yWCG3Opceu8J/3QUGi2
SXYW6UayQCV2RwCqJNfBcBN0GVwRK8JeHe8qPc+/irT9/b51Y7gC2GG8ZePQdc55IUwg70w7ds3g
DlaHkc0wLrtbHyfsDcT3TUk0/xm5SxcK+PlDtMjMH9pQxPqx/W/1KPYeJInVAWKRBM2NiKiWLZ01
NgVx2wa58En2sqR5IyWw9aAfKizobsLDAjIN7/dp5gzzqFtxY+PkAWm87M9ob68u/Ahd8YXAELwg
b4PZv3rc0B3mn2Uo7FpTaUlffP6kiy6kh3VxfPMgy0uRLOtLrXeGnr9Fdx1McJ0xzwned6nbWMbe
E4qUQrrkto2JC5T2vzK+tvBW2gqEy/hxnFzd+YBOviVKOXKVv95HAbj1+m7+Fic3R8iScJ6a7+4f
6k962NPeRH7PjOUdRZ7KX8psl1xAoNWwJqGHPjNq7HWLzpsv+6nsG4X5P51KxjicODNc2vxtzLHL
PAowHXSu5xSCctRfArBDaxREe7enMkXRFWOylc/AQOI9wEMOfVvoGpsp/hHIroIZSxuzNU6elNEn
FtztjM3v2ziCRQbs+oLIhwovNQT8NBfVpfK79JuT6u9fn6nG/13dmHKCpWj7B92lszzSJhZtCqn0
/hLsYyVj7/uoPoJnMLltjRzr5xb5FLZ8OHs3wNsJY6wUYIEYuWm2P68cilp4np3oZ31FI3a66TWe
FyINoBm3QMdDzo22eLP+bxMt5K3gqHq5fA9haf5c6D3PMmDGYgAbtpNSLULCOooor/z90tcxfXBy
8D5fifpF+Wzt6fUqN7D/Mp13TfbTPQGc7fN85tt6w2tzeNmWJ4yGxzW8/w8PahscvTJ/cOPv1PcG
IkF5R58qWuPN1qFCEdSkNjVXvBtmfKlxKPJ9DUy+s36FAvctpMx9s87Sy1aSG/1x0WohMF3IKc/C
4yp1Wf5vrM8KJnA15bJ95UOJ3uX487j7Y6APylDzw5bNCGm9JDjuDZGowKSoC3lbrEZR7kiaSMd1
1Fe0NSTMsxL+mATUf7SOUs72XGa2KDkkLFS2Lg5/zo9RTTkdcjHl1kUADDgA10N/xMZ+nMudByAk
DyayQPDZarH+e50v95cvuSzOrac1rSmLA9Q2rIEAPXywuLxf4zvkWaFgDzLraj7nr2sxv9waPwMA
ObExvXWqwR80t35d3xqM5hvjh7LHV1DnI9qpyJz+w+XNAQHxf0X6jcpFoCblGhJja1Sp//EGMBmO
3d1oYUJ2VV1DOT13B1q+0m5295xd0nZghGcuQjfwxkQvNL/aJnwnah+HJDxYKdmOEqVi6vZrtx+e
z0TW2elTPd8rz8K+MClmWJHAf3K5++OPOFQYb5T46XYl87Ui45uGHj8Zn/MXZ0dGiGL/gwpO2mOF
x3/IrzhZ2NMsekwncxha7/eL7lc/0q7tUnX+4vTdgNno61V99KEXN9UkmpAEtpDYmRxX6mp9KAq8
3nskJOXAXS8VFlPl1RcT3SwXsXE5DUsIivXCpewUn5ddsdvF7xjKKflIORf8r9sfwNMwRkmSFe04
KiYdpxoP1FldGUkM8Nyy38zEOLRUIl8ZwIrBg9yoWhJtAxRXkjQw8qqmNlEKE30GeljaXlY+9K66
hJkW6iZJxiF5MZfuuqAAkEztfLBg/eDFlewzUzm8AHL7M1MZOGxUaIjRGSQNBl/sPlvBfmrQR1WG
hd/3ekGGGqM4x/nb0mK+cy8xYTmI3JGfcTTA9t26ArfazKxD/OnNr1XJ91XclTc88FBqA2w1JLlM
0w+8GKj3u/lVho3wJPV0VS5SbkMn1nZL/Zonl4UEJOV9g6JZGAdtmGY9LVWfX4BqtUNJLc4dYcyt
UVZFDxxpPDU/LhnMDRloVEHCtckUS4bAMDPX7tmMNTh2ur6enMauzrdHGTmtSqKlhYtiNQozMVrd
+zC+Y5xKZWHcvAFWAx8PrPE4T5aZfGxeFh7mYwaCtNIa2PM5hP2WAOlVrJw4k4vYgL9ScXVQnOTl
d8+JjDe86/wO8rxyYCkGk+dOpNFPoRsjUWiO91MV3Js/dldSVYifA87jiMNsb0W34UZP2Ruw6Zp7
lMzUw+2t4JRG60WHqF/1NnV/Ua87+Jrui7AKhCyeU4hjWNPbYexAyF10Wd5YjORVtmV3FlrHLr/k
wfGa2QDRZOQBa8RERi6avPuBxQijUDiltsx+EbUxspaiFbLszcZjVHI7pRj3rZvOHVXMHfEOv4Xi
/ThlmsBOhRHeMRtbS+qxd3f6E/ETDibcz9y65ADtsLdsGobheehC5lxv3lMXVNfJBbq8m57XhGx1
F9IBZ4r1fsIGCwPbAtRSsjQCUt86yivJaq/xOXmpzmK9nvLxsCErVHNA/8JOU7lsSdo3r1or5TNY
YqvvwoYEHz1HuKW8Ri6EY8fYOY+i5U5ZxquUu5L4s0axj2dZC6dlpDdvXlX3uNamg4ptiMF7UR0s
aJmQ69y32ETnAIEzqU6/xtwhW9nAwefBKVH2mAwPZyKTd/E1powb/feXnZ0hL0F9ktGi9ZkV4EUX
BHak5HzaqP5M1IrVVZ5y2prf98MwgRGyomw3VzX5Vh0i6IRd+jRroy1lIE6kHpSiRWsuxO/BxmnT
FZxKtwDPlAyVZz4jAtXO4nLLl5uC0FpD5oKwSEPpWeBeP+g70/jEV77mfTVuWsTC7/S7csNWaZaD
gA6FwRPTi8fhxeRF9SmgU6Jqi/AAjbnjJsSYNZwABwI/la6AxhFh6sbwqYTNcBt8ueRuYb85suxu
8B2W9GBsZbSnL++X6Twb0bESfhVJdGTjZ42XPwP2VneICjLHG0OfrCFjdHs4KD9SxbeBqQVh/3Xy
oFEpAPZ0ba8QfIt48Xvlf7Dk01VrdWxuenJGi1hAshYze+pNjvcxXwfXxiUw8bAPCpO0MmB0cLMv
6UN+8LwnUowQaUIQUcFecbEnh2fp6/pJJ9zEzHi3p1NZSQpxskwvXAnI9wbwg9fl/SJicFc1sMhr
WRcdstZmFSlNv0OAJjLVc3IhD7vVw313HdtrDvCZlqY54ZsE70yUpMMme5AnfDLOMBuKl8DJZWuX
20b++gUuajUjF3YbEuyrsqZ1pwieLTH0RYtYOVEi9nL8VNcV6rIL0SMvUTPPwdiHzxXDeDWWCmRW
ErG5ZdiXr6I7U4h+Z/GenFhGfYRXDoMwAVZmHpWyJPUjuaGLT93GJIuSjDRdI12Y4+wDZbv4IVBB
l5NbTxUM9Y2bbmtzgpAqY3EKJJT7Pcj1SsAYEXA2HL/xsBtObzf8vye2XRXxntAdDfSMoiXJ7USi
doj51oRq+XiYSTYxe51HVNWY/330LXpYMymGNkzfuJvdfvv1ad0+i9b+LdmhMvpa6k6s0/vekxmO
L0hHevVLH2NAEH2HTybese61ssfLCFys7pshhfBzlyrIqkjAzBAMDd62qhYUB/vOI7GnBN6zDWau
xh08BtLjKXfIWM5x8shCNTAY01qeRgwXgLZJer2WF6MXVc0uoA0vDYMS7Tmsv2j2FcDo58JV9NbZ
bjkG4jbGc5tAPph3bVpwW6hWvSvlTbOHsiD6mOTDtrWKMNV2GNHlSCxWteigGhFpXQX//2Z+4XNx
GmmL3gZtH8wdhVJH0xjPZGm0EcCjsNB8D38SyNDWMm86hh8N6OH4Vmy3VfUqs7PO74qp7PKSzHVq
5dsl4fx3EbuXal+zDRYGe3igWe/3E+cmevJzLf4frVAp7pL0KwYoVQ9BYiEqANFT1IrX+wdxyao8
GIKxtTvI23N9Hwxz55UDYldTwX3ib7DeMl55uIcPK98WHilvwMH5O2QNIizYdi/CG4q+FrD28+7C
QWZtzhtIakIXTlx9KZsC238YDXx5m3pjlTuoweD7QWhW+uND8PSlLP3zQ8ijTSELnbWWS4gbjUX7
axA7xQKfKtDDpJDzW2Vc7tbB9JQoLvYtk0i/PHp6HBkRenNhhhTRnCSfANcYLYQ0d4HzxSpoxtw1
9/keM80Non0tjiWtsZDVS3E19XLvH2cW5PNWIEy7XAhVFEyOtQNNh+6BjIWdDlYXUVJfrD7oYt3Y
SQL5KDeMPdR7pBUwoD9UMjHsuT6u/EpbriY3M8baWY1aU6SvV3X39+Hb+FBZstUtH0TZiIeQCRvH
zpdRZYYhl8JIYQP+S7u6XAHgafyVR4zB7fnzXVBnH30y83iaNKE4VRQYWwV8u1Dg5YuArfYxU8hw
OMcaix8g/c/y0xdkzkoGy0pXGHSLK/SAkv6lAH+eXB4zuPazPOUe2okp4toMs6D7bDHPeP/aOFJn
G/7F3Xazx0mtpI5VbK1BmF120iWLdbWga1+Ce8m74e5m1N52yRXHMsfbeQwDYUCcbyKN90gf4up+
IcISz3HyUwoEvsfQvsxjUl8Bey7cP3x83lOrDHxxOHE34pQgA4irGKMSfeIjvIcAHd8spFTKrxOr
b9IqsFi1DuVtFggGZ/MRrLt4KXEP4tl3tj36dBpxd7IKIaOZQq9i/BpJd6Qud5jEB58RNSkuSbKc
rLK5J6II+F351V/oyjhmtSI+g5nKFT424kp7lca/ChZ2hX3Cx8JuIEjUE/jIfXvbL88/Vvz45c7d
k0slWdO5KEYhOQSaa/TJsaW+PCzqml7xdYMa1oX2v/nd2TnYsSrEAuB3oePnAwAEEIprP1uDLImJ
qFe1z4qbbIgTqe0FixDYew8IEkCOfidxI0Ayf77gtZfK1nFwhXlHd3+M2JRW31FBCWp/o8BQNiqs
s/Wiu8zR9Edz5NfTYnuAWPEwWTXXSpc1QNUL9R6dpDkGXA+ljmsH6/bH/RPUxXI0Wildowaee76E
cGljDxfDzPHwUOwbty98eGIEiAuFDNo+qYYkfRPeM8e6zEbOGxMpxUt47eh3fqAgRd1MZ1gHEcpe
uDH3E57R5uERP2uSCKtI29B7UvWrgyVZVgujC86Vx+WdgW9uSi6L6b3MCu80mQMm7pClIKQEy6uR
+dpKybLOtTYstYkWCoNRyOiBkKNgoz1RSSDYb1ICFJgM1mWOC92PNxcb5fwEgQ3i6mjNimlHY79G
1TD/ZfRzzTCHvSWVhYgcrTN0LaxXpqoVl/qe0+i/BAe2gNfR8oPJRRJu9ACVhxssGK7hFB8xtt47
cP4ujICA+qhSLCsj4pDk+POz9ANKkgXy8DRYF+h879kw5A1Bu2xK8Z6/kt/wGVQRuo+zcJMUAnc1
fdu54DleHVBysSxYVrrS+hjBd6S5NbyQ/OUENAh+8WV0anDPs0wNuk6ee+hb0I8iIQ7nTlwbYWp3
b2m5s1hWKHtOaTdihvlep4dshODdM6TRZVSylnQZQm2Y4ClfPX+4BVn2XRYzOFBNgDEPZ1Vinvxh
xKZx0sggZyeEB05D2EmxrUhZA5a7XHSUObWnNHOuz5O6SLdTxP4cQh8W28UYTwpStv+qtN5ZLb5K
3lF3wT16BCCROWw1juBXU+mEEGjt/F82roI/OKd0NstY+NBJvRjx2CpeND3L6iStVVYb63TqaQSz
ClGGPSty7oRA6XBC/H9XyU5PcLvMjmJNw0Ue80/qZAyJQ2K95UbU5+yp1XHzMNUWZL4xZ6wFvw2Z
8n+DzB0GOzkyLIwxE5UKfayEG+k3MnZQLxoRGJDoBK+UErd0bC0Qz2K60T3YCfh2kbSixyL6g3AE
XwJUgVLdl3GUPH/9HV6KVkN44bzxNoCWGLkBXo8QoMfieEE/N/JFmM7TbyyY92kEa7ZoZW0CzhAG
9e3HQvfF3NHXmVDWlsxVH6x1CYyPqV/ZB4zYb9wj9uaxKtGuBv5L9Y+9grgmLUOKfOndB5Sokq1U
wO7qMAA4IIcdEnbOhLVklGVGqPZ2MHdsXiFCKztUP49V92+kK8WClaNumoJHR1KHGSV6nAiiXPkn
wqwrjFRLQxrEY7g3AXSRv+r25RH94fPyWZlP2BRQrLiDGCS2tpxn0XzhJso5HV4wsR/LUOtaBIz2
PrA7JoRo4UQnuO32W/B+xsDLAojmPyL1rbSLnmpKNELeYfbKzCESCsCSctbe8E5BA74oT2SXkFBi
Yki5uKNENqXXijtMZE/wXFeovHNBVcpeoZoD0mcCrQfynsa9H4BchptcZbXcuWzpTgfmvX9gUh8U
vsInE4k/l5yyfRTvX3zxhImOqKyLLuD57XIKeKwiMayuyHmxo6dRqOUfJalGPwtblMsI5vR+rZk7
X3Fb74OeCpQVa0MU0tOUpF+BazpI/Co1oIp27u55Zh8FM3e0mjq8sw+sLNxAHVEUcNYcDk/7NRyg
42crcgHYuKWGqv9ZppWUcQdWItzoQswrE10y+G6KKRzOYyOMxzSlrScDwO6imWE8EV8lYkeG+s6z
u/a01BuhBsBwyjBHjp660Lp8cSSo/VW+Ci3867Vs9pud004j96Mxw447uyZQSDJFHMXUK04x8O75
azCWinSn0qwASKhvO4kHwxha0ZtCUiWL4GzScMovaxDgyhQV+/SakR/8LQFmCarq1Tv5EFIJ+psG
GinkG7qEi7S3M3ghavC6XwoLEyozUtukJN+hQavFsHqh9AtVBO+qs4Inp5O+Ufrhdnc4GngdONbj
6gLeTdWH4nAAM2aT69J6KAazn79hoK5PZvxl/Kq2dfD/X3y/qqqeuKW2PQrTGx4Ea5AsIjItzNDd
858I87qmvKcHXdMnvvKFEAX1QGz5wBpoQTCJCXjkeNmKYN7gBp+ReIEi7dmNhPzKs0HCBQTjDt6g
H0lDVmjNL5Uv+xN4jd5mxidvBK7puP9lyqwwxiseruXhASI4kr30JviVpUWdWiORgIKYnqlb97a6
Nj+EeWRK4vZcuvqQOIjOOvNhnFaNyMH2G+hGrh02yLuJ7kqFHb+I7Q29jhyeKUemBWn5VvBcFiuO
CGnC28D1nKQ2Mq9/nAC8dJ3oV4xK80ZAXbLqv2HLwsoH6BGegAqSNPPYZWaaeWjZriWtg31bL7ED
o1LcmXb6lXKUCnYv6FKlJ5FsixMQJcYQw0XPBjHiODrEU8xXbrR+2PR6wbqAIH6a7rMrGQVBipKU
qD4ahkGkAFzXKMWbjDK1OFkurbRdtY7XoG/UEy/atcYXxUl1V3sE+v+Gs5Ww35NymFJSG+4GuFSj
rCMRD7Vb1/WuTvY8zgLD6KVgHira5r0+pOKLaLcryUtY3WwDja9UMeuM7l2F5L9U9GZkmtT0vBNV
7xAxL7TUrg9Aif7MY9ljBrdKl81bi2KhhZ8tFjwgexC/M39yWlXmIl3prXsCIyAmidFyablxDTcl
cTGwVkmr/vgeVSkhoLiUKaFnbhxq2YS7jHn6XZYHEFTid1r0IJyhyEssTVPIJ50AXCQGWs5upYg4
xgezYaAWwBdqlK5fQ0mUsbCK5ru14tmSqIz5rhJmorA3wkTigU/nMsXw2HJs/SlhhZVnTJgFMe/t
xtJ19ytV8DERa9vLXHgbZmMnZdCqQzwyTbSWJJsmV8WN2NEirSFAGrkEOSGkmNN1NqlNwsoWlhtW
IAUv8KyXI+kgXyZ6/0fEUbZOmTrRFmD/gvi61rrJO8BKs9RXb7wHAaZDq4edNxWtiIkF0PaSL6Ti
UQulcnPv+SJeo/KGqMCUbjsQD/IUcLzPOEaHymux8BqjGEulmBoObuQ68vMZGkUti4r+Kr+vg5Dd
AKpAtEczaZbWT5tIa5q3E4Pa3llwy88iZg+Ojx56e1PemS8/A9AKhEO2lbJ56f994sXalZLySwp7
/TCkQYBOr16bEYS6dKwrtTNGKDczGH1GCU32rVpwgFgziEZNSnADG2zSiqBcFrYcBltU2+Brb+Hw
mNoDYCY/hex51IFydDq+dfWrXgY4phhBhtuMSHT4r+Ln5gK9hStrbzluXG8ZUSmwCkh3edoxXQEL
2XCqjmxv8d9MUG8SFUvuSxKafT36sycnSPByRZi6DcR5AgZTc0GfOBHANlWZMptktD9R/AWRAxjO
Ykq6r2KZeF4hXvHTuTTGYDvU7ic2CySPkF22sbRptx4YY4yO0JBwYcBFcLvEWzUYj33yxhBxcqmV
s2lXrcJp6qLjuaIa+hqmZeU301a9UTW6NPvMT7HQX01qlESY6KTb+Ce09Tg17RQ5oDOxo6Jdn2cn
ovNB8DPiUHfq3NKYpPTac2nkFa9lP2QaXR2XO5DnaOdNOIM6L5roKeGjCHUL5YH8IwxbljaloUxw
m+VS37knDucg5HZ/yPPkVrfcOLiO4SynbQdor90jQzzOnZYWyTdImuDgacqfUAeM2r4IE2sqS5JN
pYbP7UFCkNbkdmcBNFJ1hvXS7fLe7G38wfSXFhO5ZN8DbnynD4K7oPE9TXf12Zdmtr1Uaexip/rb
n3l0WjP0NI0sKb+x3QHxmf6rAMmB0e9ZbxCGjFX10brry4434XrTwpRNDdb5PR7dniAAPuYJ410T
gFEUM9TbUdbxIRIX57udlYQwpKgzh7twbtRIk/+ewlfsD1ClH6ynWKteU0A04upb7dgWJiMCSwyE
sb/7JtQxB4UfozXu+gWMQqSIUf0tmKr+VhIgI4ErUUxMKQUxKXe83genlqCeJV9uUUOrcJIvEHBM
sv1HoSGL57QI26DBiAmqymf/Hwc+Ka1646LEz/5RNYm3ycBUFQ16yhr1/5xzLNHA+cz0jMtZk1VX
zu1cdbY3N82OK9zU39+egmYokYuirU75TM30NL6aohT85UyeK5k1xAXm+3GqFw18x5BM1klRcf6/
BqtMJppFCEj8jExGzoP4pETlAhW032rKnbT/X6ZxbMaZSxoL/QrS5IpYVduVNPJhIfj92dYiczw2
9TAPzwaxdO/l1vQvFA5bzccQgxPICnOgx0BsXVr4hisS8Q3lsSeGVbNi1KS8aNp6wi37z0FF4dA6
ngF9KgaNZ54wyG6LHzEeoBqtnWRx6mYUZBnCCRDBl0j/id7SgoutmTTRMsN4IB2bFKR0HgbB310t
u/0vToanIW7KWZStJC000JHcjz3IkeUWqaIkCcVN+nO8JcjILcu9+9sosZqST5JKzht+BisjFXan
ml0CbE0BeUVMZpjyc5XTHeQcIZBxZqJ0aQ7ZfV/XPv6YyDVCbloSNiyfKFCiLY8AbFGOEzH3+0XT
PEFtWzuNk1mDqKn2G6uQZAafiySi7Mobef5T8VlgFWRMTTMy6Oq4E5F8L+raa7T/m4o6M9Ml2cHI
ATFZNBJYGvp8/MG9M2lwCKwyxGc/XJtdkA7Y9nTeSynLr79d/1wvKwbGbg11ipur0qxxlY8iy4nh
dgfZpY077vJ1DfuntAgfv/+GDSsNZOwRBri5Gw6LXHZfk7B2M75hc2OBwdwhnyZQ3VWLTNkGJUxb
hdj0Fz83zcEKkiFWbtHffbu26a9Cf6oy+A9h/FpWEVwB/ee3K2jmm8TSmOV3AAbAZg0omDSwtKBW
VSBQV8B6YM/1R9ZKjBxHXlQ/4f8iFBhUd34mia/2DLxWqBjT6USAIwlXdMhIEhqkuZsml7ELxrxm
u7E2Xx94b4SgCYK47Oje3Y26JnefCDze4efU6kobFA5Qkau+T67Jop4KCUh/I+MMRH/I8VdmY6kl
oRjPwcBzt8v2QB+EAnsj+Q6yu9e0M1atfpbUWYQFbsFEFM76rquLHQN+jNlsgAzR1irhXs7mTuR8
GcpHVqvmBOiK7NGT2gMKLlHaaqKnXxsJDx/0qPnhv0lc1Ff1enLx5TSt5+N2Cge614AwrLXXSaZi
xnlMsD7PU6A/z7hhxOk2swJgMylWsOkxcKG7ylmNJv8ygxookVqR/Q89vS3KjHBn3REbquu9WBlp
269a9YBXepy+GJP82Qg8xsfGwc+mlZ2Sri7aArMHkgJUYRJ37rNH8yB7eZ/Mb1A2wguKPifyIG3W
wo1Ntlf6v7WHkUulB9n014YnR8PpHVlOBzPJFbGG0RzguR3ooT813Zp6lcLFO2TfPf6DkjCEsjei
PrcyGIOVWrLRwWHod0n2DVCGras/0GrwhNsdCkvW/Ads2X+4Ibw3FGOhqchafPNd6o7RVlMPa6KH
EZ1CW8nRsa2RT2q179bqp9QwbTiE57e65NI/Fva+FUPn1bVlNyBDnQHUvlbbWVLIms3YrF4sMX2X
fWhQu3H3qYG4t3rUau7nICGl0Bm5E7N2TS0aDLnjMk041y78AGs2bEJxfhf8PXPn/6xg62I/N3Xw
ZNW93rm+s5lnNQ8SaWL1I/JyafEz5pDFyZbU0AtldGDS1ZMbsRXdaDycd1/0HTy5Ov1Go1cz37HN
VHwNUd9VIdZol2Em/xKThP3YREDjZEEfcCrDmceWjBK0uT/tvkvI5P8+ADfA4jae0rgUVQkXEQas
bK9R9ZvO2FrsPZ8WRSMOaCDoASaFTWgRgZ5sRtjBNgmHLosY9bAsbuehhGl+gFWXyJ5ifDnAqGfM
PBjhX71Wp1Snre93aVMMq1JrL7MllwnN8BSrUPJ73d60lx+OQTE/nYEKPCIRATCUhWqp92N1yRiw
1QYPpqhr38Ik+S8KJcKzRb7/g6fr/PiieguYqBw5nvMxtywxAh0+v1zkK+NFABkRONK8y3ksOl6k
d9xMuBBoyMcfUjFxwsS+quQ12+vR59ehbEUi/COylkDIylZTZBJnbJXLLiuY7QNG4ZeriIK/MJm/
sAe8dJOCXMhv/NhzTjrHTyfUo2ACmXFdcIiZLij3oYGnYUprgf7LukpW5gDsx4ry/vLe2LFvjoKJ
EKnjYoy4F6nlUiVpgi3CMQKdcaM/Zvt0wxeDEL0iFvS4V9TCaamrcRbxZI3sQJ/FuxqvEIRVdPNi
e4PFP5NkPT7SwGZt7hjGafA/qngQprH/bFjkJPAihBJ6HB1DmgpVN/zRExDvHPdxSLlxoI+7IvWp
/RyJlGvW9jvXyo2hhqrd6orc15iAmjM3t0d5H21F2ZShWp3JBDKacSv8yAxcA4LaHxxjesdynp/u
IMktxfJ7Q08CTSJYqvmE+jvkobpmIWFwO+yxMmZKvwJWVjcUQ+VD8uSP1gYYm4x2DdyTviY/0w0t
oM0REKhm8Z30dURmDv5skj+gMPvXUP9SbbHVG4EzWwWfiFaofJ2IEu889x24nVBFfcZM0rh1z/vL
Cn3u/qZNbOdxAEcYWu4gLZMzBevdiNVH7vYMu2/AyALwJuxAdKhXNHT4gQY3tm5j3rwXAu9JcQBQ
4Y+7MFC3SW3duM5kDbV8VFd9EBLAOrDVpQHODvsAwPDu+aE1yzdf/+aIT4hUa/he+L71bFr7jzLH
1i1axjbxkDULV07NsUu4tv6P7/IbVnC2isUo6lxpyozE++kgBG96onW5puB2In/XflbjI0BgvqhB
cz0c3kw8CjVil+tufXkg/yB+/NnCtuLAq0x3cYrk9aAnId61xncTzOqsT+PjYGQdgkzdIpJVjWpK
72I2QUHkbAcOcZt/ZJkSq2dL4WgVNo4U8rWyfTcAZYm79+SHMYllCBXodDgEKBZLRmPOaxuShEt7
d8YYPVeY34bN/H3krwAKYEBtGws9ebM0wOGweauhb1L6rxFGjojT50aaLWqsmMjvI33EghsasSgz
L8MrUzy6XaVv3ZNBpP6mnSf1J61usF1pdBKUFqxWBBqnWxWOObzP0mAhGNgdWZVIViRJkkvaV44G
tJiu6mk9ShZTcFViYQgCHNd5UwQsG2H+CcYQ6IUIdEqIQh3rEf7fiFFhhLy5DuUOADt/OfzH8tlj
nkLbNC7XMv8K8g/3FARiDeuRAj0M1WOzyEF/2NLPJWuNi5TJSLQxGLVnt19LTthxFsb/NkHIR8L9
hgjsZp88yln0X1LHUJT8zeIK+uVBA63/Risgc2svUpGGw8regSPUnFMeP8zBtdI8o/2jaKqJmCzQ
QrK652bOFdFabWFuD4vTzuiAFpwnGQQciJ6p2NsbZ8uRBnCvoVYQ9I3WN8fRI7g+NfVUtcZ2EoHb
KDKK8Zdp86EjC3wXj8B8VObFkpSIURLtuj6kCYipBtUc3EMKWliCpzR+22Dcgxz6gszEN2ByGRXD
QohbXX9j5DfRO6Y9ZEnDI2q8VLQuYkpDBHVihySFos0ZAsHTq+e6Y1l1F57s5E/4m8gs+mWsRK6f
XXx3QoUZxxJtwQednkeml7sg8cURIVQiV98+WjK8E0/9gaJSy+Qe9Ew8yIErUHMF9BTkTgSbViGN
+KjHzmGTCIH2z3j/qyPJaZ9Wa65avztJNNwTiaV3ED3sfF7tn5hhsLzu32Qz2hqkXFPYxHZff+oy
9rbD9/1vs6r8isGMgM7lpsTnc0m3/nyWNEkVMbzElFMWIaEIrXDAeim6VbmhNpD0hpHyIjPGg217
VhNmBRwiJ3dytIIm/qfleGp5lf8X0b5u92zK8q7vMIIMlgdXXCNC1NGhrdCfTnWTZs3Z/o+Ie3I7
9fI/LXWxdBhZvQPJhbPkdPQD1tp3JZLarOV4NS2p2YJiyv36cIGbm1hvxk7LkVE/qdruvmQLZq07
I52BRktP2Dr4La45n/cF4SoUsXzSc8g9kdQIgYbqEftlmXRFC9946L1VKXrVmeUCKENTy91OKM1k
frk6EQL4t6K1IWtZAqu4uZzicHduPRTk6SAjm0HfKdeBYcwAIL9E8WHw0JeRMBATbRW82uQcwd0m
oJMa0EAv/P84oJN/0m0WSzf4FPWDMEg5jB/yNzEOi1mif4pNuo7OyG7C5FzFspE9uJTKKwGDh+Jb
ZsjYaGPDWPmr1f8p5WAGL+jkbG6A21qMpbShNmSgn1BGBXAgm43DV6GOQKnR8+tKQeePTLWQYi4F
keUrFy9zMb+R9/IlVDCQX8yZrRALCIVSIxOjo2T2O5+tprF5cTDXH2YG9OhIXC3FSf8K+8V2kPF7
El0DugBkiXE7a5G1pvqpuz0A0/0SJSlEp71NKq2/zoplc8VYJ2ThMqccTpd2ai9krI9vf5Hb5HVA
RkzJRgnnCSqWwUslr2NURQiJciYkUHx0TSXUwmsrTz+7HI2rlzDxddVLhHYIsumWobtpgCMF98Rk
9mPhFgyUdYY/ANEGmKBZwiCxjDwDbYRtYS7pryg7j5ZLlDQj4SRHXC6+wGj1OUTQ7wQdsCoIJSFu
N763fkOtSBNbWA0c9msvWIoNl35PYO8JKqtfNt1k8tOPdHcc8E7YQjeuVULKMtB4Qnq5AgorqW0w
cwX48XBTcQVblyaF+vaRF8Tv/UgtbuZNvh4s/nr3uKEsDUqhn2wq7391JbIBe9vZrUfhgybO+DQj
6TldZSrEQcMq5HMlcQifP0E8DQvv6AXkrVbb3C7WP3SoVaSfAvtFNFKS2w/YnAmiADZJjYtEZRpc
eFrW4LtQtsJ4fjjHb62vfsHXsHqtirTydGkjJCWWRDLK14wmafHhcQc34DUbms4rOn6idtM+bmPY
9BfC8BGGLy1SuKloRP5PIc38aMfvmjbvjQlYxT/8DStI9nU574zK+oXru9T76b9WgD+DLr1PV7vn
h/KvIx9U2BlfN2bny6npb8rB0SWWxMGQ/Qn5jJEYaniNydAWFUEigflxJ9sP63HuFvi/AUuPFxGE
tIdRQ9R7i5ONe+1xxBV6Rrs+gDX6cV1Jwj0agcxd71MmyK6kxEzFT/qfog8EsXPyVlA1V4XKKM9X
OhWgst8UshW0i1b/ze7rhwS+0t6HAO5mpG3g9KwWLEkFgNLgUNtCzogYCIuzXJ0LLM36AjUBeVAJ
4cEO4dFIB22KhDMoK7lPcZt7+xqYz1dGNhiozdYXokdgP4Qaqoq4tyETv/eg4HMUyJzjdPXtCD/6
u5MI9iBOn0bRnJB0T7PwTXKCL6LiBpCQzPidkv/msfhCbQS0cTaPi5idZbGUShMRkbD0RUiSw/3x
OTxXaYI0pyKtl+DvfGjgvis1wBiwVt7M8pvOB+IhDZg/SMVpVjYEhPeXlDwiPw4170xIb1aBiQXC
+E+BsoVAp9T5bweIW9ep5SterrZexLyoR11fxCNszT82WN1tpZZ98MF5XTBSB+9tz7Z50KrQqaN+
ZEAxjKZSG3pjFJ7KTgK1qGkZB+PkmKdPyGjiZFtVh8zG7mSVAnU5ariYXX9AmIBEwoaoCXnD7xJl
WHKluqr2gbRlm7jqcBeG5SchVsTrOPoCQ+Fb46VJ17UGfKSjVi0pra94/Umwq4Iu2+iLhLJxK6jx
wf9EsrmAh34w9NGOkAXEzb7PkUwJKi5Ado+Ioze6F8XWtirO7mqe8lj/ZGSdw1fhawJWGI4sRdZy
jYrhPImLRfcJnsMKTbC4As7Yhokr1F3wgvNXx2GgWrrr9NDm8sN7GIh3/TmOWiFSkrIJWRd9dTnO
X/uPpAMtMoYOkK5DsR1J8mrUY2Ca1KS9xejQsh1DEzTYp9iRRkIRswQogVvohRF7LyKWF8sJJyp4
S4qxv2Nvsb3OYirfcGDTDuL99fTpRHygL1jhg3ki5AKpLrvcRrzT8qGFfCQZaqiLew9QxWBVGKvf
0LnBATKHn07FrrYzvmcL5gx7zqg0J/SXiQNtCeFf8jBi8aEDgimBc2o1YDa18e9PZ24SSLuz5FRM
Nv2JUNit4rHZ2IFfId7ZibMtemWKPqNZvT5div9REms0Vsk0HqAKuUSce559voLQcx0dDBHIExEf
jsxgf6sRE3oiA6qrQmjibSFR2f983i427S/WHB6eYG6zZh3pddZDVBwB2HoOxLkDqpQNUWRlGm7X
xMCnPlNqxKRsVTSsxP6Y6DUTD7fG0AjaQE/skG9Ud0bN3GYSYXsrVKYcnfS95WKd2BC6XcNT5Grm
ppJntNBLfMrUkXDqXxuZEEKWx7NbcNY3dUojlsvY8VegdSAOyrH9NYd+1cSIKUvZAvaAsXv+jdLd
CX5aq25CakobgNdu3jz0Q7BxaLvDtg35wIR2UGkJlSpa5C8GSSuUsS91mru3IHp0S9R98ReD7gds
DGicwa6KdZkegpCJGC4AH7tjquyx4nxG0I8bnzXswLM0wek6woLb42IzBZn/OQfRPJ8qlHeYvwfb
J6pCAYRrlOOAS4o5IQGlBZza2WOSOxJQMTLxDbr6chcJWpbZFCAh7XEZ1YD6Izi4dxeakuRIxp12
Kz9CRR4ZWgCnetdrWkTJTPOKBmBTzDPnXxSMfSWbw/hbxJSYX3Som7pqkCoSWohic7xJYOIyrYkE
uqVaySZyjnPfyAcOsiQV/5C2qDWdcIVOBYUJEwImXSX5YZ28yX9tzAjzcVD5l3Nfsl2SbR0eeLIK
gjHBXP6tb4F9S5rzxKYluCwOdaoBFneHM/Ym3wvdSgkCpmBIJHr6nj/7YhYqRtTB4ERaI/U19yHj
gUaOM+7jaik3x1mX95z1w1pNh5Jr7Q3nXumGnYyi2iPwz+eyu78u4wFd6N5uuIVjZZ29+t2HettY
lNXNI7xAwuFZ78cRuAUWwnDvUrVOw0kFoRsp5UKqKG4L7bdtD1Etkc1vT8XuvZMu5kD8IoY02XX2
fLPLaZhNxtL5FHkuoJL6EMXZ69YTplNlZNhHbPOhFjOwWa3mO6QF+PlG9dMFWy4iqVq7E41E6Xid
G/vjDU/clJgW4j7qUYNJgCjtOLV9NDDaXKzGlJ2fhPeDdXddjlwf0V/DHQpI2uR49g1I9Zg1cieK
9rFZolsCsX7OUOhl0HjCt32vQ5k6wqLkhOM+myi1/20UTpdocz4yDFGrdOTIgk85SVREKGRG9b6J
uKer4hyHKGlIV3t7uEXtw1N72CxaZulMH+MIueWwvMKxF0Hx3C4Z2d8nES3INcRvDxtVRLlMxTnS
dHqvPnwktzgcc96sNRxzKhtm4OAClzqiRERGwPjmYSQAwUgh1PF3JG7NhZspfXDwM/zUaOZP5QaP
egKPmgwiDh/ikGpJcUIJFnNAtHnOdVXZ2j1QTV3cNO1JOFXBKsC7ziLUi3xoYC/1vPgT/Suv5Ixu
W/LaDEW/dVToLuxOV6wawW/3PizNhyY1wcxzU7J0szSNQhnzUFPVY4SXxWvVhOogqs3N9nlO0IH6
epieJ0YuFpXKIjfv/hOQxdinsaf7TR5jocBTSyP9+vEvyftXl2wEiBsXuXlmS26hfa0Ln6LkY3JG
P2t5sf9NT+i2kxKvK5qWxJb9juMKiMSWH4EqLErNSPi4Gn55J0AtLsJKmHQqErygthTkXeagFs5F
FhlX/BRAgysHqqajEK6QM06kACosLCH8V6poQQlo2xcaoFUoQXKBZJu8Y67Iaj3qdGqkuoxPX52D
wbb7uyXAWBQAuIWUSOHYebUVyFqhPPqvawY3l8IZOMiEPQ5lXB0/7ikRSiw/PxQMmVtQKYGMEMfh
JVQZG5c7iSvutecGCIuNwv7ucpt8C/ijPp73Owa040fH8tyHVOei9o6Tfku5PBHGFMmcpQhy5Wh7
wsqHpbgbI0xgoSlmkDbG6/xC9Egv3SscViQ2Zk+g1wF+x4qofCHMuyK9XlX5mW5DjxeJTdaqtnbZ
GT5OZjUTVeh8113SjgI9vzKThQaMBsZXuSG1jm54XWtR6pmhyBF41Hw63i555kl9r4+E6HI+GRpI
QeXcV3zxoOWrMGyPxRZOYApwlsuZrdSxJnx4vhxAfpUJPSOVPoOAr0fzVpIysmV5rnTFA0YM8gZv
aoixJ+PSeF8KIzHNRfZXHPpMo6oXz4p+PAp3Icd1fzfTQADibKhavBdTvow3bng9WnX7A/BTw0cb
L9652/EBGGfWmrsvqIoASepA856cs3rFA9C1Oq66boYY3E/ZI15E3B/ENM3PoFHiiATUZyyGWFQA
h4PIXCtYp1aL+pXQpHzZ3DKcKFOXv4CM8irrlPzsmmtqTce+ANi0Dv/iM/pvHyW+5vP2t6B0i6Gh
xq6rWfVw4XEOcSxikMgFGZtW/rgxi+lnJOAwuReoudsQVUjiqx4xPzj6XasaQyb1udGt2XeghgDq
KKccI8wTXKVAqN4x4/vqZ0v+0dJPz3N5CJOGLdxfLVlTjPq3szx0/bk3c/ZorVgihsBuKtT000/L
U3vbMM5MUOqa9+VvAnsBWzl2WyedbJGMmvkA70uILzajdZr69Qx3OQkjqmS8gNePuKnn1UsiSQWI
WMzwNWO7it0GvVpVxdfUM5GFnAyisIJmkXmWJML7Shg7y7OMsDw+lNThqzdAY0IU/4WgVJTBfT/Y
fsqjqFVL6b7Jc7xA4i8NY6IkXJzVVJd66LB4vr9iVvNUWabMG4LVGENzVUbnOb/VMK73ULv6rd46
V4UlngdI4M3zMnHpXDnLHC8nB3jjwHYObAcBGpfxRYpbVGzNLEFeQ7Z3mC+yK7a3TyMRFr9ucid+
UEoun5esmZcDUaYve/tjuhro55Bi4u5aM8+VlqcF8OXdFZaYOdnWo8UluA43w0s7gEq0yM+N694s
cOHkg4o23dvKITHPJFx7e/pQ70uyW837bs6t9njTTi4urKborPUbak4GBX6rOwZoKybARgu8aUzQ
0OWI7CQZaTPUDoJfcOXFVL7Ny0HSFgf68V5mjWGHNFgczRubcwa7TvsvemINCcWYdiUCwlMBwEF/
6i5FMUeUV1DwW1GCkkcdsstrfEFEDguQkFidRORDhW3c7I92Dj4p1FqJ4O7nXp+JG8ATeFJd8DwE
bYA+ddYhfTT6JNhDBka3iB9Quiv75vZR3Keb621WUnv1+UROoAnqpVs5Eu0RLkorMaIMtTTVoeCU
Gu72m7u9xJen48tADI5VWU/PsdOd5fnh6+n23NR/LzAsOnkAo7Qs+z6pkgXSHsXZXMY+OpFRiVMQ
yhQNUm2YNk1IVG4GIjxRKsFCaVeWOlJMyRcXT0Vpap24pl22oe9bYjjWIZI2uy0RWEn5MRKuFIb/
gPYl5d3iXfhpFUFXY83IPrZpJIATlKt/vl+fHaQdrpbLXeLayHuM0a+XYVL/YcMgKbOMyonA3o2M
JNz0W2nYnZkiEQHN5/4dKlYIsxxzPt+yASoKPcfraOpAUELHPNJt5Gdq9ffPdzgqxW96yHtsU9+0
7sdcY2vzb7FpjAaSkmHX5iNKuqm/YwgWSSqR9QUGAcWJci+8yL8ixRZyRaKZGpKCRa38urHc2EJg
RBDkRfJ0HypTkoArR0xwk7/AFCARUT7QsYCNKN7xQJhavCyff0Hzeli3ExYidetA+QuGZYYPd8XU
kPs2InjQhVGS42C6zEDTEG+YxfZ1tUSeW12HxyUTSbSucdISXseLWIkr8EAS6pVPAG5KqpAUiGhF
CREpIbXYte9xEK5SMBqjubREKakQi02/07FJMHhVB0Q7/KI2A+TF+DAEEOfMkKU/85oi/aFOW7+4
Am3sBttz7KCXANDvUL2AKDR80r4CIgL6kY757wtHPEIujCzcFPnzbnC0IktOZoUzf7puizwQMi1U
fRldGNAfggmg8Hu+5itWLlG498bhHhM8MutT8Zm8I7scVdiG+1DrEmXCUKpOffZ5+pjOUf25BRa7
5n6MCip/fUR9YbrMJwIHQnobHq3WsF8EeV5hOUIj16L6F7h/sQxM9nmMtctoX1OVQ8R8C3HTYQaq
T9I+dPcGY1vHo7SjfSlStY/y6QuNvw0ycLKO4ysDBWHmt/8mF9+EWb7Zfyt5g6SPzKdhW/vQuyKl
qxOur+gBl/0M7lgUzgyXtbmeWv4tmIf8hirZITxmbvbiRZh4M2+tAXASivsbnT9wj6NgPWsIzB8/
YWd1kFBpaEheACLx/xrUF4nSLSZCz4nnsTppe8O7qSHI89jDyW12F6pEK+S2I6NMpkh0nz53L433
/3aXoDPn6KhuWxb7p0t40p129Kd7P2BETQpmPeVbcDsEnZ4juhxre4iDaYJ9SGbOldJLhsuICt8d
G3ymvgzhcccWhiJaFXK1HydMOgLREa1BiHqY3qdMlY8o8w9HEHoi4QbkeUMnHJFpIE4IM5ekEo9P
q5UcIsd4t9NkJ4Q4kwsvLoDRg8+aqRJfU/qIt2Gs6aBW4n5faEbW6+Hu+h2mAZHJz70xuoJqKral
WmdddzTzGJ8CRwsnclepVVykE4dQbHm1yK8HA2CXCUcPtWWJLf+YRuBGIY4RSNnvXLl3km6mVzMT
NaS8dCCCyhKmL62pfOrtxiccwR66byzr88c8TZp/3LSEdqpzj5TkUHRQ0wdffO1DTKJXkL9VPaaH
eA2JEWrAu1fsM49zDhGC0nA2Xxc8ilP02HS5xH38z5eh3+/AvVqrWYhUFFXyF0/GGRXty46s3dZZ
pkcoGFB+Bdyl4kpi+xBbwH8SY/IEp20gbXyhph5m/jhNc0Ciwuq91N6AKfpItIzfc03XKP0CL7bm
YYyAJf3qc2iv8GFyLhdHJwg0n7nUd2Pp+P3obh2dZ8Quz2/KlZzNYNuXBCa8D69Td05Axogz5wGy
tSu2xKGuCdez/j9jxuYe325aXLgg3kjKxOAEmI/i6mNVJ7pbTxJhIb1SNk5Gfd+G/dRPZFpItwbd
MRfwJFJFHcWdQy1e6xshnjZsiKBv/j27yG5cZrzMFa1U3kTKTpQZUNwkJVwWYEJnLTcQHxmuRS8/
Ikv0D1JhUoS7Sh02dGazpGiARxdCSQS65KeeO0jR0ODXVBbcqB5SNQ+J/GJ4ekvZip93MsqY765a
+9S1YKBP6jaHpsPOo/Ed4qF2LxymQ1o+32F3yl7OUCrbxX0oHnhWnUXwfucOoN+WjTiAB6m6se+v
TBBtUeyz183nQofrjpdWy4xsy47qV9LeP99UX+RZSl1cg3e2VXgAR3duCRD72uy9NpUZ5ydout6u
Ag+TweTFyyOLc7cZe5qtqtnr0LgE6Nq4JhnP53G1SN0wfL8ogJ3E7JusHp0LML17vpmg9MaB5s1x
LxZo2qb8lreG5iJqqXxi1Q1x/DqgzOKotavOY83tylXLvPFs9SFN0/2Neu8CsORMDseYPs2eRY8m
Cb5zHDzQX9C/URl1Xhd6cD8gnaQ7DGZtajMISFYYA60m/JkrlAizf74Xuhm0/JTXYTloby0xetth
SlPnSvGhYKwqbbpxtTPxxk4Y/R6vpbRxnvD4cX4IwSi+zfAorkEbecBQDp0TrRUOT7TDQ2WWWnBb
XJfFSf25Xw7NDhsUSVH2mLOBwVCG0NUbGDk+pojZ0eg2+mhMhpvOSAr0QyKE/7qbLH5EgjXr8aa1
2gteTy+jmRROGuZHdwuzmu7W1Aqz6teAoWWIVsZN5/T9szQUVk8CviHFbNb3gwxkbsqCcbGCfkkw
Qzp7i0ljREobXTYSlVRcW9SBUPF88tTm1Cikse9D7JKmsnAyh/vBEY1pG6eJVYM21iH8zWhvLfll
Gz2CsvKkkqV77CckD/bcHURdIRKwz2SPpZUTj4OKqedGBqkB1huujRiAGbEutazdOh2iW8U8xyRs
h4OcpAh7qp3XM4CWHozqxstI3jY08aqCrnJR5xbBza7I9wuW7bsPJ/gGgTSUgYky9yqW4XnFCuDy
DMaZ43Q9nHpjx2mLBNWumkYwf09lNycqTXKRidXTwCnQeoTEZ+qxVLi5HhEuQ/UDY9ikKld1zahc
Ce1f/3rbzbf8p5gg1FNsBtWUsrII5qMV03MZZFkc/9ksdAoSD5XAbTuO7qEqh7pcuC7IW+bHbp4V
yqTbmC09mMxBA+Bd26FteGQD2cGdZWBaGKxJ5O8pnRFdXNOIvifs0He0bshyBF11ep5l6H0emojm
fjrvR3gfqUEK8qlOXPdUkSzIJ1LuUms63FNAHtigcAZ4zJs5URhpYX2HZPqRghZKRl+Bgbkvmjrk
ivD+X1njEn/M0tQDRa71Usl2CIgWyC6svYi88v7nhkmyCv0/oltZBAq2LZs6P1E47NoSIZquif5K
RDGBTB4x3Fe1SVjGQZuUaQq7yG/Xr9/33gZxP5fOICGK2cLPnCihZibS9WWA9Z0pex7JnvErgjc8
aVPaEVAPYF1z0QeayIJy1+0xm96qrfl89GswdiWS10B07raQJgcj6gc4F/ahCspVfTrpBLzk5njV
VyS6MoIsA7Gjvilyaoqz/uFZrtlhLgHiky6cf93iB998NXPMoegQ2aIYSap+pWN3fMGLwon05Msq
e3PMXoAWYnvDfUP45aNIIBQ68QA0s0Ia2r/A1IdJYwOSdeVF/p9JGIZXHP60MmIPQJRqp4Dsvb7v
ys2Btp1Cw0xcd8JfDB70Yg5zFi971GNGt4cZvQYsaZPQrKsJSIRECbS+tcQWt1UX4YMd4YEo+LG+
Yz5yXbYCl8ooo8Ng98AHmhlx4RRMmu5tTcpPk92F3C6p89HUNpdH/VLuee8m59ekbKlLk6ihOF13
hXG3Dv1fsKLX20B6vUdCbgyY9SQuP6SPHAOO4OE2HTBipaOCjyjeiOqMsWruocGYGZnrZJzE8yP7
G1Q5hesfQoXGPQLN/xQn+ILn4UKqTjoSDco/B7ZRK4q9sch/tZd/wPyIVHnWkm74VqosMvWdGdT2
w+jxOVcNOtvQWVEFW0xIlKfMVekcqjB1yIKPu/HjA93nQep5+SV1gjR6JxhNoYZWGHJWdAgifRc7
aOLSZaNp6b3ZR0kMMLgDQeCf2bqTk8/1R9xohfstEyYHrpcIUfh5MrZNlls/xGqYTRD1/S39QLW+
BHGpxiKoJgDsFiDWcgrKffT8284FxlksdA9mnZV2cjzzB42d6U1+rl57rlksGDIvXGrOGLapnS5c
rqsBxHw2Ot6s1gQ5U2bx7FMKnEGaC7ZaC+zh34aDvrpBk3zzMgQhk5RXl4AM9T7W78Ng5Wp50KkE
0VMJ9budsTJsuaGJO+m1LzcDPquMD7vK+EiIMyH0LTCP6qTtCMQW+od5G36SXXxIZxSXgS/MspPr
q8d99MnrlgKuaV6jtvbcuH8SX0E89Kz4SEAk/2YRuyO4fBYwbUFYA9ERtoR19g82LaQkrAKcTWwp
8dmR0xKcCXccz/6ahtLGGvKPXlic9XO/rXZzpo6SieCb5vfcR87KwiCv1gOvY1ayH2d1lpR19Xjd
3XzgqRvGlbvyLlLJhXuv41t1UfZd2fIZvPZGx4fDWWbw8W34EUgp3kmaXvayPJGDH+VbzKLCm89k
+rHKRrniP2I75KZUHRA2Q/hIzXO5oj+syQ0u4d4laWWgIRjx1K0APW0mtZveJHE59GPnQ8jw+DGH
csHpY/uaEN7xmIOMdxpIrs0y+dgxJzOFlOjnpVmxvUEJtCt+Q0t8cWL9upu/ZOKzbzfpS/vHmaSN
houO5B7yAoFiiXHK42EUGivO2YDnJ4EZlWLQSzllyaZDPcZecIbyctyXcjVCeiWhyK4mSdIoUWKv
ncSLAK13KvxPhX1iuwOP5CdJ/aZ+62elZa3AtCHi4hzKMe3ogedXkbAm760mlvaaiweZzLBgX2gQ
DRc1vRE2hhxoWtQsSz1lr0mx/xiQ7mxjGtXO5i++e6Xc1gL6o+aSx6Dw9LoY/NdDRotm3hXZXuO6
yIhqUOtXnLNINdfxZAtM5gi/4CZwyQ4g5+UtF3bB44WwRgF/TenQy3HQ0P2ft3EkqubA8DLr+Zx9
2IPlK6cijj5XQ7OJDAdl04iK43MSMN9K6A274690Sfig8COIkFwIX2TYgbHE+TC8Eh1YTa01WAw5
gBD3LmjAC0QVrOixHxZiVw7/O4HbqR9TMYPGAnaxNzO1OOEuHLzZ2W5D9n+U8qN4HnAyZO6B9Tw5
UWXTsROccFAYtoAJlUFdn4yTcLl7T/vzU7Cfx5pnAcq+Fnxc/KhAwu8UX+536kunDEbC6blwrwIC
fojyga8ht4/SbJXYdUlEuRCpW3QUa6Akfyyct6UWisU55S3Vi30uNdZI6h2lrYYuo1qXa4nijacl
NDGTZ5wU9ANCeUL79NEQjGs7K6TIlnpp1/iculTerxY5grXHakDYCTpswOfj5smE3k4US2Yk/IaN
ijSG2qWtPjOhSPKHqVpylzAwgrrWueeIU4V/MSZ/k/QXkdtyDFXjeYCeVSjnbD48VLMl8RLlKdYK
/VEQZ7PpTpalrH2/rUoYVRi6WJLK2CCtgKKn1yrL8b4CEBBo/+rjXdARwPih4IAQXVmmJQI6QhCK
yLZN0MEZpe+NCMMPvLbVa+f08uPyuisCiD3p2tQe4eigPMjVAx8bVr7w6QuDXPM8zTtObh0UBsYP
Mpwqc5PoKZKcFT26a1pUtpgUddkFt7o7OWnnaCEf1o4fF600M7Yega0/90ftugha9YNB6RpDpJL0
Mk7Lbk9x44q+SQs2wQW7+KsvyL6gXIFTylvS2RIBPmbfsMcrZecAbYvI/bv38W20/cEbqrwXOhw2
MscCBMiOD3UoPAtY3SiX3Ab/ZdyB/mb9C6NLvs7iCxQkhUDGglpJP16XUvDTTc2fxHpP1DxhtJDm
h538seG5IkL0L6FghVdMwldtv2Ipb/ZITl6ID1HgFyr68e+dLjw2z3VoNnh5VhAGKgB1NsMUO6Uk
b/kBoeJSUT7dRYvMJID2mXbcetMX/iDlF1zbQu/cKGGdmUf+L7XcBx/QOQKBpwGP/LiAI80Nf+dA
+5fRyNoAvLu2LQjMSzfZ9YglkEkAYORVsFM7OGSm0QfjS3o4ruGPNQJ5sOUuG650BB7QaOG20y7i
K+rE/4nHZgNpeDMHKpZDzAiwezsR+hHrkytUyi2ku6fkGnPC3PIsdiTwqzokrzQt4LNaXKRj6Kgl
bFKmKzVuQoGZ8DIVPJPo/BN9h2q3redqNNoWi0Vp9VGNyyyFG7bRkKD2YJaDjJGFUCUAf5b2hZ6v
KjhKREPXHxPI6gLsvpil0yGzrFN5nEbhPJX5d1Quz5kTMtG4R9rdYIXraNfNW9NuKDYfD/YKTDE1
JEnimRSwoghryPnTi4yGacUVqyqOYAouR4y0Cfm3Ikyu46tPZ14pem5DgidyEdMEaT7HKxFL1Db7
IjRXEFjma/IYj4V+Nszwf5XSr/7YB8eSDspqnQGoMIWqc/FdG3duEc1emUF1ogEz9X+cYiQhmLyI
bY4P1xmJPHD0UU6/4085YRdZvzdjtZqhzx20vpOeIpoFksMWDIPDB7+SK8r4bYBl/yhpqh7xXIpU
eO4Q46t4sr18UFlU//Xvws0pzgzgWC+84BoT1UDdeevI4HWYzslOsWF+j9QEF5O5z6bULCCSYEXX
9SsMAhUi93aMvCMGJ3E7ppMs4uWnqNLc/AhWTTfoeumW8HTpCiSLScOV6la6pzquZPIbdt1F6Gtf
/Dd+qbQcmW6tXXmkySOCx641BCukMMtc5VGlliq2We9Blx932JIhhVbi0iuvPTWcF3daft77J6lx
icG9ZAa48DawjV2cv3UWEvu0Rk/P1RgYGA6wydn5BPVVSLE6djDSylXx3ppHsL8fcUtVS6MyKsNx
f7LP2eMvVeyRTyRP+S7G8dbvxZpmEx3rOHhwt2eGgcCXTiR+s1n3KPhPQ0nZS3sSnUahf2ATT5d7
Xzps5kl3M+hrHCgP1wliot5MD/6ycUXJG8vfRAgOGR70o+mxe0sUYl6fSdJWUVcfw7E1oNSJVs/k
GI8A2MUj4/ceQLv8jzJ1r+lhSxdIE3uVCICegtFTZHStyA9sedWoYDH2F/noQU9ylfiFunp7eCFm
rVoQSk2X2kTXW/RXcSR+hbF+dOyU7R8t3FGA9zQYPcwmK8c8XxM92tDlQ1fcFygmDqQfSz5A5rxi
1rWcA3Qbq38+K9qWDJg/y2vYIno4/wBJRO3fBRen0T1/2jjBBGvhOqBaqbcfmn/q+lp/qTiOmoMP
+Bypy38VRtudhRk94EeLsYEhWib1qY2w8PaFLPyz3Kscqc72+NKkN7iV21SVEdVUdwA6rQBxJOhj
ahrrrVus8QKOcEcvE9JUp1Ri5i2p9kB5Xn2mRC6z+SkwkW0V57LFcgvTpKDOrHNe1b8ipm+AIUYh
ZMr3YouuUmhkbFxlOD7CdqaEGbAVgoGKRlRArDPvYrESvM052tiTsG9vyO3zxBT+3DBku1PXote5
DHbK8xekQT8xWrBnP/AhLBFM5KoeUq94EU6rlh1XcCcjYTkUl5SoBcIGNN57sW/K76MN0IF7V+Op
TNIa7vulJH1coWmUNJ9hNLY2ckHMX+KcYJfgptn3bJDovKOyDp5b1m81JBCp4uLJtGZY9SFMr0io
5loGFFBYgtebotRcdNXRvhU3ycu1SHjfRyN6SrX7Pyg8txEIr40w09/yv6bbB8ExFW5P/OK4eA9I
4xgoNh/IIW9pc01UesAZa6J4QHWzQc1lJ9D6Y+oLkapgD476BrFOxA4x0TWYSKSaQFWFMLzZ0d/+
znXg7XL/Hf66o/R4knsHyzEnbgItVhLNaVAMIhUNwP6Lc1I5Affdw1ILuAcEaKXMIr8aoRodwpdJ
c40/XhR3fOGcnROQeEqtMkYJulnWomCXlAdq8Kg/rccZL4p8UQs2h0VE/xtoQO4XdCFUatf/ZRFK
l7Qd6eboSorI45No+iUS7botrW2+MTLzsNlZ1wcbfYhQVe2we7VYPSwiIT72b3lWKuohANs1O4TL
7K/1y/WwZIECLnM9K3XsoDW+IwHJFSH6h4VyLpwO+7Zs6/LK4+OqcMmlipsNC+oav5HTbsbmlL3C
dL7sExXTeOsK7UpRPIfgPJrF3DJDcuY2Sqb855XXbEQE7Tbkj8c/huunKVXSyDlN1GiOdCpnX+O6
56RoubG37NFhkB+GSN8EKf7x7FhnoIU1XB0r7WvDOtwOjzijX71pkeDkbMJcf0Cauzxx+ssXhnjn
hac4CaLxxbTVjaFdXdxSWmi7ydXlSxCDPbaPqNswsuNwxcfsjiHxOCW9dAZosOnCaXfMfXWLhkM2
TnPuAh+a03VF9xsUD2Urc3WvNopYAp406cwjGR+RC/tNGSVVEC4lZvEKhFAPtkz3DtrD7K4ErV+Z
dUV0t/ALTWGv28k340gY1n5vKiIP5FQ1b/q32HtotnxyasUb0NoIRA8rCnH7Cnon9wpxq8hJahst
l9CDvFjdmDU03RURM5G+7BODvd4of3H+Mn6EFRZkKySmUw6hDwvMBi2KASYyg7W0r5K79Vb2IgSM
wAtP7b6H7lXMyPm1VFdDj0gd9tRhXYrgHqtT2VviImrlpxRrFpif4NO5TIujikZF/pjONtX4cPyT
VsKhowt2bZOTo3VSYNIcb5ynJZivbFOfTU6hdzne61BtD/juR0bm0xPf/xpFD3ttJQDuAnquGUdH
Hm+RAnJK2Z5pXJoNqx1gEdDwOzG4rupjbykZwKzjSgi5Quc4//ea13jo+BYtGB/vAxBD/I4J5jB4
bk97j5XidBaErw+jaqrXL0rjx2Upx8U/W2WbifzqnRta3Lk6JIby8r9uzPcy4XSgSsSkJtyrNrYf
eXNO+3OdyZKtFy4z5y+I48lHdU2KCFFJ9qbR7MoC9dw2lBRWQ9VQiBS5Hor/OIF0L4V0AHZXC9lG
I0oKoqaJpovrP9rGURV7ZuigzP/vBhHN7MrRGz+Qr17Vk5K74b1+0pA79fL6hZJDV0fjA7/DG1QJ
wmUCWh4Osy+k2MMqsqTvjh5sHMT90AGacp+lIuM0q/TGQ5k2cVqdi7QjAYN5TYGHSM67iwYnAH+5
SSU/Twv1k1hfKNResaHtkNmOBXBgWeLsknP9APT+WQGFBdjApUQk2+Wn3mf7gsdFm7pykZJDJikM
rIP2PKyaaECSH8CTWZRhJZT4C3RCKbf68Ux+2LBfP/TqwgQTwadWnlUxTGwlP8jAFomYrKUw0mON
c7laJ1q4UhbzAdoSO0KAUmC4PrZ4Q1BUv8604AZOd6F/+DrMF4A1uUPMlvvLlC5yEneXvmR+G0Q+
yf5pRUULUJVbiL0Aizbzm52v9TL1OULqDcgWsKq5IUxWavDU4nTrkToGksUp7lquLeYeo/Gq2R3g
PBZYFglhWy0Y3EJxeY0qHuUSGWBdK1CRX16iB/hyQDP3pm6jJQgGUurrz4cxC5F/RGAdmA3pRUdv
iTsIxFZQhhftSO6QTjbw1YEF1guqjnFjWQg+vKtWFwdbkYHf7aLrRtFcUo7xqH+1REWQwT218n9p
qrEGEUTd8QLkTuvHDKqObsWm1Zyt90P7aBZRvWNxur9XO/p+IFRU1PMSRgNZGw9vM9haM/jmmGeM
hhT7K7aDlHNh2B33gUEs0KgB3v66nz39IzeJTHH+cTC7Ym2WQGC5XzoGI/cY8J7AjqJPOPq3FKlf
TjyCe0kOQaseFeDmISyc6jjcgAj6KjwN/wWvxzITimRBkxz5IyctR15OIMXxCJYmP5nbHWgLHUyC
VZH4iC2X8yLrEq0bkHZ4AFOBIK303rUeSZBws5+YQTH3BLthTewVd+euOg/zdtNZvY9V7NJu+kHw
dbuzIn9OJpIe8RJ7BISgJzOWZ6Bk0lKUhJzkBKoyCYLHWLvdVqPfqKSJLjfaB1a4GDWmGQ/JPz6W
ltzm2l+1fBuJQioQ02FKKzEdqfUjydln3rsStF5PvH+QfkyPYESJe/UJUjJd4p4RShD67aDfMerJ
tQvMt29VGAIK05Mmzm3EOhg4zVtyOpqQT+rNgX9/MRizl8AEci18TA5Akfhri4FiMse+/oiuu0tO
SLj6eO24Z+4203mrDAlFTsErrG+eMJPrZoMbuNyI6nKFoN9eNi5WfKahXpP3JBGDBK8WWFg9y+7a
l/nE8rObyCZsu48nQeWNG5SaPCd1ZKGklDGP2yo92p/9dAi/f9FpAEfOmOqBwkCc81okRaqwm8pJ
PFS1thYLGbxX4+wR72dxuUCIPUVD9o9fai49obbJNTB2X9aUpMVKfraV+ej8BFUuQCphK7MIrAA4
djHvVPqZ9ikObWqLXwDdvcTQvjsvsE7stmFlP+iDeBHIRTDC/APQ5xd1n7JlPTcweqD5uV1A3Tyy
lzNBsWuX4hMc6cv+44mOFalHYRIUgaT+5Z6gxGfZlANvy7fySK+U2dMoSXgMZwu/mDZ+tysyV4/a
t6fj7DvEsoAnS4H16vV3AU+HIBbo1kDpo08xxO2yobcyFrW4tygh9eHk0QcXAjdu7EDxJ+hFO2ZA
yDmDU7y0e7nKGqY2/2MNr70UUtOEC0uVZUJjisVfbS6q/2iZV6MsW4Ji+AR343DeAC/z0y4/ASic
z7iLgQjllzxxbhYT/V6h0wvHqJgeRu/36f1XtoTrOYamb79+9EY8NfJIqTscFe+DXDtSOOSGOUQZ
QZtCZPacN+Wmzk+9BqRNwcarJpVu+yIzIte80mYI/Ff5mZIuUslg5JZlp1XfNtWEXnXfoGehD21Z
xqoNiu8ycymPNwnvYQr3YX3hDLR6vFZJzY06k83pBcGSm+alHt1XcuJ+W3NGeJhh/gUIz4C1p0uF
OGEgJIoFuDFJjeXmJfb5AEJ+2sFP7hTPd7VN+xkVMilfPCD7vBeljRC/4YtrWdJCFZoqZgwhN3Sb
14P/KbqCv5i139lZ+5o5bRSaans8s7j45wXUcXcGJNQpqJEUS3dmck3GFaRTky9bzEgsCkt8/sbI
XkRS9gVQrK1tPTwTVUQCpxZiGp7oueK9TM3DXqSDMb0pelxCxtNvYn0pf8P/BK94m6fLv8kObVN0
vrMpr8mD4iDJfAIk0jSZ69tY6xt6ePt8ladWxzkGRB5LlHm1eL9xjadm2U5qNukntbteH4JdVQt+
wfyfYNMN62Ge4Q7NliieUQZiv9ILxnlyBE2nmwWEaixkYWT2G4j2tDQDUwdEct12EUs2+PgcQom/
yKTSlBr6vKpgNm8i6aj025X5JmJCSHNhlDHUqSS3OPTyAn1zgXj0aL4PkpPME0dg2HOTGm1q1NL7
I4ixEmxQQ2TvdL5c9Idu9L26w8XfZ5v6Q/hdIZaaOUIuv81rlrJnR/Gxlvo+uifiOey4PaoU/++n
dV+BBGiiza5m5ripL7TWXnOJdogGcMj979JhI2P1eHE1q0CvJxByPxIT0ChM6brckcgRcbKy0Gkp
5a3OE2nSxIQlNcsHbdHHxonf6lvgC8awT443bfTmYvbPtjtthdYmiz5bced/NkbdYBm+BW3DvqwA
uhFrilPAWiNaQsQeJlfxODlF/FPvuiFr2deJFV9Wxt98S5cB9rKrkZ+u/gx2RdsO/2lmJ+zDnInI
TJJkPWtAUKY580nEx6MSmWnFP8kLjOBWHnayauNsaAhRWTfdEO/uzSLzb+LVvxTTn61HRLN+rg6B
H/8JfCmV5npby6t2hczMQBxchB3/VmgLcZMRw4yhEp5OcGY8jBkewmrT7V+NsSB5uO3+uvM4va9w
beQGwmzu/aygDlKD3tpHQ+xtmkWyRjxSdrMcxkadvQfYePS0kcG63tqc6euNeF1oqLWmnswQSOCA
7LxhuH9cV/S9lIcs/KtwwStnQdK/i/yM5bSWcoMGp34fU6+un8CaXUuKmwvJGqfMfguZ+ACmRNDU
XsHSG3zR/Sib0ZaSO3jCczaWOjiIpcyc1QXu78wJ4dljXeNaLl4kfzHWW2fCvl6ybDoNDiVWseaf
9z3D83ebntEDqUxHu65P9V68OCaXHJ1k+HRLiq4l27sXAQAHQIkbex/S62oFsVFmelRvwnmPrs5C
wTqKi4Cm0qW7gcKjEOqqmvPxzm7iygzkhWJc3z9WNBPmr6BT3TZsYYTESXqoytgAHih7TfV4yNF1
hIzN3PgVHjCgn4NHYcS998aDc2UxoJ1dTfy/I51HI4IRcNyOxOhmy5VeAg6FijWBAzyFhvfof+Sy
0acvTHhH36Cr5DAEhfZgBt1s4DvjTqL1utDutEjF13t7mKiEP/OYJozBJ66hC8F1e5vOzIyTsipj
jZx8AH/MJHS/SoDc1n6uvKIpuPxZWFZPoBbxxDrYScpffOGLVfBFNrZzF5HLY8YBwjnsLeauT46m
4YKyCOVcLNMgN56iQpbcWUj9Hip6NbZ6QqVEM/rAlMBJDQd6MEn+pIayUgJV1Hkp9OqrCKQ7nDrh
eBGnUPXQVA8kqw/87b8PzWORXLciiENlK86KeeVdqwqrOju6hJq3yqUCxbrTwmYmC+xLFUkRrQ+Y
PM8g/nKi/InXd/XB1PvFncssVvVU2lmUlM2RXfdu7pM3w4nJd7C2BwYheEQrec2BMfHQG1fxuOK8
cOkogw2HEB0Jvo6ozn/LcJ2A7KyCT8P0FmKCWlAz2JyU9Q40cNBjq617MQ+qLxcJBLbCSwETX8p6
LRO0LCB7tYfekTmvGThsxPABpTTd/nYtEpOMy5DG8DFGWxt0DUoaFtDbU1pseO3ll83ctYklVWH6
wy+yJXy1H26vzcgHIcU40WcJPL2M8yiNAzsWL8qLVQEWrrgQNnaU4aSK9OW9svE0wM9YSM34Tp2M
jHwJpngruDyxdQXr+TVYwJshbXNFoFXqEaHFKpsk9QrIoe0Kwyy87fVHoQNpkrQ7uj3p3ggqhVuT
TlMe+WVR8lUn8nIxIeHpqSuX061q8T+tq+o9T07fck+r3e0U9JbDqizvtSwPGpmmk6/sLRCds6Vv
ArOG5p3wbHOZa6zAlGMk7YjyG/FxV3n/9RttkoYMOsLwVWRHHi8+Kp2fEGjDaZfgRuNJtYJ+rmp1
o1k136ETHMl/5oZKN//nJQiFJD/09OLI92JNxf0Ya+tGOJjUz06plXEVAwSQTlA0IL3TC4UvFVk9
ZVNEdYRt9oc76qgLv7aJOyVqkqWJ5folnmkMrmSjVD4qL8jgql3SMWzw3b6EjEXG1lb5Zg6VUp6I
tvvLSuAmvnw/aBJ6wquSRGiUSuiynO95sZizUOcFCTTbH24KBqpnjaMP8bCQIsT8SQF9l4A2rPh5
s066ONdgRr7IdNesp/w8eVHaweDreB0ZJ9OS7JMUu5UhWqdoxiOoi+aiB7Tb+e6sFXLjZi0SCI+p
p2nRHsbNLrOtlGAIpEWG2gl/S2LDcNUwX+hNNo2nia4nVK/plxZj76wvrm274fO/2S+FyBX2Dyri
JuzuAK8vWjiNTcYtSKAjX5U0lZL7VPn60r0avuv2klRNyZhuV2N4Lcgt/S24sTZjQpWOVjdMur5T
yj+6PgL6uCdtDMRkKEVoVPyKZ8b+FhUkvaZNQ0PdPtEoePhPv0xhwBb64HDDut6OkD1iUMWOHuFu
JHqxftzmExsU823Gbyg7MCwlTmem5O5CVmSVIm1rIy0HF8IeS0fkPkN6XIIFlEKy4jV4KbaPuIIY
hDaRRn934Wee+qinjrYlCqjoN2W5exHAzf7um7Md+/F8MYCyAvrBBrsG03+8ZuoZsZmJu0BwjwEb
htjGQs9FgGr3K1xV+E6e2skPtqbCbIgEzOP2+FrQNob21JkHsn/ONSs0S6ju84wqocxIY0idGVCw
YLHfiNVQeXnWWNGOL4ITmlT6ogYZIBC0APePMh9dbt38JH+1D6TYjBD7keJgBcYbyun/q+hLk+Kh
TmB6bYaK2nCryatrs1BxuTVoMK+JLNl9vZJwdPoyuAbMHZ0Gn5PKeNq2xa+ZXPXD+upXf3eowNxd
n3kZUkrxevcliECF9lV4KbQ1fJ88hNPowTUJVxfsj7J3oPsZ4+msVas1eu3R9QOTGRvByu2LSZ6S
ZPpC5QOUVRis/5nccfzgesZxbem+FVScJQv1bZdOkjkkRESscb5fAW44V9nR54tX3jcV7Stl3GRD
mFG+5J3QArLGa+4I5QFsA235233xrjQ2QJGtz5nLpjRIoSO0u+rCkvh/xW/beAxa91LlJYI0ifhi
S0vHbT00RrZByVEm1oTewaLOK4N2JGhYBwBHhpZblt8DrxhvnXuzpQH/xKUcUrV+sgFZ38tQ20I4
IeeEh9gCjg/ssodaPBmyGCjszGiM+XFgBPLBQuMMO4ThcQyFA46lFN7QMoXdpOmIgPlGzoHQfug5
RY8sZ1pNd1uDPEq2wI8nNv5eV3oefRqre1dYYKGYinVrgnBC0Wr4g4EXUt6qlez4VZN5AjEp/2gg
64Rl3Q4psFz3WFINH9fHsLwjpptrkJx4d4VLVsQkshEl4xm2fSgNX2xq71wBlUhwF91UA4uM7nGI
gd+Z9AVKrk+C9sQrqeoxVhz3KX7zBttsbs08W9wbvCPBqW8WbA/XE6d+25pUVO44hWwjiSN/8vZj
gLnsuZ156WrAtgjqE9WAkI0oEqLR8FnpQecwP39hyOYOWUXFLqc3OeSfwAWbIUdjW2tKTY2dC+SW
g63YXMEZox3W8Ib1nZQLQeevyBgIpIT7QYDXXFYDOOjqeiV/n3lVfPEzeXrFgRPaOS0f7Lloxu1g
DUUSiP/+b5oWtyCcG/gpt4r6Tgc7BTgnA0LnuhqbGytzQdran/SqFEoNx7lb4HnRIDsLQ5hSGmj0
Ssi3J8UFbIJukrcjMHVkPI++gYgQN0UnQygvj4F6uyodbHVhRxhtvl7cWv1+xfDfn6aPcH359V3v
hmzCRiwpgrtUowUQqUzRc4ucdqOS/1KuKevT/EJhQEguc6uV5zilGhMP8u4+9aKLTwKvetF4EyUu
YHkuD+ZLwvcpi1xI5LcPaZTxUc4dWZapVKv4/cMKgT72qpA0dywxkSqVeOxShekOZe3DTKxF0cW5
wgo8u1KyIrFv3XLlGqRPoFgE5R/9tJC+YzoGFaLUhFM9/Sm37dGZJtHjJFEiBXsVy34+RA7IV2WG
hLAAObURvY9LNEG1W8DhQWe3zJkm/oWhcGB5ixhYR16BW7AwHLl7aZJR3R0M8reFyaRYkQZGfxea
OjqM5Ls3L6fRhi589yXK4E8ypMXFTHUBN6S69URVt+uyYZYQmSF1IsI1x1Zr6C6D2fF1Nq5qoclg
EJAJUue9Vgt3hBdTZxCPbgyEo6zBdB138kBA/LpLNbSavuqCOX8CydttGY55hI/4+8J2UEQHUW03
I4/3G9wJiR/dZl8Qk6wobNc35AgSqTQUIBbxWTjKAxaUniZBiix8DeHXxtjkb8qF9vWmC9e08vbW
lHUe6xDELNUtx2uOfQEruVjSDinjur94xqjDiLzUouRECb2JpU3DGfCnOZXR7j+HFD18bE9qb3xW
nRyXkM+L0aNG1xdbniIwTAaNSjefOD3r5iyPlfCaqvrPwu6G+HFLDDW3Gni45EpMSk2jyPJfDuGx
xT9fFAtlfIHALPNGMCUiB6CnyNfcn4HbC50IgsXMBgwIjqzSWme1z2SH2lERl9jFTNrGohbIWt4W
ADcPm7fAfmwVfiusRmtLTd1Z/zTQZYlcrgT2TENDYaV2Oc7mKRW7ZP+/TJwwqb9fq9glTeikKYIn
ldTsrzAxX1oSghdcD8BzEWlS67irBrPgHkQeeEOBhts4c340yJ7woZXSbTYxSefcshwGy2GmijVZ
WBbxxAd9saOg3S1w8zCcK0AtvSevP7K7VpCakSDzaffRckVTV+ILM6C8xobcf3YQAVqdZSoBYrPl
9gzUAEdccizJ4FfDGAmf3VUHtznU7OgaP4hjjo1NQG3fiwUITRi1tpFtv190ol58W3w2f7cjOILy
0UKUOtt6V3ZX8SN2xjuQufoK0MU3eg5/f65v3qshwXXsTMztIDjzNQLmLj3QTKHo3cBFuNWTlxze
ELht5NNb+uZ2uVPRsbAcR4504ZssowUa38BpnG0mzrg8Rd5nY2vc7z4KSDirHx+yxWu7oxBBok+u
k/jP0eJ5lxXatEYTHTuXKm7I2h7nXRQRAlBK3VqgOonmxmtq80z1XKkEtf7kdd7St8o3hSqs6ako
vsBDgxEYH4ETpS0t171/Oi3cP4JH+FDdS0+iXbtuQTclhA8FjvCzIXvgqvGpAAaL5P8sGR9pcGn6
VyPRmkyXOflxBy5vBBLzwEMR6cmkIBHAW1LKdlmn6zW8mtbP7LwCI4EJ9E0u5AqMuVVb43wfN1Zh
aPIjzC6vKr6KvllcdY0yJJmXw6CGfBvB3HjX5/6dhKbGE/rOvhXJ5VtTp/9yNJ6HjWhCSht38N+/
9oQY5D/nt7XXD1iIsBQq9oit0XVYLQBH3ddKU8p6qRFfXRPqggrAHPUrIOvWJTLLZII3Zx9lpIo9
Fxr9/eVDQPgiyoqcTss5B7A+vlREB76KypmRyZjtQ37VctALFwOl+4Zu5MSF1H80sUfZ76zOFrgv
RDJtYxy2CFvWxQw4SRRyQ+L7syalaDO91jvhBHqlpWemrSc4S6WNFAKhZ+Wi0r3qs2zlrhNPFuYa
EEptqvv6H+d5qXT2RTupIeRmHT96gQ4Np1BOLjasuzg5xCKesO+svOp4qZBkn7LKlBupra4EKnKd
tTxYI9gnvKxF55WPd5UUOnfebNqcALT6aONzX3pSWsSKx+UlxEWXlwhouYdksk8D/qtqfzZF2w2f
7bZeD+/HSDMVkRhaLy/MKIOQR+m8iT9UML3IzPwXeQj3tyd2W6k4wo5ZImUgzBTOQo3Q5IHo8EQu
CKqYXt8X2H1XVHKCKkaKO/zgCL62WphNGKw5zFcbfu9FCW+nFTgzJBEdvr6KcqEQd+eoYxtZ6OKl
YZjRit8n+e72vfO3pNW0E/LnxmFIqQQWg5HFwhYG3AoQB8w7CrKYUlZLbQv+kgEE/PYDxTDWCaBp
Pjlk3nPCV0cipmOCgoc22fcaMFKeva95GsjEwIOfQX+s7HXSHjlYo9knYKoKWiOpbpYquuPVHgrG
/J/K3oe/mHpav+PMHrTeEIFHk1V/hx1ZyWxHYYmbVMYAixCE5rrXUE83kKAQy1wGPpfZGZBR2Vg4
P3rXPBuohMOfi+W9U9wjNeQM/o78kRUpI6AUk0IDkitEGuyBIyO/o78hAYjmqPdlwJV+zyjYeuyG
HQH5dzyE+NYYplbwCIioOqwEIAD1EferXGnzQ0ZZ75mu0EXkTMAVNvdx0GGOGCRYeivu5CWUMVds
EL6U1dsLaKJhWQo/AuymBmfAECvGN8D40TWdHufApWmQ4HRuUHaGxw9BF2RJ++OKzKLfeufAXRXe
QN7UnQ1HBdua591YUINnCQrb7AP4BReI8QmXlLE1yvWQZwxTYPS5MraptdqLRp6xAM+s2/v29eIX
5ZZ+JanDUUbU2QHn3tVEhkAToT7wqVLd7CUCQZVVloe1yeTTldpZKXkvIAz5rObcgqLxiHlplAyS
OGVgh3yKN9O0ft/K/WYqEeST2i7QI5ESivDSgNC+N2Eq4N+d+Xc1VrxXCkQ4koxJdTZNjtIlr9X6
CrL76m5c5ETT9+OZMt/kkD5tftN0agz4CEfCGuuSX4xPdYRur2k/vGGzLiBBf+rI5+o5PXw+LCDG
W3OKxl04TGD0MwxFHUnmXpCPjWQ7cHW1hYuCzMv7gsH00SA33s0+ly3y6Fwz/C9Zsyvbdup2n8v7
bt4EcV8bNYFKMqhneFliVCZwy14/DbmkWpBusAx716H7UmGbRnkkgNL0aF16at9HpU+YmhRU+XUi
DbfOIF3lsMwzgYZOrXpEQHVsrdMaDa+gvi8HflfXK5CA1CnH29WT4TI6XHrxQQy7INNy3RE/G9VU
j9IpVdes4Kk5cXGSkvrGXfWeQ5062gRJbwttdoe4Mhr3s0ZcBPwH4w4fVju4eUtVlkjLpJd7kdee
iVCFF1uvfz7kaIM/SauphDu7qEZuWjtwNfbVwK7VzZR3SUGHPRxfKT4U0jQwk1FQOzY4T/BGHDQv
laeaYJA44spiGb1zTUF6D8YnJQFD+wLoGoAn2w5QTN1BrFrUz0KRkn1wwVGriulhCTeoqZg4u43y
JUd3iZ9/F0IifDsp7Tuj3AUIh473FvZxvFu4Du/USP7L+odvAbI+aDEK2GEaliidFEwH8nDxvMpF
Izayb5ot+G0a0/F5Di5Rv3wnSfhLsAO04/RlfMkXN+lbeBDj+uVGuhi1yrtFZmI+Z7+Be8CVPfDi
Olofp+bpF3QMymTT1iByfuHHV6s0TGObTDIgb5dV+/mKtUbXcELVvtByoNX3Lnw9rjwvsdKV/CQZ
7dV/6ISgtvDOXWPk472yRnqK1ctJegosGPVORlXAyMxEwBLuVgNx74WXYLiT7MVnlAgD0tVrKeAq
utQy3BhIdaBtSaMqe61YXQCTRNERHoM8R2EQGBTaSXdqyXlfou4S+HpG7V9FhTOY16TH3j0TklQ2
7a4uggMsSMcp4+RwmabhSH+t5LFc4CniMhPflKggVN5JsnMD2e6Ym1JIKUv+JIlf+Xkf3kdHSZ0X
P8dMy3aZQTOahD9beM4leFJ4MX5+L3EzHZ4LbJ2rFiNHZuWTCIg+zVqxwf7zbdoxVSfKj8S/0fMa
uCiy0Zx1SeIBJ+QS6VlTPiEx+PZCuJWMtJPKwLoQ/EAE1mlyEzBh1J99LfyiHdV0d84h1lhUky0K
UFPzLokVb7pQBiB9NKI25c2V/JWYKviSlhzPAk5OZA/dES5LhWhCFZlW6cciigAZNUQqGUM/eBma
/EIeAVsDTk1FmFQORhE1MU4hUvu3OIaDZUQpiEzavMso/9Mz2SA60ZfpTd2Lw9RkSXpdsyaDvalB
9QGiBhKbEnzrhT7qAU6m0q3QhHx93W/Q7ERaaEnvR2DydGeZytBgtDLVmeSO+Sf1QemaA6kUtz+F
Orp8EgwVXxK2iyX32jATAeO3JufKTIAdl4ZYu3t/jQ05iFSavMa1gaJdKYPvYTGdQdIRwx6YRNBn
+LiwEkQ6iHDZDF4iwDJMelzB78qBogkrpxdsIFPGX6tuOiPVh0lbVluqWhtZzorGcMdEuPBDypCh
F0fJbwXl490A50FAcdWrlqVEPNGMSomRiQJelxCzdBX9Kc54mMzyFDiLQ6VgxF29vkii92LWunsq
IKA7E/BHa8o46ekw0rncHD0gqC/WETOx1lHc6sfMI3sFOGRJDGqluZz8gb/fhed10kjo8gQKhysy
7C63oPChTCPItdCHUox/+lC0DgM6u4OpcE9ai+r8X/K0avKnhbttKPZuoOI4mqjW/7bP4pvPS8qF
X8QpVQ48Boo7uGwZHERGQDELn3WetFa5XjeBAHmwbNRrgqvgeXVz2PB31iQJnTD6zNdbKSZiShHK
x+Y1CD86uwMq/BXRnXdEAkaBz6DnCKXINhxwyGmGWG1GftQosUlzP7aTjTYbRLHcBv+dqx30unmR
/MHAeG0IsMgQkWt8dE7m4WCJHcqGqOTEkv4VRAOX1/VRQ4c5jHY/C9p4n0CwngQc/LkrGZsJL5yY
xZdBmrcnTyQdYTiHJRFP+wHBFynEObalCUG6uTM6+QQdR/R0xSHbcKUqxNe/2CxeM0wLWUL6Ho0r
qC/7PymOZGwqpCtIqVKeIBrHUjUjDax4I5I0bHmD4/NqGApZlEZGvDC9HeQ4Hdw/qrWoFSZ7oYRU
Dc1n/nebpM2c8/6B93xHgjwJR8bgi3ybmnngmXtGvN4dO7aZBlkhanMgxgGKCGmLq3shHCVvGCGb
XKXdaFfKZlhp9rA+tM1uVLuNmeyPwyLHuIsk67wsANxc6qlZpJ8X4NTcy+0H+xFL2dmjO+47VHnu
Q5f6gk0V3DpgkTDTr4UAkeoTqtout4v+lSVsTKDe/4JTGkKeYQj5X1udtc3jbMr9Sfi+k9nqun/r
exkJswed8JMwZk2QzNuN411OP3GUQIhGhR6WdMIQqXDq9FvwjWLP6u5cRU24+SDNGGiikrcN8AeV
MvLgRkqWseZgO5AcG8N2JspMLIPDgxB48BTnBzN2by53R0CwSgbMrBj30MoVAfQp+ZmpG+a/5cJD
Ky0DjG1aKsl1iZe+jTpiE70n0bTba1Khcf0x7W28qpYPXWqhc+kicdg8np6g3OR58cPeSfavtFMy
55qwcgXulQ0wZtAHNoMsT0g32cgjN5oOTeYLIWbAO7Na/4pEitkBGL3G7SSpIoFAc9HVpKS9FEki
eMgoLjPNTfFVQq5Slo6kK5pgqbyyhjJjj6+kEdcCwZDrQTJSA1YMqLB2OMuToPXPRJ1aUjWGDBOH
lRT45upJXFQMJcepYpPNlhP0rwlnlij5RwJASESdyoKqIDwGgFxxx5b/Cfcn6kgn5ZUK7kNreR50
RknTnMQLHLinj7nRjpvtfvk69iP3HLau8IpLfP4lt/dT1FjpPnDM/I3Vhxu2rBZhEy2TNkRgCaq7
ZWsjgY5GWF6FhMqDcfxZH41hph/eeIE47AhNuEIof1lH5Sx21LNSPxRWMaa8/4rfl8P2hE+YVmGb
wXij4UqifYOEQeUp4jgznXuxEVWX2bK3BoS7u1ZRsjB0uQKcAOCywhnRZrPmyfSOe75EaJUc4695
hhwcdBCquWjFRE16Qmyok51xtzWtz+y5H3V2pYi1927KAORD3abf/PuF24FM+Mc22nG8EfMfmePs
o2TX+VgMv85z+e1ynEUzWB+d41N2stiwC7POg1+U/oHc4CZ+YlMwkY8yb+0GMcSoyTmF62HcUUX2
UPBeVrN/bQT0CtjG4PxfRFZau17rYaVDWNoL2qlMctIhP/g+J++uoEDW2sbiXqxHG3R79uq1FpSY
mmPbpsrVPbVhQasDOkVte7LYILKdxCLMxeFooBJlgz4azeAPx1XOY0AKbYzmzhVInjTqGRSFQ+JH
h8yn4yAa0jMbALu9Zrgq9WFMC38/+2e0kJ92ISBSZ+LQmML6jq7tuYiKNrz73bI193fwcoHwv7+z
u9v7bcs59wll3S60RBGpEfgf7xq46mG1glO6+cAECP0wh+cuJAOFcajYPj7mdv2ZchpR1oMXJ0y2
URzRFsmLXdDRQyhzGqz/HZcotRdPZFhSH1NHaV6uF3UNKJ+FC8ayqZzk8/AZpY/hMCSXS2sOsH10
19nHMKeDByFhoCCi0ZQaTmgtVerFFS/dp0QWijjYbhLts2XofkGmcvRVdY4Is/cC3senlf0/MRhD
hzDqVuOvvvSKuw3rkZXfsze3OBN+fu+eCk+cTOHIgmhYBcRfJNIHqOuK8gTUJXKzFkv6TEcbcHHT
Shw/2L2PRCQtZk24+N7tRm2RWDI8bEZek9RZnO9PUCQN66DYcKvxERDilIADq9DxjpwrEIToK0o+
OPGXEpFWl4qnDxM8tsD0fgDIWU4icBmEFn0kzwtj2/NiYP1cRrFGAXMoXfFmmER0KfY3XBecp4Oa
UCViVNSWWzCPN6QRdkxtn+bRZZzmeOMXSS3GTFy+P9zCmFtTITkAFb1TNLtboXia4vvgNi5IkGdR
4U7xKlRh5OsoSdwV9ArB52FOmFkpNBduEpRIOvo1dNfacWNhCE3N/5c0iNJ2mdpYmJ+8uzEcTKXZ
69AAmL/qhsBueFAPU4GbzmJJSvEaVjb59hB9GPk9HHzyfGv0tEgHZWVlP4/ts/a4tWFHOJU9o7xw
TFwZvars4qaPHQW8Wx9HLTQQ+kR7RjB9GDfjimCrZ/UG3dKAx5dFBfuZvTNUvbVPtOBbkT7GETyq
W4pg+ljWj4lG2Dl5tinTUxEWPXt/Q5rH+omG+7rvYb9lc2aH8SVCR8FVUyMKDbweGhWxvRXVwSvV
s0/zD9A/aSy0Imp3I5pCbJ8PtoU73bFdcEHKBytij56qeL+p13DIe2lm+gLLIFMF9jMfyN5GFKMs
l6+5uMRGoIMWTH6UvsEyz0s992YRPiQ8K6Jov07RAXtTMjJxq4gJRYe9f2nFtUW/WwuUwOiozQPd
foOLV7jcvdQBE/iKeokjRYCKe8+HDcFhiTDppzzXk9+1LDWvKnT5tyztpaVc750r6ADzlDL+UKJl
BQO2iYu8JZ3IRyCoQzsi8Z0Xcn1MAhZwqfyyX60qW+yViqxgb1qybWErg2rmYJk0aYBmw40mm4pg
PVEjip6828xklkftYXM2m/1hKKx1NTVQ9jwRfUJmeRXZRHtHoIKE4s+xXoyPu9QpUuec0Q2ir/H4
ZNemdjw0txAvsadDJuTcMAgZHQe9orp8GK8DUxjq8yG3bJeLACYdG7QJLwcjYA85WOclDx/UfTcU
rxJCl1cADZuBQD2+Hg/6adZJcWY8ZHM3Ct/oPh+cLh9e+nTfvWmz2QYeXeL5LVpFkQEn60hG4Jx0
+jCbv1nieUbavchAKPzWF+KQwnPcCpeZJ2PfjcPArLhSoi7yfkgWJAWTflBflNWh+fJPSSrXwFyq
WJXLWZYTKcNeZFBv3FXNcDzhQJJdCxvNBRiMaCjgPwpBpCjJUFCsc2xF3vxD6nMrbdf8zRqNj34t
+cNeag4aBfhOzs1BMQDbRQRJx5ugXDJQtNRue5HoozIzsKdu7k8sDAsh4Aqrx7JJePHIAdzTEGle
lmWFiRMJa4QS0vpGfypCzqlcxZ901pQOkPUl33TW75WylBOOOzUKiGhTdeQuB99+c6Km9aaaInxh
g+bOhCFBPRGMaggwa35uXVgsTO3mrPRd3OTUFpOasPQLTSEtEq2YdzbOMnQkDIrVl2Z+KOfIYmgY
EKJzNup/wPAHFM2lovkm9ISPCjFFRkAQKefdFOuvvi9kCRPjvfl45SB+Mt8Qo+oqrvoTBh1dl2Vv
bDuJwtP78InQ8F1BBbcRXJUQNLs8Tck6gMGtK2rjGr1Rfi6oQQQyudMUiXzygYwSIZNBscQYRShw
vzB+JYwcQbUg/6S/4IMyskA+RGl7M8f6kWYpECTGu6qyJR9ay6dnqSScW+aOWGY6QPnI2vAydjxr
9vKb0uakLeGfe54i/T/kjvKEB0j55jv8XWG096xvev8BjdRhohhR9AAOcKQs995PDHvs8ecwbeNA
iU0T1R4Vm4gvNMXS06+qd7fcWPQ9rPZ4xIJbGAaE+ER8bHNsAO98JVyfSPpHHqEJf+xcOrjRcLiU
QRshcW1A3XoqIvuCdxuoLcQIzC0Q0PQYSrRSx5zAhZi9YIzvPb6EKpw6EtAmG5txl4vFkqw/yTht
B9g7dgtXotTxJs6IMP5rBkpcNiXMqu3wIuX6g0SJW4Ez6u0XtF/EUIZvoWYIrIStCpn85DPLGn27
pITP/tfiXuhfxsQUG6iTkq9rhPyEjGGSeSPaEWMMlC1ofcNKRHjihFJDDY2AKjnaKf5rZv8p1i9g
SvzYflZOGF7uAWg4UbZnp5A/nxk1rJ0QvXscZ2pv/ilKupIpzS6w93wATsyHVvsvllbpq1LkGP1A
v34U6TWJcysXDq7qMbEDw3jze0jLNTsd13eTMCki52MWpjE5kamUS55cjRBTCK/8+NTk+4TBI2yA
Dfl9oyHnyxUJRvzWaaAmA2udf0zncGBIp9/kirgiMQsqp1ZWCxGLwrrLnSS7/1yKYkCw6e0zHdga
auuLGng4s9+X1WC5y47LwdzizaiUIzQTwHtc8meENK9nCr/2Q52ya8coCY7fRl56rxb/8SuhID4Q
oCVQztAsO+3KRVhmtjhJWG/8T9pwVmnpuFBGjJav7YFk7o5mRM48qyHBgTsWsQpIZnrNEWkc4OJJ
EZfysjoSeBgboVT5w4v9gFfwxzuoHA8W47NIkWqJ2ss4W3GTlGh9dFxVYWrogkg9E3A+yvEEto5F
ey95yYKOVRqD9xhTta/x8J5hgWBWQo6CTM/YzG9CJfbhA4HlyOF6TItJGEr3bi3lT3rU53p3x8ge
IHfucWBhurANtU+fuFGGrxs42p7Bsf0MrMNLbeQLTmMHjyE3sYZpOwK9x1vYc0hpy1zhE54zGl5k
6iCsRwm86X3ET0IaaS0VL1fr4qusoSUiU6fVUVkfborjdvOrMZF4QnZGoatb6DobuVw3rn/wb+SK
DX/JnjfmASRPy5l/idQkmEbHZvSmcyfIHT1OFbSf4z+C2nrvp2NhcZeVcE/jRx/2cHLQtLnwSZLt
+1SOSyNWmUG2EgYEFyY4F5NPrPt5JlQivVKmuuYT7B+kxWBGwZgTwFvtwm2gkAYg7orioWk/DIN2
pc8JwJYNQnkbJI0/Tha5uoG0BGXLxgwblJ8fx/MhSK7J00PPvvUN9PnYEBOdWTMnlpwgOQSPfarH
SzK0AfXS1RDKT+QZFqBEmp0kGvLucHpEBG1pWv8EK4eKIIoHUbKBZkwSMWdfvQiWl2CGmtDGs+mg
waC+s+59WHQYV3CZKPj1oxBThHcHERgkSEr7kuR9OQaFUPRiXjn1EZ+AInB3Dsx2LI3/VntnyM4d
BWE7V2qbtGSTBM9AT764H9BDcZ3EUc8mDXBTUG7f/XZSXGD4gRRixqqy7ygSEL0dzS9IuecrXpLx
Bry8eDTcnhJZHagU6S4GciPICXAxAOioyB2xEQ5k+Fm8+KvyOo6jmIuWgbN5N6GHLnb1qyNrp8Ch
4O31npLBj3K0SeKYfvCSRpUcqh0IeJrV5LNNxUrqoklo5xXwCVd310XyJqxVjAd0N1WACLSb6nIq
t9wkDUWZ9REBWlIJelBi6f6JAdFpE8SGnwsMT0h9e17LdHqYddou0SXt6I6xdQQ/JYZnr0YLXCzF
rSH3DHEQ8vWTqZFrX7Rclt3CHpbWFJriFouvmJGsmhRDSwmhDfOkQakGiqn9uAS0OIPnY0CK5jFi
uB4K6CH9s/pEcnBXcyTDIL9vvthPuOH4PcXhLyOnIfg35h1PFfoQYFwz02wULkifKC2m2+2w1Vk/
SpK+jhU6KZhlzr/v8AT74UvGNLngaVmMBwrorOSsu3TWrbMxta57igC8PGNLyNkzxwpOpli7RxPz
46iZOyvt0UyojcqpOy1Z6eW8rmF2tpi9lXVN9cm5L/xhVJloxjQ0Ok1IQP6iy7+QW3Ppyjlvp+Cg
T1ro19OVVJMoGQFOzJXa6rZAhPO06Am8O6bt0/ZEP4r4SypuHe4agBDJ37o6T6vyY2YN5JYEKyqs
Xwy5WVKx1488Hdc4CC/DREiClusSNCDozl6npuZcfBL7EV0vLFpeS8BNICwmXQoQxcfJn2FUfRv3
5qVrJWfhWOvPDRu6ptu/X87JjdsTVIxV1qBxc+qOyQTUCP8eufxvyNAd5C/CtLm/Qs8V3YCuOR9o
FE29cFITEVHuPTE+4VLrDMXSwJCgBqgOtaBVtSQ9RqXkrB8/ScrmqOaonn0o+GYNo6/WDTPzXck6
kvPnDTDBeJ6ZXBmZYTm171zeWMP7oGZQwx47FuEQAhAlR43X0GDrAwabcartq7taw6y6EfALfUZY
BNPCL2UNkx+RNga6skVnaZd3M7ZZznzqU9igO+2xuk+afmRGxc2OWCw33JwBy6htZaITaoPVTVUo
Vvbbjuot59ZCshM8bc18LGTQ4M1l9hwlUrRiBuYxK9IGBQONbEAkCfbt+p+tv3nNxum4R13Urn0p
U01OMnKkVQrIHphZPWS2sT/6pIky/BD/XpE9V9NTesqbKMMlnfUTnoLxnhejexTL3ztIMH/Zvc6z
vymncWmP56TwC0Rt5KU93xkCUnsEn6xi7S3DF+TV/UKQQfWiZbaOIs5VpEv4Al962IUxFt/uBfxZ
QuWTG2t8dr1hk5jXGpva5OSvC6uLCptQYorRSV9yaAWiBpmTkQoORwgapthOtaXC6gnbvtkaWTDf
MmlZGWBp26EkyILvpJsR4XMerj14aWTYJeMETYT8oByQlsdzd9eiLXIgLFuKFEmDIpUHpJgx+a3f
kdFCDAQsIa15q0vITABDQAVZkMXQa03pvJybbr5ydDtFSH1jaMCdmQi3UB273w7Y9wy0o3wASMhU
kZmbAqzg2KY1fkIkJeu/AJcKFd6S9ykH9FKzIYIhXwXkV6z+7ZDlUUMFMDTvkK46sA3fe7QcBSWm
nylPjA8HIivwJPH5Wd/mJ+Nm7cfL8MH5kH3eJjK0dihLlod58f6EmnVYcKqhvP21Ax9CtGcOr15n
9/Ch2ObTe/9WANWn8+t8JQ/CniPYhyPPSbfBSnWkhKbLhUSpL0DnvyLHhifTkJHD3UAf3zReqslZ
cq/XGTiUQvDuzbqfFAbKquJjR/CcXyK8nItaemfnoxx27TEJQEvvkDQ/3ehuLDcHkcmB7Rc4+qi/
n3b1XkpUWXl6AzSoJAEe8mpzs2lN9gHI1Eh1y9IS2I0qE3GwQgwfknC1khrdhZYJbht3eqMDNZ4M
t729+aIidG+LTFT4SnQkYl15mycZBCkSRKQM0Jd0a01TAJHVFdOXYPAnLK3Ji/Z3+AhGu5gNzaST
4/AXxUetda4qbuM7GoCJu1iUWs2lLsF529QJZOXxTNDo9wn+4KQ6nXE5rQV6x98whTmYKXRMV35R
qgAbGIbn7e2ambK/WK+PrD6Eeu4JmVejigy04eoinqAuMGfb1BrjzS1VS+oc/YfVjik2TF75+lWU
6ZiSb6RsgzRMvLvVP2SqSPJupTRRML3D8sJ3Fq4xl9VWYF1GQLt0G3t0LMGS5K0CC/JRjrAvq2f4
RHDV8ZGARVc+fRjuQnkZ1sj1XFtPWwuvSJ2zPnHI134kCSS1F4GsUyw+s7R/VX2FcNg0poHuYXgr
VfYPrJtMwWyIMsIsvs2qigQ43mRAE6PRmHjFS7ePm5GAmGu62d8/RW+v8BIvJkXTMYKyLJVtIiNP
/0RvP7M6OzgOORUWBYX4g2R95RtQbIUDXulZfkfBWsUVtzwsiXI8W4LtlsLe6isV8obTOHRxf9q9
9LwpGTFEw/tuhD7dGCNPvDSwYyLtI/xclcMRiLZ+j7h/xoH7UFxFoZ19iFNhcvej8YiNQtU6vFw3
NN1sZOs19Wue4npvd2x46yT18nHQtZjoPp5EhyQSulqPBK+P/A0QndxPFk5AobZwQEGRIImHNbgK
ydH3g3+YpjdpsIDFm96Al8MUdiQAwg96I0/VjJNCXf21ANY7PzMvPcg1yydHBRppz6VwXR7C3UCx
V2ebdYUezjl28QHwc8qFVwIm89gB9rkP1o7XKWhuMUYM0pWWJaABqU4IX30KA9gcP+UtdTSVNzLD
RksebucBDXPIRlNMgohLZnhRdZaCAh8fBSL0hWUonyMU3gvddZB+3M9k1p0yeKRI9rBddgikMuOT
VeXOOTjQVbvdSVGHE6uEMsUKsOvWGvWx5LRiM/j/oKOHGxjJGOmwPzJNZAxuDpa0YSUwWdVVBWl1
qVcVwkAPmor9+0bk2/vRCKE6qwWzPthyi1JHOJ9ZoMxtfKVF5gkuncj19psUj0TPfw0dMoVfYV0n
Hfzzpcz/f+Qq/5RWs8KM/CMPBt4kuzMcbPtn+8jNrk0/Sx5f2pLCwZID2LGg9DhCeGygoo2TxZ5h
6dFl0MahJzXv7UawG5eIZ1HVSkq4+7tY5q9M1hd0fApMG9ie+g7X8lGP+CoDkxUN2b7VOa99JnOA
9sk2vxUSTTxWaRS2clNQOeowsveQek9fXB0P1cWE2G8sgGTWwyKE9zmxae+92MEXh0Zj4JL7XpXG
APZLMU6QIzxW+TsmmNIqd8/A1Z8jy6yaaq9HOqU9/mjIMKP70lYH5FhY8l/bjCajMC85Fzx2AHwh
+Vgz7FlM/8fMhrSynBAwnv+JZ/xVmTYU9kcRxlEa6R85BoN8ccaCwEXnBiLCmWYdxkULPqVGk5QJ
R23Ll/2+Sbj/I4DmBFQLuH2zeqEZAXQHw7sEfB3zEX7If4vNpb/Io4sDeGP7XU7FawNrxrUCV0l+
+T3OMdiKiAhWUI88aHrq4qu8EDeOoepX8IToIbGClnw7kkna+JOsg7rof2a3f3m5B8JKWIF9ZrZZ
Ge7iK75MTn+yPNRf/pw3nBij4USLMbuIlMJ+2OHsOQeDyJoA/BYjo7hbZ/h4Z3H86vfKUZ7xJQFI
yaHsCG/Dz4BvxPS7zlJ1aNN/TyGBmVQikIZcqDihiaTB2KfYt542q5XoCRQOf6oW6DRCn6lSH6hz
4xA4VTJCc5ti2ucEfUJESL/y2uZopFV94T4wLqJoMpsDXHG9T470OQhiIM5jueFgXwcELsWr6LCa
oTnMOL7paoRgXEzmid1eegfN85OYK6waDiXogrL1LmR2gbdNNh0Us72k4bSNzqPUPPmMbV4sZuCy
QYEf/a+ukzbYJuCyLdGBfNcjbOWtw/kCk4odhHNluHXuZz/Z6C2nQ0JvxsCgthCqThjMGUfYuW7u
q0oCSrN+1n5WXWqZldTViIatOJq2Gq+8svAyzUb88NbhoQSjp7lkzrbiRusx0owtbvyc3ePW2blc
F2ktdRiW9vNsPp57RgWdLSAVVEELa6h0weiko7TYPTwFpA081uCQP9sKOnmlPO7eMmjsfDTk+uDF
EA6Aj4RStTjsLIeilUQfBCbhB1frukXiPeIxAPX3AHuQgYPNEbTDml9fwCln6xa88+bo+ZPl1BgQ
Yz8GOARU/UBBmQCVo7z9Zy26UFXZ+u9xrycV6V2YlUCHUHiu9mxGYYrEWYsQC/k5YqTwDuNVFZEp
4/RlVY+pJI+KkoLuKcPUzSbRueqH5koJb21XNj8v+P6gxI7iQ/bgyGVcFImdI6ZM53K9Gw4el6wa
zZRZU279cUxq69frXmcuGtfyXQzZ3q7xCYcbqPg6kLeuXmhiRhsGG/1a99Ti2vMxWM0PfwTdC91j
kuERQjO/x0xwEhqC7r6WSHW9ZdAmegex24M9S6OrEe9bJQwntx2hUIlL5WqscOE9weJT7WksbwZA
Le7JG4cVg7L8DgflMPgQAPZMJv085/dQPqoUlwynPXTXkgtKCOHs/tW958EkXBjTZAOdlHN4eMl3
UWx/CfvlIU7/SilKKkVtSRYSm/ceISChvD0upD+GvX1NlteWqLlTOMmRi45WIsw/t980JN84NCWg
dCZr/DC97IbVYj8r1cq+n22QZGoG8koFj9M9yKkoi6Vi39xqakama9v0240OayRRkl8tSJNqEBhr
LIdVTqJLT+FAucpGB0M3+FsKFOdRKVk7c9fO0QCm2xw2lsUE7KF40dD6d8hZLtgJtghdDNtLYeuE
bAAap9jwPDXgFcGhTvZlLUVfHS7pgTDzHtYE9ITuCJmeDYno6CjLqtnVfyHdHL1hKFH89jtfl2cP
AzNyUD/iqhIObLcYMFWIacxwjkryK05IMePY3cBd0Kp3neM49CQfFFEiP1fz3FxPZd6EXzVg2bpK
7eyNLEsN9aH9j6yBb0qZtYej59WwXTCNqB6gYeXCoJb8iyTJ5fGF+ceUC8xv5vwlNyXIFh6CPyFu
KeoUQ9O2608tEFbss1Q9sHTebrf2G1TH+Uq28+RWYHF1ZCw/z0d8BZivt0txGepU54U+vqtW+CxJ
rgoED0ernyCXDMJbFB5Td/rz9IuxkhHBjnMMRRNEnmAzVisbcPfkx/9Vb8jZczI8fgbaghTC+/PA
3mZ6Ueu1wJUTOmJgBEw0BpND6zQg9hRtngWRFUiSA+OvxwiQs3qpeuyzeWi4I3btr5piW+yYYJdE
IWTBF1BKNs2i8zbRD1/JG5MA+E4navS63ble7s/+lF8nKs6fNbKeryXxagPZVBm+Qqn5dvDjwxhm
u+RSD2cLHo2snB/ELuBSV3AQ+ndDxJa2j7D1tHz48omXt2RlrAGL/iwJ13kjofFu3j1L0900H2cR
NatncNhloBEb6tj/yqKeefmjtbnIGDppqpI1GXm43bVLvDfpHNrsRqpB82eZBCQbP3WKLMeFqp68
22rPNzecJKr58vEtghWntdgOIb1hPHMGTlEswgpcDDwmCJ38+06yZ/UcYO016wZ8KUr+Pd6jCjko
2vdUkaOS1asK6XYaopgmCqKM5Zkqt7+ZfqUZ3qC/BctRgt6md9ZFRMWqmLfg/JzcMOy5heWTej5U
mzyTQn5GLC97j3st6Z0zBm1tiUdTVC4hCUFPA7DWOBVHwOy4mqBCtnhJsU7AvIwC3k3XQyFYSzTi
nyycmlkAPjxouYWzlWkWusbMLjYyXeOnReUQv5DFJUWArBiPqsMXreJPmjckEZuHtHYXZ9QwwUh1
06zU29YvLT+xEvoOZblQXs8YzycasK7CA02ZVxo1RVYoUtNPPPRqxURdzpu8r1GcF9CS85ycUzYF
UbIaUoQYBb7SwfgHKdrcTBe4muO5ZGF09iv9uXUdY9+QVkL189RbIDQL4G1ovaAqEXjLmMfldpuI
xub0+XjSmW4vqJl55Mpz7D06aBt8pA2eWzwTuTHTYx2J9g/8mVU3+KZb1wx6qHLtVu1eO2WjOKi5
jD/gCh7lwFxJzHH5wMHOT4btNBK4BtqQF2DYuNdrTYioOlGDZ0l9aM5tdRbtFcQ05QonBd+vPgn5
e6ovm1CX3ATyuleF5YAC7vwAG39ZJnx2imQ8sqLkOewuE/NnQFMTEmPAavcNvnJkzlnASMse1+id
Pm6v+2Z8hYRUPdIxWpbWUU4Vy/AYZ6OAFl9V9QjPhe+Y1xAovY1dwvtd50dlTC7uPZD79MIh2byb
NRvKHBIlcHWQVUEYTgHpk8Q1kxk3DFKpXAdOhowp+uGIQeDLJuZxl/kof7gFDCnmeiQEHX5tFu1j
Krr98KotP7mZUbbjgkecq0YRIzJHjoDlMAKi7HdNwbuB0f3EwMC82lcKGNtSMq2uqcQygbVZt1Eo
8/mXor2ixHbHpHdV/RffNXGJuBWOm8j79PhL8nLDlFb5C4B8y16MDM3YnWs1C9OJ9RjfZepiJ7vh
Q1vW7fRwu91miWheGqrKuJrBYxfxkoWQKNaibBNysXVl+gUfYBOvvLj0K/GD0AR5KyTJBfXxoSpe
aYE5dJfIJEexB4qkt7O/sbymm3bgI90Mry5c2amD/WyhRPelu//f8/jzhgP62n35UrsiXW5d+3uR
X43+F/v9MpUfTM7+5XApjnAuLq5vY8AJzqsWujWRdoy2X6uHpP33uiKrsO6ja+Q0VT+GGe+ukKNA
UsRYJel2ciotKCCC8KzvUGLOBlTTLc0mZ0U8G8qrEn8mVmLIhG+/i6PAVWNDxM35iBOn/h2ct+WU
cnOd7/eI82A8IVlEKyXuAZLXA6JJ8E40qTorrJ/aSZL+U9DuBsxXfOXbfGnbh7kxKvJFLpGGq4OC
gavY2xEoZ3hWIcZdvJTpQaZuZJJWdtdnp2m3vzH1EvR6zHR7Eg6y2KJc2TvQ2T/jxDhOYkbfHlMv
0/qhP8T9i6d9Rhe/O/By7XiOrKeGH5okIoMHaUrz4U0NHR91g8cz41qRqvttYzFfM8K2+gG0pdo/
yx9FHB4FeCcWeKb4P2b7mDE96MqQxFOv5EKqa94cyLN8dai9KkQRROpFZIXSWaR2Q+sM9YlfzOJ/
ayER9yFYApFL+DiO3G2O2Vkb69fkl4k/IPEgtS7u7u8tkJEfRoNJojk+4Jh2Ob9zftCPH/9zfT9Y
YxXc+KGlBisjvvhmdKYXwxxsGqMBVCXQFfZebzCvSJLLrlfDt66RB8WxydWM/0+L15d4lWmpBQjs
0ASx/UYG7oM+PDt7nQvL8Wf9HUANbOk4KfRmtBEFCH+sIZowccl/fMU3XbmhrxsOnFpOt9Mw8njV
Qb7oDuLyVCjYU+SlGrmui5mYJZSWQBABgrDKiPnZDtUzayj2j9FmHs15pwH9mfOedKih82D0caQh
bQLuEQ10Qd+nPiUZf7YBrsFpfZnosvgsLTv/bTUgIp4wIitGdtCrq7ukVK/IxZZNiVJR16yyYr3N
f50ANlU3XTUrKPfMgjEFwnhS11w1YsYBB/V/hFIMOWvMOVg4DZr7CDcK64gKCyeSnlCGNFEhoPM8
IZS7P/tZRncb+Q/z+GCnWuv6CdI9uKIkVE02B+PmQvmD49YAdYzC3aCuG1+fBZNU79LLsWB+fpAY
pq4eQay+cavGI33nq07r1LmBN4iwM1UaMp3IuH+JX35APi3EUj0e9E0Is3hnhPd2hKGZCxp5GsLE
fyPorag5GSg+k6hVJkfPa1SWzBPWKxpDIRpPUAwmtjSsAdH6ZpgA1kByq/sA7jCcejGcELUGtr9z
Z8OS93cGn35ra4uM4UO46zzJJuy36Zx0IZqGcQJv4MItlLFfeWJD4K8eIbYJL2ADrC6mh52ziuVG
BIXoNN355xe3AUEpMZrXxQIy439Jwy5Dd3z3GCK9LBaIeXIj6LRtJGagaETJPpkYKeHn0MpWrBsF
7dOoFTtgtSJ4nGfY2XULGAyJcmOUqjndNW0+Y+KJqt8FLrc1pXyXNaBZRa29SfvJgOoI2PVyFQ2R
Y5Ms5DHFbJNk3cAoIt+50s7tKEOZKNOqswaQr6YtImH0ip/bm13Dtm5/GsnqXBCsPlPsR2/vnery
DiVGUACi6QOehkZd8GEbHJ3g6Huq0HnQHSfBj/pHVplS5xkGf2cub6ef+aWOm3kZ/Uu8pVXXjgD4
C0Mb0YNiu8Tmi9beSCU51e/RTsqulwlhoONX3fGGppSdydsCtUgNwkVsTctEzYuLs8BMC7LgHtjl
L/m/eI4JWHhyosN5Y3qS3VWbOuHqqjG1HA7GA6fAHSFM8oRjHG0ywjmLKUXZqlFD9ldbD3z265rx
NSUDfkOj/6TFbYABFkFF++RXSyLukjt8pXdvZdjUEXre01h6be3HlCmyBfQNgvXSzfxMDR8B+kF1
PKeYoyoSFae12EdSnKViHPoyI5D2i5YhO4jP6iBaCPznjqWQqP0j9W4OEjnO55zJbWt9cn3t4nvX
JSrUwSipfiOalapfEAPa/cIztG8hWW3XAabpJ4Fc+KNkqAsESmKn5jE2pM5L47iRjV+Seiqz3aX3
sPMK2mcfYoYFyWDm/NJDOIQvUwyq/87okFUBftc741o0WwBCdh4Y6WUsxk18RPd52E6ab3QDCaa8
B27tP8Bfg+podM3WGxx5Jp3kbGvuZSlxdXW2PsryVa3sWFG2T+0g2713S50zp6GeQUF1O44Ipe36
RWwDCCUN9Qr3OazF2oMxW5Ndc963XdkVAcro9c0FUPjCKmmM3N3nUVTtZCjTPOXTvNd/gN9orNRS
4MC9IcVpc/5zXHuE6J/zM2rVCRzt2TNgFa6r6yk/6Qro3xc5HVxaKxwNJcX3QE2Ko8R3VaIwFWmF
YR3awY1gnASvxbydzBpHpQbRbJjGyOnwPliCVK4qe8xWTtWTbFyZwDnS9Iu3l/VXDA7nyQyXLAAl
JGArb5jd+QctOG2lS8guhRHLPDdv+V2VvHY8QvBRwwxBQjP5BXwBEW0BdtmXBVuT82Fj3lLRjuT4
cMVRzWNemNNIctYWC8uHqAzKLFjJT1YtLC6WRKu69Ul0gzyvVjdWXQyRjWqJb9Bbz5HvPnVkfjAY
WLgQIy+ro2evwwM0DLbvPZO+GhF6E4AuYZDY6Z7yvwxV+ZTRKBDKv5URYaCqGvrdyx2Oh3ZhZzf1
fSuT9rRNjTnm3ieR5ECyD+BUUsEZq/Z1ZjpUJPh8MmicFnWMIYryrraFbyZzQroTVCbTAj9JgPn9
5eU3TJpEO4EXW3JuGsLViatiXA6Q4aFBIy97W/VgI7jDR2Fxaq33fdkBRiCLKXAm3uvgxsYBiKai
1JopnN37Zuu/E3zVprKQfx9F7uSdwVxHw2BFUy/uHneY0vvjtsYUGPUQKMVjFEEMry1rOUk84r+e
G+sdBkVaSU1wBL9mwHhaS89MfW6QaH392s9B/CapwB32ev6Hreq10tk8ZQ5sOqzuyEro1YE38EU9
APVc55p96joHy6mObByw6GLLRZe9kVQwMjzyK/qI4rM4xpBwBCDPRo3P4lk1LBA2rL+ZAXp3Phaf
NcU4PZ4tO6zgky7fxvzoO8eFD6MRwAr6/Y6Sa1xAiO0oKPxLwnjI+6xn3qXUGFTfTOsnnLf22rp5
POZFsuT4oOG2hN6327YM8kNGiSUClcMzm1m9vdBvzEj9XFye0xAEHJ9K2t2MA7WVXupQTq9NjuJs
6jS6XbC1q8rkye8/ze4Y2xGJ0/1+o/xb9lN/q5dX7tDYXNi5LaCbbKnGkMGWlv/YN+XzFXLpuBdN
eSpZjP4Ibd2Amn5gAtH3cHq6ca1gYSJ1WDG0PFEO6+E00qVM3zmAH45uvwqkJfHo0DeAG4TZw66Q
6tRXldOAhv57kS2nmwqRKuR5g83Xmz9wYOhKR8ZpLzQfuK8ZyWdc3OFCoNfUO9sowvkgSuEfo8bE
I/4mNbygBR3U8ZltA4UppU1KYS0xiu6UBUUqP4XNRgPlp/m+VcvdDbFJSdDOqxE5WNceb85gTRLy
MBhnT+KVVdcI+nUzCuBsUDCp2tjbwWUNuuw9SWYA1pyXajf+FUD/HXxT+Mk6+BL5U5VnwicpFkOy
z50HR+uBOC89TQG5gSs671xOUEF0iSScA6tD4Ur9pBmSmq10K+Bu2yjaADues3gRiH56XdP97sw9
EgenrcmFyGHqa5683fjKElDl6uWn7CdJ35QlvHSNJgDmZs0jcKSG8eKZqxlmP9R/Iz/HEQ7aHR7c
cuL7qEaydB8sgoannP75di5DS+5cUnQ51IMKaDdQNzAJxqAGdd8IX/54rlx7m9ZZ2gvrgzNqOGVA
/veAAZUOOE0+BaOHjlPZ6mcRe5e+/uKyit9vIbZJYmsgf5z++Sc3O28DpZBmY8cfP2hWjAPZSSoO
VThiyqfo5KWcYZSznFWoRqVEId2qedsmvxK31IOcDjOpfJTpq9i3adaFHD/y8aa4avTxsLeft0sP
tXMndKhjVzuX5TJcdm0+AqPXGiFq3wxSyejrqFupnhfQScgWAIT97xBcZXm3ixL3mSTW58UjGcRy
U723gSzSfNTUnMISKxVJHOGuBlrSt3zvu1K4rXIyanfK+1TXLQbaXurhzTtw+K+wpERUQyXk641d
F7fjiDnPkrrO6v8q0RM9jVGBr9V/ni4mY34/t3bIQ5ViaLP9QRt03rOCChKl2KE6oZOt+v5Fs7nT
5F0wT/eddMhfCdBhdM9H/TfdnEorNSdR4/MlXBJerKwURBE0HHt+2GxJAJ7315VgR271aqJJpDHP
xFkeYrHqFb/olzKVYBtA6FxSlG9uPMxgnLSDqXTI1zsJaJAlWwi14Q3TF+9poEQUJsO4n9iXMoyl
M4ZzfumCHP3cPk8RZJBZg2bcbbVoLO9S7DXTsSwC902kN6GzRgustwL12DrkVHkCpRkhCFhyffqf
S60eM5Sr1l5QbL38syOUV5G7ciUV7MXK1T1wWLXhyaELjTp/gx6fJJhtBnsoqHJFI9c8wBGsv8tn
7vuwvfi1Rgawes2Rev79rxWmS7EgzOwbBgJUneMzaLQ8G+BEMt4gr8qxeHJSau0iUQmALQQTalSQ
96x+oiu3rhG3oD3TEQHQtIU1LqUVNbT9usadAettK7zZRogDDmLtfJiCxKdHgbbUKMdn3ICqYS9/
n+ukIGoyudgqyRoGMnqxyIu/iBccOvefR5g8sbRWqG75N9G6qZbl1mngDtuwa3Xtls/aLIelYXN8
7/uBrzzpIhp4VobSNDhHhdf3fgZVV58FYTE7JNfUnP+zMZcuT4jHA4Tk2B7g00Re30FurJUopcn6
El7RmkGIDiK2PlWP9SUs/qhA20sJ9ATZaEN4gYIktr1HmJQCAHpMjOEG5MlgX3M6rp5BbxqzfK8x
klPXf6Ixxqhr/m1kf1ZDK9BDV1df4xYQs3UqY58fPZ61GmIUAswBaCtxFdy6/uoI0VbX5li4TR1f
YHGf0aDAHi1v05p8UGRDpDJNyKiW9CvgCxZmNLbz/PtREZIZBvunc4ONJi8u7OQU1KOyul8Mu2sk
AxRw+8dWH5adkM7zfL09jN1bgXNa03g7b0nOL/ZpEhHcgUgauYxoeSFwzx0DpDAqlbgFQgQ8DGnr
J2+qYe7rsoFexIll91Jrjpmxm3ZjDW0LBc+E3VGrV6eO9+UuazkwNIyTUkJafTctSY5ZfT9l7AIH
bUSc/76jVrbN5K0hb88u9uvj2W1ba7asO5DwrYci3wtaGuBJEaImaCYyxKBxYBo801wTr/9JJdNw
IwoW0HQbqt2gTI7naOFyOlIGGXg+kZBNrHlEo757SAPH9qqex7He90jrRmhbiQXaNqtDTJNrVes/
C0bt/VQsIYtfmDB0MJcz8OlaUjOjnCXm/Bez0qkILMUGlT6qUp2wbITDYuDeHKK+lJcqf/+jWz2B
qA9BousGJDS2M0XQNiaf28CTiBKJa52bu+uZQdjtDhM0T/7ODpkOp5wcD7fbUVAg0JSVBmkGhaWx
gYhcdaFNuzHg1+uqRdgm/h06usTvMAkjoOZDLctfaSP7gxUa27QeVWM9+z+YprzsirYjhJa3wksB
O6TeuS09RAeDIs7A/M2nstL1i+Q3mON8Umu81hMBbaUXH9gmnsukGzs6qo/NTeek3OlqU2dxch+Z
cL27oFcjmqJBkHchiGHMatL/LMAI9EJquEkAZ9fm/Kp39fdsr0RcxG9abR3QlyVixRnYpCziacoB
CCd2hjytAV0gcET6jH6HL/5l1jVxnZSHRLPrP40my8Qqqs4fAFd+o4V0A8mbIvnbmx48N4cQBtPv
k7IYwxaoAFqDYsiKURMABeT0FgiDIiWZqJYpOwADxJtue0+DfVd8jajm8R89m8ROISEh9WNIPJX+
zDWf4j3adPkqxdP/z7iK3MPxX0tWM1jh8DlwMdwVFKXLbTVqbFQkFJz+CCjdNgZNAv57BSNuToEk
goAQ8/PEjPQJkiQXRjs8hhBpKitB5O/iZrZsTuQL8WaJB6VL7pEOpmvtkJ5B+UWjoRC9oypNa2+h
k5QVkSBh2lnLnIdoSRIP5ahYkN/a9DpeShdCdBoL3OjZSlJtrGzjjSPMmab755kfGM/wwRZUJc6N
axOHzfYymA6OLuJzBpOvaP6tS2P0xgmU3c+TQ+ANqStexRzFIW77Nxx7zGLgOjGePBNVuswKc1q2
Kism8r8ZhV78JRKxNyNd7Bl1LN8X8qjkNIbwTh1+eOWiEN3odMB/hS8Zm0JePbfd8fbQagZQyPjX
kkB+MYrYYio5eUYTDwZHxPXbk5ynB9L8Frd+RSbKrvNA6X2efn8TgQGvl1Orkb//pcWYU5qE6iex
zfUzvblTRJ0IN9GBvFqwiVMl0+3fTdpDOo9L4kI+6mKtQilH0oQ7O1S+d6/jG0GknG+i9WK5L54c
jlB41lwv1DViQRzknxf/8d/2iWlF9Q8ZZSpFg2s5/CY9ogRRbLL0AEloS2OIkcWDtL/ql1Ak7576
8Hn8epp8oZqkvpAJkEmg7RzT6lU5ek9DkwVOtEdyRpI3Vh0qc8INvv6pBw042EJ2stXlud05Yy6B
QeYNfdaHaMn7dVD7cn7r1RG/kxKzaiodS1Q5KAv/I6I7j+Eb8aJR+k2zOQoa8weRZTyliBgJ3240
W+Q24+aNk53ZMwI5aj/HEzFVxXJwutlRe/xTE4A3uw/YwYn2mv1orr35NSqH5kW4iUUmIiB9A8NO
Q/8p0vqV0siapgbMC6kLnvPr+xiI6h9NBEmmgAOtNgUJwz4XDEbr5LxrVc9+p7TT1FofBo2g0kjl
mNnz9+b6Y6jO++TIW+flqAuhvQ6GqEmXR2dyppUFoBGq/jJVp2ljp2E0lCd/BUYSrdomSstXlpLB
1s7345cllfBdzvLNOl/yWxZG8GFbtBVID8EMU2DOz/07Q08iZTJQJNNlKIyc8yS5nfLW6tpbA7ZE
kj0C7xhE7facCTIH+GwLn99df9FAnt7dB0MxfPQHOn7BxQIKw6or0AkClYTjVvuO18t/XGoUhTtm
iv5KDEPSHA4lpy3oabAc/qvHuQatmN1kYBHngFs6Lk920YWaGtPIXRnDDjW6QnSJlwEh2eKtCHPH
KfWPXYBgwq5knXoZvwmJ2dAiQeZ5ufzRqXcTX2WxAyWz2txL463ilak6OnFBmxPjU+ZiNmNZS+ig
Hy2s8Qf8ytyw8CY5RqauoOg1McwLdw6WemtJUHqm+aDKn0y7G8EHSAzkpS6W15Ka6xTnTcw/ZuRx
AuG85b4cX7V/bxTO9ZeIbV/kiXuGkijw/9cXcWJICk8qfg64R8gWZLJqYA7oqV3DpTRY0JcO/PII
a88bnMfRZcDw34HKK4bokj4DOaPTiYv0umwOCIOL9JnLhHm+T9iEz8o47tX5VtIPscsG9GhFnfRn
BVrSImXw+MW6SdTz8hDeiAqCaPbgo/YKO5JLV/J5kcZodirRTPR2sFDa/TsDU21Q9ozZ2w3sw5iK
F0ztYz+ISJ/G8V0XPdvDBUMPe/D8YW6nI5saZsRXB+P5A1u7FJ3xdpyDuw2Zofc2OMoUCfDWOrlv
+KyPXt4pkUDu5dX5V96JJ1MTeffC+rU4wh2ZK/AIwQGHq01wcFlNT2SbJnnnEr0XO+rcSXxiJyGc
tWg+S2WbMdvg2aQw6TksdsRCGxhVHXId5PjRxdspOTGMlYgtVF7RvniXXpa5xr5Q51D7VyLUBfAb
BX6dP42Gvgvubk/ziC7fImjzae0A4n/a32xIv/ZpZmNb7DiVCHMlChLsTHyUmQX/YWidYTrRPRuE
uEVzaRGVRkzV7iM2kpnwkzLaVJiHikUBEaOEJtPRu3XWNgINKPSAk0kpb7NEHNfUttPKUVJbEaf1
e+81wrrkPBx/XyNBnX+EChLcl+AViJXUi1KgwhJ+e0mE5YqV80WVOzNbwvOGUefNQmo5cCyasTF8
6nximTBqL8GmAL3TO1YFEliECsU6qVNXmA7eyL/gkikzQ1R7dvUyYph/8nIAu4hkF6Js3/xVMoWf
cbnIQmqorLtgaF6QE+QjROSytQnRHcO2Lh8+kOtUaZTx+OAVGyRQUsk2gYNbyJKDvKc0EHBfmyqq
EgLtQOWeEfMaMT2GoABprVuD8z/940EeL/h2LrwJoNXzWk0XhB8kfCECtA0IXGHG5sTx6OGWpkbj
dlcyaoWS5k0Qca6c7XDtGtkrICmfRNkewNOwnpLfMPzsn8YLkCu83DMM+04Rd51glannGoBNiZNV
qfVNgJ0vRxyO7afb0DaSNcUsqjuC2fg08bE9UyYX0ucs/t/wHVlSrYoTUheyz+miX+pakZpXCl/A
C8DvCErSD4CR36x2VZ2fRQGaHPi1ivUTIQUyRgdByr1triLUkRYk4bw9t/SwJqhwyqMNXKtA3jsE
D/Vh4vlAeu6MXSeSJGU7vAwz+EwKPF9KSi8PuKQlOgueAlaezMInpBv5fGp+q3PNuOqH/Lt78J0I
z4srEvUOCmEcK4MSaj/jJ2+LgIhUjyEkCBYRYO5c8+iSljQPiTkccBh9Oi/yJr0kPJlKiOl7IwwW
Klh9n7Q0ODIzefMRjN+QBFLQB8JyIScwwJ7WhspFnvQWgL8ipFrVOHJkRraEUf+lftd4zmDoX/lm
4DgO56IKJk0vUYIBYxqAb4kXwYXa3WTn4PBrFvYcEssuIiW714XWvyUd+s85ZdRqR929IaDuXD9T
s6yOIxpoArUOJgy0RwcNOUEGFHjsjlTcbpu12YPbh45Is3+QVW/xcr5DiM5AHYFDal/gBJPHs7Zl
WhwZKWABXAUXTkHS7JcIFyvRhGLoFXDqXHG+UiOgjbuGFdIKBQWHk7vu+tgoGALzkMR2I99yNp0+
S73JWqNDSl3veP+ShVrMprh9mb/IxP4ndMJtfOjUbMogBRwg0Ts29sCcPjVw34caz9KLn0wjz01j
sXdv75c+qW5nmM9Zc3b9lUJMxjmLKtQYAnbOXAROBFxCRWiXmd0eA2mBCxla8I+ZySTja4bVQe+O
ujfEk056Iug5fuaH2leolTr0Tm7+xdkXP70WWFR/0E4SXrmSHElIXaBleNN/fOSHwdugmTmtnx83
vxXex7F/tRrJY+A9z7n2k9vxi3S1PEIQn3J1U7tqoVrCCmBcz4w9XYhPdcGBEaCjR4HZzuXxgfSD
p1tjvKKQehHviF5w3hzdEUv6Sz7fulggjHkZRcCLxmiPz6z3Zm/xtBb0oqtxba19yJfSg/yRpcNz
6Rpt3cOERk5ymiC0rD2R3vCUBiLdKAaqE4fcO6ZuDSnqgZa+eg9dFk7sHDlYDza76VsAei5c/dDJ
AhXKb1y4zbJNSHr03X69BPcIrQLZeB21hKuXWte/Yn2mD9YH2Eu9VXciM44uojQCP8G7dRwHSL0Y
GAv2iX1VY8hvVm4CGnxWNYKO4C6MIpYnyrePVhZvBiY7bE9IlBlw+17k2uq5S8U0SD7qcu3QOLvp
M4eAeNdbiJDUuiFpTRHqDv47ZZxof4Zy5+8IruKMLDmzkn8R6HHSQOuUptV6G49kEX9WBPCKF3fe
bIzq+lxIbL5y4KUaVW3ynfPJ/qAODELrUj2gtPut0HiFcMAHPCgTVwCrRmShGJV8FQZnqeH9gGeS
ExqI9arwiSfwM2EIwlTbX+9qabOHpm6s2cJvHKdljq/MUJ0QY6FkUk7WYevYHS7DygUHGgqlF6AY
okCb2ctTZvI85c+zb2XJAY79zeiOQaLBxWfBCU2uLQ0WxKloqEkF6Zw9LpqpM7fYsHZtWMLa2LeT
pl9fqN7ZBAj3WiHZ2UJypbDGU+1nneCzw//gesagIlDqE22oRE4LFmf7R70tmxHnl7UN1zW7sxYQ
IR98bqA5/Q0siskfQSpQ8k6b0mmTnHUSYv7RA4hpMDGDu1hFP6TkbyTeKfhpXW+m1T0up6XtMqSB
WTEZVYzwXRobk2EKz3B0YLO7+c+LSUfLAYgVx5upF7YxESm2s/2elYXnVNfsdU2vee8jrUwpSvYr
6s2FIoti26KNaQ/W7+6A3BQBibVLiFeil+inJyNYmUk47xte61t31WIJaaN2fF8Tebedb6+bDhpY
nPy54OKzXGHkma7IUW8uTh2V5zAZdx88ZUrDKiJK0vzktTfMwJt1ZupWR4qo9QPmP5q/rjJcZehk
DjBUk9zKNKC5TyyZAKtQPjol91Oo8ZRanRw0P0j87UoEuZkz8gd0CXm3ff/GBzfnshzXNkBpXYed
VYTIQ4lnVYKUcOe2ozBKBnlLioGNbZjvIjYC6ZrSiQUPJeCF+qMWYOqU+FEFPCKhILYFy/9B21p1
CU6fb7bVZKXG7IB/LieT1eDV6b/tXafMZ2wrOIJovSvGLDhXrCMQTCLnHriTdK1wzC4sWQaNAKsF
F/nURBWRB3MlSdI+vFgn8HTekjGIVxps5if69eY55xTHsP5wpNIuaEpNgoIeWuQxcV7Xcu5lPZ21
aPMrf+JYdpoSUaltw0awhlRZR+npHLu1dpzHSfC0rCtNyVZKjxnFPrxv/tv85hNP57PJ/sZpiAW2
pwOPpG/S28PAYwwzwsN5at5bKcb3odbQpQcIXIhHtJJO+gIGkTrbkkafeLl/tlbHhFt5mP3ccVqL
xNNkrZxXb7n7BGG8xEG6kdSMlmz+BUk0/XghbkOovDBk8TYNoJLrDiMsEFm2GLu4WtaYUF9ujMoP
ofn14eYPeBm249LZgWi9TgmONe9Wwpa6/l9aw1Ad0HAH7zIFnemBMzuRHjNPbbxoHx37fLwcYQP3
fUPF7tmDAr1UaS4LKYVFSW0Xi4Rbh+234e/a75SLlyXA6pRANlym4pfn2QyCOCcbB9tFXW3vNBOw
V2aZgW0r/fZvQGehSmsSPNURloV8lcdL7sjWWfzK/y+XPdfM1IKAiEtcoLHngSgn/NF94gp3r+5v
SRj6UDyVlwogbg+pT3+aCIVhfpImWNkymDkYOnToaR5JEUjCScHZNbF8wb+Ci2KrMbiZ7DVI2R6Y
LLkpMgqdhPodobt1byitnpu2xWuI+l5/+s+YvHHdjXZrDUAIRKvlCASj1e6LtOv/S6WdTSoufgAZ
HK8m5+Khh9iVdb2E/f4OfnkMk0cd+3s3pac5bXEVxwg+RB3Mz2iblbodeAvwgoF6BVLP2YuPm+Gp
H6WIv6jgPRS8pZNBoxrHZI4LWOdqFWAz4HKK7v/pY8t6kPxM/2v/OfRpMSPB/lfo6BWwNa8+dUNB
qJLxO1L+rBT6Pqvyzedi4MNkBBjui6NToBL5icEyIcgYjzV5HZDY5oB/G2b7aZq99MGwgeKG8h3w
fjx86H2U0hSa5p0O2dnaOfW9m+URwSww51M1oFhQeSIG5tgAKn57ZGf2+QevkUduFgSr0XVIdzce
+dAFbsa8K2xm+WyyBvwnW9Rg7B9QSpXrA7bLX1L7NUBCM/YgnOs3z0LmFqRfyb+Qej+WwZq5Hftp
MbTbTpkNqYoO0trzIteA/xKa6+BhzanydCO0bIucQH42LY3R/15/fgIKZnJDTdFZx6YNwRMmOlze
QQzsujY71ynRrAJaZs27qnXOOEOcn4Pvjf3Pt1omtcsmujY6c2TcfnG0xYk4dHthTU3VrSxL2Lgd
NsuLMlqVuOKlDEm+tgxu2eN+BkZXKdBS5tIFJ2TjEreaxJgcCeMfaAgx0f0tQtsyup2bF8edQOmd
/FNVHD+vsvvZ/fVDvbOtjW0W/hmyZvr58F/9iaPR7lJ/yEhheg0yDxVbaA06cfmtdL+lQeE68CrY
6Ov+ixuzQJVi8vvsjLWAKyEoMYQ41/EwCLRBEnmE+YT7Wqx3vUDENwqBFOeZdqs3Av9fM1AYcQjf
FWcDYGxGvIaHB57cQcdnsa0oGPXyH2DzaF1r2atyuuxawbs2xp13Ref8Z7rri4LrTHGZtNnUbyUw
iskmL7bVEhcGVMaF545G4BB3OX+et2H94l/c39oAGOi4qWCFGjkmPwmxBWD8wenVB+1Kwl+ykEpL
fZU0RS1rryEaUZ5W0jvjANgMs8CTysvVtTZhOG0hD1L77cF7o0q3c8KsjeG2vNPBUleKWvmhcMDn
Uq1WZqDvdXvlt/qrvbLZfQMWPqfTmJ01Qi39pNp5H53CrkwMl85jQXs88sVXOzwsfPho6CJIeYRm
xtVqnwl4Qr+/nlgKe94n9rpvqeXpoioR/WIluEtwNOWqOfPvreH0dSwXDQA7UR9sZKsBBJRvAkY0
TdiTdtJ7KZszB05Im9WqRcfv7/R+YEE4Pp8DcUO/OmdKZfvX6AcxazPiJPIs3czdDe6Deu+Wg6PT
QCQLLbkiG9Akdqzn7sfK3e0YUDVku8ooIU2t6Xv0zywiWsMxVhjNMhhlHOuhPdW2AzqQbQIu2GZl
jOeCnOoamM7TrnwEu2P/X0MQuxfBk0jFd8SjsRR/H2G3M/9nuAdDSITASh/GrVn9aaNvaoQilDUC
yOlatDKthyo/BZ7rKHLrmBexs1xLCX/HHixuuv5fKlODzjNJGbCfJclNIm/6u4ULsItpUZWs5RzI
UEWxtNCG17ncqDQtFsa1zPjECAnfCRcixP6idylbtodBzv1fpozuHscefBMFqr1/iHmNy+8j07Cd
w+RnCEUAZQ9E4J7wKpTzSddxALrsPeA+ZSOsxCrYft1I53R0Bg7i/3ns/pgT++Eo7lPc+mlyDLI2
oDJeg3tOJuAUBCeurTuKfdVoDEBqGlVSQ2mJcIOaKGwp6EOFPQq2BizfMdzPL3GaJGJBHVj2U/D7
wX3sqCj4xBJXFo/WwpH3FRMU605gc4LWadGCfy7AsxKVI1VwcOszssFcIktrSiU1lzobp7GzqucU
vw+azwo+W/vMJwbSFCNiwOzzoRKthbEQKlHHC2W2XlWKU2zr3c+pOVF4+NlDhqxlgWr1nvv8aqVP
m7WHPNyBSftgzO+AP7Kqf1F11ghYF6m2VJE9qBub4y6ygeHTnTLbcX+irwCMzlAQrBld2oR6+IMI
h6gJBGqA+sxt3dn+JhcMLcquOxtOS9TF8LWrO2MBpaL4F6QmuMlli3b1oP8KZKWW0CzZUB8KC5V1
EGLPlb1bMidut7x4e/efy7Fo2GYQD9kkqO+Yij36TWieRkUWuGycFJDoEUUvqkyAtOTmmTtbaDZQ
Tyq0GkI7+uQfnuVAPJb41z5mENDUnP8K16np4JyXKYyfqgywPqqObg1tGUc1PklEjVoy3rXe8tJj
BbXQb0ai/VW5kJT61qU1JUytrUC79Z84EbdJv7izfRaq81MdbyMmaiAQcWWULtUDXfkp+yBsFOJK
ovEv05+HjaDoyLh9L1iWXqbjtG/1jWi5F+06osa32Y4SSonicpHxHRk7Zk2pv2Y2jNCTKBZKvg2m
QywsklEMlHlrdPDVTko38DfHlozC3mewqQDzb8D9iyOolf9zdOyvCpQo0TL0TUCrt+jCjAgexcf3
fQT9TvcdrnhwL5rdWicH1drmAKhOuw0Fb7Ctuq434u5WGjj14VjMmkcsLeJlpONXK/45bC5s7f8K
eF6NgvGzTZHjnXA03pUXzXqQWP15u7LVNvZCbyBBo4p8qGwIAhBwyDNnS+9ZzPPU7CaoMnwX6E4q
/r2QllkA49+ha0sBN84P6sTFtfktiIDCv3d+iHPnE4xsl4TCJGuqxzR13it06mhpAYoxlZRLub1k
lRhNpivha9I7eDzOewBxBEXLU17TLUkm/JO3MZ58RU+i9L1AYLKjSdXZsBb3D1UvZnbF8tLNIOhm
jFMTIi8st6Z5P0JQqiAhetHgu8+rqwFhNu23yAyiYt2xhZ8Yska7e6vrhEVgUYFcVSQ7hWgsjyWc
cEd4OU7sj+gEvq+9QPxMoq/ppogb7XSWcLw8sVA5hfhLD7vFiCbEd+9IDfGOH/c3tC5axB+HV/Ic
ByZnS6127VB1XUfoDovSd+QX1O1iTtJ2vvT7nS/bHVkzZn5qUHskOq8KS1GprirPmN+43v2jj8Cx
qRMvHPsZ5GNDRPt8Eg/ATi/NtVlRnZLRqZbkqRPeTuBQ/EIHhi14CRJlGqx1xusAopvR4iAouD5S
7fTFQmsuNX8YlJN08+zLNYeArcsJ4TKkJvPRKS8+pMhsIOKJyuWpykV51Bj/6RA+3hlW1/jsxUFL
h7nnd99XlK08sqokGgrRdNOCeExaoYMfsEkgOt+FJ+aZKWBfpVc7va94iONlYYhmgVfYzCqEm/jx
F+Q7d6wYnLsLOiK+maBvnkvLhLkdjNL8R8xfL2ONW9pzEf+RcLNKfaGF6uS0WUswDDP9xu7PXUxb
921XnxABpeRuFTv4A3YmZRqTw68rHxu8Zaa+EkZaKiO5IhZ9XSca7msZESuz53ub/uHfqErhzUPe
xG7Zs0yddioiEv1AZdAMeX8exocLD71HqbA8cBggZjhmnIDLVb55StbojFqXJrpZb1feghq5JtHL
Uu512hpe2tdMj7K+3LykDCy7OcA/iCVxcmxaL90w/NWCT1ugOodFiP7Z0b3hcjtt6pWRG6S7o6Pr
BMUsHArN7AbgOEWzyQSesKe7ypCgWow8p3rZ9adl1AI+gWBjH+K2+2nImWf9RR7GmsFTNM63d/sT
e4AAmcD2Jd5CS1IrQZsBbdiq3PY0UILDEzXrL8kwUq02XyYuCBUrA0a1xF909fYPAzQEwNCAFwhk
euYJiHE7PCbzUKpz1OtO/Rty9eW0TcI7uh0jfTJd21DtIV3wscXslJbg2z8YdmTCsCRbg9hnZViZ
0TqGlOYWqtMlGW1/ZvF/mMOg+R+Pv47F+zI6tUpkbaCQZ6mFQIXQE743kYwzNzByKn1U7Yq5SxFf
QQDSDXbQ7Okcu5C9ycydIkS0Su8GNTACS+rl3Kq3b2eMu+VV8OFdj0lMkJiyuY74/LyqKW64pov2
3+9jdQTsfI6K2ZyLqMm1kp03GoLf3cTwYUpfZec+ZO/yH4ZcHoD4gtzU6LbC0sFmkNHDqJ63sE62
esUifa9uCwNA0G8abtlcoSMfrXhIT3lyqlJh9a227mhhYhs7E4+grM/yDpii7nOLLuPDcZOK0ibc
l8NNf6hUBRZtkm11IZMxvExCocnbBuMhO0BPsrxdQpOUHaCRQ8be+ilTdh9UwWelaL6H4f87WYNI
8C+d9LYacfv5i2Hio8EQ3QY7e4HtkK60mTezYLWrPp3ipnoH4uKEGCC27CbzEiNbSHzJ6QrkVXmT
79YMCewU0VDfseIx4dVqhweuv8h2dtnRjgnC3gHjrEh/E/ubfCKlOu7SeXnbNdIEu/fSA4MPKpoG
7+G3o+GH4agOF63rfKhVyliSduzT85e8moA9x+MuC8c0kI7NaxPE9saNTRyznFi5iWnSUByha8pK
du+DDunl1hP/EU8hlsGsCSpmaONu5keS2D+7sV8PTN1nK/8fKAtF0QsRjEi2fQSSVX8m6spf+Q10
xeLiFxAFJKaIV02VJ8Q1GjHONp2CuQJLqSlrLCdTRMkcQrZkyXoJxwppB0crY+zrkmDtPDhrRZQY
wHE0DBjWZoPdC9kPk47jUhRJ2YJItTEl16FRcuTNt5ZPdvF8XTxr5Tu0sdkAYx3WUbxtsxXRUA3Q
gg81C/cExdAjFbRDyeQmKvt6xfG8BjYGE0yhSMrozdOHz8ffOrzFajCIWonSVOsjqS2odBNwwJR2
JUe/2PqAV73yFZ7TLw8WfWIYIZfZ91S7Xi66e4SJRlfK7BDmXxd9PggoXglRVDniiRJ++u1AFO3a
aw9mhK1JtwYoENTpgWz7r7vywtlAiF4fe8k2Ze7xxDZxIQ1uKS8GOxuxgn3nlmVihTo16DjWvcxC
0L76FvxNBiUi4CxqsOjfo6EzVaxtJK/2tMfHOe1SZSKq20+iSDT6EAibEGtHr30jDDfLbTrEFeI5
oOehlUoYRKkumL7GykJcSHLGYz5sHsIdqJT92UBbKY64jSP02jvhdrdrKwAl78eC5bxxecE866cr
aGlt8Wsyn4EXBH+FxtRMxRN0HqdPtoavlpLeUjKf/TAvmmcYaJilbehD0CNEruXWwIIlTmfvb9IA
IdLfMCYcYGuMWqlrcb5W5iB/XnYxiTtAX1kBKjmHPh6hGvHitEkDpfOsNygZUlyps+BELd5hkPm6
fBDsMuv/tMF9bfm7gmNXFyhRe4s2d5+e16L8zRUMkSG/h6yD4JnXNNg6nVzOOFJjqnQ60HJ5Jfvy
rIzYAEw3+5oTrLqgv2NYGS+znu6hQFGe32+dPgc3gaKzZ/a5JWwt8Uh5BegOYTK8i+9e7V7EBPkD
zDseAYIxhzDgRwi5xMz3EmRNRy1PC2fr0RqATtFWfePAuElQeKefDqsH0GrIcuSQy/KbIli0uDOM
6xYi+aQY/FCnwMhfCbDuQnEU2BPsd6jGrTX7vGOTE3/BuVUIvOFE8fVp+6SJEcWCkN8TFUhGo/FJ
QRKqRrCnPFcknsDxX8Rm5EvqoH92zWQ1ayAZgZd5HI/Pxkx01LWGrkLfFclhYyEdI/cLUy1x32WM
56ixPRT6OXa1yynQpcMDaIWXEROfb2tedBVX/sqzTQPWlsYLm6bHyjtnw9hmctP9fgpUC/b+YTw8
Rxy5I7ysaDNy4tmO6n+FFRLyaF5kGSbNUZcWA+s1K6CPu4TT691GdKHvBstlf7uPCzLWg6Gs1P8T
OhTqHVYt7hZ6EhMJouh9WKVZMbSM16mrk2xCY3S8wiZXgXBVZ5tQZaEQF4vkLs970VCPfy9UVoxt
iQ9jUjzAr8tjl+CHTD9UEs4SZCAWwwHEH/8vDAUbpotBc0r0IweKvDSj0kPRPdYaKss+fVSh23kR
BwdEr4V9osxLLdI/iPikza8iYu63u8zycIes0/tHYRgSXnhYz+RjJxu8rtqrl/wQvVbKz1RBPkfB
Y1IhTZGWviELC4K2DPTFxkScRLxpHXR9JqSZSX88scUF7OA9ZCSLa9lL+FFWbOjo38CVvbVzL6+C
eHCSx9Xt36mH2VeotftAkKLWrnrnDZ5KPKSIZuUtYQdKZJ2NS5H6VD20DiuKOqutyVfLIvEDY7uB
kqhG24qhsDCBqyIzO+rQA4qtpUjICwbvpJGjS8+aj72x9limVsEPbV8c88NQJE/R5uoRTMNpH5LL
jLeIjkwCwZ4r1TwpZV8MqAQp5PBcVVY7xlbXnXa8WBvjEvQ3xlzRxaOygWbAby02XL1Ux35Hvv3o
/gFaktB2EYTCzPQmbjOyZVBrJ3N9W1T1jYu1a/c5yrfTjYLEVimo2xkzrF7oYdy2jTLniPBZHnmE
NS+01L/ewFQgpHdBCeK+MbkyQ7QE5u2Z2Ej/Kv5zM8JC2IdWGQ6/O0QGyevWonjrjNWwuaYWcL0F
3gSoGwp++7QDJkv+TSCIfFtjOFyHfCU6pidL/xOKARL1G5OarCDyjQ7cpAZe8DHBvTmmTTGDqzIM
1bEk3+HZBj77VGwZU56wEfsx5/HUSC4+KxmyCvB5H08sWYZ2/cLe7Y6jn0WXuR3eh9cxK8isiNxS
oh1/vMZAFUv8MiFXSSGwXuUFPBVA8+GpqLhuyh6awnSw3c9A9/4+AkSjTJx51WLzfJn1CmsBph5Z
T0np6kZZ6TTtgIMvOxU8m5XgahQQtYRZqW0M/13BO32E/JK7R/epBZ0/2B2uyq+zvKeWncv3BqUe
QFgeBzVQJ7n+mXv0fNlDUwWrMjUQnjjkExwkIe9rULiar0RUyOt05Ef07XX2TuF+l4Fqbm3Mvfze
0NIty5AAm02XzAC7407GtqJ+LLD+IrM3Xz0K6dQFQt49NY1fWJ2H7iQ95S8PifFXaqgHhaArcqDy
h/dWioJgy+EF69XJTyop4B92dHyWj5xbptyI3VIK0FhmIMABhXzyCO1pK24eygjiNSiDXOcmIa8L
WsGRoo0wuPto4oQ/Nc1uVX5RT7/GDkUHkTxGnUSXjTGHRb2b3CcI//H23tbe78rOgiRRHMI9PTuR
93m2XBNUBzwiI3whP/smM9xmvOHx9Ui6d5fzoYgbQZvXRi3G5vZHeMihzEkEEvedpZe9OwrrAXTm
tOv4FGceyXbkir6UjTosFMD9qG/Q/De4TdQThmw1repDrjjBqUnm0hM8THI8J+0hE1SE4EadLLXp
SvaKsaqQq4qXED63xxV7L5iZcjx7uTsNEkcZthpWT8TQJJo2lRKcI70Hbm/JJOi2+xtPDlwJRtrg
ibnPmTFXm2VRZ1ZWBxUFoIuBx/wZ29xacQOcGI40kdjqpGOLo1yfQirCRqvg+/evXrD68DJ3TGQX
AnKtNkLrhVAQtbFFP4NhbK6aOxFBGl8o7ysEHWHLfrnvrBbRpQ+KsqLFvlPTWkgihvI5Vf1Dzf95
x0DQlh28LewsZKfK/GPq0ffd5fmURuL0YFWRJwjp6wq9F5EwXvTD29vTTyEKuCqBrQ9abcRTWyLW
OkFtdnKNZI7UfmcwZfT8+y10u8Nct/18JtnWOR2qgYXlIRqcKyF72UqmMwuOM/4mbYuWyQ21FRAJ
mszfdIXohSdObryrv7BtuSYAJho2cAc+En8JMJPkvMHDZcFsFPYI8Bbj7/wfhp1V2KK/C1AeJZeu
cBCtCr5ovYxUTAp6vF/WlPYfC3AGGv1zLfh3EHx3BzeqtRcnoIi7FI6On2OgnGZGmSJv0BL20t78
wtzi06s5vr1cUc8ySikH3KeRECWqcRc5CreaRzc0V01dELBEgn+GcMc4q0hEDm5UD1dGS0VasomD
f/xA94eWPvSu93WIHp37/lmkIDSFcBR4xRYcZzbJKIA/7svjmJ9fK67Xxu4nBmRj121aOfIeNHRW
C2TukivD0UFQWoS4tIbVHPlBZyoED7qFYoKZuLiMmK2Vpzv2MhuIX+PGkzmbozOtkoFnZZS+AZsi
bmr6PVJTNjP4EAXIfShjfVzZgM0wEJr2sea/4feSrg/INve7jyBs+ajclN3OoDXDzG8WoJUiWty/
l3jbo/z2qCOyaTBDQ5BODWJB4/AXZJIq6kyiX/Mt/gY72Q1SvZVIbeGyFycVHjxhftfBn6dKcHpL
ZNytETWow+2zNFE5ChIA2Olbv0RpZxiAQ6XrwvnXSNizYI7ngJefqm3QLn00FDTQmyPy9x7TN7T3
OicFwXWf129DELwJdtuN0NOMkdUdfWLFRGEQtrbVsuBD4qic+PbT1df7ol1nSWF3sEghZSUhM/l5
CiH8uw2sqh101nDC+Nmwh1xD2JzswbDbP7N66J44nfaVrPfrbdlr8nNn1eg4TzMz7U8Q6A+P7Dyf
ngCHOdADemOtTVaCVyT/B/h5OFMFyHoypA1id0LobnVMJM6WtXL6Gfi7iyW+0nrziUOVOKtqCzND
FiEVQrbArLDOyufrQqIkriEGUGEOs1zwIXQkexn26tx6v4OK/kUB3yBXnj3ToV4T2/Bi6LOrChY/
gMlhevyOzARwzuoS0sVIwI1pdMdYhawyYwHH5Wb9XAUkwsDomau2gEnWNBIgKYl1XnJKhoUuvGzE
S15Np068KXcly7eCgp0dtVcBBaF2xuKfi1K3FX2/Ir6+jAExySlTSYRKnbbjjM4+vrRc1WNPN2ot
ABtQiBRFEXjMEPTcoWYCKEDCdGk+UTlKE8ovggw+aT7+ho/XkJToNIm4hnbbhQ9RBH7MBHEM7oWy
Zw7w0qomClf9vUchSO3ijST06A8yrLCXrt5nBKkcU/J1NvkPXlACM0qSAhd/nHL3SDg8EpXVaFEn
jGYI6Yd1JY1BToVArFNmAmwoVI7BMua9W0b8/nW+mwn86ut0/MwAl7Q3oTiXw+HEJgNmck/T+Ipj
MeWTAt/ZakEtGsfzTwskNO1gq/9UPiAsNPuH1eH2RVTVCdXZCcg/bU5g/vVS2UmnJywGE4wzEzgr
ftTiBMChnj+L7oLP7WZ54TBkzyOXh1c9fuQDdSdjyfRDRyU5RkDJ5Ct4f7ZIXTNk6jghZO+Rf1GT
VPkmfxU2pZ50addSRs+tSyI/m1HwajcPILraKA2k9vuKXSo4bOhRM+ZqHXlI9LAjYLv+Tm+0rZ1r
rht/56IZfZWsli9h/n73zT6F/3EpV8JVz+uJ/++Kfc7v+qw5TBWEBA/z9rRQpcepJKle1YDXEtQ9
/2ivwXLfXfiKnn+km6eb0CNJlpRQICtSJwysc5n7Kzpc8/BTFKD08nQEHoBO5KGrz3MdrRs49a/F
0UYfWMFjDQIdNYBP70Wfwk3BEnXbPlcPFtOT0oWVrr7oEV0x2vFrP8PkpwQ39j+ZwOZndgQp+LZh
5DTsMox7qdW8brYRgnD1zYav6tlG+jrYa5muvhdLHh20bUfAubue5qPDpGbewbpTmKSTbphu6DIB
O/qZl0FZrLW++ngJNT5WGo18a4KHgFLNtCb6h2BrRIQsJFMUbJPDuW9aZcfc5uF6IVAKxuoHUble
qeSYMzSnIpYoShFZo+RFNYU9A+pIR7P+H7U4FoaeFV0A1DF0zh80NHeMUHei8SwP+BlHGMIziXUw
S/8BDedjfxJpgqAippx920SmG3y+og0XRj9CEwuV2jJuE/wuEfZVqVPL9P53xg0BX/Ei8D3jtj/e
eov2tzQ+8liw+I554RbfZy4g9P+iFTku2P11DGB3fOJ7vVBu4Ssy4vEwzSGVf8K8lE5NLBAVt5j6
FGo7swxQpWeo1s33qp/y2gbyfGs14EK5OHWmQ//f39DGxTVqwpptYup+O+84wI8q/C3ByJnM7WYv
mQSM2Qm9VO548EZ1yNecri+vw54/osCqMde2WsLtQx0V1EbCRlgJDtXRt4JdKXlPKdWZN1OuH9EK
wDdg9EtS9qKDsrGNeyDz09XrpvXRm9QihY7ZPD8AHJqZu/Tgzz3Smvl3lbxxNv4W8nkte7FKztr7
VJMzZTpbYiQqQsSHG+19hf+dmMSpx6f3eGLvwcu6iHrmtfu9CTdZKiwwTBR0Ju7rzSrXdK/6Mkhq
9Wf0fGlyKrXTWjGYAAvLYFfOwmC4XoTusVR6luLOQZJv9vCUBbDwc4e12DbMG2/m7lfJSNdSoM1K
5RdLVcKuIc0uvA9XG8ETxC8hNvhpkc670IruBJXnmAcdPlxVwfatykCvxRUcDZYGxOeX2aPsv4w0
QTAlolMEAnGAmBmhmgqCXT0MKqpigE0nWjjveVeLFbuptDSOG7rsXrrkepGv38dnVi9FzUdCOqzn
36V+vTcE178O1wgVFnMsiETbZEpEeE6qYGdXNG/vxsgeHHAHo7iWZDURXj+/qYIX5znFy0NsVZbN
KJaxlj355P94iLEAsRFvwKhop8oAspQQxCnePjkMn4vrHZN8loj8AjoM7OIY2QaF3V1Q82kfBi+5
du37mOWzV1OHtjzaHnQaDm2/UrJmhCpRNKz9qvUCu4+WlX5k4+xy74GoJ6LfKXpid9mEoSO5Yt2B
3xWyThINXD685W4CgRGrA4iFf44jpD75vMKFgHvHh/WiY8E2NvcU+Lff2wBXNs2bZrWwL/HuKx3O
xPJ+akmYEgl9kcXlBBQ3Fo+ja7lvrAZ4d8Rg+byazoA02YVn1sFixEQ/1sZoAWXFfCUH/Xjv8Dnf
6xb0JPIB4/GcDPuqli1eBCqiefuC+B5YrCEjQWIhWv+yZ1Yd9FhQ4BuOSM7LQ7BSfI9AUCSfXZxm
RazOx4vl3x4io2SG1WadJa2fa2vGluJHrdy4moM7kyytwTlhKaq3RFn5e/qkboXsfk5eT66pIr6P
DPsL3pWZ/jmJY6XLapdzO+jRK0POgFmv99gJbOXF2rX3xlB8b1VUDtsQ+xjeC/KxTTxG6Db+ZJP/
eOmami7QzYf7P8trw/Ec0VvaL5SJhWL+eo3DmnP+ebbzzG2UpwGPnSOq6Ir+cT1OLGvi3LmnaNfK
Kw68TDduTSGd00PxcMevlTTJkYe3ODu4kiuiZw9a0leXpjiAlSAR4X9I+YbPocevQ5VkB7x5SzQW
1vuvi7kQ487Nof4gvx+u+MgxVagytVQbXsknNE/KU7q4wBKzgf/CP1azPLxLzTKZ1SS0MwPhTB1s
Ww8MY+YbUps9vCDbjWNtoiiB2fVEADZccnjdOq9W4q3Vdv6ovMHfKOA45QkEcO+pAQHClAXMMazN
marBUmRjAwe9oTQvMLBprZSeOLhKuLr+NcBUjGIgLt+90GVSB1IRuY7jTUtrLj+LqJrhZjRl3PR0
PzGYArItJda4MylyVFg6L7MJARdmi+LF+2NC2h3QJeA7SJyuuhUhn4Ex1WKQC+37fr3J9udpeUvq
gc3Oq1YeveE+hRiJpJ9ceGCrqmp+CIxGNt0E7H+8eQZPbIqoTJz7SNME/t9XFbVZ5tKu6lvbQ6gc
Rf3CgOYrZCQfL0vpgbPy047rHiH7HE/ftRgdMBqQNTq0Y6IGPszeSl41bJrSpcctOfU5bz6w5Dr5
BuwcFR5tOjeYoi9O+IEru5xvlBAVVwxVizZltXQV6WWMXGGtS86Urg2LVWbyw0nx2RIf8Y1WXGHd
aknoGUbrVr8zVXR97Ox4E54WekHOzvUzUKLKpYrWpNNcyLul+eixTxcRH8fVM7gr2S4Fknx9fuyo
/Xi8KcEsXr0yo+9fE0/dmzHpMLhy8RJ30pJlI2/axK4oRh/MMmnBXRcLKVbYqo9ZkSGYwy1bEqAq
iXg48CEDsfRDSeInUvYaenwQE5oGr8zzpvvi01Wt/zSqOPWoiSL8tOAFBlMH5CjdrvlAEcYkK5Jj
9te6umO9vZ5mOz8/zpcSLUUNFy7vn2afr9zM1OphwOrWRgekFRI/9JKHdA2IvUrcibm4uh2FgBKI
upPg+Hy2x9zPp5EZ0ccM3zBDjXaC1xYehViEpq4WPgOzoJfFa2MFKsnTmzCOKns2kJXP6FHjFU6J
IVJMpU65X7xwtydXTuZyRo2ryB8zWGQcU3ipYD1Njuhvow9k3WhuhLucWSqvGDl4NxwhZzPzmYLG
rvbSaN9E25Y3mfWUgTmuQt7Lh4+rztBlDPI/53Gn7APEDYzyB2iR+tfKsRyTufpQ8NrUWlmyJ0ne
W/bl6odmd4ll8Rpfoqc9iX4KXLCBd8u8pveGzzSjji7VGyDm66HGtYU+kjH/COO+3oUz096eBviV
8pc+Co31CypxJTypqeUdEovysXEtXN5bn/d985eE321RQZFNAsdGzE71AVB45ifzX/FeYtz9wwrq
eBTa02Whhy6vpAYTJx7VLLQ0fpK7yqlbh737E10aCAVLlBIZGniPpbCC2U/z24Ktgfi3rtaFxJIx
XSJIWmDI81KtSDeP0lSm9I2MSO0f1zLbEg0aO2IYxChlS5EgS9XV5QvK1fAKu77KkOlfmXY9Uj59
BA5vAOEaIUqphgM3jWv91Z4G7MntkjTfxg/v5bCVq5s0HGLgXdTX2LX6F+gOBkXiyfmdLeTRK95J
qiVoVdsi0NUejniXYcJ1E1UqASLII5cGVHPCc/q/JCKGyBGMZzGKFtASxZGoQFwyizyvA9Pq49zi
Jub5asdHgF2wYnUDyAdabrgxoKyY9YAji9wLDfkBwPB14eqooizuiGv4eG3MF2Xg5/UOJwVvqDxc
MCjun2qR+k2456DhbuhEuFUV36QYD9yH6Ejcy1msq4ooPN/WiNP++urHZzXeC9wjfhHpAvA69+ZO
kEimcs2uTovV8HAPc1oOfOX229X7+M0Unuj6IbSQBJpsaMyLcJ5FEbxfovy99MYB9V7P/v+evKYC
lQ1v1ybCY6Y/EFVSeWUD4unFiY3CQEmzySSTBnXZCQcDNCOqWDoGRGkdc1JJ5Zm9kb21DP8hCBVz
XRNbMCWf3SelfxKkAxUallzWmZ1DIR/XmXHDfSdjWTSV5djqmb7i0ZkmrXiS/WAke6CmXzO76ot8
JyjzhB2fTDrVL/3PqtdZlPeaex5wstg63i9xgobGuzQRsxn1Ykq/l2sGU1WYrc9yT2O052XqlI3f
jMBEy/UG8+CtC+hNAmKwX3H5CJ6d81DHrn2MjUkFm6U5pjVTUvSX7t//VcXQUbexF1vF8BElzOnY
041c1cBVjhqYEW6Ux7oj3yYU5wLLe0B/hHibhWM8uqx/1fhxkQG5vMEZk4G5rVyXAsVkMVMBrx4f
IdaXeDSwVi7CbFcZHVIQv4Yuk3IXElJ+PMYSlpecfi7rADvLne1Hxc7WdEEeGzJmP/5dcU3vEIYR
2Aw/T/RC1O3E24JSg3XNC5eQW8ATjE/yEORLKaeJfFOjG2oavTCLcOHb5IpKCfYmocDNDADYpmJ5
EAktXndRj/n3ROPdF7yS0CoUhSkrgeImGrZMfTirUEtbJduzi5fIatjyoIpC1MsFkYxiBe2Hbj3E
5bVLDw4vySKwdW3mV5gK1/cCSwva9KlNb/Niou12Qausl7kcDwdcL9DNvtviBFyKgA/bQK4y8TFj
Cqm6sDBUoCMpnlNIIK2Z5DsyAj5OAyzUXUn7zYC2oRto7E6aaSAX29iyO05QmLKI+DnfxQL5IyCE
PYwcrfwh7tOr77ILDGQBcAdVg5zfGsSPrPt1Kzg4CYnsPLCuDjHiXOqn3Z2trWJo9jinZ1uUm10W
ABvnYl9mC0VasO2KBJizLdKNce8Ey+sml8TzSUu2uZ998189QIVnHb161uEHQ6FBVWbsb+G8c3Qg
FJB4MEuEMv3bvXQLQOhARU4UhGA2KOO41ZTqRSUqUe0Kfbdnj5Ye8exHmyELpvDBwUuuxUwWVKfJ
Wwgh9ysGWE+dC5YwK8KiMpZbD+E+ZhTuqWoqQVo5CZB0lKmF2x0faPsIFX5SNzhIUicjrYezFPwP
9IOWYN+VSWjwt6vDF4Zj1pUKcDN9/ZrIFe1fGO23SNoZtaJJ3QG9/TaeX0hVmB1ErJHUAD4dxj40
eNfcV9neb04Blfuot3SY5zSqJarUrzIU3Ut8jPvWs+Y0GjnV42jZZ5kCKkqrLhpG5C48bF4orI2X
vnTpl/tAvQVwqVQQTThtDBEcNjnSWQTHmxFdsSKQv2l8jHWuVqfcPRG+FKTlCsQLXT8+9LQU1c/N
dG3XCcJ9qDhDDwuktU5jWCUgz8ElWQAusrhZJhvHi9oAa/UCFWQcPLdWCZ2+upzL9EKOXWVMjY8g
KzCHg8tyKdw3iX62oRn8r022Kqz0hisD8l/PsQSLWmbW1deTaz/WZGrHMzYX7JhEmcj3szS4RG58
xukSXohtkvyJxVAIapleSZNarS36DjlFjTMvfhCzvjmAG83p8HgMF+DCGilJPmkN+d1Xx2PIX1Le
pZKMDhCRmBeMy1gjNzazLzR8kIT8eSB0f10skVV5SOpbyTW8fim8R/iCNXOnCGW9xASOCOC69mmn
aWDg0TGQOVo8CjeQ3REhvU9AqPfQ4O5fJfjDwrwHHAwXtHWCzFtph4rAjgD2s93dTb2wJuuvojAz
AZes5WcJLU3i3Vk4eytrNbP/ZCOUoIK9VRhRt+qa6rR6EGVva73EjiHE3ac017FTTx7LlZBagNiC
nc7WGDtM75BnBhM+q+SgnBbQvxZLykNItMvXLSTlc+IK+DGhAOFWNlx1MlmVEZC2KdMzlAFN7QFJ
yTwUfddO+DX+Ko9tjgkJqziZzwXrvbjpizbdzIwVm5x/zWq5kgMFhpMrRPk3FEls27UHXDrudJJ8
HXPHMXJS3BuRGTRXVIwf6lJe3O4SdvU8naUdkUWqWEQN7wYX/yMLtnG/3ojUjdJ42ynWhC1CEoLD
WvPsRldNmc+ORLqPKr2IuEnS+OwkFRUKn81qXEJ9tQwjqcs/NEA4vFzVDiv8RhKSeHctqBaX2ztC
GVpgxETf4Jr2+Wt/nhgg/mqRol+bABrKELlAEvRxUUWQltPzXqi7VaLX/h3WOvPO16QD0Bvo9Il5
7fuH4q4A4eYMJB0RUKoAb0kwJcx474GX0GO8wWQu/zzkgds+uUylsFivX+7XLRCEOlQ0lWyn168J
7Y95OLJAKbCE7dRJiiSxDRoAWJwdINyWr4ATipTsgsArsT/3X/EQcg3yqtvMV3HhcoW3FzFegtaz
D4zjbejrNsU+DyuFR1xIOIZGERw45HEQgE92qrD6VKa0VayrjAAXvjMgCggh3lPVw07sp+cgYtOq
2A4bHVlvBbL93cpGirXlRSjgk3EaXZ7WeiHlqBomxjnL29/1DnPVTlW1V2Y0E5VZ5VVOd9yECHLy
X890JK+O854/XswVeoehyRJsc5uob8s0XLi6IMdqNgCuIBhiImgtdQT2k0wecRQQkv2Z3Nq6DBf+
yRlTIqOAPmIqVxyuuhIRRUl84LPURUZy5LqRiU7nHV+yPHk/Mebc6vvsr96asPprZKu/3wgTKk8X
T3bpjwdDs+u/SFAQILp4rH9nBnh2rKweB1uaGZSxuXyzwHxaAkE7DY4qlKCtAmY/h/FZHTwZwfYN
Uw28K3ccKnUE/kPlQHknYcXw52KcC7GiPOlXVID36yXZZswRxPBoZuvBBG75+5m6/fB2ss71L8ZS
Q83XM9biiWLNopJHmn7Z+nb0eK2sdUaqI6W7z1ASCWJbl3nyMDshfYlO+dPpiCikniS7GDndLf+o
gq3S2xxPTE9oabUj46bUwLLS50/91uDRTPNNQbcx6gLeCzXmqr5MUPD5w6gXlfGE6TM6JNq9s4sR
37ZDkFbbf2emZyAqTorwnp6YgO472QVf69LwuRzzCL217hwGF0IOdFEQaCb2fjlkuVJ7AZ0ZiTkR
OB7sh9IyDIXXE2uLiqCu4wl8ELeTPra/A44CCxy/Rlwu1Q64cec/ssbk7LWpI9dZeBxSv6809fSn
Bm0p5j4dSAZF8WbWWmzq0YiujcvIbHRzP5ztMcYUS8zZ1qsLsoUxPEcpD2ozdIVdByf3Okm7uZqZ
WXONhT1K159ENZmd5pFLhvDyuTKUB4eKtmF5Yg2jhaMqqlR9d8qKXlCYBszbW6ZhM071rGQ3uaS8
Cbg734ARSaXVENo+D6oxnZF5XnTDWVakLkqtvd3/bQNYl1Lo/SrdYXX15RerfmfTUVeG7ZL+XSCj
OlOjYWuNhAK1qJyXachHMcFfVYfuekdG2/zRwGmqizogaqaVa3W6eqXJcbO+Lbd9uocJlCmpruHk
2F8jWlLiBNEJmVHv8OZtl0cLgtb/y/1BHls2twbdHoEKPzA6wgn1+KrjqVd3K5GwoncNaZncvRoM
r92apHedUOuY0102MfihHicOP4PfjguaY9X/ShAL1xiOTc0OxiRvPNoq2o7140zj1iuOPMhEUNpQ
h59kGwU1Sve42VscQzjhGDnIXoIgxihOJhf7eNC7mNIQnArlVP7rg6xK4TKQCVBJsQMkDw0S7bNw
3egbVcbt2kMbNNSWxBu+fvEJnfjjCymZugMDg7yNDUVea6AY6vq7vaF4EEVXWzUsHz1v0Bye02dE
0OOAatG032yuOU1CPbBbykriB6/hPDVMwZkS/wU3fL8Z1WHRMtTFhD2gUWLAUIaZdoYRBcPLlD+r
1v0xbdR1hsbS5jqtk5lD50LeITLwovm7mqZ9Rpb4uwi1DWPAJtxpl2tnr3qvoEefSZW1R3Sxulmw
SRq7w/SKX/OTlj3R9hqmnpBiBlYEs9FTGvcm1sPhQM2P/UfiqIvEL4DZBd74MVUEa/g8ex9LzHVp
9a92zyzZGM/b1d8wzSW94C/3WRwSgRPFOciZMCMlI1Zg6q6/sOH1iW7O1WnFkrPo7qdajSRyiLlW
S+5u8hmuQx30VD/s1b/OxsY3CLUF80uUAckbp6qCi96rhdZcch8l6TownqaRvioNpLPcBVCNl6cq
l2mKkV3Jd42mKaKYajVN8rd+ha4TgRzTfIUF+WyiUWa60B7bJUTHV3hQGqK8pdhaY9aWBnSyMwd5
qoWoxFdfkspdVAzfA4M00g7fmWNd+qFko3vTZnVpnRRWB3aYHp9oDTE8ml9U4HlA9cH00KKtRwze
cDOFNpJkcyV88D2g/NUQTa9uIacFS2l/Rb/7sNJKv+tMjYvoJn1+4irIUM9DsHGNatkqoATcuEv5
ge5+BTLRAtTiazuXs6Q8qCBW/WtM7lp1eoDGnCw71SLNxnqC30MZKavFKwq2PV8IBYT3a595jRO3
VeDdpxJZmCEKT/nrUnL81pBtLy/YYfFp0xkXvQfo3xLCKhxmjcS/JbQsw8BxVvjt3lq4JlAqvjjj
BsDvQpyujQ7rOlx9gby0WuICjjJBcxkVKqFhKpILKmmUtXL67IZbe9+r1pyhQVnxCpUOVXElpSBL
5TEa46gdkzcNzw+/XvWvx5frNnnkBWnDls9lqF9mJ6nVZ0E7VOpLBS63s0lwxd0/WfjH/TlajQb+
gf5DkiIoT7iJicP8RnDDSI3kvZ+8fUrkkVYu4/IDzRS50NemRaczSycSPdNNjHk7UvkvBEA4aBnR
6FY0Hw7xQ3qtNNijbJoN0KXfBHrCQ/kBZgz2os3UIm06zBX8u2JEwQQkOFU7kEOuGfVf/+ZkjQzd
QMfe4vkZ5ev7GINXZM6v8PqOGnNQOBwcJphjlMuAlXx0mi6qwy1Q01OJKIJhGmaE3cbV7MvgGwmE
6CK8CDE3B0Kcug8HKRmPV9T0uPkOoNWBozuGk88TniQ0bnMJEosbl9vfEkH5cyooL+nq8nMt9+CO
jIIo/OWIDQ3dZSZEKPOTIS7tjd0CSjyJXQfg7e9b79Lhd8VoX9VY7o0922rChTKC1bFabISVPUMD
HxxWJJKghongB2LP8e6F2EFQoT4wKhcnkgnXz51vYY6J7EN2XBQlAM5N0P1FwOjhHWpUhXDSirqB
qBTsTYqphwJwsokxvRkXR2oOw+8UEwL+S5oFdzystmCzQqxOsI5hd7UjF0ipy9YdDOIv0uGGWLr1
ODbmXkgSYcVaCKOQ+UZrVwN9SyKkfESoxAdB8APaAyoPpYOvwPJbG1+gx8LlnQaw1J9ajDCVSH+0
2iJkAeZMl/XmAvkjvAra55IuDcNRVFTLF6l+l+YK6yqIqMQxXAw2elsbCo2dOxpH/eM394vBPu6V
gMut8VsiHacv344ZmaCaKRK0UOohmQjHGYtTvpp4f2xDYTF9uiaArubfi1UFO09hNr0pSR+YRcfg
sEOct68DMdvkj79wq3fXp6aD15DRD/5slUMwp9k8Wgjlv6NBROxyUX9x7oq5p0FUljXtPISXplWs
5SzLxdIeIAtxk6bDzd0z35aF6Lq1Q3tfTXqoJmwFiZdau/tzfK8BeZjAkxgLS/Ctw7wYEco/Uhcs
jmpv0LcrPU2z1FazaJ3H6nWm/XJex0tA7z6XwZA9dgdESBESyKL/i0UAzj/85PuVSZas9OJpPt0D
oSAD2m9pxUZpMZUW/M8aF/09rh5DLCyMSFG61Nf3YvJK+yCVjIxyrdrXzqTmY89zWamLS6CVko1p
7PZQblt5Hz0Bbw8mz5JtvsvPoUCQtTffiluegdzstVTwyXFB3YmhXieczQegTu4UIb1RG49/hriI
i/5mBcYjwVZLO8a4YmBE8YBWB11sKApOpMwT10NrqwsvWFwV0DqvjeNt45Q0+ikbbPphn706zf6F
bpPr9yJc20/GvCcfwueQJ8f5FNCT+guQL8A4amZiFL0usr4kPQUt42McVGQA9HvMu1n5d4MUczgf
CMrTAvgXVAaN7Mr9Dh8QVV2DNsA5PXGlx1Z0j/ywP0R3wsKIhIavET2vzbcjyz0eEXd+q9GEr4Mb
pxBROlSxzd9Tiw6baMYytKWR+sxmpKuOhSwh7GQAoEV7Gu+R4g/mthmKjeTCvzCZxsQpC3kkvVRM
coCpfU95PuxkPlZmZDHkU8gzn6s12oDBM2C7CcME299Gbkow2pXSys4DLewxZqm7UIhueAIwoeWB
3hDpQOWAJnaYI4zEa/OSmTe9D9oUe9HkaDLSbgr61XpigiVZRMJ1FY9vXKOm41fyoMkftmNo93UW
xcdNfUqBlacj7DB0ENyypnVqtJsKHSMQoVeV+I6fjG9vRMyrV2Em3gqqNPVEz1BixsjZa6FPHgAb
aY5FMerCPnK4pP2VWHcSpyv+Pbn/vDQJBykZFSAemdj/1I5wqxnFOVuGX4RV8GefNPDrycvlILfY
lkrV5qhGLkhjxJDKq2Jtl/d4OsnbkYuToHjrKvH3LBPm/hJxK1CJ7lk8NlvC/6KX79pgXEdKl4Yc
rVl9LUKQE4Kzo6XxfjqUiJ/ySoGAUSeJXK+heJi7pl0zuTVroecuakD6fKNta+TQJWNRWdUnk+pJ
Trzm4CQqF4vMG+jCCw2sRXkjl909LMxyAElS2+N69Jnzhw15KXahTe0y7Cz18GTQHggP1g/scWlf
6SgeK1ZmRytXMlXh20jp42X/+Y6P/piWG2Gu6p0WHLZGsjVb+f4mtzVbRlFoNfAtmwr0u0uJaaAy
w55QfSjMig0MIbQUH7I9R0BBTZkIGSaOG9t6j7KEeEdJb45HFOp1L3GEhTlpFiihRua109Igh9c/
EESHR/M8bQ+fFdqhuadq9qobgDD43voTygbdbJJgrUfFr0VGWRwZKIowGrE9grApedmtXDLcVIK4
A3ednith+Pad6qnfdPY9WiLGXHSENDjzOdj+Ms/8VjSE/1+h6k8Yokh8XezXNJBJSkpBx/nOgHts
k5Sbwm0+CL/9Omx+yRBey0zHHjcZ9Gawv1jbcG5mwFwXWH1LhXro9/ZHZii5jGpLlRTmRlPvR2Gc
OzpOvJKStKZ1H+GdTq6JEEqNGL3BuOzC80yn7KmNWIqnZGHgv797FvBE3/79TQZ6CSmrCxUzSb00
LT/IVRKaarQ8wrdN6jrEGU0kmsNMnjOCj51suqxjvJmKWtfwTN+Bxl5qZ9FvaJfLTm3g0u0cCnW4
i2qRiM5nJc5NR3geoLE+VUnXa/M88hp2b+i+VvUAFeMTC4ULnNGR3fLE7czpw3WGI2UOeifRIjex
HM4cMjTVKUSLkW3YOrr++7fzNljSPWIApWh+lL96sY+zSIqJlXLW6zv7boMjQF58MZg6ufDuw6rX
07g047JRK3QB9A4jNicblaDa+hUg0zlrDysgxApyAp7T1OEpyynWpRUd2/9hqyH1w+7hxs6fI3wp
PIiMkrRL4hLGXzlbsLRdrRZsC8l5xFL3V0CYEdEVEsbjNUhEyimiF81pu1Wmn6yvTvnOqFLeyfbS
AOvSbWzDE9+yyw4Dld6txkKniQ0blfLOPF85zHtfgSBXjMVNnv3GMV/LM7sLrjWVVBoDCpwbtrQ1
79qu5IY0nt1SHcyOfdj/NJtr6IadKd5f+ftvFrvD7yHFK6ewy0/SWwKAC7qKUr5W+m7vhDJ4dSKu
3QVeAadaUMFGKJwhFILKXDr+Pn4pSvswDDjoiDZPui031mbwfAC5JO5cHO3vwIUQlnttbjJ4+kG0
0VNUrBFBYTNwDU8Yr6ar3e4KJnBMZv+xNme2AzOEKNox4p5aAGousfu50doWJJplaTMOBhSQH7Ta
9bWRKqKnqM+XnIe6w8mlWypDHKpQg4FigPNm9F3/OPTrnhA54XY69zFV1mCbvZ6r0rxDYU6cbk3Y
f8KrKj26mKbMAPZT7pEtMlMOgjG1VmbnGrXWsp/PiTcHzeJSrfEYWI80g+FXaxZUNwm3uHeQXGC5
ByyZoj0cktOtREcCbkVQiopPlPq0qXP/JI3CbX8BugBGKalCXM7pXmrwyjAWG2R+m69loZVMYErb
jBCX7r7oNBwnhbDAlw9xHWk0zB72oXAnMoxzDR82h5QBVoZnrFswHzDhvm339Bu/dqFGiF4DiUuX
mSPrJickQQuEusCWD8oDER0hNoBhQgN3mfUZt4UBkpBNTV8xQ9ouyOiQJ4lERngBY07xvine1VfW
RAY5oa+u7MgUNFl1h9YWsf4lXcg1ErQHMWhWIfNwM/SMitXRmq13CXn4IRXSyIpkpWGG0SX6uogL
gwF5TCGJQhBa6oPq7vJO7K8v2qBRu3jep7bgd5ARPlmpW4ocQp3k8fL0B3jaoyg/+EsS8wm/rsCB
tULn0r9/Kn/RwKgBRwHv51jEazkhwLGbPKAbjWs3u2tKN9RAhCfV0wJRDWQoR5yY3CX87yCVcXdF
jG4Rkn8+jZTTgbi/W+9jJSxVe3OjO9zzAGH9s9kOaLTrGTdDgI58pab04MfLMlUIzJnUdw+XJkpP
q1qeIpJ9KIUtsqYsbzqIC2YKPweTW0eZwzEZsEIns7T/Df7EZASiS4JlwrkafuH7eZEc5t1gPqtv
F/3zZuH2nyTAFBH6Kv1/mplTKQcvQpc5rTBxI1JzJ04hhNN8hfA9OL89QJtdT3MPPir9ypehl40m
JFYrIHRkGSnGAxOVEGz6jCPeuX8a19hVQNP7CZmSuJzZ8pntvdZMSZ4R4ro5p43oJEStpVqLFSJ9
cnrdVha9MVFzdoL86b2qUVMDpP9WcZE431mG5VOgcYw7fkzV+A+GorzxWw88P/eGG0xPSOQZUG5v
xQjHqGma2R7vsaQkys61poJnl2Ol9BsOz4wF2tGq3NOP1ZUqGnc4fGj+wqn6PKi121ySr82LGUBq
VcZy56M+nx3aEGteytytmeEknupx5j8KeiFnbOp3MPYKtrP/n4vWCKS1TnaPVWsuxdcCT1QMCpoy
5VAa0FVsU9ZRM/kFJuv3i9T08UUfQkaf9w8EsInFmUUXoPV0hsPjUAtYtdySZtX98AmvMMZeZlhS
c+boNKlbS433scR15FhrExfxouQdWhCZEV2O8OnJL1u9cQd7Pafuwy0vhOnuObty7l3av8jSz1io
saARVQZTZ/CYchTjGVeaSShHCIAK2amn9StC14s32U3t/unTMXu+njtodXA/G4rzAYNaZtJu/cd1
CrGdUeje5/JH0Pqxl1oQYPqZtPTfgARzRnjuDF8Cscy5ZAtVQyU5KmLWHK6jysdcFodA61GbjqCO
tb5OENjRGOdRYwLKzvF5B35+t3ITDUm3xD+zwiKUfN/nQ1idJb1HGZTSuTe6RHU9hYvIQ64lpony
7SKnK/HLcj3Zm2jKIz2Bn/DmNnY7Pb0W3WAKbKya4JJ9zg/Qf/RUAtIvUYqRd+D8JhcQpMQn612L
XSa4dPXR+NWTKnuMRTPIA1u2QtGpvkqSrJQDyEbxYQi9wiNKlN8N80KxRdOKD1sp6HMBcw8IncVi
EnXQ9m16+XuLIBoZWJuc96eAXtjCEt/+I+JTG6VrZsMAD6b00IgBaKekbo5w/d78FRstkFIKy0N7
jun39GKK5GShQfZqZSgWSXTl8f5IQFrypQ426ZrnnONKn1ZlxY8wjfM5HnEHTUT6c/vnvZoMgthS
s9/yTttCAV243MY50P1A4Wu7zIHzYWh//Zj68X63WuCq1iaf0F8JkWg24OW6FGFm9zAQKVCahHXU
5x5vjmb/U0hBkYvDh1HDfTz/1BBrnsC8GhFcE10OqEYbM9AXPrn1i6pDc80gnZvobIusD4ltVOWl
QjQiAP1bb8kgrXu0CViuOrPZ8UKpGhjxu6f7iJxj9Nbv1hxKOzRW2Zgp7afMuA776wXtuBA10Yi4
2ZCTNc/eUbY2s55Nt8PjAeZESGPuT3aFpwZT6I8/LyrJAWbovjH7gncDpZxB3/zPnGdMya+Afbk1
2aN2sZOw9CBbyKf15nznFLyATMRnpDef8AV8TUrGse0Iy+/1Ab6FuNJbvoX6XHkKQNBS/GZJrbS1
dRvCjqgwrlJ8ynMIWh2XBUfQPJaPXSMmiB7Cv3hrATPdsSqRD+R+PUl9mkMuEE+WISUiXe8eEqyA
TnKkxGk9xT2ToS0ce3QrBf2fLH84n3pRzN1PbsBQZAGZiaCZSezGh8GArNJs0dL6QIqwD171AQRH
KfIIUP82ueHLHZzZ4cFVToS6qeqrG4WBAZYNqk8UK1JIBdHPfdv1RlajOVgxC7yXBwFaJ8SjG8SX
m4AhgXzldL/sAgMAlm+NTZZ/1CyOXIAfrpZnWL3XSHgUfoPDBFe9biu6sQh2FINLA7olhQt7HmA5
Ti8UYesoWsvp5Qf5ALtRedliYwzma+gqS19fn5zpbqwLRt65C7SULTkqkQvg7BWvVpnLhuBvMPRy
unhh3/J6EAIiGqvIEtdGZsChWxJnsZ048u3DBVg+wdsrps13dkTJzaOVxTAZchk/Ty2zjyrvnZW/
xE76C4JReVTICMFkmuHD7Kv4g5kHNANuNTTOdoUQXD1HGZVEnQCDKjZ7mGn1bzm31wYafZBq1tk5
0suZSOWOP3TsfAfekJ18QRhQBDdyQaH/BjFBPU/5pHaD+2oW9nSSc65lK6wa6A/F6mlmhKQB9roZ
k/PiA5ULQ+Hm1mHiXqyNtiHtMMvKDVgsoDcMAqpNYnltAYJSgxns6Xr46oa1svuFdeKMtRB0YQ4w
XE0muetO1PGoOS3FnfGhHbqlpTA7dX6Fs5EuegsSRZuoZtJRTEFgZhrmNS7ZU49COy31/iqmcAX9
mSH3lf0ZH7j6tQ+ooyw6C5a+3H7XetxIHKdK00Q66qjQtLGDBqvKEuW8aNgdL9OLnO1VmnmqxGf9
yDP7CIuXG1FLLBSo75Rn12qYvv7+yD/kNXaBUjMiE9Fken1oz/c/rYnmuwJh3aDS5Lgw4XbsxxOK
EDwd7bGd3ssfYc0VA5HXWueFftN3EihssafWBqVYcAYHSrgKw6w0k5pkBdu/1yjv6Q9Vn6ju/gfb
Ad3ivlmrCTcrfxiXFuyg9rAcsmhDOEB1iEzbO5jd+iWw2lq2na4DMryzQRV9Cyu7sUBqyf3Ca2T0
OwMjC21TtU36OecqxamfAKjb/dNoOiwk/oL/Weu03IqPiiPWT9Z1nSR/7hZYMgMPiH1S++ak8d0V
WaRbAuykC79qtZKsnuI7Ww2hYyEtX74G2dBpqNLnkKGaaPaeKprEHtZHYuZYEiiNbXsR7Su5HB2a
HP4Gk380wqs8rxS93rw7UlTiSbeyEGBDmCtCRSp86Zve3LX4KlRqOz23LIUe10Bu2D8eJ4RT0weW
aO2BZGVik6ym9ndaRgntDdtwVBSSBSVRbnjklyCgO25ZxXCp2OxqzEGxzAS4zY1r9BjIhjVnJnD5
Y1G1Thwd1mdTN3UVbcWapWBFkPmbXxv66PU26D80Z9mrYVQDNCocjaUijrB9zU6icJXXnPevphvw
kAz0fmpH7UcBYSRV8bbdHuq9b+mXBj4+LwqxVr3OrkO+PTT6Tr1ZEnh8JaeFggaH9JcgWkhXqImz
n1FGnAhrYaIEvb9VluuBwknKM/Jkt9XM7/oqCNjvcbbrBqhIsM1nUtiQQzLfSrHYnjDSNhO7ubdL
EJ7TIh729VQdCI4OyHlw0MLifKh8CJ5nXyHo0FubAQTYfdBJixxnhwLFwOQKELmfEultv7Q8lfqz
gn4fHQ+LxHIhLsFnL6DYcn4tNktoduH5FUBaNKU0ytJ4gxS4MjnKXh1/ppCvTtF2y7SXZv9u9569
kMwmOrpQL/FmDDjCzk6ogQ+OSTMBtMDmHIusvGdieJPNYZS2im1tjMLSOrMHKet/D2pPO/XxrwYF
53B9F8xIAoC+6gVgzAPzJGwmtI6aae/lBJ4pFrkMDB7HdXGP/7+WBiYTXnexXS/13h/rZoSa9FcQ
HDBh7FCAgVg47v93jAo2X7t5z2T7UkmTWTrk6KXlsKQc4rtKla/kzkfHqLc5nKTRVwfmqiUqyg94
z62prHDSoiEs7xx6Vs8fPHQkY51WH5KheH+Nln1d9lAcA86wD/fP0Hhi+vLKPpJdIHBoWPq7dxAP
o5zkWGmWYToO+NNY+s/cpoInPG3ojmVTCBlYFP2ZJGfgiY/bj9vvSaoP+rucm2HoQAYKH1sT3lRH
usP0g8q3a6Y7ECxtmO6YSCrNCgDpgspECA8VI1hpBHr7L4xGDDsSLM36KNLHiEItH7gFsxX3KvDz
oHGnAvKsTmX3cNYFB0Q1spCv/cCnzDemKSkTpPAax/c5hGQIpmvZUfzfkVvpjpW36hlG9NhWgdRB
ZYoI9BUG6IMal7LUG+My5HJQk4cpZ7C8JHLL/B/Cju2llTqRKbRwx7gSM5CIkXD3qdhfp2B9nmbJ
U4v5qA41vtr56cQ3JGMDqdLHv8jZc+D9GCgFuzftCwPAAJMyCtyz/0VBA3tYN/SR9FRL1aUAe49r
pY9P/A+zPwirqg8mTDnonmAPQA3VV9DoK+R+Kn/ITXx9YVkKidQ8M/9aBaoP2vM5V4Bm+NTxjj80
znsWnS08XCecmFGI5vT4Fe8SlJdQooSoiCaykknV0p8V58mCQwcjS/BuZoXzt4cCa454o5p9zlnp
+4VBJl+79Ok0mpMCh9VSdgvO5NhvLYgwFbDqvwHRXUqsQR5P2TzEzEulwnLzvGHjndI1qSGEIjxI
bPZqLXXhQ+xww3r4P2a9G1scfqqjeLCfaVtapXaRU9XsU2j8rO520q+d4B6iQNIRXq7QGyMfB0fb
ofWYbkz6k0jI9rvOgzEGHShePkjHzRXWGl1SVl1f7+pyOv53rXf9JgwF6UPdCq/klEO52gp4+Wci
lCxZ5CA/Bx8WLZYLbxoIwBvMSLZoE3x2K0nDHG+uctFVBgl5XaHejRvbk+/dBgJqeXlHveO+dwOt
qHFs7hdmxsX858F7aGfcxY8IVj/EEmD7/UCXVrZcaMXdWNSCv0SFiSqJNNICxfymlPe0HDmqQcsP
3a73J4FVS9crfaaQVYNDvFUaQXptCjPN98SyX5vFpCHvVhZQRItLflcrWYekUynD4+OgSAY5UbZM
49GUKFQ7Ct8ji5KGV3HxfNnu4BIz07dVQFVOXPTtYtohJ460ylmZMZk1aoj00kTxMdISrCPqXMNe
JCXcPoldV5QGhXEFIYvVNX6wZxvRUi+EVmC7AXkMI6qD/IlmFkvVQpp9wZIpFstQzBizV88YzZu7
Lk9Y7e1o/mbFdQXl7pjfmJ3G7FFdqlmezRt0ue2CcKYb9RRVKTVWoGiJEUkVXgqXHud9zqjMip+D
mJecGpZ/Ntwu8QysrqnblNpfZS7FKFVo/2F7OoExqeKyv3yjYKTKrxUa9k1rdF47AsqpvBtbmMnv
7B4d4fgErgd+cPh3Yf8TZhz8JqcdyDRfwKHd2iNU6+H+bl4TEwCfrMda5BfVBy3M7prvYIP5c46V
rU3J+6AV8bzVl5lMVd4d1kT9MBIwfgRORAisc59nHi6cNIIXcwQBcEJtshE19nNDLJdCnxGy+fMh
0erjnGZeAzzZQJ5lByM5rNr9DXYsyQJuh2vduZXDk5QOXJNAbo92hk1LZ+Bul6KeMeCGu7Xb5a/Q
yOj8auSmv95ecUgqameJ6ttNR2f7V2VpNIZQ1PVH5I2erOR/Pa6buRT4RLcfR+5fjWqf2DGL2rM9
RA/O1jqE7GMw8E2urEgJIGo+FUd4NGP+uPIgwwr+4OIoY92R3LOUjzhiKRD0rLuUk9EywAlPpvE5
CheSDEb1X5Ibx2p4lzgoqsggyF+5uA2TTY4qubC7ltDupBPNQhldBmtBYZAlxGclbK/LL/9dVLFq
stTPibv85abzl+a31f3ZfCRf9Myc26yzSucLrC4B8ge5RdTFvZDkE168v+oll79i1vI2INTpIzTS
tNcJdbyJRYeywDBdIOtPRiuome0KpocKtMvxd0dyMTsclGi97AtFoMF8VAltSklKfKg/BqtJGtPk
e521yxBI+hWUB0BpTWe+qjUumJBE1EwU1PgHh7TuFSfE+XefEUdSZZw3swwHQh2a2MYHEExmOl3R
JhiRKWjDCrKL7kUUxjMY/CgjDqJYE+XYoxOkJXwrCG8ut0wYAEvBIeJypsoQEsyIQqw/6PVuEaUS
Qt2i6S9o7EsSuOyN+MqpDBANoz0RfAsxPapccnofBPcqRy6VfvsJYqalm4pt12f40A8PfmmzzPf2
uqryS332IPad6GC4wQFFPhHl2GH0I5ZLPekL0nL7aZZvOkvGEfNI8SICl8gYfe3rEsxpxvOKjCxn
WOtitcO2aaJYq5ugDAxhgaMXrjLUc6Ftzn6GMOpoBuIibHZKeO80bIZqKaX84GlWLMzxbA6uDiH4
7nzfgHbWuytrc4YIJKFIGJd214F+l0vL3Srru+Lbm7mPHCx0K07DmGpJnhWDxq2FGpBrXYBgLjyT
HKEBQn4okgqgcn6CkLnXHG5yj0qqJPxdOAzy4Al5O0QESivXpniznDrHnlYnDPNnL+qhtgTKGowj
z8NcmcnFBqGyJpFscqbh9fVszjO8iMkNkejxP19EgXQpPAGKDRfFecqlXpaA6aOwwB1FJsRtl5UO
gW3DMgQnVQE5MJV5oGtbmtQiEr6YFUWZVt3YA7hnopzEGtfpEH1YR/T9mn0mStsxiLUT+nwYLXeQ
2s+u26E72VSa/sDqu9eJ4QHSC3Q3EAp5/bJpgxVJVQ4Cz1QKoMLcOhq/QaQB84aiDQUC4NReU6U4
zhSrJ28/m/vfJ3efflL+vIrBDril7S4wCRMUgH7FZFYrr9u8GD2ZS7Etks8l3lhRsH+HXbRms2Zk
/R00S/HrZNRriTPPyXOc1FeDp7ZHwpJNFGHDvLg2r/vIenUX/S1ZEc1PdCRlye12MSwfts0vV6u+
HPSOjd3e85QaiMSnO8kjZUvkxBb8TSBL6uYlzj2w1h6/BT5tanw8e5GTvFv3N68QeMWevRdJW0wd
G0WnUTULa7f2VQNiGj87C72/3TWPOGtZUX3G2nzinC5kLwRklEak5XdRwqR65kuAengCf3YnhQX1
xn5OE+cPBfkCKuaukC5zfdjccTBCPQPwDfLRTecTRaOouePUMwtoFA23LGPNKVwybTSScG99ZeoU
BxQFC2IwYKN3qO+NprRMmMkYDFNYk6EPRkj8/b5uvYFqFxid7FUTh/4e3FoBFy1bk9jqOnQbrnuX
+UcHmfJoJMCWgYdhFSw/3Za5rmZlpV8JXhRqTGl8694t+rs2TfNaH9KO50jwr4iVWri3OxBhEX75
ubnpwrzFnRhbWsFQnQqhed6coVwl2Ow72+mgGyH4C6sSZC4c8ZNx+niGL5TJJm0JGP8tHmsEVrSl
DI1cR7CzgucuSMHA/MvEwJwPiU3OxuqWyzzRbwWmXzQwK/OUmoGBO5w7pKL1pPR5WR1w33Mdax7y
SiQ3U9rbzkzcgeBv70biWkUtAv+IjNcqNVJjY911zgpwY7PQK2CoP6wcPLTHucl8m4raRvC2q898
kOh5ef3GGLxdFqsTFyN97wfeUPp3XHtLuz84C9Gtm39ng4PzsbAftlGzKiQjJqc2sgYEL1UxEgEk
E/CNslLKG1bpzSo57SGAypk6nvb58LrWIQfRW3mFPZKB4MxyxamQ+3nG+c6JsZ2h2ZqGSQJh0/jL
P8UwHow4H+lisp4gjmytLaXVwjdYFVMyWCi8ObSZFctC17wuzSr+Ff/Xoqg86+EoiLzIWxgGr0p1
xtIwTCXMzlTLZo1QsS3rzgBMYrsD0JURBhVpZ7G8eQFOtq7/2dQ1s4l28Ytfw9pg6gHG++9YzGyP
OBnQqk9x6h2S/uGj9JkE+BzlCyrsn7Zj84dR5V6ycNhA/RYIH9JaYzTcQexko70WPhwXhCyeq5h2
SNjn9DCalgx5k2UNqgZxyeoit4MgJoViIjoVGO1BK5EhgN98a/7VoXig0XWGkgX5J7mIWaOkj1aE
ijaAfL3PWY4B0I28qLWeEAGcBkwVggJeGmy7cbHPNotoAuD3aJdtNmpYtYh7l/POh10tRuNT7tH+
F8juMLhylQIOj/VLRrzJILoS6xtQWOVZE3f/aBUEIlqTMnrYF0rWj4T8HTxIZYlxyJqnDfwkOaMV
WfljOu3XRgGT26ex0HHuCCrYFfDekkzZZ2FkeekeySZVwZ8V3KyS9tmyvVkZKtxYhT9dDDK6BBfZ
dXEu5LBpVtc6I7V4mjh0daVZJZuZW7xmrRHZLV6bdfIgI5ahr0RtfwmNXvdF654IOGAsRfsJeI3S
lcjD4gigaROe5X7+BCFSnWwlVHxxSwuNX4Q7fK3w1OzZBf9VRRk5+ZXfGTtBdVStuMBjVkmVdxIb
ZhSr8NL+FWmFepDNTH2tTFIwCBjsJoE59fjC+U0R5LngQXc6Nk/dHO2dZ0EqNNWi7bkXzzS/db+r
UYmWugEiZgoLAlUgdpcR9P55nMDzCywgwVIfvAhdsSMEffI90hC8VhEtWZwT6AQYvhZ42ULhHYYW
WB2lWQ2gKL5O7NMDm4+oSKdSSDCfqq89VrxJxexJtPhN8++pixE6BO465lckFaV1u7zSqCmC2fVq
euqo9JeMybaGx7s/H9ld+MrO6jrWSJzSZ6Kj0zxe8g4Bj5pxntVcRUc+8WlxvBFGwVnfbFFA+hjc
WoYa7AWMbFhjgFEt7uiCOpMLQ1LPcilAztCLebqyGpvLgBpA9HodfLSMqjmIgkTVde1E47OHdVR7
7VE6P6Q7j+WMtDZhm3kM7oMQF3otsUF/ahSGc70NNQZvMLr1vbKbQq4oOkSv4bhDkUPhgGbWBkGN
HKKuw8g75cL98dL9TX/vnrxOHi9XFFICQwh2C81OPBLt+9pCBQxdP3hNy1abv0e/68ygH57eNSz1
JjBONvR2rrnMaXOmgG5G5Oon1f5+T0srC6WI+yq67KEkta2DNNJbkJ9PG2YXwlnPs5Diw85NSewC
RGLxl2lsuzKS7oqx6v6+cGrRlDuCvPCqQ3E/o5+daH70J0AZxCvAqHKHyyZ9zaHXdrWzloWLKCTW
Spx74sz8LacKVD8sOjkD29HET/zSJkbRL+MxFNPmDCgl4tvIOGdq2S10F6VoPREDcW/uZFdWHo0C
EHDgMXx0tzppOYb4Yys852jRiTo4Pqa1OLJTOnmSS3StxAeeAKGF5kxNkEc4JLgau1Y+82N8kSb2
ugDMT1UySZz3Coz1W6jlXwnbuePmmO+pvZdYRTMkUqfCSO5QGxNt1W1mWOwmg+OMXXD2WFq7wMat
Mpcn0fy/fLJyfmAFSgQ/7d82apUg4s6BBVvt014todK1nICdsia3cOdzA/EXnOGfFaIJOkKwu2MI
Yt+Lj//qh18+91D5xIs4gEdnIVgefeyD1/60g2rReJ64m0wilcDZR2tCZy7EK99lb59m3PUcp2vH
TW/ROzAZp2FW8u6tzt6a+mlNUlLtpQjCX1/Eg0QkygUiDVprG6xL83VCA3Od3IQm/50i8p973Tqp
/6V4Y/e/UjfwjKHL6lTfQbH5O94AGEfZpsHXpK5UvByAEwbof+ull8iDPngm+Okp759eOcfHorkR
vYBAPaQX7Y886JWib6MItQ2FrKma7r4qpqD+WuSGLaaP5LrAlKTBYTEacF3tY7FtazuT3oPb7NBg
fE9rKFzKE2+5lMF4c9nz8XOb0V9ljfp1dUF1wJJUV7assJ+By1OCvs+6jhkJLRJGcrYYkjoWC3Dp
DF/LhrG8rEVlJ5kNxNox5ymKqn6f4brKD/08ubwFxgX4dUHxGbyEmr/OLy6S5QYazoLk7RbWmtP3
x0tsYU+DZZYBoRhIpoc+9a8bkXVBnN++rUpJcxoSw8Qwro5na9Saxovedbplu3VQxdqsU9+ta84H
Ua0Up5E5Y9PJ2NtghWT2RuXpbaGCvM2gd2se1M6mG0ttl/ni06hPcZOiFwk1qxsqrhbt1O/Yn+4A
iq0t2OFngM22T0HQtZ16B3cz+NCyjwZw7qNzR62wdtTKeWTm+MAVqei+ruhwRCKMNf9f2ANzptxU
G1c7fDV99O/b5GV7LjJtsfcZS+PlK0UM8MK8SiVkuXcaq2UbTjKSKkbpaDE5Bxd1UH9VcxzxpEX7
hlJ3mCVVmKeR0LOkKTNQs0biz4g9ECIQpteTZ2vqeEQL5uCxwCt7u0ZyF8nDjp5y6XvKNmATr4HK
ybPOQ7kv3nnV9D3FbZeGSk1tj8KsUfR2x2nQ62S43Ktm4SLQl3NBTyV887Yn/ur/RxpsvqUuK0LO
wVsZTvgXiJqNabYWIeBFoBN5GuqmnsEdtV67owmJOF8XaB9pZ//inMjQIMlNwrWcloQGTdv06PxY
typrMPT373BZXlwM1w5mQ+F7RnMBUWkccjVVYWRmP1+9jGtiN4Nu/kgeE8LSo49uwyMditbSmcUd
7ZaqIQRdwbYmhBwConcQo5j5kqKqKRj+pyKaTtvJyJ8raJTpekUnTcHd47PN+OPYsdYIHHCGJWvM
f6rmuWErR3kW3PQqntlg4loCxEZUJhMGS0TCeFtzNEDAXVpy14ahJPDaRYYaSoBL5i8c3GDk3uxu
cr+93kQ+l1oDT0oE/e+hAKsZiMqaydIphG/4qxLiJ/n5Xwe+ICTM9A+R6OwpE1e7Jjqcrn6nE7Iz
uwHsPVOB/+N4dVzmQuws8VfGEM7ySmJ3U2fCT84tYnAZxnMTd3+rEXhWPHexTvk2OtEE3HTt1eYI
ETDg6JqPg1eSR5uIZeXtj7XJiebZVv3d5jJAlAI8DQJaMyolzOJToupzsjim72FfnA3tpKLyrgzX
CqXSGT1WGcBOsBarWci1CtQAeOT0LrMLHf2wNCWjqnKRMIm1ty2M5uZxl8g08LMUGc6T3wIJfp92
T0qViYLqCz23KdxPD2QKzD47gQ9mcoMoRPvE0yYR8wgFGrWOKVNMdeI7tBr6na26QKksO8FmwJg0
vd70T0k7fU+4zdudhuWkkgyPOKDEfP8kYlsLJUKqynd7MVCfYUKOn/xs3NVVeBIx5STP1poxyh+l
2vvfVue7HrEF7K79xFMKrOu5/+6FmXdlCCsEP/g2F/INg0FC01ay3kvxRbM1Rs5G5lvsl1ur8sSG
gm40ok1y90IsdXJBUr4h68VT81Jt6YL+LJgX+ZGJ2VkGcIXCFJuFwlLAOirNarO4d83HfTjd01hU
LIGublVwMvzNO+0YhGI+lynqQaiyMuxWx+pIBz4I6Ez5ycqUoNv2hdr05Yux3DeKhjA+6HydEbgU
RIDgJ3alF9G+5Am5b6qX3oyk66aoEQ+OOBYd00NT/jy3OTq5OdajsAkrwpMiNtxGmc/+s+BFnNHq
wz743wh8L4TcgHmN1nKHLqwwtI7/YdOYNYGLy5ZlIIsdHpHhCBks/YVdUtexNv/lyOvXY1MuuCCN
xWD5TRlfu695IC3d1M/4d5MtliCZ9j3LxzWH4rtd8DWNwk7egl495OrftrpUXiw16BKGf+Su6RQE
Ms83t5QDhIa4nLH/Vq+eUykYLp8LUBCYZreA+mh44Qd4MYl76F2zqnH2Q9z9YvGbCVZ4O7MTnM5l
htNr2Ro6OEb970g8S3mKfXfuMG9jagVYi/ltzb0aMKycq4QA8SmhLq+ph2vScbq9v9ttqFTQrDaJ
F3OZA+PIAalYBj+8BLq63Ht0a0umV2RUtPv8XmFgHebs1Rkly4HOxaQ6Iv7IGy9QMaT6mJu4Buiu
uWvrBjPHo9RZriDPA1ST6cp6yE0smqS0FoyxHrmYKKybj/0YXDkxSJZDj8XDlCbE3VayhA5sGdwJ
qRf5qlJBsqwAgP7TgXUKq1kI/r8ENj2ZYe4LI6qW7rIkZCNlUce19VUukSHItnGAH5h6rbhehY+S
oHKEWHexLs+DaBOjm/J5uvK3UL03Pm1N+1QriiSnmSiNK7crGU9UAFfnT4pSNUm5Y5AMKu6oygrT
zT2c5u5eOd3dcvSl61/n7yriVym3HRh0edZtXL7L/iot8EpMmzPdlXb+IGxSy9Wf//6PsR2SVBAG
co6nV2H78+Ca0llvnyPJs30xkbKA+UHKLAIqkONosxi6sC6Hv12fhOt+KQwItTag9mpwt2JUuwXL
+20izBh7Np3HH0LMkLaAjAQu4flkDtro/yoyws1f06aoIX1L8kzhA3ciIHat8yCPXMy3HCQToxTX
yIDNss+lo+fhthylKYznenDTBnaZwAMQDoE5sDl03cZqmQMPRg+wxoP6+xl/ErYtKyAe1TeEs1CA
txOc+s4OX5pvLgrtug3bQtI2gbBZiaGnLysUAQeMBupliLDHxTaSLjZaF4oyKCcL0zAaKFo3wzm5
oub5yFCgY3FcitO+ypR+1GDcoMR2VU9gtBzU87Co2i42y/xJo8abQnzwHrhm1TzU5rFwSt472Vsu
kC3zusg8MjxavqZ4hzEGsH1sLt09wIlOoiXQrrRnpXEf5rrW5bBWEhbZH7UyIFyPXCxpfLkJDGlK
srKE4bbkd2xHkLLkSXZ4EOO+XnHiNDbz0p0fGmcJ0yMM0SkJmW7RLq/YU3tzDYiKQMaJzT1+j0kh
6E9s2nG63zT1l2R5cUNQP9+whxxVa33JwtKCWQ7wkRAnbmoN3nFFh7lRqHx87OTNqUMluvHjIyMD
kgnmLt5DO4aKJQxBGN8Wk1NNZHgUHIXOmYXx20TGuziHGJeim1V+lD1TpI27974l5wnMCy/B1GyJ
4CaWjo1p0LaypwtwVrJ1uVglvX9W+KdfQRx4nvUWdmvGt+M0yLpvle50m927XEt7n3EyruWRkcIH
IdUyEfnCiSiJfXbW/vn46y8EH+TUzKV4k0E+Y+RGCo/b0i9DfPUaVlNIeHgn98/7ONR9suifRGvX
FhdU+dtf6D37BdF0UmSPuH62VB1qvgjVgG7HVmg9hmWssZnLY3w3mKPDtmMwOo8RfYGJTZ+y+QpS
yMslsJ5HkjXIC2jgWS46OVBhbpzbHAB03jUj2TaWdHo/8W/q96+okaQFvuRZgr5hwL0JooIyTHMa
poECVpYLeQaMLiIYtjv3vfBlGNShN8Iy+kBDLgngegJjwttDyirWOFJMxJvOdKea2tqk5Kfu7XeH
CTR3a/2HtoZH8jX+AvVx2eZ/AjNgRRFuaw3Bm0+4lVws7dm/BYAnJKU/SjK4MzMtNs1HC5iqT3De
yTQLhkw6b3nMJUZ3CUJvT684eTT/VZc6dHWX5THF/80c4rBUd85JWYoFQdX8KmK4bN8DWm/NEleb
gnpIZ+944KCp5wNeeCBLCjJTzmsrSsEZeWLuhcYhazDE1Msj0sW3n/Ncq9s2grtR4Ay/rmuxlVGF
Op25Kl4O5w0e9Qxl7lUWoy+MZ5M0oG+zlX0qAXiuLkDaN2iPC7x/Q2vEghxp8hN07yMeTJ9gofSx
g7vqke8BrnL/49fm2MQp9Xx4JoDT2jgCgjPTaMOAJ3rP8Dx+7emCPA2PJjywulkO6OYZUwGIG+k0
jL+lI3PE4Yv/gXgidz5938PsdQ0k1IKg1IaGBI/X8/dcM7vqvJvP+Sjd8HaqEPNCnETHg+6f2WoO
2sqmL+DtFhew9J276HmX99YAVhlFWxhitcUYZV2hFk/z3SpdURxfzDT4ZhvukUCJA6sLDD+SkXVt
RNqHMJ0cOFREGCG8So1e1mqwkzDI4pLVEU4XIK0+/1asmKGP7ZubhEM3iX9elh4LipfBgbi+FDZw
n9cABHkURkAWrQx14uctI7fmEqiJvT1+KqOOZrRIMGmLT6qyrAQNQ2WWLUxns2B4KHAmsIFdQbUr
Za9eKOOqJTSOFKicuHStokNZZuaLg2bjT1IfVIgTj3Tv3QZbG9j/3DbPGTW1HZh5iEZ6YipeYdfu
GOCHtmF6lcA7IoY0Txxya6jVLIGdbNfhmtxi52iNgy2m3GkekooPkiRMAPbpqli/3JoanI45hlrw
LkSrF1ZePbxSgqKkXCzOztrZ0qHuFEKKxBlzS5NkIfj36dnguYiyTpTjPfYMczwh/+i7mI3mQV71
PDiYI7aUhJLCyPbB0jQBI2M2PcudvpPa3jWkdQgo24Mc4KsZveJojWohAywR9Fh1axCDU3YOXz1t
xGVNCVGLGTJdRdfmhRmnMpVWdXFsZG4eqgac/Fjty1jvNHfrbX/zhKtg7jOYlVYiOfhurtLeM4HX
Ip34+g13lhjtFbj1bROw8RGx6jausNX8blpPHtoS0txgrVKzEPy7rjCHCkUm5O7cApRDn9uiYyuC
0tp+bwI0nGWadjUGtU/gOUT4R04KyDWjTDglzCj1it/WLC5BDVc6vy2lHrML6GQacg+OQzhn01gF
Jol1xKaDDBz0VVussMRBZ7PAACVUXoUelRgWnEuWmzr8deZy/tSY2NT9bujMOjPYsCBInBZqkEgn
CbZJSNiqesWU3f0GCGF2p1442nUwDZAIfj9v7R3dD37h3/QBE96muCi24DJA76ooIG5IlOkcDZaH
liEC/EdvMlWY5mMmMt5ljjoXlbE60yNTphyaBjdtSpjqDdBThxwnrlIlgVj67Izd7v4dpULvo1nF
OBXtYWDvdsGmvHkDnIaewNA6duMUvG6BOz2mR2iemNdgoV4Tj12EKtKqphW1e71RPkxTT82XAIbP
hTPmUm3NSOztO0uZ397C1veWLV8DGbJiVdnCiDOG7rw7ZzNHdZh/zN5TKUgfi9QT6eEJqyWullXP
YTKx0bFwomxNL6UOm4SoIEnAxIXmFnphudcNqHe2Ou9lCOI401CUVCdKmlWB4CsQI9V2XvK09aKa
/edh47SdgQUGluWthUu2NmIHGAYzdB5sx5s3rWgCROdr+LpOWngS4JVybEZlNvZEmzpzuER2th+a
2s3vngKxld/E/il6kLr26gsNupOq72p6/aFNzcjRjHlEcFwpikKJGIJ7sttK5zibGSolIzx8wU3q
64VracZByLLVN+AHvnIYixPsA5vzxAaJPfCprUdTA+lckFvt/Fvwsa+jIwNaFYCeRP7AlobiI7bB
Pbh2XLvB9yLbzxo00mtnZzVIRG2hzZTn/g6bZTxyUsMUGxIkjlb8PhQIxuC2TPAozk/cIN4eGLH4
010YmwPZSORghXV7+oi2t5iclXuAUSFiXBUX+jdZeKsSZa78k67hiufKpARUOOwbwkGPAJanvQEC
mD/JbJKRorvQswUXo5qqpy6Ua8n7WPSQNbcgeyP0l7oAoxeqLTeTonGLdPj6E0lc2zDXtV+I5AqY
rDcOP7Gx5CeZPjnlvrAtmx9Finp4twy0RxFmqgi/svYHn9FB5umBrI8bL6xrl6JXzeIzLBo7POw3
RccjgZOizFT3DJb8TMk0lgAlIsYaobb11nf2fJaz/ARSTD315yBw/HuUTvNCo4ykW6p4+cNqZng/
Eroe/afcGkEfaZVHU2FMrCTLggn+mqlgs/Y01VpsI8ReXSiqHtjtTFj+zKhDfTk+SZnwUUQjH6Ax
vc4fKd08DApWoBuyE+Tfh9DFjLRMOguzEaI0ZrshDGMbhhOn9QRd+e6vahWy5/3Tcjt7z4XBJ6aI
iV25e7xpu3Vd52A3E4vf3X11CsXk1xkpdvKIW1BMtT8DimbydzkG6qKrGe5GGhx52M0nZeko0SZq
W5+v2Dlu574Tm0Buw3H0d1hiS0FD0W85tA4u5YnTU9paTcZ6OXctBxEBvWCiE/nE8YNw83ilioWY
gM2PdUzzZdrrtKPVDa4RrzAQe1gHX48XGuPk8t91UNdD6rNERvu+4No/Sy9ZUPmW9tAdpDOaX4tr
CiZs1rK62XwsB3OqJt6Fctiyuc0i6cpd3VC8MmBGHfY8tXgnT7fTlZZ2PlewlgVlad9h4U//GW/a
v+YMpI2N3xMw7KvxEFJUeFOHaV/HSSR9mKg0vtHoNlNN3ZHpnF1GZK18aFgylcRE1j0GHIQyvVmZ
tOG7G5/PeFpOObM6yWOw6G3CRNpaY10H1C8YwM4+5RedLmYYy069uNAiO5OGzjFZCIwzDUKDEYk3
+DQJL8cKeo85ho7NT1CcVfYv1wTDdCjAG8i9tPi4QNDRvYMeCvbd1eChvwIclPGJd1HYHwqZ2Lkw
j1JllCxYzcQ1b5eHZbqtl7Dc0GbdHU9Iq+GVBZ4WuyYJ1z8XA9sZArcjTNpo3kJMIUexD6J5e/Ul
n50zfudDHWIsg4iXSiXUQxbnGps/fm4PfNo29Lk+Gj4aBAGWT47/YefxU+y16fvH72iHzgMQHZ0W
QpCkaZ4kvYuXRC8pilJNB/96enXSZ72Mwf+FQt47l7fElz+//Hobruf5xmjyg5rJYvNUsEZ7OnwM
e08dWCZQmBm6d7cxDh/M7MgX/8EPFt9LUA7nHKgTR34mTCaZPgECCYXsaxTal445oJjVY68SCdRY
r2hO0n6bFFw0hO+uKHe1w9dcg5OnrZv0/9KNBSxDG8vuPwS5OgmGAkxrqrGYeiBiRLWDtvWMEsDC
W9wSG2zfSy296P/fs4KeCun9rpiIilxu8SfUy4X0FOfJAXoaKUYvnQ7glUJ9wXQx2NmN4sLH9nJd
Z3YCMrZQqTH7jCUToyKbbFeIfoLHjWu0uQ4D1/x+fgdrnntedEUAIf83lcGEavOiMyBPYwKV6ssI
D9PI6c+RlwcCh5Hqhh5CnOtL2YX0BcfbtgE5ftUN9qaX/uYKg6295OW/vnnD9shm7tQp83UJdhLr
N0nzEwW2KvZqMzMVoOTB6C9e/n8iN2XtPFN3R44/GlmzWxDktEKBCdZcPjN5nPOsxO+9hy9498N8
aM2umAFlcgt9ZO38J2KuBIph0am2Ip+KaGc+KCL2CwtV9xR0KUZyuRnf71Z4pZhT0Z94qSozSEJ+
oV940FZDXKIeGcA08GgXc42J7MjsfvpW8tusnTbstmYBiGC19ukejFBpJC1AHdnvpyjeNGK7ZAU2
Z8Q2fdAE+DbfqR92qxpKzUyU/eP7hpHa36z3Xs3FAnbqwN50keu/oNvdRlJg27xv4F1PM8sH73M6
8ISIreSnuDVYMmRFftnJat+tu2CYXXmA6eVCSl5YzInvmExy4vcxWAp/lxvjW1S/J/gWB74pPos7
lnaX680o7V82juFdsnfXkX+P4Ki97ihKcsdtc+JP81NcLc7GSuZKnir4Zpnx5ocFRJzGsM5hihB/
OFqUqRE6nxLyo6cAjH8gidRikFtG3D8FPOijli3bN5Yu6mBzDQvIMgxyQrClgTPMJXi2uWnIjhnI
br79FP7phXtZBFl2ljfZSjjJtEin8HaBY89YtxETnk0kxheMfNooXLEGvfFvpmQ1Xq4UsRt1YI/o
qA0j0rKDVT7fKWN39pqS8cPbCfZ1fw2H2ZD08bj7lbT/yPHYGvAV547pZBkmpqwfnrIIHPCzJytn
T1NkXXMWf2TbQdQ4QqPQD9M4WxLyTWzYfEFBNS3vCnCZWQZ2e2gfEPSgQMIlNRTQYLtdpOu9l/X+
88WvNglflAgn+7uma+eTlFqp+Ey6SqPZlUUUz1IWpVmJrH0Yfzoquhp1UE1bftTKfBWOyRjCQudQ
6RLpveehL5ui9j5S6XXmKPcQtNmheRAxITHi2LgyVzDOUSOkBZPBGYfmm2LPbkWui9wAY1UcqkeV
2tTK85GJMj5LnQof0Su/ULUOqbfdDGFlbzkvlxgcbBxOHZbt4NGfizQGv05EbouCdwk2xBFVgXTw
a2cDDw8DM5BuWvasQz+evhaemn8m7lH6FHKEzGsQbHwQoAmEOvusYlhoQ57q3RvWksDeQG7rd+j5
bKIwPNTzvqAr7ZEC3AG+N2S3lPYEmwtT/q3IuZSTy0ysqE3L7uKHFeb7AZ+ArMrVwEEQTXNmdffT
qdqu/dGwVXVg+5qZtMY6VAOlgieEqFjMvvlrN05gvusSDxptXqzBcTGp4518YDxdqOde314XOgvq
kckHZSSx3QCIpaGlAkarRdr5qDe3tkbsNYVOWLhlukuafywcZAYXRG1U820hARTU303Zj1e6GFVV
vBXcgjUuEhpQhbkBnFaINi0+CC4DFrC9xe9T3aU+l8ynueV8xNRqufZ9ajuK96xhXBzcqWbKZXH3
8Ibk7wjsf9Dp91/Bby+Jgup/NfPYwIEWYBHwxb90w2xVQIE8JBYUtFVyti8clLQAv1ROrdJsD6Ir
NG/nOOcml1O/ONft6ULTgoKXCnh7Cen4yMBNxdQ/GWKzZ4iAGJw7vEvmkvDDZx2d+GXDXpR2i/Vc
XXJFJUoFqlwTYQ8N/kiaQa0CZDaB8w85+zxZgSxcIrX2re8kEwsY484v0MmjgYpnjJnS7qgwSxaT
RL4uvbC7C37EO5ilEWiHa1dSdYPnVTbYAiKITASg/ytixQFFZixbEEdq0AfCZwUvJNnZP1LEuqtO
azNUHjjoUCIa18qkdfWR1u6pcZ831HcIEiUVUj6EUpjxGz1vpnBt/MZY+6rxuK9j55vZewK0lz/k
b+0x6x4+gCfkUFFUdqoyckV+dvV1sfs76n8ClRuO18Uh1oncjDiHUCK5C+zw37US5QT/o6k7xI17
G3xFd9eWy2ACScNLL4NkhUVqI5SoVhJ7D4UQw9Z+GHzmLvtNhdf7ZyhUdnXcqq0yUfONfl7Yg1qh
TRH1R4Z0nDjYkmNGj4x+Gk5K492Zh0lhmKV8RGXQGrZpRJbK/vSCmdqX8Nk0kcr7cdgi4h88b3GZ
PiOsA/XX+rJTBwVW6yIkIl2LB2OVrlk+m6Xz6uitBzDPHTqWoT2vDZ8QHt7T769h8jFvqVhILIYT
yJASh6mo+UApN8yIR0hMaZQFL8KJqdgPJDGlTwFDcSosBLXPmPwRrXidUbYKh4XuCiTsYcMLVxii
Wky6DoHfN673y/j28BIQvWD3/QWaHN+O3xwRU7MqFkhYT/wpE7jL23Ujm82poLKjRcIqB423dSdO
t9i3eHxyCAzyT7kRRUdL7XXoJoj/HQRftlI9lEqERlr5zAbqIQ4Gyqsf9Uy5L+anWDKavw9zGO8P
xWaDS4MyLV4rQLjF/v0wBX6DhA0yrdGZHXZ+52a3jptCGXucotvWA0za8w+Ie3A9CwXPQ7Qc9ZDI
vHDzNGPRTlS4rtIEXKcTlXcKyR7bSvRrJMZHKq1vx7baX1toqi1/Z8tQD27fNRHiHYw4xDlvzV9K
M+5aiBdbrdthQP7C/7qON9AA36CzbnQ8yMhZTFrr7kFI5B3b89+RZlP43jJUlvAjmQH+FzBjJjON
aiucC6h+s4JggM/oRGWVuWOLwioq11GBi2iOiI8MidQShPw6hOGUmti7QGLjf6eJUbvClRh8pykQ
HFEjgnpuYi0ju5LjcasaEySgN+IZkXN/XAGp+T3PqB2hpHD99176dbEFnSuNoqr5zdP1q34Imki/
XtamNgLnq7uWaDWT/bEsShYF/BQlJwSMkUcW8ORwO7l3zPBHKEhUvjebZV9CdJyTXsfTxUD46Tzt
SaDDkhsprqX56ez5c6jrwEyJtCM/vJprQ1hMmIX3s0AK2HqXkGKb+bOMz4dYzBZL1kWJGi1WW0iK
ZvUtfoaUQkwPKvOBCQNWIsnLOqbknt6wDLy96AEx5Ygi1HhDBk+V7KsUgT6T31lxCvkWKs8Dqyol
6qkkRG+uFpBrV/XWjD8TyrCvRokm02Uj38L/sU/u485GarNcrsyrw0jMlE+kwBjZfDhraPk7BW8+
W2nucE/DloAtMvnAlfeVkMC8d14+ptL5uqFDyeYUYLTdzDpg7Xp1M3K2YpX5PZ+Iiyt5CUwkM1ya
1abw6WcmiEQyIDYjyqSpIG0TXgVMxn7MWcpLYVuco+pe1HXo+cbQmTQQByGwa+3W//zH42FbOwE4
YG/BeAS7cwqPooAxjYkExtubiKlCo7ys7onGwUkV5RpxQUqwieCzPeczpjquYRbnJzV+tGNqWKU3
VMuO9dJeH1W04DMbTAcyxHm4AkZCEZaaCyZ000gc2LaCAyYjyIJ/2gxHnAqSgSdu85dGgnn/fQ8+
NwEPYRBLXcPiTevRjcUuW+PhM4XUBItZchAD+RIij329epx5Ri6S1Gvzg+UNqHBgMGTdz88T6PwA
K00Wo3K0In5glhqFz8HnlaWcepwMKLdCw3cICT4YqYbsLLmRfG57W40bXWQo64YpCqTkWzzUypSY
OJBWKj7zsl++JV+G4d2VkqRjigBiGchL/yijwx+ItMoWTjrZZWKsf/+dSjcIWYb4iIAhUQAlZasv
SPmd+MY/eQpYRg6ACxjt1EeK1vfWAk2NIqxMauk+8zWf1+4WhWrIFO6hBYyJSOTxzBOpR7GF9JAz
0dbNxWtm6tP3V7x4z+vCGaIXtjTFMhG1RGymp0ytUa0YLE3qo0ee/TIOkU1f8PAryarmPgBpNVhY
lEcb33EJLMOkbo4Xy4MtxaGwa4DSfo40iiBDaAtJ3fA4X1tFBiaNaDffO0JX1CHGMto9b01dEKNO
5FYEIn0PbB6hexNQy1Vto8ZbmyybaFaweHNVvY6bHUb0F/U1ABVvBfeuhAorrhU/MTyVyROMNMWg
pGSEKIE47jpZeba1j94GkmYbTCA5517HD+RTkrRXpcXt3auGKswFMuf1TubyGBIXE/US7FkIfAwx
4lL+P17x9R8KwsEXEB28lImS6uH1SadfgW0NUeb1Z87J7l8MZBQ83CB/2bZXdkLMtuHJn/66SM9d
7Lze0rJi1V5v41wzgH6SCXHssFpd3eJp/ApoI+9o7S03pqHAMok0dPNhUHHqScKxJkkN3v8vJjgf
MmjL0KNnw7nGuylNJlsElTmUjV+woCi1Ab+i6M58HysTChYcI07oM/ovhvu7OIeAKkrgGuRcG91Y
YFLmz6QlqyGiNgTK33TzHU0F3cLdW3ttWzDub0lYczZ1cW5mUhQDkhoMbitUgroRU3cBf8/nW1S9
CPC0j+GwMUpzW2nfaNP2nnQgNGgfbdDy0EhrhNE4Qg1gedeh2xDb1S6T+ElMATvzelwMrIKbM/QB
hKRJqnfzlpoBYmqBS2yShSdMlpxKHesQOXG1LbLJvaXMMfQL1Wq0XMQO39n7PrK7iVmBzKQZe5a2
HGbzLak3ZaBDUjdJ0IP/GptwFDxhKFF1wHZ0RqAgjnkWNwoo8/p10VTx1oJY8H5juiO3g+gYq8Ze
eXWO91c2RipBN46GYypRt3LE3hnbgCbv9Zto178zU16pJ0y/4w62OvOFWbXGGXjAoJdtTVE1nKMZ
0+MkG1SDhYjGxY+MiF7QWLP9NAFzawK9UumSvtJdkoXV9Kevb1IkIkhTJvQv1BXC7RA+GVVvHf2c
T/cN48a5/p0RcoqfLeZ5jpzvlzAJdHrakNwduQsFuL1Sib5UW/bUJkXgeW87hMMad8gbYroC7Gu3
tHaVFK4JyyxmFKsvlC1sJyX82y351iH/j1ZiWDxHEdp61qttz6zizb+6MoazALbY2N2c0VEnF7Sm
jnXjumsymwimktXt0L4rIwE/zSXvdU3xjvNwy19kDkTlHQUzmDoXJhhCNpuaQm+SASjirFtD/uGM
TCLpwvtJu10xccitNJxYdRprJW4I4vKCkZbgt2Sejod/uqI3S0ViaIxEnvKZvYS7ON48Dx5YpPhC
BkWZSujArWtUmiagmeMaLhPYXlW/TVzwM44l9/qOiZqDNSxAbC+m2stEujfAsUIh0CAvANaNndgf
ehw4Dviw28qYrU04nfuyfKa7sX8xC4GB1dgF0hMqfuGB+On7gNSm3gkzVxiq50NRlSWJRFXV3cRT
JEsY1QuzI3yC1u+WSrdX2zKA7rOUqhThzuPsfLUZL/Bzhap3hGf1lI55AhgjhE9fz2ro7fUc9Fmn
K/UssYsRDAYuW1tlEbxEvfZD1W5quP8MCYS4Bj5p7OQCqHYsMMJfkYn+nUSzLg2T7CcCbAeZ4Yyt
c+08uIqaAIhJ7uPlMxK6KfytjEvCgvhf/eCM1+m6MIDwzOlvIyZgJmV/ZpjuuX3BSZ8tVcQUIcwJ
CiykY1a358UuXHum4/qjejhFEFRogHikDrczlaCxVj53lu8E/AUhTxbx4zFs6t4K9POm8ls4bhZk
nV9Wm4mqFoVm6M5XMPUoPX/OldffB3DSonj5Uvi3jKO3jyqQRe416GrEHU9iShQQTXbfUJFcYqln
p9BSYtSRj8n+uU/AFdlmrqHdzKmARrXzlFdcx131OAQFLB2y75oJRhAGPORo0iSJnzktCcrJ6vzZ
ifBZxaZ31Lapi56B04B7NSjZGc8kvyVViwsUIh56e3qyeWc7dg9wm2Fy8sd2axvqZFRMJCKEjGHb
4dIU/DEJrYc/h1p0f+oZj9es4SS6tSGnQedN9wGkitB8eI336QE4bc8lf719xsriry1ekoTY6rTo
zu3flHg6l8t7FvqVn01/jpe5ICZpux3lRWp0cSRKyvOVn1L3zvoAB1HvhGLs6u+st7zwOazwyeDD
JrYXyM/payZo3lCbRptAThY9EVVb8h6ohP0WovJ4qwD2H0h4XQV0WYeIRdfUE5MxRIDl2DEsN02e
pSHeRbjYTQm6N94g81Z5edi7wKBgHPQoYuco+cPPF4jJfnHOghagkZXCXt8O6ac3+66S8a2RLVFS
wjolc8wC7ch0qSDBOBTWxdVd0z27p6bciGtUGr9eDwpndkvH3UQZHHYARaIlZAl9nvHde5Z/khBI
mLn/5ymSwctlRNbs5Sl+TB3+TRrbTBmh9tCVdHckhMyW0qvDftAusgGa3zgEUFVVvhH/jwWNLEhV
TgtuXOTUqP7BaAIwHi1LgP1bGuwPiOx6gpxdn2ImOPQHiiBXpNoDcQRnlCpQehJ/4dIZRy2Fl9cW
r8KLu05e6Yqig34Rudt5kriA0+J9dOwmyj75zqmNLPMkwpzJ/3lRFUUEdioY4PU8hC9Gjlj/A3mB
D8NmZRS8O5jx4jhtNF7Qh7HuBmiG7vEXKnXrHO6gxYFZHEjW8P7NelXUk3JcRu6olMyu5bVyfzJ0
USC+CKbA4i4GF9H0FndJdvqm24441ob6Nte9sdKX9aRRTfxH5ZeKF3Dcn1e592kdRTQsgWv7ZZ0N
6ctwGF0FMRaqkrzTvJ7ldH8D2ivEDbBKig5saJBHvAr6Dun5A6a0X4AzSv59T5dhRJ8JsA3Q3D65
f9VAmQD/9xsQbtfDwRpxEBWL4GSWz6nXhsFZ47Wpy/Nf+PTX0zQKt+/llwyu6meIdodnVb4LPty5
sV2yv3FrHzee3lxwF/wAu+4fcO7BuLZ+YggecMYtZWJlJbhtdPAvwltf7Szdpj9V+OVWWIYeABBs
A2T6vWSVbdAElv/BBLSTrUOyGWpCiO342N7JVtzVPLI4qhEAjnTmsVKkbEbf+pEbn0aPgsUHcVMi
lbHRi1wS9KTOCEtLhgZRozeP3KJZFoA+1fJUY1uLgj84ISRm3PqpvDTrvGVfHFs3jXvwDC70HWjG
xTjAkqSHLHjh6UfWYE01wnlYEbYlBzpijLlZFeeghXORJKAp+ZOlnycCsznazmkdT6t6cQV3kvMO
DznfL0BRBUa2fMS4Gbm/2zCv5+w66pjo/Xjikvb/AsEVpXpJXgHeKe6xlk3piPCuZnQ2gdNRUB1o
Wwiq66l6+yglgXL1w86nzgUl/DE6sbnqIAf7WCh5YBLM9G4z0grdf7tXxLBxucjH2UtRNZTeD2p5
qEYY8/920Vz5TICf+yXya/tduUVRnaR5zyn7UE6to4zfjKBisnO13Ps6FhRrDTQlMNSD26bJNXmC
ZptGzrcr15fYEzPCd4Wk7RIiANXkpa081F2R+y+9lMi7LrJywqucmaUuH4iQRG9raxs3oDFWqzsr
Xh0l6AhQ6780YdLDXjpK5qEcmwPs+0Y7HYkWpaMIWWXE6K8IzGy6bf/pYRmpKIuBkVAsgbpXjFcP
gnbebGPphzlZa1sNyb94uiewiyBuYspOh4TQnqPgOAfq395jiolzsEPuIJNyEc8+NmOrVp8RXem2
EuEAmVStupsUVdzo0nzGRJ6GeWl3qFSA4F0Wj7XObYM0FsgNr4LMGqRKjUNFbG3183wAmAt2Xxby
117xdeItR6f66UQreVYxACK6EW1G9h1o7BVyISq8OlcI9hpkAwqGGhPSzP9wi73pU6RqDyhu9ajE
yZoc14nUs8WKGYNdJ6Paxs1/1IpPg+NqmFPHgp1T1hdOw/hgKXAX0WRqF2GuxtrwdVXp76p7IhgW
Yr6CKzBPRNtmcCt2dZfF0SVrSNkWvXGQngA+TwGoVwEQmAPcxfUMp+DbZCQvM314writ4c+GqhfD
AWcM++8C/CZVBuvpvHPgNqQIxKx+yGEq3AB8AIY67Wdp2/bLNddlp+orPBmWRfdPv0i0m3B4t3/S
pQGJKXxPxWy0seUyHMUvciKS6TLTclf/GmzOYC5mUVE9N5SDwdMGGIEUP286vPYrJcYzoOqxCKqb
fGUz0jccIt+CQ9l/kf/EW8zOG6rTRJ4GcUHM5r1/LYY7sPx9R/KAqTuMXxbHDHlH53GYixBYG/EI
2EqhA32L9xU9ikMfKLeIzmHyNlgqQpd50JWf0qWBsACSxUYKanXdx09wrp0I0aRbUCSBUBdNTnHS
OPRwWnArMbZA4GNbn3BsUhHgap5phLfRHQcqd3zmVEicB7CnvECMQURiT5RFmFz5TKjBPVmzhe40
X7pCyPZ5BmNfvtQXyvauZ1iso/MH+ar9LM/i/Vg86ZRtbKzPGpuShQGe3OFEdHEdMdDZm830iWkE
ajhHG1ygSuBMWL3jAyGR126wQVZbFbGez8/iiwnOnpS2iPHNGbbKaqLGPtTX4miRPiCYQG6lL6lE
xm8Q6DJc30crjkj7GLbuzbY+aYoE3hjZ8u3oCj4OJjUUHmI6mnjSSv7oHkQ4Q6ri7rVos5suCBJ6
AbaW23/FY09PB7AG2mh5FB/OWngCZ0vUJEw/BNg0OHe/iJjs96TniH7eny+ooDa/R7EvPzu++B3/
D+BcBZwXAZoOdyi4w7zabhAPL6kzA9kMZ3NtjX4fySf5MSYQPUF20MOB8jqME705ufiQkZdb2hhT
aKbI78OmCe1alxDtch7k5PrS1l5PR8/eT/DGDtIynzgjp/bql7ioOLtf1+EpsjQ/coRjXquPKOzy
S1Pa/NS1vVBHTkvIv9K6yp2rZs+kjWeuzzLWsgQZDVIo3RwSuRdi7rXTVTBR2dIcis6ZVa9vSz8M
OlMIbwmMnZOi0Cv+yCwcFwkAB1bAe30RDi9CeOmd9uIhhj8Nawopc5yhlHG0HifU5BUhSupvy3mm
h+U/ilObzStfvRhycT/dlFH80pDYqln15CVYwrE/jA5N7kkwNI6g+IGjSpBnxO8uLWQ3OE+AMbPT
YqdSX1lgmTDmDV61ZRRn2EHkgpkGS5lh4izlk4HjtyV6hihNPoQKyTv8Z5JsTzQHDTaeUN3tHbYC
5w1+YQw5Gy2noo3Q62pStNijpp8sHkXmFuqYTJ+zKyAjIlyMuc1n9hbrl/jvKC7bJzSPXUmYn/hD
Abps2X/x16yOmtrwX+y/b2zGW3GcT/VNHqNUnV24Rjz9lLX8MpUEYMMkwzZINB//Qb6cj+4Xzk55
RSdJF17v4DeZ9ABuLV+2ABlOk+T9xpePShvXEXQg8VHdyIrTe7JmR4fd3NiMQONG1hdDCI9dxGPt
IB3wNCvBnenuQ/Yt1pmXL/FvRElOXn3bRcBnCIpCgiZ/LuJA9rGSb7g5rEFpbslib3rn2uuxssmk
biJfJQ5HRK3s1UBYADJvP5ewCBSh0PZaDtMhb2CC90cneTG9SmiEG7n4NNXbSOOPLFROSZgGgJq1
4FE9wTIPNYgvMsPV2Z+c8y8NIyT7RZ232sjSCg/eXWaekWJWIwsmICUqxjK4wYSJwc1Q0s9zfMds
9i3a5WdtA2EzBjPRU0lJV2dyDKQvtQMpET3P88TO7WLwqVD4AqSM0n7DiHPy+h3qv7ZQYAx26BHw
JNvPlYthedSnPwPFugq7dpo62RzViSM+B9mZ+Y8kr0ZBCegsmOwjsjxwYiHLqWDVYeFkHqpnk5Hh
5OdJXA1Lf+lhiFoVT/1WBks3HyX1CPtM1K0EDLr2A07oT94Eilr1YE2HUgKni06xu71pVGFvjeif
QM5KOH9K0i1fnakKdpOrTuHO3FI1DkMgzv7OcJ97wovECb7RyyKbvc9ymo0bg9QFd1bi9/EoprmT
ZN/mxPkWyrPVsXyMi/P4x2HgRM53Ethr2C5j8BPOQL7w9x6rglM8PViRyP76iitsGwoUJsbkaBs6
K7dZ9DZeUqB4HJP8qAu9to2lrcmQgDQqBFaJuJWnskoz8qyJEQ61uMYN+BrpvmdomNNNRhjtV5rp
YEUAyYswFGCs81g9sAqLqaT8QTJdVC76ztwcSzvaMQ5lVjN20E21huGe3uPRnZ123jn7ZbFF3qmD
ycRfera5DpWgW1Y0eXus0zcT9oMNcKBqU3EJOaCO39V0qX9TTYmFUSwJjjhlhzTx4lqoh+f1qoDt
309rdZNJewlCtS0n1GhrQKs/awtDKLLpwWmt1b4nQVX3xXBC4srHhq/wLY44Rl/3CyS9+/f6AENX
TCDu6U7F3VrsSdiIJH2/+3F84jZF6HVyjpymUSBD13brb/wf4l3wM2STJWLAflrrt5m6InpMMRkr
eQCjYZwy8SsQgOOfq26GTvVymZI09lOYvhkzw0xyS0iuQv/6jL6J5i6IHIiPZnBgFQbITeYXSVup
rRxY/v4lkn9pdVcNUAdvl1hZyhG0TG1W96cOUW/SOWXMd8VBN5m/hW4Dm68OIBwrAli8AB475wsS
UyptM8kBWPyOn8OxB9+UjHghSCEO3W3VkCMq4lZKegaHHbJ3ludaMRN7OR3BFXPDaL1DhuQ9+211
KCFEvXZ1kY8jn0b/6l1OOvtFz6t4dZMa1h0SsqVvy48pq8F6dSQXrAEwjzf5XSJij5BimWtdFLXE
JNL+kLi7gEGSgDdOs92GzaCWoGqbqLOa/5l0OhopMxkIn2SKS12DetMIQ1qm/RW8ylubA37XxxnK
qhIeCR4rQYWKpuPsZtJMvqeQQNVaEfAzlyFmqmaEupNn6Y7V9gOSIV9+cWO84z3qX05ureuszXwX
dATZ3XXqrDotDIf9LyQ2izF5rIHV1Slal8nh+A5YVme2FP1T7ZVATfxApcAlHe8qIoQ7n8r7IU37
E7ZxxIqvSPTBrin5fH/lBvFxG2yhLFDETfeLcnaXrdruMwuzPwyBDbzsUIxhGqotJ21SOW99erTc
FSmYAOs4hUx7OqWJC09rlU9IX9Rayo7wDf5KiAMY9Xyuqj2Q+fheEFzrYnNuKVpihhQugHzaUKJg
ZNcQWdSgbiOsmfJ3e6+bb5ibR/pEIW/x1HeyJgtlpyiISPfBmPlsvrYcmsvyyR2efCe02KY8Mbaz
dVMdOd7Qbj/agybOdIw708gcLLpr8dJJteMfXv/648pbSWugXlWXT+YSrgVo0Tlv90NbB+MxeTbT
iU5Xyar1WyW3rgFnuKkNfsqAQs/DMYQM+rA88vhQtgf/AfloLsD+IhElUpAN0QjUrHJipmHqm6Fx
MnSPYGnsTs2k0zkSgYwtF8q/pN7iTBTL55FdtGfubwQ4LqjSuc8+TlAPzVPhp7Ir8oU8ume0bn25
x/nmZVzAbhOVX9cgmR9roIPNPGdQB52ypZatTAKlzkumOR5fU0qnza5xk869wedwgI4vKJjGCkzO
l9nLGzie1VAPh7XORAvX90VUIOgKMSJIkzToduM3juMR7NZiYRpeaRZbjUqmAzGYkToMazXk4Vca
9BqL05npIKIaZe0gvuVVgC2FqYeYbUi/sRYI+PSPJs7LReNHqUnlZIiUBXy2w3PSw8Cau4yHp7k6
ruWmLh7GJ7KT/RabSI7kszAWI+sG7MsBR6h6bEe4KbV6j1bb84eLBmoQgv644YFkhJF7o8iaaqIG
ZfKH7mletDxC8y8/FP919mB3NCapyQ7kQyhp/87Cdsw4siLYHYNXP6AYTGB4DlkfAtINxOjNNm/c
QBizUus/V/jTMMp+VWBK1WS+31Lh7SCLIK94FqqViGU3Yp07vb4GHvJMe3TPHHX+Lg5gdfbKiSMe
sHdhCsXjZJwVY2f90dJuuo+Ei7wUgUjljBx6PqRnxR8x/qL6+/YtytOEjBx3U/c9uN7IVeyOizZx
W68cc6euN9kpqt/9f60c2Xc+02ISjwlcrPLhtyOXRwt8Lb4t7hhA4uh2mFIxRqTfwAO6cDkUXZS6
H7W0FZNUbV7KX3uNJ/0VQkKTdtqMFGUSKjLoPQJeKD+PnxaoLFQreLSYLYAAMrtqIbMY+BhFd5iG
LekmVaNDGWgerlk6P8bMwezOwmOTWk15dF/SvixV9m5cwqKcyq+7IGTE0KxG6CFvw9uzAJR7me43
onI9GFmYdqkp5vRJ2vLT4sdfC5LkiJ5mzhTp2wc6V4MIC+TJx4cFi7b7qikRUMYtuxEBUVI5+oGz
8QXHaRRvEFpVlzCGmJVIuM8Nj4UKSLhmpL8SAuJ9eCrnk83HVvE6mXFVRhwfEOXWoz5ROm5ROX9r
p0x/k0fsUz95f5frWYNGNKvbCNYyyKVKW/JkbVeH06zotMJ7brjtA2jN+5L+f3ToMLWgCB3jALNw
aN0ekJ5szT5N5HT7GPLfgbzJ6fHaKTEfWi0IWmLzdhj2cs1Us/pRCcubacIkXWGkwwQdUbG3Ep+g
/uPvdYEnsZT82aPg6+Vav9CqEhDTDbNHkDUDgoAKWDmbB8wpieA00dN1dwuX9OypsJGYgLI8UwEU
x/KuBjt15MoA6VdwrkHtp9eV2Pgv2/Xx9aquL/PCpnJYwN6YOjiovQ+siNqmwN18UqdUa2QY7sQD
xH8LPj22qU0z2ArpY6Up4ryS69HZFkM6Cd6ptrCsIMSYvN97HXz1TurLfCGpyHzi3001VBAcR75N
jF/zmj/9mtuEaECvF9i8N8J4sDvVpT6dwVjV37nTopenYxuqAcsAaVEEhoJt/LuvhQ15N7Q3EM6r
YSF/DtwWwCQ9Pf5QgN5kJ/hroNImBSJ85krEp3JrjHl8mp7zWE+LFOwPg0S7mtaFAtS/PPLxK1tS
vjAyhkpQX6aRel1aOswVawK1mUCEMjuyBIjD7av86ynhwyENHfAXSwdYWjUPWqzemjfi8w/JGa8F
Q05XgB424Nybn8/eHxVgj5Uq+CLoVnXDm6QwZ9dexujPB/snhBU4HnURxei/EULHMny9jEZ57joR
ObN4y+I9OZZUw8kq4umf5fxCUe5DijTkPS17FzF5p7rcEC02aTSYyDwl8YgXBRIaxtnCQV0MEDZz
7k7oC0DgRLEy5I2eq5NxrVMAtkg51nGjLKfrf55kl5F+wyk8yWPKhQWTSmQx1c9RnjzY9SRDRbip
wgkt5OYH85P2BTIDj7prI5YD0sKi2YszIQt1H1rB7fckAr4B/o29fjrncUmkefinyrUmhkIQXWB1
BdiPyNZ9sbYfI379fSSOGhokb6b0cPN0zqlZ+FEQMV2K/ZQ8Lqp6d4q/KIp2xS0ZMtqVRTZTfwAS
armL9YGAM+UAjgFLv0/ErFXnxytmq5AH9gjDVVyROHilxWKWbKy58kKiXWFI5+OcDGm+IlhbmqRN
LJLBhobKePo74+9AO0FzUl7cxest6afXUc8dR5R3LhdNa1MnnTGwdVcMrvV74ycqIYwUV7LdTv7/
NSE3uCCkHT2ZYrsJekSMao/PQvtHcyn3pTslHsbYOvlnC27C5bW+TYRZ/kxYXeX9VaNA7ywTY74D
y31qQ3B6EDqY5FtT9kDfq+/0P6cKMjFn+wXFX5/vPYmjmOZwn8tn1rXoNGt5y+vE69SaPunX58qx
hs7aVSaMhIVs3R/UM3XAyxLWwiKufEHQfg3U5m6V8b5nT0P+toGHk1GoQJAT0g7cDCd5GwnnfoTz
9J6eOGARbvJvtQSJHjVnzhl59fB+aFMG2h3lBjXq1kQIx0iVbhT+91f3ULvSt09lY9nGgQa7FkKb
Sa7uNRKd2ndGCTmS2jeN5uUevNeWgcbiREzKKCMOKOrPhNr9NyqUAo3eTEs64cHBLB3yVtv2nNa3
znMO60K428oMWKOlOafU47Vy5Z8wzNGnwawDGXKEH38kR+Mhnqa4CKD7OJ9kdg5o2DQ6t2P0MdEL
fdhL3ZQSKX5tjQN6Rs4+JHzZju7hqF37PgFyfeSO/xsSzxN2+pS7Q39LDo9/Jukm7xLEuGMd6pIu
MzZVsXkXvdZIiHraRRyJakB71b9kSR8J5bMGjr+mlVCLwz7lP1MQeZFD0QAJx1k1BTbOnpm89EiH
g0tngWx/LOBpOA8z+Zn4XMdKbOUxSYqNeq0WhfBiz5O8mMMdqoHSF05Ekjgs1ASmzzsmrKCs/4wG
wcB1Ce+Yfo498eOnWP/+tmEStQg4fyMMSaNLBENX7ORx6HDXU+fqTgrdCeLSQE1rKS4AVu0BqVWi
WzApoT8db4dkI+e1532bUwiHIjgADMBsOVcTPc1jBee4pGlQVnxOi8wlT1gziMT52WHoT2GNILMb
snTZJm62tuIzYzZrRBF3GpoerOK5Pnip/naCkjtHC/D2bre2vuqgCPR+mVjPgsSTP2xJX+vCfYlk
0ZAY10mwLA3vZySRExOQMvXsJWUnCAPkhCCrL19nHXR77+UFuHdK+DUhuRhYCdf3TGelZcy6eNI5
7u9wkoieivu19AZNdn6mKWp1Dvfj0jtH7c0vKwZvC0YjRT4ybr2Fyw80Zxc2kpBWYkZ67WkmkImb
5un19NGx090PMWBQYUfuT0mY9xD3EXrwwmN/orDsvPEj+JHeAhJIsYojRFAnQCHRca4aS2g8LJgi
LnNqj5pPJBptNTkIpOOj02bSjQbJuE2/BL1UyzINCvTkR2uLUY+C2BsHDX6OkwRBQuvMDzH2TFsI
DjRWQPEvdMydS4mlb3FSveRb68n9SohsCb4xW1p/hAgIVkpY/ooOo99JRoKXLssnCMVBb3f0h3DM
iM8QQGLa5mKsIylcXHjcspKGqlieZEWeVfwPdDcIHOfGBSVAFknuxTEA2/UWDfPb0EQJ3AWkeghv
C1w/20w471m2FsNuOSiGjAZGl/3D2GqE1nYVAMIbcc8362dfaM3gS5rJ/ZP952fkoh8YVguH3AVo
v9UsTeNZAr3yj8wj8qjx7lkL8ZyFPbncYdPPzHnAxtHhhKzS6BUKd9nvXdJGy9pcsa45N3L/+a4j
PD8X6Xhh8dWuW6a/MoWTJJf2yB9rCZYbz+yM+z+yfJDHq3zGlNLRoMVADehKaeAmKH2EfLNB5m/W
f4zpZO+Hlv7iAAXnOb2AInCXZPQ6Blvffl8uEFgIszHyCtlKbQSdQpT9T1fReWdYPLCNRbD8NMPw
lkohZ9qrx7OFX5e+GKmC7tN9kU8ZqJrFfsgytrQvtzJtGh8dEwAz/a68nQB/VmjQud8xsDhEYmAw
fWzohpW7uGukbmlq1vO8uxRmhF/ykxHj9Rjl3r1DlXerfEkll+wOdgq0y85cJuBlLzgtslWr3vjP
kcXrHPbUK9jWkKENNgE9oaenfCE99/0utnGeUDONfjhK2ERrw5RQqaV9wuu9zKb9M9EAFzlAKqIy
QaWxXHeufOv/hkw5oC5hjiJBDvUwOuFNRRzeOP7SBQTyjSeU2K1RRNvmo3U1hVzQmrYxnFwb5v5m
yTrxUYd2MaGXZyt1ZOv/R6KiJVgl/xgDzihzA+HV6dzQFDpDo7OCe1CRueHiKvhKfnOw4KPcYBjD
lZWZRNmL9u+bZiP5+mR+gJzRdVV/h24iWiVzlpx1UXMlLvYUqM7J1xaFdzY4BSFn9oBQwetz4aHE
2I7oiQTTRH6rLWQhGi9OV+1poc6m8e1ySROqfQGsr+w7QTsw/nbPuvXuO/rv7HKstc5GP8QyNqBZ
uepLOKZmnqGOeMG5wdMlpXVsWkphpl3Dvaw8sYBMf1CaUIJlevd71/zWkTQwDVBIFkSB88ekwEju
csAvU+F+ix1BsL7Gg1OoW7bejMahMKEInXw4x52JcF+2ElnYbO4qsxJswq9YcOjA5ufm+qiLnzyc
3O4Bl39dgD2GoDa+P2L31g4gzbThppFweAPue+A1y7kAEM4RpBvYWceXxNoK/fnWFuPYyHFL7xhw
flEjnY2kVBpilrvssbOnodORI8ksxXgWDrGFS7GdTJGvtlitXhBWPN4w26KRthimFSrDEab49ylu
D9s4vTC19q4GASAkqloYfHaq+MDGfPrHZut6iKhDkFh2SvTTdF/MCwqvlVsAKJJxWVdzLt7133Nj
/f8py6fzNYP1YMax1uMzdEiq1ar5cPHlO6VsyizHSTCKZVqfvOh0Tz7NdurgCaxkWB2Q8fAkZ5hQ
OquHPiTu0i5M+e40YSh2qDf6RIVLqIisGjeGaKPprjF+ohugjRkrFZf+Z6Dp34jkSRKc2delSb7t
y+uYc7y1sMxO7gXUFsDoS3/k/N3XPUAOt8ryjMg6VWQ24vQoB0YkObE/Al8fvA+KO32a4ABepZyj
V9/ODJ+5yTDH1EB0J1HNn3o9xzv5PjIl7JHXCYaC0ybmdZKPQGmpJ9knnoExb6w0KPioCZpOQwGG
eO0Ho+t+KxOdEZ347RDg+ShtP/q4YxdP3dUYNhprVSsa7mMtLn4SwlNMDN7fMlKM/5wBOmmD48gi
oVCmzkfT99E0mQ6QjdU33ltwSu2bJeTsag4LLbKtvlYkSZE3GNOaAZauxwXTbfOD+A7gRJKdad+l
acfbN5+0tgu6N+GWlWboLYLTIiTE4IuPYZiSq55wBpUijGzQiiX+2hfUbk+Qh2/I9FOARdEL1D6v
er3TJ8TPmg2AdLT4bLDCDEj3H1k2nPk1G3yiGCvXh/NIdc6r4EBWSfa4nC2iQoxo+pP9q/dqs+CR
8MHW54+bNMWm7w2KGAf5gzoE9+KjAR7Tk+ffPz28hGKEZ5nYMegsXxgJh7i7ZG3lLm12RVqrBasL
Ow7BiSZsQD3Vookmb7ukLY+3EKLgtMoVev3IjTS+/y9JngC+7kkMUJS8qJn2UYvDQeQh7s1e24z1
j6Jjsg8WUx71pbgWQieuurW/j/5Sz0r18SohzrlwGRZ4KolnkbRLODyOzCXm22/gmbaHPohIXD8z
ta9V+B4NV10Q/U0ap6/H+brrzRIdFv7cdQvqUPAKWL3P5MsMlDK38zDSj6lu9H4sjXAcBHN3EeH/
TC2EYa9ifEJJbvwCPS0fEaE0NGzeQbco3Enk5GeHfbugBL9zbCu4gRxqqWIpNb+XvH4LUwqFgYYW
oMYZb6AAk49G1SsiLP6hA9/2l2N6coZX4zyLikcBLvh1IYtvk6aFCy5EvcZfbiWExyMFgtD3xRZ+
hXew+hGAE92L0kraWK9HB+dMpb6T1flBwZo2UeSib1+t6qxRa0wDwIZv2mM1vzvkr5BstE+f0lRo
/yrCxGV+fip8dCdikBCol5fJvALqEY+Uw1jaPaX9PZvxPQ++gMockk1Ik5alpw92XyfZi8dxmPBp
/h4OJadTyaANC5NdsdUtpgXjOH5x4Sbh6ZcR6Hoo2dz1TwrBNEqomj9IxP9nEyH1OA4nRTYsJUSY
xR1TjteVnWjB8b3xY9alJSDoJqmzg3IY39E6g8pD+PXjIZhgjW9e55CL+87CNkGtzxwvPZtK/vSl
/hT0Z256IaNZNTZzmWDxmIXePQkV8Re0jWWdKhuhM1RUokdRdhPIabSx0+VquDLMk2Ez8mrxNDIC
xVM7h7Io72BfMeL23jvSbmMvvitZ5H0/96qpfPQiLMxPV0hdN8IYlpr93iTisCzAp+Ha9zanmCC2
047hza8+o7Ib96DdF1GnhyZ/6yKtKfIX0n0ykBTZwgOkg94T9emf3Af5SUUFBAXKVynH7a9E3C2Q
IFlrkwZdrNx5WNIvmkm4boZcKqj6qmZEVQaUJIBTMhqNplCKR2v/x1sjM9pO1YuDnqYv5F+IXpJt
4WjDZ6+mVrWa4gz70mZPIYSqgU2LBxEsTJLaCJAqIW/UH1Q5kBZOal42DjEUaHTkzbJ05CjVjn17
oCyqMEiTjAaAF0Hqkwxt/ASrea1xvOiSTkHOFEnK4Rps4Rwt2Ci4eRSuu1I664m9vS18kfL1X172
DdXkJuQpa0963DgMkOq2vgbHTQYgMaDdSuF9W4RuITO3i59u2M6G/bPlQbiGq7LHloZMQod382ZD
XNbYYEmkNz1/2NOECGQ5AQw2yIALp5DvCcnHAXnmF0PiW4uR7O1acFcaolCBxR1BU5GWKx612NN/
csXPUtd/7ymwp8XrZs3twhShpXzNdDKIU3RvZm1Mc4d6I8taNRFt//6geIust92IuNrq5ZPhPCZO
IB3s8wo2jTG4Gb6Yp6cHF0rJ/gNLvpgA84WieUN64+DabcDGp/I7ChcEe/7G7NKkXYfstLUdNxxQ
P+sSaqfeR4j+BCXUU/zzKUUI7VT/9XAH23WwTmpmGtL/e9jqgkg2s1Q/gWQbTwzNDAYnlN/uVaKl
asdHOfjiAVbHTuy1PSDN89LzT5Ire9ETBu7F4y/KggeHnhoUFCjU1f6rUw1AHKQZJze7cnBVli07
WqgIpLiIDxEiMbb2kEWhvEi5elYj4JgLJc8Tqaa370FDBGgJzWANsWhmBuVSwRhuvAVKHX4CCUtN
bQm913DnBghP51sc6fnc928nZq8tY65P8EizBRQv8folWzAvbrwGXIbLyXRGiz1gpsR6ZiLQTUnm
ynpXV/JI8dAdky92Vr5L6o+PL8bQHotNMiuF1Ldwxi18ZV9TIpHQ2waR5f6o3SSedrv+e10LT2eF
D3qUmv5WqBmuFQuoYTpHkT2ZxCj4HDapq6aZ2h3eFOqQIH7/GCYG+vwSg7LCYNEweDhh66Tgxa19
ax/kZSGZ+i/e1CXS3XSboFt6Qg9flPv7YxPbyLgQcGoTPaB6vz7rW6f336LNZh7ZSjnIpCpuU+Mz
pPJ4lpZ563jSeMmsHhCGDEbHadFcWPCa2LvSpgClrP8FXlqNSPRJQ0iReJwdm1Q7fRXkqO9f04+A
uf/8HLT+ksSb2E/Z38EWP3qGSn3twvmSC10kp4VpuG6nHJsBoNjuhfO6n+M4wwY78VBF+fT7dIey
UYuZ6r/EUbdPdeuKzay5P1fGE8tSuaG0KwVLi2U807s3qcxy9xxFMP1GNa3AsHpKr6XaDaNpzfxj
Si0ZmncjkAkKJMx5WF7CcAYfvfulHmRyVU0sD3bWIlhXB7TEOfuSA1UMWcpnlxGAowHDoVC9ZIH2
JWOJs+KGROxGk84gGcbIuxTtt/0SYziVOymvAKwTpEBYdnyR5PcjJumoQtEEKqGExnmTbOOwbXUe
X+a3SV3YBSlTyglcRTjq+F0gJnlQdaFAIVlyGeCLXMLQoIT/tPgmLVp9CdnaRgDLgPrE065FfLZE
8FyonKtWO/Vc83p3CDUL4z+bUZw6x4CgaqSYjWEas9N47YB3LOLMiVB60SUlv3um2y8psC8GJJ+o
sgAyv0T4ykKFcajKhJKmveysB+lukVbedvHBemb9b19QgakkNN3NSX+eYBqAqe9EDzNACGMmitpT
7/IdlsOlYa0XIaFqfGMVtQN43MzPr/y5mEnOTBewuK84M9LnQK/JgBaEZDq1RkPpWvrnV+ElEc0S
8ovCUNOSjQC/SBBFfnte/HT7hgh2mJ4TKTKYBlR5RaIQoZw6WsmtflGeCUVFLETTsd/mf5j3IsQe
WDGHw9dqtEzzsSLKg2KimOoMP4rU9bbPWjsIoUpRfT3rT5JHqtSKA+FDDG+VicQGqFQ23COOtPzc
RXN2fgGzsM16CetQS2DViaV28kyl8jmH4yfin2T28d5G0O/YFfJWDUc11ZPdwTKnpIe9N9Whcw8V
yU/9hg6HgI+DLQ+MJ15Ds/ornYP3t1bEiGw/dPbEU3hmdlmpxFM87ZCoJIeP9EJclOTMlR0yLZeu
6LOmj7wpl3ETlcxDsxnI4FIVgaeJVkZuAKAMY+Cp0EcXAVcs1DIkHLUEESnGzvBTQVWnphhlM8LS
DhxmOeZ3KN8tfmNrUGMcggZe89mBgGSlRx3FpRhIuKcnQsDfIO9f+lkF8qhxi4FvEbslV+wl5mpM
3mSwxDjEVvctX5BqPjt/anCM1fcJe0s9kKqyDJ7bd9p4eRud5o5VxojzuC+fqK/f6AcwAMnFgKSl
/m6LfjwnUhWYnZ632LD6SvyVb1uTDysAxiYT0O10SDzUYZ1Gx8DmB3ijWIQxtOkAs46S3qfpYx5H
GA1BVamgBJ9iyNIPLQJJKZEeo1tXwItuempScuGvE8CfY/SFlD90k0CFXOyR3tn3oB9hau0mICO3
lL4cyQwZFKOijOTuk+eJz3wlqtjX/gsU5sMNLPHHSGkqUHGvXN0BP9MAblh8MNmFKgQFU2SMn7UR
zG2JFp4G2KZ9vFnba+7pj7/+tWr+pb5R3RNKOsoxww08w7sOb46I2c7UsUfPY9ozetMKiydMzY5j
kimSiCQMtjqA+dnlY0io4D8VkK6hey8yklROblrLe9BYvftmPjDOwCx9UOO7O+5eT0JD9B+TLXDb
2SeHmaePx81uYG+TfX6JLBTM7PuvgQQc3Uq7GVQuSD7IkmT8zjDjBaF7gwq516iEevYSquVs+tFT
M27L3I2+BynOeDHlFD/FB6nnvoBa00s0IJJU/h9fS/fBGHu5BSm9UYvLF9EJKMeZLUuf/juSDCv1
Ue571abQDYkiNP9gI2wmsTS4bMdk+I3qpEq9pM37yHr1G/R39+7iffobjnS9oUEM/K21duA2eoAa
zq7NzxKzimqt/LGjZyWJtDAQ5rF+0EG0TJmsBUmcf+WXZXMhLW5P0CPjSwafVo3CEFsFJ5rkNW6N
PGcSyrikDJPRQ1KM6bIsjxowKIIp0eDtIRAFqnG6DmF4zgZvmCA+FeF92cNYrS8sIqn8aWYSfm5Z
LrpFxHNWR/siTzHkribEVm5U/jtZySwe4AjyUQ0z1OGiAWcazzRX14xJjMAwPA22d0ojD8ve+L0H
b/fcW8C6+0dGHm5eZFfKhFrPmbVJWtxtoXNCACAdFvOVO4qPo8fvIOao4gi8hR60tr+zxN4c0pyn
iOgsVYRnp6kYtteXTT5+LXe3H2kk5wd0aEC+Ecdg7sWEPcunxO4Ixs+Qz07vkVATJXW+6zKYUTWY
zuC0ivig08qsLW4Up2LupVBkjulhaaVhtlqXO4+WmxHwHPzSFAQknTQUCWsyb8Yft5c05/7k43FF
aOD9A69ZzYRJAVI6iBQ6pzkC9ePpIQuBKsVkXDFvLIiOHVt4omhySrakACiIC2skps30bbXBfkRA
bRoNn6CRzFLdPdS1eRoig0ZMsK0aOyW0L4tbzwoIM/BLhRJveFw42YyvipRzDkxmBKjv9DfaRpXr
N4g4buJYKAdrH7s04sOgv8ICZ3gVNYtI9oCIEJWVrIrN4IZKjSuH1kmOv1VoUiUyNcj/r7qq7vHT
ZR7iHNRDLSCu6BcLB9l62Ng90ZBh21WDSTA5lsWYT8B+D8sAScIy3hNU/RsIcZTVbzXpArinShTo
bmkYgvNU/HBPuQ8Vbcp9AckvO75xTNzkvegC8GQ6X41BZfrj5sMdFu3XtHuMSJLm5laKxonjZP4w
f/V0gV5EK8lzD0MQkcv7A23f/ieWYZlmlayycvEgO9wui9b661jncyVXMkoxmn1z1gdmYsSL+lt5
qh9uSqN2YxCYg8DSqeALDOganPuA0KBxUsWFtyAllgbb+FxV7DWN8SY2rsz5ZDnEfp4xYXWNy9S9
ev16CuL8Z2O2gcwZidzcUjGn6sCgVIMUAtqUlkw+K4JNObBKdwvWS+fptywRl18qbJRmG8dUi1Rc
ARKBoyJYPbsF0/2sIl3ZRZdaSiEfuLZf7fNr7h2rz34qiJyNdsa/T1oQpv35doiyJQdtOlAXhP4k
TTP7wDg5vLnfjzpCtaCGjz34YFdpsHlqIAYXZRiqWjbvzOds+4SWjvKPUdcffmez4zQy5fBSrtRF
jOr+/yy0/VevDfdu5Dl6n3dtlzdGhwFfde0W+1bota4nlFxrgzIqMgchENO7ej6BC4kfeAHd0oiS
6n+bRkuLJ8xD9uhAX7llo2W77BuKvLE9RTMWmS7xoUooIKDpOnIRIhJCwcMVen7w+/rVu16HJep4
QPeS0mtdJoSgyWBV5ZRfM43R1Vq3Gn/cPNqf9Q8rooaDyAmQlKRD/DqSPAC1GJ183Vouv3ckXb6x
FeYvrFYb1vq3ihc1od34CAkpj7SzBqCw2IZFZXdAX01JzHg3Uv9T977vYNbpEt5k0yNdfsEZjj5D
qRpA4CGSEiA8E6fIbqTmyDNhJGo4WN2Kzoq6I/PQow/t5jTsaQs1wPPWmgQYCdRngLJdM09f3ZB5
PwN0uci5IyHHoXi84sD/cN5yUrkjTZVM1/BxVjU2ruvG9bYRt0S/DuApOhVGzFRudv0+ag4XHEjb
EWV7gMScMII6pVxKa5TT+M5EXFwYesWZSUEtLRtTcPH/j6dau1XMmTDibn5u7+1QkLQqjwf6eeTN
ztHhGsPkY8WXKzkBuC9hWwLL7hsMIVlOkQODVgs4/9i6TEN2mCdjufgIpFzt4LKG+VUGZOuu0+2E
pxicXyjirxFJHcwiqQRii9jkHqheO5mQXIlLDxQZbSijVV343/SLG2ma6DucrL0PhsZKYwvMz8ql
lbDLQmcTUyzCeURNZXO5tmtV1ppHuKxasApN7a4bHQZagxYcasLOyEgyiCexbnadSzL47JiGUeCI
Q+LNl6CnV3t/5n31G+ergbCrOMfPqNXugcfzRlNQAwlRuTb/bOY/shtqpIJQ1Fr9HiOS9fsVS37x
Q3gi/35iF0Znz9rc4sio7Yw9Sqb3iccllkuYpl9TbqfWAAnzb+PVPJtxvxlwSo1T48QESEth4zFB
DVzOeFTsXd+Y6V8PZS9ziP5ma69Ym0nf2giNOX8cKEmyOaOsMySd+fJpanFdov3Mk/aLPRlToYXx
T8UL/RIHZHmFijK8wsADUoXWc/V4Hm66JSoxQ2+1D7N2tOYQ29EYN/wgXztdj2WwJL3w7E6OYr3J
j6Uz/3a8yceDjbH0ydXgO6KuYIb1tgBCP+cKWxeKHW1+L6ra7Jo0Nznh5YQs0OYYJ1gMo5KNTpFg
scUkq/4IWDPfKO2uFdLKtO1GBKypG8UIed54wQbBoTEmHRQ5092+EW25Sg4rAom/2rcafHSyoUCM
2Vk1bHOEGAYF5tT1Qy0j7qp+jCa9yaEDewasTWxSjuvJWyfTxKYSYQt51ZgYuzWkJlqFK94+pLrv
BBJ5ExKxjNFBxjIViJpsblw8Ab0P/reNRf3SduYy9bxQfDbCS4Kq40khd+l3/FtdehrdeLHeaxB2
qLGTTL+sZfNwf/Vj22cnX8yiHNE9UH2caJnsV8fTYMqw5dOICs8rNDQiKNvmq11DE0+QY+ZG60iE
aGPJWzpQfkjz+SCDE4ueXltKU6NRyiwHLL5wY78uL32iCUoFfi8KZu3xDkCpDtkzsXf6vjDOAWSL
WsLdNIdY2Es2BvzUeLKEWJue5lo204AgQNPmJ01N8Kj3ljsP36Mpr4klOH6GWsD+sWAhAKUZFXd5
N2uYzUv/As5UUw4oqQb1voK2vRVogTnqaepk97JU7YsaxgNPuM/YyH+by0d6bDHz8iUG61ODWnOk
/0iu4NPJtqTXZfSGaSm6SrdTcJUyKeAI+ty6S/uXcRZDFJ+eUr7qQ6+i5Y48ShZi5+4SKUMAYERE
uifM0Y9GGa9ZHn60F3HNbVF1s1e1+PH7fty/KE/b73D9FjYFXA/i8Ci5/v4AdmatDMI7UIdSY4Xl
DACcxuldVpRdYuTdOzGcFxguUudXRsvZZ/s1eUiqWA3WIyc7Hxqe+tLUnoBa9SC2lBQI+6Px6b0o
Z5ib0i9+ubXrv4LmCtYJgBb5lOGuvXYlQnagEyA+0XX5C9IVjfiV7uA1WT7prQWH0tjkZOJQeKSp
z1R7il/idaey0g1XgeDUdIphXOVJAsQkqbF9T5ZR0JLLm3fSZTmrUsHL9AE248nbAL7Bsml4ud3C
rDHFrFwo4KZfEacGFGr+vFlGQ4kbUYTLK7niVuVK7W50yo5U9HtG/rUDqnSfCcEz6gJC7fcDNjnb
6jOg1HAG7YRb6+XULS2bYCusv7ZN6gwqZ+FVnFgGHEzRME+Z/+5VVoowvr2DP/Cd93b71cEHX2Dv
0fC6ITaHuXZYPvPhFz0ORthmVnFHfv7QeWVQIQmLQrN2k5EUet8d3daUZudtLzA8scv70NjWcOT4
hc35865Fy3qT9o1nABDgsv+rAxYNpua6SFxFG9khI/AKpo76mPsOiNUYlcVG2xxku5aMfEnTgFWG
2h9Y8bP5+R2XDcaPNLururmpLaRZsOBBithtX5WzyXQPJSAktZasmFKD2AcMtC+f7DBx+KgsvgRR
/Rm8d6/u3KXgdma3ZjjWaZLAnpsm3YhHXZm/fj8cvVyxcpDZrIACQfgFbezMElhFkutZTJ3/JLAs
rtvk/EFAWRkg26+iXcg5fpZyYk3lx0wr+q5IgVvpxKPspOCu/5BsWGXuLLq3aGwo7S3QpDdJSApo
TiYRuT3LJRs39GNe+RBnygTgqW/fkxN4T6uAiQBGN/+TpyfwLchD+SsASldh4/f3QWeQcWHutQMb
9rS9AK6ZwlQsAbJ7VjohxIKpRxb1sMeQsg6hNu4xz6Mn4AuAxluZM6xW0QaZXfBGJ2OWafhabbtq
AQJWO8su5Ai6O2Z+OTds12WcK1bC01m9VqUgGQXWg1YZYoNsK/v+GbUQsM4mfdy5rzwVr/RvMqDl
+H4PHFl21BRZmM8PQJVjIPgD1bnGA6QevnayLN20nofsgXeUFgRcCqf0VvzTh+QrLk71fRldoi/r
j5CWlGCMw8YMxqLTomB0OF7SyWdm+jJuWaRtg+PcZdxmlZ6Be1ScM0JHe99UqaGvLBBQbC7cFij/
p+nyrQMbKwZuJqCPjRLDWHcCcuHUI/FUMO1hnsugknCjcyPgp2wgzAskorrDBV+ZaneWxNyyV74G
CouDsIUsOv8V1z6UqJiF/f/cy23BfUVF6BnBhP/nT0WNTSpt0ffmqWH4gS0lYG4dlis1nCRpdkdy
WAOhfSAjAIAIDNd8gwuuUC0AxZVeiNWvTBk50NBwRjdkk9m8c+z8ntX+mXjlBAP3jS6YiPya8+8V
dJPOyfjOCHES69nXz1eXUywluUk2SVs9+JAPOAiDrABYYDEc6uJeKhPgXg8Wu0Dm4Es7JhvUuoMD
NolJtn400rMNv2ZXFP8CQ7i5OUBX6WABoaOV0W+6rLO3jvAHG/jApahFjCHZIPWEM5l3oIFuCVxb
IdLIsWuUNXo8J3oGTKWW039umvtuwsqUmKNa2+ylopjvmClG/h+RYMZjkKdikIPGc/NVOjnnKHCd
W4XFaJJySHr+uD7hSAyP8u7hvNOxJS2QWBwJpRolIryDdP3S6MX+XxyfgfzVvNJDcU+ZJ5DNrAKN
X4MIrRPNPMY1yGrh5ACXBaI606IVdax6l4SwYDXlRfNHcAhhu/bYdGKDBK80ou7+011FbAbPnoR0
lS1APqSrFL8e37Kw7MquyKx+mFxns4aFxLPMRDn+86KwlHtnGBHPJY9eOQ2qAsikZ1eEQKtK7u7c
cNGZDOosAZ/DLC4MqQMnO7n6eCYiDFYQmuE2XOJEx5qhA/mF9LMyeFlvjsd6fhu3YwKHtAr4rZXk
Kg3VS3fOQsMG7NzwVrGiu3wfzpQiGq19dg2Lers8reOpbDcbrVwuaW4r2uNjU5K9gR3fymni5hub
FbIot+3Zl5zhBW0ScQ+I5UGZmhHSdo8cReIo3ezXV7ZZakq6w7INl4mvFBk6Y/qif2+bnpZ5pE6N
L9gU1qvAiB8hER6+QRtMghhw/U/oKSZKShnJ6Jfqj0/r4Dm+M1pFcw9v/36dhybfAVUQj8r0X9xW
hFGl0hCf9ubK9JCLBMM92BmCuDgsGYyIH5jqGt6Y39QoYILcI5HrT8Euc/lywc98LsWF/pKUx0ol
Ogx6RupOOrztkL+oM6Tble7khBiHbF0QMrxrPeP+qLxTQ6eqzjxNik9nsUhbHPy2JF898i6brQK2
LNrabk+qcBeRdfQ2CA6qr9IBBRor1mM+xrHO/+q4CgDjFHOYjk8V6LWZOu9uUkuY1ogpt1IXz02v
CoVHIbVAau4svtK3YYUbSiFrBoLIz29En2aiW7DKe2VsGzvYNE92Ni2CGcTxJOSL1ZdULkBE0N07
TKdLuUoO3AGAPp6CX/OQeTmDig4Wi+n+L7vIyv4h8+ix2IB5ESsWjAB1IcUxT3qaEWH+XZRhIeMp
BFs0mFKaZKC8/3ELXmLVOBQAJGIzGl2ReyZWqVj0QjyP8gGU/7YnCjWchqtaMGP5TSAP2P4AoauL
mQELVaACTXXVxKRnBLqEVYSVT0310Ro1UKMSDsf3PQQOCbDp3gt3rOjE292ZUYkXLmwX361AxXh0
SCmN7x/gFulyAH6TMkoatj4O8BdoUoAd1y8i3llZaFHF4UHl80aPWkf8JU9akMg+1HbsTO0xy8+C
dxNbE0Pl88bXo2T5hdX7lWexEuLZ+MGAfyrLEBn48Pi59tYQIxphs/C4+kZwLQ2lJ9coCEaR3OhS
0Gmzhg+PSRYR32ofwfGCyNqQ8zLjEdiBP4dR5lKJKWWIsU/kox+vfwjYK8dU5QpQJYamj/e2bt+m
hy8x+kbquJJiFfUXfSPrUBwujPplSbw2KcxIjXMGz8/lUxjXQbvSKbIv43e3cIGVjGAcmdAkb9Bb
CVrPcNsI7qYztKOJoIdmJEX2LxR2XwhKsXZ/ObSpwbG+FLViOMbu9ip8TXy2MNsC0EA2QFeCfLUn
opKCeo/T1bWSvv0LUpwlCxFAqlKd0U8K/TSZmVW1O3DW75W+hbAI72CifvPwNny8UUQKlG3M7ycj
9dU1SBXDbHvhxkgJROFcMWDx+TodIZrHjjfVlCUtgicdJBm226GG+ACWL2vx3Am8myUPC8OhmhbQ
epaK4a/QteRl3jMVT7elrgLTpZGB1kJT3cj9+TeU+wha2/ZmI4LFHrkRWxaDn6B9/qhV5URIwiKN
G51LBcoD2eSqtXWO5SpjxqDtJkzLUwgQXIfr9V34PhvabHqIkXAP6xJVZaP76hLf1PD1bxNYSxB/
e0hc1JCjFnxTX0O4F6wbF1srVeS6EJoAaOTvZiNoRuUqsg0ghw5FnR5c0baEj9QGfHkbGXrUvcQ2
5/SuCByVbJw4bPTl73xW6ORUggT5cmbMIuJMWEiu35Eiyw0tLB4goLVKqISQvrpJhWuGIc5+nK/d
8fJriBPTcPi/v54Mx6FsRsyFHEk849b6HDqxU/Xu7cLKFj8kwcgQJTPF3cZQFaVHAvnQVWJ1WFrO
lLp0yI44d6J6iE6EzS68v2mHMsGMTC1BqPics6YlX1V3SQraEHgZX2hlv5+inZJ2vc/c6HwMlL0n
UzZNc9PdHBqrZXmwdsdV+nxTEFsAWj4ciZjnmcE8bBUgjNaiklZ4Tm3uazv2pnccQXg2VJo8el5s
Gft3ZTuvvoETHH9taGd1zMJwaE/frJjbAwFMw8EWlDrO6jet9H42R5X6bIAejw3X5zLtJJwaUg+X
tiA6k2u7l7yc/eWDS3hzf2Kw1SojQhtAA/71LGqXceCapi1BFxZikvkOS5jAWV0nMe1ELh2rNwgx
HFQnFGZxmQKrcFeE8hrZZlsJ4OJNNw+KSTU5fqlUaGUYZRbuxi2DlOncmNoq1Rv7W7PVrZjgz0I1
pT8SMW4sb6CuQ2s9PevHktLsZbTWFVO02MNuYC8D9OpnuX3Cq5bczOgEEeLgjwEZRkkZ2wNPVXgJ
UZxHP4VKR9DXVd13Bumg+0ie2zEgSECOFwejfrbC16bVY8GiJ0W3jYu8Lwrx1wOfQ1XvW7fv3pKZ
Hgimuhn/oqm6WEk8o2sPQxxJQx4ozRAFHTxsLiH41qXoCl8FmDZvsXI6VaKBagcRHMAq69QFrejq
BPCw4FXvZQEy0fj9LtTQfalCxu10wbU5b8714CpmqJfhDsLqnoJZqDjagQHFCyeJ4w7XuWSy25wO
Jl4wVxdBoW/1IpipSFUEyd5+z7g7pNNfwYDYKfdGsjL4tlX3gQXt7m6cxICndZ+PhvRN604Jn5Sn
PkGj2NDNsiEp5UeLBPFYjnQiXNlFq6OBPeaKt0XH9LpRkTyAP85JtwxpxLE7C1LFy6+ny58bc8qX
F/2txgWo3ho+d6pfA5JwV3MRLEJ0BB4460EYwuNa5b+XRTrfTB0xbD3ZdkqERwtHgGLY4FBVBfIm
F0bXFVeDWfD2XTtFYMukJFtpfdBf8JBomyb3UQtd0C6DAMATjQbrw6LgZdgXoZozom91jrhn4Lpd
3Zr7M8cKS52t/Y4WUlJGi3+TDxJlWX0lUIMDBNcqexvCwaRMJthhQnt/VqVzSGdO88mhZh1zKxW7
pH+qH51ok9uEov52bY/RulPRnaRCdSNx2s3Ah69/z8m2gU8Gqgb2Nr6Kypxl7sU+zjHifGzCA7wA
8OQM+baduJwAJLPJC4nWMV//3qj5ATbnCuvSY/X+EVRxpWH6HkM35QY7yyu+Q9jgH+WJ3LkYBmGS
3mxlug0ZwE6qLAX5cnH3zUwt68E6eMyjjsvMlh2VjznZcPav4B9bqp2vmVRTSw+hf0GsdE3aU/nO
7Mx5Ca7gTCF5jowwIRMtvIypEtpgqFaI8nKZ3FpdzcaD9nS+6kSntZvE25+77PqaWcFWaH+e0nuD
nz500khr9IQRy1s5y8OsuKmu0fdBCq1VrTTn+TWgO+6qf0ZkdpdDZED314z9rzJODhl9POpC3R+d
rgjKCoWhEcygsAC1sXqDB+liyAKVFrRmOmc7Y3fdDzFjfjr9AUhmlDv8kNiRBjVzr7hkuD19cyBu
nOUBwyaGML27lUvtu/iUsQ8/9odgV9jvbW0LyAcTGTB4lLtpqegc/l8/W1MFmHJs4J8hSG+oSUp8
WFCuHgXiuRD+2sCXNSgZxangA/TPlgr80FxZm6VRU6lsoM/+az0AKjIu7r9PiFOZ7q9E3D3uwy5U
NQxCAyXLg3Nz0Upr8OqorAhnoiAKfXTvT/rOOjNdcbJOXTyIjIdqFHUDeODJeGskQa7fCe9wCnFy
7Yig/9q7IrBUBJIMp0jCfnmb1NCHrBLIybbdI6NVqVqI9xVqi9FypTsxT4IF1Y+MdyXr4hNFkiBa
cJ7lg72SR84EB7WSWI06EOg+vZdF0V544uxcwVcc0sIINP4gxakXLoGlLsY3nMmbokKzR1jysshD
GJ5YQVuVjLG0kSst8U3dizGqsf6M+iECUHr3uLPNNBR4hzhJlQG/d5jhrdtrrKKiD2mhbl2mHzKN
2WBEugOSPdZijyPdHYdlg801Tqp2PNUw1E8nqq2G6UDSOAbqGr0FbZmewq6CN5x5zBMRx27YuKHE
smenNfEsSMDirbuej9a5jIcLhDRCSiUNC7KkzaedtpTjtM1WfY0nyQ8GZA4FTA0ufI/5EbQsJt1K
uz7nrErIJeuDIJXzbuy+B8qqxeMRlHCfUL/SjAEl9WZW87r5+hO7AYoliMByDrg+YVJGDbw+4vTV
v2qdnlV1d/oX76ql7Wz8V8/USFgeAVe4JBn01XDct5z/vs/2Uk2V3OqadW8heGORXctmWMhTs2v5
uyJjAO8paCnYaa3TxssyOVG8C41SEILuf4r/uYQvwHiBv6UFHZtppKJZ+MBg/Xt7MBk/+w2G7hAs
LEmY9eFEJzIcrWv7csfqKHYfVSXOsRImvl+epdjgNNXH4FNWJbZfqI6DgK9xONIXN/RsYYdysefO
9+1P2iIoJ60HI70FKh5DXgUr4mHbwWdjC1TimGp8addjBfuOAUlbY70ZdH/jsFor2bvt0b18IJvW
F0JxUL7Msxmo3FZuUD3helVaWseVvcCDnYGHAto8tuTMEl1UBJCxGU4MYvbJDcMXKIsUvh+iliYj
n4GjAhjV/HSeEkiNgcEXcMVrEMcd3FeN8aL96iohUbqT1MyLYljK8XfRCIzxnuI2qzT4+AvZYJst
b1uLvkTdXzUdvYWCwUaUqV4WVdiNMBid3i9HidvGpkFNFM/qZbSOPrIfk0Ov1Xv8aXBOzwUnE0QT
Z+BzwdW8oF414+DTNfpcY3OegJo54y6L2wvuiwi1rv3niF0wLprec6g399qPuy6ABSds6pqeHmMP
UkDmyVaPvfbQR4HonCBNZezbdySJ1bkmmMtXncDKSDcxZYSU0W+tdvurmtjf9krASJd+Vgv93PKz
LqgAhslIWB3Uxt/hyrxJsDgExsRRi443d6ywdx+R24OFRhLCCB5DlXWN/IqWLBHvIxVWJW0NXzxi
1uIDNOx/UatLj0J1sfepwl+MiijlMKqfE/m7zHVmS3xcl1D6ErtBPnEl6lALgZRcdY1Zo+OmG8FQ
3ytamjncU7NicOqj0NwIN82gofckr3cgv4CVQtaNoGvIRjgjfwgv26oH1vvoLT6EmfujJkOWJibg
gzgVLgdelfp4DJcntkGeiOgGKdE+k00kmyMXjiwiVSDvBzmJf4mB3C01Ys+oL0WcIBPKx+Bm3W2K
yPCewU+yRV93G0P3HsNUOiFlIpgbgYHLL3rtiW2iyi42zuoOV/ImCRAdjGPBDtfKVRO0M8+s5w1Q
CvYKSZWIZBnCJSMwU0r6oJbiu/AMVNZYKX543FAvYnVWIXLIIYi/8/H0D1W+UABHAD1gvhwBoVs7
cTrOmVyffnP/uxvhFrQkV1BKa+ZlhKs3owD2GGnYDCWPZ0c0lArbxutwM/E+bCf4ZozSPmRAuQYo
0KLGs0s7My7t07sdIupC5Zs/xDzEf8SbUDt7kB9fLb6y+CWbqKuCdNblbe56RBHDjSrIbQZ1sb4M
VuAMLO6bhUnNN+VhxYCJ2HuMytOnGnxc6hh5R24FporEpSrnXVyJAoh9jK1ePcNx+TMsh5AbLim7
JDl5u7guMdhGZBpXk9nAE6egBj0Ca/lteoyyGdrEQspPf7FtOyBnQNkF11cXbibmRl3ewvP1B5cB
piVYPdybrsW8GO46tjMNKnAcUxMcTvAiqTzGifmZ65Q0zi5mJ0u+N3NhiV7OtdWiNeM10VcT5iKu
77J7A4/DsIvdbioxd5UtTIVwv2Fqgg7YKIKf2MBXT35bvyw2W7X7vOipzaZS26LiNoMmLkU5dDgI
mEzwB6UaiHSQWObZVKtQfmv9q3UgA1FPWolGHlEhUuNidoV/VWPYONgu0TwR/oQJNSkatagrfW5q
4hS/b9Y0vGck+M5hhKod2gA0AMN21xt6ktavSgXIdEiFvBxh4XhedRhLn9RouHtE32J2KSz9KXOu
716Lcu4KyZIOMe23yMZPzddoSN9nDLcNU/rmGpCm0j92iwudKGCzQEMlhkU//NcY7ByKvs1N3q5s
hZCIZ7eavytNkefp0/mstaPzT+fzfshSHxPulGMqyElyu/NhlGpSr1Amm/3f3chYoR+8l6PBGJMl
I0zclQqNLKFTvZPYohFsi68f8BxiBk0iYhFgBYs3WlajFrukRzXGtIGGLS2zdyjIpwyBtwgT2VKi
MJQkWdq1hPY7guRzEZbclJSEbuAGIvF9W+5Wf/kWuqFrDwRjycB4nKYHslsmj4ZNIbf4N8N1KIz+
R4V6YDgeTW7Yh+u16YKsIVLkMqsjLIho2ynzoHU5C0jE+Nf6RqRgdb5GtaULq7d4Y2tpyynpy477
CGjcf1lnw7jEVXOqhSe9Dcqcxy2f/N2o1rS3af3bBo8HG/ZjefuFwkQD1+u8ALK3DNW9QCUKIpHH
tV7bNBjO+cO1vB6PX0CoFVCM0iXZ/mnvi50B4OtrRPhiYPGu3uVv5XfomdkLES9shPwLkmruLxFC
dgvVmQyk7lHMFRzpPzLo63fDG/buvRfcrZkOpfuH4hjOqQBlvXO/kG9B7odhmfm1ajhdV5JR4Tqo
1MMt+8+wkFbZWh2iXl7JnvJPKqHURfrPc1+60X4H+HB+OUEWZwMt75fTxCjpf+FkDyPWMuXoNOaT
DmMjR96bSSEWN7rf0J9Xq4fEk3VmlTTrOIV+lOw3y2euipCxx3pS3CsFyA3a53BrM6ivfHAtYon3
67fp6zJvJreYHNlJukLGPYrG4gaT33gbUU0DJGoSIF6dTiVgFKUr8tNj7Nlrp7Y2fZPqs3cF5C5d
MQ2dUjU+r/wUiqR1pBXL4xqXq0rkw8izIDT/bOMm1Vwzmk3tzbgoHIklQqq1xO8m3eCVpxt5DldN
dKlKaBkE0TgYxqlfzUnqqBCpya9lSb9+ruHnjGi4mimjUt/SRw/jShU1JfmJSIjqVJAOwYaZH23/
nGDXQwt7gtVwmXg+k81RvhiF3V7jEK+FjDiV5WRq+xWNXEreGANo1FzFSXA+StMykAbp9x/ZUqJs
IcO8+Ei2ooTCqnVynK7YTXs+2IDAQWUZqrdmlAYc9zwPX3Sa0uzppOt8pFjNHS+hkA5VRZ2hFIP4
wzcEAK7YBmkACFCEXgNE9wQsSIXgz7MDb9XpdBTlbh97khJx84T+6D7U4Y7mthTvAwoYv3dP4i0j
sdDiOZUmfA8Z7QIbgdHe3N8h7nQwk1tMIT0Wp1wYXD22B4UJaQApM9MwxIL874rRR6WqVTEdEUed
/SWoW5aySpZSe7cgr76hdsi484y9iNrWGJOhQ9g6WdSrDT/wIEpdEiwraviCwLElMsRwbxs+6gbS
1WltNZouYTgTuyKL/q+O6G4zGPf/AjVMqW7RfN0u5d3gUkDy+Gt5Ei8oZC4jAYGRc7uPiCpL1wHB
QYn3uDRxOkTp2jFokKHgX1ZSLi3rB9hLPfE17EKpJKlK79R939V5ulTrMZ05aba67BY0VVLFymPp
zinM0Wyv6kKZgnfEM34OZmNytQR08vQ9JAMwlHB+Pcd7adH4PuY7pW90Rel1PhOzC6gdPC2Go4Fy
I4L3QaCQeYZKnDeal80sl10cfgRdeC8sFG6enACJdXyhwlTTBf0jtvIW4TPuV8HM5qTDmX/wmKEB
hQRX/pnjd7aa6j+UE2VDUxj9w+p1xvTF+XIBD5O9HVHj9eYDhfmFBIbZpP7CIejwGqR3oE7m6RmM
GYDDZLW6E3B0JVUqGCGiGlLV5ioucI9hYqRT/fZyqKXL5Bh7w7ZTFDbik6ZxKibujP2JE4XV/Xq+
aUNcTXWu5LzRbKEUeZV+uEvYTfnTAxUV8GkgeeXEqkNAZi0/2iOZhVRTp2CwkPRdP479PkXsbNHL
+GE4eJMn+eW8dnMY/YaAY9D8RxrpD0JteE2Ag0jpUPhUrTo1ve+0zJAJEDmJlk/MezGPwM9wrl0d
dxQFAGZHvqQSzVGmusWmK2AnBvNtE081IUi/e+kMrBD18U4M8kCnsbq45ARlfUlhG1s/Tl3/W7YV
qKT4g4e1NuusrTkjBf6ybY+DLCgvNvGTvf1KY1QAnvgC8KbaiNslshT2rH2taZJxZ3/oYUYBsoGY
L/hE8JMc9kXE4VXQL6WuzWbgd1uKAG6P8stxaa1ybL9b1zpsA8bEFhJZMWl47bbCpOdboh+n+PVf
8Ok5xF615ogNB3QGVcpgBmNVKOwF/p/PY8pmal0slfg5shfEpXd1Q3V2p3SV8DIX2HmAq3UTLP5Q
02kUH2E0LivqtMHxNJNfpAM7RER+2OOaj3zvjSf1OHs7POIvxCmy0q6w6O0yBTgxIjUD+CPY9POX
wezsed5GJfXuxjlRnsIsPp45hgVG0gAfK9PszcK8eeki10tokTMVKiLm3zXuHA+tUwYGP3ccIPgg
s5xQr9SyHHNS6L3kOsV/ptFWd4JSEGqKPLJFynLy8Jh8fFFp3vAA970jschXoSYv+KYrQQKitnpZ
rpu807Q6jD6XO5VfI/V9qyXHC2I293V+wze4xoW2m3mI424hpAndXj/7N9dPzEu3MwdIYTPIZnLL
7MTKGfOZy8RNm7Gq9GTy91qfGrW7Gyd1NoXYIPZCJAme9jBkGShoUxBR/pU+R03V0p5YDUqvvPva
njKjghpBMdoNnSp+CKQt5TcyvRsFVI2Juu1JBNwfQuApkqJe5l0xgQ4Q+qsCw0ps1ckjapcFR64c
AfKatS5oso1VHW3kA5pKbUipbOBgoEg0xH3RGlrGYCtbcYIUzg9AMcHKUwsMGKAIFak4yXE8QyuN
hEedM4FvYgn37EwRAsmOCJXmQMwCIQffBI4YkSD8YX0+cqqd28PVbVwF4G53uTX+ihDxpnlKNBkJ
ETqwg3racGVVhnSFR5cDPmDXGryS26m869gxhpBqhGpnuLCfM3d3HDLlCH3nHfSoG7UyRkWfNolm
b6So7yWEffBS0fgSiSA50KljiuUZ1ViyZ0TgqIh8cdtoCxTJTQFYjgdVvV8v0/eUCBxL+2/e/iHw
T61JsDEYWZLTFT3S++ZTds+ale3Cs3kRDf1Qaw+2NG9XytTaXKmsrzK59DGhoEXq6pVkSNSCHKdw
8O/ebErVAd60tmYPmcU5tErm51cA4BmFo7aEv40h/xevQF+ccRW9uKLWrV+1cXwrhAY7C8RXfce8
H172SwBbEiLM0pKahralHGhUMrPDhIccy0wkkLQggSttjXfRmbDopebQlhXMC8tEoK+7Tq68enPU
XLCMOnoRzpbgCyQcKDRp7de3ymKA1hYANjdOaJ6LJdIykDSUIJYGXCcY7HdwHF/slBDIJQQTm1VZ
4PpQtfnUjBRsqqtAEU3O4AozEzyQTRet0rNvvxTJxBzWBrF6pPygmXQP1kv1lXJXVNVVaHnvbfp7
46cu+FthEcVGoFH6QtoAWH1kGoJcawLzcgbFM/J+EHhwptNv++2QjkZ8KMDyTW1Rbl2owKCsNmwC
jr9N9ziua+LIocgG8GKMbcVvwulhVmmfiWr88xUMr1FoqxySDjEvE5doWfsLm6mnXC2JJgmy0zb2
rUiEhPhaugcm9micvyddcHwX5djCvHvPLREAKo3EJyycd/ynUnZtxSelIQyu4ONSimUDfOs9w0ft
UgFBbm0Gugqq7JzW5u+IhuS9J85/De6dZ1YEjjR54ByW6EEPWKfACv/BbdobbftyeWZJ2HKiAjq8
j8TQ1hvyuFx/BcOb0OuP+VS80facycuz2eMuQFwBTuZpJiypEM/N4XizAr/a/pSGW9KGOwsjSQl4
CAzePcOxmFvTn3dXUMVvQj6m73LSpHhXPUuhEoQdqrapP3INHcxilz08XcSmEJ7SRklr+tRimeyt
S8Mz4/CjowPOVSm+WzKrLsMEFHcBzML1JCVMoOt/ejeY1h7hsDDl7WHXDZ0uOkVIXK5DIRXKOOBX
VzXacrFu1uyumOtvQaJ4eB874Jx6EEPWdWUR8Q6CCL3IfIYII2rSHh+/heUQnKEnpXzV+4yu/BpN
qHWV850a6EKl+2ThkDNRaMf+yvOivCMUlVLTNZOo1fCxS0MuLO2ZT3em23KFGnBDIjGZ6G3A5SR5
Wge6oGVe3BJ+xoBY2IsryynwUwEVQWQKtmcoo3sF+yPApqQQ6k4Zh0bIOakWuVThUaWxv3vmuj1n
k+anIbKCTxyj5JCnbhWUZSxDemEM/Kwl35O0QPRpF+KN+ibRSNdwz8cjdMmJz9o5AoQhUPDiAwr5
wyKXxdW0xwlxVcq9R2Rk1KL4sDNSPSFqRVUnhZOLXHC98mWYa6xe1+FzjNoK+Nnz6xPy+C8MtEGa
caS5pWkvjyVPLM7BZVssVo3wkNvDRotxPdHXFBvRBPuer1bZ29VCtSa9usjG9kr1BhwEXikZVkw6
3GUD/rquVccu1CptgtGw0DmGMeZ3Om8cozoSq997MzsshOS+KOq7fdykE6aNuG1H2lDkrozNu8o2
tF6GPc9xForSPiJLm5ObsAWrtHEHqFhKW/2shtCfMJEMCDO+OYzzsRD16OTOpnX4E/kAIg3qbLsM
RZ2mPD8aC/+zOu84PbE4B04JKv7uI+EuqjVShXwNkD6e7z9ZEuPFKTXX6QXYzC3TTaRMN1Gr35L9
irYnXRh9HbSqhbXjU0BrUrfn27dPrjdXhKTTSYYMf2/cHZcH9iVDhdjqE7oYY8WAILfYxablhuFw
ZZhldKVdrumlKDsSoVbNQV5RFM0YdiqMWYg37hZG2WjsdNHl9uF2QyyVB7DZh0n/+HyGiwHxVzz0
NEJ0j1DTwyLSjKbSM4U8BaPPCB0jCYivJITyt39eN5kkFANC7ULerNZzBflO+6lEj29+cIlcW19l
Pn0zzXrhe0WTIjOgk5fCjslDd2DDW1LWPvZFY0rzapQhIfompYl9LpqqkNTlzS00PDuQ4Oq32RX5
905MX1paOESrnjQn00wm3oelBYrnTjVHWEjj504Yc0NRGPXc9hjjj+/V0MF1iemVMJiqtMC/JJ5h
bOIN1S+x1dBGYltBgmflccQ2REhzH7UeBcznCW3hn3HLiI1rY52pPVIj2o3tknQqxK0PJshq1SZo
s4eQ20jhVAQAMIRUheo1Q+MZ5FrGpMAMTE0Fod4NBxEymlP9huaE+eJR9WElrzL/tBTu6b+DvUu2
bArRt+9dnSxPlnCg8zB7p6ZSkC7w2CA4br9gjZj9X6c9LwDwd7bIATdnSnlUlKV2yKFhBv5UbeP9
s9k6Up0+uIBh7mLzswndpQnRzb7T4DyBGCLsSzl1xhdQ2DdUXuF1WMgQ63/Oo5jN7o47UrAzurxz
BeOiZ5yzTNPwi4aKcqY8E9sbDZnWL4nQYUDYhm5YcjECXdNIBn++icG6knIrY6jd5q+vaDgE+cW/
5YpA3hGyvrFOTFDINVvfLnxz0WxCdP11blYpFPITnhSvmGYcau7SJV2/VJxWgZ5+iDTXath/grT0
SCf646YbyFOrHUxRJUtBCuI1rVuV/kzndADAcWcSZ1cQPTDnTsiYo80FWw1fzn7VCJuKf6mBjwiO
LTgrlsal19X0eK6keuGvIboThyZXDPo0A/UiZpWFc+4pmXsqjA510ZlXYuSARkyUp1SYFT18t180
NIIJv2ysMHeTp63DxVpudjN1PCr63QzLsCw31Y+q62StYmujDuAQjISfTv5WhSQD4ngZHwjva4D4
YgQUY5y8Ko5NqdWddXreERJ+6cMMhE+RzB7rbSShBcsh3GQJLqhK4p++vdPKnDUzZ/TrTGVozqxQ
V0KmBDWWNjPrC36/Ih60fsJi7/BkPb10aOPn6BWKIO8sLK1hAcE5l2QgAh3UP15u5zWoC6vHb7en
ZkLpzMT5653mxijmIi8hLmRsqnnrNnwl34i9fWrwZQIrMt/hd96iX94do1JhNA5LfndZI9kzw1RL
nwQo4WaR++5lU6sxI1DCA2zgIPsSCdwYMGqdIUkJgiG6SU7147DJvFFMjSzT/PTgu1mmKkCxfWbN
a3r/QMKEuAxnocGToPnCqLD8TQFtAQzm/2qLbJCUdaNJRB0K91gI3XVsBW+eRCyzK7w/xDU9nU3/
JbkNVgRL4XW/rXdTCY9qIkF9yj7Re6jehZNe5iRvBOQ7ASsW1Esbl70L5lMYdx2hDbvYMgKdZsPo
tQmr7RSSoLkwoamaeK37+eF7uUIybn7BKDqF6C6NJlVc4Nvs//2HCKAkr1D8/+hevlSCA4mhPIlc
0no5ScLuQsp0PCC7qRISfD8aA5/5H30pH4HwYEEZXa2B6x0ZQcDukGUC+PtxLGW+1wmmxPLe/yFo
BoyjbfSF036Uzv9YcE9obY1H187XFWCeATIgJLXhrKYAqFJFGe4SQdZ8PcxHlUm2/jOtKHFqxkuF
Or/Nzcn0Q9T764o6nJhJ+92NocDFcGqCLWt9MTywoQu3/NC3Hed1YauM+/7SApUfbLeMEfUCGlwH
BX5b7TbAowM/P2tbJOT8zY6wYtYqOIQdKb3jTE/n2Lgvg+s74DeYNzkZj6AH7hjXSt3/iiKLFs6u
cFfY84b41AvUKDyJMiSz9WKPeVQbdyWhgWQbtaIzw/cHBjw++AKbVHHoP90pzXf1jkKXzjLsZc01
rVPh/olgu/tnZti5td/b6eYJYd/Q4jVtI683WWPfFYVd/EYHe8wwTxmYywsgAJSHBiOMeZri5xWt
UBG0qXb3gvKerC8++Svvtt1cH3/6M6BZJftzNCem+258J2sMGVXsJwK9QQFNDH0XlQ1wz4sHxh/5
GbFADXRyFyDf+6pBcqJgwp+QrJi17ItFz8o8yTfRpI2QJt9RP/Js0IstFMEJSkejv7bJura9B91c
ZO3+lzHMyG+zQo5vTwTt9gAaNIyYyQxqCukD4MUPlDRx6t2HQ45dIQ2HIeZrAVNgs20ixRfS5pK8
5ooBfSLyDWKI847DzHDJeWebTrHA7IuQiBnWxvsInPl8mC3QHx6C2U7Ka5w7OV4Cw+f1cUTL2Xsc
Vuq4Er0zZhbZbZQroPqTtftW/cZoBf9MFZSILU/9eHlKvFTTR/jPCHsc9R+k31d+hCghQcwimUrB
G5Wpbsnuxqtmk2SjUrVjBCaoCcq1H2SI763/l9kVgOMLQK/I0UGSyJsBtLqrNsXAMtfDKtnFxBuX
9QU58jdbfD5RslGbs6arcbt31kGkwOQ3tpThdmDa8sd8iinav6z853Z9AvGMYAX6bohi3I3uR53i
wOLJRmt8ackhUShu4CUBjOmOnL7qS9Leo6Khcv+LJgrOKD2uN2mtI3kaobVyMp2oEfvy7NEmjJHL
HVKpdD8fpW8pQpju99bVTEbZuVL2movrMWhu/os1LszHEXI7NE9knshoCPucSb80MfGt8PBZoHer
jdV9EBzunwDVDaGHZJqzmXApc46QYrJ7kQPm6vlALFLqqQhYWFfQ6+OXm5nfMn6BnnMbVLtlC7x1
cr+qQVlWf+toAh2ihoeofOeVCZ/MF3/0Y8p8fLXkmLmfaOveNl504diOXaOWC1a/6vATyhIZDdkU
rOHm/I3tkNm28R2sTt5cuayCmSMlSCH21VjINXVSQM8FR3WzuJ+ZE9RnKzw/BRb9x7u2qhhLiulU
AtUAH0F3C3JadahUe19xA/+g+f6KfPBIYDz64BX4lPW06cE+yiUUHGr2gerE8keYLQgfOwuSK9i3
5YsrWZXxfgZxaVKsrP0CVmnuhohMCth7wIyMRvXDxaZENeWfRlESJKNO8jcxsCyiwJSJvHY80tlU
bmAQsVVrID0SlwxPb/Nqd5i0pZAlmvdgHad/H8WLkxMvsl5DYuWNQnevUyE+drk96gk5/yc+Cnas
9D9ELynVTn0ZkV6KGe7hf0dgq4mhS0V5ED6hbxhrksMV7SSdaCMcQJalSWgvn4K//ywSdIx0cMQb
ZIXVS4HSx0rHcQDTp/53HpGLxmy+cwkt1r77xYSaKPiK0hrzOlQOubX47avl06ce1lyBPcVJcUKC
4/tJT7FcrXQBcKcEtIKpHi1H+EzDk5J0MWWcPSMJKg0/wdIoiJbmLvXTUASBkxcP9MZJm9N81J6z
miEygUuXVVJkMoQ79Vm9V1CRVerjdO+kcDjfLVEArpxFCqa+qRLnkqlKXi0Ueef3vHnfyVJNqx8J
ajIGtAU2vLmq34xpHOVxe+v+VA7qfOM+EDjQPM0gDxU8SrPREsxDP53dTnWmPb9LV7sn1G0u4Sm6
4ytpbbtqu/fB5d+EBREz3A+e59tAnSG+wqGymyJdsS2Ah9QkYUADn7R2zQfIuvcX4Oph9P+0+6HS
uKf73+loAzJQO017S/9ZnAuefDygqZ1Pt7AWrJxvdlaGKMEdZJrjmpBUMySVfCImwzCflqMNyTRe
JF/ZYXOoJBwPGxC/FpwDzzbUWXoxvLIycpFPu1lGqYY6P9fUFsXh2Wd1AQ4dkaavjKVV9XF8gd+t
Xky02+NtxHOHr5M9xiMSwlsqHi4G5WLYa9gxUYq4q6jdQgaecoX/auhyF0+nLzV2Mra0iVwDWi7w
sF5Jp2ZrSlhfIIrka1My7ANgYl5xA2czkX0x3oymmO9EYJYFOaUYThMWCrzi+QT+l5T9zHE03jNK
k18GFAaV7aD7/o9I+0G3HhvT8xJhOyRX9Sf24Lu9oFZ30Xg5XPs6Az9Y/RLZ8a7uAfNmEPEblhEO
lVPmC4/seOlHTsiBuvUXLAnSxyW5SD49x+7v4bwdUrh0CacH61GZc00oMFsyX8zFp+hbaEloaC2p
UgIfYRCKzbu8ZJNB64pBP4KOuA13E+pJLbGzxbMVh4+eui4EV3ViG4qVhyl30jQ5TGdv/8xCYRUe
dYuVXSPSwxR4VTTihAsj8wp0dtGBmOsPNTI75HD7/HAbjXSlE8Fu0GyZ0l67KChhLiXoYI677fSJ
7udrf3f8OYR7GiW4gAsA8fjTnPTx+JtF61UKiHZgJALts2BQwx5xfNY9upcS7CgdSYoUejlUQF01
NMOu2QIUK2iU1jk05P+Ruko5WQJfFWoWoJEgrBN63stwvtREh7+UsUWJfSxNm2RTDwmMHfsbNcQq
QDHxqfug5jPBminE4fgE0lAcjfYIdGTRDDuUwT6hp9XxzygkMmy60u6R5EnjMOi67G1fwYGv91eP
ag6QYZa8MXmTD+97aGpppymcK5gdtTjzuTctX/JziJ4c3oIk7aPHQAh59jKqqH7ZUSSkgWP/aaq3
T/ZSlOFVUlt5tBChgal4d207o/ntHoZ06hxhQGheckb+zypZCRjGsWJlQsO7m0QE4WQOil4X5oaA
KHEcZSQ1d9m9TDcgEAYPjqBIuquvOFWj3iwrIIdfd9I14sds3sPpF0wkBclzYMBwOy5tAzkNWzlI
tB2l2GQZ06/8JuA4i7A67Gf8XEs+NohNqq+WC8Swo/rPu8PA7QUFkFWJbIPdkASnYTnSkW+4qrsx
h7qYwzOv4+zULCubojDs3E1ZFBskNs0elUNcZpVen69JfKvJ8ny3ZBoGcCiuMM+C8q7M9kRwbNQb
XcsJCpwyYU/FEkvDEcvyTR2/kkNpcqRz4EXlPt69ClayN6a8AE1bz5983wsjDwp2mSeT789U17u9
/jWfUg3xNBkfrsFvrIDcItYpS7h3StsIiw/e2bpBHPPwIq65xaRJ/zqMzlBKRWXr/rkMMnAex4tp
p4STXsoAFN8wqk4cLEUK1igeMb7allU+5HOzgFu6NagW/Ns2fWdSSH9BqKK3ws/QUZXe2ufEXBpe
mVVK6aNjzAsB2GX02PZK/uCKRsRxtlxtgYAdAdZnjRjxoGM1K1uDWxBJ9U1whl9LNOm0otZC3yBT
bKjC29T/T5xaWQr9g5USQCeadFMA8TfL+thi9OiooNTS/w+86wXUlSQb/B9hQf45NqlJJF+XWsw+
vSsJH9EfQoDGhAilBsnT0SdkB2Vm0v+kRqiafLPzIkYfXYuHW67lxlRAu1ZUgMi2pLEzWjJ+pW59
P/5dfU82ZccEcETPpY9XmVXPT0LYIN1oRKYwKHrPEygFAU8s8lv9tMTfGgSFCjlLY/H8H5bhN5Tq
8tCzKBpo147Z+8WWpq5akTpElAqTfxWlfAkCyyP1uv8y3hy1WXTOYT9eg1Ew1MPbWQEUkL2e6/KH
mmSCSQLONkakj3lwlZ0b3Yg0Xr06RDX3IbkaA4Q2VpSkF9cBQFrUVtInyiyyLmhd39ZHSFM9KZOR
3+RDk82NX2Oqw4b29sdVRTu1vqI3VkJfBDssrYILoNF9Zm7Gjp+Y6KmvnCV8eNpRNYFNIfksurej
gG/3KxCHrq1rBRRsJ2FjuQzKUudVZE+dWEW0CMdf124nKkq91YZ+K+hDpS9NC5zoLHjs1fvNr80g
5/eXOcbO5PWgHkFlzFwphWoATytj+nEX6WR9631U1JiLuZNwtjcs/7Rv/Ue8iqtETJ701jQaKB0t
mfTbH0vdiu62uJJ4GakYiBXKuHj1RsjHc35XjJQt7SS2AGMK7OTkQMwd4yD9VAWTcwbWsM3ExqOC
YOvmcqiq9UXW1DIFT7atjWNg+TZU9Awi1aoHngzcSZfX8b45S5RV+Rnu1cK/h093sWHlCToxF+xQ
+GdhYQeldXRi7ez7hSzXy0S6DGimgdJbrYayyO7ehT61VhLLkxcI5RFkFL2ZXHrJ1XaQj/LwaviT
w5/CbrZmLkBvcXRWDJTetL0t5jOFKBBdxWnGJgj16+xM6yB0s7/HASw2Ctqecvs0q0o1wXW3J7hb
d0RuSNClFzErUtmtFUDwfog6w9wDeiVWA8FALi9bFDLBlSCAaNG7N9Tmj1Ciu3auVuj/n2M9E80W
n7/9is2BuFmCna5rq+cdapKtCwjfaB6PR/vbnM3/3aYefOgBedimbuEZx8OdOplWsarsL0xE46J+
b8AcLHOxBdpJG/7iZZFKrY/uB0z0OBJFuLDcHNHiPK61Hbm/rCTWgjLiki4bKp0w87+i0dFCTJvd
GGgadMD2t0PNYQe7dCBPWz3PkWCL2AFiPDAX4IpkK9jjBK2bSYe75HFdXQV77uEsMjMD73OhGCTH
S/BfobB+sLIvj1b87TT3n0pBGjBw9z1o0jUw6uXZBFJmu5L7BCTk7ez3CerxgIweUAaEkcucTgq0
S6HdP+S84EePUG2b2ndFkeqovzgkO9Wojzod+PcWjGgcm3PV7w2wyYmHHMgRv1ZYpYy78JRsa7NQ
wF3MeL1NsifqrkLeCM3n3Al/O7cyi53Rx/C67wAszMW9zsQoMema+x+tIuaSEQD+hO3ezZgvw1mr
jE2nSryoLSkjEHy4BL4FxEFh0VQM3eprXQR5aZ2IUloYxZU54oK9XbFw/374YZN4/yLLAhy9/xPs
dsjODvtZpM0s4DCl4h9CPVOxsVV8H7q9wpmCsp0iX4cHm7aUUdV3tANme7i3AT4nmNIVMc//+tNa
zMayL5X37TZf0ndFV5YOWxTXkJxCsXPH8NcwSjnrf2QR1xaFlW66CWWAIGMvhG9Sed9V/s/ofxLe
c5GfT2+RsmODh159nBi4Rc9x4RW+FgHknFUWPOLDLxor9c6wux97cQsLDXhCTnUTBNtNlPdHG7Sw
Ag+2uzuWZdh4TdNuGGuh33D8kKsoxIdsjF/kWovIE39HG8DQm45MRLpoePtKJ8GWyEsx3lCm2KuH
NilyB4E06ypT6oKWG0D31aIx51EWNRtQ7PvONcwZGmWPrix1fYu00ajT0RmT9WM9FP4/vds+Yc8j
Gxb5dh3TqQ1qhihXmBYyyAhvaagq9TcjPWvrDg8cLA2MV1i8tbgDj4A++9XuLTVf180fYPs7TZsU
sXQoyCNUdEqRFUejxGNOVbEEX4c0tDTCKUtIvh9Lq981zTv6xR76YtKDxXLRoQVVyL2JW4I9sQW3
8H1Huf0cNJHuGI+mK5I662TwTjeYa3V2Dnes/VCCvPzD8h8r3sBqBTBFdFf/vVG/ZBWSuj323PmN
URS2cfzPKTuwIO//xyrP1lxGktglyjrUnJSLFPTG7dc37izArCJOZJzjg2GMMsxuldgELHZU+yKq
kbtzlC5Rz/PVFTr4F85wpdG/x2TFB9NtthgXEX7B7YZUFSEf8ZSXwmTXWpEL21U6VyESNqwAW3hZ
QhkKQR6ET5m07zqfg4csVWM95BNGIRtNWJS43gxLZSkOR2Q+5QiJ94f67bXBSotlURAFqfPMRDJ2
K62gePgoUn4YccCJrIYuxJFbE3osbKIL33xTImcxPLgQG8A1KKr7jvO3bOlvhQ8A5xMu4luRefsO
VjejjQlbRHZCoV4DmZRvu2o8UpQlfHU0Fw1z9kc4sT4Kbb3luCnPdGJCBkU3M3N4Vwoza5sDIVE8
WqMMJ8mVoHEAHH5+Pp72zeh+/duXybX8dT8dT8sYRqo7dHTNM7sIuSF01CtWnwBiE2DsLjKJ0d1C
esx6HbGlefZb6lLh1OYBaX8tcgWULX2a4oWxMOdhJMqmD+buEwiSHV54nKGtm4cQya6vt7Q3SXla
YP4QN+3+b3ul2OyvZRGc1+CHcTiGzDjTrDtkRG2kOCo+mBokA6GxLtkTLIP6oSvv0ZGBDPSZHuUN
ha3iqvtXo7pMXc09r/ls1azQHM3bWEz/Yc5glIMvuGlAUBittaBoWDN2aXo8vUgbmWmLmaeibxDm
k/iAP3dxcqLeVIFH4LQFjpKhY/zYRd7tec7iEui/DeebtUya0+McaoPm2+z+Ax7mqwpg3Yo++DGq
vdUYimJslGjESH26md7XrRAut9s5jgb0zTPvyhEVsUyfH6lfT24/h5829q27R3T2Y+2OnakSEkJl
2hncpxf22rU/fuhAp5wcYsQJHAoEzfJUyj7IrkKCo1ZzzknpO3nYrEKyfqs2ZGVssdLGT6x5713+
OXR+u3hnnLyVX5Y0iegboCCdSL6o9Q2zSUL1BZ8M0+fPLdz/+w45UvrvVUOadF6zD3aXJtjF50Bc
x5fELhg8FMekL+oJurZlsfruPw2xvkhXQdd8C+cPsMHuhtAJtlgircDl6l9OOBfaqQSYYsV+Q5OR
y7KDSq1q9nS16fdDS5qkxvB7UhSJEVdgT6sAHTgbYK/Xr6oTOxf5K1tgsB3X+PrpKILCy3puWJAd
va0HO8RwFzwSyxniSwla4gsOA6+Ce8qPu+/9NxFvm8lC3Narld+hcolTGB8inVpE7iYzyH/kJN4U
jH8s2qoeDupmFW4gPnyNAvs1rAe51fZRN5KgiP5EAKQstwcmbhzMVvJXhpExM5SwNk+Hnp2LIxOm
tuCSqHoLeD4V9dXLZpboJk2AcqTXYMbhxiNFPF1JYfqyYAEWEA1AZy4SaG3ucqwtbgFcAIz5u6C6
3T7P/qQvVxizse3/XF53Y+9TakgWIGzmAwP467/znYJrcs9MvJCbAaxmcQNmWNQmBFbPw2BJjdGQ
InN0nB465iKG7DIuJsaMPVSysSYm3nnxTzId/NFjYcXDUU/3uAqa13/xvnne2Fc8iM+zN6dSYySU
pZbJ/plgwEClktq0L1YDgbrzq8rKlPy/tlO8nJdI+kg57GeuOxV5+5mXZUCrWZRYx0GTs9wVKu7P
mxlvOy4od5RM3eBqBKTfCuYxujIg5e72EyxGlSVP63QddUNks2faUSKHvNAjYMnKxXVG3VUyWLtI
iL5nXwtXNji5QHiqV7hW83garxZaKZKrG+B8UjezbnyxIq74cBNcg9yjqoCfK96QsRKxDW8R/0Ms
Jvyx4yxCQjz3SS0BB4vDJltO1yq65iGuUR46Gvr0JZPIUr2qoRMj5vf7fsp6j6E+gVesd8viNTMr
w0MhjNjQYdhguE5/gS7BY6WYLrx9gxWjIno/CotOEVPsodC1bbX3qX0Ow8N7EqBLo3+h36sPK5jD
lYkl++75VCqlO47tSiacTaWdL+PzDeSVT0yuod2s5rv6B+2kCWTUtYRtrHLm5AmiJuNgp9P7+Cs1
MuzVlQFYrP6miwCjnqwklKEc4zjSns2u3YWNkIN/0Iw+QxQPrDaHeYIis58Atba8Br5chCbzEG0U
nG0MAXU0SrAFSNDVOO7vJjwWlmjbIvxqv36pfXwo1UROC1gTkww1GugW5Y1pkEG/WwLarBBTCJ6g
gN9ca1OnQpSxiowI5oTxNQ81pWSohoSsjnxmXgjM7oZwD+wbOJL0hAe2u00cmB0M+w9dfjqz0woW
u+axb/+mzx7WF4pSsGCR5P7rKhM6Z0ClLhr+T3v9TqUZDWQrY1H8DBYfxNoZTa1XFL2KkvmekXwp
fVC5g82dbG7DzoFTa1Bl3HFGwcXDE+bibMallt9qJsivjIVzecjr+UpuT4E8c0maVgwC5cULjS3q
BQXs9G19+jGVA+DuHHwJPjkkEllNUt0DIUZJLA3rsRZTFKuHAfLFHGnlro0omjxpSeQXS8YMqhRJ
ENv69LlHChOSRoDaqtOJSq4l7eZxr1jwhKZWI7xs05+NzqV/Uvqa8OhSZR1EwHUUntxek8Q657ve
0r7iVTy8cuJEA1WS+chh09n5Dm03elpkzZ35X0sxafTkIqP6l1OOwZ9WrO3t1iiMISK6Fp0t6dZ+
ppKuVhUqe38tTw0vDR+L2Y8JbrwMhYo3VIdSAPrHvZNsOhjg+6mr0xqmAsqMcjeRz4xYJ5+cM69x
SPbQcAQafASuJNfRdK5VvVlYehqWtMjigbSuNqrZpO571C07POtPom3frwsSR6H0b2qWxld2YaIt
IFhW7slOqRGmqP5NCiKXdC8+xHo4lNrMqVA9MgviNG4r8LszvMVIEEuffo2mhs490+3fa8oT+68S
B/6VB1bS8jKkOAfswqhLTzdQUbCpw8wQEyPlggwJSzEZDBUvn/s1KC59YAs35XNCzjM1b87meJr8
HkISHW9qTsCUpotyK6nouK3zeO7S4mDNhL7A4oP9iT6oFW9lY7t0u4cHHdwccze7qIVq0H1aTwvj
jaBSuGnDwVcYHihnm1PvTyhVh8qMH/JTtyNMuK6pZla3XUWixlsxnkLOnTFFuPservVH8Qm5LNaX
mj4od7AhHlIYTK2DUWoJ3TR2YiUoOiXplcCiS44THPQjy6xIvF9FuapZ60btXsLEDcSyUHg9Lz2Z
AqY7OrKCvgxArST/KkhFBFkmgjaoPYmnW0kirgnb29JrZRfGpyxpTEfQrwcJDxYgSftDVY7zVs2b
5AE7pgGieRRYbULnzhDh51l2V7NGir1Avh9BVdNJMjxab+HggBXV4H4qtd+ibWF0+PcP816dTPRH
2Le5ALWpjPJM+Z2w2eT7BTgG7gv5F3v1TBsVbJGKwytqBhDrXOXVZjbAtltxwBLRyytpz2a8s187
WyPawjiHg69eiWrf1ObaPZ63GmX489r1/edxoeUd1bRjI2hzv/NGGNwJyBuEssMb+wEs9ayx5uxp
ww4SHiEx5sC6HeJS1du2x6lt2w7PPPmUvGGMimZyl1vpdnlxXQtODw1n96KHLChZIJ2YulHiHhTh
KD0xXrHqE6q/qd4err74EeHURucsS/3d1K8ONN5PLRjr5EKs6iT67zGLHrGnfcJ82wnCKh8DKf2h
OCfnmG6m8YOOpkIELvpJNvzJH6gqmZPFnYGaUJ10rP8vgUQ2ONWLwN7hJQn5seQ8A6aEXganb99H
iETWeK8f+FGhSnPht0ziw4yugDqLUPwZP6qsgGlNBNEPMSUiSb4mDprQ+PPWca85tcCd5qJgAELt
bagKeDVykormGyel4fuvT18l2pGNPxU12PIHBX0raFiPrIz7vLVrpbrUAhM05pYYltjhm18LyyHU
Kcd08kQ2P13cBXJxYq2SYHCMMxfWyBoPJbOdbTzehzqf8iGiUG8dhlzsUXaitpFkx6z4Q7jMzSSP
KCgKvgphG2GLQ4NA7Np3rKrBplxmxTEEmCnhuiCawJAgNy3t7IiuTPHMqc8mc5LLXSpIFzKWv3XW
6i/5x80hn2DXJBZeRGApDlPikxtiyuE5usHsXX3XTQxo6tFOeNgnMJ2IWVl42j5dldwMS9woVtRb
zAZ96l781jSiI0+n9cNWDnsGlTJEOLkehQHkyF9paqKKcRyf4l6iX2MZqvb6BmeMPlQyg9qw+IWB
Efgd/jYuVq7nkFKawjP99l/BqSQpvEvTwZMBja48dI94DQKK8Kz1W/ekbDxKyG36/Lsn/iZGFkPK
UnWiM3Fe/L94GLJvTxrL9c+F0LR+yp0uNW8lW6ORArqN5gBuTS6n6XhGLtcyX+iJmhAhxw8R1iJ1
varY1nZLII/Q2I8HgmDTYksDAOVRaHA6PDwiM9tVwuEFM6rcpOu8yby62GOSrOKHm+tVKsYSHNfZ
LTsmGCbQmhvnsnGQhAMGn8WFFQw0PR1fj1VFKtbZzJd0Tonuxjv8KGzFN0BlC1KMMAZEhuQ5ytaX
ViTTdBlmUdSoTOf0IGUvNe+vTiXl4h4ZrQ8hioFj/HL6hMqj87hHzWvsORDgGQy5K7bVzeGcxj0r
OWuRv82qeOzXOBqdeDaeV6FrKCwN5Hq+Nn63THEGOxB6/MXxY+nLJlcGMo4mFK5i+gkxYzfJzv6R
Psx11lFFNdjnMKYAnXzAHcQ9N0a+MnsI5xFrYeaL8o18sWsGCN5i/0hILJUxWvBBdHpxCDwZEt01
fjLUClkCgnq3DERyvtQuuXYZwfZu6kV2vqR8HttAoCJD9C7Q9/uO4A0Ha1X5BeeWTXXKy7JRCQBH
MkNWiIzYcfVS1uMi9e9BP3p+v347d47U7S/jviRVxhlQ5Iu8AzjHaNII42SVYlgUbw/X30g0LmsZ
Dy6zAaXzqMp8oLBKSTrvZFajZAak2iD1d45w/WcSUFUUQfQw87pcnKgY+iHkFV283kksNmsDubXt
yO3umGaHxwgmbetwYB/MP6Ln28ND37S13UR+eJlqwwpzMANoTdgqd5w4Uefmt2EiZ8lLewN51FRn
IW+V6tdj+Bm+qhaCf+zjLPsyenID0K2mCzaS1g10WiFppAPK8QQ3pxtSu9XsmAvwikJhnDxjHykH
DNA1dAg7GruiiwoR6Jibo6xn71zUWHZKorIKSQRqA5nTRf7o04S4UO37rNGDBIUprf4zaA4ilvVl
jVj+X3wHBWK4oAHHEVqLhAfBvVN/so03gVHp7xfnCBqlVLWRxwf/5h3jGaP7u7gwkpiTvCpBuOI8
XrG4+n9RDt0sk3dFiqEkjPSrdtla1AkHIEJgMNAkqElLgqcyNgZXw2Znr9y/yBM934LxvcwCU83r
r/QUA7lqh4Ie1DEF1EvmGFZQLES/tqzokC8wnHtDR8ym3zwW15dni5coekdPa/O1iWkr/QBEf2tD
AWSxtU6n9zivk8FikRzkB/RGSjnlyCwRzddEaWD+3lwBZn/QyreTJuHDmNN9y5UDIno3SBpRoKys
DCCBRVEohxflrC5j8abvDS6AaI+KIcHZqzkvTHt0KjL+baZMeWyxFy3z5CkhgMqp2tjgHSW+cWSx
a1S5UFBNED7EgES7jAqiVkjP79Ps2CeJcD9HYrRGrJs7KQqQ7E0XXS49C9Uq3rw9Lm8mMV5oHVv0
79Moe96CDQ8AqTLwcWHCpjNk/p9zVqOBChSChIJm2bKMORGx1ituP0+EVPqOdTpTq6+bxxSD+C9v
JuLu3Qgb7b9r0+8DllvhjNBRecC8ELzExPK6qCjIMpuMMcUiw26wONSh0RST2y5jqbCKKKIzUNN2
kEQZK6hAH6Ds+66uy4IKa9Aa9stYbkaYFLspkusO/MATfj6WOpXU7dUQKfL0rCUIH+CaIyghKLNE
XS8Ygnjqew2G8rHqHlEEmJR/VnOUNNdBgu+dH39lcSeNWieZhZF69go3yadbke2GTjnH3W89LDVY
yDJ7xj+9lYbAOdJfdOUkQx+hC/0ly0IWJGZ/Z1gqJaNSAm/XqKlVPSWG0oCyDoVG4W25KoDfZsyx
F5h0G7nJor1r/KhxtH6rG3JzG0p5P/urotKeDAUUiQW2yU/EWqIxQUUJjPJcyqsKqutbPR908g/X
SC4gJRTSFakpPkx8CLoXjICT+xfXmx1jU8JtlhMaCpgwWcu0r7cYq7F8MrlXRruyPPF3EYi5x4q2
9M59Dl0lXXqjR0/2sFV9sqXVj24CpkXvBtsI/FFgC7UK8aFUHkHFxZNaTkShhC6R51t1/HnobBC3
JJK6656UFDfXSDaXMi47Bx2VFawjGkRBcW6oduy2zCQnO3a+0RfsG406KZbbDFLktgO36OhA8r9r
ODg3H3RBNp9ygSElqrBnR0e2bxQYWkmCClRd3VRbkggtQte+83BAf7sKfWFbT9vTSq4HySDkBOjx
bovdjq98tbwY1n3y4l4KHCXHwPuPeXZka0JC+ZQcmnVDr391LXZ/JMM6jphkvINj9EYxMrLwVcdQ
jd0xT4jFQOuqvgiJ1olczhv0tx0FjHsUKoZXZLegcyMT+SAXjPPEUcSpDH+GBsCMjOaluvPSlC3T
8tbHgmchqjD9+XjgoztFwycptMMnhN/zmS8xEjQ+kXy+zsLKtJDwmsjbtS7ByWV51zhQp3bggIbX
iwAWINNjGBCR8S3P+msnzGouA9HNzewqwKpSOxQgQUgGgFxYxdunMIHZjRJfmCnbvhck9daCQhcR
CEg7jdUw0kheDDQVfGcCYfLrYqfVA0xNFjA79yzXB+sqmMS6MhDp2466zPa4kY4PUcOMZrJ5Uhic
nDG+usRqsZ7uZ0DuFhsQ80QyIvAzDsh3uDbRFMeMe4chaW9DP6rWJmxg8Oom75CGOMqlKEbY8Peh
HWP/7zzjqxUQgOr+zriDMgK7ZWEucdIYT2Ys+RTZjqwnjN3lz+7FM4aI/y1US5valzhYgrTxfvju
i7TkhB5FlBRGCktrCozVkS1GW1zqtzfqS+hRo1HK9LDl3ZWR2HHOKs5Sh09pnD+uSG8U21zZ3DFK
tiJX7jXJBaPDAgjm6vfflNt+9BmkDvMsEupKGDn77Mw1I+Odv0BturKseYyFsT0elYn0jNVwkFFl
A5Mx956z+jfCRTq56aKRj7rNFc4YOslSLmc4EzwGqiDd0WQqrOrd9HaZL6Pm38A+0NxooaV96C4+
HQbKSth8gGG+BwOU5rZShCP/G7lbmWnHcON1h5ooyat4WYaLtrpiwQdx1y1G2n73wH2NPNRsZZB6
J7F3WmnCXrTeAbJL67owWMd/mfQ6kVZ2T36m3TRG19WkEF4QdUFBy2l79WBFkhjfuQpKNGItBdy+
vJ1puImYoMbMGScf+5AyjV27RxrqCNNzP7HE7Xncs+GiSQHwWQG+pB/OLgz4rIzTz2+LRI56Xk1V
1xpO+EQUX/8EImp0dhdJ9mGMb4xsdopjxxggK2jyksDr285LATh2ZxVRTAEh/qaBZ5lMusVqBtD9
WY/tspJNgEq+4g200IE4HsIpkpa8IrNCshz8AFb8nwJmtweE6hUmuXLjr74c4icbx9+Kn51QV7XA
teCR46O8bFNIrNMmfpXPlseUVlgRzqWiQ4+CMoHNsdNZqfP3lQD8RLUh6bwOuOXHNVmqq7gSUBAV
zt817gU6UTmJRoq+v7hx/TPhU8RqFg9HDi4mKYrCBk/qouFrCaWYl3u46ttMBv0u9ucjKjwWvu9r
zlMD9CE+HZxWtp41RtZFcxYTsLY0rCbAm1agPPm3VcdjATQIYJdNxULiGLcZAcRI7A9/cEqjWMW0
Sg3Tm0s4GE9aRjYR9cB9gvGnVKXAhyUAAMOezGQRlxIE8VX+02Pky72EFjJrR1ZJz4EWI7u+9GT2
Eot3ouTHNWLN7qYyH4YFQ1qP54ECp4zxizJXN1baYcEKlVPaoQRCWCrV62xXQa2esS/yq0W5Cr8w
C9zBBQwnnnorikX5fgK2JtK21jcTaCIj0ywPSxNw4PIThnYuyyG12P+ozKOPVVpCDDH+6T2+B8Wf
v+3zBXFRWReBFd2GbNuZewZH7WZ4JHJqcWYey9LWlOW9lI4lwDIvaVfU8PwgqwbToHaGm7vOldlA
B+X436r/EH8ScobFledv4RImZjt9kq9NjAkq7aEBkaMnh4I7JeXEyJN2DwQVRRsxBdconY7XspKG
nDp4m79vSTfXGrcyDfVfM6ql3DEkTmiDNvwvLefeGa5+Ov4LF+bd1P3ha3sgDK3Id0K6wCdYBO8A
imK5KTz7c3UZFqMKZv57Z/NxjjG1pKi5nLXZQU4vAniuHAyrcAwpwj8+jueD56+F/1pRIrkM0Tww
bpi3ImarsHnRQYZ8OEyDXP4BhbEBqkjK+VQ+doymeXcfbT+mm9s8mkQMVc3MElVSWLda4ARXAla4
FjwL8C/wMZJaSTA2HCMCnBSrLH4A+sRX9IIo8eNVpdAd1SrKUk7Sxiffcv1Nj+u0FFAT09GmmQ7k
JyQOiAuUdw+5l1ucPZQcmfNx6TZE1RxpA+4fX0iYskMONaL8jmhastXYBNmF0CPbj1oxkwReoyfk
l7s0hqFNb9ImWa00wAuhEG7PEALYnMWBqz8g45I/j9fCH4ZgOV1ZxlDxDYoPp0O4lozxVltddSFq
qgTNLrAIV1Xm6+NpTpguDMPRK7ZbXTatnpqJUFXTgjSOwdcuG9jV/DpkKHiaawRLzCH8tJzniFEN
WTv8Esr0Fwcg+xms2DJcWhquUnZ4F6JL//yLBVOusIsNtiihclagjw5psk57YH3vpla5h0loSzUe
B95U+6lTPtUJg4XFoktdEBW+NV2J7gAmHmtaD+ZtGd3dNr/G4hkCZhM30+/BBWR6LXfZRn4LJHsj
ob5drBZ7CE9ek5KjCFfrf3ylCvrNYOyUPMnfgdf5zOpHCqatRZ8aPW6JT0qk5NdkKXeo3DfV/ZTm
uDoWzG8B1aXnGL23mv6M8lepKmQ9qkFgJvXnV/KyhJ1uSmygpZjUMF8nMnV7UAas8t+h6xDZaBri
BvnJsrRBuJ6ytFAbRf37mZ6A6fQ/ZKvT/nEYNo8CoQbcwTlfZ2dpwM5CieOCI69fB52bFx0VpFaU
C8B6kQZejAtzItKm7LTCtZqelIbNkImt1/pEpc1iucJJ4f1Ayr0H2u4M2406qn+/Ug2ezWJhR6sQ
zeqBKVjn+sh3MEDH82sU4W0LGfIHNG0YIhbCiwiVcirSBFePv6HsyWjIF5mpDAZQm3P4aVkdKiHZ
D43IW+q+Lyxdgl9voNDgO1w75bjCTmTsRew30Uq47sES+4hdT4Ft5Jko5T1W1KwCxYZiefHD1Hy2
ev3Gu+FCWnNNwW/V2XEAe5ihwvdXsjur8dL+AagV6vn/zG9vZSO1/Tooj1+PAGoqehUkUioGlAbG
NClF5zK3eJAgqvxt+t5OFE0v0NUUBXpWZuzUG1z+9aTOkKWUIkZ2yV8IWQXy8jw/fXUTUw8q0Yyi
L6TGmTt9IQwceIVbJqFT0wNADo+efWmEkhQODXg3RKGBNFKxtab24ob+8MBzN+x3sad67zaU0Qsp
S2qP4v1xDfmYK/e8V159FolmuNQNhsbdz+CmDD/qeeIpb9kuWwmW7FzY/LqMbO4WMFKikHkBGS6T
upJrIY6rc7laqYLyBBHtLRtiPZq12pSUDcg6x40JsRN1FW8NehwjA0FI38Z+JwebQcL0FdcPrFuZ
+VTuSGup+IT+7IIqbKFfUv3I2JCS753xBLnHbhQj/UNspuNvyn9f6OGsSCn/Ic9t3rBWBlw9K494
3OoW+hH8CpikJMYElRvFv7H1hi6lZwAHrJEJF7HuUNAYpuKOW1Ed+604VkFZs0n5JY/GMvbpj4k0
QLUOwQyc5slFLgAzc/B1+icrKdDTsJVCk2nHPNhxegqiA2n24W2uDXwrx+lDLmPa3UX5enp6AJF4
jwdKxWK08OgpvbCnH+JwQ2gw0xfBdTJv7m6skOItt/TExGqQmLf8Ds6o6ZzA5Ib73j9UJpw4ErzF
vxvOeeKpXkvVZla1ia+pTyJng9pUcvEAQnvTTWkQQOwyy0sMkBdAobb5Dv/Z55SU1paxN0evkvE+
KzacK6dqYfMgsot5/OaLJpwbi+pqHQa2jfgQuyPjJk33PiyT5FqhQ4rMu4dQwlvnkwAv0j7wRf7U
ESwi/NMLm8rkwU5+koPJkdQKiH0ZqY7HClrjMI/NY7U+QWjbCPW7wdWhvpPTHuLo7Pnuu5ClmyTZ
ba6F+3rE0UfXlC/SDx2V1JLOhnSFr8kWs871jLvRIp2gXCeLEuOGOr8Zk0NYlN2PAswPPDH4cDFo
AVvnnzdlUl7UzTDeeVXCU35iDuJYBgl3VzvHAfTnOcNqdTctIxSFUS8FpvPW9EegCVqkf3OZ4e5r
qSm/ox4/sA2Bc4fcn2ed52Z9PgSaA3xEIC4NZOm0YvIHZo18NoZomp6J9RtwljCNwovvzrP+pcle
a7aCe7rBl7yU/n1efdRwoWFc3nSerqxCNNb1SoMAXAPOmGygY58othJDI4Q4/UvFbOhVu5wUNnhf
lgWRiv58mpooZz6Tzmi+rmrPsOUXl5f4VwmPDNoMrMMKF5RgQUxa6N+f+0sFBSV9eKUmOXD9RCJ9
pZLV9bCREoL4esEs3BWhnxE8NVtH5pGg4tXPiovhx/Ln6LYNshhU0LOrMBlp8CLudL3jS/yVFtAR
TgiMGYMeTkLZaJzDCa2k87vXZo5w6SK0UHzNUzARfgDK3KO8RECCqnpIes8QZDoC4DS9bdVRot71
Fv+SrD57JpVKy2Dz7znZzlnkMt+OUgVfB/yBbfYG38p3QinwEBM1Bn127XkXpPqu1sFbpI5S3g++
5cuE3uFSKZr+ybvDW07thr4As6BYSEhHukBeBT06kjkXzQW7yqElLtkF+VrazXz5sFRdWMb+357T
rOM1YroeDfHuG6zD1FacMukmdJILbCM1Fu7m3uRpX5yP8xS3dlC4jFZVRxCBNGIlPibPvG1ahQfO
RPgpVxSBMTK+wrJBmIZvrv69n29bweShOczS+mdFQpNIdUafKWZgMQwM9wFSTqNFcy9x9Y0EVfQB
FO+Msr3LctWNWhCenUnLb4GWFUUsG7MspjA/FBBDo5ycm2Yqt1ZuNVzaWpsA75pI+1ikuwpYty6M
UCQ4DrqHM1nz4xwQ1602dhtAS0Eth2f+xxHwaiCsBHyodhFIrDQjvqxWbAuZa0zApyFMUBGdGjRM
RjToPieCJIlaXDnAp3S4IoLbgbgM+pYo7j/Mq8SWOyMzHyg0/hcUTb4IQLsM6dLh/m0ztdrX0rSe
ojc1ndST4lmgzyMJR/5EqVB8F5D7zqLFaWlL1TbrhWtTkNSrVpRbHSPEIi8ppOOFqMCnYXyz2okD
yT2ejbgPX4rT2g9VzhrQ7VBNzUMCWHbp4HNHdGX7u2Ol/3dT5zHpCe4Rn+Es0JuHe7J6dtMIvqWI
RDHqyZE8LDMNk4msuLd8niRyC2r04uDt2N1nFBCX3kSCSzHKpl5WhcpprJve7XNONDw8NIc2YxNc
IzDJk/FvSUJEEFiZ1DdZHFGG3m2cAhxwakFJJrVuuHlTVy4Pmn+QGtXFYdShk8PUFhBppWiQqAxM
MXtxTPtMjZ5sq9XQ8vVRmnxZQPnGUDJ8oLHgEpjA9b9UgWNUyuYSTpPeN7VAn/IVRXyHDYUyk0eR
5NOjoPqD6Dgkq2K9qKYn/Pg22zIFfzNPLnPUDLY68DWBfeblCdx9AtcrJGjZxCd8HQzYBZVXf6Gb
9NccGCRR7O8LZBo4mnvTkN+9r/zT7Mp1/93padver1qbYojtUUTj/n2JyvNbXm45N7IquH14s49d
eCWr3nG8xbVT1HKEePFAdZBww0ZcJtbkNzvj58to5oc1MTrxprK+L/czF/khjihOAEUPsGRfyUTc
SmB38GBJaW+OAoWRq0R+hZC3WmOkO/laiNfTby4LrELYBt/SIRDvXlWJLILjr8PEmRVm8jHEE2hD
h5M0LNItGSyqKjZvIGH0gykhCv0gDLH6Xa/uBhB11UzOJINJZp2YEIXYXexBtn0LSDn/tOaE3xyT
KAkdi8G7sAAZtfVZuTnBa8exq49xOh9XbQdmZ3XrM7ek6DjhuHhn/A9wcpi1WX/gaw0dF/kkCAOT
LKozZ+BuHdmfurtAbc23DesRYFBeiibKlFZe1KOBste8ZDrtQ3ksDEjQWDxl6EDVw1XWqNEVegul
D8xPQL0mnHDOeOADfp+gKn+vpMk5A8K//aMpEN9Y0kzCn7m6iGBeuq+zBr1WBrEQYjIpwbYWKp3O
UALhBLQ8MZHR0LQB5hT0yUR0J42I7tRk+K8tWaDtEeKNlFAy35G9L1IaVm3f90oZG86zaDsn5oPz
aUJhuRj+7HoSsMm6e2YKj7hkRQxyvJgBWXUIVXwiL0vsOpwACAhMQmsAbQ6XzUHrnSJBQQCneDZ/
X00sYtWufVklr/xIePTs0+lf3fNOD1SW7DKJDjvHz5v+kdNIMgOjVcIm8MsiUlYyYekmGJAqz8pE
wIlrR+0yiWjj4HcCh9y/S+kXqaN77WxC2VaFHBDj2i7yZ24/3k7MY74IBvDYywmw92q4AXwYMH3k
zi6HwPczQ1I6aH4dzWh4zs66c9nvdEmfNdsA2zauy0v/zhZNMrrXjTYgIoFok9cEF0XBQ4/VpkFV
xslIDfN4jjMtoFriivJ/c7aV9MTcKDIkWs/5SQNjFSGV8a8IRrfVimBs8z/ukaqAFYSgFKaVFEuY
GCz4pCqbZtkF1iGZqlc2qfp7RmrGc3KIP8BYaZZSvs2yI0XHJsOB2jT3Jysqfj2rTeoejRpacuWv
Tz5eY4+XFQnOe6xKzDZa1pDWjG/I5NiPY3nWMB2DGyjVS/nMW59D2P+O9qJYqQauMXFMYfEAN5El
zlEsnC9deGC0bpk2ukyNoWUVJE5qR+qrWoqD9e98OPfrvdnPxbeZ1kGC065RFlV4/0tuWIMgsMAO
cKL3chu2KQT9aKUHT62I8aaDj9XD8u2azELF8A79Wy2gIUrf493MoueKUdgrB+d2EKG8udI0BfNJ
MXioPMsXnC3MsYV/dsWxUnTzFjm3XTDq2utSq2f62xEb0Z8sY0zp/18a7KKIUrpJMqORJKrfaoaW
C47VwkGl6Pk5KRekiEg6vv7sk5ctAhMMiPg4A7l8HcErgb1ZEOTIiDJX0CjrvrCVH5kxaui2qx74
lEUgK9Ws3qsFFXmEP/1HTC44CezBmzwdbcN7O1ms5oz/MDclH56RJiNCi2W3fzx3gslaCabKqw4d
CadCejV8gKWy8PnDOpYvhSAshpl+wWIMSezNWt7WmMueIleY3eaj2JE68KR5WDnXd4XNwHBGC+nJ
8hjgYcKFG3d1Oj1Oc9pTwd2HMvpQleZFNs0iTvO8vPKo+FOWU1OmcCLVn68Ne0xGWTFF4BZqGF5O
AXUbpUc8OhEKtsTa/mDDxMH08bUEVxCFlI3NPDmi1/b3dyvxIhjR3HeCQuVRNUXPu2gRoMBODNGn
WfKvoENsmah8FJXHHdqjLr38eVSDoAAVFVJgCH3EDGFypZOHxoXXeJx5HC8NwpNWJewHe07jN5k6
MDLIS5bTCE7C0mg3ks7/+dnECo3sfsMvIPIJ2aOlNI53WJjZM46z4wDdN9o8LFO5AkeYwDfyKv1d
jiVz5dOGFBIuzAt0EVeOJnevmwep3UormQD3UVdWb7cGTQ8AvDnoYX/GxfYI9K3lWnLUNlO5FMV8
vL/qnjrbdi+YMYxXVsEhyXkU96S/p0ZLiW+FfiAkpjuZcl02dqo3TfrLTiavKaA0wsuSxONyp5tO
zaqFZPzTr7/13NoWqZ9725f2NCCHU8YaqZDEP0DBtY8p8ZTQxvh+b80tqOfAR842i1yGHEQQJU/F
hLsLfY+hWz4nEOITWHo5PQ8k/CvYh4dX7NF9XUztEBm2R37B87cOJgmHl0+zHOHVE8kmYUWtYY+R
zEMXYaa8vOVspO2/nNsd6iz+FBO6+H8KKbnklYabHRnhm+TNXr4WjyR4Msm5C43nFC62QwGVXtJf
i2XMI/MNUJeAjO2nThbgyeNsxTPi65GEpPKvNhWt3PaalyqgI/DrKKm+AWAYi7A6sCrQ7G68KvgY
+PGd3vJ8VFkMnGtCT+uDGY/pCtU5o5p16ZYo4s8vI1OLmHdWkce0qUqPFds/sMLsOHcyV2UdVp6u
NuZWRqkvtvNp/kvOvlu2I8jNoQRN4Tz+ggyDxi4QfO1YJD9ZSt1iF0WB6bXB7Irq2G5Ad5boXWhS
k2owOdD8XYYpZH9c/iNaohXiGr9AUSgAylDPXMuATe3Gk7PtMeyJf9LR5Mnx23u+Mf8yr5iy+6lk
5sFSCHKXYSZJSEEAUIui3TXmECKQa4pPB+UP0rE1OLzKdZVzy143KPc8oGtm6JpAId66FjUXPpOm
OEP2qGFHxKl4qH2jgzwl8zpDkKs40m6oxHRL5jCNFezjT515XWajlsYol20D/pcz5w8LqXRZvlVt
bHcdxIj6MshIPlnHojBXsUzKEOOTOgi0iNdcYGeLJNElChQSqwtxa1spcXKiCAy1fN6eB6PRffan
bEmjU0GwGHL2Q8vYlaTuBVTs+ztWWEuI72UkbaHCm5bdc+wesGZwKLY05DZnJN/odxGJ7DCznu9N
jeOjWHjbbAIAzI6AmoppC8qUuV367ginXjCZ/BHSiYb3yY5fsRKpZnD5Rcvr73CudEbX8y6gZcQ6
9YU74Xo+KbJ2iXfQ9KLjBvTM5NijRg7HJmhdLcUAEVOYQaD25GprTEvNM5Vmg46Cxk+MRlArIplt
VsUfXdv1bvJYJcxM1J2dZLWdr+/muN4dXIGTOr5NmzBNgG8SSgpuWsbs7HBRavam0SxScBgyJbjK
ZUIWrhzCQ/iRGd/OFzQ7vaAhTRcuJJpqMoVGRljboUHLkWOGgfHm4Kne/kh3wvuXK/A3ObmPOhE4
PYtQLPzOKBmtb1ezyKRb0N7WDrM62199c/ljkp7SdhHGTgb/T7LsYc2pkpzeREFIaFGihhKcArdf
a0laDOaMtFk17xO8a/q+BKzRjhe3zDlqLe7JGfGPAFSwJUx+RuvXBUoH2uodjmxvqKkYIPCi4hrN
LKlqbtlpq494Lyf9fhOMZWdqsvQrbMHbMOyzjbbbbaoXxhFip7v8VM88YGEBUaRkXkEJoKFELm5X
kbmb/pG68Y15f7r+Z+Q/MomcpmcQQLZfzpdyzRkIfQ+9HDD/SPAJ720De0Oi/9O29ufC/eZerLm9
+m/Vgzoj/ZrkcDfsVGqvtFlKRJc7zHC4XTqo8rJZ2qhL2zIj2Tuew/BY9yiSpNftd9WT8noIh7Rp
9Rxt0H55whykkTRmSl362OQBxoX3MFxefbE5CWzNr1ZHiV6nOU7gNQyZeLWHQMh7NfGtwcDFi3n3
tRKA0o8wVMVP+im0ELWGdT58R+WGVFpUeSj/fV/EltiJ8WMtl+lKcw2sqj3N9QtGkTrRjIFal9NH
I7P/CY3JfgHzaslexj5VZjwjIqlLW4ePYRQD/3ZXld0D2r1MZOtz1xj44AOLHm99tBMeONE4aWt8
pvCJRgj9/Z8nGyLHDElghfdaeM7T4KDPLp4WCUMJCzgRCk9l8ddz+KXYu/UQB++XhVas6j8dB6XW
JVdSluQP7sBxauTBLpsugMFCeOxsU+vjYY//+JwU1oZHYk38qFh2cq+8kOUp77Ql0YF4EUft2Yyf
mpWRY5VOIFIvE8Rx91DQUi2/6DqCw6j4m47gJ44J/WvZ3DWjz/zaRpohwbjJeH9k1nZJgoaxQ7xo
525y1sE8y5q5YUo5pF/KrbrAK2lhbOovXkxYlSvt3xeHqTsA9N/Z5tqSXfhJm2iRlytjZspFnbNh
RdIadBcb4dZ5PKQUt3aymoxaRVPJ6gbPSbQD9Xvw50MdycvVatR+l62kS1BungqZxXiyaEXAvPFe
exsd9ftl3yP7+aQH4PI6OHKz9LrCu2/MuOkcKnjm1SPHxZuOFMJDz3lz+WY7FwuC2PwjgArxJvrG
3dXAPrrkBbyKF6uFFt5vnvCOdoZaMVFZ9UzD4gOFzr2zaNV12TZoh80DO5IoyM9y1HfpxI5jyyXY
TeR2SUzpTGtDqqkN0DR8USvbdNrBMf6vZ/QpLAop2yVUvQYNo4BRHGn5Kr3py7A68b7hNGWBo4AL
Yacoab11t0u22YWG39dg9kuzhj6bCKie7Fa9eYzAXOHrGlMVWhK2UJB9+lOC//nmCuwHuVXd4fnA
HlbVhlE9IAUlnKlZjp0Kp8fNVP/lF6+S4U07OxD6N/6PeGeIEGwoNOiIiJbrtmCV41/V45NVZF9v
uwnKZf1PXDujlqIjjaHWamHbJOWF1trQTtqbGVEPjR7LjiWvywgzY0dRUj6t+mcO5zCcfGmFe38r
dYUlOQ+y40ejbW6U/w+arAFpP6Qr+q39xKNaoH5Tp2nFV3EUlIEc/F1+3eEWJWRNAvkAU2ltWJ1J
AQLQwdXIIVXWIGM6CNeRIjeuE1JRNAmUhv0+5MFKixhYrYm07cWZx8ROw+PdWhH1/qDwAopnqdvU
f8hey5Apx8NxDuibnjNuo5oG9axtrEj71V98jWm1Eienqn0VFhpcKuDTy3z5L5YD0TFTTJbT+WNh
maP9ngIv4TBSoSTnNXC1ykj2ma/aDONjKzykExVPOq383nKjbnDtxWQtnocRPOHbDT7xHTFksGQr
Wo4E7uWDUEJPUq7nCRWJoOFerGw8643Xem/5YXbkxB5n5yVMrOYUBsXzjqJeb9Z1Msil0Rxh3ruP
qkySWELMcb5UAUUY2WrsPi+u7nRJQ6CROT/RaSlQGlATwvAdJW2XMtN7l2WeFIPEXWsO6iJN1Y1y
o8n2L5S//oRM8Cu56enMCQw06N7gxZqp1Elgj8GSpc297BrBbSOkx41yF6wGs55N8kv8ZWG0O39/
pvPNO8p1zth3JRzsSsCaw4Mz77pKFyBvM9Cq7dIFLU5xoXdcgofR2fEYnImexFq+pzkHQoGc52uS
FNAB6IyfPW7cSFvenon/DF+JYWVrXHpJD+giASypzOLbJ8WAK+KE5SBPEcM3qONeE98vtk6oHzmz
bc7H9AU+CXfG9SBzDHlY0bYXoEQG4w7+0YWDO4TBqn1YD+KoYIvKXOwdq6SJeyHu8QlRHqfhMJI1
iyB72HPpBZ1Cxbxfs+NWr+IRm2qfWJ+fgR99ZNcNEn9k4imw1qsKNYaq6+sVdyZ5t0MfRpJrRBj1
6vOUq9qzwm7wdKwBKoKnU043GlklFovXx7soGLRt8WOWxq8arNQH1shKjgct9ouvKMGI6bPHQrBx
ahgdKnoCBC3qDHa76CJNVMIRQdOOCMTS0ZgZ5hkVIL/zBc/s00sF15bp8LlcpSS08NyVbA9ZQ3cL
cXrdosB0syMJkN5BlGspe1bruZX1eh8dTqzJKn7zIs0vFVXepK8EWr+td771BM8VXvxznlBY+aPR
eii2dELPmdIX57qrOmZdZVN/VzEsOh7tmaP9fEzCbBKgugTLbLqz9QrhtrJfG1djIWRHAXlRm2vv
OqUJjR4yyxCCiVN+jYnPrrQYI5wSqKjhgA1Aem4OywDj5iV7qfbs26LMOOZVuQhhyh0iBq3fDtr/
JjuWPRBEM/ny4+ts4oXfOLzK+L5522ghtqbFTrZARvOLxN9NXK9oamnC2ycnlmO+mafuCcubedN4
qhhdRLV4vhVhpNiMINAtJMk1OYKvKEs6w48V6lkIbZR/Rx+NWX4DcLfLUojDqbrl9R9mYkx8KASX
YQVi+IpUMUy3rFAouzkIW7fSHdEq+DHpqnjzNFJ06N8gFN7tRJ+lJZn8VQZtvFVGI3RavT09H9cL
Nlpx61VnJQuuXrj5r3snIX/9kNOO5tterHG59sKo17tmr8R1LDAzJ4KI1DNaj5QzXTCYYJzZ1bB4
+Ox5qVdgX6nt3jxkI8fbmUl6kMLBS2a88BsVZwa3ZAe/cCFF/DyB4t+0ojyoZ2U5Dmd4T6p12J7P
s693f3HZX3RrAtqabgNoE2GxZcRiRNMeKGYT4VRcJ9ltWw9qZYu+mwEHIw/14an/v7FRAf2VwzPy
FglOUEi9X2S1us4Sp2f4CWAWUBgm/AuYGqgOBTPqv/6RNMckVyHYiCPTx2DrfVx1lwI/7GdLooph
NRwgyPnvd2sNUpvalT/3l9g3IG0Uu5zsIfw9osDBYgc9FpM4pWjbCtrNQVhChmgScuPlzW6x4vOz
Y4TFu/YM0gN18+n85u7ZI08n4NaUgtq+b7mml33VVnlFcTiVn1FnG7yep6wNymTkTwaKg10OBNab
dPhTS48DRwHxhcRAHOYgWKh5gSN+OAK7jX+Gz05SLL9E3W6OdzSV3VkMAJTNS3/2X6gE2emMUiNZ
KAC+HmGhWZvXNToNfvQdCUkL8ego6ApG9XXx/C2YXCIGJs5m4TqEIvBmH4PQ8wREfyRH7DdByUH+
N2qJZbYxbk6fftGLojR1+ywJSdIuB5ojiFK2n4Okr+rYWX06yiGsSmtwgS1GepjiOR+6/eV3dIX0
2AJOgEAzro1DYURsB+sbLzXIFKPM3s+PliLeXs32SBR0TSO6NAtBHAMh3Dv4yO5p2zGQOUzHp0tr
L9lJpNTdWKPuBGZYyW/r7yAFJSQIA3CXRjDy7RkS6xocoZCrxlBOD4NPLgWlWt0SRpuxUyaV58N3
EKNNIrOuLA+fB/aadW4FUt0cPFl0qduSJi2RNUgb6is0IktnfVVoOW86Y/cHKZRgLUSNGq1hWdzu
W25o4zLRH0JqF+dLK0uUxwa8xP8VJTZwfDvaDmmtLPhaTJ83aD9a4T9fGRCBpmu/6Do83EuHVqjQ
8bqNW59aiFuzRMLkAvDFzGPzw5lGDJMDjDLBh5bBl/vPX2UaEDY9QKyDWyhNHqFAyahU12v1TjbL
5zQgQIHnlSGe0A5/g/nBGT5qSHZKl3I8kxTisq0azs8e/OfDCNqbOHHRPB1Ex7GC7IjXbs/a/yUW
LMhdYk+E4kgDS61t1JC/mkHcuYNvlniAFhUbpos746v75fs9XhobApOjbMQnaXM25ZBMElLu9iPl
WBfkrhBLD/tTQbVUUiQFnSm2t8bttlBZ2VeQkbuFBh90WZXC0AmTNN0bp1eJPO9nA9wX2QrKhs6h
fKZjhQUghGcZzndjdC/6gAhbvlhH2NRYeMo4fsUa3oQynEH/Zsr0TpDtBJR/srNSonlPqFFv7XLL
Fn5XrfJ8+PgSvDk2jAujpKaKpA0b9BPh41888ZYMes6nB/ChihlKUBHXoLF+CIlHrp7wnNXXraqV
1D4s98j95Zu6pu4CkPeXqDYndzGPdXb5PpUkB2GoTkEac7M5pti5KOYm6pzBe1h4V83+B+ViI5ds
A6qW7k6mdL4RlvGXO1BDJaErvxiyylMB8ajKVsQIkzK8nyOePI95lK5Zv4zSuNkerof/mM+MXsZH
MwcFv/BQafKslDA9D8P2T4FCMPa3zZo6YmhrGuah3ZinqvJvlntRx84+lgj73h/jYCs804mW2KEc
M7vwY/Wdlv2FjzeHCWSN5To3raDk779irjPJhXA/CMnlenyK++UdFNH6pPvqH8z2I0tutdIoYrPa
3i6YmI5Rpv2EtDjpqkPgLG3BtY9X6J+rJ47dC2NYT8PHdaV2BE357WFqv2OLUuHcW+bUIJD1lAmS
M35dbw0hx5/y/ieRbRxK6+5Tq0s3RhdfquqqHY7hZbBSqtz4owV81PjYVbvSQKtc3jpl3mR2Mb7i
YSmxrMefmbNJgmktr/wHlZ1fnLRyQncArpFvGJx8YCiy0IiaazLhYz3LwJOq9FDSe5LsN5/Zj5TM
HpXxbU7OOgbg4ZpJYxXtTUO/ZfWZgKFAU8iXS1QhVSNITMdy6tgwbUxaFRR9aKVVS/LpzmlzetGT
2/oYG7Z9lsyFARMEdwAHksedxEmwetmOvdh3gmWN0yNxScWfSoD6GuRSgoKrpg7bz3Sr0XwSk6Xl
xkidiUw4eaFBaEE7TyPJm1KWFVkR/a7zzr/ED+ZwbgWV11Gs/P4f8DUOgKAmWaFzp0E8g9q02mlo
/eepLlHv6PozCjnGnCUf++2NRJUtPyQGgi3Etv/GJUC5JIugRoWEJnlO2YP0IXI8J6JvUHFI7O/h
exxbOD38XvCKxee3KcL3S9AJwjBWidfGYfi6I4LCANjrgAZgI3ih0qDVKlvV+U4BIWvTcn8yGajQ
O7U8S/zdwC/7zEKA/11DX+nYrA1/JzQI8BkahyQcvlze9gFZmVCqCLiWvitjAme8tSPfz4H5DcoR
PxKz5YONuDun1d0vBun+XwTZYlHPrnasxbJuDluHEHOVuu0orEUbEd1ub7f4HkWRelPZdov75bjM
sAETBlRdMs5/K7whG1A9gI8wqVOHl5DHK9U3CQwvfWqXjnhKrZalLn831c3MJU1iuNoRwJfwlsmN
PlpLGCLXGunW8IGD0oOC5RnGhY0FGpPkfyyClZSHyft9pouJRHC5U3QzXieZ1tOb5o/cCPLcbyLO
yYvMhJoktCbo66zDTWkBB2cznKhs07IT8z7fvP+z0AvRYugvmCevkWwKZgB1lsBj/7hy1aFp15ym
SpZ5sjUV0tSNF222dIcS9XU48OASRNy2Sk9zB9QHMbNlXSRDHyJkDFu938wKp/dGlTOfGnnp12Jl
TDrmcY6bUaPBs+ktufAvoWtFJvII3z8HYi71/3RcFLvAXrW//nTAveFY35cL1QhmRqGLWP+CD9I+
2UF186TaY5r+z7ag1mJdp9MSKi/kUNpjTfXlRrM+Gwfp44b+ZmXadUimA9XshtvAcZFcTjmD292z
Sk4vTpHmXe7ueqxyNgqu0SiLD0ClC1ehuAs5obo08YZ/0k/UvZ3Vw0Z4Blg7b26kDY45otYkHmbW
sZ6qfVSCRL9RF4LnSt7BR0pXcWw83rh21pUAF+wxEE3pxbfUiS3pFyYflO/bw42ard/wwDpTdgd2
j3VRWILA7ju7hQBBGGxKGPO02rKxwNppy0WLjEJgqvTVm/urBTr3BAaHSjY/fYViogCMOVPbfwvt
kjCQtTmyBB66BcsKtwRA2awlenSIg71rT3z1EfNYcoaYB7+jaLDWix5fr+T3YcauhgCUVu8awrjZ
NDp2VqR+vd+v3+CmBswna9HEo9tlBrX2ujfWvyQ+7wFOOYeA+nxoRcKeFLMpCjEzRrvmouvem5c9
nGiPzKFDJe67QtBoWgnq5h3l2jd60maEr+fQ83b0yqgwmD4BXofmrO2+DGPciapClK6pp0FeKzVn
tMXC+iG4w/0ySISpYF9iVIWsEYTFHUcyKP146I4gQ0t+YPXSGHrkEtMGYv9LhyZbKyrlGlSzyeqm
FjQY9UvwUA1AkKC8yg5kv7s4Vi5gkrU6LZpFoLJTonZ6STYjsk9tPNoUSbHHhatt3f/6Nt/kPJN4
P4LYmP1jbspDv56rwJLWGZoClAm3UZ9CCRThV0khqzZx08v5XLlAbAkT4giIOUKxCOtZCvPH6jcV
QKonpDEEDBLyWhCjQlmSPJOEevLTxm4V+c4dg2irWVQO4++C4xhZfL8+DbxDfUE91LWIUFMzv6kv
uei13gtqdIKXO03GF/3k8tzBrcjqeGGqO2Bu9B86YmKnd375pDJc2cNjeMfs4mcMvydj+yAdEd13
GSRit092MN8np8eker3/IMedv/OBLPJ+Jb1tCX8K0N3e+kHy7xqS6MSVg16s9hBHrCEQV4t51JkQ
kqHd34GHvGI9vWYWqH5zzKbZxpTMYeziOZi/RAyj6x0ZKxPEJ6yLsl1yJ4BPiDLjy92qbUO9UuNM
y1ndc8S1BAEWgSZHTug1jk7V0Cj1459HHWaBXk56FzH2IrH8p/CHGiuFHkq3kvaTCvb7Od330HcH
/LNoXNZ1FpXl+JL0ZEhmCriyu0E7J2Xxw0IMIeu1Nvlt8cp2CwLOTuoFGjELgKcJHtwf4t/oMgN0
e7qo2vy6IFI5yX7vNUzH0k0TJsWGqyBi6xGaaulVzM5Jw7BMBaTrLqv4NPyjxnJl6g212fPtjYIN
UFx1++C+kCKSxlTDHa76c3QQedyGjRiW8vN94h0XAZl+prow9QibOUq5LIGL3ST5sURJ/ehDSSKw
vOVnsiHyjQPnuXhq0gDCJHMT3F+mbx9y0vEDcYz3PWDhXDv63cUnV7Y9y4ss+PvcJ6xJap6i8z1P
MPJJgF6atwUR1pAnOEedNwbLPrcyQ8eVbDD8PXozewGF6DZ81uAigcR4xXfPLUxB5/hKIwvN5/Sc
ZVtbE97RVF5RSJpLWPcW4e7WSt0lkF0Ei8ZIZGJgfEBkUL84xpZDc4fIydcDNSjHYMsx9CaZBpcu
UkbcnS/l2vNjAmI9jCj+0FaCjYwL678MwvXVjwdKA0HBWU+aKBl2I8zkxVjDfI+qZ6UMRhhtWLsV
eigWLXWUJ3Asb3S0ESUNf7cCm1fTSCDICTUfwEPWcsZdfIDsYqSfKCyGhb0NRiX4nz+1AZjCuVw3
fQrAal0G9NJ+JG4YOT5+y8fnI0dV0wpQQC55L7nlY41lTvSfTPvO/irm5rHEqicBa33L6gMmYO6J
WJ2Ib8mcbH8pK9eTM8hk2WFxqOZAGqU5el/EwSp70wHrCrKtEZjNr9HQ2zNvCvGPCUDJxK+qV/Jx
bp2vXdYEUCnVzQWT3FWzhLKuaCu26vq/AZhhVGLNHfrrdnwQNURUQdW6xqrZ8AT7H0//2sE4ilQ2
G3WBh5yC256APUS0/oqfJllOYK1p545sm2rhK/7vLTPwEhFXDM4qbDYD1JbZrv8jO+W/zkd3O/Dc
BQGVeWkoQAftpqte9LFtO8rrS+7lmW3OF3x7A9Mjtbbc7ud4V9TydoaVvqoJ38wAH6UAi0SIKl2S
GmblzrBBeEt8UYGSJiWJeoHL08S7Sn7bLNy1hrcPrNBN6gTuwSacibuahFOTHUx30HdV+/8e4e++
4LPWw3nGGIcqZvz3pPZfpTibXXSV5xIR9dDwYlK2wxO/CDHzWx2kKN2xzQcTCqSeENOki/sZM79R
IOK922guRfM8Y2je5dWvC9ziKxMuVo05u1nTvJ5ldCGo8dwZmMFxubr5x53YMJDSruLCv0Zpg42Z
81asOygkinObR4wrddzK+IA/KsicqzZQpjmqdOudPITP9PfnnKJc+0Bq57l7ag7iX+4AvRbuRu9/
2zVNdit/fgzobIzbzDbeEkaOhRcD3JAWFYm3RktgYHeU6jIeTvhGjH5+oGUP+MES32y/suTHRwDD
PWB7UvJsmTprTSUwNXqxJ4e6b3eR+pXDsO/M2LzDHTkhRL77snObZ2V9A4NQOYx+/7WEDllTRaK5
0BeobTVW7hGH+f4rjmtV8Qg+Vy2++DdwVrvY37D5B1GK/CAT/g+qeXH3FPdUGo1y10m3n7xveBAv
Tev4EmXBcuHdEL29p9FViNRlMees0SFhReO8753pCd52K6Ahl35wumIAWj7FD/vV4HyJRnnqVnFs
ep7cdJLJYmwk5vaBZetZVyfQwJdBJbmlPz1y/+BpRe30uJHUUzOmrb+nARTEqGxvXnuP88HpSKWO
ijMk40cIdTjiVJZCBntV1OLVQBRUEkP8sHxEtU8wcz5sSzRr855/QqVllOmbHmuv/Xg67py3vOjf
k9/DUr+AYp3bWJXjFi+4A3I9Njz3oadQmFt3V9ODHc2ErnAle7niokXSp9kL3a3911VesUJm7c3X
2msQsX0ekvgHOFtVFJ43zA9KRRdVRP2ZyVDZ+T7dtIl1Tw3h1JFVX8CQn5r/e+oQOUraCFvz7W01
XNj7/v7bbq+7F9/WX2zqoYT3WaaYhTQP16AYqp8FIEFAbnompC6Ul1XfPBbBoyVO4lkESDWI2hyS
sB78YYWl+riF9Osa3AgoijLw6X8kzU3zJIX7Ryjw7EUEUHYw9UkUtO3I9YTdXRjmpbMopAPKV3aS
lzNVo/YXkZwoElX8u9lt2i9lq/EOZg+DgThzqx2KAWUTWGl+KyIPcy5jQ9tm3hR4+USo6AkxXb1g
xceQShYSdYEKVOVz3TYkROlw4Ztddaj6ojfbD5+mHDQ4/FdVDGrxhly+mQ3skDoBRO1khGxsHccE
i7gFp3KciAzRGcdRdC6W5rsupEfWidIn1JZijpeY0T8G8Z3bNBTvPjLMDKiyjsRuLKv+2xTGSLY5
0GR0Nn+WmWeSifDrsFTzICdyV4SwNcBYMzg42Kpd0xCgp/+p1rX5s2TEGw03UQcF6JlGzA+QbbVb
1Duu99NJuRSX3z25+yI3x2jgTLDactyKUoiCWm5VJoiCpQBXDQ61CQc0gIU++amAbmVdNLbZAI5E
3SrsD4AWpdUX1Sp/N8Oh41Njq+tmtoY7KujZAwujvkUOH0t1viXGkigS6DovzL79o2VvlKSbHeHX
KJAOllDNgkBzKcQcGMSrZsJmXD5LAPyEXqkxFxKBPBxoob3JzvVvYk+fO4rFsxEXjgUnZLuajjIS
MS80uuwQDHuDVdlCWrjzmTaxB5QQb4IKg2MEdB64czYIxMBSvlqw1EEhyWeeFBGnZyqVV31jj1vK
S4P5/RETpZS+dlffaviEBfbF9IlhNl/a4BPr87o5OqCeeL0dY7TuB/VCKPnBoz5KQHKwSvWGcWl9
YPUAjKyhStJv+ww4COmcMhwPWqhDmQiAJK0yN1Z0KTpWqcHGRLABCumThFCWJVvBUFbnvZ704GfT
32gWYUj6X4IvkgJQuPGlz9tga3T4Z75pgdsMGiMTN8iEj0ylfHVqFjDBRQiFEyH5gEDh6F49oxqd
DooRvDYB7+hUbpxy58PSfSaxRUSSh2gEy6QWqHrsGktYOwnlJ8SevYs3p3j1/b0kl0mH9t5AxsS9
QdTxXS4jn3HSP8eg4rbYgjVkzMEaMgsnJYPFS05h3ow08OWeKFrhw0Bo+H4OaJzON/gDNkbclilH
A2yIxj7MLS8GFWMQ90Mp4rCJMJ9scJwkJ882WBLCSj2SIr7d4xu0pP7iFjTWzFV86BWt0weg0YOu
R7t/qrfSR2UsDAvitnnnPDdb8JIdQhqsPibEuofCm3xZ4Duib+13xI+8BdXqSFUhffYgh2Ktx7BX
iwwa3lSq6WL/bo6V7hh+XCFiWToLi+MYIPEhw2cXJn6dHM65xPxD+rqogwA0ceZ7Y6DS9vlc2lUh
nbaS0zAM9zf0rrEGwW0JymoCrjjD5wS0PZvsVGpsjXaC6QfJfSlVzIJ/1KepIe5rgQKCMT1dn9cD
XUi6JQMku4RNai2maep+AMBzt6jzZ4mYtkpn35qMYwzPpIqBPldr/mBauabMT01WOKMWIaDciAjQ
Ky5z9ngWPdGDUMesVkj0f//WvCE6LbVZOvOnTivFxT96rn7swIti2T5Fxpuvkxgnrq2h8X1OgXDK
0skrUNlSSDNQxS9UaUrgc5wg0AnX7odTvx7kUiFEMjo2lNDK0YE4RqSg9jrHzRhhlij2KIe5kROm
GeMWoI0tvx9l4Tv42v50DATnX6kMJZDxe5cTROq1klyfAG/mjLA3HHCTT2RNydvuJTS2sZimleK2
gwHwz3oU1jBBlzEbpJZWjt++xNieM4WILTBYYvdTElJpwmQf01Fe/Q+fPtdiCHOcVg3L1bzvUvE9
FlLhtCqui6Ozq9Us5Jmve2ZbYd2QbVZy94szeqzNx+sYD9UMCieGJZ5fAHhzYwSm18kztW9H3rQO
T2btntKmA4a0AvuqNX035xqO7GCsnbvlE2gVcMcuqkTYEdi4RFirl6qCj34aETBSJqx2uLyIzMZc
jVpMSDNIfD9MoenJVeC1hjx/IToWFqnbGuNSTSxaSV9JNYWtc93KQN7XS7cGRLQKNxxNL4VlLzLM
5eeNoMtu9MsMnp0mduUvV3LZ4ZYHqYENRSr4vVeqhCHLBPk9GDM3fJYPl1kk8QhK0np9bXmvaDsJ
MHliPOX5o0lLD4xv2RiQNq+YGXeJ0C+yhNREtmbZQuZ3yCKlu6I/6A9kQflG5VIOFnwDSxytOb3R
ex/EdTXh+vc/iPcY0u4vIvPWPpAtwESIP9sEZafYeIzN/YKGeIokTvT5B6sot2ra2NtJfuwsioGm
E9fXN2Q2eGSfg4aaCfSopeSMIJyCxitTvA2LZ4cJquqwlIDxWSOpGKCWJCIFFQBD9FChLcl1iMKf
4CIuGs78of5RTL+eqSkqSGcwbF88olej3K/p57Jc41UzeMDj1qHPRlpaXVvAreYDiCyL7Azpqr2D
ZJODFFNQQEJeN2xnLP/PwcfRxHg2BFTL6W9vdc8sSRz7vQvJ+9+wcmMeoqTeLBAf4X+o1lbML03+
C5T/CyyrpM4lkZqDqOe5yczmcuQV2l/721/BCSWNXDz+q/RgmOZ4RiGtJVd/HVA8rN8v21nuirSi
owpqJ3XC9C56H8vHIDhUIuWAeuCkzh4J8uE4PB4KoDLK9Jl/Ag2aOFEziWDR1pBBHNMMBB8iEav0
Q3DTDxoWnVQkfBPg3Bga4RBM0DA2XwRsbZOGQego1TfMLIyXVUjcyOgCNwN6B2um7kdEdtXPT0Xj
cEEHi9gxYz+CgmACMfR/5HlTTCqVPHqiPWQu6TDFuOsnJxBxQcv5g8Q+eh0bPxqHvD4rQlOYwpiX
CVWWPmVGiKF0GZcdK65PGKH1kTQN21L+PdDM+2t+Ow9u+cwY3M1qzEgR6YsOsvtU/JaeijdcpdNn
v8xcyDumfLC9IdOO1n0tmPb+k5/hDE3uN/Z7Sm3d+5EfudPSpcRyor3Tr6iBGodjIkNDdPBOm40/
RhgJcSOJtr+YAWHnX+PZ4zMRiNLndP0GsdPQQaxJ3Rv+Xp4jmc2TcrQXrK52Omsw5VbbW0BVEpHI
jIEx0Wo5oEaRxwxAc4Vbs6S5kFIGXgDBONL4TbH2uyqmu/eTdanDmMj+ZMEImvZmyzfFhBbfW6Yq
2VPv419+AxJY95mV2FSk/Bbx9yguCb+4EsfByHnNSEzzLT9QTtQem03Qv4kbSWhMwlhU1a+gS7li
eC3hNlA7ChupNvuThxcqNWOxEJlQPBKvAkdyCCUgoCRSh/wFS9Boz/Ls7OxDQUReRHiw39ps8jJg
xgj+PYV91HG8hvw+LiQJxRue9QvfwJpCqF5KKav9rBsNOxYyRPmxPGDUvBcLQrvD3yEu78SxgrUI
FOMxWObi3kDCcWZY/+6NqAv5LBH5zQIZfhu7atPr+6ZkenRkUvUMGIH+lNyo7GKXWR6oxvlGmG7I
TmpvjYYFifJb/c9p18DiwYPvZQxObYR0xbjwHHPbPieU4NiKkDuZDy8X5WNQRrR7GBCvWLyBxNLh
haJm6nfgz822HUQEnTTup1skhJJQMYBX+AqFI4jBeFUqEc8rx33kff2VeIRvyDRyHBRnF0JyChY9
+9xq689J9fp+rLl69dBcuPr6v05dIK4KxBRxWjbQ9Ke8uN03cEY+PX+XSn2+Noyax7dEUPo53xI9
ydAp75nMa4sU29GX0csS+w7PmoGA02iSPt8TPmcB8ysgg2wctaFhVaWNT6R5fQy0gFOPyA4Bi4jx
xVXOQ1yOg/9Du6dJXcdparYjkiBg+zwB33KdPNDJCCU2nBHsgPSX97K4sKHagu+EfLbkXCJspWh/
+LieMUVUidDJR9joMF7UoXm9++BPohwwi0J1FpRWpRcVCiJO4vUnROhpG7FvaB9J5MZoesjxlCS+
14xgd9Vo9gqyucCXv6IGPNI2tHyTBBcEPoXtIUgv3ZT/Sg6kibngpsRvSXLjqLuRO3RDFolZk98V
nYli/m/st8SEMrM0mlFt/91npiwh8s9FVmiFfazkFx5xYQSSxk7KAyteEm8f3w7srxMJIPzRjHaF
sw3l8VEGzZLf6ZOzti5Gb6qvNQFgrehPMIb3uoY7ct+VLVDA1IXX9bYMNsY27t6fEcVgR2j2I+KI
Hepkj3PYESJUIp92o76AXvZ09y5njcg/iSRGcAb4A1G29/IAN7ofsnQz9eNqINpi5NHLDV2O4A2R
SXXi//tXe5ca4+OkwDPk6ZsZtJqBumRIZrGJrtjSZDaD8/S+MhV2ig5hmR17QhXr8F70/9GqoNyR
Jg7+tgC6wX5LHixq03+iivKEFuiOup0xMpSWp+D9qENarI0Yq0X7FfXS1wWfJ5YkWRz9o7+43Nsv
O/nxWEdJN9slk3A/H+x2TsS8VZk2lWA2ofbtfJ189sNZHAiLjO0VVDTAbZoErgtDGxnkeGMrtSqJ
k1GWsyR6A0deH9yAwifyqFAZGq5DQqDtyaQ61x8Az53i0EI9SEaKpOvTUEZQ61wrCxkM5E2769MV
2i6vpf9fJcgKBmesxe8+S0S5o8sZghCdp9Zb872PwhtGgz1udCrXemihSsIYkaKokKGO2U/VEdXx
mbYX2aJdAVQjWEO5Rz3073f/mJM5F2mmB8+nLw8wWtC+MlxGB0O2msMzp/a0PczIFD86T79T3/uf
0ciI/rdgSV+T60Opc3eO2eoowp9F+WEpbpQxVfCi/3C5V9te97OyTiUgYsSkhEXvyAhR2DLF3dNf
B8hdjHhCz8JFMUR7Ip2YaYyA0hKmI6xDNHGLjdrEi3KvlgfKmsRH9x2Gjo94vGHnJ1x71U1nVdwv
LxvXWt/rLDbl0LIg92XvlktBLElP27Is65VSChUr9aoWC7lZE0tRU3NfbWX2eJVEGhhD48Gn/5/r
R7h02HAlUXJukir7g3HzJeMzJvtHHrm/8AprqGtf8VTwHm7IlQkFT9FX941xGhMQiw0V/ayrMfoK
vc/89QJPEVN2M+tksrGeWCnfp8eCbM+LWMxbb+8cU9wjDX18ryT1kQpiEtAOvRsipUoOZwyvqzdf
cmMl8Xt0nZA+goS0hCXWE4V7vJfCn5sAEV0GL8VDX+Yzszw0JV0tA/hAOc6rj8+Wb/52p1KSHued
rn6ahrwisss5nV9C4Nw0Sp0Vsvptp6kCFA5SSunXAR0NpJEAiZL3S0I1OzFt6uog8cqPCD9WyF4z
5CTw1KSs2AZHXljPwpXoz0mhG+jBRxhZA1SQeiPHtXkaIgkU9BmEu8z8ogoIs60Kj/bybOvrnt2n
Gw3hYCFRupil92t3jRkEaQp3OCI1EXEvWp594OujobbJkzf5GGWIsvk31fYE4wCTpECuZZYbGLjn
eZabygZOoIU0gD9DTE1mm++gD4nP6mHGwryBIpAKTOqJSGeoHos6sIJ93C3RMUeSxB+5eSfEV6t0
QELJSakZKj66EFCPKzfwLOhQ6bA8nf1fLxuYSKuHG+Ow+5Zu/QQDTr49DMY3r9yjykX326NZsoRr
dzI9TbiBBCvzWoH00gnPxUUDa3b1SfZCf5p9LtfZe1urm1LozMDQAIGXV+7uKA03QRWeUrQ2L289
cB8ECp01rVlK5WOf4J9QEMUXdR++LnAFYLq3XWPJEHMh4TAKgfSRuhOPrNcNuZSqRZb1SUpjGNOa
nvXK+QQ/MBktyoNYvK+RtLDnT92XF7EM4t2NaFJdXjKMFmWqnI3oeFJGBvCSEPMdsxoSqODzZu47
RxHOrR7vPuYTu1K+9EGlCY3nDRqYAwthN8/IT08H/Cxt85+ItUPJyYjHaGB2V6PU2TgAkwmFtkHF
UR3UWsLEQw1iYm8PW6gd5+uOBTlBFjrdB/oNPqs9TWANxZkQNBnSpVYwQEuqLel+BhIqdq6UlmOY
7O19u0fW7Ai1U93lRAiZsb1fOSOK95eCtOuMbRoyNgBIDzvTLxjzIymrPYWgpoY9alazvxXtXq3N
bOlFAVBrDvki26PueYUdLL3tiS/vEPOqix9wCsEWkPZ5Nyv6+DEYEnOMGmIfOzR2xviLz5BuvU2W
msPiH+Bt8bqurIueWl+sIihxTjmLdeWnvVzdDqxkyUuKbK0LjSH+2wfXmJD+1S1fYStFNMYeShQi
YENe+63yOBK4GdL3JAl/afsYDG4I2zYJNMDVei2KWMQaHNmDk+yHJ6peSit6wek5lgav3NvMOJYn
s4BvDyGpB4O93V9obJi9fanuC2p+VpgyvGefabhb6FXiU+GDzZ0wkI1AeowO9jR+w4AnAKJPS5XG
N+/5jDioKoQ/M39t8zdGTxHPMpTcb7B+xuHbfew0BcsIMfuYNOP46FyEBwRVXEEBxsMun7uJIrFo
Y0AyUaSIYYni6KMxv4KCInD1WlGYSEbs/OPYTgK8moZWlJ9XMXlAapes132cVjOPiK8nW4KfVWqj
1j0xfKA3bTydNNh5e7ardGGcLytM93BLtQcsHb7QB6zVGv2HK9n5zCPu9K/vBZrYRpOVp1u38Uw6
tV4YklNiepdofwR9Fe2JTwHQfxKSPAbwcuFlmKzW7AeOfhOHtEAA+wOuMc/AODQ/FPQYIENf5X+m
y3Es10IXyNWIbWLyip//fdjKBFfSmRdcnFfW/LB7zkX3UzTAYwYsZ8f0BNGTPLHlLf5kQajRIib6
echC58+pzgIuV30i7SfFZOeTGB1277mm3cI2wOJO+H759t+0wjMeiIlkZNl+c8fLJ/OCM/jnQ9zF
HPBQaKzM+y1Jl1Z5QUy1BJuWTTi4nOQnvBqRBQ3G+w+y3fnlkP5GWxvWEHEIGIc2lGJypZteLHqy
ayEuu0VqJJCbQ1wSIYgI6q6hPaACYLDofq05icikcVCC1A7xK/PtFuJ4iQRT+nZs/kPUHLwAaOis
KiZqSukzNXQJH9KxLhgiQm8xY6R08IptCA1036ct7q1vdxxHwM9Zsu4z27Go8kOZ4b+TV3VUze7I
9X/qmec9MYjpb/r+3A+K35dG157fyKUVxvYw5nki9jsxjskqHNrvOVOrx2daAgNFq1IpjQNO3U7v
auk5UeKAcmaLrcJi7euVNXcAdg0zXAI3t1BJrq5WmnrCF78z14LKYROoh6ta+8T11SI8axTjiOD2
x6XZ7bSrb2JtUVU+lwrQIeMYUWM3fYLN8GOXum9qWCzViPN1ol8g4EdWZZWMEC0nsSry7NXZMXh6
zpRM0W9XgApCNn/ahghNOG1QpXsXfczUm++kZXg1iOCEqZt5gHjsWnrbAdE8c+t8ptEq8yBNjXTx
ROuVYP6nvMbnMi7IKUEjGxR3ZNo3IO2bz+I6415yl2Q+4LqHZsMSskNKUvfEFc1BvW/d5ctie0wo
Me0X9I+7Ofq27n4V/ytZw5IFnJ603hGZSHXP0ZkrvF3aX9mEtgYxwOkaoB5e7zMtU2cWzLzNNobE
4KkuAUjUhpG7ERae+KhYno9cGMLpDR/8ofEg5EIpr/ztGzo1l38xUevKOSo3KlUl2GYeiwWKKdAe
fhmMrDU8UlR7ZXbDH7PIiRHgi/necrG/SqUN/RPAMwWsjPbiqU/wS7o6rR1UHpowXuNBvQO357O+
kqO9JjTuD5xWmtf/cjSE5x6vzzoZfM/gCvPfgZ1QOHKA+TdQsl8ZUgzgt55Jy0sheSTbqIo2ZCI7
B13cW+oGJE/JwD+ma4aC4gS/tVhIdtERvTeCAHdV0bWhc5tFkT7fUrg8yE/CB5nkV0V0P/GN/qe/
g3G9nc3OIQT3izFwuP7QPZ5KzwN9PaaQoJGnsICwp0gnVlnxbUrL8ymAvQipmdE0HItvhk3YYs15
rcUI7hOuN+KVogX1xDzUHIELJdiC7BHKOlVKYveKBWtRWuwb/sEUsF8OYTIWqOGnu52UL7UamcUu
NnJZjRIuyiEMJ59VC1sZMxvBY0U5EVSiVZzsj9OFPI8pw2uRQGnKF8nL7dtXKa9FnTlSawi3rZLU
HG967kKQtM7GG7lxAhYYBHmevXc/xA0dISzy0c/EVBfacV1wlhOpMvmYtjUhMmMtp7k97tgQtryE
uUzFV5znjcke04QaD8EMh8CceD2YO6PFwQxIeH5tRXwH1Z2HxHd9OkjOYzr9gJ5P5aMyfEh81mrJ
j2MLN9ohGbbQj1PCLIx2b7/EqzZEjDrNWAGMN1NEKF8FNX3pS/yM1ke3kEQhgNIm7xb14/InOU7E
h6gXVUgsv3EYmoM0qxBsqAN5bDyR3dwk6nRDy1tr67xqZs+xRUsaUbivJEhplPfxdgYY0fNcjOkC
8gCkNxnF8kEA4wnzuos81ELvED5z9rVEdZgHK6MW7s5rYs7f6KpKV2wR2Ag35AmbleEzi3mGxftq
lOuh/K3N1pCfRGPhelBBTFAqkWICuwQPbMZyNNfVGIHt5j0MlHK1uKBgSgkPfGCUbiQwjVS3t7Oj
USoa+p7vRJX7ia/asLSXVJUeupKM0AQohjiVTlOb+RSereywuGWtvWtz/c/NIUGcw71GgbtgDPnp
5gSx9X+Gx9GF4UmVKp1EV2A6LSwYR/IrvwhYx6XeDzoimHDoMheuJkTMZ9Ist4DPhOlcan92y1lb
IA62ffedwgUMNZXNCpMSRhpxvfeUAi54EHQl03P/kXN+kTI8vSu8ju+oAR4Ypn9Dk+YFl2NOl6Nk
oik3i4alAsg2RemiwsRGl3/yvoY/o1gaLQwDVZU8ADnRqqo0VIh5Z6QYvUi7/fmnJKbXwDchaX9q
2DL3/sSs3bC6Zg4X5Ha/cuF7eVDGq8D4CE3QKhhw7ifd3rY2GeSfwkWrIKrd7GgaRj8pfgYp2Cn5
tF+Nvvlc4032e9sGPNRfJ2zcrIBiI2PCdf8nriJKxNLtt3ynkO0OJIDv1Fw429++E1o+A0D5w/aC
hWGaiTjfK362HNh/o8En2PvrKuwNiIZ4YIJdhz7W7hUMeOTa3vCJ8Ceo5rDOuVX1kyph5P0nijfD
Uem9yaQJjNOU/Uoud+0RpWeFvPtW3MkHvFlOp7B0Yvf5uCgfCz52wXHJxSqC4agw9anetmy9Vn7J
HWbHFCELgamdT1XIg5RZZeHtnThDrnyLMvkzpLcZjR8pYFO2Z794PsFsQ/5B67nU7xdIF8w4pyGC
gdXIwpCgXQOL+FWvVLgxB20LOuHnLF5HscjY7cLwGmgZnkHiQ6EJHadgvIUA3q2hRNKT3msv2n0K
Z8JrpMP2/8yezjAXZtZ9D9sN5BGk3ennm68iZ+ahbUdy4hR0gvu9wldJhKAaOl3ocNMLa2TqJcle
jpWPaq7jKHzOvrz63wbvkQ3pwE3wE3VIC7Q1/tbcvwyNbo5Y/kB0qNQtnoa/Ld/Ax1SwKO2ApGPv
Q5xHZeT1S1Eg6uyxbG1eOoL3NLFKsMXEaOZaCdSBGSIxfGC6gO7clkwFDOCNcvQ0i2qBtzlXS978
iVf6y941zA7lBYo7xHwKZZoxCCkGxbiD69dH7Ic1h0PBqjeNNKgBXThExc6zl1Qs6WMnhMFpect6
miorL5Qfmri6o1DKgOoMruY8fioAz2knVNv0YHlVLkY7LmDBkGpqd0m+Z/5YdI5/wq1O4MjsK4uA
n1GhZg5bgNhHJKNFxpecRCdQ75LOncrLOV5oBi2VmGTUrfBYB78uWCDXuqmNAZH8SkGQSBemZXnp
oXirSoHSFEaWgcrZmT1LotvJu3toqHexjTfYkO+MJLNy/+Qy3evwNm/QKYK+qe0FP13GjRRG5ULg
j9c+ZcI1RvMvJ5hyDjUCWAsFsY6RmpVcw89JszrYrwpJwQ5/RHG9qhiOEe7zZjcIXHXFPBnsBJaa
G/uEVDkePP5D5LvXY93WcBfarFt4tyYehtKE2neeF5dCL7F3LaQ2qyxO91xqDRKWd2cNGHuOCLmE
dy2CKVy/DEi14JMvCt24A/8t+3zGSuFfyP1DyorcVDZ+b9gcmcUQ8aX2p+NcKX60JlUv81p/ivLL
5HRBVZQjpLG0ANlBR9/oCnnn6Xejhjq7UMw2HlUupwQSrNfTEMLf2p4RzHoG6Qp2BsukJyQNjR+O
gtmBmdYijUpOlhiHfDcz1YQebUFJc8i9jcbvf+YODW7ah2qYwr7zYQfdrCsTgoljNRelQp6SOLVo
8o2qZwmnBkFlINSrm/TCRuS5BR45EDfs14il4LY4ISsEFs1a2s1z+iE3n4q7rj1Z/LLXYDNMS6ph
9zK05Ar4TQxg4otSaC/1BBAzDZrU5bg6m2S33K3aJymoREzsMrs7cX9bOEocEtxMdp719Ii07kxN
bn+w86s5MKGQPvPl3trPAepbkeT/kdg/xDhZXFfm/b9jZkswUeGJSvTYwomMLi1zHZePAJatfJgs
78/ueBLwd/Bht+XxgS74FUwnMyjGmJaYkzjA4Sk6XkbJSpR63jKE/heLwQdiUnJBXMHEIYcqQFS2
RToK3TXEDaJ5np9icEco+xb2sBFJ3uIbFiSl+aSOc6891KkSE4yFFRhkQ3r5CC4vlcYUipz7b/K7
+uS8HrDoGodj16G23YUeUXXhXeaMiWEjl09TVXZyW5c6p4rt/4Uzuj3gvQ9YqfoBv2E93FYXsKXv
I2kV5BJzwOHUDPBKnTl4UMWs6xKBaLHd87jPAzDjXCqtcuOfx+wIO75MHi8yJydupxL5MScos7mO
YrtgdZxn3LZKNOPISFeJrZclbWlWJqh+RY6AoBr0FPx9wPiMT9iGpIj7trYSR7xoL6QWwKmSLip9
StW4B/4czCAs7fn813yD10QsR8HjMdCFrivZyxrFH/B59dJiuMzhKFuldVHtSIIiRtoRtp5fTKw9
qGT8aehVQD87z3mDJqPfN78CCo+MC7iRaQMzphg8ITHRYps260RZRk+OA3eP4Q3SRa6VS+9pkDHb
xwwo1yAtM4NaSfHrhXAzErCMiSHxW1O//NimRKe03ViiBNWFa+RrOHRzGu9/9gGnEurg8Fc6JSjZ
sjo7QHRjyC7wCZErYRh67rvSNVmNr+kCqX9rYo/EELrbKDU3kjsoO1iI7HK0qyQfvG8AvVv1sLl8
+mL9qWybi3KJg+cnwKYPkEfUw/WWIupzYgmin1BV44eWJbn2yYa7Oq5R8LcjL4X0l/j5+Ly4kgWl
DVlL/XcXJxXIQHG+yjM8NbyH27+nJ4EtAvC7bXVzZUK/6v2gmT9QFEjgi7Cu8RoZLJNyWkl+uVZZ
kqA+sUZ8q3da24J3/AcM0nETieUrMZHmNf5VUW+9wCDkGog3PGStQe/zVPoshsAKMTWm/iHNykD8
hUERMBlNf8N3RGX8myd40gNT7O2oQpAvEZg1d8/Q00RRhBDIubQaTMN0r9ANs0HZwYzaaIXihHA8
mjbIqYVmm3W3gDvzYPP918CNlSxUst4OJTxTd0eEBggK78a+PMp4ePILmEIU8AeUYdiNZCTRDEfp
/oQfGiztX2ddy0qZNb4QldCuord3/b+ko8GDUI90OQLNPmum8zU57VRbGL77fdbZgo31gmqEF3gb
9RWf5ZKiLdq4a7LfrIuR+2MC5d+H6X0WLqSeatMByyGyDbjLZtYiAr51XRsw18kiAz+MlfAqwAK8
75SuzHtXMc87VXjU8tC0+Qu+DQ5ihD2Q/2s8t0lXw5eCBJSqulgu2D37jF/Tjmu7JEKsMRqfmHND
/+Hxp7NgyCuqT/EqLoI9rO1ml1MB05f3tUaOFE/oSVAOVtstC5EpTU3Cjb1GQIzxhSPrc3Vu9VBW
bmRIMtv+PHYOgNeKYo1op3/l3LlVjahYOdxK9wOwVfOtKleEFHTpbwoGGcuJ2IlQQ6qYdt5qD3kP
USTnTh5NgacAeOhAZlfVZqxBN2GC15m8SQcDwAys1c/CHNgsL2CThinSlurwNMCcxF9tzzVWAW/S
gAd7X11TpJEdL17A8yG21iIesvP3ju+yyUgAoYHL1S85OFJFx297rkwCRsPuVRFrkH/kuAobsa14
hlNlP89Y+xBj/NN6oY2e4U58PrEgE5SPvpC1VEOSwJslXfh94CRU6uGdYYevu4F6oB+ANYJ7cZ0T
pv9VeliPxoJ5IhnES5Te3sw35zkJTjrfbNv75iLS11sItSeVok1y6WkL6CQQfMFI4o0gPbGWYVYI
u2PHu72TNjHEYZX5upRq92mv/DO+loaNiuTpmZo4FWDQqC5ymMzv4STjCmtW7aFto/5+qwwd6w19
x2sB/H+SFR6Pdd7lj1SGiCK/txYn34CcFwE2ut0a6bX01Z0iT4f1UAuHqU1UREPKx4t1qbi6JkI0
aiFmQPc9jaKjgcICRMKvEyg2i8C6DQWfnvN7wR6or+CTnVgWManATQkCy7EGBokdVA7l64Iu+mbF
ylmeHNA09Lsxx4cyBR27POZ2YjFvAnRL8qbUjF4Nq9i83rPnS0GUreCOVdnWu+PLo5G+3vaE8u2r
6Kg76GmhaK+UehvYgYCODrxbMPvo/5WEdQPfBOlyoHaSgfNUwruXN3U6aTyjjqDTHvFlvePWJ1Zv
WWpqdwOx0n+2PAmvgCsFvdlWfTLCXfSgmujf5rqzziqn+/nY/8i5Hb6xR18tipiaXnXapQVa29O1
fJuNOlgNlie6anhz4FCFLSwNwhpreT/3Xsd53z4zHxpVOLrcCFsSdCTreTCmATJZL6e7akiMhji+
MdnWe5nYJjDNmfInV4Eafl1MpUTvAmTrbObr8H18TyJNvGzoU+xk/iMZkK0clQhiu4iCiORlzf0+
onxTweZAqJhYNG9w/tV8AdtQ1RvWnnxmxY2Oo5PWMjQ8YYBSgvrsv3F8thHl4VhjEHVrWQZ98bqi
rwZZoOiYkDWCcMGSsZSdjgl5UttaCsDj0WHOFX1lPADbo1zUGZwfGak2uYJqIU9S7m7nCimDPl8h
rUEhnH9Hh+pXlVpiay6+s2UIUU0TqVmQjsw3J5uzzQ3oDWmlatdhDLUm40/JaxjR7kzq0rY+TOwI
8Jz2iSikghy1jOlUkwJCDPi7fjmsMk4UYl5DCbZZAJUiwxKrI3kEqbHUvFItO924X1W7bLhpxznh
5JCt8uFUTK2dTq1Za9GrnrtpRVi44C9sk9mvI7oEkbbHqBwhe0CtIexYJ3Rz5BBZGW2Qp2nFPYPa
JjzrIRnTpBAN+bFgvbNMe7prwLgqUljntHQUiQ5bv7c3ChxxztltdM6KShrXQmHUhjAxyzEqfWSO
QrcIRnP3qxYTixfKD/oH4xek8DFdhN3xTQuJUh24TYm5nVGPWOcZN5CrciV2Mgx00TB/mU3E3Z9S
+W091Tir2NBhe9pCl685I/blfHTshqdOYZrnrw8DgZzCDhq1DF6H6J4aSueBLLDx6atWyfwBhCrL
VrCBtsNi6Gw/pURwX8zFE+1ubevdWOvdtJx/9YxoFo33KiBUcZhKmrMDM9EVOl5CLNDzrSXXZdeo
N9K5IYfrIp9pJovlB0VI2SsH/9Hmy1Eg1ApVPczKcEDH6gLcD7yCn1z96tc1HKqxDZw+zOaHQEef
AcXlrO7yBRfWyhQvmzZI6Gq5uL0vpCPzIQf1Vm8UitbE1DU300iWr7cp8y3yb9xgNA6jN8JQyQdq
Lk1g3pzlNSIuUO1N5EIfifL9fhoek5lFGHPblJbUR0sX2Z0BTiqV0OhffBRyWqUXoWnjLaBzJ3ht
AFpnA7LNrerFtEEWyRUmm2lx5sWj4skajc8XBEwb/oWhKVCX/r2yKAcoVsMom+QFuCUsaa5bFrTb
diNo/N6A4zE1VjJBm3qLtsj6FiP1qX6p3vQx9q1OLknimdd2MTFJmWnI6Kus/5ao89uw6+fEtVDy
c0GjSrLziPf63EZYQC4tRryqETodKV42XJvv4oEd6i5z1wFjXBI4vBd4/AUf2QL1jDoXbkJS2wQc
qT2Sdyaj1ZYhqw+GAABzcQuKURVXio5UNQtM7RNo4v0JTW6qIZy+jMHnUbIA116HA2MaZsO5fFrL
dNzJ/MARN9rbCb0I/72EKqrq0bfzOQzBx9nHqEEgYApoj49TMS6ZVA2I24C1QSDPTS+gNThj1tVo
aVE7XFINI5OwKVSGXJoh+FR48ZENiqcUY0ZniO0I/0lHOYxLCea8cT9f73hSFU85zpaQk7a/0whz
xTODr6hrsIcLMWb13ol5nOH12WoV/uXXzPl+TKz26nhHqTMc+lLEZqXuZUuFGsnKkkFfDBmVR4Q4
F2qh3w7RS0vH60LDg7gX5GiYe++Nsl3rtu+e71h91+kZmWXxYNXW/+iYuRw4zZ8LhvzZD9po4eb9
v9ofJVnYcGYSKfNFPsl+n1vAzvmdOSQpN8dF10slr7QFKjqVDkKrMtdYa668ds+LTU0noVrsf3jT
Dlw6zvxL8sTLZM+0sRugy4G/TQcY1oyl3S1NqYWI+UuCf1TAt3Fzo4X9gQcZb8zybUCyN91rlDaf
DRcvPj0DhJXCby0vlgxcdEPOAjxccni3F1LVxORrddB4l5vdgzw2pznUJO6/f300L9q8g0/xWTOs
JNbyAhiBuFtehbgABcIPoji1T1/u1+Hxc/vMs2Hs/+HgB0E2h/LcDtam5yTeVPa2siGs10JxHt5J
DJWI8JmVGpyCXK50FMDUYFZ8VxljS0GHASikrjqMfpInY5gMH9AqRZ8quNM1VBhFzTKp90ZNqhBJ
WwxsGU9LiGS/mG0bzLl8ZMDPLKUZNEPYIibU5VplfS9lJWyNj6Uv5Py7FloLjl6VVM/ntPi/hc5A
FYoHujXHt7k6X986Wk+/gyM9ZS2vwtykzq4Swr5UVAOfNVzLvxd6jLr1qcAW0xdklR0O9kwiLoj5
8AdRW636kgmRxlsMu6B4+Gx0u9OgLTsbj2jHZVyEzHUnZsA3bZxxxLYHvau043+4j9Nj7umRKWDu
Ix0191xxtJ85CFWut2VwEfG3GIbvTKR1DZ4XrHiOdkeo+neQTzfd1tu9duOKT4hOv5Hd/N7KCkrl
QudbhlT2yhXh2C/vgLB6lNLAHJnXCUTSf+LlmdhvRvSUoYCzjKObHH/tkjj9qIAC1klMMETdCYEt
m0Ispua1GDCCK1bxrlpol9YlrllFeT4V0uAK1MVWAgYaKRK7fHXt7eeVTZES/TxJnrMXVCkzMZk/
OPKwryCYu/5mT2Vy0wDzj9rWeBmGGIRoby8OX3L4iufzX32v9wdBByQ7e57bkmQk64AXHKJ7qbe/
asGlDcJ1pv0BPQUhj22G12Cd9Y4BXZno6YV+XSuEgMiPujGv9Rt/m88lbxGLbykO3fix9Ih4ODg/
3MRpYh3yK4K/MOL86FhXxnY0Keh94aM+wIVj9X4TJdk/Nplf/j2jfwr5dn57tcYFiuJP3IaMCaTK
0ckSSqv4aAkLSRLdEAuji5WuRXzbOV2UvrEP/SzylBGzQeZCNFEHSOH3gPCKDawrDwHdxz1V5xxf
shiHWz8k6EVAnyPiGWjPd6q/JGuLf2qPyrgtNjR6cHoqCFovCsYE3yFHdFwyhZWWV9FNFHPiIBAt
VO5iwlGCFqfsnSQ4KAUQFl+jZim8ewf/jEg/p+Ga1+7zCoLazBQtJlTooSF3xXikIPu4DRH9Ynvq
24Bj6TrtYqibOd+I9wtyBBq8Gbx6nQlDk6TvFNDbcEVP8oIBwTeOIfp6Srle6vIXrY7L6SbUJhr8
6tBqulX0upSCxOpJZnJHnNwb1Y2lXwkRs20eGeSKLmYa3n6TLh3a2plQWFZDRPkgfGXleR2Z+0S/
guiAA8YA+spRACsWnlkkwAq0W0/kiSV8esKRSiYhojsyropfMDRYmVYwh5iXyFT/+pT1wRTQ0C88
dXyN2vBXh/S9weIuviCWi7dQqREGvOgysOjJpcgqvrNqzaYgIbgpk7jE48wG+rLaksZn+G4bTgQA
ImXkJ2fFyljFkPqFLnTYDe+JVYaY4xHpw9JcebL0qfXeIO1wt7Foss9Bx4e4rQZ76TqRrTUigHNM
JL/bTjTW0VL+3QhSF8JnxC2r/pDmkWWEm7Nj8+T4BC+dxmCAJO5oeuAPgaQZf/Fwg1pOAFtAWYZh
N9QFeUKwWP8flO9kPiIm3WY476081zQU6V7y4tswuZlHfhs7d2yhk3uPwZBoXzTxYKhENXmwCBMb
9GxemtDLhrR6/FglP9HU1z+802ujKwD13SSjfCT3xoG+Y+dZMteDOHhz44R5CnZLy1coAN2tNg1c
pnyJXEr2mdc1vIkB0CYDjw258/+5Hdcz8oLR1RJnNpbPim9lpe3dfEhk6xPT3lii5kw6OitGNrw8
E/Vyfv9y012xCDaE1xg+eyvi7J3GJTD6dKD0xgwRfpi+gqYWTnbzWn2jAl4vEmem1VqkH0GOMSZ4
mn554ZD413UyT2ZBgfGPSS9pqx2xtHW8keITXgF0uStpzziJToLfw/piqVVdW66E2m8WtPb48OeN
BETBPsWMPqlwOh7JzgmcLe3903iAS36KZWZcYuCAMsjreoB1wnr0iQutWXkoRzawjQlYDwVCu7UG
j2yg3PC5xO3CcH/ML19z6edi3cLkysMZC3n8pCD25o54gCQWaftvF6aYR50/jrwTOPrjqF8FD0xq
hl3/1x2M/zKzkSt1DkW3gqoopCfzaMVkqmiP7lvRWiv2VhRta71fu9WbJmfiuBth6W/WHCrr5wW/
FPsHuFY9tuFmFwvKDJFd1FTq/liMRFZDPsGUGWDRFHutWdSec1nBlXSS1+P7aB2RRxTGL819inms
EPxxnCUIt9GnYVDIEZuwaRad4pD1eVRKPhzg6zZw4KWsubljbLUmvU88cY831E1lwEMKfdJGotd3
FBWC864HreGdOi/vpr6AW8Pk2r1966QGr2z4k1uXawP9zLCMDQJSSTKBB2v/5ujwSAxzh4U+DXH+
Datf94N/VlaHKZl7QIMysqTQ9Juoqd9zZSwAsvEMddlShwNgAl1vAH602bZFEOiOEFiAa5ib9re6
QmbroVWaA0hOBUGY5na78ry1/Ab0zGpq9UqgQKYbUEfk3u/qkh1jig1K9E2gSFL11DPleBkROy5R
ijW/ZXce0MYSyTOLg8tSgGBsCgcdma+YHnH9frUZyYDnpm9cuJq21o1vWHzDiR0sHfjeCmYht2cU
hmlKw+57fEY9qvGJAoCCgiXOmh6O/PBqaRqca6Z/20j/mU1/ofM6JzdDz6vh0DP0Q4P5YJJaKIWH
tB1uqrGtIK62jITs5HP+UwuSq6zwNMawx7fg0lOJKS661/D0V2r3RU9/sauwTFcXvdABgQdv3vn8
yfeUAEb7IbXzTVyofuV8ZVyj7GlMxqkYkhqqhXucoH6f2ZiSCfjWMPrDL7UkPwEzYOW0x5J1sspM
4KLpCrOYpMqwee0CifHsIX/b6CQA8VECbKMYxDwVdxWfWhlwHXS1+l02/Iw+5B+LP0TNn9udWZrW
V5EYomzYGLbeyj1Zm+IyzR4a8mDfV8O/XZ2GdmXr48GDDKomURJkdUaj64pvj4Csju7XCShAZ9qu
kbi7pnOcTIYoTbdKe0/THW5OIxQ0oEizr9Zk/hsrkjhvmQRBBnVZ2+wMdzlBAfrRsiB7Cs1PSPfM
TMnOiWVTv+MJ35RTsWI7NhM65xKLFuU7fBn9Wd4XgrflDzTyvZsQ/N7IHHnReE8/KfuRcXAlTZjB
5iDV2Jif/9vup2yyabIJIoVOF81M34+aLLuB5ADD4oDKsuK1+zp2cHFOFEw99izJ1AShEpX6DlEM
qSD8aFDcKCx3C2O/HAqjMbVWy05bz2S0ChB3Vk1GBGUKp6Fn2iEL2cLQmvIRuZanFwlp4pmZ6vV2
vjTpPUmE9DAJ60TBs+lcZCyYpqOLPUTd9W4pupCbhsm+ZfiCfaA5pzXlF6IudWAj8oVZ3IYZG+3U
zQ8lDK/3Xfk1EEEqD96vj6h7leO0N7bE97l4GcAseIADP58A4c8WSGovNLtR9CLZV1QzJTX3kr83
3xwSyIWUMNWyTqfRynnLDC06556fBo9z99d8ZZBfedJzRU/AyNLqqIq4kJ5tGZ2cpRChAnDChTHL
mzvgCMhe+DyHLXMvxnedqwmcgYoFKUOG0TnGNamCL0loYSn29O6NBBTCg6EvJ8gvFZCGw1cbbqgJ
VXnNvm+qyNwz8jCmAt5cIrX367Sp2HM73r/uaUaRtMnyLpL0jS5aFLOOSprhjiO65ZXKbY1oXabz
5kOTLKQhF3w7iW17Uv+bXzGZrGNglhOsbO82GyeebUxZdmvMYbXLOtIZlEeqwz8aW0Eyup9flAKj
QBUBP2EzJ1GmK701R9NNAF6QGg0j2UA+TJyXmjocbqDbDOTgcXGOnG/YbeZnKIlnd/QYQRwWuTjy
O4VQalTls5rRDfW9yyCZiVR1yOVUxHraBXpOAdM2qpidczCcyWpw+bMTPEFNa4AfoaIgrLPbJmPW
vY6hoZm/qqRrGdE31yXkBnqNXkIFUnbiQNm/oLHeGa+0JXMy+tP/xq/+WyVp3VKHSlsTMZh7WkBj
/qhwNeSZpXEkJ8livRIeWRRTYNdrqzax/wBQ96eHd/vvMSxeOkaRsXVIQFqEUmb0bhHtaHojqjtU
02BPCC9vFyNYAmBi4VzyqAw5yJO7TVus/gMpg9Q41VIdK0jsRvrcp1cRlMI4h1h4XxAqbfrk+OZG
8OLH+JfUupw7S2ae6pz7RXa8wK041Zh+0wxx/TP9tggDqIP3VIrEH3UK09Uvru4KhOefRp8sJrLW
I3eHF6q9VbraDfMUrOZOyL5kyA2l1JWX0T/5XjSeNDk/kK4gPtRo7iRO9TvAzzbIGrRLY4+9N1sG
Loeu+TJcp5kXUTKNBRX362q4lhBqCmNRbPTIvxFKHCZsHwtaDsHDQJrS+iqpF+kLT8RFBRtq6i6s
j8/20IPL1nN92NJieBtKG1QOvqPdonpYumCfXCeTJxUHfkxYN0ZMjeVnDSmzcOym+0MBkryx+guR
ep9w0C6SStik8Rwy/gh/ZzMcpBp1vgSHbSAnPv/59MewDOOW5gblNOpTRwSBbblkOAX/7ORbrGde
roujjjvwEUnclx7pPikuwCw/VZZPC3/aLNskvKJP+tGOnpjQScaAPKS1w/aH7DAg09AXw+AE5Jd/
PuWCYhEwWMpM4UQr5Ds7SHlg29cSVXxGDT38K5hD//oeBCfNZUGQUdBfIjmURyJ4IEtFi8SBdmE6
3KgSVqQRawdtVd1t5gf/heS4GRaJ6k1f8ft7zeO+tkA3SJLiB2+sCRwWDDpugwNPIgMCA4L6+tZ1
JnSvkI6aHug0RDBOahB6EWSAfxY7OloGNT9/i4p5Np9yDJwo9XoRaNPuGz37Hgpj9EfGfTv+DXZu
u/+ulFsRF3UYnxTMMLxN8raarbrRHAgkGElFoVde/HrFNKatu8spZ2kPnfFTHhHtAS6U2f8ZXC02
PEYPTWPc+bPhZBiVAK3oUKVjO+dVPvnb/WzRpNYCm+FEkQvWHmURse7N2yIyxZVSnmsS0JzIq3bH
QhsjJiGIRsY5xITFDtsUHoeChlkgTMtPv0nAeDqM/8b9JX653haSsyjpnc8SY98NF5hFm+7A+GPB
9A6gApnemf/tlVljeeQY/Vk2SPywVqR5MbcoFeLeTm6pyIKHyHhhc8NakAQM7MhCHA5GZpCPTsSt
dCOlsHd/6vBgzuHllJvN58ThKzMssgIOJTe2ein+9Pn0O/GSEhvumUFyetUg1d7HPcYhYtZYA/BG
5ItuMwLLWS9WY9wDBzv/ijSfiiKdQki59Zl2QTpcG+YqL97JZRLwsTwh55tGkpBsQ8roOlGbTr8Q
Wn9uTegzdAZXBOux0lk9bOq7DMYbeNgTDHPcc+R4p++RWR6ytVO6Sfi4lwY44Zu7hgMQrg5c0t9T
DSSSLxIs2qvaShB7dgDUgVvmdJmgzz7V9YUkgNVV70vWtm+/SIKHgyACqzuImPyF1L8xXdkUeXYq
wzCZrtOl7oZoJY7dzuwjMG9UAkKxcr+miBJbwaeNo8JrdO4gn1Yw3TjQJdaW6KJlAkK9x6eMuihH
Fp828MIPDIXA5kr+VDVXeD0MYcWt1yNzmqZPB5vh4mUwfhVTN+HdoAzFVQ5DkjrgseNHk3YZvRvb
7BKOgiEAvaV4fhk9Lpl4aNZfW8IXyNT4eD5R27Ec1NnQdGmbGj2tKrqDP1Ag0KGiEQMHDRo75mcX
GFgtICC70O9yL8B1a6xaX+ZA4sqG4XUj2HHw5SRB/Mw/W1g/ub1t0swkNFc5qNpDTyWX6nZnD8Ie
sV3VVdawSI7GJWtZNWJcYz2neb8N+xeMW2psAy3L7nKavPS20ZPSi9Pk/iGd9qEXnuHiUevzClkf
YdzlmeDbDORf6H6vSQuC3jlCgs/Ptp6iSg7hIbPgqzTrlax5BK31YKbZiJyc21oJHHmNvH++ThMD
DWjMt86M/WCWlKqYdvEkggyoynNcTVYbh6e5riAf8ALT6EMRyTVS+3arGN+k2tmQ0y8q1FHPm1xJ
1zvD9iLe7fa7tln2VO3HipyAOBwGv2svs5pfAF27HWI2Hv6XbGtKmPWCG/c8EJXKNO3RzrsH+uh+
CvJKGBgOR6flTrg+3R/TB0MLy1nSnKmxh4RlILcU77VgpXvqFqxa452bXrM1d1RU0sLOdpRGoT/k
BYUdNsnKv55eVXc1xyJiugc2AuZylf1OGh2FiPb2bPmdZxwqXM7r+oMa6QnhJURZY/kH2206TIAp
CGg3BdsueyznWL2wkpksgtCaWS2MpleJb66J6wyXz7Uqo/C3DXj1OoJC+O0u0ff7b1KNtMxhcwpq
6x/IEWs5apIKs9/Hcuq3IKrfYSxOVg3LcB3jFtjC9fvaEGGPO3tOrcWsj7r7755Mg2bpIfHTcL1F
IZ092DCVbihUbqfv3eUgC94huAhjoYSqxJhLFY5zmng8XNgTH7CijB7ktUexTwHA4AUSH+MILc0x
kJk6q7NltGU/pXxqTOCpS1GyR0eE31gKlGvy7EkL33LNUm7Lxg2m/k6mIYGHhJ3LWl0dy4YWtX0I
7Bq7+QSXPn3/wAR3IWHDQpxOMxlqz4riRa7goTNLmd3q8qR6b0tPJNyBNvg/P/4zhb67CEdfFRTl
X4uODOji6g2hWg9lOnZ4zMf2zWQXoxzRCBwAOIuj/I3tMAVC+xaame5+oDoc33J2rxSYytLZZ2L0
NAH5Z8si5InwP85R7Htz6qksbfNP/9Q0bWwOaO+j5oF7jopb8JtYT0GVVLyPSxE9/PnXmsQkCF3D
bXzYACuQ8uwlD70F4aGaLeAWhOCwkQeq8Qfd2pRzZgO7vyMbCqGrgXC6PIvB/5EmDHzyoqYoWKy4
b1F0iL9+EgJYTunCbfVKBhN6W+XcEHni+bDTm7o27Yj1maZKyQPABWWnAbYXqJP0yvhVkanYoylm
eLzkUmCUjLK9vOQ02EeOYr6JpWgOB7ai839q7dvfEWM6TyuRDKhXUhBrPSKRQjvjxSILDVfTPo3c
TtPxOZEzLXG189YxPQb95l5IjEq+JCx6rO1Afp+IWMTnpwg25msdSyGdIFM6SygMFCTm/pap0wy+
zkLf1KUHRiRm/NDNZZ+OPKytW2cxFHdvn+UkZysJ+Et8qV64b6HD19LEJfRve1hldFL9K4RQgcla
m5N7fcZNOX/ih6YDh5kPe6ogadtPRafGbKN6/df5lAw07TF+l/zd9UFTflhLv1wwxGeXDCUYV6Po
aefgLJjkoQedYH39EZUVg+3l1VOZ+djYbWWcZa9taxM5J6r8FwnYopZef5dfXSH0AM2mD6xEVuZX
EUT2fmLlMmoKUOVzUOjClSII0Y4qxin2CCNNKG53GUI7DHAyb0Qmej0G6rdC22QPkW6AJy0P4P6G
5QyFd0zjBTyxhjH1FB2pilmxnX05H0kKffw8OZ5lNLA/quhGrK88D2VgiztpyebjxBAnEm9clP6E
vW096xAfrlVcV+PF9He5uB6kceKQ8CzecJjSeTfunIscVBIvMRi9HaHe18br3GE8FjuIIMl09PpK
Vi1rAWIcOLEuO+kM8bDaBphchCAtB8xo4UIfwVA/nEZ7wsQh93wvEBktl00FEh9BMlkTFJVVtLi/
Ii+ittrwnoUPcIavJtvv02cWUrMY76pEW11xbr7zNm5iZO9f+KLDcao9LyRMLgGr6onW9OxDUPg3
dxx3FnyBer6F/GC1p9gSUGSfuHpuV8N89p1G+5PIZVghy5sBeOkko1i/LlKdgzwOfgmSM4kgr572
MW7s6GriCXb1bJi33TY6b4xoTP7vo+X2xpkHqhz34Nmq1ipzOrreCSe/0dnrajxvKidC9hHPA0bO
C/OaKtDHYsvq/Cj5dtF4eH5uMmjZ33lk5GHAivFtlkLayefZLxgb8+1bmIiS1tfMqCbdTPapvn0I
86ehJNkWmTNwTnuN8Vzi45myR80s1AYJYxGtXGnCmAcC2Mlz772nN4M/5P9ARvC71faDVm97Lman
2KsR2MYqCdkIrlUIs2iFtQer6X2AlasxxyqlIy13brVVcWvhrOXqSwFbRuonzREdc/8mLzPuGjMW
5aNC1RNyECgQfTQaLvgppGkrkWB999gFArAeLRkJcaSRc/ALkBT7yOjYx0f3/YiazDxnQDKXkU3Y
exoBRfErDDgHXt4/D3MHF/buUoIvJj3TVOuAmVFWCWYo8y5NHSIV/wj/wvfc/+oHZR/PRkP/irR1
7/B/7in4una/nnSEuALl+UVKLnbh9SEwBD1AObTOUnWhxtbPqYXf4hvYAUUil2HADUEfaOzEcr2a
cXpd/5G0GfflxcZURuTASIPpclpvwKklHM9ChhUoHwPUumd2QKU2+yjK3W01rje+4YbKikqtvBjN
Km31jPACKA2XZ9txP9kQiQZi/w8PZs4EKLmm9UZX8vQUKZE2+1JzByWGthhVn8elB6W4LuvRRVBD
8K2vcgGBEomKii/AfmXNSuLOmri+dJL/xx7cmQFSkg27xc4Q1Dq1luFWsRhwsZbYIZoRnAt+Qybx
1P11zOd0V61YZKdkfGhSZOu0Eh1BEOM/KcRXH54lAAOYEGoZjtsZU14FvuAVe8oURGCEh6EisZ9K
IC5Py2L6fUKNff8hS6fzUAlcCMhy3wcEt9KllLpaXM1PfWtQGA3lvouhnLTPjrYtdmdUA6OSU/lu
KDO9XsGUlhVdAx+Zrol9s9l33Kq8hIhz80dgl4B1NuHyT7M9O0RIUyufHFlL2Sowbuj4b7MF3sSp
q7GAuj+BvrFPYD5VWw4EwDwhCCW3JIOLjeTep7oTvLEwpS1LMBT5tX7l6C7vhr2n+do4yFognnS4
+5bsqqk2pqjogn9+mAgJcISz/XKk2QgQD0Wz60Dkiw7SnPzKpQ10by5oTGADicx/jVakZfRxhtIO
UNwYMfLIHHBJb1b2mgWNn3Cf++s+ZPPOh095jxrmswLhGu74C0mT3urvKtlYG/0uBjV+ePSszWsJ
PMDfMTNNEkDp5hy0fOiTjo+lOuPu2qod3HD5FrgDf1xz8K/nHbO3JHR071G2VaODQXva1M5j44wN
IIiGw3a3kKVkZyWltKurYMTP9F0t5KehapfI8+rKg2nyT0yPbhGMvVoq6WwMHUv0RYVMG7XpKNJg
ZXvFhHJ/HJ2qGQIdZojTpXROLB75CnPaloRO4vub1JIrvBDkozUOV6y3RERkQJgLWG5o4FZDa7pn
FnXF0qYYR9tZMPnwd36iBEolHOZ/OnUs/pANS32FYnOU+4KtvwmXXFUGOjhNuiK1JuYSsuHf9PCn
8oaQJKEXr9bE7xLiTThClSrZKDfnX1sKH/XtrSunwxz0Va65B4O3UyZGRLFY3TsOEeAlzuJLlsHf
UlQ5Ow1fs0tshQtabVc3UoBiTdDhxb5eNXXqGVwCbgVtmP28Gv/YBpHbNqYDqxsnMNU2QKs0EwNK
jRsvlQkLJrmw+2yy/tUEGDAb9LSniNZiAcWFLv4ZnvQUNTcrVMIUMrwE5+5yynCTJHpEaPt0NmJq
s4zCqONMVTqIE/gW7JKtjN5ZDqbIHj9klEmw7RaRvDrW80qwy1mbfBctTEOEgzRWchibpVQahtHB
3VpgfFaxJmdd32SVSasg2rYvz3JpJcMbSYx/aTv3XLhB2jDGWMlN0V2TH+BE2CIgZnYyoTGquUBp
y4vWhkMVNsa4GcvbHABO3Lnro6U8PpzSkAlaYKuM5G0f6lI+4SOGpwsNy9dfuS1jkY7rIshlDpYO
6Djwyxt3bse3+N2bZqvWJOEehQLoDG2UIVoKpzRFAAe5jYahwdYDhdAeJ34Gx4u09tp/cds+XfCc
nYMNIt3SjtpcA78muREguHjSJZ05GgD/KtF5n0fQ1tKxdwLvOOQTQx30ETQ/yfO6LSDPZiX2g2zt
+u2nWdujbOynOAVT6wjN4LqBMeFvAxuARVGDs0S8oqazFZ7yZGb1+8R33w6EXHCqGNF1/IFI/gt8
qIngn1ocz3Up34KBb5KHbwlEh25D14ATmZyaNzTycMMX1YQSZVkOXcDAV4iky8Qfzn/HluIbjYe0
EBsEVkKooyQ7fGgZ3wOqEGanH9casptNlF4D0FaGDRmJlMIX1gzUnaJSTzap/JSUKeLSd2TbLdd6
7d2gJr8OkURueWmSDvpNzIJxcopciRS3Up1L+SP/Ou0gO50C+tZIir84GwhrkI412QZgWFRK17bN
Cg/x7z4bH5E6cxpkVDQKbC9DjZXtJHbKpR/5q0QN5hcK966JNTxDi3l80CMLsWXuzqBT0wa6Q2MH
7rmFCIhv7uk3cLTZzJwhA0R5nXS5FWE3ccZXdm/XFbp5N31tROcoZCCN+Sx29etzOMQ8lS6/oAZ3
nhzTnqU//Bu5jkYIsUbqbAkfjTVs+/XRGidBnfC8ihSUow2/T/OcU/9MCCzVHVSAwYuzNDvRvLkS
LhuUSbz6HmXSHZEfSq5ge4VjZSbqPaj7SP5wSYb2iUisCAA1jXVgHZEy8drmgWqV9m1D5gu1x9ZX
8tJspwD5+t84D3Yqiqr/OvyGlKyUgTEog/510cCbde+0EJ652b/2If+VGJWwN1GzAsWfhOfF/3ot
ScT6UX7N+hR4cE+fph7CFPel6a3CsO626TpL6Z0+e0tPi/YZqKWvSZT2vJl4wg/kbdWmIAS8G5pf
9+jUG4eKpcdl65+bceAr6+8pnGwvV16ek6ym/6KLjZ3sqPVXUkkxDvv2cHcDXeh7zDhz4MW2jNjA
oLSek3FofGpSQQY9Veo2r2d0j/167dKuH6zuvofodMGaVe8JteymLCIPTjUB9rwWWwPGtBYHCahq
dwS04TmMspNK+jeDamSxRNuRYD7EsN7qumxjy72zB35yu9GRtFlh8IjQ0c5Yd6fPXmgxg3Hm2Aep
NJngOS9FK1wXGbzeuROX7Wk41oav263nxZ6J056ZAKN/06VI5oboNwHCuu23VvqxpviPMaAg4n5C
sIRkjqJT59X4s4d4ro/aIkEkmRs1tRi7NIibS4uztWFZQ5KiLevA9iplP/eAoNOneY0KV9QinErW
ewzjsNBsGktjI3ZwDpFZf3nElOWxxT7qnwrwkKblak46TCYb0kP2+5XFfJOlT/ly0u5Phmp+d6Qo
vQCkGCz6MSqDnriAClav8JQlELwGXhd2O1Enwo8Ryc6ubgY1pvgmJ8EtY2yNervKOpi/1TmJUB45
1tlvqCJTCchbFQbhA+6bwivyt2wAGp6LtynzIkQr75kR9/4+HM8w7dCVIC21gJuNBKiNSkPbCh7g
7r1O8kDNTJOrGacpQ64MmfTlW458DMVyJWe9N0NB0FSIC4cRaYg9E9uTNWSsH/nVo9W4ilr7lzUK
S9HUHKpGyVoPGLrGORP9bozq97JbbjTbAxEW22ztkJZ/KCQgEMef4kSrmGRSLfLUs3tb/wWGEpxA
jhGkNiuf+9VTq+twZqV6BbpqI5sLajx0gyQeMT0yMBkmWDQkopXjYzmxSdmkx/Uw3Ht0MgIA+g0W
Jmn/2ktwXoEvcF+iv4/ZrbFkOfOPqB/esybxWNI7xvJzcHp/5bDOF95kxpzKuiyhAp55kw5/mfWl
67hqFgvDDYqxpVZIkyMM7vEuHbDsxl/Re+vo6jaZZgD1bxkek0MeK1hQ+LQDJmXWh+x7XACyqUTG
Qe632blPpIPWN3C6ZYjthWAgM5lDcNpydc2Jv3pEVpEOFJRS7N57Ky9nMQqOeiuQo+icYxuoTSCQ
RChQa/D7vVLyB/FiSaQraivo+x5rh05J8oxIAFE9LQCwVltaDureaw9/pEQMp5YrogJd1gjtuka1
faHr5gdPR+SgR1TDUH42GLOciIyNQL55hyMrqPaikoANb5Xe5RHDUJSAZHn2t3o6QziyWJk7OgvN
aqb1bPAKXA8aD4V/JKu6Lpq5Y2j10/+AAtJQP7f1vlvVgmYlF1XD5wZumlnIHzCdyF01BTXkjg+b
gqsG5ZDVmYQJuzyrLM7kYpMUVesyoPlSKNwbR/GE4RelY5weURbXyPt41WCShgurzKwVIRs8zrB/
T1ERoYrDOEJPU9wPAruKiqvh8w6wZQW9vZohNPda0EwZpcE5dwnKsg1HcbINwf8F5/8L45ZjCNpn
T3See+rC9teTGjKezqWh+ptpv1YveM2AB64Q1ZZFucVvRusdPGKUEWXmsieW6uQyGpyj4jx90fdP
jfqo0nxtpexyeptZb4Zq8zTCY2+qPqE/azgi3qB6bymavzw1qYyjNkKU+dtHjhjdrQjbPKAFRXZ9
o4InIqlayk1cKkChaH14hbKq9358Kacvz1y0JfKT2SDbJ2z3thYkSXVJEzhbxifJt7iuun2RaSnP
EMleKAd3NkMhDX6pMm1iM2qag2MDI69EQKI5h7opq2XhOqtEcNMOB29wEIgtYnLgq2NDuyfiw6RE
VuS3zQSeCkTIfWYowjag7Sfz2iTK37n9cFbK/RYEoqvB0qqtOZi1LHSa18YsKPGJOuu7tuX+xBay
qtFtWExqNvug6ehTM2idt0OjP1onr0mVh+rk1javdOdNq3/YSKuHob/FsSvD6Iw2e2rWNRZOkJFf
6dEnMU87p4XVoLOiq5/3Fi3cuKeNT1iEsRCvielygOoFck01F9sMRk57Gd2hX0nJBuYH5GFpHurF
D1KywUb/bKoeKlwv5juolJKEEVtb88N4oQ0rQ0n3r5+GPryzq+y8nz4UwFLVlpdiYMNImvbQgUqC
s961ahYU4LGsw6bXGvLbZ8JtpkIY2zTsdkg/1PkKtUVEchjUjx8aQ0vNyveIxsoxDlXW7/v2+TUk
TGzkjlLFHNy3ycDseFcJ9CyDJcSOH+0E+Nc9UkdabawfuO/zFVNoZMSm8OhB8oKeG5EYB4GiwiwW
dgH2Mi7On0/n1hVeaFMNsiDpbqPsOZoMJ3XUa1ovpkYwbIn1Y5yTs8GEGW8mXhZvmE6FJiX+ss1I
ri1Lv7eP4IapFBcjpII7aFUw0Bs68+QAw1qpeBfUk4Rc2uoPxi+yObtWMSNBxWeFVP6Uo6EKm6+5
mGDLs2g6WQQdz/Y2a+QApfL2J1on+tZGXUKR1BiaWdOYEJs/nIG7YqlJUGDCGQIFjeOY8FLUscga
lKvcexrvaOJMXG5iyPZONOJou2YfEm783SWiW4UfQmw1cPFkU9pjmCZWsvoUQlmVgycR401B3cXM
M/Ghgb99iT7dNeJNPLkUuI1Cxs+QDShMOt9ikdgdx6qyfRz1zQQseQov94qausvaRBvD9lOaa1G+
oed71MgpYkPOwdUAnlQzlrNf10JHNplq0SEVCKId/IbpURyQ2V5BKu8G+5YbBYInomOLkcMTvIm1
QpU31NVoYjVCmn4oSLLQSdojm7PZGra4N51y2RpfkjcIDZ3oSN+TgoWQwRIx2Sfo3PcOwKrMXXrq
EaBi6v1SvNpmP9HOXUMoks+hI8GifWkgq2A+c46bg/JNbk2hfvcXCA/jo+7Zk8rKmwvH1njRjQTz
88LCY2Q7clS1x61STiS19RrPJwNsxc3OEFsi5EhISvuzVoE6l8bS6JEMT0n2oxHKIaepPcA2rs/G
/wgw5ClEbmhCPxgp/lpNhCeiUavOrrtuY1rPjd48gwfZsM7U5Qfp9+VAjEDzAcNanN2vtluicHOP
qi3EoSLxErAln1j05zW7cmvFaFk1pGgSFSG6dQa1hQC4gBD212hyHO1qGnEC+9HJESH+fgnWa3nY
3gt4CvtPiyrNJisP7Y9DAX0kgx0IjpFR8sWGRLCHbHLnQDYnh5LJDJ8ME9mU4RinSQRv/Oo5rIxT
QIisonJ4APdtV4VoOLJ+DcIfpesLdHbYXRsvib7OyvdagoHnszynoy2b5TCcMr9ssHnfLUHtTM22
Ugo0hbX/5pllb+i8dSc+VVCFtASBsPRStycsuJKHR6iLvfYrR1x7iV1S0TUEXg9c0qN4FaGB0Zi7
QIwmv0IaDOhedYuSduNJD8WOdk0uLiyWWoz8te8mIRJP/8IMTn3+5JT12XUzE7B/a0qO4uaAx4fW
ENvDhCKANpz9VakB2tOcJMyBcvwxPDt1wo5uC6eWPKbWi6KYSHXmiMqPqC9rJWRfzb9Cju5oMjEf
bGXYv6nUTLotL+eHqnPkws/5KbUgnQjpTsIh1qyEK2p1WRjyO7gkfhyjagGdTGarafV/yA8xxxQT
mmswGZK0pSKPSh8ykwjEcIAtoknExpTaFkuqKqRtjxAkZXCs2WnN8v/AhLUG2rbs+NjXqpYfT5s3
Iz2UH7wFjgNTO4cOk5QBdtujajShK7x5WQKUTwHYrVBmr2ZKMXdY09s2ErRA89WTcLwq6kztf9nR
h9uGy6r8qFyJ0anpmV3XW/7h0H4qxluk2i/JMzeHCkRY0QZyyABfBDDNF8Z77QNwU4K4hc8G/ZTz
NtqLdi7mZNuQjIsy3oJ/sJL9BnvQNJwXqcRBnG5p3QAGvMfriME0hMjMqW+TUpdBvRZqFlkI1CeQ
xKIqNQtxNCjWcs4ARGsn/sGlKBUBYRA3f4IIoxWFTfyR5gjl7Z034KhrNrJIE9Jt9+s5mOWhjj8M
YvsPiReuyOvPKZEkjQVH/RYngbQABzFaKCW4lp42S6f85WR7Gb92SOoUPxQyyP7TbJ1Z1aAGrXmn
rg32NPdUSW/xGp7oJQ2FLZ7TDkaS6/x5Hmd/9HRxj7jsh7tZKwBFeUa0BLy/o075FODHNaUzbIHF
/qnq9lgbQ7frDh3014qHmZFi/4yPQx5qzk7HUVljFpkb0OyQjudqLBxdgMFSRgR1fMQ1SmtZalVt
8v53k/ykocv++ONZjf/W6xQffuEFTAa6ro7evud57sUC3Mronppv170Mf9gBZvefJ8MdzlOdj+Ow
VfJJkcKoWCWO6pGYCfH47oATOoZRekeEgeBpio15gc2vTsr+VolAqYYtURTvRgCL7mAYhRPkq8qr
XTiY0EX+IsNcf9eDUas8j2X2549bAF8Wjfzg7mc01s/0JObGrdOIxVK/LOB6yXH+PuZLK6bgTMdF
dkpdEDmuKA6K3U8OUTsn+sBMjD53z4Tn4J/nfVgQmEOcp6jChAAo6hbqf2Ymxm3j8MladwZ7gaBg
gWIfptmuG6Tb802ACuNiVuGbLwi2Fl3pDWBkZjkqihEXyhGFcdOTl0sKS0IhH3iBgg1zX4GMqq7x
EYv5LOsdQM/xiKhwkAXo85hj+J5yW0Vbaz3eXq0MIMJmkDwTvB8bxYPs1AhUnZF1BurnrTTU/8eg
Qk/lh0izkEAERGGrC6vdTgS/AwfYlP638SS/G1RaE+Q+HFY4Z7M6zYOtEg3c8cus+QKGTij1VDtv
fP1sNxBdg8cOeH+SP6YWjDoYBBXOqA3oUGLnXNiBpcBLpaWb9foLv59pSpGQFso3fwvWHL7AFRG9
j/FsENM15S7Vz03obHIpc995oFWC3+KJlfA7TUX7t9n1Db5YG0wkL+70Gmg6nh4mgTo1rqddYU/8
nLeE+EXxlPjKZsgVuhGya7OwWgF5xngT+UF+rqdD/BvnH60hknhSx3kmwpcQn6SfnQkxNaaDdYg+
J7lZKgRfOXFXvEkDvE/LhduxICU8sNvUQRHUNWBuLzrx+KiKDqrxDvc1JNFjhngAEUfIyGu9pwIz
SWLguWj9LWq8UfFmiuLpEA24QCW7czmGp+538NAtH9G89vvCViW5giTPsO+WSY5vzkbned3S74K0
eCgrQ1S/XAqMC1dqvFSk98X4XQFAaAxpZxaOqJ2KAKBhWso0H64gH68cMlPxmsqyLLRIU8N7O3kD
/dOo/GiI9kXzyiR7++fQNJWgSquRnYqXZXhKIzm19o/OMV7P4yNbHrRZTq4pVLQpb/+HeEoat/+c
cp/RxCjCC+D8PV1vNaqTg3irBaESSwMNSSygIU4j0EmNTJaIzk9Jc9/Mft1yN9I4R6sKpzvDF5SC
kzvV52olC1YG7tRgY/QWGrkwF5xHZSPVa6Tvk7k/ZdHyMGVIm40qHM8GcXhNbukUGq9tlDlckgEV
F75KUL+CyNvW+oE/Vij6BKkwt3uPh1AO6/i7WjEMkmQLIaVytp0vbNvfYMQ+K5+OlxNChPml62bW
bfaoZ0vqKq3smF7oTW61kB762Gs9FWjC+lCFWS9ijFRDkR3wMmnoOO73la2iIxPzBvhAsDHHeDWK
/8k/BiP2P2HY13GOdreEl/8NmiRGtvTUU18/MBy4BtfLIRA24gyMkusKME/Jt5BotYFS75Bh48rr
d2w/SzG++e5j/YE0xG9ZDya/zBh6A3kcStLMzRbOvdiSU2Q+NYlISD4Q21srwBfZeW+MHi4ysYp8
N/XMwiSeI/w26yuwkHk1remsicNzl5rFPBeMHGgiwd5WfWF5rWuvXnbihifQJmOcwdgsZLyRkIeg
PYbu1kXu8pjFPD7TIa3MIbD1CX9qAN0EPAop71liobliaZOpWluCuKX5MtkT/gsZtPdAjdY238BE
lxxWZcCLZbFdJ88sh1FsTVkfiICoEGGH0H5C69ZMAVZOMZaepUi74QCW+ZCAdWY+a+zw8x1AMJvG
pb1/colQ6lCBXSM4BxwtavsjrW7BAc+heYNV2k6V3yv0JSP+OhfKyLJHXsvC4jMoQgFXdBB0dhl8
NzPnF51qC3a/5ZRDyxF0PaehInjSDy3j68S5CP4oIPqycdp5x6NLaqP3kRBD3nZMWPw9QGYJgbRF
oIAd/9u+8ZHjSEA34sdlrhgr85EISIbdm6sFZB7+YfIUJbCoE1s9DrYsYy3ZGzrgu7Gh4wBoCNia
e4ghvRHImJX9Etp6IDg5PcFqSrav3qh4evmFCV3b5H/OZJU8Ux27WACULQDnJ9LayJjQk19SjIhI
9JAcfiDYcNogT3c7tIiBiQOQtFa+j7+rfE0G3ptL3LIezCQzY9Kb152p0okeMfvWxmokJSp57oi5
NcxRUjfaecpUMp+PtJuvYxkRUmC/ZP96E4JuOSLP8NV19IbU4RmHNjX2WZCLJ8ekxZFINjcTNEgG
T3VQc/xQCpCTH3kN3601BiPsjMj0L45dmbpHfE7PMU6UrsghmokqdC2ttQsbkL88xpWi2O66qXZi
DjfUq+fVDxyfDTRm1ASpVp03Zue2ykal1hFIX/hizw+doX4f4iM0Sqf7WD5RVCfLZ3BUwFhhq8uN
X+zp984NGIKmSF5cK59aiRd6+Vv2RFQ6hDja1WDSuiqP6cUpa9wfiKzZYscvVd0jSBmBlFZVQR47
uRN8khEUthVShtc82pEd55RHB9OBIMAJVDdeDGtXQWIhUa14SQkzy+SZi8B18+r4Pv+qCixwHTYn
ETvaaWNGVnw/yz6pQ2TOMRiZTMpjZRd8O5jEr0tGhloi38h5sLwY/3i6MBvQxygZyFYq9fjSRR/B
+M84sd/w7kseo/b5xxgcYKR1v+aleXhMD4MraLvN0goMR65w+4rXAwFdJtrg3S/NQVr2Y9vGbGsc
2IZhXsBB4/67dFRCPK+EGMfpYXW1QDIHIOYrGpSPXCyBRzaCSrdVo7jkYoQThoN+X6DCLWLWErOQ
aBhEMqnkHGi6aXOr4M9885jrPf4p4HehR4UB/lvYfegm09sEtcVk9EiQRJlbc6WFHU/7Aw+XSd7U
J06iOGUd0SwlCYSNITm4gRy0AWq90FFaTUW58S14905YWSUJID7Uk+IeJirpjTHlPlg/18lSHTNs
U+d0vge+uwShmijwmuF3St3PCtojoVdBbG9HchLJQMla2tIImkoYI4CcndQpxTkDBtSgDmWbnduW
LITK4+GDTfPtU0YLZ0qKCYcLXKzrej+pKiqkbLOsdA1RarfLzqKa9l8lvYGXS4tMf5IRHH8p+3Vy
uzKEQhhOLqeSwlkAYKpTSAefLffzUUb/veeAnAImgSuABvvDdqM3BwkggDJnQQaHe7dy/gkStk5y
HBowQxavXg5yfvbjit55X1z4WK480E559VDKTYtrmBn4FjPthbSv7WbvvQvaeKmgnWTFaz9oZ0tU
JMTXE61Smibkr2aOdIIkIktU8R5UxL2w9MVVM9A6Biy//TyYu7PcXAqP6oHBSB0PuyqY7adB6CyJ
uOfLfxmqbvriikGDv2XUVpHCe2A57MJr0S7PFgb2Y70YBKUPCJDoWrzaCXTWu06iSUL+XO6J4sj3
q9mtegJfoSjj5r5K7eIJ4lJlgjFSLO6FDnwTkuRfC+8L8+mFnrHIO4vERnR6dQoWqlhoLRmeUOFV
U+XMg03W1zhLhNPKgonEzxh9l1ECavjKCKWdUKl7ykLKpjIEOiz4Tos6yXI7ZmdsgsLWMq1+eLPB
CNcdzpUUAZeIryRKC1uPoGThcQ0Q2OSa11qrdZKkuR0OsvuQw+1E5Dp4NDXo46hfEAXQbSMQTfKI
B7RGpOgOmRhQn4eNpN2+IrkIlpxnL15HdxTc4Bs0Txfrf6BSALl33hnyMsI4LLyN9t2lbh5fgPvr
NL5SK5Y0VcwJIy3CVIyHNYp5cji5kR6AJZCu1jUY0OO1nbJQKZnlMTdEQ54UkWN3r0eq88SJ+Fjg
HfgjKnIySDcPqzKgWFdJxn81AKqmYIW/dXUSkRQ6G6B220dMkSh1qabNiwfhHpFs7/v9DELn84d7
I2NhMHlmIahs1QqNPEmNb1TCqAgX3JMcI962QWWxN1VIF7oeLmZwQomEqC7YfFmzEbRD4p2QUipa
URW0hQ/aLU/I5INvv/PKgtZmRFwXxJTojFDou3ElF9rOoSYDqdW3KiVQRbLzfH8n1tqdjnpVI72F
tcONndNDVrIFfFbq521imHpBv3rGIX47NnSWY/vkROd/B3wqZwpNu+h7V2ryWWAxUdPn3pMDZSvc
xQFtSYpRJ9gyazvNASYp8lluf2Ncw+iLcfJWI77EaBOkCb0IvNFFsMKNebQ8H6oElL0ctfojCwgD
JGYy+ZnqGpIBV6Nm5VqAO3u0B3o9dCjAref9CCjErsNLHOeZAe7Th8pHb4lcYgCZbK0HzrMqh4hv
EzJIy71JThE5k1SQDsbf72Z80G65nhRXrZaaT/NfAE0ikaKmhPadto3OV6j1SshfgnhKxcCSD0VV
WmTMpaGhe34BGWQQV0ZuzoQA0EdNytq8BUkiPgB/nEjSXtfh/TS0ArBJ6OXYkSY75h2txYJKzqGG
mgle5QhpEKXU0sipz7MDfMqZjKwHSyF+QIok3FSAsO8Qi/+ma4BTWLLZv7uXXlZxq7G/vpVv1Q3M
CeVvEIAIVF02QEaOovmUSYOn+xr/Kj8HfFD+3ZilyaTgxdF3uEzF860B+pEVtXCS6FIzASPqmWJr
MaET+zyOAyF2qBVqeKmIZp6kxIYAZmnChQm+ZOJIw9V/jQx7DcopsIYTl9bQ3LiSW6VW8jWlXxjU
e/mU0WzpmEYYC5BIr4X5Mkds1KWrkEaaPbn/87OeAPxsFmNMoiw/FpXPNJ0u3Vej56MQJ5y5HEro
14c/4j26k+8IHIdmbwOwrKMmjy8j3olPQNewWreE8X3pXl9h7sh7D0GcWvqbfCyeuSk72815K9qN
+Sqe1iaz2U9nCFdx2ToKNA4o3yvtlhVZq100BzxheCx/PPzavCdtr+gvdwCbOW/hYq9MhhQouZrh
DpQCG5HqrZOsIhotnivegllRvn+nZLll8XkpoO/ohSFlfSSglhZx2Vzf51CjDMc05fPQgQmUYllo
obK//i09sryYJsgokV6Bl1lsVmQ3da9lnxJ36bfGo/3+OXI6BPjqRlE6wGH7lTo9sUDHAELg0p0n
/3g5zuN1WOjFh4qDeAYonEWo0b80UAyvN0ZOLxomjjEF4PVfpGJ8S0sbvmCBnnvE02OBOayiPdY/
4B3gTr82Qgnsv8p008b7UayXXqWRKUIrOMCmfFSwAXGJRy8D80yPL+nWooHUU0P6z3t6PZhN9/yp
JCvkXMDCPTZxvdXQqe7z4vfSARYn6HVIb8BYETLIFR6dOxFJZYtJl9oBNxTywxA1KlFPJlAGN3FK
74qqsH5sSsl7XvA8oQHzCeU/TD/zAcIxwQ145wnyzX+7uR9WdU96MgGHtbAX3ZdFk/4/xc01iqCI
+WzANtUAzr6PZHBFQSowuLH4m4/91FEDAv6nxGoDirBhunTzjqOPYJHzBRfcJMbxk5DzCAwATCaC
25WVf+hoVXlBrww02j5WOQRPMeizUEFy2vV6i420RHHU6VwMtgU0sKb5UgCPPulPmWFNcCPFO4kM
cRaB3u2T6k85ykH/tDQvOwyryKmUp2s4aoaDI4OQAwHOC9VhOtstBMCs7FYK3EepnuF4dWKuj/1B
A1RcCwFWbe1jAqGoYk5lgharNro9gahhZp8Wb0P13qWx8k7FoQaiy90kABGb/pVf9SPlStVnmzkx
NMOIquXT3ztYwYMp42ewRcaIiOJX+g9kqA4Crx7pBaoTbjlEqiYczUI8vvpQWFAi7niASstA4EUa
lLDMy3qarwQbmITJcFkpEdPd5+raD4asq31bXuXK7EL5sXBuEq2FheHwo/rw+/C/QReljHouiAt/
X/OCEx930TW0ngbCFKUa0uE9ntZpTTgA267LvfCahLJ3vUmP5KkioaFzHE/8D9obKl+/eQ/1mdbY
uAVXMygsHZdUKygtTTnd8H/PHA9ygfKiNtOxuVBjNVv2aDAZZ6scMn/PvFjRgm7jbRSItdS3ggMK
zr8BdQpYFHA+TLa7eHZjSTY8PUYS66IY17OLhWt7lBcAstlvBtwmmHZLa51J+PGSaw+nFBepbjwL
z1zSNs0Mh+YNO6dVqAEbD2hQvYSg8MZQ3TnhR++YHHtuPhfgnlFN23Fry4aSvf8roz22K30s8dtj
yD6jOclH5aizxWRzzGhCbTet7y5cySBcCv6N8k7ELh56n5YNU64SOGlZcMZprHiER81rYpnV+3p0
gn6ku2PxYDW2nK7ppz6xhFKE6SNRPx++2+tn3Zuqs5rvR4bkmrwRwF716x/0H8LFnKIrCLghFxen
yomdT+our85jHaY/nxazudc3by7c5miOFCtdzwxVOKljf33UhzYgdBbZ928kLETe8m47dSwSZvQH
NDQl/p3F5I6FA0v1kzHme/neK/dzilaB6XfxaIQCeW11mFbpI5CP80vHiPC9hlOjv3eA8GefWc/E
r+lSaVexDm/dgse/gssYn5KAXcK2qsm9jJBg6UHxDa80Ma1v/+HvvaRysKa61NqAvCzisw/nS9Qe
mDFsBfPd/NpjHXUknQseDdpscVJSkkYCB6a0NxSp0EJ8IwcslTaDHGAL9KOJk7oyUZubDR4kg1T7
rHhR2CQNtq02Se/vC6LIFM9I9kiRRtFQqHKsZiln8dfqXXo9xJzKApYlz2O2OLPqb5T8yxsDDFNN
ubd1oIsPx5RggbMrVIou/ts6FnCo+2+HywUWnRfv+BpGvAV32cBn6uQoQbna+2YWfzyWpRAyM5R7
xf8+chOvlR5xC53TEAgELQdjhRPSh6HIhN6VD5ZK06tptAQNGnHmw55I6bcSCRyvo5joBy+Fzj8f
zMyDelKbvxCNxvnfpKF4zEuJHxTJhSYiB12sRNX7q2jG73UOJMVKM9ktToHKnuDlU+NiaakyP9LD
MCijBMAbG1dAPLY4TR0vdvCgYN+9jDbtISD13jPHoUeFvKszoC06vE5DXyBhejvG8KtUesOVhBXB
AFIdg/6dONpgfdjb1yIVAJcgEHXVy6gFgXqYnQq7YZHReJ4I+4l1XerWxijT/ZQrcX1zw64oes/7
cNUoOMv6tcKLRHrtV7Q2Jo+ZPCReTzykLM/vpLVgPKtdaSeQDETPf2BwSWNJrLQotlYyFZAQJTjS
TI9YuNcX5F+Db3CoFL/5h0F784kNBD9qYRx/5yuUEZo1jU9lNqv8rqGUA3e1adBuNCGwzSLXTBox
6AY8Aj8zs1t+hHn9Nbi8zNG366KlX2bClLbIu7o3mQUammzLL9ebvstBWn0ahV5rcsTgzzgdXC+S
48aUVImS5XvzX1RYze0r0piYUxybXPmO8p495MniOe7jlLshReX5HCB7biJWFCX5T7yerFDXoBtf
nvxr/aWQBcytyOPJEGomnufx3/BjFug/AFNlnwp3uIWWb0p4IG1td7b4J0q1h3Djz+7GICKwv0jJ
PGkVZU2y7o1HqMu13liLYSPZa4ehypURheNVvsDOgJmEpOv5psl3ykxBPPShU4Zxb1mGXOZJXFCz
iTQcFHWg8iYoTLFc4BpYpXoYXzH1ii5KS6/cybvFan+1mYvzGDVA3qTMzhq6mBY7ojMpd7+T0mVn
voCAsGp7x1+mlTdNTCPZYROYANCRYs/84/8Q6NCNk9pcERHzguovZF1POjSHbhhv4F3ErfkyzIjV
qF15OaRs5RkdMMoTpi/z/uo7DI5XiUVkTKhz+3ljfOX5NN2zJ93USaLa4OQmxop9uj2jTu1rvDgd
FaKx0U2BIDMvtAQM9BJoREa9RyAwn+NU8GrlGqO2RV9OLhkaVkGQeae0ohrio+nuQcDk1Jw56ek+
npm2jxq7UmpBj1hb8eZhkPHXZiLtJqRE48SV+LafaylD/Y5H6ysOPw5p9mv0z1cBJcmBG9cqi8T7
tMumaCICjTCZNW7nFDddeeJREDj0/VE4jLwjo66hMQ7o6K3kQ5sJfEzhMUAa1WnxlQnusbO6PNHm
m3FzQ+6lGqJpSnKHjIopTq15JCoXZKqqIXGLPYbKJOXJQ9qeM9w8WakLT2WYT9H+Ay8BMp94QrYY
Fz+Da1jP15dIn0z0IWrmW3pvGGSIj7H0j1fDkP0MjfzO6Uop18Dc3zx2URyZPIRN951WWiKVV319
QZyuqsRgnDfTwbU5B7xKVKmFWKGrtEHqxSMkdJX1HbYkOVJ5RT1XrDNR8xhtAvezUqon7PFLELJw
+B4EtGUg3MR6yVr5U4CHBKbczDn9nV1i7YL4MEj14qVr+2kMZWNuK42cGgOnwcZRAUH/duIqazx1
kguNeAZjecL8fGAWdpq+V/sujm2ak10vtv+B80vi/MFSlECxKh+q3IiabNk8S9AjbcZA5vJVEfFx
LKTuFRgMRErh/zQJwTIO7LfCc6WM+xEe9ImsEMigSMA+CQEKQgU1GDH9T2jiZlHHuc6VZSmu71B3
tdF/+7Era/0BBKfsOzLT1FzUcHcj5RcN+ylFU3PoVuVoBbtfO2UDQz0xrL39DWPnGq1QznsxR+G6
PMeVaCvB/qMoTxhGClLMfI/3BfW89wegNNnmKaxIcUY/WYt6KvEAza9g0ib9sezj89k7M5mPT3d+
6e41bzSfyvYiSYQxnrlOBKeaaja7RmojvJmBGzFohnG+uO0UwLjXJ+lU4iEI6U0dX4McNS+PvoBF
6POfxGSOmBj+d/XfIvhKayggS8DZGczjkgbjMtfmSgk8b51MzAduMa87mjRjXpbY1QgN4ik4RhQV
j9G6bbQokKayQw6tNYgY2Tb74hf1WhtVT05fanAgJGz3d66ChTLfLa0evUi791gA7qJlOz1Mc2+X
b/Z5Vpe+tX26dXZsEQjx884DnG7K/1Mywapl6qVmUmliWszMwMR2CZfhy7P7zz389X3l/sdoPx5b
UkU48BqyPMosd7cLZdEFhJP1Y1JfGH/Q27v4MV2ZPBrl9AW1kHssl87POWVoCQmRULPZmpRFIUG1
d4Q25bC8+dkguTEtLQFsgc/Lv2q/B7XZDs7I69/WkjOyulfYmRGvJt195h5yacWlQTTav+Mes/iF
48ftvxO1AXDNaObILBTTQjv+e1XJcei1TT0xMO2e56pRLAUJbLitaurEQyaBGYwUaoIlFBPcUwu1
M1WM30sGqc4Qh8fajXdLWN2IcvmUkeAV92W+q22cvfpBjqWFzEAUawPuzJ4qV3K7ipxQqfHHkX+u
Uovl/JF3wMC5IJBGPh/MBkMMNFE3+b5+mCfXlCj1f0TSjnKBTLk4+bNSkNP1s1NGj3+2yHYiOjJ1
AfzMrivuXsX9lotnoUceaEEUyqUZ7+MjbHbFmJ2OFXwybYL3FB0WE1tdwKEdCsoCe2fEZbgxzAUf
5BKrwtL6XOGwq/3kSOWwfUHB9dydr5yLLTc94jrxFiyFFVFBIq00JeXD1MAl1ZhveI3dB4RlAzPR
EPeK7c5RTsTBpRVc/MV4HUL6XmOZzv1BTsEPAStqOkJW2ljU/JzEQ+ia7i27cy95I1jgvkpExgK7
O0Kgwf+Xkw32d2zih69oYzuDR6s9E9WFZEjmNJgt8pqnHbiAYAVNtA8OUHW0TqIMqYwM3PfDNt4n
OadWGNzQGMr3LxKwdW38sdOued0DY8ZU1wSX8p5YGmmYLBt18BIBzLTAbmVSabG+RkBCQiwy+Vbx
8sHzYMkWgzyRcaSp0a07oNDUQFEbEYZ2exN1Dd0QSRmZn9WpQo4SHPhhzlHUpgu/KQRVGxszifyr
zEypw0HAYIJq7yiefN3lw+qwVoEV17P/Aw+eqV+gYagyaLhukDiVo5ZG1bJanzVysdbrHntVgyy8
kdGDhL6aI0mgpCh08015zpI2Ur3+JtAyuKPc2fLWuVqxuwOmm552SUWDmNzjSb9q18N8ODSXvRJw
cEC3wWN5TA8lLZx6iySTNkjoXkAweCCCUSkMtBiRcHXDjY1oL8ORQhQCxYc3Mt45b8jne8eSWBdk
jlx4xWQKM95rXTGMAKUF38NpJ4PQHJMtZFdUQLmBUaw1OyU32cKXsufw7PXUEJtFmTZklLC96Y2f
bY2634sLnJKsgXo0z0vhDZM2TQWQvDvygU4xS6WhVQYe9lwIycWvsfJgBIV+Jlbj64U5g1xXggRk
H20GGa5D8eMEIDw3uSDrtJL7NtFlVvMYuPeA+Sl8ptO9esnB8Pw3/hE/6KTC59lw/lBK5QLpnx2H
G2cGYiZBWXGZZjEYM79y/z3wikTyNsKMGGC3Hw0KriC5WXUGPq/sYp6KQwQadVjJUeLD/RXd3Kwc
LVTKOvLoZ6+w4bSAF+X7f/RLRQuXOc83wtR1X2G94oZ1E6waGDO5OwRpKnIjH47BXQoHCMLHGSk2
jmCMCc6sipXUAA5EUG+V30rj9r3B7/0q/G7jD1G2iwVrci5xRPrmS6L4ElYqRDqxhoqbLT9iSYG0
XzUP7ofOi8kLMgjYS5aTY55JZaEk52PnPiUk2fnt0i0qt4zILU6n52D/rhzZepmx6RDOlotnhWZd
rXc8MBahDoRBpAQgOB00KgVPOnjJ0eNiykyx9DYjFvG3hLZSm+27vhlTxC++Cg89VEq6dn29k/iB
yVxUV0IR5I76rTfOJQCkC8LJSPhPQafp7XMRDPVGtwdSEcOzDv02l2L3Eqak0DMoSC+uLvNLUmvb
6kp3cgwGp1li56P1NPkypBuGu6ZuX1AnKzZNk55KYvBCFKCvmPJDcxiqqnK2Vr6XjPyr+sIWXBH0
aqD5b24HNGtMomQnnwaZmNjKh5xg4sAdo5MkM5tSwHLHEmvs18pvKhvgRo2WHDZ7b3X0ZbUyAUhL
N9csUztF/woKCt7jz+Yi+qdHHbupQnaftB6csEQbECEKTyD8WQw2ECIKxBXCERcqBqWO2ruZSgGw
XrxL8L1LJq3xtkSV3FeBxFjLHqDkw51zwKNBAFx421mV/O+Xq8HLDC7onO757qXzBQT9mvjUOOYy
ByBWNURXic90/ad8dOoBSxbfQ38Xuy7vNuvSZnTT/IDcdoIle8CcldHlcX+zKF9S9NIXgTKsFNdA
RWdyGpi1POv5/TDRbiubT0nnPFawO7hQ8FvE0zYKEC0ni6LDVR2DEutpBRej60jFOxUBL9qk3Y5c
THjX5hM9/vK6XpvO/vSPd8g/Ha1OYPj0s908gfeWr1CzwhXwLDQpOdhOSbJmk5BRhavGWbNDqrIO
RrWOH+GqIR2/odN4FkV789bBeuj/HD5L5+J6kFaq1zpNC1xvuAfgJtF5M0qX3BKSTXSxVvHE+ZYj
9TtHQraqtJPedMs20r97W9SoS4E3vllCA8axxi4aSEbSQbZF9ZsyO8R2OZ5erdtdOSssa0evjhl9
pJ3gumA1AQiRxbU6gJJql+20Yacugtr56Og3yQy8/UPDb/IUic9iQkz6t2nNl2IeQWtUxXASs60h
sBOkC+AGAgP+NczMnMbaMm8nOKPB52f3O7jzsLQGoG8hp3kkuPR+sTwJj7aAlMnwzJkcJeZmgTOG
8DckaHqMXEKuZhQ/v7jLNQlDz6/n+6yy6gMRUUjcaEx33H0Qbt7msdyDbTMi5ydSFKH6DDiPvasb
eLC7l26o48iRVlnaeHgzpZBFY7YAX6YBFTyspD5Nka4+YtSKNXISxUlj4w0ohW4UKUbXZgrBy0Ck
ugtzVdSsaXfQaIrx2SyZivZHBIU4EZsOCeXdhw5M/PlzKgP4PodoaOcpe68fLe1Ug7EVf2aqIGlc
wtcxi2IMlA2NSsk2vs5gWtmbqJAvMAvOOYlfb7CCdFCn2f5nsDmbPzlrLXzXAd0CXAt1sC9kU+cX
x84DMuBpbBrXUusZrrw/6ToTibYWjI1SaYYZLwngi+Y7XFPfSkOyMHQEs7L2pt5KrRmj+xzyD9CD
cqwdohMLuiN4b2Rwnfg5v08rHzbZfbLpu8MfiumHOCAC3qY0vQvgu9zHbFX/jpFlBYEWxGtsJlTf
HiCfX4Qa3joq3RtdCd/p39tDv8KqO5pLvkcfa3CjVTJvThWgYq0EiATzkLQjeQ1iqPTRyCH0oUbF
HB8u3nVnRZ+CCwzIBzAtGWdNoJptbMnqf0fXRzjA1givt4G5FrDmS+U1Nc1I8bIy6FnWXyfIMoYh
OpzUbbRUKApiKKkXZ/fMP6JwQn4SIEmEX08L7btP4v/4ttR855ZEJyJPl3kCFc+jwoRqu3ZsQp5x
2PAu65Md6cd3NUOaW8fOz5SKkTHgCCJFtba4qGjg1NqA4U0sXNwxe4MtoHUL77Kr4PIqp8OoNXvX
jY1s0I/Ds1O+emenb9yv2gH96dGTy+7Y9BO2t85wZsFDWB6UCEhnnfgw51KRfgjobMwB/vlGfza1
R1iXOhKYu98h5ss6nlJSdxLvcXCjM/stcV/c1NModhkThTuHxt0Jip+45v24JQm4UqZzfuc9VG1w
vS0+IauuwaOnh5uLipXs8WnI3QD37LIIjVx3rfjRMp3g9nsM5sAmO1mhMst0JggyIGh3I9xAeXFL
2O653RSt3JSnUEv2HLZonYFDEJD3OKe1XGxYS9BNfDkMqd40AebFVPt+6XECLGHQVZvpsJzpzUm9
5Vwegan28s+iAydMzwLHKiOQMog90A1c4qwW9KiNNUEF8Rjgu3v+v/4qQni4TtZz8fXSZvFwjWF/
iThG1csbjCanN0d2WHIqoe7wiLTErRvGDNAjivgeSM2r/fwciuya9BW/HP/uVS8+91tJq9JH6aQN
+ih/RW1Q+Es5XjjH6KzrvQzk1oZA2TOJ3ijeV9nn+rDlFWTd9VpiTweF1ERsnbS0YDqxW8DWWzn1
nHdFeltHhsHfu0helgeKYAadGAToO8v6ZUzgOlglKfMiHHyH4xc5Yr/nb/6yfFg9nsVoi22qCqcp
gjr+irjHOnsCoUqkprBP9gMm56L+4Ub3wM/QWxG/QxJsA7PkxNXA/J21jAQf3JX8oUWF6mC5uwae
QxPESmJrLEoqUIain0CwV2AbNne7gVLcaqgUvJMSWhAuh6PoWd3FiXffukpv2XJPkueovjxaCgTg
FG7FODYgoDjQCMC49xg8TeQfFnqAbbE+7ZoBkDyzLqIcM6Hqh2lPyb6oqIHbOcsbXR4wLUq5z1XP
w3sEca6+NSJ9YpmG8oasblwWa2rdoxCFZp02gmwHEBmDRhjYO+XVL1jiYQ6J5DmPGZftnH8jnFO7
LxswbhLYsOQeAi7+Q+Rv1XmTNE/R3dZXM/lXqNIhoB2ODFA9ihBc5/y5joBQAtYl10BCQCLv4+f9
2IdJ3oZ6WQooOC4/mAmR25S29iXqw/J3msdtnA9uCNx/Auza7VbaF9pIOcJVJqs3zUILmG1i57JL
ocyNPOD4xLvTvY8nI1sGWSwA9BKKLBv/0TpdzK0yUQ88K9krjH8xqAbQ0Z6GmWE+dQSIMXa+Bp2J
AfEqWAb4Xec1rfUiqTIggKhv1yFfo1B8+gwxOVF0HizwjbkCk80rI9B2Pm8uyNBenCVrGWWvhsQH
sNptHB6E4Og/4orRJ9tVFb3l8id7vsIXNMXC1kvT/DN58g/oMS1Fyr//JFzqDoHhSYvdp+AVDlH5
qyAPJVZ9Mebg3DfXZ9lH8uSJpz2CB9vjo88Fq1B52eO4sL60Abj2ACcz1e205+cB8W706PrxM8CL
Q9ZEv7famuo7i9ZQv/tu1QTBUr7DidzIfP8248vNP4GR3faG5WfaJwnGhdhLUCRmcD47wplVWWPe
wFa5oVfkroyXwTTpXT/KUWlojpEDY3MKbiaug1CcW2ehgRljCfj9poEIM5FpJQcRzJj0y0PT8/dT
FO4jJ1MTd3rcVTHCcNzqEt/PkCtqTvtvNpZAi8gkgwkqKyOugpho8KYip0MZtHjGz2Mp4ngEg03Q
ld6mo0LaH2JlM6uwNMtdpS3zcm6AUQ/vE21ShSapVAvq00wq8C3WpUhO7Ql9aXdgno1QLJN/fIgI
VNPKMwloEWbis+uTgDcJEUJYew2Pa3QMc/waXseX6wJUbgQifz4mSLHg41NHJpUJSVKHHgrSNvuH
UEF9fMEA76AKlMsNIgRolp4lr0fBakueejatisJcjH/UEGRyXpFnGYGGjXsDAdoTd+zTxDpxtfyH
XTZ/5Bk2vsqohbm4qR6EO6V39iQDBwmoSsT/GP3J7hg2GfwKZxYrNxYYQZCX0ydJaU6m+KHH1uMW
8EDjvaWop4yZNVU4qhKLPaTsewePSELXPk0KLGRVwCSJ5YoJIty80f0De5+VTxHQbz4vjADcMPMB
49QDH44w2PW5chcm7f/qcaNpTMWrPaOsFcndIydZIEsJdCz9KJG3VxOH0zRKn05LUD1n2s4tbI7I
6fXwFF+2HDnc3T/ift6uON0lmLKG7HAcHe8fE/l/5zgdvgNdmYL5T8c0dm7eYT0TjCFu6t6ke1o0
jT/VKPJ42913o/tA7wrEHo3jnJLJbz4b216lW48IzpApJ/myFK3tCkwHg919A0dI4sWJ1nqG5mUp
1jbrhE8Zl8FeVjUfYMPolCUhk9h7bGz87/DQf0HwZouctWJHZ7zQlQcb39IO25kX3oLJOpfcj1AV
KhTaWNUB5a1K88tLLZ/d1vZRQgVgnuezv/QMrpT7ZjtGtr9ShancVNSU0j9UhGlapMvCEZHlJJUq
rpt4UW7zu9pkIdMVuafY1bt/HWVG0D/2oKj5Te/ifp9U3FLtF872fI1Ie9etJ2f/6VNIQMDts+B6
KYtLkdVtBVwW2/cxW/DD8uSspKR8tZSNo2EiABlK4JJTdrIG3JTf0jdk0CpqsSU1HckM7GSMffOF
OBE51XFss3oNZuQZBcbcnIBo9AfS+vE5ppR5yVZpcjVVq86p2FVwqmgw3xxcKOWPrYpEKHsSBKw0
ZxoCLlfnt2pbnDxogcqgHQv2/LKt0qxZvfQo1waEm+63M7awGUvaDE8FR3l2c1fffiGuuaW3VtHO
c6HEhopDDzt1CiziFXu5xaWSSOcKiyKHul7b0GI27GjtBgDRWmtAm+JeeJYpSYVAz81kRXhU9m6M
p3oQmffk702NR/IXasPAKWiX7Did2uwcezupLr0ZKUisLkp8ed4I9czXZhEL/T+IxJdnc9es232M
Yt8tKMy96dggRYe2eELuxcGiVFARdZXXgXMavCt/B1Cyi9GrqgEmj9kwFCmTdsvjZw5YaarNZVOW
zBAEi5KuvkLmRE5imMQmIyaMfAGhqFBzFjyyGheTK30iOSHgpGAw7gRvjn8ZpWY3vpdBYuzco13J
o/nJRvBu6C63EuRiTEVELx1gjhxNBcRnZH2m5OEwq3pSyBEBNWFcXTVkIQOrVjsXqdHy0cJIYf4Q
Hl3223jWZwWYglt/E1U3nCAHeDIxQUMLDlQygWRzf3bVwA//JUU3hb+s/a+kzQdWhtdVKtzP1Vpp
cBQZspFKu8PV1y+oycclm7pxlGlL58WHniPVbFiij+bk0d7w7C2ZGOa6dybA0DkZKLUL90Xp9qZ1
CQ1CFUtJx2eTq04GV5KgWjfycWiK6MwCXM3mD0VpnvMCicwxNBxOPxGM5YKz04kEWqF9yZe7J87F
s/WQ+G/WFKxolWE6woWcYqHNzpahYuZ2DJ9ryriJqNXcftUPPXwPQ71cMwP076GIvVlGNW3GnMwu
mHoqUNNuk5QhO3C1uOtAQAtbIjpWJrbXt1QjtJJFaOWe5Ct8QUkOpb8efd7z88pKeuyraaSF3W4B
CBFpEGIp5RAK8zdprlhYfn8YrVhLo/saJLwn0ly5SzeJMyOtadqV4sGG9MOLx1u8HqNGHwbywhl8
v/+93YLxlX/52CvG/2Vpyo6e3csVzdcStzJrYZHiiRVASF7rU4Q2xlizc5W7INMTvIEHjJfKtucD
D1twu9Qu2tuymlFJ8AIVez98z3rXPrr78REf4ChY2iQSojPmVWtbqHonxbktU6UnGgi7/WhUHCVe
fVhJIX34++QkEtJ+PKvLZDn2vWHXNpWzQbhtbedY1rG0g7Z6ggp0aSR/SohB2PRzLsgV5TDksTWa
cda4oweOt4vpUOFryYvf9ZLNYW3RH/HE+yt5q1HfqTWiMXeqETO/baBFXgTqiwaY8aQ31906Fwbx
ONbbtT9nMmtifCno4O2tsGnveR/kxIcUV0o0B0BTgSkDb/aLrb80WoKpJ5JpE6A6IjRZ5kon9Upl
Unvuxpaj5NSX3NNNc6pTEuXV2H+yMzCdHSJGMunWNCMN3qIgpfi7eptgfrLgPAIjszg7uTXVV7nq
Vc2o7xra01zpbPnOIZwiVOXY2Ie+Ak59/0vHUPqkRRJ9lyvGNeMqAzx+HwJDmVU8lMv2NBAR4Eps
DJaj7Ya6M9M2PsSu3WJrbACxZHFySSwyFsClQY1/p5xSTNyEcYVG26n9KFqPBLfLaktO5cLh4LGR
WM6cUJXCngd+vE/OykOPaMvtYdJIA8RBotyAmK1QMclOq0m2r51yPVwlzU4p25mPfEI2uVqjY7dW
IjoonhDIAt/EEUfbAhfMyNMvqG/HWTnZRRgPSvK2kQE1PfymmnZtoyi4vWOZHCgRISC8BNkWBi2d
8zJSgKI6Om8Vm3DRuZr8CDUPbIt1/efwTBda5yokgaVM+i9cXQlLh+ocn2QEuYO5gPxE4WKQLocr
5rQAOaqEYrctKJI6ZMnt5vc/3Ey1f7mkdn+gmBjH7cpYga17Fyv8MgBM/XNUAkr5rV+pq+Pd6uds
hSjIxUqofEztQwef7AJeFmwtpO+sS1iV2kR6/dhATWjRM3gsaJ8mzx+dKP+/6SkMA9gCpHHJHETY
ipkcHHgc9alryiJJmrzKkEhIy4pXMw5DFfI/eTB/0l+BKtX/vsyf2WHI+jipdLa4qdO66HQ91601
vnv1mj50t8kIUNs0f3BTYatN0Xd6vBl+bU9TsJZWX4HgOmCeBGRP/syuoVoODam6cAEtbkUi+5MY
uGqQ3b68NStNZvvnbc28T3ImXsvyAatX6gEvOWkeW7pCPD4vBVqrWbhkG+sM9ekRA93+5qdnrgRN
D0K/iYD4XT/l1cW5I6D6Qfwng3NsGbNUk+aXVFf/egZ4tbZT8JpHxdJjdpVq5w2GvBNDEPJbx4XR
wfboNzjLsVKyZ2YjkL9JV7dUHIyZ7cTIozgRC/4qkrvWM4tLrdcCvEnlDPuxTK62f4GczNT5+lh8
t8TkkuufpRZpaSfl4wZ3rtk2Gsl0gQ+KjTmGe4QicHmjBn4krZ0Hb5crgUYDXRMGV4RoxzJ+D1Qr
HWH+nKXwc/vVc959UtAMEbZaS0ushMLX8cxTDLmKithZoTXKMDG/nyiV8d1Hc3DzhLr1Ur4exWGp
NhTQAi1pfnhcMAzMVsAXd+mdLUIqQamaceosFLnVLrn0ybpsLZWPmDYJ93jIjrMC4q+VChwkbYvA
SDaHM3iuXOGwwJvY87mUmRRnj6wZ7fDN1ZFFrkD1MmVpa1kZ4NGIhwNzkhs8mBiG93j6u7+87Vax
2EqGtCEzvmvp+MMItd0V2vgsdTxJB0wH5x3KHKkVBRcTuxOI4honpZJqWi6RRcBlcVLyKkVVv3fM
KmjUuepAWK8VcLilUXN74uWwYNznaDckO3Hs0ik5pn1rgQafrq/RfLHLL9u2aFMCP17iPd74tTtn
4N7yjTHS0C8g019Vqx2iwk8n4JpMJ8VKgVCMT+h/3BDwh03ZTynmAcqMrUCVYt1OY9CIfI0pLouX
nWyVxNkeZ/23+9/8BBreQs8nvRNMHk0i4EjLj1v6yApIUlxq7OfqT8LdotlrHW/w0srIxvJ0BDk+
afqV945VubwBOpGlFYoBjAk5wa+ObDf4MLk076maCwRM4yUSGoqrkxb/zki1AnnG7+GQJ7DoB6wt
touA44WUxmfa33zvrBn+/i0ny68QuoAw2gLUHAScMyCjSWOvggN74Zn5ckaaZI+jZR0FjWn2137F
K1eLawZD95jPcpv5BrjKtObv1Z6bMBQP3R7a83BVQKwPJJvc5qvFdHN9NaAgWFaEerL3RzUzAEnE
aQ+28onIELOL7hllGmI7btU2sh8RGAHDkZsMYRXNSd+4Ehd56IfgCjZHlRgrm03t5O5AOD95qhtC
tajIgDEvYJ9yOgV12okn6nFNckBXmKg8rIalcxYwWgcgsE4zbZS9wZxnYclykSq2L2YKGWKQ0Eoz
57ftRcd0sMHUlBAHY5sdND2hYTJAsqfquXZfnuDGAzPM6f3EgvxH8TIH0rdP+/CjlkA4BjKorOc2
063YwyCpiRuGzhi1nuBXZcWk6VFnZ/PuIgWMF8+yUz9gL7xCf1SzEc0pg34k5M0DEtTgGIlszxCz
WrB9HKKLbUwHv6tSTDc/Zz6thesP1EaV6Ffjk7EOZ6rnL5+xnI65AoEebUToiZYUWWnROmAza2hl
Pnwmg89uUMpj0iii1VbYNh5pCyHfOEDsC9ETjjfkYhykncktvzjk3paHnH95rCdssBiarho1teLx
7RrjeWlkbMXh2CoQNz/79dmPds2sCMCOOHDOn/6UG1QVqFyGgVV27o3ZuYsQh8Rinu5Ag3PdTg3h
pjrSDtLzUm9fj3uQgre9swI07kAaTylH0zgRHljaBSQofq8JGlZzqrr9RTycK5t+f69MjF27p5Bt
5jQQH+O3ydF/RXSfwyyYjBLEvjYIutNAwul0mayjmesHHDYRrCmgKF+tfJkxVboogG7NGfycJIZE
8VqIzIJBCSoaQayBfLjYgb3QghfW64WRYzf7N4+fOW2AozZ+ABUm65W/lzsXBXREhPyw8bfMw9GE
SM/SFcMqF/9ET52dWgnBvFNcEL9zLdAb1Xd3+n9U1wwagTe2Q5P3FJa3ZnsOOiN7YUuCFG+39Lgm
K/YufN31k++24xhyNxnKsvipH8bPSKSvKQIPJtMx377GN5jf24gforBQhV6ra65BPh5nZhMiWuSQ
tsJIbFqDfmZhLhm/cqm49KWnDOofw0z1j3Tpz5wXb+EaFhSZ8D+HjvIUyVy91UngishO26IOE1u7
6bGXWkWUHsqITcYTGuxnbpYC5JDxWCXn919KMBCKJJgi3fFmoKoR+T7P9Tkp5tMAa9kscml+wy2Y
b+l8Dg5Hi9QCZ1EC3ov8mNS+DP+zy14kx3UTOpj08UqKbPXyIEsMto7hmOhCdLZ/XsEmS5DLcsE6
PJx0Em1lTDIo/W0ZywvY5aOf1eLMmpTePwhlqC8aATA8PR3BrQDN+QOFLZGedDqZJRa2oH/DkM9V
YRN98i8aWwAlpH4IpA16jM+EjNTeq4Nc2e0KclryVe1axQnDjeRUxPYBuekiHVXlBafXTbQ4Kp22
DJXbKsZIEzPMI/i5WJk/WjWVtQR7PiyY8SU8BWHjfNwymhwt7ZSJMSBmr3syH7ECpHWp7FiIBujV
ENAD08y3BVHhTDpGTgjJuzwuvI5VZ1zLoJrW7Dug4EURAQZ2Ovzm8lbdv+sqeNcD+bfNK8LWYIGq
76eU3O9oGfwyWJ0OGnOJ+aH6ZiZuRoMCBGb4KcSWHNzxeVCZAI+RGqHoJ57pEV6Tw4v09BNcnGlY
pUhwE+GmobPbKDeqTR3oJHSKivLz3zH3B+gSZS032lOhuSvVZx3DL/PZbFD9+c6qhVMCD+zFBH3N
BCRCO5jAIwVORlU5MqNqOO2Lsa4vNY4LhunTBycUOuXEeQsa2BK+XewC0uSGovUbBrNlG8PqBimx
DQ81loIpcopXG8t8nHkAI6tkSUZlt0jOp2WHTuL04SSWsua9DJzr7nbX3huTQIk1wC5xIhGiKdPC
ANW0Uk8rRTZdMMAcMQW4FdBjYWtkE5XMwaOUGtRRiRmC/lnapBSgpPc3lhulXOKQ9rmUIL2yKDMN
QEvPSWqaA5X7DX4s8MhjPdFTSEvjYr9bhHbOAZlyXTnMRd9XlsMaZ/3ZSuVKRbss0q6RX7ikghB6
B+majOnyhmjxBCQ+i7vpslUQgpZ1XLEt7ru/UcWxUhx8nMnWSlPxP08iWRiTkpUZjMDYzzwNNLfa
waZSGvKajTZJCq66cAZJ8m96dIQziWhUJpjD3/F70eZP5rpsHgPu8/3RvGlTMU5bZguYuEaG/BgU
g9/IynGNjzI/58obBgqR9oJR04fmBiBFwZADKKCCSFTs8wBU+UsQkzFjBm0ZKyEtjPeIXuljBwub
fgyFmd5nTTVKkUl8tUIZjhxDO82f+igh7VacLlbKDDNLMahFtKYc08VPIALGez1pKsmQRzoMcBMh
nxA/LnqDVIbSwqFXMREIicZlkftUhZ0f8yhf/caI+BoC2Io/4w0wJIeQ+LT9Gv+p6tBwrBPEvy1R
VooMrxiRydAvLBXPGINOASaz9wa3S7vn48p2kY821VrvbW9qxYsaa6bWD6+BO6Wv6saXx7gDQ8Jn
6Zjvi6hTtYRTzdkxjWDpcSSOkt3Pv1DotqAWxRy4oqup5G283Z4ta4p0ksK1BW4W0OiUSyrFisDU
JkCzbwjqArZlw2/SVvxnUBzYukH5BXZcXGxsRnxtEa72pIYwxT7SgZyml3TfP7E1NUxyllMUrsVH
Lym+QogMeIt/T/UcEri+jZpJb0olZwdv56PxxQq4LDJsCFmrm5WXAJQ9Q1lQx9ZLm7aOeFihawhN
HY1ZamRTrStJwe5rMaW9zXuNFL7UpTd6gw1vIi3Iw65weVukECEqojeC7bKbgLikIUqyc7MXERGa
nh+hUoZKMxDqT4KFEWrhchp7/RaOnGnigM1fnQOqQIRypzt2ztXszIm8YS2fAmaeA72P6iyK542I
hvSTgNEM8TvNdGRbNIja6Ozl80qRfEHo4dR228uhEvq6enVpGqjgt84Rb4nFkXzr7DQKM6dPJWJ2
JrRWFcqmyHuN8okGashXYg94eGxOXK5CG3seEvEi8pZ6IifK+PGAY6ss0GfBzCnulf6F96EjpukG
+thi7dmC4xSoUs9GAk1QhIlhLhYbJu07LQoNPLNxHs9c/uikpwE0WS7JwAkaNhnzMXQKI7Y6seKQ
4UmFUOkYtop+bUYCtqSa9PXEbg3CM1KTtaYaLEcZIYLXLvEL4yDPhsKZpIrgziLXQoZTDETABvfN
drzOy1rKvD/OyQkiQYSjtr/MFbwFOet82HMMyu/uldW5Vn0GxPaFqxfV1ShOn93B/Tl4N6vW3OUu
8sA74qLb9/F4MArZF7dMZ5LsxSJsXdp2eswk/T9HYoY6Ll5IBO1VLtYWbn05OIurL9iYi63cDimt
XccxVdcbHoWNkwDfybkk7Z5BfMKgri3ZQGyhG0tJOKoqZCoDescYiBCCOcHX4fWW6ICLgjJSBJ57
wgnsuPxwuNkkdgcYbdi52op+Hthsm3kJJMqgSynoMS2kvaDkBeiSGYOivzt5b+Od2xEu9NkpQb1k
tdvgfW0u3TkF47qj0tNrj/EYmJ8+SNsEn8Ss0gUqOoaSgdsEQ/RzAsyZ3Y6oYESh/sNHbReAmgGq
mvJ4W1jf9M0/fCVLqST1gqR1MOR0T2CgqwxI+vuOjWysQCdbddm77OqsAsD2bx3DWKKyNyaGkwX/
9d9sh68vsbIcbBWUJrSxITCTFddZ6l9+REBCBwDz6/ueU7/WzdsvWUispREbb0hBwmrvwmTAIH9j
35fD+AkdYGG9HW58vgHEQDNOH4dWnjLFPMQWtG9+aIRdiaFyIrC3edU5jDQYleZhvWmYAEcVjcoG
BbyzpLQVtbSGhmoC9NmQSXG6OGMbeOS8zxwfpiCIMyoH7thUlCrtw5EX5TGWGiiZL6pyeRJ1XQZw
7pcnfD98KA0bs5xEjp0fZxt+DEZWB+RCsW/cGvwnmGev38cRVVJwM7taKIhuAnH6yQEFZDBXA1k6
cFF8u7k16doOyb9VsUxy2s/Dk4NT/q6DpzO1LplKzx6x4Q4ivnV+uzAkONDUst2+Ho8Veb+PxsI1
pINLXBV2ad7ZT6+B/tHpJTN5x1fTytlrqLByy2uyigVfdFPd3hzPBn6kRurNXTxC1PyIzct3LjwL
F8dWWkgUriROtPRbUgNnhWX0nM8NU6a9kvVAprQhRNYG8EQkTSC+XH0mAxHWEyWuv+MTWsf00Rh8
0/DNZz9xQRsq0x96jaouYn+VUuV9MOTZXSJbnZpSyJDK1D88or/hrYSSJr/pknJbIvSMUnC7gnTw
vbBpf3gVokP4fe1ZZzNqFtznufBw8yZTyDg//dNT2RJz/8TcMqBHml6LamM9I3tfHd5FsVSe6YjC
oOxi4YOa3Xvvndy2CKzMgJCJIhWsga1SFJusHcS5UwQyCfS7J0WDJVj7NFL/ATQDPkQX0G5wGC5K
9dOFlSKbefIGfXdCgAsx15lSzVP//VUH/zo8UFj6CEpGVxBBD6YCgnnelFJUW5iJGun+9CHqyqSv
OJL4KQfhIUiVW+ThOFWdGZue8qZZcEL4zRbL8CYBa448pieQWmf6RX2l3e3DDkqQMsvCuAavrK5o
dVeZqZUnHwja4y/GmucWwrwxdTYxj8UFXRjstB5Hvaf244cvFNeP70LmkCV1p3jBwcun176HauvS
JpVBhnnJPxEU/7nEkon/F8VK+zX+QnwyfJSScaFQTz6JSMlW0+zq70sK5Wwb/gJJqQvQx4TL3VPf
5dMcxKuHwHzAXNfw1VBRCFT6I5ohiTQ2fH4jCpAgZCOL2xx2KkR7tF/oFIyfna8uBRukoy8tKUi/
b7ZUVOA4ZDjcYir22HTJkTBmkipqHMCfW4b20zlHhgvpP+rTIqkZqfyVFMoKyTgS1ZuzIuWBo/Lz
Jev4gWdG+Kx7BVn4verHKCR+dTjantdyjQyTybmjjmOb9RCNn4ZgxM244ndUeevYd9DJsBnPBp1h
/2r/6NrhRXv62Iqo4avSxd4qOqIeCzw4nI/flBRrFk90/juY0L0sp4s3uG7N7XENcaiBXykdakBc
uyBuN2wrN6waFRxaPl/fbhPQmgyjG6cg6U6dU29qfwGD+WbQa+R0cg3+/Eb1sQEeSu7claKpB2mF
pLTJ8ZVlYtw9t1MZwYUTHAirJEQAYMRo1jOenyVyT8dHLKvmn7GTdnCrfG2GsugYfD4MSgCiuncX
7cdSXequSJtIb4U7SLZRd9VdavfXnuXLTK6t/Q3ERmmZA8iYwkNU2JewTk1DbiZCfx5UcFfF3lpg
0PvKmn7xnPeUpIixLGn5U6gjrunEKTVhTI7Ks/w+KhVVEwrgsIAJL0NFAG1Kf90CETWKmVn6lQWI
gS8s/J1O7mrcdWPnLB9K1qqphdMhqIVmVYSroRgiztxwy30wg+pJDvWjtqqWXtZ3li8fpU7VrdRf
y0zp3VH3mnk/uFhkQafN6AlqAa0gz/U4YbF7uY6qHfE/IEnyaoGovoJQVJnvDSUn8aGo79RrVSv5
IP4fHqjpkPPYt65fiUbvUyAarmd8qr7fPcrOQU1y7PgmC8CtkrFzac0cXyOgk35WY25/AeBuaoOu
TvYUhkBp9NLMrivuh6eFkdjnJ/VwGl5sDRwUKY9+hossTuIdDTU4dyEEy9ytdVQHDuOFHdu2HmBj
A/xBLhYzLjuiAeWAm2slbBJcbskFP90uJYuFeWJhc5xLTlNLthYzvW5erIGztGM9ntc7VILX9FFm
xVRSE+bnw5d2U0zy/gyQXgPry7amU1h99swyldiIEdoGaUoTf1BrqDLcx7aFmhJJ3yFbfllfehuR
w//u0jBEBI+y58a9xjKZNJHPClUVnBLhz1ISdNx7+nrHOyNTC4KaSdcxdkVXPvDVLgk+QyWoa1Tu
d3py0UkzkVnfQiyZazCeTSGMi7l78dHWNb9goRHG4q9mdULqr/0Nh9nTPtU6eYjBfznhAGu6jKPW
08pXzvvPintC0mTJ8PE3vKp6FhsJbwyrCX4BHil16R6l+QgWa22odOhvHVTojVVVnCigRibvN2aB
P2wgUX4P8609dJxV5CdN364j0WeXh7sr5Jrkok1Jljjztyg68Hl5fl1xnMV5T+6SJgmFLyqeB+fD
ETF12X8zfBcVjZHE+wRQWK5frFHkUUmwkQ3SgEZnE4j+elJIGws7itICPGHyGlKjJry9dpYt9IMU
o92UWkVYUU9LARUJHQbOTouTu2xbmC8PlqVKzwRQCQgSQZXB08hHGz9XgMy1LXShAGFIQQ4s70O2
aqTH57GO4/WVh+gOCCS4SLq3RvqHTcvvh6smIRbjAOtSi8WJYxCqGagQrXkH3G1AUc5lJ/UpbSAd
95LWG9RdOG4jMdS6JGQvBCHQGOlBe2tsP3MEaHNI6nGaLmGfxoCqXi4DH5o+9/DOopDTuf22wq8B
+z36abZtrijYEaT24HAJqoFY8Gi77gtQ/29oUv5IBtMWdwMA+vVkQ4ipBN4NNNVtSAcq+cwofbds
oCmJKjGVr7QosaphYD4iiUsSRupaMKAxbLEoTIUI/L38j/mtL70xrU2mHmIEDtqCBehcFMzcIwAf
Ki68Cx8A6uoBpOy8Piat6E/mZrcADIuZBVkHyJV+UjqfqodL1Z+i7kWziwJ7a1kojMjLDr06JbY/
ACvUETbFVciUiAKHnQq089eidtW2Gbra1cKHahSBAhYvNmpuVnc2+xQB9tnNk9C+nwO2dqVBQdee
amZt3eo5cb5jHZcMnBTdmcFZDTfvJnuewyFVI0/tqTkNn7dc6iYa6Ys5jvWPMFMBlO7t7PAGaIqU
xswQwnJvJN7wXFcSGArVTiNW0sqgdCv2+BSw3WaMW7uT+owudrfkXUkEPQoIejSmFKM7P53zfcKO
Ia5C8iJEm1vGbZX0kQ1pL3ADAQsGvHN/YqvaMEUbQKmbzEVWPA6UbQzlJCo/aWAIk661MOXL+5d8
yDa/GSYMur4jPf+XJeT0lbruvqoFqtF7wG3M8yehK5XgkT8pemlw8ofBZwPVOtyxk3PNt3bcKatW
oTXYlekKWCPnKpCI/Wa36YnNexBToDhnnIltvcfxAVTUy+YUWJMEUOzZrr7Iaky+Zfweg+L0Go42
AeE0QJWALlbYZ+OFurweD02glsZpYwd8VcvwvniROiFpnPGXfNB0+uFpJDyWVOCcesaAcjWSYg1J
+PZeumIGeBtnHT9StVVYTSCbYY5X42XqAhWtr8JO0QL8j7ewWnKYANiYky39frmda9ZvJZaqVse9
WaTPssu+yS6sk4TWs6Pl/gWN+Qf07dGZF6FGxv047PGOJRt2QU8r7VhjTlwXW73MGFAP0GgeLukB
omdCC++hJxQu401KjI3cVauknuHduHLKXcOfgyEF9tlGaXWovp8qPsZRo/TPsGny/i74AM5uiU+E
Qh8wl+F2rr6o4pbqg7Ol9ABpNjGXRam5Wuc3HNGhwSFga16hR8UbHtmZb9nujvs088qSMsoM8IUL
MttkQ/iCX3dpRSjhTH60YUDNu1ZqufmrmTnVxZtymOlIppKH0INPeDyPeUt5hluwVvRRwshCbcDN
q9a2HVywopsBbtXGft3NdibvnjEdXVEnsBsVoyFDBrcaLRCVZaphqw/ehhHq9nlwtFWLsfvdLOJj
Wk386kytcWjJ1z7XurXTDHGDwHnszNv9/xzXj1vOgoLbcq/qBIywj6MccgbONsoL6Hti4/AB8/6L
Ir96QQztovC/TTkRRbiT9gyOBabsvsR3KAZ/S48ENHOy/8K8+jI1b+vXOY3KOduew73bsy6f5tuw
wRAvHmAEW/X7ixhZbROR8YZyvlMCKgjPJmXPdiR17YJbsDojkeomEw1AAMAkanGnxEIQgm0SuB1y
yxt1TGRa6fSYm7b+HMh41/RikI+ISW0/nJUtPxTbt6UFM2SFCSWMGQcM2XDjWkCx8mIXUz5EgvRw
QN+tVG/XoFYwSZRDc+zzCRDzIQaFys1l5/klm2ILvInY18qT9anINP7ihZcCtpks7epQJwexpPwd
it+tMUdnfEsfmBdx4/DgfRG2/nrs5SXpRyfd6HOMaJgG+Ku0bnhqjKtGSYYpiPsSEmNOoCF1pzQO
MK7L3AlotFzJfbCZQVA0yEKgNRKUFttqrDcnXTkFEM4iY5bkMvO6wT5us4O/jiynxb/AWryFgKsh
UdxmVQZM4fB/XZB3DqhhvSNGKFAaXvrf51XXWSC3mKQB9dMsf0O8CwlHjSNKfQs8hWlFyhGyJUJG
bGi8xkZINBhqGxHzeA2aZ0yZD0wPzz+ZDsU5TwKY9W040L1ExN+gIIxOL6QhB96BKoZi4wOZi44O
OBZeD7b8pHim8xg+YDdMwD5J04xHgWbeSiPwEmK9KxpvczO5nG9tP771hewgtTNVkuCIJA0/cV1h
khijI2cjCjhcrUaNPL67+GXNKOv51VONCPSXF8BQscNyvsCHZo1zG6PMlzjBQOA+YWazVNPYJ9bs
TUXf1DcnzXmyhp5kd3vM1SyjWHcIUpjYHIpTjLSBo7vH4LHsFdi8p8HXFczfUFuH9g6yQUCs5XWi
Th3JDjJwU+imr7Afe972WCBMz2sp4Zd3Udo+hgivygYKqQcxrcihvkEs3uJ+N0PQ1O/GS2Zk5LJY
pTCZH2QbX54vLSyQFgYe63nxEf27/UJLGzoqWi4uumEtavFqoCzU7aRRpaFzTuy/EpwHPIfPbfMn
kDWZKpyHNF3qKad/Y6/uid9Wz+lqiX3fejPDtyP4G9GPxa10ZspXj+s6MdVPeuFkoxzkFIaHEsJL
1/NV3mnkxHXLnrTTAdcxMkKKsiwoLlejpOWzTwrnXMw+nPmMb9fBSsFUL7o3QCOTlVoyUodDiwXj
N6nS89/DuJHDzF6hXEqRAsF7MFCmrN4QwXxz0V/vxYsjYriAcN2WGWApzSNX50gYeSuUrqYMKQ0E
Y3r96IMfCAnYzl9WYE9uD/OwtBOgHeVXcsh23A01m8VF4PMDtr+411w25l0VTQKbfnat1cl5ekZH
QRad9h9Y2PdzsFv4QAuf4C7CHKquzRtMeFrTR0wWkkb3Cf5fpnzpi35Ge5tOKL/cKWAZ4yTHxVYc
PGrhsE58OFAgUDTZ965+YBfqQJ2iNjKggH6MP8XChqVFncL70aWwokmYbYio9ZVOmJ6g7fFkm0Lt
tN+AdBa7pcWBLeRf3XqIjQgQL9jb9zgaaxIVvlA7YggLAWRXPTeSYeVEaH6Q5bLsybIzPL4ZCPRL
r1ZZkNwCQYXwFC4XSZXK6x+QG26EQu5/ud7pXYg9F6T6wsKx3QV88PeanAtmdJv3NiO0IJhKyKHu
7GAmUzFWvVnfDbDLPEQ5S04Zz96tU5k8a5p3fWs8qEQubBz+pBdBXylEdxpPU5XhL1yjg6jdtNwB
6MClxsVxjUgc6a+mkXHw585t/QtxAHI/BN5Z2JjCuzjy8yL8ixPihLOSWzF84S3owEIoC3CLpQra
CQ/I8PoXVO1oxD9extpumKqEo9vxeawEg4MBEEnp7OMASwxyjiG7PUsjf0p55iwx2hRlt+nKpydh
VIdn3C754eALNPwfO1PLwXTZhSMMXdkdrD4vUW7tSVLuza9xh3YudyDUjhMs6HU1p/Lzlivv7+HH
aljOrkXlTykRVll+vFgeKP5xfscPA4kDDkH8ou9itZ9IWUtaW+jFYHVeWqSgFm5+kuQY/1o39adN
eBlNfUnjLCTHfBwVYC0qjnD24MWVbygQ4Mlu6c+GiHyLLI2Hxiz44r6w4Sq5t97/mwJ1JEIUBTqo
+5oekbqBiSRLIxSVhvhLduRX4pPSX8TwvL7Boe0jxHQfKBPZjkPugEq4kDfQchAHd4cvXzUTJhkb
Cx5NHrPljVtdQ7Re0Cle1I1adH6zkGSBPd9dnJpzhdASUZ/n0z0CL/N4tHPx9HwYd/1gJKk6NqhI
JQ2civC23Bm4C/wj36t7LZnReuxDU8/KFAd2UMCIU7o7rB2MUent732lO/lj8f5587ZHkRir1Uqt
YXgifF7ll3OXwie24DLQfNnnjDpmZoSXzwl2FBZMYskW5Re8hXZgToW6Xo5qiJ/PQ1CANmx0jrwW
hnTdME9oey2tCs4PUL+Kwaj1qvYdZCb/WAq4/2ce1EWGdAc/U9egiZLsag2GYeoRXql7LVkVoSp8
BANEeBv9z80aoTOoqxqsDarTXWvCT8989Xw7kapPBQR1WP4QzfIFI1YAIECnCW/FRt2YPbYZkiV7
REre+3M2DyKZE/pR3nF2jAXnUrppsxlq1U6K9EDA8dnpzJlToZHSA/C7swsXY8wtPUTL+vNiDjnl
SeJztg5GTxchtWsWyEOC0SDTXeTXTQ9J1y64JEaFhJBNPKDWNyy233wLcQwuIXu1ta26aMwpbbq/
q29Q81iGV3SDfYq6ddaVgrZJrdJeGDSFjcwevzihtOxa8/HVhTwtIU9XpEkMYgV7BDd3WcmAVBpL
+gBt02Qiifgb5zIOKFH4yml8CvA71gpIexKgwrhqY4D8EYSAnugrzD2ZQ5s3+R1tVPvnOKiVDlw3
mTXkUFucmiTyKvE8TKrZ3L+I3UdadH3lfHT/VzYe4N62nl0B8td5RnqabL7NIOpG3ghXJWrYU/6m
lLZcdtXKGhDNrnMihOJr8Yn7jtipLtXEtAR0xalznPCN5eNQ4bsnIOpaLSGgrwGtq/0TnUH4ilb+
6y+yVC2VKSoBvrKXE4Sprkox1RB+pxBiOiaJxZlz8KqLABw+haAylwi+QreGYNFh/WKNsIPCXkhN
mPo2KPd9DgWZRzAFc+yonbNbWAMpMW3esTpCwv6ndSsH+sd2imT7ARDjh8ELkR68pVRcaLCo5TQ8
1/lNTL/HKv9tmpbRqFvtQ+Pm9H3PyyrqR0LqdM+jTIj2DTMsCrdMyeQcODnxrd11Wp8vp+64Fq5M
1W+5qiaTYJTuYsJyYrGAXtHBHuVAtbpt36+BjqtLpuUVVwQHdg8jxQwfVyZmB+sNSL3loy+QKryr
xv6VHVs/oThC18c65avnRgcy2cmK29IKmQpPNbEm/oB8A5SiO4iyJ9FQ5cdRs2BF91bYyOXxhtWh
KzbDY072UobePB3AV7iY9cHfrrOuhhwyMZ8EI+vQCNKPWUczgR42rCTljwkQfbcFwrYPMAukzG61
g1ReelF6dwgTNmgpGejzJ4l5PCel8RARTooTJryL/pysuOWcDhlqviDTW6hEmkU0RgoFTfIEMSY2
68zACyTqjxzOxDSaZiCyTkkmhxbRb4X8pazovW3m/nFg9RqrIsOmUd9yl1Nb9Zun1Lg5UHVURhjN
PWZ+cd6nhgW+wN+UIvHFbUefmE2DJ912H7Bkk/P1J5jIvPtX7aFeugkBTKIA1tezpdvJp7KKSoXz
RBovLKQLHE0GzkEGOcQhPKzB0fr/qwzCnIdltI2Vrw456VoYoDIp6/KWoUbbuo1IeXh+IHrrF/xa
s951KhY12LGH1D1Za0GiRxQGaapKv52XnHMdV9lQUKtNEK3pEqmkkNOoLy1sZyyoIjhEvAP/5Gcv
1KapDaxAjfEBlCzuIxahu3BVHfMJL4FmUlC4Ss+NihlCskeaAWe9S3OlltLYUWHSn6LNJFqzFIOB
dgUaU5p0rz9bIAZAY5HY5HB1R/avfH/wQ7hRL9fx3MCpQVLJqlMgwDEedW7KtldzpZsRuSUcILuf
jmYeIs9swFkunwdjMGh4KfZ+9BmEw/zM7gP/AUx8U/IyKR+ksF65jyCu0D7O8IJnoIWiVIHwT1iX
jcW77WWcVyo4URO8eaZSfV06y6McacglNTrMWGYz0ClgPfibJN8F7URhKT2HTKok8nx/gbVmLv5U
2CRqTaewTyz4LV+TEJSp8G+tOyrOs3KTpSFVRkUd/S83IJpgMQ6eW17hOgu0vpZtP99Ggfsj1Y+Y
+AahhsnA8vxsuz9/hQaN/PcEzxEa/5XtmWkSHQCT0XL8UgfAWaymVhwe0mWPFp/t83yXBKBKYx0C
41U89Ta7RdDkwMPeZ6ysHgguIa9NnyxP61qQOpELeq4ndoMnDKTrSWzPFEUg841+kqJ2vfH8FM2h
HBI+uXtrg1Dl4QrkZ9oQnaizCx8zrvzSMllamKsNbN4hPtA8zthJeC+J+0S9359zQmMUx838R/LT
NPBnZr7GegH8XmZjmXUeST73WV9IPJ9KIkHbfIHhhX3UaVkB/KQBtS8dE6iAEEd19MYBvBpVoCCU
nV+5YKsET7q+xLmd07k9kJbyjjLjbsVAk4fq4CFm1g1QyQPqJblmczMPOD+E1NfI4wx5AW04AuUf
Qw3VUhey0T0LIjaBCyQF7PWjX/9kbJ/4lLcGiS/3dnu9bCIyiz2TR/1LGpPZOslXS7B5WZT2EdS4
ON9qUG+UwsaZVzGYnERYo4OSGO0oEqXUjMdaqZuNlWmCmPSoGmLnZ4rF3x+XB4+7QP7pBzpwgXwX
B8yZiNVW7H52VmJimrrydVe98Ul7TQrgvpX2cS5Xu6/H5ToqZIdM+DdXUGEVq4cWQh4coBCpPsmP
yKAZIcpEvDBfLq0Y/Y/8sMRCXS68Xbn8WbMgg1l25OBwL8yLWRKKGGL5lJqStxhot46QHt2WBiM7
AsH3/nWrJZhLHcQP0NMrus7+4elGMpPJmAnsmaPgSEEW8cunbIsKJ7m+3qTN6rcV+xzC3v4k/NKr
T3mQQ2lPkH7CwFsUlX7moyOCceKfdxuLwKPoJROexqGrMZ6uPfRIIugX4XNLNtULCfGd+d4E1BUh
+JolTpdyj2+eCDJKENeJM8TAVF9Q/C7IhwuKYiL8uN0eYZVe80nilyvjdXG3N9MJgBx9XNQEbbT6
lPlvEJ/VtcQ0+ndMArI7sZRpTxE6nOCSDJPpel/FWiJQy5UdsqHv0dnEFizxGX7lX5RM1u/AV80q
o25Qi7w5o1ZieJ9nO6YG/Q+LdAjjStx24cDScKEJpa+wMYEbczAj131pFty/lFblSGYQmhlgLK3Y
tYGURuRe9GBZDvIhR9MXV4V/fWtCcpkgZnsFkmc1bII3BoHTbOonkDTukvCkGJyG25952AoH371f
0T8Ov5eJy691iq9LsKMjXk6kQI5SPEknsV+fudvord/I6q1uk0KqezBtytQc6L0qlXaO7r0lDG7N
k4LQlrAZZIVg5XTdJfHiNssbqHP+6NhSjcSGDIWVOgqo6ul1vRxD0NhcTTqchlp3zfmFCqhiNsqn
8UwDjqxbKEbn9sy7HPTTdfROidjP8PlNB5kuKrR3jlWkCCu6vlPTFxKIzmqpRFoEvHOvqlemJ+c7
PiZIsx3AY/9hs2L+Vdfe4rLuVgPRtE2nWgRKRJPcc4M+1vGUNi6iKVtCFeRuB/AdBdqriHSqEHro
vPBByptlnD0umseJRZyDf35XcL21RM92IZ6KJojAVhk0Lg0J5wAY33bqB6Aez9BGi+YhFxRPo8pY
25JbHeatMMfYLpocOwZE598SZnqK+bSH+q6zzKmyVBHhwIxoyC/X5bRK3zDFLmdBMUchjS2T0rF+
Bv4JRkNi7dcMAWIke6sL+cjtTF61a5zDF/Rd6qG+r1cixErTMx1ppfdzHqfEF+bc4Cv/ji232oPO
m5N8yThA4B8PQ/oWBtCCXHExrW3EvRTCRFIIQ49wmkMoAxoFcsj+a5kuWrCLAcFmoAcRRPd2iDDX
jiFqUbkXeAEG3keJML0XQ+2dw7+/ekrtD1n6rFqe6owANRsFJPWReB0gAuAYuHZ/Niw3uYuPRSY0
bItE6YDEWqkkv+JQTaaRp8hv0G1ar81n9l8ohy74LAdx2qVD9UPOvtjSwCRGX0juUmKtM+hH2edP
ZOKocaCuR93FxHpKmwRlsmMsi396OSP7A7WQuRgq6B/g+Z6xFzSmaMyT3V+zEKAMMMywMNujkeTU
aTwyRlHFrpnUQfwSVbO0rGnS0Z1AVM6/tVXhBrisGavp1ybVUp93chdC2WP8c8ngeFiC/ksdvauU
hOO41+REqW+BmrZmsmKdYWoA5wD09CKqpz9hjOgYdw+uhKrbpXmgFWCK4XdDAo0Lct2PCd87ZmWz
JxVJgK5Ozk+cH9ytWyiymw8c74RR3CfTPZHCGXLBup8OitTb7btsclrjIVpnCG9roK2hijgXSVjt
5PX11mAlkI2onnXF51BkCwNxfi/5tm+rL+WOtOb3i6snpZqnDuUYZbKSxlnrfwUHrRm7aOJ3Qy2k
+0bC32Z5n+NmK8X4OYJ+3adM/h4pltiYUEF0H4QeQIpdoN3tE7J0KntRXCayR4VYcNsE8T1CeWJm
+Vz8nqJzH9s3CiQuAPqXE9+H2H6OeFKXOJIFZK+dGb3ivI+W2mVQHBE1AaQEnRRB8L6Y3x66dfV/
rvi3b+EolFeyJVjIkzowsHmvuCuRH5GGQQrHqzsTySipHciz1HJC1/H5BxMK9XzK6DduNPt4O8Az
+dF315r5H87itx/OxPuH3sGQWmKnxFi+NAqkgVCGwmOVDcg7kA62hagDvANiVUrPdXB45xR9RpNs
LJjA6lnQfst4GG+CunBMmiFYPxFRCuktItp1QfRqxusFuSVAxdHo5kaf4eOR6VwPFQXX5/l6T3uE
fU5fJuYp6Ktdgt/pQuHx4piUyeJ9JhqWPnSHwh0lTBfQ7jnCPnzlyUerIOBUeYIMif3AhWiGOA6v
ZohB1mx6Rbw2RlvljUfni+bBHaxPDA77i9CfgJUjsK9PhUwTcC2NH3anoN932WDiCOrIFPL3RJN0
MOL71ryLD38Ds85krkYMI3Si/w6SrZ8CMCraWBPsVSnJ8UtlY+EQhbbo7ttMB3FhY4hI8D4/006L
hk06HjJY0Aw5Bvr7x8RIGHHwOPU+WBuhPo07vNVZeF9MGIhNj6rNdBLbE812ZiDKl2+KN84Vut0W
3nbvqdRcuyDpiAmFcU4jpXUCLzHp9qxwn903+uBwX54L1PcIS8wBc00nKM1vAyaNMx9rCzXpt0Zw
zyOKPPtuSUM/IE1l2uXsnpSvWY8O4dgSyer5UUrwumlCihu/GX7XjDQ1rMDgfHgPySQgM5Ei1QEX
IVBhZ9gC2cUmOHbxVkBazVjXgu2ZFv68NJXYgy8dRqkgz0v4jzmii19aeULEhXz8w26ENewVD4iG
IJ3HXev+kxgoO6ZFe791oOK6EJlKjOXJ/Djen1GwuC2nNPNgFbJ51gznAK8E39nsJ7mlb91L0NmR
cgNFOObjVc/Xr5FJ4HuS6XoZ1c+YCWZWumrjffkw6BBdYevV+vT+xgBowWD2YRPeL2TF7QOTazU+
XnUum3MZtkZYg9NfhcBBr9fEff6gC1rsNXeTnoM/vC6tsY2Szi0l6jRRZ1nY4BHClQYwUE28mT1f
CM3E0c8LKoWB6y9xLuM0VE2jIJnve7QKb/8C7os67f0F6ocz89dVbX4g4aFrpKTicExK15Y5xl0I
nNG/51ztKQZ1k0U8+28xIjR311h54UDtDYT4u40cfu+Ziqv4HgsLdeRHbF5cMB6phBBHoQbBeHan
Fz7nJFkwFRzRkixqdxI+d6Kvwmn+QNe3UY49xicnU3PRrbMh+VrIH7YH0Z71xgYilTXNaaXZ8nqV
fak52WFbaQO2VRRKV/9+vD/4PXQ4Lf4yRBphYj6b6C3+cATSkd1ydBh6txSvi1El22oeeVMo14VM
pP+77sp2iEEzxhbRYVi5GtWVtO+AKZVQ8AqM0u0IJzMxEFGWGn8GcVUkP+fXh6jOZaf07Yo+uFk1
FTOCOttZ7vFhgu9miEjKnY/yycDKJ82ZOWE2D6CSoUlWDUarbVW9sTteREZgIgjY4jX5rDHgOLBZ
5pFry8e3fOi7xn3zv1A1g/gJWlU2nb+d5OoRS4y973MKHDJY3G+kWTD8y/ND0Q/jp3nJd4/bQnrC
Wqy34kvuxrKTV8mUn+m0cNZRmmVioXx1A4vPlwvew8nxioezPe38DqSoqw03wH5SvL3mZH+FlQ9y
nsuxYvO1k01zW0KK/IiYrXJJUOeo6BZ6ykmeCQz6HxbRTI8k3t7728Pf0XnzEdi7vWYO04wy61Dh
P/uksQ5kgg9ElTF4FsTqAZa+ZoJjx/tc4fQXlAEu0o2c0ZnDsQgtZPVRg2i+vZ3KW4azikVk0N3b
15Po6IhRb1C23BpEqH+EFGaelFR/Fsy6lwOvBpjOxlLOg2DvV52TXy4el3SQQ4pV0BfhvFctfAOr
HNAxF2HB0EtyzoH3FnUl08jODL70dNlvyTgRGbLW+t7vnuENRi0tt7wTX6aDfeiFciwm8cILyjlL
3Sjtt1ToH6D6hO3ao63V4rxmDyNZVDTn03KdFbYy+FPTBWhEXDobkCn1kNhmDERhfY9sZfn/fbgd
87ewuupyXnbnHf0lEEnSyUN2c6H+rTeis66ZEbdcZHADcIrpmm1hyauzUPotb5voN6tXiJDas+mv
svPmJsGDpg3NjY8lhZ4oJXVD27g+NW+uRm3olNQ8Tu3VwxEAxd2+OnRTzcGJnYmCx9oRLJtMJOsc
3lHFQhIf6z1EJ566LjSxza+XLQt8zvG34Psp4cAU/6kjU5VmS7K3TitCXqeXhjRkjwThYonE9QrT
2IhDhbNeQgZiUMONwznQ/33/B4RlcSOMlpKU3/U4uGB2VlXFT0ABj6sMRWqAi3S6VlOztZc/3pGj
KBxaXqH3dIxD4uoKMiqlW3hZXBJZ/YwqBK9HhIXheGV0orenydub1wnEVTK07mRNvtHREAite/uv
ujjueTq1exJopuQsGbOFRZ/G0QQ2Zh38q/dIqQmDZyGEj3BH4C3Z+PC2j3C7mB+kLJetE45L0DoK
5I0SAsiNVRCJbSvKjwYjhsfEz3JTmjHX4uLvDUvhTays9X95njprKeyFg6DY4Sqv5YEJlYC/9lZ/
1u4Bd9zP2Y07mW4dwmDTy3lY2AWU0QjLp4OQhyWbs5IK2WZKfGcZWYPehDSYX1vTEPO/KdFHSPfC
WQ8R+ogq4DizTO3k6om7i/VIw44Pfn7JfSlWQ9d/44X3BW8RMAETDmwKt2J3z6UM3E9CS8y6aAsu
ouhJis32Htv52nwvOHfZTvLKS2Qp+APNpWg5e7fRf3fY4ARWUpVcJjueswS3tV+5V0exk3cHd9K/
OQ4Oxv4oy/oS6QRfUxsqTWqeIx6mGuViBvD8r4yfulgL75TFPmDcD1Cf39ySGf4mwBUMUm7i/xOI
i7erCMEgaTCaX/f/libIMRCuBgKNI4jpSJsBThkGJ2sYD4MSycxF9RrL9gsN7jfjO0kATZwSzcac
LdZDgguwLysABzUualxmZgmxdEuNVOr6ccC+giKl52EdIyaeume0esaoDZ1nJ/IIvyjYg5avNbPH
8Dd1yOUngcZk+cDlHcd2U6Z0YU4sUKjIIT9QS5RLvdcJymEL3pUHUDcJOieGowHuy4qUppFoaLZN
QCU3fLDNfSjHH2ABeLiDftIZdyFNG49ZKiqIsVzl9wLt7Krtced2jOealcCYHJLs61iYXiHReL2M
KOzGV8hWszn94GrkVZn/sLzDJYr9OS3XnZnnDjfPmsMcfaL7sCORbuTA1cqNynYfQemR7G6UUKCF
t7i8dQw9OLV1NNAgj3GkOCb7UTaxwVWOqBEQ19gTqjLJviSNhAlByEXD27GwUEmhU3ZVnfyBbNOm
UCdXHcgkLK2E9bDmoJoWY8t4Sgc9ADN8A2F7ZxDY+AhJWtWAnJIiwnVmoPGY81aIb1NBqwj3JQqp
73EwnjQsBVezKo5V+qVqKc3CJIZ/O2PtnZtsSLy3vNbZvadKZTlI8pu7txEZN1Hryx1uWNI+U4HZ
9XRqEjhYirljSBi1i/SR1/ULIsdNlN/OHlxPDAH/E1VzGlPRgtwhHwPbLdDyUBaLVTcqmmQIwYRk
lxVXV9uDRkCohOFf6uu5Uwc/9K0vubJzgufEGFLSAapnaW56bCZQ20MSN7ADMT4wkjQI15uzcgdi
ctwhX74BD2LLsvYAjb3p/XagW+PhxoKSybFhiC+6w34aSlg3igqRNnlfBS+uihvj2on+D38Ngd+1
42mkDGZ7q6PVIuDSawZhmXBMG27ElK2/5A2eqMMf8rqaBae86Z5oHvSVur/rQEAjhB1WiYRNTbJH
26073/CIPmsbkK15hF0yMOaysl5un4GcjuZJNGswHjG2VjnspfyMRurUviVu8Rsti0eTGH0DRFaY
8WjWae730paOAfNUm2yrsPWBMYqaBcY3422qXhy3k++Cok7H1yHgyFnHPE3QKwijcvtnnnzFz8FY
qmzqAirrxtF6GGSnhil0zXl6yv7Nk47/ALgot599+qK2+4rS4Hzc1xg6mCJB5b896kxkqQylp8k/
r4z3GKTAbQhtYrUPBiatHNO7xxBMEACOucCmn91LMDK/MQRl8rJ0vQ6pyp04io0/bi5ihS/l2Z+R
/B+CZwIxh+EbrXcuooOC5SXHcxMB922up+Nth+40C/EugZP0/q7srfqnjBZEioJZ/fQPaKUauJqV
EI0daetmNSQCcHLahxhrcuinZjqeetfb7FHGOLgRhMXvKPabzfrbVbZx8QxkjlrAqy7dHbXbvs6A
FPLpTo0BjxxGU7onLPwYEE8FTBkOHesqTLX7veF3L/KWWLhO50T4FTg/hZBFNs8GKYMVudoYbt02
KspTgjTciJKKCbaaX6qS7KeaoYRQNBblNo2dzax9MIRsvPZgcXBhQGvRULB8DszNFNBi7VwPK5Aq
c7hjMVi5LQViet1AyNjjemtbJ4vho6ZyiJyTM0yPv2mQolE+9Vh3FzxNFMSbLAtUNkZiIm/ruy1n
+MgrmKBefJZEjqA4KG4sgUVFjgx72ZMvo4fA7qoHl2wiJttpsLNOwpiK66uoGhnwQeSEEnMmFf4+
3eqgGZ0MIv/83BlnSlpUPCXOZiApySQVg1x3LBNEN7hXCtHcRwz+ODbJgHlA5lGkwPi32BjPosCz
l+17/ivipFClWRMpCBgPfxY8AzZPAc8e1cj1mOWWDyop9wsBNT061g57KykpjKNR1JzFuesysC3n
hu8X2y6w6IVvgi8bLnVV2FzD3MCWduitdZ70cHPgRTKl4CmC2ZtS8BliJVauMpABRZFpWEAuVw8v
6gMhlaHlIF8WoKWzhxBi5XoZOVc7/WvO0nfwVJsI/n05+IwbSl0UcEHycwRxLnymISRzZrltCptP
kwrzenNek6AD4A2IMh2pbbPuOCRjxPJtyywOXDTGpp9WeX0J3r41xMlgKBUz6rb+zDhBN3fo4NUI
Q1wcxFWvNvCyFkVOUfxYNIy6uoWKISAwb9zjPAcqw8y+EkP/w4EnwP8k3zrFQ1jTHywJbaiCdHXP
mFPgFJgBorBjdrBW0tTeW2MbJoRrr3MA0IQDkQSIVgaahfEOT2f4sCmk9oEVDXXr9EfnX8LjMYKR
Mix8AztGHGVFKbglh0pt3wwCGsTBd9ieVgWnACzmrW6Qmuvl1D85Clcds3+bakfW3ZpYldrw2ntL
RtwTjIBpwiP5E3B6x0s8h5aWafyXO3PnXa1/UqKUhIrzgBFHG9sF0IWDgHXse8kPLubmi58TDVaN
crGIRLncnMz8htztdb7cNIapTnURXXUyCGjk4/4ZFwyJBtZQkTZG+BU59dBDrtF7/mwGy7UFULkU
GaeeRR/HQd+4aybX2Z96QGBn45ughzGy5zxnVq2PRWMEpfJAsiHJX0qtWZzyo4pm/cPXlzavNVVb
AgGXrajMD/4kYFz4rS0OYNbhkvH5/NVsfKP0oXS2hZ8enUJyQWzIP3th28pILijhcjXEcvY9CEX1
rdD5cZhRqqb6Hix+AGoHKF7DkgLUpWU4iWtVo4qUIi9hxU6E6cU1NRxlFdlDu8rW2QVSripusqxp
M3utdCI8eFxnwLQNtDjnII1YXfzEWtFD4H0aSNMSkPAG26mRpUsPxpOS9m9zZyCNWgSdwv2C2t3C
XuBVBQNLIXSmTYeF6rjJcEyjm1N7ps/vMVDfcUZMRnXKviUXIeahRtwG3yArw+AohQpOJjbz3WmR
MgN+RMtQm7k6qfD8Xz2lkFF3qaKuH+J5eosasAIDybVe1yVFCjaoERMt3rE5BGI1ALSGhTrWfOBq
Pr8zjMX4AI8RsWV0hV7N1NcR8vGL1ejuanB6uTOUzda/QkiAwd427iKAXCIC2OGYj0DAplTurmjq
wj2XpDRq+52uR3CqV8xNEt6/MnzbWFqVm7q4QBzwm++UF+NXipyPDZvg7SukZmIMLsB9hJZXtScf
7EgCywYEWYKV90cESdhD56MIah+y6OIXt4vt9NT/E026efMRE8EwsqY60Nbjp/DlfN6mYcecuoMh
XqHEOD299BTTxL2n3XH8QkjH/QX2y9iJD9plCcktIp5v/TgLGzUICKg79e635xtY1E8ocPLflmTu
qRkFdffU6LdXDOwuayG1O81vzeqnX0yqwlwxxYn8lazjbd/wsLma2oQAE10ykdPt7CA20HwDT9i1
58vXcHrnNnAr+PpnxLuSVxluIZax6Be6yibaXODCjYS0nzoXGNrZfZTHWmkOnjowQCNKCiC49Yft
X918SteCEl4Jy0ci0Cl5RZEh3OEQZz/hsO7GdepCUs5HXE+/5KRM78SLAauEn7C/1UL5OM8wFLtu
aLdNfuhXX+42PzBN/1j8Z8yuV+x7VOmn8wK6CFFr7mmWpmzq44ho1JueJkJf0hNijAf743Au/NvK
vgJ3s9cuFvxUU6oNDIVNX5toRFeLL13GyCKW+hfJkuaiTosc7cJAloUFU4M3L/l99Gz4rlA9ECdz
6H0LoG0ujhrS80yf2UzJ4GiOznKGGhx+EKJcHg0VTAWGI/OT/JDi3KlRqNycpmFeJlrZWeDocpKk
mnfhM7NhsqEZlbpP4zmT7iD9KeD8w/HOntjxC9HMxbJeDLSqxdmIxa6vrdghoEedtrelLvkDm7Wb
9juWp+VITEuRnWvdJ5NT28tAFhPEp654sSuvyfwL+NS+Bnlvg3ng0rV76txDsmk3C+d9bUpGcEfp
PF/CfMyNgtWFgCV6A2Z4E6BxJyn2lPe7nT8Bg/kD0O4MDTG4BM2PekR8HzmOBfyfUdpdyY7XonAS
iKnoR7j8ck64PwCAWHB/6Yh4Lm4NxfwSJ5CPBttVagIaPH9k5d6vrP+KPTQDBp/EqlC0bm8ISnan
cNca5+al9HYpNxXoAUrNY0z7N/UxaIdAghANhjrHtLasq/hpMGmmMlsXtI8C/acF0Ol5FHnYtju9
PD21NbECfB5epkztZuds06kg2tajHnLrBv+1xRobJ6xCCOm72Wpf+sh51aKp3n9ZB2vWTX1lKbEc
HNy+0SJ/htSJMiWVU+7XuuXYXpjWF9w2YtIANspNUHMVx6i4mJ/dkPdmuyQ0yPKJze5npuEyT9kB
W7ONjoRL1671DXymr6keKHraQDPKDwjjn85cXT/tgmzi8RuU/MiQt3OZGESoflMVjJrpS6NTgQLn
eRJJjNVVPhX3GD7lS5fmBnNr8Jovzjw1DQh0mpZr/eUQlGiSNt0g9iH6HAyj/pWcA5We0f983CH0
LlDEx2ly8RuI44joCy5F43SoEbcjFup2D6/4YPGrG38PnLKFTGblelPI8GpFnLkEGT5mxdSL4Wqj
Iv092pVKnqZiwlCPgKuJdODuG9y2iSbGiPu+Cj2FMdI4vIzBK7CfS3DozkOTb16YobjvSiDdvvT/
HjRw4pbemrw8AYvVdm4C23GZjghJ1YMtfucX4RGruHNcFDuTMQ2sAEBIkY01cQNh05wpsopDK2wA
LCCM9TubOfe3AeeGH65HU0OigVKa3uAJUo9i5MrvLkD96W5JlEbi7SmbYSxIUxpNNE7I1T2n86cR
xn8SRRXjGN5IAb++LZROOQbC38vMm8lIiPi4iIFPU9hCcIeStTPbt5n/dhwki/tmBXZfPsSf1YFd
pwBiezDhnJFmpfzR37tcu3CBDxb+B13VgKp7/7+o0bR7gNRkJ6ZRqIfI5Um2R9x0BJdrJlof7ERP
fAAzbhVKQdgdteKBItHBVssPJWo4nMMVnJvD2ZYHzSFSn463nXp5uRhJjlZAE5IhIbOYX+mRfyg2
+t7NBbeRjq+oCQysklUSvOvjMArLNy0tZjamdTxxumCqMG/Bl42Hsmsa/8NxQfV7YRf/rxBjOzp6
mtqdstYLSCkdeoCF3NfscQV2rHny5cLyfM8ZJbnxH8ejLLSDJF9+4/Nk8rDW2EF8hOSo4Jd0jRsQ
PUhOd+UYC42It2TMEYTLYeplH0dpbI8aElp7VquisGFU/qxfKYj11ocW8tP9DWcj/PEf2CvV0yO5
J+I26PmhUBmQ2YFDEY9spCbbabGph216QLDcYbEnQ7WPY4Gtzl/Z2da1fdL6BZS4Oluee7aGoouq
JHMp2Ce6oL+yCF7A4m1Cb81rx8DgG4F6BalaJy+qQsA4XTTEMM/f/kh64J1+c05GTC46IcWbAg/+
FfR2yRyKmOitwzsaWHop7UG07nvnHxFnlg6b5NtTMY1Jcw3jR59M0bDl7eunEA8QUqEQVpLoTZbj
rwree5yK47gM8mK0al3wS9mZV+J6Tdth/U7BFfGB3t/vdEQPqKrR3eisT5Dqp97Kde2Bv0BNT7rA
q2o70zBudhxvNzMJ+ww4aKPjOVxn36xK6P/unrnFhS3pgrQn+HYcrbuS2ifuhNfiEFnX861UjgKA
mV9xEEKcL1IZGFQGwHp3HCvGVDwvZbqHf/kpRDyRexpnDasqFKGmzDxUztIVaPFTiBxptXnrulPB
0Zh2l40bjipPn37tvFKgReqTy4/nf0VkfJ7SHao3SGsCYBaoLqm79U22YwDkh5FZ/FIzeh9DNh74
C3xVIoZJ871qf1E8tTupiB3ySE/90D0Hr4eznmaJBwuYp08lGXHMmAVQnd8t/9EDBjeYMQqy4dKw
5o5tNefBc1MUmqA7sr909NER+/ix4TuNl5uNIl/2YkS76hNgNYAsMnvoq3GUpKJwJfjbbkuC706a
2kDFUjY6O0aA3Mk3bmXdIkL+rCb+zWMP/MQd3tUs/M9zAW4rE99xfzImVS436mkbHyyYr8hGiiuz
lDULfEw4Z6O+eTya21Abk9MT8F+JzVgz5F2NZeHEWb3VySsCyjJAbnBXqSakXWFqc+3o7kCXHx5B
wIDGqCv1EcGDWjyq+T9QHBdAX+Rtw9lxwNApf6CtrTMaPbg1yDg8DgfJV+Z6dfDHQkAWRsW+lo76
rUlNVFk2lqTieHA5/LDmnOC/1xf2dRItbkbQDJeVHTGx+JOovhT17sRo4TNShvvrFDqzCzHQgWSA
1muYwDO3D6ZGUwwKA8+4W52aArs2OIithrft3GMVR3Z1HtTY0BZp3RttTHfUqVRJD6Re3V47pW4z
xAWEhIKhwFhKEsqctxdyJHtemvTysy4b3s2kYjY33gKo+jzvYTPsrBFIjFrjznE0bO+21TJ11QEM
FN7yRJl0yQSozcaIxFaeO6i32JcCJhO0mX/qnHajp6dlYsFLTVuSvUXwHP+pU4jTHOmIVbOA47RC
Q9EzjIDHZCUT8hoUiXu3Y5NwIa5P/E8UlgRy0sFK7L010L5lrGxsjzh0X2hIYWjLJsceZWgXP7Q0
0QUs2SVx7SZjCFscEIKcXClkRNXfzmV1Bs2zUATrENj0cnX/yVSOtKHIUFzxVGRi9PQgUqaf9xnX
sFBiB6r6D5+VAq1MYvDdTj+EoeRpkLsxn6Ap1g2xr+/14QLxA+ZtdlQGT4y+163Rb4bML6cqPr7a
93+eq8u5KI9trNR8cL32D5ovEXT8lHXhYSKn90fFvbLnsNbAU4SaQO+PUCX8w/2IUvnQxvIVmRm6
l9Wl9PzNlMcZSaBjzKTq6CcAhLMyoNfToKhCwahSBub4gzKjz9F9JjViIZ14Bxa1qTwRSqRJjYuo
HcChQ//mS3LtzdfDTtM4cU33qXGR9wQiQSq/prbfJia++c0KgewnGDCJ6o30rY3YSRCL6STYsu9/
p9fJWheRJP9Vc5u2cS1WxUtdJmfVichAI3LRlfQkpB7oeF0ZkxiVUB3WcmxH/m7oc82DyHYqoCCP
vI2bEmR1resNHqHAXuEl6I2LlptiCqLuCeQHpCKLvHN2WtnA8i/MKdoCRjsDztv75510fzel4DDw
uM5Ec8xojr/SIqm3tmtJh0vEuq5WkfmtTNTQRvoJPUV8WswRuD7WrmeLVS3swYhpFUoMpEQtioym
E3YnuiqRzhegUkOkTj7F6rMSUq//PBsihNIo5/xNpUHpRBHjTmm9lr8giSF7qsQgL9OGdLKdVVH4
G8eLpu0yv8l4kdMNFiAk1BUnpT5TuOgDDuLLj+f8GxDQ54vv/kwxvQ17kDmtIaIlON4Mki8BhLKZ
A3IPJolK5XSRYLHli/SpEv1UGKRaXGKem04HHRl8YfRdOqRiT4/ueWnrmTO/khEj/O5KRrBkD0Lx
pl4q53QxptxRlO6T3NcwC/rQTTX+mgt/Dy/9xA3sOfDvMmyjFAOXYzZrXyA90XGPTMjMaHkPrjNA
4luSsfmMyqIYWJBEyCfxtSZvwTClHQz/bo9uFZIb+B3t6Twc2Yzz0Fr57DPsUMYFuBA1Q5IKDyws
yBStQuxFBjgtCmaf5G2YuBvlHzfSFKDSsYq9F02/fNZBJWl3tLEdK0oy2nb7UA3xfGGKB06TpaiH
UyEWm6W5MzCz1CBUnzMiSsDjF6nvjUbkzzbkbtSf/+dvzFbEdbd+q/V8NGYVZeAKAhi+cnHrWrn2
A0cRUXdfwgbUTIxU9m6VYS+c+JISsK7NLLuabcY9cCu5SK/+kzVHU3gO4zz3QRVprUXC2ETRQyzP
v9XwA0QIKVLcMSlp8/3EVRwsHjfYff7GgSN7dH/X4L1BzRNqb8OZu4Rboj0IP4+6dieUV9ByWYoo
0TQGGlqUoMCQQxTAy0GIEqAE9FHVpe8W37YHfCPCy8JvQf6Jx+9PmUyvURNa50h87084xCVpBKsb
kP8huSyi/ueL9jkigF/+nczJNrhLhJNOc25WvJ6NTbFlE6IGf6ODFLcA69v14gklNT01tmlc8/Fb
aCJ24s3ygvp0Jmra8TajWXFOlqmy0hQtyip+tIK621AFdDiTnlFyYX3rKQ4GcDaATSI2jO9w9o+S
UAosyNpWNpH8VWkP3O8Gbw0R+hrb14yUROZQylO6TAh0TI7TfUaT7/KE3oBozU3PTOxRiY1U95wA
ET6ErQ+1WjB453Ftv+fOqdrMLqHL6YHcEXRxD6taNW/wcwJn7S9daBJOTbWC9lIcXvWNj8isbLGy
K2C1PVnKLr4Xz7V/25MhLReTOV9CkBTd6GWtULZfZi5xZ9jDw7WmEfZABGByenm7T0ns2iYY5xJV
EkkWBchiHJnyJ1sa1+J4/HDh5CgtIycYQP7TL36UGeDLSAx9+52eMws4qIdLo5dDnwyZDnjN6qRV
H0xNpvXl5hMHALBRnAHvS1DNruXOG7FyGAYAfL8lbpK8vCYNRsA9LajQPQk9ph/LwROMP2iGod6S
UE4Nmwb9JNQ5/OuUqab9V6+h+DQHbpfRauxEoVh5YRHDCE4Pm5NLZtX/XdT0qn3O9evHqHpNauXC
ed8Uf2QB/Ny/jkPOUqvurPrqlam4xbztGLq9dfOKlJyhD0jyEx2NwPaDYIFLvjwCLHFBV2/FLpbM
TR7ZPlDkalEAe0Kr0yFLjwHDzK6HxkPQjMmgHI9nXu/ByXyEl3bfShZk7yDFrqHSpKWUz/dwCJFd
C97KqFQ+RRIrPffhlf6bj+RwLtRv3cjFrbVKpvO+AxzZspEj4MZhF3jX4qYHQD9kXkld0sTqDdtT
l2VTk7NGVyrsrAf4+KrAkKXWIiaWeSiAWgrAV0/ty/NzMF/YLgi4rfsZEYfUDulOuUq6ZnboLag8
MMt846RqnBG/EeK1nwn9/KztbdDJka+Kg8hP5qpdHARX3imRDj4iXhZU/eYuEJ38BHYOKW1mfvN5
mfYQG0H+4EwemGq3SddO90m0bTz+m0z5GKQRiaWp6Pcn3rhWOzQ6J/spAnjVGergUY9KSb7b1cRy
BUtZKM9XqthWic+x6okMRJMxdt9b/kvU+i4wDgfoh6peAjRIucXhGAEzv4fL6oYcJYIwUPisYLzD
F97Aw31Od7peKueCCG9GTvA1NA+4oDwunQ78vmCzUda+mMxewEfZHeU0Hnxcas0yZYsNILLh+doO
vHBqcwFs7YtdLWffxZooRHehP/E11iiCDEIlDQ7MdJM7Hl4wTw5s3CMQrCFoRF5cqFE7AYTxxX1N
WRyry04/J/omPEDdmqAKCTMm6XhF8XgrCHTcxM0eRvnBgJyquRmdJhAL3AYqziuV+aObztBEFK96
oZ0sLi5RRmZQsRMIQq3Tp9BZ3EZ+WYbDxiVwAJjL7hMC/qWpGcrpGFhK2LYADPQytF8op7deQVXp
ulnF+mIvAqrshs6qiD2DCCGk3zl7xCv1dmGHPFTeqXisjvSgDpHlNiEEHqG7/87tdcniDJc8RNen
UNoLw+VYK4UuW3g6ODXstjxXv3XqiuSQplwRDazRaCXciI3kIFvRAEV6sVClGK7J1XQuXGtxEZBr
UrZwCDuIj4v/s/+nUNQhTOhN/EYCn6TspF7U+xkO6usVJyjWj8KhAaj1nX5pB+zQ7d7U42CVQ8ZT
1+8MIHgVj8hTuqFvKSnMX7MVKGpFjOWNWzXtZk7mMJ3tKqCOkfWS7GFMJSHl+T0Uf9IKJkXAkSvo
aBvYHlXZk07H7ZEcLaPSpKJhtBFI+by+F2ETudTDHkr37R25TTMNlQzBsxv4FJovZzfH5Egc0HmC
YGEjkYkAgbAVMq7ig8tcylpmVp92EFe+KIRdY7GYuw9M0ZDgsQYL03ygXICidM5v0p6gb1+atMS5
66Ahlr4Cu3UlQ9vH7aUyxKuZJhWQ8FHRGWsdr0/AmKZcJ7KiPTfvBiESCwdiQJ5es1kjJqlcOFat
5bORnUqEOk1lNUFvBsO2FxPkGt5vbtCkfIYAYEO2AG7TwW0ApOCgBLNtynT7ENLCoFRAQRocXm5i
ieeIwAkhY5PsjQKGjvOnAMpVZlKi/xDFZwYcuxAckFgIA44t8qPWZZMGYnNfMKI8xxpO6v6CMunl
IDU3EyvAEUnokczuI8JkWRp/SZAiEFSMU1ghkJsFNDK7llIcqWBID56McV3zFua9+VKAint6nRte
qp1JxbFuhdPY8Ed7h3RNfz9Q1Ore3fQORdLVHaLLjHt10kwdgV/CdqOpdRnzZKBNiZedc0b3u0XZ
XSj5yId3Z8jNczVQmU3O0aShVBQb6eDKRBnfVInE+lxqYjLF7oBecPvjsS/g4Yk/DZbKangqJFK7
O4UM8FIVg6pr1LMcV375Gl4pWqCb8LIaRctz4TQdbNU5l38Fy7hbuKuxl9NxMYqAIbbigOQ7uABp
6S5IVX6zi0ows3INjj9RBu8VvXbDVTwcVG6PgwvH08vUur4h25i1X1q5yyXjOyJ+yTphaKCQwBHk
fr0GpUsUPXiSMy5f0FU7mV7U4f4dz3shUR2vBSGq8tIVnshVN0ldFPcQzWKm6B8/E0K5015p93Ax
WoGcZ0rDvwA0VZmQ+iXkLHX5J7FZyw6Y35W2EPvt5foAv7Q0zemr5/aEk9EN/ric/dTlws1wbi76
78Puuqfgm8f2sx1ZTfIwPsNEhe7cHJWuXgxVFNCMQTXbtFMrskibydSFxrjykfMaR6rEi1oKrBdd
YiAfDaUNjVdukfkMlbydfb33zsZWXFnF8dAZL2LrG0WyLHy11R+4Weit2hADlPEgQPK3x8R0s6N8
pjHoKlSnRZ3MGZBBX7AYzU4YWMSGSRIkn3QwDCfACtTamTJD4/+lW2Ze1aLhfkAsm80a2hsl37Lw
pYiGF5X5QOtBKmvwo+zJnWUc2d+AFjwM10/JW4AZq9Zj/Rbc0FSzAOv10TdwJtDOsVyMXbGHlDiz
qvmZdCkfpETNiQYK+xtcNFfHRoC2ek/+FBlP6//nPfVFvuPKjmO6xoUgcZPMgIWQaSnsbqufwYuH
vSJ6U6DyTnK6NVhisB5DKhhJVHsuYONCu8udcpOutke+8rJqNiSjFiDwQJ5xRpcFj1X/SfRUKIKE
glswP8sHyjV0AZZBZIc8MstX8Hkdn9sxnDeK6MwNC8IfjHLnNDsxCPwUs6V9aDe7R+/lg9vdnJZC
ji5wC0D83qD2wUadHyLd2T1+Cdz6afDX9Xtz2bSVrrk3iRvO8ZToag2mykPKlWRPd3EvMpJPc+Xn
6ZcJofO71o7LDuwtwseYsVkzLlZqEmkqix/IDKXn7czvlYKUu8JzhmwScueW62em9+wPjru79Wb0
TNm9ymQSkmFL1Y26QisnU0YOyPK/WHJgkkLCWY1fBtqbx+bkfRbVHMd4hWbGBeb5YkKhLHjEboxv
7hsrV8T+u0Qq0KQx/jl++M6TtsldKZJy8E3GZOtFWrc49YgbFO0YUjmlldidZ/5KjBtbtd6stZVw
JC2py8iCvRdNQqByRaLfAwefPF3R3vfQwnHEWS18PS0CUQAqmEG65OWqVTARvOgWKghrbuQ21mdr
a03cSDKaXQUoes3gIpcPVngLaHZhEtm5mb7ZvkE6gqCcBq1H9bbYK7djKkNcasPiRri1ZV6+rnmp
LWrKVOm8aFYmHhPRH/NhJS2d6QoRFr2vxxu0L3vCE5bBf9DDlbU/jQy7avKcYsUiaNpBiQtKREar
Nm2QMSQV720hPkTFBOCi+AIe9KeHQMGP/dMVwaJ8e+fcmRUL0AR/UnKFL7t6mYzxhRDQ2T9Buwuj
7V22ZUtpk+RdOm1KHBuX4IiSXQ+AWQ1ti9/6KzlTy6kmRqkqFx8rS0Yr5aWra551skvJJTvVez9r
qok64IxrpN2U/2cwXPjwpzNZ3N4WoniAJ/P6rhCW23ChkJUyhOd93iLGljOCgMXbU7mntg5GHr7m
NG+Y4vJG9oomV4jg6c7bO0bA0+KxORzg6PBQTOmWn4bxByIjLZLwZvRwB2AAoq2ALRHPWvlz5XIx
3yNk0ef2jBWIgPt78VodUoCjQtETWg+1VvKnBSDcO4hsBipYiBW66IkDLXK/cTjrh0RZLg0/xzVr
ei8nTFnu1+tmQVlyKsZ9rh2eb4vp4eiQZdTW7X3bIbe6hhzShr7oeToBT/WPih0dSJhahxtmQzAS
cxfm1PX3Mjdujmgb7BqlE1/HntWm6k/tQXQKxaC5/XFh2WcEJQPPNrmdkEuuWEq9aEyRnt1eK6Fv
PtZ7Vax5qq3bEmPoKG7JFJ84CkXmT6zE+6R8QXHIYbZJe3R5k9gBKpR8IrjFpL1Hv880CO/BXaHe
gv3Ec4x8tNpnxPf1lKWQSGyLjANYgoL7bgAz4Qi+eRg1ceH1WdjOn/XWgpMGGlUdUWVCpyT8qI8F
42Xb0URVvRdiqbbIhXfz+xWiQY9aYLHOGwfkVs4D+beUwADkm8ipIEq82Si+e0cdcoxOkuUqMK3u
jRt0Msq0UxdjJVShiRUiSc9dh0bYtQDOwwDWk/kLFChmRTaKwhZtlsfMMW/kTReu+eIGil9Pq+hc
cHynvcjCAa7p6pQRHkwAl+KRNC2/rhJ1wuUSO8eVZxwyfZEpklT9A3y1HZmrCF2Y4JGNhdsN+uEZ
rId4z80mLt1xYbQS9h1G8Cu3cc6TX3Z+xK5bzPPH1kalhPP+6kZCuPfLv1bwoa8uJFdfZR+1KBOY
YC5skmxG4bd1Kcah8MISnvaosSYdd6QQoebxi8IAXUzr+0GB6gH3UkokEfW8s0Trhy7vkUmWh85L
J4mbbWtR5zw53bRwpxQnnybA4ROwmZO86IyfvKMGwaxzeCYrzpcAlclQweYaMVGNj0rYc4oNw+d1
GmgY9aBZNP4fNkswFh0rDSPnnaFomevSa6ZdtxnZXH+KRgxSp8m0xfvTJMw9Pt5HG/3LEh9VtgXc
anq2dPVsSr/fE8WIH+ER6dM9j13sNclsq/6fQgQdj2qLvx3lrQQ4kLsyNTCRdRZms7MrgE1iYso4
EXpydPj+zpmPcuhreYmCXWHs7EEgDYWwYRKld6V7fSPmqE35hy//M+YgeDRQ6kxotDQfO+CS5tOg
u3sYw0+S6NvQtnS6V0M13XLl1nguxs7fnonYPz4Cnq5HYkTWNNA3jv8975L0n7PiQOnMVajaFsTS
mKDtLBSA6y6XrenuQW0+TRP5Y96boamjeoSdw7HBv5sNJ6+udb44zlc8qQ89tQPottFeJ0SYoB5e
Yw0uQWk/BCl6M8Xb+nNjrn5z8pXlfmBerqSiSFMvJnqNpqqLqZThq6VwWB13IylQVVyRFXSnCI7E
2JIkmgRS6WAdTaK0veRQs5NGEkfnmd1uKntwnPJ1Qnubp6EJFNZGduAW1VNeGvFvi5SWt7SQwzG9
dSCuWR0DEAtae4F0xi5ZyOAfUoOa9RFYJC+epGecGxKfR7jJoe1MuwrkpGEFrZ5rgZ+nyeck5mQ6
mo7UcXz16hKigk8BE83kG4s/l4NkkUHq0xch0UdEyzXOe4Kdpa6bgL5j3MD8FE/qfGxXukn6eIZ3
wg4nXHjAlCNte+j/w10dQMFqtKwlkDouFeEO0dse/5HsU1GFRvA8WE2TjN2Ay6UVmalyzLS3Ifxy
5RqhrMVdYj0AXF8itLg1u51zYW4razbUwfM2KMUHNtEfFx7mGmnwH/4scP4BpEKfhTR1O1ysP0Ry
M13AU4q02HvMn5Xg/D2Mgpks4X3Ztn16W17QcmbMqugIKtC6XBxwPnRufY4d6R8jU7FVsqpHlsiD
0XA+aXM+6ecv/ifmpTId0dWw8haPM8EfvciKat7QhUwM8dFm6ggtB3FzJpQr+rscT7V+1d8B9NK5
Terqx40shkZ41JkevtepUGHLyWwoBi8PUBT289FKYNOYZdfIEJVrT00S9HoqOmsBQQSN58wPEKKB
EG5R1b5AXKQtOe2IBVIkwyr6EDwFYHki8/Og9euHqDDT420V/u4TsB7oiusMNvegf8p8ibwUexRo
W/1ggf1GO4+eIpQDNxvwpoMQIC1LhH3hZ/soJNr2zQ3nn9StaAhaJ8kbw/YYhpjTnKTpCHkp5DCu
bdHqqMMakcPcFCPqhHNEHEON2AMvn8W800aBDaQtHkVKXNEkbvISDf8fAOLEf48fBfr1c5AsKWXv
9LSLwTih2gMbjoLl5iGAbpJBbjg1iwXyCf+5mJIqBSf0VoOR3A63bi62nFvBrbv8XhjiUTjKhX0/
xDKHuCYZHhbaJvkr1wQSvUzk5V+8vaO1gcp463vFJ5YGtpG6gZAagLfQm/xD2eQxWFEYwJbwlXb5
TytUAp1xpt8MKUppuJAdAB31UstKsMCfM5wHB0wm62wh+H0w+Mxzu/nbYOh2NoB0YljoVPZyc/Nb
bM7FfM+akTZ+waYIUw6es1nU50gkGl1rT6nQ+TIjsg7nxiX6zngZBXcjcHMUG7aNkX8mULd/FMfo
WMdG2TtXiUuSIsc6DgTjKUU1VvOeoP+LPz5WglesiCwC/uFGJoXAYoKz+dZyGm2Rd5lepnSy6NGh
BrCJZ+nbIwegFIu9APFTfatKtOF0ak7Z8PrIYDph5vkjJm/WGHQkSOu5YJTnwtkdrAshbmzaqulr
+IC9o3Nm0EGHJfem4mJ8pdSCwHAHR2L1DDjp1r6gFE+NNJjhE8JjCe1eMRLNiPYJ+KIFd007fb3H
BebUa1vLpnJ7EJZ7hBsxv6VXJs/yrym8jt8bj0lKbq5ur/p8tNioIRfWMeNRpv1dftC9jYfH7F9B
uUXCPvCdk23R8uTS09UEoLnmrNDUSrcHIUTAkahirwv0yXL1oPOhUsz8fjeFKkeyY9hSfZQGIdfl
nTLTuKgSqWX/Sg30Ja0gFjCULE+19uNpIbF2bTAGGvhZkPmN9wheS/MJOYHAn3d/6C7gO7ma5LPq
pjG3CT5j29XhAZbTU1VHKTfcCEBo9ouMxneUBDI+I1KFMWqYq68cM3elKHDcYRZA+83UmPOxOKVn
5wfLjHstFu6QqAoaS7JzF6KmxNVdjA2DfFkvByNWfK78WMeAnnXrskWO3Fv7TWw9H9oMajlKBYFw
HoaPo58n1Awnf96IamtXrS+8zWXXuqv9OAXiTI43iRi0/yCEugCuT/HDcJ7YYj0ka7hQFcTj/5Bg
pt6Ic4vh7WVA1SfEmsp24yNtRPl3UJmH38tabktI2Vj+9vxjw0Z26YtAu2mzfYswb0SOriRfLdt/
4ICA/FXtltS2HHETnGpvX3eLyFa/Vp9n2TaEYpG9d0RzfOwxWoGTFitAWpoI5sa/ftyblRYQcySn
Tgoaf7azILr9SER3Yo2Egyny+vpMFk0jBugslUwaDurSvRHegzlLeRHJt/BKdAEzCPQAmX9suy9w
Amza+DWNQCnwfwnyXVFf6Vy6DP2dfKfkiMKirG9uQyoWXcaYnExsXtaJCDYWk11sVrIhvmEsceSU
ahcwyxV2CvhjvCpmVu8T4ag3n2Exrbw/Fs2ojAOCcI5Xycc6/D+F0WXs0gnWibOXEteiey14et5r
6cZOI2szhvsXfemZov2/vOT01Y78U8MTLY8ZHnef2dh70N8dKL/6Qj4pMu5tCEqMPK5JwBeeknTj
q3WRxddUr3ckcSaOBnB3ctaAkACmSiosXnOxejZ+6BhZVlYxkzjPZq9qaxsbqTfhj69QBvbDNO/Z
zOeEhKTC2eOBY5yHr5Kv3MM8kWNSmMnemDRzHp1DETJIgRKkFTB+nhNGRlD+6wvOzpwQ/v8FyVRL
GMrLPPCjbzdCw36tLdv6QBAXgjDNQ1mMcwRLqsRUZRsXSuXpUY5o0gCfvjQoxVGT2JaeliQnGYUF
hqnUF0M2EiqisH+d3CDIp4oaRP7yTijBLjBlqLsPXEARcSON/lWw4VM4qiaH6cXW678y6LVY2ckG
NJpy9PP9tY8diKnBiiV0jkKB06aGIptFt5UjG2vVb5jNl0+gkdPK6KOG9RO0AofNMrsYsLKrrqz0
gsKSeusvq/ntI0+AAMq30ajxzhgKjKjlIos+IFn1cp9zpzTAGOZ6YIy5oK6tpaUPpCzeMnXrwbWy
FcCgq3WGX3fDYfrkS0IvJaNHoeFghcL/kGqDqCSk5E5UTXOrTtkpuSJi+TWKxggsp9NTvJ+ps39j
9mE5XMy6dRKOOqdhe9ep/c44FMfPLnInXWC1YapXvERnKKVph4O+J713nhWk0lOWsQfARqkt3OmA
CIIWs9m0lYO9PJQEBaa0cUccvm3b6tnm54Dn7TiFj9ltdGaGpQHJ/OIGma8vxoaTIwkv77IFcMe6
dH6O9JXkvF7UOyo7Xe2bQabuW4fppBhMQxtFVdzaMsaRl2tYDx8YzOv6NJUfmjhl93mmxZgxlf/v
ChZ9YMrExnxsrt9YuM3kTxA/kawv30ObaXLnd00g2Y1SnDRkPb32Q9Qw22pze2YXbOXRvhMPPxsA
F8Dao5smQQ1RB6DluJae4157L2xWrHfuxcMfsVmVhtTIfYraOCFEzTqN5j1XLQWz66ucCo6UWWdD
F+qwfQwAhGJgMuoPUvY9AHbgtT49CMSurly/ELk33L9hFVQd8KjfOZDmTFaGsgIa8SQOhdhp1IqA
pffukJwclDqAI+bkVmlihj0KvHDBuNvJbRLHs2NwbIcj+rrlh1ryTNjnuzMEZJixMv9wmNGTansf
wq+Bg0r5J+6GaSlhoCn6qqCtbLcUb+7opLmUIjgJgJ1GpV/k5cNCeBoRLjk56mJhCuvKLtsZHDtC
TdRIcZ1iOb4juyH5xZG4ISsDm18WwkuzLU5D882aUjNBC3MFkOs7n7O9qjMdNuwHpwwpQbZFYrCl
3VWo0KQwHqQu5Q1Dk8hpzLv9WNO+kohCJIgbHv5TAnSXmRrpkXKeO1RSDhq9h2LqNL3re0Y3bGV0
mCSZ0jx0eiUby3Xa7vFsldgubGZ0Lbp3ACHfdJU64ionWgzy5SgM6WRQbsVPTFGa9NfmSG7Ibh9V
lhTTiRRa1cIkjXGBHNU8QSVuzSLSyq06TObd5/A87kKYcuFWnWZuxl0i7n1BUdaxCZ1JpYDWqxC0
zJ+5GtXoYA4pIvdd7B3yGQjyKj4Io5UQpBii6H6FeeH7mE2iS1B1wW/KSUKOTFgv7Z1u/5xlawdr
bK1r/rqbACV91ouMRGqO4zCFa/2E+LtA7acdWvXMm4XeXjQTotswNAjwvZL89ZHWDY2oklI5RirR
WmO7B+gsswCtlOu8HRGSYjvCHN17Oqi+YWbec3ABim5Ft8bEAz/1KcYOZs/1D9MczI+FUld7xKfs
2VBgJ2nUJuOgeHvj1/1ywLMxa3/DqpOa1EQJEnBPWWUS0csQ2lYVjvpMutSLRWYm9j7dowXznlUh
PL6Y/gnwpRpftcx8CFC8z8/JHOGkIEAak1U5t9jXLQCcQYHo+wY2O8U2Mt6EEcf3GFe20g4heGVE
2hGyvv3DigjLjNwtU+vYOW/t2EIlK4sIuqyNXnVrEIZYhY1sVcilqVU73zvUYd4QBts5fqK22qnv
ENJka4RnOhTPUBQ87MH9T7mgXNwkTPIJk1j6gHc+Hw7nyqzuuzoZ83Fp9BKcR3vSEQgTEa8/+9Y9
GXbQEQCHvxv5bdeslL70U00hquP/I7PAzSaxW5810qKRokphy783HGfM1DIlEvLJIbtoqjd1fJ6Q
+XwCgvOSvweK0afamvBr3XSgqLFmyEqKfHKU05OW97aiUGByKMakGd9V0icL5LdW+/OVVQs+Bx2K
/wGRR220gj7lvCRE7ztj4QbPxghziUWtFPc3uXwRJlPQSJbnmmFWVUGV8nCIY3e49pX0JukFIUk0
BDmcX8fgs7yNLjloHSiKkklkwmnGXQqDRwyPLR8bAICJlzcIO2UDgbNGRW6EvIB6tO6aW4clpZDJ
DjIwYUfRN4y0+3I+ZYvKNAVoTM9MjTxAwPYVbSQSA3vnXcHlry2ZIcFYBg+B37cOc7CZ/ju3wpdn
8uTj0hUPBsuIpGly5a6tiNdq148sNWyxErWIePjyeW+CyiEDSywZqEzE9lIVaL0qDCKi+Jq80LiD
S4+VHndCkxvgjMII2xIn5I53/WsuAwsHuautwar0ivfsSjXK3l+DSG97HKogrJmSxN4xmDPRO0r1
NxsqOydm3+EEAOqqYHZ0WAmxFN8Vq07hlJ8c+BxeEf6nwOuX9vX7McIxY6/ZJiowsGO1FL083hRe
VxGHujyuZz/uqg32mXhTSopmRXfGfBkLGra2YnyRICQBppV1f6E9t8VtCwLrbeCDWJCSXLYby93B
IoJd0gH4ltWvTD00ra4AMGBxhmYciqy7LGe2MpdKXLn3p4juLSee8hlsa+xW0ajKTQqiNojWX1oA
jXLAa8O1MQcuJ4RFWg+lqTj7idv5DxN5KHKb6yCzBym4mRfZQqPwv7+83+bhEA9xMyc6TAo8LbdO
iNjDWQCQifMD+1SmYwKx+bPrPM52geWLG1g2/AmVI7WdO0LohQdofCRRm5bvZhf5IZDgOyMT1wzX
p9nKbt/mLywD/u7tE9J9L/U7VNnO7E7VhfeT/XRgG8XzDQf3cfbp8jBXeX+mpf4+FQUrJ3Fvais1
0njuRtVAkIx8hqI5lOn2GmuybNyu+If5rOWZBWhnjmEhfmvUhlzoajMWaBn7PxnXKlscueQqpN5q
wJm7EIAomhzAz8qjcpYqUqfClmWi03bWHK6BEIp9zc6SEiYrkgdf7nPooUHR6p9QrW7QgbGbzrgv
MRwdb6QJ4j49X42Ofnr7iHQ7QWo4SmxQYNFX4uYBe/qEMDIwzY3j6GQ+QC9RydPYtBTtYXjxVsBM
t6m1tywq1frSb0a/yyCm3lwUYJpNhUgwUcYrDXv0LEM3Fj/u25p4ji8ILvlGv43CK2pZ3C/M7F8N
xrHxFyUnDwWmN1GWBh7tMqTpHeFI+bQXwVz0husxXfLM7kmh4VRnCU4mezl7moQs34G5TLQ/Kj7b
4JnTgIvh3N/RpAiIZlbROO2sk8CbNVFvxivaTuiWyB8lGzxFKu52aAVpdSmrCwMan4jpYK6zletl
SaNTpa+ZSy6/MXBv+aMorQYPXdN9kpEYlIH30e8+Y3lJeMghzexlQL3GrZhZs1mpkYfEVOXrdYSz
O2vH9Vqou8cS222+3tG3bwFlesDb61bNbZqmOA8p92kItEIVi7lEQt5VNezCMvQ8yw3BV09layJV
N3VIGXKdQH1ItxWbDknAVwAAZZgMDtK6CYL57TrGsFwH+7IEix5wGyPwL+vkqZiUoKRwBP1qgQsZ
pOlp4Ih+DqeypkCPDQao9u/MbOTVOUvL2xGa1V/VbMLCPFW0YoLwd6S57R+XUZx2bgrywNOyAgdJ
gsIDed5Qse/+OKB8rwuEBsa9Car6yoz1/3zJZWsc0CzW6v/WRF+RhIsaWslgAvjiWdZbYqzOtWSn
sNkiXsxFR/fZIirQLXdsFFi1n/FRLXMD7Q8kkKxPl1BmWw/O6rZXsKJmblM1eQghQ7pFxpAdMWoV
G31CMEYSFMmQr0LB57LqPuuBc7crZYtTBzlbtmZAlo9tSU/ZfiwoP3REEkGdwSTlzgT5YuUPJvOH
7GLUIrNMTeOJ4k8bC9q0yYj0spHkE/Gr4L91oQTTVJnpQKXyddsoTSF8C1M8CyZA/dOg5fglJuRX
153PQXWs5hMuiOLHZudlRnA91VD/zhTj/2bkppLCwzpFaZbYge8kXgurz1AzEuuf8KHqCNl7jCzQ
wAWmcfmTZMkK9SkOUIDbS/PB872i6DXSs41mxOeoa+TpyWMSbFXQMyRaCjVsfcMMzBblgHKFUMxg
6aj/3kEbDqxBaL72+2Jviy51tGFbrig1oavqndw3tUc9Cn4sQUf9M0IXqnkb1JjpN7onnuIw26d2
Y0uMi1l072HFHAPVXEMxhxxtf34ZMjZJsDWsAAq4OS822hkR3ZT53jn7uKtL3idc7oRo9GovY/rg
qBE5xz2XLLaTIOaQMUmrS5bnz3tCbzaXCImcQT4OXRoh5KbSM0H2hxO5BY3F38cp5xk0XyGT5gZS
JVg/vNTyRTyEC5+BRt85TRZMD7zcbB5HwsmjyinKvAlCzF3OWQ7aJ1gxJoOMH/XO4juBdTZvEYEF
jPlOSF5X2lwpc9RfDQGplptHI3xSYFUsuExEUiJF299JGlPapdnhJRNY22oet0jDwSs7+C+4dtMa
4XIemJ1LmnAOkWGJQiHd7SPMSYIJwrDDO80nD2pJTQQFpupYZ0zFJo4AWGJhstGBzXKvN0jVpQ6r
1S1kZNuEEasNfIGKzRMBVajc9+NQVULtKm+nGWH32T1zgLf12xolagmdgd89nUxEGHyLFQs9xYOa
Sm5DXOyXirwAwcLtgzBnHpev1/1VFAx0/tDZZdmhUzjmhBDD6zBonMt2cAcFuG0P5Qlz3hLqOi93
5o4/pf7utRb7mhx+CDI8NksycsnpTrwFYxcgmVtqJfa3uSwDn+4xsYN7d9/uwCZqwrhbVFb3h4uG
et32GCyKjEQOUAZFkZLZNODE6SwqMTukYJ5lZAczFN/z0QHLrxpPhrW8W8A249Gh8mSysAwfG5i8
OvOQrxM7gBqjtNrkziL4oCvrZBfPNo3wxC4BPA1Fnsq3nzv2wAdH5DVj+/YEoLve8cObFwL7Uecs
gdYWWPS68SCN/MwTuGVng8LikDaMHbfwdtO9LZJOcmYeAX+ioQAsAnypFv0zeCmdhBB9mpvMf2RW
1khj7E45g4nZyhYa9RBfSerO/hFy34zOZ+xkUHqZRhYwtszezWOzevwNATx5B4IN5Zd5wbu+Vog1
55rDXYjS1hBB9Ylj3JQUPw15IQyFF3wNgSlctBaszhR/J688RTV8dBdgNsY/huTWwEAHm8dlE+hE
D5T//kKXxOoeOS6sxwiEFGSwJyYgbyo0OV5R5eTxBR7S89FJVTw25RAJ6+juOmp838m6ecg5X3uo
lJ7M9ChW6QKLI12FiSVZ2vfmnVyH538VNn3MMvCxYxu7caVrwtRfIb8kumMJe3E6y1zRG8RhYl8u
z6qYycM5VrAv3egI9eYkq4ZgK5BiGJ0LFSiAza2KYOYXjZPS1At788HGuLIoet8812nNxMtfxqM7
SrFj6rdymiftmV7V1O5nTWShbzUImEqTMKbpr7sS925aVvDlFzsX/EM8E/WFwWOaVwKI7bsfxktA
223yqBkVx9X6B7D0Klg+x46ZWYmKoQEfc9ZSR1KSqug/Zo7PtXMepxTzHQKuLOjLflz1zINIAbQO
9F+1x3ZjrkNTRUE09FPGw41jwY6rYpY+MLZANAAvlT4sVME6zDzecP8r1hSZ/cHoHrzffvtJXibl
szU0bUjFW3tF4wREC30fbTXYTHc/V7QF5nCI6ghz+S3Wan4VKdzEQJiek1TBZqaFjBYqVgVeemvz
i72f0Qno5G3N0ZzMQSaccXFNSjk6Max9OzlRjr8UbK1+hJKXFOVFRzv4rWGQx9DP+U+cJH0Hti4q
9cFDdtqF7GymFEkIxiAZDcTbqE8aoI4wRAv76TQIvK3PdgUDIVoOZGdWvDp1qhvTG98/B+YOuF3I
4kK2DUwakEpS5rvZTtKbL4JdYfiA822eCarMts8uuY7Q/N9G8tnIyAVsshoEkeiUCN5PzIawV8gn
9eIeZ1zrGkzdj7KB2SGiBgKb+Vl/MUHqSUgb2CSMXjV8/B9Fh6ZWn24ArHHZ8aQGoa2raO1+aGxG
fdC7LhyM7JhTT4UoZYdCEXgzDzcZ2PqeGHDsLKt9DGjwj7xw2OswxDXcSicTXC7SB+6gNTBtyeoE
SfWeQQsRk42RkJij3wcp00zv1uEuucbjwr/ahoKA5KJNvqAYl68tX1foK/63n++VSd8misiE6mCB
JMHzrg1xVTolMAFZKRbutvBtfk03FUZCqexQ8vN4udnZlcGbMG1zwxkmBe13tT4pgLs4pkWDbd9V
IgfJ0XlrZNkkv3yWafneo2TfeOXbFaRC2I80FIMTuWovh0vqm419isAnAFZeLIHcB4J9RygQd4Y6
5u7REgjQit6cycYfMqh3bC2C5UZcXI2lP2XdrCqxnnV44EXnlZua4ZdbJvOSHjjS8f/oF60tsLmX
kjWqy3fpOE7Lx0f2kpjJKLUMG3zX59EG1X3HLp1nS7R+Oz8cy334zaVH6s/AkywYGMvOYTN9p2Sr
pMdaqQsxEdhOOWzFoRJZKiLj1jgFdDFJClznELZXepyvnYd2TA0/Ya1rM3Q3vRq5iX/jHPcandfK
PPPTAlvYU8ECr8OPY3lFPqH10R/YpDlP7B5BIW0vqVWw5YYJckBh7v6Rk7w5VKoIt0P59wTir8dh
4M7gS06/q4yB+d6uVegiMo1MGJgrm3s47dO11OeI+5Z/29U5yqUr6HrdEmyzGw93P8voaEtmQ1KZ
LArqHm+lcBjp9Kq9lrFTiScIT8+9Exx4q9azqWRsPp9CacsR5TUw0OoyPBiBLEWLB7Vj6a0sORQy
ci+nhUJPJT9fezZmvVu8eu5L0rVa/g2vZEKTX9BrerAityl/y5abU575vzWRIBdGBT6SS0f7edQL
iyNeUrumi1Db4RYBIlYXaTZHhgcU1FyiubFUlHTxKJReKi4xy/NeSw4prjpbeE+3WV8hcFt2H6XN
7N5qBA0jSBi+mCa3A/57wZNLhEr5YoaLeGsVxqVLlj21NOny2NF9NhexyVlJYbz/4VmwTGK/fYUj
t3aeevofT3MPNibSiXJWOZb4W1kgwG9fMttZkVB2iUT60rYAveikx7/RO3nLwiE4r6E+9JKvVunL
4eomoqrgwl5Ay8kY4B9VgQ8ZIj7JRew1jZAG8iQYgyRMVIj/VDqU5RtILC62F7fzCNQbS52BM2Zf
1kCEvlKPpz6g6mC++l/cvo/xVeijwWM0ggbwydVtYV1xS0eBsv0o07v11m6rpgw8tivKJuI36AfR
wc18gS98L9voowEEl/Al0yuYG5LChE4RKl+MJc5GgiPJndmFAMN7Jb5DYUWIkoXJwyicqckLqIUJ
DxxwAbt5rmaEDz3cH74sUVODzdGajJgrEetFRVRN2dJkYxwx3azWFTAinmONq2Vxw2eJv34Ja+S9
pyy8wtReUwrGEuPN8c4dSCqqXgSsLjE7c3wKJaNV7Oyhx3e1TXDOLcQUk2zvAJ19cr+7huvzgNq4
yUkFlrBJ1BNiQ+3m+d0+Hdhz/dA9KNsBaZhkEIQUzEE8n22D8PfiSAUmE9xrcbRcc6FrVTJZbOVR
mSEJbCJPGWTZL5pxa2v1RX9wkYG0wLLIYn63Xi9dSY5nfYmYDqgv6V6GY/lFvhkgXQ20xypxZL9k
h3soVAjwQP9GmEcTUSlInfWHAdKUy+ya+YdAnSkwqtkvFhcaKG9cag81O9k/570B4gFJ1QcmEYxY
0YYjKA3tPlIxJYsxg1b+Ne8P7SkmnM2anC+byLG1eNr7oC6K1PdRNDV26ZQOO7AWZOX6JiZORkuR
QspH/y96DynntmTwYKn/CSOUSmnhEFpY1AKAECn8jBmoJTLvJTQx3dUoyxWrhPNG2WE/mc+qTD2S
Uox7ri+3tidYA2Hcn8/G3jWxG4isFijRkcXrnLyY0Ag9GmwtjD13nB15wbvFKwz/x/9vJO+BcoIj
/babdn9KuUnxs/86XhqDJ3qOCGjpUigO4ymqXZzKk/oeUmBsA/vGM9tn//Q7PpWutnhSWiNM7RBs
MNjQYFFGhTca0xqyPozZS8KT8+nP+phMkLFX8OkKhlt6bU3hBYZzWcALTrsU7xE9H+XqavXShnuP
zejiqWXPEgVAxVsZhbJ5A82QzZpRqbMIa3R2di8sFPkp6qWIkivqTLFZJFqFT3Gg/h803u0/T/cZ
Ux5JkaxEiu2d0uh73/Llyvc4wcU3nQfzkybsQRMTJc1PicBXWr+53ZMBkXm7KAD8O/7IuzBAIy7A
864is/4kZjUn79ra4tpzSO1YvtmAjZo0+9VfhMmm7XjR5VqMLCRHZC37AddfT1nBngt8s4a1HTxN
LfcZJlPl1jOWLAznKrIruIqFDgTk0stx7g1Qb/3bOcvZIDw4hZkL/QImuUF/0hRLCXU7+J+60y7B
hQ3ndhQG4gg3/yZIp1V7/x8GtNoVtEnBWY60ZWFO0YwlsduCtRGKHDGOYSOxXQ/jxpJaeA8YB1Sn
cdMdkOmwPfOo8ZSCJqTXWcrV7L3OGdo7TV76rnCTgMFSohpNfJIxMkMvx/2KE2l5chNtnFCcwYYi
IRiCYE5+8Hv+F+mQCpjHqCMFR+TlF3gkrodmVHGAHJPwH7WbUw5dRmqeG9M+IrC+kbl2I4Yg21+I
OSkpr6MvtZMIpFmDLO8S2Yci3q/RkCRI8elJfnm/aPhezHtQazVIFLxyGiR9rKerjpBCfxJUEWk/
ahUiGl9psOjDGSNBMhwoYDosivF+AM2BYbuyqhHEbW0w6wvHpdI0Pax2hy2ZyM5h19UyCiFpgJ3w
o6GaRKz592rCsnovshALC74oDqMQ7s9S7iJv3AG3dQDljEKKVJR++vgKAOHLRDZm5Ubk2FVK5iDZ
jSwAbbdod+04G05sqRdv32FqRvXjQju2OiX4J0yxwsuZedrpAGnNu1yKY+q6nCoZiCf6ZqlwP0i8
9WxApRk9VEu/d5lMMSrRE6EbpaVQsYWxetvUVxNcBih/o2LHL696TnHsOZh/kGrYtwjo5nHDFi4M
SZyvFDLMafnxEi/XI4TeXVDw3hzRnbx838Cxq4j5n2Z3HJ0gPWy/cKgYPtQ5VxD+nwRtblNprTnt
7R5t814WDbuLrmHeJ8rX8Q/ANaxHfLZBStquMssiPd0X/wfW7CiJr10O71FUZFlMWQPm9qo5+hmC
AL8hpix1WkZzg3R+uw+kfx7jCLe8rYWJnbLsdy8W9pRn80B8qI9EVKdX+XZevm9SmC/gfCx23HIm
ipzUT98glGoue4fOrYoQibX1vYbdjQsR5Fm+GBZYzOukH/A/BlJMA9w0EXQbYhYKnTlmc2pBR8gN
L37trypuWT/KlabSFu2wmRCbupCiaihhnBkonumPzBdZwpNrcd4YkG0KS6GAIxmmRrCdQ8rveLLf
kAxaSjTcjFtAEIhQ2tiD64dU8AOZZFxkjU3nBouYmYHBLxp/5JXDPdr1SJf8RHAubu+HDi9SvkLB
cxJYrnod7H4Vl83DwVCl9rySc1KZcus4ciH5og3WJymFKI6SCdUOy4z11eWWrv4uX1/r9Rr2fhtc
iZjfsl73PNAc0tSCWbT33aIE47yNt/QZKgvhivp4xORb8EoxuPcH+COzHn6RSIQZWPBZn1TgnpB8
+XD+d4PizjnpaJkguuH9k/lRFw3FGFOEhjQDyEn9D18AuIoHLJ3BKoyJ466F5/NUVQ60T5Okn0iH
yBP3Ge4Bk5Reoh1I8CJbgSPZTLggcVbpDD+LieZmPue+XVpJNPTwS43kx71NH+AvxXNsRStZt5C1
hnLsUTIKSyw0PtKq3Jb8vXr6umtrkNUgftvuzJ3z3fx7oOZqHXIv43kM9DMad3hMc3whAPAIBpv7
P/GTLqaV+sFRoYD0XC5ODQV1aOMxr4f3FAOiq0f9AUx+mI+Cl9ePMVG56STW6+f+ipZTvoXNchk/
ey/3V20LNzWihtdlmp/57m8d2XwfphbFFrJIsC+luyfLs5qqt/Je6Jj2rlHXrgsYF0+Pw8KC7kmi
Vewgnm52lzum0CQ6C5gSTKzMIdOKy+1HDNTQZFqloQpdG+j2n1Qm9rnqKNGo4JrCSoAro9HAjy3I
hNZcBJZH7PuaV31IJgqLavK4C+cgNK3U6xIuVK+relntduR2CBd5GO7LqcL+bViRAj/mTt0FAiLU
zgEI4iFvyQnF85rHso5zrFGimYCXmHmynbHhuuJE7jhAC7o6B/Phr+FmZBPSUfOghfe5iA9EkeQq
rnnnjUs4gekcU00oBCJld5FAU4UOB8zd3asBolT6UQxC6TeBtq6QtH3e32RRIv7iS9GdVjhXdUYg
oX3u5bGZOIigvY5oJwTA7RQLfjVKBrgQUOOKUgUb+Ba+gWb5bpG3qXezONZAkfbG+WoR+e1r0Dyl
0DqGSpJ96hYyeBBinRlI4iim8+4bi9OpcyuVbGWBj2B0v+S7kJYqg3vd/awjl/xtxLV4xmTATa3z
HLrCeA3d2vPj4/lsgFPHwtOqODDPQYqcR2Hz2LQEea8OMFa8qzqxMXVeOA3qAYVCgsrToKH4r8o2
OmGuvF00SszjrAlzCAcEbu8cPnWmO3MDnPg+gaEZNvZW0kRX+NdE9c3wb976/F0GBL2kk9FZxoFt
O+7sRqyh9/NYqNPMVCBGc5bNpQDLIZShguzDctkY05C/uzTvFkXx6s/zvK7aKNIn+vUlOtx24xFu
I3e7uT9TLGNmkBb4Mq8XZFZlvtYtcjfFWWR0X8rkKmxHImG+eDxaJrWY8iZ6E0pLiXJKPsPYxWRH
0GsBuNLSGCYGwrQoehXs9TBtiJhtdw2QVfUWpOTjfS+hxOojBvLAYe43t+L+Xj2YlWkWPXCcPH90
Zw2y8Yn9v7vM4QfeQhKB+MDTQeg0BoKbgC+SWtUL6VyemVj1NCxpanV2c7J3xszGMfS5q8ACWqAA
NcIzqok5kXy3h110K+Qw//lZbjF3cpdDwGYGlO7nG1mnxCRoNBVkmlGN3DzS/wmEILuwoZxnOkVm
rnrcHQBh/orG94XGDhAnP2yazOXPcDsnslb8b9elojZtANIPR0HePR9ABWdSeFNZkNrqSVu2kz3o
G9JMxoIOnJeWqYIr7F2/+a1xKoJ0cVCdX4UUqBrx9UMUj8CEYyX8xZY9nj9L4OJ6MoM86UrDyZD0
2VNj2Mygb1aB1FawIsUIYQ4S4US1LELYWJbMKlR96H5ZwwJe9PaZ3j0jPsGAnEekxgibavEjKENR
nV8705YbfgfmnLBWg/uFEhv6OHdPq2lPDOkM1tX7/op5kfJ8Gk5udK/p7ybBMnbknUadiC9HFqNd
Zk7DeGnhC1dFertkx3QLnx2LD9rn6Hu+EDbxaAVTOLNHtCo4bjMbxKyp8ScHUbRgljKsGriLzaSz
C2A+ZMbt/xQGmWpxerJjPvdvFx8ZK0FYgQdDc5jyoPzwrt3RWhyMfmVUU5n7HIoWahgYVKpR5cFW
s6Fh+u53Lc2/Qk/Dozf+gMzmNTtC4taZ3tvvN9bq5KXv9Fc0zo/dtzaAp3npJGkK8BYMh8wbp2hr
9Z7PcbPdB+osV0WqDc0lE7N93GUrF62DtnEfNjpHPLsAyegcKu1jO5uklTlsJ0EZCKHRgBL/T5+K
terFX8yI8mXY6UFPmdTgyc+Fl1lXvLlEfUGQ8P2HdmudHlMMlbLnuq3vz4P20lwgf8mptWJPiF6Y
xC3U3mScBui8EWmnhehSWhJ6fo884c0plOeueaQaSarfCzFwv0Zdthg/rqWDG0JTJbT3CvO482ax
4qULSBMVN2hBi4XZjOtfQlW3MCLac8nLZ2oz3hA8n7H682T6pzV3yIMhMzt0Q+H2jLjs4uk7KvW5
jmfXF8IGc06zqyexJBQ/5NuSkv4xCVJWSb/ZQq5vTM5ggm73L45CJ7hRXKErn9n+V+myOi4EoqHk
hD1IwPq5FzLkIYGjXw764UuPOWtGKVsW9+dGtQgrt4kejRLgduic8otyDEyVyMrXmGKKxiQcdnCg
YFddKEG1T0+KMEe5MLIGs+TVpekFi92f58Ws4XP8wpPbeGKsUO0MPXEF+uBOvAyHeXYaweNRONww
vVUaHyttbe2FOXNjVh+724KnmLGcu2PbuxL0igESr1KJ96HYuXWbraVgmnQBqs2jIwab+IKZICZ8
VHjZMMcPWm3hEUtA5BB40+DSKuAmgmrOVIOjPZxNv1WIYhdiRXW2Ygp/5Po6YtZJp+uwGNPYNBPa
T7YpU9dMoA/5qpgljoYT0Bvohk8TDRDpGdugLiTOaNfEgTGl/QeeXekFvmnlk1BTlFH5W3Sc4GJe
i5W4DcxtHAdd16VRABr0+rmvbiIWNyfv55O1rV+dOpK8QkARHCU0enkXamZFR8N9uhCooNM0Q0+E
M5ZjGrBH8tjQvzMyV1jVFhFnYUgZ5yj3m67GaNBAkMnAIwyeYSs1evIiBPF4Wn23CuSfk8WIUPhX
LuoQbqwje8FdTm0bg2AMd73VbrsFo90i+/D1p/fw43TjzmqdPRC26pXIp78lVyZF66kJFkSNVWgi
+vGkEMPPIuujy/KwDKD4BmCJ8joHhFbUKYEsyKuZs22/P2OKvx0woJ3OqBlvYamPx/r0wNDCmCRo
GgArfBFBwP7ByUURQismi73gGvGP9fkjaTwEGpyvVDhucGNWb0dLJszZ4z7NP4pa8n55AtDnHXTn
pJODvWaNJf9OhAFshY6bvLn/4YPsvhIF7w6xYLRCesiUvvQIQw8AEbXBnSkGZ3aJTzX3B1UDfFXw
pcT/vIkQXi7tV8KuJ4/FiVGlpPPjF5ozKJbU4jq6Z8C6V544MIKbCMGFiEh/Uq8kgwpekGfVFXo7
VReCU8GYKXgqporX0RQJDKGmeKzWIgZcO8KBxRYjJRLCV2IgWV2abU5nUMwgQNM9zinh4rcM2r2Q
jw4X/YMO+W3lqlY16rgpx5sd+9u31N28ZpWGFDDD6XObAkuuDC40wb2qacngZaNQS26A849h2OBb
Ptawxk6gRoCnHRxQSeDShY3Fduc6DrliJvoAlosEcGGyDB/phn1JjkZCvQAQdlMz8f1lO9RvbSOV
vwP3LvF/TO5z/QKxnRiQD6RCCTGfx29N1h6EnDB4O9vvz4UKXAD7diIey/DZjbXQQT4RqA3G6uVE
mlvKFAPJE44xXFwmk0HxTjHJAMNRBHkoI0YrRVf/kaic8x5UgJH9MGUjvcY5GSXWBBEkNIF38XCY
l2/X7fjIfWOqG2yri4Al9RBsFHo0NHIqRh1U3r+tBG49OnuqrH5/AYtXRIeRGZ/LHKzseypOMMxL
A1iY4EJmkNvP3tijXpuAWGC6wSi68f4u+L2jRz/ZMJhURaiUOD6/WCMP6xNJE3qMOkuAeOjBJRIq
AqjdltsEucbmaBs1HjwDFWczTVkV0I/dYJeC95zNut4AgC0ZkqOK+47moPUK3eDnWJRoUDog9Bq/
OYhWHHDxTsp/71hnXdiNxnq7vEz3+ZVfP34P9Pav9jXPbLEUqJ1gwlD24Sr17EUcjpVEWRo7jwk4
MwHnFj8PRhCf6U5wKgIMDLGByzS3aPjKwv30hhx/qvFFcsF77AtFIoaJRqToDpxyfgKbh9psKyvH
oR3ZWnDs7oH1sTb0epzGZO0NZ4BtKo0JVybtmZZF1D8gSkQyUjFSFn2BTkOxaoE7MGmce+4aKHci
UsQvIoBkreVHhbzCJq9J2b1m+k6ss2O7rBNgtL+S7m48deolhBZMUkl4lmoWfM7bzDO4J9QoGA+H
pKzrVuBYMSqwJKeOtGKzzELw1JgxbzFPEfbEYNOppCagdfKZjr8YT3yr42SFbB22NZNdV04qY5SS
ehQOyIcJadWPkI8P+xT07hYPbiR/0JUlHOmBwP0xqVqvsRKiiTf5lwKtwPx8+y/ALVxtSzIVbn8U
9AmgqZTGWeWmBy92szgVC9cgDBW407XI1Sitbn9ySbIIuN/YLzET8dZ8p7P83Lpaf/LL3F8Le3gA
tiBpSUWp/+fEFFCIk90+I3lhXWLixJzGSU32cVUGg4a4xBg6hXiH3j4+eERmpoaud+bpST63z/+T
HKDKj+L67AlhT7UMDzQoJAczpUJ9Gukqn/z0JlVMTwWdM7WCekZJBYb29zx0vFTPtspJnFdMCH1e
QnR5sQNbIoluFAzWAmitw2dx4v8+QpXz/I33Do5Co6/QeZrd/9NYRALCcXT/TJ8dSSQBotD8QoCG
Fp6Dlb/MwCZgvs+I+45n378HrZIZYd3xsQ0VQqv7+UTgEMzXuJu7FzZ0R6wOFCWJnRSdH3uhOi8K
kFT9yShONflXoacfQvR76Pksi332UJ1s5VEGWibsCyEKcm5yDZZn9J5Qh8ejGxe69Dnoe/WKH4ba
NGv96Jh5SXyv/TjIXF0ups8K6L5ob06WD1rkXJeRQePhYQDlGrHKBTGzNQmDiBO9NqlwMHs4rfEW
9PVSFPggBn4W7mm8MfF0BdCuH4wagVLYwOIqjsJOAJL0CfOqd5Z7uxRQl0HUum1Jrj/4U0FN6vV5
v86eNnK7mO88A4pRbmhEBMttQMoWbzz3jr+AXf+9FE8BoBFKFRvRJKzBhX3XoxpyaEsL8BHXYWos
WZS0hYl1bPtoa0XCFC5NtYo97eZHQgyd0HvvsyPWolfa1DuaBcTOH1/poPjOXlAt2SdsI/qJe2Lq
prUh1QDeGC+QP1xrmnlrIdCLH9rXgxwoCMgvoGmHT1itfZ3VbE6akt0ot5kkUH3k1RiDTyaVWDll
HwzEvEmuhGHs3m2veTWIjRdiPVHhzmcwyWXcR0p24dNfYAO6MvzxjySq88d4WxGp4z5bA7T5QIZ8
DWh9jmWVjBiutOP5BbOcVdPcT7sfRkVhI2MW+LH6aXI5/4vCjb6qCiXF/LaBIKsWzCGyve6I8ff6
yRtc7asVlJaPSoya1de5LW9kOBH+bh7vzCdba43WL34km+7/7daNO5x2cg8BH6xR2htCvyBBlkgH
etRcRD7Vyp65pwW8GhZrVbwPelF3rKERcFwbPCx9Hyq3pbqhK6nMuNi3GOj382qnywcLbnzgxBuL
k2uipjyxk6YzketCmYJuqK23rpCQ/kzvVs8wXoJYJCHJoXsJVji6YQceu7q/xMpCkDh+ZpxmSIyb
TBYxL+xouRK+fXucQjVc25QKQU+nVV8ym5gRqq1GB0NpupRI4B/YslnaaHI1CdX7fCOCYZ8Ko76P
lFT51wFRi2oiZfDvyhtHLlrBmFrAV3fqqYoi9g9L/iV6NSbhX2WOis/f+A+YcZLTpkKzhVZqnXdq
VjHkAzY+9p8nsUowArYXbNLK93Si7LR/9DNgFUvdMJaW/6E7DFCCxbDCmuqDM57pRmMMU3D5mMQ0
veU5mpgeBx5O2cDVNAwlfMNMYMGeoXVuTPwH/BchJyxNkGCQNHcn/7PMSrBDyT1vABcWhNxRy0wh
5VppXIxrOYlAIrU8WnTM2Hz/iMWQVslFdlSo4UYl3PeV++4Sb/PwS+BYZ/9aoA7/kDheIbB7FXt/
tH0dyIxP043ggb5OCznkYp3OuySIznqxg8A1xIbx/VPaJHOC6eldtRujONeWKjlhc9lVRiTyesgI
ohBUg+bc+ydysb2FRe4WD2gix1gtfFH1QYSwWKlhSq9wVG0B7Dnt8Wmdov7KdiBwzPQnMWplIRIT
uVOKeVLgDJapi0YVMTsyUFmc1ZDiV+Jth/m05OJ+1WCOIXOHvb7Sfi+IO49xL445i5gU95xdw2Iw
0i/I4M8tw8cO6/XX5Ey4SzDtPHZfZ2k8xCuDUCV8wA252MHV70ZiUr9caIeXWvnxiSkrAQmAHLYU
kjfEV0GwHEWPNLzSAhNr96xZ4/gOn3BydAXBK2a79ywgynTGB40Cu6SPHTnmeWi3JgGbwjb3i1kv
ljBkPdT5zUjUC4D9FCT30AsY9SWMww7BER9DFRP6+2U7zRyvopSmQnB+PsTbaI9F8JAoJxBnukXh
INh7TGPNkMB5O+Jxz8e024jkZLkNGYqD9Nyv1IWVamlAFPtb6NnW8jmsiRX/hTeUUWcnKVSbOU7V
R3qVmhRpCTSIzt/L9XqETAYpCR5aCLOgW5NEm6BDE2rBAJQXbywfLBlgvJbM4WDP5BFdAOOs6JHk
wLH73uLasD2a2TCFmKL7cA+3xl4+6WfqOgbRLK7cGsDrvX9rXf7GPyj+JMsqCMWj2Ls2p2yb4uJd
tgGkU0JHpI2HztuK2YaTwxGoAGEIrn2drSUAUo+QHDeXXMRmUIAlfp4BCwzYdwlzm3W0d7tILy63
80oA0XKt1gPfuWf7pI+i9YU/KPe/msHhNqT9R1k3nmM3OxK5fAvms1okp+844UTh6LMLA0YmKhcW
ATb3yvSlvOG5c1/PYnhHKM0u7JQ3J9oMQP5RZe9aCKgpvNlXnD7bWZLeNlt7GQDHkeW4pgAD4wUS
j/XoZurXRwnFqN3+H9NCTpxJ1DGsyBbTYzo2Cwh4Ug4fQa8Ylkwar+ffDexAn92QjjcP/JMrLCVY
UktEdqMi2Az0NmMmIbHVP876wZnD/pZGsjFwx6riNH67S1awe1VcS99c13v71xoTqcCeFuT15p8w
F5cb7mR2bTRvytEmc1r67FPZCFOx3fzCf68tEuwA4XTeIttVgtl5cqE4WFl7XG5ATEebhzF6FQgV
W844BMsNCnfGSAp4tc46JQtU8khzAnJDYUx9nktCqyQdT/V6dPBPbUDC6CrjioKJZ5/7t15Log6J
WmL+q7O4jfcu36e7sbAWQvfnxOe+mY4scKCLn/57Jqi4w3KVOETU6Nvbb78xcyxdHlXcGaNZoaTw
2xr1PUMwZIpUR84Ncq8XqWo6q1jkCB7Y7tjnSltlIne/bkeE2zE30Mm9qi9SqAjir/L1ueRRYYYF
sgp9rDwZ4AaHKF4wbNR//NHR78sGoI9vBbRIzd/jPoxcxh5lYW/7uweaKlNY13pITxpT2f57oqc3
/KDRVYoMuj/Y0bxeWfPR0NBEKnzv+EoFfWVyOdldBcq+Yadqb7fOJlQt8z3Z1KgzhYUP8vbnSluR
GgZxD5cFLxn0va/9niiC5iJ2nc96bR+Xjj7AHMuYeWLk3RuSLvzGVxu79psA5OrbJ3G2EP/apkCX
C3RplH/lkWSFhXeXEOaGAQI6fhs7/9aVl1dFonEs+6sOFc875b34R8FyO3UfN7BsINW7r9XpyFY3
ipgm6wWJKt2sevQT8u4Ce7/ge816LT2VN9yDsljD2O9EXOcawumZSrkwOhdFj57QahY8HLLI++4f
o1DmJ7C8ALq/tzTEDUcuOLrYS1IIWIbkyAvznJ69MvemCSpaQBSEFDqPIYvWVgr4XofN5zD4MAuh
WuRR5zfAY+efw2A/fjy8UKl9zI63ASrgoWFUixtzeD+ssiZ20IScpQB+5ucs+ZqoSoe2W6AyPsV+
CZ94kFDj1rcWVmjxEv15XY6zQ0+TTb6dsguwsr/uiCeHLX1O3+6Aw+oqySipJkOo/NW0H9r2dsl8
IhzQkJfSWovXzUhFB8h/KIykK9d4sRgtKM7Nd7gFeH7MSxYjWW8bEP/KPLEe+x1fkEnDia/mn2LO
Pz+/y8vvudoBTEMpWbKZy5n7JR2Ooftu3yspOc1NdKo+Yyh1STZNuKNFgBaa4GyU3zFe0s1ObLOm
RAC7/ffqcHPuq3p6vgJQCFBG4tjlWg8en4SEw5e1lrCvvJubyHlEXnN8BNOsX2544LW+Wl43P+Yv
EPU9TbRRbFQRk5mau7VFoU1hV0ZRpCPMlSqvMw6z58t/Nwf1EQ3A/Lif/N2QOF5pN2w68E82uFHk
8215zSEBNoGGNACODyfww9t6oxpskrYtVWm8JSMYVFnnpuCpP59Hg3vE9+HKQfYBamZtKxNlgYY/
D3p7pnh8Jz712abkjkLwsaQoB/VmBobWLESyQIM0AKJEstD4fus4T1MBaIvjc25dbROeqPkicyYr
bo9KYpsyM8Tkfzjof3s5/lgHxjPumXOLI3sWBpWbJ90yS6IoD64mbBOhfZ4gzpHptrHiBmSm9krO
0kckPXyjVFiAkJnTA/EKIjpczr2seVRg/87kYNc5yj2vYv8Wf/9je3i0WuojSGBW9hSwTNRPFow7
TgjkIzhHUiaKAlzP/pEQ3Dy92Llv606m09Mo9l+Us5Y5hJ8F26SUm3vpFoXG2PYCbVHnd4Q2jdfx
9bWCoQeXifZ7CH8Wmrtxo6FibCjEkqNcVDAdCArKT7MIOGRcFYMLMCqkiux1fWYDji6AOv2dtddx
tHHn1D+lqyOHITqLJhdWKCsAwpgJ18oQhHyYgHexeou85rKDpelghk+FYDnGhyh0Dxw5fOXtkOm7
wXMjRoxvCv7Rqz6Z5HtMS5kt3pn9+/P1zBSd6WsL+5uS5oLm60udoFRcWu9XYZQAz7HrdKw+TeW3
uXzHi7dP4kfEreznxedz9JtOFzTlRora6DEaxYAF2x+eckr0R1HwNqRYw5rdMbLO6y7dkfLOL0/h
evpyGpXTmAsDfMqONaC4sWsb8/js5dDSP2GN1iSI8DqVs8ScIwF/OaMkom1OtN5NFihd1vJtfPvf
1napR3CRrykm09InOzx8Zopt0gANKYSgFxMNYZEVEkOshJisiS2SGkaad8xyzcj1AC9sCuXWLFfs
PMpvnm1rVT4nUwRg0eILCB8ckV5zZVdVnvppX8S9VAw0Mpn659zhzK88Z90gylK6nr4aMvZmdZEY
M+IYKEIY80/3b0P7/VfXzfw+/Efq/ZmWNsTBTMuCGTyYYTd5zeRPXnTIkrlb0XkCn309cYrWWLSq
du6TUhNo8iIORYPFcaolqVnB3zOYesvEWxiOjt0GcoGACnnTlm1TcELc+ch2P4C90VrSLp6+cEZK
zyy7j47a4jfzwiUnmWbEWGiLvATD4AINU/EKWpHmxg/zfHE+V2fNFtUlTRdKcDF+s3mltojj2gs2
3bk1cJhypfNN18nA0d1xZAZaLzal/laFXegtQp27TzdfwreKSgmKwmsM5wES612iApVOhlEPr7Mu
hS1Yph9l7YsPA6Eks5C1rrpG7wjC7nxLZbFBGUTjKe/vcnDsyyOW9rErUv5RpkMJvc0r3KsayLWi
a/M3ujoX2BI7wJ7iDu4fY3anBkxa/HbVXiTWQGOvKZNVbQsCtmk/7BesUbbw1C8M04Rs2+Y2+WUw
TxJLyg4wr8Iz/ZjhoJOA+TdTRE+BrBxC1ixJzzPh4mIDAjLmDGI9p3hrOeByct/ZQg5u3YOk1CxS
wlQrbXOAHH5OqhDvQU+Ts/g3V2qDxXhb/geOadwFOKMNySs2dLUhZkUkQvTsA7CUc1JazMgKZgMK
tir0FHZ7vg++Eq2XRlXCSFqdKmyE+E7VKredWxuk0KsEHvbxiJcIJ5vcbSpvYOdMG8MQtP9BZ4pb
2ZHk8mulo2WCr2tX3BBV+WVzE85lBAtgoXQGHvSuftcT6sAbQiTj4Z7PtvxUwmq/yNFpYg3u3lhi
EwZlxEcVCp+wHrdIijJmvBbVOwPfGdH+go4P1zoSuPl+0SmXQkxDLcQbTIxmkDGg4jqm02OKPalD
++V5zdElm+B2EvGLEEJXIxYG1691nggZyiq08VM3GKH9ig+dcpRFyHozN5mEEdIsmNyl7YMfvcWl
O5xQit7r87rP/viD6Ron+wf+OV91aE5USh5S106hie/Ezh+4IMoctJxuccfUR7q+ASez1KddkvOx
c1xXQroqTrcpOdSpEvx/aDit2Tm8tsxNskeQucIwqnK6U2PKHTGPn+MPRv6RFFWpIYAgtPQtWhwN
SfU1BRGUkang6jbL6/obq16skYGL6cIaikbx4zHogDe1S9aw+QbD4qtsLUCJLogoyhreO4P0oUyL
pADq7A4eAdjsC8tgkW7St+Tt+KFPBcOUS/8j6QSK9zwjV9caq9+ywhGICLDGORyCzhfyaXKLUYSS
B8vR9CPd3Nc8B+BVvlE+WBA3zu0rgmKoONKTJfOHf58RAioWOH2Qaz7sf3GTKvvWInlh/NG2/m3H
gxZnR1JEuGoa8FM7Esh0Bc5W7hpVM+HmTzCAe4Nv9bAiY1lzyMiS/Mp0aO78US1pWPO6bUUrO3tA
Ocu3wgKpKG5S8g0UHbz6pxSNdlJctVez91dGjjSJazwlpRRgP2/389ZWa7EAGMcRaVsKiw4S+XEo
wWKZ6rNatGx+Gpa0JZu4bI2yKzd/ZIiIlr2QWYR1zdrRunZpyhp92v4uRhuDLRWjtVGesnYEf8qx
fIMQQbSc4WdvBsqr68dC/qSday5P5iQPeMz9E0PVSrGizWnjmKYchuEQLLGmgI+wMjsA1g/5/GLt
tgK6YdrLaWYW80n0aWoJX9enmkVE88MiRrLnlVDPbArCrUEAet4jqZH9z839HqoHCJE5rXShL6SM
nw95CHYRZpAsM9J7d3pLhpDxXzrrQsvFiOZxmzz3oF1mczkFeHT8lJLJ7CEFxvqmKYUXygEwvPgC
MsqtOS4i9NK2fmKVZ5GF3U55U+SlH4kY/v/pipCiuniSN42m3plHafAYRISfInn3Yyls4/zQVwcN
C32xfY/D1EAVciL6PyWPC7i/U/bolKFMsis3XpSk3YMkgXdY9Vu3gmGXu8TTA3wUKJDAkUA5Og3o
QSggAOh/gyQAmF6gjJXoihF4YYr5udyromSPQ4gIuaoWsDfA/fObrb62FpgZSrYahM08ho7vCs7N
Ym7IKz24pDC9Zzzvm+VUQjyw7v0q5MTF7/VDKgT3RGzlWza99YQqAqDWS57dKBFjDIR/NmNPsTrl
j1mG4O1aCO4kWTUevfa1C7RhmahPH6S1MKKMoYnAVRyPhwkJdvx9lQNJCOr8CHj78JIdsZWWcY7U
zWyTUnH0klX7/fqTyIDNihuXMlPZLQxvCHUDDgGhdgIFibzqQExOhlzdvwyzpg25Ns+5F0ppQ6BN
7TQAklTUZh28LirXpYNWTJw4BWOslxiilzPz8+t8ahGhqIju/Lxp/woPGGY1hCRWMx1FrFtwZu5k
gLVI6AUz9jYNJ+EowxaRJmU06+EwMXjZ2r42vylhuDfs3rTEmf0h/Zu59G/TDPY5OoS5DgiF7gWr
PD2lkdUijRPgUxX01IMPI0Yx1gY6XubdR8EZDW6O9A3HVfVXCTTJndgi/mRFr4TiNxdNNIzGP4Js
QKZ2iMq4QrncXUBm1pxmnZ4hDvnau/i6eqQgKRt9C0UxHNXiJZvau5bAHbuL7YTqRpCosdn+dida
k1x5jOqZSK/s9bR8Ckaqc91DzCxyY5armkWVJDPgLbbYHhXopk1YqJA8OkD9TD2yCCnkiGnmfLoL
xxtZIBTiwmVHdcKX/OUYTAPg31iV0Okeyh1bQb/sKGOxKNcLIILE+W6yVSNLbhvOjPIbWzQ0/snt
zKCwXQd9o1aCWeB7gN6QuL4kel0psvm/q8SHtw5uGmyvOdaI+6gUpUcNOnRcgHiZIxny5c/67aVF
BveI9fubH4PBBFp4vCfhbTqp3yXPw/wAhOkLzTKnCuTInwLs/ly01idnmqQpxtHsptqJQsvVGyw6
/4Gp2Su4i7pNU4nSyfrT5RLzgMVXSFS73/5d04bcw4By7b3zGINd8jPUzY7rgyj9MFPb9094iv7s
AiRk8HUYZ6P/Z/8mcBkisvqdSyclOUmr/PDR25d1O5YETF0AMw69KByosdR7QuXw/vAN8ih3vBGM
R/e5W9KjPrbqw4Y2Iuc+Lc/IKUob+tBZ5n/N1YzkWPyAawbzPci8u/QfrYtUuD51j5oC/MNIc/fq
/AaU5vaOr10+334ma+jGmKOkG9j1oe7NFVdbulpjMZGSlxyTJULhpB6+pq9ogW5V1XPEYz4/DXBS
sB4OfjzdLWHBPeTB1jzFVPzHhL58RuYw9kaDplb42pFqfHJ/YhsGABEy4XWpCkW9LxR5umfOe4fU
W3KYb3E0Hjqr8OcsuLBcNYiT84I3ABLyEPL8Hoj/JkOprwRInqqc7HpjIPi7lwk9VDHVdXF5twak
VaHdugtWBWx1XIIaDnBK+lzFZ1PbwduHzL2fEGffeKp9DvGeBI465m0R/mWKUVHnpEWOOt0b3ujM
m1Vrs+RyxmV0mKSU5tdtDrwDs9o8cGu3dU5B0Dedws3NDyFAD4OV5GXNgbXAP8kV/cwXC8Mp4Ves
eBLfYDsVx1elefer3ytflqpSLjQek6Rtjj88YZ1oxaOWKBbxzzQXMGRvZSLNIrw6hkWZUUAqN9zk
pC8MQDuhZau2+S1SjAIRVzglDQTW5TFERLhLmx5qUx/aoNZCLsBVaEFhKLL0ypkSSppa9l0NAKH+
0bJnmzQbPL7jDriPaYVJbK+mVFt4CpIcF0y/ggPvlmGSNlToKjxkdPMyKXE/MHeRnDqWsYcb9ZDe
dPFv4flsdkw3JH+GpSx7xiqtITvG+28+trXL+8vRb1VDhemjAgrjDEKwLwG4cqaS7qt4Uaky7qos
yjB+1qTk6cPvtMNgjpoXvl1vPywdFBuqzHb4F48TL66rlDlf/CkhHFXFaUZeDtJxm18j5mfMeAoP
Z7TRphthMdpdYQH7Uk2hKNi3186+TYrBu0c33Tqy5R/cD+avA+DNv4neJY82466JQBnHQE2qsKYb
17uU72KPS79VhgVfo5+HSBeL8dCHCciwFjQNSwtpwa8Y88hpc6cCsx4MpWReuK/pchX1OyUFbyyR
KhyaZqnPlNaEoac1WUXxpAn3+jRau+Iu5b+PGnam6qR9N0KahEFCPLsJ08mn6l684c9lZKXppfDk
DSX8GA8uXPk0cINnPNgrGf7T6SKEk52rNj+fP6vbsuwAZ7ErgoLuLoZk1I0jhZRIeuFeiPjcfs7A
f+kCrNC6+9aVqEAzLih7buCL4O9ZY9R/TA+M6+b8uGfZwIT+EsZMKdQxEI6yP/TiaxelkpOZt3QA
7iahsHgAHpFVKiV+n3MpPV+WV98iah9NXfWSigKM7ulFsY560Y7cuz0fXcNzymKeIQqBJMZlSGXp
3TOztjwIkOsHNr6kAyse5gPYiDeMB5AdzuuZ8lg8mBVQh++PF4PwMyLAx9igaJyJlsXAM/rKqWOE
28WVcZIyOUqNY3TkVWKFBR0pzL0lgL8BwkB5VFl5C/NY9nltu/OlLm2hIz2vZSNCvDYAk9rjtvc+
flIF0nXM8G4q5KJv7RY0sFIv91sOZ909b1QtUplBre2aG8TSjQK1bxJBFnhuHuyS4h4YjuOCYv3Y
trywsy/58pqSgassRxmc+op2sY6YnMqaBCvBhx2InbkyMyIRFbRKiLQ5Z2K9pxJdQn0d62kkkDHg
+SbJHnQzG2j10wSzTaabmbXFHF4ex06eXaV8yZhgHs4+7i026xuEwSBAvM7g3VkBIv1lw5iQqVea
WOxfaGcvbJX86OBTduLBbxfn8wAjqz0PPoLdfIw03JNzH6odq6ALMdTBW4FN01xKsxw68uQGnC7f
5ZqjRsy838QPBUDNGn4JJi2se8sA/firhKO764W5tsDsWx+FWRTrP6/6RutfW3TqOEmqVjPhH3+D
bRRAZEmEe1pen7lmKuDoUMzh1IAs2Kf8Na3ZoJ0BocIMMDOyscDaFXfIrSx4lrdCueXo9GY7nRVU
5FaTPlkeQfdIyQK2MHQNLeCH6IF3Nibnl4nVczT6HCY17H6/F1bs63rAbiY9RbyxD9zVZeR9dXg7
PzdtkznLIfnIG68XS6dht6tGu0gRmhmlZZZ30OacT2irMmdybiBi5GYPGfNDbrKanaVXUqYkiUAN
UepVpNh7hfiVKPa7IEISoCBZ5ygQWXq8sYPhI0RlH7xn3eSnvQlsjVFj3LlKJE6hcDUygB1Ixnbo
wZBldz90JrP9e0sp84jKduE8JmTFHw+z51r+5w/k0RDcxwJKsIF86fLeV9sVeRHdE3cUdJu04I3H
a34wL/FbxvPPlW31V+dH6UyWxyqqrlWAwXN1HXI8rh51iAKmCpyE98yqOGjeV+ynobjPbTrlecPL
PeuMUbEuKuNJ9knP0oQQuOc2dpeaYBOfFoNSqD88WP3Nhxr81BMHpB5OYz1IK51tMgSLpf0VbABW
6L4Yo3D0SCynDKPEuNPludgXHOZiTilgaa9BLcmGxFQR7VvgQUMDypuARFepyBJNmfkJlbvbtlVE
G0JdwQFehC4L9BhDG44jRhdHpAhUo2m53U29uLec5M4l1kQ9XQD2uX7t9ohdmYsFF65E9fIc8i+2
C65vqvdB4W1CGw66kBqiThhclE/yUJG6BQ9Lds0oFfK2PXROdgv73zGSXX8fRVNgF//0DAYHkBHT
mFgK885Tjxwj9X9q3aqR1MiCnNJaVn9ra1XzgCucZyvktMHEBfOqsUawpmqT2deHL1bd6co1rvTc
tq/UAgqmd+VLEH2i/RO0NXj9nIgkHsLTylaxLbLXohC7D1W9nJXjaD5Ws9DceQ74/unjZUhRXW4b
WutzBwefFBEv4gGIgVFSey5N1Es1q05+BFq/o+lg+PpK66IiDBsx0HonnTJiNS/k7PA9ob7IeTR6
kkPJMAeO4Fp/4R/a+8ggUFzavJw+4svb6oOUWZdKX92OTdwZL7mMvT9U08HU5uRu9XMd3IFY/Okv
pFm56FpNowZS3xNoLz00NgtG1Gjw2LxCNkSDJbFerSlXDnN8zMYZAE6wIEveOy5gUULE4i/09s6Y
6VVBFxJm9pVZ9YD/JspBGhE3LFik2nijDZ1s56W/AQV3pmzOomKOk8iCx+lnP5/JO40SN8PvU6h/
pV/fzB6gOXWbFkJpnLH2FAjdvIwW2dAuCCrVWzjMdOAk+WgAaY25fa6VOZZ2QjaOxbmjEsdcacjX
uOAQCJOSMknolZXWQUcYqJKs1pEaLaJSlIKYwnoqyTxhxDSHb5Nn+1xbpoCb6VoQUTK1iYtP1G5p
IM+lqRvfG7947eVu0DcwjR3p7jmfSM75REYCm7yEDP+P17ajLpkN/GxJfVRd+SNnYajlt0TQUwRX
mM5maMNl+pxA1iGWWTi/tH7x1Idhb/q6aeB4HHU8oOsO/pIlxXait8Zz3i2vfFRf29EO5tQJGTQc
brkIkmUdj919Xi8FIiyt8nGTUQ/NT+AO6REgTVeyvZVDWP59zYL//GealxcP8Dyqi/KRFucTbAts
0PpaUDLDsJ/YtY7/css2fTMpXb2gwhC9TkIO/dCCowEw6dvgwCgu8ZTp7/40hIuN5rtx6iQivpJO
MzVim3VhU+mYbbu/baaDeQFYlq0Ng+F4C/t9ERrpRYVbIcjKSrwca/bDpiHtbgsJ7uWKu0tL0k1x
evy/kvmkZclSYF3MJUwGPOhlzniud2Y5/g8c6dSpMKBOQSDT6DwrssmlWkI7n61qov6S2jMExQts
+zeUohEEntE6m2pNBf5J8Hi4zmizuDPY+t3ElEAlNsrAi3MhTtyLQXSyO0MJVcwwTK6ibo2hJTCW
RYBWBmwz2OaXlF4oKjIO3KzP00/wYqYygZO2Q/Y8nDx4b2hGl3ZfdVlRynb6cNGblfFArAnBJ7K4
cR3rMMsb9JPB/GiQqwugBZ74ap8wvn375dvy8+QhWknxjmEG4ovZW0BAqQB8J93qGY95tJKjdQHK
vPVUAtjXMpmAdZccIE48VdpcWNrTz89yN2UQ+tceVIyxzY7YizICgdFai1ZI4QHaFyPjyxyrcy1M
W4R6pIW/tyNglazUbFlY8we2Xh3btKZlTBFUpgFZUHst04O+U8Ny8/8FSyppH/6ruDPUPK7ughNV
df2AiymqBmcFoR3Cm+6ZTvIhOCkiGpaVF8r/k2jbSP0tNksXePIt8eiKrZINBUgoSO6xY66vFOxc
VM12t0hwM5EppGi3k194YLREEJ+FxCZwNO/j3uIGUjcpKYo3NRBlr8n27isZTc/IG3i99befw72i
om0nwVccVWAe099m4W+eFtYDVGciaIoeaSmZtJ9NTupFyNlfbKOex+yYfLt3qMbVCmugkk0mSU4X
I0eKa2rygUOCCOOwydekQTBY+k781F+jxcLvDw4M+tJFjx4Q5Npw8RCXXkbMF90SGcGHJNVTF14L
4jnOSj5aQSN6xBTcKGvczhXe+RvMH1VTz1a/0QLGcXhrzTLSDGpeK0vp4GAow6oyN+C+Q4D96Ul1
drMFuuAUryYcXpbZRSwhEaNp5bo6zHWoPIdKvBOJ4XJypzsJ9QUKGcFjIeZ9K8KHt0UApgnMgR0s
Rj2srKR3ycVLA+cbAZSvAqbFQe9FNliGVREJOo3vNxcVXvVo41ZQnRWMR9WjNjEQc0RDo8AYQAPm
GcSFleTF9mSXNIPTvOwzsMse9dtpOc0u2WV6wYf5Q7yVLtO765gCj/SKuzU7qHx4QFrxfleluCo6
bZzjF5I7nth4MX+G02gws4pwC1xeCR09L3kIsrQh8aHkAsYhluLa9rv3O+uWLANA4OJWhFxQ+N8F
CZ3aLak/+LpAyPgjF/kkZZfMA2B2wF7JWT1VJxbryyI4bOxgfrr70Nnoaw/BlQrJEmMDhXLbvQ6p
ViQiWJFaEASOj0VYEJgFWUisUdJIdf0efwZAOrVepMZuNnbq7XA5wrUYeXNytszQp0Dc8iSJUjPf
Grbk6lqbqrdtOEVRU4RQ88+kL+Bn4CyHjABWEMopkKbRGTDAfO7NZhk5ffuT8oYmFlxBJy6eQn2b
xCP3YzhVyOD3y58jzlZvOER7O1ozN8IvO6cemRfH9m5Dl/hdWZVUeTiA9iAgeQO56X/B1poctcJI
E8bJqrKb3l+mTMt+Udn2AYYyhSU/t3MIs5uc/d51Jp2XjMjxqMmFer71ylL+1Sz7xYnEFdVcNmXq
zOgF4pJE8Z83dH6YWmjLFVO+9QjDCy2wgrd5BCvpByja6kXfYdM2Sc1EuFBFAtaLuVff2nEVOiaZ
njFAzbchXJvV386oRtRvE/U7uOd19HWXBHVWvV85MS8lqdCupPL6ZAv6b9+p6apu9ngni2EqsX9I
7YvhARj9Hw5A4Yf1MMSdyUaaSmFNvfVPVGbvIgCoU3EStfskt1vtzZX3yqCufvvwIuf4xunoH/q3
XUo9kJeW9IYpCjo2pAzTwKn9Sf75+1InvIuUAcBhuXXWSywouwTo3RfO9ETzHomz//YrMjzGkBbX
fQE93DE+3hsoHcd8BvrQw9Tt7H/LIvqBSGoE91pgSa4T26UqLHq+dYAlRj8o8rGw71Xh7ARc2mGo
M/JUMtT9WGrFnoXl0UNVoVsMBN9MExuXARtdvibp1ACT5XKw88eSJ/2DjgGXRl2FbxTmCHTOSoZ5
bBc7c896uYv4SAp0+R0foAPdpIXhOdOe+JKVe5OFRhh+8PvRp5UshHJuIptMsH8qcutkaNDjoitB
3jgICgyLmzhn/LuhrBE41E/7sWQ7RisyyNUQTWs7TlriODOQGRoG2AXpPwa+17owWpk90drpQg3w
5Q/1q3Dlopne8Q4EabzoQmRTjUOQeOck67k952bvNSsZ0E1KWb4MlOMTbMt4buCjjhut0KJarlLw
GFTRHohkQRHiJ7EKQkGX4HfGgK+a0z3ObbsMz62e/+5UoJ7GSKDoD/9jKnxxBcyWTQktNgmOAXfR
XA7odwYFtRIqOKqzNxfvDGv8JXGQj2czN+2tayeRwerhI1T35wHJPN3Ry943NWpzclSYYESVsv+L
OXMGTVjpDYcRFCUjIDurXA+CwGlWTVjW2Vf2OgWvScKPnvA26IfPhXBcnmN+BjvNVAh47tZyIuAX
usBPllKHOBpUnkviXij7vCaHKBn/mVlACZZsAloCNyAmqNgVUtaY7p6H0k0ULUoPx4cU4nOXRCdt
Ax+d5U8iwUYtmlTE6IupsmOg5NUuvL+hjWKnp/T9WJXjYq/jcdXgjuQVgywAPRIOKiZsdjktgE/F
o0Q0rUm1TCui1egeNzPSUAz9e0Umm2R202ofUsVmiQzaDWTxKtna31GlyGGAUCTwiw9rDD1zBr5y
mYY3RwEJbiTBXQnXCcRgGn6LxhH9RLuZpq5CYGb8n4V8OSECF62dnotiU8WwXCYpW4VLdm56qCpw
vAniueulVLqPRxB4gF1d/EE6Y6nrhMUndzY3jjzGQNHd+EqM6CgRQFScuNA2dLmVNHnstuZrIZrv
e82FVCUpLIDIDWiMs69zUoExNh/FnWpx5IMJuTifVB54UBvN4Ntax0CCJZZSe9HUetJQ905NLZrE
HNgkgpt4RDoxri1VKernx8IM52P9vWd+B3bS2NPiLM/t6YMbwwVUvN3pPsCZsi61H8kYOvjZg9xg
H0y5wu2hWDt2UPkIDxFS9hyDHAsnjcTosD3xc6bffMzUrwQgSWhkmOTvUecfk2WnrXwf/DUygd07
DS/yi9uEaGMPga3NOcbBB9g52cnnCuoEno6TApZWpeXd7g84suBfxDMaMkfBgLucDTTKbnJXExxL
x57JX/Bj8CJjcnkIOKmvQq7zS+s5SnDXXK4A05ZAotGYZVStpUXZSGvQVVrlHOIdfLlUhBk+w/Th
Krfzqy0O/zxALgYihToX88JlNBj6wvTuAyRxMMuXM4CohnCus4Rph3Ia8xZ5rWPTpXyE6dht8If7
ZugMnIsmSczjuqWLlb8ns9KL51JWx0hinQ9P4cAWLDeVSFjzRFGvCV0s8m6/mfWJOG+nb0dgn/EC
s0/paGij7mFKJ4hTPuhV5I4x3MCBM592DpMRLeiQGLZFzV1zgWZIR6JAxYNqySnIpYhPFJGTiWok
lLPZm5SHHLb1TpaE2JhLoplTemKwwMgKbgh1/K/eAF2qTS09xkRG4Zpm78ByS91bWUvKgXxmNaFU
ot/gfcSlneSIuUg+c+tLEErszJKauNGgBrS/oHtixVohuTZVzI+aodMqTDYl69uspibF04rovXZ0
0lQiBLz2mmCdSyz+hJRVLbKlG8NfUCuvDBOHeV41+aAxOyWhwy053tTfqpV+d/fQyEwWrJUgw/GH
ItM4CTkOSAxheNqK0yQeYec/GBwclG0i2u7t2V12/gW1H23LI+PHw880Qm2cVM7MJ/G8K122lbHE
0BacrutXtWA8DmuN3GqwpwWrvZ0kheNfwTsbY8Oa1bDaT823LeOPyTWI/qXKnu2bEWYfPeOC6OUQ
3sxW88mjMeqzZhlIfeyXCZdqjHaBNovigwepEvCov6RBbwIXe3Z010OA3MMEPDaXSsAwvOKlC/Si
DFhR/UusGveSD3q9gCnExqbf0CeiAOVY9qkoeMV5lfoFIf+9E0n3zgG/a/RJ9wvqMszW5i4Bv5j+
1VTYY783YQUrn/PKB7GuUHQINb1SykBubeP8/hXfiNsOf0/Hocw+0dPOkqLEoDB2TdRfvw2zh85c
8VTm9lVOkWqfDCvoqg+0gatk7gfZHwHPYAtaVTr/kSV/SLyDSJWm/JMFJgU88+zwlCkr2qtJl4kh
4iqmpsaM3w+9itfA3ManyDRjA+kKfD9gjWu8FfJI3Vo/z/nPQrrnp/uOTMq8H+M7w/L9PMFP5VrS
99SCP8htuglEjMJnuvOUV8aJfFa2Ho0czDQPshXsRMRg9CLrj99u0WtVx4et3gh7fjoGOWCDE3Zk
hDxQtyC1SvtodKU6XPK+PdrU1UctgtSyPP1nLGbA2iOq/M2qQj0Lmf9D9oljHwspiQLqosB803VS
v2NIK1oeQTCGMgUuJgOrwgS/QP/A8jzQMK6wMqhUXd+baJ0mcsB42koRPSDZihdNfs9Xe9hy898w
rBOA7eeBjf6XIQRVJ8af3JXtgBl74c9xMSvySxN9hJn5wWiq2lM3KwJKZfaQsjhPQ5UeMt417D9j
gTBEKQk1bB/8l8KBQCTxQj4gs9BD4lx2EjWYMWJDrXkfWId9f7xix4kDuSWXyCiHnR9zGM/hal5B
nS68G0Fg5g/TOpAUKJaUnPd0TcgC9dn6b5Fp+2O9f5DFszFpVn8h8Hbaq45VgmmwnrP3p48DgaOW
4UWObgxzOzkvV8hdUDxEh7av9qY83QPmQ90DJnmAy/KeCkN6lo323tl2uO64+RNCKGEZDTAslDC/
6+P/2nQLigTj6CAN3hKmF/DPDEc04j6AYtC9E5re+Ecg/i0iQZ+LfDMZf9oyAJZuZZo2YOiJOPX8
D1ZKqgHFQsTR91XGgcOol0s/F2GYePYD6pDfJX/XYmhVCzcsm/vpJqHtAhyz9mZh1Z7MKwtjB8Tm
874+4Jd8VW0bOhqchJm5qabac0KlWVL5OnDCsHTqiRstS/lnozdPJ1s+p2NFjH21X7hbIQuYUbX+
zsn1XrH7ChB/YLBCj9WDgJwGBWCFgZuX2EJI/To7vNpMGlKEyMeTQCo8LHUcY9sr1az4u3q15vYM
29w88Dg0OGznCkDXRm4u3Cc3PneglsyAhRtRp3s1PrYOql7RS8C9RS3fcYVz6hllTDHF71kLQj8b
s0Bhr4ojN+oqG5g1jR+927T9lXdWxUsCTVp1wjN+Jk9zf6veC8F9o1o6HXVwq525vzF1RZztyi0o
ulolJHF0Ylz97UP5SgvLIetc0mdHuIarpfWDxEvDxrThIlOx0uy24Mj3W3Co0xCTVQaxv0fn1IiU
Vbnr2QwaI5ZNGO1lBa7Pewfj45v3Nt4ShjdxtUt4PmBQo4c1W601895vLd0ELDRw1XDIldkXtei9
qdyF16QuhIOjbDYbhFy0wHY4Q7YnHmN0rWLeK2qMfYz0lDoSR1S1y7km9RpdzRjr/YTyhgywDkU0
tsJdIN5QRu21g7ZCUSeL8tolbcgS7pocrKFj16u3C5es3SlSO2el5sT9x/BiU4Tb6V0OS72CcGTa
+n1V5FiqwYhu6QL6DdQAgeaZk+nLJDPTQhjQPPZqxmVZq/J3HjtY/iWx+6+0sKDr+WygjiekNXO5
qPvl2DKq4XfVY74841IzWSirRDmG9ksYJOLnGBIyPInbYVE+EDtEM+chDzqJzW1MpXrIg1BbPkP0
TxIX+mixCZ12Tdia7003qCsjl0w5oZe8kZ0bAC2KWntmUXLKCwuFWNeJkVhZgnkJrkgI8t7ebV8m
+zW453SOGPh2ia/h8xN56/pYokKYVudlZCICP4j7+amSlUzJqgoiB+eIFi6wnSopIOd157dP1eN/
odMiNlB/16X8tLpQyDMY3tQHIMhTeTU4HV5pi6XGTKNOThrUy8CPKZ3CmiqDcSmvgEQELQlAoXhS
mxaAkaxisthfkZQ7/dioPyiLp8ZDlJOmMp4noKTETS3cHwmnY0L8KfA2fAiOfuEDbDcBlThxyT3m
AXY2OsZIqMHoRR6hoZzh+bPjYk+xaDoAJG9NV5ZbcxIL0pfCeOLHJYTU+KRDVBBtDzSoK7Oh5xJw
iJsKwL3hIAHu5U/oVib5CxC1+ZYHxG/a1OPVjLnnDZP+Yd001c6BTLqq8kCqFui7gs577A34NlDa
adEmBMnV5dfQxHjlNVaK7MTYytjpclOdDjJf3XamZTx5vG3g6OVcCLO1cxV1hyAm7rVhO3a7HQmG
Q9TQpMC5weutapNxl7P+fQ2k4TxTOyuH2bu2UWKdIIe3cuc9x1qQZ1HT2GwOvZILMnuUSwbSiPn9
Ua9Y76RrkS+dQC5g/SiYjNmeOjxgMoqr8yewUiC1tooq+ILAZZpd5EDzQfKFP06ygfIiP5vY4cPh
TbcfLDy/Sc8IkslrR6KtLqsLNtEgD4e/RHUaWgNxatIKsTYlHRE03OOQ/GNK0YAoAUqMqnbYuA83
LMBK4m1fMuuHy9qydBLJdctr+McFirmn1DLVsWxCbiQXcylksAly5wLsOWrGj/Gm+duFAdC3lpoa
h/DTAe4Fwzyf45povJ/gGXzA0Cm15Za36yj2rNsfrFi9rJjkmJUla7cUytL8fgomDyCA4bRK4/CJ
M7d7U7/FCmdM4tdbD9D50DQNHUIf0vMblqSqMCrKMZjMaLaCmPz/B4J7pdVUvcCAuWb+EBK/ZQVU
Kp6HDm3/dyTDRa97N+Yl+4WKodL1g8P/sBfrkdEr5rE4eRnWDKC9BekKFT3pgs8Zrzd9B3ojbn+N
l3LyjabKthRHigpn30V6mRc6r02ot9gVtU0Ng43QVMpuTvusJ0XFr9AUx5CC8f3du4kkRcO6QURE
Xg8xK6YIequBy7EqCbcI3aT2YKnfiUFwrInwV08uCA4iBg4cSrWdBr2kTQZTZYkheJDU05s4xSE0
pfRBV8asPIr6gy/3phbV7wZ9CrMqBYOTwXqZrljy+W/y8CvNZhMEOXV01CMFrITffPK/kCMjOY9O
HNXfyUMGqFomHe62Xy0k2FmMP7i7IYOsW5dgpyphW1RjAncvDi+nTcPS1cBI8bjz2Kqtgkd+yABb
ZpHvE/jiBBZaTrdeiJyQuk+68ioAcPiyNdQ1G3BttkyScUaw3ZZRQ2JN6FCimp8y1RPCR9/VYbO7
xJI1MVUU6Hgzs3weU2Ku8V7M5kUFi0KzDls9KGiWameQJJD4DWmbAJFuqWLcJz4rz5g+lJ7ZfQYS
bx60B0jPLopAUR7UFKtefZcn1Ao3OS0J8alqQHT4y03YjlRSMI8TsKHbI0DxW8CzYUSBwnqv/DWX
BOe54KzeowQQGqk/iK4cdvIQ9wwYJeEHonL8xmoBWnhG2GAz5w6hQlqkgXUEHdTBlJ7aGZ3RdLb+
xLyvkxAFtzaxYE2kL/TTts9FZq2kFBHHpAzdgegyABFj6CFRHsuatRrW3qkocq/Jiv/706J5wxIl
98Q32cY25q3QgSM4cR5xoLv26BuEyJPoi4iLs3nqS6UG3oo5R4zvnf0PyaM5O9b4f/DBLR5YUyqS
oqREe978Q100vAYHWiWtxebz9kb0PeX56L4I3Uo/AAT3QdsgVtqmGy6aACuEbDz68AC3mVoP36tf
wdOmlnW9jqpQJGKFJ1rpn97+gTI3q0AcE4UOqf8/gF0eOR2QAxLlzb4eJfgGs4LHRNW6e9+9u2Cs
XTj9cXlx1aNlYpxsrzsv+7yeGeokP3UGrNYLqAo7mSS54rbJf9DrFfVjr9rbei4WHe4l2zBDZWN6
8D90WaF7EcR93Aw4E93M/67lNZc6gxB1Lnnz+CFIKw+8TjAz+W2ke9G9M6J+2PIF+pRzrb7sA+oB
h6ylLiKOkPgZWTpjyHo+Rg8FxBAX5bLy77qrF+rsqWsu/C7uuTZ3dQS7oB8BhOZ5Y8a6M88mzSb9
UP1NchVi/8vO36DlEwXIo+/vIy/Nu8RjKX0fPDDm0p3MBPoiImiWGGEKhuYwefemRCu1K9pViKQt
Q/hx25CWhMaBk0qE2LgFWnfGX1U8EZTbE++XNdJOlfgscTS09JL3ptFPlla2SYjbCoH043Qj+x8P
4B3jAcIpr61HVRgZGGSmpEO9+4JxIlePQ9wEANdKmPlEJpMBrOS0Mh6mNcYret87gRlS/eczJPw6
UC7VDTzz4DWQ5uK1jwehvYHhnnZCOmQqJy0WC4ugJLgVlgMQDHyL+V10X4LxJlAtoTcNDHH5mkDk
OToYozAmB+c2MM2VrHch+JjU4QEVUBe2ePxJg5mFdvp2/jXdzHnBBqk0XwViPl0/gesVyOC085G5
s7DUbaf98GByE6GFS7hPfNWr/AbyLli2tq7GRF346JFu4tKxhs9n/5mRA6Nbcr9Ze9stWc4zlEed
L9EMGlwMW/cdfut/xv9dGsU5O5ZErEQAXp2dXmCXHeBIV3Zp/h4VxpWI7D76tzxWvgfXfk0fdzYo
hCj2dNt2Fdd3YtbmohayOdWOrkJOCgqYEHKRdGQOIUMVvRMmaidjdEfMWx/ZfZiZIkIX5hA4ekI9
GMvr6XSv+pCOWpqgIJufAH/cQeKPyFNSdvbNSE0DFApl4Gapwd7/6t2xTy3wNwkErLpy5nfCVqsJ
RjP+meBESS5rwCYE+d5Wlgt7LZEAvk5VkVmQf40IoY93z3bC6hqMCeZlVIgml53mXicFpTkFFQuF
HcnzdWU/ATEFKHfet8HyBJiCuQGndy6EdBvuBWiU+Me6QHnDoIIMXuacwZvWAodE1XLP1leOo75H
7Y0cRC/4U5MJlqozBZlMX1iPVZODm3h2oe3pNSzZdmDUx5KHEMe5w73AEhQshQRpZ7qewEyujCec
UDACO8UyZez/DkQPfqJCeK57kijhMxHI35l/k1NQVR7dJd6NrOCihBpCYe+zIkmDsVIfQyPsJISb
M/hojpBdPQMDEvqO/rd916+azCtLINe2mT6qMN7bfxdfXI7WjUxhmzWKEEdE3czIYSW0ciUpTB7Q
wKaASO3/wHqzs/UvXqPiPu/bRpguDmVIloG5fRsEmp9HmgpVZdRo/aqzcgXZnn6qXJ/kCTiSdOEx
n/g/8dJfbv9r3MzF8F5v/Td+38iaiIgblaEio5kKrKoQXylXOSRxA3IIFbKCrJTVUt6ayq0FfSgB
D3tMEESkMwJAsoQkC2OOcCHJPmUftBd6M/bEhoTpDwi6eBiBx3zBnRdLp7w4oOUgB2DcUA7d4fy0
MXoG6ydgjfIXFbRx8GJ1p19+0zyyX9E6MUqMqBUP2+pAgDDYz7TOMj3Oe3XKCcrYKq12b3/RW6mB
ANyS3lQZwaoiXVku3UVPGNhpHQLgDIBKMkVHoH5ocKQYirLCspsT922tc9q0nPiPPGsLl6iXd/M7
7ItHIZxBTA/dF2D5gshIqoPMAav+MikxjSix5/8MldYowRXvbdioLVx7JY/HaMz3ab1mqHf+MToC
abssqP0Qrp+DSwfnXjLgrO5Mvh+JyJUeE0WeIQwdayOxGPc6vlcKrrEJImENP7wZWj5o0/dUI2ID
YZnflPAeiDnSDC06Ipyi9E6g1D9EI6lQitK3zciIQdC0RpTnlFknosEU2yt/SLDtxuZQ3YxZCIu6
FfZA7PVAGdjYC2XFy1AaoO8Mw3gaUv37qGlIEEeNNPeWYV3785Z8AU1YOfAuX5p2VsDvcwjA2Zmm
iA/WTvxq0XtPkLvsdIr8IWxE79a9DT5rNIbONjqAmGi+uAV+e/xAoQlhXZKtmoJ/ytKi99Y8M+ZJ
EZJLghzfSzVCMhFlD6pIYWmjoWMRH20vZzL1xzO1vy9/0iNQHozqL5bYZ4bvi1ZWWDbFB4fKkKnI
YDqTXDCcINYlfJfqFEvCSR7L9CIi7op/2ZQSIWZ5Nnhs+13gilsXfEWd+tyelhIpzo2SbkCJ2fq1
yzkhfHq34prEXczJZnE/RAGtsILnUlVpeZ9HWlpb/6bxxU3s/kZoHZn5Xu4YRuyrUrom0Qf/2vxB
0CEeSmyzFYr8C+KD06Jal5vGuH7APSkTO+T0gXdC1yAXyYUwXjdqZvWBqn2cqUMXF+na1hmcNhNP
BZZbzm+XxFShT/iCkfr9cjIVg9wvQ+/auUyl+ueq/T2jvunh/IZsBQNnZhWFXwTwrHa2SN9Z6D3c
XobuaVk1zPid2Koepd8fyj73YGGAthX9aPBjK3DmPXTvYZXl125UlZLiODNaRPgEKSfQByQLaDOv
FcoO2QDIUHnrkG1R2eIAMqt+FT3/GeicqgQOBEQzHWIdkiPP6FrmzHvZ+Zd1q3KkPd5GhTi9bvQ6
Ry0BQ5571JwaQdgT+RvrPGsFtD9asd8bWWRuJS1+EDm30b6WwkKeQCl2eo0ANZP43zoARm8hQiiY
mGFI4Oa3WxDa7T4O1PzhcytRdBL2vKwakHOJGnKYnIP4GiAKRxvfaJejAiWZGdTNBQTuV90RSZmO
sA9o1/i5+6qyRa14E730nzhNrfu+m9lm1wHtJmyywq8wNfzrmPwa+29SOk/4eOpISsxXqHnZH6+w
NXJ30AMC9OTVi2GkRbfoN8TAt7jTWb1tu5O4xJNfL6XsdCEW2WksyyJqN93CmvOPnbQ88M8qJU2n
cz73nPXi0wbzFg/q8TnpRvsHoSsateGRWVFDJVuzUS2voiDEAzbIbL1XKtqnugoUkc12DtCZg1xJ
pdpkAMFMhlx9UtfVGaskLwNqqCqPckmqOXFUUxSDbY6f9R0R234vt3kSfwR8Zh08wc9eFYkIOewI
cKrpWnLp8mSvVA85AthEFXQf43GxNXmNfErnp2k2HgbtDyhsLLxksop/v3Nan5L+B4ua3NDmrx7a
wHz7yGuN06l9iwtYlg43otCkaI7FM+0BS3oOD+JhAcpQMCvyfB43telNi7czdMi90Ds3xZkSerG3
J+At+1D5a6h+FshQsgjSqcZnw61hBGln9uC6ioAHAHH1vnyt7c6ZldaHVAlDZq8KNN2SU5/URoC+
rv1tazftU9mLiwfx8ReWMm8lnkYSxQJenxhD/p8m3Qg8F5vQ6HsOJnrDCVXSW0v4McFIaUHIGfn2
lfEepHVTvlSNc+aOHPGv8L/yZuB4NUmgEj6VpdOrqcKh2ti3o4xvzY/N4D/zuiCuP7KE974aX/op
RtgpvPRqx6hChLH4OsWbChYCqmDQ+NiXrJyat8AFE7c5tCtadH/1aFszlY0l/gzEH8TEw37hdciu
1KzvGVbRVvR7gVbr4SRIWYmr55nu8jbWKwsoVztEjHFu55xbsiwhJnpmXwpJkDpy/H/Ch47e8Yru
GCRWQOjuW0Cw0Y1i6azwvDKgqbbmwSrK5c2xxMSkN0NCF0iQ+ArMFio/G3xaTL6a6LmuLRGY9k1S
3s6ca1+qA68wKwHpPnPGQRs8A6COfJEoKfcmCONBIcTgsLlnxlYXu0Vz8GOaIIn+AzKLZaN0F0HT
9Lrp066tt/Qrps1gnusH623fXMyMY7IOpCz3fpKYOAlQbw/y0TsHo4tu88mEvsm5ZM3rVKuplo7H
Ll2joM9SpUA5J0IAcjK1VEKwIbm5b0u04YtpQ1xManLASSGLxH83rolv3J1hC9/gEhJRPeEI+O2k
udlWNX5+kQX4AWV5QjMnULxOESi7gDyTIi6brdgq+05BYR3h7/ld+BHs3Sq7akS9kAgZEU66kSxh
88qFheHgdYit6LmgYDHF8pToG1uwbOhyg3KMajznNpiCAezawNG7w3TA6Rs0Cs7WbGcZoRURrm9S
IsyoCgsLSvx8sxNANQYMvUWE/0KROngjVb3VdVFPXA9hXY53UY5wgUzkAN2Crnb02U/dJwNQUCJd
kGZjJPAJaXYdKl7pGg5wcs8Kk5XbYy7w5vRAH6KLsB10DAbYS1hgnaxtFUwmtVg6QjKwxkbN6CNw
ni8hajN/EmVOvhuwP9bwWOprRjWthC9XAGYivG0c3g5uzpU0AUGyOoTMYY8sNRC+WIZoC+wa6MRX
9R49lgOMRwa3RSTFfCKpf7LQEsmswxGLD5ZCGPcvVg0KYvtAP/5OCdffevhtKsrwSDjcwYQgOH2i
Bq2Gb6q1Quottvm+ffDVJnR2QGJvT9JnokvCRbyIikbZPDppnDQLreRFO8egz8EVspECzu78gJPu
99Us1sQAwPaf7nr5/9YgJrvk4uSzUs1l6q/nxJPMSXYij8gVYcpSD1NUJWTQkH3P9ZvtWytbOCZV
JMrsweAERa8HFDA5h74GlEikorFovihSejWK6IN9YyJmkB/3cZJRDxjJ5odWJipzDV7hDC7ql25U
HPB/3HW6Bxe+V63UtItQHVkcJ4+gFFqWHEDXqTVTYrvpG0bsH89j1ywdpn3V+Ezz2C5Qj8geEkT0
9hKGJ0FF8hvbKFLan3w6GnVUm6k0L3f4xPeXvD4XbDzuBU/gvX2mO15IrKP3KNR4qOQhK04JJ7BD
4pwNpGK0c8a9nvim3zS78qitLHpt/OeDLMHJm9rf4N1ciTSwTDJZ8Xtfow/DDoak5+DxXcqpzti2
L/Ly6DISb+/d67w3Acluht3A/dNTugLOcSxhMbEMnibgoxWlzrl9s1f2KPe2fYVcVsCkAYx2JDGB
8wAHTndZJbP86UkGYloNyZed3Rf5U78lcXWf+e1bDGzY/a+UIh4jY/f3w8CiluWJsGE9squOXLk3
30UprubvXOVbwZjXEo5Ihjph8RiBcRKY0m+znH6bLZ7Ofa4Yk7Lv7bZ6v8bDzrN5v9d9U+Q09Bk4
wPedF3B/N7LJXVWrU8ol7Us1Xp5ezaRAmRB32gd0fpOiN9LcaxV00lR2GipH0Qa88SQcjPVWI6YM
273HgBK83CXYuZBbx72WTePM21uGFgMLsDyWGHZbDxDvXLzs7/qzM0RuXk6QuIWqd5cmARUzhMUG
Jw42kzF+Ir1lfLnhnVmID5h12wpnkRZx1LWJgolvshqm2YIHrL3FEGSS++kRHtJNhjmznVC86tFo
PfpNkPz1N+1OJuIWBQNuHhjwXC/r2vvzjQyMGj44hv94d4CJwXzQFLss4FJTfURbgj9FyaYnetOG
bv/Il6eved71Tw4WShSSeT6wVpslGNZk0SYF9Zb3GpeHcwze0YQW34f0U6JvnyQpAsL10paF6bfO
OVfT6R7x1Qy+9nJs02Tf4ko9Gp74c/tSWB0fy0DK7BQ81YqB06ILSRZ4n81nXEpJMoKhak4bxl1r
f8MBj1VWzAxSUQvoznHCtIgpPy7yKZKcDOEgeuKq5t8Ho7syh70fG4FAlKBYnVHhDMGG90bz72Ew
EMnQL5ewhupzfB+FgWwcsPoM2vdEu2nLiKavqNsfqufA0Ia8wnEbX5KXVnHSdVaQlj3iBSWPq3BH
6fBIlP1i+4tJDQZhl0etnfopNT8zxIING6Z0HuLZss1+s6znTEgAidMUh2eXFUq9W5d1Lba1eG8r
iAm/aP7Hvc4be7tLZS/nXi/WrUNQMN68olcBkgcH39+O2nTXTMhDM4Q3Vcao1Hr0Oeq/9joor0eb
EkdrN7RJz54idGGL7ApmfbE9u4cK3Gei93irdPxTn6A3naUfBCAycqPXW8PSZDiuencXu3H+9SBe
I2CEYGQgGYoEURX0qgTyZUnyXkcCKMaya8zhutGzC26jiR2shLrjsiQ1yWYGTtnkr8g4bZlT3cVH
z19Hi9XeabnhW8NJMnoJbuUhIrsbvMZdxwyjtIAOrkbJWsQMe4Uk9sYlH7X/6/MKs3o8iR0cUqU+
TBproRMq44YpcI/1fwm5tSEHxeFM1CK7HYpWBncsyoo3Qy0g1slQAFvs4HozZlbQRXVor0Y0p9nY
AQhy5rlXk/xHZsKBhliRC7KBro3lrVaa2kkmLxwXbHdH1Q9LOoFctZ2Gz4KsdBoyFDAl04J8ZhDT
EeFf4cyg/DlXNttHCNePvkPLCKoCv/1yXjnEnHy+RnpBKaInDyKOlc2js3tHJaHRspuFh3gt8o2W
EuIpN8H7pCrAX0dTw/Ct6cRloDI7y9an1GzR3kNOrPyMVEj+mvasbeLvLLQpJ019mlxpAts/1u0B
1Vs+V2iJuyPXnooRKDMGpcYKmcUUF8+qr9ld8610xUN8lCKiU0tgxGDIoy6YtnW2N026Qk3gwxTX
EbgOR/zxGq7gkbYSM+Y+bxyLFtYaGtTwkiVudDAF5oKUnxLsi5SxYsGMe/2H8RuvNUYG8Icg6FVf
KrKq3RtEjFwpuVEqHr/5eZX3XCXiRBduZs9YrlsQJBjrJqNfOlw5DasrJUud3HbSQtJbCtcGIla7
LlyMpaKyH7MSHs26QCT6UkKjL77EtBRe9yz5jeYY0cFibl1jd4x/d/zMWl5qev2kofnRy4MSGf85
QOFNOlbYvyxdA05VKGKiEvlHCRechHjX9+Isus97gANPPOy7ORrbBBLXYZ4nUjiv6XY7mxmGbqvU
zd9Am1ruNoGuxdhUcs850AURwFiYHikvuyKFnsIEFWMBmdi0JQwUs3NzSxdqwKxiWDk9SENCVTEH
ItDkVtdJIk+8GQkvZMyLjT6C7hmJuj0w8D0xlglfuA/YbHEqjAEzR2aZ+7ku40BRVpwO7jpFZtxJ
j7vVJ/AOD5mTz1QjOc5uullckHXMTFauh8A+OkrMwliV2lsupee8e6QluSGYO2iDSghvnOAIRWJA
9S2phBVVK3eKoOJgNDtGnT7nonHIOLL6GGpnadJhs3F1jVt8lXGt/RmNGnKKII+pe1cCV7m78XBU
A0kU/HPSb/Bx2Aec+dSPpZF0JWyuLVdrtk88WIUdaBwYth0LohapFBjTb+rIsQRqCZj4ASVjGrsy
0nApnPfat9z99Yb411JQll6Y84QFnamWUi3Z8sOBlNX6+Cu6j7vbdvEflGd7tBarcVSJ/ESrkWjJ
vFE8yOiIdri0IfuSJ4JQ1W5cokuOFqKk1pJiKQ7AFlht4wtzX2gvvGyvzznueFL0YF709hhvzgsY
YlYnuPT/HA+MNLvByARKU56N+HmlpYTikPbQOPawYLgXPMTMmJlW8wIV8ZTzCSirofTBW3tWPwJP
ovMjS6t9QzC+O3HqgvpaFuLNRAgzqRRBqo90Oo3a3dt2UEeAr6Pd9elVpdQZVWFDYoRo+U1simSf
pZ9nQRhOIlhqEOPUW7C2AUmlBvueonF3cUsIqWI8RS187+mNilVLKM/din4wbjm3FdkHlVnOA4A+
csl84I0JJRYo6khZ+AdHuZNk8LJ86Swf4llrCAijOny4T5rQTGdp8PlHbKSbYJhqjP9DwOP6JoE+
4uzjt9PZ5x7o10SOsV2ydKcSIgn1xY+uSWUuwx0FNY3OCLO5n9rzqTqKgaR1dEegOTNX/kj245Fo
u13RdfofoHvQqPt9IwbCkDq7D0rwaiEN1pKqRESlQ6DyReOpYu/dn6XtIzUvTdk7xKiNdWlaFfFK
wstPY+GjdDjM36ja9sLWt2gcZMsCJ5AMNdnRXvPcObU/8bOjAsoxSq/47ZIBCBqQqo4y+S8zan8l
aZKi3HtDfurEhzwMMP4TKkyKDgJDEruFhP86x8XlbSuJOpuFJPk8qGIhWskIgOrVK8Y1wYI+hU2X
nh0qv98yMoOTmhaZA26DhLFqgJFrGz05vOmtP34SBJtuFK6uNsPpeeBvaC2m8Zvu45F5bPpbozCT
KcqXIJTL3kIVbkeOt1z6vyPwbXWx99DcclPkbqYxToSWUOvaoem9dFHVpU+vauvbJD3VpsPYT5xs
ylFAxDXMMbjZWy+u43POHG7LmNxk/7T5yipWOEdwAgQOGHas0wbJ37eZDxGBcIY+265FggHosf5/
uloLZk1zBGtzLcboJUsi1jc3bcsxK/Aqf8wcIxgBmlCYDIVmTSl1GKfCay8qF7Lo7p8yY+027ItI
vIu5Txpu1cMnt7Iho6NKrAWkBEJIsMTgvDFKf817DzAyOVRwNF51MFHDJ5Gw/pOc6NJ5iXlp95ZW
DmMdZmd2cuYSA3nEiep4ptqeL73RtoFxNaN+ZXu+xwblnVd3MJfraJhRsNjsNCsnLDOuByfGi2RO
CU92jrH+YSSDy+rkTKy8yxJxWdsc3oP7LpESUR4ot35V3cFuW8eTZVlHGH/rWk/yx1eBNvcZwVLR
MiFJmhu4TDxCMBmw9W70SRDlsVN7gJtuurYatDS+F1oP5zSMz6uDspN15A7YDKUy1qQrx6PO87FS
kDDYK1wiTVThxzxBUiD4aaKqQsR8/SpKI0hJ2gN5bi9NziPVVkQP45RcgcGPhS0ot3hS19hl/Hhi
mb6x/8LjmpGlVUqCA8MV2endxqRIRFjS1SYnQ+Z2zOg0f60WVEU0PceQkjzAeHibACC6jyyCBGse
iINGYFJ3AL5ido3IQnwuBsrtflOhQtFZ/mTFA4nb9YYfZCo8xtAjY81sDflkohW2HBr4YG/anIqd
+srSvGH9qRbhHaJi6715u8rahVgjPBd3FTx1TChI9usmobL+PhbKhZFQ7mwCcZou8dePlSJEJfLf
l+nGonnnKi1/2qVlKEF+AOq8+3q5n3SCgiceICTRp4r79O5pqV/e+q114D7EH13gZDsAKfvJmSyq
cpbMQemULZVtLfN36xMupLie1psd5qMeeg6MDs+5BS9kw1hvSSv0oDsbX0lUYSLXgbzp1uR5UhOm
5sdPdKbHzoH8dplujgttKdeI4tkFxIosoI/qHIHDVqzPCoA2hmnYDBPfHJT5hHG/a61aUdaW0x5z
8zn2PeukOS47Ac00anvRyb88Gk8cFZPg/51TD4xAbelvAAJGeapREkclP/HCZUYCmXDSKvZsnMxI
W0Ns1SPPdfYg+I/ANZd3JVCFoDKSzUXr64TP1aqC1Bub7N24/nfAxfichjuucx4/dJ3uO6HGQxnc
IBSJEG2jlshirZ2P1LSsMncdjAIcMgaBevVt8W6eX0PU8K4p2+N1MeXuZlyXtUX8oI2eQZvBClUp
q/b9p3HpvbnSJS4rYLie614yhkCBpaOyde0Zhf9wvYsWE67UBI21ZQedSqykWFu8qKkISPVdMZrk
C9LjUZyLgn+e39Fu0RgW+jIxSWNyHWBUt9qZxcvg3UJxXKqI7wKzRYU+j/LXsx4ga2EdInnqnJ2n
PZ128p+EfeTdTZmgx3wylPdjKF16DjH5enRPqRBjbYpvs+8ZBuuHlyhaVZc6aCDspCUxmlT7WeLk
4sjFA9Hz314CfO5oZKvd1QF0hPm2UywgT3u/pgcg6Op+09w6xlZ4NjfGTMnz93Ha0OuN0Z1+liPp
dynk8b+36Rk1OI6MJlHtNTH9LIqgoIRQMZLb+GOVW6Oumqk+l8qeyBGP1uV0FzhBZvf3IKCq+ZXv
SWUy3d/faH++j+EVH2xKEgMaynJR9gOjBUQFIeswUiEDpfexJDsRZALFPnWvV1RgPeyV+pN64taU
PO4SSqjZD5GMh1WrZZeQcijFAtH51BKYxM3M2CTaloOVKMTJYu4m/IEn48VRWuaYX7DfOXSGyn8d
g6OXdszbl79D4J6VpZIMiOZ+ddf4Ma1LlOgk3cs61vZHT4PNxpGgQQ8bdH9wi2dx1Sh5/Y+PcDBx
Q1v59B9FHDkRp+w/gE/Fd6UNkQPWqIPpgLYr7tdjX67nIw7aU3yHsnPZBLXFb7ZBfQ9wThK4R3II
5BUET79EYOOk+OoaI8vj8NBv5p224wjfJWIu1PYAylVurtjvvu16mJKMKCwKzIY94prRg5N/5CJR
G7dOGbGm1XgWQJKGJ76Z7Imz7wXjTQcYznRUmWj1du+N449zAVGdrw3NhXVsJvre64cb51yoT6VF
+E4VmOxXH65GT+3sBjV/DEbuKvqhC4DIGvSSHcphP8J5tgQUDeaI9wFXK2Y3Q3qtJWKsLEgGwDvY
1CEFIlWvnkbNsCJWA9RV+Uwpuy95muB+xbP2keh6ASZA/RiNSjIgnCF0pKoQKQItAB2Lja8S6UNo
PuaJzZPh4RqFEnoc41tnKRIWkigMj0G7cDxav5vQCQxqVHjfaOSDTWQCici+mphLaCWG4Wmg9WFB
c9x6621i1dCX00iU5tFNGvKGButXPunVj0yebWnzyWdPAktotQ+MFYeLQYFB0p+0KbshJOApW0LE
AvXWllGuYRDMXcXGwYjYp0OVBHnDYqWBQy4lP5XYezIKVMwQrASZmzS0O8r4UOLJLMgeSYR169GX
xrhhOGxKCBwi/M2cXZi69YvbgXiru+T7kex7nlgFlFuh+5e6Syn1itQjKThz+mklrWz16t5uRZzn
/hMqo8XHeUgVJuvoRtG+q6ojcMUoLaC0Ju9A9Z4RNSonRZyUEr+bbAL0XkJzjGnOrsQfnKtfLJDF
ztT454Nhw0ZgQ36TyaMvzzivJLq4wqT+uh5KYA/qOCcibKpZG8Dn08rn0kbpFiHw9W2y9Ho09okT
cHDV1QqyddI0TDezSYNbyguKVcCO05f6QNVc27I2RO+917gu+Ht5ukCaJ3lgTVE4PtPO5w5XtpDf
H0U/ppwtBotnjUr28HbnCihVH/3CQ8Ptu2XM3a22zym88/EesQn8TrDIjXB2tGMNmBmY6nY7UIfN
PTO8kTRZJaGYoEAtSVyH/OFuoS4nhTATDhowoSQwT8gV+LdLJShYsjb9R5YbpAEE+ks1SdpuQmzr
6ji2IQGePIxB4lhbR/zNpSD5HiGJtTUArOExY5GDuUO10U41PhSuGvdeWLUDuV81n3dya10bR++r
zWHpCwY5giDsqPNtyIwOkS4Wxe8xvz5u+fGTOFp8fnhFmCE/EdkD3HU8IG5n9tAi5KC1/TxyFQzC
0La8S70Kf3WjtSI20UxV1WaD4m4se4X0SvaXEECb2aDrNjLGuVVDrd83WWG2BZTUadRy9+fG3rml
SeRI9mZ+AicmEJAeG7CF3u2nol4jlZ1pGM2/ixgvL6wj1njk1yd78ZMtQSJLgE0PYZsuT0zoJKVg
N6AKbAH0IvqEE1mIhG8RwoW3K27rkKIByXwnX9sejvJahgd39PUjiph7Gfc2kXz87yc0t/OdqDbQ
vrL0kssRoVc5sT3HpXq+DuK4+gfWeB3y+lkA7Zl4VAX6Hvuf+YaoIfU116DkbL+Vx6aBdVJA3Ywc
xGpEV3eM7KJgK1/2MOmUkauis0chgyt/es7HdzndEfC4+4isW3tFnmv3U+ERRj4/rmvTcMAvcoX4
/cql0J10bcTQeVeJQf+hxNaa4J4TCVT6wqzKp8zb1QaGy/HzWKl8olFNMQGq67E221iDAzOmKN7v
E6Kf0/10biGDTQiams8Mwl4VP+/EmMYIrvUAodeo6IEikXB+vunAHklU3vRnoNEvyNHESRzKDzWb
5QMuGQCRgEKtoJWQQvKrYfwGmTSu6JZPQUKh7T8VfAXf6Q/AK3qJ4S4438L9Lf5clYPly1O2Ia7J
9zzRop0ZtgLCp6YXc40nYzqJZTOZdHZTFZ1/QeWlW5hN+UMmde2bDTvyctHhOSKs1APM4FmM48Me
lnKEnnerTCVCwaLB0QQRpWyCcEDtRVQW8YPG0wGcKaTRMtIjNI5ioODfedB1Ue2ulYOT2RRy6kVD
cKILOZ6rC8lFkMKzq3jr24gMSkYaPiGNXX6ozLhhq9Y0d3Y/w2SAhsDLwzkoN9elxFKCtrBkzulg
+j6vO8AC7YIESPrWS17Lfr7ee/96fDQbzAg+TLNlfOaCD6aNGS4lFYeju6hWG7jvr5WLzYeQ/Mix
apORTcpxhPJ/CafI80d0hrlOno725iUmsH/NjERmZUSZCViU/Qr8CVo5RUMNwBNauTcOLWRUYMNk
Gplod85/GqIeWABGWKxUb1DHCzwU+seNr5tnNlaLsO9gO8iZ9fIrMJqMQqV0OQWC2+PSp6dsErUQ
rXHRkATXX2nIf1LTFOxmrBbufQfVkQUHbetkWx5gONXZgtWiYU9lVRt4jSY+QE68rgLTz8+yXxBo
jjLzwonwWngqf2iAGkP+QRLwHcsQ2NKjuxfQ+1/XKbEfPlxA+awV6d5/pxsr7Y9eEQas+/pXYgHH
l+pPHBR4l5LMd9c+zmTQrDZ+zHTETMMYqPOKoYfcItj57VyTCTMXmGxQND7c0kj8IkLd9tHhRD5B
DKYllSKl0jDyf/vN2pErKAe33Sy81FRnMQaVA+lVzxiIF57t8x4mQqgnySNV5LP9xiyNca1/VpJP
QkAdET2H7zp3R7tEybPsX2JEfKY5axeWqDiVKlJOSkOWZ/4Ot/FRTWqwtrrF1uA1KfNywflHQGFp
VW35/YiPKXgAcmgqyITaAQgHKFwVrmx2KKk4epsZGaksxtQlENMadWhfL0izSf5MNi9opevDIpIG
SCAi8535iEteb6oR6vQqp8R6MFibw6MtfqXxPPdqktEEFcuBjMgqCAtwGazQgMLRa9YyPId7j2QD
IyGGLx220MlFzcoYFR1EA7wVy2DYpc6gIvrc/VPaHs25TIuF7y1LzSfo738s5VSH775+ozZnceMc
ObFJEWOpNAWqghJsxazv/BdUut7Ck3Rzi6dcNqDuMfzoDrfYt+THeej/rqqPzPuhya7UUwboYOCM
P58OF2yFGf4LQRK7GODtzPXoDgbs3WFoM71VIqbkz/3YZNKuHisrdlri5q/HkDFPCTZGyRR+PtWE
C3B7vBgV4/uoemqCEJsezQGudLwXe+LpFwmT8xsaiMlphJZ6EmV+Fp0FH+Gp8+53M3L+PFhXX2No
nXxRgYumg63R2HnrdPgMVGMfiHAaXH1dc3SM+eviKs6uL3Nu6EDbHXqKMggRrfbWLpH94vcxbx+m
rYRk8WWJ5Er7buYD+WqL0A8Ql3PKBURMjbsWdRLJ/3N24zOkrQvz4a/9Q5FDrDYKS9Hsg9rNjFM9
vIP+F2i/VcrlSayG0EMqZlJcO7LU2+zinGYZsO/gQ7x3b8aCHIeJCkgXoTnTSA1enzHG8vpXlmYb
ixsdPUXTMRAVgTKTUM4zj2KmQLGrBPkgRTBt7tQiaFiUawLc0yXrcp7lpYr8EQsteYMAXTGil/9l
7SWFM/hfHqf+4WihSMBxp72+zVBgOktGJzKTpPAyGHJvygmdQ6P6SS5R3ejcjOBotXhzpoGOpQMj
VIFX9cfIJjk/HYp6RcJ8dfoAgZ52THQYlmIRlLLZxcKa5FX+6dvZITPTub6DuO+MrtasfEOcF3gI
hNxh6VR39omh3sWIh9w0oy/z1OK3u5CtkVgKT0XCTKolxnBDRaf35wEIAjmUGSrZsw4eqEf7gxMS
RFAiPwllvum7q/s2jsfkhvZzW6gfw0g/o+nwPSnuqZFt/DBlkA1vPswEgS4a+jCRk57JZQf9zuRo
RMlaokmhaHIEuCHWKxz9yVwIo0zmMeesvgF06KDOgvHScz1d+dxIge4rZ4fjFtXDTM3HGmO3WE9i
Yb0OVtNc+Fms9HdTF2/xjSjfRktzCWeLWyXEuEWNeL+KtE3cOv5vbZsUHC1cok8Z3t7Zh7c4fiPp
OJHr5f5Tn2qMAfvd9SUoCq8KeYxvpxT3Q7/YYhRHMx2CETgXqnBqrdre9SE4GqV6NyDfq6AaokoB
Tt+JcEAUvDEi3midiUl0s1M8uG74OZX+Q8lR7+ND0bMNJE8ZYfRvtd83nC2QUWgksXb/oW3osV0N
GfNzTQqv/HX6FuLrJhYjWImk7a5hOxWI7Ls2moLWskwHuPoJZx+E3TyQlepILM6dOjMMeNCLK+vO
UrGKAt5nl3N1L2ShAQ3o7LjQiZ6HGvLcWYbuPMOOEE6ysrXkiWn7MVh7Z9vYa7wXqSK6/eqONSFs
NLV7v2bWNfw1a/R9eHolV8YkwiZT9P3vCYni8yZRIK4Um0/387nQtaDDFd/htRnCkaL72qQC139z
N/U7Yy+ylOO9/4n+tIM3NL4O+PTbwfmyyQKia2lV5qUfKOE176vr2JUzH5djMv1Y1RuCLUZ0cYVp
eDrtDzOsmAWiEKDvAsu+DhmqNsa8LdwkiO0IUPHktdb5iGGWWYYpNku/AVda7ZCd79FNA3JU9Uw1
4DvGq8xi/QEZifD7HE2CTw2YBzhJ5/IPVywalFBaHueboHQ/VwL5vb+/OYJUkiVEPn9qm4aCdPKh
ghezg6LN5TnW3TaGCIW3XKHyiQCQ+F0BFqP13uPeQkUu9EauNZjnVkYBlTxrdh3izuvGUsjOn18O
5Y/hv3AROpyK7QWMWv3TByRV7p1CKA3aiaeqeOSAr8l64cCoHf42EMEn8qaeUBiCW4jTxz8rs3gY
Y/cWSndtvrAFv+1u7PYBuH/Z/tCP4T1sIb3cIx6QHGYwxPQkLtcks1Z+ytogLDYN7JSPMyRCscGr
b1HTpn4EDyvUO0V+Mzi+zmNEoeJkh5Zzm2BDPn8Zq6jH7zq4osWy1gHVy0QjoTDMIfipzP5gqaFd
RPjKiwx9AOE+F9WDS7iA8p8/84pcIht31BHD9u+gjJe9ISOzxr+u84qRadkWKifQGH55naKZRotD
R/lYAA/1nOVQ13Fpf9iO4M3HSUnQ8HQ36KNOn9Q+yV4M6yn/dEFbFYJJiKVhZkhpEaoSOEDP5Rdo
2NpI//Fs78z9YrYbyMB/3Y+DEiYj2gqlX3Bb83fjlfPs3MiyE0V/mt+JLzkCAS0qp/4IcBOH5wRB
zIEhLibt91lkCieYA4u2jIC+lAn95dFAuxgwnsmx0P85dZU4ICg5V7MvDtaxb43KlLVDnALOLsuo
ZQdaf4uSc57hgt84o5DzPwHXuMzx2iVj8hLAzUwcAmtb8lixV/iVgj455EHPI9VEJyTPq9gUtR6N
5nx/sHjYp3tv9f6u0wOkk2oG9eLRxHXAubfAR1+vIaS2gWYJXOKMeE3leaCj5BAW2CN50cCkYAqE
MPKTKKqzsKq1+18AXvBLJQt5N46dkhoc9RUJB0u5ad/DvnyKgFQ400XjFf3Uo7LtAhLmPFm1jWXv
3WvEQGzoyhGGQOi+I05/ORKPeIG26Q6x62cmDF7hfU8VrT2eB4i2S/3qjcxll42gP1m2L8M+s5P+
yJ2vdEqGmq3+5Zf0BU+DNMSvg3VXUlVcIL3ZUENY1qKQI9X2YeR0rKqts1y1MtNSmwbJKige+LbY
2+avQTaC4ingmyM5AyGrjhKuwMWsHMuyPvxSCJnq6S6cImz68kPmH8JEC8bxFMW1P5zD9aFzXUps
5imc/xgtxCrAn2Vl8BM18YhCjLdKPzbbm1TFfV1DNsF6BaSfpwhySX5nIndT8mMFvE4ox6zjMI/3
yZrg3uJuZkFhg0J8CbORmMGDXnMDSH8/GLYxvx12ugCKLntfhR7Nnh9OJoR6K5wLMwl6nNUM5b8K
RxQlMsBxX9u9iXXt2AHE6txhx5YcfyBxaBsSbiLpwdV45gJTByDW7dyeZsLkPo4VWf6tV7ib2vAR
qIAvMa4SW03cm13djaDBRiKyk6qwTg+tBYO7dORaB/78DIpEKhAf/Gm3k9Aknkj3maHZyrULzqG7
LIOReIwFLqPalwnG31HMnipgMW/Sz8NxV6IBhB7q6iJDljzVXxIm9BbS+83G4N5Ni5CAuoNzBOjp
NF84LpyUmo7pvrc99U24MbWTsoZwa3h7CflPFH47cgmq8Ai2FEjVmhF9qhcO5kllbHvKgCusb0xC
2wBA19HwSV9iDKU2qI2ya52uKFDgkYpE/Ey0tMXwCDFOoEFORqqLfEl5sHPbgz8lhvTOuHtrjClO
Za1PxXWJW5sijKs6aaam1ZV01u4nj19tzsuAKzhwScjHE3E6+I8ZOnH80FwN5sEiFNjk/SUHhv0v
zK/K29UbOJRzHWHgz5uJOVCGAwY4RzrHPddtSbLpg1fcwGRoVosVl8816VsRdmFMIWQIc4VhmZkT
LMWqud2KitfPLtD1veonaJeOpA7N+W/liys5SF3r/XQCOsI2nH3UX284YYx+EN4Vd54L0LK8abmU
cxwfyKuEcREFzGvoBbhagzAYmZahpB88Jyv23iEfeWqFVjBi+bk8Wl/s+/5tWM2ZuR9FdGmIXRS3
pg15zwvtm8datFnhI1Ztj1Ns2Jh1HhvYVFFJK+YBtsAMamBMaNLbbLNxzYKn1/0E3b3eWWeoadl2
UmkupH6DhdxKVAm3pci7VD1E5D1SUszbBHEgVjoo3l2XmNeYWavUlrKmgYRGS6lS4BDCtLVWRYLG
ihEkqRiaMAEBtlZIwTkJiomjhE5DEYWXvjK48K9/iB8zcTJbL8naKXEA/eB/PH8jfwK5OU/ZbK8n
smdbdH/XNRjestjf43wRTNo0umC0szdXKHTyfngHMG9XqTYeo++yvUVDjVdDiCWC3wIXAYIKv8Qb
6mX77l7+CjyOSB07wr8TGJr3fEuOLAD3BgSKyZTlqDSsDSSudlH28TbNd6U/+9LJrKb0czX12yuL
7g800loe2LGbi+p0uDmIFnvwyWj1jghf7SGCsptZCqEOLHuRB+mJkI+iOUtSOh095o1Jvs/mCpEz
8vgqcd/HTUDKZ2c1/3QjuCPV8a1nVtcVV+H+mHkq/FR6Rw8j6CLWCYKCEH1O7N55mYwO7f6vE+tf
mQG8SCGKIPSQ3u7fMnn+00hJ3frydhozoq83tB/5Xf81qUKHnE0zXxqkF1ShbTT85LbpKDbqyk8b
mWGMlERlgZo/WEE2lQ7w4H6N5LznyD6hyHdlXSkWh9tN6Li/3+ahoYaknZZD4VBifdTYvHQ1DGhY
8Rr0KrxY2PPKCJO8OhmdBf47s4403XqCGHrWGgo9kuE1G+d/hoUlNemr6OkG5fwgdgYj75tI5koE
lGUxkNUdn5jmIcOLdMJ5mLra/R1fvT+UVHazuxd8w3a8rLA3LrgtVuz22hx9qSpZXQOGcfoFgSNs
or1P7B55gTgQ4TmHrgX5viS0pi6gVq4EwT7kVG6qHPzZkF8BwWxppZdvCe1H+jNQhDyw7mTd9olW
wHmJYsZiLww54hrjWQ1WRQ/uTqLVX71uSzGPoANmTbPois8CmfxzQTBeI5/U185WWR6zlGk2Jo8f
e/Cl+AAlRsFyNOm4WgYMWqwSHUYOFnzHEULjSJtIUq/g4aHLmyh8ir2UjoKziIH/8ewGaLnjkody
4glWPWmEJrTEO5j8E64T4YiqT8eei26faZZSL1FVMJNZZaPF5YaD7k/l9DWlp858RWexVzmyBqj5
Jyf+krqYgSyGRCIG3R6+BOWdxEZuEvgi3Zb0ZGUZBk52PihaJl+F8Hk26fbvqhGUbRc8nvPn4qJL
4u4VZt2U0oyzE8CxrID5TiWFhyKWur/tIxQjpsOFH28zqvlmou9xTeeafgukzMvjBBUeltqNHTjB
uTi3kKONoG6XeCWqdgEo239KB/o7PWE1f+MPleAkjyYjlKcLXpwhkPuZTV3v8Yy3vTMmszYQPrZO
qhowI9tAqxSEu3dp82R6PN29yyecHkSKp38nGOoUm5HWyTfhf5ZzpngASYf+0Pdeiz9JB7oVZUp/
kLB80g+IPeM7dK9jVXyxB/SUBibppbp2P0aE8bZ45rvzvDo9nLGAOT1ie5gmREpV43O5bYXemxrE
U/IxmKxORXxCi0UxkIunIa2IpsF7aZmaoZhuUVlt40NOzpqVcqbx/pOl4tAPju3Aej+eetv/PVj3
3PiZZj5VrAFvCleHtBM2doWt7feZN6aiN22uVLH7R97BN2JG1naWe7r1oc4W3sp0o4qkolTHvB4m
wwmZvd20U8kC/DqNbgfitnpUnD10WYSQZ8LOXgaFBY0sqjrlPdsoL1FBgZU/5l3zmfcaeOxgp74u
uyxGmFHTM/MA5R7pJ5D3Mhi2GsFxtkQR/h5Ud2d7wJAfPfGdyd/EwCQhru/0G9UiuDeO7ehVtKnQ
zV5zMaW2jnLdELhUEvxfE1JD+PYlMQ5e3aVNxfKi6xImeGtouVVcGYAEJvMelhzCaXMBJo03Nz+P
VUyNJu+UPK5GO6G8FowajrN3J0BaAbKmMAjTLII2RrtQVYSw8mciY3avqhrt7HPDI7+qcLXXIoS0
zVH5XQ99hNAuPVI10yqQuOW5Y8+AVXUBLwP4fdFrVG/ey27UEyxURFpmIHNRHfYLJ9R4L6+iK7E3
+gJqxfF5QujD7wGxObT4wnBPmyiWa5NOZo8yQ8nwW9Flcr0gun+lL1r41s1PMriECPk94R/CoPLV
/f1qQiO+uRkgt+YwCL+SB7IwV8h3myF6bcBaI+3mcvzX2/JIE4KkzDQHO+3dL5TQQ4zbscv2aHoj
0p5MTGeSSxUfZxGYqxXLlsiv8Ia9cIu4sfDrHql7asIGeeuqmnjLrlNBtrEOkKhFrNHeIIYKP5Me
2WPDqANNSJ+cfAQfbhb7uh2IbWnWXyH23VhUciyqbW2Rll/25j8M3KS2e+W2SnJUDSlVtOXBDt72
y7egJo6w9ureHY+cDNmpgBXxdcrTPbuaId95Hno0asfN2q+4n51prszpjL0nWTkBcgVbuNvTflY4
HHGEXhTLh7REnamVZxvBJEBWJgGc+Gn+sXZWxqXd3FJ9TBHC3atfd4Oi9qGFZMji6qSceG82axY5
a78aIc72tW4arh5KaHj1DeQBe4Q1edLrZxoSy/h41junvDDmC+88dD6ltga+aLw5VxIGfNYOc/9v
ZJ1/qOijIJ5F5y2GaLZIfaSMXb5WR/HbhTWyY2MGAr1ziiqNK7EAi+Mr8He51WwRqP0iFlBmDJZf
3wEOFpTreosj1ax749wXSRWWJFkA7D33gevbEIys7HJI71mUc9pfHOT/1hzznZJFV2rZw5vZ/UMp
kLOGRm2tLbCipsXXebq2xquvDr00d6JLf3OKMr1K8vn6+BuQ5jO+NZHhCJFCh3D7hGv06iupKDMs
HKilgDdglqKKHj4ux3wXCbZ5hN8fw2Liy1csm+3NUkTkSvD3753FHsSx9DnHaOisk+jF/Ppcnphd
2/qbDjD2SLoetFF7F8Q3mcwlpl+/cwwrW5TdpyD4w0m1ORa14i3urC3bT+L95A6spy02rBX0uOX9
BdMnV2qic4uxt50vKlVTEIntkoIC4ODw3cyKnsnSieYNv0+VW7izH0aSc8f8RjmUOV5LC0oU17wC
jj4agOQPBoKThc69u+NSr8S2hyLir6Mz5sa6HM8fxz3cRvPPkSBxjNUoffl6gRf7JtfkRDErr4m/
WII2iGIZDOVejaUphVlptW/Of2/INgditQyBOhVCosrpoMELaWEL+ES6P3c8EeUlXxGLAD+QPqzQ
5C6/t40Vluzv8sXu5iuQHVGkYLBb/QnhgxHOV6VV0TYTbejZDMyl1x+5AVTyWz0Hmo+2xJxMhXCf
IvyMEAD6cmSt3XfxV28r2WqqFoPBlJ+tLLkA47ushjKcI2crWoCprRR84/3AZimRAD2o8Rfe1gZw
T7Kxa3jxcpC/D4YX3ZoM/xl87vh6wKVnaEN700mCTnjKl3dMbTDSsoXezEcNymZdZvpvTMvQY/5G
8YAt+LZduVBeQNYaj1mDx39AFlj5TbjFr8BOk3rz4vEtJ7oZHMl3tLP8SAgkomjOuqEYYx2GARYb
S5JjW2FS+7YdRF1AE3gVnwmz7aS++dxn4LpCOXetx0o6a4Acmk/1oMRx1Xjhl4qV8cDnKiysO7AW
6j3vPA5KuBKAYeV1Tx0oG9WMqm/HOXdlw0m0ecZ5w1nCVuiL+Y8022/+bQVzHL2qkqnXtIuVeUu7
w4HBxyIs16VPPLpY2DqMkqkCmsnNW+bCzXpb9iy6yGJfOTgOf0T3OjWhHLTShhTyb5JaL3K9s/NU
dGBHiouAWs1A6POvo0p385fFGbyKA/vvrg0dGDECA0MIHrXHwvWZp7S9AOzMHBMw3IyOfOT0siIu
n+HCqj0bPxuulMoVEpt6ZERGHZBwwinVaomHx9rVCpTZR3kXHvBU49CWNrjaof2x0wU/ekekhAeE
RTP2n05I3zpUVOa3ftRKEULJOSn3HaVxvY0rZjtucCaX3hjdB6muHvDe+f3tMvmHpu7Ai+u49gY6
okMczEqEiL1Z9/aVZm1DB3mLl3uFEys67HM3xiaTFLIeECjVIR+nQ+8uOSQy98W8VtGhP24TayM0
Iu4GTw57BhxctajPfnIk1VKOdo+d9EPuSW/fDi6b63gfD31hA+oYOransIkXlrZxc1t1Mx9xzPfB
U3qSwb51P7Fs69zoTpLMaD1WuJbDDrsUcoCYsAW9x2LSl9DsFZeN3Z/47HyfsKePA1QAMwfgiuoo
B8M5UqGsjc827wEdfC79J4GYJvgIxfEHxdH/qA7ff1ydObMJAZIZfOASdpEVtcLkDuIdmP7HWbCp
xQtbtL/3VSXa7M7EoMQOdv7MK6PdY7x3oH2uTUXdOPq6tQ+57Tkjq39tWhoIy2okqqW+vA1qsnwF
Dfm+KUZ7B6f9DnjnhzNOu1g8DDdcGsi+W9smwQ8z44lTlAWUhO9m5fnHc5Lp1bhSIU/uFElYR9Y5
DmGwLGMaXONezBe0mmJwlOtKLRhpj4r8nPhc97bvkmKf6XINugeCXZbIrKzwjWbPp5yN1FPffJgT
au36Yh5+2q/PtYrsUG+TdqUAcQnWVGiiKWDAKyeBSDXSdsNkz70RsR43jEkxhTjV4xpGygfqkO7w
fNmedVKONtIRMzRM4A4m/iaQ726DRNh4U8UYKH2M1Z/srSkigFtv5GcMA6fgz54mn8buKIsVx5RN
eAKCIb3ARZ4rCT9p/kInT41cjbv/fdHJsHzOc6Gxv245NF6eaMFOmbwc5yAPBY9tNFXNqZhYInb8
hBLuFIzLmcNkfIkJvYa8kBKVQD1dGjR1NRj3LtNd0ETUOZA/iu0ItGL8og/DaJulcIIUSS/5vy00
Ur+WxBpSrEVqvQRcItwujTjxXtRrFbxAgxZSCZO2RYpyx5rBOHpq6v55NlFZSofmKuwrJZ1fpC5b
v7LsR6wFOfLCM5bAuCAmG4OYuj/u16B+BXMPOAABSieF0R6Gg36CQgPlcYMB0Zruc0ZgAlDZHBhS
vksddnIvnaB+llhxSP+Z6AwlZfyRIwLhQwKdEazg4nrTwQlBfDgVjayyDEvVuniQq3ub3PMswOZp
giFJSzwRUUJ/VeFXwf9M5X0S/m4iy01Is/wccf+FJ+CW6rWgahWDB5fHWxDi4bkxcRsJEFxZLW5A
EOpXBVGbv+s5nGef6dNRBIH7bSHnJQXVHcs328w870W2HTbfHjlJOK46rOClh6TUXEFwFTFxLA8U
zz8YABzXpi39BjQuhy45aBC/jMDVNyYacSsCBYJ5GkNoSPoTj16/ThMrZMRZeCsjig9ghvS5+LU6
jIxXYs2qEJl+qfN+gSc0dPLhVHmPzqSIz0+6jVtjlojQgls3vy/JkZlTsbVSBBiIpCRjNJHEkWL/
/KGwsnS7OcnkSaAmfZq9JdrOP0v9XDeoD5J6qHnetoQS9F+qiFjuDakg5oylpDHps91f7awDvF6O
fDCL4NyyJwSKZeCTfjCPftkMmwD8yWLQNQXd8Oy0SSNh+F5xcB5IKk4ksthe60fTrtvSjJDU2Ebt
WU9XcKHSdIMl1g9GOMPGZGP65qOOMTomtaPQwwpa4O4MTCO793di5NagPGcEmULl+EdoCs6G2BjJ
/WK9mqLNrBQQW5V6X4Cs9wfO8aPbCPEFRq6V3MCv6zobvPA3iZFmeF3lAMHtfP+2VUkuK+hSnRc/
shj1jUODDiR482KlnlfTVxeqy5mN7tgL4XtdO3zc4SseQDOmIkYjGzqvBEm/Bk5yRcdEoTI2NG6x
6NL4GnnAKvnKrGMK1If1rcisc+DgVt7RdK4l6FL3R+OdLbhBbiVfun8Cm3jnQEbC2cyiBbGE2CJi
dTWtA+Gtmg0ZPkiED0M2EloHoTEKbiuEDIxFs0eqO+q4e9lhD1ClfjKNybgui4wEFjmJObPelGGm
x4Qf1qF4ORr26qX2sAZeiz2Py2Ds3oLcr6dF91Gr7QcKU2wFORKAZV4sikmfcDElWTlOzpWC850y
8PqGkRJtt8KO8N1yMtScVIeab4o2BBtOljeYjcLHDrIvgk5gjcVG9a2m/DKSYYbZEG3ZKMqY1l2P
LOJPJ8cjtjS14kiiku2piuL6Jz3IvV9WxTIC7Y6Cw2t9roweSHkcIP2IjefqGdMy5riP/7/YOtDg
ymstoPL3DDCjW39jNaVwUm4JInDHTO+gppDndddEKt17a2SPTAmtUzQfyUG0pnLMqACyWDgZpHib
q51zddJY+vOdFrej6C1x3l5RWsYFwrUDJVzIURTMqBUuCc+nU0LRZHreAxZpIKf+avpCthjzS8Lo
Ak1j0YzQ1FuwiLNIsAhDb0Xc3nk68Q9Q5APtzzym7gpwks3va44dvPiPRlu58E4Xg57Nq58xBRuW
ctKOpnmAkeu40mvl1DkTAzA/FEV7ostuH/4tS9qgvxR530wu0hV6H39MlVGmUDQz/0kj1jYWp+6u
yxrgvpgNEvJFptJoPt7mkRWymRX+2zueNnkFIigBVsoFCtdHAqKbiHUCoJJeUKxIn14HGh5dOCZr
95UljLjkTOnGyOpYXbu5VpXvNfCT3GpZfozFZqf4mY+fbiYNF3P1DW6MNdHXR3mO/dNf/hnjBUOL
D7vOKJEFQNC7RNQxXkkgoMSRkjymB4VSAD1+6v2dkINROYQE84czfVbZfTGasdcka/SBicV6YhQx
ldRgYZv/I+3zbuFlBOqiFa/mfLvle9zwSYYHO1xOx6dna4uZIx1wAyOZjxZ7OLmzGHKbuecQrON/
449BEu9yxC/C6yvUeMCC6qgPt3wLsNVKmfX3oitYgNMXAgtZYjkFBNUnRuA+U+PIkUUecX4fbXbF
NytdSSvciv5rHYBZJeC8leW/wuKgUW0HhV4Km2Bjm0nunaZ8kCoYL+8sGpXeYyHtmEDqRn+zAmGQ
85Y57HfQDqy0YevWQLkdkLEhdN0RsWNvPJg09ZV/hMkpxa3oVBi/BduuRfKV6gtznVVzaHnv+Ar5
TmwemYa/38pR+shKb7FKtu0NKI0o4c/Fj9BPsBesr0+WVj8PMm6aOH9BvuhpXBMiHgitpsZnGzlc
6nkl1UQtx89X6NVS99St7jhiUmogvczJZZnbRbh1X8IhcRRzT95CkIE9ut/0JuL2IhZF3JC/AD+X
5e6X9u0A0aaV8NRkzLr7F4nAHFBT/yhCoDylZNclb6g0ywDNlh55SlxDBdlLoxV5nUHWvg9DXyP0
IOl4AaNy2Q5jixnQ6KAX4MFkrsa+ZDiP4OrmzSW2Dqe3AjrbzuVgxPAFHDBbPXGQf39wbEbpNFMN
CWidvB+OUrKY6HMPhE6csdheQdsNw+b+W9S9AUX5Wq+3d4Eqlw9eulknSqp5dZnDajPg3seJfCyz
nM3Mlwl21OlFL9az9wXC316dQqqnOU2ETs1dEWXWcu4IIBPHIPnzIwB669Y0gN0NI+zLIJUAceUM
TqroxUdzJSkNIXlqL2l4pozHjglcKLmh/Ly+H2Hqe50WBOx3Fqt0ckeVHz5nvOb4xFPdsaqEY8WM
m2n29I5r+6JT/m6hKWVQSPuEb/VVaQpuaP1oJRnyArbJbf3ThgPFNSgwk5QncRVi4ldmY5UT27AT
l2KIqbBwC3EE13VAkYLYbns7AQ9ZnNitln0w1GMHRSoGi63Z0f9BxHrhinGlJEZIatx5as+EnNnE
tjlvSrcUDVQUojVDTXI+kEaEIkA/5cNb+GjYmdlw/fzpkmM77bJB7jRIJ9CxhNEhofq/Mie7Pqas
NiuFCpoTyML0ZR10RuznDaxoOCjSOIz1utZuF58AZjTaHlT9v5gv0tXdwfP9pXMC3fFVtMM8016a
oFaL++uHiYXaexTX/0ybLUcdCRD0HnGuHvLzFb2jNPxsqiNQkxKweui104v+gFhjAWmlj2qpO/tK
yN2Z5SB9MUWjjc/5TMK2fudnz/kITHqd44irSuPhaT3Wh5i9CXep15oTO/I/I43gFhCkzILM5itk
by9aiNJJAA6Ur2xW6ZaMiaCmrdMhMqmJLfLf3C7fLLBSfitb4VMJqTo/3Z3dwOiOd4FVqAIoknzR
2ha7RYh42y1yYZrXb18id+HxCj/tNpWC4FTetCVRMQUgpYlbDXhAtVeWAY0eaCU1FH4nYx7LEH0Y
rlKYlEk2ByEsUL0fPzKawidZSrEjz7N5qX6FLYuhMYHbIe0AGqYtQRfA0VrLt/fbZVmQxHITKika
ObCRLVhcaRE1FubhCE1LCEG6kntuGmw13UzpXL4W+ofd5zUGgQiS7XqLU29fvoVELD0A5IO0mVw9
PxNVZpJ/hLgjiX7NiIqTGwYjj4Z9YyKV+UwUFZt4KiFCLu1GTppD8PXPpmJ4wlfxj8MzxPgFZi4X
q7K9mshxO9vEtoLMkPxkRo8JoSeSKeNiamlbxMzaCVKVVeAgu46munPIoIsATUXq2iP4TlNgdNxH
E0o9OrafC29ivjm+mTGdPYARoMfZHN3PMMMK/C2I7+Jzlr+oWR3Rl2n+pBQbyz0IzJ+X32kUHCl/
0i4+we0hbL/b1W3j5HBU4mXb/PGT72sGwv5N1nqfcs1NIHDdzisGwAayIf0PjoMvhsT099Jw0MoF
3y0mA5ciyXrNE4vgwE8miCu6/0R9H07NYqa8MOFTqURBFhbotv4zTThyH5RCZHKrZV0Jir/LF5x6
IHqDQvTziDn3bKfRP/USirqHbm451j0r5dv3AEfMCbwGLPn62IiREau2dfiA7xzQTG/F6h/fxFD9
Sk0Ml9ddGjbi7LSnCGGAmhRGFXqiYgsDSjDhd5abkhJCyFKC2X5E+JFKJb0WbFAF1TBbHvCFkj3y
7LzkkvAMGWGd9+D9ib21wAgxPmaae3zBQ8cq4rIa59xtyFGuVrAHR6BQE9RCyrv3qJSWPQAWihMR
58EhA75J2/ZNE4to0mDQi+3fe5pfaqnbPpc6IlBxzPzNCT1VuSsS2At1fFtdMPhgh16MVSk02L/u
+p3fpTbH11itGXHSaZEKGUnskImeo3thpdts54LzCPj4tlAdCs5DM4XHZ5O3qgQXC1AZhxGzG2Db
yr1S/ADB+7kDn1mrlFEMS7rta0TydzyWxRrT3vntMTUB6DzSJcom5vLlgURR0rdw069wcSY/F4hQ
6koQZDuCgXHdXB5ZIWdr/h4aRAhR9vDx3PWK8jvaIOSZB9qShzBzpMkhB1Tqgyi/A5rz9rYQ7XjY
rxfaSllrdtJEv7TtsB7fD1tqS2Q7RM/C0YQ+P2PCJlKtUsONkiv5NGUQRA/DZR/JcJcn3uo0QvkM
CGGpeRb5JCDv9/ROE56HIcBM8B1OCaYXpNPHMeAzRwtlFuinOUPKJcKBaybt6/DhnMyiCH1pirbj
J2pRnkBjg+JFWHzxJNpWupJuCt19gr6aRMbvXafWT+QGscK+/2a/KhgYPZ2zrZwr0VVubAx2LDZK
3T2Vk/l1nvL52G6iJ519gC3JmO/dHIP5eMJLP0HnQzOabpuRSIOmWKEFYaasJTfY2k7SV/ENDnDQ
/41pxrydWqJU0tWRqhJgpFHnXDH3W5oub2cFaAWbntyMHa+XSjFbUgTxnT3kDfozzeKI9Gli8lCy
QjYVp3hKRBWHoRSRccOLH4dUByCPhRWWA3CwYqCXIf+T5ajkUujIqnuSv3354psdFrurO9sioe8d
0oobrxm3ihfGQd7Qq0nRzVwHlKTtu/yo6/bMgXG/MlpuTINSixDrVM1RxPYafh6mx+HH6foYRWwq
Bhzy1nSr8YI/EDWaNRERsONfkg/yQkrg2Sg32iH/spKM93I+2h2Bc25ey0+czEmGICtxCZFULytu
tvHBkhg+lKyaC08vnh9ckScJphAwsia5OMCgJif6fjGNxK9BxcySyxvMRBphzndgQYmM93vk8Oy6
7iP2UL4p44l6qHlYm6aV+GFir25V56rwu06XYNnZ8SbFdL5RAjIMaIPPPMQ6eGay7UHOJ4BpwWXt
vOTjbHzwlAaf8Tut2b+mDpvU58BpCiSqG7IWts7aR7mKX0T0nypMx77JgIjtGtqiXt3ne2KfJ38i
h9eBETKfE1GKA/RDf21G+DtvC6OEpsdzRLgd+axhjedS53ftHJE5DGxqJ6EZ4DmabJY3EzQsimBj
d3ZBKa8qfb0s5BExKsz1oyKJKkxT3HAwQc5+dFj44q4U6jqW8iJH/gR9gpW0CfQmEKOExHHarfwd
oDX44F3H/DF0NQnZo+kyr5LWwoyM576b27iW9OjrodVkzuzQTq2jYSkO+r08JpQ+a7s5b5RYERWE
WngnPaoA7DHAheHqsYXq2L5EmuTxgi7kBtJfwURUA/CqynrwS95N0HXAiAJFbr1EYz8a2aJ7bD6b
v5plk7fHgeJ0namcmWv1SzEJrtgZZfgbK06TN58gtpTOwDocpy+gGmEfp3P0z+I0e7FXzRXYZ60C
fQq7/3AbugxR6CfNSUHHwT77Y5KGqBMvmqilvL5UleIqYAYGsbOoHF9pwYEjQoK/+XeUjRYImwHj
u6tMR6fqeNK6Vmg1Xh0niBUoQSz4rXv9V2+9UztKGCPlVOAdYXzvHM32LOQ0Xi35b6O9+e73PhXn
ZALz4eJE67jBPO+/my38HaXFPfsp+HazSxvTwv0pXj/bOB+OliJqHzFcvn1b4nik29Rn4UuZE2SD
8NcLZq84Ty58X4tAJVjrc13UnlXofJcg4D0gNyZxMn6RmYgUsLY8/SAhbKZmrD4pUCHVWZsNW8p7
jFTX1vXmVEmMifcqx4840rA/vwzmIY17mezk9i8iYtoScQ7S2YlUe98YyaEGnja0KUTk8zCyFPz5
ANOMpNVhiAyjORirox/2P0N73Kq06cxkI25LYR70Xq50O5OHm3qEEpI/FG9cKzBOw+LTViB1VO2Y
o2KbV5YOp3wwiqU3TEcWG5Nqam96QSpDWEX2b7xJFPuvp2Kw3J1JEwZ2LpHTyqcasmWvWxd3Lywi
n/qaSZZ5zQ6hXcQEK7r0NbOY/zuVyFLDhxYuyMXzM8UAD8dVvU+iVpIP1j2AmbwmqnOpJq3yRP6P
MYZg+BvVbgG1dDLKRQOBtFW+UVyzPhco+XgxFQiIN/pBckmS3WS9m9op9CeT/H+rDu8wq/3sF99i
FydEIAHaEY2sS/cBT/VZy1MG5G9Jl3xOJIDxV5MZjpJq0lBxjybo164qQb1iXb2acOeETDBJX9wx
89tBR+YMdZKWrqVRxn5rpuDsXWwKnj2rbvJUB3ikHp80HQLTQMGotxdKBmtLn/nKec5/DN8gg1CF
tL1zrNvTZz6gwRMMWGs/1MoYShMpP9UeRDnsgMI4c6UGAeTX6YiyEAhGH+HeziI01QjNtsP/jlC3
7wi4CAjK5guP8ajSt34aOfHzxe+CJ5cl8aJq37rFvLfSecvljd6xOriDTYrKsmon7wPSpxHPDDpK
5b6ufbOvuhKEQIl48g26UL72xpdQPD8BYEX++7poOrau6TBeOxpUN1VAU1c0JDWrQe6eSD8GJAG8
uM8CRg9uryyUlvM/W5Cx1DPytbkAROjh4XMDfLr86HcCPRti1GJWLOhwPZePD5/zGdY+KN/3QRr2
x0cj8UflRWmL0WG9KEJQSkFUHeTH08BIvwd7NVRSQXDlTbDALAXg8WBAP87nU7ZuWJbzRRJ0/dez
BoNjOYdvAV5Pjp3arVtlFjtqLa+YDGlmZrQ3MBx7WG/v+1WbrCJtrcmnGKMlEK49EF5h+VrhnZ3I
Cqv9zzflTgwfnD9g/0NP8d7QE4nsLtVHQIl63KLalduFbq2H/LwPCMiZLhOU39NlKuSRq1XqH0Wo
ix1pviK5Cdz3i9K/aIomd63+bbrFSaFj/qEqWSR5E7j8VJimapZkLDs28nyCGIQTKIjEfvUSU6VB
+vuNe0ajpYzOZOXAKzbK4t2cloVpm2O+PsXUUfd54DwJZkvvC2t5K7Qb/P+JJSm4TOxXhaYLmsRj
DSYY7v5ymUKHUhjqd1QYZ6kZyxjVkE5Sjs2h03LhGQxTzSxMfTEdlyILVVBrw85WpgFmeaFx6U0Q
OsVr5Ha2np+3uIAd/hsyYBJd0v1YBykL/usQUs3sYTCWn0/yGk/b8fzWtIKK2V2qJoKb+WyMU9G/
7uciJeedAjHLi23wFzo0ClBTjPTe+Ukr+bXQ9bie+YRdYCnsSvqlnhLqrWkyPz612NHwoj3VA0JK
G2guiK6vy0gUip6jtkIr+3sr5t8f90gjw4XetmxjTKp52TtKZsFJtnBmgqKZziMZMUl8SL35taCy
ixWfb687mwu8OWFTIexRKBbvBaXAQpa/RD5zJ/Cmt5OPtF/vqvfdHovzXygwAs+U44tD4hLC9mam
oPtZ9botWzTneSC3AHijIuzcZbg9kWVd1gyWZJHN9nVk27Wzly2IfDQ/YvvlR2IYae3ecicKrxqH
bOpABTYOS1IOgELrResajhgvmYGm+uOesUSiNwkHVn4af81oaAT1jPhvhebYXcIRUhjydOPS6YTs
YIKjwJ5mVRAqPvHNRNxHmwhEhM84ZXoI7WrbjFiLGOv1aJzjF3TcYQwcv7AhkjuOLXdP2PwNlj3o
7DKI4p5vsbpb4IZkY/1RQRaaghm8KPsGygLLxQd8dpbaDERV2WuSFAJdfOsSMbeYyIb5/a0Etp/B
mtEpBxqHJc8dT+JQNBgGzBd7foMRyEKo3o75DyrI4YnBDtIErKBNYT9NUpJErolnFAE+dkTOu1NP
KNZNgX4ENuRXl+YAFtXyJvzAWtR2Tt38dRcqttIJyMh7jYZNlYnTEyoiHRmcM6yOOHAs7IdRkMVE
IcAmmrEuB2/p3x94Ur27qyihgklMiYN3K5aIamdDxsPq8unHJOUzHkOBFRGuQpf17uW62dfbWKs8
9smTAVprnzK6DJTleMIGO/U27GCIzzsJxSkZ+gycAPrV5fUVo9YEuaUH8RSGX22fA+FLvnhaaxgx
uS4YU1mCy3N8AGgUpRvQ3bt1YADds95Z8uLHHNN10r5Rs3crkfVLR72gVokg94TneFIgDZ2rEni8
n4LZufFdulhYRQ9f0I8K23hM2gsE9SDu9qAmLyNZmwjhRK9vhvX0TxOYQT8jP2ZU317WEe71gTuG
5aytQOcQrerPDUPt/091qxQJFA9HcfAWmqxUYBxuPYHtYFqkViayQXL/sj3OGB7KZCdhknumdEJW
PMLevkjinBK59XvDU7OD4QhHj22Pz0rMmOp4Xd3YKo8ootdEvYxV3pNJAuGzUe9QefK419pfY9S0
Hvu5x1WqubSaKfvRc8mQ5yi1EbJRt1Yz3KxhTLiQTJ4VfjDANvSuG22F/epd5z76tBQIJgQcJpyK
31izU/nvTJHWbSpgeDC1bBgtxMVWv3dLwRscmxVZ4TEsJqgP+UAwEqBoyw110oxZA5uJyJXyTsIb
yIEre3CUYWLO2EiXJBHrygrKs4w4j9lcWKCme91TTzZCu5Xv3l6uIKFTmX+S1pPWvo5AgVi9+c2U
ku2d+hfxFg8TCFwwTjXDVoE0z+uPpxRxnbG2/AtuFmAR3ZFEnuoqpS4evEwCpr3G4IHuy9LHxF/N
AJtLfUb6eceTIryMToUShHwh0Cvb/L2hp9JOuTujHkCME9+W1l1Pm0IA2Wb+2P/AW8v8C/EQvhVu
/v4FNqKBeumSz0ODk5Wqj0VZhG/43UAPWuA0bDgULMXWoATVDMuBq0KCzLQjzv2KmxG8yknKS4mE
hSw0T7pLMCrcfHAoXSMTmwbmLFQQsMnmqXt4q+Hsgzw3PiutnT9wryZjLgMcvX8zT4ZUvdotr/xd
EceLUcNAxXEo9iw8K+gutiAUiTeJ6jnM7EJAKBOEmZlPqOVXgvR6fIhSJA8oRDGSUviLR71uao51
M4kl2Kp7yKdfLLXOmmKE255r4oz8oXrVxs+l9GZ6riV+4WgBEvycsCc8kfRtj019PKgF4sTAGoLx
NUZPPb6K4rVHxC1H4F0U4Jifdr+nWTKuYnXsuCWrdZYcw4E/Ie1z4PUnTeJdvQ8xegVm9xwcKqNf
y/8SgV/TZMnEGp2lAzm9tjJPmTCoKfvY79lS360/yPb9s70/fQptD/Og6+s4RYNfC3DoMoNt05XF
RwPNL9khoq7RvX9xuSVgkle6lZ63cMxg99GCAJgXuMenjV6/nAjv3MhUAC+yCwNWeK+w4uaJdXKq
yMtZLtCffbjmq9tuhxJstfyqHnOEJdETyxJnjojxth4ZEomVx0Fz645LLR2dPB7vKxBgoAMWK9MF
grty7v0UGBc7BP7LwM/Cu9T1CmwRDfSZXeZ3PsKmT2M8NTwxzLw7VSJ89iNDKoX7h1C8j0Jg5lxj
tBZWoclt9SOqhJ+0LJeTGes5UYFPueKp3LuyjSl6rhMVIDznN7wJghOuc/9XBWaxxB12v/pQw3jE
LK/IGaEIMvf2SV9FtLR3Csz+J98qXpdDj6h0Il+Q2jfJZDDanLcHRA4Wdj9DfQWhvZuOogaltalj
uKGmiHnobe4rJj6GDkn3nWmYfJUg6/GUXNvQbjIGOLBqkpct6exUKueJlBPac7iJwkJjDDWsAu+O
eBekTso0cTlgibpevBDvTl4qJb/rjiCQbtatgWRmCJqufiP24d6326TiOriB/Uii3xXwYLfClZ0P
YZLpxhueAn92liY6DRPsPYgbbG0Y45g91DSQBflWMf/v42GVcaaeEyW1UdiLLYbd7d8WJi6iHSy5
HJ1FybtXQdcuBlhyIhhSSG1wW+eUl51oAxA//PkEXIVfU/JlHHoDjOgZtdiwK4F06ZvDl0mKLGxA
/s1fGrFR4EkbWM8dk3mXkQvBdDSsziKPgDwGF2vT2i+UtY6C9kXOMpbZqcZ8DTlaWK44WrooRW8c
1ih85ieZsKj2vk5DUk5gIGooaZIyJiCh+aUUOUpE3OiRWp6ROCdbjXj9e0IUTQyRe+fTO9JRWNxv
m+Jj8EKCvjeSyhvvNON3o/W2MFA8fUNg168JYjFW2kqlT4KC7CVClsJvhQZ2zsMz9rlG6Zr6AyW+
rpU7nAMEXZgZS8g9vDx0LYg8y9hdDXttO577Gtk4XKyszXBw4LnZZDjdPI5rTGYMG2SKsgi1ak2E
ywOMFeFm0c8lm4KmkVfkndhzm8+mMNLGRXNhG5f1YwhYa2lG34uapX035FCewPUCeuziBEcMxE8v
49OFhkYlABB/xCyeTme2RGCCU+Y6m+800KIsWmkKG4d0k/sNMG+uooBGWl0e/vD417spYPA3htO3
uOT0r/XfbNezHwYV8I5XtODCWGoLnt7Eucpr8c7nidOyXfq6qoFdY92ZEW3J4F94NQxSpgwwPeFe
3JOwdihx/9qa6Q7EJ3YPFdxRi3FrvpvN6PXv5MVMOSr6aZE6Ls5/x3yIDKm0dCGLRt43Py2iC5Ij
XkpkrV2im0NF0assYZaYdSVEruq3NKxHltsgJIXgfIJ1ZxKuGzzZMfeV5g5R5MQhpl2NJ6j4oXGA
jNDkQRuIckrC/8+WE0MhcxlI0peP/tKqUvLIBRDp4qJWBbL1VzEbhiTe99hm1+kHFhmTk+h0FmBV
gegPrQzH3Lx4BzlGzWdPDbOVfkXOpqdVhvClZyl7n1fSXwQvks/LxC/WokDpBM+rx7jilWpciWdQ
sw8tgjZdazbo+dkMOD1fiA58muqp1u5BYSA/3p3sMbhaWA+XtG1DzgexVDvbzVd0uy7wLu8ZvF03
7pnJqFxiPxHGhgg9c4N+AuAKQfXIn6W3GAIGGFRrizDPyn/3B/0Dnxsl7l2QCrCLaw4/NR3y4115
EltEM78ZwR9xzFZJJaq7z40PCQ9edorKor1uX2tiFgkLXE2w7JjyVWSC52fA7RtCT4g5QfyG+pJR
GOQvLLQZLjMw5bdQJYn1FxJSr0IO916LHgS55V8yMBFA/PsPWXbcttF/yFSXGOVrjWs43HgbB+Sz
5wclvtYzA71SQUhVv0b64Jm/PTKjvs2ZdYNYzJX6Rmh+4WoXfBL6emEl9d3JZB5xC2XQda9KR9Nt
oAnJ1fGPA0APTh+w8Mwx0mp3/789DCAGAUPxtffKZeadlGzfcTDdS/o49ywgagpKGUqLCrUNffC6
jjCp9B6hl3pWuazXpPfiWepi+e9p2J4ZhDgJfsuvu9zzDdSWdIyQplbikyXJ4E18TaUlMU6HSSgq
c888ra8v3K7N7UdpD3+eKbjBviSXx26ZlIOXh/4sowSoEcTqL2cDpbxcXBsYEtm6dL6D2tUojb7r
2sQ89PeVQkP4/YGU/U3stHQzaCSHjCXGieSWkHnn/e8M1fefLAhKjjYorMDWNjKInSQHt/C1K79m
vTZqNBQFz0n7EtBB3Tj/lB4/FK1UUNA3Re+Z+RiTSGy8bgW9zTaZ2N5HxY5fBeIrfjWQq7Q9jAxP
4BwHBGQezcNc+C8wdAYzCIrb6rDBEGGCmt2mcsr6WGFBVYH79t3kClE91cRgYJb4znZKzgOszzi2
4v/L0f9KaqANpUhMta2de2r5SpKRWXhZb+hgwzrrgsUwhoabxXXAE82VvWVReBuk626r98knCVSd
fyXfUrOZ64gmBKfqEERcqebgOO0pzxn8THLXzz9vw07DFgJezEH1DbPwg2JNGg6aRAwpxTr3Scq3
eA9TlYOEKdPZFjIQrjEBP67PeIHGSfnXkRMzZMnhBOYkdTP9pQhiOGgun1QGXjG6joaI+8N9W/Bw
kqSi0a3Kw/mu7h0sbQoi+PBISx+/aYyuYdbFmzv5tomk9WWL4y+SNyPLLKsQfmgr82f18NsrvkAQ
fAiTUepUv71Hh4E4rYeF1+E5Xhxa0zSJ1TJTyGzmqh/Tol18OrZW9U7QCPz2d2rJ0d+K6ghEy010
CJnLBgo2B0Y6zc7RyC/6RlKCuYp13uKp4JG2M3F43UACOnZuQeskSp3xR2C+muUk4g6vjTyMdtdW
UjIYyIhQ/ddz9WiB6i1yfK6wWPPVVicwv0qMfCs7XArdq9aW9doGnaBzEwsjXkzyxFfrAE7nxja1
c8TQfn3xu55vfdCKGd4ugGOV8qEkEmYg825oWfhQVIy71KntpGeM2w65SdjH8JcfyNJgTvpGHt5i
GRu5P3EMTrbfqVZwtI4e03BYwFbXsnszx4OOAkGBYFDnSMFXTxZTI6RjF/C6c7jb49LkLlGfgD2m
V4X+2pj05IpeS6ByZih3xRfHA4roIWDj6ygqVyZ+OwcjyQxd/JefZ78s8jmyue7klmwkrhuynmDO
UgIzFPjW1W1N9fviF3sWju4mmOxziZ2ebk4MBksa2btTJmZmxYyrHPbXrjTWfIo6s/jexQkRUfNj
DD1XnVVgAscCLtk4QaDwQ1nC84NxnzGSOQttgWwY90RzMBHy0muBBl5FbyCifwGRHc1qwzTh1JsL
tDSimuavMQAoHOFeUcLooddlk98ZQNeUWtsddCWZxmdIghwAQarhyp9y4Iz/w8lTxsBWWPGX13Va
g07ZVazZweIruZdThq1Tv3W7BBbSYAqPImzY43uKEGaFrmOQmsB0mxDu4Pk0pD8/dfYDR6qhGtQL
Ve8Qrl8jhkrka6DjcvRkafGh99bz+x6agM3XVcWRWUEMeWrPgeRRCalJrFqTncM5/bGlFMY07/mE
XFkXFQS+kj0zxOz2I1/qrplmNIQYfbQsyTyIf7Udkz0b8twJiMgsQsHNI0NA3ThtlZ3SoIYRlKLj
cVa3s/kISLGX0X6ewdQIsLK6RI0d/r24RqSP8qxuGb8P3ZW/51zkUvmuIccHC81oeUyXMRzDjJbQ
yyPYT1+I1Q4czMjjyCaKzzXcONECUnfmUaYPUPqCN8r3kBKI00VXD/itFEwyPHDrRvPvSl4M0XuX
SClw1OAbGQTIkuiCmCjz1ZzKeF2bTwxfWsTwwUTnlKlvpiNqXZCTZ1XIKfWCoRyi/4FDrxa49W7Z
NF6dNkrm/kAv3CJQhexWq1cl5oT2tkG/xGixz/4NVh0yvN/G2rF9VNWZd+8/xNRH9KXLaZFi1Lra
Gx7eW0RQ8cIf18HXdFlyRABcGFA/l6H4AUnUmQx9qzGtEe3OOMv/fOFMOtGzbW5T1TZWNNReaCmc
WEh4fxLgYHpEWJIaUj3TvU5+FZTlPldNaT1C6DRQ87vPtZueBbUI3aBOCY2FVraECKVWUcSvAIcl
Wg6VCAqXyFInW7w/osuA79vP5+UglqzK0h9w0zIAmXf6EeAMzClaRvKOLfPhEKpLgpqCDtCLou+q
5doRltZ2qAYljTLXltxyBfNjxfjKnvs0urvOz2R3bBMCpmJYFgfyrpE1bSxt8gSv+D+dqBS0g88u
18gSths7MpS1TAzT4sAWzLtcJANMHIAqP1mBOAhE+gFRhUsOzkOg+29oR2LI2LrvuguRUqYr2Vey
xiq+4485I25YOF1qKFgP8xLGQ6asYUvzxAXxaEvI6ngx0u/x6juDsEqdcMlfYWFmz9aJkTt7zqLP
RSYWp7kUl9engCo5mVJQ9TtV5WP9MnVYQFqpGelSoOtybYofDYbsTCNiV0oxOX5nbM3dDUgX4tca
zK3ntuS0IpeZmR3wtVUo/IwJQEsmbdjCkqcwfQ4aVfjW2HI17ER3h6CsWA+e/60smA0+Q76yAbc/
5YrWp8rz05DAEiBbie6QVFAORos7ij5LfwY1OC7Z1uqpCD5qpFMGcL09azH84ycJ5ndywteEwud8
HzIpBhWy7IH8GrJYjZQltGcf763tvnWi7wC7PoD8Nfkuv6keotELg3+yRGevbRgMR70ccN7GSOE6
ctQrdexwh6/aRMzf8evEe4p8HQxilIF/CsS5ZdIpVqvjoDfHqsGrUREiNWlcTCitb1HHF1EckHQQ
+i0rjwMnglcDuhEU8QkUpBEC7E6Cb2iBsNI3wnO+joF+CwsSf6ppjLpZb9RlobddZrCcxvEuGR6J
fcWhXUm2rvIEoyonq5JAy1ztv9KIoapP+WxzmTpuxdB3rvU1jVp7Hhg1xnmv2G2dIxXColD9jbpG
MUbJLMVr+XkJqN3yLFTaRMs8ppYnBF86uzJxdPHpCvvmqpnvbHHgyBzJXOwYkS7b1emPnFinW2mH
mlRrO7OgU8ToL/ojbrT+s56l26/iScYxvSww6hxAuA4Gjoa/OYSVvixwEKxHzwjcdLMYjur8Xl61
ik9Ih1C0wTu6QTkaaBC+nrgkudfPdyvbAhE7GdMdMzJOKhqAkRem7dbpGHfA8oPtwsLjbljsb8LA
RTkdt0KvF8oMg45Ec3YzT0Qc10s3e2AA5VWuSwZ5zR686yK3wXkJbI1QhSm60e/9NTx/roey/hZf
BgbRjpMhmazp8T9Y8K9YjURCBc7mMQLTBCSqhrWFkT5yjlR+TaYicHlqoaOFR6u/vISVQucu/njf
tk8T5Yv8gnwyIe3OX1cNb/diRay9WcUK3wniMQMne5MeH7ku738cSxBZKJsc8JSwm6UnFoIqw816
ABdQ3FRrop1ppoo7KyON0ZrDnaX+nYYgKhaoyg3kPPWAZPOkimGC0aj7O6b/a+z3ryYS44RTWxS7
5ppouKVhV/78tu1KAmFqv+m0AFlTjLofPoQZMll0r1GoNym8Bf0Tf4hv1TIq+zS/kn5Zt4fNX4cr
ZCgS1coMI8xVLIesUwDsZKdzba4y9VCGHpwxhTRaug9QNHK4bWKXTqa6RLAHeRoM6lwASH3cNdmp
urCg0XyJrK7bbu7t7eR2DEJ9vBynFERg/72qPMB9UxrbXRasZecDitebxArogSQ9YhLs/z2Yk3id
yxiLHOvnmo1L/eubKPI5m1obDKfunRg9c67gzffSH7YWbTojY8wkl+kXiWLtyumnheoSp7LmRezj
uXiIK5NgnahaPmY5uCks7A4TFxsIjC2FMciHZ1QdgZjeM0Gga+nET89qRA7UllBdtc6WuXgTdiaw
/qad7ZxKbUC4nZt2hr4PYkpZ1hpujKNOkqpqG6KFJ7h7VYndjA6gjSYYT40dgUN0vJ2aiwYziXuZ
OLEIdT7SCxavKvsrK5ebiiC/INWPk2LzmK9H67XZ7jv9jjTjO0xBnrXgMbKAMNBvNjQ1mRgcsDSt
kUQhrWwvAk4weHz66jFYj6ZPFZZ2vGOGcEjLbGYVDW3aRrUgAEdCoR+tXeNyHvY4IchrDCLOno9L
HjTq3+saWj5sAujO70ChYf5lZr07nrZIDIFsbcW0ODMNIpzQFncToghuSCFvK5EoctS9D7ohFMZe
HuanzzoFsFvRuFofB1JPnL/398mG4MM9/WRgF7CdrhGgfwx3Kap8R4QQWpisSt9tQ5tMq60B3VME
EvbvIZVoT6Evd3G1hLv0rErd3pGZ3LzBTF47qd4TUB7/AJJ0NtWEgSo+ekzb2+Xlr/uWekz0AVaZ
iLtHlil1O206KvwvSwIdH7WWGLcWAefZQ9VVXy3FgdYt3CN9x2/Nyd19TuTjcQMepB3OlSR4C2Vl
vgyG/38+IAWOge/l/fimzzXMkw5FIHgzOr9TvqZuOhjRgIoTUAXddBuapo6dNmMhpvKxuK+OPir/
Z/pE6I8tnxSSJ0+zthdusAgMKsz/tlxQbGgTF9sNGh2bny467ZFF/2lkapGy+6LvD8AFvUDymeNZ
A1EoxIpHaDEfwleJNyWPoZTWh+cbNWQqkci8pRB2ldgz554cmcIxCecyu2+eV+PpzcqIFST1zvFf
tZHG+YIvHsNgi+r4HhwVp+PW1M8lxigO88q04JqTK7PwVXN/1U+yyCgN8QQtYmxB17F8mWVA6yUG
aedRhWfq6xVLu1ZrL9rtNBhL9O/CV4sTYjaKvYiSqhsE1QuLPajAsOVnNFlUKclU+zSWvc7ItdyS
O4fsd2g8T88cOGl3cmqgH2pIwx8EtQixvRERDlvYGoLzmyZU36OLuoEN6jZc1a/mn1WgeyoIIiwb
2QnvmGtSzQeCvrC0qNn64DnApyZLnm/gz5iTvOJp1c61H0UKfYxkyKgdl1sjFFp2Zw7RpxjhfvEV
saOMxvAOsEFEHFX+6RKsbseZP8Reou9X7Zpb7EGUPVYu3hR5vDDOkREWyVyebrL4v679ko9ZIiDC
qNXPslsoJyiktrScoyk7euvtZWsqOCgvl5Jttbjk5WrwDX3X/vlpfK+7EUtcsHtrw2WvG3lAZbNC
KFmGVxdrYRU2jq3dx4PqCq0SBbdpyl7N/0fgSX6hck/LQvnMcI6FgLCupbVzOa0wHPFG1tFBc6/Z
EvyRB86Uo8HuMNQCxUEwHjadqRCl4cm6Dg00fg5iExGHfm0vAXQ06UVsRg/ey5/JZP2Aoj4h56IE
aNN12gHE94lCqvVscryjPoPEioilLJHJoP3OwysIyeS5awoa/NZ3ymBaTQG9mNZSQuoBzyjf6oEr
Ye3ZaqoPgpaGx3STncgu8y/eNnmyYI4hqeph/5YgTR3qDgOW63Z6mqlho7rm8JFO7lFs8HTIzWvS
fNoN68jiKeW5FORt4eUNpy1X6lnzLfUM8t+PH+pJUmqq8RUVzWgVKqnjPXssbOgBCgSUPCyVJ+Sb
/27d0BynAPFT5JP+5Igd55CZ/QK53MuPVbWoPMKn7lOU3ESPbOv+zPQwBeDMZM5Opmv1vSIFC2/0
+EjdosOx5rl5hrD+IRO7Epk/WDWGE5quF0OkVrIqhFbNOS1zTWYhbdRP4ll2lt9SS1A3SA+tzljq
j/d939xWMcKBoTWivht3vRjae7prpTQbj/WqRU6lKFl+3gvQu1jkceCrt3chyAs74DEP7uEElVTJ
chOi7omdV9Qnbs8vXYRgvnv2MILuDMVBJNQh02k25yt0OG+fkT4ZWpD/pE4RfO5EiKNMRIY2vuKk
aF1pvVO4HkJe53c1zLlvvYIEdZQyFhR1p9SFQXf8Ui9QwL4UJ7h+LTZMEr2aN7gwmCChKBezWjuk
mtNB5kbOtvpPHKs97lLDptFcHAzSlTEPHz9ftPzpUBXWw+1gCfQXvnRr6dMpT12g4XTv0rOqjyK5
rZzFnRjaJe8A1BDwtirJWyIkR5CBQjA0Ixc+V91XzTCJxr01vvlFa8U5k1V37sKexDSs72A9BslP
M5nWQJxYcL5iprHbgo9Td2Ay6JmLLDb9Laxm2Zf62NKNRSr9r33ihaDmBRdacZ99nyV1bBEav6DZ
To25giALY0unK61uKd+7Tc7LYE5+pBHFiyrs/qgO5ugGLrTNIY7JuKEQwv2lED8kkHf+q2IWDcx1
xZisemFqwBFZSN3pbYrbsh0V2LE4aZy9/EgO2JAIZl82LqtG7c4ZkAP9iFctq0/TVu9Z27WFMFro
9BfOTcg3+GoyxFhfuKbL4TeuD1nMX6bQy3rUYzUYwLpQ47ICe//aV48Al12RYlXVTl4lcsjCQZhd
IZ5GJT7DXvAdmefVmfVIWlHJB1kzaeGVvaLiiwaicZYIOFgRXenOW7JRiQ9S7VUco7VPohMqereG
jKUODYnhx1iIb7o/7g+7Qb/1txoeleVPgOM/79Y5mvA7+6wD6klA8qlRHb08jRD1lfFSsEwyqlQx
DQOtq5tvnAapPMqR6iMfwyL6hEbVr0YxOE1tOnj26Q3SLYZMx/SgQzG/V2OwTzcU46jjAhzIEnCh
g+WDUWZ2Dz9GTcUoEDPRVGe61XGmRMALEhNtGzXRemC+Co9XEYiPHFHRZN/vbbYE+zOZHWkzFHu5
szJ+i5hJ/wZWIK5dRNdpDcJVFPltNQVYCZbH4aagkkRTViqEILJxbnVpvMzXCp/AyDgJmg+GBqTb
rp9sZ98wsDvx8HvE9iUN9zCjx8tVGHqO+8ci84zQWI+LsefD8ERtZa17k9O8IgfnELWu4Z6+yvfI
pnBu6Pyhu9bF93n21uQS/zfvjy7AXZoKzO4/mgcWO5LoYDiFRoDjdAw0a7qaxt52VP7NYq5hj0xO
qzfdTAqOZ4TtfOmeaLT4uQxuR4PDvPsnVa+GZxlaWuOY9mdp0DimhgqOJVs3i5dsnjR2Qm8faMNl
CPXDtAjUHIRuVPxr0S6gKx77JHihWj+8zytu6FY1LH/ccRdYXpNh+YRmHCPKh37nQbzmWyAozm0+
I3/QLg5y+qUVt0f1Fj1wVIRmu88qiAmDTa7hUuhkYFonkCenMR3CTcCf0EwlFYEpQKTtLRBjziY1
9YeFTmS02tUEyadXuhr8aMh92OSb9tp6cHdIvEVCGE3+IN642KqWYmRS4Lp9QtwRJC68epTeVe4w
YXGe7iXlYWwVbAPVh5/a880+cRM/TiTApGPt3jNB5YA8QITzN9Thl7KaoOI+HxZYrSQx3VbVRv33
KJeA6zrF5GFh00y/sxSTzU+BVYt0/g757AkRiWXAXLXQrtI9ENSsDdwaodbtjIqy1vNKuibBmyLk
k/K2DM1XxnIxyoG2o3XO2XBQuxe6XQtwQcG0Di1VzzVWtLrGdZHfrKP9W+cub53AHg2tNBvGra35
tJvQnkreEpop5Z11jsN0cT2wvY+Ytc3lThzSz+lKe5reITHiEwkQiYSABzNQlD6RTKrxkvsHCED6
T5l1i6YHvr9Eqm/IYKGX9pfGWgKMo31D6paAwm9srHDv0twh2lkaLkRoJzOXUnBZCjJb5SrNVVeV
N6piFzW0nKjTQ5Ui7SQZhZqEggoNQSJJ0MdrnynZmU2iTH3djV3OyQIHdHa5xkvo4ucOiYjV/h6e
K28rX3D5GkjG3d35jdq8/3NmJinqvgi6X+Cpq2lzgbIjQhz8lSQ3o9NWkwce2CpirJTH2L15WJbY
+Tp+ITS78GQ0UZX/R78LgCEGqyQcCbEnpixQzM1ZwpSX25pgoC/oNzCu1bm2Enp9JHQsqmlK3Rr5
1VhU+8Lwhdb0N6Xq3fKZpDVmH3sIV6T4IEA4q+3waCQizm5q4yDJoRLpXZzZERzJuCkdCLUt6TkH
44JbsEI9gJdc+C34xHwttCV9GMSwBBKdj4bh8dPNkpX4AyngTGMOMiVmBKQoVmH6HrYNP6pcWMtw
gAt7Xx4r2Vk9Z7teCax2NMVoEuKifqx5r+FyRIEHwM679f8OwCM8FeEewH3+hwVnRVt75if9kLu2
wvi+59nySBeQuZ4EfZWVJurBHtJ4h8w0trbUQ40JUH2qYRyS8L/QnofAeBUAFL75eDqCedpa1fYn
BQNYP1ZxM5+tzlo2LA7clnd0sSCkxSFlbzt0UunAr8+WvShe3lC341kexcJBWq1x+t/bukmOS21H
DFezERYE5oI29rdOkV7E6PTGLE2hloCcHSvrt9SPEKUfTQdYl/PEQhCxrHDpPGALNQXF/uyx6eTW
1fDLjBui1OVhcupc3xiZDIVgLv1wxYEmb4Cgd+PnAYBi3cY/Y4f8c0tedg6yMJXKHNxmbaZ303aQ
71n4qbhYvCRJ7aRSqZjwqGuAOZ16BJHfzN7jXFV/KHZqLlTiqFkpJG/Z4172aiFOmxGjYbp3xsoa
zMFhtQmUyX3ZD0CcT3Q9zN75rdw02iz707dARJc/MhGW/pjAnOEdRmNnGdtkfpgo7zawy+7wmFty
jPhC61+bPR7ezgnj73gR505dpA4zzjetgQGxFzt9A7I2Wabn3BFjfLLXMfYJbtK5tKYuwBLSQJ65
kl6THn8e0ZRV8vcjxPnZYC5aldCuLVp3deH/jkr0cKpHucVDopS7sIFxnH2LP3dxoYDEIyftUGo+
Ds1dI0FINnAuESK7JpVm9PnQkUHQsXIYY6E42lLFBoOEFnDlfUR0lgGoUS1PC5++omqlKkrBLlhR
dSF4NCekDnj+Dwg+6Bzax8BrTXudRXQXeJz85I78HCpM00H3ZNtOiBism5aj9X7zWsERKb0qttPr
yeosvvTjKmmp4xfJQgWoT2Gh5Q7nibWPunHB+llPuQO0/1g7AmkNOOBvhGXZyQLyc5J0rHF0yLNu
Wo0dhH10K76/I0DHYZ89gc50hW2p23+OAGQhRAG0nM2ndGzPEE0v/eemcpy+L0OVg3vfTKDKgC+S
sG8gsDR8LoL/NBcEoKcrexD8bW+JVFP7vzt1K9OMj4Ewtw9hsIjgKExrbu/uSdtdCrCmxzcydkq3
5g6bPeJj9uVw+pyRZFgZaLL//mY6g3HxpcCZQl6EVSdAK6lEzUvL339WvueDQPak2aqrEHVZi1sg
6L92RWwFkaklf06kM1Mzdu8GGfpEnPhGvEwnxL7kiP++mH36Wt6QZXiv53yCU5UwSLdDIS4Z8KmO
TU3v0DkH0BdRjubdtdNUnnDBA8ReY1tsKD8CfrIo/a+N2s7L4sop2W19EFleHJMKyxZXogsahU4e
pOZsrY+jaPIwUJ0zFuVPxOYLC0t3LhZ+xNrV5NjxMTVrPa1C/mjTVKUOqz7jA7WiPQXlItoAGkzL
6d220JtWri/PC773vvEM11agJzj91HdaWGv7tZ7H0ND9lQ12iszrIdI+BG7/OpZGnnRdGA9mdRHm
OY/xsZCEOg07Tp6s7hWn0N2uc2kkLwfEJKSTjN8XImO4kiFqR69TMTKi2LwdajPMlDIngnwOthRD
zPBWJAVoucXQTU8sjijxfa6GAKy7syFLXxSojEH9p7Ed7t473QS2WcQCCfIeQVs6SyWg8npjcAVl
zsCl+xn5iLsp7FDhSo1yapYp2KCZ37m3PpYa3j9L07uCfBFRvpVSsl/a6i+YyssDcbZM6msNqvPj
qVDp/PBojOJc/U2vYysLcbVw9WgvDW3LAteKN8OjaF2ULjiduv9uuPV5nIdeFofHP3HB0vDzgOnp
pV7McELoRx5f/gu6n620z3zZOgfwgCiEn9mrczwflY3Q7cLEvdXKcd2lVoeCy/IXgC9aNaBEmBXt
1vy34lmk/C2x12wbLGi1rnvtyVsjb2fVLaJPg5jQbNYl0k5VIVV5HIDlaw7K03O7IlK8oKtMWVoc
Dp7JoGInHUADFVHSBKNz+qreNVd+7VUanRxtXmX0j+Di21oTUcjT9Z+OJEaUFsJB9x0tHuI1AI05
WR+WultlRnfnIuHeoVVxAwnF3UaTuWJhPzdqrnUB1OyYHRuV6mFeCCE8mhnG3rqQMwg2TDKt+AY6
Qf27EyHEBzGFN01VQEfhZc4pHzIyD2JIh83FNVv4bu8qsBClScafgD24ZGGfJMkw/v2GaHVzGfTE
kraBjdXT6Bg6Z+dKDUA6o14FZKQxXfdJr+Q/Wjx01VwhyVpOfLb/B3XJdrO1j77MYYcBkyHVbXCV
TPZ6//ugEIXg14Qnud5WSyHrE8zRsmAh3IGXpkazLoLAEZ5OnW9TG8k6sKqvL/+SYhAYYfO1oKYL
IcMIY4JtcwmoU0mvLdUtbsuLPM6xHxzV7+K3AiErxMEueLOV6TWzBDsNH/NGPEBZUGdixDHawqfS
id3djWim0UfuNdShWBcfIMQlm1uwA3HBvYooobUneuB0GPVJmaqwpX1yxVNHMUbxhZPN/eTuklFl
OWbJTrk0EQOVXBKMAV8vQb/1uORmlojiaipd4APloYx5sEM/rfBmM0XoNsZu2W81F6AnpZ1ObawY
l1fb+UiwUTqn4l/Rb8JkJY5DFb7GYaOwl99eoiNu2wbf6nzbezN7JPJPk8nFbhCsA9gA1vwDeif9
oLMEnboKESbqoVqXHTSWl8zyMBd6Ezb6eomnwZhvJygACNvS3HWCXABv2QRa0X+nrGM0ga8pSN+3
LRZ/WM7wIQMAcsjWOMSHRrGyoNvCZkWYSzm2cc7kOv8mbywBjpzMyRgcslTccHZxjR8gePSmk/V1
w/ulPbhbmOV9polYft9fW+Lwl+KMVlCbkDkP5HxxYKIInhxv/+dWFSpipJmQfrQg4ldu+t1gz5A7
W+MYPdKPiTRW+nR+beGDZXw3ZrnZYYjzfmQf8T+ANzd+AmHNy0cjyIHOubaD4ewas8qXCZcngwDc
0Afoyerl1cSIRSKzQYCSnj8ASr3l5M0Fpzd/IitV3Bn+qGSt7X5OZ7M9IXt+rix2SGgFjLX/eaTz
QBhlh1b0znRURGL1Q+g/uph596jnR2XP+DlwbS9ilBInsz8xsrwjfJt017QRkYWEobIDZrSHoAXd
IMS32z/D1K9RiWKRZdZ6Zq+4jA2HUXwW6/4uR3MU47Mrxij1PFwg447oz6IDfB2O75LqHB/BP7aH
H34XN9J6IBgVIGfW923ntQuUaXJXbz8AykwWmm7rBzmyCJDqjwRthPDS2wI2ds81wzUI2Zm3n6yt
UHe0QJn9m5a1VCbY2y1x+FmGjW5eZAXMHy4t3MUzMA+ylVAB11EKXlWebEic02JYI4O1m0tByaHd
I0u3QaMOrXDiGsdgZhvq4p+FmdKt9xTX5d7f/mtHxaiiwB/IXplFPIVNuKudlTMGQPrG+XAA1d2M
AlwIS9XtRJWFbRg6IpDALUMNfsigYYjFKokM3/MTFhHvZL/w6gz6w7+HXObTh4kIkyp0g+NMoSMR
rmjm/ujFEPhCjpbz5Gi1YBAry36Ei0jjomOzJr1F0Lj70ACDU2JxwISJPXGnmrpJmlvIjb1TsXhm
nCwJbPvPcYo65ycsvmekr27oapCREV2kfau7z8HgoafRqmMFzCHtoyFHAH2iJRBHgP+xpXV9//U/
ooqmAStKJFBErOnSO7xhsacNMPZc5OjZHZbwev3WmponOhiIIldvM3v+bi+pefRmaygJkA8NOcKD
hX+UotcWH3Nadxhcz2VyB3+PMZRvLqcRG09p65gYC1X/RYj0vDTH5SDa9X+xHQxC4G2H8MM3jCUt
JYJdd/4Ejc+JSzFi7QUiutgBsq4dAcGOGewzojKNhtzFHXB7/5knYPC/C5lDGdCmQQ/Nl3hE/GrG
WqEu2p4N5kZlOWdy3IOqe9r8t3Uj+zAg7DNrfO5F987yaWXcY+4IWod3rQfLX2bw8dl4A5f6Bpd1
lUMYQtl/AsxzsBFUCb037qOmRsRuY/w10D+/aKirXGmxNlG7mJGLpq0Wx/kHrDpc3h4t9lD0Jqx7
qMBSEqeLvpvaZL/9ojnKSp1Yduv/EsWghMXHdtuf31D4hulm5qDQyjZ1gH3iGK6dktOIBQ/GKj25
JyjGzhw3oCe9MVgFi0oln0Vh7VZKHu2WlhtX8GCJhdmhtb39cugpnsSXUqRmjr6dJ1thIS1Rio0U
aEZwuQ3as2854KQGgz/h00SM5mfARFtx6Vx5nB6qC01zBsyEIqLlYDGXL0N7PAkviTIwT3qqVWkB
BZbOCifz3PhqsRRlcijWZ6rdVK10ABq/Fa+UYvay5ywwhMt59DnR5EC8oDAQS0nixYBWYelq/rev
U2tBD2BnLLwgUONCvhnUFfBpcnqvJZ5+d7FYCjTl/c/PB5t5lH5cSE09qDwxuyKNarb0YtWSDSYq
hYfYoSegDK2u6inYuhIOZObwVUkzCv3cj5nGCHtVmn/U4+3WUCg040FlOS1CV7rrXTQUqgxEjyna
QB03wc4Tgd3sRH1yvmGHI7GVPMgSY3hBDykiHVpFiAnhrxnKWY2hBg2+4s5l4FrB255nTR+h3tMq
OWpYBcd7ZQZszafJhWPfMq9o2mUwoGcvhrPcyVr4IRGeaKsB54pmlJkyj132h1rIKTdQuOLzTf9M
Yq+KHUOKx76ANgVmWcBbwo71PxdDtskKWfEfKy96publfWtrOJhGGeU8qgv7U7p++23QB/awVcMX
koF1Yi7w1bs7BINubsHYTcs+IblYtKB+ayyYtRdt9GjzovTzF6pOP2uA/7MTS5mQPplZw+fWT+Gc
4iExBoYa6prJ0F3uY+xS0NUOaU8ovr3iTldfJL4gZhRvYNoepiqEJxsfK5eSuN315z3TGwYYBYlg
bmHs00zuwUZAJiIjhA49C++9Qy+nBWjzhyok+QM+FH/upI+d+L6KfbjEfKfInJ5mXqndVnfXOFfa
MorQdIpV4TmTsZvmwb0zVjzGIbbsBl1h333Q2jNZ1lQ5NyThzychTcpc6CS0yL+8/ByZ0YlZ77fG
UPEdNAzmW/qAABItRzKV6JHBvLt06Rw134YwXzmqCrHhtEZkFkA6jfRKM31MbV5Uh00f5/DV8OiJ
O8UEQltCAVUIniUHJJlUP1AKrR4J5mL3/3dXEHZPPa6LIJky1miZY3AoEpPASKXj17HEGeaQr1wM
TFbHO+RUhpGZj0ChyJSTUdLND1oKfWQIVnoQ/5332v4Rz1uUdCc9mJqSb/ml9ohmKahleC3zTPVU
VSYK+574mx/2phDLCIW+lPfMxn7YnhUg/maDD/+X8pAW3QI2ziue0pcle0zo6ITnEgSp1ZsyXM01
Q7WrwLaGIzYzh1kyOr0iU4TEYlpPGHej4lIok5/33mBWKQSg+CmpQq+yUk3xL8klODTnBolD7s3C
y6vXg5sx/8K0u/hUOsTdzL1icAptcQxMlQS38H4x6QFwjdYDXKpx1wH9vSueYtCXwECIAvbPblBB
wzMRJu3qyYVgtsOPkjWU8G3rRADmYnE+maXTLXEOQLHnffed4JT2g+9MH9Ju9rejSRiUhs2fDAjJ
/vGQpkkDBHgLCVuviCl/b9a3138C9kDqCnHIzT78/krHlhCbAjW6kRMDL4nA1ksy/9zSnn/Ew2rs
NoMCY5nBYHrvKNcoZN/5iXR8K2psxKJ68kD6FM2f7M1uWdHz+mw0rm2i9E1y6oXKESNUFgVCU4NT
KH0+YxIlj1JOkGcRAGJSQC5LAYl9mz+7a/yWyz277ANTlv+ZjxQ6migKalhQIpyuicP7Zx4WuAE4
B2Ud0m0WB59Hv8geBAzfzjFqpegUF0tf6iXla2nIht2Mh1u74h6KPbBmpSm/n1q1O0XIQpRaIPyT
wpRwJq+Y9yDN26ioFJzxnGCVN8JtB5Q1qlfY9Da5K24+ak/kCvUJIk7eruyG9NL5t0CTTMwA7abs
TqUzvmJtgxKpOiK5ihqj8eCbrVmipa2wcsqyro68WRBxZoK0wT9UWhVvvpzGm5YPirjHB/H3Q5+I
wMmRvARntk2ot5u0g4GysxD6zhm19TLvVn+sziY80N479x7OULNQaVZZt1wA3pCN4HG5j8HtcY9A
KSkFpwDS60MULSG1sfFcaZ0rhGVfYZAt/SCdxqt7k7GJnEpepd0V8gFzeVBDsS/rXZ7e3hF337Oj
Tl15weld9hg+RJRqF/I1ZSLAyj3MPGs05M0u0GYg0iD1B57bxtrC7KBiQ6vfXsdDLYeWzfCTcILK
BlEZQIkBxeC4KLhPI6FlBy0Q/GfjTsHayber3b64c/5878oze/q5kZlaJTv6GLU3Dzxi4kA5R7hJ
AL+GVySOXtMs5IwdvJd6AT/NJscQIV9GP6UuQfLFo5SeALZXdsXGjR5K3AlShPNn0VNlEGwkTt8a
a1tqTvLVFfO/iGfj9EOYkhFWT7i/Yi8GWuOzUzh+Tf4RiAgpOWChtnGcTp8YK8eVwkjRAbkLFn0T
c4uZeO5YgUqymudj6TDUG/Kat0zUPR9JRQG5tK+UVOhYlFmrhG69UFqtZVUcTialyn0d4jr7eqk/
HnsfKWtmPciYGwpY1rrqG/z2pXfcHbaYcI/L6eKn81Z37N8RIl132OmPu1/w0Pgz4D32vXuuf0ZL
uHGkLMt/uwV89MyWc8tSfcuKEfw2ijE798TqqfnsxeiorEw/oD5jcDIQKzg831jc4S49pZB0paCs
OZ6G/GlNRwC6IF+h9Qm0V/H8nBwRensoD2m83KS3KRqFE7TwPyo81jsFYzqkB5TdDU+25DWIYPLt
ukrAcD51Z8Zp4NtjMfrKh6sJcw0tcXA0vheJA8tljsCYpqyGApPx+4Jv6RgGkUdBLG7DyJE5RO2a
7nlFX/ZSrpCpB/eX0BEbvyMSCPSzSAa1U1DhPsLbHMX9qGS9OPnwtEoLGcyDDWbsQ4E5cCgItAZK
pzIeH6YxpI9O87Ptu3XoYcy4pYMxpRxFkv8liXiqR2CzPPd2rZySptDVUJ2VGgZZqdqt+ZEyIG3v
HihfWWuiIBocAK76EPVaYaBXC0uxQcr+jHLRvnXDHYp+Thdhj/GaPMmExdMGtvbzwQ3zAWXPHBno
g2RH8NjLeudvwWAd73ZBxUgKUM35Ny4wxTQ/TWhA8OYmoMxBNGcDMta+jArXQ2gU3mTE/IUqh/dn
4Q94oKHrW5ntRkUiFe1K2+Wph58OxkIM0/0yn6IrgqrRbdGml/qJKB+D9EYYQVOd/1xF7qeyvLYc
lL2c4IQrtx49YegNNaikBO75RLdRyDtWj4mIJy4ER6LitILT0sY82CATbiQBkmDOzhKRjl/oOah5
exFX0FgcviH4+oT7XfrJNhJRMZ37fL6w1I+F8CsRJa97eJpP+5mnTZ4n6QyZjIMTxHmF76+CwkdK
PqyPa8oewN+PKXVneTC4fl8R3Yf4QVg5FtO10vKmth74Axnl3O2xHkTCQvgOp4j40TvrjbGdIIW3
GDpKsGmDLD2801cgnZ5aAGOUvSn1ljNjrga27ifHcdLCmbG0phtwwyzJbww3C2Qf60TyW/ssbug2
y9lZvAmx/bTxcxgW/HtS6ER58pDTibjkwzfmFAa8LVujtwoWxgv+521jByU5uMUmaW1mxAv1xhu8
9vokjrpBWQZewrl/QYs53LvQ2HNf0DwKRuY/SCZmjkR4MHjdenGUlaBfkH6PyOmwO7LkkGv2aVIr
BhvlGdklnl5GpSTr+6Ny4doOIQjy5EOxdflY0bbUN+0++P0kXduWCjVOFvq2csVOrblWF2rHZUbX
KKo/m5ByDK9KOZgFt1FY6TjAI6wlXL/HqOvihNmsgLFrgm1AaWv2VweDnES05GbMwfd5O1PaJhfG
Z5qVnPwfznIkBV1jbcWgaW6hhjuW2dTXzQQoZSeP3FikD4GTtz0oIBD5GACvApRdR2q1G/WN33Jf
h/LCzX+phcPSrza+rTvmVHFYG0bYpxcCk6fOCJGrsttGKggVsB9RWK+spVdBeL97CzgWt8NoOH8r
C2gkPKEMMzNpC0wWNt3ph0/eAVfi/0uOoiHxh2Y3zgsFW6GY8JRWrixGTmfkgP9SEcT2gxogANxW
8uSFnRlqg0jefx5pSQnf2Z/Q3w79F81tDymFqIlHNfI7QleWJfzUXoNa9GJNMPSYaggFCPxQ1My7
YaIBuA7cIBEl36y78jCdeLeSE+42IdEZoteUDWynV1HxR/XOhY2St5sFWVM+CL2Pmzauqnn4qwJR
sUmyYB8UGO9vXNyAy2pKK7x06w0g11ke81kYJlpf4Gy0GVDyCzzoi+QLzW1AuqAriNeX5yFHx8MQ
P5GFJfPUaG7noVii1Hoz4f/gICnTRYrmEmCeoGGRjrp1CtxZSt138M5yPJ6ATZ4dMrfzv0aq8Za2
b5IfernkYieWSdvU5xNFkQEBsGWd40jG5/PpllUFRqBybP2YL9KsNjkTBYViHixQ6ANWvFOsdudS
6rXJbff9h5gU86cvOOLrv+q9tsUH5HxlyVNqFvJCvVnhVhadxI7UyS+Ue/i+LbWyQZFUB9qTKgzf
YaxDWCHhScHaFkMjnVzQpWsBFSR7u+K1OWigCqHzadLewSDlyGIpJ9YtDWGBtKHqtnL12a0d/7oO
fp58ew+6jXeiuFI8iyQwLtFXdyniIrQccSsXDcOwzA8Ss97KUVKiWVtQfmTj2iGK/aHFYWBBdI4I
2c1aaaQQ+LQTVck/ZNolbjBXz/YN6RApc6ARPodILa+AhTa0QlOXUI3sh7ceMkhJwQAeiUVapvI+
TV1zZaYrkL+H0Wd3X+AbD3mNgkwRw8C30jvApfCFOcH8e+p1YU4Zbn3LVTc1HDFzoWnzLlQqYKs4
+1sCsvODq/APUuyw+f8kBZFgAEulJBHjlWSWrEJ7esku/wb6ZFEg+y5VFCm5um9eBn5vkK0PsO0H
9ysZ1CVFB0IyANCgCLwIW5ctk46v5+3eSJxZ976fXY7rd6Gi34MU5XuSuhepnyqHkfa1yYq5EULl
kVCuaMkhPkKyliztqT4yF8TUVSOxQapfCS93NCf0FJPtkjzIAKaxHR6is4ThR9+eWa0KWiSYxx5f
o3UnmhOxDxCDwD6xEbgiZClq62RIIbTFP1EibJuzdctia+vlriOo80OBGBBxxlH5tCh4lv00HoPo
bLuFALV1geZRJ3PsUAqUa+zdc+7F3LLFA1b6GnKmAsadr+G7KWaWetidGh169PkO5QelpH63Q5CO
upHiC1JbNwHJZsYb7Kiy3USebKfXP2GYk6SripM5G89Az68RH2hpb7Bb6FSdFIy0X7jLJ5J/97fE
HpAneZyxXkKqNrNhAm+3ndVdERHxlscBkeZXDftr42x4RqrRmUOk1qxVS3ZH1RxdamVvsyjjTjNQ
HzPGvWcfE0DNQ8r3AXzvP1Sak0DFDcPcPebm9TqTUEQo7gXetM6rirZ0BOzzFSYmpwXRTl/ai7pn
MmPzsAg4P9PVZOnQxRvFTVsSap/7FBN9ha4HuzGDSyOHK5/116H0vpjbVn4hF7F/t1EIwnPBLSRe
IcyFY5YoU//DmBYPefdWQTLtUQmFa8GV0PAIz0Rzp6oU7r1k1YbxABVgPu68AzD3tJkbhRsYOHSV
3GUtGyHX0xuFo7IdysuorVOhGke4akTkUrsjl7T7AW5zpXU/kv1gdV6RwbwWrS9hheaHKU0IjuGL
Bf39p7FA9bU0RYGZH3zraJnsRofHpkKYkkLBcoJZV2rtnEGODZfLKN5z7eKFDdeb97sdHjxoJEqg
vIZgO1+ObRsEq+E90wHf+13bVrYWs7A6xf+FL6OeHmmWPuPPd8lKttDgiQ2O9G1YUY76V4yVfP+d
tdcWnWP6s2KwasuX1BM0f9dNx9AXleZ2fW11Ioiz+ZTrNE9dtA9JwUgyThRZkmaXq2ZCagSW8aV9
hWpE8KK3a59BkQFZB+E0FW8yeAo5oF9FKtYT0ruB6Hx9JS1b3E/l6ACDzXtqrPULm2HEZEO73S/d
jiDQiYwuCKAXwzUs4JFSE4yxduMtu+H9A1+8OgW7Ra4FqU7qS2h23YbHWqlwD5v0vD0FtY2thI91
oZKSloXlZ6g/mywk4V8P9voZx6OFUMYFkQynfln2Xxnlcu7zlqhLDfXpzBnsKj2M3iOyQG8SlQxA
nLcWCEHt+HvF5D+TuyvWBoH3c3WlLxqBDct/Ho7csVaw1lBbPVwCgrlm7Y//n4e1FFiMcNcKAoXE
lBlSLs+whvsjsY6tCbb7xh4K91GTAgcyKIMCtSC8cSMU02vj78L88lxWyOYjfKvc2Gms/rf6225V
PKkuNZJ30fqZ+o9OywDXKae5DF2yRMs4PqIUlQd+WkcQAoVlUdAlOcoEv5+lznmooS9m3wekF0xs
N/6AjIDllUmZGqd82IJo9Vjh5WR1OcU2EpDQWtbxXkDW2L4i2LHuAwUf24zhkbPGGiswT1FywGud
NqmCat3wPHPAh0XN8xuoHHPrkpZCwdOvPHUHET4I7buOQaQOTNgn1ma+LKks+DUjVtjy1nK3m0bd
XGzCGHwTbjegDddovJ44AnyeHUIii4LR2ld0CIyvAo+DBcrf/m2cxpSNHujntuINBYCs4Ld6cKY5
HR2VvJ1iB0u8ibj7LLe6/oHKvEFYxM2tWVxH2HbNua8+3re7K4JUSLTEw2iDIXY17aizvJe47tCv
IlN/rOZy85tODSOdETM1KsyciD8JObou8Gsb/f8JU7sCqsI8J7bhRPMrCRj7v/V3rJA9YJpzytMo
KdO7AnAOErNpj+jlHdghFNX+PAuAPMz/mYrwtE4hYKCpr8e76S99y8jROjOa605LJ1leTK8eEpaO
yEgQRrP9RS+4pBewDeVIruDX1+St+Qv72euvHjOknYN/6NrC7uHWtGS5PlFhnQ2QkCqYIaVWMPE9
d3MADUjEGQ3ffbNPdEnpH23JwqAV/IlwpoyX8diedg+TWi6qqQGaHfPLv0zqQRVoscxJemtmwkfB
CikduxF5omWLCNgwjd7vze0j2XKn/hhFy9z/lD5KIKoNLw9M0GAEwODPXwCyV88JomTdk/CpBss7
OUfJG9POVAo4YktraUTIymDug0VU19pfT+uZ4oW4AjZZKEMtNgd6piS8UyI5YCUpxa2sIqTQ1AuW
w0jbY1/h8SG4WyTZz1otveKAUwmKqDD3thce+ZEkfHE+hOhVahTMuJZI22upGbxjrd2Bcgy4kXz4
/QFquzT7fP9d3YE8VvgLh7BFSw0zSkwdNSeSx+c3wo7E+cgxuBxoZOORd6R2W4tSs70+9b9AVB/0
4LYkfZssyzd5ZidIGM2z4gi4KME5zNIjiWYO1Lr7VSZqtVQpnjYsYKBdyM0Qg0Ln0ABT+axOjfpc
UjAyRQ6rRl7UtltjQFXtYo7N5XY3rJDw6uu3MJAhPqmcnOmzsrdu6zXhHVGfRUEOpRCpg1dW+lXt
8MqhNGyLw1HQ9awAkz229JoO77iEFnkdvSrNV6iJyyVCFmgLKZhk188A5jiyLv2cPXZp9k6fAT9L
jnECi260NtdK4HFslE5dUguaHgz8zQcaqEAbYE2bN85kStS8NMd1sB/sNAIwSF1u4H6OzyfaD7Mn
DTRDho6o6EApascu/FQ/jgbmXYmhqnooCuQ4nqP1pEVQW2WpH3niNf4aR+bx5IkGJ5agQMccuxc1
wji1kFGWmIOqq0mqFLp4JNLuW+4VF8jprB8AnqJaeiOfRfYzVoA34dK0MXk7x8zCTrG/QiHJoyeW
yRB1d+QVQwrRUaTbrxZ+PIqLPBJa39eDIWVE3Hv0KWXSLNeIqiwUlt78odhGJLDeTqgs8lJflK2Y
LZF2Vln86TWKWbTDLH/9m0tYgCS89Cx617xzVwQRnrKiateUuQqMfnwb7LIASKhYUonUOR9/GUcQ
66I0kQ/E0msPo69mKsh0Ke7dGLHCwodSxF5yE9Z77ho4F7r2bwTak3x0TPQB7HzRvovdn3+Y2ZkG
gQnoykVDLGUv12JgrI7H25fDD9ZGTmv+1kWuCxF2kyoUeJJe2ftYTMcBlD8iSDibCLR7PBBGyxIN
Ji5kq9rvDX38Rd5ZXgEbLJu15NxvQXmhg+2k7iO8fceabkfdD1A0iKZOnzSi2C4OAW8SLtCw/tM3
94IgMJ08iYB4QsseOOcLTCmo4BALRtftOEIJD9Ll1TE3Ga1NlwaOoH1DNJlMfrszcbcPKOSvLYMT
eeXfAw/NhjN2DpR7/hnAdHXmyJgO5pcOML0WSG1ntx3rO0yv6n7TV3jExDwyLIODwlgj9G0cJ9Fb
oFX6Ue9trzg09DP95t1mGoxMaHAdwpSa6Y86z+Se8B4i8DFnQQbASyjSUBSGXolwUDTeipe87Vdl
JqoHFcxtlmF8CEIZMYApynje9Z+ALmV/3pr0SImkM7pePO3f0OBAVDjIEx1XgFVYeKUVv8STaf+j
zP0TVQPq/NKFFD3Xc80TnKikBx2O5grEPwdqZjJ6c3f2E8fJI6PiDriDV3KSBLrVngzxvjSlwqkD
72fDq9LBNaH/Ya7OT2w1SVBvdd2PlvOxu9rLEKTiuOYu03yEi2wjWsJDlDtK+BaS0TrSbVb/0vJ1
06sby/QlNVyzf8gdFUORKS9rAVHDITFmCUfa0eyn7NQKJ6obSyK8hW2yatQMe1o76Gfq8YtwtPlx
jyUNByhUF/tHfWsjzO/qrx6Klu7UOPZ29a2XwEV80Uh+tZaKcXpPFsbxsxSFRYagMcdWjpEuB2Yd
tJhqCitW+xj6X9ZVXrLy0yqIjokjvQFStimOUY8rpnf2mMUsPhLa0oNQtYCOukjcjlFi4ThDSTrP
nU7O7h/dIUpl/rNDlRRWB7fkfi2wXS2g6EWfkrxXABdDHyrWh+aHIPq8dZphS1ohkDBPMxnODEP/
X2MyGz1wK6CvpFYOFJxOoyfjqNoPfg3bRLNIid66Vf2xgARPD4E1e4plfUTYdACnomzZyKIWo8qE
iaP0/XMHn66lKuOyDo/5YlBElqUwszHalvEjlWWbHInAe0B2Sq+D0wBHQ6m1/VUMSBs2idjPXwNL
wzvRqhbaUePS5zn8E5xiEA16KQ4JpdEPp54ngEGmpg5UlRU38S1X/Xm2LXxsHVMw5PaGv8yhJX5H
2HdtvfRhnivqW9nZnaD85MbPK2dpAKT4ify1lJ9pNZTrUKB0YEHXAJfhSFOV2aQygF4AaaeTWNk0
4WBHi1aKmj0bMh8Xk7HdaMiq0OOAUbPrfysDrg01pl3A6E9U1LQTFhv3/JMfqCvY1M1au6Z/Ade9
u9SRgiZtQP9n3THX3qRP2sidqSZqh4q6xR7sumsF+r5cA5a1pISt2YX2lnr4J+hksP6g/0HznMTd
/UK7oI0QqyGI5tudouSjT0RBMxNmj9xvAxhOqFeuwTPlBWyyiiXxY5LYizvq/fGsUhNWH2q1hZzy
JzrGI5Z4K8Q+LTZOYvfrYbHVDJx7hsTl/S7KxkRbR50Awc6iBU7G98aYCRJlmLP55MKk9naZOC8D
QOwzjKg8V4Iws411YJB2xcBS3UnPS81hRCUKfEk/kOyWB1ui6pXP7FWlOHFbjUVsJu43Ja4v9TdJ
REy8j0Qtgt3WVqM0nWBAQRN1yDipQoOXY8BhKBmHeqd497z880uYgLilU4cQpSFcWsl+AscpXhYW
xiMJyVxGv+IRO7iSh1KwZGDjOLKYFVEXY+uMH4dX8gELdYkMW8F3cp5nZYE4lkEndjAWiDlkqhgF
/XSIPXePj0UWTcRTMOt1aGPlHjEo6n9D2gG6g7ZzVqssCyMMk8BLnVzI2OVV91GhcPilXFTIv2C5
AAqum+Sz9yZjqMAB5N94+o1fJXrhbnV4qMxyX49IKfyedbFehPdijK50c7lcXBW7LIyHte1fDYz3
YhVRIeEpVJyEFBLKRhw3rbJYiKyIEEZvfduSFy+6PVV8G/oDPGcJ0Gm8l3jNCiZrhrtxb/tuwFFj
E+s/GX6oApW1jc7mUKNl69JPes4fg9BXahZrVzGLpPL+1yRQs3cswHGxjTSY5piE2i1pdeLFWevL
densqwDGGpiTcO+UIQHEb5FzHxBlA4gDG8t/xMpOHInrJRXfIKABn0GYXMKakVTshSBZx1rOREzR
N/XGkqA/pzFR/tytKNoJd1217k3TG3MNcnxZq0AgyrR/UqxjccqLI2uCOkKNVfKEBCrEObAK6mmr
oxT4Nc0uFsyGhBtU7+IkyUR+p/NlWE3lDv/14loLm4kd2WEPKWc0bSt7B70TAUeQs8GSzWESJ+Ou
TTszkh1rNp5XrIccHgQmi3bh1K5sRGeJZ9bt5eLr6Kl59BN0Hg631NsZ2nM9vQtJpMpIuO1pBH90
wMGtS0WAxf+H35TAARzXwlV9NChlfucVsC8Q2UppDGNJ1dVnX5XHR0iUMGLzM0QqIsxTt5zJIp04
ZUa3rBpl/thL2XBXrGnZtjpABgsyIjaUDVewVhpvn0tf+gK5gxtNOb3YMUH1jEBP2N01TReQflVu
y6QNKGzxlcXQskSpoBGOQvN1EqLvmZ/zOruY31H89/Joqv/xXQTKq3TCCT6zy9+BxR2CVV5AtDhA
Iwrvj6ecifckNHfYVa3ARIp62Qn8ZGt5UEirch9IYlnPZ0PdcP7bbrcdmQhLZtPKt0YLVZvK554q
dxOaThDOyb8zJ9cjjqHS7gbt/w4MKeFK9pl6vUIO0k+TIZ1EcXHWNPOYpZedT64icubDXDurmHeS
bbPcLB2z3HDj1WQnlIPBkGCPTPWdXuaHBYjSxamE178uw23T2Vrp+9TgRnHyFLDclT6Z9ESqio3r
zRxId3jGP95dMLDHrMZKh6CUfcCegCIGPPRQcFYoplWoUkKveC6+Bn8ri46Kwd9O2sqck//5C78I
vWI6R8Hbe63LJJd6o7ZxcZT/MCKG4iN0ni/jD5uaY6eJtdHBqZfP1Ru9CEmIYPz4/oRpuFijuMAi
Kc7x9ttp4/RCdyGd4o1TUFRLAp9c7xxfL4Hu6lEflwpHsv5aPWx3e+V1jfClrpTHLfFuwRJSiNzD
Kkv+vsqbQK8GQFF4A5uWzqfJYgcgS4vDBTPiX6RYwZUzVYYr1M5yjQ2dUI691+Qt9mAe/dIALAA1
y+PynYGeOM25eZ+uGRTohnu4PSBjkWVAOX+RgbVAiV6Tj4TKfqyYQh+nre64674bqzWPL6CMBD1a
6o1ap1xkdxjNZc4uy94BvSz4/e9f5+mYiXWxmwIw3liI4AMbZm9WEk4dNzs31x2s5jJgabsE/VgK
YP9wip0afcsnpAqrx8Tgrxnyz0PX9RLV1dxu1qfhtFIQR+Tc2IuPyfCSkwdhPbV68sKRq+oodux3
lW3ESqBphYbJM56KTsqMVETkVyQpCDR696J3WCSuQ/L5urXxbi4orIbtx5Pxj4kSP9oxemMqi7WD
dw6TGrcsV4AMB+OhIViz+gS9cCHilGTd+hTDmiQShx3gB78NrmaEbxqaOcro04quak3+ZLkw8qiV
UkhHUEkZyHh0cj+5Eb1X+73+iNoc4Z6i7AeNM02AJwXlkjTTQCyFUoizC3KnMsw17sQgEJVUqIhS
YRXt6ikXbLyQP3H+dI42ugHcYoNOYjBSERg1S+xv0bgrmPqtrPrCDU6m6JC56uTOzm7+C0bkT6ji
vRmXuaTA2zTyMValuD003bMcxHnI+/CG4MTnh+efXmI/306cCfWbun22MolIWBEhVb95rX0Rrxjg
LyYJkcfuIzbdgRj+fOZ+EGzTn3w0bqjDDYvGanvrpwTrZP5nN1FYxOSY0tA4wYxVM2wIhmEKDRiB
9VcL0VkLMw3vrGT9ahTWvbipim0VUgaFO6X/5XBYbZdVYxTD/49Scf+zxZRBXwrEgTFhy/481jk3
lM2NWYfGKc6uW9idF3VxKrPeqHWYARfxiVWW0IArHYv4+4jxKM/d4+/vXVQLHEl8kqwHa9iDg1S/
mm9be1kiPHugZHLc/aGbnMwLBT97cIQd3y360107jdfQZ/ad6WztHbC4FB3OERvATnSKtEtzL8N0
wDSblXJt7qdcrlJVbTREZiqWl8APv+i5xyKFChkv6Tv4mTB95csf8eFpBf1YkvjF1DjdTxaUFGIX
PSGJEBS7LEyd6jKRsnb8GC98LAo47Ru08lzdFo674wvJSXTRi/nBUe6looawgpjeDZv3poXZ3iLf
EnV36XWdPloGP2cn3UswpIX0clDrGDGXTIH1TqNAXEetAoMdjgbbDVMRWEn/ueeeayyeIFqqpbli
YY7vHpIowrgPoO464IwDKollVR/0FW6YunjeLMLjcs57aN9/mpZh2zxZhpQNtsfXmxwzdml24isK
ClCg1jSab+TflyOraJlCFy6Rrei6pySABNB2Eyff0XliGKJRhbQT3YoOtgJVy15n6HzCsh9ZaG90
Ew+clUP/oWmjJaqQA7Up0dK48g58Dw4vavWUCGHrIlNDw6sbM+7wa5ITrfGWHHvt+K/gQNkhFSB9
GbLfItm+dJ1KTScCgIOlL4clt+aeJRUnD/nHwNWQc0FFG3zOYQqFcM5Yk/7r3+Vex37cEgsvB0Gd
OsZcPS31pcyaR1zLUqMkJupGR9wRsqlRJ5yQlo9aDAwUInGDcne7Pb3Jbp9FS4LMmPFvs1VreVZx
GGMRWBOg7RvQFHSMTwsMqFCGoHiN75FbKTtWKQrI/9Xg7hle+B1m1TMw2ZrLl4/5IpnwdSgermz6
JzP19U7wbw7cDfWY1l7BHFhcWxGgHxLnroYzAbMvcLwLh+37R0zVoz/ZvSafUhc1AP/wRGlehXzE
WCcnzcnRsQe1coHe2w5GZHyka6S8LI4M9kL4T4PxvR+AvNqxpsOK1/XLiy+PRwvTa+ltGi/U4RYX
EIVi8pLED1s7CMqIKLxhgn+HcGcLaSQQUGg+cRt04LtGn+gYS0NGMF3/08h6/tTCzHYxU19ryTNR
6xcQJ6GA6Im8DO1/5wJenptc9/ycYuYMMtRTebC22VoOMYor3PgnvjMvf5cBMjX+7zvDx9VNsLET
VrFk2ntUF4KW+ON7IJ9JoxbEntERaMcOrIzbFRnl5jzHS/hsp2uJ79qCcYmvHvUsxidPSyhCAeba
yXScUbxyH4wAt87Pio3ywZxBpQ3EWZws0WPYQm1U/WM9v2WAM8OY03KEeSWJcN/g4YnL5sC5f8FB
K2X//Wcf+IiPCvcW1dJcdPcCa+YSPvdwZgYQImXSHnQytiOM8MSZ6uWqCraPF7FTjgdaiLE1VN16
N+OaXF7ezmbjHfp1RFnkDbI/OYP5OZC5tF/zxONF6b5b13GrrBwerzW3NLHGP4t6s2t1lrthCx79
I0EeJEmSFGrbDW9qKwN5lGX7LQRfIugKHgYgASIv4r6veSA9GmgQI7g4K8D19rjHlRI2G4F1ucme
QJ3ijYZ1jQ4QoPW986SFioKfc1quRXIFzyhui23AfoPwvku0w90QAX4xnfJXq2lRmE4bGeNzwx6K
klDdCsfKEGXOD9aSnarotSBVHz0ARLpn2K9OoOq1FDl2aIAd0JETKxOTt3t76NpeAnfklW/7JRZT
iJuZ4OhgdFyVxhMSfYGhgYDLJiyriPkKepDBytsK2/Sg/AtM5FMQoDe3larG1PWzXVgdRme+PrnC
Yrw/4uRrOIHHmOkCCJQS3E7c93RTNfSXPAcmUyV6ekG1G4htVX8gxRowMIj8C9pq16qlU1bcbAst
mmNFd2PHVpxCwGCYBu86lqDOhe6PXNpT85BrqyKNYtT9TmQ1TOVBc2/03yYMGT+HxOhLNKG7kcWF
C7q/xA4wkEKtyHVroaNLY2G9o32Ss2cBKvaqwiRecCL2Y3BKhIghYmNGEyZ4L85BeAA3lUIDKZd/
kcwfGnQq2/vbfMQ40sX+9ULQAe76vrCJ8xPTIK4mfyDjKjFykvoAPvHePP1PaTIQOdqGhewC1xBx
ScQTCSJ5K/b9N+KwcVbAFpfJpnPZeD9FspfNFtNYptrI7bRATs1K/+ZGvrnp0ZsfLZw2zbmCwp9m
6gAK1lbRRR/keHpaGBcPp+9a3yaRiAnDe0XdXYEdZcLtEjILSrSbrhYxNzfB4rEF0tuUzd9C7Dt9
n315TleBrXQJr2/NO+MgrMNK1FqppHEHj0ZWr7viK2HmUZYth202vPQVlUaIQFxG9GvkYNqsSXbt
ksC07I+pisGkvro+VZ6TyFpSag1D9n39O/iqqHFIYXHmuCgGF/8x526jRFqvN2K+YE+TyFKdp2UZ
VaVEW9D0iAmzhEGb4bdFk+aXJIk4Mrk0Io3zKn1t8ewCTBYz87q3vckhtDxKTZ0Mcc5pVX38w36B
tNDg8HJ8nyW0gKDzXU1cCfs5TcB4hi8aT4RXLiXkNVNyI82Fd4JStxzsyujuVkE5pIfKndT+kpCX
J0TEY7A+wIGhoxDsXsSenjYmQfFjAciENrzb3Y+tf6xy180pdo/49YNzDsKkWoO5GSuZsNo5RoQ7
EImsTYD0nbLCsMMgkD6YuIc1Qu3zC276Y/nH7IjcXLvcaHO6RccWhNurkMINzpqnfOZ5xhhzCBRk
6k1qq6IcvRkHqdgRbxNu/EQjm5/+MPeQoFYu/5+wiOHAx4Bt2LAmlli6V+TtvLVZztHla3ZgWuMz
dwoXPjkxCeLLcKOgBFZmWNCYAxPKSkhoDajRUaPNGrSe7lnDPHyUg17Z2cPUIDpdBU9Xr1eRNPVv
GW3vDEWNIdw/4W0ioy0dHfWSu9jAfjhuxoS1eQbFDqZAW3D1yzrISZTdLpcLfJh8Dw6S5OL6XBsy
Ox9336rxYR8l8GxL1l788bSE2ziXv4AXR5oOUmWHkknAkTcRWzQhbGKw9QTB+gS1oli75M+fojcP
dQ4yD+tU+aF0o4uCNISS5mBav1v07xSskhwitNHulTfdMXwpOldn8iSrq0NFE4xy4TDmEf6Hzhg0
uNP0DMsOVMPJ76NM7cUuAsfFfl5Bd0mq5Twrcsqw/Mj3c4sUpud2GXuiGMNuctXIAzDCAVBOpbRe
NdCgx0yN/wn2yShvCk/5DMcTu569C+GvDs4uf/Tr9v6ONuYKvODCdxWGawxazpghXTckIdYGGVTJ
pFjr2/aZVq5yBgA6+1URG+fodzrgMMfvTDGVxIts9kDpElYaU4iv43juquAwjs2BHaaVpMsscNCN
tttwwiBOl9WmrqHyu9a+i3rM6ZmUTX1y7iEBaBwc038+KShjqeSrZXTtA4HefiFs4yM5UzOSn9uS
C/nuQ/zG1lSJ/3nlPMt0Vy0LJWCZMBoriWsqvaaUJuoxI7oD2AV29OxywKat4A2Wv7V+abXkOXN7
ykBeVQ2BTvxRRfhbxzrCDfx/XWBiqx/w3BcI7m3lkUY3FQyZ1qY51ODQecR6oXlBDaUECpVEnSSp
BX09KapGDqkCw8fKvzF+5m2hj2BnMRm0DJ6KUUX+OrStTtiBVD2lVdhX2BqZ1khu8QVHmUPhEzAh
qTVALj0A40417JVtk8GCtzpOQTLacWkqqII5RfFO661h8IyUcKuFQpFAIoQYfJXjjH95VvAvAKyW
+SFXj93YdTVdKTNhtH1FEE0F6iNWFi5D4SD5lKBA9sZ2wxyUbqQh1QiUkv4sNJLH0WE4ZSpBh4eC
47WsFfaZCg/wQPZuQF/wCdZYXMJyYUKBFCx3tbGZqdIpFKptWb8gDncLmYLVMDfrNSIDqslpsi2I
MFNKFKV8HFNEL6P1OfwFdT9hzCU2iYZpfxP+72r5giu656+NHczXtSpSsZ7DQmb6mmEtLGWwFWop
J0wdjz2FeRPalIt6y9zqxm+k6f1msweaYtBbVRm0bD5aBuaZRTDZiikAom+2lZ7MO9js/B4hT7qF
f3ScMCFS/th0oN1LQGQTpt3VFml7M9RdK7ZnHzmfcEC5oWavv6DPrn2JAx8GsOuFr5VTkaRehioM
g7vwtMNy2MObu+zaShXllTv3arVqJwZJoOvfRwR5nLHnJ4zksPD5SPuhS3YtW1s5IDSu2Ce85PZn
mzRum+2fIerlP9510f2hkgFxkIfD8MIMILMuyctAznRpXCQddVLtenMS8rMpr3HHoe2hARDk/Z6x
OcQtslkvA9yH2/2Qu8oejAyVqyq0h8ehRMzaAH2NktUygL04nIcUPVwRppi7u6BMxLnoJId+zmEx
ZmhC0byQ57DpVddsd8uscxEvQCQIH8s3DGffaS5+28cnRoErwEiZaCn9741rE4eYYzIM48ZSecpv
q5gBS0GBkkLfs/hIQeSKwZQEl+kGFzva2G5CTBiHxRJ//2lngUiLakUoSLnhU7yi/npuG4P5+BqG
jVY38kQ8z+gzpy626MCwl0SS6bgvkhC0ONniXjjsO3mTpaCDdBM9+IIIs5TV/8wn0nfritc/HwUC
AhmVZTSs6mDtKdhDbqXYHpiEG2Xd1+wTOXFUZpevAP1Qwi9VDXsJf2ZPj8Inn6tv73HwGE1vCofg
gVzvUAVF02EY5bw9gA2ggkplTDxbYH1eV5YLHZA0WS18QqcloTkwQ9XU4rIgT+gGHAdjyShXCPRd
LZiVdbD7OxihpClSxoyDKBWPR9MJCkVeekvX6OiV67sTHwfRtVfsNyLV6jUnh7UQLitu2oZKNafl
HbKEDNa25tlo+fJV61VNDW1uHZ8nzZdanGZKP3tJE1L0P5Lq+65DyjnaRGdXqRfaQ32JY+PBxMIa
Kb/DvYp5cxxXP7BdWfSJcPuhV/CNPW2HPNRQRUnqMH9Yq0nN1fauyObWhKbzOWw5WvhQPhJnfna9
W2gI+bNzpciEcjsqzzeokgNObypbzO0baf0JDLuqEk3++BFj9KVOcWGgo8+K1E3anUixIPZ65y+O
WyrAWVclbHFk6onqqa8Q9GQ0FLbO5J3KyxAdh7zlOyyw0EniOmOAl0IhsCylcYsofQyb/gKacZnr
ejOUK0Or4HiNd5aD8/u9d3yUcucXtjLQE8oNMK1xvem6ZlQXJ6wKspEO+1USBQZqVW41UzeZyd8+
n1h2988jNA3LlCq47s+apPUDNS4j9RP3oLx3Y33R0oU2SFDg0if1cbjVNVm2iBDEPpiFQZJEqjvt
bo/a3YyRhYtwVnQHDqbSS0sNp17F8zvIWfIvpacxWyGMAIx5fdyLCvCiOBwMVezPiV/4eJqBdVBv
TMZH+80+UyLHHRRFMOeIsoUe4CuCTT9rU50QXYhPggjG+K+HaofGyreD7elk1B5gNuAXO8Mb7Stp
kzlYX5B81dGlydlzyUpje0EBwsGh2eTZGDROX28z3bW/sf4TMkW9arJ24dqvn0v0pfIIYNT6n2MS
/Jn3nAmBo9kXNlpO40siT0Qoq+VlmTf7RrId20OhIIQjVCjBEZme8CpYE4fnnz9J/S3PU88dENbk
VzkZ7Ta4SSvMUeH+iUAfDSUofo8u4/J4iXRuGAX12scw1uU3jRVzEkyorV3fQtMVLL60MARoW+Vz
KG/r4+9eBhp1ORMfNaOhzNcoz1bRZy1AhCPei51DKhH9zeLtMfYkFc7+wIO51/ds4IHrtYM8y6+c
L4uedvR8knJ2nirdevpn9lA5wGSHu6mIbx4BIwRg5dZ8R0YpMv2re7fTxHvf83SXhrJatqdKFIEZ
DoRvYmWDD6mTuxIG5z1j0hfKOg/fOKdU77wtTZ/vzsO/WC1na0UzjTHSyyYKVEp8zptrDp2UIG5g
faAmlgdhPdEglk4/Oxo1NqT9/4PeecGcP90NLIS6cdvnj48dnBhKj2mIcn6VFCdqWA+1qqFcYS8z
xYwGvGHzdZ2n32lLc8X9+tpFZ1Ky7SZvYPdE9h2eXB/6eS0eQdVaq8Atl5rwotCyw99cr7v2vhBX
y7sjb+galR1V5CqkrCIO/PjsT/xbwiCD1EsjImLvjhUQac97fpQvaRfs4XjdBFS9rmxDsA92tP5t
EVG682yJYGLUmJutzOVtHPXrXdZVjSFw8D02sKoBLZVuJgdexOQ9xQq/7lzEO8U196bbcm675il6
ycDW0JsH46hVPzN0icyDKCyoBF4ZEvxZHuBZW5VQHf7nAtxw6fuvTXLm4QRWyslkfvgwjDGFEH07
wwXijl+Si5VHc5wBHcKmX7WqSs6/IjU9FTfwtZO8WbZAmtan4EB/BOzH4fhKgfuQTu4N0+1/1VjP
o889rvUgeqIPyB6tuloaNcNd+PTJj5M/99y4ze/E0YmF3jb/ug2xm70xnjDKmS2gZC47dsQWe9tF
1d/eUNlRQW3YxJmVt0JHCRRy6JstPGW/G9mafsMxFPkI1lA6xpSNQa2V2/ZGWf3cnYKMLpgYWTs0
/vvni6+ktP+K1dYJLI6x34N/pqfUeCAB76P4QLHOrELPpW1I+Mgj5aQAikOMPLrGVncdG7Ujmtaw
zkQLrJQP9wLqWdMYK5+b2iew41zRbtbBCwh0v2ZuVRKrYipJA+sG77veHGuOzDfDTbvR32fwQT07
H500BULn432nvEURIA+VWRI233smPAcz0OSmUdTO9E2NCkR57YEtAkz2Q0PbJjG397f8PoTus4sQ
PKnrw+rPVo6gdd7cm6rmBC2z7sLMJlRy+AFeVM3ykirNax/jBxSpnBuDW+prA/OanfteudFpF+7b
MFKHG5EZtYlDa5lIe8VizF64pqfAdK0rffATYteWOckfJHBercmBfkwvennXWNpDH3iIqknlPCuu
yAzUhJVFQAR9EuhwTVQobvZoMj1omwutQTT7iXfjUHNnrxGupSS3IXJFxeuHA8k9uC2ZAGowTbnI
tOdv/YaQJKbW7JHiyXpYrgZwbB1DI5Xpu0V1HjYKSLO1GFQXg7mYPRvBcM3ssQEzSQvn9NsFrSPJ
M/ZFvZs7bwSKQJeGJalRZ0nVz8f72m2z4jidy24YioKR4urphygpenNUk+9l0zzgte76XsOPtVnY
HfNQyHM+hvxzytwWSDc6TPg1l9stAvn/dOzMhRc7RIm+k6++n5ZbMyyzZPVUwTm0EIhmk7wWAggY
X51lfl6KlsOFuEmpafk14cz2/mH0ihUu5Gx3r9WLwvf+KyM+E5QmF1XtefvL2yCf+ugqXyKEphI+
G8CCfIVih0ssOCoXitmsCypxDhxJyyZ52Hmv82vCAzhCmeirZUZxEZNZuquVaoqJQyqm7BALOv2R
l/b0muakcVNognoP14H5zLHABelVqZAs5eV27jVqejvCuQ323nV6t0ANRcNwNu74fS+93HJeRJ9f
XLLw5cY8C66HZuqNYMnuj46+Nv/FEYynaOLGDxIJZHQD0xRBXQtXwQ6feaHXVVYnuJ7MaJimqMBm
mXG1lODkOSCtsLxCY+Q00ewdKqdfLxf8fs4ZD8OhzeAtLkQ5KXtPUYLt/PxtizblIvtItG9NG1oB
34TNkpI6qfyGl9ATgIqmQbpEA8bWaLV9mG8jvo0GwhjR5dJOXzuZ3SjP8Zm6wTM5q7o5H04E6800
zFb3lEcm+lOMCyT1id08tcfGV4slmTVJ+4hJRcvxDYoOiea/PtQGaSNMVI5dGXvJxeKEdTJuAhXI
kEdaWjcwGq+9CixbLKIwaSlLbDtwWiE08wRLmah//iOp3LnkE+vUJhk3wgHTPOdjPQGZUukgHsD7
aBg0QSzkLHoAjiNqoekmGFAjxpUSMmhMl45zkOuuCydpKaVpYsYjh1aJ0Ju1FSk8V+9gJOaO553X
7RSIj1KrOal9cOYGnMSIeMHQG+jBeFiJBWo5A5L61GfjGDf1Ad2++xFYs1KsrMEEsz7F6bkaumoE
gTus9M6m3R+rp+ELIxnag7e0UOxBH+kipio+hMtbvEdY4jyb5/t7lBzwejOsDRpulmBl7sA01xuB
Llzm7qafpBF0q6ux+tVFmlhte4iiK4gopyDOx8Vw9dl3zThfxVk9xPppyuQXIj6jcxJvsMz1Lwdl
uKM8dU9ksoOv3GstoeYKSN+YbfrrVzTr3/QgAU3jbBlSYZm5kctrZ2q2VtvKG5ggu/OyHGCqI8v/
Y9YroEL82vyfbSuIL5GXg6vOTjMUg3alc1hYNVlJoXLCBqP3YZF4PeV8ZKB+E/1klN9uQE70SVT9
+8mDN74B7evYvAyrbGKOzqNO3n2dGhcqiSuMEqOcC6cdAs3jkm8/U1FoHK9bf5kE7AtSmdVYNHZ4
r2pSL1+H6StGPMgLgVQibA5K0meABajpC/mbApN6lc0EcrcbpnkF1EmVGNXRO985YKzpD6yUXXMh
z6FuwBRkF7f0cFlg+AahfLQiE3/rY1SGFXDqYlmpJkkH3LMBGdkXpLvJp5lWOFX5Zx3GOlNKf09Y
6RyfN+NIZCPCJ2TnPJIC3rM9fNeQbRATiGZe/QVKRfBOf+YqCaC288+qmq36DBeqFzEab3t2kIKW
L5+xcDnyjIzn8SCmbmTWFbI5FuB5DmBZXTm+Y8rTkyzxtkShFyO09El8nZU65P33F+KaU6xRCt4/
qi+gqsojQfYOvEWK4Z17oWVq1hOzCl0DJaQcLiQhOYNwgvD/5rGFuh6MFqwxwo/7NeJyWxlw1Kqs
YxLg154nRqLxKC8y9VUBKb0cK6itvbQeDb50voDx8JXCaSq22TpOhZQez8E6EKqe8Z2tPTyvLEgt
m7204usjp6uLovp59zkwHY2HH92h/Peh2vK71ybtmrYeno31rFSAy9B8Fe9eV4bKTNcJaTc3TVQY
OY4hQ+ZFLluRSL/D2P5hZ3qb9DigllVvfLE3L7Ie/fJcM52NtN1+iJurHZFgnAqt1i3W/pLsaBAm
lQ9vnD9L1i2OLqdGqc2Kx6LfxYYxlJvJ0Q07/jzsixDrauigxkQP7Y6P91ZOzHCxaOHUd0qrh57D
cjVHMn5PhuFxVuYUicY6hbq5bfDcG/BlKjJ4uyhOl15sWEvFBbg5FSJinAEORKYcUPnz1zypFdyn
UKHQ418HNcaSr/hKVjMN86u+FFfNXBK3oRbOZlGIiyEHqxqigwif5Ly7cOO6sC/y35NrmYPavYBB
RxVEzJZbGFYWA0ch4H5C7n8FXbBatEabIGeXIwazBZDda/Zzfp3mCx3zDziNWQz4el0n3vuaD7W2
b+zsBR0+F/Llx0OD1u6k9ruLlM1VF3zzytQWcuLAT/ucg5iOqRnxsFjZJ6oQLyGQ27jsUgi9U2fA
BdrfJCS7ruLu7eZvkbJq6AB2ZjAdfGwJiKWNiSxbtwsaYweSkYdKwtXs6YXw3X02tue5t+H6sExn
u2rApAQwO+G7ZGh8+/xzIpSLUIFcxG5Uh5bnfjYnDfP5kfOdKlOFqKcPXGKfB4NZYijMZI8RGd+u
XDab0/kOr+t52Uf/i+3cks4W7laZU/SrWgqx6IQSKDNAG9o3OlErsq3bf3oJyL7/JbUgUxzlviMv
5pCU83X2adE5zXlFsUg9agvBpjkFwaO75VX7l9c7VbZdZMcjRQhptSSwZ+NEj8CxOjwWfXt+HQLa
yzISnDN0XKk1WWUK/9jps9Ib22tiRbvXWgnPzyn2HmtjvAcCH4cF96kX4dvY0HnZRVXuJH6f2138
0Hi3V6t5DqO6U3WpkH1FKWIarXpU8+Vmhgppmv6KPRWlbWPZ47oks6Jn9oY69nCiOr+pmfr0qYHM
zroVWvkowx9o81ps2jROFHVd7YhsbyGY2JiMewx9lc9xSpPfvBofZOyo4xBmjst9fpANlEOtCfdQ
f1ICj9E6LYUpX6ZC2ws0TCc6zEDlnGaLbmXV6sCJcODx+kiUgcSHCVcExBG6ys4QrGeFpW6TutJo
1Xc2J/9egTk9D4uWjtOE8XepULxVgwmO1ET6u0mL+yQGNNi7v6ORmz1lFxlhNQzHn7AtW1Pp2kFS
Y4hsZOnWRhfB7+Pwlof70FnVJuBwIeHXt+NAyU8K4kri7gTKmvFP1sp9m9KtaZ+4yrez3VQ99wK8
Pi3vR2a4dbmlDPSLNAcJpZKVubzEu4GAMg7hqm6Hzv0wowytjtL/D43gm50N+TbEdUA4Yqr7kWih
bvdNzR93Mjs3eUPlkIErt2ddXaBfMYlZzo2f5f25J2acPxLw75Mp3apVpLUZi+C6/X8fho/29M1a
APjkvmx/qEkY0cio4r1GEarTzrrbkQ3G9ugd1Cu4XsdldAfi++w0be5j2zr3kmI5U+DgKG1ClnDD
1ju/QW6qTzDSWn3gcSohzABiJIZHOwxloMssR07Zy4HvMt01meeklFD614MBGOltIXG+Y99kDYHN
NILE3KpjGHnEd5Q2llpypq+AJgGywwnOJ17mvs872xzdECQyDXRGVKuduJjLyQ5yBe1AxDAzF5m/
sRCu0KFXQIwscxkJjWLI7BpMp3oFvjQPrxnum04FAbdi4wkWpfiLpU3x8u3EkrQZ1x1DbpflNR/U
Mwrbs/6a2DCdTu/KpAd3GkUG8b1407wJEtLK1Lk9obeH9EO1yO1r+HqSyfEbq8g17FcIpHLrpEot
/voyLUGQrm4DMj58n+xQYeLd23moJtLtmGKgowjuY1UgUMKwhWDKP1SP9RGv1ZfAtmaeg3bctwmP
jw9LVT+mPN+dy9ToYhzZTO4wOoTMm1KZoBcwL/hLHhdpVY8ejnJq0mspVnoXlqBZA6dgToIBXDeQ
j8PnfWD7CMiBJbD+3VelRBnKZOEy0gmoCeDeQEyXvjXbvp7/G8a5TYo1u0hVW7W/GlNwFjfOV4ja
dqyLFIuvyu9p84ywHX8tn1AleKrG5a+BIszSMSFb3XJqVyIyZJoP2lRUgMN5kQx5tgaIVQ+nsndw
cFMpG/2uzQg61P9FRtGwd5gKdukVZ0hj+tB9/hAuYZTMxzRKHEQ1An2rkbJsxhNUeLdfVii3AC1D
1kR0swaEZT9hFw07Zq/q8P37ycbGVTOr7UU24vB6FO7RlYVtIiwK8SyWfCwi4CdQbAJxLk6JQ87u
dorlWYKI3pfEoEEeidbZPdBtgyVC3+kp+rt2o20yXZkhRzJTLEmCBSgYw9RX4QfkmlvlzkYzcysn
UaIJ8MXWz4oYOYVgSgL8BGnqJn5zAXZYC67ThYF/CZV8XNEKg7BtYxKAR9qxFBBAGu4x8r6xbQHN
YfaRwTiPIRPToJ6SGd8rx5AR20Qz4tlPjh4G8ZmvI7kqF+6giKng05UEZkjapIC3+3gwOy6fp3ga
/vge7La3cY7943tIjtMNx2haLhqv+wrBEE+CiCt/FW5d2orDJCqvP07FmQTmBtfxgm6czgxsAADI
xykJhvpJFwmwOeTbhGBqvbIDcHRBrjKPWiS2vzPJPKk7vk0V318FphBdvPj4fCw2lUN+kzER7SGl
dEzGKFO/phA1FjSeOTalmDgN5kDYzoD8rpDooR2C7lyEGrDpj9jYm88WP90bhr2R7dfqNm8q3OiL
CDR9MvuxO77w89Kj1/miNGTfR+XN11qRby3/QIzmRqbju86Fovzc+ZPV8BcZluc4yQDWM1OyghyJ
KNtRIijFs1L9bBtwuX9/fLQhf3fmrd6Bs+8q23i0cO5sFo48XsOmX6Lj221tgpmlVPwfWua5zmXo
20VUwO7UOTWFH9NZNPcBZkEqZ12HuGIA46U0akXatdRnDG3ip4MgFiLVACIiFYfZjgmkuQBXvmcQ
d/h5gY09G7xFLCv7MurlefZZJvo0F/6by9Ax0jSRjfQ80/3eqzTYCL7CrcMMO4PxGHTotzMkuJ3f
9V92btb/qHPv3hDO91GxqZLHV/IlDl9vYpryk3ZIRKCcjxbwsjUJqma+TCBMYJcCMeQPQTRbxMWI
kpaETCer6Akg0Z7X8x1bOxvt0ImoF2kbTZ3uc/qX90imS6TOHaNAg8iWRGv7hQmrMY3iOUrZ8V/p
TFCRhYZCSkUlPY1GcC/suG6oOIY5keDbhbTfAatMcYzOXQzl2Nr2fbe7fwEoRLRYyPETiJ3S2pwq
mZX4dj0gt7t8inTp8aaf91c6RZrlu1gXmOgnwHY6VMExRivlPZKhoHpDsnUp5MV2vGV/t/+IVYSd
oPS2Zm90bA9KcUuKeR418zIpG3Cy9W8RVfJHqLNVfXvmCx6iduJMpz27dMuZTAsZziBmBMkWtJ4T
+J3hv9oZJN5CSUrRsqoMVjBPuzvovz+1X34FtZUN4YWoJYjJlJUClWdOvo0i/+lY0Uxpg/jVj62k
ro1E61jzqBRWvmr0sDjD1CDk+HWrJYIrjuZq8FrKeXkYPDA4T/38gkkrRXxkQVCkAz8iNhsWNA5r
TilD6jWFoqfI60Rb9/sW/wDTuNYMVvzE5L7wIDqAgskBw8qPWo4yaRw1Wm5ofV3v5XpHj426zMKH
3v2RN4KL+uguHeyYU3VKFFxuDV2lGLZBcx2ESk78G0EsrV/PSq8OJIq0sAHhUwxCGlMsrsMsvQu3
/gimVaDF+Xxl+ShO4F3Gh+hc0rKVqw3eU/5iUBhXaJccV18/ebOWMzuJ+E/6zBJaR0FB21qBkO/+
uPEHhf2xcfXOEJltkDJyQljtXJYbLXjb84H1QVdtqsdYh32stDo4wWVdJsJ9T9wHdVMwqLEDIQFA
8qx9pQXn+8ihJUvGTLs0gfy6KMFkEOtxmFSfaOkLbYfDNs2a/MWfKFP8/elCBB0p/0N29MWsS1s/
cNWKRLaPYORjz/uzXJz6gVpANSAwSX+igCch5xF41jpRevY8M76xeVxuhjf5WxGj/Z7JVOAEGi/G
SBVJ9JNeRCnvRJ2AIjQzFztksF/efDkve6TpKzO3hHmAteGj53HIdFkltr5Zi1+QLH6JPI3Bx8JN
JEdqafTUkw8iomXZjYAQAHiFozrbCLcCMkjCkaikMnjRyMnx1WPVjfdCpeTrvnjGA/MxClwHEW7l
Vf0zuSuL9eSsj2mgIz1leiQ6FtqBlqOiCdzFlL3m/hnRPaWdq9l9X7QM6bc1SuIlZZwxPu1AUXx8
+DdlpChymKjM5XlW39BcFlKrXa3uNv2Qm555vjkb6wC3iZZncjKNh54iUytqp1t2c+LJiw7E7OHz
8PrtcqO3LC9dO4LXMSZpJHeD+q3cOQWd/321cwR8DrfhlcxkQBtIK9HnjYnAwX5KzUOKupBK/73u
lg0r4rvZ7MKrze5sbp4+SkiWOOLVorCZg/ODTXqMdYrSIrjS94kUYUZCDPViVaBiBjlYZ+7wGsft
hg9j1iG/n1jVB8hju5sFZ9kiHavGVvZ6Mi/a/Ac/7+M57BM2ItLx4KG1cSKqyEv0kFt6L0S+5xBX
dH2+wviboYYEloeYE1sxijtKaU4F/QwhFhapCRq7W4qVVE+VbMnTA7wHZLPBA7MYPMQdBFvK8tU7
tvRHo1UoV1w7mU/lK92Ki17HsJnujrUYzHjd6Iwdn9LaBaJlb80ICaPfPe7fAMtf+RgHH2EDiTeK
On6h3CvW37XeNfEUMbgwOJD2ZTLLF8AGC8GoVEc0oIhU9yzl7CcAxZVGqlMkg3NN3Ev1xw2Lu75E
IOObDUu2HSAgEEY4ZlrUF9a4UdC+fbN87nSWfZKIlLdY3h5+M8hDx/HBgjwW7FNWwgPR90uA1Dfw
tJQEBVO9/bVMuE+P8X4dOvgYAbLiAs0Gz2h32bsboGvadTKf8u1bXgJrn5VUKf1P8qcAQweu9NnX
ifgK5UHTTQmJkO9wRICGsXiYzZTBmvZchdjP1OjV1SMJgZNp3eUTlp1//6DDlslU7xp0Kztjwky9
6ejrID+Kixq6G4mWRgtiAHK/1GWNAW30vMUwF1fl0uYAWrZ5SNWGIWEX5yrwhNmjx8lZe4I5fMtL
VOoqGG+LmDAuw1AAbJKnoCNtsIu/hWYuLh3UTd1u9RKn/XAwBRWPKDWmTfJU0JneQ+/GhTzopTxm
YfTFdyvM8E8ezhWK+VRGBazmIB5YP6k5gvmXKHce+gNN0Jj/rIJiTog9nmUkZswkFGnaQWQa2ixt
2M466JpKGGh/VpcVhh+oSpSMHTelg03qm+m1jp5CmK7QPqfU8GCnQ9LBQ+yrCi5z3KQK38DTmkdY
1a7HxQurX8eqWeDFjuyn5LoItSwq2nVWbpDExw52Mw4IZVh58ZmtupOCyttMXPTnrkBKkBdzDxiI
6arBEJYEIvmrJnVbMCx3c7q84swdkr82hA8hoDBwimff77x6RZ7CUyW7iojohQHT8tIfNCqsFpWX
YGyQzMfU1ukseN47jS8wxdOSwci4jWKlvJlZ1MI1F0vO6LmzxohyZJYOEeKi9+jXwV4vnARiz/O8
8EHiq25VBsCB0gNCXWUSyvg0PcoZcsgS05sucxdZrLUqxvzYzniPhfPs8asikgJd6Fp1ROh48CQO
2R/5e1TSJ7USIrKxbb7w64MFpaj+bPazNH84tEPmNpR9kfwCej2W5btKeaP43j1o2+H7B8vdrsgM
xGfPASg+Yt7yS4e2eQWkH38pW8yCGTAuLlE0Gz8oZh/T4td21Udcq9SuPLKYHJmMT6upmFS2eSQG
rSHWdV5PC4rQTGu/pxnBirv1n4xHDJl7s/qYbvh5lXh5nJ4zZvZTdfcZPMthpFRP4re9SFONXgRV
esmk1hUgr5HwmkR7RtDnGiwtR8dyyBfqQjDmxU3Ut2S+c+9KreaTA8GRrvBbTGiw0NJnfqemt+wQ
ir3sUC3/Sga5oUrCbx3jnixtzkZBKzgQ4oRG85p7OSytV2j3XBXAfZgNixCWwM8v8F7+1zmlZ3gi
dcq/PUHjr0/sZ8Pqk5sEcVQreQhoczL3fSMqjz+XH4nzBFM8ZhKIgOAN59GhhHGSQ54C0VVVJmVY
TjMkU3yQUrAxaXzbaSzPmMWeeV60PgeZZVblEB4r9GsbbT4EsWgQKfAXv1LpSw6cToX9YLzH89sZ
jxZF00ERunr6SWjrmKchq0UvHT6+wAA9asBNGSyeWVrqKYnfJn24W8stjORsMSI/Gt6PUcCQ+zzU
EfyOi7z3Z0YhkOQ3D0ZV4cKXwNTHLJn95T6B0RsbM0NqGK6B8jovdXybjpavBOdXS+1Ii3jiJ7+V
FzrBAesMmc9llmRVLABDV3yHfCkWnhw5wJ2HcDgAeiAoFeKce4uF09tqHsCBYbezXav5BkYobIPV
eN3rhWEE67ZgbSU1TUw58nBBghdfimZMqTa9971v0K8Psc2xsvwMUu9YwzR9qD/ztyeCOCJZ6ffL
I93JJrRZihwXd/H8BvXeDGs+EGFpMCiFDoKe7jrL+0x9ai/4rHmORlwSjjbr1lTkgyBNiT/PsJVi
pS7DEzAGR1/xE6fNjJ46IDKWnk8D0QEqO9mcC6FJeC3su37gnJpHJM/Ak6u6iR4AGt/rAPXFhS01
5hilTrAZrpdQpeDV0zcNwUEMqPwI2NkL26ogYQzrFSAEILKKQFBECkPaG5qB83rSzVdT+gkqCt8o
SsbrxSr+HD+aJEW0RozkMCLQt6c4kNarV/E5XG+eP6Iet5VHEbTSGo1LBfwIBSxOxdQpSSC/HrT7
3Php6vhbrW0U7Wx0WAZsAgKatenLH9fsrg3CqPmpl/OmQk6BeK7zD5QBFBZ2E0JflPViUPWLa/h6
upHP93eQibHvjhKo2l4RLqAu7NanyWn6j3S9M9kR6kDLqx0lsTvIOEYF3YR02GhLIUnGHdl24Zwp
+JCMnBDLKipFvN5xv7kGC37x2siRZ8GVP9cHKixJOKT+CifFllMt3OYomB+Jg8Bkn8YYKDD2pu/O
yssByLh/L4OxG5J9qKPj+580MA1O7jhRHEdv94I1j7xMVyskNK41wmEFu3pCf0CsVvKhCJXlqAk4
U9tecR2H80le164znibs20IM8vW/CbrUOst7vkd09A9n60uIgAuzj8Mx86wWC/EFlZ7Gb4Ulgp38
wkHjzwd6yO8MORF5YMuD4F7crNYvw4p6O/kRiF+VmelBa3l4fgTZ5KUKMMV5QF99UJHhxiIsL8xg
ue4+AoLfoIvbP2xoejo4GY+V4X5nTudipHS9Fyr058mW0UcYI2iDr80ML6Fi93Srrtf8j67EshpR
x2gzhlVm2pLXQ2ldgtYTAAz/wFeaLtUHcltL71l5Mt3hkJzEJXWo5lVtRimS86CKUpdvIl1fFQgo
zv5bimzwR9Nuw+TEVm2tuES1/8m5JySw+z3kwbNpnfV3b49TIHWf2QTaBTqH5eKdaq7T7OwkID2q
BCvCh1XuKL5o08qJ/veQxEvYhseZgY0jpmAbvNkZpOrEYsYwfQ8cMXDZrBnodh6AWDzNQSwmsw87
FEDo0GSnGNdX+4FuE4XSQImgBqkFfBucyVvl2cTeS7B+KEptX3Uxp9EtbLUcmDB1TB5edSEnH+EJ
bv1oKL6zjiCtJBvHrIsBqejIOBIfTU3Elwg+FYCron2tKHvxI4ONjtzUZWorXR+BL3N9+biTjsYp
gqCbFmMeqG52qxxFPWHvfiOBvvbS+4UFaUEEyMH7HO83RN9Rkf/w5jONzcosrDUgT6FwoGh44NlC
Uu+IemUMwExMQ5qdrETITr1CrFVpDytKpwRj3LXYO4x5qxzTDioRxW6kFYAvG3qPVvUGeRXzr3dA
l95V7q11LwdGVcRP+UbW+iFdiaspcINNx1YqyAwEZA24k07mqRlTGLE37JoyOlLyfNaWo4rEyN5L
Hg8ndjX4lsSNTuJt+IaDoQexCPAJ5NOjClOH4dn/hLmhT0k/VJG4MEusKCGlYJJsqSs2ZeO1miJg
fBj0wjJYwRddaUk+psHYtmTKLbLnQ3I198Gl/ci7uSN4hhz7+4oJRgqjrmbRxoiMLyVGox62AVbn
4NyYOl6EiDtXQlOXomJDYC1GTweK5FP0y9qKLoQ707mHLfpt2kOSI5TwSciCq5dp3oHyew35/sCD
wgZBBAo2bekw95CCRzR0O7kIgefnz98F7nRIsl6fo7xXEF3BoBIF33szhVr5t/Xkvwgeo+AKm9+2
ge7FRMNgd07QioI8uUyXl0lxyc6bckpTxb+iSK1j586XTj6wDcRy4ZkNE18aXJ8gQ/L5s0kv4ZC+
b8qpvffl4LbRs+YEWSaaMCc2Fc3JAV57m03HZrBDub1Zseb4m5JliETN2/A4Y0lnrg5go6BU8vn5
0ng5CJ8VOlhv3zttlDjnlGwSlbI+uzCNT4dmUjDIOJ4wgvXmFhKhrjBp6hBhl5KDQjtq+IVoktn5
eDtoTIAdJM0OnGJuVnyeQ0uq2txAD0aS5DOEqkC5vTX33Vy8DL7ioHCKNNu05uzYUnmq2Qx/9OwV
aSk/GKqliLWy+clbU+XegucjbP5FkYZXoJkHCU/CWmmziYZUVHCCJZ0ESzujQr3XzPxZ+vfNB6oN
XhpYleTsWt+atAupPRp1GigaD0ZnJdBJCh06wyz4Fl/GpR2SmEhv7nr7gYHp647C0bvPrfa3EzdZ
4WKX9Na5mNbzARKtDeg69JEPlOX7uvZrDH9SLPF6B494WiN5tkZWoywrtUox8O919KozAa5cg5JF
SvL7ucm18qoZrrqHc1zgBHpI4s8jR3UiTguL3VIp0ELBot751UxruLn0x9o5/GLrASOZtex51qvh
neWO5jkHebOnIgBWoqRvMkDkmJD6jRLHx+yboOkK7wNsfqTfWHnwdeywPWQxS6ECuG8TuzX5hl2/
8B47Krmmjqf7QoVNYdJkPBQzeYilnjp1Ii6rxH4tKLsC52HCNtwS+jc9dFFE4Uhm/JRO3ots3pBh
TgOqBujPy7cbQTbwmHRf5Wda1zAnRQrHJFJrmRylln+GYpY86fKn+2k1tns9nSdk5/FMkWUy1ixz
nYA/GOrX+B46KbjMsmwkzLT6PFTsQbOfa/2OvA80zd36KuoTAKl9hzfOcQ9ozUD+vsXWcNWKAIT5
Kbn6+VQIz+r28y5xzLzVAWEMFQBwtx5WEjXE09RWvF53BJESQzbS/uHIAeFt67msrpzZJBCwaEBr
sZ0ll0dMLFUfm+CyKhl0S9NdLCmd5K1pUC7FwrHU/bSsqUZj0gBZq10KqcJQ9/4cpP/HauYLJpaT
rXmiFp0Oj97uTqJC59qsGThoX7WA1eqdtuAbcOJ2xkcI9HvkBXxhtUQ9UK9qwQ2Ju4fG5LllpkHT
0gxLU0YB0p6oCU7Piu+BqjPc7Cb7G9qLmVS+H8VyuWfAFdMFPItOaSLGoCkdARu9zc0tMrPknp7M
Dht9NbPhYg7dfDiGb1IYvL/njcCf9qrSWYNEBi2PY75UjZmm7dyWsiwmEvs1Bl74DBS1qDyP8tCO
DGixEnibXbH+qmquCHp6AFEiTMXguuZKjyZegDwJ4TaYlKdPrJlmgAjVWM9adHLO5nxQimbs4/HR
ALnqM4D4ErD2RI2NEFfCHZOUa1z9hOdsPHeHQ6wK09+itgu4QFEq6BITAlTWAqVXJfbVNhYKquJx
KuU+wzSyePDiuytnlpdp7hCA6P07DGGreZAUhiwmpPFPvVQqKKUndVrKxCcNbtl9zI116nTMs75U
IF4hU93LQsKjUzAwXcK2/UNySpsMztOhTMSXaHHxwZKav27g/vOXlwSUbYPHPQnV8KuYJOqkReIz
Y2V688anqeUUjLRzxcNSH6rUVBMXHlc/J0r8E49ZUmP10Owi2b5ukrij2BoFVExeuRoYlzIAT+ma
JykCTKKB6ePh65mlOVc8bPVjqNldI4s18g1XDedsewp0x61QGTIHULi0S7WETOXd3+01T8QkQ2D/
Z/j3Kcj+t9RrAsj2/fjfQRp+N5U5PIb12Ps6ZOX1sH6pw2pm7E6cejIsYscWyFmiHVLX+kTzALSH
s4/hKfta9ayh13IBVElg/RlbSiQTjBlOKQKvwTpGvLRRsdBtgwUGZwiaU+bjIBYyd8YF7BUcsLaP
kwGDN63HKSzHFhMzKNnaXiUhGbFVPa31AmMp2l5O8QCreTDaeG50Yae/HiAxvA3K37STdHak79aC
wegyJ0sj5S5zY7vS+Wm98SUaBHzdg1XIPjmTGDPwPsAhDXvfYpXsa7uy0f59g34CAwFzr1hhjXVB
r+CX5qnp/Tr18naRhT0ztcB8Qy13Kz6Gr0xYV/qwxNJTJxx4S7cxHU8jp1mlz3Lm2VwYICjUWvNC
2ZQlYu/BrbvlQRpV4FQQ3c+uw1i9wk3v68YGfN3mKZPliMuTavn8wgtW7M7BoBeXIkNv4RawCz6u
yHmLyxE+oMJokl6aoyR159azoPt6BUjc+rJmCNu9ohoVj27uFv3rjnYo8PpJYoKVy6SqEeIwRH5O
nnO+I9LGHePcViTDPCohGhVmuM/3QA87xouMw/g7wZ2q3ahSMIdjK29RR2xW/EHXUAtfKTS+u186
asCYBxDJhhy4m1zoObMt/sHzenNLUoVi3+/L430EVoEq/XOskHhMQiTfrG9GV/+SOlNghDrMDin7
4k8MB/7sUmAHi6fQ3BJRHuffp7+J2aq/3eCv7DyEnxBEHnKrznqV/q1FlP0R6qDuRpf8WqyCZAVN
FurrndAC5ekpNhq+ENstNxCgVVgCnARzc6HD+zN9/RRpGweWtNid9ELqFMlowMcg3RdhRRZiBboj
A7gRcgxB6EYDCGwqPh0XUKS7QTbSowBpto0oJVnEl+yHxUwr/e2wF0jTEVkqKxrNo72HbSLZl9M/
0AXujYDVldRy9eHb4W+ctNHH8BVF/8qXVlu31sVP9qaKI0x6+pykc5T5LDbryYjrrwgxMlzgre7I
OJls+36suQcje+xk2cXlSp+ZUkHxh3o3XdI+nt3P+n3POTSGlEOZPJy8pdr6T9dW16fREV1R6iH0
c0RUJm+vq+nXUFxNnsc7G1fRearYMtT2YR1reVxSlJ47PZHGs/trDaN2DXSoVYMHOFebipKp6bCj
c9fgluUzmXjW0aDYZMfMB/TbSKw9M5E7QqY5ka9N4i8XsqQvwlBATd6QomBo7OpiVJxh5f0x3YAe
04ktw7AEyWyr2DpgfrZcfj49unkRwWuJTzGVsLYkH6EwPQvNmHiStM86HKRjQnHfH8OjuQt7VmIK
dPg3untMAUSKTND3oUEf6/w3F3Ug9zHcXFAPVoAeIQ4bqWyoDYZbJ3ojZFpTjHxrnWzqa3Hcumkg
HNjF7YoxMdkKwJWmyFlDsNW339zfvCs8QVuPj4ctKMWcNKMiBoXqGkd73Ld5SHbkNYTQYC2Kh9Td
QaYYfyvoaugYxA+64PqCFEtwGdgyeDtBV6lry7daQ632zgnj+qxzEPuEj/sTJQWT8kLKwOaLM5l7
qnv9cvRfo8MaBVNR8CGMY061dAvdAMenm0/gqKIhXXMFTY1gOXnGjJ5lS5/UhoHQ0UwwZQ7x/Z6P
7EAxmH9vwgVdWcvH+6zAcAlF1iceb5Pks4nLT3sThvbbtU+b6Q6AMDl4qdIHiJo3xJKtP07kjwNN
CgChjyW9KW1eGhM9F64cexuYU+HQWko2hplhkMEeaFPAH7Ahne3ABPTkp1u89TEItMDTBeH0Ucm6
DSEjg3RvM+VHe4ji7ll2gBIb1nbOb0u8AG8sdFQTG28dEP1I/qxYYmAwmiBZ78q98dKREHLJuBuW
SHh2V7JpkgKCOKqHBkmT3J1c+xfAJIYUVzOZLhNjQEEH2YrxZbpGy1Nc32UPpVPCzviiRDQCMnQY
3kGeycjP04Lo4zyMh1RlqvNgDY5abnnh2NV5eH6yQus4m3cppUyKB4xzlg7Yduf5w+yQ6Sred+9B
1clNO7x02Ss3wJtv4XZiT9MQ1h628M/o3fMEMI+Idc5wf/du/TQXMxJKW98jP1FOoACSs1OWGB1v
65NXfO3PSMNyEoXwWqv9n/MpeWUbsPn4lSpI6rbICW8mW3gJKyObhRf+LWmln3zhk0VmdaiGZINH
i1wjmCVY5yE2r65nq5ySDewshxl/GR3rQ3+Q3GSa4fnCU7cfMMs5lAkZjMsF38q41FQ8VP7M/fxc
KfhG9B7MiRhoFCJp4H4JG6vtYQZxIPJOWLklDYMY/zrQxSK3J60ri+ZH0PPW18wAPgVswR5qDjyo
PRVrMOtNXAuk73OqjBTAn73zy6FyXDbZzz1qA+nqfw7Xa7byF7PKB5ozzVfWF2Me3DdEnCeNi+T0
pcVRkKIh9CsT63XdnoxOMhAyPCJJC6p1KMLK0UZ3gePC1jmseiSdJpjLkAunGH6YMDt1Q/3dDFt0
XWzMbyx/WdGaQIOFk0jXBdKSBQ4VycuJ1DnGY1VLp5kasr3gSH7Dc3WQK573QprmD/fjRQV18MaB
84Y6i+cajGX7eNkX2CQa8NJfsrnasCrBvucnNWbyCHbVpPUoHQva8Q0B1kjmyO2tBbx4DtXRa27u
Yp77Nq2ChbtkgK70fjPlPEfyjJDmxUlMHiInC29O+f2nTmkmZ7sAbjWEbfr07IyXTdzpMISywdUs
QYsVRM6kL1pI7L3bcZm3tr815WBZtrw8tTjf6678bUihNUgmmTOs2VejgOnQZtIH5iYT/K/ggoBi
s4j9UDQVAE5aJpBi1W0rMWfN3bX8tpUyMhJd3l92hLnosDhWiwIoxVz4DgPnp6hbOtu/6QkRRVWr
sEP0dcypKxz43k84a013S4Pc9U0rrbEDCOBoUxoaaE70RkCZ2QwJR2NjwAMP7YszfzZ58ChTU1je
t7vZIrazCQoZs5ybw1WbnUGerHyaSnygc6dh5HQPRXD2V/WBI33hf4wp1CfnPGtRjDwnVR0/X6TJ
ihWgYEp3Sx+6jEodEfZkjYABSNsd6B7wF2in61I0Jbujn7X8y2kzEBQfdnRKIFEQEiknpjMOD2mf
aF9WzMem+VBswrAtGg9CEs5XtqozE87jzBlelUpqfpPkaGDKCuKmd6fnks8NABFERoW8NHFsGv+9
RuTEb/xjY5FA9H4MLqgtQIYpnwvMBU6erxg5sntb8wMejLfePZZm3tJpITMWUHNueFvoq9/gBBpZ
wZZH1ehpB2O8pNac2MWoXqIG5roO8tYdz3BnePv4xYRkkWj5gGB5UNcVlXao4RtvchpF5k/SMOX6
+G0TEsmCyn2mMpKv5JfVAe3EYsDl42u9aRC1vNGbUuowToMKT8h7RIuckM3qDAF/VDfrDPjYNHm6
UNrjI91Z1Ahmw4Mopfp6ixP1kelMYx12GblvIWTd/qBWvvD6SaT65UXmqTxZQA919UU0VbvmR/2K
/Ad4U7lUOoHHvd0Xxv8G3vN/tC9SMoGaQGEZctTOyDdlj3wEVDb+ZQNXcNWLfsQ3+3kic1yJks9c
gWRYWKxhCKvfpwWD2th8OFrTRLIEvfMiuh5pACtR8wh//b8Kvml8GsP1oVt7tph4VRFXz+AVZ3ED
NNpZviAeL8/5kce3q72J2O8TqgatJMaH5bmXQ7SSg7PiN7UVWDPopC2lGd5XQ4nTO4zx/qv1mDjX
NN7vUulG5A3Xxt/C4WGZ083G00XaOCqRzIELq3YT60ThMh6wtl645p5n4pecg5z34/2/5qVNTGH0
yasfKWrR/zHU1cMUx2IAdpKAxhQqe07anfTIBf/wvwPnExl/m515Rh1d+RKlKWcEda14gY7VTP1J
yuJPSgoiEXmw+f+/Ev0zYHacdQIJPS3FqQ6P4vMJ9Uo0MMxf0BsxdwHUDOfYazAsQ2yef77P950y
LzYQF7RwWwsA27MIEHcFpvPZUaQhC+jCtTjTeq/f/M0y4GVSvMkymapV/a7WYe4ytv89tGw2YwVv
/zaQCj/usrv83zofdq5/+4/W49NC8HlKMT+i02lwjGgmW17mYAx9aZ6p/ryrF36RSn7r2Usp+Ab5
UOYUEn3TCI8kgrdpq2Mvc66guNxyXzPONlZqNja+2rzfeQxEVKB26dQRCeWg4huIiAGF4nOpphCr
T5nN6pAXaamE6R6Pn3Kncu3ZENlWTYugEhrg3ganCtV3mbQ0YMqG3pn8Mqx3nKuahVfRtuxp4S46
QbxtfhV/L6jnbyZ3CLo2EFrzsAgLFuA5sSHKRUQpULgucYOS6fGG3CUKm7Io+R9unCsIl8r8/7c4
fShZc6uY8Or7TZCpq4IENUFDB2yootfar4GoHeWpL7QtHbIvlcVxlvDy0Y2Yi0iAOEynraJLmnYB
+T+3f8C9t5VjCWtxL+2L3cZO+bFO5YP3Ha5Z/awLsQg1b1Vs1Dxl6jA8w1MDUMx4E3kfwmREebVA
mwigza3WRJRIW+lD8a5mugq66/oVKCsy9FvXv2iZ8ldozh9RyB3gvCQmXZz3FFsVbDIv8fUN3vOj
ybN+57Mh36voPTr4mBGxRWSSyU4UB9WvMOJPf6G/YXtZL+/ueSB1UoBmcgISOMlOXq7DqEK2VW87
ik1gkB0smlF95U3LX1jkOxVP/qCVuJ0zvgkoV2EwVWZgvOWaYvmye4nQR2B4p6P/oG1tZbjuNo4h
2UQSkRn4agCu9yLlANKoWy64gqU9XlPnqiSFAwqiNyF7pqs/d4Tv/y1/KUBGUdsVAWKbK9eAiUDN
S12SNMWj7sYaYzb7fIl+1xOx9MZOv5jYoa3wJ7Usvl3jXqoPr7gL5DJzA4vkLHg9XXr/0hyxHqxm
Zdrh4BYCX4ecZjv31jbXWGj7zLpZ3sACViJBJgmZeBWcvFecKC5cBHpqOAfTb7U7KbdsOwyuiHj7
5uOJzLCoGJqqBoIfbwAYEK3g34Y8FO0d7ECZsSBtW6sJGk3O9fG7NoEAcLr6VmgPJlSZVUHTmDbd
smFIaXNDlSzpuBbUYb1ytfMbhW6WZC4HruC0vcZruxFD0nFF/DeUv7EmMgkdZnfnLnXQoESAV9no
3XWWIlkKxX/nQRkn42/ffodJA1QDUySKA5yvnfo9ISZgAoZz282MBLvgUcefmn5Z3XEMJ97RMoP4
XwwMuHjiwn4+XjAtHW+m+C2FQFJSn81ZpH754OVD6THA8ngXm/8oTFWla7Gp2abNDPix8PoECG/h
0CAokfgJzkQ705krTHBYMZt0rstI7Te2K+wzK0bvofIKNl+6R3Mph63mGNub5JXiil20cQbJudec
OWEPU5+cmfhrNbBs400gVLFRVq01p6iG+wTkTdPmEoQLbticLWC7G559ttVsFMNl1hJyCZZIRCwH
AKM4ylERecBZkiJj0MXepofZ35bdLki1OfsQbaiptnNehgpEGgd7bJUj1SI/gUaUH214TOIGXKVT
iiP3GqIKkjqGn682ZnqdTsDWwU+yNjI5JbPUgNl5XI3wmImRs/IUgs6DlHp71cblbgGY0lkHvwvl
aqWKLwoOpY1SdNId6FfG2YLNGaZ/JGuIGtVQ18eaEYnVkMoGGw2/mUg6j+wQvqhiLRfwFb/0qdgT
jidSTnlr9GWEuD5UO8XB76dsPwaVZTmFKR8KHwautHv6rm2O8my/YD6Nc4OiX3XnQrcQ9W19IAZq
Dp3uqjfuknbOjMQzjzTwNcbEOXsfPdwWLybrnOwwA0ZPNnB/waKoLUfCz2BA3qcjYfh2aELfFNPy
Yw2aulONZFMYINZjs0ryRuoq2Bc9BdEsZuR6e+8doP5nLAmB4US+LA5loqK/PXru88tIQo2Ir8B3
h5beCheNRwenqmdd4ZrhCXe8cS3SEKBfwqRBYxtHqjHQJYleDv36GUmJ05B8EM3PxrA36sFcaae0
fvw9wbLAW0C7HQEkTx69sEQyXMhAGHopm62QqKAmVtUYhfXdiaSh2vWMo9JTVjW5UETQ/HKrDdCe
sFmbg/09AyIHbMy/BKgpWMgCLy7df4RsUpo7yLfenFfMqHTo3PiZxokbJ3zRf0e8/8/m89TQdI0j
k35KhdC4DVdHYOYYkZZzpEykbeSY/spuOlFA6GSKpgRiiKVKNAQRAei8vlNpF2Rej49vl51CyqfG
e3gCnHU/5tZbW5XqVl1OUCoPrbixMPbmKfVgcSXtkXgWbb/sydB/UCrlmhSVuS3lUo8kZlVV0eXX
dwVWbOvlhr7h/93cAnkYdaE0bGXyktL8GrqbYSYJm+S2JJq7ZUhASt7m63fgGVXJEZBAALb3ZKv7
e8lsReL+3bS+NsdRtwwb1OXC/0r3ysdFUJQUuEkJ9bouDGTaOIq5AcfSdqpszujDJwSBaOe13L5D
g0hYq+O/SCDNsZ/XHCbgr0+hRV468qZDbkFSr8C3mqPNA+GYnVo37M+uF1giq0JL69VcGA+ZQRhJ
BayYivXwVCm2OdwuWi/+x/wEwuKFAjU8FD8WaQ2QQ4Kci9JU6cPjzBIx77DZoz3NpShRXDtpwTC+
HoAhyGb+7hyqiczMY7yYscPmL1Vqgvs8rSbIfN8rjdUz4/D4eGSIisOHdn5BBmA4PfflJ1y1V2Fd
Ki9iqcudppb5HJqCfV1ac5agE6ZPcfEPHU+GoQNPHTaMoO9LNYTFM/UhsDDpe9u77qeqMhQRYKC9
H2Gd1z0P92HQwvSdLUqpEZnLTMB/TsACutrL8mbZHGT4Xx5ebt5YWeN0q90BXHw6FAkuR8dn/t4o
UHmHHJmsvFmcnNv2N8wp+O5dfkle9JPGumN4utuhsMxLQHd65P3laUGR0YRdzgSs0UcJT4wiwWb0
knrbGN9JsEM4ZeufCHaPIKxpr7WlVz92HLO4AKdKu+2qPI8yBntrLQ3FeC6LTFKGzXvspIFvL/u7
N1yfgZCeE1AYTePjoM8k079lw0mjU3/HNJ46NgM4H11f3SNdlBTmitgW51wTaJejU9UvVQj4w8+j
Q9S4btrJByMwjD0vHBvwwJkKCrS5wg7MTj4xVaI8DoHvWkHHA6Lz6R6zVuejUPfOPzIxeDVKT4kB
NL1daryelhdq9fouIOAR+vaFo8m/M9fv+LoBI6c4uRwC5TFRN/WYDLaNaF3jFKe0ksPQVd3Yywze
QQBpZLrR9E4Z3FHydaO83pJmDoXwGzbAZt5XPAdRl6ZNBJ4t47EedsFXqRXqY0sWK7fDmQ380P0F
Pw77sdL2pzQKO2oRjmgCElNpooXX7oS3Ey6s2zSc+d5g12kRzGqv+CPiPcb+cpULdJnNynszm8L+
IMKHY2IsKy8ZypN5Pf4DYPoRwEEArSQQ4y+LYIe53TvL8JSNFognKmbP37STgHi7vcQnbNDrHi1+
8aiKA8/snpSVf70Cp34UXCeQcVC44tfA0gxDU0NuBaqwL/FbQzzB01rTRegvRPjVlqvEh4Im3XaL
Gk+9o1d6elMMWRRxqPNjLMb5y7qzhv0CCcpzT2mYgIS5cxgfgqZ1Le1jVW+mvCV0UuibkOUfRXEe
ilN9SSTT7N5F7+fSe6+SEw3+a/7/CdrGNaHSdCxQeGwNIknhes5kDrd00UvjSNCBxxWup8+Di4EQ
UB0a1SOpmkskAGNiV732tIXYxo5fjteJycV0vS0dzYF6XCCfDzxbsuZJEJMs3H+w7amzP+xj9Ppj
c4S3FVvJ5+dY+jQVhWm4P/ftGXSTZp4twBS39NBb8hXK1OR1l5yIimAC7u3NrGWDRdGAGNXF68Lo
jT8WABEAdArhQgBBKjcGOxnsVn3vohtx38XyypVIcI3UvFXtp/02bwp0SPcsK/UXxk5/zXoV5XPU
ZBbisYGTwNiIiCHrsEmfEVCewsXhxzMQn0FQ603A6iLgoCGuLewhMSx112ejvI/SBTFnKZiyHPpM
euet2dVAsrWgE9XDhwACC8YMWNPzTqrPU0w/thXL9X1WB11+RD6IbeusfrF+28gqs5lYOgjTQX2A
JodVn3p4fQQOf3yLFyZdte5MR95h4i//eno3MjIBCyv0H5yFaeZ9kdMpJ7xH0I/Tno0/8/Es2CFK
wOrW0k8wdrOcoVjeNMfUK+M1thZHAkRzLCNfgqPsFL5AjlpSAVTtwEAaJJYy1g0V8jY2As4hCkrD
0NEG42KOW9aB45ED3JJp+TAmJYaHsFl5dpfLhDm8zpiJNtrqm9Kn32RKCqHj896iuPO8oMZIt09r
ok1YFc5Z88uMHy7qZ3fROzrOCStEfij/bg4J8zs5OiojMpXkxtrjxb2CPlrirxxsPcAN3v1QXZi2
OmC/FrTHv4Z5rpvwId2cjOSqr4SguMKG9DROMUKCGMtwTwe1KUswsEfMR3QW+a2/kFzMOqHonLCn
dj7zAQcvhw7K2rs5CMjoLcJH/+P2Gqnf5sApvLXg17nLT2hYnTA87aDhCBpkCkMsaJVlaUpVUxka
me2dOAuioO27cSc9HpvKEIbIo72s3NoE7EV6l5Rq8/pc09CJEm9m8r6OfNqs+1rKV8zeQ+FDvbhJ
cOVBvyNczEI5vwtsOdRJbZSN8PVIIm5VjjG6ZafUh94crqdd+PrzMHEXOuOVby7x8JAd9STKFxK2
MdreHyeaxmBHRNalcYSIrkSZerOy+U01aM4krVHQ4iGuBu+IXvvZh/7IgqNveOlqlNNkVxJLvxoB
J9GP5f0abMlbufmvYxWQdnoIBQstjgGiGvQ5oAHN4PLb37yCwo2IJ/FEoyS7g5BJuHAW+cV6fMAJ
q3BlQbrA7BIWhoV9jI4U6J3n3uAAaGL2uxCOnsxlqcJrjNLTqLRHKJMBTkOae5ICiUJIqPylkqDM
/fe+qlBXzasN7ZGIirGzcAFoeZpdDSRfPr9wZuhma/hWtZSmbYIkbW8KZmf+K9Znu2/2EAu843DP
8AV273rW+abRHwLFHTZ9Y/g6f1RFRHzO3VqXrPLbw0wm6zweafe5B7PrGytelcEFv8ElSbxkrUGW
FW5RgR+yuZ7QJApkQZSGanPyb1UdVWS00vKx2ug0RK8xQyZeIcf+hOkuHtqlYWWREBSpAhHWvGU7
f6Y376npWKm8rfLBiNEUk4H8yWkF4LTR/lavBLKejTdSWr43OTYFITDdLMbnPs6F5/gBsHdK937p
f7pUVPv5/ivJCWkADE32SxpEoWf6qjVKSdlg8/UmCUKiAXCMWTf0jV/YIC3/DCR4U11ix29ssLp5
9DPz9SA9TvEw/GiLjRoFGu64SdQkips+OBXvUgbYzTJrEQvz5PBuNqpPtymFBKs7X1xxMIL+HOCa
yEw1+uO1XRAzFgMpvgQIuqWyhoohpsdkq6G+oUdaWMPNw1d0vYPRr5HZ8LvIKV7JLHZY+ei6KcpT
JZSYVL9TODs3vf22d2yVnBVrRXkY4E0JBAD7QJao0CH7sU44m5YlB6Mne17ZBZvDUZG12M5bGoNt
lywt1HvecnTkSE394xyq3JP/kOcmF5VbpaOVksIgC78noOyKQjlak+duwpq7ltAkxQiH6es15frX
/NMtFhHU8bfNQmvxxEekCFdb+6+vEcXZUQsf+S0TsPaYsDwdd/1DjZEcKzM5oNKyX3cMUrA1JwkC
vxG2A4lkuNBFtiNAxBKbUA4S22k6gd0wm798Pdcr6MfMoF8FZD8a+ogVrVipFGlgIQFJmOQKn0Yc
I+HaAT73+UlUTjE95OqTMDLJaGK9O1nJ92CYm0sk/VRhWCJky3SrX9T78FGEu/+wLLarODrWe9Jk
veAJMNonywvJ9JeGbcD9NbgSIPrLd4k7aGT+7etLgX7sNzSDXd7u1DcIXCZD8KSEtFv6AQNYmVv8
pIbHQC1bTT+s5VbEnaDLMb/RioKRKmEj7Da1nu9oNkYb+mqLR3jcljBh4P65cu77v7xN4Edd3741
TBokfIlIbhEh5Pd6CqHLCrgiUPz3c7DTO6HyK1DFFBKkDqfY7WVrX9VoIoUuVEkN+gNGmz0gIDOy
F041jcz/lglcdAuWzQmJsTjfHXqy8XJA57PTwrUipd6YAAgJw7swBDKmrmgNC51Hlcb4goXhSjLQ
+3iveFjl8ee812RN2E5iXks8bnP8y2QvVqc3Mr9ATfsjpSjXPKifqyOeBCmD164DYQ5c456Rm9qL
oe8qZvTIj5IDj0HTVcHb+zNnOUgUZPy6OhWObQL2ilzy4NHeg2NtIGPAhTjVebUXplNTfVDAInHM
oTg64p/7yViDFrwgMzmqaxfCFVNmZJNVhw/Wacfwq8oMtZHsKHgHdjtyWYG998REsop53Gc+PrUa
eFvbTFRMGQUHjKmrVq++3sNQ8qujrR/Ofdnqz48eLAUgV+0p/fovgaASpVp3ntKcuEaMHWs+11i4
DrzmFqD6LZht7W+QD1hM9lEBjhPDx79/q3SeQO/SIsYl5nyKJ/lOcd/Usw7nHfCPdDUZcO3aAxMe
0RtZWMNsXW7kK6zIWGk/Dz6nY+RJKAzF11WfBpc79d4h/MPi4h7HwFbo+gmxRq1YutVM3UrFwsLP
1gFG+KrYISMimGx26siE1HMCbmmsTttKw99Gi7dCiNPImjP/ZWubCOVuzPHKXhgvzDSv9sgihAg9
bwuwB6epnDjrnanprSL5m9MiAZPYPnB3WCdtT/HNNjorTN6y2IGG/Z0HxEqzuSldVYtLvN/6ORlP
uqAuLnw0t431W+Yxcje3+fbhD0JAfXg/99Hrjr05cB8bX9QbJJ7JxnUeA8Z4zX04ZGRNkfMFaKj3
vAIUYeqHS9MB3LOYnwmEKF0e1sWqWM00+z88ydJ2NBvMvKNDYVGlNOQ7qQqdAKl106yQsscgOyiY
U96xmQ1PyuFixmdK0w+/k7EZs0TnFT9KioDt6Uw0uUf9A5zpcIwhrNI5p/bBXuwMpuqvKyLgENVb
XtrMXnpehB3HmxrKJXAWXJppUttxykOJLWw+gD13UTJvDS/LS58L9Zt+n8cbuE8yVe3/++D+SeNf
8ATu20dn6J3UW++IuQ2Wpu5WU3AjTFpnPtou5W2WVeyDhaRp1i04/zcPo2gSoUsHann1yfx9mAWj
UO2Ht9xr/sS+GeyMMY6kopyTj46ulBrijT4xOTuVJrX0f3ZGkRqw0+fp2mP7JTWgZfXvL+P5nnDD
B+jktv0SQjvOfWY52lLUXZ0uEddFnUWv0LA7nkrPZc7UrBMgMVZcdFV3M7Iu+U73hZgsLQDkzyyu
ObVBaiF1Xm8wnF/K/h4xi+ih0oM6DUuHNwpva0FbS0lkYHQkftVtGb8d7bJDtI6nF66MXnGmPr4B
VO5hUhDOi3Ce8eTDVYZCYaIMOwij1zaqw4BB3fyS27mUnhfrFc4rapNkPI9TS4tO/7uEnkljoTxi
QYPgrI6zJgELhW3GQpezOPms3yeIJecu7gYF84IRFsfee9s6wlQgX2EiZ5GwPYvq7w8nf6oSdu6I
bR+qINpsbmd9xCCGhk+rUI8Kw7hvbPluXoGQBl9Sa5+odQPtbuyftMUDdNTciseycYE0UpYlAt/a
jS+X1xEErb8jqvt225aDNxLoMyuv/xYXHi0/TwIZPE+t/BoFD0ZY/zd3aySNoFsHBr2+U37549on
IqPtOex0IqnQYo/Mwt46SC8qb1k4a/oXP+BcE2M0gSeFfgiPgoND4o6cdMTPcN+Dwv164Cecjf01
hh2vcwyHZNmlSNDgYAUXxSzjwJ3G/Pv4gnBefWvMKWHc73BD7qkf42FwGjoIjJxQZytxnx4Jp38E
Ftfz3RL4GV19SW3YsxQ/3gg+27Id9ZibWYVEOQN21CmDnM6zawIAs1pjExQRKfpPUzkqRTF4L/oM
0b+gOOiwp0W7u+z0nS2YC1WMj7osMOwIx6OLgNaMRzan7M9sOLbP64E3Pwv4VXq7Rr/thCltpL4F
8c54hAUKAnQ4+GMKciDkqavL6jPLsHJour/TlYKkcLez9CsDzw6zEFHCOLTv6Qa/jirZ4f+yjSNW
omlKLN4z6UwZxvItnpJDF0gqsXa+HP8Tye0ZFA+jKzVSmdNdkXxBOPkMZYGd5areJdknQHj5fJIJ
w5YUDuoAOyGJJuOC7Z9PaJl3YR/Z4TFC5XUZ4zvGeDYxsjyLoxEhfGxME4YMzsFnibI7BPd8KiiW
w8czBdPrrce9xJT36cHtwKqRZFoxGERSdHR+fFeabQ2QZ6lBmuy8jMPdxWd/j9pA01NqdAe64ZgT
0L2q832r65/8Om8+Bgi7cwLBdX8tjBER0yEtmD0ZoTIUiDyg5kJ7jRc1PWx7rOeMHIWlkg7MBNOb
zwZ5R8DyTF5HODn65vqYQ5taMItP6kpKAs9IS0uRX9qEIqPUFwA55Jz/GPdr4WE1KEtcfDq6wrZw
A6oq/XiPimWGi1Qjz6uKpzjbKqANbbrepwWMU5M/k0BZGdFyJ8YHyvnsgbaQ7wpPgO8B+8LxWFFx
m9ePeIn+9iiO9Hfwazc3kzTZEzrVXBDeK4e7rNn5Icp/AjSD7PRG3XMp77IQyp5xCcuta99NIHCy
tT5jdeGcHgim4d2W+tlWE697lRCFmyHg8gyLSNjD3Bk5b1zyDmvfAHiI+yPlWipB7Qj5qq3h44uj
bFgObNZERGQo5FofTnFqFpS0IJpu75+rNBGfHcdhn4xvld0VSa9bORL/U2I0fszmKDFL/GwVX/Fb
UV88BEYAvQX0usRytkb1fVDSzM7OzKPJoF+0xPdGAekyIw7OLuzbFJzz5THxt7PKcNT7pmHd2l09
nKT+7+GruTkvoY6tkR3Ds70rZLN1Bz2D04JkEWvOEdARjIekIhIXYQyDyzgIh5wChEGH6ZM3c8uI
Yd6iAZqLAj5RDWq1m4A9E0JXBaIkfMivesYO0PSvSR8Aek9hfs4tocQ18VCIihTHzua9jFNTVESW
ltZGiBV0naz1dcQzaAkf5meIFUY8N3nEibf+gNs4H8l0yUKzwd99n3UAySC1bbxkc6c01yWYoxZ0
nrYQnStM7QMwChoRxTlyblWp03dNckUB12WvQoYXuh+L+zsUJJHApx20CA5Xt9GDJRdTgh/g/0T4
O+QeVCUazo2t1Y7ksxsiLHuO7I9YoE5PXDqY/ZvvHj5oRzu36rQ+SChD62Emc9H1Hgia32V6ENhx
E3oW0qOrDxnP8yZ3oXTEfsHu/ofJbf/ldsQz31KiDfNwwKxPG2MpMbBpxAXg788igcaW0SDXSN2R
Z7EvAjdX6hg7oP1orknZbzt8Ov4cdusqsl/aG9A4drki/wDCB3lIuLXW+GaT36aa8Z3SHpL7dNJW
qUhb0nuIgQBGaTCrRbvJDODT+OFIUwxcL0V1gojdH2yekYk88a6kWnSJ1kAuDBQ/JK0C0clYXvW2
BcBmCl6uPU9r4M4Mf11cALPXGrDek7YTq2gfepw4kHeAPVlpNcSYp1di7Q4M8+/7+kDx0+qVcvWy
ZMDlgvEDA8gVSI90T0GEnE0BYlo8R3ASMC6lgkCPef7yD5ewc5a9pwySv1SJcWKukeiIDJUGZ0DH
6Pmlzxxafo55tkn9ffJdUXeP+yf7QqX33dzmr6O6+BYlgG+zFSeFFz9OiDati4TemSvyljAmbdAU
R1Z/DfAtBNeqwPc4MkiRKU6JlseaYRKow3gFGzcP+xn8HjKO9bJfwsKaGInzxKt/Pwdi2sBVGDUB
h8k8M6VzAzj6qcrga1KKZz+i4bIxJLj8zZP/gX4C+w7ZucN44jYe6vtaP1rivE9o3v5A6rJHQy7U
+Lec/ihqpSS+MB0YgCCCafo8x1ZGxYPgeM8lFD7PQ2SSGw4wShZ1IACnKWR9RhzbSzOukoc2SW+V
l9mO0Ycj8zLhIqBpHtrR9DcbJakU/RLmXb2HL2VH6EfLjqKIGSuEE4eWYHXW4/dqswkTV5Wg4FJd
cO0HLPIfmanK45QYG+TjcsgVUx8iMO+n3zc/ZsyayUiqaQs9+OAeq7iBZQUU87z8mXyhQN3CotrD
ATUyiMkvRY1OPsn+/p81DSb8XtOO13K1fSDY+v3SDb0eZh0x6uSOwfUrccoqoQhq7ny7IFUFenb9
UvJh4ABjL6Vt6+YJa5eV5vcglxCJX22EUVHQrITCm2CN2qQgzEYiHsqjorg0LpE2Nrw0KZz2zxwU
CQomcLmvklkkGwa4FxMLLFUz6reqmGJwu1xjnENZSg+NBKICEzbPQU90Fh8hXylejWChyzdd+IRr
wlQ2XM3FLI1bQB0PF28CjwjA1Ba/fpYJEs41UpQtORLXUstUJcwOqMib88eERhPMAw281A/crGQE
g10C+WD9knZCk9SYcN0DxDedsDTTt+T2SDEr1tw59jN3YmK0SZMH/iuEDfKrCUvoaspYpzdrugS+
/IVvN2dz4f9w4X67/TFI1IAgXzjXJqkXwr1cT/WORKy87so05PLWtz20CNdx9y1i5NgJxrpbArrS
Vp5Jo7cw8CAfFEljKY2vNEZ6RVRn7HgwrmAo1sPO33owwP+XHEGd9T5QqxlviKmohuOQLn+BuQzY
t+yclZCgmr2OvPrYaJebs4qJEhc67Pf6owHemQi9NAeEIJzBD0vJrbt1hFQ2UEyR+huC93qAmsbG
O3PkHvBUqKD2vgFoBKklIaofwg3qIBMFdRDyFhUHZxJDdhXa1mPGrfoDl4DC7F+OB+4mkf7+al2p
1q1ucoeq69FL04rp7daM5khuJn8XIcIZQoLtY0CNho/9/QERc+LL9RMhdoewNEzsoovo5HSF3QtF
ZG1+l7N6MEphguoe+9WWZs+5brzZoZ3fI6lH+AcWphomGhzejalczeb/kD9BsgmWoKYNw9OCZpis
2TxwlMTeaFp4wLeMG4CKWzLXlADHx7WaSQMr7ruZTC6uoNxGphrPFGbpJPYNt7HCoPOE98IgHMqG
2QDpdoyl8Ie2JsaMD7njy0zOzhz88d76V3jOY0ljOu46dDBg9dyo951zhxIVJ/TaMQXEmVwtz642
0DpcAx+9ikHwcWf1SnZSLibsXqZkHuMmOwrGgryYRwF0hgoKR2doA1Fcqt7l2/rR2f4WFB32/w+z
wlCvJSpmJPKnk8F0NCMr3HdG0T7KS4SppEgRAtSL9sE1JIi5g/8H/OF4Cg6un1Tri4dXE3z2eykQ
a/rUHW6pzTQr5wqqkmbEx5Jp4Qv5kYvwr0JlvSsV1kyV6qJMA1YBUh5wofw4AOZFsOv8jE5hycq7
/Sq5oejr9CBz4jpAT/uK9XhnDbNeMoIb4E7saOMtYHl88XBtLpgOPz+jAgqb1Irok+mBVNf2cxn2
dMDEaJaKUAMCyjWYYjlA9sPmdz2QMig0nfWuMrKes/S0CK5c6TDdCbc+bHYX9cvvBnh8I7A11rSC
pyJMnNKQd4SF+3ky7pY0+WWIngdEfoSzZGuvaLvECFxYYdKlkTzHITnxcJP1toO8FYjiobmE7LmS
b+oxnq27Ql7aDCq3Axl9TFXnQzivoIwrNiWmGoQIcmpb4/OjPzCIJB07WDXFwKacqtoLZaxQdVl/
waWgmpCXi/hpWajA8JkrUMqUhu+fTgg0WUKcGnwURd9xS6G+iTAZlOFeKcp5I3AoG4TpDQBkRegh
JhS4wx+uHXfa/xPvQRcQAm2W7wkcC0tuBt32TPXnPK+i8A9TeEkHfH1IaON7VzqtnOtjhGdRvU/0
JrSw1HBR/A/7asDLWjfComvIzBb9YZaWCcJwGkoN08T5Nk6SgAOBrL2XwjKrqDrKG8lOUiJDKGSp
VY7GAwQM0XBE5zYtn07go4eOxiUaLBi7wagpwpie1PI2PMbtMaWSdwD8AHaQ6SAGAzGGkZzRW8Gw
lCLUsXLBjE6VYyw9mlfhEWsbKSRxdcwVKTUGJyDLXq3Ldmyszn1yBglqHN83/IgKqUQZxoODjDBX
Yy4W5LoIKOs+oTIAcjz1JMgj/ZlDMqnIpcwR1ePXSAH5SAXaFNzFyadb2LLDYlJE3dGuO87SUgv3
h5Huej9Di6jbj1Na58I2pBrLe6l8RmQnkqxm7xfnFIS9z8a0KBxp7oPcyjtaytEzRHJqoPE8FRa/
b/wxm0WVBnpwCnMSGwk8c0sf5GzNgVXUwP/JKbAounZGyG97S32LO0ZPf9PyQ02XsMS9sYJ2O6iP
RIWFGo2c/Vk5/fJzS/8izPSAoiiY3ObXw1fGyvsj/N8Yr/8ujlUFC/eXTcp3fcbe+V79XzfKjhui
PLkJO6sqPITNOaf4svPjiePC6XuymDsVAmXEZlPX93p36nuwHIPGKvO/achbNxHhbYrL5jEPpoAR
SMJn3gowGCY4GtFnX9euXcIuP9Xh1p7KzbcOnmL9wNJh3ipJGaYMb8HJugqeLfd/dXfuaB/bWxw8
rn02gSFnIvtL7UppCXfDVK8bMWNStkU1b2Sf2j2qX4RK5FB445gKOClXaRzvkF1DeJ/quTKHlaaZ
o1PiUDnjb7ZEGPv/SeuiYKdZNxqxcn3NEf1tquxVQAcnOazIxOhGkKTRG65Rr/juYBlxyU5pj0V/
rLOB0ugE6PzsH3FxBnlAEAbdyB9AUdeHKKmqHqDR2+OoxNAMnO9AZvgrH6WWCZCodwYXy35SrD+c
BjOI0oibUsCcsUYNW4sqOcMXdXzlcB7NxzO1A+3wfyunGOUaoSMqBI6WHt7JhYVm1we5cEkGAMmA
3kcTch3A4E/pwQ6JwkU3ZCbQ8uyZWoBotZRlMR3FLsDBbwj+YvsclWbNBTZBY5PHz6Ljp2h9vdqN
lCYIszlMkeElFsMrcBuUg8srhS38vw+ftp5VQXyNFKw8gxJtxWn8OBPsGZ/yzHWcnkgVOQGG5mQm
WemXBsRljnGDq8VgXsIjfRsYvNq5hjVXvBRZ56XjaQcfTZ4EevZTx9X3UnGK1gREM6CNpAlykI0O
gMd3pXi0D+cT08aAbMiwdBVXC5nqcn2ErZNjGwp/ZtLKgemD9E3NlCW3ctcgDywI5ZzXb+Fx7lBp
kOrZIPXfXbCkHAinJWFtkt6JWWf4J59vwpuWYdsVtCsH0we8mxfD3nR+OqNOSf+UwxfkrB+KFc0/
1zqjirVi5wHVwuUdH1eNk7RsEOw0J4TVSZ7C/HBbMBA+1MSrTYNgqkJLI2CDyXNDhoIs4bQN6KPD
u+IdkJ39+hfccJQA1u/KsR2fAwpMOh3YuwdT/1iHMMCOWSxnEwksygp9O92tCG5ZIuLVCWlhTtpH
bJ/sWLbgTBUtMseTqZLv+CtYNjnDfWAe7VczTTTqBkgHUt26o9xHQUZu+vAU0Z8XJBlh32Ai+BqO
BNRAAV/gW6aHQB9yyyvkZYuhumvYmq0gw1SI3qZxihXbMLadpvJ9ugzXEtQgwuJQyy+BLSBAMNvt
f/ZEiIpG6tgtyaiB6wD2snObUKNypcRV0r1xpXuXXh/qxJ65yNXZIjdPdtfFaLfD2fk1Uexwbt2N
kHlx40GZ6Yt8b46EW6K2Stac76uAh54dvfG8f/+jCN2aWrOqPvDZHjjEW556y/LQUOlvqXJkywr8
UM8uZK/5KdGSFqdOLn+0Of6+ViqBZk++2acCjMXnB64OrvfKlNgQZ8CH/Gw8vZrmyYovoJsUNHTi
MQCDZitm7qx+QfUuQBLHkHCjlGWF8Lb+RwKkCLKCG8JQxpgdorJuNytiJ9NGahH1iooK3MrpRpBq
BzSdg59sFk3e9QKeTWYDasWxT9TKOsAFeFTkwGc7P8s/0SE4heW9NEhHZ5FkynngKj42ipGsUC21
iOkGVvM08ZLUEiV/kKPEH1qrQACyMSlX7McMuWUsgMkp7I8kUF8hr5X5x47FNiRM1i+HQrqwq55W
/3GKhi2afzFErFcZdxbUYk1XtTRyqX1zRESQ9zpUH6y9BrDma6e+vKDLsmf4lwc4nFRBrEkf1JsC
3j43TMFr8VxpFiJQwVn3NbI5vJN8mKqILCa0F8rfH/bgkd2Ln+MEtXXxhWPLVsw4WazSLEvBwB1L
kJ0fLKNtWUIEGWbgCtx/Q1teCBhFkayYzC0JnR96EDBW6yl3RG74GjH1kMyU5XDAb4PXIePRVFUl
HHSoH1+T5g5045ddy+h0ATm840/NupfPPhW/IR8v+CTP6mxEXIrzBpEMVOlSkaFiBZdZm5MxDeiG
3SVBr1/zvXSinHc90WK/SyPYiD8xxOSv879AP7iwfe5VTLpoMb3VPoJuCWWOyMjyfSMdBKo7nrNV
od766TajTlU+3SmD7xnTOuIxRmxUGkf+esVz0AHP7XUyfarQs1Cuy58dZV8BbmvuEqb3lFlHy/1/
SPJ2LrqoxGD78V4bGq8D7nNxAKd4kxj+9YVv4WQkgL7r/Ov82EqOaHYC1rp//pPqBU7NuXifbhBE
UTsKGTMEJV2QCBmJJPVhWK3SyiIhmSEpv9Kbv66Tz7QpgwiAWggr5ANcTJ5HRiAWw0vm51Xwzyav
UfKV/GYUAgJ1qQSWYWFr0TzPYVRo/UuDMSWwW74PHXGVuMmH74SCIuE/VmN6zbbhjmj5vtRelQ7V
12GdS35ii8o1QZkHkozqJrwlbmG9FpKAtDajC0e4efMv148Xuj8Jwy+3tyGUMUMu9jMNW8rta1Rz
OyynJAghLNjonlb8YqGv8SjjEJ21lXUYq4O3YqNbRAW1Si3kjAqqX3WBFlDOdN7te0wHhkysWc2j
VJ6XN6si7eOSfDqR/7+pMFt33BoDKcusKUhv3hLz1pVPXcJ1ogO1Yn6hU9sF2KHMGJoY+eCuFBx8
M7DpCL4Siq61UUYAa/fpGxB8Ub5UyrLa4vn74HFsXFEhSu+8Yvag/1nC5j2+9QW8+R8/QJHZU73Z
OqDRaNaM1kvRd7UiL9PrLUYhBn1t3vC5g4R5rc/GnySRplbq/+y6vgUC42qtlWmUQZJikdnXqCN1
rCQrUHAGiY64Sa9YLtJx0tTSwUEbWf5jRQ/uBir0t/nLgZfquwgvjxYiyIz6c3qGh9brl+38+aeK
SDLxrbe0UktZRO6Ag4sSBXCmvUHQ8N3iW5zKrdO62vS0KRhBCuxc2UIAl1aeuGcVT+iwkc2t4fKt
+PK44UWdR0s3UzmDaOhVY0J6XSifSd8ZPgbpoUmrUuYGTKPMrFmO2dVE0pApcrAEvoMl8av5Tj3m
5rCSHX5XOGdSupeLQNKodCP/A5wVmfmHAPU0gwgCID6Lca3LYDI+UT2ZMvHwxqt4qihDs6l85xc+
Ds2dndy15baaMij5BErEuoEVjSCtAtwZobmU/XXImfdikLn6hh98LHT2/Pf91qiqRGIesozW8dek
qn7a9sLWT4ZOrm7f0Q0+VWwgoCcrtFzflyI4bjoNEKW3zl2Zu1YBdzOEzpvGB6c8+Xq6/UnBWHLk
MaeKAsk447EOT4q74cknX4l7Smb9LIGsAgz7mfrlRCT2Z+y9fpSKAIzCpNfGGqaS5kW2L4GHhGuj
+tSiT3x+J/InP0SJDScUdRfcNsDO93v5SZHYDI8gij78KtC54cbL0g0gYNEVMkfnpNoc6lZTWJvr
qF2LJubIiJDR6gN2kCuXErScSzLjdnj83MHUEHc/ukSlNvm10mP3pWNfur+iDV0TR0dA6zWHTnFc
GUMDIHdhgSeEvv64ApHAQozIcOam1gtSVcDT3KKRTcZXvzUz5DiG02iBZgsCjYT49QsxO2/OCJUg
o9f57v4NYfJsVVIVDkK8Xcnbm40OJkC9Bn5NbkXEKjc8VfUooIXsvoM4TDVlariWV9G/fje4vJEB
Pj7vRy5BoRWh3r09KomZ1hOf9w2OSIVkUdF0UrqAsT9TePDAKB8pLQBKHL+bmGze0KzkXWbzryr/
nQIrh9lEf0JZGQ3o4j7MjloyG0Y9bmT5/zLjslndCHLmMwHRXvFGOHVDBLcrdlcccEB+RDkZ+GEv
C3DvjX9nsi8wtTGRTJJOaOac9/+cY6H47mglk+/dPFXQaWXqYrJUgPpV5FRFbeVXABgeU+AGSzE3
cAJd4Z4pIbHC9v60NzfVwV4iT3Tktp3HrJSVQCTQVHMFoPa3/llFwDj/j/upJ43wX6mN7aUJQkm4
VRJYLsPkFImolta7YPtNWsbANDfcqFzUqG+NEBixR3XebnxPzJiQCKrd5xCvwgPLOggfzTpvnvWg
i25mKRyBpQz8csR15CAzq6Kr7HU98ownU6p60ggzcJWq0AXWOUGYNec7zl+AJssS7FXav8l95oDD
I66dWcKTPJ59PKXGo42ER250GxLu6o82zpLiRQ8I58mzo7uL4+eTHFPZdBGjADzGbP3VgZcnpQCM
KAgzMLSvN/nxXPp5C07VS5enE++DWNBsQiLlfk6DXXBdv6Frq4t5nTWdVEfmEh+lB1CiHw825xwb
2xHBxUk606UOfZL++S2SKvOguFiFCip2iN3ErvaMX6icgFcu0fc4zDRjOQsjiy3XGKk+wxALsZcm
0TQKPTOE4FJOQf4kFAmMlVx7tHSCZWydzBccBl1+bPRTaIm1N94qy2g0KcdX0K0ksn0JM+LCQX4t
z+QiBI/XGC5nkBaP9zKQt5KXE9G8uxmPEdUoLnc2RbuMzyJWjrEyYVTb9z48R5BC/as+3+L/Kefh
xpEqP3Bj6npWSLrPZ4fB0bSvGPi+puxY1cAj4B1b5zvzwBw/Y0tiX4fDDUsWQ9ECidf9lmD0/73c
cTwMkgRoY0j58uTUYuxykF/bhbQ8HFx7TeXumUf+890ySt/l3XgvS2OEs1+g1OJ7XwSp7kBguo4h
awkySR1tYyz+sqfeFezjTMXDjMoHU+tLE3fx4KS7pLZBWhsPC46iTFsd8a2tiiVNk7+P484xu3t8
cAZUookjhMk1ztdShi6FzJEY2B6w30nKIIk2GC9RiLUkpbPLqxeZvX3/13VjwSl4/MIdT3IVtvMb
C/LTc1oEvCUkNwdCeVIRom8RkU5BcphHGuvA8W1Qv1tJlBuIxf+guphqblpCCdi51h5aTD6QjM7j
Kh1ELQsWBk72dbLtnEh8XqNQsF4IGZnaR/OzLHOfnrizZ2iB8b29mA/AuR7dS1Bhdn06IFq5MEaS
g9khQOezPANDH4cbnCRz95Q3j4iuGnT3/nE0wzJw4Q3hIPrMgTTooXiskCwbd3pF2XZCuD93JD2/
BSy5tWDU8OSSh43dSa2AE+Sxba9340E8LoWEeCkgHO7j3oneTguHC0QlyL9vGaAi33OfdSZZ5y6D
P/2eVF7Fw/VWUraXfYXWEYys323ESvDk9Fi2GQ0PNyIx9/myj8v2UXPWSF/F56lIRwvC+gHLEx2N
gkLAoCBTGMm1DSXJb7bMZhi4XlTpIvN2LSKSu/aYfcCH/FTk+RyP2baOMm1/wa5GpwPD0SpCOBS7
gTiuIW4y4TwteDqQ6GoVtkbx1zC/Eua1dpk8yLEBYRI/iP99SYyN8A1K9/B32GCsoCoMf3QF8mfQ
vsETx5x2nrBmbeK5peec5yi4sstXF5O3ahqgdlW4O/vWtuUVTxgDasjFMciPhv8aRMEAvs5U+8NC
AYc5RyDs3UBAm1kxuPszTLpsK6EMPBlw+mYAqL8h8s3Uakry/7J0ombNGoeFDzuFZjuFzJZPeuTg
8BhSfOcxWnbm53BYRZDBFcY/1iZRm1Vxkld8vmoCdI2jdsRrMMSGXC8onExeWrpFvhlRFGR6KdBL
fdP/7KwOCi5ELeDNPT6B5k4Gs4JHfMJnWe8YFWVG9FtC9p1cWrqLDYZCK+dTZUslyj++NYqTHUGM
N6skRp/iEIU38RJGlxk++ss9lfttLtAooHQuocSh3ha9Lq+TM1cQA/cjFAXdNZfWTRT1Mk+4visq
ue/OEsJYPfQNgDrs+Yc3ULFDijmadyIPLqR8fqKq1GjGgTqGxf0beJd1DIykACqAo+A8avN8JV1d
4vgj5O4qfaqYJCGtoxPnqVd9LKpIBmFb6st4cPGd1CxKvNfol5Mut9q1JJI/+UEcPC3qZUUIy+Ph
TLalb1Y2fsIWWdeQAUJ97HkXyVcr23ls31Ksc8Ly1mL8ZgL4trfbXS2f3U2U7uMnzTHBU/EOdOgf
VJ7TkUrJQhD6AI7nggAjfFiIVa0b41J7Nv/rCj0XR06XMUifRX0eqowa+spVafjP7vItNUak2Q2V
9BRpSqSPlH4biB2/+8BK5ls4OBwJbmzZtlCyiVl1YtB7Fqs1sG8lFoiNEm+OIQEIQrCICHv3xF9L
3xLRJUoepwxgpDtWwLbA1V+EaWogn201YJbtylSd9hqQDqPktLnWWMbpng4PpX08qhBMLRJxwa8i
sWTVaYWbJWL+jDwwDb9FmYTf9sGCEgD21EQJbmay3pVKgXb7LLEKCyawy5IuhZQRMzsUn3KysNcE
RejX0xRVSzw3dF1m4BHCG2AcV0EEMYZgwXLORSyWeElPVAmLB3C7wevRQy89RuNyCnBlqb39E0pC
wmE25LsLXNtjFa4OlUpEaXCdTusvYN38M2SqHquVskAIrZBPaQUhz6Z9bcN/8ezsyXLnT4L2+wVb
rbQHd12kqI5J/NyrxVEr9d5b9ILWj4JlkoYwg3OaW7W832HFnRG9OTnPpPtLVGZRygGEITqIx0Da
S/y6whBIdqSznlEx3/3AyW4rQW886nrAYPE8BVB8BffO4Ry/CFgWJmISL/jHePf7lvXa5KN+LK3b
fjA0p93ZlS6Y2yo/d5TLXc3VKapu4jE1bgj3iLo58qR1oWxAIaJoJhY3J/biBRDPa84q2xnMNV6L
UxClxDu+6TDI6/x+ZDYtVQlLhE3KSjA+zKydniqDTEyqvAhi06xWITIOCeKaJr1CcfJ5RkKm9jGT
guYS0mjlN5AMk03TDDyNEQCWcqUTXmXM3Jux0CNKW2JyeqtUex6MzvOlo5tL14xA4afszTVE+QEw
owRZ31g6WvJYeKJyplrkpYtONmQn90gFE+8x2LlwFc3ct5w2g6Lc7PapOLNNDlXQ6jTne2EW0TQO
P8TGSV8PBe/Kd2wqYCRnBI+efJ1EISG+fL25R2hahumPALe+J4Lwm0mROMA0dHdyswD9m6pp3g6W
unvNpD9DGkKZt05NQ617E03lEhfzHJDicdT0KUcWnBho0jgiQM2n0Vdf7j5M9WYyjgUidJsttu6x
6cPatLhGMUHmXdKx1Lt0EChRHs1YxCCmNkh6Ao4UvkEwGKdy3qJovvx283zDmoxcmIURyOJNo36Y
VEwsygPdaiTvPyGM5WyIH0sIZslToCPLfoizSRAr1lMVyDS6a07wfIPW1VAskm5i2YbKUuNGYnr1
8tcSFsl1lpfeR3jZI5jbybST9uPK2Rmvl0Waik8Ln3CjQD0zAu9L9iq9tLKhIL/vGAuEiS+qEO5v
fkWPe8rGeFWxzstWorP1gwVKSzIZMr5ppCk7DQVuDfzrP090SllzI0+DaRRYikuY+K+CNfA9H4A8
4hdQOgp+mnvPui55Xdc3Q95nT9dAw9SVf3HSNf5z4AwKZd1guD5fQZIGMs4iFkFjxBoWWOIp1ubW
CjPnW90LhE7gNMmjMYU1qcLO973dgaND3OlLYkT9dzZ3aqdLRHi/2Qem2iuXuk528YORnV+i8lM8
j5Gv3il2K/W8LX1rKX0Kr7DAdxSg3lfujsJNab3Ta0rXvPOMi19/Fz+7pEW5Brh1b3YkB3JUGNKB
d3lNYeYV8kvpMeYuwa7mv5l9d0LhhW6pUZG9eA8OgZZxazouM/v+Ce0/u39JfKWE+AKVI56OL7wW
FnLRGJX59MMoUbYGownI33F8RPO9jwuBH0b7VuvEvHcRo58SLTJTQsUNceytqUCbMBXg/ZOx5eIq
o6DtZpAmlnwxfq8n/JolslgA2bcuufn+JdaWy7hKfOkVZzzpH66v6wCvDW+84HzxqJY1W06omDKz
dqo8i/i+es+XgoABV2a9UvhWy3I6juPNVDoT2bnhd/iCgIekkR1ikULUULrcj4MB7jrSv18g590+
h1qzLH8N3VsBDeVAp6/zgASNall2FbJauHB+w4mBb7hKVstpqlSEd2Kh4l/n7YhvfuWp2jPguldb
I2Tb0nOCxkRxn4gZ6/OpodhQkKh8mqH2N6kBRfn+n0rBPyyy0eKdMnbvDT5lp2Il0YHvfHiTN0SO
PhvijzeXZWsNGThbFFlgBFrluQJZ1cqmI721X8X6/NlooNh2iGm21coSn1eCU6+BSYSeGNI6vhOv
AQmlwZQ/xkbDPsWJ6lX3UjnFzUCE6flSn1oKjTxGk4VVOAiQIJpaMo419+vphv32U0KU/0FqeTSf
DfTcEq+jwDA/Y1apZcJO3B+qwQcK8bSNJ1NRMPDp2DNZ0KynusUxiEPGnz6v9Fp5S8sxtZmoBk56
yeYUEDONblSKoei4pxkFESw2Zupr5Zo4qeseNvmeLGMOrKvA7suae6Que/VnrtedmBHC4aQq30hg
9506eXG7U42QSoI3/YXlUeZrHGMCsV1X4N+uqQf5KCICHG2PIwzk1aHYBqyWCQuk2QO93M10Q+qj
3CyKgm1JcF2U4FkNwineYrm2mqxWOe8varsKVLDUPVuGYD9Va+i1wdWndZe+WSpnExV8pOsKtFTd
sc8luHJuUtePk1SrEt+sntbrc3qbURb4VU8E7l/qia99cqxnnjNgQPMz4zhsHa34ktQ6lpBYG7jx
dBIA2XU8Jotvi0v6aMybtDz0sgLHwsFuUtRpUFbZHgfuWAqvdTaNme56DFVQFuG2YibMTM7EI5KE
BCQMU+pstVN0DB/W6V2RhmMZUMq34fe39kpDAIz2J1GM+IvaBPsJ+ommCpVxk6RCMIiwxlVf6t71
MIt2x/qTwQMGMizDV3BqBn7sJ+HVqKEaJEoeuBB/csIlIPZsglOChrlHHmir0FP34aWHlUo54BW/
u7/FgzvaL1Z3aWENqKe1dHQOVeHwgAA9MbpVRT/EXaectrTDerArmU3lGcFXfd0puo4pIQsck14n
EaZjfOWcICCtONfsK2yUqOVk6PcWHRXRPZUHg7ma62tUcpJl3pJ9r31X8SM/81zvr63q1oVfyOI/
W2x/THN8ruZqQkuxcwj1o8+ZFHSbVvNuPdcsxEzGKeGrrEgV7hoxDSlCYIzHuxzo6v/ft/vvZNw2
b69W7Yo4RHkUPMzVC7hwoyKmbH1JMtSM2rB7n30cQFYCkJfzQcDJbAqNXMOUE3KK74jYwVPybcMV
43/5Zancjbh0JqRGMz2SFjanSXmt7RlvD1HggcvWGrMNZOJk1/SDZ9tvpINmhfrvAh6Bt9we4k64
aYU+x7TXmb1Rdjj2hA1SWoX1JusLLD9awfGLlZbzk/wR0Xv9AjK8OTbCxyr0U1l5hLKZo+VSeyt6
WUxy2DtIt18FGaxnmPCkY+i6K5oSL/qaCuiKdgKacEUa1fx2Xq92blkrHnqDBfG3CTp9NuzHTOT1
CTDnxCOjh02cfSj+jggf9aQONGYARWhd1s04djVPlB+uDqTqGZwsd/mWwOi1F694qkc3NQe1nGn9
axZroHDwFc1pyfZIx6ONZ3H49GVXs7NUCcVGOzh84qHzhWYeZcaSk462Ne7bt1MgkULGF4GOfrNu
geWYZmFZsMGhBMrwBT/1BwUrke14+Vh5MyxhO4E02ge76WjJipvUvTJ92Dd4toaSpv9TB/y2aeuV
yblqYW8Hlv6yd3IAEnvBxg6RFpwTO3owYb5mpwiJJ9/I9X5A37PMQp9UzFDjrA4ZNVlJU4hwtXUK
a3ki5O8S9sjzYbX0YkoOiFGACIaPgKWEN736Srns8rfRG4SpxOWJlfN3urvM9CvyT4xnMj4NY0IU
D+0ZtPJjLSm+D5bKkjNZnS/4Gn4549fjVSHTofyNIZbMxA+NmZXEJFhbyR9R2GT0KdzpGKqRBh+d
QEBkB6oQpql8E3zMwNMJd7dXG2lmuiL8ZSDQoTUyd7wBxWxMBcCuisNKJr8XRCTHRwY8OCewgOfc
WR6UjYzaAc5Uqq0moJ3iOBdYwLu0R+uH8c8b66n+D36jc2PXePbkiNmxyYOnbdW1RoYLPiBelfmD
gtazBPv7/h8y/Lm8tHf1YncQQ+V2ctH9DsDsvfYqZhq4p5L5+A9iWAPK2kU2z2oXKIZr2+F6eSNU
aMZob5EL6x7ScQWBwPrNZnWJugdsKrIzMfF73aNvQfTB38tHJ4AlpA7OUypAeSgf4Q9oX1kFs0LN
8LaYfjpOijys4Qo83yjnOi1v3Jim3U939TlSuXkYUIvRV7GRQojPlX0Z0OEVYh/h9waeZdq+wOkx
ERq2N/SpHyGqQwfvzzZUf4xUKDnA6Y1a2ueZqd4RfcJnn8tMXJb1xqYyFHwwXdhJ3p/6F/rTqVVI
OpoWn12tq/1dFBXccEzJx3T8snV09104aSlOmoRUw64/Q1nOojQLfIB6oBRCzInhbXO5KZmyctya
pj+K/WqpssZT6w//xYJ7/yrrkZpmRU5uvfujE2/pxJGFfU6v9mhsTbxxYBM/2zE4tSoAmwMs+cW7
MT9EqC4Cp8VOxIdP/edgJJqOzv+p4VFPu4sra+h9XlNa5Qif9x2CoX1sULljmJUhGt6EQBIOOu0i
kgqmlXQcMZnXCfFzyatsFuG5uuH+ZvGlEwUx9buUyXuVFEkuT5TO+gdDVlVWA8wVR+KXvGCXMgQq
1XGxge1dL2lK3YnykZYLdJGTZ/3paxSgz5rRHNmPiamB9QnwRHzO6o32aWh7t86nPJuvlkrBYy1l
srWm1LlEhE0Y40Zw2uXt8fZnIQHYnxphx89pcVI0xfQ/Tj/7uUw33mx/TFER1ZqqoJCYMKZMxz9D
pIzY9/nWjmRKYmONQJ3UfVQKs/lSAZcVJMuwHUVRfbbR0zxRAWceMNSjq8b+8cee1yECH+o/GnyZ
EaVNhHubktO5vegdmOmeS/n29Gn87vJK4qCNe7xIencpdWRP1oJT62z/kzLfkLpdVu+GxT3y2QQc
PENPcKxr3yMT/ViZIGGfeDVZELEO7EInUr4sYroHsCg1lNkL1Kg6inmwSGklTafn+h7Qa/3QpHZB
DVxcXld9RFifu/Okh443xwnjX39N011APPS+NaVRnpQPIE0965JMhhJUA+Y3z3F0SZj7/OCl9iUV
nQ0QxBN8SSNg0QORcc88w7UtKSc93EwmLFnBIVLn/be2US/iaBXl57/lgSTzJp6092g9TXIbFmEG
ePZ51qNr491RKX8I70ojzsoGACjxQShHalGWbwflghMDIrR9QLEXNKMK6kRxy9ig2Zg6FrecFeyw
UI0vhSIDmXfwNT1kolJniusWhwCNjr65lmvisJy/CC4dWkzzNbsjkKNQEjlpNPQP+KFP5d/MYT6o
xQkkvJz7Uh1JNZN8xYWWrBwnisVXKwjR5zVGh1nZCLLY/U5mIddsyaxtO+NM2btdUtyRVyL54Clf
sBPnq9cTvYKeWvb2AFlgyUyze2rny6NYo3OJLbeVX0injy0xv4EkbSZqzQNKkPTAP0CKTyzhKrzU
RDrG91kjEk5dZGMh9q7ZZ+w0nVFxDdXOY+Eb3kZbnwX6UZOweYt1eulwrBsUlMa0hJ17xzF8+fpV
dKKi9f/fmK0PXsvUffZ97CJKf7TWi1tc+jYbz7gKPPlwYTvS9BfyImQXCxhY5OfomATnP0qGU52F
hHvtUQBETGghTGYaLlLw62Zls1b2eJsWjZ73YRnYBRVDx2vBK07d2hGo8YlC70jQHiZ9JUxvnmdu
EMnodvRQ2yLIInrO2n+gTYzTnRMDDDkJ6n8Mju1SHArJwAAA4Aj9aDY1zeW7T1IhYR6V+eduUnpN
7dAbzPZhaeNpVED7Vg1EqAQFwVo5yPYinj0V2jnrtiWgJBt6flGH766Ltv0bIdnioYxGNKTlM0Cs
ahDJ5eLKEyNxL/nTPg0GQLpsRhhVvGhjjItjZMXcElxR7pNe3vMWlIsS3aw/3yiyHPqeFlYfiWAo
yw1dWw6GvRwX8HJk9eJu+NTeHIen6Qrn1zoUpVsB/poilulnXQ5pf/NpzotUOB9Dj49bd91JvTzN
dHcJGW6w6/T7Bq4ZuqdOkIG5MsgltSbxTX6xDOMBm0u+XwTSHeyDuAVC3C8Vku8rTRixyaFs6MzI
uHm70npCk4i5ZN8oK86Vrul8t4EMt63ayBsc/6QxvUcKQADpkHDZGONh3O1umouS70lcxjaL/RGi
ONcgm2YvUIgcVBFkjVATObaLLmCqGruZXOJ6Tkf9Pmm+UqTB++V7c8+Jkg5jQ1nR07c+FKU4SW3I
Y0iwVl9azK5zgNpxia4CWK5UYHjJP5v3Izrv23x4gYG+CUEeDWh9NKXYeN/bIYU+i/LbYlzyMAYN
C5SBpS7/UJz1BgxFZ2Nbapc+0+zm6x0/81SQdW/at4Jvn2p23mh0crbcYK3RA3Gq9M5b2KPVyePt
Lu7Wr5A4thGx3vQ9yT8adyYkaXQVptL9FxLo+iWz305PhITkRAO+elUoKmS1PjvJJUutjGsravxp
x0KJohJPX0Fr9Tz/6PLj3GjOFuScRmBmi2Ig5Qgci5yegP2zlTxZ0Hx5iJ8c2HZrtHgcL/cJVJLO
DA7t95HFPyUDktGDbj1ceGMkiXvNeoEgGIQU42jLnfOi8jHz512BL6XKWxVFjxsn51f3is4ewAwI
sKgVnhgATnH9zdmRUGvRoVbD1z49LPbSeiHA3yPEGfLOFVLUbO3KZOCt4zpyRRpiPb+5j1lfT5aq
dZaQwYyJtJ0IXmgIJ9A38q7wJsj2Bh4C2wlfV8ARioBeQoHBuYrlWOvoIRZQUgCKho/z7do8ntdy
RwcjyQS7IXLuQIInVKQHBUuLwuD5S9JhntxdyIyoM5msEquCDitrzNi4MSbIDzYkAhni8H2tJq9C
nDXGJo0ayRwWXyf6CIP6BzmpD+pWLpebWZRzH/IMcs9aOdMwOWTl1BKDv1R0sjKX6eyv2/8hgFxi
Q8tKU8TLTTrDQFNaP/8EP38vzUOM7Dw06XYjKTottPz9QIh3McoBqf28tZ4bjEOGqBhxoU0np3e8
sZocof+oQabsnFdiHo9d2HbGvk4eksKXrQSU/iTSLxrZfVtnUjkdqSJs126IdQeuOgVitYHQYHyn
gi0zYKMl41moHYm94RC151Sa4BDFKQu7TNZ0cWt0yYEW40ub2QtdpmtjLyceX7cE//F6V+jiZdMo
rKueGgOnpdTNMUMzj+AJS64pZ2biMYwuuhg3ZRD28jH0sg9EAv4L4fIvk9j6j6VepRcwOe6zxXCT
XQXhI1tn4MlA1B0fkfJyjS2H6QSJEMFsJNqd5XMRsuoQH5hPih4w/xja5uhU3ufJhx/DqvAMTrTO
SrklsC/L93aOgFTqGltDkHF3P+9evMmGl5aELiefGCfHcmy1kpVUbuSQyUWDAEdgEAeqXJTu1FjH
RsWr3Y9zJQHurQEDSchoUrbaIdLnhvW//+6xFC7HfogxiUM+mi6ZxO3Y29XGrZIpB7D1XZnpvCD9
BD01PGYlFufIxIYze3B200LluzYXnzRewDItEUMm7VIvKvCzxcRLGad1OhAeQSkSRJ1+PHHua4Oo
/Dcor7OmFDq6zKMVy0r2ngyOY9ZzvW4rrO+as3dNfhdjfjWgS2/oII24Mgd7pOu+VPBPF8fk7xcC
fNoH7mFff9sZABSvUYZRMfb0DqloZ1WX3LaWTk46gjdC8uZfK9t5U6wnaQujeGan5FqrEtN2gtgG
hJYbp2LOUVgynSqjufZwp2QkcwdmC+xavXmI5TIfbk8l4UESas6LhvffxYEwpFbcVqdCmNPleFYx
3Hr31vjFXPf6zdgQ5DagSf/bV+qCw300hrGoMy2wAj2/4Gi49FtKe2AMIsda0O50hprJcyBlkBDN
9AK3UPHHtVb9j69bcCQPUr7Mf7HEwh4EF7QVZuwjq9YZqyfBTFFRAdDvbNNwF7eIlufx2A1NSaSF
ni0nxYjGXJHTER5L95f/WTX2aALR24bxcSxM4ae+YQ7m9Hk4dD5++UhJPli1LNys0KY4/GpGTfWi
VP5edBJ3gDLhAPGp41wndxdHrsfNRs8DtGDFmhwAI20ZoaEXjBGE+58bV4OG2WTzWFEyQTb6UKnp
apKmXrldXHZIFD1vuG5HTf3gQr9/Cjg8XN0WAp8Mlp77YnGdh3W5NDiXySFLDpI1hNZdp01mmyrx
+UcVm/ksO08tNbiCAG1bZ1SQ0D21LmLO+MU/QNq1O73QKEZmR9BeAjOVGguhVmclQHDdy+Ig54tK
dV0Hk7uHUZu2TaaZg4l4p52FD46+swRH4oY8Y1llwctxRFPhv0cRMAKzf+31EadyJWIyjI5rcBB5
S/d3Px47Cq7jIuIYbyh8yFufQqYl6cC8YaAivjNR5PJirg7O9wjZ+OOBKyiOZDBVwQ8dImQCCuHe
sC9RCB+TIWOFx6FKpikAiFfX5140Sz/mN3pe9hswQmddfhJVwfZb6ldsuwg1hjSwdO3TNYZiXFet
jqoP6Q9ozfAKuxuF4q0z9Kq97mwFHvETp4UUwB1Hv9RYHWJqD7se/eOupffwesxiKIaThfeHpdeB
aosWXpLD3ill5uY2bGm4cm2kCKya3aMNMafmm8Tj4nCA9fSbOIlSHYA8A2Xkt6rBRj9H7h/vagDw
Sd3tqX1jXDeUXJk0DUk+PeATny7v8sta0EzuzdYfwp2bDjCQ/u5m8Wbi/zZgpeEDtpFmKd8tOKdy
aub8qjhIRvBfx0qNKdlLUXBgX8MHBEbwE6lBWeCVdJiavm6z/VUNBxpSEvAsWJTGrNF4s7xug7G3
RdNPrlBEabpgE5vbgsy1k/rUddSljoAvxbd9DfAegjUDC7KcTQKyUTXgorjDogzNyT5/BpPX082J
ZOQRfw1rPVdtKyTlXQJNmnyQufxg379fG62ypaU4zb74meAPHh2gg0h91xz0XH/DfP345JbDbGPg
4BhKHSpb/9AqShg6v0TDq9qhZEvFDbjsEtG3z2WUOlb+DG/OfyCqYo1tVNE0BP0sFv4zbolJXCjl
4bAqQ8t2tMYoqJ6zat/wB1GqFXK7eoWYDe0oshUBL/4D2y7FqJAz2DybsP+oCWnrG35KpXadEHl6
7vLIYar6Hon81Z8/UCL/PFR1hDIrs0x1lSmgM3DybKX7P13idsw7q54YQxE9v6cVcGoW2xFHVBWF
ufHXv1kyMFj7RfFp2Q9PdjWrqajcC8aTych7r0iiQQ9OwU7kqDPTyrzqoliogFVjBmDURCdTz3I3
EAG/b0+cyipmfQ7Vu2scVTCmSCNbhUJvikMiGb4Vblk7kXNCGZQKQ9wPTWWf1JKrBjMJX5pZLsCp
wvEMHQeIHQMHT8qiH2QRum3Wl6vx7D6ZH8kYsS4JHlJMF/meQ9XDoRXyt5gxNyyS5c8gd8prJZ+r
N61EQmVqqustg1qJ0i2SfDorDG84QB4AA/7gLR2KskqVvqetLpq87YVld8khQGncncCvHQJRB6t4
vpjmrRUzghHCxKTvOHIUg0A9tmffhxKbEC88U2nHGt7OaCBjr7u15ulz2yFacpb60q6YTLc627Ao
V+s7qIlyI5GZ0rgRZf+DEnfTzPyxTu9sHp3fO0kDSmm+gVAFYrdXI74kyavwGqvhB5Ti+QJ1FD/w
9tWelxEfa2CV2CpoPBTcggquv/rPlGmLlXcbN8kbUu5WPq+fXS6h0abbPyAEPr39zlX9NSq8vRGu
c0HfAVFEZnyQWmbyHk1tZliD/ZVUvAq+Fs34wrQLmtQGyc7eLIdJYXsdtaC47ePtjVUUa+3k1vei
AoQ5zMWpP3qJlAyTcxfJk64p5Vkr2qyUb5yqVMkidn+8KhBPqCK847fKEmsHdFdxi/FU5uBgV1Qp
A49QJOh0VJ7NWJzm/a5JUXkNwygBNU+HP7n/F2mcBs5EPlHSUDXtHQQGXyiYMmOD0l2HvYd0VdDh
ykJmBegPjd3smSesH3FKTPf+07mPP+nDfMsaN3Rb9wG98oHWCM/0+mdMbKbQ3BUKZJgxKfU0B6eD
jpUQ1Fn0F+kYjpFLpdnClvara5L/4R5LqQOMhvt/pJGD0vjOtx8BdTgzWJbAzjDny92oqiGvU31M
MpAAmWasBiZoa71d3I5+edDYEohgMRr0ugHrbI6MsRQZAwp0k/0voNAguYbRhW2qAsNNu6I3NEp0
8DKNGeC63oiKi6Xus4la3VIXaFtIauVB5UJQNx5zZG772A+vsijtaC4iNZ78pQHSivp6iLWkWzEg
g4v9fgPNSPOYFBTEPx2gCwQzdDhTu28SgP61IVLCgvvWkNHcdyG9uus+EkprvEhKIM9Ka/LpWz10
jCQSOlDbmMhMTGNcG5o+LONUCf3BcmxjEirTFGo9gKruaPBxXMtuhF0h8JOyr8LYi2aSgXCmDhKq
v/cD1StKVayztrPBdZakGwOrvMQOEs4twXeBxbG6XRiQYtZWc96MWU8Vr/PzoJD+niDQhZwKUnVj
Etq4RBOt1ORxekAcQ3SmzrOROS0d7vLUNb8zch49cNU7nJA7310dUOy82TPsfOqFVLUb4SMEdnFI
wuFRXJj7AWwweI58p8UGvx4G0E9DgkwovDm3s1PEWDJVeerDyfxvDY1x3DODKbsr1hXZI1HcveGf
3jG7dnpzNUjHjB09aR74JERynU8dhkQbp0kl8i61654qMer6Gm8i2BuK0RJDYEfLeSzCqHtV1yRP
fzHoM8s09B/2bYyW57w5qe4QntWEnV2vc+zNNzvvWvcHVmZNOQbm8rAeUpnxRQOIEEDdJFJCjZkx
vZxHkUUqIRy9b6b8pIamVM5TuqocTa/EoN4cDbZT/3sPR/SJvtnmTVAnfCMDGYhY/NEv/8eL033E
o2ZJ1znJ1eFehv+JCl+TdVaQ3Mcr7R6g0LiaCJiC40VHsce+T7ioo82VxoZ+ehesnPxWgPj27EIu
6FX/Nnw5PoAiiHGBEhvoIGNlufENf0e+U2WdVkAVxlEDQcbRRm4ozra8ytTJvWDovHG1kUqBx+OE
XVCduhaEwZg8GttHnlqvUd0vP6sSZe/Ae6IvJ5kDjmmgIlkDLyUd74cSKx2eeoARZkUEC4dIurVN
JW/94sKhYRquoZkCtoxiJ6DoY7lh2cxNfTAzWKJUCqujMavzf8/ZS7CDs/ZAAMnKqXpidPPQahCT
KbBbCFEnWbHzHBZTncSiOs02UiPOVVzHt2hywInWA8QpD5QP07cfsJ/rp+CotFsEu47GKRQ1q31M
oyHpAJIh4eH4rjdv8YFZuCoZwqu+8zeDZUrg27pQBf9ASFhU0NZ04nZuB7g1//Y485mGl6UmKqyx
k0rZ9IP0dm6H3ppJxo5mnXNq4QwZLv7eKaeFAXLR+3oyp35/YFDqtbTGpxWtS5PXT3B0z1ODY9sR
j2umlJ63xakIeTRHj/KBcySm1TLpeFFI21rswc/wYaRGgmCIJxlvCny+In/9GpHbBTtdtp/TxuAj
rfjQA8NLkyTGW2zUI6cV9HPjvKiCFq5tfb9RLugl5xm7k749l/DKRAQMm7H7ycqSfEtlLhUapbcR
kLtrYAPhVWkfSpSE6bRJW9oblIOtXAUqFJ7Enw9ZSJ0wonYlS+k/sNHCMl/0g4PZrqhXTnf4W5Gg
vokSIbac1+YPrjWPyjoFCarKOhypchCpyAxmK434eHPIFKqrpv25eDhloDMlHJ69MkIdkhgjST44
DrDFDs04L1M+CiUsP06Dpic5Ln/e42RDcth3T7JE5UHFXlNxliaFKyWtdQVZa2wDJikR0QrKo5Dc
bIkUqHvXIGGs+GHgOY9JN2SRZwB6tPgdkWyiNyhEt5M8qRLUVSOizDwBBXM7qGbtscx5efv0dCYH
jzlF9TVc1MYnIUy8SH0b06oorjbHlmucYown9MwpX4jlzyJGfVQsefTF5twaPVvGPOtL+EAbSGDW
hKjVPDzKJpqJ/mD31HH7XWlBIIKoPJoSs6eRef0bW5BLiMH1Tvsy0AS3Bzmax6FAU8uvyRDug+ny
Qdui8K4/95eUAj6HjvgA7Stvn8GbMXBIsE12oztW/HVqM1vlWIuphaL+1jIXLH/AqqZUbHjIAxnf
4v/3Ix/cM0Kw/fuc1/oe3ZM1C3P3AdP9B2Rr+WtShT+F/tBPxJgM8KFk6XJUA4KvzxMWv4dezWa1
rA3magmMc436NCt8l2ldGNDvU96tYMslWMrW+/BswWLUjJjAquSYzZYAPR6gY1RuBiCHK4KFVHlW
G/FTc5lTD/QicgavaoekstoYnVe0rMdEvK1gNi45THwF9NKnTs20LGDtUbFsuKuWfejUDTQGjHuP
NNV6ClqUOsdWuKW2O8iqcv/kCsscdF7q93JCRTO6I8HrD3cgwEKfi9HmVgPslJEGpRwk470KUHUW
D1If6eVeX4y/ks+xK9TV5Vs73w8BjkHQg/qnnu0yXwdH+SIZoZYJxUUiqLskX4rP41dcn7rff2Kb
WhVc9o7i5e7688c9inM9Ms5/jkbbrdsELyOqulQsJ3PIonICk0JzawuKq61nXIcDDNACUzRqFnXH
JFGI4ZAXrstGE5NndebYSHRmpiIuNu8j37/dvfrlwOPM62HIL7wnG4tDuDaxP8p9WMIaRETcQRhN
Y0eWa0XkKfkQqeYDublENEMTP1GNJAequRzPP0aNvBI0wrEOnUyXlXOb/3ehrg2II5mQFp4ivT+E
bkG+/VTFWI1mXlbG1Y7QzOOO0fKal7sovZpx/pdg5FcS9UqSVW5qOGStCP7rzgdmR3iVBhPjVrvf
QofjvJjIwF8wNScr/0PFwDbKUgAy5tzqB6t5ad1iK1pKiQmpopPe994k6V1u5AA3jSOqV1ASKxO2
7mY3mv7b5GgxZgxqTB7m6iPQJnMxS0p3VcvKA3Y8vDhbiE6Ff9ABn1KuFBG7NyErT+uyTyprbx5H
x9I6pH7zR3yRzsQcRMKh+9S0L4jjzpgV2CYIFlSdGJOJ2qJWno1qs/Ub6oD29p4eOKdEWzPVnvBu
ZUi/nRY8zPGeTPhmIerRbh2bCtN5bMTGIhnAbpFy3lkbgFCaDQPo1GVeGoprXrqNWV7HqHtFHFoV
fQTzJbGPJjLRdT3GEPODWSVSeUTUEsBq/msali2838fypzVYFxYXsa80Z0a85sxWAOiY2RX+WmXs
CvDT95GF4EEC8dWmJ8BKFkfe/nnmxgugAPUS0RtSSmKzLxioZXZhgKQgHXafFLpjIV/DT2gOyuoO
FWcDk6Q85yt4HgRLRrge7a55K7xyfbJ8gtjbl2bnHazOT4PyC8yoDD6QKs7qciBZH5ypzvz9SdSL
ideR0RAF48rVPi3InFjyCzUBvL4xO4Yz7quOWp6mOI4K4Oky8Y20gQdN98DCn0/fs0LTBjJYydSL
b87HVf8AstpBiTzrli227G/r55Kb0aGC/MA54t9ewwLzzFyh3x9W+TZbX2WD0YfjaCYmZa6MtBOD
TKOih3GZqg81NJpnWOQ5zo7o8l1IN14d+rHjVZGkf8Ox/2MSm8cvqS7XbMxVeGtRP3TD1Zv+qhSp
AcVR+R63AB27B3FgYFokBYuKsa5DKnCFzHGnTjotiZdVJxPwD8Tj30XoPXnyId+RPuZhwTVBRRyp
7mbWi0jOTwIlyYDNUQG/fcfFNmTtYm/Wi+EocbU7y7BV6LkK8sDYpAcoSEBdRfs/f0Z7aQMyOEqD
AuT6HM6qitofcslkX3hP1jHVQiKMrtciCC3DLzi5sJyYvDSERy6Euw0KfbYEArAUL7tPglW+LigW
b7mFMI/ML8JBV2FtzPFxzY6qWAC0tO/0+R/gyiyMbD26YA7dWE2yC+ZmwBxdwF/OwMlRlFxGpKEc
52p4vmmk+A5A6DxFcdyGAUyQ2t6eVRWB7j6eSbx56VHeV3RZ99huX1Hfn1A/mdz9yswN8H+YLqnu
Z+AUvxAtx7FXRr7tmvSoxuT1o/Bb4E3rHgHJbTKBqe44NyoaEbfI6YmzzROZoCQfDxwe8pAz4tGc
M1EnazEUNFOXrFbcoxuowNyA/+lW5LOVu846fMRxgIEDz9ohMfJlqXggGF70GReJPnuW4+ni2U12
GwH69qU5Dnpf19bA1ABgex9sT8LjMUXZ/k2d9cWT6AlQxp4ktmYKmmbVvpAQJOMpD90hzbOeG1b4
2tfzcrVJrDXeTutmAJdQJAgLrjUjq6/KqBtaM+DwFxc3O2c+jTTrbBVvTestK3/PqMhFIgOoRVLt
CpaKRlLEmu1PsEj37fO2QNumiBRcGg8CPpRwijiAHjYBGHicGSNtuCbrvIl2yTovckGQI5eGTt8I
Um5e2ZO94p2OpU8gO0+OqgoKexWdPHW5YuYfgFO1sjdMZ6D5mf2ha9I/dTGVDKLXfl0BF7BhXjkg
P1jOv4dh7MbUMj/x9ncB5sMQVeDqMCP0g6A+E7OaguKHeQuVxAgGeg4e9NeF+Ylt325+Py3CJREl
zDmlhJJbZXwtiGupKMWtDUeI4KIH+KUXjmN5YjlewEq57ZbZMtnJypCbR18lXoEMcOVrwUVN4myy
dBjM9PL/e1J1lKxW8KeEQhyUOwyt8d63EBkHDpcG4HWu0HHYzBlG7dW7N1GCp7De6QNWSXL7Qh/x
YeY0lRyHk9XhkR2sL+N0/dhBkJBt9BtFLyNrOnAS6VaKS2ronVYnI0nRsuO/gGCAk9b+iR8cdJ17
bo4ZbgAqJgfNIyCI9R4sDZ0q7h3i8IrjJCSDISVwD6WdpvLq0iBhfDNN/nJcDDSQwfT6bFbOBzkE
uj4PzW3E/9Iyr36uAiTzc4AcFjZyH+y2IIywA4crVr3eth9qu0bpy7rnbhFYiN9Nr9a/n2on+r+D
m2Et3/SJjj5pcgbUGlvz2XY9WOSW9R3rIL/buSsSnnO3UNAXMi3QR2knKDtFRAsKMES9ToImuhHa
9S0Ki7D4Vp14hy1hyBWLT0AP5veWnho9kRHLCAgTCrA8LLox3leGlktuu++p5ZPOeCLiJxQjH5Qs
5XlbuEKIegTcXstb2bd/z+/q/tvX7wIrabPkZTUPYPJsPJdu1yvdmRnpOzQTkcTgl7gHDFLRohC8
AYaL3g08Uy/pSdX/G660b03z3yvc4E5a7tUeDs5y1TyijZQ+RmMi3zaJI2qUBrTrrsEFWUFiRZ3P
20gqCGgB+nwkkOfXqQefDi0zd/o0BlVqAxec5x4GwgKr7EsXqKFGeSED9eiYzw96Ws1IITczg9kd
MGCdjvcmLTDRhU/YDMkUJbw9Y1WmGW+9SoziDOQrG9OtfYpR8K4JTIF06lII9H7IgSevda9D/aTV
VYe3/rwuBmqyTIi8SSgw+D3LkuyweNzFFhaCEsPq5xsX+zSXLzM2TN0i3xYxpmauoI/L2huT7nR5
PDnMvcViyyPu6+aA+MYx5WzuqpXLJjCnjszPo8Mfv8z45GDOgjxMhitH3GbxQPssUr9vQ0ePPjBu
7nCVbqSyyxR0AKMp/15ShA/GUbLajWz9/wazwd9dnSWWMX+3XgQoZacQMihO4tin9mtQ9qR/sG1y
6UjFEyczM/R+IOJhTXyUKGXtkqhZ7pZHcQWZjx2Rh4gGfkbgncvhLYr1YAC5B6VmLC52lOq47tTO
1mqwnjYeo5V0BMJiglqWN+0Eq1B0i44P5E7M3ev3FRLhpOIrth4WhYQvqGR6Q4uhIvE+S4MzF3qt
TJWwCrMCng4iEE/aa8zs0Af8+VagnQ3EieYEGx+ahY93UsGZR6ZalBbI5iXh+PZszXJ9dKCUK4a3
+erTCNBSOKEHElCQFsY9csHGxw9sm4JwRucUOQUZ/t0PZNLsdratZCs/gfLgbEF6xuErSjB4Zdn9
wfMrsEi/2N5NA+99xE6oe28gVR86ozRdXqUpbqUE8S2hog1qN1DMAG18tiVIiH2fSW3AgYcB+Oev
+pSnppqQoGXRaGpkIdvPybWemZMKhLwyvweMEoQn8b0QVAB9+AF4AcChnOgzFu7A5DhSwD8/rcYD
drHbxLTHqUPBACJQjKJfdXO8Uo5tqlwBYS/qCCBiIHBMNerauyUYoHDQ63HuMJ9fAhZX6Dqog8Y5
esNqUMO4dVCQDDtgxE4vB6EHAAI1GibP22r0ssAqLFmPRKN6WwgJaMUY9lBby5iUEZ8AAjUr+tk4
RiOhTit94oFcHBijKXyyk4P8uQSAuPKYPzf9qGDGmP37UNzeG6U2YAiTx9VCrxyg6isWHbTIW29J
kVnJRTODm/G6A7eOuM98/a3Y4eEM20qNZngK582cjf01k1y5ZV1I+XGh9x/5p/zdaEZNZmXhcOY6
q7BlMvLP7VRQFypMh0RT3OoEoS1+OY6FcTkYCUHSyyyBh5Y5PwOjZVsY+GJlfOMZSoWfV1oN7KvK
E7AqCpufU6B3MI061Ys3tVXYn8NmkjQppdbCTx4zi5OIuFzL6CtwjC0yySIg7D7SVB8dp5Ja9w0T
11AmsAeczGekWESGs1jjhGp8uN4WmQ53RBogXY1GWGziISBeYEqTwrPVBcNON5PnhjxsBTEIOS9b
JvU4dJQ3jrp+SE4CD+ncshf2YadUweIVt5tM/sNhaBVCB3H5giQIG/AaLsp9Y81oHRQLpJ7BBaL/
r6XxQmg+Ng8dfoZfmKUkNkrezSH8bbsxhrJctEAv4a7ge3tI7NqJ2K8YoFSxm100G8gpVBUdJzjM
KP3rRU+6cFFB4QaeXbRT+cdeOQAK9fkqaNT9K6fGJiExHW2s2OzVf5oAWx/5lcC6RFtToOjZCsyE
YBFry4XvFdbbvGkSJAJpojsmWNjdaNVbSD2SXPEpkPOPNgF2miz1CO8sG34BnoG4ItGik0+x3rRK
KfbG7Dzubo3+Kb8fnw1jB3htez6Mz/MmKxQTM/aCaUMQkIQpmu0x4R5zfT1NtV4OPtCvmyW9MZZ9
yqVCfIlzxKDkcUU85M9b9PxKIKZdUf2GhwuLj5iDefuGH4890mn4c0JMN/3Mjrkt+ShbdEjUZnrm
PDDaX6pioNpuovnMC6Hof2if3Svy0mSaiuRwe/mWaJEaH6jyaAclfve7vSzZypKViH3JkyBamvyL
CbTls1oWwEBaz/xS2DUY8KrktDPRhlJrLcQT/nYJNBhAmKR3nL6TJqwAfgbFC/2Esc9QXbkOX8Pz
XpkUaZ/q0IfUTjypYHhBulbwptPe4GLAb05/l4pEiFJybyYBkOx7IKmlYUFtTjijxYCXDKB20uOk
arDPai9qMKGZwRCbbBcGvdNjXfXiyhvGPaNCnjFi7GxgHQnvHak6OQC66ZH4Ynn4wD0fOv23Vqmq
+Y34hpNKrUIgEDvcKZljwZq/FXW1r3dha01pMEFnW/EmYoS7Kpw1swyh8bHmG2/0Fryx8rjoRLSE
Ec/rf+ft12rpqdYsSCq7uTCMQa9fJtFdTaEkuoXX79fTdA71IW2fJTpQ+66KLT9Ljtt6Ca5njzDr
DA+Qj5mN/7PVTVOrFX9C7ePt/fVnbEfkYNR5DLp9gMnsUwLtXb5G8GgTepuFRnRY4BWcY5IXXba1
03QCCOcoo3Yg2PSaa2u2Ew4aXQ5ozvUIdgSfcEG9VSKZVJzQz7bYuY0Va7oNTiiwGCUxS7TI1ZUm
BjOnihW32Bq85nCtxNsRTuCi6XJc+9z1ZE5Upv/no66HH+bTCCR0xt8+ljC/7dB0OoaW/rZrhTTh
e0unvYC+eFA3SBda5fssC21SRKnQe8cxIMsCzQed5gcGt7+KofW9DqQYzvucQy5bshAqoXF3bnV4
qtaQzyrmzsw9t39N6J/kX4d2DaA+DOTFB422MIeXz1+/9wnRF6VtZ2wwSYcLZG2McLVreDTbEvGn
lqJpLVq8ULGdqLfqhR4ZYT181SkuXvjzBibgANQPdrBlc12G2bvbefbdoC8E/G7M9p33JjoBDVTC
EuLG47cndgfbNMagVnr9sHxNKZxLN6SknSUslsrLwsymPXoeMq3OnJZyqB+fjCGQhW7fM+zwSfm9
SfVBHt1Yps4gXfVlJYOel8qIrmNBBw0KBQXcR+7ssWFdwEkcdZ20zMywlBoZ/KvXb+m8rF2QaeIs
ztz0cJPsLHa6qAGPuxxlw/8J4HNRcBsUZAr8HYpIxatd8YHEjiUqOAf9WxSIGtXn1U0OGdFa6XFu
G8/OcZq6a4z4I0uzd2JimkCkUJ28R8m3kYdvJM4fWyHSOGPwsbZcQU/d7kCXr6ILR4M7TL9MbNAT
rqT8TN7nQjdHPPWKE5jq9kDZ4ubV3Z3r/n1xJchLUh7KhJRwJzFB9L6LuvqfoDnUl61bRqGwScf7
NpnNFqrbNUELtlW0AqYwJ3/zLdSE73IngzEBk8slq6Y7IHYE77ZsKMOhOB5fSBbOAsScO6JWWReS
qfhpaRGa/+BTBjKdasrsy2LfHEtvTzGazYIS3T2ZeuUhhNGeDiI1CyNAhYr8q9fDGjp39cqc93Dc
U8ntSfVehhfL1TnlifovDLL2iC5mDzQ3GrEUgDa63p44/TmcJjLHM2XYY1mZeej+MOvOoXR8afD+
GNSx/jcM39Glt660bg3mkU/S9fXvBvnQ2VlIQnevigY5UrYKgzazCKT8N2KCMSR+To3g/C3bmvpp
rYAMwOL9mEd/GaoVmGnYOZsQk1zOkshfo2OVAOmX5Qstt336MoDgJB0Y6hx9qrGvLHcZhEm1OsHK
U7ybB2HHaa5pM+HrKMzwZHZW0wc5IPk3Ds7OMZdMKAo8xMk/II4erVClJuI46FXhM6058XXCzxfH
mnDvPj77UB/sA0YorQTrNrCPHgaVddnFsgbIOUJ8t2fkSynQDG/3RSOhrtZAeXtw7v1vRA1SkUEa
v5aaktBrOPfake+nuFrIPrym28z/XQeHSS0sazcnG/v1nDPiXBM7QHU7XxnJmngiASVQnewauarA
05Q7BCtsyH0IAQ0BhC/SLm8flSbgFCkM1Ex2nA9fBZRxU6Dj4xQSK+wLRaUvJxSD2m6jAVypF4RK
XLdOd1u7fJ+NQQt5zqr06o+v5ibZ0KePy+y1bh+220yxq1riEl2apt4k3zYxo3K2feM3XQiIV+E4
QX5wmswcAOPFBXqJMA1PUADbDlbDsbFT5d9HQlOxfx2tw2o0Uc3QjaIt8YAi1QrZKS4NOR7TqsUT
7MvA2YLAA9oNA2zzit6SseKmy5PAVaWawjBD5y/S3bgwBuZqkS3B3txKNdsWmryDWoAVR8QWlRVM
E+0QEbV8YAVTe1mDnD6CI9R3L9fxXMi2MCuddwixe4LObrQlyU32UI/1kLSsdD4CbmXFejdjgIlX
JXUOULwSXjlTIpzZyBiKghD0sLF+os/hiBQXvCkAlU7Ciqbe8scp26RJWRbO4sR19cjwH16C857p
uw5qQrmCnxEMZYQMiSGrPNqMPcdS4jo+GZcJKkws2FxEPhW6gtSZfLX7+swn6j6LvbTlioWTwY6w
asCh9IhJJ6MvOoAFgXnYV2q4DFM0ZxHfJlLyaRzP75Z+zSElgnO+Q0UZhqd4MUMbOjYmdO+j/T7C
nf6PKngR6gRC91LaNgVavkMD+dh97CRBOEWB9RlnFVm7aPCOp3jZfDC8twRNeEJpWNtnMte4HC8N
wCWBy+/s8t4xFDJRcJs2SUxTCn+tE7B6oT1BVJGCt5saXKHofLy7iO13awLIwHSSXvsTMl31zQHA
u43nn+Q1nN3uHe4A/PYOJTnXR1gbm6ecgw4oroS53EBJIm2XC0HXxm0IcUrZFKUJzU0TeHH34p+q
dCRgVwcBucAxhtTcpa1Sifb1TNYqTkcEKQu5OcrbqScfqdNdPDokd0AwTnKxFL4xN7s7fkbAMp93
06TDJG8Ar3GijfH4dHhD8t7TF2VneHhJW9Ml+cKUYYzwKReR4IrHwnJXntIeimDCsrf5g1I418f7
phodYYGlMhicOxMkj/CalI5NJ4I/9d02iMS7ogvc6Dx8MMX7SJiGvTAxmmjzGfw2f/m4gNKjuIWV
yO23waIFsicl7XTDo9IYkdaLhnJZCHwyxVw7rfUrnuNXPrXtAqNb326GHbUByYlGwrz9QygbI/an
aMPhQ3Cnk5EqBPvsn6HqZ4bWrVfPZ6ijAQrhzMug4pIh8LOqr5EdErQW0A+5hSnR76bARsYjV79u
/IJctLkIKhqpZW4WC9IhYODQIXoAGcgmpUNmBZ5/nk1fVXKY/zBoc1fqUEWnq+LQsoYOKH8XWY2v
jc1DRVRqjYjOq4xhnOEslRqxVwCwAwnEQrDTuCijFpGYW1XQKo0mx9WY5u9MJ/M2TwyPV/7DYfk1
IJZJT3KpB9dwr8WXm73wkkBsxwn1kQmcXjMHzwpR4NB9dURGjRAqGQc1MKg0Q5KSo2KgpD567fDm
asafLAnSYjbypoPFeeTOQsLo/tPCPKs9Y0boDU+FrYAvec6ZH2eZ2KRxAX65vkn3798hAvKu5yjC
NaFmwgZX4NjXI+Toe+GmiJp5Gx7MiFPQRMGHWlFYLZd94NMqwspvI4ZdZ6lXcjkmEBB8VOWfUssc
igIi5xaXde3XwVYoxunQ0ctnKJXlEao4E7Q1CCa+9rolD6Qjrnl5uDI8HpMbw9KYJWK210+wQNC9
NQGTiaziXd6FASgKFOardmK4BiRrro0bNAr2ZG4NFhumSZ0p7NUeRIPUk7ZgezBRP1srDTw8h7Id
CYrAe1FdIxii/vJgt5Dei3pvmHG9xjeywm1sZMT9etnS2Qj0jO+yBlDnufYspa5XrzA1ViSX7h/m
Ke3O7bqOCObOl7wnWZx0pOYvi+aqiOG6fzldx7qxz3l+cW3tqGjREq8Ph+aQAWb/OhmyhhrlpoEz
hNFyhWP3v0pAAs6mlmQagbFusadQZMU/sP8YJJ4Ds8RiU5gM7p12czjAJWAJJ92DT/WX+D5ftcpT
HTIS50xRWxIhFHVzVKHGQGwHEqtC+j7m1NWzdIFpzUk28fcewe1etlP/gyM7T6SCc94XZu1v4f6w
bgPMLPBJBdyb4mq78MURjCLxMXUef9gAllTkA2ezU79WGJeT+4LB6GmKf+4sw0ce0qfczwQJp2e0
4Gcaf5wqKiyCbUl+dQhr1StXM4jO4UW4al7LHAGGEnkUr3wODJGBE4d/8W4f78teci3a/Q+73urn
S7u+52f0tMp0oez1/aSIMZEaVIcsh/pcWa3PrrU0bOGNaWcQ/VaP1/88JeUuD72ptuGZt5CU4KA9
zi0Rt6Ho84sKKg1jps4IZYSGl5YU3QiMF6JxJIkHoN1wHFrVYf4Rfu65fW5B7LR4q9fR47i6ULSx
TN4i9GD0DnYFIsWxK7sSKGZdli9VwS8RMUTqrdasPwiJWdbxQsTc6jlwE3JKg9neq60R1qOGEuoo
3avJ0G5mPL2eS/tnvqmYDjbNu9bjRmV/GP2R9s/OUPUKjWPIXdRr8q9dDhJj6LTunOH8mHrD4W/t
rlio1lbsEgZXvsgQjxIK4NT2+SQPXNLtUSJrKj5alLUwrTLOmEGpOJ4rMDQlf2rISnAvuJLeomVp
w0BUtqHRm869ika7ix3oKxQZ0/GwkFAjS3PMfBNGIq4JzluHeOm2ChoJti7E98jAjA7Rs7TTkKso
RcstxHZ3F2VhCzMdYc/OIqzys55REhcW9TXRhxTxqH7OW2+8MwjKaLwS2XK73M5+mXZ7YgzEnFSW
vP9ieZRTlORxqk/j9gHR7uR8+c9hOUUosfsO7xvlPQ2FvU83CMPV7IFujJmPSXKm04tfyo5PkfeC
AK++KixjLjj6cCUUIkUejohqZsZ81kkMign/3R+o7M8GQ5UUO+Jpn2AJVZAEHLkOQiQcCc6tQyfr
aRbs3NlOEFm9J9iMGBzhkG1va0JtyVegkP1SWqiI92UoOVAubCsmDmFKc+BJIGZUX1P/nEIz06Kt
z4iQJIQxwpI+iauNJhs61yE2S/UOh8/N/G70BVkCw5DI773zolBEOk80lNxuqp639LdRt2g4W6jW
NxyC+uEXb3Y5TpIvHaqHDvvZhcfP+mzrqVuK2GUoBv7+Mm9VG7TkWG3nLRqoZFeiSJklZU0AN4i/
i8/p8jPKsrgIGw0Z/J4FeNWAB/0DjUY0fZ0O2sA4rs4QDSD32ZVYipmFgLp8xhmSiVypAOrqRxiW
BBPWe4lA6j0vAAiPWUnKH6NmCG11NAkef/btFCo5RDDSJjYMUHNvqR17nSeZAVGURvZQ8KtYgz6l
RRUx4R5IQAbGm/qDLusujsIGMx3BTZ7swpFLx6vPXNBxDjsv9xnCMehe00kKIzdNGtG0/Ejo+c3I
R5p/28ZGXhmXY6GUO2vYmjeaNQAL1wdEIs4m7c0044Jn2JTh+eXBjNzM8yhal+zItWCQFSu3KOjH
a/vKYZiRXdJlZW7IarRhamuBAUu/szOZ7OzpJZAX5im55kqyIgGQPOqCTWTWpGR3XKrNwqNGiJH9
3sLCDLI5JOQ/CQGu8OG+X/LaSbVRrcFK6rDMEiDFmUnMOewIumtFdugC+0Ji2HF2/7MlmMTIvJQa
b7XdnXQwpCU54GW/pNudVhi9UdlF8K3aBQ0UCivsQhj/JkSv4tXjYsc/3/GOM3Uice0NUAx2pcg2
NMWGkgUf+gGdiE4Jo5yoBZhE9Jq/ph2CqOTMPmmQ4KMxG/CiHknYA632OZVAhqqLfZ9PJld7yJQO
RKyRLAVF/Sm4uvwBxU5YAAWlMSp4KgR6C+rtHN1sDrKd8L20p3BMz3uGxrFGF4Bw+5RrU5JDdM3S
m9ECLyNHeXjR54jXAMM4eTTTrv6YuK0+3j1NkII7jzSqshgs43mvJxuxPrchIAHMrYh4aKaE8WRx
JNUvNZiarYTnXjyEwjrv+Rmtf+arDfBnNtJun8vNMZ5YLLoFpcdhejBkILKwpbnNV+KqekV7MtWP
fNnK5dsnpNdqVDCGQsbhNDUbXEW1/Yrxu1/1kIKAvn9wP+y2jsZUi072R8+tAXjW/IS0ySSl3eOP
m4KSZDNVfdWUYLHyDS9qsKV6w5UDiAlviJZNGKpyt8kkf4LctWbd7av59pNCfNnJvWt/A7/Tj86j
RV+h9ZaCZC80UXSu7gXgck8XInb7sriTr8zzOePmncNpg/3osuFRxPvmUOJ1xCgIyDqpsKXOnh6x
AyNhRLI0Y6UFi5VkKcatIFbuG8+FIT3OmZjmo6kaCNuRM58zkOUJhhI0BCZMbyJXiSo4+WyZeP+3
Jv09Km2TECOkqiibbNydSyIaDKR0Bv/IxU/0srgWb/1cbr79Vt6OuNulxExzbnRxf08BnQiCOKbp
2wzJpCVptsNMi0GxH5V96taKKl+GyfCKeZCiwJRxiCBMPlHNZNlTFuOvwZWe4/rcD2IjIYvmdvSs
GD99OQHXVm5cZgmdwDhRSI6t7uPQQyE9mIOhxUvlhLu+yD29G+wk9BaTxlBd3QM3vAKsL8/PcGZ3
8mdetgFMdYscwTbdYdPsgn3kd336FrxCkNb+pgU0GuRCAQupQpZRyu8nG8XQ/bf9BVGuJGvya25d
H4jrhpknCw2IZfGacCQnhwnjMkPm4mHp7Trzvw8zGFtktaryJYLAP/AjzTVUAxh3C+dUjtwRd8Gv
/f6PkET3buJUyQGB9gAKJGJLgtzT4T9mmYp0DhG9EpB4B37xbHVkcTwnr6uwURR46BSZAvXvGbke
vKNcmd2QOdQRCIfUPV4Jo7z6953nzJLIIDg7ymBac4haUoO93zikK1LhBpgCOpqfP5CYnzVtVoI0
W+qaMKnRPxDde1u5lvCAcU45l1jC/HaqtKl3vShFXab64F7ATq9vLpmbM7diTN9OmGXYyzwVB0Zj
XZnpvYrXWyFUDUYUqO33zzv7HpN3SJA51mMDCju57fSeAmH15uAIoOPaXHkjM+ivnNZurQruiBdL
0toqDsBVEhJVDLZdA9FT0CKudiji2fqynL6OF/YogFtUGVfjNGYzdg0hJub6OLMWiWgf9olJXNER
cPxp2EQJ5r0+5onI79WmURF6pDDsCMHeInxyMJ9Aof/j0YQbRcD2udoEDgujRfH6jJpyjeQYfHvm
UuoqJaLzudnZShNUv5gv8UMQ3pM/uXg0K70hfkGUPk5OAuLF8HKZ4TULdSJUxhUjsykUHQwAZXx6
L6uIcZsRKGUSKDsrQ8D58W9cii9KrCkKbJwZsbSSyG3wRjycdtNWHfoFTvDdiaYG5S1FpyX6K2TP
H+2gQzEBzXk2yr5aCiLORf1x7jr6adDl8lm7Z3Xrgsu+qe8x0mVf5UyROITtmrzg72RJ1PFk2z8y
BIXmgDGhc6LscLe6I8bbC64sVAl7QbHoL/y7WqNAh6ggsg1r16lLy7v04IHmX3DbKwWJDO/F17S5
hCvEXzEJnQm+VzQuSjYCjOgSQJIdM9TJHvqxFCUsM7Qf4lIVRWmG6JxlntdwpfGF8Ba2/ZZHOjoD
ks4sv79IEOnuRn8/tYrK+clVFaS+WO0b2JnjBjAsljrkotNbcpAEIkINC1js1ye2ROdSTwtIP1We
uQMWdZq6cFBxmHOFV/K9zfy0aFEZMwjMW3rn3bAJj7gTqwHvuON+Ts3457zSG04mjqsGoJpp+1Bb
X04FdDzO0oMa/sgJA+XtjDymOpkqmyAg07hWv3isdRp/UHjDPR0Mj1t8tUrXnCA9rXaz1xKOd1RQ
PgLkeJr8NLaU5z3ZVJaKpjeylaquv+E2RR+JAmZ9qlIl6iiY6Z1MUstHGIbAwGBcvJhabxIL6YVg
gJZMv/rBRip5MIZquYAM+qqw8VdQohDrUMIwAjj1IyxjalLZgQEPq+kUNLLr3m1PehjIuiJQjeDq
1pUNhhcWS5FjK9TQI7teLd4as9E7as0rNYpiuKTASc4WxwuF1SF9hlZ9+EJh2/7tse3fRzsqhhtM
M7wEcJ0P62wOf10n8Qeot3mwUMCZxu8Tb4gAO/CbXjo9L0p8kGNRAjy9HkD4apwh0RSVs/VfzEi+
okKWMxXKR26PUEjz+TtyfuK+SegLxVVNpY+1L11ZUW9cBDaeDCL++1XqhtC0lBSW38hQoGutPOEZ
DAKx5GBJWhCGe+u+WV7TQwyCHU1bbfd4WZMoupztHcDfP8ZbNwj/GOHwqO9Wqr0DFmiNkidgJFdG
vM3FW1RNPC/I0xJEekLHKoC3kD0wGiA25fMXSeRAdSWlFVwTRCGTU30+DLsjd0Loh0Slxu0liIGX
Kvivu70FqwVcQ+IxCj+eLCiLsZdMqW8umvTf1dC8oWHPYzl07NVWw9fOXFeMYbCyAkNqcalpfYrq
VSRbYw2IY6AZwZPEtDkCbNxbI3JyIJWXDtKt6vpJ/6RM+aQlhhQtd8nUYwWlHX9ybxOa/6GeIInH
7JXlnWr/vPNHouqcBuq5jBxKZnexngqtAfrAhD6gowECFC8rAgmEBxkYccWJ/WgzbVAV7614zSmc
XuFDCce0dtJ5bXn9qzymfkPZf9Aq/h9EV7VPCl4xhTN9gH2dK4aocnKqNdJfq8ECpeUMUSyKAiGv
IsHmGq1t1APfYRxwFu3gRshS6evG8pTPYPTi/WfbOiJpocUWFTc1eU9af5MbGGFitJjaBzjRVhvy
cQLXTF2wBzEcNZmbwI78HPm771d3rRxjxGuvoYRj1RvuLcgOIh5csZxg8HcyWeh+SRqEcljuDN2V
9jVSUWGbTYLgyycN3oK34TRJ8cmsXK9MM7QI9CVNeMVUM32dWs81/N/YJHrctlWmdOea41C8NO/Y
iW7JjRPuRkMqFhHXKpD2zR1gM7v7dPOVnO09Map15FoLxLu97YwWPZzc7aqzo2CEEEz73qnvymue
ygt/dZXoAnmdhhQjzv9Vfw3dqVqFSGtYNuMZIDkcHjwRm8EfpZx75xGVPRleqUUY2G1BtDxpnZBF
+bCm+3VmJagLz45x6Jlbn5/8h7nLh1GghCe0OCchsaKwWUU1FT2p9c4gL+NFVzSP/UPGyoZdqMsB
QQTQRYJnldcg7b75iH3Yndx0iAOcmjJe4Lg9VWD2VUfMJ2WZry6jIkA0Xq0zK7mgCs8y/ntuSrDj
/3KGF9g0O95Lhm+QYsAfO6Xje+30qWu+PGzQn2SuGoa1VFauY0sZR6xpHp4Pg4myB0G1ffNr2AE8
aNVoTAMYcXWFgaj53ZkDIOgpUFHygEqxzpgm30Uw15ydePuTcod2D8cgBB7bGzfUNS220MscIO2Q
9+uUDAB3cnCDhQ7DWbVey/17UmQkplvEyiOuMeFMbY3eN0ly5Vl7iWNeJ7FUY6H8UKjgTts3q28C
nfXsLz5msM92Xknm/buC56lrVe7MW7MwvbcVXZ/vFao7JtRi36oII7WXmiKRwQxiZznGbYKK/uuI
mVNch3geff1TAYkbiVwLaquzEph3gFmLnjWyjmIIiPqCAKHzmIyiutessMLvKSvF1HQg+bk5xDUc
Z1Jju+YKq+KSe9O2OJ5O8goqU2jUyETQPuJ2XCaoEOYzt2bSSikpvhdprH0qvXGkvAb79sCHG9bx
8YylxAqS6IXLl857MlYRkZgyb7hlWEC9PR0AvCMrypUCBJlfLunaGrJRV4z50Lpv5WZ+M2Lo5lDl
XXigadygfJI+j+KHQRHZVuUjdpyu668ds7Mg/28+G1ktEpb8Dd/UlS98BC2+mrCiwSMGewq0zItv
fK4yjnW/4ji0Ts7AOEPEKp6iOVHU6CeW7XaqIdrM3mpZcoJem3JILK6XyObSJtGSqC4RfAP77d44
MrljsrsTc/c5meXYx5bZK4rRHp+d0ziBKdZ6ujd/plavJDgjDEZPVWVNhxax5cRMpsL9j+W/p1YY
9nS+PMcLx05lH5MES0pnC3JSsAFnccQOrNlbBdqoHi7JJCWa5p2A+N4oXwA9kg27VFMXA8qptOSD
Ut9IwAVP1tK4z8804cHX0DE03a0TCWTiQ2+/quxfokmLjc9Tw2rCGyX4yG8g44NZ/ToQ2yfjVCT6
V9a4lpghxDurKDAoenWCvGUvjEGHS/bjGo7Xs9fzPBknNK3E70MHy8maybNvBGd/ZG910uy3KJ/y
sWBf6DRXwpeeUH2iDMfbk37ClLjG0KhEJFXs0d3hjnIOMrFDddjyod+4Z+NTsTKnGHh0bBZk7TlI
/nF8W5jBXSMFfsQhzBA1QHCg/+Uxu714m+xpL+wsOoc6TGNzlFEHPqRHHxWxFqURODvmYXbXYYnR
fa7uHwRL888iYueWsCJLEha5odxWLzkC8Qo9Q3fbZykUNxIoQrm8WteFAkhKjUrMWgkZDWjTYc7F
gNcT543ap3umsuGDUf9zTlRBNEqh1mZehZQfNGp/+5IsXr8xZXAySSTRLyURFEaxw0SfZLR2jO97
29P/5Wlo1m95Nll8Ct1Hh8BpSaDcze86FyuW+SFVmFMbkLv6EhAkqU9X4fKr/FvM8cctFeSdEIOC
zkdw0e41q6T+sUTbhV/SX2XJY4uq5AlJd4RoUOPVs35QeDIGbkY8kXPyEbPh0s53Fc+JKYkwy1Id
gzrZGOLtwnUEW27+qnO2ZdHwTsP+OmKO/ECPj0snC7AJGBtEj0Fkd5ba6yZBlOnbd7OBGZG3bEGj
w0P/sy5a/qFeV2oDGnUf35+byLgWSFTkfXcyfxaHBQ6fYeEqu4ve2WfvgxxNuj5g2szeWTtrGzmt
Znt7yW+DkNBgzV7qz4j3JK3nUcmpRKulCg368o1cnrIJTwLVvD0mqb0aF6Dj6pTg87VTvzosH+xg
CajdEDh9TQ8gFJpCCAfVdNacJh8XDEsuidirimdup7q5K0p4eW/+Ao+mHYibHs7jW02cSUkJogyO
XJ0TIMrxaK/NpedQIVLGg1VA/LBI44ZwmouNiS4szaQaOQHAGrS8FeW9GiWwJr1GYtiD/N5/TXdM
JlF6qKyoYmdB0M0QQUFoCrYcEsFG568NILRUWLG/Z1yHMY5hVTQf3GX7uCf7H+gA18oNiHS72kH7
EOi72RCpr9gpf1tfWPv1ZoHktCiXs+oOcTiSU7mdw5Zy4x+GnxT73RF95m+uoSMshOItLOCbhDuO
2ZRr4dDCaZf0F5BgotD3KQdhxFnbHcABU8pixNoMlTunRwjWLbcBvOExQxovbdUb7dM6tSYWUdsz
/JvwQ//ZaAm9CZgSoGDcBzMGasJc6FDhNlxpK6BgTA4CFNA3sFoSIAQgtfnVhzXty+aCHjruUzZV
jQZpQjf3HUoVTo4fwS9UyRzg+Exb1M7S7pg8WyNtI4Mseex689mQSzZHLBsVzJ5pquxUoZTjC/5X
KJPvvTtO76tFxkI25bc4sj1SZ58yRF3HiQGElJOFTReeQ7Vm+w0yGFR9I5/bTiS49clDGwtQdOsy
B3qlzdJwr2AL80hhZoDXGYrdlgjTs6R52JLbnDKEX2geS7ktLc1IVv1tYiDuzwfTNZ9yVUVz02o8
5xKhYzEL7eoyON1VoFWTbW6aaz77GNHwm7YCBnL3obanlqwbFGksVtEllvqUSntaRipDZWE2rLT3
3FewFU/oNigrJB7X9O++9XYTj9v/0qEDY3xHi8vcnVDDHpEsV2gxEcASlyYeWLoeQ3Tq1ROmxl6U
xPJ0JjTXCA7IYajQHUZ9B3SBlSKXXDan3iEC0QxlX/GZzzQYJ3Ad9+2cisqKvWiYWu6RQecH4G5m
CrwViXAbyu5b4vUSL6MY7Py5r/WzHy9vh+9MCCRuHGr5uNVL75iUY+HJqcIkL7Mo8yoYswH0JdTX
8waA8WKhhAkHk01286t3uNqrfFUgd6yvau+JUmCpPhy/CGCB4wi58nEa32zimQGU3d8DYpekq1Un
W/4d1hGcKHykH9m76SvlzlsTWX0YK8gTflBlErVnG4NkqBI3lzAIlQWm6U5U/hWL7wqshM35q4av
AbK9hrUIujcgdQVpvzpszby0IZwqvpbGnJe04Jr09txQ+Kr7M/9vZyw+IPiY5qJEo5WN+18DI2by
H2gpSldI8F1O07d0zEIrX347mldXIcMNDobPSFlhrXGaf/PycV9/yiApku/rboRKZVKD8EuIUuCA
1MVoIdGiVoDMI56bGIwypckLmazelGurzvCXaYTmLkYK1QsXhxkGx8vQ0Vlt/rqGCT9pDGINm5A+
lJAHG2tJ3qnAG2D83tBaDLY2bMZz9JURQhgj03qiTV3JWrMomiQrxC1sg5njARJqJTfg8lScgoFE
rQZBjQR2Wrydl/t5bE2LbIECkb44WqaSUOTUS3dCXvg5KP6GYeZtFGoTEvALoh7zLZaQcvRZmn6t
8hJkGv8EZaCGKvKBVQUjQ6rlAIeLoYWIyv5F8zJpPhd0F5EWivpKU11x6WKSHrLV4Pqa1EXA9LWD
25YSgdor7HoxiEzYyNHMktBNSx/fW9gq0rCorl22Yzh+yLvy4qBvw0oZlr9zqoe3YcvCi6Udwo/I
FyyLboYDvDv9zlPnZZPdTAQonQrh/oWfOF1Fk3/8CRQyrb/j8BZlHdLeJb1vBwCt1kd+MTOMtGaV
4vcPhxq4iX19670EDGRbCxyCFOoI/0ZvcN+5DnywoybbdDXcOzGFxp9ZTyDg4yjblsnZ8UPnnvnk
oBDoxijxfXTRcHVxIEkVNyVmyvgVfF/ZZ+lAtJ+QQ3CP+NNGZFAOihCOZ7p7lSdVA5H2CWsulBgZ
vc/O87YVG+skRe9rLT6fXq8gES/orcy4iOKXxZ5SRAasLJevY9HJErvIbUuEpzF984ds7Kpgc5m9
+ziIud0uTJo2xKfyB3LyBHqMABdVO5vB9GaWHox0B4migb/t5Y7J3UckmTRVuwpPyF2e+PWJq2KL
I0ZUYedagUerTGBYMXH+Hrl0D5+S5w1yKPLu/czdC37WScdFhd1AgplMO6Qmdt/KAhDI0ywTcRhk
ijw1X9M0+CRb4bZcuGwZDvlkWRfDLd+HbWjFoVFDlnBRWg8c3X12uVp5+TGWNnMOHW+5t723p/P8
24xTrJ1eKH3eSMA/SCc6y3v7RnVmvq8OBcMhQ+1YeQam/oxsvh/Uo60GUieOz9u4QdHUE97EOsVv
puehwsXPxCzWLCj6EvjuoVvK8DRo1Uw1IDyChXodyFd2WU9CXch02yVS1yECLKl8viAzoiv3Qpyi
EH1FRDQ1fT1SDaiG5cNoVJ28E1Snxsth+/jJzo5JDq1gr4Gb1l4t9grfTxM0XJ9K9ibuI2GaKLT6
w6YyEgreR5wKswNEq28OLH+6OqVGrWUh5HqcKoim83DlAziguF776i4qhcS5CWzoMwMbEUHzd3kQ
KOLj3NL3xyPpjTiziauJyUBAZ2NtOP25GxGdPk3mcqlVxvT0fNfwYgvNraco6PYxlsrPx4k3fn0v
cTU78hlTg1gmTILFTc4JsceWe983wbAYWTEiJ5awkg8MgfUK1BKZLQAl9GIwowTO6EdGAU9Xh6qV
4k0Vm6KlHs07UPm5yxzuM9WrRiqJhhgGiGrk5itcl2mtd5ap+Qa6MVvxTnUcdrDe094gZGKPqo7z
dzk3yzQmSC88uHIr8vgoMufEQGm/NgUQfM5kMDpz+rwQSb8tYQCG4F/uu1jjQsT0JmAugtTCsuwP
g0QRKDfTgNBD+ReCKO3ODyvUb5/kp2hELzigdPk3uJKVs/YxpYabG/M7lx9TS5NOG6hvvmWjGXxF
W+n2vXamFXdhp9AULu7hDCVr6v/OyZg2EGkUzfgbmyQWNvSKIEF4bbcAuDEJH4fyjC190Od4wMwF
S3OVHbyhifg0O7QNvPssSxoEkYidots65TdCDtVIJ0vL8GWJSrRR6xncDdzqeZmGeKwA0EiQoOOk
GiSdi1JVPaQFxRKEXK0xe2As9fdWYdpiat2zbFJnTj4LUpMJNCkM7wW6XvgYZIFlSoCFwtoVnRSg
EJnsZ6ywU1j2MjcwAfrzNyGn0QT4CSEalAucGl+S7xBWQcZ4TottmJgJGq1N1Dmq/EUHiLOyfDzo
Y7CbP3jX0OgUO8e5Rgiwrw04wNB++t6VvnQx4Gj8pgn3NXqfhnNYVCeTLmVKaUuP8O+EC2rw2KK0
x5dQZ1RB0QGvm9hEuLYaRGRdoHgV+ST5NQCdtkLgRTbpV4ZK+x/qx6B+xyvXAQ+nBqdHyOApQOgT
4i30reKYJ2i3pOfLS+BPCndbLZSAMUVtrHU8H3PpiwFy8YzhgMZOF/cPpnewom7gIYrAkEdDLUPQ
8mPHZ8TJEjjofmTJPASrxmkcJewN3eXfPX9zeaVfXzj+u89ujMv2tzg2xHU4/KWiXYo4ZXy6ks3s
bDJbrBTB87i+t+qX1ovFauQoqkd/ZJvJT4woZlKsxNB4/Y0fnIz24+kFA3CSGm9QgcsB6xNpwY/D
J6L2U2NhRSDuJv4wIF/auGyRuaMFYvNt194nDkXb8EFLx0/V5wlcplph7/0Vw6ALt54TUo/tocJD
PKAXy3gAYkI3H9cXBBIRMJjRPQY7SfmkxdYh7fmISI/h/RiCFxZemdN3kTYhT2GAMK4JSfj3jbaU
mE8LRTPkfnrqDo9/OpweqONDg/Gx5fVRSoHjaBMpGzB47qrufSQlOTGu7pHhKaFpE3Ed6Za6BrE9
ndV+es7TruQXdPSQvQOZmVNmrXhxvCf5aJjJY/lU7GxAgZT9VHaW/9bVz3FM2ZkQzBPzi89ZYmyj
xKS494GsA2KJ2NjJL6cgpafomr44apQDMEOT42cRn6u9IdifsOWiqrixTDOmoxSBWWAH5skPG6/K
CQGNjxXctIRFan26q7r+EJihq068oksUQTKjbmtIQkmHl9GdnR7/yRhGZmMT+sUpn8qGMpmzAZye
xina4xTrMTNExYPEctoUiJlyZVoGJHNFbWOkKysALMovTEZdj/rsVL3ntupvahb3gv88PvtGIWuB
gB+znNdHdE+I1x22qRiq1KZNL0oVKlaKKRR2xILWv0pUsD4ZNltonJU0esIo5mwYp5jfp724aTTy
INFvXzulQ3XaYBmbMB3GTcDHqW/k/10aYp3tobV0YqiBNkiy55bzhCO1ZeJkOdriipNIYMoTL5pR
9LQOshch3tul155ZkjRXXFOIomCggYtEG/NVBm4WNLZqxFobnfqbuqVz6zg4oDyLOWkb+a63FIJG
GztU3BH7wbV/kGOaLHtKFebZiEKz7o5X0g2O0jKBW0m+PFjTnpEn5Cw9qcft6GHs2gh9QfDGeklX
IFqcwPqLrewbdEaC8V6ddpfT8XuYOSA0XXB457Ne0LmYMBhQ9oJHgjcXdNjYnsjKnkOiuD6XnWAN
YAnwM9QJ8fMSiQER8Mm9XHX+Jtb9gLotY2L4dQgH+RXRtnkovFNfarLMdvQppSsLkTTFZ5yyyr/d
PhmHa1wG13dHCBGUdYQNN54hUZqXJu0BNIcguXul7rHoaqnFw9uVU4cFFX5e438D6sS7qha2IW09
Q2Vw3JGVc/eKgm94k4wVy6mifuoDug/Hfbwd6z/1PPFadRbdG3G8YOhfg57hhm1kVyyQIn/qrdzY
8D8bGVGlxqSXOgQ6o1iwBYyAnzZEZtkEoXS8A7+wvEHXN3YKNMMZkYzxMptY+uh2dMsoKxzHT5tL
+kEuh1SU64Ol0DMVuRk64kjCDkNZecRH6KOuYI/f/onsavzq87YI66WtLGwSqCyTlUYRYL6w5jcW
5ENE+QvlBG/7m1FP0Xero+B+/TeuH/QVGJlIe66GyE1U+3noT/aNb65dSTH8lq2flny06UXOwQXw
h5HSfqz0N9IMzSiybipwTtfIKRKpS4EY+5mjuLH7H+WkBHBa68lpplbUtfme8DQWdVmYUFRANluY
NxwQgm6HcRpvRrhJ/OeubP2UBDuJvWkPkCSA9oAM0kpp80YNGhJtr9h9avDLcscT3KXLrD4bVtY/
1ETfhJesachIy/Pxtb5iFa8HvV3u8vlLQTQaa2ojDxCeORIC1xs3a5BWwyc+xrxAP+9otVd7dxt3
5sqcY9kC6bq11P6YE9DMc2txm2KyrWGRdr44OFw2O/JIOS6JRPQ3injr2V8YWlE3ACLAT1BM/kuQ
HCgsZo5STYhnO1EVmbsS0JGbZwsaBWvjsGMr8Wntvnz5rkPdtd9KHSOfxNPYdyCVAZO+3kK35UJW
vQ+LwvYKHh5Y5hBBWYzdGj3oyG7sC/wGEMxx32S305VsMt9XQhOZpZda32IyqoN8hKeiLxCcUpWW
NejVSGgCWf6QAjX8a0zlYh6obyHEa9NUp5dtI6vBbkm5yizfDDMZ9EF1DKkU3+/zCAZim94GuYa9
qWQzTWwvZHCeWea5SsWFoFG1Vy7rlPitnZ9WPAdqRtZ0usVwnviagirgCREEBymTEVa7IztfyAbS
LqrESKceTtrV8kNcN68oiaJcu1iCIiPt0k7HAd/mcsuosW9VGtSpKOWOy38/obhTCzo1N6hCjfXl
NVawB1xMr+jJpuOCXEcElE0bBZJ/xdZ40d+B0e7jsUW84Mh+ci4DWYmO90Cg4acVJc9W/LSZ9zTC
ZC8y3RH1kbX7p9Yqd9ALIMHOXX5wrHKq7x5Nk3XiFDU8tJVbi7yxeg5h7x0lrewiCI34AeZ2se+A
ECKTMNFeJFK0p8iTsLGy7KdoliC2XIO6v8H0V78W+cNk7/w6gCglwd0yRZsZGJnVY1qYCV9pcOqe
SwfTa4mXIj5V/Hwz0eo1Y+6IuQM8rjX+GfUa2Uz0lhICnCTYMbizAOPRyGXfA6O3JQEgmzkpOrJ9
KkFKMnjtM/yva7chCVYTCDyCeuO7jJ2l97dAznJ/6H5udjh48tEghByxw3bivcv03mIrzigG1npQ
EBGYFp43dJ5KHxHYg15yAEtiwEXj7ANfPncn3wKQqRIy+i+QmhgmcjM3yJVjzreFExBXJvX0nv6l
QeViz/rBA/Miz9/O3bcoyOGqnLJxkKcjFWx6a3nPBhAHRPxj4hnhS3bMABB+eWj0cuvo43FEXpCW
gpXw3uZR2fbS7QI5SHHRh+1N7+sSyQ4jCMzFnkStKIpKwiz8h0/sc7DCDmGL36mYPcrD73j3onat
53nuV102rS7CriEZMMXfkNoFoitUBwe6XoI54CFoJglN84Agg20+N2EhvhKph1nw947X+i3RlH0V
60Xql+vT8hlpWHayoeCk1rEaQytmQAA+0wFzn+r5ogX+otwunzJhXkfsXhVfCuCUJVSMpJtDFRzb
UtAiMAWjHnFaRNXGkP3NMOmmzzec3zZ9HEaxsemHDtQK92liPMj6Zl8bMoeeA9kMxX5XKueTMIER
1/50AUyM0ORahySmsnHYuI//01ILJFg9Cy6hcpxFO0IZoeAKjuahUmGnCV3tpU2EFG7RRiI9AtL8
vn1hTMxS9ejSiWOMnajZN07hVanfuGea+Kygha6Di/8do/wImfzn0KIFScmmPEqOXCjUYOT+yTt/
f3BGJTiO7khiFftCBKHzqXmXcNYpVcCvvaYkMUmy4X6Rb1cg5td5zDPd0xIwKL7EMv+OpyrgJaCp
YOo4ueWdn6FUoa9kAMBcJoIv8C6IPuLQrd1PrdbT8R8SNFL3YdVluLAtZ3GPudZZh7L1rnWPSVnY
bKA9EX7dv1WKUHD0MMHpDtj9A93UFGzJiXB9VK4KKm2MQHET08dWWe7T8DPVt4LxqeEdBVwPXSww
KqDh5pfvuuuIwGHtoCQ4MNIcKu708aLcmMTEMbzJDGlWlIFzBokGO4Cpa3OLE4b9vadpn+yMPuL6
dhkATpuO171muePcwTsgXmVT+A+DRh+Jx3qB8j8NKzP8Nlh/LCan8vNQXY8KlZpzftPESxP+bRVe
v3bl0j3N0/gY5RXG0UWky6N+7UdHqCh/0MDFNCsO+mJsJRRAD9jtTkYh1fNmY2HvSObYpQpgzbIt
+YOLnjLVjtEtNvb1mexe/yqJe7TBpFpA2XAkOESP6Jw864vbcAwfs0+ziklhx3TV1UjjYkwtjTUF
SIPtg1N3eeVPagZJVo+ky5RgU/x0VJJ4kI/cM4fLEY7WnDM4W7CMEun+pJ7dLB7+RVg8FvZ4D404
l7Z2d1Ob32qHN/xnZcbKklS4zlxdQk+LWZzp6rVGfK9hxDOJRlGafL4nD6BG49MTUbscPjRw/J+3
MtyAlDdSPLoz8TbxYgeBjgdDWo7JZaxO0Au5B6tkFkJbWXbm8rUiajY14EDrDEzrE+cBI0O1xjM6
MQ6PMVUT22fCwfwGc2L+f/hWD5aqM8hFdW1Da7OgMaQZE4XBLdY2T01663zWpYvQesuW3cGaDaeJ
xGkpwAYRMfA1tpSu8waKtaklo93cW6M5zqJHxrunEf0lK1PTYK4oJorQZXQDLMdtU4p5TGYrcKMm
S2xvW5+/gsyfjhVbp51Macn9S90AiwKi4f3AUSMbw6D3ObEXe5sWAqJXrJ4uRvF3cZKylr0bvDXL
vm2CMCO8NdfFs+A9DSHLjAhCf7OzyIKJOqDZNihOGZ/cYZ3eUKhiByCFwbUToPP66lGwxW6GQgFX
yq8Y7PMj4gKTdZ2cX65M7qm+NssjFNztuAiRHYQ+kIcudSU0Dpwhra1aG3LP1SIHQOswzl9BOWwP
hinmJJ35OyJOcZy1k8FuqsMeyNZ7G+xAr+7vwSREqogTDmrZGLZlGTZT/r9dXXDw6mInG8ZCiVB4
yOgySDdZ9NZR3tklcI01yEcm9aloEF8kU57McSutgyYButZkkFvNIo5tiRdfRICGcOIpV6YfonNN
JqqgSeXisSZUP8O9muB1XFbZw2NPq5xA+EjCQuSE3rXZ5iX4q/4/xf5FgnbsUiTq6vUG30lOxxjH
I0ytcT6AqdYJn0M97Z2FBm7HgA+RwHM0CVgy/QzPdPXtR9H1Zg0VqtF5CQL/Uzh5t4YkvpzLA8uS
CXKccb+5X3KnLWdhmnaJLjw8PfQFApQgM2Z9CEDm0cUa4igzAeHDaqvx18Ui5u+YX6Fvsy1Ad/Q/
PMEwvxAB/a59JlpttMvHvkjbdIO3RZx1j04sFeJi64gk4erv6/aqsnzyDV3xXBNCuITegQXcuGK+
cDWDFVJOSgE+eToyEQj0qw7fGFdmg4WymTNYjAg6whS7XyitBs8shhTxC9c5dXPSOFQaNuOTWpP3
gfk9LX2tCcw6OPclJUPnYhxrtOrs760BUsol7j9YvReENPaL8SHXwrx27dMPvEmvP/zN4Ti2hcCw
6UOsSPGAF0tYaBem/TxESzJ+nQQbewudZ/aE+9x+FxqL2cyvftBc3DIyBetBxnDtvsOrSSHmfzPq
7VjGT9sLF+kTVOXgyeCHZawbTHGiAZCYRNMvDpu4Iu3OFrZhCDobK2qpkhW/VqhnQK38AY9kn5lU
+Gfc6YzBETJYIokFQKGwbE1J0/y7dXvVh434jXDEEAHemOC0T3fYmuFq4lrzS0QRAr97tnuyt0dz
JmYzdGQnudwuV+4yV3YVIqlpZ8a2FBmo1CAHLWh6FwCEpjPZai5o9o7Y6dFRLvmJQgmwDCBgpN0b
LZrmsW/KQKGljaOl+j8b96anNubwdhocbDezdlimpvShnUpUX99Vo7XtZVZjUAkER3WlCDjHCJMU
RzPXskg73Hm7RP/CQHH0mog0/QGUW23SNW83hnFTVzwbQ+1C7gsrduNrCXrY0eSNid8jtZLE6iJH
KsDJJ8vyW/9iFj8Fk24ZXmM9DQgnU6W+aVSD/ZtibKBuHuQ82O7aiXxw00o72q0VQHVtn/kIlFwk
z8fFyjsZeDrVZ0D3GyhpWziodbrHIr02nuJRpn/lWxx6wsAbr2uWMVx2W9+FrKX2mNR1gA5aZYTz
jSq5XoXpKCawbPj7ujZ9jo9wjquU8GLBfiF/5exCSYyEhLO7SDNMpSMnSInMvLemRzLRDW3X+WBa
Oirqu9wkvgfTgDZUSVXa8F4MnplZHzXUrpRTj7SS40sawuG8/mngRWTT6LVLkST4Dr7UIjmBBLq0
6x885iIpGH6fF8wqapzjUFQbUV0NiFspXnCicTgB2VJEVLPbiTmIwhk5HSa2RrTAOYyJuROYpiLB
XHLDOcQDX0fcRttHmS0RSUwH7puFLXVRUySAI/WIbspl80HhE5tXutnnpKmDkKKaiY6ME0sBiDFX
YQzr0ozK4Hqjg5BAVRH8PQSAt5XpKfLPWeQD4fjqAXiRNwzdszFq7Rv9yNMwset7Jni7GnAVlul+
7/Wdu7AKhHpV4sjS7wY1ohOzpo1XVa4pmjMrGNt/jqMRyHLjfnEYYmJ+61SFcJcFuv/pHfRUwOC/
WY35B8vGltGnwhH/59jP+EgOtYQYODPW6lPCg80zKRJXYJLYavWhaa6YOjHUkJ8GOFVsA+V3XkPm
oMW7p+ieYuyvvMVygl8g35uUqtPnwT9GXOHQhomzOis7evkRrkEOdGsp2zK6RUMOGM+LgUgbcKiV
QYigmpFmd3nWNFmSA751qdtkM0t+0Y+ryFaDhoqcZiYmggQKrcao6ZasCsfXhfvHT8Gwus4dj7ut
wWG5ao39zpUUQXvm/Yp0W8W5khQyLDAvcoHNcllm6pz3aQVbpEMruerNB+0NHnwSY/BCigv9LV3x
KLI8K404aYZRsigR4F0y5eTQb7MGWTal6LBntthSPcEwUWthMCAFMQHJxgnJ4Qpr5U7cLS4IPOWZ
S8rAB6fMBVeimUA0AAgdfVx/YMwAmsSrdbPXPU92yoUa2Q7LWnmJIAApvm7Oo+26Oe/BnroqDVAi
JhgHWI7167OtRSGBT+aCCxEsQsfrBG/AvG3kT74qz5YUc2lkFVVUZsGG4rgdGOpYeU/+kiE3Scbd
qHc3zLtoO8fd0025an2wwZK6g/8Nms/4LZpY6hS5OfqHZ0bUYeU7/FivXahGnZA0a5ihspOfs2Fa
YimXEdrnYyhYNEvSru1u5QPCtrOO2LPM1Kd/tKnyx+fnPvqPz97jQsbsgnqugr1YOhzoIRsAvn9c
HVL77HHK6HHzbrJVetHGz517kXEYm1jSe5nRR3q16rli0aUBEcYBUjPQkq2zA+rzS/3jteq5t3O4
VIo2+oiHjLHBMVCf3JJ5vN4Eho418a6AIuLUKHzaShdaDSBXh1kWgHxK99uf0l9Ph3q7G0n5MVdL
IccdRmVHx5nL+2Fzmqj+nFzgPOLdaFWBqcJxs88f0tSZizuGB5OnL2QOFAtf/cEx2qX+5Xiukooq
rObFf9di7AloZplmq4nTfT5cRZZZ/E+f57EDDbHn8Q9gCrC/srQkRjz5bXXzE+eYZyRuhUSplR1S
E0lqYXyOFIiAD2Jo3lFfsBDscWHfb/4BeYy2nILhd8bXPAh7b1GQ+NDmY9IqRUudrqAwYu3zpEwd
lN7dnVzxLnkYIV8w5oudt6pcfMuSNN3IowWY2urY8YGBkiq4Hbabxr6HswXTlgspvWv50kqUNcLb
Ju9kXSz8H6MG3sKDLoMT7BMOo5KV3VInK7Uk51ThfwtagN703A7l5KVBoehCpyaWSsBIyHq3MtLz
V3/rA77sdF44vDzFub/G4x4Y6zUXfrrWNzqYoyeAqzJTZZUrbep99UeiDxaTyPdQf4Hdwms2vaCB
GKQK7RqYS2ZnIwk9VAu7DE1+q3Pps/Qs1xsGfMd8x7cI3bnQ5nuEguJiUQbiUGL7ImVRI5dvcKyk
ZeAR+EI2HYxrbs1Iwy6DiS7nfkSBUdZSPdnTR1v4m30ucn5hpwl4k5x1Pji6dCmj4oJ8xAPljtNV
QnPwXvSIGSKMFuoBZLa9WuMCnwR6cIr0BN/r5CKRj7cpDJfBsWqlvogtdsWGGeCg1Mpe2rtMmtD6
yHWhrM3oo0BXBea/3Paks1+M3QGaj4jX6f+ppU08J2BHwnQLB5slw1b4jHjO8QuTo6sfDCdocO/5
CIx6Edtz3YPn62dZGhGdfs3KF/AixX3JHX1rdFSlVsff0YjdcL6EVOAFuNh+YvxrrypC2G0CRGOd
7dHUfQQNwuHyyLdFgJkjAJ7aYEAyjk8CmCVSVu0mABcp9BtCmRyFsyxNDUdgSGjpYhu017Q1/YA9
Py/OKsOP1DRs5jNpbvZcTZBJSQHYz8PTieJa+xTonKLoRqrE9zaiOVVNeoEtVfRVnv5NNVb2pkYa
GQG7ZTrIVMflmvr4zmKpcKrecsYm9ZxLFhAGCm9ushJ03XTUYIp1JUI62PRAQjkrLo6jHu4jzxOk
JXawQHR7dVQApk2UHsaW1O8wrUMObi2pxB0/6GWOmmx+G0OjDKxmVVJDyNNXKspzbcTJdB5ubvi9
J6mp03Xku0vHIPhK1q3TEYvYupnau4kxJDaVv5KdaMCM0jXQq3aGFDJ2xw9c8DH4fWrzA71N1rgt
vT0ojvPvROtVC+SyJk5VqxK2H0PKl0atKrMJf/DUS8ruUIsGgN8yR38Y5+tzRCbt3GJ0Zlmt/iXO
lL7NL7j4s5+iX2o+I0eR4hgYEsOOv/R4+TqF0tky5vhUOele4W/cVW+nNXS7pcjW7l0+cTYEEaRJ
cYY84i7AQ77PPKdn3/FP3XYLKKqQFN3BDe70DSqRjEGkiBJvRRMFBdyDRWsQ08j+JE9IFwiIuTC1
EUJTKFqeB2CYe0KPPM//R3RYVc3H7zAQ01IggjyeCf5E9EayHPBbkN37IVFe5OK+F6likRY8HkYq
4vgNyHKrm31B402RkqxxGTju/+WdydQIr2yW7w5Ft2qmN7ZSi7/dhpxhn70KjTlwj6Iq5GP5s74G
v9X0cblqsk7kUg0ro3EiitsKMgTpKrM9vLpHDW73/SSYjttGPdZwwGOUDwDoClxuKUMfIPRNAUP+
MObWkFCv8YWwjxO1Tk0/OKhN00KAWWkeAvsEX/roDvNmcPeowxb65kfNA8ojMyiXSFMPkfLn4tQ5
u5GWZGx2djj18eudpv/AMaBjfvQOI7cvKca8TnTVkqimsZjFZ+IUwaiRq45tmdRij1uSC1TkJRxj
XLqNpqB1L0I9ZEYOZ9e2aEYXzZV1vkuEVjMuZv0iGj5Ljo+mWka2026079lqq5Bc2oOlTG3ltk4C
V471qPqYH21Dd64mBgT/+ioCW6yjr3I7P0XEtVvgSv827RFp7D4DmBkkk8qzh7JU90b1xtORQy30
/kF690VvfYYf6LzPS3BKZ9z8D1paOCy3AE61uNPX2RmA8k28IqUotiEvmRMSAZO8bfLljFf7AMpg
6NEctGXfyYchBdjVsCE/fhR/tpiv+T25UcXQAvD9cV6TeTHDPpP7Wxolgv8ldc0Ux3FF9flCSrV3
XmrHh1LOJkAkNOAyfuFl93ZHQRuOHr8gMKIuzFFB7utV1vNb3PaV7Viedt89HmiU3gVoKDsw+w8J
cfv/OyczjZZfUdb8D2Dx5kftuOelsCGXYGTb/tRXkGjkqAEJJERLbUPVzx3aa4xfH0To94I/clbo
5Jmp1pOcktVy8xzR22vrR4bFQeUyoiZjnecLm+Jf9Vn5ITjjTwcrKuxYU4W3oM+OgdruIXB2LKZP
/CcIXMLA+LCa0+cf3jkd8qlq9I8HGFgWwvYaq6QopTo0a4igimBHhRqLeOUo5ZP8NlIdndXUJLD6
8bgUw/ZY0aDKhMhNWnNV8lvfwiUdz7Zw49TIKIxR6022jkq5+iaTaKeI6o3MRjhoSJskWxIebCkc
RWOxGNhYYB18aFl4UimUKqydc7ylhqushzsmLDa7Q0K0FSCicU3yoYTeUpWzXx8Q5H2np1OCKUDY
2nrHWnyxgqazlDJoLf+QjB6S5H/L/TeSbbZ7YyYwHtBNWUvFAM0k5HYjdeVyqTXVlUt8Ps5bIS1d
6oQq/UUa6xdYugcB9LFl1sAPF3Tl5xlbBR09pkKP0jksWqLK1DfHPQkzrbvLCnR2a8zpe8GMTX9j
3ee6/eNbpFTSaVKD+kZ1C4MS9ut6YMKTONynHjtyRzxk+UyfvGu9FQPPb2+tVpqaMnpC69qx/YpX
s3Kc/TExHA76gIx6U/j80liI0CH4jsnCYsr0kfcD5l/gpXVG74sVOI+6RWaOskStR78cIVCLohaI
s5wWxcqQQVvmMXRq4IzU81rR7PnnbyBHdlt+kpLXezi+lcwN5WcqtgvhPxb/coHIP2jbbQspIyju
lRkuCpZynisDMKEpTbQ6AF+gnCmRgp0GhQ9UvrhgvyBFiWau/mnRmo1BHaKkt3TcCZLDBLVNnTEb
H7oK6szPTadjVx9+EdlQ1e5ZvhTaElXxyl1EVs5uYnfcNOpzxoeyCOC+huO/OypgIwgGSpJ6x8fz
ST1upCJe6em6xWdVlQVrkAm5xqGjQslH78bh6JdlSzhRaGRhGRP+t3N3hB6VQi0JiXdU97QLeyq1
dKVCcdHDctePNRAad7ARUg6aK0vvjjqohCSBrCEYvZNqacEcFE2ERefq3GvvzzI7fnZVDQoykcIm
bz2E0kmNNG63IHtkvJE+AqJx+cWAfpo/9mVItsqVGwt8/t2Mfv/9qnWtvwmgX8OIL6tkPG9Eh6lF
AY3DeMRUSEPLeMdNirLhEIbeUZc6HUBvDWtpUreJG+vVonPJhxAUE4fhe7leS5E/eGMbwsopLy0x
lFs+PFaJOfa1tNTeZ6werUpX62aoHUKvZDLYnkgC0gUDlhw9mBizove9jk+UVGovLekaL3acuigh
/ic68JOqJMFGhFD4ChppncUJz14AgwXfjn9CGRjc0STeg3yBQ0LDka2qyVQrp2MTiDk1o6mCmXNV
DJ4n1iAOR9oapoN2zlpuZ8NB4XZs+4GBsHJ/wkhrLxY3sifWOGzr/pUQg/zy7tQWa9TvkHbOxd7H
e4OAJSvr10Fsh+TI7wDiN68ymco8G/rEzfbpnO4/MnpHq4YSde8LnFvjHm1jmVDpMwUaEMSp/3zW
8l4tEMx3KYa42HEXAWhUcnNAnpc0sGVaeqtQzUGNQZSdrCMGig8zeewNUnBHFZQyd0ABGP2IUiXP
FT7+AsBgvVdea3tD+VaH1WO3nwu26TPuytseEcqNq7ikCU91FHC9072Q9wxByPaCIUJp/kiOqMGi
AnY79f0KCotOplit1b42S/STGoyNZ+JeZF8jGdzFIvVTJTS9QroChwMxO8i2qaTPOMKZjQaPVzmt
T6uTFIdtpqQios02uIjx48kYCshDAWpfZpHo7lE5Sukbec0qfpKM/1ra57v454kUAzaDy4o40BcD
IywuT3lCNy4TOCZblvGaOm6FYkUv+pvPe/3KwRZhhHW8lvfTdEuBznL21HweBhgs9ddjY8/l+NKp
9yclno1BdGQDY/cVr2Z/c/vfEKHtHWLINK0FOQAxKUo+0saBVjAZR0mM9xR0JrQ6XsswdGQlfLoH
08kGeQZXG9BuDN6mwYnuVO5fFhVDIDSC1/6HsTkxJl6mBzL/L07X5Vedy/58Wpbk0OhKJbv7GYjm
LPNa8V7o/NYPu5ZKFvHjejX3VxOTTY6z+/ao5YPUUFbwBDoj6OyCRm2mVF7wvU7c4FeEVUkFCsKw
I9Sf5205m66bIsq+NwM7dl74pQ5KYvYfF8deYNppVzMuAkTppPvYHY5CNnMSm1DToR/8Qigr2xlj
XPWfn87tH5TAVp4EkbTmttG2CUW/u/wDowLUMCuJyJxPKMKhWDhtvbf1qttCvTv0lm50QZMQN45W
6mWxKUh9/kfeI1fF83U4XG/JaHanXj7T/V9hRHx4y+1+VrRfKT6rvaOnEoud2rgs+oKHOajANceP
rUBqk64we1WtyRdFt5DkuySGjarg8mcvdL/7VWXOz+Zb0f3vUGflrtO6g5eFbFjdXfCeejV5ZI0J
iRNcxLcuKGMRdSyIKjNcMsjAPStPVlpXdycpEPpTWOEKjZU6Yv/PeeKB0hlKqWzdscuVC5zyIx3R
d39xtR+lcudgCmctFe9XWj4/ZRwxpVat35kKplAU6tKFmr16P8hYCBz3nPgK+9BME9d5g/cums74
J/VS/O+7Q811v1vMT8snSo1H5Iioj7+vvNsB2fwp26of6Wepy/WkNGwIsJr7O7O5MdNwHN21pa4r
TlAxPRltwSKFCBofngp4WNhHg8qIusUg4NJ+hzQXHnMHrKkNs51sDYV3UNzR+375wbk6XWuTLgVk
JbQOY0GJxSphCeAN53f8XDSxScGxusLuZMfmJp++fT9mTPwbLIndjw86yxLESMb+sPdgvEdZqsW3
VMNcLAdHaFDJX6pBYFnMdx/CkzwHT2XQLOb9dMGkZGeFSlA7yA6g7dF4V3bZWCi5AS1k7rBCNAF9
d8nt6/An1rdPgHIc0D1IKRZzjfe4QjuyTMhg4+QM/+3icGCOnsQj5BR5a1Orxk0NzBgj6IMtSlRo
gUFcASIY4bI12LTCba/e2wWHtdXig2kx7Gm7UJwegSvkrGcw2CbHO761Cc5YdqZCHxB3vWQA325M
Cw3CgGGCjsXr8YVwYNfD36mFcHrOxfzv5Dw9uYjlJehk+WozAoIh84Umonkqlo7u53e+kqcLMUSZ
i+IFNqOUfNrEcVeAYZ0ziQLNi61T4UxZpbLMo4khjKpkl/r1Tljj8Didw3g02VfAoegPUkC6dWuJ
54X38G8iHJERNQeZDISejkYemyZej8cQ3ad3Jv8klFypE6W9em00mqHdMPIleasnEaBfH54Pc+7/
9LVKM6EWCRhkpPdPLjJnvGgcaef51szqJzVWau1yK/iSwG0OMynvtYqE/yOwwT+jKzMxO9lm8Gh6
sGXG/hu7E9Sg8ZpZSKF9/ELzzXUPLqCPB3a2ouLJwrP6nnfv7sCF50DItkcEG1ajDhjkjCV9x7DP
F4Q5JFrl8ITqkBeV9SLTvv2w7ko07xWX61dqjqMk29jz6Ovzt0AwZGyKuxjscdM3htH8zDFF4CbD
o7jZGlWBqlGbCnsC5uyrnWPT91gyo8c3hylW/7wUhbLDmnp0Jmu8DL5qaAlJWdVzymia3YlmNFrS
5ULf8BrDsqIFPTRgoLfuXe4CJOqCGrHPWChrSaTJy6uZEwv3w9DwMRbUcDS0ExwhrcHiyrQOuPRV
eNbCnZxHOgvPj9amhL2DNGF6w76ojSDrbcpahGlMEzGI7QVCyguw1XBEyy2kR47bD9W5xZRkb3bW
UCOZ9/QeiqH8frZ6f0eNc+iLMAgqBTJMrnTkm2ZdGw3JWbUelWoNae08wh8pSp6LKN+piIsCknBU
HZHQC7hvvRaxZ1+LM10bkz+2wMYq0UnhfCkyjIYtsY6WffEUY3baBskgRSn3g/SnJ//MHz7r0ioD
EifxAQ9nAPnrMVi8MbpxQ4VDBrbPGjpUsuiRJxcie/WCyxWwrWquygJDJhSWEVttrdO4emPO6tlc
Cn5kGIMiOymUP4kPkKmVZ3lF77WtYPO8bAtl22RBJeLmPq4ZjBiwZTJA8hsALSd40k4IR84hsqVo
tyjSLNINWGQHfyoXxtyoTia+8sWkwSaVoKNCwLASoaFG53pqGeshowvNHq5mlBdFr+/2z0vgobBP
MUgzbA29Z/oHSNr4qLY+kKAOYbbePyvnbxtfURA9PdqeA3/wrCK7dLxPZRBJJSBCwRvxYp1HBDyU
O1uU7IVGvM/pnj79xGT9BBgPyK14rlFXN4iIObEYHW4qqiaySJm8G3gdAWItqIxnRCMIXrEkXScN
TDLwWNPym6cGIjPSR2cOKH9xmJcJw10HGkDdj0WV7RGipdglEp0Kmio9/1+UZSTPpDsA9ELQBxFu
THjNWyp3sd1KDfVgwgsXHUyb3YHaeU28iukkeLBLFU0FOr6UD1INExcmQvgEPxwTv3jSPTHk9zxh
HEQCvpkaBp5sU3ldb/0oY6d1Pq7YdahrBVCqQjEThQVPynWw8GhWdB4RtMGYEU5odVPDgFxrA42e
sgpoOhgbpyEFhRcE+1vromwKMxtDnFjM3lYdH7AnGg/N3wGLpSH37QBo+usuxiv3o90PdGq4TjAI
s0mfHYW+zwWn9VPrCd9yHIDZmNVf5laGirmGzN1DJy9mgw7RrBV3YclakfEn3l1GntR+g+kptRNY
IZWX8uCE+7knW5hGuTzzwm9EaNs3reQDDOoRZShVowf30AiSh3E/kUzhTbja9PB4BtARaBG+8bJ2
t+X7IGWWXUN5GNaiEwHIzWNZTT19uTLTJXi0MMWvYbvTZw32Vjh7V6jG4e3MVuxg2cEHoxXX4F+D
h+5GYZ18NE1pyt/u/Vt+civmas2YfDs6SOG8BYE9zK8kl+WYUlGVNGvMY2no4L9rI98r7224Oa1+
t15FC37LdIvVhOyKLuO+vodPEQq8n8vp6iLurzzzyBNijepjsqr7+HEoZ37DOfgGz6Hk72KuLmJE
Zq66o19dC5otrP5RyraDTqmybj9+LiLnPlKlBntJ7+G99tTnQCWAo5stWLk2/+Ks8wX/ezjn/04U
+AfIscoERnme/b6KuSWKkJQM+970aMR2tpDoSEowvTAxx70/hnFy7zibxg/oZKIfU+yfEsfe0cyz
pIPGD+dyqyEVBVh2QiL/xsMgfWhxykiyymiT5GdWi2aR33XRHTweivgD5pi+LmMzlZhcWUv+/YTN
RjCr6kW7Pk83YY5eoWWPUoUu/X/4nmJF83Ojnm2t7syLPkIXRZlBSxSIBwypkOud/lNYouIhSKKP
pB61HqZBs4Z8n7S1qMWVJ3V63H38yhi5LAlBklNkJZ9Oc7YFUAtK8boCIRxiec2tHibJ88YkBhFp
VjTQTklxFwsVr8ro6k7ETSO5/NEZZd4amy0UoEncZmA6FOGpi+NyEzjwciTncByckY/zcwTIYsbb
M8nM/z+izaTeHJorpEE/5PCyTJQgyFSmy0QvCkgUbjt2BOLryYcsusDYBYk29b0Qjoht3uVtee1/
slwl6T6jf3bODkmQeX/5KgKZ4McycPOuQd0PVEGZkj9aKOS3Kkx1eXuq4ojMmvuOnkIy+vqb/N9T
US5wHQm7NdVzHCr0reDxoolx3JVMx8r3gfzVaiKReggVVwzDa/c/tpGgBlgRvB/fBll0uSENe/Qg
QAEJJemUB3a5IP32nO/8GRfzR7loXqZ2wwUt77R6/hfJF96kFHGxrrUOQ2iflQcUq6XNdNi71W08
EBMan2BJOC+eAdPrU/3FRCM2OCiA4fjYoGLYwaQR4HNDfWN1C6mspfh1aiziO5zQAuZxHjnCVpyj
9dk+I6XBqrXliQfOX6bOZCTIr663o5c6pc+GyW0c4qlq0GzMZkrQl37SjJtNdpAXsmHa6JrTZU+5
MxwSb6cIqeeIipZ3mva9dyw25x5zT0d0x1obGJMQg2WDZTzyW1Pky2rVw0SQjqqCi6dmC+RT5mBR
B3Snw+cmEVFuyWo1DygfCLfyW9aESq7NyIcWPCQIzS6rArBQCJvn4vLdbS0WCW9gbwqBVpEvEJ0m
07NqSqkoFJKcFfewWTAwvJbHzxsLmlFdD8XQIkHMGVcLhS+caQBNdPBLXvZB+U5HZ8Xk20XzDuox
9KTtkiizyKIN/RKR4iZFJdiD9vP7mEsULf3tLbQVW5EEi3rp9rfXnCydI9FyuOxFUms0vbghYjyJ
3lEcqRSNb+a3MiypqM623NtzIRqESC+Pcp0p5Jk9Odj/qNVwH+Q0unjL8v5bZ3x7XwLicrMGLIgh
0B9p9QqGhu7BCv0URFprHMYTWB3nGPdN0WFPt0BbVNXjZnfIPU3R8LF7pzld6soohDF3gdYrNl9W
13Q31Qcvv0lxHA1qyavWCz+M/IgkT+pJav0t/fmU+PaIsRq6Cnhup57Gsv+/Zo++Mpldx62blGbo
8Bfs89BR2vTSYphjKJ7c63jbQ5zVaSadGW7xU0z3uxOKBOIoY1m4VWSEnV8iSI0paWmTry8KXFWm
QaT0lQVLgZF4hau7zGAJvc9CsFqqDnG211N8cDa+SqA7fc7cSclJGHKnqMfcuXeDvaK1Igy0SnRS
CuLaixBmfLSAt4Zq5VM57KN6h210/Wjeb5fc79SEVlhPA5kwEZCoL7FI+apetkfQtlYQrs6wF71q
5LNeS6gi3HvxHniO0AisocN+9pfk4DdjYpaBm7DTe63KHeSrCREO3BD7w0pnLGxmuQEoBGToY59A
LhCKeTSQqCMHOcmxSzXuLeS8Iraz+ifT1PKFO9RS+KYTFeeMEZciZy4k4T8wpdZL0IrDij2gBkMe
coy2r6+kTBiUvqxHKRUX1bpArKj7iwvEcUFbKfxoeynHKv+sNZNY37CfjX22+YdwNzN4dTBWi8Je
YzCBncsn9825rGuCJJ/u7uCXO8eoiN+arThihiOnFWEO7pV6mSMbRsc+5cnTGsoNeLpwbG1N7bne
qj2y5H4AaRZMbEIqaciF2otKNLBJmfN+I6jGz6I7r9BZ4V6WjXg5Pm7u1YPNPsLI4tJaWQ6Tuzrh
nwKp42i71IuA6VU9B/9QHMljvCq1ySjHGuvUj/EgLOmq48mW9bZgLCT2kTl3pCBzU3Tgyaq5UXKz
vrRoRnA4zIOGGQlk6aJCtL6J3qldDdn25JcrtOPxfkKqItxKsNRWo78ARA/1Ls7nFk1Kxvyx/GtA
BzcY1VdZaOnbCBS+ktkWhY7xGe+5DCgN1XB1Rsa2PYKNHDZqA5yaaw6fnks+MLLvPN7DvZitHky1
WSF+hwB2RLgW6CJ53UFJQ8SEqSRjMM+/yOYAkfFR8wSK96ucWoJ6ugEsHZDf3rn39m30Gv/4qoP9
qOmNFRWtP+at2Q596H7M4Dviu/ECRfthC4A+F1lO1YFv74KCPHwlVCT0/R7iLgGueosc0GmaJKi2
FHzo8G3+vEKQbWFnzLmNpXHbf8cklX6/N7lG6qYdVuME67lZb5Mgy42i44G5EIw0zdAO0UMl8dwV
bFVTvDyv2s8WF4gCsmsqknAWf2pPM5pVWfh+14jV0gHWtgq1YYsimrQm10LH2Y3pY09VjEBOgYAd
gWwlkz5Fbor2aqwD+j1pEz9EgsEk2h2XCoRBcYKzI+T5cOXVuoYmNPyRpORIQ1gBYUFk1y4TXN+0
AlfPi1CN8pNCdcV/K1fuNForinLTVv3etbMtWItcfCKVe2reBUCJKBmh1ETXODbdv5KrRWHq1Htz
tO2bUjgdAGDt8BrZPb3HQSTcxkC+jFGZOELZuaLKLa0oo7ItDP2AtsoJG4mVHMn5bdzOXeIt152Q
bPNrUW759XojKKwZSlOlZ8FMfJ+fI5qWnbmPYph35B9/1e3qIxStFAQyFvIBPkZhSYUN9hSy9t4i
T/LOhtrAWT3SebwKu0bcYwG7Z/67+Yy0b0OecxO1RcF8afMbcJaUtVjzD3ss/LxvjqZrKuQYtENK
23TAWzvt5fu8G2kz6vi1maf8JeW9BXnSf65qp+ZlPKXhb4i2cK9Q/eZNNTgbExU1dsoUFHLCXbCz
KtXLsq6i/tiyi9nwbrh/GVbvBGqkbxqf6+vIIZDEe+a2Ut+poH0HG2TYb7LR1Sp+aGvd7cxGWD/m
G+4mAq4e7nB+b5/jwwiwVrENQ/NUZlTHLpnb+L2uvZeEdlTwqRreOdxM2xB7oauoKAEwN8wLFO5n
bYvtAYma9FI8gonudfWp7k0DrzvXAh+Eak3FE+ubfMMwxf6EF4+GdBjDtnRCIxsHjUQf1SM3+oVV
ur/UkRmE1+xJA/1JufwAmgbpv6tWC7UDtRkHPtgDLAhY/1Mx9W/hvdfrLqLCbedVWRgpNEachIj1
ZNEXKwcVXxVrWmREwG2Di+Kt5qxNvfM/DI6d4N9YfdIkxBP9JXi6fSTO9TNKXq+OCT9/TdwgPV2F
qse3q0cJKGnXOj35qsnlPiVhYkg7xurja+OG0VAlrAgDwmHJELSqLfSCHIgK1dnR07Ab1bz28e8K
uBrP0kSTA4UvnCxY1zRjLDGnm8Oq1Jxj7ZCzMldxl+gqiO8Uua6DZmyWir77DHIVYNg32IfAqRFz
PikUlYW5l9mwRiRJsCTQTojc4BeyjUwhMdKpj6t9Y1aPX2J119FOO8q80LW/CcPKSnZL7OtT525e
K255ucvWH7xxJu3UNREDbnFzsruX+pSLllZcaoszQ8Ja3KX8myaTFJboCKaQ2j3eBVzsszv6Rz3p
oepNHrLGf14IRQAwvcpZKIqfT+IOkZUOHSNmy7tfMILYeqqmbILw4gZCZskQFFO/d96c00b5CY+0
OFWn9LOXb0IIdZsNjbkb8Q4bHPosIqNMCIiCBLwXMbJFX7oSJ83rA7jgoFdOC/t6+tXfwoZYfr4W
crQL9MHtoYNTfd5WdyHFT3+OUyKds8yrr881Ztic8EUfN9lowvXmJdSVSLVXPf5ghfRfGxHxFI59
FHYFhCcYgm35pRR7SmorT+wmbN/X/4eTqbCKcIxjYgprqYfQonmKEekTcjKHpiGfKGVCyM7mz7vv
C9ZEmvliXYaYdCTHRI9uTPfVJKEL6pAsnrXW/UBbMdf7u96pjw9QZiWOYoNoBQ5XoZBoK1xKL9Ei
0BmeH7qcuwvoBnZiwNiTd5mjKu0/fK0SMTuPhdSlUGzFrIa3pXo11ilk9m8yaKREIH/XgADSXf/A
qmM1WRiXUnUFGTsoFVhNEHu5fH2chx+ESkLyNz3ePxnMmfm2efa4zdA6GuZT8wfxhNMgb/K+POn/
SLREgE7bOAjVvMjGoOx4GqH+rZB+AxGmJjcQDRlkf/tlbxLITI1iJOjV/Dp1QSffYnFQ2n8yFv9z
HbwDljFoVcXe4wWoEYlK5ScD+G0TfZT1EF9PZg6e3Y/e4E7iOAb5K6Zv6uJ+Z0uQpXJsD62qcuJe
pdHZtpSgxImLl9VZz0WVA9sviImI+GcEETd4ft0HNmwHE8rSyYiSWo3A1yBnC9fsdr5LD/VI25zc
twN4h938hysG79JBDhL7Fe20eWgnGfEJnyHJBA5JXiSLuu5UTKWVNCZTHYDioFXM+OBDTcvhTaVy
kjLB+qqcdLqBdz9VRnBiSlsVjuZmu97wc39VjUdM1r0pqriUppkq6BD6CFURWtiTg4sMsx6QRmdn
TdR5ILTHxGGrtGFqQUm/TQd+5nkoTzVdbAvjCqriXORYsxVrCQmFsjm5FteReWH5imGeKsrF1g1N
0b3oV/d7KtjEEI9xaR3LnYRp0YAreW3m9UzFLuN99YB3ZHkDFGF36Kbhg/Sv4AYeUfYWvmHbCrqc
SaPI23UZgrV5tNNrOMMejK3+VS85dTI4EEZVr3UeQJ2Qo4FzqabnhQOh/G8J3gllDyblWgBn7LoM
173LQUWnYS9R+IsYxJkixFisQvCmi+PRuVOHa2hqP+YJXoEV8Z8Xl5G9uK3Y/LtiS88o8In41GvK
sf2LmioMBhuljpAoYa2I1TGj6yuYtZgme6StgzlOOz7b+o71pAH5CkcaBS+/8Iw8+/AjuZmej5P8
AC+qTr+Jv6kztaUqdvYH+JrroyeFZnB62Jxq21hxha8L5D8X9xnak8SjIeIErI/gqw/LK56AO1jF
6EQ0+XDErOTkIlR7vRzo3WyE6w8zzslVNWUUceYWmX7aCK/JVepJMhbub2OZkKdH+9lFRl8kDWHP
D/Z2VvxNP7GzwkeUbhldke61C2mASpzL3WVdPJTiMcgcRJ4EEin39gF5U3+aOve6kqnM84RTxSDt
DMQR/D6NeQzESxKjYtATYefeHLoCUFaLmMibgMIuJ08l/gt9tHkPzXHRFzGIGsuLPRQG00C97yat
FgKjAjEKBoJgymFeSMz39nX7YzkgNr5kvEs5LKBU7Wr8t6YS7eXqouMDwqnq88EpTj2Nm3JYGdxe
IAcurL/XLEnHkmuy71DL3TRCWRsLwhXsL6HDXi5Qg1DiAXlyQy1tjVY+HUQ7ceLRogLn//40VHgC
w0HM1O3N0650n+UwxNi+J4NwDLlx7iUd4+C1zy1J29wmON+KncopYnMy9GiIRFgX+U7XKTYMZCfc
pwhDVRBfEm9Ey0+BwHpRn2qbeZwsBheymrdvAkXSdnNPs8NK2sJRAa2WmX+PChSU32qixoHJrJRF
gtcXR99NmUPLZ+x2QnD+0siUDvIeyPq2TNfiw/j63ffuX5hEK7DXqSrO6d+2AC+RlvvsV7BxLD9f
IUUUEZkyCBRW3NE/5WCzaYEW/XmybQesePlS8vC7g+2Dpri1kQGPSMkpWGmZ8eO3S4lrd5aRYp4h
QT1Bao8JU1jMEe1DYVCKCp8ZWwyt4nmqyk4F0Cm8UVQl5SClZ6pja8lhjXh/7f9ChOeELHDHzWpm
nqYfuES5uKgJoCTOsnneRJlyrD5ao+B8YQuV5cCRMLnL3obm2lr1w0poIEv1Ozq6JCPjqF/laCsH
6rg8QyIP9Zz5CO5Uq8KJ88sTfWZc4gd8ttAMp2XPauAcMbZ2+nLj9l7WK0GBPAnU09zMCupmWBFh
cS2vHNApkheBCKBvYzJL7/M8e7PkFYEoCoxBlvr6hZ4KYrihKxbemjUrmzoJobYXWdIbWXDEUKv8
fzSepuBmzaI8roZ5kkY+y3TcK5aTPkax1qMbGZBWzt7wZutlNDpg++SGXVR8jnHE8UMROnaslAB7
/+HVQtLWDk6s8BS+QwZV7BUNZvH0n2KJANhymqDeWhM/HYDrNyc341YLv4qKaPNYDXKwG19Ywxc6
FIeDeUi/5shlNy+5txzIR9GnvyAVoI7TlqpVPw8d60/WEJaMkTMLXfYf5D1XrOWHuGXS22RxsL+6
T9bvwbD7eX13FS9gDX4a7enwYQXGm2eBeLgd0zWTDLo1E9bZnfhYum+vF5fYDfD58Z3JTphzr7et
EcMGanZObsDCT6Nt34VYs7FZzcIkm6skhlqr26J9iZNL/Y0nOQenf/SP0wAw+ZterXiXfRLnbZ1Z
T/22C79NeZp6h9//Uimorh+5vzJQOhZMjNinVbtYJAWVQzQGEpylTnemWeiQtq6O4E3jhW4fdsry
GsKNHpi2yas6jRfpGyjFJUSH++CZ72cIXKhhO9k7GTCFXvzIi+v7s89NLA2RN4E14Q18L3WsVkjC
eelakr/7rIw00CpXRLJ4L9CiKiW+GqkSYvDn9Ti8nVdlOLdTCTdePkZDzqDRabSelf/TrlSq+F1/
Qkl6bXv6icmX4kNN0m7BGDtBxVRbl/sG6BtlcL90ZThohfl0JtXoOACPT/lLkBkJjczjjIOWMp/x
okhr299qPo5Vzmg+4v1V9iHxST3rotj86oeK/7HauKpXG4dBCghBIqI20UNwk+x9FTSyAGK3ocGu
TWIJoyHnEO3BKw4OCaAvM9x38MKLXvWyE7SaY1BaFhn0eW+99oEtiznsVlB9vGkwXpjaNYCBN93Q
1AUYqrRjo+ZQwTcpZHViGJiQim4/rD/Luk+I6VZJ9xAM/TM4zaQyIdg9dhLGf9ywtrT/r3INMPTf
2LTTaWu5S1S0FMEChYf+UiIIY3eZfNBRpe2EkEg3Aw+UEZkQCKTd5Y/6mgQONEcOszsRX28NLyyL
YYnUpnFvuAvGLpfcEzk0946chGcMa5pLqDQCG7iJglIwSdxXbUVzFeyQ8tA0/EPPC1qRxiPt/SnX
J1Rvp8mSKPdWG81OvWw9p/C8TFf30rf7pCPZIYVgnb9rShjX7FN5cIEvCrWW5NfnMjXKPnNoRFkf
bOuPHEQ3gsmDNmTKRE5Z6nQewriX9xsoikRILTz3c3Bu3lGmQOiX4rz8KuQdLLeVZ5zaBwU7TFxj
f4mffh9aX8di2lYxfAW2xmU1/tEQbx1E06W7JPnuo4kuYitxbzedDARKbChEp4H+fCaJzIRti6JQ
7yrmPRxWfwv9QlVtvz8oXyNE9pHUpJlcri0RiYjTCi+Uzve/b9GxlROGNwtte4Ts8k1s3o6marIz
z3d0Yx51y3Q2wAIZYYSbmup6uNCStVIjBmfUjE/IwlSTeRvcSdfiaBnKxJTZwAcIdOp3qD2YqY95
EGlK0OUjE4vFDpay5UWPBvrf89+UGA3pJBALN0++PNrlOfrZmuZV82KGep4pjzGrDvHrHM8aNQ8B
B7H+JTkaHBaraGod3dM3QN2VeT/VB0W4hJ8ERV757dePx+y77bYKqXt0JDgw9Sus/ksPv/NDu3NB
aHz7rTDkA10wWnEKMwBgU75HTtUzeV9KC7u5MRtIAu5cO9SBP3kANIyGaj+0/l1J+2W3npYdiXlO
A3aXAav1H6luVNlAPVpwazPBwnNDpku8qjHKNFgh/5RF15ir0MWJBaIBqucaj12XbcXQ1CchFEOi
jtLDLtLNGruSpCj3q/iTMswbDWHXmb/Vnp87zb2p8GxyN/oW0w6LBX7Ht1dFP+P9TSf4Itu19xIZ
EU1XULBN2Eni7p11zkglgyHMwaQ4Yz97+BKRL2kIDt59UyqoTZiyPuAGc4duIGPzFro+75ZUV0aX
iBHgsVgxUxpb8WiGkxkwPVak+1zM0mQ9YxpZAk0BIPp71MQa9VJmq3OVp6NUBErCgv6IHMn/eRmp
/3oGBp9anM3CB8Si+2uKBam+7E51RDYsMYgMV0ffar4ruZtfeCSH0/HEeTpUY1ptRQ2tjmYSYqD2
fzWsfP3OP8BAO0tQrvWsG3/qfI0r6u3eq2Gg3G7mavMl8Sb3Ln7VOLsyQeeOINstYN4hZcbuUoMQ
ubD3+fY9VK9cQFtUJGPv0Wf7ZPB+2MJN5N3LhJCTby73rbAoFx/ua0CfdxRR1Bmak8oxbTBG6cI4
gOfXShMl6kDB6kZwHg4mNM9quB0PLoiGHREye3OFnPdbE5de/UXku1jzASYvRZoH+S1NGbokwNc5
IhZXszRa6WhliMsKhKD9mRlClqRKV3+xfR66ASVEM0ET0wuAOcpFdfzntq8neeanc4D0QiE5h8mM
Wxqgiwd5O6U+4I3OF3iwpCaoG/G6wQUwGAeGYkWQK0CHju3Wv/zvQ5y6zQNzBts5eR4ndRQuAgcv
BMgMh43lAkMhDi0y/OlZ3D9YGLY3RafJ0uGTnLRugvGS3PGc1XiGElUmFKPrIm+3KaU/75MStKJp
K8DJm6xILcXgn21xIefpPb8vOxm+hwCV2BAbr2D1m/+0+RWWe0xEOp6LvemBKXcB926IuJaInYQk
CHALZFpIsAJTc8D5T89viwUoUqjSG7Q+ZAfwWWbZcUuTZjc2inJoY4tEYimfV5wq3OhOenrRs39n
r5geVoCXyTA6oOSmAgFYwIKDSOtUt38EPsjWivbCQSA50EQQGPd5k0RrTuyaxg+Obj/R9iqsIUf3
7iIbeWxVGYECDKq/JHHPYP06PGKFSI+Y8OjakwdrsMgg1CYjdNypi03z6tg/nCpPJl3jpDoXWdSw
GGCLxk1oxjUWI6eNNbUb6EH4FNCAs2WXcIIOFBanzH0p9AKHJO8RsoM0nOF+SXBQYcWkjw7dmJWa
HJKQz/qP2yue7C/Pfd7GYZYGwwvp0UL/V24ylKuZIBYkbXqmYR35XasbvQWTL4kwtFkY10GhvzVA
3FQe2MKyrg59Y4q6kGkc81+mGv7QVFPID03Wbs/p1PDmOuPmJVoLNAVLZD6AZssaCj0c4xMMGMmv
QNMrcWre+qbRs06FoRTk9GJ2gT7KnY35J9XtTJWHmprx3eHBXVA8gG2lxwndQk/2kZ5l8zlIShoH
u9SqvZ1H2iw90fL01q5TBH1K7zdUGhyRfhiJ9a2qPkAfL9dLY3VkONzQopD4p5F+6hfNSStXioZ+
3s6q+Fr6u0HPvIw2q8VZ7Nlx/EiHR/wYAKz1HUTUKXExrSkRz1C5vDxqkKzw+Ty11AdsEvpK811j
9xW/Of497Qyv/nhy2cvz6+bJhWzd1w8Ay3rPCv6LrUOtRHO2wxXfzIwCfIOaHBBZt2uHBewobRKr
XAyyD7PQ750LaRFySij+yez5MriSgijv4MEFbDnwDbH1PCq1tur6AOkPKO3g/ysaq6igoaB+tLR3
3IG/tO3dq0t7eIkTn8fcL7oHe2Ciowd8eqTXe+dpYJqtQQzP9k4k6c+rU00VJ7ceYOilI8hbuEJN
KTBtUzk16Q+HtuwlZAPnGi/EuV2jM/vJHBSN88O8C5voE/PBSkONi2AMDg4woqc5BZ8h1fIaOAIB
Nj8Gvx/db0+V7Y7blYHgIj6rBk7hrMxh7rI85TfWp7RmK3UoWgARbfDPtIGc1ZDnz6wtVzao4g79
dRCAzFe1UXlS3L64v2ZAmR9OBZi2qK9Dm2M4atpAkK6EZZpUwh0yEfH+Zh1ut3osXGbeyswbCz9Q
Ka0PqkfIO0sdB8jOn+iOB5sEIwid2vohRq/N5Pyvnstdd+HzCFr4mEBBa/f9ZRkhL5lDKCBrM6xW
Lvt1ROI+1CHNNH1j0EKNYECUbTZuMeOKO3nQowS1yfMhmyjBcBXhiIkdccPgwWG/+/OEDcBS15LB
lojQcHUTjWn9z3yZdFaUEFXoN7qCvvV2Kq9YT+bVCjOiuO3O5XsyyDstlsh/bZFHOWdq7rxpOhBu
wL/AaNiznXHwwQxBs4Sx4sT4MsR5OEWt43W+/13APQ9ZXScWzlT3UlanGD6mj4Rk1HKbaqObwL5H
wNaKUmE33+j6n6pVDD3AipAiRqU60KWlJVfETD8Y0S69qQjx9ZccW0EbElm9meFUSfyL5cSopASm
wTEeOCX0vfbvZSCs4S62tH47/DU26YbJqvwghCj8+mtWe5qUlPD7KE+EuC5xp6EOKv0EwFcqxGjU
W2WK696UXh3wN139Zu2JXNRccvZ64ZnYibtAakxbf0SJPelaW8pt+/AYCoi+uvCmZWPNqBfCxxwv
L+e8e41cEEpqA+IAVhTllrb5I7A2qECE8smaBSr49i//ffgbw0d5Tkr8tcMNmSat+AfI83JKAOqj
x2KXxFHAfxDSoGAZoMPCkPsGLXJCufsgYr1dAYzHsrzJsxze1g5GrmmubLaX7NqwnNt5E1XC5D+r
nDgWlZzlS2FrnJCXdieOXg8JeJEfRjh7kKChbIN6ZHEGiJQ1rUpyZRdY6RlMIkNCgOgwjylr3YwT
/CyAGP/AgXuGv4pQ6bNlUjaCca3ULlY1cR0awZ7PQ4De4I0+g0DAjZy47oqvyH/XnPyNs1tWcRjs
g+1UO214C4+xW2tyYygg7R0WWtGDGEDnwLVABR4lSpIcXwkDtxg8gKvkTcPTnTOz7fP+Pjumds66
uVIJ8zc5C0WSLeMBWVB6inXXpdtgS5jChbtrfCmZoMNE14vXJd20+pg2EeWv+W1ncc+nwqnr4c1+
ejJjD3oLPVTxE0XN3tQoGZuUyNVd2i6tyZJ+7PqtupMOOBpe+6LxBz4UtqXIfgqzwOGkTjcrZDUA
IQoQlLXlQsOb8aDcxrOgZwg78lKW91/DAqe2Zx17/erwMmgoJaTc4ovAREqhAGqhTBs1OJ21ESN9
N+capqEqkoJ+smlFN8ASFin+D+IY0uorC6jrEGxtHekBl3tUTefY8jDkPbFxf9jUd331OKWEoccf
BF5u/qL0jWbCqft9q9sITMOQxlOxh4Qu+FAl8DKqsBBlUsyznp5NSx2F5KB+0ch+wLaon38D6R23
1oA2CfMtAwRNZehmjf7aqdtdTaTDUS6hfJLUXuICDts6os7iklg7v0ywJOR8q12tGZPVg+N2M5PB
E7aeIGm2ReXazb4miBkEJWGU14YC8xmDMARCA6J2M8U4WWs6SSVxKahCPMcy49Cq9acqpivRvCxS
258B+ugr1Dbe+0FrcLfOFERqIaQC+Hex0LoVNFrZ0oEPkU0Hy4uiWw6XNumplHOef5Qx/SOQSBwv
obyeTeR4M+5RsnmafUufLKVvelIWcl48MkZsAKq93kScD5R2trXoAOOI9ja69/JOH+YWP222fV3d
n2f30FLCegwJYS0Hn+6Fl0/0ycMneHwbgC2tkqiWKJ6c9RPM2app9jq3+LD/Y93VRSBx8mPDJxsx
AT/Vwmt9OZDDkFDZZy+NvL1J/ccheS7SGbo8gQzmwMUQG6MwRlqi/H9IMA/PrNX/RntuhBjc344q
pofoYNMBvIT6Da0gXyGd20lH2ZTxEHnM+U+3GjNSqqKVaPix7c5TXxWvuhu4r53LwKOCmzZPSmQL
o9jQvkX04hiT6tqpMnJJky1HZTSKphrgYufNwpOhLZg+exVEiPO+asmi9IBk5uozLgPGTx7yozc9
osZ8Niw0IE6lqcLmK65uuxaWMk5uEkTlofCkUXC72FY9mxe5YspAaO7RqMinzJBVPhvnHjbQ/5+f
J20/a8WDGHFc+cdzffO2sfGBt3Gbceuf4AZJBz7amHpdj2xIxbJhX3CCwPC5usY51+GeTZo50Glg
aipfg1qeV1Olsg6JqLWzKQD77fcyFnTbd3F8fdeSJ/SEAEbxjPmFjhomPGKd23A2sv3OsKqQhLNa
kK7eQxZDQg0/OOBjxDlgnCPjgXOarmbI0QEysqs6Csg1J9KUt48pO9iLjw+/JkBT6xkqWR5BbDrX
Nvty+DmS3C7Nd5eQVmwaYvzzgTS0cpHWiXq2MEzRxaM0xDNsi7cuzMmSuBuvRNqyza5ryCrOv1qq
scxQUj1p95zrGUJalpTC80zpt891j1eGXZq2JsvJpzzXrrpqQdn8hXc7RLFWq5/R3DdHk7GQDnAc
sGdL5mcq/itJ3HncelE4xN3NzCDT999AHjYJTVRxK4cdp+tU0i0C2aT+QNTR26l+hhmY59Ic4yKA
3WPFxgOqGouRTrFgDOiW8TMWr9KtbzbA/tWV/4ZHx5TODhjeS3NOvYqtxK1uz0xeFYszzACIUsq3
wY0bNIc/FdxfFvZGDyZ/Hotqwos1L4fyFjgWxrDhBGtoBLIUMyQAENTL4jBfbR6lNoVda+xiiDor
38Yv3CFT8JDyvOOmE7UkfvXtBUzaQyXi4qo9rxk56mds762ZuuOlgxRrZfuK3OTcvrKjX0LvFRS/
QHxxd6/v7+7BbES5aKoxikJCprX9uy7+p41Wi0TS2/7pO5+TcZjxCR0BTa6vhS4l/wZTXDdolIMk
+eV9yH623PDNXP1F+HoVPq3aff09ZRpShiOlBKBS209fkRGOLIsbbSlt5u5UqquGA5ac0iIUfanw
W1dBO0p4xEiQ+vWYJzbsV24J8IQs2fFctIJolKhI0X5uPyOXs+LOlHRUtVyN9LxFXGQcdQ06MDhG
ihKCry1muM0/4YJa8b3NFICLBVBqqHzqeYbbVxSrj9cbxYUwZFF2SkBKMmv9Ndc7/OYRkJo+01NW
a34f5aqJvTQNKJ3rUBdIQck5j2Pj4w8582/a0IkV8Gv+Y+TcHVuhIozcNrFaxQhYRZh1PbvyQpG+
7Jiyv24e/CH+It2Ibp11ijtoIFSFnfnwzChpaigpi8fWDaAYmMyDISRrLC5RAQt3IjuVNgc9r0B7
dKpDPIM87Yl6uzVaO1OIPC9oo4MxywDUA4A1P2CjXP2xMlryAfbfD8WAZ2PH8P5CM6FKqmDO50y+
CSXxxxLE7e4cj3A0M69XQ4ycJkf4H0cAwUw3jd/Q0htBQZLcLohxArCbcSF7qn8taYYc/Qkl/Zdv
xxhXwSetMZnBAIDo5m5/JqL7M53Ttuk4cnApCF0bspWSVBu+Q7oqyjBaIX4NMJrnPAdy9zmMOvHw
QTO/qEKP8Gt7SB5VmgA4CU01OG/UqYRMhhSDdc4/5twKHaJB0ZrGPIAkuHdLXm6SJPsHbfXXmscE
EFvtd9wBZFGw/dbkNfpl7b02GOjeYzG5K3q2x2+DV8jw3cKP8UmlmLFEwViTR+VgWWEyCrDw7k2V
St4yEUg8qYCNnh2psp3v0wurS4El0jXOLCwpt3VFVhQ1PnKZxZRys94ofWFidFtJa+mJZ4Kj80q3
qTu2fojqG1l5V8NNBC+836I2emKPpCF68EBtq8Irp+IQfyzBWIB0h6zIbc0U1u3fVNFXN1kKea3J
Q5BrV/ctEWWFbJHoowrcM4ofEnjccaEBASYNx0ZmsThkab1T79Ls6ivWxPYQ/hFkOmr3h1H35Cjs
NT/YYq4CKXEL+D646PlvGemWLiF7YTPFvOATP3evKzrdSrjjN6R4uh1NNdkWgFtvgq6VTevkodd8
/SGOMHm1zYZDYlkdqdNQQp6Mq38+ECXRuQJWvsYB9NfBX17RWNwWd7LhkBz4PqNp1Ps0EHod7AJw
L7Bx0R7PTHmR4ldZbH2dU7VlYZ7Jk/O5swimMCciID/ELM+LL6fqu1aJ9wrbovLaAE/UdVlX+UWW
LmSgog+QHxZNrXvZjQ0FhSaFk5fIOAHUpqmW8WKnj5Ms1Vw5WgNZciFeBzLX/6TzIPEsuovJrJoL
+kzX7wbtT0NczR9RokXtrItz+w3bzgkeTZj427ifeEgtFG9JEGYfS8DhWFdbD/wzDStzZREuuhqG
8eGLZ7aZZFffEVK4wkX4oOBMDedCPBlDxunRgMA2KZ8K+xS3AOS+u8mhdrgcfR0ZZOFEO67Pb568
9QqBhrqyAY2fHSWvkFnaw37L6svxTBqMdsuZ/tKjpCsydWjpL5u+598gTNI0hWF3RNMHg98M5XHj
Voorbq+tjqdqUgLtzFxGY+d1cto2Wg4NV4DRelkLHuqmUmW7LIaK9Wk630XILmG3VJzuMrcP7hg0
aFJJmVvl0EU4oV5h4DdoCNV1rouv37kq7gkHO2Kq8IZkJtILp6zjq5UXfv+cVwpKZ7QSgJvMdkZF
A2gaiZJUiPvOuF2hx5ztkkZfx6Zu98sccqwcCIndStpctmA519HkijE2jt12f1/USaqIxbQsq46L
50lSvUmlBPykQ/M46jeIWywHINtE7hnL9IMg1w61DjSuM20OomS64gOgA1ZVk91MuohmHPODwkSo
o/B9ucBLIL6bC6YnoPL2oVA2prmF47YrFoct+nALX6xZn81gfweMAaerWuV8sADUKYLHR8Q0T4gJ
H8V8MlC6prgS9OVo6VUJqX6qbI7+aqzgig9gJayuWuKI4gRQLJmHxK9efdPevvxtPs5FRojYlY+5
yD4t/nW7YYN+Z3pU/BMg00RNyAqd4Wpdtze195VAOn/FZAAsUAgYOSxGI0FGqzl13DlSN/7ICr8F
I4/znaPQx7Wk+Bq3+XP2ECHW/5Iv39v8hkkhwtjmNRKwcAeflLs9pHSldriy05Zr6SXqgSz1hQR4
+5MzuqdJoxJ6DiQDOEG2V+fFGQ4N6AJez7Hicpc4nit6DHLPHT+BQ/JkMICr3GX9XFQ887UHOyTf
KqdzCiqRvCwNehnlwIXCQKzFAdY6lIaIJ9Cc+VFun223amAJ3Yj8s21oubgwfBkTORzwIn1TP5c6
46qZdi+PyLdkXZV3/TOU6IweiotCy7bWOfYhqjolVmuD/5lFztfFuue9/Hd/FkntyhHJ1Ik9kpL0
L1R3gVGHUEhGotAXytlG1yTmh+bnYVA4+frS9DW8nf6QE7TnkPEc7E9ldR/G3h3R96wyMkMHXegF
XVyUDgwZ0SrVR0Ncve5W29hZ4od1No6Rc/LgFB0IT54RUTNT0T7oMP8FLXr9Mi2Itx4leX8Rv8hR
tkLrS12UbOhBjPcig1v2xTKoFgCK7VMQ0ajxTT95IN7I/l4MS5xvKjydYJa8Nw+FXe6ir6GDF1J4
Fv5QbQNKjatdAevvWgRHY3dcsMBFdOePWU2jTMoe5htMewN8yR2zg8/tHWstYQhDNcCXXHYNWZIN
ocA4YCZAruMbj5SR2nqVQdnoV2OsnlSwE/EOvIPJcrwYuh/p6LmgFXkwSP4h/kNDqP4KRynbNafD
60MG0nXsyXXZqPULsZ/Hj3Nwk9/x2/T2UtJ3Zoh/XTUBX3FphOvXnDKvve0AyjVxEFCsqDPCCC4h
FPYxnejmHVsTaXRHQR3GuqDBvQ+2b14+SfMR/0MtiJIABlow+WsWyYIFRfzbjlGwl7RaPFMLtLle
Mpv9f5zC2eM21YFT0KwoxtpG3IO3qZAu+/xsKPio0PukLXCbVo/kzfP0uUTnJMAAUR1V14e3oeOC
+hgfkny9hlYjvRgDLWgkExWTtt4HvByQo3BSGeXBcyKJxxYUKRn/rRELgjXAdp4TuLdBSvj5deh+
JLWhnNqpxmCdoMjvVGbuvw/78ca+ccJoLcUN+Zcndd+etJGb+Q7HduqBZtbzJLko6jWPhgZI+YXP
ssGEX9Q2RWJ3MQCWcG6wEE04bAyRGY07R7J81SMzK5CGoyuqkH3MK2bjtMaXNeokEAL/HQMyRf0V
rSw87ENjRUNaLUIxh/aZKQuBhm+oaIU/BitOtKicKbl2riKXmRQVABiLczW2FL3LbfS/TPhULWx8
OFUTa9IfuY022043EsvgvcW+HlNDCMc2c0BwG2cbnVPKO3DQW5C+sgYhokIwW6pvSefC1H9dyZo8
qA7EloudbbwjWGy+i7ZOnK0frqi4UnRSyBDCA5m7B/VsPOTCB9ANnMrs63oC+AcvJhp2t2ZMgiZq
bD8Y7+N0bVBH2tPLSTzhiw2s8kNBzV3XLv4Id6mLIT20/kU7W8RaFYJDrvMwzAtLeCprOAfSOnxM
7G2jEmIIv4hE+uzyIxyIpbIQBHyoyOgZ1UW0VjgKM36bO7TKbYk54GRB/AKn6FmgtoASimItTqAi
bVZDriS4FAp0RrqDPn5SlbwFcDK7xV+9RcX/CwGTK1z1t8nAhF7nkMR91JJMRIPrBa64hJUBSifH
M0igB/LaCFl5nKOGkAvNOkYc0+JyuonQOXXZ4sb2CDQZivbbWa+AVnqodRzd0DOoAEER+boLfwb4
zfk8fvxR3l3pUBJnzN0oUiBGLD6W85AVwrpXPHqOZgqrzvaL4JdhoIN5f3JEAUjDZtWBERHQMF6i
4dGadJQ9g60w7ASHFCbmtjTUu022yvKFd1Tpv+b8qJGHRqY32Xe/JyGOHp7XaE9xnaR53Vko6IZz
dxfk526Yj1POkA/j7/tNpoJJfxq4SMn9TI63uJ7wpZxG60EM1+dJ664gDD/EccMt1FlEiBNtrngV
nKowdYjLHbTbLHjB0sy19qasZju5R5IbF8nxTzNMBBoBDepq5W8r93BRzsLtradMY4tRuzNkBWKW
x1TiaxeCFQX4WHO6YeNcwkmOL7N0sk2EjMqe/ZW+EI+SIJqIGqtU2liAtrJP6NVkCxF1RL+so5Rc
IDCMDOFYWo+7zMxaiCxx8ZA+PZX7WrFfn7Q8AoIDq5wLSq+UpsqolfoDaGXClAu3aOIJsas6wAsO
XnZnlqSVg20lxz3H51x9sT5dJoJfoCmoGFu63dLCRltiK0gQ5zgM8MWH1BbPGIOcz9xmD2ewn7/j
GPHnTdk1kdMHHgXgj/wwdQfFhgw9NsEosi5th8p4ShGhvEbrBXBu059VyWIXrLq3DR9fUEQTjnHV
VXtk0edKMo7OhKDklU08OurApvyjMAfCu6h5kMJP8Pz2Cmh5woABgFLR/ovOo/M4k3ELXZmBjb7E
DTQDYhvduCjNwsC3ZS1c2D5I0jR6mqqvaciYGrgk8H2OHOqrT16WTFUD/3EpX7hk5ihb1vw2mut0
NaVV5k49K2WvX98BwMB1cA+IfajMNWKxCKUJFObO8SkO5C33PZnfPjYwbLJ2Lhu2ZTK4HSdzhGbv
kr340F/bvIAOYtZaXeUS9+SG7o01KVQA/Ha9j/xByu1zHhBGGlnmUeBqgDl+d5EMbFqCeuoccBFC
P28GF3TdZenDkumyi5tGBDiCCyhhEg/c/rbhWQ6wrv+Eho/C5rf1bq6tBdGms8llQZV65e7mYa2V
dTZbiwF4s17i1gkZSvhZobVwO0AeYIAKNbg0H+2uxStjWMTqE90OjIG2dCxxbaX3z57ds/v9hUFw
eMD8BC/YddjlR5jTWPEeOonqHI2QpOz7MVX77E/LVae0a+PrwzAusdaPz7GeWh42ffDcs0rZ23fC
Q7ojdUzk+RnsjUlTHv8nlrwmu5hg3+ct2rAjyhZu2GRjdR+ON16anxTiaZ8VbjAfUS+EibQcdpWU
+ZE0iyPnduy87QVfefWbDTXZz+8ygiHr3Hf0tQJaNNfdvQbCi6O2wSS8ejtD2sQ1KAK9Vvns34w2
VP0n46yViOrE4sAM7Sv6x1IADXPnVsCQMn9VPFofIhhfaByWfEkOmSlQiaTzbfyR9guvKgAJwg4B
I31LktVQU+NhcWX5ckFG5ggw+1jelay4oHOEuFRSPkFezsLVyTLV1Wd96YrRlp8SxCCQVzO4g5sL
U+MPdMFkiNa1odDEnrX1ukjGY40qyxo+GN/Rb4hyr3Addy3acXd7pJyTkxvOlpuXNVoChYwzsZa4
3B/Cg9iw3bcEjFubvRE1V6DeiK3Uo1qxGUCgJ0xkGoGrCBt0pBqFCBKU0wTDFH8o3of0vdq6ycsv
TRA++fnizD9D0fFeafM94TEZtf7mt1uAfhqEJ4FaEhf+D+tt0Wm9gIZMyHw7qdJrunstrvfH3vtI
GqNsg4Sur8rzvuKyaVxLi/0yXmXAQWkuXI+wiANZ3vgnRc0/vSn0PATIQ67AdjWwN0wPC0VqzFM7
Y0Ho7K8W5ALZ+Km0uGI0S0YL5NJH8fWKBfYCekklLebkxSyPCM7gf+8FdfRZ2C69oui69Q8+Yq9P
LndjcJyNm63SMkKqLwaX6Azi3lFn/eCakDa8kTjKPodQvv1xaocFe8cX8xcOw54aV9zfFtGvsBbP
Fzlu/VLzE/GBwkho6Co882MW1e8kTy8k2vJBWIFhwZeDglUhgWWIA3MKrTx6YOjc0+xFZQOupXAC
uE8o2XVlFv2XoMlTfZLtRwWpCbf7dkj8NxL5wt1PqoyUbrMkP83/RzTzBiyYmEqjpqduWHv3pqjn
XdUUXxxZRtZDhWkqsPSIktADYCHDdWeRABDBizA7j1pS3CtqsfS//g89l3mI1aMEv1gJsiHEI6y8
exFMFn4uiLu2xw/dtc2fXCq0/Azt/SPKB52UrEx/CU/ZbhkCIc92Goz3D9/Ju7ADzwbHOe/0LYAP
s6tGdXNCwEZJeyEtXtPcmXWP6iio3aIZGAAei8E5Avmy7eTFToZIZFRyjwf4gAE+4PFqpMo6Lmni
ZgpKO2Ks3Kk+rcGAz8SRbyuAPtaWkGwDMMwNt1Jh92FRM8ld4Qqv1vzWiGp5YWKkoMC24n3YZv0Z
EwWexvoZwR1QRmnS1Z2CxZFGhHiwFuC5ZZyHbtOptQuxfxUwKJibySl2vtOSOySfMhqFxhruvET8
wGdOC6i6Z9OCt0bbfsZLdOl9Rp9j4CmagiegBdDqvrQ/ky5y4Efm49r70hfc04XLft+Ar/ToaXR9
5Muf8xod34BWdEoqziwuBVBstmn/7AK+j4iKzweOsX1bH9nwAb/db82RWCnyR6wAywDHYVKEwW1h
sYd0EgvAojUbpYXjSa1Ehh9unXaL669YucgVAtog98jEsbzQw41ZQM9UYbTJ4YyeeYOv967hxb0R
oUAW+lPX7FhbPq+epUoKOiPJ+MidpKgFOmHbqJeNGOZTIkW9gVdEg4vN7MHV6eiO3iiHQxzCp1Sf
Ajq7HXyxWeqLQijJTvO6rhyokub7lM5g8KAcILm4NyR/+mZsp0CMPOndH+6unlIxVEtAmA0hNNjE
XW8sbALwX3Wo+T1GuPjscR4hfw0Rj9llwSu8F1o0avljIbxcj7sHn9CNfRngqphh5xtW+UOqo7Hc
a24N7syxM0U2Py5ZSyAYhaRVRPZqUqtrSdD0JW+2hxv9zo1B7iv1L1rl7bZeKKnCShaSpQR4rQYt
uggYlIp+3ksLKp8zUZpjDtHyBUZBah+gYKAD9f4WKx/gPgCHH1lzWWlRto4HK1PLApEXI13s+Pct
ANGTi/GhnlbSAGdF7jLw8gUXfUme0Qd3Upe3AYTBXpvSZFsd0Wa41RtoTwB6vV1qNZCIgPg4BiVZ
p5Ob7wQT+nRlm43FjIzKUsCEbF3lGetyZa0rPWe9WayAHHbMh9Ns5ANM2KjO60NeuSHSs8slkm96
0O3urlLGvb1duEjYcAAUZZ3YSdZFsKbjRpo4TYkJLpjuqtylk+b/xlackUDEFE6fJ2x5Vq+LBNoT
597dwEuoC9+yP2Rb038tuMIpixDJM7q0IseP3jBomwMg7DNwjc9MQJ+HlirqjrF+sKnZsss0w4DF
St8UNb2kqEDRTp5GD8dr4u1ymIVlU9DltiSzwecWggxkG6LMmN60wzpD8gElfq2JUjyJRodpaSIR
S7+tLCPd/kmqBdmxeNYOpu4CH8uzl4Y01vjzM9BRBQQL3jOF7LV0Ssg2WkrlJUSGhrDgNLlg9fSl
icZxwCbjyj/GgyLAiina66C0cLn7naGN/YtWc1eCX1oDqbBdbvQOy1pKzRxN9yI6tU7b/VOiQLkE
s6722Nq4X+P+xPENRypdj/Z8BAYtTAY2JfDT/DY28H5+NgoW7EgfhwO3bEV43qrv6S6W2iVC2Wxo
zMB4LaUibPpv6z41TaXeVkBHKNddyScgUHXS3dUVavKSmwAdsDMJca3cL/bjtx5WeIwHF4NUt3gC
cdeCKtWOSxXN06tcsdKXGxjiezDZSiYztgV1iBZ6Hqu3zZxRrBX6axlOcbsgQFbBOPYVAZ77YDhX
gEgMM+oRyjxVDwfMTnsdknCXZGd1wNp2yFdzbCqQ0DYM0Sy0meGhVbeutWBspYU207S3ef+WBz70
jAylwnWC1bYr7KD/SV47YOWwS1+7XVtvsSTcC3rYtpGPNFdht85PvymA9EU24POc3j2pUhLa++sH
Y3XG1585USo9QvqN+fpR554OQBa663TzMdi4QO6j7R7o6i2jsPCJBwA6BxyACwVXBOA66FyyNcCf
KY29iH+V1Y/HM/HaNWBhHig4iXbgLyhzflQAciuOUYugUXDZ6yEKH/sSi/EukivxJjlWKQ/tg7Dh
upCvnbFRkZIDhN4DWFWxW9MQH9ItL3DaBPW4NlRI/yfeIROYCtw/8/z5Yfow1DySsZMscOLsqRIy
vkac0nsrurD4sAqPRGe6e/OzoSu+J/d6aFVL6cYZdPE86MzVBNECIh0gSDDNk1UtmHahti9hFcr1
jQ1pcttUFIPJF67iOWMbHb4XbkXz58FnyXe17SCld4n2FTKT5TMzEBODMGiMxsOLtOsy7Ga+xLCm
MU2zv0etBWFx12Ryp6vGJg7xdW2pm8oTCJTD22Uz8EuGocLBLIn1/RTq4uvAwVPXC2ANuPdM8i8Q
qM9DGWzuV040ZJthW7sY2dSCdrUYhsHqxVEgPqMPJq2HkbDpYp7L5S+xDLADN2RUbB901D/EiqQr
1gGN2Znv+k+TS3WBpJsnnaZCJfX/JmFGv5cnZeC9Q2b1vdYoBf8mIhnL0oAROJDSEYteTPXb995q
dR9HwM92E+A0Tlo7I+1xX05MKT549P1djLXAWzerLuL2G243UQecFuLhBVzquNpTRtTVdwYdrh74
1S0U8C3HSdoHvp+29nphRFCFd5gkYX9h3+QPePqvcctLSNKcpHp7yxi+Zj/VXVQxUldTC6ASjXup
YVnZjazclDfVek7JNq2AGGlY17zivCtfUlRkoBGHyr/ngSNscR+hhAgXfsyMYK2VmwJMy4l8Ojib
gKJy/JXmcHNYtT9iW5oNI2cRxOjABGHpECwdjU2w5y/tDMpt/orXv7FWGEuXR9sFDsp22UX1+7+j
lX7rr+beucVxOEpXhmQeJ4Yv/X5AEL9edxw27z7mOje7dHeLxTz9fpOHGSp5MzSCcPqlRZ3uR598
/HiEtUGT6Ag17ATCZvfBLB6iXCn1vma2+USXOEFw3g7rOPbc96MvQiRjNfL+a1E3Jema2tu1Bm6J
fQFNv5mfl4pgvGM9YpsLYCpLNqVpkIMvExPXR3GvlNBKYp/+s6/3b4YKMsm5fZzawppOKKYVn0n+
0XKjwZTgI2GPwFVbkNOobF9tLWu6DhMY3V+ttA4JKuGjAMo7phmYKknLa1OjVMrDVkuZceAvN6kx
xC/9tCDoxWkgMKfLVjFnCpMMde6u7ggXbqTJlJQoBdIH5qE0uVp+gBHZofJaxVgkrEMGieWVH3lt
8hqBdHDMBuzCa42/D24IMY1S+MelyN+SPHiMhIlXBA5hNI7hmdFQnbRlQs3wh3rB0Ss5lh+PIoLF
w+F3b9MuQL3dnXkuxFUfyzLl2gP1tURMLL2Bl08BJvfyuUlJIFzyYc+d5Cec0ApiMrinizeHMfde
Vt5xoMBYq6qZkbqXikwx5C1NvL0M6l+yc/+RI3XpSaZyku8ln1PLZsl4V92oHZ3a66kWJPvwCOCQ
cCteDI4YJV0C161aOH7hIs2sfDk3GXoBS2h2eaDXbDpondXFvvjS2oOgsQOfQkXwKCnqzOvGSGNs
n1hrZGQaOv9yfxnJ4IMx5YXzbNj9fG5P9qqKe7vRJm+jjY/HwgDvlmi3WLeQ2UtdWeQSEPOkDFLi
0R3Yg0RysVmnvQNG7wKXsUrQ5gKaTmrcwmERXfYvJrn9HStGKmXpniTlF/sPJlas+60qGlBIRLXe
abS5TM1skW4sXqrbn1Wxdao8dUCj+34q9PTzW1hNKcAUlpJM+9jX+E9JjFyT9pgww6AjTS60PJzR
of0PUYOxI+T/cX1+QzAtMBuzg1tmQal1N0dsDVbI5kosUbYfWzuo+1Gs1WJ1cu+OR8y5+y4+p6TF
pATDxtmM4CxJ39GG/iP1tZ/5YtCAxJHlwwXGjFiFbLFwfAAR6/scau0+QqNv7xDDlUN2gkR9Dzs4
IIwi00bao0Q3dyLqg21yGYGW5hhk75xwKOMEw6qOPe9duuH45TbkarmB0uVYZy/GZUwzbjSGoCZy
+T+lh7pLF2WoVeKCoUjA6BL9iSPt5iOYXg84EM4jQKE5jjz2R6d/UopvwCMAi6ff8eqDoyTrggKV
xTIF18wHiP4ET2QD26wGLXwoy3NChRDQT+x+doK2TTHi3UHyz784QOyoAJWlCnUTjWtvKkBNjibq
1XXOvLybc+Ax876220ntLQUgatJwZcn72PtUw6P+CO9JeU7ALXNcXN8ofAe76/x9IGz130eCmO3E
/o0Bu75VXd8T/H4Bk3ADBYNjk1vGbAyqAst1dWLVDi7nMSG+V0Dy26Om/RlV4EvWYa/Y8novQ0JW
YK228L/pzNLVsgl5aFwFE8R+krcyDnQTqF6QfmL07G9qrrX7kf12EHzJ/5el0iyvAS4z+uUhNamI
0bZRPsBZ4ZKXOSBPQxbclAfgdqDwg0kbv+J46ixDXHGJb8cFyj312hvcWUneU9UY8o39X77PMgbS
Rsmx+VAi8Nkg6b1QMtyBbICRmbpDbuuei0468QUn/AJeJGPtAnFUM+jLRbmnzAypgmxKiJVcyFcT
QAkeTg+u8SivqjvNdyY3to9S7CVJadaNZmpnReXOmMTikiLUiL8PuN8p/1aZM71kS/2nXrfLnPqN
V4l8Z/y9cr5IQqVn3xNXIocHak0lZGU50VDcq4+N5sdtkpzfBVCOANNdD5gpsRuVRdmOA1/CoSIs
dbI3/Bqi1m8B8MWpKMUEvkKtkkJEPY4KKLajIj2zl+WoaS3d6aXNb1I/JaR8OZYymg5i9TSuZbX6
5ghXaryXkblOFfggEw2StuFv/VB1nPknDtUEyDYw/c5NBtSGXqKVcvyV7GiLPlHSPdQFHKmrdtoe
JfG9LfXWHr/RhuvPS44ohXWwfObWptfWMj3WdAM2VnE5IDWar8SR0t4lbSFVHEevHLNZmPmztk99
Jmibao+WFIPDYH36cfoygZ2yXLT0JDmBhYKGgPXr756hs2pnosNd+Jzrl3EmYKVAaKpwFYV217bH
GMRBmvusAbuX0Zrids4kXAdwTfqu86JyIUIxcH1d56/9diBJCqm2hk1pkC4P7VzeC8v/fzbSD9X/
ou4aY17+VwteTEo7kMI7oDivbM3KsC9DnrN7oaJxvC4IJ67BAdN8d8Hm08EMPru2MYIcE2dS6l/l
xMjxaS6DTcok8+vu0jDVPSWMuGhc3N11TKqmM1+/8zUEdh37v008GvXJASnJqi2/1Ybm8c5TjoM+
SO4Yu0t/4Ph237Ls5amX/822NJYaTq5iJO+TWXKFdC51Y6vi7KJiiYS3UkgRUPKQm5Wb3edCN0E/
NcMC1LpMo3iFuKHZPFZTiz3rUZhRhxx5d5ZT6YlRu6n/ITuKE5LtHywdnAT8ToxqdnULo1TcHIKQ
KqbcC0eepJzfrOMrtCHlmpI5miqcVyfwrYbehTtainS7DV9kcikNQRk1DzCqb+EOJxUnGWcwYlhu
97KNsOs1f8TvQPoWw4bOg4TViqKEMR4cxFGMldp3WTZKz40uwJYOHgz6pWljYLcmvwpwezclruod
cj0jOUIwk615UwgP7V0HhKi/B9U8ujMXYPkotcDdVbG5vRtBe3NB3ult/Df8RkBCg/tBqso9qRX9
ACHHp3PZjlMbCiecKyGi7urMbrzXV2kRMvle+lF+pgxHfolQQoZH5U3PADwxWYEQnPziARyQHP1D
j1V0Wu1zdtdDt6+Tw14+kMKvC6F64hXdReX5UZmHNe5ladalxx/VlYQZCH05ShwOHg1cbJpy/fxn
lMiPwyYaTfnLyo/X8I62krIOkul50fJ5wnpsqTXMipmeN8PMzYkzZQL18TSCPNaVsuQYcbDJn6Gq
zBlgcsFn4XYlCVV9z0BnehBe3QArNO5qutnCYWD3Nx699ZRI32SD/baLOXkc+LLu2aM6GhRo6lVf
S1wfGW5BWrODbnAlIwLC5VbajWTmO5WNDr0ued4fVJaXE6pBv23gu0E0Zf4+qD8tzcLjSaZd9KyG
nJ2mb44rHS/uCs+dnY4nsd1ohfhVmWlZiQtxFo1QyCByTZrjtXLt5qxIWintWRWFzn2dcK6NmEfR
zIZaoq7hTfvHHiBbttv9cZKPzmZt4y10kUQ6zupzPaldIJu57YN75ajiNq8UIAncQx3hm23+jJ+r
cxRzwRQaxlZJ0BokszTbkEySHpU3YYDG5oClkmCBCQGVWbWnjlYWYYvsUDD6vTG7ZNmCX3atIiAr
GJt2VIEAXzDrEftBFcbMlHAVgLOP06nMIeQaj3EzMCf3EdvigHHT8EOrF0gtm/TPQ7HfyoWrbuB6
Rx7W83gnW7bZMdEPb90FpsBs5hSggxD/AsgzOTa27Jav2NQigWfnUUC+XJv16pMV7+qXS1cBM2lN
9WkgPKw9sxZuGJSHto5bTkkkNlWznAKupGi+dbIsDkHn2vdb0hYE83yKHpTQXT7Dx6BJh1dTGZXr
xFfZq/UoBHD3VD5etmlzD/muL3yespdt1vzKrRmW8Qe3QTvgKhSuW35RiqUVTzETqCRbgjnTcUxq
2PWMOCvWd9q1hrzG9QX4eTDPlpzjzA2+Jwg5QR7TEl6dcWuQJo0dHYmYXfe7rbmzdld8siNq5UL9
bzeFHKE5fj7ZQkhzWU45wraIOJ97tMHLFJtlY3TI8uSkeuV1pdJlbLzQZxuFhWUWb5TbAkTDqA+F
J8hhtCD/X3sd2KrA95wqjn++s8fSPOex8QR2D2lNf09/B4jtnyM+3mNcnnz7OPu07pJqty3Is/Sd
ITqr4BYTeV1v2sIaoZ5jMsIWw+2LgzC3DwNTqJnwinXeNmsFo5tdGgST0bLA6nXSm1AEbQ1rEiIB
0KvK+l1ntoRkHfLGAh5KitPXowg9du4kfyiog5RJhDhIlR7G5cqO5Zq8YOa2RvYNx0riTV+wwuHA
wmnT92gkK8bcKjAxDsLXMRnWzumhbTfZ6V9hGeua6tk5tRv22ZUF8Y22bPpp5xfPPMy95cF9Torc
sm7cxvP8GRGav1FgwUilCO2MnofEEHksmoDnER98acV+bZpmaD6333HQAlWBTj5iXDV7PcI1aGkv
2zHDB1QMYGXMvEehUuDYLRAZUxP+H3tdoLK8cQaP/ZO2u+H7ygtIBkR/SOSgDdneh0l99GSKLLRr
6M+qXKCzsk9A7NC1ufau7avxesgID89qRdnyKKY9VI9/TviMU+Lw0Bi/004IB/ipiaaR+0pxC+CJ
N4iGZbL5hNONZp/dgNFf5i+CRkXM0A9cf8HE9QwJDlhoq6/jH6fzlsxuxIsQ99BRZQVsxaaYs2nL
mqfYyVyu0IrPCrFP7NVIrbOpPsWnIABPKBMcMUlAPV06AiCB8pxwNPosJESzmOOJPOb28LDNYjrJ
8Mbrq7IyaxKeXHUhhLw5UIxWqud4cqGVP2fh614PtpmDi3E5FGqfeMks0L1z+BAHowOSvBjghxqL
JPAYn6khrh+16I2CU/pF42bgMHB3GiFiNBNQUafYYLsd0RNp4ZmVKFvcEj9Qrsw4ceqQYRjtuNFo
LDvpZ1mJ4aYkNuWj6H82CsHZvILfSZ52hg6yEetArvor+bBZWVSab9vzmS1bgaT8r9rrcX3GXxrq
7H4bzdCHLR/egpqhlfiwjMdIU+4UUEMOHkvCH19gJduucZv6MxqXWhedFIx+YX8CH7r4e63zsGLk
1y+gfl23cGzZ7UK4aZDDdGwWB30wi5xDwEaBhleWg9wYku8M3awRt6wCFOyyiXOrZdKvSmG+SPZB
vlJBue3EUNWPDjgZMqmXG7yAbTB0KiREJk+IX+ZxVwPa4c3vLYbkWg48nMLzuiA8gjEjOukwQWBQ
HlLYhDf6CuYLcxmc3KGHIdLk0IPs9ZikDqwkwx1nX270SlSJ9bnt8rn7VZTy7CaAuZnAODPqOm6X
uVx5GJpf/rt/zeegXwDQAeQT8SX6W5GXghCDH3jFngLS3Bw1uy83zljni6Xrnlgt5FJMT67AIBy7
Dxtis1wPbN1LUzcrZ+eGq46F0iLDUm2ojNMcw3oWPmcV7EnszoO+lyvM/4bQK40hlc9UhjLTK9UM
bvXSeAFra8ZwEojfKq9DnIyuztiZaexcSU+5oHSuOGAzH4zOcLK2Tg+wEDGLVg4ujRfFx10dCeJl
FkNmFE9seWwB4fihGUD/HAR/6nlfqey5kusxD+eTScRxKggEcxsRIuAn15NXxTr9BLCQ6aDHuaCU
3ZxeDQbMqGzG9bmU/KLl37z3VCcUO79jEbr0CkijbesB3QwxzFHsHVUCyPKfSdBwxTytiO0xde5h
sf55hSKsClbqlpop64nIVDw1+cafRmmxDgSM+nuidW9RwWLTBPIkTIJM6KqYKUenxgobCwGu+bqN
iFW1oym/Jvefvid2iYiD5UxjLgPr2VcNY/st5CmECyftSVk3Gh3yicIqrYdFdG4wIL2lgeQhbwNN
B5Cmb4onJ7JGXmFr5nebXLv/XOJSx8PT48S97CEkLuJLDGZgZwotDw24P4L7Zz9UvxxK8PqtwvXw
wfkaMq8u28NML54XrxZY9PaDvC5z+d3JuTd0a6axlA5Ruk+H9H/s09Xn7IV1/S68bfgV8SMRtfFA
1kiuQGubXBl7Rc9XJMGlBrn0938S/LVer3jfcNbjlDWeiy+uwf4TDJoqRjg0meveZCxP17LDhFBQ
NLM4GSsHTb6s+7JBDQvrZ+pgGsusaooHbW3KtBdX8LeJBFe/pkzM07mlA3A6M/JqiYQCY7hre/vT
r0wsEeh2fOdyf+4Mn204YVx69QDL6IjgaNWa32bIMzP0nQgkxQBhxMtlxFQIw7qPXVVVxi/BCA8r
Z5qoK+FZ9ZrcZ72Ir59qze12G45QAFO88BS52LB8imi2OdxDU+4AVvGqeqOYHMR2pMtzc6h9tvh9
TcN5UOsP1ffYIZv9PbqQJuMXkz+pyEDpKCj7vD/r5wdZ+IE+Th4uNL1DP2s9fWQuu73BEeQ8TNGv
gsOUDk0bxE3bZq4wkfd1IlXE7qjRw6phNsHXti1WLNlqMz/fGmHlqIQTZ/gOmLSru0Uppa4vOdRb
AvCFUAuePW8zVPP1E+gMMF8NXUC2FSqCTx/tXp5wDxxPYMm0qzGCcnT4Jt/mVXEPccc06SKfnwh0
UOMEaQ/NAJC85fNJxFgUebsaNy2qCj+YTAGFwm/mQXKndR4WKsPZtQbr5CZZIqF/H1t1cqRqx8KI
2P9MWV4fnjGNxd4gN7MDhPSFV90/Qx1KiqO7BVC/C+FpOz7IalXa0dtQP0q9M2RQzXYVGDCa46SD
NehWOdFQtYjWKBs9DFVTweUDCi/H2CRaqcWmbQRfkXxTBRrsVqLry77GRrHDYZJ8+kpELZ5oby1b
ww82gJRMcJ3BxL02IJTAGTRkzj5SVJ3lEWu/Hz3UfjdKZt5SBtWeCg8UUT4h7zk4KXuA+zmOfnNa
Sg5iTaZguncLxAJZqUe3QmhbBL/5O6ywpKmy6IHUl33ZUaNjGgGHpr0Gr0x20fa+zU4p+NJsAIHo
d1H/lMSyN4zlGVb6IKwsqcrZQ485yDxFKt3oQZX4HiFSzTNHLF3dxHw4P/kvqvSk83tH4E/jC+/N
aedI5veRZYMp0I1WQs/KLgeNla0CUcnWq+BZQnjgEKvISXzMh0zHYXs4NptBSPt0zoSF41KHPGul
BqEryw5Bhc0mb98MDPMN/Trja9OIFkPkL1y0fSfTRwTFtZes7axYpD5us0c5pD5OmrwlHdXST3fD
cGrcFOYVnHglTleUVq23NEe/IzSUt752+bmFsAO3xRZ8nwxGtveM04UDo37g8KmRPu7u97qRxOpS
f8VREoQC4vUpn57myOzeWnc0jVG/VFtj59QWFNGqEz1OW8hN0mPtBLYk8vY5cKTgTig60Ca5D1VE
Hax9Jp764fcKA0Ck2UWc9RFjkqJdCqzHr67CodeLm7NW08lZo3ucb5/9jZUvji+mk/T+2exikQeW
uzUPgROMmVqbk00FOPGB+CmHNQ4CdUQ5al5SnM7yfnZ7WrpvJDbTDMzUkW66ljrmKGxHLXbpNDUX
i40axgoNA8jtn0JmTPIiP54rgy+Duob3oRRxNy+0Vf8ePqW8WGdbYAhyJ7Yb2O/hqhTC4tqbzdL/
cnGyOAY3HqdjgG9grG+kdu66e3Jm55ERmwu9x3clBFNrTH+bNyuG4GzyfwHRRnmeX/98aT76qsFW
/q1yLR915DUeZ5+3T8I06dhDl70u4QtgiWHTJJEUHM+rZ9eIwATgRs1jXA7QHdD1rEtG9skcCWIi
xGsC20TP5bru/GNLpgRZ2/3n43b6vR+CAt/OKa5waVheSPUJJ0Xx3O7DT7xASwniWMoIQo2i4z2P
VxYObbf1qG1BOEs5ENQrpkk0zErqj3vIgk1lnwQoXWWCvM/0r4nPFFP5aMv9vL5nRhphe5u3qA1a
iorGN0QyrdaweUq2kA0rj5hM3IznCyzK1MXHIy8eJ0paBMzYTziX4z6v9ofaDjtxm38Rdsf0fpn/
OQpFoDh029B1A+Rm8iqFyLGOEI2tG72Dvc//U4+J2nM592bfjzil00rRAvmTRF7eVkOgK9VefqmV
mDFZ+VUNlC7EJHHKFe2uWGefsNVCNr+4keRh01z3Q2T/WcqDl/vk2YKtxzzY00GpaHCluXF2yMx7
rS9AgaCWAW1vYQIwaqaWteGygP/8MUOLX463Po8eDTFmhl7DAs7jIhgI6a+rj1BZQ0SD7ezUty9D
Igq4JXaQqG55NMuaAFO0klCg+LlTCT2isQrWcEkapKyKL1gbxHjhWmO3QZi+NaAj/+e3pK+ovKix
6d6r/wKrRGA49mI2rG7r7Z3W2L7rsZysrFCEqediFeJUYj7rqNsXAa2CWaTEajX1Bb+fePoPp6/Q
hE53hd9o+rrrkUKx2dv0n1qbfp2dEITDWMOrA/79Fib5shliZfH3rvAiHF5jrrGVdq4kfsctY0Ps
4tFu3bGn6epUjrYfz/QTIgpZ7DjQi/07J+4aR82KTwc7S7hVqEMlK9EGE2s4TyzG9JdKadTS/nIm
Khj0cj4T7NvJm3OSPF5vWduCTS+LB3E13x2tzGrr+8FK7ibv1MkGHLrmL767pEth+3mAr8iB2Ufn
68PjuHD3Lu6RK3LTKElS8cf1+3Pw4vfKOGfyzT7jekwP/b16cEPdTaHJ41WCsi5UdEJk6l/td8ty
2f2xpiO0/WUSBeoh4oWTIIKF/6U3Dw4QWxJrZljpQHqI8RbKQz5+snDkwKs6osNiT0TXANb/ttGr
CC+E0SWrzEEj/BfxM1Zv8l7KHD4RuenIzljLBn1izLKXRrOoIEbnmhPJaIJ8OupZOz9t3NUZs99m
VekPPuzeuc6p5rTi+ACWkjNKZcxM3UJ9UpeLVdBCwDIhSc03ucIOOcLJEEdQxu2jLW7NA33mPHOB
8JjmSovP2bAZ+QODctUcQQyUJOIrKFXHpPAH5cI+yl6FMUrQ8i0fys7JgtxrsYprOLvsCepc++Xj
reHci5QFF9TLetphqjg5+k8ASR4S0FUTkE+lZsIhWStpheSffAcXYC+I6tzutXGIHfzRXEP5ypOn
s8igC6MsjcOTj7rXWZEoLN98NBSZ+mA3eTF731fwlNLLWxFkJ0RxE0/WJRW6SRodhfmp5zMLuF9L
oFGNS6UC6sN1GEUdXCJcKDNUTMeBf9Om8zpUnviXzfwEPUqM8IId+oXnk7bXKSjtaWIBQvFUoL9F
51GhOlK4Ot6GqhsQJ/CIbwyakRnkm+Oi6k6ziG+8Q1nESGQ+fIAFRLuA67OpQUzWSlKf6Tf1Vvic
7jztslQd42P7FocfJRs/KMiykFlbrjdAXT9Yb0p9AFBh8LSiZn2awaMLxkYlM0QwTVxw/7KcvMFp
8l8chea5oPi1Zaro2zIJl1QbHenOswZoMKb+0EHwT93xtMJaUZ8cYilKdSK4BM/85ppN8sLhqSuP
98sg/eQAoGSUIYC2iv0UeDEgYXCYXaVP36hJXzrVgnoWzcfm0wu/qFY62aThzL3bc3ZstwP1KzY4
dOXtoRdWcV1Z5kLdyjAUc2SpV7gjC9n57BbsXvOtQLc6fEGkPMp+Xa4pk/8thecKCOtgv2x3/QaG
lz/2XZbm6ygspU3m4zZaFvyQmg67VEGLsiUR+JangaecOmmvvgCi0ngaeDJ/JG3UdIsf+Fy+ZJ3Y
kGvcaYNXlANY4BTjgRpegkXdseVKpa5UTlfWbsTt74ksqk/kcTOo2QbwD8QMjyaL4F7+0Hb8JOUH
NFqdMc0JWiGLEGUvTBrnomoYcRhVvF5efdHO0Fpm7GahSnFEB1Nwgh6yRhYBRltwGdJeBSsbqU9v
KTIY1QBz1Ovjd+ha/+0WJSVF6bYsHbMQwc16+tty+SO+c+NMS4aEvQQw5qcF0sJ+RhDqBT2LhX4h
PbRS0winOHUmLcUGvGxaLdfY3O/oHH7eKH1U6MVSQoB1MJs/uyXskXGvVdKrkYr7dL3q84CBvEAZ
wjnEvv7CuhKbHxLAeBJk2Ahp1hkJnPTNFa/9O6D16EwfeXiApxUUsTXw8Kilxxb2O/Ih3m8Zg+rk
YqMqRyMXdUJYLJVaxGoczxfWcbQj5YVznxd7r7VjUqeCmaU2hjL46a9z54qpo/DGJrDZ1dAe2vJR
PT2+rUdSV5/VQnbEiKTOXY7hYQ9PayxxZFx/L2ncGEQMXnB/1urTVq0k9MFg4p5gvZRZbuEAbmUF
dEOmXmOk/yV9KR73GOOvpcy9hZA/CRLXW0pFTK5d0cqqqWS9ks5HGYPvh/0Xi17ZAYPoDGQHqpeA
nziF9+TjqSjz+vrBFbq05zadDlUIHOTW+wiMOJYGrwV999w9SfGPvwLnWa9fdVXX7ekFuQk5qNBl
/sXf0Izs13/318Z/GnMJoj6h29PRlofSW1JKcwbU9QS2BjP+HeKElqctifWt6/2pujzIcbRsWo1x
qihMw/daFQvbLsWLWYuhzuBqUiqFKDK3A96eSmIt8CXhT66NuBtGblwF+Vlg/Uk9hP49ApsAPCoa
ULlEGBJIMz1ICGR1jdyVYYrOwyP4gpA2K1S9oHCyd48xpP93655ILrlTYgb4us4Jo4LudRaPL3Cn
kKMuZvDzycWfHbSFZqxCTl8sHtG6Pl4jQcCRM8oxzS0kCbXArFRG5YLK1ZKByjqAoO0JEaRKPWE0
oteVSUGTNTZHyQ+M1fkC0CYIhoESQHQDrdj9PYf5PKIdr3OLJckEvPgcNZ/g0f53F7p9pAymtakA
pVdlbr6XBP+Eucd159ddh6tSSLg9jWEawUHxfDTk2ja9OyIN7o9GbBAd/aoGr3d3YZb74mjqub1/
pK2P0+EY6hTpi05lbVINeY8xw9/C4Roc4BRD4TDYmFLcK6V/Pvjl0lBz2whjbyYlc3IluWnPIFH9
hA3GB1QFyYFkD9RWlZJprA42w79q1cIGt6vK1fLsvb7isZnRojQZtDbKHjdGPgOyUYQ7JC+ydyCI
ZeLa3BH1xtOydSKKgqPnQ62QqXMG49BUruGiobVPKhhxqtNTDNAe407cwK9HUvPhhIJc0Yx6hxM3
0VtId3hgu4AQSPe3atdSUIJT5ePU+FPbW5c2aohJse2Y5lTOQXU3Yi4XERpqTTmDR/MTSklHZ9tX
n+43sgJNwg22u7onyC0oAy4Ua/Ru3zrsMsjXb+mjU8ZCm9pZSGdYXrcECDgodwuoK84wmHMXy1ku
1RS/bmwVcio+TPCZO/a/T9WuSPv5aMds13GZptAb78hlgdchLrxpbK6nY3728QkR8Kh1eIVZb82h
OtNDJCnc5/h3NZsasGNmu29v6zHipO8wKfF80B6KIcSW1mXKpNU8LHLJKIlu2yRPbvhy2yw6vXn2
BVnPVJkNybSBv1HUi0EBaVllACH/oA8/ZZw9+LdmJif6BtLUTgKr+AkZKwIrvf2ULpn1NaXtQvVY
mJ8WlKaHZQvoWt6aKysbkB4ESnzCWxJ9GF6lq44vAs9Wbc1gLnPEEg1aVuLRUtUzhx9UKgryPtKv
xyEJj3+7480nOq6bCGLISgTVy1V1rdBDH3X4g4uShEq+xaD02f6wUYYDKRaTPaIbmcXwA9KAWsgS
Z49jP0lw3Wat6JWW2RCZ0/pFnpOMNmW+Y9vMVcIiqBOd1AcXpfQq+ZCSX8/RFRL7QpMJuhBLwW1d
CVMNcblM6vCTChOBcUpPY0gxbl/hmaqm9kqU9OUrd6mbePbasaJul99QPAYr44HJl245Qg7WaynW
tLzI1HP5zIRFwQxHySSpskA6YEuMSr9dRDd/WPxAVyJBF0jS5GTmlN1ZI8i9YWijIJcizVi+v1eZ
nGKtVq+KH09ji1GDQNl9DOfy4TtKn/jRNMudBdkhE3Ax6c5xsfiVm285nr6DwWNP+QwZwg6ssytU
/qVnOLw9lPS/WqfzQLvVJEuuOKKNNeujcBxjtbjQcTwSTBN1Egxb0zoXinTPr7Wbg1t5f5Wzh1wk
QKMpAt/JTg63X/+u+VsSfvJRci/u6hYms127VIq+czoULL92vI9HbVNGCHg7MXWPFFzuVF/5xWNj
m0FHA70kdtEi5bFNn408b1SJ+0x4fqT3Xeh5dHliXwlbXLMrkszPKVxPImOw1joMVXkN4ic7YTU4
WL0s7IFly+XHnCjp/vokOaPOQa/79QOS627LOWpBSryiH+ZFhSWHG7H6nhDB5eXKDNdAw5UaYcMa
YPELIk1WOZpAQAdNsKwEjh877csOEHAWTPQ7SdfZGMQuMH0IPU6lIzifEuYsDcyGMNSjIxUJ7bJo
hHY1O4R/KBjCp4O3y0dKBx3uWWqv2WbPbW4eYzC6arswcaYeJIypoK4kiJTVFWpp4j5+NukkP5I2
B14W3mEs4F9NR8oikEp5s2RQsZEipBQw8yOtSbY9uQ28PE4kCEZZKT0gW6vkvUfZ7ZmgA4GGS5l2
zbHQd2xct9om6pFyjmRftoUHCO2GSeoZgCWuZdUNrdHyI2/TuZ9T0exGqp/ShlsxttELkd7syLF2
Vr8F2ylz87iWriHOTYGQcQlAtmrH84oTzgfLIrt6Ye2JhYvvVE1f9UME0gLSJXzq9838lN8i8Rjs
jgtyFYx2wWlGuXPdvhphipJMLA6WdZU5dFDitmdu/jfugZbenZ9XUgtTNsK97FUv2DYrt2i7mCS+
Jc0vvzH2f5LnjMCC3a6lqR1rhf470/HTpObhPgaBN5Kc1zLScdt7gs72MWbrbZCqRUxDnHud1vl9
p1xPEXqzHCr8KRxpQau1KbykLlSZbSxpP9bIhHMkTmQJsvQP7aECBH2ryrXt9QDvGiy+PWt381RM
9Bg1cKm9LDeZA9criAI8ZqhoMxKlMhNjsutI/Bnn5tWjBIK5kLivP+EX/ZBx7DlQ4o97kaM+vcSv
IGBJeCxyFAs/cOvSRNg2x5AD/cHauh9aYdmKD7C+quw/shAd4g2RCLCFtJ4zxzZISp7mdEC9nYv8
I8z+CX45sBGQlxEakx12FlTPwTYbmWbKjzaIBzIUnyogSFCiw65gIG82/XYl06zCAm1qYYJVojv2
NvcAf/6USW+V1CRA8D8d+xAlSrRpURaTYxPFoFboVhPbgPmfzNBbUkKaZlRkXs4msQV5hAN675VN
qjGMskzpfbfgGvH2wq9P+dJ0ZwgSwMUXJ+FeqAfFxH5jbd8SYpM7IGV4cWQo4gPpykm0JIAQXdCg
0JgiZlJ8DPEZgVnexuLSAF3IxGDLAJqVBz9iky5XmzBF3gWEuUAVZlGnASdC85EXz4WnW8avAYnB
5eyuhosxIqaMpmIExCKarGI4nenxskUL5nV4xc30KpsWVwaEpBgenGPJ6kAOjG3IfAOPfdJcLinH
AhZfHrt2LBAQjMd6bLml+KlW2NfJ782yTENWa+5KfLzNIIr8m6T0lZHcfP+hpWQID6dyT62Bwuw9
xp4Vui9owaQYmkOQCivaZ/lT4ZC0jVmpdNmZtvq1iYHGmXwxLn54buzGYmfRxoUH+Jjg2tK7wT2Z
BqLvs/fTFrFPIRqVMWS8WsUs4QJd4klUA+wG0rNHVpBiFEbjq+9iWiTXUmgwgQe88GnIVDz6zC7Y
lYeI4hDSuA4sbTZz6ZfzS75+9lcr+WdIiwJsoOQZIIvSKarPjb/8alwGeApi7Uvhf47AKgBwuJSw
OvevnSjkp7SBqhwk63hm8bg4EKjYV0QIlRHwUYDn8xlEfLSj2DJ/4VFgNVej2Jk5q7l+oFqGCF7X
vcBCpGw1bGetrPNrBUuK1J893dNq6EwPv7iNXXQ5vxbVcK32r+kY4ciRnt/nSFIUsvmQSFYc920j
17IS1CBlvYRvnFTggdYjk/piVM6wCDHgoltzfubDfCeHlmTnN2I3luZ+EY1/prkASFqEn+LTJDaM
upsj6iV8kgpG21F8RxbdNakEALwTpIDw0VM/wWhBHikO8x0KOz2QqFPw5nUqCPU9rmH27jYDpcuT
4o09q3K/jNkersSs16z//80zP/+Lux28qX3+uT2PXCR7OKkQA4oennLZCr2RzTEPeOwzoopV5z0f
+LbsmTOM0i78j0rmNovJlb4gbg8OBLyMkUu2a3SV84k4pFncfvt1077Z7cZMuTKSI1qYbIvJU5Lm
zOJciu67UgcTTajwNpMUo9b06B6qROSxQmPpzEnotISkZYysOtO/hDSQPTZUMaUfs2sxMz6HbNPq
cVYbiyX/lAZVS3Dzr5hWTuaIl2687hDHhxqyHGtEOYaXdpwRjuFVZrNQw3SD/hWTaLnNhtkRLKGK
dmTOhXusGsvhVfzjjArTJMHNovKYUJTg1BaaVcUmgPn5zkbP1MCXfNedXscA26dbovvaBhwFd0k1
tAF8PHtWlPYM8NlipMc5toZgNW7Cw1Bhja0sqNoL9BxL/edAAM35Gl8QaTNtz5Cn27Jipeh08F3R
ZP0mEISVkVwF1JIKovvbN9WnNenUhW6J0lb6+Ikxkml3sMwUMibwYj+r3v8bNbctU2cBuhLe/wPS
rMQVk+/UOGb0+W8fNCaEe5YlzLHnbPuQXSVWhx+Fh4ZxGuR6Ums1y13y0CyN0Cx4OT1J8vxjzHZR
WdyVpGEanAMR+8J6+5NewdF08teDkJnaq5FREAfe2m4H3MzFqfzsZ8ZLNYwUDp2LWGIkzAhV6jwW
0ra+xIN/A3SLGS2fQSIp9TAd+TTzpQuhuSl3JYwZZH94tVCSDN8s0e7gJt046vb2plOoasOOJd+7
kwUpExTfCIV1VKvh+URSvspCTpUxv/kad6+yXdPL6x6Uf9sb8wMPj/EYo3R5NndFwh0hHC2GxPZj
HC7/fqAxVNpez0SHd9N/r97NZv34X5ed3yvzTzChfkETmOYsV190A09BDkwMp5YCXCs95qrrop//
Hk6mCbsoEEHT/3GdFA9WyMohrGy+Q9J2n82i/l+/zmRAL5R3dWrLRSE9qqLymGxTkjb/yM3+3DTD
cPpIpoE1sjXTtBrDqkVI2b4TBe5UEGkEmOLXdajTDQ6QnsSDpUthXkyMhw6ri68L0npdUDT/+T87
QTkOYEP6WvmcebbKbz9OCl6xFoWNM/ZyabqcQ+uQ8nDaCmCuQdj5PSHt83StcWcgqOAHs8gJ9AFZ
ev4meRAceZV/i2OCguVlqydOQDg3nVOV0Lst0v/hq55JNPhqjIdJkzDWl5Fs9NJ3HhSoMuxGOlLd
fyL4fR5tdnp35N0MuHRXZt1Ve5OQ5F0QoEOazVhR6NeLKQL2DNdopDREBBrGV9NA47nbpAruKfGw
v/Od5h8BD8y23WiMw/HDJ+u5+kOOqTsWiD9cwpCXFtLx0FM7TQAGsQKOzpxQuxlVXPboBmJwLxtK
H17J0EWVSEgOKzSzPREYwERk1Ymyecxap3GDMLQczwKpnJJelBPfAgCGj1WDgBUdDpfkAFY4avui
uKvXorMvFk1WV5j7p2qfmPaSk9i5X9grt86/JySaJ1VAUWkWOJSfA5p6+kysTHRteom/O6RvXGmC
cdumw3asgAtTgP42qeNdmZwM2yzuDU0PveMlqxVahNd+eI0Zh7nNTzLPd4wCIhXC80+nfT+sUFkp
egT1KWl7EODGC5k/gKkS5XmSjC30aubmssOXn7Xxsia53vz5zQ3hb6EG5p/oLReCl3cyeHPXqrSg
d1ATjM7Q7T6JHK+EWHyKLAXQmYKUgOAd5da88+Thva/4vzgYhLsZS5Z3Fpcw8AQ8mbxC8j3C3xIF
gw8UDVaNVmq5oC1rvuBQQn7bh/oS89xdM7cByD2WILvfeXaufRtDWJtAa5yKoylYDhZEHwOCChQY
R19R5SUz53fKeONSEauLEZ/9HQWvIs/buvG7qe6zBK9mPDfnSGGkHozQj0S/YxWkh37/nkAw3zLP
cyXeCp/qNbxtyDhDDuFrMFUF1yHKxNZkhBQ/2YgjpllKqzte/C3Y8Mjw4DgRgueZpPO6fBrDdg9t
odnGAVIF+MIa8Fs9jYyYAYdy5NRslL3un+eNTurFBI11D4p+fH6ObTuj4+XfTY2UcjZVlfo0ox1k
KwCNsunTq98W0Kf90L6Ejb0cxgCD7TDSz3NDBPiKKscPNuJfh8UVuxYJOhq99qHXBhKpwlVqsDj4
iqFQ5+N4v7cB/hMgMsnTadRQzaEGprRG0pBnu+1dn6ynsdb67eZUq1kaabk4sv7XVQ7tEFqhJhi/
lGSjOjdCPu+dBAjJPNZ1X7wjiRqlPmflIgvQn0iNIMF+/2HsejVRqAYj7erD34WH/koeVj7t5CJM
vQtnWa7AoTNNXpTpwmkLz8WCBWMAD50C6CGtnO6IeJsRkLU7Ov3ZJQy972/JePZR6OaAdtNpE2aj
pImlu0UQERDbROIOYo/CnrrY8nZCYyBThsJXx5xUo3wv126FQDx13JqIW6/HzaRp6Wlfi+gq4+bR
D9b3/eiIL07LBDNJSTHQBIZffNg/XO7KpaUxhlDP4pfYvJIz2ic6Fld7f+I6JgNlERgq48FonkOf
dEbLSUviLrgwu1GJ1sbCErD644miHU7DRFW2JxGQFSK0hvp/Y9f9Td3i6Wve1+/pvIWBVK+gq5Xm
62GCEvRd4UdGvxuy9YsUVufiKjO7fPXIooCE+JS3sv7ALMhy3Ov+jK/3DjUZH7E+7euhALgp0iHs
Lf7pWKJgkOP/CDyU22buZii/gc+FL3Hipvvk2DunNCHnqJoSJMukqapZMDIboW3XiGvddfL7f1pb
K8e2ZALU2i5wQgoJ/Qfebvr/ln1csu5Q67HkhnqQaaNsHM0Ap1G/Gf8saIEx8jFnbOoLc/kDaVC3
dP4OeYVtKCxZxrr0hBgMv/DyupD+UcvPFGTDjBhDj0JgqSNCbaZw3ltfMz6jTHJ71T81eEMsRzud
SjjFh9LJIL6vG1LfXa+0G+aCTJ3M2pMuSl5sAIZwx+JJvk+BV7RGus40yfmmF/l+zU4FXfohjUqP
M8k0hMaffORW3p7sF4NGQo+sz97zMpoXQXDU1zoqZcBAKPFUNuGDm/OgWvi1HcOESK5WGdl6JMRm
o/yZkXDfpOvN2kLjTu9DcKioT2X9q3uoXwZfd0hCCPa+bB4AFdwrJu0dEeqZtyWKL2+0pm/JKlxh
fxseHyl1igze+r1kv2sWd2FGm5WkfD5fiiswEp5V4CQJxPfxII72MA3f3u/cMKUavFWL1QK+Dls0
9J1eVfLmR0Ye4Y9KAZLsumHiN/FBiZSGpt/X7aTmzjm1oIRBb4i7+yTJnNiwuxLtx95GxTs4q/JX
Ls5H0GO6f0EpTkiyX0xXmA32vY6XlSocQf1XvILl9CKrYGijzDIGElCuFn0zJ+wyFVM5cWFYJ0Mo
cS9h8SwFt/aMnx2L1ZvC8ByTuKdnLwEjP/37v0HvUxJApEw1GQ3lCiZaOiWExJNY9JkhvuSnRUx6
xn6YrEOmWnwPFi0Ta8d8HMhGz5SFQKwmN+kVGczLbKZCWmBInEcu6JwYJb6NsuT4ZSTi8xU65xVL
wsJqnwNsmJdJ3KdNy1/wyzTinc5IKHfU21HNO0aUGKPORc82sdh4jEc3MzUcjpMZdyEhe0gOm9b1
AN9/6ndRcl5zdKZmcrBhSt/ErNg3Ml/PrrO7ZTTieBqktUsVnFGVW1j6T8geDyHwjytERnepcD4b
a4AVvqTMTPggHhk4E4coMF/ChNhBLd1RrmPkZMjHVmIhMAnrMoZn3ise69vr7vBbpk7iqPnDP6Uk
2A3xDgkIvDNVuJDVo64H82tgFINd4O5RfF2MimWddCneEgjUnkBoAGhFQZEduKYX+MS6VVnc99xz
DPPnoAQQZGekMVZ399c/rq85TcotRW19fvttMIDgMLo+vUe44c5UutPN73NyDNZxW+U7Xovj3Byk
MdO00wVn+/pw3aGx+JInHLNqy2itKQxZ6LElEz+tKi05B4ORVjRwzdqkrUO1tSmUp6UhKuuBZu0V
kTvhwVcYHLRZKzVs6EQJa+WzGd2/t3Y98prM8gMMlIsQGe//cBN51kg/3nhrmhVrSts1FIa62PlM
C8NkV5YHM9BDf4G3rG7RfwSCEPFGgHwjLgng5SeDB19sD5eOS2YqEfo0gOzPlJ2RpuRcObDgVR/H
w19vQZh10pDMm+06kCQm0PEoIsGJnLSofPdzsB7bE/kNNg2mjv9HMwWW8J+JIg0rNHCkM+6ncC2M
qOBmRMgmPFoAx/VH2j4SPd69jaFkBsqNH31qzTNuZM9YB2eWDv470b7Nv8WXNkJwWoqky3sGaVLY
L3639jyXqXms55MSWc5bVnlqVcquSr/qJ7oiw8Qld8IlhqOfb+cLd/GDRdgVirZY3lsJihRQwhen
BfVeG9SV6FMGHCSZbLm/Lrrsv7GaSXLy10PmPlWqmKC6bqCwKEhlx7Ed13FoowXOQ0qqt4MdmimE
+CZpMsn5bv5GXNc+vnKsNjxs/KhmkFnDxPNxq//UFXrDUhBua5LjGdLTz2XvPxasm6WiXSYrsl6r
turwc7CrpQdkJWiy9x44PIljLLHcUs8SfL+THB4fE2g5+g2p2pNQINSRhHcximQV4bXFlAMWZoE3
1u2G2wQ8DTnXwGtShA1IC5rUA9p2Mv+wwc7caVpmIuSIO6sq4yb0HxFwZZqoX43SDsub1UvyI/7Z
uyokoia0g/Knv/BYbsjmhx8ty5Xdp4aRudqlLeNQbK9MBbxtCZyi3Rd0msc2wX44AwCdXxO6uXH3
wh+0hqpEbLpbPUXf1OvjGxFHBEHhvefTwG7sOVhvkt7Qd4xIMpiwXR7pjbu/AK0qCKOmJsQgTZcU
FaekIlDw/ZzThMG7eg9F5arGl0kNkl0Jjf5JvUN3NoMcq+AWcdq3/+gIEHGeKEFZ/0AMMEQSWp3O
6b6XZP/GIx0mUhDQbMl0Zg+a+BBPVz3MS1+O8dKUw2ITbZZIYExVfe8+bB4riqgXQeRaPoTD2LhT
8iAWaqGSIRDZU9sLJW5elVZJJuy7HODBCJ+lE6AazISSIul4mb/PEyf6LNKiAgHMPlCl+t753axz
6fQDH7/dzq17wPEB4MBvzZm+uesSRNyYrqB9MKuRWfMCcPxv56YLbKBMraYONQQjkqKzMTkmGos6
CzFWAsVFYBbdmp9Uyzf2OSufTgNjTlbLKzK5dTI48lLWfR4cYYjTWwZ32qCcCFrxKm82eOKyhtTR
1CvATKP2sww/HcguFPW8GMggDtNBbKmgvUsNUhfASeBJiDCWxbIsdVyxpOpwKdaPdRv2+MMBhFfi
579OMDMizWyVE5OO1IL2qL0ymWuehrGhoMtPlmZYPqOZGqLYU71uL8BDTwuS59B0Edd7GX8XGMZE
6HkSiKStSXECi3GinXOdZWwOExlP5ARFIBgrAsY8q/nWEI+rK9riPM5PyWjR5YQdYEf9JYdI86r9
B3Px9lrmGVpeJVR0aNP6fKkpfN2xFRLPIKXjlZ9o0im5xD9QIjtLjvs1BI/tK/B/H8RZ7dRQUTw/
pD1VB/OqA0/bryyrNVZMcAjMTsA3X84KNUhjMLDsuNPAG00MisXtud+EFNcec8n3sFcZhoVaur/L
54Edos5tNxtXVnCvbw5YHwqKaU4yJQCd5YCaRpsdE3S1Df9fLT2tpNAGftMi7F5cuhdwq1aQZZDO
iis+1BqWXH2dSXs5X8Q4cvpw1KPE0oaqoCC/ka70Wvj4po/hdfho9etVoj9UZWjD5yHBGF09wQXA
2weFwNavw0y1+vYGAxtY2LdunzTM6n1FyRehor8+sckLb9Fa/XWmr71Kz8Un9mPcX6FzX4rrhBqO
PCnxy96VhDDSywnQx6kPwY0vFsY/oIYEHyvQOGVhENHQkeU6CLcngdqobi51iBQb6CpdiXM4eFEm
l4FcwPt7/rcotyXRm1KFFBTivk/BfLKeJFYFLEoFONgpua+C8F+ajzjX5qs3vyt2qCn5sQ4eEusp
VGL9KwPlODakZ2EhxeKQRkNwzbnKmhpud+Tbg5MDuXtl/jcOPYFJ8aIBHFZAtNicHDr1c6zs0+XZ
vnW/j1Xr01UQFyPa35wWI510sFE39dQJqVuLWxRx+INO0yjj7Z2eeK2VIy1c+GEvSDn44CgiRdOO
IkkRjmu5V4w70MNbRQWyYqv+De03L3KYpJGJwsUF7qVqhdyjIZd5f01uwB4Q8GtJrugUuE109Wtr
garqDOkU5AzRHnLjyNUKq1CHLfQ+yxH9CBkjbmNGRVBX+PWF7BFJ2/w6ianB+HLoKnBVQLOCEpDr
BgLJd4yUL96Q9KnSCBY8qUqVh85O/Yvhcp2GALjlXDGK57+OlXE0ai98KKdRQDpnDuU1E9XQu8gw
EbAbGT6xAD9LJ8qjbvFiVXVWj7EZTqOobthprlThYFnyAxq4os/u0n3j+MNQsoCaLliz0akMrv9e
yW6mAepqD6XgxTCxphomnppvzF3H9iDgTjK+sYduQi14y8sPVHQWxnscN0knXR23DcHwuuGTRHGq
vACOvdxw3X8UDmtHPCBie7ACWv/QytA2GOGerhC+eA1O2mhDxS5HQJcHoTr5EnCSq6IZvMjzO22E
SoOV1BoSqbmF646+w87NJ4hc3a3hVoDhUNP4bhguXwX+2pah29b5TcxVcuzJaC6y18Vy+6vmRxfh
b8ZzYMxyNQr+ekslO3Hcpj2QQdHnEA/NyTqEBbs/LMPoQDmfnx752CEH+DCLYCney2b6zY+OKekv
V8UJ3hsa1OEHLTJU2AXvbBZr9TK0MwoQrd1FIMH4eFZ7MTl4AyczZPH1Q2PZx0QjSKr5B01rGPSu
+ZWHWONdC/KCq8k+pOktpsmNmlhjwVl0VYtEVbAS14sMWA75gP+BaYkcQJI+EjImstqwdiZvkvEC
KeEoNl8IzF8agjI1QNM2B0SewLaE/p0P47e6bpwMAkmN2mezgLbddXcMrA+gzFjrtiDCmNDdT91c
u0ao17n61V69ta4ucnfaAB6Vt0w1aynEmEF99e8W/K20d2iSEOxOiQYacwUtkDaZfE44WqU2xbnG
j1Ix/pxFy6H5voaT3ZL/iy/u4hdBgZXOkg1YGVDIcF8js89fpstG+6fPjMQhWvlFRFs/ScRF/o4i
C6EMSAM94Gju12XGxl+llJhnCaeMk0lvQHDssjlwJ10RJBdcNL12hDtWJ5bPdjCc3tYVP8A+MdPx
huHF4z5XsY9VBCK9NZNQlig8bNA+gP2NgVx+9OjdYbS2vK+Aup3nB1Ip4ynolB6Sq8SM75jzaXRm
OTL/3y13rklmSXbJ113tl38uEwb3uFLa27mKBVXis94X9YkEl9N3MCp0ryrP7IxOUzV1OskjU3B1
nhhJqkQHBdyxJ48pVQyiqizPnDdjCE9HiQRiJygV6xqeQ4QCTqJYCfFqR+A0U05hcR5ZgDuiycHr
i0Q2Hv+G9BQ5zA1DcQkMRyWgo8C9sb+MiIXYii95AY1XT0N3n/tU9BDchvUSEzRa5t/oUVaHggsh
Adly9wIUX7p1lHHZ5TD7HJ1Z8MLwsICeuLSEtDrpR+V6qJs49mX3b4lMz4M9/r+NE8IC8Kiv9yaK
exPajbEd2XXkOjUOwlE60vQhKtVd99d8XibSgEJ5NrjkEjVpifWQvWyG9ROuj5+ZcBrgs63pv1LR
8H398uELGPteLaeYNrZ0+1M9JZ1/h8p4sw1He8cxV2fTGvmqcWM62i/QhnIRoy7mG2ypSBzXfROj
y2tXheMdwpRAMXB/LFjqY/DS0TBty8+KnP0oq6e0sA6tDf6YHIFcrR2aBNq8X+rhWtIleJc7A5Qh
s/fiYLHmR5netU2wUeW8mAJNO4b79294pyb4uQ5lxcirDOKZvE2RrqvZC61FShwMtMz4m3cVzGwI
I8IW0217xRTDvfVWwwmgpKlmVdMviUZwxKdga2MNenRaMQUCY/W/70lYCVDM9tLhV1CVvNtSXzmN
laNKlkEMUXDSdSzqSyTOCq9t6rPPLHSfMA7YO9QGIUYDFGaM3Gk7Trsmt/DDMvFmjwwiFjygcl3v
OQ33Vnp0gLmCCWqp50YyD0ChIn5UKh8nelNs7jY5DkxwSu8JYPc7iriIB9Ywwrpl2bEhoGs9ZLCI
MsOz8/PdSN6xrGgfZl7AFUCEDaJ7b5S4RitxKvwV7DulJI+bDH0tlA9vWKL5iVXOpZuSjsIq1d7x
PEZwed7neBVFq+vTTCTY0TqD6tOUHuf0ahEEMzvA/cDPbKlF5v68kaDZhoxN/NdaP80xgsx3fK/U
nLbsJrCdY9CxZOSR6UEAL6k2XVWZRaf3pxnbI6Cv7kIN9XNFZeA9iFFNJYaWn9gnytd6rYPX2jDR
ZDwpOUNef7MyOeqb3Odg+8T/e92x7XFzwV/gjqz98Xd5lkaq14yTBjfsZKeUkEXKsrFExG8GUCE+
ADaSfUpUBg7LgAw5c3/FTTZeaaTvaF6Xz/lwgg+umEv+EJgJtQXr/wX1zCRI0l9aSXntwClv6Mcj
db2fSXIhvlsQuDZQwzd7JtFcOu2ufd8Jq/xa7w0vBDlcPVhbOIS4+0goa+u/WozBary4ii8wTS9l
8bHK9X1UXjO0yMBOifbWrB1V8CxbN98YGYJdHpg/QdScG9iE5clF2R41GH0yzg8WNb92L9QH6w4r
A4zOL+XN4NNKaPHsYP9fiVirxIrYmJfo6U+/h8ioL4TXHs4Q2H8/5DpAgPw3t8RVFxN1NsZW5OK8
R0pQa0eZcbb7qqqCFw3ELX4PrGjeqbGKqMF942AN+yRXusWe1J7xttX+dcCp/1wk2gxlaOdL962k
jVZRolvICe763eeKiqLnN4PfT3xHttoyqlml4q8H9vaCAUdBYRfp9xufSlYNgAaoNZkLcD9r3f53
9iJt59yL2h47WCyfC+nRTIMJWjMH1bqGMLzklshcygHwVOBJQhMNp9xC6TpsNYTF0Xji0coot0gF
4oJZdfx4BwjxwVnj1zbZYWUg/Me6hQMGzSEH5SHafREw16YwJNO+AeBLFXYXvyqc/awEaU+WS9NJ
H1S9dHx6jNyj5qSeGJAnQ5rwk85KLVmd/AKYruaQ7FS9X8xgFfKEhJViNGL8BsbVRGhd5Yj4TIT9
MPoyTxN17017x/aBSyqx8eB1IVWOzQTyCo8Q8bjf3n1CFMKYmqvX+Ghozf2WkEKKjFzkoC6fTMuO
CJ1ruBKst9z11F42DbJj0xgVjzP3MPExNilvd3YLfvq6hWgNEJq4u8ciASUfCTOqSqMJpMfXAZu5
4/WLkzHcwWjMicrBlrAUkoNLNP0c+Tgr2dyoPSnQPvuXl12wXCnyHhv7hWCIznsvNrRgm2oSI2kw
vEUU0mONwlASDE25Et7yVrrGGsnEdpxbHgCIy2q+oKZBEPehCeIIiL4KNwR114b9fPHA+sKo4jpp
As+V41oTKBv5WAhT24PfeiLURA2Gsz6EmRtcd7PmWRJHVeOjCaRpyj+YLIc7Lhc20vRHPz4K168y
Quh9UicSi8x6/cOQtdiSFR/fW2kIvgyj/HFa9YUdEEHbfo5JpMy6rhV81oDbXlhsgV6gha/2nK+Q
J20KYPzur81VE/8x9u01VqGe1kd0E1m5VYaURHdHheeuRhKmuSMG3lN0lqflO5s3CrZaCEEckVTC
J1pfTo9v3NLPaKnd8ti6uVxhHDYHu6iduXRxCGz5c7lL+aSsiz9/J3WCGFDF+EFhP5Q36Ywlx7an
wimcZ0WL/m/h6yf3xXAkN3BPAtAMYPQPjvyxUOlZ92IsoGV3BhpSw9xfawQjJxbHi00HVJwXSzE9
Htg+1dyfDIyJqb6D8mbRGxiBkCecbcF7vRipcDfS9xaGg8wcc9icwe83kx/yMpyB2ZVBDV22r+XK
EDHuR6vjyFN8WahzFY4IWtOjrtCDQDXjcYtMLh/Bp8LOQsl7xrMh9alLj2z4slJcPWHPmLpNxsjh
+X9uW/7GDC9aXOLyIMKZ6+sWHCgzVKzPqmtha0oU7pNP+iUOrBkyCqT733VU6tB2YOtneBWr0MzI
D6la3bTKvwqhyCsCcqjQyHYuw6rIrHRwgXMBIcxAHsmnZ3pZxKXmid9R1leQYqHTw4A+Oa8GlWxj
1/gYZwty1RI+HSczqlBNzIFPrM9cRd/BMxzKLhIxliD+TAKgCZQwEiHfx3QVCx6Uso9TD7GAa+f8
uO266UoTYh3HzU3/HqQkTDt+xV1cP2RL4bjGbwiLuGS97xNXTglEZWRR6GuOqtHJ1XSjBTgkorcM
0kkdKV086Q/R9bhJzHw0JfRgnxETPT72ILsBnkF66QRbPp5jj3GRBrv30v+jDhte+dTYQUkbtY9H
JHp59ojf3XXo6k4UAu6hBRq4Ii9PXHJ5KTCxwjBl8ZITZSz93HV86r9RyG/saYa780qLpQQpzjLR
AAtCkimhvxOS0qmbuA9vIpShz9yFSPiYQHTHqy8xDHGfSDvwsCaGSWnGrWXcbjqjWOG9CTeZxYq6
euvsN5RuD4t2cXhZDj31C4ZHSRSWHtY8iWOBgEKZ8/7EWeDJrTp+a7kSzLmdFG8xHG/KA4JkTNNF
Io3eW9uqYeFi53Iod8XiK1XQRC8jdYE/L1F2GdakabM67i8IwcA3oWdIG4+xIqgT8leje3kYLZY4
gbB6ebDdYxSKso3/qS2jVGsebMhuB+i+T6bImKas5lRSdZN3WJ2PtvZiUT19gpSYyxIgejq4kx4W
R/lBxHgGGLMYJnxvI/G7Gv+f52rbYFtJ7G09rvrmS/DxE46XhppOxDA0SbANiB9z94lEqOdhQBlE
aff9JyEuFJd6BBceb5cbSQ1icgHZGdqwO0tCaN/A07YlhPLuNjN6XFVEQydN+oOwL4n8vYzODe0P
lBT911GEbxcqg+s/mc/bTHsAllV9Thi2x3/Q6KEw1LYWuLHJvySO+gIyOS+YPwpXrD5SrJvXh1kp
1XWOd17s5RDCIIqhkFJqFfNgpjh57+jgw9OkCvyW7Va6h0AaMg+h7d+vdwSNclhghQVvqaFF/6/q
WbE7IQ2T1X3AXwXGoz4ZL6ZUHgpmDdZVd7/ivqqBKa0TYJ5SqGnkFLkLYPlmQvd0+Ld5+IIzWE5O
TFjb9xX40LpvQEryGjqNXlpqlHDA8j/6a3GVrecTu311vrXgpvvEAjpA59AVrZQz2lE4ogpPj2Qx
ePZldno/K+/he4uiHknet47/4jsP7PoC6i08Vw4IXeJnxNXwoJnW9Q/0Ar25wue9q5HlK9pR9ZD/
Q906+6ICmY8YGbO1nunf7uYEFpzJUztZ3lM31gup8KYpy0DETsU5UUa+yNsoNMYnfVGWXMoo/kLf
RBMWUmb5RBR7fEBTP8I08kTa2rP8WR3X5jx17gOQk+KDK8btRt1+x84GQ5712TKeyKA9NzudFX1H
LcCz6ivBPAiKyu2qkfCGBX4/ovC8Evvgf0YiZe8ebVtfNeG2oUIhzCo1Ys1Q+eNros4roeT+t+Gx
YZJrfqIZIKGQIYX6hZryO+ThyhbU9Xb6Ml6pLjHeEt7RChfgKMOIGgOFGyY6+KarAvU8LJiaYfzi
oAXrYEyaicVspEAtj9yU606bM2axasjGsdG4CCS9j23+f5ddgkZMI5cD2fhfgHCD03N8ZdDq5X3H
ERnUGU9F9rL1yHtWpV7STaaZTXe/wjyGeByQolid70dazUvDdO0EGFrcZ/eeXGBMZhljpze2mbiG
ICcQJWcXLh2MDT/mOaRevF71CdJ8qH/8ZnweXVqJNwpfNtndGaytrPB54EMja5poJ5J2qAlCe6dI
NTyCu0C40LcIFCjG1sLWB0K5eXzqypp19kdp+xFBeqntUGaLl+ya1pZW+WjuIAG9C2bOQj0Tt+xJ
tCJ0S1lCkYeXshshcibtYBRVjfKmv8kdnq7Yd+123VPy6Cx3+in11KBLS/XYEzsfuR8ub7ze7IYJ
q+Hj+GHJRIQrrcJ3FRYmV4O2krfttmZJydPYQ1bGyEa08LUcEs49ikQMpjN7bALt9Lt/bgPmoNaK
FkhN50vGrRONclnX9NuXgYKUooKp4CKWMaQlfvQSU2eiB+DUHqS1sYDRbemBJv2AHaTwgo1ts1ux
KK7udDStMoNKzHmLGFzS8PWfV40A7W5rZ0XCb4DG1IgbgWtXmjFFrOOTk8aPvvLtmVqB4YItQbVn
Lxim/V3FE2XW/t3HjbxSBw7tMk1u0YnLKjK/4qaUinz/1mnTr8QYPEbSduikQs+tdOSbPPJbKjJQ
QV+d7NoHvbbSafM4jcFwicKNGyoM/zlJpPvjIuIes/NloaliL2kB2J/E3u0fjjbfVP1B/Yi3Yxa3
ywNgtKwuiCoYQ73UvJVpHTvPUKxydLbZx8XF/dyJrM3arrpRPEPZOIz5XkZVwQnwtybY7nae0MRI
V0ww/e9PHaHCfWNsU9y4CABu2ElKlLMOyP2HmeB0Z7VzJXUKEvi0FpciEKbY+UGMHFHFA6pqC/tR
VvzdIIeN/0O5OWSIbaVG/i8Pp5w2NJAFs4oS0rsiXsJrMXC9eniikxNvfTI8XZqEO2kG7YgDSd3U
WI8S0yTcUNBVeiZXEegY9Xpi8VTPlo8D5jA3ikpANo22Z3uAxn/JhQ0KAIh7uF0R2JYFXzSQa58m
DGmt/+0yYZel2optCUj/VQW09Ib1GXF26l11tyBc8y8sCG0snY5RMm9Erj0x66uf0cEQ3k07hDyD
2R1ypUSvXC5HMSaCc4OMQ3vzsCUyBcrWCO/cbAqT1Pmix8qfpfDP68y9fTigfXgc3gn+KHAM6OLW
wG+Pz3qTrGN3MqxT9zj0hmwNjV85sRaewQdAnUNt1zaRkvhqBk1cOc7wA+2Xnj2ZQKilmzqsYPOs
Dgspi1T9X72dhiut9PRLOJZXSZajBQeVw3+sBLOUaUPSST8PWDEZKTW/AcF6+4fg2gT9U9wcB6D/
bjqpwWuZqNz7FmVeQPHWp/vcOaOJZC121BB3bhI9CGFcn3ssgmWO5G8Z8QSprcUB0FV60wS4C3i6
+IDF2WtDIkYI5VXCbN8iAes6zqqdjoL/eshUgOlW+BabWYOlRYoS0OdTsRERM//kuiyzFoTW+f3l
k8exla38xr3e68T08v8Zy9RFFFW2Pnxj9vdWc96LrPo6eDXcoeerVCB7v42NXWylY+/X5cKeF5sz
RJacqx7yJrLEl5f+Dz2vnRDR3RmLdozk6QmEcNK7q7T6f6keDiUdy09V6WEhyXHvFMBMafAbIWc8
TlPGQghJO9hHTcOTuv1+B8KvxIoy0Arb5uU+CU8Woty2SGjgsH2CtTNo1Ow4Wk29hMQOGShtr8b2
SIRaQDUI5c7gF4JvHUa0i7HRKfTGoL/qSAJWoITaXrHvpwCF6Z5SHcb0Q9eXQWaVx4t7o4Tjij9M
ALQ4gx0Fa5h1p3uKKl6AuP5kDvjzH2VOxuLTHWVTJ3v6mm8LqBx9M8c7DrS9lL9qZkdVDyA5h+E2
5lyK7g5obDPjJaD+u1G6+8sUKpGNuQd/9tl5ZUyG4jbkyW9613hyIcESEYCX8JVXUVSPgrC/PEmo
RNC4drcg4M/mVYCEx2upyB+7A/Ec9u542LFFk/1WnTEc53pnuYjmnS7Rmj/vMk6dF0vfr672JdWE
WIchF7YoJorUS8ub8FUYSVJmLwZ2lnRpu8Y027FanfWlCWEmvhVwEaZUwG0DiNzGyIyi2drPrTmq
aLD9Xi2jUDHayQ8RGWDrvjil58Gzk3TsKwGo+PluyPuODLnMgthfj2vRh9y/OujP2VX1ha80V1lr
Tx++vyWu2ok+dlZgZ9wrdfnh9JUkqsnyugGxPllBK2IW1bzvwrKXrA2VkuVs+qqxWPPa2+lCZbko
qetwVdfe6wFXtnLvfDc3utyAkmLDcpUi7q1ldUSlzGH033F3ZRXECUbrOcg7r6nXAtXswa8YQqAe
3anjRjvjF4pS/IfA2K/l8ye8uTKZZA5wZ7LTlZ/lAFC+3CJuDKF0P7yqMbrvcm2hKBbQN5aFpfoC
xSo+sJyK+V1J/u3WZwix9pBCeRr4SQAh6kxQzX40BcxKUFK5L1R/DnnwPiysU5cClUvBn7rHeO3J
T+J390+L8238fNHEMJyJr7PM/9D0lsExeAiXLovKoQvq8z4+QPgzAGRJU43pyx7G/csTcVMmV3Yk
lBhQwEij7dAtBDfzQN9UZAVa1yvejuffhb3E+7rAcOD9YGCDIG597V8oxNrd54SIvnndjDzDxuX+
ASEzx7/8JtaNqBdg6DTUxVuosZ3aPMbsz5v5I7VG8ELa7f3jo7KBrUo0uoSyREuku/Ju3e+3kS5Z
oULLfDMWrzLdYZbfgMYibyskxAhGOH2sG1wytT1XYJBWlm3yoJZuHnuxhcN5ubznb2BBmeQoQEUC
LIqh4IFl03kWosqwZ7KBkX16Cn6YyFYSos8FCwxu/YgOtPEr12sDxuQEhlvm9p7XBTmnxssyujEe
ULhWz3t2vaatcVLfGJW6wjln2FHsZeL242Im931ZEWtOOfSS4enpL552Qwixznv8MBSgiIZbh2Ik
lFG/4W0Joh9feY3vD0yrY50G3E8ldwJlgzO86d4e+4n8sHQi7XcJA/0K//Iv81hw6/3rnlvRCsjc
q4bA7fEYE87ZFu19Q8CvUBU1f2DyPI6G4ZYNW/yGSaTWgFj21ZKyT/czaYO62hmhFkdWpeKm1Brl
QunNiurT/bVCEJUXNjBYwSTkFpTykEmnkqn3JfThZbyennJ3o25VJJvIZSVTvXzsQRdfiXWDBo9U
BQn/5VPX1K2nIuRdOLUzCOJnp9Bji1k/jDDdNybh7rwcgPb7Bf6rAPAP/Ag+tJmy4WSASYp900AM
oisDdXYwX2zVBFiGrM+zVXyNIMqZSimZgJPFEB7yx3PwVXi217ZsrDApfHIJCShFiigXzViG09MU
cSXPNE09KbeBrVQJPbDppfkNzvN8EYwh1eq/0kzmum2N4x1uLB/cwndZ1dDonFLh4Psyo6zg/V8e
oTOiSup99/7cjcfyhIwdydjl/2pTejjl4fDeOMAT3p8HhKSyMLTm54nqToHDf8qSFSD4rvjzUItB
JHs71We+ezMmz/SADkKikjVHzvBhazmFBfaW9ODXCRWSKXq0kT6UMUW2pshhN/xqPOjVTho9x0K9
rXkQyXJgANoZvGtSW6uiq4lWD8ac7GPZv+a6IM2m3g2GINOaQKbH4F4bZt+T6wnadrP+Uh7+6sqL
3f6maS08MLJ5ihU9atgFAPhoPpbvq019ArZdhM7mtwEPH6o1/btzy+jDtc9BTs4X75mx/c9WyscV
sZVCHXn4kaupbV13cu3yN/0JdZHeP6oz3iJXG86qpl1LbHa99Z8okMGQnLei5YHdz1WC4WYIWyrm
vDEClvWGDHnwUTuC6V9XQ7Ffoa/fGZGZFgzg46a8XxKcxDI48NHKZxt0bI3ijAjCl4MK0YPTVQ3f
OGj9vYcVUuZ0V5Yh4i3JoGSxRgcWq/kH4okfdYRUjqI1puJx0IGWlnlUXZszLWRm+kAkqZPNlZEn
vHF8iUdFrBy/lGXZpIRe7Jqx97N0Fs0x6H7zrLVSfbrWssfbspqDu7kj8T3W+k9ChffnzrRvLnnY
HR+jWke/JSIh8oMFE28n4bPXguXWatLQQS49Yj1Zctb1RrTJQ/2FOZ/pMgnqSdtqjtxAkddJjz7L
QWIxCa+OeeqrmyT92eHD/Im85VnPA21QhAH498SpRx2LpKuqvibYhk/sM4lvM5U6c5XbwuR5cYvC
ZewXRcAQ+bnjqYv7nfgL7BCQxkf2Z8JdoiNH/5rhbZ1LtxC1d9Rmp7mRu4sXeElxEeD/dz2R+k9X
4JjU19tE5M6iJTzCDV9EQ0RmojYapT3r/MN4OjtSJvropfVEpc6nLsNzm8Px/8GecUBqAuGXoWFh
QfIf3e8DH3jy8MOIU3Aue+HMk1NMJq61V+DZZ7S94r5lbj+cB/USWG3wZSwb8lofEqo9yUPc+aBm
yxRZ685dpeYNhFJFpDmmH5hOMcq2ciYwNK50nkEfF1SByWbGee29BqMatwifQpaBvzJJAn6UkBUI
A/Lwr6sTzXlUzmvnwGWo71b9YKFUTmCjdqAv4YpH54hFnNKNUMsh8mwhN7/SnIM2ya0C2pcFdOp6
K+pNpTDQf2b5cLtG8zibx3VTgJk5A+BmleIhVnoeOn6L/PAwtwlApwX30wrfZBrUApguUopejsua
B6U/2Fyil8cDtE/NVF0P/bR3rWvr/pStWSU9916ki5ZfkJq4oY9K2yjJEex7eisKuavCK6/6KTmk
q5l3VIHvjB0gY83Iqp6Cx2OQt4QdtXbTWcqP4+F5IVmFtTCG/R88EefYVaGo0JpCghw+v5WEq7xV
1TQ8gLZYn0QdzIzSOPqiAlWDuIx5fw55YNMtdxxDGC3dtSt3G3TwGF0IjiySgRb4fkVMGYEelaVf
XcU2E1WQ7HaIAvHItHQbc4Ris8/IKA5iCilXIsVtVNB8oPJBJbkLGpTkCfczMSlo6f4nK3ssm/HM
EGpTDBcDPGRUQOSE0/r8nvNJOc/d0HmNJwI6UE4WcZmaM7wIboK//Ky+xeFrY26kDt85ZNopnCxn
ZQs15PmWgi52B7/Me3I553xld/hw4myma6CqWmTNLgy8zYSbBE/beYGa34q89X/0W8tbTRQHNr2W
wbAMzvdIsoh5eiy/264Jqyb+SScT0oCx6jfSjhEviLtwyl1vMO9M0lfVRde8M5df4nQ78AjlLnum
yMwc5W9ZGqL6qb2VHJI5Z9foxWUYokgySDmVGdHQ+lAfrGZ48CY+qb4u04gqoAmWNvSW99Mne3Ga
ZrKJVyeIvlRin6vNO4rBJMbvOJ+8HldM/UIaJzMNaDQaCXk7NdR3D4e5uxCP6DsA+74Z1sT8x/UA
DgEKe4HlNC+bE7ysKC6oyBfU0meoOL9ix5j/EtmvKXK4Cgi2friYcUJCZy+sodLhFZmkdzImTRUy
UwzJK4cO38GExztBdJfNrrW/rnvSBDa/scB8US58h1Mh6oUYzxv5etAm7pgdn6OxsldLmWyiYA7E
XsTH4PBVRbAfviezSkl94pM5FtsOuWGLRdEmJUxd73Xq1cyuguCYKpS4OV5tTboTBOgp9rHalcPT
RE6BdWKrNpqC5dx2N84z/jh0xSpVhQcVJOZtToI+vl/UPbdAv/Hac/PXSPVUi553JhZJWeayDwt2
LWoTOioS1EVquUuQe4C+gvA26RyzDXpW8+aM2oW3ZZaxknVvHpYXnelNzi1DUeTdk/OKe8uhNoYY
prPzhMxbIX+3on3+AzX+NqsxWRBKtuEwrOic6y+W62MUKqMka1XHWuWIiaUaIJcyxgIrsFJT8xXY
2xR96XJAhKG302qSQ/+JBWu1zgjPN+Z4y2rAqknJ1/j6C3UuIBX+oe3vugX5ibhyQYYUFLnORwtd
ARbqRYGJeeSaVQnz9RVXbfo01CTpHmQ9W/o76rJyUnnCy1XW0Z4PiloZqGjafLypamOPI8n8IABk
vR3v5Guz1aHtI0GcGjwbTJmcuTigFYqE3AQT8wG9mhkIwGqkwKQVelQlqGVxyTwNH+EreEIjh6fv
topgNlXQ7XxN5cEBIPfLOPo7YDwFUh1Xp66xmD5J/jApVTRGNNwknttqlhk8gB3cevmxlTy3Zx14
7KeggPpdx0cWhEYay37Mh/cJ5oI2PbCTYbBenZYg5pCxkIWM7oDahPYnu+UqiDOKdhMM5OaG5GDj
KdFVXFLVkl5cHKQsjU1tUt9o0hXgztgLkiziOm6H5WMYIRrX3vIi7YEBvrRvsvfcSlgPMIcvZ6VU
+UAemrBD26v2LDcnxDOhaQE3r0HX87byC3qy59ogo4Lm+prOFHgN+2oAbh1ZYR6LaKLqSo+8QOmY
4RDv+Pg4ZzhGMEd4PknWbJ5eWrSBV9EPbZ7NvbtUHoWl1SxuF7yfIVytX49gnwug3FYBkRY1KS1t
uDXesNq26IXoWMU3n18T0aqEQAurjeBY1j68b/OKrUil8cU9GSMjsj1He07W+tOjrPlh1K69lkNc
cpOLDU8/Wrk5fG8szxndLZpM6yeqDN6fHN/V1bEuOGATj1rm9++Si1AbBI7Olmm2ZfW582wUMT5w
l+xgcVhGvTiLT1HGfqx4JvOYwwm7qdEsNmUcjlFf3BzLi5qFks9bx+w1rC8zZ4u9azyaQC17wd41
90E4cqjgVyTjJNfnOfJMELCchuP5QA5ohWfxE9TqEaqNvh6JI5JfAlKv53cjiVTePSl1hXgzzV1G
iOXH/2rogmEyezikyV3n8tFZMdTktV+mDPM8L28bHUtoe2aRFT2Phz4uAcMuT2558Pc9GU0sij08
LFPx5wCbJpQMIO3TJVoiibHkbbGgOe6ba+jBDAnw0DO0U/lraSO8Rkt5N/EO6kuz+i3i/rKyZ1ZV
JinObTEMxfYK+NI7o1ooW6mDc73rh4hiNLJ9zaYXEo7s48qX82AaVPXXe2aDB1gqRnIHwD4ARfE9
a5JdP69g7rtW+t9pP3Yw8K/rCz/ArBnb9isEykIGo9RGT3hes7k2ioJMGOv8xh7pzEuroudEjLbb
TW0Djrio8ohJQcniXtPRf/SRaZcDcelgcb1H8VLB312tkXbqkPMe0i1TgLLr2p2iAikMbK/IFQrC
uxNTXBClZuLUEKg6sIPAfllVGrQWBi+rSR0Vm2X8KZ7p1OLaQ+m3ZkgUampz4bpctE9LfgTWJZWk
wFrt+zfOBTdsc0swyL5V3yuL5vYCLYYcHALChapGTq469YHFSKmtCG6PczlP6+30gXbOMyQ1ZRG+
p53mE3pzMY5DYmlai20CRBhz26TgRKxXlE/Se+7NYqjbqDCyq6ZG5oI7RSdJ1H79fAmxgf3IoiFn
pu+ZFmdzEPemU8fLJUq5Zgc/gF+fhak11AJeaNPdKCpRje8/6hfTrOYXzLyaWyOxYM5J0yYCMyv6
E/uGbVpYZvwYnUp9TCzHm3SkVjjsPFvy/bO+sOtdEX4ZWmZKiHbVpe2D+0JGGYCLfXxm8lh8cqTJ
yav43ka55qdzZVE44Yhtkzfhc2bRgk6A1eBjUTdAQMOZR/aS+eMmOl11ZoYdOkRcda0mRuUNqYvz
qfagnNUZ0ifSSthwsZP6GLXhdC9KoOcM7j0/s0/gAhT4OMaoYQRpmtj00riqvJlrbwMMatmOmoOF
54dz73KHZzta+K5XkMYn3DWvXaVxKpiwJLaTwrLxFM80Echu6zNBq4Dnegh5fpMds2vzfY4egdaC
YBaQkhLwFpni1yWqfPZom+3k3WuR6pxNBFzMuw1ZX8MvOQP77G8JuO1tcdef1V6r1EMSYYHST+s3
cuzmMdpMmNiZdBFuTitBAmKNS8AuYQ3ykoSlLr46428ZOrAMCjzfRQIpMnHkr7Fca9lO06PKHEdG
hFnKQSTKeDX4LE1wKshHCwX5y1bJMpRDCQcyuZjiLo1xaO4PBUJdKKBVgWk92CN7Gp7VWvogVcrl
MadICXTrzFdLwhgo1nUhsTrjtCKrHDpaxnnviM71CaMpRuL8Q256OEhNWXH35G7EjMMN3WJHp2vX
oSkbniyfZIiNcArBbTwDmLF6LpNROO/9dmsHqC58UciFnz6i7Uu440yk3BjCcNQs09klUGnbc/Ix
QFB2XyJxysePd/MmVTh5bSw2W2y/mNBCABScwbNefTrBYFqP0IzSVuznMBbon3g4QFMmyijYtqfb
l/p9jP5faUC3aYXEEOfdN5KD0/FvCYeygajjgJhDzSgC7h/HUUYVkZq3sEaRKxRgRfbI9F12pZX1
EN+1HQNK1+empjFLLCR4fOV8Z8dNlGMD90F9qMlUbQ3PgVaMgW9EgtW8sCAp9nNM9yGe9ayArETw
KaMLRkfQAV517BHN4tut4t9nViEtSnyi/WyDWRrlAha5nzeRPQZZHvpv9V5qx9EeBF9qLOfGf+22
13NG40ea6kg2qXquIZLHpLYLaQ8FrjyPFmgtqcK31XkLm6pAO46Vf7jvPWHd5WUsSsU15QRjWUsh
e/Bh/BVHen1IBee0zwQ3V472lkJlUL+4JcOt71yFgBhD6vMEr1HVVGZbCN6XDqSvtX10r09TQ2ZC
17mYFsMmEeLV3zesqiXKxU2zqJMoaLVKEyBnrKsMViZn+OzKD+O3wGStVo438/flKUbvURXDWwtq
8D0tXY87/gS0XQ6B9EVLLqSb1Iy4BPcS3ZWqyez6LTZucXtuY8IlcTz/kOBbjoMw8r/8e6aTqyjN
UfKyeuDx+KYBKT1SZka8Ps/j5sXsTfZRLucbbBPcx6neJIS14j6we9lKdaQKy997BSi8C8OpU3c+
FfRRwQxr2odHuF2n/nDY0I4vQMnFiwbACU4htuZG1NyTZeSQDPXmsiZvMqAYfJ3INpKFvBM1tzTH
o7nBpSVfZFJU7CmtuL6abB4lO9YwM69zanRacEPYFHUWYUdYnGBa0OkTxPypeCecs0NYd5byPXbK
ZvM546fgl+GuFfc4TiNW1c/cSbUN5cs6iAjVBqTqCtj4VkMCuEErO4DiRTsrWqPC+mKoDy42+s3a
jsuxI7Y8Zp6PMczyArCEgYoU5nLCN+/viUSSN3K7uKuhbjJ52r+GRKcCUkE2k1yqEprfh0ySQ88+
+4rxINRBcakHkDB1MNe7bLaGwoLnpvK1XlT+ewDAT6iPw4tUoPS2ttmmtYL64Q6BccaMEZaXeCrM
fO7c/Z3OZVIM81a2HVFRRHsuE32nsqsOBFYX0j1VAX8q0+nJiiN2cQT1mKV1s5qSoi6sXG8iygzk
a+A/60rg6cmLVh6fIOAuCZlIsnd58Rdrw8rid/ercOEFP/3Ycq9NxZNKSVfiZcv7Y+INX0nUNDUt
WK7a6XClzJVTXGycOOfPImbIvvXdN6SCPFWaSNgiOF8aq0bcDHFTb8Gc03KYTk1wY5d2p6LJ1Mus
CwBLHyGnr4JYM2ZoDrS9D6iXWI9b8SPGKZF4lbBc0P+0vVSP7nHG5ERzhkDLv2cTRCHiP6L8tuJB
aNgHn4sMJxrN19tE0HeJBkLhZ43bUP7RwXiJE9YNk365+vuVbYA9N6NfVX+uD0jgMgoqN/UkpqF3
03694tvGmMiSzfwkgiT4I/YUP+8kt1QVbfoGIhkfvYEpKQBfWltsXqg1Oq2ATyGtVLvpteerJbwS
WwBfuaWBnQcW6B+zqng3rnHxNTteondULGtCBe5Clw2hYT4bENUF9B1T11d0MJYWfcnV4czQlTkd
SWRqSoCt2+orq43ARdcStG6sl0xuo18U3PpYTMzANBPUVbK5HpqwieeFrslVHrxcxIUEFMzJJNdj
7gWVQrG9wpEz6mvVT5zWkVNYoQBb7d2bC0JCdfqXDhlsvMWxtRRvVPv3lnhWUSlQfZfJx4wyAFM7
nxXzmM+ZwDMWCOIVg1hsMOBUT4//whQqujBPW9faEeex5CfwPv4I2f2ggxIuX/6Sny+nbDVBjWBe
X2W12RNktRpTPl2jZXzKMLN7x9wZsE/K0E6XSr5OD23p/01ly/y0bDcdSvsye74xL7aMGVvq25b3
6cVFvR/LHj/BeR4tDy6OFy/cJnwtgxljF24/brZblsD68uQzdIDAXbQ1FJqtAI3gBUZNOzGb2oya
0jLgiyhgJVOa9yjIG73ybFaO/9IVsjZZy1l543ZBrX0CPNYiT3QD82U0T+EUJ8vPemSMjOU1pow6
hFL1LgnbkFXn4BOjlCIjGSS1Uf83BbpXtVTcQL/NEt5KCwuzyf5GZy+3ZoMAkVM7kzDn3MHiJ+dH
bL525/iOO5jPk3w9HMn6OUYnGtQ8aHKtD7O2i+zaOgSOpvZ31+po7+8GrV90MqdpGuYf3CNpfaaV
mFKYgi8RQ9JtxTem20EuKhWZA7D2DwVJt0oQ+b3GKTK9aAOtTfWkk6FQar2mj2iab4l0F8loIdLE
7p+flXEyBTI+rg4rRVg2elb4OEDVRFBwguRtOgfLbLHsmi8jrUgiXpwFXOYaCb++TExkJBFlMzIy
fo68OGVrcZnlSsNAW4jmmdadTr1CErTVopo4+3zaqaSfedDOWNxF8eWDux24Ah0QF4PvhoPIKHRX
ew/zbD0kBGPPJGQdRyzuWRUtPnBWyjzSPFjn4bXy+XFiIlF0ryXRjMtyrk/fQYV5NVaRafMWtAE3
i1a9S+7V96oxcfQ8o9qYYDvbZsI+dsp7QPzIUi4ogXvk2xkGf+o1YewpDyOTpnuqkXhNGVRpE8Ys
G4sA1ZbNyRGsWtHvqJKVQRtAlhFnkvp4meP0i4xuV80eXYy991//KMrCSLC3tCvxGbg76+Yc/6l3
T9aBq3TnnJu+KuUF4+pRs4M+hTOrpLsb1UK8UUYv386E5qG0hHFje18wYBm7zEWCHaUrUajPEKuy
Hzv2bT7dbqgFm3W8S4KfuKC0eJgQRBJqaeJaJMwjm4DGS9cc5MxsZlBhDYGcrjiwb1/TTbl9XITq
OlivYezUAjvGc3+VYfZuNA7PLjXEFEiK24jdGg9z5lrkDU1/fRvZai0FoRmUmBAPwI3BAKKfSFnS
9Aob8KoJNmoOxZ/aR3eq/TChK3TBRil9gA01NocQg4crVdXVEIAkAKw1JmONs1jk1R4LeBRcIyOC
+jEVGWs7A9F00G1Ms9Zk4GyLb1+5+5m0rcS21GKh9iVsqbonml2L8lszevpwQ1lYXTb0NI2EAhoG
1bS5a0FGm+oSxaL6R9ZCV8SLyLDImIywdBG/mmQv5vP+SPUVHg0BtDCF5LTAtVWzTLLsu4oO8VjL
RGdv/pw057n//Af8Gl99dPORlPvHW7OZI0B45/9aeEcwcXcIQbtegRZRxMe5CS/gKAOVI+w9eHdU
Yni0jxEuhS/wQuTQRYWdlSMJ4LaL3/C88yna/h9Fw9IPYE26x6NPeWVlvvJ7nlbnSzyLirHowEx2
9tqxinaXDVAtxYtwqnVcAqGjE3FShvEXPYcPDd1rBE0iWfBfGKUQ/sXakVtPboQZNZQWyXlFYNkk
XFFZ+3DOeZz7IHwaCFWBfH/mIGHJxp7TfW4aqA3uLnd9qiCKaklUmOgKP5jvqkg6mjr0jHtLN00m
1M4GugH/GUGh6glE3PoZ5X4BS6DZUych821RV/NohGj3UGbCfNtQ9LSqgQ/l1dru6vcxsAQDe9S6
stxUwTOp2krfpqBagNRUf+5lPd/YvL9EZy6tLhRr627W28g4KeYqG5qH926QazuHGdDQybXiOQ7H
LDhhAj4iUyrwj9sJoTV2s1cXn4ohuRGpFWgb/K2x9LDuxDlvKDcU8atQFgUiVSI4H+73s0djxQdX
uSoUpKzkWrLgSmcMhG9mZa/SHJKQtt+Ut8WDQIUgexFMWlvZdSUkLSIukS+SPKYoZjpz7NMEnJ94
/s8MMV8EjboMDcSSV0xeeeX4u/F+MWmGVYaHh0KleQVT39VcNtSbGdhiLI3+jM+cD33/PaOA1c7a
s3dyfSB98gVD+oFbouxXKDDWPpNTQSdX5NGrJEelfTSvihSX3n6xMkEjmkRXPzFFArV6rob7qZFq
4RtZmtBrF0/LMn015uUvX+8MK/ipZc6Few+wg13YYaZg5Q86luXjvg2LiDKFXz3eRT5XBAt7rI6w
TUxFf1wMw/0axZ5UBiLCgxT44fmRw0vLGEi+m79/YWAgpcFCQ2CUmrWx0va+jvKx0tZELTwVsTIp
kvXDu613+o5x/8own5f0UJ4RblITG9mYtwu4G9TTn1mr8Y8Ian6uNlG6Fn+Quk8OcWtcrMifRAA8
c0yfCL0CW+iDpjH9GI9zdfxzM3estMbx8Eb3ZHLKOxiM7dabZoPHQ6ed+m/kMjrdglskcRIsCkLY
6EEzc/t42tziBzEPBBBPZuR/NfnG9TV8pCFG8YQwyJK27/KBsRQtKNUHexJ49gxlOq7pwQaUqZoz
bpmSvMy2X5hlv5CjcCFMFt2ATsqfP8W1+pEYisxdjinAKA6qD4mAeD+yLnyMoPFipWjZwCuGjBD3
FDJTeyEIV5DvoV6SDivoFeap2GvGwEFz5GqMF/OYpMgyh4yx1hhkV9LrLw6Wv7/Z1TZSuMCl0/1r
feX96xghExAPKrsMrxARpj7sFohBkKU1wevGnLYX9guPR22LxCXmaxg7qSdYLcfgmhpiofPuuAqt
Mk3C3D0J92pZ9ezdHuZPxJGlqVN8f2pvckta/c5Iw0PYgsb0tfid6tjr/6ht142lMzeKp+A9jlYh
Wx3rAGqnTEjl3o0YMiDoPXfbcDW1HOCRjtBSxn67P3XZDG4/3suVQpblip7RCOy35uO/8A6fKVt7
Z4qGiXg3yRTP5ojjCiemL60kz4xq7XAPoTgpjxXZmVCCFSGOV2D835BXVzG8RGJCO+kcDwNTHTg6
MRrnMHACHpOuQiT/HCunkuqPvlQnfoEjJK4chFE7lYEo8EVWYZ2kv7bxgVNEsY27n+0V47NwrH+O
lvT0SJY9f43b3Ueq6ynGazKLjTn+BCQNOOSXwwMHvioPgGHG1dBfR0KO9zFOz22STDbvt/4M26nF
XaZ6vLT/QsqY6speR3H6ilsYREs5KfeNZrK1OB32TjljfJ003lKbbn+OfUGvJFWVCACtNXENBK3u
jTNWr8VnXblckP8hmADxjkfaokn9UWOH1Aoj2kVs1sKJWzPeguvojvohd6YVRAL1FF+BcjMYEULI
0ASzTcM/hk8LElEhmFxVaCXqKA20N0fDT4CdN+9+83UqBO6y0OQOeiLVt7oxCHABxNCT8ZIeA5Yk
cxlTArqrzENlYqdQFjP8K9gcNNk6HXBycDQ1fiH1PJdp3Z2hGAN0Xf9szKa0OnP/DzfXpeV4icgl
+PECLhTQCo9JOgTTTBnoDjKy2gkVS2TfdW4EbgFx1IEec5cjHbChb8mKiUNGjj40b7uiVn/wGjHr
1r9BqO6VgvSRYXnKXiQYFbbZQ6eh7OolxIe2uIPV3ITR9aO1F1i0KL0Xrkwt7YDUuNQZxM+MRCQp
BCFJa+yhdXbA9RpzUUOLKMkSlTSKIr3mi9uOlfS5SuETBDX+acuieRF2gEdwlGVcPxF5b7HgorfF
HNu91JYOHMOLZm1qT5D7sHR4yN3ta3h3RLZmhb7Db4O4wZf5K5WC7//fH3gjp57ReaJPJ0xphNDv
hNltV3yxEI4OE9eia7SyGIIGvar/ODrxN5c3+mzVKLeP+CgSpgzu9w7PgZitY6m7xR6DF0iAur54
lNqJcduf1PWpIbNyDm/q7b7KO68ZBDYiFruQGtduzcJTyHwnqWJkKmmYr4lUNhS7GJZE+WA2KTcj
wtPgtmDeRhiKoxWP2pE2rWk5qO+zbqq5Cgn8/Ujy6WzxzNTt5vx5RFjfCNDqQWrPSzZu8UocNc1B
jdQ2zSW2zlNPwOBRJC1scGYx0wGSKsZcoG2EwJZMgWReO5hmiyC6ReW3gNB/0hVQ1BrQvxhX3sN5
+utulmYZtHMAhp9DI6gaNqpp8Hr6r41VvDjC5Z2SRcQeV7t6ORKRaSpckLVZaHtu5/SLxkIET/rm
ysB1WQEWQkqXm5u60Zw5NmQFwTtpeYtAvQ1Ur87TvsMOssYFrr53ZAkskTWXnWpPGshtzLiuLtHO
HHvhaCeY+gdSP5eFJQP6LmFJFv/o4rsFmo5sXaQvYs0fqczFG+dvCTLHduxOiArhXIzykhuyUg0k
S6H1yy0K45kPrJ2bzk2SeS4RYWgvBsQ5bzMnpnTtbQ9CjPpbz2XlP2bAPifNQD8rShVGecl64vGu
DxC0gmUtGCl1TVktrog3XjFjceZH2CcumUfY1tcJS4c1pr8F2tiCStUBcPDeC2hr7JIO7oz/IKsN
1il8raEAGSilnEGjFMmGcbmaaX8wLJLEVLfRy5Ojz7mWZ5OFBE/pCoEBJ/15eNb8lryND3J+froY
17Z/c1VJNQTvLtbSdmKacIQLBaH/PNZDNUaX9Pj8ugQS+jyZHUJJBC5innbdKyQwGRn/r2Hfk1wj
jrT1XaZt6LZS/5V9oh4wjCr2mCTBd072IfUl8wFHxi3bOSfkZniypb+QSno5SNXn1KVIzySRnn7H
FG/wMU+VpaoGxOfDEH3eACI1VjoOqeZBg579nVLCQLXJ5iBYmhSRYlRN04Vreyjr6dHYVbIXOM4g
bbLW7PiY4JxTwOGs2T5MxdbQQJC4VvDJ45Z6WALJLyRDMUE4bz1KTkoxYoP4Rcwk4BMATcG+mied
0MHLn06L2MF2j/voj4ZNScPjjnzSNzYeaEO8kjOWaYI5p5GYwAcoupk+DEhlrosOkzhRFwiHYrFk
/fBpw7dI/vg0wa6Lfj/dMCBeeOTZfnXklnzbx0UHAEN2fbBN/s5Alr74FogedbanHpK2cqV9C1GJ
j5GL26GBLG3REhusDYBjUBD8pV2Qbs8/fQyQQPqloAXfnx0GdfgWLSHYktRvISv3BL6f77TAz6hV
t7nUSJqZVo5BSdquY5/NFfb1AEgB5h/pqYbwBQG39IWQ7/r3LCdIivs3tv5QO741RJMXWyQW7GXi
55YnAIGnu2w26n3oilo6Bo76SKLDnrrBEFgzAl1HNrkV9FN4AgthPFFyWbzIT9qfhqk8Duxbybif
t1xVHlZz1tp0qGKcSTG5Gxw215s5HVVNeeXSW7HQ/V6IraZsKKWUqvMBA9qNRmXlBmV2C3sIuFmG
jfo0nbwwgznqok4UE6vhHaei7fCUttkI3jAJQ6ySWrLTW0PxpqQ2rTCdLEVtzi1zmEM7Sl/Mlsvf
eOBmIelvg3Lm881Crb4OQwI78+osVuwYACrHB8VuvFNGT6CkJAjakmsrg8jm6k7FBjIJ+LJSWMcO
sOriTLErMpZcBlMYwZLwu+gEQHs3100+3OsIuobfSukNhOr6eyOGhTc1mxrvOBn9gvgvTDZV5FNO
xpmvhiv0XiIz+DVz0toME/n7FtYTFOIdoNdyLsTuapyG/hQYEuFef7nT7Iug8dzG6qHVrH4BCB5U
NofYrI2EFMKgAdgUY43iO71tyBhuSWlDbsxMKGeVF2qM5MNKTq8+/XrVM7MoaIzSWdlGo6DKhYk4
OyG3zNJ3nwJemfAFrYcUDo8hMlq9ARtDZBWonvwzXozKvBpfViZY+WGbZiV8MBHrMvTyE+G9HxH0
DkuAoStowmvjcCv7SpXGlAMhNJfnr4C9Mf3FDrIAsnB+H9IkVOBJvtFrcQCdX0xumdBPZHSkaCv2
KvUZkUrmVGiDGveW/jc2C6k8NNxLy+M6he8jaYlpqMGZ0J4w+9BUScoqYQVqypIi+F1+eFpM4JiL
1P4cvgjGvStxnahlJCNvEkyufNOQCTdPTHqTfGoHdkLo2QNow+WSqZtl9UEcazLN2WjhDJFWN4n9
2YUyJHJI9DJXWch2lK+eCge9FA3jrKWAjWfw7VMShZo2XQosNgNWUUyKqwEJ7NQKPXsZ+Qs/EU+i
uSyLp3+leXjsB1BMWLCTeXtSGgoP3s2Pz8gAMFVxZlDeVu/3Ry6vLdxD2QaRky0BqeDZWN05WFmX
E7fqxN2R30dJ2x6X5RZET6cY8D1OaNvFQ9WkLpnzLFQMDDifW2zsLEDroBH283mCrY20C9zxZjek
8xCmtYeEpExxDGcztTn/ZEbFPUO4Y5inyNogr18lZHfvoDrAzb3rHEhyF5zd8Nmp06FOY9M651jk
RNdTR9yrwKEnFDc0fv3yAu5BMk1JqgH0c9+x+YjfVkUxlfbXOFYDlBUMoggtH9dTcstfXg7C3lLR
TJBlvsqBmu1o6QxcsPYq3/lUI81oEwmcqjiUP8rjmqyu+ftUEO38RqucQw2tOouA5AbEzMhmgNLg
b4g1GQXvye2hJC+8Xo8ZUck812h16W3MZ8Z4jwXrXndUq7zzDE1UchGfmWKNnpF1CJBftv25SQ1f
gq2VX7CvVCThp9CU2bF44aRcMq/+91cTA+Fsl9t/j0Did26ZXKC7ojTOO6VCKZuWe9c4SB1LGt4L
3hsnQiJCNzC7lQc89Ilt2XBhLEImeVioPcTpSs4KxL6T4HuuPU0zNBb61kwFtMqPo9DueK8gD7hi
4iNAqfksWorl1TGYxmEErsSEnldyAAIy+MtxrCBNQ+v2PPLRS6LbyNUNBYp7uIsmQn/jczWTl+D8
l2Y61n1/NRuT96VmF1TUIJt31Xs8MUGoh1tqRjykxl2jafblhDaSAOkAGWJEJym25Lof7SidQBYZ
ja8o/9ItD4me/tfooS12gK6aqCMbx6xH3w71eTxoR8helYG6mPs4LPaVSGZTT+t7MI0nKJyCfA5I
fYBDpxhIZ6FTWnF17gRBJxN7AMQruki9vwsayz27+qNun3OQtQfIOmfuvbc8V+4DQ1NqGJakGQWd
TZ8XUIyDubcty9QRvfhuG8y+HIJ3f0m8z546oxoUPOR1/O67dqwAndjSLllO/hxBKZzL1WnA3i1P
oBELNEuV6BNISHT1y9lVZ7Y0yCWwLv314a/kuSfzLXCBIUzMo0BVc5PYdafrlLEWafQ9R3UhG4pb
sFqZV386X8WYsl9aTo5e8LXy0l3UrvOgDJgMmnGqGgtEy51SUWPBwNG16XFpK2xQTrqKaaix1Ixr
U89SLJDfKqK2+buvcXxsHX0B8p70nxC1r+dxrlhFWfEXd9NHyTak0Q9m85CROoZUCiWMLgT06Urg
zFNfGpLU/5yqkTXFmGNDK6A0e0ht5Qcrjzw2knenH6E+cCZDxQHwvR2z3xIKVeEYIuRJV8fHp55O
Ltv+u0/LCZKDLr+3GhZ5AnqU7fWtpHA2gPbLx+HCKdIAsrHNJfp+DHP0c5bMxqk6XTFwyalBX9BL
pg0B7jbOKe8s0rAPR/LcRAFpwEmnRump7WYp/M6KR2Ntr37B8CfGZOC81Z3zjWJMdgxpAuu0Xelx
ikAOlpDLWBHWwIztxlU4ei5qv6tWWKurb0RXUCYylXShgFHr9mIq8U5Nems8tL2Em9oB5LSzy5Q7
bXheG/xO/Mt3BhU3Rqmivn2/s0EQ8qAo22q5aeIXdKp3Phk7CAKDLj2TjkbRvuyEHlyppphnUQkR
A2PZhdOmGXbZzhXK3skYbbgQqwsudpgxXsvLtGxYKVJ6EuznjYOYuiZ3RsqjcdpS4biLm2PPEOcu
ntgJ+E9C4c/2yiUkE4RjVIxzO12dDtf49ZAgnf9ZaySjK09ZnjZ4Nx3iQhB6FS+izKBiOPCIHtgw
zRgeEosXZcU8NvHyVZqbJU5aRVrVRBPK87CmpI6dte+RnM15vSFL3ie2D8EMGEpH1w2FbJpGn9KJ
xUePPKoiNW83u/wxeJJ2nSUvHdfafoqc8eB9LvbTT5BDJJZq4OOo/ByCYCr3UyTOY+XMSMyY6oeY
4F27kKEbuFXl9e8nJQhJxreRj9T6x7/q68lBD+/8kTltXBnPpDsn9DN8iKnXxZO+xm/YqkUxvB52
uTeLrzcD85sh8TSk9Smd0ftv3ET1d93kPpxuuJxqoNvm2auMY8mh32LHBnKEXMeumAtQUlUmSvN0
gY1cimad6IsYN6ILWI5IJdfU+gTchka3XRx/VWC+dmH9QjJhDrh5xbyePDZlGjxCbhNbbRglmND/
AHJZctAzQtjGWWUL1EyzmKL6rhuJikSmqYMjHhVqxDlFqZdci2q6edSoWemcWkQ/Xq0QUKEm+QmE
WpO8EzvdohsYjRYu0iWBolUBP5stJ8OdTh7StpiHemZEimvpyUnroCVZIEaOsk9w7BEbNw6JlUxK
U5aqt1/kUxTxAylQ+pkVxo6lQM7LHx2JQxImT4EN+svFvZiRfEQGtJLPFOGZ67UYOByk9sJTMoxf
1KaRYJC2lqGSFBheaCtUELQao2VyQXbVUSMj44vuktN5E3+fiQmWRtv1vXP6nQe8wFIBg8DaqOCG
uHHjRHEoXLfBBecn7vM+8JuoNV97eJjAxeJeWbFsRtsV7nQjTdHW0wZ9qitA6gYQj69ByaBXtNZd
plUzz/jdD4JRovYLcTOz8sbwOYF3qMqnlly7KCu7XZ0xyTQ6Kri1dXRbNCBXb2ZbvyyZwAks+PZr
fF2OPYLx6HPgsdIY/D2vnTl27S6NYUjxkMfoVjOSklJFd9gVhztwjPeFCYhLWmHBDFa0X7el6Au0
d+UEZSA2dN9ZjGC2/Xk1kiJtjTHraSx668xKlamkEzdSEhRpsu3f3BKZ+hqpUxesyUgBomkrsuSx
S2yOpPKJrydgFVy6ZLOLqm4oZpls9xUepOqseHyzeCY+XpBXb0wIjjQlQTN4SE8LPt7+TljNE7Kl
hGaHiJ+fAlYpewgLV+R2ZZlwcbhv0xqqVMu3jgjtKWoILucYJki8I3066vkftzA/LExQOIe500Lr
jWb3JAw0s8DDzRl52biY3ctBceNaYTcoJ+VP3Akb5hrkypfKmY9TRJNkSOpqsZA4jiTBIxf+kJBc
2tZxGWEF5HL8olBlnFmstuaZz/6+8XA7c6oVH/gJpcIU2Z8pOSrooNAGhzuV80C9T22Esa6ue4DX
hx8Fe+hTKktgRAmhD+Y0w1AmUr7VmQBcVlRsDAfZsW7/OtYvzRccvKhfPvXAf8SZPE+YlFtp29Oh
lROGgg8gCXenQ4Fr5lucyPZdF1ix5Q9PiVWuMdLryQ6QktO0iGcpt35Ve166Zl8HdhjZrl3tL40F
MRa9EWl3PyDsqHWeeDLbLDwFPPR2f8TXNybxxrIFTC2ux3erAoh2ej/Wav+DL9mqUhdBslrxtW+F
DnqCPBp4MH7XUiqZdGimqtB5WeefQMCqfiuh81dPzdGAdu8INcrZOcpQb+ik7Wnno8WUChfal3Y6
DUNCmMEuztLMS7ouQ8wxAVuaJ/4Y2ZNdkc9+Ww8BBNFst4nOtiQ4jVAh3LwqwgVeSXrBJTElXGau
peL6nKZq0pVmjaQ1DUdD+2/YuYXDGZJTp2wFWVR13u1fmqyTl+sg9PEJU/652RifuiQHZlIk/dOS
wEbWOFNB6GWGko4I5Xzi2g5yV/OT3xwmQGX+/9mg05GVzKLwUnj9qa0QmsvpGDMU14x26/F49Fee
XwNav2F/9pidAUlq0sI61jJvX30/DJjykyDKRCEPbHO4s/UXUQxdzQnn9vSOyT0LGRo6/9jHP8R+
vaGJ7Ee+nJwLFWrVxhIOp0BXGgJYzRjAdOzaJ3xL5DxE8dSciqxzHMA/Iuhugqd6NvUQqVNX1DTh
XkUd+UlDUj5eWiAqG15wjN9bNR+PoUMnJ0eaCoJ0eJXwhNYsgpibM1nnys2GHbKG0ida2a273A+J
7+CRLVwCh2IGzh8CNjjcLNPebU1JUOoVRsax2ERVY2d+8saeGx9WJrEqGzDAlkw2RzNAfYFBBx/F
aFtpIWawt/uFUsVd7vZMP9U60MmkpTYeg8ZEEBKlYN3jDaQn75rZJBfNwkgF/AVWqeCTSurvfpUn
HYFJnISbFo2FLfaHa3AKPOPyDSAjLANgwkaks9NJsBw7FobQzrEKErIfZx2WG+RHfm/idU7YE4/g
Zs9ceg8QzpIZXyXpyGXCNkIdoQ628CfzajWEtFald+uIKw7+6MDeLYopkISh8e8vuiE1AY8JqsQY
dd9Yey5e0GN0naLhXDYsFsWKm0DJU4xwmZPznmxdS/pR0Vux4AZcXqpHuCoCBIsIL+50SEY8X2eQ
UDzypnV7yycF8C0ZR7KOam8w+4vw0KgeDrB70a4cd7tNHvhYxQgcB8SWAWVa1vnFp+0zA5VtaHrg
L0xHgh39Bz39fOJILxuTiJuZy5reJlCDYsxFqvOgqH+RPj9VamTHHi6akvw6KMkDPRRvWbxHULBw
qJ3TJICc7ungEfm/U8D+IXExEMV+eOT3wtKeGJrLjBuvEMwd/v60zkjQFBeU5oCY40nfRx7WePdS
7t5osTfMMaicFjwOVvlQJ2RsKgcKips3GpgejHm384z2QOZQGZvXnPKtfNpbKOfYtItu60dYcyCp
MKNdc0VLRfxG7Xg1HukzbmfrEf8eXLCyJz/vyLtDVH7/gL834ED/bLpKZ1XmxVcIHUku5h3LngP8
59FR7fjY+VxeNYiqTG5YD31zbIFUW9A3g5youSN7ZxnmBXeBXEuRBEi45zKaMufXo9J+2NTHqVc8
jLIDRFjjclFP1uiEKhzm508D/+BxjQEAgSD4RmBt4FsM5PfzutpNLUlBtBXJvNvRC0EbjH9ULKTE
BDpLgPLmefSvpyhkBR8DwuBryM3ujQNpGNNip24xs1Svrz+8wwpJAk9oUS89YHmvj5ijNXlcUCmE
ZCZ1qJ0ih3hRIl0HhkkrdON2JKzPoIDzeVBoBGjf7sp6ol24+xBg5McPf2b8I8JeaRLlty+6De9H
z+P5sE5m+ejvVqINbEysqG7erP6TwVTb4FMkJ2kH5b4qDC+CQU7bh2SjgS+JcO/77XPzpMexa7rh
z8GLyC/BZCSyUDSOiBXx47RyCIwhTlV8yu+AIcBzPi6VstA0XTSkvOlsENk+JnQouKjSM7f7DZ/o
mvGcsanUMU2CUAyQx2dShYvTqQQZdisQy6yD52+9DdLrANSuq2v9lZo59B4Mlhl+w9pYYJgRmw1S
ou9b/fQodzZCivvgRbHiyFfuyKG17BzjVRXW4o60lla8eCVpd7TAUGLpBdAWk7aHNCoNnhsqcH+R
KU9QtyQ8pjZc4FdLP3ZHvJhBo71xHUsQIj3LUxzWa88SIEJfs22Ok5SLYerI+HgXSadUibgyCer3
BPaU+ZIOjdmrQV4BY5uDLA23tYzR8zkT5QWfUTsLir0hNBCqLWlRUKLvkSU0Yd0NELNkaDehXDyJ
BsXu7qae4FtfKzgC+PDmEt56IP+J1o0efRfxDEGnXYlB9HV7sYYdpVrE0EKFs66rxTKzXFg4wLQr
4YAhqYQ8hgvsgxAG+BVud7Qr2nycAWNulvluEDNxro58q3wD/nej7SMZbK7lrwVyEDJIwx4Hkvz9
nUmyCUKZydnTSFSWZgmGQHFPg62pWEmHlgWOpsuzV0qMduoZnboV0tN1mQ+xaXj2LSrx4H2Jxw0A
4eyLEU8jvqI34dbraWIKq1udSAVzBMlxWknLx90oCWhL0xl8tPP+4N0BkktXasLNWfWTQFjGeTsL
rNR9EVGc3JwciG0AtK7CFGU2/Ev9ci23HucCfmeJNvQE+MkMMq8tNcs6rX3XUuK5ke4fPsSGS8tF
e+8LrV80mdupx5LGTm5WsxlTS2f9qB6qML6bplcYlp/6eG7BuD6eSeKRM3IJGaQ/RHzgsRNZ6YoO
vVHnH+QpZlUEOVJtRjeLN583rSpoLQpYT1PbkPPzHpXkc1QrNNpFwQzIpMhX/P9WBvpnSBRS7Alq
EMRhaUYLNTlMLUSgoRSuIwpTDbuWaIb5euvQELeflrDVfQGslZuJBiamkNN9JIwXLh292GpcegMa
Dn7AqUEZSKxK4aI9NZBCOOIRY//CSj9ZSgGVHAhk/nhoP7L8Vatz1HmnQEuQRsYP+vGpEW4V68WQ
Y/K7iSNlizenMwG269X38h86SEf/ir4wb1jtxYrAs8Y3KeeJQYazoqmjPQcYNIQW0gVYBGWi6LLe
w/9pSgC65fvv2UAtnwtViIXVXXYwvB9XdG6m0nLjfujJAZ8eo86+AqdHA7DyXTQiRjWcn9CdjFBY
ok04ujyf1/sTXiH0ign5xpoMGN7Vq+xqKh8On2PMsUiyYHwF1i87Y5tztaIiYM8Lx5NLDzDcO/j5
iIr35WvNWunMRt3mgvRblPi7AGFBWAETTnwz1mIVHR2xjsyhf2y2Sy+f1eniiEKMGPdIPfNenFeF
O6UB7u95WNvG6Jh4QjbH9Ucn4RenmuJk2k7re0zj2Imu1BGJa8hMts9faH//xcIl60AbPRwruN9f
TYQFXmi7RW4b99zrh7/Nl33P36Z8s2hNQEMcoLYkiM5Pgoy3rtdrMemYdjFTZR728NwhZS9OwjEB
xeRhlkvcS4pciwfqsoX64UZWVcDzs/EX4knuV1YuxlinLGzMD2Fiq0mnRE3omZsx977YS9PpHF+n
yHD6vBKoze589dZlwj28o7d+Jtb0qM7BQcslm2ku6Qn2s8j1TGptVX3SPRyus7xYZvMZ/op1qaCY
J6nXV1t+7aFpiSvgq3BXwxSb8q1bYFyMIoOu+XSWVbZWZJoYASOORNdTTj20eYNPrrC34F1JuXmP
xxXL2DxXZRhsALBbBS8lJNYUiBO7GwqhWbw+xnafXl3CYrNh8Q9pI8ppQD/qDlpYttZxUYFq0mJI
hdA11fGW8L5JT/WlCTwA35e4jQjMjdzhUrGLrZ3RrqaYbijoVmEOZqxVLeZ5mrgw6PFEtMcgOZbZ
6CpU+GdQ1WFvZ9YSH/Og3CwbK6duCCJThmhwlSuIbIUeE3ithkYG52ZQjfcSW3nhupA6b3k/zeO3
V6UndqCqdTuMvHdytoY/H4JgGKlQrRKYq6s7DdWjUtORyRlw1C1NRzwgIE7i/fdquAGmghcwINjg
rBE25cuSeSdVOfxvuEiDTChSMBquDXFZR6mFQ80/Ql+6EKTzqSJTtkMk+WKpqtWD7B0PQCblNEhY
ofUo1hmOjwfUCILjIxyiG4BejfjH/Rxg50GlqZq2RjRUOg1R96inDZYrxk0cqL6/KKFiprgpR07s
c/SBCZXaGV1GRFyo7+OoXo4QWV21obauUUqSxwtNAWWxVUB5xUXpuu0NTNTSmNlzcSXw+JaJTfJp
4dOSZAoJ1pPEPnSQjCbzIhhabJg1hC0RBvZFLquiVyw4mr6ptuE2zQH5Sf03V1LUEuMwmtFEbqoy
Da5IzdZuASmSGk6gDTzhcbbKV/aeHujt/dZPoi0k3eZsgpc+acGdqTEeDHaWAqBEZgj9QYPGpGhr
0xg7OuCLI0cBfXoXgCeXQjrJjvwnopuV9yMEI+EMc4/G6zSokl+3EPF+fGqlIgJSu4omDulERwNg
18U7VXOksbKgT6GY2tO8gEkrN8OQ3/lgO4yZC8aStBXvSsm6kyz0YiqxMuMerI0NdTI90/75Lk+9
9+JH5h1IPR5cruS6w5EFocJ3ZMB8X0QkRfitCAFy7bnSQEQQH79BOo4GBFjxblautHvE/2WA6qNg
fiTNg2wswVFqS7ItwqkPqyNqljVYR2DFar2lxmRmMtQPP+q2Ygg0/tDVQYtnm6M9iwW4Oo8GC4fL
qG+I2+GwLegUlfSIdOarbJR8M4s60lKW5pGFwnmFDmN3XQT2UaVioxb84cpIvXl2e4YaGLETUAb7
wGRqSgPEHUJMGrhjeOt4d5k01sVR+wZWqQujP/+YcIYytmQFqxc3mw+BjPNht2gDa7fMIk7eJk5q
wBGAH7oayDXh9Jfk1Mxfdhe45TCfcb5yRMkdpLW1NIPKHO0DWnCSK8+GRN+Uuyy7gslRvc6UXqDQ
oiL2xW1q1TYOJn3/fgDGiHuZSMEZWSkSCkGKwkx7AamBoGUiocc3+hh2jWqye4dBfj1zbSmrGMVb
MnQ+XXMi2lxusVMmMAdy+Ru5eaJRew3ReGI6qcnSOqHLkxYi/eLPwOcOv08zA7fhE+gE6yRR2bhf
5dx8j7N54eRMf2tjBxuFBboqrOrHlezGkfAWqMylWmOkJunUzrADSThnXWal1wDKCbfQjJ1ovdAw
lKKJPaWTH/qv3yk+paoYeIw5TWwH9q4ZCgPvycR7dR5GNs9zHwcf94BI0h67rz9RjKBG4QY4lfkb
qeq/VYP2Y4YGbeloM92BLfFg5wT+33mKOJulfytJqwkhHXzIiNV30a8prBhFTjfU1ICodq1mOlH+
IGw8ZfkopCyKXYAMHNTrrwrFjFHyHeof5828sd5PpZ7BJnt/ahc6cWY/l9f4ydEFvjHJotETguHC
jYy7caeNs7UflkBk5M4wfTHPDlVLG6yvKWHjKwARB4KVp0Sx/cpmEUn06TEQmgXMtClwkdEKFgb2
lcsG5DJ7rLDtpfcFg+eqq61U4eHwiP1vLcVkF6/VMAkvhbOEJ0lJoeKbFdP6z2G771eXtulboL+5
tx5KU7mgjKtHMP3VnaUuIVfGwg+2buUDFHNwBmPmoKz0K37SLqHMTgFBrg/cIiyrYHtsuGgXdIUw
rEeGKqepqrYKEIhfv0IMM+/iLA1x5wPcs8EAsuqfdgVcvSiJAIjO4f0qABHQz5tcZR9XeVQKaWfQ
ztac7amEBcGz2h7vSkFCTeG/eYufCjLcYU8V5lt9lML33rIqF8S8kVtwXeTuVnpeRFgNc5FhMmlm
a/12R+GT1ss89l84CxVGxGRaUBTHHIaRPjSyPWP58q4dBw0zVWymt5+LPkb5iPNVkTN87Ll29sLW
oh+yDvBZ3Gf0CaFiDs4y3KcSR4gsNegWikSaXAWLPMkmL2heZLVx+G6XIk1Qb1NWlydF7Ibehc9P
X5w3mSjmYX+svmlUs2YQyDgCTw9s1cT3Jk02zZnJeiOFQ8vWLMFGzWOs5PjRbaP3XKs8H1hcEaiE
oaF4mEod1eyhVZTKQK+oXLiXTG6PugXa1qNXzkJ0XT3u47pggBx4PUrpIz25riv7naDa3vmwvDq6
ei6Cmr7ra4DmCM8mGoefSxW/xsaVcQh/w1AwKbpkoF/8AOz9m9gzfZEbKv8lS+pmoIbMIe8E03LR
34qRZbYeZkV9KOw/l7GFWKMce4mlJ29OGd1K4tEygqcCWjT9hkEWUH/f0FrSr3JY2XF7WMOEE04q
Mr7XvHAn+AAR0vHMUpdqWAO5ysvoemWMXhHxLJUB+1xI2Dwy573IuFpT+QI2PAhDTBkYMq+Qwrjl
T/am0y1pXaPFRZthVPpb6EEtIFs789dHuAka87V3GCeZU/FA1g2IvMuCRrzynILFe5HJzj8MRP6i
TBzT8I20puGo3g8BSz+FAysPLjKyei5pX3Z+T0JxBYgIF8u7o0FEFq6MbAYIoyIOhyi+3mX/ahio
bdbdjVPOjC7Wf0Da71zvn6+Eu5pIdm6+JiRKI5fFORaXXR819iXZ8nnF7ABr9nEaZSH9S34qoRf+
AoMaDmvbdRQHQgVD+ONqt5YpB6liLraQsyRAL8rK8ktjwLpoDk5QoTE6WkzwmuQGedIaoemCeFjf
EG7S95LYmchEdrb6yXojd6q9/W3Fq0PjMQ06LoSHbhwOxa6tRgz0IZmzye8/jZOTsCRJAcGi6zjw
pKt0lfrEDyUXzQuVrG0gRPEzAN/x6jnEclMB4N9/Vf2ZHWT5daAwUAesIvjXnrem6+oWYH3xjcFu
Ryl1a7dH4eRwJCBguqQ8r8X2zSAve5t94bDNnu/Y8/LIhAO/4UUGLshucMPUorDZ1z8KgiaJooHU
tsN6I+nUDZcDFFpWB4Pc5pZJJjqBtwLTRn17bmOPl7141ScGcTXTKolGE0uDTuIXv6rYWkcJZDHT
xtrZ9pG28I/qnZ0RlQP5yvWkuENmDs8RNJPpfAiqNuAVYN4wX+1fwQVLyLwG+EHdE3yKtuvR6SHO
SIGmKmxJfeSkOCS9gLRTP6D0ibat2pKKJQuTMji7A7M3YhZRflhXdhnq0JnpvNCgj4Z61nlPhFwX
Xjpfw5GmVHj3wnRn5PLXdMuTHWKvnxCs/D5ZUMovXBePYMNKmk4HS2+DwUfIMNWMDuk/BTyrDxNG
hm5pO4XLqpPbt+w2+0AgjJybgm51lS2IQLNY1bx15A2LQpzDWiaIt9vXOvKrn4TwIl411JzN5DRd
X5oDYap1UxjCTA3X0bQTxYPkaFk+sBPpcbGw2/g0NghsU8HMpzQYDo5MLd2TW3jW1zcKUX/i3OOF
nZvFUrOhnr2rbcOCg+g8AQKwWDdOAtisnd1f8tovHINkHdXAdH5jpodDvGh7Qz7D0RzjKFNxGI+k
H6WRFZSObqgwoZLT8bcdxhwE5pIkjVib01Uo6lGuCzXRzWCbRju2SfIifo7o4SfNxZbCSZGvYXmf
ymkhCtyzUOryKNF+iYe3Sas8A4MszPgkZDHNU1FdB7ppB5xcvCtf1yVBozmfeVaPhVWy26PL25Rh
9QBHcpnh7MlIxjN05yxcbNFYohpY1kHD/ErVHRjFmP9ZIYKTTnJ7Vuhf2YVs+HqCZI2znVENd5ZU
GS4U9ec5kTDAPNRPnXZUrZR8y1CXGeOSopek/Sm4D7CCTE+mOm00vUsXTGyO+lTF/fEqVHXSdg2K
ASnCllKZoyQWorTgFzYlRiWWynZp2pjrLIwozcZfZy0uWnyDGguccfWKCnA3vEGmvKKX7fUAHbsD
zfJRTwrjo0SsVsCAiWWYjuKEAiGFD+zB+pzgFqZKDepHeC20RPg7sfXZSZuE8SF/8kZxUPUP1XKi
YmsmMkvvdDD9VAvfgupm8n3s75/0z3s2qL/fx4osT3x+L9rHXAO0I+lMHojcmxPaXf2Zxi5irMrf
fVK1EWPgZBo9ABP45dAj2+rleqW7dz6FB4oxvgzg+8IsnJgKctcb8ErjhcvL5c/dKP+dEsjhtD3J
XRr42RytLIvRcv7P67+/lyibp6CSy09yvq8r2WYKGdiDpzauurwPusU9MQiiAzpANQiZH0q4O5Ek
5F05TuMdycijuToYhDB6sI9C5/nYbm9mVFGVTPNSg6y6vwCyWVvbuRi/RsOxaIGeS5lT/OTmAoW9
tf024zz9S+SWHbCwGRxmCEp9Si01tZ6HHI9YKhXdQDUcZD+2AxFsaQApNdrHnqJq/rV38etYB/3G
JzdjznmzrPI6cHZSjBkr997hqtxa6c2xGQodluUWb5/o4fk6eJpuTqmrUVuSMJnWfpvV+SbKtEhy
Vic82PU64xVoRmFPJYrnynnMRqhig2EyhAZ7uorPdxL0JJAmrZACeK2cnUE1pCu61gJ+3Kuung0Z
/T64Xm9g4izb976NZcaYCykD/ToWW9IkOvMAZc5HjhtryQvRvMp9xyVirMpXJQ3exysnzn/yWqR+
s2yFUo3Xv+lPG/BA6zPkn2OFI/KuHgomxUBj3u8xUJ0xFzsZ4n3ncuWQtSbZeDTx/w3xAafc4vge
3s5VIjnMiHjOHKERQaObkHjmTL/Q1hV9EAwl+ZgwB+ImWLMB3+L5Ef/Xd0wo1+Gt0vxyT2zwg6lO
gkhexnrbUFjqaRPLi5WLv6s1aRqmZW/c7Z5OdfyhtMFlxc1ht3cheKGoqzVr51W14H0kAi7D+HvJ
8tBKQe1xXfd72M67qFVfllwBxEuASGNGTPSYbk7YpkloIbF1laN4LqChUdOUvHno/Y8r/E+hC+hI
7QM2ujWHCHMd+qVKyBoQtLZYRQUiOu9kMyzQzv/tuzBA23geWHKrdjknugXpu7tb+yWVUeErDX53
Daq2sjjZLggdrRbnSKnEvZVYiT0btAcsNaka8qUmtmbt14fEEW0qrrPdjg53B6Zlzf24WQz74cuU
anN+p2134ep0p389UoDFSkfZdy6/uNo0jvrmT6aMkDikMeYF9uuOvi1NkhTABdRTHPVfbMlRj3Es
4hdrNJ3aiKS9bk1TQHfq5W0iyjuAjEWPmYUQHCZSqed+tm+PMRnSWA2uak0nc8gDG3Qn3iNa3zba
+HtBzLTlivHZTMpxXhUzbelfTf6ID+FKM5xWVHZnc6c845+CkIhiaVv6ka9wEEYMeW1RXnz4XsPJ
jlsYaaS6YlL8Qs7Y/UrTMah/8Cn/J570AycItedKFVw1dAgJc9PcFm1oJmNQJS7B4YQ3QdjksLwt
4NxgpZ3DbHsYfF9qScZIVfoNyvmykX2/d6hv7QcqcfBiNTtHRTazVD9h1UFMKk2Hbm1tV24/iMSa
QhP+CwEEmQHQkQIasUFZAqq8SLrDI7UX4pzuMi0CP4J0gYaTTWX8nMXK6nIucawrBICQZQQmyn4r
mkMytbX3S2OAE7PY0Ifp8JNYAJFa8UvpLxuAlM7LL11woy68aAs1z+8MApzgytexmf7DxfITMW9B
McNe92tknq2GfWqbfjNUTXrlexQYwp5f6qu4oSaoY+yi+GM4tiVrgXkrwXOH99PBNJZxAaDlBz+y
dClHPmWYsLcfGEC9ZH4PnI4gLkYke/n2u0+LfH6aT8AefQf83ZJ0eeylxj52gYQdHfmVI9zVwGap
jTh1ZaqeQN37uoEZTctMs0v7xs400VuF4cGGZKeDQK4Lb+U/PHJ5dUBvHQcNpPFNI5jfYHTLo2LZ
LwkkXHqm99gVe7O8KEDpffXdhki1UzGgA7HOCIenk9NB1XUMPRshBs6Uv6lbutg/9mzUm0DmQtwb
K6Layu5xogE0IcZ8n+saQ9mCUg7wBp9eJ4BCQl2xT61hB922aQhtza7u5/ArlFwiB9IEjcGdfH0O
pFzL/mYWuVaZrhRtBiRn/HQ1z/lsjxof9DOcECaHSVe+br3EKDWLtdSNoAWga/sh3S6j9fPVpQIK
N1nxCkL/qnPpl2VzBNvDi2FW3V2DDMjCSqJ3oMO0/QiZ4KyoMvOGODRVcGotHgwNfM/M+CC4S3Zy
DuGsofNAkIkwbUT5CpN/RxmCgELtBqN5zu/RiOUkwdHW2UIlDSP2FG9BS0Lxm4KS9j4JIVcNCPkY
4ik/erNnEfqKCmiuJukfaitsYFdAgfNz2JW60KhJz1x6Nlai7E1D6IBMW3cfgsCCOSqONRrddDZv
0zSVRiZQtka955ijV5MuKzg3hH4rt1zuXDjmAgCuChB4yMLqTfyMN9lj6MYipkBpACtz2t2sM/Tf
GJuqYOpxE/rFzkJRyz6MHZ9GPUsmq1ZMe8YJuiVSgbiEXQD2OroKWI1MvP0xE7RlhdSXWB1uhL1/
HgJKPa2lid07PBLG2tF8t3bmzl5VILxY8BbcSIopbJ4bXB8tG4hZfgvYlznaXAjo+/VtAd15rYWO
OUoETLK2VJyGp+XCrNj80gEedMn+y9krnBzEDhgVNjTEhX3bvxhOTd6qolOlwc6IKCRBxNOddZ8X
yI1EJ6+40NRX6UVYnOVl/5qWp9BVL5+73hcF6bi47wcmVlhUVY/p3iyFSEIbf201H+gECd2v3Prc
rVVxgzrM/OEIEVt29R6AfwZb+4xVZ/AEx0xHZiqA/L6MQtWwxOCTckjm7x9Ulx0TynuN3MIMbJIG
z19zwEqyGRNmJccXb91W3AULte2uE+m78Eh25TqBAdfMrc/+OEoI+f+6YgQw75+5eX9fbj7KD3l5
gDiASKWWIx3ilVysoV8mE7ITjLeyHKURn9MhkxKbFId/TMTKhsZxDPLho6Sd/FlmvEJdp8qzAYqS
swYYxJhLD7mR2MDBEZ+w0AXDSzH696uZD6fwafdmY9W234Vla1trQDltfD1pv7Z1MuPNGan4s07G
vNt7ubrOnYODBwOgAG+AZmlDL8OxXAwm9rD0WIBtCJw0SMnQLPautaOqkjLE+bL3/ejBHh17NaJC
rbPvGwRw44lvub5/oUIkegU6QmsE2jDqN/dgE+D6Whz2p48MDQAEiRF2+CCbiLItRCbUDJjfKOhy
WIUnXkXoQsaNSzdDYIcJoK7yOv6OJSW/lPqlqbLueo9EZTME+BHMfhACuC3oh4bDSfdFefutkpLa
UG1SJo3SMqyMqwMIm4YNk+maaXNtQV3cqjYW/2LNOeRoCArmwXNC30p/ZclcFIj8NIPg3kEjUmch
GarU7rro92XugYagCmpC7pNIGi9VvH9B94uYcOw7ovLcKJO+Xvvitlwg4A4NpIrXS2aJ362spV1s
Qr2c8A/0tLfG7XnQIwifNAQiUpMKu1V+1rWUBAafNivH0ij9kXcRfxB5LIBdJF0fJA3qjukB11en
j1FBENCDA32p7x8uZ7SSdcnJPlxaazE8KbMMtp5aZSEgD3HbQSK6FzgOsMD5Ep7DBCMWHPaPqcoL
+x5KtfM+DXLTCyp3n+PnDMiWz6bRbqeS2jwtBf1QdqDW7H3yAZUiRhlC8RzjJFJYL/VI0fAD7goh
6V0thlxkHGErFYgdukWBL6OcZeO05YDOOIXYPU6F5th1UUUEprbIF5ZzRemYhoop+3y+c8v1eSOc
Q49kyF5e92hXqeJi/PR+FOZj46qBSzKFoI82a4iIkr24tDcx8B7aktdl+RXlimHXjfRL1NthGnfQ
58aDZqXD1kBamlPzJWtz5h1brCjuDeYNk9uZ1x5rexcLpTdhizmwekrCRfItd7AnP3vVBztWXchv
V28CwqviyRCYzsa6UVpBJYvYd/iS84MN6GAKt0hBDQlnCQvCAVi7UkH79G65rLboQhNYNtBH/3ru
6YQRawcphw/ZDTFD3JhA1KbWbzP0JB6JCGG1M0ode/zgbshe9wvm0ATso3A8ZK+jvpwTIQFSMGuZ
COxK5iS70qXUSl8pLovlpZYdVT3utpU7556n7r02BuX0MD/IMdx7w4Cjd5eyLwWoqfC5MhhAhPq/
XN8P5c+11Rtu5RaYHjlKc5vhAL5Q9yxw1m5QSxg10MompfLtTG/1EvTuslRRRtbuPfAAzoAL18iC
nVRDsN031sSAp73Rl7Nea3S4ceVnVu7WQfASTv7d17KDR5+m2cX+lq4/5lyDWG8JCWjP44fPB3i1
wfKoHOUUH2vQDmQsgaXWMBmSuzq9gUBlCb5dZ47oARDOoB7+vSeKTnF8/mHxKu0ZFn14cqNWI6LL
Xlrg8XLCEfrFd0WvPjtTSlelc2kHS1lwGr+ySuEegVjX2Y2YddqyZE8L7AwgAA2UF6J7ikcp26QW
D8SBydTrr2owUwuOjKOq94Z7ebgcShvpIxu8/mUGIdv/V5jXbpmsPyRhbP7aldRKEYXcl9vAyJWo
YMVHyUkKeBW//rcF+ukm6wh5o4spU0Km7ZtnKLyMVo+GMcWVN4kSzmoHkqmwuJl9WtWB7ZQ7jpWZ
hZDgMXFJWIp2upYHmdBTO4aS5J/SD7y9BSxdGph+U5Gy+XL0JfM6vFXezsQj7rkDQ3wl+ujtsJBu
VX7igX6GeC2Kaf/eEhrXsrXAzd2SWgCUP4keVKbUrxGp2oluo9W9+6o9FYCP1tGh/HFkugO3q250
VTGuZlP11hm8uivWla+xW2wjqZicsbG6c494lJ9tMjeGWiEaQl+dao2AVgyeT60w+SnQgVA/OKa4
hb5C8p3ZVXEdWp8dmfsSSUyJZpoj89JDu/6N0RX03mfPPRLGijs28dbJPHLH+spO2Diyx3TDV0Zz
o0V/rb21Icn/Elb7WC/avPUZz7X2uFVsTjXanT0rwfMpWmCek8BDv1ziL+uBRXauG4e9+gPEEeUf
A2TbPq0gdKLKoP6VJC9N5hOocA/aGtfpxd2MEmMeH2Y4cY5DfE5faYBI+dNzc+lLjeH4sk4zsFmG
KHkXymtjNVl6JS07dI0k8+ADKIY3gGUstCxiiEjeqAZsFm3Ku0BflslAWjpKnGOi3ffaSG16F9aM
yZp0pP8TxJI64krGV/K29HJ5cAHZ94xWMCnj00Uvu5VPUfgS4WBAsv+k84p8EzCMefkk5N/MBoLl
RmWaGKlkkTZgeSNpcaFfDHWAcEBA2UHJJyS3+IGglXrlmPe6zXw/B4NTOCeQZv06yipWjkZKiDvh
oX3UbONvYBMIJyiFtJWvkT7KzlGqLlxrBNCWsBj0r9BYVZTHjO4H0N2A6qF+TTkoas1bv88lH2zr
A+VGdQCsXToZmadSSAzl9xtu70gxrjcuWsK9SDnKmdCG6T2rOOh8OzNNNCfFrWAjpH8DhVG1pzFv
8I70y4B1f5NUmPr3xn9UVYT0r+JR3bHkLBCw0ALiq58cATWPFrmseWdZ66LPXNoIYWhQzu2tF+Vh
5UiNSI541epSL2fXPvl3nKuPVybYqQKkNGzZth8031sfNwYK1LRZ1Grcm/e/raqyNWbQbfR8+2v2
55612YXsRjg9wztgB1SJSFxk8vhZKlzusOa6huUuU0wmgtwNDp073MGyEQcT9EKw7JhUt4KZhLWe
iMBC2gGWx9YETLhYba3UB/SKO10N5hjmRJLRN0xIpTTzEBfquoaDdMbab9SF/zZPPBUB+MZ2VLEB
kmbjhUMHBuYl0lH4odqQ/owxx2qJDMf2h2YiT5gYS43zutsHMsHfHaWjaoe1xtMJewgnSpCmCYPz
uEP4N4dcEICOy/92bFQV9/PcSrMZPjcXDHCsGAlmZqWBuw6jFbyJL29aEJIODNPXMmzQw1zB2CPp
S0OMN+Zgz5Ki3WM914/fYQ6z0MlV4tkQ6fRTmOQCMh6TDdKrmHpNVVuFkyNcx/ei9taypmXSezFP
Ts2zLFoIB6Ff5XiawY2ml6vr/zUm8f+/+EV1BUQ3rrysm3j33AkIeqkf/EQWtPl/lXkYBuIJ09Uz
i/r3WKVlsG8Bxts05hTzkG7O9k5FWj/7i05nSr8sEdYyeG7Biy3OVMsPU5EhWK/NH6McfAjafwAB
GaxCZW0k3adYHcZq5vI32N+LzS+cFFDvROSpguvW4+EJb621WYEDgmJKkh8bibCe4qHKzTmkZuXH
GKfJnUQ2GNV4r+gN0qOlCZ1/lm17HRi5ZS95hiOoOvZ2CUiaL0BYxlK/RtZtwmL8dts4TFzgOUoS
2VtfK1Z2julKs94xT/oSAZx4Uga7xAwMxmVlD+13S+csOl2W8YzPyY355OVaAFMfUKZlw0FlwLjY
UEF/LUzZVPBcyLBGfGTMwB22A9P/ZwEgdsbc832jOfvDYX+QAd3YaKxgZ5oIyMgAAXoqGRi8UXiL
agCiSm7KrAdee91yqs3LWuZqGuQxplAAuQka56Hdb2MoDryA7ncKYQ0tx1JBoLFd74Yjc4pScWyK
EcgAD/Kdt7KHCN8xD4XpzZ8ykdynn5vup+16a8r0wMsKZpxbelX0NMjHjoGGYOBOXoQldQ9mWizs
qpAiRXkxDfu4iXag6q56w9lRUJ7+TgHoN020j7qUJ0p6+IUYkCHKee1NR6pvm5pNyMoOxTbj5q3/
FN47ROylewinVySg/7A8PMzp9OF2MGKHS+GxjAjs0KqYBQ72FX0ysj/S6G6IEyQIgjhELPPbKI6k
HCTiRDYMRuX8Du5Qkn/ce1QKkwoL8B3OUpjf7CvVRYUp+F7Ne6lRkPlLA5FT3JinS6fRgbtEMKbG
mgkmSk/YHajsfJ8Ku73TYAVAX9kY67v210isaxDxWMtbxS/NgctpgktLLEzUGCkVDibcLqKtPbzf
u2xsseu2RCaVVUOyiUxpB6tvKg2PjG+Ky5tXdjfTBVpHupAVWKZUq7Hb06duvf+0RHiNYrhMDBOK
z8sWPXYcIierjPyCDbjcBk2Jr+6gcXm7khe9B0sTC21nVqmpHehPVTnHzCVw8Yzc+SENh02Mqxud
wy2mZmmaRC4a1pGvFee46sU5RBXO6JHzODsrqIZT5gqQoAKX93kfKj1rrHpKjZMjkoc3mql5ofxr
orMNjLZUC0CxOjuWg5/BStsSKhdk77Au62xeJRKjGimymSV1m2LLdkpeSC8d86/QVy6hHDtbx85H
fL881a9SR3rHsu+1v0b+CPVmsVEbWvcrI4nhlzzXTpRNFzg90yTblUDy40uSUiE5sXBPWlaJ53KP
Ny/IPAJdii0VtNC8LI6zcHaxLE8RVTQdayreE9qpAWNlXpN4dO9ZZ1gxEdKxyof/MYSakg8nVm6j
b0X7xeNlA+m0taOXusg/8zmJ2Ppf/mkOv0B7HjcERzv8mNcG0ho2tSlCWHqOWmr5QXO0h5JQjroh
h8TnoXdzbSF4vKbIxJM188jnhnHytqpCEKaqBlF1ELhMMBYUdVtJatUDr2TJliGmWeUMBaNAao/g
PenZWR4aE+V8zgnBLhI/KU21s6lsyFqg5+iRBGxrhrOesm/JvOnt2TND51PcR5D0golQ3sLKFO3Z
5F2q7lp2cDTYbiompF7XadbH3o7nHutDNs3CqHvM1s5fqphBvXA84sh17keu5dxAqvCnNGTsDsQL
+2L3VcsNA/ot9xjgJs2yOmpj4bsYrPOaUn7wLiHVMYjUkUtVk/c5kKtKHxk8UK1seSFxmFqnsbj7
PtsccvD42AoiHjL0t7lIK4xRyWXoON0IEncgpfxTuiCOObGRiDw5QVJDrjvgJ6kQijjrHH3Fly/l
QEAiBttY6e4CagE3ksLrbnQXjCp4P7wxuYvCYsg4R/KMpem739uaTCPKFyewVJLw2pr8rar2hAzF
w4osepm8xuW7oOb5tsMowArMFDIQ1S76hd/99/fHjxV0wgeYS1xxH7j10ptjGmmAOiKcxXFo33dq
At7S6/4HvVt0W2ftJ+K0XGnbfFOLRzjB9DKh4bJ8JCKLd0JeL0NHwGztGftkfAES0Q2n5mBWW+Ae
JJbgqHKdpUZyj/hiUzbDzQ1aKr7TNdwXszEWBzgfi+bJwK0zrjZdJ7wTwaOhEnLxNEeJLfII3jfT
+2sV9FAk76S1fx/LUErA9GNR0dIkF8VmT6yTMKhin507Y9nk6BXQhnWYk9e6gASIlBMpK2DCErVz
+wVdRHxJrJQmoZMot7dvW0j8u8plqjuoLFn6BXC8PzpM02Ycxo/cvV2AUNoyytrz1qMKArRRhLpW
a3UQTTdbX9MWYVXv+iOCmihOaNqEwrcv6/AkijonZWWuRd4thMXcxajbtjQu8hYa/Lfm8lNR5zRD
xsct5vgwJ6H3k4RAlnf56/Ljm5Cis/39vH1ECxGrtYs0rl6WaPLO/sOzEPQsRPLy/+e8uczJKnmp
7GUXiHMFLhTmwyhArutzzjLiA7gXEmOksKqKC6vRRfMEBH7QprZC1Ne9rk8CmoNOa13k8juOe3ff
/WlJY/hgEwuAzlchOA0FNjyNXsL1JJW/TV6IkkEzmTUu+NiTpUBYvypjhj0z2J+j74pYlN5bFmn/
amoEpcRMMUOQoDLNICcLeVN/07eeZFrncY1+7BfqRSj8/sufwC2HvA+QdSXQdS5b4h2/trP9qVNs
8KBqnESVjaFZ62FNPIexR4OIY4XZd2ptq+pTKGvx/gkDi2YsLokMU3fpxQSYeaYGwS3DjAkHpMFa
nUKx63FjIip9/HTVCkMVywRe1M4CoeQ4XJipyXTZau4AFVPOamSAeT814mLkM8oHa3ALTrJlAqGM
EmIAiMSEMUnCOWCe787mVdTmUsrrQNGPsHtmDu95kDPVEhMj0B6MPY4yRsKItY2qeK1NVCoKbreq
xBnrW8ZUR28oyFWRNL3p1tPEkhlj92cN/b1uHlgw7BiDOf5Suegz2hmSoMv7Z8EaAy7FJwtIR9gv
GIBGUgiP58benUKPEWHKRH8AjpFv8M+caS09wvCkiPp3fcOkSckTJI9pPOOyy+xhdnLKIqYINGad
oC3mXSv1ChnWbtD2M3H1CKlS3Xwry3UOyBjHA8LrWG33esc3Y2Sq1mTj4/2hXC/ly5A02L3zqNiT
LMdbBoQCiDw43GGYnCTKqLJBrELhXD99TzkLyl4w1bxBjnTpO6cF0NptdPujkZN0PDbQr2HAlP8d
dcWCQUnuZ3y8meo35H6NhKIRWk+r0NVVs3ngiyfcOqOhb1AAdAaGCEmqWv+5razY0TNf611M71Oh
gnOgkWzgyPkPmuNiJa7r5WbPCJEEKMpV2grKvBOJvvonOptu8ab44jfYltY20rbckvobW3h+SeJk
u+sm/EF8WIFnpHwBtqvRomkbwRJUOiT3BvsPEpvYS5aU/q0kmJB/xJNI/i4N4SWUd+U467xocock
t/kDtpFZtKjpv1aeXrwweK/mpuXpzopVMHR5rtWUn5Z3h6ECGTQo2cVhLobDQcarh2Yp2Cdf/9lj
Khdb6hQZnaTmgapxGXZzmXytUSRWpK/SGb48X/7aaoUMCCsQ/g6DSb+Kf7qIc/H/hUfecoPHuLRC
/dCk56HMK+a45Ra+lEXusvxHnYp6qH2tbb99FNSntJk3pNkoU8tnlH2rxv2KZCjYKyEHANv7tyYV
HTBYzWvyOly9Oi4XcsTBOcy7jTbeRwnRQdQXyOtZX/gl92QCoMwneBrlKKQ6BGGcT2D/sGZVCwtI
Nn4POaEaSIljg/APu3I8jgIZ+gZ9sBZAiAwlXGQOxbrYHD87wAf3L8WAGTN76bGNXsNwCPYMNvbp
LfoBdJdZFoQ6MHBV2msHbG9GpT9xnkqbb1kqMcmiyDePaVDgJ0VhXYXZtSuXPybMKm7/iWDNvx7C
AceIR2BKeVfgJ0q/CdFAOGix/6Y5kTzjILsCK2TuWqxPi2wvrbFgzPbtvJ5cWEEVEL9ETGOrgSka
uH0CBqCWb03v+aoxjASbsEMzJB+XPzkH637OzikOB+u6y2dzfl/0YTbc3r+keUMKAbMnxnqQ/IC+
lXl9JTeJ6Lf8jsJ7kPP/8o5BxhqQkkx3ETt5N3VddpJZwnnXzSpynUB+qmaHY8N9dJIkAZCdNzP5
o3YOKH0qiv5zQ2VeuuX5736mbkXk/zDvtXkfQJ7h8B4oLemW47V0SdDyibvH67AuOfFJySqHePra
28e833NdmFcqiJw7daYoqKKnHfwLHk4r0JXglKSn80fr+Y8+R4+QDcszJ7qINMEKT/HdC/6qMMOD
WV8hvICKfAmn7k9AmYcZhgs9lBug8skdDDJG3CYfoEnjWM+KDOk873SaVgvt8p8+fgSu+ZSY9wgw
AYRaB1VOn4piqeIL8amy0iJfzBbd8PlPT0FJxd045NxBjJU4wmN21K4bo2YJQPIEzhyi4KJdW+6F
B4LHjrxbJ4enbiNm0Q1RQmvMx+Htsz224x6HOfbt46DyBSw/S+rCWRPjEocEpxmOqqGLy9VV/HDP
qnmo+p1tAakBcwGySA5dJNr6KvTovSQnf+7yBoBkWTTAFe//UCvYxQoAqZVcD8CGjE7PzzWXlXyj
hwERLqrCRKV0cGiZ2gLm844AGpEklc0uh6Jvw7JO5eOcmRA2F++PHGpghjRXQmptFp+z3sm9Ne/u
hkKK75KvXlLGead7JdrUB2TPxfjOy3u5IK89n5XHAhsUPugIJGakM1I0B9RJDYXuaWyltHRUHkxD
zAfo/lMAyB+M+Kz+O39rcCTS11YsowAHMouCenU+3Y5SB4C+SS6pPjsmKysEXW/TbTtxQ9x0IwwY
g68J4VntnFkXGwMJyeo4RiHQbKM4A3tton+v8+oXN5pJnzl9v1Hp/Ay/3mRuqfvBk0j080IdMsrH
Twk1gPCvGUdvvSpQcLDltpEX8x6Zr1CGtTsdmtEDXgODKAjcemMFcEULwK9OJyvUCrl5swMtLfq/
SFvVxnaTdejn2sxYRd8qp2gDgebQFPsgPVrYsWx91VEFplCZWrY2cHdyQsv1XlXWcNdui1hkHsXm
GKYR2nIMlECIiyoS0Wcn96J5jk9S4XftOYAf6iBaR0CNVnmI06QMTyxplSc6D8SavPyoh+N9t342
+1+a0dRgz3IPvOvTr0jKNqsW2n8zKcZrOXs1Y6PX7sO2puiuHcqQwxzvGhSWY3NxUpRRw4tG9tQu
J2wNPfPV+htAFnAWTA4CbvCC7YwHJ+qPsfndcjMG3mtADd7uZzH2NkGogVIQneNreIjLy9nhpqwv
G+Se1yQ06AgcFllstqeRpFoIp0MOSxvt7PLO3XE3lgGpDwMeWGsiRNBlf5edjOW1HX9mRXKOyoqR
2DedFJuF4fz8FSSzOznxYfprAs0y5P701SkkuWwoh6RsC4Fk4JM/8JMoabvj6o6BBKLvDMSp0umQ
bkwv0wFT2MFrOqP/86zZZnAUlfVrcl364XAyvju/WDbJ3DywXOavuzuSNjhjryDGAZLifapSgzxL
Oi+oAJz+RLmLqE9+wakKIDmw7rJu6rAyKwq7EadZ53d/kogJKNCBaGiTbguG8yf+HZW4RiPqlz2S
Nw26fehuh5ICOzPRSxB4cHiW4J3Rv+0LcF8W+wa5UuVh6QsVxOMXqaRL4tAiN258W4Wwy8LnM6nh
CAah/Uv87dz9Tr5OAKkWAQo5omtNgziq9mrODpDFiL9Y7A7lkRU+6nl3m7Zm6F1D2ezREQi53NeE
30W+IPhsa6ZML8cTi3o/dRGz7OQb+ZTw+Q/h/2cbBoW4lka8tU8OCEME6tYSWMZb/ZAxCk6wxuOE
+tP56os3mRbs1L9LJatzTTx0jYbLqTb77PneuiyF8wPDjxa19nG9/W489TwEHBHE62puQ9B06VP3
KqoYDFoiU0xmEODp1IYLoEt1tflymunjQ2FitEkPWv/W2uls3w0p1bTh9dx8h7wmx0Zs4LLOrR2c
UpFxZkHVwdg/sOw9LJPa6Ri/GyH+Jdxdgi/5qiQQMGlKD/AGxgRRSPhLzkU4WLtQEIibq+oVjtUu
6dxtaouj0Fiy7zotp5VVdIaBPeRBQ4r8jMIvWjDXwLlxqoQHDS9dxsFRMGpIPQ8+PCvnfZnU1W2r
l151JZqRUc0SNFyvNBQJOQaEKgZAzSN0Vg2j9CU70L+0POty4796+qrkuQrdMZuO01PMxiPdpxS9
4pU8yp/4oTLMhChGAaMjvgvlB2Xvx4dVGDIEwPYe2h52P+yHksyj/bNHVxVtOAK2fGFJqArKIQAe
5Qy88+dZKExv5tqwMOzhV6bvncUKC9N3w3FiTmLYXFG/WWf0WQ+TYfal5kOAWm1Bh6pYgeuxzuP8
BvYM0om7IdYV0+TmOaiOCeAGjd8a3JFk8O9/dI4q2FHIUx/cd/viz6qxWyrw63hhoXGReTP8+yQ5
M9XKVHrmbhn+HG/NXKSVnveTo2YDL6NwQG3u3Amj+rRm310efpeCBojbEBT97ELXhwbq4DlMYfOE
/tdDGxdto2gpdNkf8tJ4m7A8OETZzY+ZoaFSfxGi6IIDK63+eyJJpnojCqn+y9wekCjDp0S4V2pL
XMv3L9n/lJSUQBdPj2jlAPpQtk84HvmPQJFkyZgaXOmol5vhDpZO7cECPk70cv3BpsEkWgg4MSOF
U5Q9fYSA8QBAxAys+YXoLAERGSpsuIIJbAhAfqZEJkQkH8N5qNVza2M5P/Q9GZwY4GZCLRw1dpdx
dFUn2cmiT2HuOrdWYXDoSSqQ8vGEF7eZ/77D8XxCRC2eE4Ev+IM0e+qAGub8uHezBXTwE3REed9e
Wxkm3tLJgH0fmqRYS8FDgNVziTd5SAc9VCDJZt8Yw1Jkqjuemplz5yvrYjhUr260o7w3KMj88vBS
r3Q/EoTpYRqmI6dUMRdsYbIdcLzKJ8FTG50otyUjQO9d3PGNo0SYEzXpfYEh/h1wGky2qaUPUY0c
aR6a1ymZq4tyKR/1i3leeK+Zm0Egnjz6q3j0jBeEDWOgO09R8ABgtZG4M2Pdc18CKFaGVs39vRtl
vnvkpk+psGa/L+Ix8blsRAbdiz0hc36Uq3SWoj/WZekiMdvts7JDCpuwTouRSsg8ZT0oPtCh0SYE
I6EHtKhbtqEKZOKnzDwdLgPtamtMyzZ0bQqNgbJux3MkEfDnIBTiQtnBQcT18I1jxuQ0N6mPXUxr
tFONkKCqCVva7rxvxV9EZB3/ihFXqQJSEn3SwNQojRBADj7pU/4UFSj+KAbKq32vTbYHOgk8guGP
ReIuxQyVyXTZIXEsFBbzYXm/65fQTbXdd0vPdI92BvrsgIQ1+u7pK9a3h8m3rZVXxlhoBGiKftwl
yiONwMxu9ETsvQmFrHJEAdiiMIC3RrO9e89AIvvdeHU/0ALKPzeOhjDtcXcuUCJOixIl12bgE7/c
CHm7uOuBDgc0Tn4ex275CR8jOBmhzhVfub9xQ74bl2TF0/R6YhkWNVqCWK9VlkbOh591c2TtgvA0
HTRnM2WF0reeA4iNQSgU+Re8BGeYe7P8dbeyskCdBpfiYXxw6K0R3YBxSIQ725t5wWnMrLIowK2C
FnatAdi9lWyuAxT9KwjwOOPmVBFUPa8YqT6JvfIq7fL0oWQGNic4HFbExCSVhjttFSuzf1fBbLlC
r8Z04oB/ipkprBKNg3+FCiIPEhtGdCG2+ObXEjMhsiu/udACjrG25dQUscwpNTy/zZClbB69Izd7
iTotWs5Kk+EJWC3c+YOODjhNFMP+4P+BsPXeUJOHhaz6mJ4UzcRPqVaOvuuvcO3d2y9Bhd4h39Dq
TdvSY0g8z20ggNzbrC4lwisVxIpMkiI8R84qRbLcPBIuE1v6dD7ArXL0R4OKLiZCrnjA0pyfUQRS
PR7RzHeWUl472Hdw7/V2PITokwK/5o5L3EtN0Rw5/9sgVsPZQ3uNirSybSc4sNiRAUhWWh/dbE1Q
pBDQX4RgbDjfFgRSqqmVJUVh3rsyU1OQvXSEkWc9BTn3HovEV7msu7D5mi7uUD50ql+lQ1v/0anW
pboHiHebeWGVMzCUxr3327YeeO9w3MLxVRgWU1KiS7klq0b3/CzZAiLYvz9pNy74AVBEFGYdyWrx
E5yEKISggm9E7gxtQHkzBkqZ7TYYe+WTJ5DxpSA210T7iNyEHXFWiXb69Kmcz5YiUNi8O74fJb0m
4O/SN+Gtnyp20D+xTkP7XX5qMMZ/U84hvcsTj0ZYeTanwIhydc/OZWyPVusdYelmj07YqHYgb/eR
IC11DIRb2Io/QCh7LXk8FsHssFmlB78KhlZcR2y1GR588DKZdDjZV+Nf03lz9JB+xJ9NA4Mv+3cT
MTE/ygXRU5fWjmDM9NqP5bplt4+alKHVvLIm+2qeXkhQ9/BD5iR5bCCULbd9TqupOL603jUOR5je
XABsPIgCvrD/aW5ciYBNTGFdUcYEv2VvqWkUFWt0VydretlZDCjVJAmF3aASb16zi2N/Y3K00nbh
f7SehYGJSnEYKDnDXkE1qof//0ckJkLoN3R+VPFzlBwogtDPy6auyQcoUy9DlsVOLzqFkV+MxXsI
gx33zhkRVOXtVjuZPRqX9HW+vGtNXLmCz0GdonxuafoJT5NNx9rL+V9z9VGjSn9hiw6s8qUS/Mss
trm/e2jxkvUiiJy2XiyL53WIncgDLX19gt2jYNlEjpQwiDnqBqdFPUYOqxXB83NsW0N7KqV+wK03
ORt45X1JkAQI3WqLK8gt+H0HJm1tI6aXwPIcI0i4NpeH+X+qkRm5OUR1dB95b02uoOyDYu0Pgu80
hajnMAxhfhwJ1tnSq4Nt+RbGcHTKey9pJFvlRoXM8mR45srL8V/bvbSvZVtDOOUSN9AFneVVV9O2
Fm+O0GZX5RR5Ui/0E7Z5VCt82tCfJKSXPru6vwLYoEZQxq4+zns6Q9I1+fsGtegYW28ryxSzcSUt
L1Tsjkrhzpln9Xl/BGoC2dozcM8c9VTsFBumZz3fvFB6w9ofaD7f/JQJxDJODu53nQhsoTBGLsgm
MOuH2/OTe0xMtwB8EsimZm3uk5TlZOZYUWuMR/3bMf10lf7zo/EOh+3xS3mZh/R3AecsJost4zQL
CJuPmQ4+RGwOizQ70o3P0iIaYZgqz2Nr0LE4Ll8NH/FjQQJ0pvMxqD2Grd+8zXS7lCMElgkBYc+N
gyWPoUj2qKdPsEng8YKxxDfxxN99WELoUTS1nhRwT9i6EmgI1pQMIgCCeANqJlJ/VsZiMnFjOeY4
rHcvmgNdFAhXo4Wg5pCbxSnH3GNwbUAF7KR94pUI9fUtGSios5f/jZZXRlMJduN8ypakD0SQEKGJ
F9QmPHWTemvSP2VzOgi9FvNm/obghkM4AqQY5p5E0hiBd6G5xRN/4q4LH034FFGcnAfimenrq0X1
XoAS9V/U8+SIx9Gd57RSbCvxhsKoTCbERgAN9e99TzJEzlMkoL8/w8JZ9eriwNaiOmRHuzSN7vOf
Fd/v2VwswMWS9sM0+k9yXrWP4hn2tv87G9+FhG+Zj0TLlXPSOTMSlzJGNqEZCF5EQ6+fku2Wt+FE
aqva7+c1zQdZ0vPQwwPSD5rnKOHz9cKzQYd4r0jiqzKcbVM8pF9M4oEGuHJjkagJJr0jNZcYDoRw
76Z54KXXu10VLhEgPMGK0w8PzuQACUApFhlqSKWBTA0aaI4OT2SOrN3O3xXO7vcNo9iDFuSA7bey
Kl1R/4w41PgoJD7p/szxN8p3GldA3Bmbb7mcixhTp7zNPIGTPRF4fwta6hLBxMQHX7XgTyh3x/wD
qHYGgqECTfuAmBx6HPZdNkn4RPNjMP7+xApm4as/bb7QRYxnC53cZmFS4CQol1FpyWMKhE5PVlnE
CgvrHCZt44/zB5bUUGbn3GC50zQaPdsIMFoV5WR++9On4UNQ3WtjILbvV99qZCLd4I6qqilcPncv
whvKeCOJST1N/3gRb7E5CM/QymhoWviXacYudFtCVUH2zvizToDlp7+UdFgXxkhRh88bBjK9VAvJ
JwmZQx9JHnK3JsIu0a+GdnUkzo4wrivZJlx0WFvUKchY62bz4oBUiNe90F1q8YVxd+2qjk0iCgGV
c+IPCGuvRKBYdYMQbGVyI/TQ6bx7mrz8s7tRZZOqRotbjoEUQ1gSbZD8TUgiy5oCYJgyyy0TdhUm
dm2+sDxHYx+q1LjijnFs0h+2pcq7rxTa46q3O0WUMtruOg6uwsgdKupCfgh3yIH7zeDQYSRUrNxn
/ebyKeyW2BVnQTvgka6CIBr0Kfw8IDhuJsDAOeqQZI1fBeXR/u/75eNQx3x/UVc1bew4zLkOO8J7
El93otywfW/ELxleDWZVGEHXmjKnAALupN1NPY0xhUoUUWXDJikJzzs1k0uHN+fSWX4Uz3hnbN28
pKwqbGvCf8fUcI5ubeGrKVdwZlSAhoQborYVdh3XicKYSc1tSFeoU/jV1DTMEhZkRR8RDhD6MRHR
7VpVfQ/jDtdFHbhTabWEmBfzpvLVgTAZzz9q9R2DxEpz3mbwQDmy/KO9Hhm78uyLG+bqaDPKb1zO
93w0RRd9pzwS6gJ5wUOtp+quEKBgaXpIXscrKfgJRD0ja4ruY2tYo8GpXSCDPcXTpGXudrlTLQj8
q4ohsoVx8+jQY05XJfXxYdEHNQYla2mU20gra506xtblhRNihhc2Ht2BV8QCqKXqFFa/GDDQWnsY
tfTa1QoTCBh6rvd8dmH1ycVTMqy5GrwJt2/tTm+1zq6UhCaM9DqrPXqY5yLvsHTNT5qrjIn+0gHg
q8mqZP7HtxRdSX+YLp/PSSwmK/VAWRQ94z49QtI0g5kEO+iYSbCO6DxEyqpOTfLwwxHK4eTxuutv
8DhfhfdcBnHPL3xQEFXUlS+FtMlMnIhtj+nC5NEucIp5wqdN1bPG3UvZGTfczbkkbD5yNv84M8lA
CJ1lhJHdUml82ny12FnPROrGXwgOQT8e3jNoRMqNblpFqWkh4YzQcre9nQQ/u2YPPLmrt7bdlKBZ
3tcwngbhvhRWRnQCGvbMBfuXQjjSIesj0z8NaCpHx2t4EkVe46YeJz99JbbXOI3n+tJtoyFQJF8M
teCgj4Cy4DVRzUJOdDHrk4ZpRDrngPN5sMWyUwR8vg0Et+X6rt/ZinPnrJhMPg/P5Dg4PWIzSm44
C7t9GmkHzJ7Dm7kehvuFYChXJV/lwgYMnaLDtTbM+UGuUbjh0GJXk7IosH/hOUEhnchr7+MGDN+D
r28ZMwa+A/GP30hBatbxYB4RIx1DVNOQePsFtgyoQ3aYtBxZnzDlzd41H/Y0VDJaHTcnnbnsH+3L
LwTOW5+TUO1t0uf/uHr/5GCFjphfEBlHiQfWW37a6sQaQwsTnCGfGPfjMZIrFfiYKG/9GJ5roxD5
o27Sc6iIdYIeEUOpzqqfu0oSXUC49kEYDZrogf28HVQqW9K+5L09voDhbkx6XTBQd4lYbklKGRP+
NORdpSfyrkdRhWfZVzDLZqGeJsLyjMmstZOE0pG/HTHy41YiXCGOiJlAIXeXpOs1hIrvzkWjcrM3
aVqteXMSFVYrrG8+m7cvL+INCEEDxn8nUnxvTR5XYqLXWEb48z2269/epe/F5R3ODQ8dXOChzsYT
xA3GQbEGX/4TeM1RGExDBIio7VxPdbd7odod5gfJbxIZqNsEduisp56lNdPbRiqqGVzV+v6BxHLm
tXnJWYBeY70XLp5Cz0kTv92YESukXbVpfFfCQ5mUedOEbnc6ZNLYTmEWiaZc4vYpXQBqcNyLRA9b
Df6vUsi53cbVHPvlvntvcoa3a8bvFnsFI3QbOiz6BNLebglMzSUOjx4bRjuYpuJgwGZX9m3LVh//
mf2XvWNW4EA081q2DOH9myERartVsgdG0+c7lNOJhcqZX6sos6+VRJEThbp1BIBcAQkxqMn3T+dV
ORnTaDZzRwYMZsUU5xa8nLqimPdPpBOorbzCWb3yTKb4gnqXDxa4MWc6IWUdXPPfiNhPSQOuFnVP
7Kd31ZbKQpsNDcTpSd9D0Xgwi5qsfTCR++DjksCghHOdflZ0fd6stRmeMUU8HPU3/lqk5M81prh6
f5VaxVIAUpGbqeocAgoOqOTWRyTH0Y9xQkGAbwyKUmSo2lYwTXa3PXrtRz2M4T3Ullcmq/fZQoFc
Dp+zR3FsJKtzsBuuW7NFpyhi8if+n4LtN/FEfCYMqMnxi85oWU1fdTQnH7EqayEk2yAml4+HF/0K
mwdCSIyVpvSOJPcIo5j60l12pw+Z+SQDAyohyFBPgC9Jg5wR1vhIz28K3QkuHIC8+YPhHBBkb+zX
y0zgOpaGDr3GfjcBp5vVsrVxllNTdsjQhMcMHRVBZW+8tfSOST31sktsLTPdVMRqE6alME01IBXm
/figIRWfw9s1XF3NOJ13/JLyaIaWVRE72pf4/romJZOA8K6okzlPhj0YSknyOgATwO61E97IrHBK
FaORlUsaFsJjVMqcMUcu2ORxHFBjyxGUTzBz9OvmPfiunB/mjDQZSMvfooIenXYu/k3OgIMIUISH
eWpVGYgWgT9Vrjg8zWB/O/sAM5M7kym04kUUmECIUcQBncrMaUMWUL1B3V5x89BUmRyzdvmtkWFh
XSEDJwj6dXl7UQbLtkxmFYyvHPzaGFYk3ZKyUFqZnSe/VOyZdAAj65whIQ4T9S370n/7WF73gSS3
Jo2hZDJsYK550K7drFYDhmu+ByZvm7ZlpsWodenFLImfoemW7cWw7ssiFavvv2TD9Z2CXUmhYAaT
VY06GlzAR25kqbBedHoL0wqAFbfM9sauBkl8jRFv4+vs4yr83TGnJklMU70VIsqnrEt3GHVaTL1Q
UPYz85vjerndkWPPg19kaWIOgtOYEHSyviSE4LoAAFyfLtdK7Wrmfxp7Woqy0a1mNGHv7kJOoThM
9Kk8+Npkd7abY5LjxvfR8vqH5tDze+yLCo8hc3aXApN5VruVCdQPXfi0Ena+jb1H+9uoUh/uo+A2
J/LpXdes30cyp5a9NL/Uh2X6SRPW8FVvbogs+xgLNbYrwbDAR10rPVPJdWDEozhHEUxRJjRoK6LH
ATkh+zWC2hQA20e07ulGuLSwvy1g1HR8MuFFxdsRXWUOAU0r9ZP9s0x/1Vg1g6nAuK72a5xbc2kg
VU/dA92IxdUwwQTYmsik83XtesHG1dw5CzZEc+6afzb/oZrkBZ9Cgcpan61KDFMPGpR+SCHL05HI
SqV73YazRcnsoSZNOfv9ngEQ2SqmjCi8Og3nS9uzRBkvkN5ZwaPW9hakGK+vm/AugLDIrvD+NnZu
MzO/MdOTxK3KZdbfi1yvlB9exosTMDB983oXgvWph3h7OqQMwh3mGDAb44K4zELM4SW6e9/H0ELi
4He3u+fBCok3DomCHL+MEy6soHG6rJtxXqNAm05ENqJugPBEi5G+3xpLQ5riX6ffwzG/gUttpfbz
qkh6E3rsnbah2S4AbjyQpXiAJ5UXu+t58Pdpy3jjFek/pswx3cFw5typApCYbZRwkoEGq6+Dd9fj
Rp3ZZq9yuksd5Y68kvquQaDQWOL3eYz5bQl8QS2R+OP9QBKc5e4unh1dMzKYHmkoOPO+oxDcgTCn
vbQIUymQ4Tu4C1dsQpr/m7SVmiNpAL6DE8nCVd6ZM3D4KPSxLWBmxaLRcnu76/9OySL17kM6tSSc
4OI/NioCFiqRcz+cKlpfew8sf2K7OkQLBJARv7w6tBcoGcaNAwqX5bXbVzupX6uw+jZTEmF2IgbC
UsuW83ku2tJGlU9QkvX2jZ8+IvFZ51R0cJvArgWIKpiJBk/Xk7QbCV8mYo5T/8vdARNZ2lt/O0hg
YHrX6fr635oRAuVX/rLDDMHg6O1nDoL2pSldq6IxGkxh7FJtsKl68gnUdzptaw8Rct37rUHXmwn/
02aRRvp2W0mIw3Oyq3QhVexldWprnqJsvxNp+D2jQKtyCH7b5oHQUe2NiarkKFvR8tZXSdwKpODU
0RKbtIubeVf5BHY/F3xnHoWY07XiYv8SMnW4lDjp1lZRvAuNWFe7SUoPSIr2FIMrV9ZwKK/XG4W9
oZqGHH3TMFtqLjoZcCVznFhjydaZCh6FV+Lc6DleE4Sq3ltFnZIVS7/49V2LrOPrXbjziSLVhPrJ
BkZ4fyKT7S/sundz3PVdYTfvSaFZakrC90Y3eFRKtV0U026TrrQVrOeu4F7Syh9m5Sch176Zl67L
aDVNL+mWYi2n44dEuHJ+0dF8iEVVcsRChXHdy+dLH4feaPUnA1i9w/ysVgNSj5SCKnmvnE+sz0UD
SRqbT/XL5cx8O1eRst/Z+Zbpjsu6nx2iqYpTVEe/QvetTprV/VO5RopytVznv1osFoI2ZLjGVVtl
5nSqonpW8gYhAVttmN0meJRRKZ5VPMixffc7XfkrfphToA5t1lsSeFYM0hFwW8y/qY9KuVEQT5RS
3i9vdvVemNc7gvQ6HyTBMSEXLAHhsarKUFjBNAhIq3qIw104vHsypuu1gObpF6YtN3dqlsyB+8Pu
xv12mc7Xu7tcaDJlirIC3Q3vZLJ9DrAZIamAE85jSMXWd59kK1dF749NjRK+/6KsH2Hta8gsTuMf
4ucHez9W767d0kFjun584TYVMckMdsbxeixU2RW9ftkigb6bAih8EGyoS0FwSjjbIiCDRURg2VtK
aG3VRPw+oW02/Cbu5bkgSuBuBW5dALe432ZY/KE2GfqlvHyrXNfz4UEbdGJjYIxtOQ8lO4NfYkyF
NJPKS2b47hKyEy7Sfc9RpzXJQWDERKGE9FhH4LI7CWSvqtv7TfehB+J4W/jbDbBpfp3UvAXH9J9S
f0xejBUjbEqUgMbnvmb+zYiVogqGPEyMzA28leQuDsnK1gD6UcxCcxp5SR8NM72qUJ1eDIcOtUfh
S12lE+EhMldwX2qCR0XJrh22OxdUeTrm05bfUbTgzBSXNj5ntfQCDLiXPTGzr0NM0nV/on+3ifgX
0oJzaBmwpFiOPL2Z340l7KQTD15kUdiDUHZX4knNvZEypAs4/c4xMr1SYqc0sSvIyKqRkR8SYi1b
3NXqqsi9+66ht+qSIEYxadbnh9SJo6eaIYQHPxVo8UIjZxgMmSRKJhsj6CIDoxxhaFtUbQGqMcgF
LxOgcXEybXHCSSvyfA7EtvE33YVpxTsGnKdk4oEOZN1gCiyRxqRicBGKN0iw/le2EyJ018yOTLED
dGtk4d+Z3yr09XwiIWFbBwgtQqaKtt7rFMnNaRgrMz+OEaFq3YOLb3LnKEn25qOu8FU9PfLj+f4z
nvMA3lyzjmJ28KJQuFL6SADXGsHMwX3HiTlztRVDXMJti0hL7Cd06qO9F0sWhknvamq6U6pcsDxO
efQYTzgpLT1noR6kMI0LiglfoAWkWAXBrk87m35ZPodzaizFVysqUzFTwIm4waTA6de29w44JGZ7
l23Zr4HTF51qVNyd5zykNTbH/8L0p350VQmxdUCj0VWOnNfNe7RSIXEk/clz4xD3uqW8nVj9Vd0x
ce+WJQDC2VLRk9IbU0Ubp8YXvLplzdHc1wWZPmi+GIf33uktiLyK8XFL3+YgLFFLD0nxNuKl/1o6
ZXNP+hWXIv/6HgHW9590KtFF8FbOgvHoW/u8yOFC8FgZzwpcR7HhIBgN/SzntVDU61aHg3ThY0OF
7IWQsDT4YGeCnpsC56X3oJpXby94vPJ0QAwY5YDH7XZBUOjNLKH7ezu9FcseNvrg0Q+D3H7a/W2M
3ccxvTfo5mv30l30ynLuqkjKCqp4rh7qrCFlPXsrWrDFGdueT69Ehut6Ba492HoOIE5alQpkA4RS
c3Nf9Yp3USCdLPT6flxen5NUoDpfKoRjzx8/6GOnbxmcMDbROPuBMAzSAMbByiGRpN+PksF5M0G9
nT4b2OYjaczXondRDT91Na40pApxlivE6nyCmEvyxrClu7d3Xs03m227jiLgLWL5ZAl40pkl52eQ
JvIskNyS1f9u3OYLtQlvK2s1qsFmUEOix1uazgR4348VWzx0O139YHlnemFwf9T/cSzQiauunMPl
3RuVluyWbJlFClRrce2HJY+OsfzH8WUUbJ0DeyrsziV4xZAsEMVPdMl8JGT1gzeYYNCV+/cvPneX
rAR4obt5kFU7MRcWSbw50p9UhesyC1rdMwOXmycH1qn4Cvk/gVbiYDLC++zdC6TSKxT8DCGFWXDi
LTDtU41RQhANGU0X9xV2JOPIztePxEzBsPcc73GQJ9Vw7g+7g7HrZpzCYuSIXSq7PzWPecFTTRaa
U/8vSl70uIDTkLb45p/D/MF6niyAzQD1Zlx3WE8rqBYVbPrZSEfv3AXmTKkCNfWiR6DU4lT9pDH9
18bbN5IoXhfahHu7ANAZDI62ZkVuImg33knvaACs1St0iPVCpPonuqabhuj6kpxkPr7kaTD8x/hZ
n1dmi9FRRhxwA/i5A4iUIVni9oBm9no+UTvBWV7edsuc67UvnY1qpP59miTj6ZFYcGRA3pXJ3khS
75P5E9a0amMgYhs+SjPVMyMXIh/aIxOBA3JY2q0bnImZzABh01fwPgbBLuRZ17XPAExtWKsACrH0
FHBDAPD5UwmLTPdP35yhzLKKQMTku997V0iiDVWw20zMae3CK+yHk/Q1HkrKlsZ2zeIMIPz1r1KQ
LwUGQ2rAAMn3gwlSvoZ6FrVXoc+3IraRx0jm0ShiytHfZjedE5C3BKMFSluY5Ju6ixIkZ2f5UlhF
YzfYQIgq7aT4nj2KHxkziuScQYUfyMHOTto6Heh+OHoIYBbth1vNoBJcunNBMuFcAHAnsecGNwNT
OQT8bzfVaVDieD8hywsw7Z4SYkH3CA3FUsC4BtECQKMP8+msdf+1toDuE2WGUeIgJfx4uGZ/Y6B6
N/AkEBxlyWiEciDh7mtqdOJ9BN2AAOW52vW715uOFOWAHRrcwgEONnRn9MRWXE9NcsuTDUzNnxuO
lZ30AEctfW+geeTNP3KqReacK2ZkVq4kltsNkWs2zBjOxeyNAiB9qxDz3N9F98lrBX74ZTT2yCYR
HfAaEyX1OIutD0BR6Oi/WXA9uU2UfJS/EL154EkKdEiSD8vaBIDArrHOL+NS4tt+J70vVQAo91WC
S9eb5F8TooJZ6POocDBPHL4AUWSqzAEJieq6qsoOjdZmpe+mj7ptsb7t/hBY6QiEjg4v9H0k3h9U
v3wUlutSsPJo4B7JoEXb7/e706l8vKWJR3SjworKGc3VO8vjrkV1LmxNKw2Wnz8qJF1ATtuPKZTI
eFQQYRgUURoN+3wIVjY+qJzhI5ZjJNdeV6TbnXjlLFz2kWQAAD1VArajt4gmYLxKloG/WZB+3oEj
FpW90iVjgEYf4lxoHUX5GQE8qjt4EyJ5gFL32KiT/7ruzjgXzd9l2JLUY47ZOZFHchTjCtxROmAW
Peebv+BgF5XmqjjxW1nwqkSGq2zz20TCxd7yoXpUM3wew3yth+kbBSaXTUdIdNR3Aq4awsDmPI6m
0L5tyIpS0kYvTt53GoLUHisjLqmQxGbxj3QH/ZFpp8QnDpzBITPcydA+CFHiR/E82aZ+QXElK4FZ
VQ8vOrUIZxcosK42dSTxi5JMuGP/zjQA4PKzqGFrCSsp5MhD7uP+8Eiuk6TJkSztW8IS0CTrY4fH
bnkBV/HLPyigIh2gahA+E5v8mDbZLAW2gEeV4TmiKOjqoOEbFVJFAR/60bn5uMOauwVbeo3Pej+u
P7+t33OAUP7e4lgTnPLpRI2kuX4h361vY/BCzfgvQCXFuqQVQ4gOcIKfdH2A4VycRCxy3/+DlgBX
I9zB9fapfvQNvxEBCWe3CoU2PrLmu7ui1uwQx8BxjLpyjPFMKBtX8Su6LjxVi2EWxdyphCDIQani
s5YJYtqRakax6ZtJXEimbd+ckus6GMqOhGnPegIlGWVsK+mQ5h7Y/3nAOcV0N/kFytuKIsbJRX1w
nTcNnY44zrIBobLQl7BxsXfh1OiOOghyRRPYwMtHwFV/A8Du/C1UWFBs3XlwVlPQ8qbPstznpIsj
a1hBaJlI7TPoPV3pX3Q8YUCIQKLjVwetEkzJFq1R0Y5fsw/YXOfG6gqcRAolNWneqwlF/JCAF22c
dwgFcl1yWuJJ/bUUxFFnxkS03k7Ql59h2Ebbf6JZ1mKq0S5nm7teUBxly721681lb1mlAb+0an11
bYt8ne7j5kw4VHcc0+h33j85WYlJMHnG1eLxZKUob2194sIu3scTUyVXqx7GVvR6aWjJwWf/dFe5
wDjqsSWVIP11gUm/vCC/uy5cNAQDeKpvN1Fsjbd2FMCJiFqlf4dEnrInLQClL+kjZbuZu70671yu
gSQb+/enQ0Ov/C+AfaKjxl/MY/xP0yH5jYD5vage+KPPO1dr62S/rG//uSS7G06jlsW5jwSi0biu
Hi425JSQdUxvepxjSWleUoQyqN2tguEABygmhagMZk7rI2a9BDKuml5D/05S4DUR1ZFXaSAatyZw
mdSTnqg/pdMzBEd0mA8Om8RSDf3T3dhSIszKga1wgCTNVYVIZ4Az2sYQJs08LYX3yA2Olei/UJIM
csWUlIAZLJd8dPaapheedPm5jH4my9fj7v9PiEhj0kLPyoLf2WnRqTAUMsNs1rYdmJlXB/Ocu9Uz
yS+V7q4VObOcP8pI2tyOUgKo7UcfoqcD/L2gULwVjZ8e72xjcNRKM4oVJ+Fyxn6sLD6LpWO2MfIh
gNnd6iXtdJ5U8McF5ZtdmTZ2X/UnFVxTVyUdlK1uqFerQu65lsaymXmRwvIV5fLxv69wl815Il9Q
Sk12nU1ylP3Q9Xz2otdNs8cD531PNtSrB8XUCkkVjmMohl+5HSnYKsDXdeoZ48SXgdEWioKV4sAQ
Cala3mtfNZqInQhZXo8zyhDPOtEmOA5uF7nAFYZEHyojt8a2WLZL96WRfRcfG0WtzzDZ53yLf5Hh
mV8hGQxmFA3AnUN5+Tc9P/AXzvwD4nJxPxEvpu6FWTJxn/Zog+ONLy3rTnsUkhMccXGBQxNM8VxM
yEHu8bTFHrdnc7U2Ojz1zEIk31xvyOB3LM4Q1LfJbxbXnNbn6mLojvrkf1vG2yMllem/iQkcVEqD
cBi28yafmvq0ZeyxpGXjW9uChDn8Z+8sjvakgJWvnxmhpOM29OXOS8UzLe7mzs5MCsyUkYdJYkM/
OLIxIYJJAroOSlKxVMQG6BjciWXV+aReLobJQO4yQKTaju/C6lK0M4HImmkTRSqvKbj+9viuV0y1
JEnGZJPz+Yr+x9leyta4g4RBTmKJuxi2Oh8HBtW1dHLviAoxQdYlV99IbVEoqUAa3h3pE+/JnFCF
PMeVb/QIOUW52MahvMVzl8US3/B0+u0J9IKFFrI3o9ODx/hsD7A65dttYv0JabQzcw1zJ8JGrCLB
/f1XQ8Q12H9xHxdjwCT8zSiJszN36s/w/Ms5tYnbRFmtw9QvJ6HUaJNiqhHL+Qz/oc5pa3dIWaPw
9ulM9NlvvKs+T/CP0ojgewEbSPDpSemPDhgJUnaUbnnLfk0RAQihs3xFHTVKGN8qRf969e2FWo6i
VXtDSraiEviRsUSDFN8vcsb2fXA1nqWcAh48uiJ14j7JCRJ598zAyjAaJ8NoOQgxnGuica15Op2x
WEFHBSBai5L2lev3zlYWCpAj+gPWypPhCnW6mpEeV3h0sIqHZwewpd9I40KnwE27DWMtt6mqf6hA
3tXEEGosuqAUgJ5tZsgxhDkBF+ec2U+Py1A5SnxuI2sx6j9EC5OKIqEObyIKhbpKW6eXgsz74LSw
uPxNvDT57a/35Ni7lgWBmw0eE3Cbbk4wCxz7rYOyW9H+/0TBy235e9acmMCqWp7kacNSWGj/WkMP
i5PhFuRtq8tEfZb4EWSPZhj8WT6krJeW0jsLJVAQP/wna483MpcTPvX8lvve422QO/aoJq2ls9GX
/wPdXe7/gi8TWY0jgDyMiUO4mgE91Ee/cc2CnUJ1RKC/HpsL+0MyfwZoBXVFcVCwJtEhDyUrtEzL
Dj1a5n4IX0d79hNQCd8SRIbNX8kg8oxbbNF6LAki+PbtgoYQuI2GsKo8Rnhhoro9Roa7CMvwmTB8
5TFThl2+QbUusU32r15iBdTOsg1n7CHMrkdzqGf9PtLftk5O8rsNTsl9osv00ReoaYJFpU7wmn7k
19BO6SRC2FkO5g0pOrzxTQ38K5UF2b1SoEVatbVomDClNjFERtD0JIbvZ1sC5HzdJ2cnwICTaYKv
l5F2bdM0C6bfp+NMpFGumLjoLbxzOxx85bqZglz3nvIX+egIM8F/hnOjLw1PQHC62sIc3M3pYRhZ
M73WwS2KtheFy3JwuKL3I1+iNsVHgHZahlbMRLhTo4EYeJGUVVKjasTieEpIVrm8p8Rpqx9lLJJr
Kjz6r5wSDIktAsWILDoSo0uNvJ72rbrwJkAHR/h7I498UffvCEIggEKTC0GaHmendeSXv2DGjXPP
w26pwG2mIj7IZdDMwYYB101QbBihdeQLHSvii0atS1s32qx84TSZpKFj6duNbbS3zdTj4iZYterv
anrCyuU1i0a38RkRsvjaWWbMBqClhCjobsbJjA6W+u/io8Yhup9jmRwDqrLoIjdsrkcQ9/OFv/w6
GNF++/Hb1ZrX1ugTfzgJ8y5i4d+BJcqVidWwuS7yTW5/5VNO3rkSAyhLCAOFRWmFo5MaR6b5Jlf/
94bXECULpq78tLDj5RKjMe6+Aa11lt53mD9yW8mPkJw2l0IuJgG15Pg66+zqAoOMb0TsMlSuLUzt
gfEMRKGoxq0TbgvrznuG5+MZEkbsFlD3f8nIMt9FHqiutzna56FRGKxIly8sOasxT8wooaNoVPq8
tvNqK4r+WJLkivg7cNGhxHugM2gqLzTIpEKUI1Lv7jy8V9RSt4j/w/wOQr1B6+n6ZAD/Ov812gE0
D1ygAiQtZpwQoGC4PHIq+UQnDcVOUsvzDHt/sh8VDqp9Hq4neYZbI+ZJmlkBxiqrz0Jnc+55sSwS
xFJPk0rWoYNiC3gAj+Wswo6FgmEpQYy6Oy4rMOU3SFc05sW2do6z5w3psif3w6l6rtd1TuZE/2bi
w6hhSSV7RXw9cd2K8v5AktuvE/op4tnX2sOHhMb7f07GIue8Ib9cVICX+ZG8dUHQvrBWFeayzZY2
YJyrmf0M6XzwGIW2nuk2emY7w0yuZqEnDbC0rzzb57Wmf5CL/lHBzhZJtZfuJvpZgu3l8cwcy5oX
AhfGLJ/QrHbJKEIw/1czs+J+LIoVR7Z4LX4w+aE0wqmqBMGtwO98tmm7qJ4F4ElY11QeLTo39hkT
V03dzXyANILvNWDp5/2c2f9vU2pBwXvgaP5YqAjiQnXrqKe2MaL/K6opWxRRmdHr+7yaphIjKSTI
wRQVb0/dlf1rjF+jP7xO1AS0/VYnuiJF3Xr0K+e1RybPIcS8Mjn6xG/YnxX5KcgxMGMY2YUjIMmg
38cNvbTqPjKjXN+17aAEIv7oAkAQ0s/iHOLAFVyWzgL0t+r+IjcA/x4MWhP+lRb2WNWfHb3qI2Jw
ZZN4meVAkrRxUW+IZCAxKEaTWYnwGH+/SVvyQaTaslkYOsaSRkOjVFzuD+TBa3FZTpkMPdosDLkC
VMu5VaG1UqfmshdBstRyDaO5//pDG/nAtMk+eZ4lkkC8iOFyPCxxf9qhwZ7bZAcx733JiI6eqxVd
2w7VUm/aRSVyfeRM6iGvE/VBdaVQk6VdjypYxovMviOXYyFlycxk/FLw4aYozl4KWen1mSjWDJ+Z
k3/jD4HRWo25wONeB+913f4k4m8yMeLIdD7qf32fshlnpZh9zr6hQVnsHP+V0w99RZCvV/MB982j
lZET8CwE8mkqvRzEwfI/cFjBNqdi6Ax/bkvjqzoFHTdXE2OxLntjKgKkzsU3iiEa4qJyCrGHfi5T
VAqlsf9DhRr8d9IqVcidkUgrdtvc+BJD1fj8jlHUjRwoLqmRNpNY73+uwdVyBvVpFgPHyDIrIHpr
bAphgv2FUSbDyqY8i/G77dJQ7bODTvVCuybeM+Lt2XT4oGCuz42tl0/WhaZn+ZK6kZb6XRCm2zV6
UqFeC16a/+GhgM5cq1ov6GOhiCkTR04kyhsKx3WVtRZ/HvEGXI1OMTO3Yy6w4H2HX+hknbrq1D7i
/9g9MJpK5hlKD2xgQ4SL3KX+vzKFL2tV4q89mAV7ebi1tbfRPeAFTYZQda/3mUdzFSxXjS77kjsP
tffHJBAIf15Sjp+rV6gC0M7Y4PgMFMy7GWwyPR7PFaLACr2/zcmsJg3BCtQZ+iZ8rfBwVPZ5ziSF
vIenK+Fs5m5NpjCow3JWUmb4BKnDVBVo20AtJ3ORW/vhDg5CyozmTillrRsCc9S5Wk1QUcHLLYBW
j11apCegCEI8Y6GK4waN2Zeh7vjZCmA/mb0BscHb5bDFCCYtqABOac9PDXwKJ+CGKIn7K7O55VGG
4G9eyX3rfZTUwX74rFlwwz/tjbk3qhjScyMe0S2cx1OEzdIC/N0pqs8pHORqaAoHi8OBMMuMh7jr
oZn0j0q2m1U7O5JbdEGZGbOaRZaqzddphm2x1JwUFwjnzIDpmfLGnzEREM4DPtplUI3fzVYrXp3J
QyMQQnuTr3kIQ6o+jQPaz4i9GF5IHaYTYTXNbMuyYqOgaLeL46zQDcaq4+qxOygUorzcG0RiyiAK
iEtk97eZYd0IpVOcYIQeo29CkgJpJkxxctOzhEaAUDc2PC3Ni5PbtrW6bduJCjtsO30F/oIyNlJF
ajeMe6vz0DNZeA3uuO6ZyBHOPpXskNhRSZqiFkDVdq9Swrz3TNpOc9GQIFlrZKCsh2mgxjRY2cpx
+cWnZz6IMMYVj9f8U6scpQkROy1qPdZM39d3LuMmTuwJRVAqsXHK2VesLu5o+VIWfbq4rJPVtBZ+
rLpcnT6aqyJPC20kWqiCvpdQf6tb/N0i4FtTJ9OuYY9t/Ocd1rYDCsn6+RVIYXtcQVkgagw1R9jx
fyINjaCmDKSPc9mDepmNDRDERqlDksj3hqheedOfYqGV7Ao+Xr9S9mahw+uy1YTIW0ZGc45Z0EeO
e7FJD/sT2/eEBk86ZWIoN1NaUj6UQbQYAAFmFULpu+008pu8AuG58OYy2sHDXqdMt0/A3Q61a3NR
EjrvvcLGWLLwEzm8pWS6kqiSaMlk2OvQoUaL7UAhSAMuT+wzWGF0GUcmIjblcoIhcgi51UwgYMqk
XpkCMP2/O6c9MdXK3DjIQyFDWjDgEIdz64FJw/WwMasj8OaA3REwx6wlHH6MBEZq36shlIPqiMby
zdt+K+sv4dei0AlyGYfp3gMpNVnCxYEPjF6+ePJUogtKhsZTGuLB96lKd721E2sr1TyK1fRtQemh
p0+PagYbjtv3ilAg8fW3Mnp+etvO8MJ9ovHgV0UzezXCdzEbZn0x9+4GNmhesPRmUVgt2ry3mnyO
pRA7mvtcvlbX47gILgt5QVWjJovP1X+9oVbb//ABhYW6jw2VSf9CRjLCq6/uwSCCaaqXW1Q3SvFZ
+cB4POxSjcXnsukeSsjcf/beeTe4cgQZG6cZ38ei5VQYOOXbFMubdNS6+kGf5aEET/sEz8CO+tXs
FVuquT9XCF02MhjID82A8H4tvZOsn7l8ueJ3UwjiYFW+i6DWTIhiFtBkV2zE26T9g/5pOeqvZnfi
0yTL7Wlh1mEomkgLraslcGeqiCmrsvdt2aOASdZ36W7VBLxmU26KaXCHJ8ap4KggIR6RNcyjzHt5
Cafg963eHEN1tQxmoYobt+lbCHG4Vs0Od4LVoiFtm+Ens+bp1wVdTIC5cD7ETnjq102zR+h3pPzU
6gB2XEUVYJvb8bftZOudDWv0AY75moqK9tSCDRmgN4HiKBS6bUAp6mJKotxiUQZZvsBBA4XgucZw
gSu/lm1Eislh9kt8f9QJ5l64gg3l2jWS14LjW5GIBqZgACBZTWQcY2+4cHdog5miyRvkrrZxrKrw
cbgdlZEmsfc0x9Tf0GEmCOsKqZBNEPDohHGK3wW30N/Gh14/vKC7b9eGlrqmRA/pLByKGUqRa4RO
EayBgbUaNxIA2lKvjVxjPCyPTQUGP+bwp5/6JYD6TFWhlxehnKyJlppjKJbqWbyGQzsB9WncJMWN
/hpSv6BgK53Do8+HB+3KP+z+GvoM4nFx9JsFmlLGAtnpl/Eqa9d1ppD26OVgeP5MYQHiD0T5a6wV
JCzLlcEoV55alOlk350wPqxZpC7XHnbkkNhg92yVyj3m6VwlkMNZiWgCWu4AY3LKqQwEjYTi3aUO
Ey2Yq/el/0i9unRbnoE2qr8YvC/e+l/jhi93uJptEvSdWOtnMRvvUVO3u/8ostQ5eExcmiT268yq
iztqmfOHg+fHud46jtoMVOrvGaSVHuxFVejHcWpteLimx/gN9r1BDr5pRHtgNyGUUR3lGdvLr4fQ
pPK8c4Zs5j6l5RScl1UHqOAsTOvSe5plzGu/1aAtyh25i8dLHVMYyQVjvVjIlr+pbhtPfJK0YJ1l
1ZjrW5bmZKPTDvWk9pnLrFKpShjXszt03F+MJVNFMo+5vmPcHZvshnDMqfs9X0Bleu4tN163cyE6
fVCzJ2k5RM+F45x70FMNg7UZpwnHMkdCRZUJTBPfe9meO62miKrmbaJt7E+H5gNtgnW6U3Xb20l7
bsAKZcoN3CHCqSsv65xE9pzM4hRpmXxhbGtvUNlm8Y8R98R3PEDGRDVie+ml8Qrm6gGW/LWjYL//
jgcG3/FVIz5vwVVpI1Ac2WQcQbG71bqJZJvhkaRfsHl2jDkTiwvxZyujWfA1DORiONnwp0DHnuwJ
PpTIasDuh0rksmZYRxDZ9YBrUPVYDk0ljegDKYoO74InphF4UediA+O4i+kzeXmY6ih2jWuM6UhV
7Ffd8+B0L7aoc+sBg0/uepefImRRL9JQ7yjaseERRsdbKzV1QPyt/C0zFPRjdW4wFPZMi+LfmfVk
/Qc/Y100aItF1oJ82T0nxb9XH2BgV8w7zzhHi47GD5k9sOOvtTJmP17ouAu+1DNnDPi2LflSnBCz
0tSa6Aqg1ISYTGiBNMQVv7++6vsJpD7IyL8x3ALgmVTBa5WEt8tJJLZxW++T09pZF3aZcX67xpVX
EoRhiXL8lBmTbkUNf5ma4wW0dVPvkcVLacSFYsbLMaD6+yslgTKQ/NcbxuK3t/f9CL1rqboUB51j
/wj6nkMw0lbxMQ+HR3kb8ngyX/gwegt4bdiD7v7m+okxBdK34o5sEL8Cknp/GGpSGcq+WV4wKgya
MYrnwDwUMsSnL4jojNFvJqlcbpp/N1C5woWB9YJK4qtJ9AoVIwZ9bB2/e2y7DLna8YSet/tXPBdZ
8C34Y4V7WTZkGivNluvEheaWG2DHGKYDqgeWOPRWLRPnCu4l6y1a0+DKfJpPlw/dKQX0Xqynueht
3WgQeuKn3rJCKilCniDxvr5VXNnE92n3mGOxSg/tIcwp+fkqfvoq96ieelAia1f9TeV/ypQlqP6C
DRJ82kvuDTZtl/XcDV7NNffrcS6qyKZ2LCk5RdIVN4jC/6xr3xApu74n8ymdtGZAipS+ICTc+pX9
gY7+KPA9sqp3AP385wJcXGE4mFcxybraW9otqj9egIJ0e8Y1CZgiSx7U7pTT0AhqmDpqE5r9qMhd
FccXCWpo5H6ZwyctHGEmfcesNwDZnsxFVILfEkPVvuFcGbHXzZh8uySENFelYw/WKmK6i3Dy57oi
lQHM6MODtRySsg7L2PhdgGHUGH/Vr0ebeQ6sgJ5h1Vt/FmpIlEnI2KAjZpAG+2KGCi3bXxi5Cwef
P+M6f+oKc+76NHxcb98w63Ah3YoA9vJ8nFDP5SfMSFRG+jQ9COteARdgkB3a3wlKYajYPi+eQEAI
/YcGj2dhoiOoNRe1T3zoLpCIPLxigydDhO0cWxwTu9ry5xLZP66xUlbKIlMwMZSTsKXi9j3tt8DM
B3xI4EpjUxv98X9Q3oqn3m+1iL4VpdkkjPy+s6Y1eE/TEIfyiCoAb5JtzOP7eNzvPoxtUr7rQRQd
WaKXzQu9AKc66EX9ze+QiG9XgxdC34hgnpY4yEwcc/HQksHop2RnZAGOo0URigXfEf3tEneEWMFK
eEv8THHqRHviL+wUoIVw+QNh1bKo8DRjiEWYO4KICIMxTCgiTQEb9aV4z6DrdpTPlIjZeuWvPV/e
twR4haDYXPZZRYPiJr9rxGwaSVNuCnjgENdzJbPQWVR5USEw84A19XCfGGnw6Soo1iQoyoN/33pL
LsfyfCV0lgkT3TUWs7ZpXGeQPP0w5VLMs6VSEQBP3r0IDCPs+vKYGYF9AAQFxbKJiOSUlG2gVigy
h7Gawvk7NQPfg+2BxtpxpepPwpjq5DmqVfrPP5/trl+D3a9pEwAEttjyGYsSMVWuhi29gqKWeXqz
BlTFN3hdm+3itCN6RDQ+Pp8CYEaxNV2FeUBy0zCwRjGCHC9tEPPzo0d/NRNJlQFFil/WbpIdh15J
Nj/3WJb0GzlgJh2RKDcGRiYSmxbBhpRKUX3PdfLIa14tt9AnUWAZoC4MErr/YWJVMozOxbnhSb28
dgPTtWQLCV2Nn8c223VsxXU8K4rLmeGGqetf3hCx9w+QRqYHFo44YQbPHaVZCuexei3iXkpEuahT
OIY4uYmfsKmP30Ti/hieXUEj54hmePvl9nFehZi0/TCcyztiDxDOx7MPGMkssoYsAGH98QlPIljz
ncMqP/AO6hqnDBKyrA5+DeO5rL2LSZk6010orVkkTr66o+liAs7Mwy+XT1LIae0UkTLqBCwH4PzE
J7Q9+xwNdYlXIrCifnezvpXqMdOoVsRWKCCiogJXz4D7t4tjlSueVrmfwkRcG02L3geH/HMrDR54
ZvfkXwkQxc2H4dA68ul5Tu8smZWIN9iElIrpQl0t/ujZIOK8L8xVTOBwx8Q0am9AzHDcxUIfIn1S
e9s+DresJy3hDj9hVDLfYZ5h48UXyOGucLUoVXvgUZvJz84d2IZAWSXicFHLgimj+eZ4YGvnRfSr
XY9tFuadjsDJFCrxAOq0BPQa1wbJPJXd9zvx3oLhRcAsEx2ZP7iYTGyJpwTTHsZBZL/6uqRgSBrG
YkpNKJD10O3AQRJzQq2LSDfu/mUFY5D5U8u2MKNnDd32cJNc/+waJDarrjcw61c9QpcX6LYD2rH+
z73ib09hu4zF80TrSrthSi5OuUZNAnTbh7cyogKPCMHFTDMwpkdZjXfL6vyTduLIczg1Wf9j5+oh
doQ9/6KAXU9Dmf6yHZo3ZDzXipFm5YgvnLOHfbrDdx9AYLe7+Yf5KII+gcww1h20eE36nMDcrCmu
75cTMkSBISsps7mPttVGKgLp+J10Rmd9BMXmmQ+hQnGt4tLuw+I1je5yta1e4yKYv5ZdIgbL0l2A
bt7/L++07d5rDo4i6dukhWP+TwgDatNcOERf193rjY3LLQ7aC7El9I16Biw9nx70pMtlpfPo0HDm
U4UnM3/aUSSDGzMfNCGcGi+gTMViY97dESjitXHuRwtzpwz+kAPX15q8XZG7z219Y3V/nRwlyw+L
9q9kN+EBCEof4gMF0kl4gE6VoQg55P/ZAjzjlnnjMFNyCKeIEDSgnqkif63SnILxRS0/mY6j1zQB
dnJV9DlAba8EYBDkWwLWf2n1+dYrm1QRJYQkGKKCUThnc994ACNIkMo6A6gKVswzelAaYyevHil7
srtffa+OGKZWH/jGCmd6rmVK+NK3PkPdgGCKaAh3GCDV1/84BkMcl0J6ESwilSkkYDPLkm3VbYK4
rloOQ1k2gt1us9B9fm4IwWFUQJW417BjVxZKIsJyWrpSqnqO02ZVE6h3NoFqDcwIcoPM2LQ105ev
8bnVyQY+JbytaQggctElGBV6daNc4vRYQ0Sr+5kCE6XZ5snEbeMixZKqMpz5ER1YhxPi0C9fRK5T
FXzLkDyHCmR5Snaf8MKcsLfvX3bn6vJvZkfFsuZBr8OBr/1gFGXpjWH9gcfZOYqCFYDzAJ5qHm7D
Vy0Y17rKWm2YwjOUZ5lB9+3W1CUF7v9XGIV9kZt/gLjikwWG925P0Fnnt6g1R6eL5CRKy1tL6f5Y
nOwZmtPKNRUSDwjs50/LNBC2UOwho8wYJ/JEgsszL1IQKBBw8pYSY++KkqzcjKVRlzqQaGP8v8um
EJTsaHcv2szm4LdA1j4Hr8syIfKHn9KYPWtm3KDiIIUag1tCswakMbl0ImivTm0d81qrfGryObBs
hGJb/WZnTHJYA575cjMsQ0v0XplGrTLNVUbZX2/WsnAf19vmTaAxyDVjHgSCT774hXgmhcqdMhg8
/N1BqSz0+MnrocqQTqymueCoj8mZSBaFdMmjnyr0SZsQvmY6udsMVG/EGbJNf4iIzIX90RHn2BC8
Jer4E+h2rxV5ZRE8TExNIYwv1Vv1NQr3MyZo7yarz2xo9pzfV2K9xlS3eLVgTPa9uEtxhBisadni
g+nusaXfiVBq5LyAvOOeUC5ibhtq77NbB9mwkSR84qPC3YqdgNZlV3WCZnggkU7TARMZF8j7+VF/
fOMuDBMJDqLOlkbf2dBCFI6MvPip9tY2LUWC3OuTD54JZTGJhLbLbvREijxGtkeYWUpCBsgQ15DB
j97sgkShwcq1I/H7RrFA2Sq0DA5YI0M7khXRXQJUOHoquLfFMN+E9IE66IiTmKZK92vGqmKuOZGy
zPDqAmSCrneGY0WWuEVLGdwqCr1m1o0QxW8RV6J+enYIWeIBzh02bw0KYNLFFpALsjNyk1w5szm2
qlXlvAJ1WnEH3qgMaEovpw5aVn7j6IkP5I73wTjaacahMBJsUgWzhtMxdr5V3c8QLvDAX9cz/+CI
e2qRD1PSy4136DXoK/iPPh1hRp6lSGh3VqDz5hG5ukeekJHJWyVscY3LKzU3B3SAr08UL/L9nwUz
xXTbsXkVyAHofteuvXB83ns9uRAdZptRKQbmc6sy9EF+R4Nz7/nJlD+3W4vAkrU/ZNk5EKnvvcWL
XTFLGjzLDpFDSq3E2u26TE17jGAs4kIxxFYZeTcJKwTUJPNuU+McsYYxbHAD6liChoWiOzrUW/eo
06+ZkoTmg9VEBnQk8ImLKB8BkPbCqKhZXXXZP+TjzMPMrbtXg85F1ffIrMdS7l2uUDuKpILo+vcS
KwkBx1NhZd/a72AjW4E5sfS9iKwUZMsVkuwdvCCAfBhdzeEMc/580M6mYFudlcd3bCI/Df8JpJeq
1ZNk5BxRVMrvBpw5thkKALr1apG4raNUrN5GgHwM11gMOq2CvSwc4Qdp9PeOteLju06YOqLYzp3Z
+hbIB4SVSWSd5TImEv1mxL60VrnGXdPEH3UhQvL/KZwNv6Yv3UkdxYkWG75QCHuJyTVhh27nHXyb
vY2sjpo1QAkPi1grMSTmYLOVM6BIJL3GMph7eZt6dI5KKtiLx7QS31P/2EcbuN5wcCS+nYyLw0kk
JTm3IC7RsA5h+NbE6rfD8gNWi+/vhi698AhT/dT20y2nftUYbto7C5HNk6Rherh7fewWxqIYK7tE
T4QIsX3rXdkOd+KjAJhZyyUzj/v8JSnf3vnXjyWqpBWnBXyuMsVmPnTgds0jIRfc1H5KgWPiGO5a
VGU8WqZsIjOzebn5iyKkNaNW9USWro4+McqYQ29VsM9CQ64JatVnKTtuVMdLHP2DJUXWPNgVlZx4
hHmB4qMVEUJwf8d1+pDFpqJQzb3u09pdrQGMwIISqtSHmruwipK9AgyM+zQ0YBK6c8gblDp7+P7A
U6DWt/aLTFL+inP7XSfQw8xQUIeX7mdLVVLalF96O2o5OR4IXWmx133f6U0lDn97HIl0fE8oC8UC
oy28KEWzk0wcpgtS1xPoFlEcW4x8ZAitF2cc2KCwoKpYNT7ZSf92LRuBW+we/PIO/3qiKpxCgkO4
RxVxIItkLqHWhnS2+zunTAYxu5zFRtUUVWzziU1PR//FcfCP+atpvaqp+YDV3PVkr0aI7rNspgZN
ebQiOm5I6U836xZntYOLLsphRMg1aMBdtC0Rtv+97dJAUrBl3GDMgoTSL/wwDdF7w6tgac4J1dWt
zr+kP5W9VMoFYeVb90eDSTgwxmGWVMzhjVzDIwOlISZGN7ZJVqyCDAWpfgVxA8XEtJZZJNdn7Kc9
bspZxiBpyRsFQSaoo90oQO+WfwJsbGXAIM8RS2Iyl9QbJ7fPQRxU84dtkrijLy5r9yYmmi5Dur3s
FbECfvpLfwbBXUsMH3sREkUrHhtJhSUyOX8JaCRLnL2vKGY0TRXIAbfZpf6xr0bQOGjZ1jTrRjtK
jmTrph11jJH+XeCNbhTJObnWRj3Rgs0lVWL5aXnMVSR/LlgaWEDyO7qJe/m9odVNuFyV0KZhNKPl
MmR0gfJiWoy2Pm06TayCu21WDzTVXqZHCbgVtxHjRF003G6BxHex6YiRR/+AuC7y3fJifPmEQabx
azstU6e9LOrr53/C7t9TENrz/KuU40u8VN8SdfmnE/v3eS6CnDsSyTwC2zW9Vq2f5YPNGARC/gRE
aFA0AIDLHdqyaJJqtSwuufySqbLa2me+MIYwKDdSwW9q75lCDihfX4WbHHTV0wNxFB7EAvn584Ph
eJvsypVXDrcyLE8l6JS1cyqzGtXnCYiDK8OO0BGfUZBkrSJ37/eFGVwjvvMubdtGfTk0u03Fwa9l
0vu2crSayOpj+44tGZe04JW+NN2VmbxU+UI8gkC41EJplurY4v1wi4wX+k48eTQjbQn0dlFM5IYk
F7PFx8JK012O4p0TGnUWGV8WI2CPLz8e6qWb4/kBwlXUppuYhN4CbbxJT2AbY4ygM3tURZCENiHj
adUKaf3y+GfVk1sNArIkl9CDqXxCUlZt2HoaU+73uAz68hDG5k+/tq3tDYx0pL/uf3geCvaH3JIM
vE/51Z+lLDlfOAAWXkUQrEgR5t3alsmrYh2VZ5k2lTCDZbGweCXI2xQyfdQ1AkqCpeD0dfiMwAZ1
vHp9kYNx0ovx3JOraVX1adnrIrUdfGOAhMj7md6fUw9RUKqL4uQN4p59rmuHUddaAnW1VNWEsdbh
agB8GKCJF7MXIX/yCsyXHPoTcksYhqma4J8yijePMjdyKxUYw1PcFZ7u0oRFrvSsATyfwu1/JRKW
KGmQ/iGvsYCkNchR5h+tQX7kVoWl4G+aeni86yQELESOsMtXVl97YCsgnn/Oi6ZvugnvJRZzBJ0R
26qCNvVUf8rUVq7NzCQf03+3ALydtv367iEnrooX/UWLVJu63+Ekz+zsDtUedR7FHV0+aoA5rGia
M5f6Y08UXC8JkjFm56uY+MYlBfi/8U/U3XQRQr7DHC0EnNd39gbO97lgxAFrqGqfzjkiz34DRi6s
FL97u0Ar+KZzjyeZQTPZVY0maHTrAMxRS+n0vHPseJgm32RidrmJjgNvy0ucgztrgW20BA9/H5ww
XjBZW3/dYjyM5z8DJ4YkhsmkxPkYBIUEPx07GAiydV8kqFIHZaGMHLYHKDxRTfvkMQvQWI/Xc7zN
PUr0Uo3xgu7QTmw+fTwuQyZzULrQeV9fo2AxpuJGAcqEsFJPQ92ruu76BSQiatm/80DgaqtUZrje
wSPNNTejYoG1nsC58zbAYFgVxj8FZyfy5jpOyDd2a3KdCdC8Vtppd45WNVmG145pTKWKs0IC4SaG
uEKb1vQh4SY6AXUdEvmNbL76fAHMfUiZd111lFxoQitZqCXW4Eu6G00WbXx08E02tNzp2BB3Z47H
/EFYd31Iqr3ToMWgp1lbIRc/62T2EnpUmXDSLH9iFA849fVzSNKg6Vf52iHlhRXLuYfLtQRyO0KL
IhKA/15Nd5XgipiPOIzYenBqATBxN/OFeEr/CzQjmL+kPOuENzkAsOhf+6ZzFP+YjLK1qcZsPnMF
PyHMvlBbpeCRuIkbCqa8MAa5zVOmzYxZb7UHTiDCDXNb4cwlfsG+1qjOZQ57GRhK+vfFp/OFt2q6
R5CmPLTDRxlLl3qphKUMXO/0Uo46tZfqn/0cHyOSa7t9ssSTqWsl1RgMWzOQ9tzoye0tbeLhtw6c
e97cmSY36LI0OFIWC57kcuyeTnc6OYtGtHTwGH/UbQPafzwVQR+9UBol/nQXi6712YSX1iw+ExZO
3JYOrQMS4K2BixKSh1AejAoCEbKzwOBIzIVpXkY8bJQyCcJfLJJWfs1Bp1zS3a0yqj47Wum5XDe+
G3+zbI05hL/H2jHUZEbmk8E5AZcTke6tSDp6ZkxSgA7u69x1D640XU8il/VPeJknk/1e8MaTqIef
2XXT7RBvQBQ46UHuSXt8WJKd4WGnBJMPz7YyDiVK6SN7E5tHHaFDLGN2ldLkxsFQ56gS7K15RnfB
d5kX47PkNPz9bu5Loy8PUNxm8tQ3OdnMac5FP/JNa5VG9wNBxSBf9D+LxAh/OK74WVzh2PHx2EaZ
5rKwRc0+TwLmkjJv75PvYiD0tqOXOI5LNFqWF6RHYKEhB0yZMEDBeh5cVkXiEGK8PBqornXOva0H
Q+QEYil9lG9kpnmdI79OF0D3V50SkGeDBM+AjRPJ0FZt3LYglVANiEzs8ys7oUuSIT3toKqemFC0
cZXeb4HffWMVuNsSXSFKtI8d1liHqx12B8GsAOJKqRuHcIEsIX4Yh+GHOOYnYKYt7+TEyoJhq1fo
gT/8rZBCnObbEHqWFkt0T9at17h4TfBDewXzeLcx3p3eXrmZoO1I6jhP3udkTrGMiplT0y/qDe8D
GKgNRWStSW8ozaAiHAsdzWgme9AL2qRMbQlsyDydXrUUAMpmleTAG7T8h8fD2qyJbR5vK1grbADa
4Tu1xwadCOhsC06zyEccs9DSzrlwe81WgQtQhH/B9tQmpTp9Y6pUhTTBBBZCnXPq+78Cas7472Jn
DlJPJLmj1nKC5r1FseJasGHLEpqwp292KsFVlyT8B0kIqeFPBTBttIuCNJRuo4u23SfCLtiQZD1R
lxtIZgbFQHqK7ULHv42f/e0/DE/abNEKk8gYqJK4sFpnGu5bnhvtxX60eXs5WKRQUc9T8YQx/3kD
UUpY/gcsV+UB1SVFm76ioX+igveFilHAj26L34F+TZRfvzpOaChWIQhMYnxfSSVqySMp5Pnt1l7Q
C6Kqt1RicZuxohp2HA7YAeCkemFpwRQumjqUcJW7VkMCnRzssyc6P0KATkCKUQkYPSdTnlhhZMbf
rGWS2vQRn1eXNHx7dAEyLcccJyJqZqeiKAL2NJCcTJX+FAtQcGAnXaxwu+HpU/UdtLo3vFGTKUfO
C6bvGmIa4sM7sU8+qnb9aPCk7h7VKj2WiRaaOwbFb+VTd9YEiXgKk0uQfb+PSCqk9KJqN2kteIOX
snPYCLhh4F3Qo5qDPip62y1HgC1oOSVaCx/K/9kadct9KQ6NnnIzQfUmLwuFVo7y5vDmyQRG9ioU
hjnK1W3V1D8JY8Gl9JyyAkJzG3leipUi2P5hSFxnzRpUrOf3S/3hbebP2fouicOgShv9/huq8AnF
YXXo9x404rJfLsGBFiVETJstE8Df3iG+PoJfTECKtwhxzoEHTsj1qEAC9eTOUoNiTn+rWIg4ti/p
pkAU7Q0Hgl+EVw4RVCyZEFcVeFDICwK/yEHzzWrxpzzfl0P7yJeooraaDA7lHZPlS47n/mfq8a+Y
4IzOwZiX6DK+Jkqwoynzf5LtHW6cJ6Bl+eHvnpRUFldmNccODZiEyJ/rSbaK8+dXNtL8ffUL5Lff
PTNiQ/5xeHRBU6E9sQBWvEUkHdAMlVYG6UOOlYQy6hWcuT6KPn+9qgRqokpmi7F810Z199hQsfo5
GMmAfh1Kj+mkeOXa7p7BH1tt1B6oK6CscO9epeztW0KpBGYya8sn3Nk3AdccxzX+h3b4jY+issZZ
Ap18pueFDP2uJocSSLBVH7C7WpTL6+au1/lkfvstl6LscOyt4Q1/AkAVMDx/kA+FaiHtotQjmEGL
s9fex7D7fzucRrHb4Eib4g5xbMYW1Zgss3pcMm1naSNZwVrTarbalAH4Lc2bmxqavPgA6LqIMgYR
uvHs1uxMWuLa9jKYlhPPOivh8iY8dESfKhsNICsONw7CWVLQMbdTLHZenRkFKwvmL77O4SnihhXg
fpSlsjrCH6CCo2PJ7oUGAjpMSIJxDCIShSwQ5o2rpemGKHcuGWCQZlwAtNBbKiSlQ9/Z/rTAEjp5
GaDS6X8sjZBtk6jlfQ2i2aGAZIjHsqPEJhytKqOn0ukKbqwK2NrxrzOgKyfF45dhdMbT968CG7di
CK+lTscOLDKYBm8aOA9cnEO8yYyADQTcW1mSh9qwSp73ERr71rKWtzHfr4YI7Zg8G2kYvw0akBYF
P2dTHlcbeV0eAXx3WwjFK+8acxO3OKnKAsanzb3eLVHe7mlAtbbelLH1RS3/Wjd57DObXuiLAqeY
M4igMSV/MnYyu4T8kENdg1eQvZLyAwUqaM5byec5KS5DU4ZcBM3lfUhdVpZuuDKnr79ddkUiM/1J
A2oVYRT6dNXCrywEjxMV6VTjzbmIbJvaqZWIU4LXgKjpMKSIGR6dx2GH81juklWS/zLT5THk8JrO
vxWI8L+E3RT1YhHLbUr98jW20uOJZ7CTBClzKpQxiYCQV/vSJqc12o4vgNRYaDDFlBM2croXT/pn
kqiyQkZw38eyloUK+I/B1+q4E46mTs6XKH8Wabgk6tm7q/B+tR5CssRGdrPI9vZpm5M/qFVJyOxV
98AZ6IEy/7cgj2omZfuGGFk3rPRSQRcRlLepwhj4kPZkqOk1mcmVxrrLj+VRC0BjvfaKiS+wLIJ/
UJ5lY22YkgNHGA0juv3TnpDHlepP6QnIfO8lhIR8kjClSXpu9WKT0zdSpe3zYokDggrnhT6QU/2k
9re9XIYD++jFefGmbFExyFZoVckUs0IB5QV5mQGhmw9JJZUZs+QTmINzYOZs2HlGehZA9g3Iw8ej
y4CjJ1Bp3d90RTPvm0fC/zl5QSXDG8Vw2WwVTB3aZy4s8oG2N0o7dbjXAelOGA2uOKS16g8TSJlc
hNHMV0Dxg2XnOXgxOtMNMaa7K01nL1jypi+MLjmqxUrnthTx09YVfxYa6KPYOLllRt16QDM9OBji
sSK7cONkBcZ63Yogr57x7oQDQOVbE4Oj6SgDgxG/896gL/uk6Ynjz5ZftF/RmW0B7LcgX/I1EOKn
a5vGwc0vHrvJPndo0ODTCgpMs5xFjfAuwvmlVL3WUL4PnaDnM+lP+aWFk7d8Kpu40C1O1SGacCWh
hEiUl8dIYAG/TVeQfYouhBF+xVRZROgW9Ex/zsDTs4JqZ2E129S2ZsB5OlMJWDhiNxC9BH5AKiJv
EQvTd4egek9+TO0C9FZuC0IsfzTiPs/L6Db78vaWpGesW6hbphqOerpVYGHLtTsKPHkm6a1NzMvc
tp3dY/B6uecypDrbnGyCfpgEEeY6XDH7Z8LLieodRwzlDhekkec0zb6JfNGVpA7xGUHChNv6yYpW
YEXG51y+NVY5Z3vYBHbtWf2Q+qO6ZETFuAU3kIXQH0slwrxRK60thzxzbpBjU4k4eZDpPwp2ofPS
n2EfhUaW1y7Vj7xlhgVRUsI1dgcKPWSqrUwHu1Ipx94rMBxP276QemYLIBLz9ZTfa7IkIE5X08XH
MWU/5xwFU512iTiYJcYHWFFaoLYIOaLjp1PH+fovm3sxMh74I2MKoP/UKY+Cyhj/MKMj0bRrSESg
YFGB4Noln8wHYM0UnZSQ38XZlw44hIoHa7Q7l5BAsgvJZUfGiS58oDZpFWIEqfNO7hvT08wA1j/P
Mf9h3Kba3Q6sIEV6AilXK6UMmBfhXSUyK7uJOhgCCmDTWocJ4LikzGc1Wqmm8HjBIPW66Zn/K/Rs
mDuSxobKucOgzBNC/7KJSJwtYD02ytUVruil5dbaRVQIX/FObbNZshYWovogheFCyoBtihobqrAL
a8dFvTBxrNwaHiwQ8VSBVWlKw0rW6VG/NRcudKFtFYJOCmV7l54znURi5ZsceBDwPS8Sclp/MOvR
Tphdd+MD5MYtZAeBB9a+5PW12LYYDTOGC0d5vaFTLOUl2B51e9NciyDF+8BCKVAXCSJWq7gSvOeM
kX5cHHWHiAeSegGVeprkZdjR+Ft2Zf+6QypP8n2NwyZ1jobJ94p+gFNzJwHyrKwy+S1X/htGF9Ti
SMNkcqYf8fWGQnjYJ/e+iHex1332hshWqo52t1ukslUIGNQACfkULEsnYVXm+wROoENzHx1UWHET
HxPAcyPXpUE0A4Biyp6dHXduf90oDo2UiYINpd2xLyTrrcgitTtSHjJ/eNC5b9g0InkAExVxqlEV
J6K805lRcIMeJCODW4ijQr41mGqoOkIQjRw039GEtXCHIFjpLllbEjD51jiaw+Su2Ylrp+ulldj7
GFVpnh+QLTAawmLSJgtrMTGj78bgkRGpCer5Tk5sqZFcoYT+/Mkh9bSJY8FZf9eGnjEecYDFDcz8
PQnD3CA58XxB+CaWzb+dwIGkzrWVleIToWHqrg3THbFPq92UE3nKtUtZsG5LQ/gpgm3iNFcOxVJ1
cdabmuis0xILyDKoNbtpNFWAs7BEeX/+bUCuAQM23khuzwdFf8EEsmRr3ncaCIBUTWU9G94IOojr
kAAjYb9DTra/imLFKY2bdIEnGGfEdt3SJQPI0ImyeUSAptnajgheM8qMJeIlrMBKMF7ZASmh4G9H
hzKM4hQs8WPxmPNLLBRx7EvxWnb15xLlAoxel14cwmwySi7q1DD9rojFInFmudgT7KSXn/UD+lyO
du9R6g+G+VuKcPqIdpGKtvvTEwLMwE5vy0aa9bDoIunXgI9qrGUZGHsZnXn9dANzBD2Tdjkg8CwU
Mg4jfOoydOXffBiKT0paPtE0vIGP06n12ttQeCwZmR4q/WYYlaxEakRUaMNCt25r+Eb8um/u+4i+
JmM3rIeyRzaY39Br6mr6io3/PdTcgetCaesoII+2+wEGbP6ehH2Py9UMSmTNxdRKMT005pezAddI
8V0mcBq0r3vi3mfmzd9ncxndT2U4sCfPNFk+BsZww6y4j7iZlAKpwpwpOaagB99gKasosU2oM2CD
EJJUwLnb8wLRayaGQTPVeLmO8ixpvzKObmtMUZSQSZPEOxEKg3yZQ1T5SXx3DLX7205R3tZwH/nc
U96qUWcqxJItoZkqBsNKF1Htz/mD8z3UHOENJpUcpW45btZvK6qi56diQJH8iyWt0pTn/419xfnW
x1Im53UYY/el7tqCE8dtiCALfDq3jgOlCymlmI0xWXtishynELkTwdtiche/zmcr2Ic2A8DFujOl
Dxle4yvAO4Ky+X2HEnYHhudp4w5tcAo6OJplE1c67NfjU54OuNOFfghvqh9bl/XiX7N5POAuDiaJ
wywN7cyqySoITHVEVaGKwDn1yL1UauHbp2YCQwK+23jOUiCJtDuf6r3uUGhLllemsYNGWQp+ofi1
dSwfJvqWCyUhKZD+scqU86T7vqR0HZjUames4QcNPPniXwdCcohha4yl0/wttgv0iiwF+Gb7bbNN
8A0xDCfvIKk5hMqBKsnXRLNKaWyfdE1I1W5jo2FvXQvGi+Rbbq2upAyYZZmUUlBidcmFss+eg98h
AXWPD3qtgvJ6mtFRKflK1thex6kr9dyo2XchUCMkgJVq+txMwysSXxQ1eSWtmXYe6Y8YTmf9zd6z
+gm7cVc0sK13MvVq4iaw6YB2WszwecSaPVqK4tLGoQv/66DFlkFglb1q3I70OZoKZv9NQKkzZh2e
Szq4Bn73rbgOVSPvituBgE1SKQzUVwfJPmCPt5QlDVquiavwoMwPOandfue0qrSyQV0BGaOWTrXF
VD/UClMT4d5g8tPvg+CNY9KXhP/8v6X10OsTqTI1uvttUQovZHI+OG3PcZqyKAyCdrWF9JFnLR+K
LVqAIeLzFhUAtokJTCDP+MX0wBZrfdKOLlZNGtOP4614E3fNBwOsiipnpdE3iUVBEXywK/owCMvA
YRq5neTjff6Tks6sES/+91M82l0s2vsuzGvOqq4tXxWhuN/3KuG2YVr3ahABAILmYZ2wmWKIUF5C
SzCyWeqGNQWd/9srV8iyHyxOyXnlNvVTknlhX3o6xWBvosxqxh3t0Hzp/MQdiCAms2OccKUIP2//
2Gd1G2vQ1tSgNODCz3s8cLtO9MTFhW1N9Pz2Nz5Wy4fCMA5H3fQ+JqTlFiL4cXJ6El+A9nmf9er9
eYC3wbJ2QZYISij63oLqIhauYhmZztlswQCNxYkN1yqMArCsiY/bFMtLDrFRnqgTeKM+mtdMVjqT
y10IViTDFbGYshV4JR4VsXryzRNjb21mSWHgF3h3ArmKuHP6EoujiEJAhj0CPjShu0BuocV91KS2
GsPn8AbfNGw1wSa7+BzQF8P9UCrI1XT4sPNohfmHw84gXxmmDl7ngFzhcYxR5Y/EsTEPWsjQ+jZT
lniCdPJn5wSqNSustWJnuDGQxTA/dvPo7Wf+9VoaySmvKIX/X+6ghA0STOsJxf0ex3Ic1cHdcGPU
4Q5oU8MTXdX/D+hp5FNeVlAXLkp6AWcNdud3a63gR5UhyTIW1F1KKDJncoZWW7MlNadKt4F/7DRz
Y2gArqdfOIbvetQRr72VtDpBH1FaOCu4JukRll9bYXUrsmanCdyiWP4wKk+Wjtqj/Eo94jdY/i12
+/6tRZD+OaUAjBZsP1DqthjHiYlDqCq6I0MK7SYp6UOHVQjEm1d8pRTUm68j34v0vkKn2rMWF7uh
On66UIQBK3WYOus6Yq4stjgfQLOWqLfqNRSqlsW5tZg2MH0ceDGjpbmVylYJO41RnD4WRgcg9/lm
hXEtIHbwuqAkGjuXSCB+KM1DcE7Be7tcqeLPcc97Ohs7tgmgCn+AYYlaG8bSfiHWTDnxYWiR2cP9
FxH13f7XzK6MvPe5ClPRxA2PsjY0Zk3qlE4h/9l0WuZ5/I7GXj7ArDF5bYBSHn3Ch934CQaGhyA+
LSYApaL22pMOVyzTyC/JbpSED2IK05rIZX7+yGqVUlXHehVUe0UKYHOd2ZeSg8daEDHdfAt8a5Lq
U0hirybjXb2RnR3/VBXtcTcsbWJW8cPtGvWGgEUWqNWKMCLt+1pWvW9ODoDHYqVl6MPuDxQLXa23
xpUJ0Hhc4cgS96P4lnfRwNFvaR8/2k0wF87LpW8sScvYJaxj8vWuRBH2nlV4b5vidUOCOAN/ZZ78
lMXmz4k8/qGh1jkUBu+FcTemWPbJhjl52pHqc9+npCejfHhhjmONNoRt8v03V1ae48JqKh1FrCRY
WhDrYzX7I1fDWaLiRf/KA9qmkLs/ZWDFbg30Ul40NoGEfE5LNkMb+oO5tsyYjArrQXy24vLT0kHg
aa1zIXE+bvUaFsZ2r1w0nxT7MaYYTTU2oUe7+MihonrCDg7evS8LqcvuCWo+3o4vlFYKaRe1IPWl
4uw/1aHUCeyb7SXpCI3qDy6p+mzXMclg0fVQOFGdA62FZfzS8KpKBEFkaN/OCPQq7BajRv84AWfr
1/8Oigry8lMOGaw+lWmY3S4a53l1i5RqZnw/12lrYQs4NNhtFRrYpVMg9FDqEonGCjnGr4mxgCDK
+nUYP2j7Sxfb7GGFotn2x7bneAJdbIfOsn68wyyF2Nnzh3Ophss7JgLZdLMzzRlKVErv/tp1a4iO
mZ59ponDJj0syVGl6iQix7ZlHH1Ar3NJV4SusGHzTMIkQ2++WO+F6zDMJBeG5qBiUQ6+eOcfyfTJ
f0p4t7+EvlL6bh27zSf23Se6OyDtZMfovbeCeMNsWwUBnsC/8HHGq3ojjoQmFRvXfMOEruTRU7YX
Xv3qiDM/hqtBSHxVEkyWMDtPPuou+K1bVxKFnoWfLVRTJo1UwY/4MINtk04z4/eHgj2hk/JjCh2W
6gzu6x7pRLW+mAP4ee1bJ+NAEVTCz40/IEjeHfZdtHkhgptWru3kvyHXChBIqKxURtzLDmkF8LHc
LNWKIZ3vIXOQrB3jSdGkTh+rg1bamUfdSEFecQZPtpIlg8w7OgS5zsD0XB+1HkfGJqMi7r6cObe5
milHQ9DdSn+voMzN3D/6ldxWJ2kOXMO3P7L6uKvfDrmbFpnMCU5fel/8UDeXLqh95Bp4BUTOqJnM
dRvGbLRbxq+H2uXCFFHHSfsrhBol5LX89PzIOj/+8QQmbci6pM3qazTTwEuC0taWZZBgCadwdlfj
JOfxfnIXwK996e8aHAquolUbl53ZUdSVzXJAMNe8K2HNxf5/3HxsU+jydReW3UO3eDbZsDPPG89V
simXdS2gyU0RoSvQUywkiyI6OMhJ+qkQSD4DZklwdLTz8XfHArj67MGbU7s8T6yqNOzHcCQ/HrLN
c1nh9LZKUX3WSF/pTGXadV/yBOVwZC29w3M7WrReeEUyVxs4O3xhqhe/QRvNXMWHWQCV3BEJT147
9dI8k2D1VVAk84ojNfAJ9TE/IMWrWDiHx9QKbmEg/jpNKuU7F7044aTNGKzE6zzLXFtWBHS2QwG9
mCuf/CG9YO0lbLUgzIzAw4BjkfvndNxp3xoqrQ0h7Cp1JdS1K8M7PPprCaqABoAxPMJoCPUNLuY9
E6QZN39Yw7igdYbd0g/VJdLHoim34dEORATc33TfiDnRHvRRNu3gPTyCYeQohTs7sU3WAXakIhxJ
7LsWtUnE8nWTKKOZsncHo7QzSMAUHGQBGtu8oO8RbB5dhD2VMjJcWjymETOtA374DABmfpePC11I
Y2BC66Lpl/rN4Qii+49U+cmU9QDDpin3eIjJmPdoIQVCbDSu+vc/uNirEeIAP30uh4yZVDIcImz/
1DekJQmsrgMAFhw42/MzjWNynWYlHcF2S2mWMjfZTdNba86qlVhoN9Tjm1uPMBAj8Fsh0mhtr6sI
JSOjvF7ejGxVndpSFqJJE6cFIogqDPwr5zTWs9aI9sPjbhzdY0sTZyJEVmq0TUxXQBWZFw/LIJGg
vIhvWPXk03UiBIoAG88QYrKgZ6XyxKtsqnwEazC4Zv5Z1/BRHXIPwNopWcjliD3tCjEZWS7zCK3a
MdhbE+5pvmwBd79b2RVBeWfT39J/gmORT1ygr/GGZNlL1Es4eR3M1sf7bDWPTvCSLDGRX03zZ6Zr
cqjDaIXbGFIpQaYhI1M6VWFnXMCPskvcPmJDr8rd7bpWi6d2TqBVKgR5mulH2jzcFZaz17tfK28V
SNSBgTS0T8WiH0/To7bsjSWbzpnEhU2WXCyxkHY/LBikrVhCj5KoqkfKF1fxiGGhn9xwZs9nTBtl
an95HihgmbgeZJ2BIeAxe/VqKp15Vs0bG32ucdIb/43LrQ/TPZH9EN9xgQxcVSYLeWR6JjYJwpE4
H25QtnLs1eZtAf93bOkLwiOQNnsuCe59NYfRKdGPWpkcMoOdrdKoncApwZNxGI3FJfbUWqw1VEQt
dKP2az9y1VqqpV4oylu3l1CmdvMeqcjyWwq02KL4vXTyDnmD3Ti/5xYi98PwNqCgnHCTdBT2CSCQ
tMu1enW4Re3/XyDJFHi9NMVkgr6/8h/0snjSJGdWsjl2Dut4Ye+V620An3MO3i5CKp+vvRpZUF2S
TpFT23CafK6YPU5TjLSslqwnBuQ5AZ4Yst43F9JGpIj2W2SRit/3PQKgDwcgp1Vr88KEnXAYcvdY
VrTlHFEQI0ELyDGDcR+ZffQnGctTW0lLEuqvjYispw/raZOt+syAckFQraI6/4b3nfzKpCpvIY3i
1f0YHPlp5+gMlx5Jo+NLupm2yaH7pyPx0F/KuXbn8X4uBVY5StRMPIebe0xpjLk5GVDic7VEGVGi
MmF+RfaK98XgsolLqRNGf2pU671jtDr9TSE1WtlkRuQixmeDFHt6WEZrJNhIj94bvgv+nuQqPcR7
S0fuqsgv+mJJr4lFpICtfqgy4A7CVgMgkMWdSYE83MuCYzaC8npLsqbEUi5Wau1o5it9BNznCaAH
f9lkc34v+n4zmtqF8vvv+o02B/RxZNtKfONvZ4AMJc+bTMhY6qk/f/1aoZpBPecXT6fJhMsu7uw5
v8aDF5Q9VGA4v7xrSsGiCGhAv3+Eul5uYj+uDXUC9V5sBw/OJQx04YK9ONfAI6Y9tBlFpoV5rw3X
s6G1/154byIJ9iyc6nFjZzhCjQsGt8cNEA0jboHF4JVukCXTNuZ5PMlHefMrJB2ho+rWUDcqftWp
0lT3IuRAmy9SzSeZTlVMngLeeZfnd5mcjLjAmqOJMiP+iWBc/130YBLXNOBzZ1xXCiDW0JF+hsYL
RsvSXSPkvXyoThi7+Tw/fS3ucAS4WwiKCoOfD4RkUrAxAweXL8/0SaTvlio7ZcBEouJ31UR0dRe1
hIIJX2mNUw8aj4auznBwm07Kq99Wquy1Zo4Sjps6i75g4HQt0PQnUxCJ/aPgudt5sH1JQbjPxk8n
BDL4nhlBGrbRUo9qgLKqcEIbOrMJI/E2IXW3/dAWUQHVJZHcQyq74xz9G2V6u3ixaI3J1A1tA34s
ej/tpfbfZSUlqjcqq7Vbo8vRxWGdX88ldupR02tLTQcg61fJNJK0zxYpKWYBzgLzd89foNdsf2SF
gUg2OL4cBGHzp1Z2bnUsSs+9K5xVAQskezF6L3Zz07ZNr7jkaOBzrq0TMY/5wt9sHA8ktmHbfGIk
V3PpKfMgv0FXxOiFHprBcVY/5mYtEPZNG8fWG0peBRg4KCtLlMibkLX4U3ma9dxjAcBqSIREiOqW
V8AV+MdklHDDrxeRoBtk5wu5kXLq75xM0LxuR0U/SvjW8Y8UD+Ixb8I1u6ApQtzM8E0dT4rGQuFc
ozNFdLoT5JZhLWtvKr+I4jx5dFWSy7hmPjgEAD21VjgKR0+4ugN/25dxAIhk2nA60CAK/mR/Mlko
qjNncY3CLlI+wt3i9meuqahAV1w3eohai56GzCfnkSIIIlulG1bykXqS6SYv0FiYn/qgiIIhjJWB
I52z9VsSK2HxLzKgyHPcbx+Rz5AGOfqgGwUoEpuwKMY+MBWtrTHrgtQsaV4AVtI42wf4+Wku/As+
wwK5qjAjuEY2j48QZZXmFuTxpzCNnqBeCjF9CYkWCsor4Nglu+pxKfsgT0Y+fgjmjr6dm89S94hL
KGcv9DqN8sPLnR4q/GpoFKgGkASfpMaOqzcPGG78mLiSCRyGzFeqImpccL4pY+0kVQuqiGhKDpzg
V0gFJCjQoIyj22uuuH4oIDMg5WLViPd0YxXPOhedGZhIKQDNKxupAaYoc8GDjln4NS9y3JfxXeoD
+pPj29wp3unZJ/ydKa1MPBneqBpKTSkdB4kzi90a20TvnVRfPzRwjFH4fzQgJE+N0kIhKXcLxLG2
6NJhiXVJuFTwCl9/4Sw41QTtrSJbC+KPCtMgNT2bU8mobWN2i6ksz4D2Rx+/9dFbHtJRwKSSal7O
EBbk0tB7jPMttj7r+9SY6X8a8le7m5zU1mP2oanQwOHtk6klfrIov+tq3ypUaXwAQRLBwgg9cZwn
Cg2DOr8RD9iYb4d3PfcnZNPs6s8zWQrqofRjcC9U+TOREm9ToApXiwbFZGNUGVXG/TY1bKJ+p4QC
2AIJ0msKHbF78ZhTMJJvPQACDvBpsdGaNxTcShCVHW7+gOpIS1OxcgZkhLr30OTLUEZ6yPaE+2sF
ZabGYXFGSzK8be0bUEdcf71NlDJVYU61EWowJQrj9bg4Ti+WI5inclAXnnSOIYeuHXPn7Rekh/oD
HwoZfT/mt/LlUKsY8VZ+c/c9n3K8QbmJp7hDoAH8Y/5Ehn8hZk5C2FNakLJ6jkKyILaIlqrkwwWT
W4BN8F3oCzs4Q40yFBdHjlYV5sGToOomutcjYPsnBIliDxzOHWEpJAEDytqzUE3uhzzZg5PWJ4n9
1TnXlAgAQZsmaSwll3ozN2GX/W7erthTOuCFfSXBGzXH+mYbr3iuB40JU/jbUWIctH5+7bhTAt+j
6GvEwMKF643qebERtfIGM5bFKRczOcsC9OXJ1VHuAuBPJw7WOZmXcd5XpRiE5+ZU/FBFarq5rcQh
fPzznh8WJvHCfsz6XojEyQJRVg/vkFBxnJlTfVwVIodzjErngmeWKdPthkWSBOzKF6Q/Qe39Aw4o
AXGIpiTe/5bpfoaDJAqcqczjOEtYQ8rke/F19IuPMlmmh9/v00EksocqvzN86f/ZHPEbkqMBzQQi
o9UHpL8gX+XVNlPOdhCT8TW7/oYmNN5e991sfwh4QyBjuFAJN6krq/u2WIUOoP6989+Oqd+maH+0
VtWjGGmDdQpd0bzVmwv95lCvMN9d0wmS/R9PSdemUDxGngy/eDtJ9ovpe8C/CkNINixykKLDgmfV
KWgnghR5L0GbrhAESlVWdDYvlseAxtxHQ3Zg+gZaEnxR0qYXot7aoo2cWuPDHF19St8AgU85bSP+
w4WHHxATALikkfiZQoRGLPBzyxiQ4cKvOYV0cTe/P7p2XWhL7HF0H9xjjiEl+YLNWIUgR5E0gLCV
PHRBfZjzMNUsgJAKkuCxVM4z1yP+9Te4sLp907pmicTQAftpBvGsJGNDY27sIZGoVs+Heok1ORfn
XTA2fmDee5EYXgd+oOpKCD/dR4qBA9dbd9MCYVrKy2LVnNh0niS9SNY6QzuNLSSXUfy0uQ2fBqtG
V3+PlTfmFC0S6S4NpP2TN+7ZkokABH/3MO7N4Zz9GN8PedC/fAaCGrYJsObk0A0JSnOV4wkFILRf
1WxwlZ/zQZLdSTt9W0B/vK1RkZ/8MOg2qSbftJG4USyvyD6WP3qP2sFN43hQz7MNm77hPkhkjMt9
EkbH6sCrcFbcj5dNZiZ6eyUh9ZO4Wew3CpvHFt+LgA8Xafmr5BKaymBMF1KpcfHkzZ1uEZlKdrJU
V4rXR+czoCCuHbfByyXBhrgN9TFTOApPd1cQLuxeR7VOJEuiszV6MHbEqN6XgDSj6/kgpNX/zEjo
I+62ohVVFttouiWF4iRA6B0/6rC06EWOvFxGo0P0zuByaXjYdTlZ5b9M+oyXq4Kq+BKeBFppMnIc
iMJiOyaLnxsgocvmPwzpfzqYBxChVe2UfLv79sNkIDXk2NM3DNJtJjlaYs3C6E+zo3FU5FwsW+bs
cQ2d7fE3gXp5DI31t9yUJzc3CefQcSLoT5bb1FPYgUjWlBd7eSfQbuJZ6B2wUUIL5K16x3ykgLRE
uU5jA8RDiOjBOXKpUGzZqy4tXOfXA7+Dn1RFcWOJFOdipeTXq1R9GBcKKnAZUzhIOYCUx+W0dllE
1nRMKRItDfVX7YZlKx4c5/B+uiY3pgGq2U4socR6n2E2F07256wG5h5abo3Qs1kspb61uQqwOKNf
dC69lhFzoDLScoMARAl43TlS0kHdaizn3vKOhxaejWgP2NzDaqE7gXN99re3YzkBW12gnWV2dIf0
IgwmYorFE+nxfxAW8hmTErx3qbmoXePcsiy9TpDKgrksO5Cj/1a16QJXzdZ2OGb6h5R0Jt2oiE5w
RCf6jUbu7bnRxADBkXs0pg7leDpOgMqtcAZqPFrGCBiSVSU+YJv/8f/Z5W8C9Wt1iBLRZh+rzCkP
YWn8FmoVkAtDPf8m3tTq5bkB/JOz0SnKHk9ZpMZNLtXjSzEh0XBf4cbplt8836gg9+M1w6ry9VUL
3XM5LYgljL6I0gdgau0y0vrC7xCxDwmr7fhdO4EZQdskzuFLpC3DcUjRU3kLlNJmrtfn+R8rr3mO
PyWc2hjJNOj2USIdPJamvT7nexMQVXOaCDkk+2xwOBgYR6+t17t09qu0w9cwZDNfEkqGK1ywkcZc
zYrv3ZULbd1qb96JedpG7Eje9JIn8fvz8I6wgq53HUdMQwJnwjt/pMXFuplw4u4wZ2lCNs/7tXFX
2L2D9b76+VcQNDEP2SkLz8KxpN89N9afYtiFPzMug34Fxx8vIA5dcBIfampWsocAJWDlWaEYUayz
NNze1eAKZlal+WTXGRghbt4/926XuM1emi0CARukTie810yh9ReBI+9HoZwUmUk+kIZi5LdrUDHH
esYyXZJdAe2RrG7mPqKqrfC0m63C0VpfJBG9syt19fNaP16qXmwRVQ+OWRRXbGLS6neJg9Ft1eAQ
D8wHFyUGbp3AWchemBTlzC9IGM1HfFkRlwBAmznLqwqoG0S0XqmIwnEDrHFBmLZg8pu5fopgITo+
V6xGlSivjjRWyktEE6DahdqvLnYoBljAcJLXlViLJhY4C1wd7C1r8B2ZxTJw/B/NYUBUCo3DperE
t7h+VVGZfY7EyjOqO3j/LEQ5RXD+EhFjSagXXfBsKCvnaJ0ceqwg4ITzceZdv0h+slvvQxIHmZMj
c8+bGB390V1HT5QSNMWsUHYGdRbY1T+9bsgvhYeD2jtuA6rr5WHM0Qlpq3lVhabQlUgtYF4iaREt
OM5LmNBzitWgYv4AUCgYb6tIUQFO9+35XlzAPKIWAU7dgztexklOfjOhaw5NloAutjfR+HVqChw6
IrhAxeEKuw+H3PK/7VcTkarFnkqU5a43Jm8HRnRD5M0D67u2PDRB9eiYqQV/QdnmwYzDDD7GQW8E
GhUC9prZ47yUNA/hjqzwGd3h5SioEVVuRTGvQ1rYvfjjnNCg59loFirbkXcWukibu2/L0UUN4JeW
8oTuWz+eqaZlzcleNwUWVFOkXv/qjLy6fVrbgHZE+1rS2Pt4UWV0jIjs6mVCyaOCg+sKCK7yLXRY
XbbaNmEK8OlPeZom7YUxn1PY2u6TMHPgUTV1Gn+0WetfZF5y9VL9l6z7n0TCruXi9VEDQtt21iDt
12zL8Z1618VxDW0x/FCZAWbRuDbNFRptb3VMn06C39yOEMTB7ZVoXlmFli2IbrNiw4V9f97p8VVM
8MfyqeD/qRIZ3hpK+22zxBLW6jJOz8fbDJ3sBk4RkkiQRSbMY0GVs5A1tV12MpSvTzY5c2FpiGpU
PeiFZuzUekwu1OW73WLRohWoBZYY/Vuzq3rRNp9Fu8C+4DPJYuRK+TGVo4vncSwWesCe+wnxUjA4
omvcjPtk6mK4v6Ok88vLU/MqyFnvBzJckmvUZ0zsBe+1GbI0LfQFrrj7WQdQuThCKtgFpK1gkB8x
99Go/nK9D5g9iVKSYKwwXcIbIiXSyIDKawfT/AlU7TZLA4Sbnwbt0o8r0meyV9kWg8HWT+X9j+KF
rdHOcEyitKUi8sx0Al81FQc26etOdbPFLONj0/VbqYWPf/lCUFpJ4NcgEhwRZdG8ZX6Jj3iKpxlX
o3u3sYQqUXGOZtjmME1RrQSgr3VeHUuvOuty7BkyEgM/5YHr52XpHPAVnCAE++gP2L4QkTKPF9GJ
HzEKXDxudIp3LSTd1/U+QmunkBKU1Lx3eEdEUIWKNZTY0uqmKXOq92842VxK6eF+JPNHdO8ISEKY
Jmzz19iTNJ+QSewdcYBtkpv+lzz1p7zVrT9n+HNPneR6gwBpZvRkWURr+Do3jH4pegpqdJ8KEive
zxaNpiuTFc7+UA46utWyMTbjYe/V4o5lpzpYRbg7/X5jU5WDynp0XK7q3/oPbd4r0L0dVQUUADU+
QhYWmEywY1cLmFs7K0t12jlYYeFiua1KvUOPBn80UK/UBJVnl2iiDVaUEWLncMrKFZVgjtSapJ9g
5v9HM8Mke5OU9LwPw3xs78FkElc5WOYdDXr3ZBkoWTY1Z65p+p2oBvaMQeEz7YDqlOu4XlEeGG9f
ZGqa3jCvqEVLYRGjOG9Ztu0m18/1K16+GWUlXyOauoG8ZWgSHDo3ci9MTPmN641n0LAGe4LPdoZo
ni+cmjjCV70bxH7cvje5cUTTBwSjBtSGRym9sX3y8WZfddDqa0v8lqMBLsbpqgZLyd99uAfW+ZzR
Z+Ld8sofLoEqsIb/TnDCsbsofckCqISpzq5MnOCjfkiH+8UujRk09LVTN/zsRyq9ojOMzhij2LMn
HKeMbAXbA7qfMq97jUQGfKa0ByTEE5valmy39jhMJz0JRNpMCY5XHgo96YVZRFv7JQBLBhGTXCdp
z8lhCXkSASHf4MgNKEAQdBHCEjun+48kcnmbw6/OIXcnnHCbbv6lTPU8Le5Oyxokme+ITdXmpU1e
oGaoqxZ39mw3YyVhea3ZEoBXW085e9jNw9kaWcRqzOw6cADTH+36fBzI7jRXnd8WYRkVfYA6yvkJ
U32ibUCsZyZKTManlsbkaP49alupIfTQZBqwJafSAwUxmSReqDz5g7PncEvpgdtAlYKEBwVn3kQP
3cvMC5D5mZqLhqHIVh29yCCPhpwnH6AF84r5gE+M3bzlZVbXTAdPwVokBKZlxu3W454UxyzAcalE
Hu35TJObbC9LC/vbXmqDb6RmOWcFtJehxeX8po30STHH+uXzizXrJoOFzHT6y5Qud3tebRpBGjp9
PN5ILjT7/d8ISal4QXo0uhkSuQtM3GMwkIieQlJTZngC1/qXpP9WV2XDp/oGDl0R6VNgcRoffi+w
MgMCVbDXV3ZrkTqndMFWjYn53kDL7gSatUW4qbphDKLpuWfWJTBgB417vp0G9DnsSdRoNOSRMYZa
oYh0FTv1HPi7C+Uin+qQJRu6NUJ6Jxls75unRWvNtLlQH7SUnlNiyLd1XVoHDUuk/M+sKLCk5gFP
xppBLEcnys6OLN6Qe6/IVXMoaZHbXDNvDQnHhg3A4Hrg95tesomTP7U3zGxARiYtmywl8GpHoyPY
GiQegJiIM7+SXPFEXltRYrbAw2qvYjjP1+LiXBoeifUaEDpOc8dpU9LxeFB59OqiPyyT2EQG2zc5
uzdY76VU4eZCqIlwLkODIzHnAjU+Z7TVOGcX3Yvp5+0ENQ050Mvg2ZmHG6RI7MKAIZS6IgEKTaMS
/Jb8/tLf2tQ6bYkCO0xWfCJE/jyqVFqdrFbX2kZjf/tkGsBJl0cc1DeJ2iJOmtNYvEFet6yn5cfd
Sum820yUHzZrUR1Y2BeNe7g4xKb+wxRadZ97ZL8k64rw19jOcskRnXYwBhQD5ayCaTmzqP0+Z7Mh
F/MAwHscuwa51AzxaRXy0N0zwlnZpeHB7x9sWWlmbXkz1u8LLzkxyjDKR7MX4mccxrtsYyiLxg3j
D6EsX2wCtxjMFgPrbbHcweKy6EO54xXQZcPrDg6IPUt4OS/dd/dIpmHsjpfRzG4Atyngsbz08h+W
0rBSLcmiBgKOVeay6KYl/KftV478zo2p/N5g4v0u8P0iyrXUNPd1wibZRv7/eT5KJtv5OZuZCkNk
aV0MtWzy2cmwPC1KS0nUHyo/v2AvmJ2gzioDYsF8l4bXLAQsYp6mfKQbOSUk9MdhJU/Y4q7y+puV
m4P6hTkG2z91Xb17Q8JzSb8V0xONVlfUGxQgxcgAsOmro1camEPXIWR54s7JAcip4t/cSLNKFBUf
J/6+bQqkmfF4jjT0RSajMPE86he1osZFl4idkoQPGBIMr5a1SPa0NTjvoPxNo75cSjgxzStNzkrQ
UeNz4wHHtv84Cr4ETkCOxHKzgp84l/3Rcj3R8Wd3wwKM1vHK4IX5RDOZX0b8Hf/ymvxgNizjYuII
P87qgL+JwmnUCjFBhcYH/7Mj8gGlqGwB288oy6tWN3hYIt31qlLF3UMPN1OopZ75tP+nqCbGBZmZ
hGdqn6mGcAGiOzCwRwpBHj/2i0B107LiZoyDyUFQVajJiUijFeOHeS7beSzTJ0LbOOu980Cak2OW
+pwD2rMM1xynyxww3MyPPQZ35aoxgd87pgEKxZE0pj16OiwSep30yCigmwy350yluyMwwl2k6BXb
v+kNELW1YuJhll7Iv/xe4sRSeAq4XCC5XJHsjTeXo7PltVRADT10d4zT7+UQoz9CM+Po+WDlw4Sx
DrxaBssbHI1sLjMB7Ivd0FcsiuDC5LHusTBwM99QeyOzLNxafBNXlC3i6sm3c4YvNhl2xCleCpQ/
VF8QilrxCUv8o0/cm4WnT6ehSV8tuQiAlRDcn9UbbNWfKd9F+kIMPgugJ4Hv6rZ+fc1GpMV64WJ7
VR3kNzCkmaJq/qxpww6hw4omHfG5U5uDQ8lQZRFJBZXL+WrCL98PPuf8hLn757dg3NwxXkPinNH3
RMY2N/TtFzLN23FkUNQuCpJdk/oWQzaYQYHI+zB5OlQxZ4RNvzhAFVTLndKQBlU1E968S98KhWeg
wQNkBTqX9NqI+D4LHGo9hY3Wq3IKzY+aauyD+RoiB1/s/3kpUYnvlosC51bRsD0BuKLSG8H38D3p
T2M8WFH2budWgqs2RLj/DTRdCigyQnJzeb07BNVCrhgZNJ1pUW07zTmbxwAluIfdbi6NwsdqGz4s
Xw+c1B+XKnvYAmKFm0x70Db7Qr1l+KJzKUolnF5DYWSl0SmCuuBvd+umVsKHCPaG9UA3WxUFS2UM
NCZbG1AlIqEw6fqSct4ytDF/Mu511DD87GvdquPnzOJ388YbPPI5JYv5ERZMZn2AxDhV1epw4im2
J0dOXqGQbQ9g+TJthrsO8lJlaStO+/XplxVHsH6eBqD9XSMYLHs/76zZ7NJlaTo090dqszbPnphC
zhqHKdPWIZhcuNMGcuNLErFX516NbT9WymnpkFtofCf6unWTcIr8umdzS7/QV17Skwb0XBCXP5BM
UxutJgX1g1K2mGCi91C7mV8W1VnfphWi58ic10h9+dxA3cXpzO3sKC+58YbzLoCn2W29KjD66NRw
YBw+y8JTzGTy0YbDUpp0Z1nX81zRvJ7nzaRJLorSJI1uuHVLK/75YQxbpdcQ08QNC7B+Ms8Ew4mp
EGjv0rQKdp8srEHX80AyQ2cHH7Gs5tSoxJCYexNND/jSPC2WFcQJHRl7kSzm6XhtqU/QejTR7iI6
8F7c4rPdO7qrRXza+Bl1XpDDtjjJUVMNIC+LO4qeBHIZklM7UnUhl+9wRl47I5eN9TAWlQ7BfT+H
BNge/FO2IMgoGsM5jZb5TjkM2QDBYpwypP/VJHt4k2vmqGiEYkdWJUEUtKMFIT8jxx0U8o9Geo+E
UCX2ldpO6S9Bmr9ff7WWmopILp/gnvn78JuH06iXAVz5NfmNvnzSM2La2PMgXn8V1xkLpoxTx8yj
kyzXkCnol66KyEbmJS49ezv0Ewn6NMrjNAOeZFxrXtSVLYG7SdsXGf3CFxetISMQbNW65kXgXHD0
AoN+uc7oHIJaT3+nfFZBt9Q4I0waYH9IRiBqZzno0mubINpcl4fp6mlzayAyPbX/TE6qL1nB+SHw
zsNHHCVSLCO58x1vC2uO0ZgwZ2Geagsxc78OSd0bbyzlNKIseZnLyfDhCBKzyFmZWFZXBbb7Z89a
93BIiL+Y9oqvLUW4XhRP8K0Vu1tBJcaTJXZgpIgyU9U7nYhfYUwd+N5RyQOIIIXM84czFnMf6NDb
ipEUTria4uttYEH1AvZ5TnXY5b0R7zr4cvo6wIQFVK8I3qJjq4177L8nYJqA55y8L0y/jSP2h6iE
DC0IPEwGkLAYSJ8cnOK5hoCW+TiZ/aB/eGq3hYpD4jz6604+3TqN9gl26uDk4Ssv2luEt7D8TwM9
Iz0WJHSslT/u1tmMTNeRDrS7uem6kpL4JEKS4Lb4M2tqtjLKOE/5KkUB/3kNfN7uaRKWS/bNKXVQ
Vrw5Eu2UVWncV4HVVM9yb09gLn/9t2Go+T+Wv+376w9BNbNwRjsdVjQ050rvSGOAotYFwh3AaZNe
0+6KiIRKbk5gT/6uv1ceWihhWy7+bhNnrRxQ7Zy/YwXehHWySs8mmS/Q1nHbNdQ9iEOBpT+Z01yI
zzg19a05FKlNr64LmRMyBWyiArxlQSSPf4+di7PQRYj+tPgyXrveFwZaPa7yDYWwlcKcPThiv3Rj
r3Ya/4lsChRqLB7Qh+bHF86OOPcDyQcoupaj6k+eLI6/1ATdECnWhrijQUvor/htAmMJ9/oOlEHa
JT6D6/vNRDp5R1bX6ZvPSWkkVw39cMMHI8J6nrzcJ0y5/7qlGmpAGdjlNM3IIa1kfLwPBfiVVDaQ
BEi5SUpL94ZCXBmMpcN7Yuy2/4ihgDZ7lf/jYSZCyj62swslNF3kphgBszY+uRcCs/kHDgOii52C
ktbSvBWl+MuybIEKA8Z9E8x5cCwATKdBlpUu1NdqEX2xRy+ym9kgOFJBAnSr/P4FB1bgM3iViVgv
hpoDqa2yCb1OMOxhoTUnoAES5iQ72qwM+hKZ0fQW93WjqxwgpaZRU8EyLO+rDhSarCp3JhoEX18G
o9FkC8jKT5HNx/TmTQvtZ7fp9HEnbVooVvFSCx0k5BwUSbaOOzogI+4D6/NNChK3LczoBXlE3Vib
L4Wo7IbAB8eAP9rqWguBviPthBDvt4GuXxk9qfxtHcWndpy99o18iLVjoJL2WCncwYn181o3phrv
Q1FLteRKIFPgtufvEtnGPDtinrAV3hemohQ6oq/ZfPl3Sk1PJoXhXGE/3K5Co+02eLIVE4fQzmZv
ddfbU5ag3WmzoFSXQ1CcSytB4bYsWaInBEU3Q6pN8TzN5hOyCDpAgCKX8QFLOocULIgoC+H+D1Ai
d1TkOH7j4sDok5HBXKCuKF0UAh8SLLDFrCuASNS9fPmJnVh1OrIXFM8NxvuU5Sc3XtCVXTI6nrJ0
37TsYLhdHuohdUtkJyQIL5svNkq30mIKfQvqazumg1vqeAXfoLQLaVJK0+CGa47hXKzpSSvqulLL
HNENc0jFhY2nuMuNm9cghio6myLn7K0X1I4U1HPgi8Ep0qUk8xWtuEvbOzGX/BCJZ3oMvNzf4bCx
HZNcLlQnrZH777e8Sjz1JoxwPU6jg8XfYvDsPVnrR2uK+X6F8paR8iUSMlcmLdyipcWGsXfaBHCt
7DeCcFGOVgfHVMZ9LVy78/j2+vqWLdarBb5zE89q2i9p4A4Mwn8iFcX5/45tyypS1MFD6OV0iCG4
rYw7XwEcBWLBxYWxsKtCHdoYM5b6mXOk0GxvRd2M0rDIOMCahkZu4XawVo0ZoAb4jSpFf65PdEZw
1CGNrZ4TwYwZ/ivlO7JfrEhpKnuKL1WfajMCt40xjH5vYvJIadyvHSpezAkazH29N+Mc0vhUAlJN
9SEr8LaEiK7qe6qRpKU2xhcX+2W2O7kcOH5L1ufMJoiNYmtJ4CuBd7of2afgD4QN15HJ3v9OFq+4
HM9u9USIT65oiG+SrL8yDWEX08Ij+AsPwkznBOQIA5/dAjGrUqik0rJIf0WvBqNTBGsjKuPIdp/V
5enyb2Zh7eeoIkaV/lBSPLrzZfACpq3mP2qhpxStoSiDx/jQvQMjhK0owg5lY6etii/Y+IEvthZ9
966cT2NwsVpSwfheVLVJ6lUycbriPj/kb0CTssvlEOe5Lu3dQHqFa5IwI5GOQG3ee1AxkIrwtkdI
gov6dlCkxsd3iOMB2tWo1J39Bdh25LFzO9aQqnFocIKF5fjW2PY7lPK+Xnl21r93mweUYyscc+7o
0GdJtPFhcMmZOTd3iWIsGQWdaxe+G0B5D0e6iIiAznmqUi+xBibPKiTi1fOKP5DS3GVoA3nesXgi
rfEXUK6ihv2YNOYT/hl2yyogosHd/ELauAuLcpSJ1JD21FxYlOK1tdcWHhHtuAMj52NQNLfwMOxr
mf+zz8vHYVFr5eSqJDbS5DGNsVlANFa7q1mHwebGke+uUCZzHMxdpCdXHXWylwvoniD0rEpk+gcg
aKgEdNQBYYhn6cRTraBjW0qNkTh5jyPPy6LdnL3SQC3G6EAlpv+yUyQdO6CNDKKK37wJBQWPr5gf
6mOtP0y4dhMbf5o00u722MyXqv/HJ5e0qrYUcv4r8RH1d0Kg6mNUXB5XeCVw5BRnBUltEqfvvShW
xwJDyUh2332JQSAU6kZaUgTPRolk4NbpR8Zx8YPMGTnELPI1wSe8b1FJbqPGU5RonFmXVUcStqPs
800ngGxECZydjSoGROWhYsB6JrBjNZDK7iBMHvxoFgR1RZNiB3gDLLLjGBBr3DpcXKhLab3vvoj/
rJqOz9SeFzUYgCWLe2UV0ky1fFGhXae30H+JzDgblXx57KeuRTIkcCuioqpCC8/MRS8Iy0UK9uqU
kR/i4aaZSOwhpTJXTNcYDOw/EIV1tATrRY5FVSCtrqrjg+NXLoYAbFgilIESG5yfQWR2aPnOvABo
pHmdMtHrH2CplFtrjNLL/td1KFgwO0imjedn2pgAJQDHXxLel8TdN2NrZCfIJprpHDllLtW6KLam
Ypwgpmsmxjx2Gv7dIRP7gFYS1pJGU11LYHMFfTzYH1WmXho36t8l6jrO4BwiqJ4JLqvdYi3DO3Sl
eo/9S8eoXwNSbaYxc/PgGwfKRhgaboOO4bLYrteQC08MwlSMllk3fqrvOXw8oM4jY3MuwMFQ3pOX
5fkjbrZxvm63CSSL9QjiBo8lvnoZ1nuWIE1uITx/MsrIh+OAc6+CX1bnYCKfTqBOpYmV9UtSs8Zq
TlmsPhvBvjvEzjDMv4sUoMMUXP0A87mpfHMndED8d23FKZjDbgcQGZWSsKeA3cLFXC9W4ScmjdkW
LdgvzGj6JC9+8KcXNNMl+C2XX3/BR7+62cxwlLWfocRzgYr/4uVDX+CClSUaua0WR1/HPi0rKCYG
IyxQPM9qWmdWKoEyh7jP6uFpChIoVicSEZdBeDTk25WSFiJE5SCtiCLVdkKw5+CU85h/6K/u8K/P
PczW8uTwMf+FFmyhfGKP+RZgvGQW01kHwAHzEt+pncm8IZi9nmrZRWV2mOe8fjo586Umnu/rfu2H
alDG3i/MMM9qox0UDcapjUWQ2npHiUObVSsKBwLztWlsqb+JCcB9QUPtfxv7VKQimb4MeedbNnhf
WqbZeL1229/4m8+2c+stTsR1lzG+MzB3d06OYS79r26un18+DDGvVUfDEQ6+KCtnum7hdPPziItj
VR8UmmwZbjmwFty0KVBHnfLfkA7250N8rR2uBqREiwCI8cT+QJIV9QI+EQ75v5orO3mzPRJ6HsuP
7FDYmvwzUwPxEeAbWYFrI9VPbvCr6faS5PwBmKpyxO6sGCm41e6ssWyy25vO/bJ2RjXVrr3Na9YS
kXStarWsHdmiG4rSo/IoPQAKFJd5+CDiPfsz5oFJCZkIjygihywJ9nPxm/lzY9ZaR1AKd+hJszGr
GQoczS9Tvn1H5MYhb3Z5uNuL02gZq1EWjAkDp77j7EF4VnOOCHksTCIwuFstdce9TmXSPy5mHT7g
f8AOA66MJZG9rbk2JKUjwnnpw50I2nr08i++3fDq4UaLdP0HzfktX0R6Tx30+4N4GWRzsc5HgiDC
GupDAE2yrkePZ2cHNuaaaiWdOcgF7JawCrfWAK7h/ppT834bd9qpnrVOUj1TmkMS/Id2AnFKLZPB
BdSfPlWa+AHWir9YUprc/W+XntAD2J2DlD4NNE7AI4gwUGDnoVDQTELFsu+677pM1ce4AIOhJnaS
DgKob5+kaBDcF6GlBFWHjbry04MSLso/RrfGjQNlSWTpPbC2R7CWBnBlMYJfl+6gXZyt0EIzsMg2
ZhUVuSwviZyPhKzYmTNR7s9DVwcVeSptpeKmacBRgkD2gQknL/yK7PoHbUw8C+zZ7OiVbvFaiiaY
luIgBB8lBPHSqKSnmyMi77alfcv00o9Xw1BpoGp6GZuvV2tbKHNsRHRaSuVrYJ5Q66dbeiOI1uoM
f4S+pdFtzK9YYlBe5Mvf9sjiYgQSABQztViZVMbMycuT5XykG34/UmEvIjtL62gxehZeKZcyYPnn
otd6zPxNGnLVZ+W7xQvEcWcMzY6sELSSI2qOgyX4QurfvWA03vU4GqRsHCpJ1vi1pmluEPicdGfs
THL4Q6thgOPIJGZVQ5vg6jZ/ne1GVumtw4P+tl0kFmLUW8GlSQqQ+rhheQ7jha8OiCjpfGxrCxta
Jrk+kg+F0YMkwRVeZQd3605o534WNjy0L5n5lbJGLfHO9l0SLffIhvs6W89apATQ1EnKPczgZDC6
4cSD3pLm4Fn/izHPGeXFATiYc9zNynRnhWPPp91c+4/vliwc2HY94iH8tzChRyTySsbyo4rX5W6t
T/TjAfJIgY3hqryo+3T4A7xRQePaz0QD8uPGFAXmYmAu5M0oVhaloaCMJDkqPUj/e8k393v2ozUr
im3PPfcw+4BwX3SLPMckLmXVRZS5I9cZW1pa7qLdojjfT3vSB/fcKjhwYvGduXiYg7+RxQN/DrjU
v5XWUZlsbMEVB8kZADUNixsJx5EdxNt1DxmD3QPhVdtL+He2LnnlSJvCWbs6Nvv9CxUq9pxDW/1M
M9nafuzAF3DLU+RcnSbLu84j6/fCNbNIBij03JG1Bw4bzq4yPYfwAzSumF4HB8Aeb3y3yyOupiJW
qoFgq6HBRW2lf5fTtwmOna5RmZM6VgEjRgagwrnXHIXuCcRllQNYlf3pXsqHyQDmwgMLcgBcZ5Da
Sjoq8+k8N2vb7IR1LWLwkQmfM+W8Mgkj7SjdDR/7ZXU6IHx3OPGyYw5cl7igwrWiWmlqjLQwUgLR
grwSygH6N65CV4/kOz0Zijla7B4jLGno6lJKeNxZgDkSvWrj9/MA50wFm/vQdZjTmm1PCVz02Bjk
s1SvKp6e7gI2hSjSne9wuM/cAZG6G3hTMnTTcemxHkr/vmemVpPxCWYodPqtSZj6XFXJDemxFdLL
1H1Gte+H08CWwu8CPE36jsMmFKrksl3TGSofTT7ZwUZLW9bCixODwevVcHUlMO7JwluNXvAvXqF0
t6lOtTkztzcw+UxYnLyU9bzN67f+6Z+gavv8DTA7WslVM74lTYFRTUXLJhpOk5gvXcXtcK6LB3CH
Z3qbAahDN910+z5t0DnMTKmQ0NTfzqcY41Gk29XIalFX8nPE147ibT8z3FT4VsdUgzOotMq4Mol0
G8XlatzeekIGBBNlBBEhQBAXubZuZaof3/N5KHD96j9+Lb+9Kk6oWTFTUhBGnsqUSQ7LqzGMjrOm
t6Oonor5G+UIG/AG8MxtyiykqefTRIgLXuxohvWKVp3q9XabJmIluoy7Eiy/6oAXZwWnvt64CQOm
fxXQVbFTleRg63GxEW4OpEGvWwsAwAQsszcXX6MGHjW+1bDuGFPfc/dV5mcFoNkmlSS7eixz3eCD
uTZiq9VIvVzf0qTGIa3SOGNie61YBx+lT+t8h18stCzxY6WCnQD04viPEivUsQ/W56RRuYGRWtuC
NdXSTUTEin39Av7hnhFxqWJvWhshvVvvN/U1ARwEGOV8rrzKVI2WFUYMfhuYgFy98UkoyWiDtE+Q
XoQgnfXNY73P3JtGUpLNNYWym+Klrp9QsUVgpoF63QbFG7jinWnUkKothyh0RnxdVSI4fD80dL4o
IaeykH6bhcVLYCnggzC+9g91Z0EYB078a0jfqxHj0v46MUKycyPqJPK9g2tI9QZyivB40eY/zsDy
tfndbkjGcUgP7ojQWzGUtmg4fMl7rXIch9HaCGSN0Islc2ihFwK+HP4wUEuKVPH/9Fadj7ZeaeS1
UzKhl6WKcB/1bsHGcl/kS2P9TsW7YJ7BGn5lvAFBdxu9j2BgsKOUSVtCGcWsvH6PdLzKmaQArZ8V
T4nhFC/E7giutjFgnrglWPJAp8TP4D79SzLNrqAA5MRUko1AzaxoBto5FcvFg76xjGBZ5Hskn2eW
//kGk3ZekvFgE0v8784TYg6bWDHd1wV/l44xw1hYIyOOJjUpb6IilILMz15NexoFBfUhSOjHS16S
QykkZqa2vCytdmXsCTkZdZ24Fh1d4cs6i5XqsipMvh++iIDQRTmumqCTqZlLGgjI6mjEdtNMJ1jT
SpaDjUzw4CnWeSRTrztboPKuQDpGMnPUC5+8q9PIILJwiIL4zpNNSk+VqnxbeosLbQ3yy+kRdYUV
WYi4muyvSrZy+4ARwTKKlm2SakoluDbhh5Hi2XDR5PQX8AJo4eO+ngzGM3Q3kd6b/7cpDZ4/dtc0
/22djg1AkOtwahx11Cz7RfTNz0/4fxP2XvxtbG9704YgShE4SUct0cv3X60KSwZ5hMLP4D0Xr8+j
weOrf6BPitzcdAmaVgpnEFOEXmAYp+1GdG1TNTy8/93Ewb6TJ5Q3ou6t93cuTalsP8oIrVyIDFe4
S3q4A9qCHghl4UjT7XkYrJ2GTVmwEhxHdoQ8wxGTkXTh+li9pvaMqPOPVsUXJI6oGhg3S7EoRZAP
/GTxL+FuJux/SALSHy+P/V4MOew/XyhDrun03d97x/OmVhzXEK/tK1sydxhVjDClSBrH56KrfFs+
XdbJdB6O5OO3e2CT1hNWEMDrXSWSViUqjK8DQRkKQPMxJcJl1jYhBm0AEr2q4VNWfMxqitHj0qLL
neLbWu/sIBx7CRPLG/kdd44RVFYNF90uJkVk4V/AXK4cg5IeAPl8+OWyvFyPib7jRb2stue6j74a
U/qCKb5LYVFU+CWEw2lL+LIJAdbm1HakuTitAHwgBcSYam6xtrPiZw4fad4HnodlVo0/+RLZi/i7
jB3ZQA5wa4UMZiLKm3yfj20GjNMpHNZODfGOz/RotL74UNRI2c0Js/Hh8rqgHdRBTZYvwLoNISKg
V1D4LWrwIlKgI+rIlRbCMCPj/ov972SUPMBpcj72QHmWU8o/DA2aTY1yUbxjbxVVASzJl2peKWXC
EcmdiVmox2LAkjPYdFqBEgh0cFSSuY3+eIg/A0NjNdV3L/Ro8IEyjKSINyghJJ4OWaMWrpiKL0+o
lp+JdZC0C1CztucwzPR71iUC71HGAVxl21sgvzz8xW71CdfqEXzsllvfekd/eWjICVvhc3adyZA0
IQYfcb1srawU23FusOptjSa7KMFNfLECu/7nOUTmhPW3N7IKvi+noNNyf4gET45UiRtuLkud6Lpp
ZZLLPbZSFN768LaccQ3vu8cjlj3SNascsWIzJa6qKR0uIkIPiLomjgWYm5aFPxpbh2EM1STdUFgs
5tVOsM0VSVF9x7dGmjsq3gbudGQHX68dksGlzxgw6K+mZIv3P0gwMVXXPy+KIgSTx5iVI4SmIGHd
BE+D0GexLzIB+63TUALfLplDyEj+Gz6q4WSQXYQatQ0BQqaMQuJmFFwjUM1hO5V1kIwOhfoKtzbB
a74cmWs2YwxcR686P7QCbwK9O1z0C+5gQIwalr/gvgLdYNTK39bbhQvdMmQev8muHaWurPvuzOga
dcmP6jeZEqBC91yqQx/8IQjdwp+GtwL9D6gvAHOnIvc7ObzR3Hel7JjPTaCbmLL6SjX+62sRKAIl
IikfCtrnoZXxpILdf03pCgO4gogagQ6PsmZ9lbKYIqVmeEq3zKdb+rkgP505HAU26vUc25P3K3NF
7wC/CbmwNh4ZWzYonGQhpAEaEdZhleuMYCTCkMfvCMZDiOvPUVQVyjwwtFQxJdCgM81CbB7fYLBw
hd1IO5w2WuExJ8yd+bdeXqg+bQx2izolKMuBvaBsbd0VMFwvzQkqLBlrIlkujTHMVQzs3H3bInkr
NfzWZj4f6JlBKRENT+9C8jSdevUIENZRrCKWPBF5oMWSb0X9OPizW8KZ18hd6N2urXzg6qxkTHa1
aTmK9oSa2LT6C+VnSboa+k1hpGH/fTjdH3Up3TZoVp9wVVJljH27FF8dt8JlZ0z9HYH4iaG/DpeQ
e1+GiRp/p/TCAwbjrOXlnlZ0mKg1WbIsfwpTFo0TidEvSIob9OrZexqF4lTCUOpu5lz7Wz5WUKFS
l5TPSX/uHL07cM+J1/56pHS/Kg7bgxbrU2PC9p/Tb242pHPjodhy0WLYdQC95JXSjtcjpFsHLg/f
Yfg1CuxCbaPcFNGpjlCTObx9CLHlaM194DPeiDq0J+v7CMVS2igI8chvTdmL+7SS01n+e33Gum1H
hygt7h/2ZcA/peJCvNzreq7N5m5t4e9cd1bU3zm/qGXHpYWKmrO5iS6qm8l1qruvvvzuOBeqU1mO
ct41SvfUbZy3xOZMMHEs+LlARf3TeqmX5TuX77jTyIKV/ND2XR157ZFqqlwybFs8R/hEMa2sp2Dq
USv1ZfjVoOSZq4TmsMTOlma/ZntrHMJR5nCppQ7OfOCAlehHYxH3EfO1Iemp+y7chaa25IgfkO2K
M2tWevG0ce+WjGU0wIjRj/f3X5CjFUyeSlyoFaobWdvOAq/tOelvXxZUbu7kk2ceHSdBwGXpPYG1
0g5P01CWcnFT1zw/W8/urG0cACatLZseTBeNcT7wLhsPH04gTPaODOaR/NxfG+QiHGBrw7KwOxvU
E2riPZqk4YfqRwtoO3bHSLE1fs34KDuddmVFZXIG6dOJoJMyNF4EgDI16xkE6WQ8BK9A1UcGw7Z1
5BdMI5VOT472vsXJ0ECn68J/NjJGsQ6sMnslFBfO8xKB7N+Cy73fHF1EOVCknpIjqdWRFSqJ/6EP
u/oLUlUdYPrT8Kua/uwz9gbJxPXf3XMXJqOQLkjYz0FdpAckH4cGm7PwW15QpE52/jC0JhzbVmvU
uCSq86A1dMY8m9APqNaYMGa6OIExs9z2wigqRF8dW1tx8wwnKB5cpKwb09sXVvtWZhDnifSRQVVH
lzqL5oyu8wNLtZ5TL06tKk5E1Iv9xvNFCzXKMkzLHQnwL9qmog/a4ZCNU9gO3q6qqqNKXZ2YQ2ai
Zjmm0W+Sk8pA+VIbGNLbB5Qt2md55qwnW3cNKP/Vg0xgu8BHxoTSn7AjhvBJJy1rPiwhT66dE8L/
wHrtwMa5YCyOuLmJVymBAgKm7+Jr6XBGVV9PSB3A/n9MpjwNFl+zXRqqOKxMpg2rSwSpkjQWaHi+
hibS+Dt9JNZw0PKo8AFW0ni1kwYvH30QxYvTiEbCQgIgFSw+a7LJFVwpcuGzsAGYoYuat7Xo9n4+
ZyCKpaRwXl0WE6G6Ta/xCzikJMxBXdYnfWSy97EEk3qOcOoX5+gektWFzC2gAnhFJ39bEL/xJEXm
kKgqKZb0cdgrfP+uubwAphtSfZySR7piJq/8gfzDzabkzNHdvTy0mEq2B7DKvrpxFio7tTSMnaXY
yN5DJcfN4Mm1agcDFYnW7Lm4gWglXcvNvtwGfWZ5HGyQ3KZjj5XbzzldM0Xr4984kMsYWTatEbZu
5mDG3Xk1ODFUOscNjA0UoitBV37j1EbGtUMsgeqr6w85RCIPxRjB+xnZmwHAF0S+7/Q5vRy5CBGX
Hdom4tPJcEZJnSzegUoPziRuxTEb/SN+EzPMQ7C7siakInIVQphFBNXU8Aj7QDpt+ufeuUa/n5Im
O8d0xJp86a/oPeOzB63G201KHtQDqHVDm8R63qhMRRFZA3daabyhwL/iwS1SCytqRJhhX1HA9Kb0
oLWkn6XczBJYtqA5ULxsqeONqa7GI9K3WIyIA8M9PboDCIJdSil9FstmVujSnfOMrTYHAvnMk5Ox
31D3X8/bWj2uhWkn50/oNyLSStQSj8+3FP86K/kUJ2xVrtxvEsUma3pjuQl9bhXUuRkmzhDXk16U
oiSWeQPrvTA3y4e896qTyvjapOyORza1kF1XwNZs3iOGPEC7gLSxYTm9vuwWXcJ7kLly5nsCZ4mm
cyJuHnqUWvdxE/r7tzwCEdeiGqd2LlP7csHzXyBaONjd26MhCHRCHzEvEh5zpWb9Fa/pW3D3AzJG
lhd/3n7Wkdv/WVxUUZVzStuZHndbjENJMD+q45QM3n9iEwF1E6wP0NIqX/dJvhwYXfuxdIDpYmFZ
rtTz2rJIhANGoCzt4uj5fSuqLtiJ+x1BgoACmM324h5GuFt9GPMScUslNxLdNPpK28L5lriQ9UWV
P+4sz3byImM2WjT8K7kJMcl/+GKJa9eMugiaIHbwu8dMGfEn8f8A9iYvxy9ukXxDeKwpXLE/I4fa
/9v6aNNHC1mrz5de0a+dW2r5mpIR4sfZCxscfAOtOEQfpEdX9Hjs34XZINCNeW2JWBUiyEh1enb4
SoLkGTYCErRx/thh1nRz3kLIDOAgJiCx7oXdNIaWpZWDQghKbgtirpWZtR0sJzikkZx2Iu6ugg3q
y7k/MfOeCumqVbP1efkKQXBiTybmCro9/RxrzP8yzJN3c2n6Yl3hbgsu8Vyp4OXhMDcQB47VVT65
OPA9Ke6Sd2AJumO6cGNHqTye6ULlfOPfC/POipI40gJUyr3YJP7qMSF0c5sXlP9Nu+lyzJtL7EEq
oLnWvuYRUNtP11vRQKMdKbv/VjXxKVwoyKwjOrCYIVXywYu626aHdyk6ttz6py4bc5jrPG9dwUoU
sMCRXYzmQ7j5XiLri3XUMYdd9wxyO/lqXd/45AQR4peabi0kxTFMlV9pWcyrHKE4arAw5ZwWGOOY
o4JTmzgseav/JPBIavFBz4IlznTnFdJAh1sqCLEnLKHCyo60duqm9pcoQk2CUuh5vCtLJ1i2qUH2
hsjNKXcdPXovqCPw+Y/Ox7+sKGbi+FvqY9syHQvF+UPfOwHl2U7b96WHVBHAP+cp3ALkbiSfvEez
kzdwk+zM0C+zedvyUUOzheN46kxjvWzOdpWXsLESwT2wXhPRWYqHHOvTSScbZNmkU39j+KEakUfA
5rf8FFV3C7uAV3w6L8V6Ih+LGo/GsnR8ZHQBUIFSjEdXQOGGCpMKaQDZftUdClo8mwquZP4NR+S4
bKrh5yxDu9XBMOVpcN4qC4KMmLXyXNPeF5GEfwOPaRt8b/Ww1ydbz7ycjpAG/uwE6yozqdTGKprR
a1DbyPYR7sV/bM8zj2goIaOzLJKHu/inc/KQGE8ZNJUTqb7iV5zemhfzmSY+4PTit6d9eauovD2V
6CULwDSlQSYXTHHQ1P0jYaeH89pK8w86LnUIl0Vxo5KWaTXId3I56ijaX5/uD5LftP383MBANceo
g3ExTZQ/++m9d3P89X9u3uivvqE+SeXJfiY7fsR/xWyDEg3Sf32QIu6XgLtqk2SBbuuqLBfn7ur/
c1nlwXkFRYkejH3FOohd46L3pgeIE9YAhxJywYtD8fTR3SBMvrEDgHoj4+HU+xRvU+0pwY4aj0xF
HyK3TNRUfRagDw/mcyX7DLe25tKA4exLZN1V7yEHmJc6pNUKxsA4psz57z8cwyDLSUmKoO9lwui+
w45vpFtJhang3/z1h/4+ItEPsZNIDUwVNFnxaETka/zt2Xv6std8+aKRRtAEyJR2wecMhvAx39Tg
GgHGw5mKdLV3L2YTzffYoveQM0xtTHR4rH6SqJgRrSOBQPWfSQ+akCpBU8ho0Oo88XYSHJ2IRdFi
lPwxDzNL2UjAVepcmhvcrwbg5ZAHApyO01/QUEDY/TfzZ5lKK5Vp+FoYdzKEhfFW4jlFp5j7C9fF
QeZ8R5GQkqELT51kwtES0C4m5Zoy4s+268EZ5ghBDG5Y3lay9va24flEvfJd1RRIzC6zh4nS6E5x
WGsg3Dc3nOsmCTovrT11BDM5KVoA5ssn7KGaC3+HCji4DhaoWTHgYYsKB4+G9zdng9J1znzNKafs
r8BMuoYkHzRfUpyLm6WrCTsZb8gtp2iSrvQycF8XQbefX3K9edYydgXg5fXnvnv/eJY7EDzJjZjd
pEOmSYoZD8iSRjt53TAlvw7hxFg6Ga4VDP1AtHtOLYOMzEWca2fkSK9aG8uGomSX1Zcw4jZpwYLV
V3ZauwQ3H6/nyS/3DFsukuehWAn6GUVYJ9RQV/TaHjvf0YaoSmqbjM+kUTfFHkNe8xIVrN7+CN2Y
WAxHHmgpDhJgw54e0zGAx30Y03Sm1pSabmeSMuKflXcwf6hNAg7NCqqJgHoQHFeqRwfN/jrwkAo8
SjXiQDsZLUfII0p7HXwSiNrP6jUuWnggxdVWtc0kYhP/79oO1gHvgqyDpMUr9ua5HjI+6F5E70no
vY9meGmcmhFrRILywDrpR8DlY8wod0YfIevvkjRLGZOcIH5vBOGHplw78pGKc2zeavxckjyPiMDK
aqzNGRUzbAQXC0ACe+8iz5IIDtdOUeQR7cKh4AKnPwTtmBmKfFnjWIYOGHBXZLF9N6NAYJc5IV5j
YLHUuoZEoCGf2ZekHlTn3+jnRcffbs9BuDBV7HUZtMhh7u/qN5GjkSZbK+OVWaaiScPk8eBXHnep
pqtJ5LnCgYoyBF4sSo5Jb6GKHP8rTDgyy7Mix7y7ULAUQOixpEsia2t+sX4U8QumgzhcZNKPwIbr
TXYqaAbA0fIICxw401NY46z+8QeHpkRZOKNCG1GeqN4YPMMpfZ4GfWBWfS9yRJnXybY4tZeYajp0
qRpoV/DvsS4lmC84b0k/IHjwkh4/W8xhi2INHUedf8/JCkMXj7e6hj4ISEJgbs3wd0PuSGyjjG2c
R/ox9OqSfpYV4p889PInZoC5/TlG4oIE8nqDQ8lAiob3DItaVvwR1/FOPk2Vx8SqjxmOb4PUBUgj
ohBaaX9QtM3TUbk1oyjuhFvgWD2PwgAhSXGW2lHV2zsJ8NWKrkV33ARCAiGHhYQFj3/9IZ0u4TEe
Dn+GuZvq7lUM1UQTosaiGlcY6zLWPlEogkyyaojw7xldZR3COY4Blsv5lonMwQGJ/rxgMGA3UrjN
K4faSv/cE0KArQ11bna+qbTACTdfETaU7JFWogQq1FmAPsDSSsyjxMpRELqM9Rqt8B+OgciP/5FC
5ub+gNvKH1rdzyOnTzU45fq15oxnbrM9tfKJYzlhpjXMdEPEFA4Kes0ZW940nhnJbHYemWIutUea
BZVOYobi9+yxaLGvOdJjqCxFrtdFF9J/jQASyPlE/9+vYkh0EWA2tVqKQSzrFvXc+xfgNPKNq5yL
fIUNujS+hsyty2YG+SCPrAUPtlZ8Mcv7hySeX1slS7HpIlCwRmSwiVR5Q6klLHK2xfIJmlf1GUqu
q6hrmSXlVa0G2w7jp6/rLznbCQmdfT+ny83iI2frCJAH0KfJesg5YGChbTHBcB6W4+eM79EWhILn
oA87cz9EM8g9BrNHOi2MWAsT9wXYvTVE2jHuPpidguLUKSyrVzJSa5PfRhubrObvk9OyRPCxW+Un
wNxWrirrFj8x6IMhc7/5l4cyDgGTPjvRg22ZxpNg1oAIgpXhcLAiT/S5cola57Q92u3vPhuE+6w+
6xq6VUvuA8UHY/A/uRBd6iJTOSgRSjC0mvK4bIcYyRGj2mZmgmXekHBLd1KDJyHLJfMWS//TYtUn
JILYk8gspLJJMopQKIfAX3dxOxzF6E/L8MI2LO7U22YXfZpX8oyX3e+Vs98C1sv+e6OHOirO8rom
bOdX4qlqgfKxhHPh167vJohzW6iF5nQCnLME19XoMBReMfpj89aBxdRYhrIY0TpuE2WnsR6btXJz
tYet+hlNXLISS2eqXaSi21l7hrdpsP8QJHX5Wb4wZcFtqJL7D90E30Keq2JJS2jhtuwjkVN0IEur
4wou0bcntS+VYgtiLr5yT5GxseplYVS927buk5VMkTMjbD2EPBTuBibWSuAp83qVE6cb5zhjy/0A
cQIzbvDHJY+qmkmUvpCsr0wPNrz3GM+eWAqf0BP0KB8C9dBe0okIu6aXNFkYy9eYNC8b4lJDYVT3
ulAOHEXGN1nMOqXtqm7TbZE4LacMAPTFxjNV/Ansjg1EFpGL3mECZVv8Z4cXADK1VxL0I5lqGQTZ
g9REk/A4VHhum7AsKlHjq6vDsNQhjockcbZB3Hf5Oq7pji807v8N4v5NA7qFHoiLRktoU5TwqR3O
gRWhRA1cSbxkjlnDjhXY5CTsb6GkppFJPI+AEtkHdSIxQqySA30J3bXrfiIHh7uZNSz0EH66MpwX
J5mdGeqSbd0lyjm6ZAy1CMTrC1HC/u6G7L30PoZcYh7dOxAd2ipbOWrdnCamJc1lAUQcDjqzSDN1
utVM/H0Y6ZUHvBBNSa1W5HRTt2/4Uq/5CK20Kd/Ducvou90LooX8OXHlzuZU/1GatW/7H3pLCNMk
pDP1SbFrbw7xHIsKaGM3pheEYsQ0PIYU7k0m+B0zyN3CTLw74H/d9ZdykCllMs53rPibWsH4kJeC
NdoBlkWsCXhf4346yeWZg6du2yuJnt+EAiGne39aLVeR9gPLKDasXdJjBrdTBcaYmsb4d95aW+1T
+bKXHqyNps0DT59EmGwTTf7rVWWrDosb7RRzuErmRxK7MAE+qwRhTFqdMfS55bV8ri6V/3tsReJ8
I/6IPdpS8ikPNCpTjYTEN2KES4WN8nUXmzOqftewk+R+M99cNG4ZAKpdEvakdv0hKKq05USEnmXb
k0o3MXCSE8eyvcobXzAuXm4wrfWa9ORO/Ses4893EBehGWpF7jse2AP1RpYtO0W3lPFHqL8/gmA3
85cFSi1IKjIYTXYqlRqpwIT25yRag/4Hv1P8L8MNwTAy6tlf8eMqeC6kMm4Hd9O/s15Pwtp3Ziz3
DSg3mAy63Ba8HBMp7q4hgOON0sI/GIFG+qVtqDFwuE2Wj92KXSo4RsJV9//3CjVvyS0IxOcR3hhi
fipgKVgYWkPbkpHeflsUts6V29mBFlKUScgv4YhRZovkod3Gz3x2OOQhE4piP6C+HyYn+0YdN7Bh
qcLdpoE88dmcthJp8pj5b74+mDl1IBgZRl0eVDCMAR6xbxU5RcchmlcfQ5ng3gZsemXXbKCTEvTB
n1f/4tI3zl95g5aEIj54jEgNdvaRe1kRDaS8G//c9KaLtFvtedltF6jpt3BdI92kob7jgbRrKlXe
9Dqy4mHOwyz7u3PxqENXWl1G7jMpaqGhCeKBeQaAEd4DpDPSfYUh2c1aP4pAv92t4Vwo691ruc7R
p/poMlrBOSMOsOIHIHaThl576lKpqysep2E0O+wa6UN3pGxMK49mlOicHwfkKWwZ7WiCA4EKXUic
u7uQmtQQH1MFNyb3vzkYT5153JJrxpfQj4KoSgFkAOrIzXL0FbB1sQ9CYCtDBZI4IFn2LWDQsCNa
Dvld3dzHg1ZxqSEdrNtum8L/7V/WutZhIOqzZVilmA5aLnpaSTTTl59KD/Unv6OsXOfTbz9vNPKD
p3m8cu09hGsiDY0UccJ02edHcXJbX637xl3b7SzfkfFvEcDTFHDcOxBGoa08XGCbo2Ap07xpjHHe
rf4Ri+ADM74zRx5tKWxS8+PSnmIODmdzNlQH3qQvK8VhcfImJyYiiqHQCgYcGWlodkf9Vcxg4sqv
sWoy4TedQP23PHGOQomZ53N/9QkX9XA4wIAbvaH6w0FAOXA83NZrakQYIrn8BMNfqczu3/fyGo+L
eJvHsm3zDjI2S+2UQMhO/nkUSNfIm5GaaCPr+CXLhEOebtoWKAnlULKnd+O3ZTiU3rtg38mnw6r1
8CdFWtz/nbai4LgaMb6YIO47/KXP/Y6DltAyzziXFngGbLacCrHWT3BGTQLPY5MeCobK0hDOQ93S
og0uQVs25YOT5/YHQlrCnB/SNvAobIFoxe8Ok8SvhGFQGeFkesapjz473IGdwG22Zaxv9dk/T9mP
I6agC2vpfCiQRWuXoUwR5X+qTRZIMU+HOQaUhCMWvw1J3TiyvANb32VEiZoNck1oAjdXMoB6D29w
aeIpp8MDSKzK6v0/Qk1Jm/a2TOEf5QGsLER+v2Vx8AZ9yeHCFxX+TepyVfbq6d066C7khd+FPhEf
SyxekinhEcTeHY0Jm1kYDBd8IvxNLSXPZk7yjWTYGZev9IMWf5hBGHhVotlq1KxkGWaNKLRxUdOm
Zvn4M/7UbzqpdQRjkpmRk2pe3IAOZXnAunZxmZ0aVS3hoav49ADdAh+JjwcSODd4Q3i5+V0TLCz6
LE4j9uy6+3mJyEhzBiTH63LN94VHLaang0+PbapUynQPGY9Nsc8Oh91PauBANynBtMvjkUIqS9+d
hKKqStAZDi2ctUkDQ2E5ao6U2pIMwxy7/G35aqBYFaZ69eaORsv2E4RPTGP/qLwEjT/f93f60w2r
2MzBP131HFGSSN1BNhf66emU7JhsDi9Y2kt5zMX+BQMizVCFCnQ1gMtdxhFkhj8xk2gK1Np8vF1d
2YTMip5TwxmNoix78x9zd2WvD1dbttKmfgumNhGOt5Zc+WP8s7Ej4/79HBDpZoj+5a+pGD0/YrRu
/jsJFDDQmsxsoB/+2f81qKqcsF8Gmpk7f6xYv0Dqj5XUcpDudrU00wyO9yqjIn/4GMhLJ2LfOBzt
iKY1X4tb+OL6Gtob5tLWn0O3lHnpe8VtZnfmEN6JrPB8IHWoIygSlLkZzUnAQhHJ4VAD+Gwqf3Ot
/XcdEQPMAd3lua60Vk3JKtYAPHbtTw3LR72jbGQMiNpEz15v4fPazie+mzb9gKDDbUZapQqHFsQc
+9oNZaqs/jS0LGWLMFJxLNotmDvp9PnMxe0iGfrA9VFKlH82cZ2FhGsLPfSpaLZdG7uMC7ujqNQb
H4TndjdOdvgg2uLvh1ekek0bylvt/PRDPVSo6inooT+YLAjKocRdHJnTRNMH0yWLQehjYnySdJRP
eUg+ySILD1s0/71oZjaglfy6XEJyTziKdJM9PaFmPf/nwAkQERrlKr4Eh7c8KMdNSZmEpU8WykFY
j6XmQU9YO9VplQ9Vou1/4BSZaUTwWA8vwt9esulPjxVAWd2pyRAiDoGbMeEoKP5vhdfvJ2WQHiwX
gUnI2O6iGPjVlabu/icLTinZ/EMi/9jyM450Dfn1oyCUpBH1NxeMmFKPybrYV/4G6MS8QBLhZzGY
X8aBE9HMh45/FjJ6/cNSKM68EZL52pvUcQR8SWtDKftivkAHqGKUX5/sp705kHb3+aMCKNlbmk6E
x9nvF3qvaGgHpYqJXBIDzD3iSIaO5yAUgaNSvyFTpqtJ93i2JvCLzyQVM6b1JJdR1MWTvdwvLoST
OyWBtUe1wI5SQa/lLPqoUdPvDFdEihU4ig1rc5iEZz5qpyaXNzDLMYT895y/aC3+GOSTjA4OJCJO
9VEq8mUgYhSY5p5MggLQSGEMULhDgSy7EEBRGlWb7ZteH5c+sWTPJbwU0W6acKvCQr4PLTvbcMpe
8R0WMwGuo2sGN8uG1nHug7pbUBGE5xzNjj524vtC/o26Ku878mAfVEzMQ3bDOUVNmJhu7iuknlOn
DydQdII7RlDQlLlNL+oHfzQGbx+FrGV2R0aAx5BImUVl/rrm2tUg+ZfyYe+DCvsnoAtduNnTf4vA
yVMsXNBmdFqs17LZJ33b12o1OAmvXwiQeSRUbVK/D7KAxI2xw94Rk7/qfEY/IvQNXuM5vswFBUc7
Y1aFp/a/NY3rOpgqYh/0PONn3Q7EGkMkJksr6dIGyYOmT1YUD/AzawA2mjogho+/KBzkXZ/1P0Jw
vo3fAPUO6m5XWofJ7pdI6m5K9SJHVajqPUkTrZC+zJcnzwps/Xw3dxxXaWtMvtJr73WfIaaNe5Ic
u3QSof9jPR9W+Qh67wHD0w5T21vbdT+tUSi7rc2rmgruQ92Tt7HrsHNgsBl9NFBXS2tQgznEbVzr
GO9VwC67J08jBUzdhditK1HWyN6FoAJYVUGNhYk+z4+nDpBWP+PQDypeJQ05Hn0cbw7ZqIxBQ6tE
Q9b2NGnGapxyD5+qoQDaGtxJPM5cUiCEtU8f28vDr8ph1AOirGGGL2nEHI40S+/0eKTF1qVUCFhf
k+nNIInDh5qvtFM7jZg63k5lBXm+gGswbAJ187zWqBOZkvSxJccDBM52JVkpUfxqVrH0U6ObZFum
WhV6a7TkNymOsm1kBTtDTMhZNLYF36pUMGkLoXlWwPdl42y7ltTidI3TJXKfKzTwZ0Kt36joVpvb
RlMRfAoJsmPVKhJiWR+K/jO809xFu3fF+0y1ncm67C/xovd06g8Gt8v7F5Or41hqr+3+xIrSisZd
IUf3uemcmuQLn6PsmejraFeqa5cEu3F81xGXgMFrauOGq3BZ07rUCTkYoBkxMx7VLApP9bX9NHiu
1iwtWQ5y6A0XbVEZ5KhVkP9sh3VhgzA12k8scvpX33pbLzNAGZfkivAXklAQM9rl5a8pLjPhTeXW
UzUy1XTmVnv3QKdHC7gx6yvLT2Mb80vYQwSddbEaAxGC2u1I0ix/zm4IplKYd/4QxrdOkfJuAt22
QbGxCyKgbjBzg4Pj2I0RV6XWUy4qQrYM+DWtF7BkG1XsrxXBc6FJjYM33c/NPVNwXUMiIMrv3+E5
IMnFU9bXoBvD320PE+IfvXyG6LwQ+P4KMHs4+Pfzch0g38TZyWrkMnZF7rSfqEZIKsnEkrMsh1p6
5nsa/InUHQczEQOBbGlrkaVubVsln6gumt+g5QjPe7TzTb2mmX/tjzj8oIEciK2U+QweUhcuKRTP
Fyu8QDfhmE54tA1nxfRaRskXrclSQitEwAP3wawjtMQyjPZvsV9Ct09q5JbzyDaVCDMNFUzp3k1n
Dqaz6gLJtBt3W7zBsXMR6NM9aTLV146TbPIRETzHEB2hadGq2SprlGCSIgMTWbW1F+h1+7kLY9Gn
kEj99FJC5XKiFqGv74C2MILF7O29z6GHGcArlrPF59l0mF37e6qovuA8mLOKsDpXaM7jiCrgmMfE
eihT/sCvUKFQQ1yw/uiwFrO83Aa0+q6mCDvrqVQ4cpPKUzzLHVLMEnuCsAdHlg7d8t5A3AA+/qsv
HNERkv5b3QRrEXPUBdnod1k23qSugVMnd/EVnOGJLZAp3a+rmt/rIZLOiBKkvmfm37aMo5zFZx0z
W5sYE0L9eKK99SVACSa5/FrCb+NKYCHvyMJV2khyfWZ7zWQRNu18xekhQzWzHoD2GSEjkCpJFfT1
cez/YYFpwMcojyCL9CHt6ulHNjpONRHCPP+Xha8Pnuus3TALsyUUJJRuL5910JLoWSjIgP/URePC
AHECHlpd0VASMA/phLzWUZpvA8xEsLW4WjGTk/GDfh90zp3YVrito7qqrapzU8wKQufTR64cAQey
QqDx9nUBPob+Pqc/Q/Zn+9Xlc2V/cyKUSer0PKaOIfB7zhKpCRbk7lDPmReTBH9QVJVLMfcFmqDa
vGRrgtsuFRrPQUv3/lFzNy0Po389GPgFhtbNH5l14oSaa/DKuaBWn81x8woz4CM2DsABXtQxRQXV
N4yvaZudDbxspr2BKIUdNaL4DdM9cAnVJ7LUtQalwI4V1G98Q3wORCv0iBqiNjqVynvykNEBkmxG
cNQtIOWo2K/I9ghQB7dQmKCoKDj3EDx/dhSKGOpho1Bij3eXil3OHrrKWmIe2/PNrolAgU52sBoS
LW+7zJmC0buQ4P3810XL2hAIZBbQIAMB4LfGH4JpNR/ix3a/Me4/LrRuZMieOxO6yf1fRYHqh03n
zcXtfn4KrwL6rUYCfusR/JRhJk0FRx0YCAvvw2+mqWoHyj8k282roeAOZATBZ5O9W/kTKxa59XKR
WLsiU72h1MahEMLbunj9Paf4V95ea9eDyLQedn3k4IByskOpJVGrecrThynOL3lEhwPiiVPUo2Rt
pk2O7skprJeHjTwlBgFuGWEE23Ty/kjuxWjG2rdEWC4LjoAGWB0+UBPcLA1XKvid36qB9kEymji2
gsQX/WIcDPIfGmoWTu8lW13mDwTPfuOy64lm57II3V3a4uUZ7dITAnJaVawNpntmeK0EYSvlDbDc
Bvy2M+MZ/V5+zqgc1FV2Qax3wOzGCwCz8NWiIJSPfSnrbmG+8nNfMW9D4JA0jlZdp/KWmMOwNP8l
Zh4ibLk2SIhSmKj/wTUaQUc51SyPNWB2faQ0bcogh+vTLSmQxvupoy4C7Jt8uJ8ZQYwkJuL8zAzE
z8W9zgiDYgvnYtiO+SPqdJQkidhwFVqgQjUovg/UX0IKM2WnF9rB9c74GNnErHNfjhq7rjPkKGjH
koiKMJENcIS7fuua2NQvI8qflEH61+fopfWCRAdLiQMNPLSkLqwUqx2DveO2g0JigTlG5VOV4T0s
H3uHYQJzuaLQR1y/qcVpVwvyvTic0disOOJ5f57gzUtQtepssTkzLOcN1erS90HnAHXMHomPBJFT
MzSXMYQM4mrFkzmyqeipvCg0gJbzLu7NYt4LUB1mpQ3dns4BA41vR/A6ahopxm4sRuio0SZcrwJd
2QGPmRvhbwNMZHh4QDUWD/Y2hW/WrDF3oZ5/dhAYNKiTKce9Cvazbr2ffkPPJqYIF0lIlpdErev8
3WtZSg3b4xc3Mb6UlvL3aNF4JpLjoeUfbY+0KstZ7fke03YASO3I/66fq2SScPzhXPftJDvbXYT3
+Y37RsL9WvOwoEBG+33QRcw3Jn+DN9gj7myF42XXSwaKqOiwgtwhQWJgRCwHrXAB/z8nmRbnRzC0
UZWfuE2ElKHYQa3vfmCOQ+HB4GLyY5Cngd0ZXSIfBE08XSt38BJUSqWLhIiQrvrdd3PTVoDSF7Y0
R5liILYXWJfCv5r4pg/QTtyNvqc/xojGNJdJlHgrF8bJyJBpp6frfkopSBPYYGShtdCEFz1W9RFZ
xjXh6+AxjpzsyZsklyYaz0NsAU+k1jNXcOHI7g3THpuZ61yQeQGWZ1A7pgKeEch8yzzQfmXvIJGb
KMNAfADi/lwWCD/3adnnLUO71xh9aNCgkC6Xxan2FTYNWmqkTCZUvYwOQSW4zgokA29lj2m3ZYic
AuX514XzrUfFBskw3QVXi/vWASWnCRSUBrCXXl723sEH80xB56Fz9agVW1ThnQUeMif555o3+8MI
PLqiSerbSaseTbv1XhLjDU3r7qJqHGZYuy2Ft3V0ZtaOXqXrt2MPiyrKNUFhytIa6EQgncgYLYTJ
VJbZP3wQqhj0f4oBqaessriBE9+tTibxU8A+WAIUKEZX0MSEaV4twV7p1TjKv5Ja0rvqy4ZKJtcL
sfLCErgmkmcM/PYGH/aazYELbuTfQXyiVJm+BTnISL84RaoW5PWTm8wkGeQySOloyjpbBcLwotTG
koscu/nmsZFmPL4AAxJI+NEpAYktowLxiEZsCHnDo0zFrJvQJavEO8kFZjXtS+cq/QzpatL4/iwT
eqGCFtTR3Dtlipmg2AwMw/jWyOQhzz8/H6SW1R8icfbeYhcfq6h29TYhEHMeYq0fflL9owonLozx
BXbyZIokkYuQUfRcV68DZkURPRVsEQCjgKXMdtVKsPHoE8rx5hqAHVuwvjEbN3D/yJ0yagYnMLen
PlNW71h5pbDjJFrNPAWfbTGGxHdeYp30cIMDbowwaAWUCGODnoWmlh4D7DSaigxxLpGAtt+vSy0W
H1tdBMWTmfQ5OUcofECGdGjrMFmUYTFS7fz4fcGDAng66kK3CehrzeXyJAs3glM4BOFpnMVi7NUj
twfJCtPAC5eUlXdo6dKupQDYinBzj8f27LCCklAjSaEySaXtEGpR+WX0gpsX926bPfdmlfNSDkBJ
Q5Sy00B3Yd4I6B942xiy44zzm1HHmcUSHYrapFNJ/vtZfSEAz5A/pP/xeRgYw9YHoiXalQMS5nr6
+fh7ujBwz/saM8UhWlrThSyMVfwNNx0qT0eO7klvzojlNCwnBKf193363LuS9yBzTbCfodEOjJn3
a0zjtJ8705ZHNbb25WHKEQ6bghO3kNTlGmVk1Ud7+ZwGrd5YDsSTvv5n/MatLCSuNLCBHOB5zXms
bPTJT6UrSnv8iwtd75DkzGVQHl+73cdHamvirb5jPsloMu0QuQym+zcsD6pLuwRa0DcvSu/dKAZo
sOvHmSzd090AADGzLwlnYJ5MEDeFzRax65YPd6PXU3QjFnExxrqJpZTOQcqzPHVqh3i5ADos9KL6
Mjp77JbYFN2iTiMPk0+irtFoTkgb8UkOdkrpiWptO/v4zQ8ESFSZEE3DIWP5KeBNlnfgs1E2KdN7
PqUmLqGrzb4uaE9ieIEWi7Q2BwpJrGbvvzhGpXaiRx0XNw32Bk7+0gLDTd9ABJ2Wy4NM/zXPh4Mb
OnNspuE42L0Br28omocJvwlgLDoYqCX16BkKsISwNPR2y98lbD/TThn+ICAJLFYaAZQLe6Af/Ukz
1QiIJNKV58V0yWszAmZepofYh6T8UXNagIHhiKP6Noat3U8L4kEBoxgfBTvElH8j0707YOab14uL
YcjZoGx+6LVaqeru646BHH651p5yaA0sz5QaRNAn+sYlwcvbNQm0c5Kw5uIuekVfjjh8KEoPUg2b
5vDe5uejubM+aQAiRO6hpd6H3q9UTxGmUIZsPDW4/cPAKa9EqStlsOC72VhP+BmjXItSVJ0tNWOE
ebA4A9tZJlYWFFBQkkCNL9WLCjyqVATKi5Be50onbt6CDmxsJ7r6w+aJwwD3fd7rFGmgKT2WhgD0
GuVsWalIOKhBYJOwE3NdeQWZs4khVLEWc/9LMSVGwWlyNf41k0jt6Ogqq2bVhMh+76Zl2NAVroqx
gnsWSVMneEk4HrDTQDFUVHbfa3s4FIoFxAo4QG1lBAvsJV1RGxL3XaJLaJFuJ0b+g1LKrIubnsez
AM0q17XH3v8DLXvN234+fEsBlaaWornmpqCN1qFciTeI1/fviSdK024zJ1qVWDItPT/0/nvColm7
MWY54NrR5zTYn/2Dkt/Y4guDYpbg9s8sW/2co8n5gt52Ay9+l8JZg17G18RPWRbkO/HVLufRyL4q
xLRmeia7Re8CT8puWTjuQ2UYkEjh5ICANsNNAik927UlX6aPNP3ZxXhJZqzB6BwhmIdFjAUQ/gbR
+QJBDWbVzNwe+UepptnGrjbhpP/zjo8fjf1u+vTlImqEscayHrqV0nKabD1sTBeGm3FrZ+GVQCnZ
U+rnOF0OFtdjkdwl0sKRn8txyqpQpkIwENVhGTalsggAbopph7QYnouIbWtNNhV9alhq54AfhseJ
RbFTkP3th6KZiretFS46Oj8qjPvhNBPRNP/9opIzBKUGE2slWbin5DZF38Y2M/n0zRclutcDsUFS
GuxEdKihvVNv9yXh9fladt6Hhei5ZaStlRXQHjjGHca0KQwHTJcVqgUWvBaE8K8ZgOgAbMAHpJbC
eBg1dTekE1DRXeu4FHQ5Ri2XOGTCA9ywiE4iXLg/RKT2292ESa0hx68hkgJS6rJIK2YSLb1Z+vgW
2XV8ZR3dBjMsbX4oQ40XxNquOP3bI09sbGMOgKvbouHRueWhhQgTtSXGZG9L+fWmUTaM3IkRSn0J
fb2yprdoaqrK0juHd9r2Mt4zMrE+NSW7SIsUTyyMZmYyNDhsnBOnubKtEmOALq7x1OWBjFsw5eoi
UFx17lqVxM7hPa19ZaANHmPBwnlLyjhhqQl6gH+LORTVI9c1AndET2+v+dAZVJFfRDIuLIWThKQN
XndpBAMoQi7Iftjv2ct/e7dqTXj0lhq6ZOfSwMXQ6XW/U/xj8R5ps9D2aCohsduhKpSyvf2zqH96
04dZcG+z9bNbYeiysM9/BcYgiWBRNM6AEICJfsFh4W7qfcqzSmwA3l3qmJ2ibZCpQ8KO6zSFTgWX
ILeZ0dfHAJRaA2wD5U684tGVP1T78awvDV384LyFvvmzMr14JxpAAMAu5kdR6pVZNLIAaVcNFUPA
bTDXhG2w+aHrFZ2HfSNQe0RNoaoryg+29cUvnhN6Q34/KBK6C+VrNRiMsTlycnjBf4kKfuTTaucb
4N+YDubzw5MToHVnrr0g5XY/n9P6OwKzicgZfarQzvqXxe8exqwbQoJ1JQQAOEyYGBHHFXNN8ZWa
THj2eL5agHAEN+BQFZnV9uBDtUgMB3t+kRhA32eaBNO0YN01dfxlKL6FgrnR/4yOGyshYhFDWD12
kvjlCmsVfAhmJx/hA26wFL5liOUg7g6Df7Ar4bxXZb7uBZYFpSmxJYdlxI+wRBakv64gkv+4BFC4
7OImg4pB0jfKDTt7UNK1Dqno/hl/Rdj8ZhvhT7hHZMqRmPfzDnhGPBWR1sh1aFO7ku9IFMQQCMV3
CoxXBVbEBZbQsfyR5HgHjdr1xk6px7EuVwLTiowdCv+qCmbOBNsHhnMvFanFGN1VMM9sU7znkr5g
chYZ9x0N3KI38uyJagolaEws9bDl4QkPT8lDDL2uHR6LUxTF+fFCkYptdZo2TSQ5SucF5oPbxO1T
L6EAtEUsG+Dyaqf8ZJVseta/jPP2noKBXYuUTQ6FxHHUPRjSKprRQWJjXKo4esYQ+4arDzJ+zLwt
OxgKYcKQOAl3o8kQd1eixwK/sMFOA/Uh1lyXUNnuLRCUjNydmsBlvaDFjOgx3ayDbqn9Qos+2o9O
yrz/dF2PDH3XnAsANJFJB7Nyx83HIHkjqwVgzRSitcakhkGMEMdBsFtgJrtZS7+u0E+20BdSbnPZ
B9I5qhrN6XEYlSb/IGvGqHsT2CNbiFa2QZTCaMQii6DK1uhXpRChiajeGmfyN1NiZCMCP89EioW4
3na8X5ucOG0puedVm5UqWffig9a66RSwOu7Ru7vKdNh7LKDbhcLKz8j5Ssz4/tdqOEoTfVCKr0ce
M9ENsjrHft3f+5XgS6YXmHTWSRlq3KpgGEToQio+7fI7wTOfhnCo3HPS7jMDf2FwUf/IKKKmDhbC
j2FqeDM+jU/++AIWmcC09obohQgIXCFpiLS0PeobBhiY5ldKnng89dQRjGp1z5jeps4duLur8eL2
FJ0w5XuoCRtMkq0GfM1V37HwKo8vVCGA6/offoqKYSxfxVvu1OBvELvp04w3Ex/gpqjmh4OG78IS
vdhj1UlLocO6hOhJphD+OFgXFsgeOqow3HDSDWjw0Q/PKBgmOEwEaKN4Cj5q7eUDP3fBJw03G4Ko
k5Etr6Fe9fTuRrIdTDn+hC2ejaWsZyozCmAFOIYG128xE6iBLF2EmN0tTnlJUx48nhiFoynhGVEh
HB3Urpmc0ERU98U3vyTtm2KApHbGUiWISySGsLKRqMT5WwGBx8/VM/xkSK8RMS1sTwC3F8ct9yda
1P9nEf07A2rfrKc/W8W80mpG+INjDaXZ4NW5YZN0wfua+Moml2OVucZmaBIbAW8sI5APyioem8By
2e7ZRp70Bo5OxdB8P1m0yCvobhNRyGMyDir9mTg7Zq4H5Tvk0PMLTMi9RPb84OQHu83NEyw7Nr0F
nA72DHPRvVbuzoqL0SwBtOsPD+kXMZelcYKw1RokKbK8pPZsOQ106UawK0gVxwbk3NJKx45ZX9hJ
z0id7vGxsjs5V1nadi9LOj9QS3khyV/ln9tAGE1IJNj11cJo1F2PieginoJUmIYEOjQuNPq4+2mU
rlBNvnilFDO80eZ2Utv2D5eMKL/6Y0rQXbuTGxIVlDH6GV/mshw8fWsNGo389H9njE1LP4FHgxAh
0EG3yJfP+x0E62Oz8AaWDvoevQVmMmilARLquWiTIiQPUIBdLjVzq3RYRQJ2q9Zim1fgpjhzHVeY
JAMXfcbOVEwv+faoEq8uut/x90FjpFaVUukk6lslY1VS2cLXzgPRFOMKj0RUL5Bx9CY7KVAivU00
KbiMxyZquKMjk7mWhQ8oak91b8/iF1ugPKY1FrSfAWgpO6xVc27fGMvPHL8qUlyHoKhtt4clVKHA
jT4MenFsNGMcP3IcfeNUsXEH2NE+2VVHG0GRk0SQSk1DDqiOoUeMH8N0Pzjmg0Vl29EH88WCjhrO
EDu8r8Ewx5M8bT47zEfE74oH2K1gZkuhfZoPBIOUffgRaZrb4GXGMsiiPp8C1Sr6Rx7IF7knrou3
QxT+pqh2NgUnYWDNkJRrfunPLrq/7nVp+ySoYDppxUflsmv7xb41RKV7xY6vYIKLgWASunTOFiVV
hN+pCBKZE0CEl/VFCtsl3XtvcXg4UAatW90gRQWQUzPW55NXoo8bu4YNaU4wZE+GsJPtNOnkLh+d
GLnpv5tKBvqSF27sC2pQDBO2V/f4TpDPxdSSvCluDIowObgDoiMH8PE2nLnXwMF2tx0JkRN9ju7f
V96M/WhQG4RrEIyWeWJx1yLZuf5XAZjZ8+NhFozu37D0SPIWHsjqerI/TcHOkupdSUt/GCh4bMHd
5Dqe0jU6XjQvZROn0NgJNZ01j1tFQiwias7stKurf3eQDvZzOmZcEZPf2VxcEmBJFOMDp+mimbji
q4qMG9DpTS7Xdi0qvM+vqltqHuCP9ZicYDTQp6Vur/t/FYF2pTWy62k6nbLnJpvXBqryO8DWKmDo
Y3NDYw7b0RSUGQ7avYHcQfm5sz0VrTRVtiSblstjC55TnSEbX84y6iyPd6y7LU2btRiVtBXT8ZYY
mr1BAc4V1PbaTWAXqFoUkbkdMiVoUO8JqwFGFPfCEyX/j0Clhc0iFFPsavkrhngYXONfQd2iry5d
bfmS+zrtnRuCDc+VNV4SCXK1YFf2DoQPTL3A+XlsEz7hnJDkra6lwJMrklXG6lgs/AOvjkQ655pu
HxElgaqOJL6mj/dMN/nIb64oBmz5MBSvuPBkrDrWIsZaA40cgqMz90c3lDSk5p4cCU4zMbDJYVc7
E1xqSSo6RVYH09qS76fwo+NrsA3b3UTTBbyJ/Q8YzMiarRj+rauiQo//MSiZxycl9+6F9guIz9YD
PPjm9gUZ1Kx0SrZ0bTMq+XiwgyFzlatIaK/YxXLXP2i+E6xUj9Bn1lCliPJWNt+ORwD/bjgPIr6s
N66QZbVmDAhXZsX8ZpazWuCO7EgPLMpt0hkcxvdclf5GYEH3nRg/ClwBRumUPfnxPKTdy+mHdgBj
K90aakv2xAxGmC5n59Bxaps0AQGFb4BETU5WM03iXSOnHukvZYN/BRTHzC8uMbFsBGZJ960GRTSJ
fw3XxT9KR2Gs3yfzYQTQJhclKd4hhfQvwYq64H4m9ZoGkveSrXEVBYGb4RjtEoL9Iuwf3M8JMUT5
aXtr5oIfX36KQmrceU7L1q37K1369wsDluOMMXX8O2MDOSxptBRP7gstkhX0UndBKO7G0GWLb/cY
b/15lN8bgm0EsvgGkG9t9vutw9BY0lz5TIdIG8O8y2mbi5t1O6XHSrw91oB6Lepfv8Lrc+7pqSh0
2v0TQ8+bD2NAxM26gUPKIHQGBVLNPtDrBXgtRMKKEDBD+6ZO3ZtUpOC9blpV9Qqvbb8tV6ybhUDW
y7q1ouWkqR46XwWIPOwx7/z/N5GjFhKYPVBMTSElYwwuB65tEm+4k1vW6hpSstdo7/PcWceM7dCm
DP79PEACOkWnu9U8IDeVfajZi9Pv0Wc8omhXQv08akZSTb6g+yTN3jSVfN7bKaLbj6gMH+rzEBEL
piPjCcgQZb4kkZ2jzZ/O93LLoGl+SEyZMiPwCs4rMkdKXnEjyya3etgSUOIyLRBagQJevyuwtq+O
wm2HvFKlraCDNkiakmChN7XEkmXpPU4dRbtvtJ4DksFSBPkmK93JjAohiNTUkDrRw7sF3KQLdVUT
MNVTy8zHEFCqqqgJNS2SW9A4aIY5VGGjIzhX7EcwuxaUCTwjWpoc4KXME6AukdVBiH/wd/9SGv6x
C8Nqh3PnOtAKoaAY9Sz/BC/yaRP9INJUCANtENe3NNhF5cbtyNd6PR16la5dCDiEH2o3l9JMAugX
RhhOLppmANUhnDryvX5/RPNGrTBu20uuDFLgdERQSsj3L8zC4KHNDNyh5a3da8OJDf/Q4kf2iPdt
INf31BK+SAxUDdnmX7rnwQlIH/UDQMF7M/dcSlrRG8Kf5IhmP/q6ruxOy/XTrsOa4esZtghKDGq7
2O1vchNPSMbA5I8sgSYjuBxNZFgpRYIY0+axa5xtDE8ZzEr8syXDQBoWp2esmI/GjQFib61+TTu1
Ud8PtvECm2tQdzqvlpbjd1O1VZAMQDrbguoeRxTpevtOlrrNtJNxCSA3sYgkMYOjywpQ5KYq/Lha
h04/pdNNXf+uDyh/zkQVQYr/yTyAzvYVG/Ve8N6NKYjZjiY7EmmAFm+FE+KLeGHkeY0jDa4q2EgX
VoSoi8j6zO4CEwfioPR4tK7DuKq0A7/09n+7sZWWb72FbhatbCrhddVCsBHKFwqig7NyB965Fnyf
FuxgmElV7k3y5qOh2K+RMuHlUXXM3xqqY89hOMBjZt432zKmKs7dOZJdwKLrZjWf9KFzpz1bf/Oz
YRU0MayM4pbvrB8bGoGJWcMDKYtQx4SlmmQZF2tc4YDSU12lbKmwqNKYH2vc3eiL211cnnYp6zQp
k5W3G6dhASih/ELqYgiOnmAt3dlNnTI9XNLSjdFqjqz7juKtfwuX29fdZExJWsKQ35JKPDNVLKHk
ELGunGGnX/PdRUjlRaS7T7oYaOI+MGq2eztHNXRS7ySz+zbkkLRFhFvPzvXwlIi7968Ytw5fje5Q
eUDQ50Ifg7gtfCjZ9V+idkmrw0orHE9aqSVe7B7MVU0oiGc3ofatx8JgCCTElZ+C0qv2ijoBQUF2
/iw+75JJx2TOl7iix7Z6EvRj7J5HjACWFK+lWBka/NZXGWJX24rBuVrtakgZ9l4Uxl15hJv0Rtrv
Yf57MfCpZq/bF7bHbwMDudAQcz1ZeSlJGYK98ATWxqJtOJuco/uKEtgmlvfl2NbrVxBcmdXJGuot
cDOJcNchGIenCFlQbrUVC8PzGnxdoyuoJNUQMjYmLSTcTm+bn7Qtn8SfAvWwXu8Gz+Y8JQHVxUA7
TVb9MKv7b3BtK35SL6TOUwK/HTv3QWIBLfUxnvO6p3EenOuaHjUCQsl7AxtZV/S/fZLGmd9ebtYD
6ccG1bDBrCfA2MFxfjks9xdjCpvFg3Iu4OMOGBNq4kUcKj0kXexoTxkGMjEFxi+hVqQjsECgucan
MFj8Gzg9j3/GomMyYokEDfxvPJjdK2Cki5op5ivSLG7rEkB2RkKMvqeQ9jMAguXqR85O1l5Bgyx6
X2HF9u0HKBHgo0L22xjqz9wUv1thQzPRV7neI/1nDLpTIe3l4KChJcrlFKa3nYedE0D5tZ1IRZi7
kR/TVHP9gwM42um7ispj2/77PTB6SbWy914VfvxV+iYa7cjLAKTy3jPk6NwD8W/WC6iweVTNWS0Q
f2cEHGi03MP/fWWnMEm4IytWw0cE8nLECyORz+eJehxRhi4izo5jQ4as+Hp9aMR+3t21PpCHyLUI
CP/Imz/saqnq/7XLHv6g8BuXILOKCbTcqrwRUojWacx3oOpJnMxsiyeDkhTXU/HHpfVYWr7YJepG
zHc4teqRatG20bdehxwuqAOJHv4fT6XMc7HADfPMT24ymc6a5QK0WPne4A7t6utOjibaQroc5TNO
bhPvLlSrY2DO3wDOXQuflTWbJzINlfbw/UQ2LiAo13SNZsbo13zRybNQ3v7drzyweUi3jN5gMOe/
oSx1ho9qIMvSWor5aCwS5XQb/jWNdxo837+8BvnK9FsXORlkMZLvpX0Oq299cIzZqeape639cJIs
mKj7vp/xvgEIt8hBhwxKA4La4CiiFxcnzBTxeTcIZMpfD7XScKmkUttQpZldIifllbrYf3h58ful
iYnZIX6CvUzBQiL/kNiTr4P5rVJcnGf7nC/i4g+qIjYVOJi/E+zcIpkNbXZ+hrB4om+4QIgVToXS
rA5j5r/kCZ2v1HeA9bhh82CYGmGL6O+evSdO5b1rXbPfKnToZeOTUNCOUq1XyOmPc6ok0nP/asIW
Hg748TI/ZfzOV3ICzY52Y3n6hI1yATCNAiywaZOyDJAzKzspOb2rRm3lAhzm5mbp8qI3pYui1t3d
Blt5RH0bZBAys+1vyF+L+YZ1VVskPoQ9wDKEJYpoQ1atDeBZGoeYi4dzUB+u3Aw/Tjn1uhRvY1l5
UeZqdqxIWn07Ok5GFW6B5OBPD0KEv9YDk+A/z8ZQEY2+LQ6JLpCdCsbCMmtlCRVOyD5d0B5voIpt
y2k9+Ni1aM2NcdD8/lLnxdQigFu03d0W+8jjnJOfPGVJFEyVRAJVg6g/P0vqoFVOoLjSh/a2KrMF
0sLGcjn4Rii5YTOxSfRzMVVX4bgCOER6NVoym6bumKNbRMMyCK+D0i/++xpErl3qYBKmu97JW4wZ
STPQVKBdVfXEvax+yUJLvsy1tFJpFxOodqeAsMCZFnH2fRNKNGn/0NpGRK1wF5HKaiYKEk4tSZ7l
tPXmWyoEpecpHMRpiZaEMKzHmacOtZ5oWybShSGPnp0FTHueUjY0g0EtgvTVo+xZCMPygfbhCejs
GXMjGtitpJo1U89fhiMGFf5gtT/vqjHieG3qflrIbi2fSJJZmLCa9s8C07qVTlTSRe4NLEyOu2fn
UiSZ9MYFkp2RrJCUKA7wM7gYPNyAXvQaAoEhX5uCwWQkPAtCZTJPMIxb4SkANvljUbhDnnDJb/Aq
2F0zEFxuQZEaByBCFYrA3iw0py/ShfBhfXo3x03am/aRKhrYM6iEkcxIl5dUhFzQvBVYFaCh5BrV
PKkQqlAlV3R27Kb8rqfiEmJaqkpYshjzpg7muTufVogx7v35gm+zKCwKA82ru1IVhAdaLSfdMD3X
K5dtlRiLLFTR5kAtkNKIbeeVvjox4W0N/rirb4C3CI4DRGwmAUnR2fD7mYHTmymA23OKGy4BOlpT
4X5KNWRcNe3m87+Q3zprzL29O5I7BHCZAPxiyUsC+57FDAaNX8IOUPoaSv95/3x+tZI2CXMOMeAl
mQ3TrzFO6z3mwbrXCzr43UdxzD0OnvfdmJESfUD7Mls8/Q20Yx8mZizScgn+TdBG+PQU6h8cpGWe
ETmWuXhdTzKzI0dstz24xgtOnmt//wY8ud1F6su+w3iPj+YzYgTxTzf01olVebbHFxa56Sp8LFcS
HZMbu7sU8KVFATKpdOCFHTGAyBvl29zqXLaF3lyyI2dm1q5kXgciLiNuwuIjMcKBzed/ehhEYqUx
Uj5z6vWo8xEM9plc3hSB8EikVc4RnX4gbUeRmA9wbdzGpb+3EbSLnKJ4emLaHox+RkqiLOQHmJfx
kahdRsuOs1lRiPVYHVWc/s+RSAYr9hSqxxVOgvxtmlD+yLK5k/cy6duK9zlr4CSqk8D7/UE5Oh+u
J2i7Pxhg5pW5cKj0xad9O1lC7B8Dr2rygWRXzZeD6HHmG+NmV+1DFqMKjlsVnRwLr3WezY+jjWhI
FICTCXd/aRKE/KVawqKqrrZfWASbHfX1rfCABZyi/PNmWxDO+NsgFB+FsKOcxcSrDTzIZFtBf434
iLUkF1BKbfwaS970JLbNqzkeF8KL2MmSMCZwzj4cZGpA3mNdbqiqL6/c+vOh8gcRkSEc3auoCRAc
lbr9hIgHauCC1RAHdF7klxNFfuODSZ0kKe1fSjNxdoNbry09JLcieJsdKK/BC4lrkg7MPTpdOUYP
4ADxutKKGYV1AIXArACsbYpiQyKYponLiMod/lQyPK/+RWnUL3uOwDcXuh2KZLbaKLy/U446s1Ba
TXCB5NkkD2AZKxmJkhatGWGdvkwEqAUSW83nyGBWufIMcsAgiBuDJ6yz2XlieY0IPg1j+a6ktgss
XTCy4jTi/ko7oyeHa0sjmAGlIDO1NuN1/mUK7meXpIRUka0qFI5w3dSbcu7SkV8h+F/+MdFyaZVr
sooJDoaxJa/zQd5IXSmBWF98poyM/Q+7VK/KD6BU3qbY/CNyE6PyHv32iF8V5ctzxDQo0WWZkmSa
k3TlEKWcnReQoNToNEsdA3dS6b3pWU1/UkwAuCIhuECqQXpOJMqtx4n+K6hw+fqLQwAHbdaJTDc/
b9zxy1sOrCf3qi5HFaX54ojWoQ6lgvgAAKtK8KAl5aMgGaUjL+DlsXttNqixTPbQkJqsq9fNCXxz
TSWN1iW0xpOHLNq9Q9AV7rV5olKN3lufFOoJzIvnKz5LkphTCUCpFtkx3ELnRNnOXWopzaMmWmN+
kpVxe0ZNHeuEwVYvKfWcMERMgvp0X6RQSvyTcmoA+kU7vhDWYgHm1vehR9PvqyuC3TNU/RNly3Wh
hBpibPx14NNpFMusli2+8Ib91j4+SG3G0Qp4kX7beDPvtxb0qbkfUx4Lw7D5X+27Y3PdMvfkzwmH
UAVVhjgxhlPjTrKr3F0n8zCR6o1uB0FYsMGmctoTa5LYy4gpxeP1j8SVWrROm1cGHLxjqKDPA7g1
BaYaenNmLlBuCdJ8xOIYKYchyXk80PPa890odGj+ZpaDfOMNk69yu8MmJbCFcvhbF5XUT4HO5QdD
ynxDg7cGrlabD6mQzi8EULdgVMtXE3eKHsYPaqrJ+8twCcxOQQ4UeFz9CCKOX7NMuRXvq19IpYOM
T3tj/c7+doFZfd2BxnQ4KQR2iPLVNg8ZsCXlIgsx3NNYU0zzN+V3wZ5JDeheDsDsT9zfLq99CMhl
/WdZ3lYCz8NAOykqqrl4JBzW4e5VFIdON83hwWUm2iLLn7MGMP3/OII35WtQQUbOoBojxhKdEPc6
+OyPA8+Y4w+wtFVjtEdzR0izL4KwDPwTWCs4J7qvipnWf5aFC68aB50O0MwI6ynG1K5ortLz35rb
oFrxfs6ROqA3iJOs32yuDAe5d3qEEcmpCEe/Jg75DsFeXqdiimq0QAK5C2YEoXq4w/uLsSKiHN62
ku5Wp744BPcbetOJUGJzh40i8W435dIz6qEgPxXidpB6hXtEXKXnQcWYtucjfgccAWRWJpso1thx
5ifi9hfSsXUnr6XcZe1ynTFFkONRTSp94OKfNxFd0RA8iwNBGb0lAeZUAOArFOZSQqkxoAgnHStt
M/nklNQspji4Qp74FFZyLCDz+2xEMkzPLPH1e5r/1eHBiOtCqvHS4jygCSg5X4z9i/hPeov7DOqf
LubtQJVulT7gow+4kC3fsJ8ppNGyxUTHU5AVHm1TfS9KpzCnXy84NbBxS3zcYFhPw0KXdRLB9MoP
czv5Co0E3W4v6Kgb6DQ8NpDBKqwQr+7h6srzXrmt6qxfI8QoUtfGOmfTtna5l9DxTOQexDhaKv2O
dndT4XfLwyNVJU85zeWbODVxp4nfVtyhaKmMqTS+v9CHF/kGyk/WIUQnBjGyFMJWY6kDuOhmLIn/
4ZyURR6JMa6kFU6Ns+ksxSsK0NGIN7NQo2ZChHd4hGwm3ojuKkqGhJpGDywElbHao5lNu4dw0M6F
y6Qt/11jJmjh4zA/pqeo6poORhqmLKyAFLPrdHev9Q8zRHlPPGGvluG3uC6wuDMKgOppkqV5DABe
cmfagP7g8ee5HPybN2VdnJxyEIotjkbKPvPO8k371KpHibrThIfbJlsxUsf6EUtKMj4bgNA2Aw2t
VVmXEbk6fug0YWXKR55jVr7rhtWMvYdAodbGElMnLLiuJjBnwel/a6CV92riKbSWGG2Q59ZD9Lc8
LbgwJX2GFuPGaUpRZVw/ds0kooi/MmQuKbILdmcrnNEXMr4j/SsncLpImhan9mWEzYu8iFz1mGoI
bsBBAMGuj28YIso2nmUmD/fEhpJYr1REyysJHEmGpR0bsorepF5v5WTvJwCymf6LzbB3KLnzrFIx
N+mCSUvJNknxN5vvTqJ0GFhBgm4+fGLDiw6v0yy4NPqdgUE6+4b+PxOES4cIin2KNITs+12NlFR6
i6ni5pZF9LAgzjCPRI6skK5HEQT8jWX8W7i/9R1jk30DpQntX9LGaYFhhoZdSj7szb3PdgO54oTX
TyBwho/HDiKjsAhx9cSqybI9kv/G5vmhugz8oBJa30Z6Qwckd6tA4TQUbQbhTkisSilpf0CReAzt
5vxlp1dXQShS1frQlBAc8VgKx1B6Z0eJJokcueshSarVj10bWn96qz6jmPUjitNvSPlIdC+ttxmv
+g0i2j0ARRPYonguIqAI8kbMDsd3GO/ij+RvhdgiXDlH4OuVw970rojoKVvmLycNG459q94al55s
ecRuCHctX2IGb99TrbE9R1aqrdtPFTyNDgZfnoG2nttiQT/+WeL97aU26qES4KQwa/GHoloXdtdg
AykfKoEvLX5FD9CMDD8s8yQfM1KJtl2LGARFgZJDNw+89yvAx6AZx/f64KdCWCaYc9CUo3ykxT9/
rCevEOy1qLM74OPbAmcbUQUU4mpBCxHl/vUlzTofGfKfVsyNNElDUS36yx6Nh+k9RE1ImTedgyps
Y4VQanIeZHkpe7YQmZsoY5eg8W7SoGT77Hpt0e8DISyCyy2lJhlneh0YmSk0NnrF913oqJN0/Wnk
opn54HfRHmO9rSYy1eaVPZ8SvRc5ass5ZB5Qr3b6QlhUlAhdQUEO59Z5UQoL2plsVG3W3pnZ+VU+
az9G/lZguF5ZTIzohBQMGQo0vVC2NlWCflF/6xHdROEfGF+24ixX2KUSFqngGlclwecnXpfQ+u9p
IrlOLc6+MTi4qFmsY97U4Pv5MgVehdvmXgdEUGolhGA6xbNOIqAswmsaVzlALyuwMt5QlALGFWl8
Knj2o4knaDCJ+73HXNA4WVBJKW7cLK9951tA2gXjjbBGBJ3G6gxnnBQ0pxqiHtmVCQ6NcZxK+rFW
Cj6WOLHStVzCUai/LM62i58bGxQRhQoe1PMA49wDrqxrHaIgOXX+KkwdRJ3XbPXEyKsi29M+c7km
asbalNHkH/A4nrS90tv+YpwP9R9u+vldRL2RYwd/XP+3Qlwb0fWQ23jkCRnvJncmU+k74uzUSWMU
oTBeBmMc1tj6mBby76VZSRDIrXkrVIL4/FFAOEEyGwJGlZ5SS9uvIl20ExYpMCwdiUWUx08/sHjg
BpUSEln4A2KZsUOa+GNVSeeitkjaWcm6e0jtpgCHXIHJNyHi3qeFtFVUJKxCgcFHjiJA8o1EACQ0
+C5w3Wm7B3JCaqMuJoeqns+dCbWcf/hWg9kvw453iKymfakt8d+M1m8RIUPrnHRFclG2P1XHL1PF
vZQAnTpuNqDVIlWZhM35uuiaspA7odcCAkMcb6e7f3xFianK7cBPgSDzTXd5ffMs92g/RvDH8KUs
z5udlVWmoK59HSKxrAtW1NSbnMPNuDZw4NdAv1KFXVFOgtGFmF5hTz1vERyWxzojbahk78S8iDMy
GWYPeCUBNnL4DuYdzuo25jk32o3HQoaJTFgX5RdqDSBAcpgepr4+6HkKAs11JTaYeJnxgByfHpy+
Awsy+LISKo6vIv4hwgBZi6iPys8wSCz/moPD1sLTldp0MYrGnL1OmgGlilS8rck9zgKFNARUHWPP
oOx2C5bcSx9GWZ2DpSYUeI7yXq6tD2VZevpifgQe+y3SPek38HV4f47ZfRoed7U0DenYoKuzNn+H
7Y+ynEoAzX9BJXKSNJulcUL0MnzvoqgvV9PCtEVpeDh64MYXeHUJG1jxjhQBndTFuyiBYVrZY1jJ
XNckPJ1UJwPq3v4mnZPZExzsTDgUl5Oc5Z3cFDu1ulRgYM1i5vC9Io1n9DdLBg4ZLt7RgJ39S64v
IbWr/5n8758UBgBCIVFyCuWPUTO68XbMomlGvS4TiMv1V7ER+IHXN7G1vA9u60Kb/tRdL+A+vj/3
TTfb8zDPZ6WN9HHlKEN5/su5YYIcIzxq6T+TUE5c99+O6DFE+HOwFNmQtHA0daXEVjFss5YluT86
mrnUwkKN1MdjWxg/f1JF1ytk8N6jRaZiGmcVGzXBq+QCVapmaKDF4J998LDbdjMXPm6xkNpU501P
d391ruIci/9CCUz+J1jQHFe4tU6zrLv09RDwJcytXfUx4CHRM0HOQes70a7HZuhtYqaKLl2Z01FB
7aDbxqrDEAcOQ+FojBTQnLdWxAcrTcUVfTjVVYprzQId0WKO1H/g9CIgMocVd2ULluU0EoRSM9Iq
KIO8ufnxo0vqwy9bUN8f0V4QktCb9+PgNiUBmRbKswQ0GDBQ2DuEmp42QYTbi29VsS3JTb4sUEsW
g0pzNstFgc0BQ/AWPns6CmV81uzHBUfP4JmT1M8Ewq3RAexVTr9L/J4IrlbBSd1Mv7te7AhZ3oVf
3FADvRe6V2ocQeuNaa0KKiGc2Zdy1Ba6xEmPUYjjjCVJT/HJ5TvnomQeG0iWec9ZpVEvtltd/qL7
q3R5OZboDROwEvDvfaZnuEFq9/w/mGdm6dXw5C8AnTGr/OEUVQEEkcrYR316xHIn27HvIupG+/+a
cA9nVwKZuPK8UhkQlClI/dZAFeycLY2E8QUCdkivn4QqEYHSKrvqVYD01i5amN48fSJCwOFeuu12
/8D3zcLHY21QOHjJD7crmtgYsfHqnDBr8l/VpJaVGmhMtRe4cQZOGNZoPaUz8FHGsAKsZWrfh9Y6
LAbAuNr8vdMVTJhKll5ahGll12gvtbHXcml0ApWfxHW/n09e2NUxnYnbQ3282QQkldU5ZaB0knvH
J8x1tz1ildtXRX59PY4AxMQ0jhuFxzW3/E4kt4huygY4nTUCm4jchNi5sFoauA5pDFUZqTc02Ivi
426t9FWQtqI62xVgdpQCXHKclS4oerzUljXk8dkhYHJ14/qiGmxHbVnIaJEn/2R9VNkoarl/RPDu
hJdmz50jJh3euxhLGY5OiDaL1lpRkXGAp6Es1ihX124S7xsoF8AM38RxCZUTqujDihFzB/qjrZJb
hy/5+d4UoGvB4iU3k1V0VvDyPPiCsxbB1NAsKmCG8TuVTwlKrcv+t55YT1V7fcCn2v8gRQq2CmKz
QFOMrMoAJl0aXA2NCrZjfcL/bhmdfQPLQYxvWL3ZxX9+UkIA7mqGWqb42tKycgyvIUKSDHzGbn6M
Ak7xPukl/4L5/WXSIZX2VdPT/3UgA9GCQcRsEOD1zamm1PmD5bi/gccT1EEj07ZrJm99Z9BBpJLX
bSCobcUq19VYe0hiHXGuuFPuIMjU3KpyrBsUaD4Y289UxrAB+W8wE4E/W7ExeP1JYxQN7Qh9EJZe
1FqeL4JwCK7GpUK8Pz6Kq0BRn7D15ZM3H000ZY/SjyXp6Jruluo8BW6kkKUREZQTEzLbjVX1UKRc
ZuWmXMn67+wyLbx5Kgvpg18strfpwcegWlvX9qTlmig3OuXw94cmGj6sl9XDkN8aaAztjj6r5gHm
tOblfCJauSevt1WHdam7TJdhir4zd9MM6JG3bn88m9RXO2ByGS7dkbWWgnDsnSvn4mQOH+HyR7Og
ucM7nTh01pzeNPYFfROB2AHrIgPyy5cNgcm/nseFZc9xWmroqT0muD2Fz4GVWNz1CmReBWsIDq+n
oiZrkUCpAuC780ajBqPjLdduMJahOgFj5npssB6VB1KgGwTgrpF/KCkuGAGC+iLuJ48dbLbuRo0r
41EYaAzk/hcGHkVftwVZq1ruZ3tjeJOEgY+8oo/yAmnlb1sDvUZ2pYx4HtIbF8orE716kbmL8yC8
eosyTkB+hvNnTRn2L48C1K0/F9gzzFZ46Wq7g7RQUaXmhrJfgV08LRjBU6109ziNFJ588wGcGi17
6ODWr3GkEcMxLCDUdX+y7bkczBw5hlLcLgyJy3ReyTh9cJngqzw6FNgSdQyKPYW5hHi5cmTaJ867
e7qIZWYBBrkffpZRiLeAhKAxUCoxNZHNTUJYiRTw+zadFvGJScGfhjWzLT6mTv6YNfdHW6Bdy7ko
BG1U74g6jxLPQEVdKtohIbYlHlvUq21Sv9rnloirOekgF0caMAmLDu14iw2nn/HYf0tsQ5+hAEux
fucq7DqVh/qgGp3PA3eI7/A/fS5BJnrhz7HSXC6i26zH8TwoUcKZCRcuPU5yRFIDBq09SdDbkHaA
ppV6veduWa0F8C3gyKbmNCRllDH+jIKjcK8HuIzwT/GGB7tlcQH6UlDNmHD/HkT2qTFvnWRGO4ki
9E66Pxsyat1NM9ghOHLq39zLO0D97sBTgP9vOONSIsVMPl+B+VVI/6pZaQaXSsfBJEqhYkFMHukL
ytloomGZdv+N+ceHj0V3N8yuRmgd7gfiPTkAsf1C51eYmnjDTo0uZp2Lk1v3vBhi8sWoKHT1oX3N
nap/Wgg1dbkp+BQxDPbHG8ZpIe3GOvYOb/BPkFgBCWuVZCqaIi8TnlT3JoNi7hJ5x5i4esm2igng
pcp97cuFEL2Ljv8NUsQgBd+KEbEuxZk4deXTI61voMNb4Azim/W901KtvFb7d+NH+7BD2Ic33Z7/
mWAZwytubuIMXgrz55u6MWhgWkirG0zBgBY8sWWvytk6y4ZAnYJifTVF4uvH1L9mxpITx7ICKcXY
TMnPPC2af3KhFYwpZauOoCv9Ya7wvpnl3KLsDkI4J6vCnfD/E76vX4rDf6/VMCo/DbFTobOVb9HZ
zUYKRyUgDC67MYckYYW08DJIbkerweMn9O3ID6FamcGRWnuBVi7pmUiedRBcWclkdnqfCRDWXEtg
/ypkbIU/UCAYIr5OlSZrzpVu2Gk7Ktbk3JbXDPSXDJ/3Tn9+f3dBGqciRLZg4uuoqhD/8RHj4RT0
xS3BSCT6l4XUrkmGNAEf38DfWNGlILB8RsmnrHcdDrWYdKpINQtHO/R6Q/VoOWtz6RxIrzXuodSZ
PP1XqkZEYLOCVhsugX8d2a8hVdI7Vd84dnvDMlss8QWVDRm/bD13pULPSKOAS+PdyuKgTIbh6jD/
qExj1uB9jfawRJzpQP/gBr17fnJa/S1o9lcp2UsPxV5tduuDpf6pjSBdVlsMosVtHTdj1JAonigG
UC5twhC4WK/GQcIR5WKH/8agi0ohsCJCrrCxg6qadbBZTskVt3JwUfHGP/XalAFgiJNrOfd/9JzG
7fq5KIf5V+tHimWYoEtRGdjswBI3x+Kb1AFpr1sEV2gtDEwlFUT6nQftaAPOPUKciOyQRbAXSGmC
G88YCmoza/CExxy+444C2d/A0cYhQTykJm95HeuojcVUB4gUFqXT1m8HY63w6ly8NuwTJ17+Ib6K
2Gc0dyGKfs23HcjDnDX3Bgchg6HCqhs+JVkhOVq/APAvQzhMwhD6xKTU3cx6/pTSKy1EZvirWcj8
zDyfHYiXknFnSDdS12GPLMCOzXAUglu9sNKb7NzR0FvzPZoKLSBRsI2tr8cYBJcKUc3JrfM+KX3i
Wz/qysX+cfwWWME2dK0harYw7R8wrhSkKayajWSCphqfyNUgrB7I1a5FzEWcVDbncXdveQErJsAE
he3MILlQPfCGMv2Lerh1zr59Z5YA1gJ2SBMsc7gDUgwvh6/FZGyD9w8r/Z3hiEYDn0dA95vzn9Nd
M8a8Mk40kD9C0P3lBg7M1+ykpD2yfJ0NQ8ut4QzIOJjF2uvAe3xZeMRt3vc3NxYG1CJ1d38L2oBX
U7hDsFK8Lv3jkVo+GCpjKBVwOwwuuMhER57k0hZv4Rfijb8EJpKvPP3/eQJuXiMSKFrw1aKL/Uob
K/Np/7pYUKnh4GCtcJBeKmXJfBffI1ZvmSo8aYrH00QkJT9d1/sARbbZSX6imVQKMwFCXQVQZyef
fMt+FsjMUlOwfbFz1e4v0+dthVRoD1jCn8F0A/RvC+l8xWdokWW5dQtLklRIubvPCedb2dl920Ce
rQzdS834ySysIytR1k8XfoHhx6GEy+BiHvdesSTLIvIldWV+3leItmdpSKUp5k6GdvP4ufGYxGjC
iuo0/imR+rsQX8ibJJ15WKbxPk48IrOY3fbYRIcgFHzLy9EjqbK7qRiearp1rNz/Y8feCTlElce6
ejl8zyDQFo8S0mPnJUN5eZlWiJgZIZ7Iv4sT3RyOr2PpNl4y9tzhjh27y21F8fcxcTzOG7oqLvRI
IR99SjFHQIDBnfIuX5fJNBR+vcnmFuRSs6KXh92GwPgO14NAChKldSv2X4c+6fy+OS7RS1xt7Wbu
SBQZNjiTzysG35uQTtJYKeYAsJa8djB4tR1kx86BNR21TFAJcdv+S27Mt4XiOG3O9jaJArA+7ps/
dqWa4REkBaTEUTghf3pAs37vyn6sXRBXcg28+JKOHwJiVuowjWmJrAfxsHcERMdaSSudWZqQWznf
J25l3isiofBwqBVz7AFqgTAyzfvgQlftVdlGt05IMbsqePcTpDvpH0ZcjrRj09+g+4r15ivBTeBR
+mLUCCLZEgCkbEEPa6QuNsJR15lnjsFmHT1uGhet6sXOk5Zflejhwi/G2tgrRZKJSIFJt9ISbsRG
+WYNX7mK3rzPUvRsoaUA7lUxTVXFo6n04CDxKztwZxMsS98VJSQL3R/92CPdYtfaLrHG1jr/OqMc
yBLVBDGTAc7XqvB0MQRYI+FJWVz1/+nTMQuqIj5jzmsFtrkpoVfsoWOgDjgRPju8fOGkuUbW+LCS
Q07tWKOpRCTRMjymERgE/79PYHuyVN6KUgSjAgUsKV70VSYeu/DI7Ix0b+1+TPDL7QbIIJnVBp95
foOt6eKDaVvbJznweYaPsmbwZLQF3VfHUbXzTgeEfyFzD9jCJg3yAnqpXCUqSAAo8D1yjsG6jtZ8
NUvnK5sNsIxOF9MEB5+MEDEF4FI1vvhEjK004c4+Qe+i55tAMGNvnBj9GpapUxQrfWNfW0j/MSeY
mF1XwCR3/39h3A7kEnx08G6M9S6Wn0KlXAW7n/XwmvyqX2GNGnWrDg+1LHCZ7vq1De+IpwfafDzU
S6G9KWJ4/vKRZ7ss5cp50t/pDVsCMzn/Khc4oWqdfGgSwfonPjbk2zL+r2PXF5+CTrRLBx1cYR1I
VUan5hHeJmJS9SYJW15OUCKvGqG/xnYt4Rt8XFEVOIc2VyaZ218LSrknS5CewPJYymSZSaGxUwzr
gy3Pfl8o0+lMNsYO8EsiOhmTT8nDlrIrSpOhrQErLjFLnMIEzHZaPq2PoBM3ntpLkeXN7A0CJ17V
+aa4jeC3QFzbJDiOoDPsE/G1QeZEbWS/qB6YMQ6UtwInOKwCnuFCujhi7w5slgoiUqHXoNmkhQC/
2kDAl/ITgl1UlX3V9I0y2CAuVCC48l87gXPfBzEN7j36HVf5mT4qQnfVHE9j2K7ENwyWOM0XEjmg
dXe9YcZ1U92KGV9A9fjr2XIE67ZwuSrb/nRP8Nj76ftKwrdOxIF+OhWnW4/DgmWVAGgfyHhUklgm
0R654sKGFmz6BHNZyDI2MIZmiMUnP1iZtVcSCKlldflYom/TS8yfhdoUT5Lwo6yzxGIp0yCx8MVm
SZ7nbQUYvjeAwgIHu+Oh+iGVzYfHOPPq+VGEPQiIWeAaOFwD848cjRNscf56tHBPlD4ZxnTBPxwv
Vh1lAp+Y5fVwwU6PsEfvaxuXMzWtQcOHTHrvkwMTqX2nhcWHmqQtwlFfPJvWTVU5hacTY+VAY3/m
CIE6NV+3cEilU8dKFfJ7Auxf3tXdHKM5QNGHuPRUfbgq6BOkwkq4Mn/JGqzNqdtvHDIeiO6+55Ng
rXaXsvjGOx3NDuT4hWiuozzi4rI0whk3AGqr1Yc9ZMIbRIpfitDdfl10aU1FbadhGFakpyWDWCU4
KiiKPWEMoKdIc0QGGVEqAbh9MuCCgoiYTKCPdGqseyBmIJWz2w7xD1yjh0+0k/q7PY2bCcBwd6HW
M6cNoS0BLfRmLHF4cTb3l09tlGLREYEGddXJ/G/0sf/bxQ2QdohdbVK/ov0KKPQL/OYzyO1IvXtz
fFxt3pQ3xQ8atuHhfopY54wSFuUKoIO0EiJ3T9sioOQSTLoHr691WVRxE+xI3zC212bnWPwSRAYW
QcK0aJXXA9+rMJT4yWkStx5uYzcteGsEUGsz5bv/98mMWBVE/OjRvQWk6ZPBWk9DP+3LHrGUfMwV
0UJLKg9kBlY7QcvcBe9R9gs6haU2yk+Py4FiHjk5dKTEkSeUxCEcbGikD5ko36ZXglXLdI5I2Iw2
ne7owBk7fvvNC41gf+cE5qndcVeQSuBx3YOklzCpRC3BZ9mg8iMxo9aTL5Tn6RDL3F5GgkLmFKaZ
TpTlHV5KRUcTyOGnC4ysQc2krqkjKwtltDp+6NZ+2FQ9ZV4DltOWTWDORLKU7q96FR6r+itUsCZI
f6D++eu88bDSoitCWgw7egFLtym41q/etMxfS6/vtuOkt8X3ISsUqMuv+1XSz+cJ2EQEyh4Yu95A
6fZ6/jUtHbn9dvTD0WJxx7ODHuCBzn046YhMS5n8tkrpPJh1vr/ESpIOlaGztxX6fRygdl1C1ObE
RPt6JcTABnsXks18rhpknsynt0nz/ABwwprh0VwZidLViOxRjVAwNXOmCXbRP1ZNtAJn484eES6J
rsxhKHxtgOqP9xKOg7D7ng1Qiy0IfGBOj7h7qXsvkSNZgbK6ijK1zhRyWF7CcpBiMH0AyVFz96gZ
mq6V3BojgEf1v085gqcciaftwn9MBAEajnQECsbYG2cPrxqykisZF1gELCJV2WbgCfy9zSLGH6Tv
ZQssUzeWGjwIewhmHNa4yOGOZdGqLn17p+xontLAIMn+bbuR5SjCWkNEECBPpMn9q9L9VaSTON8x
nzE3+iA5v03E4ff48a1+G8TOF18KqtB6CRpx42GH/M1omEmSoiafHpPpXZQBpeyN1oYIyXa5sRtd
dGlhijBRbFJBWBek7In7605/1mJSd2dAFhN0rBuwDkQtFbkLwHqtgYehpabl2FPsYU598mpgEFHd
sCXHdMFerTS8Um0vtQyENex67niL44HnwUe4aceXgPUn2mw4uZkCtg2Jp3f6M6jqL0YRcumBK/gS
ITSFI9A+dlusv2faz3p1TznC4tm+Kzjdhk84LTmWOgugtN9aSYEMlWDU9dJLR8oY6aVGnFdOnDhf
Darm1DZSuzZ5ovEwHJqtoFO8VwHnvZoDe2B3ahpjaFVV5pPjV5UTxEyZwFKdG7LSZefoKZuKMyhD
/aytN9iWsaNzZ3UIQ7bQIZ4PHzdJEkEvy3RuZb8lBlsqeM+sQZFj6hlE8EGtJLsL7bAFYUwBgEU1
H+bDwvVVjuztQFpgGpU9uxe2Cran9E5n2KAlzcn5XC/BmQbNKzbGI3u47UBIQ6O+7hPyr0Wq+LYx
Ro3VEVvZXICJmBnWvBZYcVRYCXxKjKG5FGDkUvEeULek2ziGIBT12bXD1QcG0LP97PciGk/T1H+X
/R739U9+8xCz+SnD2arcbqUCGpnUVKZcVmscpOv9D53QzjCqxyXMy7BcBMeyYMfRHoBBvsskjBP/
2UlbWO1cfbNqKgv0d1l6Vf87XNaQbmt0PuwZjCLJUxmXtwVuA7z313C2tXpuzfq87MYrcbSjtkQI
5TSssSxdHe0Kk1b1TapmzBsdlENVL0vfDgqP8ONmUN1Vd779aFaoxG5ldE9QsXSRXz/FJwapvVNP
uA3vaAn+n7hcUY7ac+LREOoLEMnL7pc6GiJEHG0j4DTrDOapCqrAnVgj4q/HrXt6oQmE89KYKfwA
fxmvLsQbw/ExH93XQjygIVxQPIfsg2QrPoBrv55TsVOTXwbfAjBEVu6+4LFgwx5bTffw8j67pxHK
Ld4obfvYGtD79H1kLukg7VDOs30TTC/AklveiAgeiIIDN9XwLnt5RIJXeT/VCdPboZSdrv4mW7UY
JpnrLnGRRblcrADbCTfsIkccdCQnO259IQPK1F7GvCOhqdipyu5T+1+C7BKikAtFamWwbZnfdetQ
gEjzELxJXaxLSIlXgPNDl0iy/RfSqw9rg5lS8qkmbCbNmxiQzRR3QO4GNxnzssCTA4G6CT7WeGmd
7m8qfzS0Z6NnIJSY4Q8Zn38T5ZfsbsMHgQDgYhuCAOpqdcdaD3bO8s5g5hjNNHi2iVWxNe8m8dR1
4DE2PQP0m6dGZOCTJVkhyoQl2gLm9AXjwTBYetg9/LPt9MlBgQxUV33MOu6MxsjH/CXwDKlLCH0g
nY9aNLpqYJR0dLAy5+xeai5/bRtAiUolGwvHYXfdZDc5zD/sdSeV9wvVZF+GmcuZlrLU6FuGmsK/
n3luz/YMvnXDFJItnWsunjnoYTkCb7ILL8rzdntkqqA9B574iJ93qR8XuVPZJ5NnILWq+v2kLPLP
MOzfiaA5qzJbvvD57O4fheqGhq9Xws6N20TfgvCJWyi6E8bTFVC95Z5KWl1UzcOux659bTvb65dH
tizhC1jMZoA14yCQ24OsBTLEd5aUyHQRE6tKn/3VetGsTJuCRMxFzpltv1F2qaa4F9vmMv0SzKRh
ibvCoXPc/pcDc5+NYsr8iGjLNCrNqOwY/gV5j7UhWSVZBxcjEqwcyZP4IB8+uLSmgszF19Z+Vfqu
8IYuh3AVkoxK8Ov8GTYtqUUoXEyKXyyWyeY4cYcmyBwMUjEJOCmv+t3+qHgJwLVYe1mO7XCxUlG6
kAf2IRwcRCO5nsN5hfaD5BNLV3QKaenAhwfSgkr9JDfrMpYlMovGzGJK0diOOprfdua+UhbCakz/
Lrm/pWL3vvicpQMlW05/tVqg8BKEbmZtwvzQ3sZ57Irx83+754Csy7IOWhlwNxUg39egqZaqn6G4
12jJ3xHWIVBjTtVsOXdCQ1yAPzAwwq/gyi4r8TffibgMrihQUy5yWj3KWMzuM6R0WSGJEXQ+bJFN
Cqc4mxoOMZflw/TgVklGAnOz1/LrMyb6amsmv6Tnpv9Oh+dRpArpYO+LuBosIxWLZknmt+NK6Qkl
DG9Flh+o1ihghV9oL9xYSbcPjk75P++Qh6lA8QwAtiwGiFfBuWRqXx4cUrPj63fA+xUoLNngLBq9
TfVY+TxUHWg666pZqbXSSs2C4Dhp1gao0lSjoUjv6yIp+ywsdSCXSuY25gLTZEg+a9TJ0+7uRa38
0hFMA/PWH+5XvPeixjg46DoxgcyhlKRWWCrzoR74Iw0+zjsnk2YiCbaY/lZy8XrRHh2x2JJPXxkl
RxE3FFBk+x9xCh9YIAo4/T4rePCQHWA5bi5M7psxkAZC/bVxUCurIQliiUGrF6cSo2DOfbfRB8Xh
6kiT2K9FZZh1KqiwD+7eQoRfYRkTg5dgWgz2HHnmBJzeE0P8wIeIqpWBBYY9BDmlPUlg8TsJZGn3
XG242AESvDUAPvd4129izQPltxs6CLIFTxofxEClxn3uq57Dd4igoGRgOIIZSwHp2MBptb7bHF/q
DeKlC7FwzwYDkh5SQOK072O/WsPBOp16I8l/I/rpt9dOs1ZotbsLbp0DhS1rP9qCdaIBGyDkDzL1
GYJwSKj77JzBtTuMQ+7Oy2UVRMDxLmV8Tk64qfZ/Fu38sd5H+DF7SPGYddSIf/g/EYNbqUdoxvCQ
HviqQTa4GrrxoIQdLSSb8GamULes8DdzjXPd1QaHe/lL0ZsDSztluT6aXZt5EGy/I2QbxRFSXxBD
6A63tbzHbBLDd7rNjQCr+b751WRIl4IvIls1ehPMyvsG1aORdtNI5SUPl3hhuWvbY44VzV90LoDu
GG7a5RyMuLZUMEeDXglTihdrh6if0NvMcN2Tca3dq9ckxrgAG5IJg1x7W57/SOZApKlFcJ2bWC6f
8d0eg+r1XpoYLPbBNxfWbbDVq2HtUlzWvUvKZyIW4YBzuwbxltEfNVXhcek7gSYryBasOd/HuquO
BUzbVdeh94NDMEgG0zHadVvomAaxHNskv2dnp4/yJCkScHPOOj6w9nPLPVO1y1up8fzjw6lpQOn/
oZdxDO7CN7+phhHrJpsdbxK/7EKYmybrVZetKZisFRvm+Km39Adq4+M8e+BoC4LAtx2jRMv5Z6r8
S5e2v8fUsTRCJVd/Ocx06SYJW1AtW+rnPoDE520p4zVbGwZyjMrx/C5DOIgueKrUdiWr3+K5HZaq
ccGhOOrpkdshNl7NOGC7Gas/OfcAkHIcSHfg+s4ZCVxEnFAeXZSV/5ACDC3JUYm5gE1qEm0zCDV7
YV/HjFH5F2N7rLIxcQdrtNi6OWwDCrrhsZDE02gM19I0D/+KIFyC3c496ROHQ67IGc3mC/qSTGqr
0ehS4KV1QpfwzCp02wTN0IW42Je6i1llVphbVwsZ9MkNZmpp2yW438e3kZtaaMlImPYmYCMyR6oR
g2gTBLtu5uHAIJzSLXwrc/i45nohFbXVvgBFif0MNkQXt9hVHpHijcdg7ZQjUoZ5q/tGxnxdNpVq
miYOAPyOjDGQZtwrjMHGzp7M9KXbsqxrU6y6nAKihhBTJAgNDCWqYwSOqa2K/26/Gvsb3Z1yV+L3
lwJedeTWpqO2W2ak571gxPjUsivIYtacGNVwFRaCA+T/IacAK0IYKIC6VCpWmhKBXUF+Gk8zU9Dz
jML6nNUEpy26qSRjZdzELZyHHw0Au/JLx0etUSV0hW/CwvwQ8UmwS7H6xh2DHPpMsAcibYbuMnFm
ICsrzSYP1fqdi6kJrggwLhnWD4UOT6MPWewh66gznymu4/Xm4PJxKRsF2x/FEKSmRDmseRXWhqYU
6lv2Z/dSkiMyydGhEXiM2J2LOyO8sNEM2x/8bjw4qhpMIxi0EnlZf54gwQQNABK+IwRWEjM9tbCn
T8kiKq0fwk/aOki3d46JkF2AR2cfNoLmB+N9MnCUaFLmUUk8cItFd8uf0RjUkzC3DKZ3klZTvQP9
uATRX6vDrC0kNdYAxobkd2sLTNcLd0NZcPWufWRqL+w+A3f2x8N07zzHhKAI5NVrJe1uvZrZzMd1
zlrSErNh1JQ+fRoZ0dVoSZh8uLcQo4UjkktiPl7+BDkUxRNXsauD2nPPmSzIR/H5mtRPXu+Y5zCx
Jp8aB0whBi9/6/U9cRKNbMh3xKH/FcMnv3v9DVJ/aE7GIwX6EIttGqu2yXOciHhKoC5zGTtIOQ4c
1p3cTdNClXDhZmqs5NYLjMXYv4SmYeINkp/fEg67i94N8LWYZ+EPCXpdc4zfIt40b+X/rizs43Ut
LZaechIeIMoe1oEABLwKpkRANrG/WRLPMwpDRrmOHTxG8OEw8tejf3PcceAgTD8jlxuQRcdILw9j
/sO5+UnRW9wUZpXA14CPjTaLxcirve25Mp5dmq9HOnBE8+4Ov0vE7nz+3DIGhZAA63E/cgXVgTru
+7+Oy8WX18yZW5ZfLRD8l6d3oCD+03TiEhi9E+JBKRC9rNtUNFEf6tn8YTILPTgYeFKrxEG4n6xQ
WOifMP0MokNqISpseiloKgC7I80ts7eIhz6MeqV5D9Mp6sWG2f8ScdxuhtGj1221iUkI8R3GlrVR
4xP0fDNJAzUV86LA+tAyVqv29TJXLafGDvE1sbdMwx/Nzkk1uryRorDgzHq76DRwPs+BZa+KtwtV
vf7XSUwMMufUx4m/V1PXPGDYhU40Nt+72fzJ+6blr+y1QmOujSBmcIwObpsvZnt+/d5BjGhY17NF
azWERiztPWq4C9nfzIhQYmq6djlgrq+vmQX5v6DAw/pTrZvjej6nJ1KXgP9XeiELNmDnJ77PiFVN
945LxHttymBiH3kEn9CnVEPfgOOV9wMvmB3eUGFPTHmWqHTHEeVgn+gxqrZG08zlK4A0BhrKuBvb
pET0sGAcx1hqfjzDioxUwWD9CT55du8e3TrjttVROWzowx+Oj6zu1Zw71JcIpAaLq2ucjoxts0Er
8vYuKGhJkV3jNDFrx51pOKfHICM8L/l8gw/73Db2DzZJ2Oj29O1UlaZECCvDIapfdBvOyYEtWAWN
EDmNLc3o8Bu3Ztp7OSee3iX9EtJJrcdSrCQykRNg9Z0i6IqW8BhMZlabnQnCwmkPSRJIMlFd8ODg
u2hW0SfD1YVJvlofZdUKyFnfT8OT6HLJYyQDSnmJsOkhkOaHqumbHa2qBc+/guLobi92LXWpQ8Su
jzXtHwQLR8nUZxl5OEb5BLWk2ZjUakyF/yDhp0UvSFEFKTlRVpaI9i7XUx0FpUKwm2oDGDJE6N5a
nART51ar5E07LF8gie3NkCLt5ekmAjoskS6M6/l7+icVNBoAdViHctVNS54C46wLF4/EwkqrD7uF
yLBkvAy9Z7zVrbyL6n9965t3aM4CrvWF7PwvegdJhDyY26w8ErClzTajQLvAdrIoS/7FMZOctT/O
pPrXfX7ZOSchNSUScRqe7PZZdTmRMX0UctY6a8OSpKqkqO2AdHimPlF1KkQzw4bkuumWBFd9345e
+BbMw7c8BTFG/qE3oQvfxq78bW9dkI6+v41YJ14pBc3agKNZDIg+7EtpTcrVTHDNQlR9zco03luT
e2yh8HuoO/UHsugtaeEn053NjD+By7PEiFMjT52aJEp9cUu02eT2aMfbZWveRUxBILdUEBWCUvjq
GV+43d1MvpptKi/D9F49XyvbSfmNqemuIHiXg19bpxaJdn1aW27652dClY/9uc7aUdtDr4Ngm7h0
/UBgHmgD1N0o54lPwbJjo4zXTiNEOVrE+sZqWD1wQ/tobXVZEvYgseGt+4SDvfYHmDKxXtBoZEMd
PMbozvXUSF0LM3dL2k9ntZiMLFBNdGB186WkE0BTJUuQl4/5KqAHXabSjpSfSLXegif2Qckuqo99
hz2ry7EmX8bdcxdpP7uxPP29S59Fho/lC6jQ0m5ueSsZC/q0mqs6+K1qAOwYSs86FRyeXfOhsoEC
wm/A8mjH6Z9LMuUiTuWIm7vfYXWAM614glN2G+bSQURMfXLS2WA5erJsuHvSHmqPU7/MAnE9WbYl
mkp8FuQldqs5B/5OXrRnBpC13/8Lt9e69b0Gs5yKWfdhbp7vgKioyfBgy8rIB0CM+qDe9h6HCBKV
uOawVkdc9RtVezcOFnam7goLYBiM8j40ywCtMBcuDAfzIkx9/ZhkoID5COBeQ4jHdZ+G1QoR0e1b
SoOL5cfA4wWPjiXfwl50IdMwL33g+0CNPtKhRUZAltG4N0BXC2hKTNaXQ68IAcR/YipUJaURGEsz
UJI0av/igUYsWKnj7yvw17jjMQpahW3dZMd/ShPqEQB8Y/6HYFS3t0qJfGsUvWEkpLh9+QHQjBRQ
+h46DUhUvFKf5E9RJvVfmW+rGHrEdekIWSIFtpfDkui3ww1xBBOB4Nn/Sf2yyz5VtETEHzvo21ka
PHkVIRdkAyN1cJuip+XwE2PZebH0c8Z9ACeAQ+KYP44lLZnI0QfMAORsTrG9mpRbo2spbS+fie9N
XjHV00Y2O2NENlOQDmu61z+ySqtrEQLcqGipLZnBBeoCOEQjl6Sb9BeOF3/nepOhkm+EO0GC++oi
3xY3yK4nTVv9uZfpq/wJQ5sR3TukKh6/LDyyDzFQ0J+CSRRTOqq3kff2gSuYGwwQWSAQ+VZZ8+7m
Q/vjDTJfenhl0vobArAwcbf0pl1ezuYZg92EMqv1fKCDGDvNwvZnkM4izPH4YrdZWbqQJcxBUg6/
M1ac4nMpkwLKiuQ+QHewL7zleJRw3+Q6vb/Ga1S8XPcNTUVwi2M62oEYekwa4TF/8S3T/uKcVTlo
mJqHCEOqZTj67gC/7cfIZln7iaFQb1aWxxefOrSda49l79i8GO75q/vkE5pkJtSh1OcjdQ9j7I3C
ihsJYakNItVfJXpTAHS7D300BNrttljt5t86Ys82TAN989wJmRj+gK4vZ1ZBq808+QYaVuFCIoSv
M9yOVLOCsZz3/CWQ+IQ/AlQ8N2CmIEOjvlnUz6CX48knIADiHppujcLo/B1T+Hy0n98WxXbIxgM9
fY6nvnQjgGtLMp1aLkjxMfBtZX9AXN704flB2ImkPf1yD85vcdYXt1kDnQAruxwA4qIWBSICu5+S
ETxlwshJq6o4+0hGxPcHjZ6TG4Q6pqyE4j2emdKS7rnFZCPjR1uTvN/+Oigg9FUH7AexkOw4to3Y
pSuKoWaI61fU4Y7nhu6IVeqZ4QUW7WDduXaeUmqxpQ4jVPawGyFWdpyWL4yk0p04sX7oTu8Mc97w
1linOaF9ty1HhtVOdK82EjqJ+xwL3G1b1ITh11jFsTiCEIQz2FVDiY5TUcecuU9PNamYvU84+u68
HHloyYxY2zObdb5bDC75Po3xBarRMCb2diqC5gREFMv89FVHYxqhxVSY0tNmOH/HNsOqXD3EyZcG
O9Nfyqn+yKeB+rYxal/62MVydJ0utI8IAwFLpE+nI0wuqAKx2sIh2UHreiL9HlDaOQYTzDtv0yD0
q1HFCTBTMeUgWbhkmntW1qFxLkDhGwbxSbEJm6VcZj3hFH2uYrO30smKrk9At8eB3Xw0O33Foq3C
sg6jgB/8/wvkqugkv7k3odAw1oiOGNxffkAwcneg0ig3fnD6f49GkKLcbaufLm5qeRA5G0vplC7N
v+dbUbCW7M01tyYh6NWRWbTyFUFwWQ6WvpdnvkQexAgrgAmqnCHpAaLM2nHEj3w3dULp8303W6El
muw013t7fpllAGfHBL+jYp4ABjKwWrbd/lvuSo42TkAQ2LyG5u70akIOEam7P5I41XDOfhFbgM7P
J/BWOMnuyDfDJvWBRQCRHUk2GmkUlksLHhCgy0qvPRcyRZB5uU2yUx4Y3bkAag+JftwK5rOp0edo
doGepsefEm2CTobJ09LrFA4UYW6gv6nj2yZclOoRJJbzzjOD+2XXxRb6gCO54pdQgh3Lu4dcj7zO
HktRRVGFc1PWgXN+bv5c/peHcJPKni8BvqFx1c3dMLbo3wOa+WwErXtVY6aQFpaSIJYbKrlOZ58U
4RUBEE0MsOczaTY2SWjgW+EX60nL6RYPZ74G6HSjRy30Ge1q9bGftcKP/DCdvjeS3sGKej7wNOAn
JY9zeWRSBh51F9Tyvu8uXZAFb4KeG2nk1bK6KkR02Rp2hlgskv/rlsjfCKCTLJFHIMjxvBY5aGeC
2LM/JX5Z8bzWAe6sfz/kWGVnm6tj9+1vOsyrPsmfv46WK4G3lbj/0fD/hy/ZOLmloc80dsuHGEbY
Pl2wfY7BYRlQzrUYTucVMH1Df1gBKgA2z7zTY8JMEjGIjCvXEjg+hljG7zMo0aaamJ6vKtKuc/ru
H/z6kQEyoBNC+blp0E7kFef3xA8KSkbvrP8s5c04JKov8GwfJdyRR9xS7iM5p2G7DUX2A9eDfl5R
cOnL7DQj4pwiublNNZTt/OHCTQ7C62nUCV0XkEAaIknYefTRBYzbOXcZGfgLiIJHcyjobnBhIH3p
olzEIe2/eU8uz/B4fsaPKisJjmyJ/prec9sTr2MtOlBgV44ZEfnNIEko/eZJeQzxpb6tFrZdzlYl
J+33J5eFd3cGsartw1+ZX1BixZsKWkV2nm1LyXGIeKOW6ax3+vPwMdkynIbvjQVm+GFpBmUoxMo4
MRCQSqRak6JDr0gBstMl507YcGWW7btcADB7vb5XFxv42z+S8S3V12pQSQXrTSMMEeRjEdpfEKn1
YQA1zhParpbPSB4BWcXlD7jvPAc6Fa/IMCJSZB6QCEM2N7KPx5kkg3yFJBj69VMtd7CX9w8hx323
J/NeqCm4aA6rB5l9lQiwd8tCeFXqrWktOkhpLtVN/KSPoQWh9HImqEsy7GSIxmVxxNZs2ZvWddIo
AmYXMtFkBHLAAbuExAVu8/F1+VOiTMuu8Xq7tgNvFyysTdhw4oSOYHrLOx/hglH3OCxYbqHaz/qe
JjyBGDkVf6E9rlp/Y9wHWICUvc17VhWFxAg4J8kVuFemKJkJZc5TDkTs6fH4jaxnhu5Xbndyw6ju
zZqnchFpaByLI10bxfrwMv1gaaC3yBXMIkC96kMJ3GlxgJN/DiNM8n0hbnnkLoi9r4YI0QzDRClp
3XjA5AlHmgUjR0rvfRPT/QLcz4dGk3VGCZIZl9SGYk+lOpyR1t1ocC4rdLBiYJtQc41vqDPtNQ2k
QimBgrNqIgx5ij3cqLTCjgOAuHRM+H5CMtMmU4HSYewzTorGqVJnq7AYApcrINsA2it8cPVkAqDe
9e5qJAHmwu2wJIcvQlP5uAWDzEQoXP0OD2o0iKRG3yc6alFipb5pIUjxyRs66sxcr3qkAFR7o8/R
B2vz8sCy6UyzhW1xHd3VTKpbMvqyaqYZRwpqSAeE9SPC1JKtiFvedqYw/58SVOeIWsDZv7DiqMiV
9M4vcOgORQ51RGUvXVOWliGF2Pe1wovcLKfso7jHviHcKGCZX2mMp37S8LdK0vQMTSMLrStdxE6E
2Fni4VM5gDqeibRqup3rRyjL2LuOeyQsuZDtMkDLRcxC37bTOF40k19u8hI5MU4LE+0x597w+onQ
Y2M8F7YgrhPpBG76B0ECfL3pOyqkL8JdIbDaPLKITRnhD+s8h4heq3pec8/g1Xe4NOdV8gkgHf0A
LHQuyF60uAx/aC6jZtJZ0/gGpQds8IxO+r7i2h4Ee8o6PxysQr04QZxLT9RF9WQF6aTxY9gmMQMQ
cfbzVjwjCLY86alkbroCqR7Qwow/Ie/dhK3AIVe6kFfioTrTzL4rDZw3h6NZg4Mv6VvVcoVHRF7F
ZX5R2r6Bv3nY9prLogJVyel+LRjU438frL+p5LqUOKQt41sHmifSa6e5ou+lyGtNAkNxnCnbkZBG
sVFrzk6zplo+w+jipEUhxxX/RtvMuIxtvTua1nzUHgJwKVGZJdk24Z93ctG+sGHo+5iq5s7PtRU7
uM+VP0MeBBu2OojIm0/8hjaZG8VIcIuCSCblrBvVkvH9SpgaTDXritpdnDF+US5/HZ2orqaQ+rDQ
pSGp9qLvaSi6UfyR0ilfidoMkB1/quHdeRIfeFK9JmNyWJhi0E2VPRA9NB7gS6tN7O01WKiFM2sy
6AuD+RuMYIpJMjveCAq2bJ6fw67QSWgbgjXulFQwWye3x67gPhd3QJSQngAn8FQSIYuQfMeTgkYg
HFZyqB+j0Pq3Inm2JFAo8CtI8WzrgppxMp3NuG6ug23L8VMW+sWdj7HBwHgln9ddcThcLENQUr8z
2rE/tJf+iYUZT6I/71z+ZN44u+B0G0w51WE/7quI/eR2V1su1kLElv0stm0G6iQUS9Lt2DY6R9Pa
+nzktrmy7c4Zp2ZFrkXKxic2hWjJAFGbLZJwJiGnUavrdyMKV9s2NczlN+3UBVTqiLXHMqapszVp
NlqFPZ1AEMBsXOrXRPRExP4bmufmUkMLIZQMakppFlvh7Q00yhH7me9xxf+09FUGZqZaO7SfiivO
e4TDbInPYeagK6t9hSc7tsRv1pH8frEDsm6357eBRlAuf0R+9nspctW0n3MSOc77YnKW/lIuR08x
ujyKCV32b4KlRiKMAR8WbiKgJ++4Kp1JFfh6k3FLf6RbFKLy1hVURH++z44m3T/KaCCYWoW/vg7x
RJvwn58FZtppc5qEbW/aFrj1dB5EVVDgDJMb0++U+sN1rw8OrpGFEL/kByGJBMjeMObkklnd/yoG
cOXhXi0vvLxHt9HzalehLy2RoWJpc2xmpH+hG++XG4HIcrrDOlfAYIvb9NlBJ0/spqRmzPi7zNV+
CQjrQelL9dAGoaW/+ACAgGgoZk0xCrb9MI94UHcU4Y7beypi2vINjdJ5eOt7HSegr4YHPB80jnFm
rzWjOchTDYm+5iTgnIZO3qrYOsy3rtGAI/puTJ1oFhJIMFNrCFc5VekIztvx2rLoFkTywDJ/lnne
Syw+US2YBp03angyTvwN0JO2cbxvRsoLM6uDoORfWZL1AqFPNAZBBpHqxgcy2fxo2xU7gGQ014tf
V7U9jtx5Q1jwK6i8lTNFEPR7bi0gpPUdXZT41EGiLYgo86MUcbnDskAmV8qBw1PAALv9dJAQc2xP
t+RESO2uzU+GANbBGDe8AdcIJ1InnybIZJ0rU5aJjR56fOAuA9zqLLxv3IjLhdSTCyejt1qTBizI
MBjsmfqM0IXDSLmeJKUYea0/qSTHCnsISNqO9Scj7ZWrUfnJVNOqEeWdmvjuUN0/iLShrxOoGZX+
lTrj9FU8PvOiITvaf7o6dhM6LBr1c30n3do67odYvv2i+dOZm2MJ6hHq17HDKcs6a2BOx26TlVcN
+j+eVKXH5UhIniX6lqSpJpRgReMcuK5ToYFklIzQQROM0r9qgitvcExlKsdJauHGB4T38AfNO344
mZwvnnlr7fuiRzYuCo9VJLqL70k5QxfmtHC2EYWt9YEYKhOccHSbV0YVNxemGA2T40w/j2nPN8oO
HXLAkQUABpEFGniZRv/BuyBxKdeoR4596zF0E6IsFvziggzwztN9qPzOapkDMdNTf29NObMAuhhW
acnDhni/Hb+bn3VcIj8AvwqTCrYmlWFXEksy0o0Tzzoyr12fIKtadqZfkwxE6OcuJ+etLFhzzJwr
ORDyG9HVE4+vfvPFjQ8Xeq0AA4TQv74EpbtxARbC7Z/RwVKpWwCogcvEryVWoOV+J9cz34/NanUQ
QI1ksOsaXUSDjYxUeVHiqCv5GOE4O2TfB35KNx+va14yJ6P/VvQlFAERq8YgbKwJCGgcUbC86dMW
PtQzcU9uDsood68MZBtHK6HGa/6xrGuaGzClDO4itBXf1OPMeowwoHQ/okpCYHHQSQXJPgSwYvsg
A8mI8DrFLj9Nk6B3l/Il6Oup5JVbZS88YPzu3UbpQjYvT9GPuCvc+R9FLbx6h3hUHpkKXZZFYcu7
c8VdtUsgEBcu9g/EUh7oaBPRNyT4MBvpiNj66SglqIAs8XCBJ1uM5UDYAXpkXqnRf2vtRN1/v/1L
vfRU/hSaWCEVTFiXZIfC8DVGXX3aiFb+slxBCLR0cj7dT0y3E4aY307d4vfrUG9WACN0X3DM5voJ
YMJtPrJZFbnMeQwhMgYxRgYNrIYflsmkTQv/xOydZu86nbCo+trNnJzaYwJe28oJ5/DmUJ4d1g4+
5Aa4ZGt8540GcRowGITadZSM1aTS6vD3oz5pyeJndLALX2yG6bJ31CTJ06pYJ4ErbM4e7jvpKx6J
nglioOR40pAeKZynUHEI97P8JAG97G3dNcNOiUym7EAyTs+tjPYB0Xvv5Xt3gBW4L15Rz4RLQEA0
TLA+BFblQG2Fvk2W3FqBZ0oTJ9Ei9QKUR9Qt33qBdqEpW/ZlZDrC7+r39MmALW4PCHBGbbvUXlBQ
Bt7OJJomyBeCO0sZsq7RD8FsU8w7fZXBD00bYLZRJHuguPUYn4QstPpTp1HnXOB/V9tD1BM58n2v
xdkBD2lEkk4NCYAr401D83CbJeve3+rJ4pTkNYhpMNMYmJ4fSn3S5+ZYq9mrX27nGrkEIPenVD9b
FyibF1lyqY7MbTmMlXwEAIGRQubQqgxA94+JyOtXCCD1mYf6EO4L+GCi/zo3trAXWIZQOpZM5+7V
ZAjJEV4h3xxLY9603Fz54HDMaWvc1gay4GJRrUIAo6Fna7eah1ouwMCtGUkPPv8r86Xz60oyLRme
vHkN1dC96gFK6KwOGbeLXpKNUP97RqqDrU9vudddSdBNyj3DcxA6u0VEINsim0HJ3XL1rOebGNVy
6cWx6N+fbbOmzqNelNy+wm90YDrfmjEaMJFkMlKqfrXGtMM2+L+nLZiMjLM3QL5/RDRGJOnB+YwA
i38P/fIC11bsoF4+wgKYrtvNqGuFV8TUsmvRlmn9pALV8lqcqH/PXfLrPeOlos+jtQg5nLhsM4Pi
zRN4qQ7kfxQaneHWeEC3LgcoQpDmINQbFYl8J/Csxi6eXVNJ1a2/Kjdo8db1sKi2X3Idav5Ub6+k
pZIeYqNHhqVZqRF6tpoEiSddqrglv2mYTFQqayRnl1kuSFhWJQYfLHTqOze9ey7eWSdphXHJsCxe
j4RVz9khk9QM1Fa33mcVcrRqDFs1sLmS9Bru0QzAlqLZWnzBfeb/CjJfwnvRC9+810cqD/NLkbS8
GQoSDY1QHmxYX71F8UxlxdbLD3I0kVH8jNw/vgMRiq361njR8Zm5qlWYVdqBKTeGeI95el/Ce+rB
MRGfsJ3E/Ux4dFn/BLDrCZbBeU5Y0BXccJ0oLLB0Pfo0gE+uIIXhVbq+8LH2zeFuhJQpCWrPmy5f
Yg8iJTk6nifpVCvXemjHastTxg7d80OC1e457c6vPaIVoSZNqvy0+gdebsNI1d4pie7HgDqY9d5q
lBzo6iF4+rIiXbC3Aq52FupuxD4eVChcXq+tNWrvwvVmNqrzThqlJGPsD37aLkX/4udBtJkic/Ma
2n/JzjeLFsrcee+TRkFyk9mnzjI+c6MyGAyjmZeTme8PhQ8ObC5g1Lq9zipMLRei+/UGyW+yX2O2
ntx9bxvWPqyVOWRKRg394/QIQTMS7AjI14B6Fho1c6dxcIzJ+aQXG+qAHa3UI0lwjH4B3YWeOWPR
eOmrNapG8FMNcavWmRkncOKFsPAvziFvnZ0wwXTYUpWZ3WHKGbQDwk0o5Jc5FBjqHcP9IoE++NUY
SaIa1SY5nmYB8IuDe7zKMGFN1C/JVjvxxYLtYYKVuqKX7x2tbOUKPD1fxKjz5p76O9cuS/yb1VEd
qok3T/mbkUkfb3AzbqQK1WV1uL950hSiZagUxlMDionjSSnImWLkFJSirPboQux7l1rz1j9x2Kw1
wiH1v6dkk12OUOF6HyuIYzQ1sXff6TbDNAD2CVcmK0e+0rI0a01DXgoRel70kF+GvduDZYCAuQRN
HOxQ8aZ+FwQC0PvIzfQ5S6CwJKhJLxGACZfk52YM5ZbLEEOmOre6xxW8SV0UdwaVbCeXTP5yqHPq
VwhxFgSP+5UZjn5ZaLR6DcgpQtKhOZwC9TOfObsdMTSyNriUZi0NppO3/Lm1pj/xpDM8gaqg4Stb
x5JxsJEWVWbq0y134Bsr8oKxei8MNFqETBxG8jNsGY8dqxOdqcHc7vaiixODZXTG83g5uYszdihm
ibjbNxdmEUkEZqEZx/0G3u/gByc+GOgsnqws0KRagurBLB2TXE2UxDs9fSN2yjGJfTj9DXq4uLS+
WvxDHXi93j7oNgvsX/i7hsX1oomZRLj48HoKbLmpvjS5CKnJTZTxg/W7zovDCN2ryKs9jkp/psqW
rLFUAVUpskhgpkHxZ5ADHtZSGnFfV6nmou3PAByvmFBAG5EN75jULprsOzp2N4iq/MkXgh/uIIjs
So3Rb1XnjRkmkIuDw048ydNr7T6tOUpiDwDZDcJnjPk2pea3FIUpDtrFVCZhbME7L01X499qYqyE
ZjHW6pqWTAoS94vp1n3REqcqOn8LcwmWM4FjScOJJB9tyPBv6XQlGwhuU51reJGT4Cufp7xle89I
eaElekqwzM3EDc5wJC7CiY9tTaxjQdJL9O50Qco8XP10n8DQaKPbz9Bvep6JIx1+5UZJCLO0Y5jW
neYL9bI3quLgvZgF13Xga9jp/uxpIZ8ScvVVHnsK5a9xYvT1PaAuZ0vqp1vRY94D8CevtuIhs4g0
8wlYn926Q99Fl0LZiSlds3nyTYmu1lvthBJolFuf0bWXfta0Ih0axNF8D8t3ooBqtzhz25CtWhyY
HGYMAjvSRyJrJnLa67gEXkVWCbLOM6FCagxxJgG4b1uZGHC5AI5lugwuDf9w+rVZd55t8lAjDVGd
tnyfbIdN23Ey+Z5dpXcSbYVMZKW7c1ihO/v1V+nF2iJyV/zimF9Zx5ONS4J7UfwAP1DTfjCtOjtR
ExgTuTE27Qz1eLMjlJZiSrQaIR8d6Sy+4gPc1geGjdziWpRd/ea5b4Z0ACIq+kLh3WRTODUJ+ENr
I/i2Gb8vt6Ol5kI11tZUNTaS2Q4Tpyb7K5GF5eqBCW4hRN+siENwcv/d6kfGlyhYqKigCYv/DaQ9
/f3vJnBDGsyJSkw8Njd8Bvn0Xn87Z4qYq79NkBt/ATwiS7Wa2dS+TsFr6/Tlgg1p8cvb+vIZUqQT
8tl64cVVKDKfdU3B1Yf26U1Ik+Em4IbiGl3ENEq+rXSgLKWJrNJ0/lONQWjndO2Al+PIJzzSy59r
AuVFbEWOuWROZLKtF4A86cvRSjRZVkAFyhn/Bs46XH0oZVK49jrPN+oBglPEK7f4Z7VD9Vy9S6Zi
B1p8tEYqCt0/oJo7i1wCot9ZHWvfKyjkhwsLswIotL8IV7a+e1IO2O+E2j/60JgWN+auhcv1FZ1T
6bYnpa9ets6GQ1KX7f+p4hhuEZVrSiLIbbYAeqU+DE/+P8/A6o1HRCuP7zBlDlNEGSGV5zRiOsTS
y4G5gEf8oxbrHJI5MUkwcI9tOcAlQWQFRzEvrfcm30DgYUQRvdeOFv7+x2n41MVjLBnyHToMMKSm
h4ou1VYnUeeiNoQpKqzt3PNErHt1y80q3dQ1WfNHdRNxvSQ/4vYL16z56qogmSarPC/7WtPyUWZq
p9gfG/dUs6hnnz0Y8mGG0K4Wwht2noAv8X326QIAxWcnEr19Yk+wHuowXFFkX3VjiLLL/R57j9Ux
TljMHhPfixHYnULR89d7p8V+k93tCSDyL341Vanki8rsgpYMIumzjK9i2EkWwoL22cVuwl7C7Yq1
0o6PiPcA+cKTjMcqqAFuLH+XoZYh2sSXXLjaF8hPmMA3Ha93ZfYjfcDyGwFaPvulqHZGMKqXaNQ0
rD8xvWVK8EO+FsgLnLlChpuzZRXTzpw1pLOotqWc/GG2DjRdpmRNQWfkEyiaKIq0Rp2jjFtMgfTo
FBEA6t9dyxZVOPYMVuOml4UaJBuJkEauksOMpYvmPRJC9QcmHpaZQiA7GtO810xtb4cTVJo2QU72
mA1eZIwFWuL5AaYpchjCmGK79ifEKYdnYhZZbBoPu5UTUC3jaNn/V39fme+P7GYqhLu6zWCyDzOw
o1Ip28BT8ldIFuvW1rX1ZXguXD+L3/sHmHTKMoB5mNSa115H8VMtm8RqFsrvED/DrsyUMBgTwFAI
XZCtMrc4TuwOlnN6+7tXUfNchv8aPT5UAUWDhSAClW2bgpuc21eashbC7UzXsWaMqVJvMWr9/tC7
wwkPSrQtPYxTwwgBVznp2ZMjU6IB5Nc+eyGojZwx15gaK9GlCcLt2tWS+B/ftn1fWLF0ueX4KRjt
JQebLiPkbtQ/OAXV/FLxjPCX47S5LB30BtQ2YqVVmBXs9qHwLgiMJ7LsHtwiXYsXcWPrLJQ/iPQ2
cwdGpqNTSOk4fRUw/4vBxSKpuJC88q9Jemwe7S9206GKnK3QUbyj8EGmkJZgqvOoUrZHnrN/Bz1T
N9X7rl6gJdXaU3ZOjlx6hP0rm78z1yjiAtOsn9oFVQgkPw357uLk4G0HUDc9/F3xGlvPWGuSNamy
CAT2EkG6GJ74sIyszQEXr5LpmQbSaN4A2ieVSLbtdGWFQR4YaX+IMopiLm361/O3KmoUWLpsi3AW
azeZRIS6wundNtKTjoh7pxUyX3XR0py6g2/Fi8m77Pcx7Epcuw7WirWsgHte91K0kNaCHCmLa8b3
AR2khVYe4nj5hGY+0EVOWL/mT4xYq2spZ1AQvK0uLzIrekLXh558HZ3lwZlgxJSuuhMcnKanfHmM
5jkOFbUvsxUIVCmn3vRDmbcS2O+wASy/b2W86BmIOjxWzzl+N4+kTrtYjYRA0Hvnco9KGpfBAuxv
4FbNodRrXX3LDwKTaqD56DgI5UPzUx63vj4Nli6N9AsBDA7FNEdbWSoNPHwSzurRAiYmfc7lstv7
21IjsWp49pOoJC/HUk1Ch19NkCczCRRe5RD73IA/5FzUM/l54oElz+KpST/FwSSV5fHYrOHmEJHF
9YxWgjhIpmV9dR4A30LpoSBsqPte0u3rSFcppic8GFfObvm4LuPdVGcQV1EQSoD/3b6YKT6xTeU5
BvaW7IRdUJ8SvFdkHlc2CLCUx/om/SZcJpR3ik6j1G1gPBVW5sqRj0pXUqTr3hahZ22uPmO4W1sR
mr2G6G1+H5Ye3vm4OgTnm42R//Xua+T8Fdg8ZHA/GgxwnUV8C0EI3GFMZTO3NAjuaC6vu5b9plCI
ch1JKDdsJAY4Gj2uWJvBhMeYgDmF0bOcja2SNnVBRmqVKyyv5xnNZSO2M01bWIniIRLOQNAIDFmd
iLYGkD1rj4e8hebtEGJbtgvoS+r/LV9DbyYaONI0Xcai8tWaIC0o8PTgQz8HKuachlXPgANZ+zOB
lkMVeC4xBbStjNaK/u8K1ifj3RrQb6VVnOjV8a6W4OX+8QAl5nchpB8R3R6XV7Y4lkHHrQaMFHXS
kf5JUuVMnzW2RMKfVSwqq23x98uEaRqA47S3NWcBEM7cftjxkVy9f9IMJrAWJRUCLxvfgiG14Mn7
JTeQuEQd0l1EQ9HOO0IfjG0gwY1DtSU4xAyhqtIET4dkOmrm1M6P6fdPAddbSQhKvKHfeSHSa1bn
9u0KVHjjuG8tUaUUYQbxzofQ5b0K11Hr+YvWaJ7IWujrlYyt79nmD6SV1XisCfVUWKAZ5wrOClGC
e3JYsi3l42N6fL5iMtbspWolI10mu0A3gN3jI1PKtq7IcpDAjWojGHVi3RMM99W3iBIMoE4PTD7Q
+3kpwMTbJfc1uRtnEKxb0mDbBvNbSet5kwtrQg6QG5F7lCmAdtyCVzpW3lx/EdertuJ+o9zj+7Wr
jDoEYMKJJPvjRl5xsn6Ta1Cq4IjFvxeoMQ/bJ1X2+jl2wjJKY2sRmejnzitV+91yIwEf5mXz+4aK
XxRgatnA1k/Spg4aI+7YQx7XDZQVyEp5bl9eI5neZRQdmxmTIZ2gdERGlz334f7PPNyzIl61E5RR
VBgn8wXEoBqqocAu8V61JRN0iq5KqXIvax9Hcsa8je1XYAqKKT580AmnhF6QLMM3N6RkDkLv0t/H
ZMQNmLj+K9qsmm6kvT77XgBtUHMv+K2ncTO+5zv5wlZGBTlnfxM3AGIFaddMYojPZNgL2s+X2hMS
DFSlKwmV3m2LcjnRvn4EAO7KnbAX+G3e5sZbqwcwAMYjIZmcsSy+LLNOd0SSImHP5njWlgShTk3I
obM25aQenji13pU2ThDz7wNQyf02Th2PN900034KyPdXe3NKPn53ib3pfA20jvikxoSXJVLLu3GH
BZ3Kpdpn+kpIMmdrz8BAFfo/Ai7QcyCQjcV5s4eD9GH0n4ZyjspHJkF7I5rElnswIcSJgMHvuPPF
PNVlLBZ5zeP33rMFLoepmlWZZpLn9w5vEKOpQUkKauXr71oj2KgHdWQHH7xX9o3bNf6FpgOr4C9S
KuKLrOxne/I3+/wt0Z4IA7kIMHV4tGc3mHh95TW1hSJQeYYUaW6GewA0BwwGYZgkzU39gDtVvqD4
aZ2pxUzCOSNN02lB1ZX8u6zfqkU5D+MsNUgOTDSJtpxKd153Pwo4W/VI0GQfhhhqIgnPfw8n4ujW
8+8DoXmyJsfVjyAkWN1B3b0/KAFrSvQ3IxeG4CAfZo5E2ARpmxqD1s0vXx+7q9GmlPFboDHL6wdR
RZpdCQbo4gZiUbzNS6X6GcEVL6KbrH8GWs9CkDZMekcBITJCv2cY4iRxl5o96tO5fpuRISZcN0TL
93NTMhhuUaqxBSorv2tEHklKrtsEoG2KS1ggRsQZJ80DLGKu8LzyfqsTCV+oep9ApCCadevZpzXf
CYBd6j0QD/JIbcZWpocKrkhd10zz8u2yEQiNRPWmWZTUAl5an7SWUqYv+d/1iLt4BHS6nBm5TYte
sJb8dMlMRBbPur3uoa5+RMIQgJ6hR/2baisor8FDP8w2ln7hTX7EisilcJmi3qRDDBYIAR6wR1nR
VdbTqL/t+hz9oT7/YbZYRlquAPHzqShJTFuuOtjEcxBmBWvUIJW+9nb1udRiRHvUMtCBojkHlKdg
2UP38KCZgHw5/l/Sw8Bf/IcEJFl8dMSfO+YLPkFSGfxb+UkDJj03XbATKsClFRAc7nBI7Zf/5Tly
iy1beHwr49TnVvgA658X1S1Q0KBsniaPkKQ5fIsBAhTMqAxvCHAV3k26fIWyNMSsGy+QRtNiAEuY
TUuHfyacyR/8nJZjsWEsTtBrjmAgazMaYt46Rh3U/jxtxv4G+JmwAIF2LBMsAkAoi5GAHvPzCMxm
EAJsjqPq59rse12v+dWNykPdNrjHM0XsNBmBiBbSlBHjKqn49a3dMr8h2aucRjris1qeKgA8dWUE
HtOWmJi6KLj8yOywryzLLIK3pIj7Dxa/FtgoOQD8bVXZ+kEPWj6AU+mYDVHWVQAINGBCYt8c0Nt+
p7woGzWQtgXl4bCbpaTutOCYYmvzPvf0sKmPL5KSbJ10E+ehN3V+6/DGqx1dlYJpAdPRbt2cMqCc
TMrvZNhkUWIPl2M9CFPpea5bLk+E9qNLe/G1yxVqxiHuhjutjeIGvoGk3+OmA3q7YFwjrFrQ8MLz
bNDxrquFMOaEbfH4osztLM66F+yr5tgB9z0mzFS+PI+Gdei5PvWo4oZbC+6Fv/gFI/BgZytwvOzA
rUmnqod3DQpgbMyNxmKcv+NG+mb29kn9iLQ8bTLAOV5Dw02Q3yXXY35ey9dOwWCBO7lhoZvrxwME
+lMsNfKWy/zQ7E3eWe1G2PzJ0RI+7n3VUVYcnNdjbGpgt2uAG/SCH9fOrX+uuJ//z+MKQAI6xr+5
ch6f029jlGYMe3hrkTjkat2/bRHuyNVC4pAahP0MwkSoIx0oMEGSmz9YjkQc/DoZq/KN5Umieq79
5QhtA7LcAs9136r/XOeP/7zFeGe6wXKQ9hNpezypA/cXeg/9PdtHdvrIrCO8nG6t3EWwAFhyaa8P
cNFegGb3whvfvtNdNBO5qXtoU4llzGCkaid9HfmG+LLOrXCIg0Z9iG7ZxE7lwAaDdbSh/6uIByCb
jq2uJkatH6fD6aFpJe6nhE//vA26GLkNlPzm1aQrJWy7tiAeB/o+cfJfF1xGX+fBYlmWAjvhYYki
U6FL5L+knzLQ4st0B70V+c6p88/2mz1S9Wx6jhGA4euQKUehNvdojEqsa87Gn1GhnQ1qPWz1UA0q
jhYWiRZmoMROEvjxL34k4OSUh0Zww1vy88Gj7U18VXc5GA+5lxoWBPOVwWKzYMeqbS1R4Esuz4Qj
9+Mzw/Mda+jk3qot4a4fBWWasgnZht12fhz32eer88i2eB7NnCqkPdf7PxbIyK6J3RzgGKvwYGrd
yRxKRQyv1xXlIvESoVA4ZnTlMe+kb+B5E/oxvdD43PW38LzzA/V9Ggjk5yadPS0hZ9RFDfs5qV3M
1ikHNI7GJCRL0CalvEYshShkIwKcaMJ3A+FzvWzlbxTX8CS99ml5VM21HZImv7xAMjtufv84Y5ab
sAJIa4NnpIn3SV1HfUqCCwHHXMhGFh/SO0+vWqc8SLtFbrHecv57uzwpQBHxlM6jMjdjj0nrE18p
E5wjD0L+MEObdr7WHU0ri5O3xWm5WkQ/aTT6cNKNt3Ti7mmBh0hGdyE1Jr1IP3CSO82qVRqBqjUI
ppzLNW2l52AMXNlpimDMvyLQvk9NxIRXXxq/h4d/h6c8wJCXfVCF3thu2hWvNEjYka2gzYrKwL2o
C9T+T6EBy+gkGBXlp2TT59s0KSuX9zTK1x3KV3t+r3XxcdgcaVGpCBhg1Y4WbSv8gIsh4n5fFbeJ
qHE7RB1KgfLaZZQourbyVzDkzzLegnoxYFrQbA+RS21tQH1BUmlUrJmOZrEU415qYLaNU85nwRhb
sOmuAeGg49cQn22L6cRLi/MkkvBu1S5hIM1r7Myuif7mcWpbwGgdOBNot/QCM3NhVD8iYYpbHsSy
kDY6PwLZhfJ4Yot1xKHSpXzBxtgICnfTkdETRcVd8hMUnd03HgsgfryGyuox1FZqHHUhSAlH+eAu
6HxcKFZKL8hbE+/EKnh8SXzug1H2scemlTi0KNBrHp/f+Qt/gBfd7qVnkOJ5yjFapYsA62DCjHsh
FanSxz1zepzVMFpsq+rn3mbgdqgyA/64i4gbUTfRQ0zw+a/c8dkfPyfulU6azBaA5/iLHtUCTmn0
0G7Vat4VaVNkeDm2Kd4LnJteIO70JAdCHofgxjtn0Qi041gF+HzxxD3QEXBeNCbD7C5dDrrkIdn4
qrCDG7YW9sueAKotfdZa5ER8aq/UQnCCCj4InXly1jQts0TEhxC/HMsy8Gm7eMa4Hzyg7/ercQvm
TAApmI/FoLU8DjKul73w5BB3tlj3juU9a29nIKM0h2uknfBZFf4x3mMMfYP52mpyLjSDtkZLFx+I
v00guI4A/YeT4v2tLs02gsWl0zmUyPC7JxdKlY9T+oCs2FIEBkTjeyU8dUIKvpShkBRDuKMtWrm2
yyM4roSTdmS9SWh4XGObIai0nRWL5dLkjS5fBO6KBpjQ2v6TuGA3iP0wc67DURpj+7T9Vrdelpj+
o+JN/6DuqtA5UGzfOzAqcaQ3oLdu2bB4TgdOJLfDecc2Z/PKU2BQ18hXxvQt2icWmqzzZqoig507
Hf73TB4OlLj3MiJcrhxlzi01Zgl4b21B19yAVEWFA8JaeB9xqwzFpaZZ1zBA1SJMedaQpn2eSfEc
qOwpwVpkKIrSdNv6v1iON6kb9feYshUY8fY+8qusMEKPKNru2GHVpFUQ0RkeIsmMYL31s2PQHgxv
aFPDMY+hx9TxsWZPJD0qoL/eIWRMlN4eGlhodkEdJzf8PXa+vyBttSlqlF7urexcMiqcDOYaEELI
rV6DrZ/LsRI86rKkSkfLtOno2u0US5GDxqbf96EfRm1U1NTrt4UDwMpIrc2h2FKVlS1UkceiA+rb
Oc7ODNnTK7E7UeKBsc9BX462EQmxUNfRgOGybI8Y0JXUUcj6dzd/+iAhk86RdT6naPstl7J4YE1K
OHR+1Ezf+Kc76StOnLjlWkO4Zrr6oeuqKFrDV7a5irhFGA2lxVmzGHa3hGl09gvjFc45pxPY40On
a30bl+n7O3tZXirzUx7GtQmOIm5cH7AjULM9p/LS2E9JBx7yLpPydhqt8QXvk6vgFvGSBSuJ8YBU
HewwayMzP6DMSHjYzK1yS30janYObUj5V8icS4ABNIKpImOUg1xH5pn9etHte9OwQJpI5w5ceA1b
u5j8W9b7i7tc5yfJw/SiSSeF9Tk0bjOWy1yeMT3NHP4+umcZSl2cqbomZGeZ+eJISY16ATtLgTMn
bGjap0Zn9bTxGSlxv+fPvikdJcPWXbST4jRPJFfYgSBqCDE7v7rv+IoAfoskHTbQ6BkUBbiuLzsB
S4JW7/DARhT+gVnMqVY2R2aYMSrhU5YuiUaUh2uCFCRsmeMGR527NNayemxF9h6CgY5q8Q1tW9XB
21XFSPs99NBXPePyB8Ib1P6Ppsn3VgH7pdoBUMPY8tceF5kWeNUGNpHVk8MlECp6EzvQvfJ/lVih
fBhEWTR8wBaDKCuuiZNXg1XITP2Y47k3Qa4dEumKIy6YQFG2W9xz1v3uWHggDqRSgPCthizHyC7w
ptJnIX1YKCK0hTXbOaT2BCAGQ8OXNqO+6f75qh/plJqT4avVWIH3sSy1qoxAjPHaDseLdhPWaXZ1
vpnOH9yX2LAB+HvJDHq2pxAsSio1qQfOsQ7OaapuvP+ZgbLdjlPt91DqZB8pv867/Csr6jcR6Ayn
YcP8n8ehT/dpunt6iJgEG6IYVzm+f1bvwLy8QbYctioRIKPQCORBsV1gpH0SvuyT9VBDandPaNAU
GJOXWxzzx4afjDfOa9DHDPYytG6TPrpHdVyhpn7S4Q/W/+Ju6SJ2Ptvtoeio8AQi//bAoNV/QFSJ
7neKangHtHdJLb9fRSvQRC+2t/EoFHgLmq98M3OmGu1Irote52jrQdvE6flZ5YFL8KEBlIMo0OWQ
h0qS2HHCE0GZC1wdJH9CCng7adonbbWx7fMvUq5DG20kQ3EvQ4dg65XSYgRtItVRE8lRiTR4qogP
9rPsE3/wu0H9JIM3Z+zIui+POfbGYKbuEtLGfAXYUn9pY2PAg8iJP0aqTmLp1NjG3ytd91nU2gpP
oqL2nz6T3E0eAUITYiMb4bSrj+rd6lVzJj4qXS8yOPvHuJK7byAIfvX6ILJW8sCiCpzaQT2SF3rl
MVrqwPdJh4qvzJSSLkvCHsTc3+7MU8oze6k6wyx7Zm0PlWZRWYrp+1UfAhtN5PFX9sVuDNCpcP/R
DRu4GSQ58pZ1OotlHzZ5O4tUpPTenw27rDMS76L7IEQtKdsskweFKopTPXLGYOrrUPQEMm2c3WdH
uxTZv1AgnGLUMzplMS/r39hsPF5RzWyNh7mMgH9E6tjyQk9sZRA97NHUR3VFxfOI5aYpnJdxggBA
iPwoVm3HIY2YuZcAGfK+pBaN8yArMPps2N9fWfAdBMGLoIRzZ8XMxshIPVK/a4WaLK2lVuzHd8i7
mA8mhsYKphePbxQQNiD4WMdkWcInkj2LwaPK8IVd+TZ+jomX9627UnvkgsiZrtgc0/EFu5hZ4bc7
CK7wfRhK703e+zBbH6JAboLy5dPm+L74fQ7RpJhT2mfT8T5ckdBQk5Py1mVBGeK9ZNlIoXDh6zs4
6X1qdxVDCIvhLkkicEWtKTvVKoUgXfp13h9I/t5nH4U6009u5NUHC6NDVqD1CwVGz/9wDWRLWDbl
Ff67oCg/8Zj3wuC2C+bcTXCFuEqfylDi+MA+Trc1FRzccUJ8om8/UtfhpBV6h3bVLKvkcO6m4KYj
kOHnNExJZH+abmn3EjC+VzAn/+ErfL7VSKrff+dBlt3275AKI4wG7UL+1H0fJ8brMlE6S/WPuPDx
1vqd4n6DZEoUSPMTJ0voBaFmoxRmLZn3ScxsikITYUlKsg3ngzUb4YA/bYvcqGMKMdbCJyuF1rdg
3NUl6M1RExe4NQb+r5lifc8J7t0nuNyvVhFDYTOVkhB8g00+xGac5tUPl7tzg5x12YMCsBgzfvet
Y0RY7QFRaGumnZfnX4kbvcdhVeodGFvqAyrxbAF59lwdnaSF6w6jXz2EW2rhEGUv8aHvm8fdL3/+
AGfA6zgjF7DgJ5Vn3IknUKiHjlqTGqy8em7H8gtiJnK3ity5ddQRPW8iz2S+CL+8ismVSs82HPGl
2ante70KoAbkDA9vu5Cw2OtGWCXnQyKcso5cnrLsELmMKylkFv5uq065m/aBMXfJ8wxELMWanSon
n1F72gcJ7YCGGVqxsfFDtgx4AqxoqUZlgJK1iabO2nyyBDCh3tIVkZFzG3deTlLCMyYyIIs6SEmK
LbuEZK2JQ+beoTG95Mjd/0bgiKQT5valfulQ9u2NQYoldyxiDYtyAD4FlP6Kgle+GfcRedMf5lRm
9a3Cwxy/AdBKmjSkDaMpaem8tR4dLrabo+acT3OWVCH5/6ukbK08WbgI8HEXsj4TPpcw2k5J4410
uzCa1x304JGyCqS0N+V6yOBsom1mOP4Ul5WjSuMHINOjS1nrtAWkil/oOkNJGiQICguoQP8jWBis
G1ry88s1t0G2cwQkzifOX2jjIWUHshTeyuGq5Bn1pKE5v95hkEReeJBDKh2+WNNrGnRCdH0rZJmr
f8fsgBVQ/9xGpB7/YW01pxTICMGzAxjAEH/VKpoJOyrcUvZe/cLWMsMcyikr9ay5xNG3iGhX6m+u
tIGT99qfxbUbQy7220qkPCqpi4OoPnkMWLe/19IPHcX+/Cf3HM0VM0x5H6skfiWPi8VReSPwngsa
9/w1/kddVpYTCBVT653EIy/eYg3u/r3PvVdVMXWY1A2By+jN/12UvC3As7Rcst9VE3mwdwYATyAj
PU1oiy6xSdIItxFGk3EV/ST6MbEu47abSHl5xLEqTSXCK0ejoBu2g7oorZ4o7v92/kxXk9XeMcAx
715FPiUdGwNiQqW6zls1sUwg3pkRtIRGV/BAH5I78YunWNiNDuvxvdZAOlLme6O59irSdkj+DK36
P6K/oBpT2S5MSMFLztoTlRntY/nSGmQ/bkGrfxapyZAlb8iaMYsq4i7USLe8+Q4z3xiVloB2w1Bm
uTPpr2TqYtbKeLFIBjIhCUaOApULecyYJve5Ctwdtg7FTobtnkyYge8O5+icgQZFDulprCZkjAj7
5cT8mGwwgNZKrqieIUwuF4FZrJoD0739EhEb+GUNAECfL2BCBW26ffURdST894FTBrm8+mcTaNxd
ZVgHOT81mLLHQtf0fU9Zxl8cq5PM74WdYcSELUhsFCHFHsEDWxB0fNBj/xXg/BbdQtiRbHXPb1fc
b3XsgbTpNebXKh0vrnoVboKqx6GtSyk1EeCh8YeogrvPIHi3c8rBVGzpExp6T8sJigCf1Zx+G7Fd
xr1wWYAr4x5s2Rq7rEdRYhrm8Wfhm0JbeBmiEKqWQZTN6amZd1CAmnAnmBDk563ACvJrMKVY8f9/
43HWYDCURMzLxAwZy0GnpijKl3x5L/GlnlViJMBGodHKClyMQ8+2y8avsPsv1K/+D5s6uiKdIdS0
yLnGLRpq/w5qp3K2Hd+IIAXZKVCHm3/2c3JdyThnBdaAwFvdEJfciUkTTTQs/2dSwQnpoW5O19wr
f0AjAR53Xj+Owz+j9YQE52I0HZozDo9bgor1+fDrbyFzpgIKTqI85MOuDV6bSZq/0yMY1u8EtDB9
Ojua9/xZipBrqzQ1+v90CBXActFHUiBbFDYFdgiyH+McAYvXC27ds+dqlACpFbWPcdyRSnHCP8de
VX5oxYy/Lg8bMKI0KWM2g6ArK/8Wqh+dX2ISfRxOOqapcr6+PHbLZcHdDyA2mtt8E0dFuIhdFo8C
cbNNUoJr+dbDJGAPZ/PXl/h3WK5Oo9jmhCOWDtgwRccB4eOz7ywjCiYFZF+uDf6lGMkaExhvBAby
xX1CQB1WZOGFelzWoEYK1lmRED8v0F44YjQlLWM0DhPKKmZgAhRJe179D1HDDbTsgZfn0IxuJqRl
Is9VORgaEYNLJd6C/CrKnhIVAJDYx1XHbKN8StbobDH7gEx/CR90lRa7wsRXUQhcvFVlkdlGKQS8
b+eBwWxXw4MojRP+OhcLNQAuIY5ZOgyR7xVe2/ki0aNdHdWY41lwz1uh6isD+U8B7CFMtH4dwnwh
H8cwf4pFPQC90DsABDj4ndwrq6Htw73aZ+H1UTBvSVC4GTj7LOviB4Tvk+D2/CaZZpGGP+Dv77Lv
mykF44r2bxB1qhq45HdZNGpPDnPpnQ3dSenp50A4m92baM1WWgE+gE1Vjjr/Qd3ZeJFydjtUgUZN
4dP13y6+9+5OE1GXdTmpz+nW3E9o8df7KwjoGbCWBp5ZGX5AZuE3mggmB9tWGzvmMd32Wv8Fym1c
69JCvk/HUpG3Zhm8reaJt//zSJwFuBijXrMfJ0dmkRL0NotjUXaEjQ3Hm0K46HnmFIwt2f6zYYWO
w1di2DIIwcSr9i44HTLRvmqQHiN5daul2Wy0dIjQpHodSKLDG9dz2z3mrn78VCD2Kh9B6hYkhEMp
Woph4bEnfFvRdvLfU8fnhFaEeglN0JFBGhuHFSyzWy8Z7msajSTiRdaYvjtU7wwksrF9zehGiPs4
bxzk/UysFCD9OiYk9lM9pkr3fsVv+WcjnyaeRm6Zt38Jn0P8Qk3TGUtqz1/kJIMBhUp+bTTik43B
2FzaHx1xkZpXAeF5SMngz/hTW71c7/Uw1mm5vAo8kUOs4hq+liM3ieSBFrjhMuGvC6WCSTmg1rbB
IRfjZOsTIT7wEB28nJ1iY7OUg62BGzeggnINrNM/sX2m0I7M5YU85mozk1io/3O+3imHoDz7tXCg
qUtJHBsfGTx23M7dmPrGVWwZy6biUrFmJNMXNUghxOBrS+uoJq1L/G+R2YqneZxykkA3VPKl5Bug
yl+m8ydCycfiT4VYqRi9FGoubiL+DIqiS9G+ovQ25NCD/KrFM9/8ZKxY4CiZR1ivhkiYPth1WfKm
bNjZgYIVYcPHOFYdJWTxoMZ96aJLRchPolV6D+iqtgzpPUlL4UeJP8ZPDEzgZAG//EGdK2PDCJLn
fXodr4knz1mLBB1/pNuueeZS8Oo/tj23rqZAxhhtDdyQ9t9FId5bXLgY4ptGTaGDd+2HrmxhREtK
ptV2hXWm0j272rShBcVj/ni/QxhF0Iw+nPSnxALf0yCuDaHA4Za9qG4htAlYe0sGZHC9AbdIp5bB
6tug7lniWAv8IVM0evDv9x1t55sYIENhk0RIQKUbOEn3Xbirb9hYNGmwG9xt1YbBamO3gZbumxbc
Mk115fWMn38nGOz1tyQmUuxrIf6hz+gEufhInvaBExn1nDYNkxXYOynzWW9/UiS6fm4j/FoarIoM
hkWfNuQni79vh4jneZsN49//UqKXiyG4iIUpOKc96PRV9bebinq63MPByekR7X4QwgnrwnzJaQrx
t06KeRdxZ25Al6gtryfmjUdqJGBb+T4wIlYSftVDqvrxoKpV/JGEV/4jiCcOtAhm1A+uj3dTymdj
H7tut2ixzqfTl7X4UoDSMiB+NqZDGtWAIX0n58ReroFYNHKhzaGnt7XigWzXHha4bql91QPH66CL
+DyPSwR3BNZqW8EDTGK5l6qel9lX8uUnBMnDiIfQvCDohmVJYv4hafj59ZlBq+ugBriMHyaEbHNR
LV7uziKLhIeKTPaRLWttyHGTJgb+RLZ7NfPdarCVRGHcDCnhtzBiLhHvp/hjrGp6YEN/JESmtDBU
aWu/GHWFj6aSxx8FVeuqhevhFSgrsiYmsxyMBbk6DQ0TgWLkk8O1puYv22hUa7ZXHRpmuOeaYqnn
aPBzewYVfUm3vXOQoV42/UprrkoEpHNnrqrSX3qeq/JE00pI+op8a4LQUPWM+SlUqwiEw3mWBY29
J1b0fY813I+PT3pzko8MtWN8wdItuhqKBDBAiHyNcl3vGWydC/1q0nFrhvfbQAvqP8IRxTHumpoC
abqqi7OOSpyTQ6qwWbI2K+l7CfeorQzu88eKMxH+tX6A0IJ3nkNyp3abVCWVP/eja2sqGkrs4o+7
EDL075jTkypGXiqPLgHh2qpuWBZ63qtRcOwGKKJHlAJraV+ULIi7+UuLxZK4PT2o3VJJDZuj81P/
oOEQdFhJLMZ43d44l0Uyw1MFT2HqEPg0TxfogG5HK0B9GfPdkeSUNTnjROjWy+bdBIO6CbEivJw7
YGVVJFAAVZcOhBH7okNhpamhl+h4s+ymW2S447EXDIAqIaQwfbZvyS7f+vBdz5a4yPt+4xix8IwL
ggbUxH0jFBxsT76L1qOvEsnufjr3L90Bytx9fCfRI4oCNrqwBYJLWHpfNOxq5oADlCxG9xFop1WS
xT7BZJS+JeBzr/NvK0gtujRHlx4R/z/mDKuqY5Ge2KvhzeGMI40tGMftIuqsPnH7W+2qaJMnMZ56
ApifHk+V9XxhtZxUXGo95GDzm/sN9csjbl19Z6leyftsf/U651sJANExa+nb5huzygW71cgQQBWx
e1nRGgrEfJCIajmQ+FnAjTlK9Vpu5OHQ2zySGiRkTGl0AZTrRBjxq7z/IjGsrjK4szGFoWyU4WVH
FBaGwUrWXtLTMoSreO3ZdMjXjTEZ2JpqPRG3brqEVhZWPZCX/UgkFBsA1IlkM50gLtzfB4REl8TT
zcMj58sANRDoX/xrJnDH4+FHHKSXdtOeEXkjO3BJI7BhwG18hZVzTcefkJxza2VSE/YyIS6KI3Zy
YvMdHhaEYfRiyN151yfTEOds2C+dppLo+jHqYCsqB8Ayo4dBfTNMKG65Dw1TwnB8ZeNFFQLAEuq3
kLnkkTCoLu+Mh/mvZ+2FVZwR45I2p9ve1Blk8t8AIdukXpyGydLo7gfK9v2smYoeoC8aozZqXIzO
WmBSy/Fcspz7lvu9JcU2uKWoKZ/DZ90Ry3g8Wc8n8jrZVA+jXybRDvvB4D8vw0+nmNuw4RBOOHbr
zny3oPf0i8JYUzrxx08n48y7IlOE5YzcW8IP64SgUv3amcoJiD76MtLMIs4wErgJQ5aRdOFsMRXO
5kfoXk4tHKasIWqChXjt0GfzCc5kvRbdl0L8HtnfsXKm73dzhC02TG3slxNRj7v7uQXZFWbEC+nL
IRHK9yeNkPMpVoQUaY9v72bzKliTV/J1UdQ4+4HP8V6M0Qns9MEiZZE7XELBFcgDKNDH8hoUKp98
dY9vvnFIRolA6HQlRSaJxL4zL/wci9coKU6eQXhTzoKZE2OOlSJut8zkS1AQUz16LWLklhvX2KXe
ZlCXZFXh+qziLGXAehgudwQY3en7bFKS4czDNpv+uhYnIhXZqGKIw+q3EH/Bij1tUgUTPkcOcpfs
XE3Ehw/G7bdujk4dKVtscRI6uKvlOPkBOUreIu07AFU1F9VPd0RFGJE2NpR0TSHOymqdiWndKojE
Jz8aIpqrCfvo/t1Uea0e+JGpTBKBBwV6vp59TRHCVLQIbkwjvbqSdg0PhxUyh2T2QKpmBwcTwnZW
0ijIZsn7ts9StKU3X5NRc+k7wmPJIhOMgXG0CNDSa7cBQi1wqJDLf3D8uB1T3RtV5Us91zwy3BJs
Z7fMHBSO/bn1Vl8VOV95bePbzEQON8GOtys2PknGhY70EnK8TGfmO6XAI90mdVaIx1Svza6AvuIT
mo1/+E0CGNjxDvM2EQ5ioeBACmR7tfLmawbNWdArQo+0psL3Pmm7O8Reqxio3BMybANsxKWm+hFC
ZHEeWTxsFOHzAOdfhGtf4Z5JT+mJfXIrce4u42JJ92n+TWYH3dM7xmNRLfq2SQEV03XiGA2g1SVf
z1onKonKSKyJkoyi72/fGGhSh5laeAMlrAzMNwTOLCB2TY2QXrKjMM5O8poY3mfvZBn5WCu/hKs9
h8gN4hiYFxXfFwr6Lu4WmU2LtGlKhcAbsOOn0yOpVaXW12pBairRQX+MmETlAM9BaB/91M1wwGZn
o8U8X573lmSClfxaa/78eckAJ+dUjs8vF0StK9lEwyAQwzgPdUqChFRP08fPPXjwdsb2b4Wn+lqZ
LbrRyJ7AxdptWwnudhLlyrvgB5oFvlIEjw7hkWAw0hlwE0eBgcKtL9haMmqAebCU3Rb5PZITl8o4
NMu5tWL9mCbhX+8i2hb5F6Do18wjsFZ/vRAj78v5RDli3Jh9ABpQG1H5p9sd9enBq9zIIYvuVoGE
/bfx0KPFxGYQ2HlZM8y1GJb8TD6lzh61IF3KG9HoGUer46At0Cig9sk/7ApALFLL0YFMia+Ee7pJ
0AgN034ciakbaQoVPNeerPOnN52ew67jGawIfwduLfFgG5VDBBgRgu8+5TQIE6qVm74ODZt7Yen9
4/mP6UeCJnDdDfcXIj1urg+WLWLv54G0+boNnSfEZ9fPhIqB1e9FSEipNmNTyJZrDo2Zmxi+u4z4
sGru6dv0wjdhJJUsGpyjlDekAAKKeZ6VEVcMM/8oqwe+/vYW1EjyfjqmViC2GU7t0Z6UjgJkH0r3
6HGaDP3oSkmPAtKesYMSikbgQtlbhA0GI3l0zJz71IDZ9m4d3I3Zh2avVOVco2yYAIRwMJvddCJF
hDMUxSfZR3z/9KbhcExNG6ykoIaDXIW1wbMGeFxMNSbeIhjr5cUkB5hEWcogKTLKJxupkQ+Wg0h1
siGEKeOg9+b/JEJRWzerOl2+e0V01Puu6dpG0eS+Psuz629dJTvjybLUrrLsX8nBDqeJ8dASaYY7
eFnD/go45vdTpThD6Wjmi3gsfsSOoHphULsF5tkY2EEB/rmj5uehcUiI/L9amaG8Jq0YzKOwk2AM
4rFhcqH4pPc0OuM2ljE2JFz9l6U21TRxrWaxA2a4vMTGWaebJS43Q8TrxtAnIbHmRMdnOwSNzC0M
xP4x5e/v6Ae8T7RnMXJb/8Yr5susI37NPxhAboJyXmVCAk2B243iOdFIpvAN/1hqkQj418vdw20p
nQpaB6iv4cmukJzyHeEjkzsq1bwHM+hmvNvh+TaWNqKhPbme+cwGKzvztpVcEFI+NIKpIto84jj7
QZLkdpSLeP9P+dAv8mcsik0YHijWwsXRblYd2Q2ckK/wvAk3z5DJ7fx8aBHKNaKsD5CmBsEK4AXl
hnfcJEQO4/V3GOqSiCvQlTvY/tq6tbSu3zNPHOHnCOs7FSTDOhs02AY//y6gMxUosm4vLR65Qzvm
rZlsaj0/029vZG/EL9AMA1c44UijLKV5/W4x6YZrBgtcG7UivOE5/3Ud8r1j6Uf7zL0jsLRcoC8r
zBE30qR+xtXVY9SIbkBg5xPkcP/2N+aWH+/CheKtW8wfut3npEdl3S3bx4JncNtwtbbZSdMBLkKH
1BDFQ225hnUcQ9sRxRbngALIKNevsrjpsF5PYYPr+c2VKsVn7V/altYqyWs20fxUx70a/t85oezg
O5nCQ0amgRBAx8ccT8th82v92HyAd/8NgqUsEySybBXxIGUHyKIffU/of4xN0+OOZ6Hyevjbcoe7
O1mScIvUU2fZCfWfeYvUh5o6pTS2Mpw3z0xlh5BgedWjm/hL8fMWTDdWDDb0RHrKrysQG57sQvJQ
l3etMdz263m/F/743Fvr1eQI/KTMSQFmTZoOa5EdBZ5VQSAwZMtnQOEwIzVncm6f3JpWTv3qDuit
D+RFNP1So9jz3IwPRo27HyIxg1yFYunrvHdHRt7PoCt0PPgaA8CA1wmYtHnj1gX92mhsYh6sd05g
0dF9Kj6sesUOSHeAjv+n7v6VNunRPywcmxR+FYYrnSQkMlucHsUzgSbNCg9RPtQ+D2r29eZytGj4
907s70ryi1cg0bvafDJJt+qd/0WWINVVb0Ve/fpFzMepoP0QJiskx679xbKtKxYzV1XJkmYxTMPO
g0zBeKm9+SslOcyhgyR2Y2VPYFP4nYDh5b4isHryaOJQcHJvm2xcBPBTtB3MNOTrvXNspS9OlArN
gcWMS/0a8RgEW1JyNZQounFbehkIWE09oEPyF0//FcnzLl4Lq64Gh9PwGQa/0/5QVvXv5bfgzqhQ
bNXqqe80Sh0yQMQMD6yPsfklKvoeVm+n5R3ZHawI7kVctY7ez7KTyL4Kpb/B6YCrxJ2VW1iZb2RB
sjleTuafPHoPYk3L10/UyodK3GHxDgr2i3tqNysw/qsFEv//VlLm+Mj/erzV0BGoBZhDkZgfuTbM
AofOezifLrN6fwD7MNlEIudzNitwSQLLYl9HzSRj6+do+YI32aOBQrpusjMzenxzOk1aX7kA+pok
P6my4XuOtc5+c/Z25nojxduFGfpm+XNpE63AE2wSt/CcJZvxwY6OMUQ7hSF4WZoR1m86t38NT/1m
dNy/4Y8S2eI9VOor11roNvLYFS1+PnhZxx+BQ/VhGmAas0E4qHr+JCHPIiw8RixaqPvSH/9fC/Rj
lhxVljxb7odIML1XCX1PAXtTKYfkE+k6LI+x54srGzJuhs3rTcsE/JYqPoRgf5Lxp9XXJbwwzB4X
aFiWBzQUUM6fpVs72JUV7lpIrSeJqpAOolX0dlBolqnwyC/kp92Xawe+I3WOB6TI9rJ4lz1eFeey
5TDAxT55XboXny512vQtWUBePk/RZxStLG2tUZne5PV7JjSdU35NX5UGFtLJBaSObTgrXVytcAeo
6OWiwDYiCh3Qky2uG933W+DyrCqMj2ipPY6KfUiKtN/cCri1Vr/zBynUEuV6UWwUS9+aWYPqCfgU
p9XNiJ0jFply242JahjZLRbbxoHCBgYncyLrwOqhq7uiJnUqA4+Te3HtcUGqpJm3Qqp5CZr73gJv
yzNslpjWISqufMhew9knNPtNORWEp1bFYOi5TW8IYkUwxrAyYnDxcLJiiewK00kQ558IsNBLr+Iu
vVhzwb80+ipAAbBLUlemuZyiGpSUSIre5MSvFzJXGijU86qcsUJUbV8lru/LpSQO+xuTC8CQFqPm
3mvmyJi0l+hob9uItuML/Sdig6YyVoyLW53+aHLh5aA3LoqlXj/jOVw3MDaPyVqQPEAFy4QwRep+
2lwAHgtznNgNSERt+3vfOK9ktz4XQJBOiGXSuxXIQwNaEBci/TB8U5WjL2BnOE1F0BZRKVeYnmk0
jVs9gTPA8nnI6h9HnuOWX6nxCbhcaA9ikwv/o8YajIHX0/kK7bj9iGBZ/kKy6VM7AJCk35GKJWfY
p53p2T+5PBtgRfctuu/D1AwkxXmjH/fKR4k99CCK3dAjEm4JkzKAZwBwCe3LRZf1MeXnrK0zuyND
sjTawYeI8CZm+Y89GUU1gHw4MzHI4TLEVEbrpstHvK2+IIchbqF2uJI5uwbYzrlWzZGMm0jpUEkb
WbloHcpyznL+zq9y7yKBdzxaYoQ/JReWFh9vyV6NfmBT3UiCM9mfv/veuhN5LOC4OT3ta++GhMpo
DMXYXbttBDqAQjjAe0qLqhx9amUhjGtwzVpNXrJBlgeZW4dTAjzDxQRirsIbfwxi/Tq4PwrPRnks
tV/u9XTAFPqjQixeIn43dvvMlN4L4TYGVa2hP8+TYvXOZTQsDmW/2yvAz+3hKJIgker72QgPUpxM
IRgoM3QI98zdLT0ieRsd3q0dXkr5h68m2ufGDS6WGWEubn4ISh7nkCdRA43bjsZguVKp5yajfMf1
A6595vT9/Xpw4Exq+KBsHNnyuchKHAKOGs1GZKQ55W5CyPt0T165BvhIajEp3tKSFQFTsGUy6er+
fGwxsmDiDc6pMFHOI/GLabt+B6VDLvBRiv6NVjVOqmeyf5CfPVVkwsDodCigt6duSeSjCdNobQSc
p5LDt2esFOHBI6g152vw1HZ+/Bw7BO+iXR1Wi3RisgrJZT4I2wQAt6JmbW2C8n9jt9PAafU5WYyR
cL2aes1lgVjhFGV4Ow7rD5nlkAL5mT6OTFT/IzXUcF3jr8uUarCIIe2XmujczA24Du7oQkDaYSp0
jpKXYpva13+dXqoJT8A5Lva35mvzy6l6giShcrUQjwbV8OeEUecvOBxt/dZ0mdR7WsuxmIT73MLM
t5do6GDHX8vrrwpiut/ikfqL4xiOv9yqiuuitb6hU/bf2VxS6cQH+4VqZKMMyudKSmeiSKGDc19t
vl4y90gY94eSOYtHvhjJfpX4JkHIaaHnGdxx+fn+LPW4l38sA+NRIeWZzxGXSsMvYHJd0VFuZD/e
IYWLmQSmrojWI5D27/iHWndw+M6sCIXyr6/1m+nxDwb+QkGmGA8sVhP8V1aa2F2wBtHSZ7Io88l3
YW4FZURTA5hPNQxM61xlugU+vNy14WxFkUwwXiMYHH9VB5vtmD1VTSLP9mw6OgUxE/NrhCKgKajf
G9tKH3nhUgVD0N+nUvryWbmFWymHmvihgNQxddOpu3czLoz4S7TtMoFqxzMt84d7ho08W2F53C9S
Bd2vj+pO1v6Dy8n0i7GTaxNl1kMgZX86TVEtFvpeB0ZTId1UMCDutB+CHcjRoWlOUP2Ijkz9DVwC
ksegvwU63CWXFXSlm/0oOwDNWhcK/9xEOunUDgag8KYgxSsRrFY4cBLq4xt1hHbK+VX+bVQMesyt
9d7WD2CXwXbFsWbbN823irsD5PNA3VJmWUoeuKqGapICZHZWpESswlwmihVAw+8FGJQJJKWjyyw3
gTUa/JNYFh/0xF3lJX9XJCvEb4+4WstFxaUi4I7oGfWWGnyme5pmv8dm2jweYEcbmwmRxSj9nieI
konPL+ciybvzvOhmhc/3i01nEkmVwkmVl7/ddzwlSSbtJYb3xoYODNm3Yy+itvyzSvAzYtsXXjhj
sWV0S4p4Exz/0H14uThCFf6mBom5jXUHSW9dx0okY/F96Cy2LXrIKJau2J3yJuT69KKZA9xPBbMR
l47mdgzpMusTNG7fY0hoYnyp2FOFC5hNNmhJyWLuiKC4rmED7iSeD2aN87iMSH8xaILRUjv+vBEF
AKynTkCbkd0lo0jQbNgmT3qZ0T64OXk+e5FWe1hNbYytzRumeFzI2QAqa2deIESGgGxuQgLb3bAM
L7/Czvp+cSBvMFb//DQPAMLd0ulFOSOLGIBRGXqOYavtc2BDrwiTMkdV+Bz/yW12GIr0/TNUdCzo
ZrW/qoIFG5G4qz0BpjHRMygoDKLcQqNE4Ire9J4Rrp70+MfdwniUayCyoZRxfDsMehHum/hQLzjh
wWRVTwxD++ht9bLlCdThvtZb4GdhZsBbSD2p++dU2yqQlrIvZ5ivDg9yEhFbu8ibx+VsWY625ZvX
jSU9P2iO1SC4lKKxge0EJr/0ExOH+Pjei/RKO+yVthB/Fwd+W9wgum+iHQHYW8p749uwwyhWwrp/
Vo2j/gbgcyKWQHJ9doh57yD1/NJMaMTx8p0e1P/kcCEI/qTtXabpwzS4Zo04SPCyM//ZasS32UCi
/9QKzoz/Gal90qViVDLcyhyoO+kyTA2T+UEpTtTJ0LvmRUEpB2r67+agxFllj+EMxtamSfE+dSnn
DobXRdeRn6QONB7DG1gKxCJ7IgQy4PlUeOBm73CMXA2ninh1CQziXS87JimKXzs+E3Ian9guN7DQ
bbLVUfwknVaT9P1ogKv4d2ptU9CBBaSZW6MdrmLsKea+LSRfQVRQNUSIxHI2lEum9xWhDWRCW4Ds
9AHT0jCHpVsUvsW0ZJEt991kJwWqe9Moj0mXgGvfqe+iFiCBoWBrTZ91vvr8B9SEyRgdvnfpDDBS
zPSjkHr96EcHibQKqwB4BY7kc85fxDgBK9QvcZaEkV5MazJK6XIJwAKdJCDuTgrNsN5ho83WxdPr
OdXRUglz5TPjB/UN2brUJZLb+vPOEcMjOWnldTVo2/53604JELus9XR/IrohJO5NMSdSMzD/LKM7
9slw/Bqb9ooh48W3hBXx6MhzDNss6/FURJr06vGhJ208+323gqoJBoKkpUFo3GqXOTAjKz63S7Y8
DV4WV/aV5P2PoTVZRrq0DDPbd8BY7rMwSLdUUH7kaju0s5SNfrPWmQ31OmDGKI+68eqRaw/N4bRH
tVEXyymANHGsMPChHN6n314LMhDuP7ViZkIpaE9sv/mvVVT7V/25aZ+iwAXaxeClRdNVfVFvpt9c
39p8lj5IFAOfujNNXTsGT4YfUFCpDOJ1s2h1Gfk/+khjXjPJvtNnhwg926zmp3Y03eM/hbaxeEtm
1J3eUJ/LXRX3iSf84k18FAemnR5TmosSQsH82b5o++U299yJgRNhjU6whxmWAnczZPAkxkXYoiFs
47fcpiA8ukeHdEVy2fFu4kyA/Tz6PPwVFqGD3C+eFxnNvyE9G1bsp4edvKisXNf2qirB/UdmY07f
4z8on6a4Zi6tW8jE/qtkS1SPsvRgjoBDX45nzbtKHKUWFyKXJWSOUj7DqmK4DXPHMlkh8Y/rhjvI
gGYg6V3d37IWTMmiNjeeNx7YNxngnk8+ZgO12I8DhksJ0pdzT4uZUvYfQP/MpPcaR4Lig9KMlq13
6oiUQ9pe04pbeZVhrneQPG8PRvuGv6dQm7Gq0wtI9zj05qgHShLbZ85ZSOusSMpsdDAsiHDgkMEC
nv6urrEHGGBegkGo7vITaYzihhi5u9iCzTAgbwS+NkY9P/FN9y/KQGmHmZhHFMImTLKTeP8KWCyb
yWKMAHhdQw5SZDoQdOaF0USG/C0b2pFbXjVgPNuXJbNdlka+ii3WT0uLyW6xqqoemr0oSM3iSWVG
iCO0EUSvlDw75d1H/zZ+1O8k8xx5v7pIOg9gldW/uqRkfxCvhXoaMSHLPnt8JQzw4Z08dctCvZMP
OnX6mEQ4hk/kX0/M5pCxxLhnzyv9VdIlLh/EHUspi8CdVrytuYGkwMvcBskF8+uwtHeuzs11Ed7m
sj3wLa0/6r6W4HiyomniqdYZeX2Fe4Tcr3m3NpWDRUKv9B6awFPMS8vfXrZ/dUwAztL31y0HcAIH
s8phCK6HfT+0Hm1Jsd7AJ1RebiPpaOa7VwgnYzFKRVXdFxX0wKhiOECq9QU71fqIUfJ3z7R4FGbf
/kBFCkzf20nSOxx8kaxf1Irq5FS2lR6eLY4vZGSXsbZ3lkKOwdHFIbj4dUt9CdL5XIexSpigb5aJ
8ty26M3QuPlY8uOP3kUKaDQpqqbNo2mEe6EWKSAYLmkw/R6NUbK6KSa2aVBJYuIZAT3cM4CIEWs1
9KsV7hiiQ661YkTf9rEaLf+rWtiQuvhXqqI9y+tBHPUBXvvPsTPbdCZ1vBP9gvsbiARPKcN/vdi7
A/FLsepeAnQfVE+mfp1GEgGBB1lWic9WuGr7DLJqOQlj6Rqu6Gm0evSZA7poOxuHN8UCjEcRQw7F
N9ui9+uhqEs+p2lKiCOqDYQjuHkpuEXJDutqOjrpIba7BqBZCJySmvc/kxCydOn/dQfU1CfrKAeX
Yl638hCCrdMfx+WzThkwxynjtIbJxSrBKefpmlbryj4398ats0h+pAM2AsTtZD5hW0k39iEKR9w+
N5cJMu3BE71Q63VgYyLcS3doRPhpgR85kMT9djzaOKeENcNuo8lPe9kal7rt8q65E5mlnj3PDgxf
ycPSQB2XDRpl6jvytrAhWSxeOQO4OgR1ikKXq5b1SAh/Mw3P64yf6ZX4FbtjSkedxrbFtF9fJSFB
/XUQrMRTYCwlHL4TBR48j888Io/8tM9GHNxdzr6HUhvnttY9T1YmbkVRl6O000JdOOqcYgaJbdng
MjWHUCMSaJ0Hor2mM/44+/yogeKT1c5L6BhohuZRtcuPQLXT4BQ8yJFYK5Vza+blPs8HXC9Hbhx6
RwIu5c8pXqdwl5x1jecAXBGeLfKVq8jKVDccAFhrQyWbqSmwve+5ZpBKYGdr3LzLS9qanZ9FmSKX
ThAtkwmnnouW9lKtv4XNdcWjIhtAkwkqa8HI2ZxtL9tjtqBeZ2tsz/xS5D5TPYuMBjltW4vjwwon
9MCzQM9YvPmza/rADjZ2jajEaVAd3s9N/g7eiuofNsowRWgDRwobH8qivtGbXG9/ukVibrifz7tc
gyWDMwAvskgsXKoT+jb6zBvZMa1bS8tu6ddzHbwETroC/K0l5Dd/wJtX061PdszZu6ckh4PjsJc3
Jrk0IGENe+i4AYAt1/AE//DddV66nNPDdezU5hF6VJpQlHbIuarsjiFDRD6G7n+/0EHatASEkYRx
nyN+PzNm6iOo4GMt3ZHszROXkgfSWLJkMIz/3sb21qjXBzgGwbMMlXI8692F9U8JoYEKMCpZh9jF
6wmUxq3aL4veY9yP+AhcVS2Le2zFHy9QQZkVayc0eGu+ik26jFKrUDmnvR5WSnpu7rnOP8afnx0V
a0bsN05xQgovsFmkpFc4hdLLJ0hXIL7hlWHXM89nwpmrX+VuJqfevgy79pfiuUPBUEGtpu+kgDUA
+cqjMEPjPDsGh9KBn6zC9lxxA2XpBwxghY59oEXJQo38BH1k82pwdry3cSl1IjFCz40g+qFFTnmW
Pn4Wz/lpuc3fSpXJZTHepw1d7qp0LqX5Tn5XAgwl8MNfSNKoJj4cq9XCG2V8EcZADr23DDM91b8t
13Sdw3Vq9inSDmfS/VkVvz0YgHj8RDpfy1RcaxV7ETJ6vB+GLU05G5B/9i3aiwUfLiA/uU4JpFdp
qkDf9DuF1m3cvyF9b/qu+NgYfI4QRPnMXk8bf0BO17Ez2IYDoZuPiGlFcin2BTArtXCJ9DLljrkH
A95e9xpZas8vRd+KBf4SaJrUuVbFSEA5H2Cfj5rTrG3oaztrVOX5aFA+sOO5b37GN1b4BAa40hMB
9s/c0TFHwY+fo7kPJrMKiXX9MxnmhYbFQkz7f6vGASn03yQeU29x5qZ+hC90dOGKWc8DG67uM/HE
b8XAwdH7SrBRc2WoHIFiso057vMGi3ACS4dLh9Dwd07c39XDr+jEffCiFg+hU1W3d21SnQGFk6I0
pG8qtV8aslH5VOwb32vDRZQ9n8vC4xrzAVFzkHRc2rjQDh0fP64KgPceI7DW3uDE9W2kAnRu/T+5
vzKhSlMGJURSk6+yjlDVH/mIIO9O12WJeAujQVsbu2QdxsVtqP0E5w4xnTObe8oSfuEBwFQ9omIA
8zDhFjZViMD1mTV86UNwYqOjUMKMY/Vd3weR0RvYzTu94q2D77We0sN9ghFbSErv4OaUuJn5a1D6
gJ4g+79ICtUhDGPD53HFdFd6FKLQanm7EABH0AEXHRXYpCyExxiHfe9WJQk1qC84qj373oFE5kdW
d7yH06VhPe4EYtLHERfThV9wKnAp+wrhrPAhSSmx4IcgI+A3ZBq75MSqa5axylgSQDdPPW06Vs1u
nZpAlarpBNnHw8x1v2xZ13sRFj1JyhGBEvZ3B5KFTWtHuU/AVslkctIxPhtFnns66E8mW26DAUXQ
3Ty58kpNzBgTLVLz/2KEkRRTMHkHhtDfiZWBtcDO1He1AgFyCjzwO1KP/bZlicnpdtDDExqE9u2n
rI5UiMkiXqro/U+HTN5gN/Y6mo4x187KBMynsNQmqhYKgukod67Hfqh2pfTUqBzPyfP7kEbr95JI
MJcaV99kqXBXX4mEu9rP7KVZe8HQ99DXT4ISKIcOD5FZciQpfehaC3kxPNKioDf0mgnaGzdB8Og5
wIPLbB0sLY0iRuJ6nhP82Ekq46lBhhNn4IWfQz050UtIQS67ASwFOrfIrkur9ka/q6xrpyJlxa3B
ddroyaTW0VokdcEH8geLxErfgFK24dlmqtgeroDSHXktvBunmXQ1tbSTYYFKk2ku1/wgE9h7g5YQ
zQI0mHjiMrXrpsZqkwfaEhePmBZt90LBNyw2A2i6gWQrm742zRso0WgHpu6e6R74zjbNFwOqGnmL
p2cunbNFA8QwHe+Vl8z6H1uoeNJqA09ZTGfUJeIXtAQtUfCLFJ+x7bmz6kyax66TF2f1nS6AMJ7e
qDxh+hVCQg0g8jGxf39zbuU3K8M0mlUwxZVd4XHDbjvsMg11TLvuJzQTz3mVKMaRYoY1VLHiLcZG
T3Qa/EkvcgfFKdZqAOofNQ+2FmbHEYhQGmC7cuTmHlmZdRRhMgwlpUn7DD5RtNCnxUM7QBHRqjel
3pCBgHityDEgurf5QZdduCiljaB5FhTdN6qwcFhOA0EjsLjMq04hX/L6wjGPTMQmK9X1OvBmGmyp
R0p1Dl9lEEfWgoZEFQZ6/RuAzB5bI3C8rBEgN5rstPDHGVDsiBSP2We8zCITucMc97Dz3Kld7Srw
NuV652iz3PHDTSdq6J/RdtiT/M9m1jDnVXdTemtvbMhqNtHSk/YwchchwRlHFNpEOjpkKcCtE2+1
bEAJyEKkeqSw32A8hMDHbvPyp7tPKK5MZggu1/lRsPTD8zzrC/4jadDwXeqtqLBDtb8+0XnIvwcZ
5nMNx0HM09NFAJc+2OJD6B4pGo/IJYEIX9sBdtGDv6o6Y0QrBgJJqDoibbPzftGcvkt6+tnndqyi
a04ijLQ8MrrEdxKIWiA/we2Bd0xE9LOh+wrsQ8A4zSaFy04Ig8OWJ10FIctH3vWROfa1j6rzz/r8
B8syeGLWfhRWPNo0LsGCwk8d6IttDv3Tr3bkFimukEY23EtwPbsdoC5VZ1cFM7SId/BcTpofd7a8
EXH9JqbezVF9C4k90BSjpXUtLSooEBYPq0Rj5J6M7hq/JERUl/hEXT8ALP8Wo9bH9NbxL2ddX5+R
gcYkQ8Pwqbf1HogAUpbldCK6uyhlHSRxO8hJA1IVNsk3axJobjgc4VyHESQLalhWZ7zAC/6Iqtzo
5jMxUwfbTKDWptWJVk0B7OaKk5p4TqUpmQJoasKHsRfvJkiLQ/Jpe760AdoyLt1vh3l1xIIxhNEF
9X3qkmgOVvx6Lo/kcG+n7RHfvclQpYLFgmCpyrMEyXzX/EuYCXBsSWSmckcwa7d0rIsQ5z5ZGTpm
5zuvR2Lm7w3o8BVPYdZ1t7xb01xKVonuZ+Y4yi/dr3mqKF40GwpkCrZxnkgq/e4zh/RPAuLrV2/u
snql4je4+s6444+tAAjnXdZX6ISJqBj/Ocn6IvK28VdCZaKYdB6Q9iBhQQmceoG336Ao5ZHXXZW2
5WdsummhImO4OFNezmNCK7eua0bJUPgYWeeXxT+arkFXu/BM8/25EImLOyfrWQe4ki6jUAFECkS2
pzgv96N/5pxBt6f7mFPkecu6uLX0n/YfEKi3DEbFjjt7PI1pYIcC/gUZxqW6N7opm7QDwkjZG4uR
ghv6XkJ1PA+OhwGeXBGWsP79qe7itiRSfnMWBfgD9hg5/PlI/b5sLksoXJgqy/rg7xURcZmG1iaP
oz40JDMV0Dw9E5IHrGINhAUxi2KtyYg4R8xgv4N6lofd4P+2mdgo5vPzUKni6xfizD5yIZ4aggRc
Ua6pQakdayEvIeTqoGk1p2sWhPntMb9DONe6MAWJeqHzHonJ32bbd0Ul74qer8MHvFhrv9snCnyf
r4U+culq9ZXo1VfmqQn89sACz4NfGk8SSN++E1AxRSN9P6FnVZoPN4gw3miGqYARjp5MY+C/ijjg
5HA8J6jXpXkdyz+E5t7NqKVCusk00YJP2FsjgeAneCqo/PA7ELBlYm9r55JQ47oS2ydnpFwhtdKU
GzC5A2Tx+1I+xxf+Q2ctFYLP7hEdWEQs9jGhEgrhvXhziVDR/k8miZM4J5fagg17I5uTaadvNjM9
n+z66Nn/cgsOq6nYR54lYhK+EkkVL86UpKSMxD47bNtBAdeBgYVlHvd2VlL6l3gmu7UUr8NN9lMY
KMdjKGTxax4JtYm+7XbUZb9H8AJEn2k2Gyaw8DPxkI7GX1PNSfGaZF706bAWUim2ezALLydHTvHR
YSDkPem7uXI4ORVpzG3M5DNY55jmZjwPmHmaD4CVFtXw9S48d6gO6hgtR2kLzBDh26+nNWKzEJcK
ccDFcljSEExaTNQjU2YqsbBdu/he6DJcbkfTRebRgYxmQm6Ykbcwsrgy0Lb1Rv75OevbI/XKCuyu
vMyERABcfC0k0w72w7VPwGFxxRxNQeqRFcSQzzs+mEDrH2ia2JFunaQKwmXdKqDx6M8xcElUhjjg
WQFvM2EI/uoqDuHD4SGjLyVKyz85YB3SfAJQRUMMUjYO9UQlYAY5tKXHoNuoOQc/rW0oTkcyixOC
9EQz4FNxSvfZ86DoxoYNF1BKVTSi/82ofoF/lMFs+XQTiRyt41NA2f7gTKeZnCH06BwvLlhzsJAm
ICkx3V4RhPFeIpO1LjWBbyZx5YxWPQRLxIPAa3shoOMr3fh6RUV/kyuqZF05NTfI7Ghjih6+ucyF
8k3qQbArHV+mgyl8Y9nvNhEnYSxvBZc9/yr75jex/MtR/J13LKGB+NOr2VSPmq89hHu+kSQKb8ym
qff5K254SR00vBxr196DbXOeeX+AysODBFisvjFnhjQOJ1+WLrYyIt/nplr4DTuEK+uoSRQawGMS
vL55+etYF3FT40yomOlSQIJOU5OjPvkcuFdvdz5ngnN2wtfFrAJAqMvUGcEuWJPXmDmuHd98QHVL
MgRRU7OuQbZJRSqeHGsQEWofEc/JvzoCDdQ1HTK55Rw0MhMxeGod5iwYdYI8rmhYWJs6hcAN2BNr
WucXCqIhoH94Io27KIlEf2sWhbWPfBxbQvqNKXv653PSnPiJ+A3FveEZKvi4OHfTu/COU5JXv/nC
NeprjCupY+81jVd6JIjyjSXcTulUVKIz+FaOKr4RyOKGJjHKD2Oezc+vHWG4ro9qAcJh/oo9Y6Vi
awjt39qgnrMeT3DqoVYNH/KZU+jiEGnzFZlJ23a68DwVf3pSPwKnB5oTi8Pzhizqm8KPaY2Fne6X
aRK1aFCyBaMOZA3dtCy8GF6MyGOJRUfI+N9Qgj8DvMjYnMgp4bTlt5CW7/voSyk4ENzXDve/x+2L
X0C5SlgxJgYl1kvjToZxosTU8+47x2ogMMQvn6qaJ/aLnFRXDDwiEOW+G0ebPA+3N9fAj3DoV6JH
TncXZNfzJMOY7hsAtxHaAyzAgAFwqjfz+oMx084GX4MhVZ4AHO8P2uIObktLCykKMnGvfEVlXDPd
Ag4A14INdB/MzQl90h447s3NFTIqwHSawXtHdnaoUglkgtF0AnV6f0oZqdOIIJVBXoJoH+Y7c54q
TM4yoGkZIFeyZ/jLUXt/HNIwkIYjVfFME/aFmnrMkZUCIvIW3ko44ZXd395NyQ8A0JhQzq5vcd2W
/UU6VFlokk0eW7uQfpQr0Jo66+l2plAo4CARGNJiwbMTza/SMlfckfTUCxeKndk+b9kJGD3lYZuf
d6lu0udUwjXI0GlS7erozxknMPj7Wg3rejoI+4den9aX0dUcvHLiECXswrcpE7acbJfxx7CRB91L
j+IHVm2pK3mW0T8XY72JFWZVRzFLiy3W8PrBD82DA39yEVjxJsb2P0pzAob19cZhLwLe/FrDZHOa
bhnPJNs5dyT0Ic+NMDyp8ykX17wCZxwCT+oWBGTMvhMLEZojZ1pS7wpvKveJddTMe0Maursxz6UN
+fqXmKKjPCIZ5fEt1nf739ufTUKgL3cM7l0eYqJrrhtP6JTjlKy/yXvFT02KMAlqJeWnllXTwxFs
p8zhEETHD1PG9b8dxjZYrhNAGoL+3Td4hJrFH070YisVtkBBr7LsqTxexFrpaRdhnQoiRrivKxfi
Bk17j76KRP+V9U0DOpCLOb+b3ZO6X+9s3kPOcojD+6CJY4ZMO7brwYQTMx3lHyL3uoo4zHVy13md
248GWfWD3EstocHnEnokYx4ub4ZLwlHSrvk+6nflCRinzuwC/s5sBUkbXyMnQG7k0zHwhNfTFy80
oKE3kWgvVOjjxztiIQLsPJ41RDpVH5x3w0MCGE3jfPzxbmPha747Ea9lHEXs2nscPgCP20+tUGck
sUkcQMnyOtDAnB10vXrbQkEElxYCL4WAd85txHokYDs0o3p20sPEgLYCSgYgKvi+iLpJIjOrGUYM
KmC8pIaTp7go+HeEuJRECtkT6949wOIotr0/Cuivmg4QLDRgWWjisvPQvbb1H5kh8Ibg1Jk+dZ5f
k8Kr9H8bnNqBlkV5lom+l8DdKclg1Qo4ARvy43k4uYAU+XavFLsMTt2BXHJCVp7sxfRe4l74hsdJ
v3vNRGuax9VpkwkIdlEzQgvMuVS3ANLap7xFjzyAX4vznoDJRG7MSOTyE6NIysduRV5QUk/NEeF0
GtSj6nnqrSyDWFBHgD7ZGIjflcb1iknBFviVH0usklBu6nZTdJsYyqntL1lesD7qwHCGodBQip1R
gSpkyf8jNe6jIW0WAeaqduB0gLa+G/gjLZseEUZvDUMOU9KTbZ7vfZ1nLWqwzNaDZHPZb5TgM8Pu
1u8q/VmHOGfjlNMvpM3Qm0B7MtCAuucF4pu0gmMA5s8aqseT/BcubEONTKXbh34AQlh3yfZqXLma
chBehtOWFnbtemsT3uh3pvi+omTLUnAOdMsi/2YYmK046bDxs9EijMqfRqWsJ8zNCaYWSsFNCgwp
KbFpLjB1vxPd0M5pbS487njAQPEjJmzXAd7IjeZuo8RWDfgiwPD/vZP/wfwlyy1MHDKG3jqzs1zs
EJ8w5LnPogKlAKc7SEZ5rr3Z9uQXqHRyCw7ZYfAbgnX5p3tB0dh9244UnUpl7q4OArZWYsAHg6q9
vRP+RTwOD7PtIU0/Ei0Jym+sgslhh8GK5Wghi5XN/NkvtI1ZaIIIpV3GWTXvdICqSmzdDir9FviH
yr4U4+z1Ol+ZVQj6Fz5gj+ZGPGgrvOPUiZv/+rJLctvXtPTK/UPmjDH4apnv2UstNoyqrLnePVpO
u+SBcKV88Kwbf9CX1VsbHDAtuWLXPLavUGxciig30UG4xADjZ227VSsoKQkvRoGNNaHRiFA5rN9t
J8KieKckukEMs4JPWMV/en9iU4v+F5GP1d6dfFrPV1kp6lowl3mGLFipsGg6qxJqlyJnrzHSF2BW
oL5sougHO+fIBUkPt0GkZyEjf/mDeLVqcdP7vG+bVuRqRGdm8ePQqTerYyTxwPDo3q+ak2Er19N5
+aiJ8Fo9dQP7WAcrSp539DPQV5eqS1tGe40NpzM0uf6b+DCulcYcN+1KQXMsTbRRhbUawrRFr0Bm
EFuOUKmEIbGw6BSPVwJIDsyOt/r54bVMO6TCCIWuZlytjWeBD41LAPuEvBleG8rV1c5gDk38fnSK
y9HVv8WLARt196elLdv3yFtctG1q6uCT1EAEck1df5AKfdDauQc5dLprBiZuLNMqpjkKCRX3qk+g
lSk4xalVIv6e7hg/C5jmfnlPidNA6ffHGfsL3Xeher9WwQTsYapjiODtPsEPzy5NbonSYjn9gUo/
eFq63tcEjqqSFd5cv4D5eyvfYHheV2/Fmy+NxFv2ZiRZeMz0mr2rpxHITJlLw93i764q5cAYFRDy
81iJ0qFVLbQeGDWGwaKZHMMASBQYNlCaI+dMXYXHw4aaoSs31DTRCdnyzOJMGrGmr6buLCepCAzD
8kNcGKcFaH+a1MwE1xYVTW8fk7EA0MUHSKra1rq6zmbCQmgCgM99SRW3ov3ET7pOW5SvIbd3e4zQ
j1qSin39K+i5f1Yrp+2ovwqQm5p8BYSLWAIucMI/am7zvs7HUS+rUYInHaZc19/Yga4sPKcxqoaq
Cs6tpRwLAJkFE4z6v+dMikkmzLop9DxTySKbfH8Nsyyx2pWPRavQHZhny9KUEh5/bfECsm3qYPRZ
3Y2r2gm1cmJj3L7aXgUmCbX3fIC4Ndkpy7epu3WbvSOWi6/L1qcXHGlRp9XuwWz7p5VDuB4p1lSO
Cai3NB9ijfwXOElFDeTBoxyMPxJU9UkIX0Qb4bdu2vr9qxR4khjLHtTuVSvjol+JCqPiqZd5jd1i
I9Fa5t8I/KgLx4XQZT/4B3g3TG8LcrOHMnVFCFCXDLkYbp9HFAA9ma6Kspsp5tq+WsvP8CxSZu9Y
QL8XYi0+JDyh5pUql+hzJjL/MQOeS0AoG0vPD2QQKJRDqu5iT/OZ1CZhuwUPbxW8s2ac2gavr6CA
SaT96ybN7Etg4vYjvHK3m6bf7AXVQhbybBtfoZVmdV6LKJUa2nsbXoL8Vfmozi8mJH1RL81XC4fY
PgVXqlRGhVPuhDhhP/+lkpvBuQJD2erJtRI6lTtEkT8gSTtSf6ZEsPLTV18abFmCPcnfEJPgU7mG
zWaR/qcpRnA1jXVMT+E3UiL360JkM/4i52jxrqsZgBHiz5j55oZ9/XMxZp1WJOI+5ad8GAEGPYCi
glj1DDXdRz/YqUOTvRx6R24bdG99yaowguQP2H80mjjB3zxZ8ps/ZE/7+O4mp5nnBL49U4tGLZdm
z4rIBhxG4pego6Q0DsxBuNb5wTv79IpH4T/902g60R6+VJNs5Xshlio8ST2IR9Jh0O+IfyusFitC
yfPPQfGnDRbzQmIbWk0t+WiSmk0+Fpz3xlGTLJN8EDnVwVW2eC2I2MMAhSO4/rAgNssZWAoFiB+x
ptGEMrBtgpjp50TVJCTQc70L5SBEbXISrIPCcRmViZjrwnK0HHlQgGhDMXJY+dCvn2tnPkmkYhhd
6RNLF7LqKDjY/cB0wAU+yaqKmbB6Hasf5AaSAcF0zDA5mRY5I+nR9wznpfIKC6StZ/ThMiAHsTgp
CAU3CIy/TpWy1UIhjj8i7h+/gMeesLfSrZadUvtgkRlUverH/fkl99gri56zHJLNfMl2wHiLYuAt
1mCnhFL96pDIsD/2+cN8mRHLjO1+6jGsp0jlZktCYfkbKyDTVLy/5Z7PReey/72xoHrmZDH+Xgmy
mRBc4kEz/usj1yRE63wU6HY09QtT2kMDJ75Bozc678hSU4mY2Fv2nRFIfILfGPPUuiE5oGyzUKvR
vHCKBY6SCKXsGMb12hbWDkw1ajWUs3EfwuBVlybwfuRb+vohqgpYQ54hKgVbks+8VWyVACvIwiOz
VXpreDPlt3tMh/cUPkiFXIP/uQdyEko54x5LBnuDB0MmIFMYqwGK8SArsx/cdfIIS/fJk3vJB+DW
myeaf5AYqBy4GIIaupT8shgsvnU6N+x5L+kK1f23pzDB60Gsf0hxOZyFQF19qq5Y+8HDMwczvC3+
0irvlELr/EYwo29evkHw2Jz+YXVTaXHEBLIwujZcCtB7P/LtMiqPjB26hGUwZAHA35NhqQxozmau
oRmFmojqhalz+6EeNIaJFgijZ2yaobDupkqLKL2h2ZOtlVRIQCqVNw5p0AFNQfOECgXbyVoo3Xt/
mK11Umej++/znxjQEMXjc4wQZmfJZ1B02qahFq8bBzYgShWlUq4Bg722ydAv5/YfRXCByp1qQKnM
ZH9BbSZ5en2McJYxBWNSFip6+lo5YdX+eigNEnXo4Mi4S8RcORSYh16lyqkr4TVCJ8v4Dgal8ACv
7HPJU3yku2CUAVJh9elRZDo8qVbijg1l8o3lyXxC5SeVJTSCOS+aJpFzrkKQ7yiYt+1OQu/xbcdt
WQCs4XFVhbri02Azu0d2JP8nF2hIbKEL/kp0M+TJufG4HxakV7ziIl8ZjaR6oln5mzQJ/xKOG5sd
bzxQY4ZiNXoUPrn0e19IyNh0MvP41m9KFxzIiwKvHq8yP9CkOMFV7St8oV/zgNr5KuXS58+8SnUF
8GZRbiNdfhJfs6xsxoLc+INsjNx68wNJsBb2H7acy2V0tiApjPOGN1ZqFR2ltmXGXOVvabVuHk8z
5nEb5EHIJLgN66KArK5y0eFi6prRM/r5TJ2UiCWktOmCNlmrwKobnaxP53frhLbKKoElh8brEKMq
0Mv6f5iGK3LwLPnrABTKLWsLEeFs3jzgib51tFYK7gqhVMggpHYQoB7ejRmYDpJfdSR6cQ6L8oN1
dNXEkPkHl87Whv61MIxoj/aWjHjlDPxJu0Hbu0R4VSXkcgM3NRSAJBYkIUz8UGelOAuc2Biuoqhe
MX7LUG2tkz6VPSoWJBopy2oSWapGDvShyHrSmCj4HyH1GfG93P+hl6rqTuJEQmftieUa4Q2JZrH5
cY381jEX5Tb+XawA4mhDEiRKtYa+8INzRXuvLPtH4AqMEtY0zWt21cc1fwit7wTGSaj0UXpu1DLw
9BNeLSyg4InCDFO0CPiK7cLblpq5S48+C2NalnDb1v7lPWcf0bEBgC8gCoMS8qqcVhMq/px+0MN8
bY4/P1bIy3DzK1a7ynt2s3i6xn0BocWVAvTtHkAcxWkO9RLwCRA11dMak/pmmEy9rmCIthZglUVj
ep+ocQ66JvlcKWVlDkP072TCvEZaFNaV7YPCzPxJYK2Pq+HwL5pS11B6OznuVnnuEIbQUhBJhthp
GAg6Yu56hfxtHvT10jnU9dy/HDNKERfHSxrw3v5MEppR/UA8pWOe18hQKTCLH3+a0hfKYpGpWhN7
d7onSqvdfxo1NlGjGTWIKfieToiNfMWUr3Veu4puhLxKA96mgB65q0f7tq9YQb9IXtT40NCPJRsJ
Ep8PVbOYFNcfducmcl1ZI8oXkpj6m3WWpYGMlXOVqiMfxpgOGa3o9AGuYqNnuUuBSaXVjkJEfYcZ
GbarM/eqZ42xJ49Z998kAs3rcjKb9dTu1FUxxWVC6FWdlTe8QloaWtvGgKJyU+g18CD388pu6RG8
pizIffPKRDsjAToE0F+tifGfdi/0Sj51JLgPfdJRWdLJ4/OO3JViXEBCbOi7QCWqdqooH82efz/l
eywTF9etCONdXqH2DHbmHX7KAVGyyp22qFFv6XQkA5Y417ZCZiTBe7+l2LdEFxKp2YThQkVuLNyv
X3OzfjWetPi7UcqRYH39vEe2+ISUPM8PvEyka+k6N/HltkbtCF94sfTEcZopcP53JK/7tqwEra7W
GfqQElvgLXJExTiuR8Z02naYagp2EdX4pXXPZGtVZA5ng/kw7T89TkeDDL2l6FJvJCvwb1N2aPIC
XxQiF6ZXhnjp7SB6WQN3Ndxutn9w0sC/FBTs/MYz8pUHf3LyOaeamJtrmA4dFfhFsZZKKW7xvbCh
U2D3Qk39IoOc90/38V44gXs4h7F9k+W5nub2P6VPDu8/n85a9BVxsXGX94yM6DQ4fecjgJpKL3x+
h9g5hfMN6uFLMXBIGfJUwg9n5qAPOmrT6IOWKPB48Oq21z0QxYLg/OMioyHpL+JSmQh+TSz+O3Xc
71FHSVmMYk+WhBDW+rSaTtop9sMwlrmCH25ruIIGowwB9IS/7fCTr35wEBXPfVI9/sMwrQUL1MFG
8MhXqIo+QRquxS39GwKjW+s+TJLPZzSlqhjepjH82sWiEnxb91FWAGDNE6oCR5JCYd0nvAHdOCiM
HK/l+P4tNGa+uLjdUQ0Trdl2pRdKbdL8eKjaRpPV9ARxdzMNE7QoptZ3eYJ7+u4N8OAyq0bc2T6w
9NqIXeAqEBh6XYemrWWZd9ASTr/NU77C6JqhtyECThSon9G0fTt9DAbPXk/GqycPVAdQQea5n64u
2ESxoW5hJH80778jeCzBia0u4eu77QXFFwb3LR33AygJavO6yMaG5fJXY9Z8AiRjvVSPdSThg2Ok
jRKN59z4A9Zvx07dy5UjGuYV+0dd38n0uYp1fv3PukT94yfvu/z4m1QGyDn3OwaDpp6tv/rTzYfz
oNPOrWW7JkHbYEfYEK5LLaqx2EB1XcB97WjW5kWxarO8XNgCnB+w/Qu7o7qA/DaMAM9GIKugnMRZ
0rxscs7wv0IgYhdAkFRLgMJb2lDzhhsGC3Ccy6+iHTds5jN3iqmTld0924mlFQUUOIpz8qfYZKmk
3zS31hfU7jFCKA7lL7Eo+lIOUwGmrphy+fkOb471JZ35ImR5hWBoC3cpMDO9A2VmWZcAIoWqDdfu
LkUOs3dPjYEfFmtnGNJ7WylbKYe2y6MrI5W6hTSN1wLjfcrFui1uUflfupTQSL9e6u6xVEeAIBM/
VKAsSFwGRuyLucm6d9Fk5IGTXdYecuDMpB4pvbzMQownuquwv2eeMLhQMDOHbFi2jCcuyNN3Hb01
JxIt2gpKRAfmGP1vwFFuGOfgWvLzrfjglNedm+pUoNlVN2Y31J2JCyfh/tP3UKHo31ubczzHPBE6
mSAXpjkTN1CEVnA9pG0djqzEMdH+qHSfgDujNodJFPdwlnTQ/OTyX5Vr3kDnHfcV80KJdcDAgDa/
chq4hMM/y2iDHBaKmHrzlQo7QDRaehWtdKq8zTnkiesHQdi4IpY5zk7PvPWk+5O+22b+s9vv51i6
9q06ZEl6itKkiv7/X9Y022bNsujj/xl/unoq0L77aIyIEZxKdXbBZb5c1CrnXnPZoarDItdPs10O
WnWDDlD2y0+DnZnxVNId+Rsz8R9clkQuCTPtl7h45TcgmyfnJZ8a+baqgCZfPzhXoi0rf5y6ajpZ
2Ns6hnPPjCM+aAvh2tP1fxcnvgQIUUZIGuN4PMhnmvwbiujTsBMcvSCJ8RE4Am7/LAQneJNeatkr
rczzYHqTLGoU+gns+9NAIGPOC3Y2kRKsDymg87CHOevC+WpNk+VM45ADuUbchCSuru04fwr910xK
Xvpn5NmlQD5EKCwmVk6SS+tBP4tlz6M7UyB07akIeboVtzAQFo4JQ9KKd4+XD1hJ3hqthOFnE4sR
7e56BV7Y8tAgqmFMut0PFBnqDJm6q/DmmsLN3p3aUg4Yi79JZSbHYYGs3jf8pcwMTvk0lheoOoV/
f0trm34AI6QLAv/4b3rWr74acgfZQSsbESRLpvgKyBMB2DA/IhzMb3yugr0zjd0cVCO2IqzhzlWb
sVAdyKiBDr3Di2ZkMc2ZpY8aFJwhWA/G3NSheTTed5ymDGLCt8UatTdmgHccpn4ebxvUUwAsnjfh
SA9xVsNk8D3lmEqTHTWAeO0iGJmelKqWcYpmBxzKHSO7A4qbWjLRlHW6A+ti8QLKLv9RHoEFaOxv
z+4nND83vHQByRPtBcl3Kz2tRqEM/uZP4AQGIET7Z/yLYOZj6pgdDMs88w4PeKjv6udWyMFtR79d
6onYDzOuMHQEG9hQwe9J48VgnmlDV3aBEcXBkTy0mzPmJzBF3q3hTlXFOpwRd13CTrT/Rhi7MsQF
uNEzl601h8DosjB4wA8CiFQqXORGT3FUMkxfXhHDFKmNsPA3Fa3lB0FDpPAgXpc1/RWbBAlIBX9Q
+bHgdopvfAgKpEeMs1vJ35wr9JlEcnnYf76F+PpgaTG1+X7e8NKMTI3ZaEZVq+XmGvK2qF7tmJtr
2GjdmrciHBb0uZaoi+yLIup479nS94B5qG3p4DXNossXVro5+IIaTm0JqokukFvy1rzSk2pXuBnO
0tzOTC7+HnoRm41rB0JZfDkF1EQxI8JweRTfviG7+3XXGlbmbPHSaj2oBWjem4TP2n9Ftuae8O2H
5MnSkoWbPe2fbf2bhz0yKSustcDfliupkNeKOpp/dyooei+UJP5r804+eTz9QzsQLQvf8Rpz1j4c
FNa4qqP4zY1W7T38K0xM0UnpEBRoIHpveu5MPTaUStXHHI1RIS1A+WlCcn/a1mesGWuSxLOZjRUW
uRZX1d15BJY2BIUkGq8CYUq6P89tzq6aFPqQyJBZDZSXAlXMA4n+mnO1Q/7WRh2JpXtbldYDDQnU
EKVcH8O93QurOoxGuVIF+q6hYeZ6+ntndzJA8XzdcuiYXq/m1emXN0uPu9+miE1KqwBYLX80uBNC
JCg6EH2du8ecBV2wm34VRTd7ilBPm9EmYp7IuJphMyU0PGyOZKCK/w41Hj5XU6p+x9KGUllTHpRi
eGULbgFco3X12BJTVEghrwRjZOnLp7SfRAJzpKjlUAYznKWkWZ0vyqogjy1MIZnjkV8/JZoBdTmm
hhTCYIvzRBSUizcRQekBM8KXnymGmXNVUwcRCnCOeLfzjyBBvLDsPzG7PcfLdlgRrLVldWUQlX4z
VBBNyPfcOJkN25zLLFXFokekdgZYVfXKU8WJIkVMwcCP682HP/veBzMsHGwE8KjTk1BGigKcG9Ir
06RBNOSfUD3EMMe+/PwRVDHxmipnXgBPrE/FCUMy9kMxiS5C9Dpux5xeAUODNp3B0zqbX51WenrZ
4DU1uzIWURYvXmYh/ciYC9l5BHCB7GGDrtzsgdkdMP+pzWoAx9X/zuRrtRYWx38hZ6pPkN4At2x/
cyoQW6Zy1MqhaiomN1Mt1CXyQr9jt6s5L24BhM0vUsjEwaiaBOIit/IIc4gfyvOMqEJXqeKOKmh2
Lc+6fBh8zUevBomD7AORsv0yYNxNXs1JSTS/EeSzIi4SsL3fVv52CaybC65U4gSJa6zGlZqylNkA
/64LjZuUTN+5UtB/KmV8+DqSOG3hHBcqBjU6pm7X9YEga2P/0jtRbOFQqluiKNb4QFJTEPsJx+BX
UA9/Jw363jbshFI39/jmPFt28cbMhfq0n3TF4DxrS+FdQo4YdDW+OqdJORQzngapaWEMomlY8/Mw
03B+3xPsLHX8vJ6edRkEVfJ7rD0+zv/5wVAy27dGtXeyr0qydcuSdoRRKE7BVZFpy5mbw0ryKGum
HGQbRpuxtJSRzbeN/5zezkB+bYSKH2nZnUtFfhWoSSjoPBR+Un2B9aQVCI8gyCM5goEimnWS7t54
8LwqIolWuz8hQmhxopY9RvRXNQEWl3kmWr7QZQJ1gU/5VhHl4rZcFT828iTlKNkU775eTuGG+RBZ
p5YVqD5RsOxgudAQVbJSSBh1x9tmIRCtvxjDLAlYBFOZLlaneuCyUbpObMCQFmvIw8syH1vURFSM
GQkZhRO+d26WX4fobhaCziSsrBZgYmRR9qT37z25Vp+krMJtEe6I2AgoGq5vIyZjZD3UO+5TGcDK
cy/e4XVfeDUAsEWeCRpUs/oJslk630gGOraVZfQYzXGqzDnCwjGJlzeIEQSNuZqTbliD0WkI5jU+
tVSN1Jlv9ahqn2DKpWjpHSGUdH2HkvXmCX8xRa7x4P6QJuIkZ8hG8JXuygzZxRNu644Zy4f2iPsO
wWfxHjuCLFUVXy9hZXTSppnGSSKvEd+ExXlfb/1NZ8hqtQeryKlacXnRoHOx6AG5lNmqS2dv2A2Z
uo9t6bi163I7yemDOhjDWe0UG/wWr0NPn222T5q1Pika368gaf+hQtgrQmbn6oCX/wDH4ul5H1Wa
lF2gHZV/EidKzabBF/8jfOpa0xNHo6rEGZtuysTI+FNrDHCu5XW0q91HWRv9Qant8GqEDMJL4PW4
4pDYh03Jc3JlWMfmhfd1H5mRQcSEd4dJG0407nHLYsLXdX+bXD4YHx6joqchTKMgfmcQ78fbzBrA
zc+L73MoVQ4dRisnWWkpnY+zvXV7zF4fjyfwqTOsfYHOPqgSUv1bCc7t/Ne7h2Nk/qp7G4qmq8cX
ylKQSK09kuT8ffcxrOGVU4dxOovNa8q8/KkpPvK8x3eOGr4Ios74POM0YFgprdcVNFpvYIK1ufsa
qDJ7W7jdnZJNcROre2HM2uw9/VSfucuq1O8tg26sILRfIbmXrABuxfhQ2PNRrt8vfMH9cdxPanPW
eYQQDdPNiAvezbsVurZFbSrxw++VXDGQflqBR/SnW/KcVHol/ft0G6PsuJk9XAMB6Tqx/X3RZakf
j0F6Mc5l/QyqVgz4dnK5xVeZdUj8kLwXB/573M1lwFkvXsjkbMOCGSYMACnsmM2JEbHANgpWaWWc
wTvbHms6DvsNFsT2t/fNEhikqthVZcy9zX09TqiuhIu1mMDzCNih7YMut2yktTX6QfENJfgNCzFs
sjmabgcVyf0rS/eXNFpHOG3IU6pl2Xw1m4Xxp/t9q/BAM+4pAbSIX7wpU1ZbZeBHi7dq5FEJOnik
dNaBUPaXSmj0ihtMLqKzfeKWjp60HRuCKwpO+V+Vy5NiORb9bSFI0E+Q4OobhlQXxYu4nRzA9dQW
/7W8SGhz+eTFmM7WfFKPUvd0iznZ2Z4IIG0uGrs2qHZSDb4zl4f02sCLxsnLUmJf14af4FSD2qEp
a9ig9nLQyurBJPStglQK6I92n7NPpWwNT/Kajt7CB7TWHx4se1lcaiuBAkzn+q9c14lCtHyK61HX
2NsAeCyEveqAdWAf8gUXkt5fFF8pcq4c4kA7qKSa8Yy5FfGbMBniN+uA1Csh9Rq1ooV2aHjjfv/z
afWGYQPoA6XTOH+jREsW4cKjzRen+kxk4jQU/mXmmC7aWcT0brSEdrdCTfPOEsnJ4bg1UkT807is
yaSeP2dAGVmZtjgVIF5EndrEdDG64IU9SrX+QULkEo500rlc91aUZfllhykJyYCoNOYA4twZ8Aq7
uYAXzTnPlltT5+8qgwPp4SqPcB4PU6R1G2u8DQyzC1dX4KrcCpeD9OHhDDa7n6uW+cUREgDQgh6w
xK5dnijHIb/xHRujC8fILPBMfu6Qubq5aTo4+r82ZH1zsWQQ9uw7MYtcMOPdw/EcaInGKNr9sl0Y
lVi1EF4vZgwFEnSNu7doNvhsNdvpiAy7Bo0d6ORmBsA3MXZlhNdCRoXQv78LscBSpSVqaJs7dg1u
qA0YAv1qlQfxzhupLN5EAavavJUtb1It60/L4wSrr1Wn+DsV2+I0xFJy8Tpdb+OWEplKfG7cU7b5
ZWJoJL/E5QhHAjZ3E+myQ8RoazlbrblrZKPM791F6pKSMHIVs9Mbxwbxc+sw0UONkiolY02g/tlV
Dzv850dqDJWFvd+BmrtmZv9mMVGvFaXfj0tV6J2Cf25XwvHfO14Ao7KJdhByQDb+RUaODROHXPyy
Xc1bNysRMdmvoaQOj4Pc63J/wgM+DWfKV882afBbFnhsls6BrTXS3TopgOCTbGxQGVUPq+LxRr+6
Nr4JvYuI8Lj2OMN71Do3H+qGfKFHiryFnp7JyLdWmok2xSfXnW41vVjQOc/STA+nbNSNk/ycK0Vs
CzSds5cFRw8Rdh9f8jkw+K1fu3YYmnglUnWvEPvf0lY0pXtqS8EacRvlCnx7aNEMTBvVP7yQArzF
e6SKx4oWcGBA/bn+zjA0lc9EDOjgyb7F5FbsU/8nf8HAkYPEK5wEXCtGP855kUyF6K4HhidJOhpT
XxjM8lx5V23szsN0doCUrzKc0TZiguKER0+0olDihUnP7roCHtgycX9rW6nHf+0oXKWbh8i5TSGz
9TpCZUa670j4uAviN3HlbhCk3FzTkpXNRGYhG9pkrBPUPnHDeMPanmse5E2tBjshm62T+2QEJkvi
8DP/TismLfGXlkv/BRJP2l++vfsmXJLl9tmSNGw/RmTVY2b0T++kB0vyw92D3YWi9Qr2hvgqkmRZ
zdHrUewp3Mp/NdKxTDeccHQX91U0V6EmG92Bs1WHRyF76OcCK6OexRd1cjUM3M8fDHUZvjuaQw/B
ojOSLEM4jq7BXDAYPi642QkdF4N0u8G+tKQ29bWtvgiO+MOtnRZGeDPKhA44FF/6bz4OV39KUkCo
qRNGBYjOdrhdorlkakzrkFRN85TkxOwnltYHOnj0TNhX+zi1osEk7Ggz3anLheaUjV8eXl2U3sm9
kMvfaVpJX9zesQraQJ03I8lAIw7F1lqpDxy6hz/fx74J0Ofh5lemutWCVWdwmjD7FAJcIxFQ4dVf
CXm7eMcGpb434aIUcqCE9MLSNsAbS30Ko3EM7ioGFvieKOXm0zZccvBdGudrQMkcC8fSwomRHB7d
m+UTKgnX05xvnx8XLGnPvptt8LabVQcoG82nEeomk1xi0A59GOYSPpvnTVIPdRFGmng+T1XYrQ/u
jPu8v1mF84v23XsTZaVjEswfGMnkybSX8fz+ha63kigH6v3MVaDhjZDAPzf1PhVvmqtknhvRi732
v0WZn0I3UH8hHw5VlmlRX1e8Q5HWwoGtgsvs9INH4fhcP2PFxcz87y/n5ZcSRDJ3VI4Zj235vowh
2Wxy63B2VvJZRxQqnoB9kI9BtXs7dLEWErcizTXW2Snu5V9Ldkk+qDkpCiQpeCFi1rdpg5njZ2o9
BlKyQ448BZuF7ZOmG+K2tSLLLxE7ybf1Bt7Fttx5+jA1Fe1ox42VK9knvR322HZWNGEZP96bxCYq
3/u22xx2CO/RA+tGRQyaCfdZnpkPGyNmccGzMLfZUsk5qIz4rGH3ZX9R7GifQoKY2FTprl0r99Kd
xCs1J/Q60ob4dOOM6zOnIxHzV2UIjFxLONOMh1fV9+qCxoIo6BHVvvYKiK4bIOfylsPNFymv2DCs
lE9yEJt9wYSQLkmevc20rhSuSiAadMJSP9gwxpsNO52N+gTHBgzlgivp4hEg9p0l7R1M3/ry7xAt
xem/Vo8l9IfVF89RKYWFUCCowlhepd3RfxXzuf9y8PvSC+RzIfmuGeP/7kIlanUcme4PAxhlJSGJ
lWnJ62P3Ntxy2aQlFI0m66td8Z+BAylKzIUBjGW+tNKsvT8IwqyP+0D40/dMRO1m4fe6TMruhKIF
qiPuke2fzDCCC2HL1E6X6BH3y7QARuG7S99jmLO69/EWcvOKG3jsx1zZiKNHrs/gciL0RrhUTkBl
tfkYko6uf+ERVJ8mJ8+N8foA6ZAo5hK1QrYv4aNbCGlpvhjThbnhdOxUr/e09N1TcGt1ZkpchCcm
ds+NLx4ESQs4xePZZvygcstx30T3pa+N4Es3vrvMm1ur/10j1PTei4B+mDQ9fZq5N4kNdnyDc4XX
ds0+HOn5lH6KGiOFN0Z6ywSgzJ+mMN2JkrLbPmZLZxUSohDJKgktoGXxENWUjq+pOQNSWyX9a2wW
akFxj7RsLrQWUZpZd2k1jHn3CIhsOZI7D20gQFoRVcYJ8lwYUmB8pHbWEjE+f7LUC+06UVMTu4YW
si9WfK2tXvWXFhknyTQ+BbuFBMrWBseHH+ZauvS8G6pNIOVTxyAVV+1RgEbs0f97r2l9aEZxqsZE
b8SzjUPrw87mJarWUFQslDDk8dKh62OBlIkw3lNUexJ3h1SR5ks6oRXqv3FJljh2U0qs7pGuUEtk
E7wb+nwqsAWJp7MS61byKqWq1UTpcPv92O0h9uEmpbwjxg+uA6xehOtAcA+q8uKui09DsMxfMaEI
zMB/8azhdlmRvPxkeWesoFsn7PjtiSFij+V7cdXbTB//+40b66QShhy7QBB0gLLZN2Udt3rvr9X3
0LjVORnFPnQB8TPEGIbBd7yGVFBVNDdts2tV1wO1V1WpdLPmWSlTtUdbAyV8VBDS5nyMFu5YqBSc
PbcoPiy9pftCJbMJv/ErcvY2fmO82Fu5ISY1saaUZhBRz0I+NVZ9WqIopAHLL13Q0xVKzAw6krgn
7TmHuSCADqA/GtyuRB5mj6J+Y8BEc2ICg54jqH7MTt2Lxs6m4pRcHO4kSUTkVD1R+3ow8AaeRf9P
e1es1PLpRA44UNejY4YvrC0JyaRThiMvKzoOdWQK79iv7YVpO0VecDdEsE/zmH1JteUH20qyCTVq
8HK7oqb2tq7lXGi3wd6j5duZi7jitMfupHJN97R7qqmsvePa7PheGdD8Rh1LmjN43DTHNT4ICBM8
NxPg/9N3sRLB3SOfs5jtKoegoUB4hO01PW5e+bnqIPXkMbmo9zjFel8qrzj/zU4GjNg2ExYhbYY1
Xn7xLHIWTs7yIsu3O78+P3dy/IhOf2bypfhKFloGgmIhp9nu1xZ8/nXjxrEeCHkrKOoX1p8TtAn3
FeSpliNwDWVCY5dyHNKLIpZlE53L9E+4ePFC9XrTEZ5pdo0jfwXNbkyD3cT71mkfoo+Pp49N9x4I
8dyllMT1Xn/EZbI5hQ+kLSgYBdtvUFCYUCIlq+iyjV5aAdjY7pyff8KGuQ7yjtIw5AxJ/Lez6dIc
a+Q9yBFgzWNB+o1SWYr9CzEVzfzf7X7k0/yOJ0GiAA0hHdtKq0zGcWRqaZfCl8cCMPHulm1zTV8c
5PDSxOVTVWuUv04dciyydPQzk4TiyrN/xg1gnBRkm9HnSmhGnKCOveqhiI/9kZpzCnmK1ncx/6fJ
HT5XRmLZ7re5ccO06lAW9RtlpRReo0pdcnZPYxFds7MqQ04X4sZx+0QiZA0nQkOBz8269ZdWJg/Z
Wf3E6acuk9mW3KlhWXDWhKWDDpZ/ruZmEfbduElJmOU1rZmZCuV/9sFj3LYMo+EKl3DVMG43AJpE
SEP/xdT8Dopv/ED6cC55VLS6q1VAcRVUm50thQFXDn2BQBHnzL/LgMJtHIQbHf277jqDjnUT7wW6
Nyy7Cx2TgATAM6IDw43aACwmgBElYihdSLc3tMPTqOsEQRWuBZXlnUplT9g6fPXNnOk8aCa2AFKr
ouxz1ShyPeYPvc007GoDcD7eWmOaVQ+cGUZ+zzLMyu5LJC/mOQ5b5ExyLVZQwq5OBTeiB8nYDWTA
V9qWXv6OiYt2d0ZsmTRjHeMp9JzfMQ6ZDxG+vg0dDewBwhjnq0AePZlSzLwNlXKxSvdwjYNp8Iym
aX3eEzHOuYhYbByspBvbxoU/otwuUqc2IS2ODYTsqkfn7Xo9prQH3vnwp5HjOffsbG1cxrZu6dbb
fTxbjhqtuPQMepu8XfyXPPv1ehBoNVYFv7IsSrPgVUQopims1D9jSXcutG4iNSr9vYivd8MEn+V4
wpVdmq+5F42kK1jIUomu0K1amGtRg9Nzm44JTAvgwNcK9+bjgiCt//onvpE1QOcBJvRxdXQcuied
zXn0kLCp33YyaoC1xFNLt7YTFytVm0rxs7pr1OGRc9CxU8+980lwwSirFwrg/f39gBpiJXSBiVbS
KkILBWVGEJeweb53pzFhOZNHftp8q6CCDD74lHmnFxZ9L4mWWbydKga6Qjx2HuEwaat/Kx81CXLz
5LXgWf1wM5k43NP1CT8bqR0iMhH2MlEPcr5BXA7ZsTpVYy9oXo4TqbMH3mTLk0h5f8Qt8s02huN5
ptEAqGE5IyoKaMMlm1vJZ7tujxFZ4TngP2YZ+QP3QkWxCT3l2+QeW8SFtS9DVaRhEQOTnlv570mv
xWjKxT5ayjtThH0mWIDWQZNJuGlnKoEe/5SRlk5v8llokX1tZlwZKcn0AopwXeQn/9XIlUI2N/el
/HSNePlK1natS2wZHXVNJTcbtTmQ/yLVfqPQZFMptT2m9T8nNb48cxORrEbH6pRd/56NlVShcZtX
P2Yw/g6RSKMXHFf5cTxOcIYU5MedL/n8aEB2S00fQqNJ5b0J4HFSv+Sb3eYqk3Rn9U8XeHQ5xuHb
6w+UQfHRFGQlc+qKmCHA2S1NL2ULvPKYAg7lihEE7QUQTNFm+ttoa9rCABXOHgnu0VnBLqiSezUB
VxiRliy1ASbnpqYtmqgRuLbuLFU+f4NMpD00YSX37XxzNJ5iaEnwBOZX4Df6Nrlle9e00Phuj14/
zFRZ+/t3d2JDpVFT/fU4k+lJta4NKmk+5CFBlusTuLW3u5WJh2OGF40LzAogz84h62Jvnw4IGMfm
/9WNUn1ZHd5rM6qa6PLNxijZCXm2pMKEknk5EkwomBP+ojKOP9aT3VHLcfk5qoSb3W1nt1vVoYWW
3boNksSfLNHcfghdINoJdNnqIp1nSrm/iv/WxgmpD3mEIVUmu5bHlclvR62QkLRpAb9wZrmNHlx2
OjmftvfGaZsAScSpONSBPNQ773dUwqjEoLHC78QDIDt1BppgWhJuFMSACru0m8KhutLDAK1lvq9S
lozk3bq2VSk4XsvwS13odjDDtw4Qk19jcHcS/18wp1L4czSVD+3MhJMiP5qeOmxsZXs/NFCW9mHJ
fdPZeY0avMEo6RqABC1O/zMjoYtzAzSD45Yvo08UfdlgmyKbXOgYbDN1QJRS7C9+9iWZi+NDvEqo
KcvoOboWd/hOyQTtudAPPl1S/IT3jUa3LwV4FEHBNdiaYQCqc9SUytm2Qkz4zDFTmKiNTh9fUkPX
erFPbY33seyKrQ5PSqPuu0YMTmwxLKcnBUU3Db1V2ZSpOW5ub/BEO0GQsd1MvmR0caWqzLB0HVxr
YcF3qdN/B4gshnDLA14v8ukEW9JZzE+mwRyG00A48eFHnPt6Gt8NZlHis7NK6wnKd9xF7WTEZNqC
KgxFZ9Hk9WJaIa3XYUoC4OpOA9j8tw/rYo6BHjlX6ME4Ap0Hi339Q93Y7GE9VksJicnNEaw1sT9i
SPHC9wJPnIXOVPyKMyjBd7xD5dMjVOUpSR0VYgBoMXLf5mAaauksnvokkQJFPDPlQBkCy0szgMLG
QJVTMAH0ou72pxJ6YDZJskRR9Yq09eN/J2gQ0tpMTn0KgXyyuiNPTLf8CC5AEiGgYTP80E7EbLEP
xmUh3qlA1PEbNFF9aoi3+XgW5wMj9sqfBJJp3ypb82/q8Swpq7lQQ+3i2LGmhgQiWc7kByX04OId
GXZ/p+w3dU9bb48nWsb9kFEZi4xEltM6GoQgFwLalLhL5uMbd4k2dG+gbboc6qaIZsKEJIBuUU++
5x7k3AoYlohXpHrt8u07GP2yab/qxWEHlrAOf87jM3uxgy3q6wSiKtFMz+RjDSznmvEPjbHjL3mc
JlaIKWim0BGYX7RvwK/piVp3TIXfmdD1t8l2IYCFkqlQMpKkV/g3lLtiKU/RxeP0YpdBQOynErRS
+8Gaz+eB6FxvaEqjimOA6tEmnoVyqhZpLKt13DMtNMFrD/oF89V6VARch57GOtep26qTNXrp9Rql
6A30bsQH3pzOBvO/stA4YKb0ZBNmuafYfFsLaHF2mjWG6ffyXa0I8JjqYxq0IpXPU4AB6z1A8+8A
yIm8HB8LxAVpSONNJd38MExC3TV45iQuuvC2D9kcQxM1/nXWx6nCrY4VTpwPHTIyXSrS5WL/TkEE
ErTIk+Y5GGDVsWMC+c+CsiNDJ4AgT73gCi4EL89ZMw9B/xc/G4kw6AjuXM15dzonNokisomlwk6I
R7S1UBm9Kt2iaaDvC6gBQWwvvPXsU8vetLrJoPfe6+oPJjnGMegAXCfVI0HHeu9VljxGAGq8dMj+
+Bk9UOfQ5eeo5DmysW0tgfqHqbXeB5NWWN1dPI3qAOOPdv8Q+2Faf8AUWes4aXBqOV5Bo3pCCY1r
bewf7W8DRg8EuduPxf6dmNJrmNUrmJOiaGIIkGkKw71R2JxCJeuk0cDgSPHSxVRX3cbDBixkQpg2
SfGMSVEGakioeXDHlPA8lc1WqBPdoBv6qdENx519xevfzuvoy2lqYW39oqQ5eNR8Q6D3kVswTARl
Eb0ayASsgjukDWfIfyYghU/fqVBnTdpU7u6A5DpQ1mH6QSD6w73yeynNpzg3CeeICbrFUn4eov9q
r80cg2i2Sqdjsbk+xmxbSeDrnytBnSBn5scNFPikwzdCEXikLA4Yx/QOfL6TV1GZ3RxI+vBHmLCT
2vDNSegPyS7XDuyQ/5ha9jO5tAlr1COGYawtJ3iJamPTN8CMkJxyqwbcgdoHOneY9Vn0A4MJxW17
3y51HhjFaNBxbPlCe2cXb7K/+z/AbKg3cOdxYmK/naYk9Aeai65Lkiimy26KqndrCKcALee3FwAQ
2e1pO1wOZW91Xd2PpEvhvhp1C2eR3TSzCdJIxzRFQoa3LJdsMkUsmzoZM83Y5blo4+VKA30m0tDN
3YabSLMC8yquttq8C7ABu7nid7JSyfg1LDRv4Rq1fS2Q8eC0DLJaA0Noeqclb+gQ1T1+uNCPWOPR
uI0WxZ+7HsbRMNj0Hy4EtGBuaPKssJwdbTJfpYfqV5XawdfpWLBkGnSF8MAbBVVbsljhTdpcEXgY
IWzWCUQtBUqCNTMCo4vrC+HglMmXBKhJD2iMbRWNJZNUKNgc5ldUG9KAmA8NXiuhOVyOFPNkQIf2
0hnClWWfUS8MiIBdo22Yl5UKIOGAyyVVpyxzcuAuHHKe4t9e6mNZUBdBPDZk8+y8HBNLPMNrQ1cR
T8qiUhmsfnwkE4bqGxlWKDOUlB0vMcirqg63WORP1w4e/fnvW5h/NzwnXfIC9lDV8sdqfJlqkO7b
KwHCc2MqRc60wezSjaCnI6pCmHXPJxUZVrZyO5g4FmKf65YXjuOwvWQyQ0LOEsRzQQkgD1S+SmCG
VDFhRhaSpAE+h4p5QCfd1OdKgMsteZlfFy3LH4CT4mfIKS0uEtsqdeiMIc4H+ipu21ttfExSCchQ
i4Xeq0zPiovWixYXl4WPh79LACQ7CAbOQaVpzscTUxTrfIxFO+rPwlyt+n5p7jLHGKTYBUR4z8Ar
QZ8+nGfZNX+fPAHaibEp3A66VTn4k9cwleUYhTrfaUDt8vAQXmP3f9rUQpNg4Izg2DZtrZuLvahd
Cav3ydzKWWzTDAY2QDsLcF9CGlSeSSBKn2dk3t9exYHkDOwIXNVQdCio5qc6SeuXHDxnK4Pck5RT
2JptlkCys3NHHsmJlEj6Ca+xnXtBa/bv5qNWJejGjnopmn6uE1ziIUUzCPQoiO7p5zJMjdLgXmxu
9DmxPbvVjNAwY+0Kcif1pixbJzfqwqO/6CLAOi7SwWm9DopWE875qOhN3tBFYlrdLthraOVsgHr5
nxrzxWqdvZpnpKE5ebrBwm/3A0d60Himc2GAiI5iGtE6X/WGkKESYAkv8rSNvvg+x0I5D5kjZxmQ
x7QD+khNqZdL0aEXh6SxR7KvHcn5wKc6obssQemNNPKxmGLYUjf2aej4FILG2VvT3zfu4d1ys0Zs
D2QN3pkGyFpjL5+axE4DDh+y/vkCWhDE1/GNOazHAGNV/Yz3APE5ChdXGqdTmXp49b2Iec5bXJT+
fuzH+gRoe7MMMgOkzCklMlWuG43IJxP3JktUpI7U8lW8Y54OyouDwgYRMSFhL5vK3O32xSMJFydt
gws5e45R278+p0Jblb1i0kCHyTq1hQhPZlWpPXhaVCU1jnsvLC2uslOOguN9SS1+gcfWNKQyRVxT
pg791kig8+uIDZjdNcmeEVRArhrVJeuECVgQV5JjKprZ9P+kHWV0fCHcGgB+dfcKR61XIMhCc09H
YAdSkBIz0A/snyyaPBVcs9BE6b+eB7BEVLKdQRwsoLOINQRlSrTb2kbD4qiZRS9cJ9x+BETQUnuA
H0qt6OLnv3AhsMzpDtrCrqyj58s2o2CGc+3RGjLQZKdCoYilx5inJyEZyO7CBQ4UvUC/PvvqaZPm
CciXhRwsyBYfYSjuSLAHPNGnpq8m39QuBpm82l9GhA1NPAvcgMDYj4Z3Z8XSMx/Od3KmQyRuNsvc
lLOCB2bNSmA21gTGdu5f3YeAw8u4eEyF1rMyCCC4QGjf4SSYj+Q85xGzhg6Qe+LBAPICSXLGfHaM
eeVvkPvbpmTDGNaHcE3GG2hpf+D5UnYXd3/DNmJ80Vcm4B/asIvs8OzVUA+9ygNYDIFQyrWrvDel
aJIfCebcLmtoh/325flj5Io9g6KuUTwuPgDjSAhPPYxT5LVdw4mHl7zmcIeXHypwt4ARMvj6IEAL
irAVY9TbWekhn0XYr+IvhStCHkFZb7CX7qVukgJT2GNq6paIEjyhx+N8TatVHdmLyEZGat17C3t9
4iIkRnHp5GWUBWccty3M57NKCr9ghByqMWs9EJKNLURe0JkiNmJBhgyZAX09PtQNsfuddGLh1K/X
wzX3x96M8J8TjkBv8CvEoGrXGb1GLZpAB/SeALm5j/gZEVCDavBv84QwWzYPfEb8lKqDHl7urYf9
XKepPqlwm6VgFPx677nYmLnUNb7YySYS8BCOmHg04OeHUAPvbviSMgN1y8A4skA4dJw1TX3gz9bN
ziJoSWvq4D8DTd0+hx/ty2X0sAm32bhGQsrYJoTGENYhUVlVxB3CXEMFdit2QH3UbeZxMrvZiSXx
MOV3zlTbzIXuFHtqesc5oWR0d2NxmHrz+TBVR7rO5Lej+OMo/roAz8/JX7nTULPKczaZQmHF5BGW
wkhfqCe0JskWn+RAPx9zO/7jrWFzaLItntVxcQ58B1yHVTm9V7HzUM7vHJ1ErbQb6n4dJqKD0Fi2
In8w9Ulh0CZJ+36n3lJo+vEDkk0S/gKbzsHFnWhrwuXzicISJ7jlBjuJ9Hkl/T38ux1KyRUUHeDq
2tQLRsXX9BdXFflwVDqyOGX2H/iH4bCfxEnDSD12vWEqzsbjczjrGqoc/qKEmzYFITD739lrbXXF
PcSAsL6awgvWYz7M8tAxgoTgvE2pD+7wnxP30juhRwWO+OhvfefEBXjMlEEu4EpcZlg5o+CpQDhE
osZtqdboiq9Wue/zVOW5RyfeotmzArB0wO5ciady/5e+j9iRhxDzwFqp3Ho135jnZASiomlZw908
2ngSqKs6aC5RAx7hNGpNZiNyNTh3LYptK9xfdPxBIVjMbcms/hD5YVIrQwl0JXJxFsjpov2I0wnc
hi31Ekm0cSmQeVCm+kvTQo0JimjizjB8pA+zjnTg9mq/w/lqcZKLR2GHPy3VzVZ9q6Tmeq2r7UAA
nLk7SH0tSY7XxUYGUZbmHOIVDu7Iim/QiBIrD/qdAAAagix+txgtuz1tRoJEeFPCV0MQCEev4ufz
uOSR0ZCc0dS16npBpTyFEA6GaUCIe/3HX6fNrTG9AHFtw+fdDbF2G1WHcynWkJv8OJPuKWuVBs1e
rHDFMne+sf7aAxX+SExb8oema5UeJwTpjHN/xG2pK+knMeGMeAIqgu1V+7VQ9ekwaF4Hq9YB1UhE
ntiuT80BAfvtPSfiy742w2KtOzK3Syth96JfolVjKBQIter7CgxaC0tib8MNEFvLVWRAxu14KfIf
Vw2q7zyYD1WRlGVejUpdXwApejsSSOjWlvDI61BTLR4W1kMECt2nzMEN4d9zduSazcYMLQdV4Xvt
c5Oxhzefi2kXPlBh33QZd1yb8IWDXOlHQwROMymD7f5mdYjhwGScFPaHxTNfEhxMAwv6l2LL+Zsh
jsFYNiTs3jNtcs9GbEDZSnHu3tfjhne52yT7bwssZ3mJIZGU7WxzzI2AIPj0hbxTjWVqYOVt/OAB
O5fYZrR+tNWvrSFTXfS1Hb0OlpDYr/+yPPRBiHCpfKfBbvGDQ1ndmBgFpSEMFRZMrYNaBxDWq1BM
2EzdJ3LlCQPUs2txkN4N9Q26rdctrTkUqsc96dWjwJKXRK8S+EtIWh+rzG83ZOpAaMHQPGN4DA78
E3F0gpYZVZ/fCSkbgQme1y3pk5bOokzBdVRd5wIQiRUF+MCEMaixSKW12RVTWUJfMSdkESToL1HO
VLLi9ZdCTRmgkWpYEqqE0wh9Ho18woVw9tU8kYBgk8NoiyBjX8pYkYQhqXYTBInRNKgsEvHdhB7G
4VwKBmpsHZLTGpyF9RO71zpVmb4JYL74VkdD8E60Ke2baOnp4f6O/teYgORmfboS/RlfAZXaWlnr
bv9KI1S57bxRcjomhFu4jeYI1kGgP+hdq3VMJ4yG7jFxjCu8OJUDcljXjBz47ElL3feHg6qPK1dU
QoV6DVPEx+R8VfDqVbPsIHDusrePuuCd82h1zCqM4TNxapOhoi7+uup/f+T1UgDzmGREzpokxlct
m3QzINAUU9eXl75j/+NB/gkyZa6YR49I0hwVVGV/Cfnikg7tf08EUyhIgupg6Ur1Z4vrQH4GhR1S
JHqxh1ujW7Iakw064NAcnnx1AYn+oBy97Oz+V3cF6+OHKZOMvF1FH28TH+RHDl0obiVQUx7jUDMq
fDg+VjZ6NFcPE8LKYPRIcaON2pGNTDtfnJjdn/RD2aUJVd9PJrSDl8st9N5cdEtpIGXGz9LTdHs4
Oo/ppx69Ta71bgzpmJW9sup7WzB6hfZ94Mv1LNdjA3bL77cQ3XcS7KhqLsbD5yjNrF5obNJCPZEV
2AQF74iKSOCKeg1uzSQgKWnklUGtLXC5or2yuTF3ZS93jX3EGwv83f5NJsr34NMbx56Bg5n42GDd
bHkbhtaoPMo4aZ2/jb7rmdLUiiytBRSST9ub0xgXu/KemzZGkeNQ6XiusyRQ69LUNBAj7WaAb2vi
+iEc0S5BdTOZMkCK4el4ToE/rKqRD+LBONQmbyTfzzjYOnuR39c++l1LVq+8BmwxImKUKLvhyvJE
i0NV3LW8tNR7Le2NZWHElmRYvmur1Y0sXf5Aqwn7y9Xbq/zWw3Vtu5456d3RIRwmh/7FjeSJaKfV
guW6M1/vKf0ZlsEEe0N3OeTVRE6bWMgM3U5Z0xmX01KfvCOAs8AI9UwqzySiZzmNsmyIniyy3/Sc
qzgGuHw9Qt9M5G4JnC0+m89xyK69/j3KmBgGLvUnDnwjD5x2twZm5D206ZGhYj/s5BSqfUZwya6T
uuGS+uJDHBjwXXsqrrqQl5dvp8Oye55QieffuXI0AgY0BrX130ubI0kKRlKw76JRJpKW3Eey7/f7
qTqP/ka5W5ihUV2X1CvzRFHRgohCElcRC/xaFbOb8+fvgAcVMVFpIMs69LnL5E25YhKMAtqLNDq7
sGtjblDxD03VwcWR119suemCaDUl2To2We66ZTcIZ7iMTjLU9J8lkysc9T4K2n3S5DZk6W4PnqIQ
m2NaRTbniSclT3xaB6lLfxvtI6jKFNOSzo55KhLSkbC8ykjbjuJiFReXlhcggcnzzzve1iE7c5M8
EgOyXejcvhWzZ98MepHUzcYIj7RkUZARjsJoKGoAWmc38XvcWFkZmAYTOm0MNiUI9KjFmnkET9js
lx7IwfDg55xj0i3dZK+ZSc+pt9suwvb3vxqHQvGE41aNg1ekDs673M+K9xj9kS7oJK2/v53riCJN
rEPApCLMemZHN9PuN8cBSJIr7RbwEy6xEu+tCoeNo6vPtJkbhpAPt0Wb0IOaSP4Kji/oXEBIWLej
wOy81ZMdVjzLi0hTVPLTZ79TuCYFoHM7bRebjt/VGruGQLwzZpUBsiyja0xh6uRC1v7Vdv6U2ZQd
OuZIIlIgT6ckhhteGlfbfpXiurvWVCAywQnGCFrJ/+pmUZ+W35Yzo0apzddJ7DoLU8B9wsIVuma4
QYVzDzSyNdE0v6QF/3beSN+bcsdCv8FIpQ47SIqmQURxeSjGGRYfXDbOXSl6nA4yNRtNJca88jmf
iGXr5j+pLy5kRbJVJbhF4oL9PC2zy4wAUfLuWBsqFTeji0EIaqiynzgvpRrUckdOdjk+VmRoXWjz
vJ4BmmNCuVyDNNKedxbkZ6I+7lueUxg1PEjILeDczOFtfmRR5+YBfkREM8D8v6x+PF8/DQ/m7nYy
4Fe9WwO7J6AAT7SF/+u2LQnR6pDU3zPnBu7i4/cezEBrNhFP3RG55hB94kjxozI+E1PSC97T56mi
SquGhXXM8x8z9hnd4ynwTlRbuXJoILlDtY/Cb6R8pLwTKqwotXLUIRY5FOpNICOeFQUHJnIxp8Bl
J37N5pDeziYFqxCH9oiBN7JIWv8us1exKMzGQWntEBkRYoOJUcIyw9UUkQLyUHFvS276BIPl0O7E
QnNZPgWgKuPwWRYCqo/0CzjRL6C4szplSEaMAzsWWy4jX9gAiMfrV3oBi/H3cDbc+7bW09wck0mc
xPYGlodmwgbaohgNub9wgme4jSbFQgSy92sC+HSN/JCXL/oyLrZb5TcNTkds5HWE9mi52QaLMHT4
IHgfgil79z7HENm87s7Zgj7w+qxsm7+nyqfHPx93OxjcRU4uvkNENEUZikA4zM7+oYdF+BqS5QSg
PYYk7Q4D1kQgIzUL2cOF5C/rV69QaWKdm2DmPIzF7wSJ3kzsQl4tGHzYmNd8U3fRtAIiMnSYuHqG
FtML/h8UaQVZfpVeRHgfon+KNZr1B6mp6cAruLUZd/97fYYv069OwaYH11HGu5swOMqXVmW5xTdW
Q2P4C6sDDuYTQp5I77x86frJ38puMXSdgiqSHYch6IfL/rJiA2K/k1mPmj963GrzItE8f/d4gkXY
Qp9HiUE2U3LaMWZoR4vOEzo+PDMSyWbEt4BDKZAEcwFXJGv7WmkgFe6MRu1Y2LOQmITfAiTsW1BK
PACWJQDhCmbEsjVWazUzlISo1LLJC8L7O8HBA00/fAkzPogctGecjGBNFLSAEHOytAOouCAjyCzt
wFhkwGsxOeayvmiJOCuviazj39WnZll4yBFqmeevKKeA/06Qkp2hqVF4rRsDi45QuzVImlZbBYqS
TA38RPz4yyjZLy0WEOOlextPxR5onDm8cQ+Q5RgxgRuxWOrBYTK0lR9aCkvMJljKhO6dNVEvIipm
/viw3We9OdW6Vk8EMvvnnlV9F7itpgjNS+fCssOWgZbHFyLY2T8HZxaLO+ro2UxwbQSq+tOC3fW+
f+62/eLkJeINRYQuaVWW9pPG8kxSmPALTDj8O9NPaXKNDgPpHfpeF9MXoYv7CNs0BT+HKMn86/TL
wWLBG7AiTO0eym6dkCI/GicFJ6UOhzEPN+H2s3uK1orUOLXMjutHSjEkiAYslfzsMFgkD/sTqhi3
RGz1CammF1II6df+cnGHT90HzqiPVMrEtfsT3/I+IkHRfBv0/spcY0376LqbFWo+hGYAmK14uH/g
ZWsfhnuSPWrSZwMuuGyzVqAPeZpQ0+aJmRTr/+LHCjLkW4JqR7Wqa7TanuH0qHZoJW/udg3suxED
Y9Ah6qbyOIhvYTawQQJWirf3kqa5q8hLYylzER3BkhX7gAV9L8J5B/B82eh3BD/eXzzZELZPqXSu
DnMTN63Y8TanMpOpUHFBhnNRTDKWDemP4fHutlaSueJeMq+raa1bbXGdxvTR9paMl1HrvfDq5B+S
IrOZql1KfuxM3o6i1rXA2U4jpUZ9scr6mHOXqYThKis6JP4JF1avaVi3UGEQaBwDthBpqwpneMWh
aFtvO6mRJeC9eXohJDFVk9kL/Fqsw5BBJJZ/x48NsCENUyM4SwG6Evqe3c51VxW8fnXIL1Fxj1XN
bVAdgjl19BgGN8/ii14QMSVeRocNi2wh6AMfMyh0bfAikCAbns2Woxq83bsWdhxgHDtiaabO0/07
csh9yNt41jLW3meKwB3LLyiq+leDHWAKzaGczU+Ifj1scw57VmvP8K7kfBtj/J3HUlEV/ghgRjlc
RTGFl8dzjGzaxQk/jC7azBhUSlXTICNmzUW9pA0OOj0ZwByRQ5k2qGJAzB9Juhk3Md6g4COkdONi
DQ6YGSpIWrzwV/fehQxBtMSQjPrT8yFxzargHvj5czr1XKFgbhdECGZGjtHiAVaXDGCzwSPkPMCR
nXo1AOajNgxR73mQ1OtCAS4FuRzuG5c2eedsO7rzggL5yTEROmhRF/BnXHMUmDhQIAP0AIEtNj1J
HWqm6PDaF1aOyCJvbspW4pNjrEddpQuE3GEvVPZVHvsWpggZfajUM1TxkAalzLH4MXyFy4HSQ/x7
/DPZ41IofXQews+fM4aY6B0mt2b4999wFVRFxjBsEruoT5kJd0DrY0cJPBSiDLTKDz75u00iyeF0
mGIy9+J6dA8tyEaD8dEABigtw4iu8yIokHIL80WCwe91KQyxouSXO7E7mKFtIiFf1pzB3p5Y05iO
bYxMkAgvqsn77o255xBzVF2ULIkmllV90ODPa+4fix0xE6K0vj9aZ9SbQZlDma2gfOOdyuf2tFwB
Frzg3QCuZPuiRc90oRRHUxK9XKj9ZwCFmaQtJw3aB5IUnCMz48qEXjkTLxpZdD0BA9KoMNkVdjKV
/KjiI+t90fA5haNhyjetX9nvDnmLkZ+gC7xhBPpIBJErAP2xsYJ5t8SpOZ6JPcBD4RRY9exKuU+q
UkR+LK5Kf/5UwgSR7/h9muscYExfqVknijwXfQWFq8uTouZdbbmSjHV8Q2+HSAG+uvGNrmgD1hQM
QZ8Sdn/u9XOal+IwQWi5lH12/toEYMqq05nx9A9D8PMG8KxRbzmR6mg1TJCIQQpdNA0eom8XSq+3
v0rMnBO3gC+bRJLhD+8PTUd2cCWEhzajjwrDXBtW2nIq6OIkeHw3spESCM4o+CSGwFb21pp10eTH
lSsBoYqq8C9w9GgMHe3I73L1wKvWllJEpRp2hZeYyEki69AnhNs8Hz0GJ4RsEYLiefcz81ebcwjA
+IA009A3UrP5vwQEK9UZQtpjihvyMsy3g2a09YcsELoy0iM+aeQz4MG+0B0rr1jub6TgqCywaFCN
BCYW1QBp3B80dCpKUNh5jWQw95K/HqRVDWiSTWSjzgOnqGmLqbDVnaR+ZAe2xUQEwURO9DMGqdyB
Wh+vFWV5hGuoOeJFOJi/Ku35W1D58WbEAY4Uo4WTzs0Rrx0EuW7+eaPcrYhpfkG3FVr6lBR+Sced
0P6T8D6TUtigm0dKtEsKa39KJVP1FvUWfuXvH7ha72L1eh0Xig8f/gVL1MkVLq/oColahoh3JYJP
ZOmXU9FuSpynlDK54AYKQoyx4MFf9bau2YnC9MchDS/eyvxXmLfECDcYTsoDAy3tsJHitujt2VAl
+nemMl8gNUx0muhfeacPPZa8XMKsnf2z43Ztpzv3zWCIjKgDk33W2/DmhRAzOJDXnj/cG72A5myd
npeBcJofecIOo9NSuA762jkOCUHGWu9rH3vVmg1l/IqSl+96UM43wlWDOcbrhZomxUkSRAWD59t6
rJOVKeaeR6dUEWJVs8ZUd7tK7XzjWckL/kzq8/J3zFWHhX6U/PPEwlAsWf/S3o6iTtsR4ciScp2t
r8tnXxXLVxQjZ8vPa93daf5H0cBAnr/RgHxwBnFXLI5vZJPX0UKjQYLRYR4iAUumCSZlNZucBb76
R6QxP0+zdf4jDCHdH/coj+gDQ+9wiTxgSEaPqL6xj7/K9PCjqAo8bfan+UVAQPRFmKIFipumLfQh
31l5D+brzYd/UdPzYc/ekS9iu7ZDou2ouSFkaVF9dyutyDtO5wd4l8kYnAL5zbw39ov7uwFyemYW
NCbLi/1cx5dUtW1004GXkubo4I3YpS24eGzTe8hMcs8i2TdGdL1CFATyahc4xuZeEzxgTuaudM5K
k6dY8qbtut4x1kS95i8/gX4SzYW7Y6s79yvvtgnC3xED5M+LjZSNJWmYLIe1JeuapRK1v+tINIO+
Cr7J6FL+whFvzZ9Hmoq85tM+LO4XKsulEgObaKFM1syo57Y4AL37FBwt00xHRm0lrISDVl7RghSm
bEDdNtMYyzhVRB3YVs9CM2v3VUynug3nB8sGgZFTKA7WDctOtPXKyJdel7NE1Y//h0i6PJ+SYCzA
cH0d0WY8fPGgIYACXqBylavwVK8E1hUPE2ZF+WtNCa8yO/QSUDtHx+aW5KIDWdvYr6SjnZvSy5If
we6e8vfpqILpc9gqtQS328+gUCvf3ph4H5VdAa+vmOZ7v+ulUzQ+JxzIIcDy8C4OwP0NtGWKgMQr
wR7vsPXuQymZ1KO0RznTHrUIoo3CO0utn98XfqvT5r8XYU6ed50eQxPg+YGg6s9SgizAyEOAEP/d
bieEtUCqBiD9ihLcKpihD2F8rJXToDCIfRlFP7smZhm45U3FaDC4vm6f7ZT+q6u2LT5z5kQzcZ85
i9kHxuB1/LBdhehkG0szGGHFFFjX6jHWFoiYhYE+pJVA8CHrUnebXjFy9eSF8qDTj65VcJszAaRe
InQuy84FJqJz1L0+RVm36WAj4SGMksmEhjex0bhcAEd9GmMLT53SCBxsn1yEbgkQ4+oQDNYaBg93
JLAkfnoUpb4AiIsHrIwtO8GA98Q2KX/M1pEawbaTpbFf1dXOoCpRN9/16ZwpUgnmqJronflXFb1o
+O6MX/nduWnqELTI0FAbrESjLYbjgirqOcS3Y2nd5l8Xytm5Jf41GaDGJjuKviMhckNjcBZIyDKh
gZVBIF3dwx0H5Bx/UGZbwJHGhlg7/LlKLwNca7sKZr6eqBrhu9iyevuCXJT4GNHC1qTFjFiUrhT3
JLAG9hLct0LoCFzM2uBZQk45Ug8FKYQ4iukeOzocVuWu28mHM6J6KrTTo3AxSUtdh8AZUuQC00dy
kbDABX6rVUc0Oj+IDIPh4QTt9ScbwzwXl8keOPOD/KzBDfgfwCMGFvMclSrUeTMPAQYDP29x3inX
l23cceyfaqhmV9crLQjUJsSx60B9WIeyF08TppeWmvmmT5WWPman1sMhPcNtg2Zu6uF1mqYyd91T
K1dQNzrLqlW24iSsur6U0NPey5t5yAASlsbWL0bZLl3/iyqgbCeaGKai0ZS+jM7wM8uqvFASruBr
ixNskjpfHVQX/duSWoIYAsCqGRe1GMHVVDdYit3EnjXhX0DfKPCrLT8chDh63ocKrdohzQkQVqQ0
s8oCxaFzp4veTQr/h6tqEh50WOxfQmOZDaV9Eem81IhlVavES4/AZXRmRLoNkoZAqZR5kKZ4aPIX
JkxtILywWI3vuE01V8Udq/KCmMeHZHNIGve6CcshIA62nHAS7SOF6p/KJnqEE2t4+7kDIVPQXbJh
5ZoJIYwAwOpEnYNTf+tVBFYsBu6pqoOgJ+ooUoi/LHsTBHo6vzhtJa91jYOLmMK8zwh4D28TH2HO
vdRokl8pTegl/04gUsdCpw+fovfBlH1288O5kehZOUYVcdH10qTLIJxjsYwtQ+B1Cs/ge+Kh5Mfj
FmKZHMkRT0DVmBB8G1dlIgJbHOqgVZVQfYoeNzUXkByZK3jXp+R8ZF2L0/6EBr2IkxHiR3kgiKso
Y4iKft/G+4/hYZjq10xRF5VAZrH763lgKZeGjYwvsZuRiJaeiOIgk+c7rqrLl/z6idduOcm30N7D
0g9BL69RizCIs65pK8HDmDGYS/fcd+ItDhVKIsKe05WdoEzf3tMJlb1eK1f8o5sct3GKzzlIKCAF
61NRk+XJ2t3DM5t3dGoWziTh2waGgna7jgr6bhQKm1vZDXzNVsQH6YdO7TY5Uysi/U7qRoTlWBQv
uNEfp5+KhTR3HGVMYiQl3rn6AvyFivI0Vvf1LKIOKIUy1WP4qdomSygwuQd0SyGHbLFYj8VDeK6Z
hGbLK8D5kOA1y/tpEf68cG+3XBgwL8162xrZHW60Ie+Hcv8CEHhNobu4moQwHqNIWuR7KQNCq2hl
k1yf5oiY2OYzKFB9yYM/uwxJ4p9QjyNuoRqssHRhED96SS0U3R62lgw4CS3IJmnAEVNbQLvR0F8+
CRE2/bX8n35Y19eId3rfCINGnF+vXxg9MrcH1sz4pReW/OE56iOeMQKXLODLHJmKZxylLbKHfbOF
x28qbbzeriT3R+SnLZ8viUdk+w9JVv12HlzP+vWHov+g/t1PzAvxDhlWweV2EwvsghQLP76/VIcG
IT4jWsKOakcpJ+W8rrKMcG/yporTALVOBK0MTcJmFUVJ/jhndgSezqF71dDEm1WQg+I6bKR6IH5h
0U0DOiCbLhWj2cc/GQYyNqLu6Ys0g5sCZPIvn/Xd6tuZJQCapvG1sJ4ncOJtuES3R5QCVskpk16Q
sAIhE/lis5NEJHWX8w8/kPaSI+vHXOGwW/hVJublXpWykWOa3UVwFMI6CYiRJ4+TBQObUBwl1CLW
qqRao1/vnRbaG52AR446lHuLLZktfHnRJYtfqnBhY5t0Zt9GnxVCzxlRVIiA1j162DfmS6yzRhuy
C+I6kNuZVgDgJm/Qxa9Etn8E1DBXYd0idZYSKIdqFyMJodIACLbO8jU/mN8nisb2Q2OYNFbavAtJ
CAcf+qFUv022sifzc4LUZxoHzBIAU9L0bluZQ8PMtsiTZeCY7oYafhw0XJ4NHWGOqju9n8p7HUJY
gRCHApmAWywwpzGLd4E4W98TVpwfSf0BIh2tvOBgFQVdfdqFZ/SO2WCrgnuZpwyDuA2gb7ufYARH
YKXU1p96vw8Nk8ipv8BFQ0LwyEnEjyf9NdsJOCy0wzOk9QjUb8tNUpy8fbw8SQVMpzECOpg4YbPD
2DxEY3fj4Vg2x47hHuj5aiklzQYElbib3Yti8tS3SnjVn84lL25VVXooZPSo3B53vcvgtV4o/76P
F6uVsQhK0V6udMFyqgLDm5DNzNCgSlTNmxJanISmNdCdbo5j4I+Rcs9xIIwiH1KJf/Gd1Twhe9mE
bqDOfSq6aMplR9dJXw4A7bzeJcN0S0RFoMSFr8yyVI9XK3Gk5Zlz2BNi4FR7ixFk9MIW3HnLVywT
LT9uCoJJ+moY9QPDhKGVmc/e9zZe0Ed7wmoL4PAw/kOsHUin50tGq0Dschpcvgc0QCXtIJg3ASvx
g/RYBVUcyNudEh3D/tBHguvKKJxgNjP54B6nBmDQEEnLxYUYE2tdvHcpNbr2nDrIkhbex7lPdbC7
DK9qwTMMrP/B1n2lPHDqPW60DLtqfe9BINi3jpuWIh+WXiPTQjt3kuiL3p9TlFUCgXYX8YNsCyms
eNXAO/7BLhOVJG6wd2AgPE1N8n4YEChpXSFGUsxDxCGmrJL531+zrv3HXMZvVOPWlNnUYQgKD07/
KjSlLYCmCaYWFXHymx7FzE05H4Zv9/q5e52Z0vDwS4B8w5TfhW8zo4xZl/ZyQZ7qdieWpNYu9KpZ
auLJrkN4elGi2Wk46qL426ObbjaX+l9mnxSwV/nfWdEJ8vCn74Upo2SBZuF6f1B66IVchKCegsnN
Jh1Hc9q/E1pK3AceFsp6FfPfx3JCln3Tqwjoi9zyVXeYVKl3BxyLuU0kkGCQ1j6Cnn/KQcCTJIcH
hHcprogjdPjVCbqXYHxaGr2G/+Ga4OcsGqgglrAiSTAgR7npVnPCqoOmMI23AouKNggXxJ0ML1Nt
VNVXYWjxqGGk7KB9RDlp0jg8QO+UI0PCS4mQINDXl/dA08MaXTMdDqtU8J+VVM0Q1kZhk6GeBLtQ
Z7S+Sj2H0zoA+Lt5ga2u5nvIdiMUYprM31ziQ2crK56eIrO2ZXMtOmKdAZEDZUVDZ9NaIBfCzxU7
1ixz134Riv2GzARuhZL9oeOygHbagNQCdzO8DzuM2UnapvL40dhVg7MTUH51+EJUg9W+IpQGGZZR
QGzFNjSPnYTT23gpGIpYWDujV+Mb2SE8hy++hxT+ypSkUuYjylxr34osvLBvqC2Q/UcB/JiAICTg
JLsUkyP0KBqsFjTH0tKlpJWkQLOYk3i95txQuWfWKeSM/4ebp88KrDppZFE1/u9/GTgubM9+Sp9V
lfjIkCCF0gHwldv2a9sgONM3uBhA6D9Oy64+95GyDrW0fJJOaape/erBX/wmPOB9h9b5WGfuM8iH
rFTkNo6ZexGvfmhZsrlvMNQrs4DomNRe77AWHOa+DrUKHN3uaoNZP/d5ypoMzoRwuEMf4ePFVPTR
uj3I6Xs0MNc9Zo/PktM0yokSC+eJ8qS9G50J7NRit3k8RqEIyUcAUJV4YHrjuwsuuift55GxDIw9
vsfuXKVEiRHcY7UvoLJoDxG2r4ZN9QvhABurWSckhV1WGD+N1n1sBB+lJdIL/xD5WS6IxZVIISqF
JlGy2qLDbRLp0LyieMlihYSPog5OhecXVLy8rvgT2YD/W4H+oiCI3haE9pMczkVUTAt+ZSsIXyI9
rWVsIiOI3rr0RksixMT4aEHbAIfJgKAOo8orn63E/Yl/8CqDwMFdHleW/NqKDQUbeQlg2WcYE2G+
u+uUtWUXZlPkBWrG/nFfSqW+wSCgjyPgzr6OuS+9Kav0vcbJholj8ey4mI85QwR+FVzwoVo8bFol
AQeKE97CU/iEe2SE1Wl15YyO4GOPmUaA0HQBhsS4XtQs6WlCYor3Wog0mnFgyKJ19ssWb6kAV6DH
oF8kCdh5bUsl6/+3hGIGTbTGvp5LW+oSjCOVgFkzsO1eMYWGMHvVhLlPYB2weKvLHTtVyXeUqCMT
exZHXbJ1IiKdTDXnXWMlrepNarzTxn5z805y+JGP83RzmUFxRjrZ5XjONzlcZBu9nMA0+s7VQYHs
hexAX7A6KcLa/2IVeSfmYIuGyfitRMePss36G+FjJZbwreGqE0qi8B1nrhbUGb7dMoV6tBN2DO73
ogCa8LJ2TGWPQId18mpWhZU4yhOuzbq1NKIwaFjjn3fzJO+b8yKAi59JL9CxyZ0KnJSEW6B4URXp
tRXfBLU7teNGRMeVC2L46yM/zd3YhWnqh+1w/JCbqsYTOxsaD3o+lYssFubVvgaCeTOARoDHAdYr
K1ldhoUee6wLk21sBS5q2w/diLV+Lh5eEamhh6RjkV7Ju7HtBmWS3PqbBlQkrO58cQToDoOHro2u
Xu27HBzQ+TcKuZEvbegYD/SGAuRYK2lgaYgGIhogX5KcOUqq/lDyuogMqFm/PKEqeg3q0f0F6n8x
efNqCKDxj5XT4uy2cKzkYpyEoY7TfDNlC5qBeZbl0rlcVrBOiBKwWkjKCBuUPpD1frtDYVeQEnNW
gGDC/jDP1nHlCK8YXFs9ONxMFXu8S8uJPyCQS5PaVdUzMXYAQQfY68hnWhR6r7ZaZ5oVkYJwHHvn
1QIWvR77jeAohjkWDEyxOouuInGq2QDJyMn6jFFQz+g7w8oVUX3C/eP5UT1tJfkP5n8Z0EvxXxFe
JPOQQcd967JD+3vcVG2IDN+iNTrrGNxFgic4YdDDJv/kqpY2d5+34fNezno0cbTuM0cPN6l6+PE9
/aMzcV5b0WRNl8K6IpEKMiuIb0rKWnB+8ZZi+atXYVW7k+UUO89fdN4/XwTLan4XF5ZRyz7EHYkh
Vr5jL2kx4peRWhJVXkOIx3Tjmw44+CoTz0AeENLVAn+6iXQ2iBY5zTMyYls98YO+mQD2S5PySncR
0JW+NLQ0H1W+b+ZnkiNTUOEggZ+36I/GvtXXaLwcqyZEiJgLzq/D1Ly4qMeTiyU/4393lcDhklK/
fpuZElNVJ6yBjVc9biFTgNcJAOIyLvS+z/WymCaMDhR4PbTNv/iQWN9nCiTzwg7BjkIfcTi4QOsB
0wqZQ2Jn2Vc/qCsJ0wR0/ftlQYzKlsRJhYjBKE5kJoyqc7qFCAkAqaSvwIXzqUKPiWgbszI+M2Ej
3D8BRlC/9AD0j1dE88gjUpjGdn3iipO5Zao6wQWczB2NTuWTPD5ErVlq6zkLuPhTLeGVldlI7Nxz
vKJg7JvMb4kOZwwfMca0FGgeUwKtxz6gKmoQ+qKRA9jrD5L4IXSjUlkGkX4hx7sLFZxYuX+4adMM
rR24OyiwDQ9kSTVTZnnY88Z3DohgtlcjvbiIr79VEKMcC0mY6zZnOf1W54SYmNgnihnLKPQ88NpG
JxLBUHVk6sh6EputHbsDJyJTe0BkRh2NOEYoAoR482H7kVNtj5FQadsYq9qBs2aCi+I0LrpWsf4l
J/ofOh5eIyClGkvkx2UGSWvey99BrHzk2+jCjefBCcaWuNxhQO9zv02RH3ItmOGeRJHAu34ditjZ
eozMloSgZvY0mFqJkCw3q7TaYFYrd1OY4brFNeFywAh+/r+yLbA9a0JalxI6L6Mn/11ygR83RNxc
6vs9E3blp8chkxVs2DrXMJj+AZY97TkVxQvwpd3ybRgRoTZJ3Nzht6D+FpLG2p4LqO4+5xfmbx29
btuvPaOFpEF3jEvDkeZcl91uIJdP1PD+j/dfIE9+MCujoxT0HEsmeUBt7dTI7AvEGEdMXrxOGfky
wYFQ63kZJDMwzxqGjrUzKBKTJPAhZaBmId4b4jAvv/nf0s2RWiU6mgGw1+BM28hk6W7LC77fl2Bt
zFQtDVkVv8LvcxG78i3ajSV0G1KxjAdyVYfmAvKPa4V0gKgCfZ+sHaXi0HpPPWR+7oCRTqibrkoX
6jKRzcA+cn1tf23bkMWib3HZEyncPyEWiRLriHmkA76xxlZBmlrVlcYVppgqx8/fbSqs4q4S8/jN
4JSXE1ZAgW7zxXtGvqte7lEcIFQrn7H1re7yHVvw44L+As4QNWCcfni+Qp+3ppyXvej1+zizBccy
jqqCVDwLRyujkjRBwjHrQpzWGSEEfaAVtwkAWhgU6tiiUG9vdsQ1AoJFQqCVDmGC4R14Nv7B2MKU
+QqyJJTkC8q9+IT8OoQ/1G+WT01BJp3YWIqSb5Z3GEOURHegPJtnmKLnhcuSD6t9t/UP4cUw4R9Z
isSSIiLF4nHQIo06ZcctTkZdHm5ZYHSErBFL+LdPE5sA6/XaLJ5Ol4KUo1vG+S0Z6zzJ0LRJafnR
mdjK3oQW04lHRUFt+YgixrOfDKG+R5mV+ct/B752UOT0/Xox/rJBvmD6ec0uBCppwL6SZiBdBBsr
NX1GZgn38a19+kIPLjVSGjBrCVAkhSAouYyJQyDMqsobJE7JUFrKfZ5f6fiHHvISU8iogsfpiO+c
fOqqQvLc2faHj5Xx56HyJE4l1dOIljtOpSVwD36R6RouO2WRSW9yBILlrbRzYc2o+LC9BNgyLEVt
u+qENIq01t26CpzxPJDxNUFL1mio4WYkSXYZH+18ZoDmSn3e6+qNfO84Ul3+7gA03mIuQOcu+5zr
CKMvi11wPo6ks9u6FCPv/gicstwrGh7hrUjwWCJGbaLM6rurZ+D+z9QxOSu4nrpUrGToVEYscFDL
Oa6SWCSOSFbgPLGhxkimBJXZwGIASFYMjFyzXzHfpx6PgMUbqvq/1l2E1UFaqoOPDDwnS9SKMQf1
81IfB7eysaUiE/sX4xTW0ceAh4odC0y1KUEuUq2447IfzxSc53zcsP7T5gO611GKW/JF/UPcFY2u
o72KT+IHHQN4vQFSpUcAsAfN70RJ9l/z/LenTqkwbXFAKnWl7fRtMnOcHe53EdWsAtgGxR2iaS3T
GuBDS83rFtdfnOjaTD+uE84noBi2ms9uFtnIrbwctU4OpLFyrtfU6oYeapq3vCnxal31aCmHQBqQ
xtRdYJBoIpqjpJsrE0YwwjOSKKGTpT+O5H4GMuNoT86XmArRhrFfNqTHe26VGfpt6M9j1NugxtOd
9M5qVQbcz9CtJhvjZvCMqMPc0R0BDYhM7XXzqEEBUmJlTRRDnCQguRj3QaGs1ljihJ/MUE7O40h3
GvpXYqK87NxrJGG1YvaGFVtJ/M4yyu+S5GVoTxihif8Nv5dd/Wj2eihJBLLoaWK16Baber/YjuH9
ZnbsTKAFYNrMw02Hpc1jBufBYs4l87yg8PfAFZzHJ7MRk2xLjo0CaAIryKkHoZDrsdlWMWRQSAam
F9bain4B2chuXV4AIJI/Ho0QwvHKsbuO7mKtlsXOi+yuS6gX7kvTN15x2UStT4NQXhNk5TpD2AH2
KqoJLSMYZqMg++W8aKC+GGALb9eX64dxbCgieJiQgf0f5jc201AWQd7IaieYrHPuCzvGuWeKvrmX
Rr+04Yfhc4h/m6OGvVT6gZZzrmYkto1xcg7xuHsP9a5UGc8pdGTviIMIdR3jZcjSB2x46SUT1Idu
dUv6DSwNIw4PcHKrVtPNGUTYF0k3v7n3Nz5FtcX2QtNqVCA0d/vsNrV0BkLTLqq769i251l19UuU
SHKYvYDGkrpsxCyTTe4jrbrSzH8q3yxldmo7vWfo0+lY8OwyAYZYCSBTwJWxeos19IpP3ZIUmvuW
5p9SBq61wzljr/6YOgiO94IjHSpwA2jLM28NHEPZMNWWt08UZ4MIuCWZwDoVJOGXyUaZUA9p7mFk
aE2a8v4dLIQOB2RaMa8CVxRYMc1oZzEbBCb7jLdIwJe3fLc0RSVrDA7vjHzByxE9h4rwt1iSgDJu
tr8GYc7R3uTJrqNVlVzM9S2X2cp18mlIJKqd+N2QLvAT65V9RHDrkL235mCRrEuSJuMvt9aot0UV
BPcOUKbaS6bHGaj/T6765wJqh+jXE63EQ4Ly7YIhcIRPd+c7SoLnpYiGc4o4AR33EY7/AwkCWbjw
H68P7Jh7NgIPRmbb7eI9w2zUb7cNYd8Un8EtlvHhvuzm90TLa8rKQctxCMLPPobkfzc6kPOMkhhM
48wXXW+DTbBgzKceyD/bjtXA4URPKOgag2atamUg53j40br/0Oy34s+bvkmwRStSPQkvasOIm0HC
c/erKi+juzooWm2iWKKxcsrhGiWHZEXllK64WGJo2dAlLoRJMpqZWyS9HHkBlJ8omuyB5gDFzFUH
Vx6AllWijGCpII3DI9lUeMYtYWWOHwhX5m+KL80V/I6tqazQDYGekLEpSvcxm1Kai0vnMtowPz5P
tOVJLHpxCjB2Faj9nuQ1oajJUk7o4KdujHjEL13EU4s0Zs6E3JtsBz27hRaNZtisC3srkNW9cYJm
rEf+sqwJbBuMYnCXNkWnEtZGse4tyUAUXxr7bsWUq7DLVLZKNuO5sAfyPUbDsQjlaEmfTPgB1sDW
rDSTVk6exTtzFLztLFpUFLEP/19tqpbyQtvc5o1s7wosjNm1qclRT+dlfs/AIUjrk0J75O3OUxAA
KtipOpUL3Js91Z5KMMsyW9mHbo1RVo03eb9OmwAwV1ppsxsbHmG7UP76Esj41yNWWDTXzEp2bd1u
AMj9qXd01PmfMlWdZMpezQLr5dCy8msNJROha3GxqOVNgfitlCVWAcH+LeV38KK9fpu5Ui230C1a
TFLkFlvlAEh5nKTNw0qE9yvHP7YSZwp1xYrFsZfWvyQ1ugmXy6AcFnBbPzZ4mkojGZzZQMOMgBmh
UJVnd1C3bHNjntkWSMwih5Cf0c6Ndg0DsG7GPlZVNKrSK2icHLgoMV26hFSx4kts2pT0rnwV7out
jc4hp+BuKrXWPuWnTSttrWE856a3mSB7xuhqpKq0LMFAsTgYRaWHkG1pVlHuSN8qA2vr+xakENOl
Po65Pw+R1IsDMNsmqZJEU89yGv+drL/bXe9SWOo8rgbz5ZrRwl/5PmPt5++iHP7yW3s27KM3jGAb
tnCQcV3HvZgeFCFm9asqLxUpGqQL8C3vyeKYiUDeEAsbRkV20DLxVbyr/EqEfrMin6eqMcrb5veF
V2tH9MxITgGWg4kYhQ02ouCvDRGHJ5oOuqW1h9ClwYWV3CgYKZDJ9YFd8q61fpccecOozNN+adjK
ND7e4qWgUj80DG0JLFgEGXVS0NTJwSmbgx2nfVt6NP05ebtA+v1iIw4NoeJI+pIpwIOwro8j6+AX
4eiWZGdo5WFxps9nR9Pq+I1AOdUaMn+TpxDWzLD43ZoRWYJmVm5pj75vPV1WVIwq9KChY3A8yVTc
a8b5c68wrSu1kz5F/1En4awNHeHX75ChUaJt/Cf4AR66ogsyQ6FVZczM+RAmEPiysa5dscJCt3Ar
49lSIDl4/ajsiee3ukkUxUKdt9r/gAPB+V74K3le4U33jR0VTH0loXn6USSycvYOLutE/UzSdjeY
urMUKF1lJETPzcQJ26WQ45T15uE3J9MyY3e5O3LVm6Z/p8sHGGHAckOEW3/sEWhbLRKgkliS3VxQ
ezOm6SnmiTdOb6EQ6iP0qs5SnycLZFcTt5E68lBygb1F9r7hfOPnQVXlJyUUM4myzVE4RlJ8i3Xj
mkP4KXlQJ1LX/yBBb2+BdDNNqCSxzfmJI7JWHOmDYgOjSsEGXeVpfIfKCLGvRykltjEfBPayjk2g
bMvVg9kyPHLY1By+Y1uYjJGNF3g/B5H/EwCHyXCckPhiseGAD2ZuoBZq94DyxdOU6Fa4U3rS0yPs
llBDl2t7SOJqcpQtoVKuD1qvbUIllTQx/695mGvXnGddVlqYG54scBfLLHHrH6nTt2lGEwee7LFS
rTFz+9HvWPvHcf8/DDVN2X2G/s2JeJjAbX643ezyS6gUyKLvgfAKCXo+C6hAC2+GEMkFuyc9Y1F5
PEJ7mz9i0QZvrLu8zu2gDarxVzJ8cpBoseYb7zfP0nhu8bfMIXGUJFTmSvij3JWSM3HG/M8TpbSR
VsGPKu4eprdpiCJ7BSeEQ9/LZdEoUH+yFRuv0dZayzd4VOT0yYWZNx+L58Tp8GiTtuq1l3bsvirf
4cnq55wLo9q2DOhxWB1dWuKruM/BnRyHJ/kjQdr4aQhk2FiBz6CdsC8Cl99xwC8MlSisKKc3DAg2
ZlTFiRPWMwgL2HpTcib8Kz0YBlAiM3COkdkEny2AA3DScRRg3EoPabcgITvVW0kcj3u3NODT22Kf
9PtOY4zxO8XBSPlI5wQiJDeKzf3InOZMNQFA0G5j7ReGIG270YdHSaOz00RuhWkJsjRCHgOfyWt4
1MiPfg6/l/DwpZrVIOxwUWUv/9rLn2QsOvZn3jcZo9ek88VDdpV33r0r72rV7w1+VmRyTMb5toPc
QQbqtEfunJE7AvgqP/AapUpKMsAWxLPB0hDnEqwsUixaLzxuI/LlyeIzGsU0VMx84uO4T1LdFzJw
7xuLGRDuvY1r/dTygvXPlGSnFcAOA+kLqN7mVZ3Q1G9auMjahvxUBFRe/mwcAU/qD6vj/3sv4KS6
tTwR6emMf0oU00ItFy0n8yx2Md1v2mHjqxL17abMK2+kne7dhuRyuzoFpA+l/agexXwD0XxxX5cH
+dEOFpN7B7xxEfLPwFuNVLYFXei6KOB/sfAq/I/vFfV464A2L3MTVL3NdXidAot7DE7hsKLhWVQU
Du6GoJmfNd0fgoSp1cgQD+spwTiUR1BMD6q1rKjtnCZMJPWEJKQ2pHaBhlaNCAkFm8+51+Zk3OPB
HE+FqdT7xZR7jc0nfwHF+4PCixQpa1dQmEAjDxA1ziqn3brTvRnwowJiCeGGNnkPh4pjks5l05z/
3dQPKXhvv8NNY+uTZqD1IiRQl/Dg63n2LuoUaN2k8M5PbZvVqJZETXDDIGd+QBthna1baCcRbia9
OKGhhBFgEzXIACC0rVMQhNcTEIz/qWTaB9nOmCCnWVFf/dNkBeJ8ift+fg2oSF7kmK1wmauVZd4m
jo6WHxa5ZQBH23ZwMLkV95kZLokhNQ9+Qq4JbG67nP9uCQ0QrFMtDSh5dIZj0Uyln9+aJCUr4U4v
Zdt0gEUC+g5lBt4KQUfwKEhmLWl/oT5tPg8KhSD1eB55caZUauub5asI3LeD975pApnO22CyN4/N
vRv9wbeA9Ndl/kC0eP4X0nP6HSl7UbzBYE5/iEBRmcV/O5fMIY01bjUBHScIaqUFARwJ7/cNXMwQ
x/9O2sMWltNq8MeEhDONWXdfl+5L5Ra/nI8Kukelul65IfjSVVHrrWPbXpZjh7uoKfluPNPhHZJe
gR+a7lrQz4AhkAVOJ02GC3w3G/tPZ1zl4ma/czRAi4Majkw7vwhoFlL530i5NGYWm3NV09KBlNIY
yjYb5bp4jJkgjob4Z6gUobdncyhee9JNBoYgBBuy2EjNi75qS61a8wxveJQ3g/SIJDMjnrMAeU6M
RKSiBRr70+B7MuqaYGB21pNLqdOmcHPNaYDq6fIgepI8SgBmssismFt9RiYyMqAX+4GQPbmhmKG6
FaVGHMonxsSA/lXHPf0F63LMciLy+qx01rir1kCcsaYNlcjnCO/4ab4SrdsSDOLECLK+JPNFKJUy
FK9QBly2mRe+tKa3SUtj5ubyIcyq9sLeyeJJ2sxO+MzY4CSd9CBaVUmfreaibXGXfpUcmDOwVsLc
BJDKwc5Xj1JfZaNnIj8uKbKI+GRIXUCPiiSAFWgqs7oTngkdKixsewLpPVYsyJVNriKHBFKt1q8G
JKQWtMHmiVL9a6oDcX7V4Oc77DmQ3IZtyAnNER6cN73GptbYjiBUHqKc/YnlwXtozlaeqstAKg7C
VkR36/DqL66HHzQoNl4cNHa1PPk0hpRubhIQPMFkE1X6xf2vSajeksoKBTDpisFhAlcT/+Nsld3d
J3/sANRGuIo9hw14Vnsl9YK1Eg7FrXbPHVw5IfS1oTN8j2TrVvL4no4KgM6piPWJ41ZGE6LoGoo9
ikoASQDbYb+LWm2eSWJ7RqjvHrcD54t50qw4Eg6zQ0fs1t8DrievZDfcYzVnc8zzKPRnaZCsJlqN
2Ah/yB3guCby3KX1IQHI8H77mOFjasFmq6bxGfuxgee3zSFwPTXls024pXGdBYeVLycxOQJxhXzV
kT8+5wjdgZtfh4LRmzvLGh/R5LjdJJz/H/9cgJ6WTrWb4jQE8Zeqnifd/3QCWzZx38Om9TOmpn0U
2jhbauQfMPzRTHgR10xjQM/VUKqhBAYdKzvi5UOhef87v3AU2zF9Ua/Ba9hRPp7oahFKfgXdLOt/
ZMtizn/2Jr9Nwcdd69I4tRiD/uF2sjT7hm+N8JyTDRCkrkCb+HeFWGDh+qwKyhLDkp8k8ZCtNx41
HBZGc73D/OjT08cU2h2PpMnVUuRvQNtlQMn5s0QlOC/ttcWH8G0QtHt5BsM00BgLrRVHwFWWKzk/
jhougc40/AJhj32wO7VeZkCsRYl6t2kvR/nRrg5SHt2kGmjlwh84wiZKSGAEQQ0Y5U+jpUe019vP
0AYZks1mpMq2WqjYb2/3pw/4DRZOGHC+ovh4X7diz6L9y8NaCMGXjCX4AqVni7ZD9iSs58tsIYQo
nthdYwOoQUyFZe4Q5APl46ajoFRI12Hoy0F3PIBx/i5/sgTLYhi+RK5xvhrpqWB6bIjy59gOoUlN
iJBPiRxmwdRjYpyDJBQEc/m69NjFMw56w/XHToXFqq96jyQHjQEFqeJqFzLee6RzJV2g5uulmjfb
UDKAWsMnsqPdcRObMA8fSgZ6WmKgWRZokUnnP/yXni0lS2nK/huVywa9xZnz0LeW0rAf7iJ0ges8
3lGnHQkhclNPJpOv5fELOCBuDAFjq1YMPvKq813fDUMvB86dnsf73D1c41uZUPczCi52IBaVhBNr
u9tJU/W+00krrbhyaWxxvUZe3Q/od5X6wO2WkUe8xdeTq4xxkKlf0hL8u+RoA3K1M7bDM/mlung5
CzKf3xE3a61ZehVFsQUeux1ALw6o/YeyOtREEq2OJFlhA7NMg81a0C9yD0l1s7zo+Bw/wl0eIh9c
GFy0gVjgwRJB6NvOaO3kbh4hlBRKq3BnHVoWIDzMuHQDFs3nXIgy3T3vAnqI5xMf+DRz2TKqB5f9
GtmjZrVrF4+UGMPmQAN2nDhGjWcIf4dCTdNTLRjVfwC/b1FvsIOmvBtZdd81biXkHGOkW5oTr9xW
QUuu8m5bQsjSyqF/9089zAPXsMp0yHQAjT0E34UBW6qR4loMHCn2ZG0tDqI8Sv83KPirVCr4DyiG
1KwyGi5j2r8l1Wy7XeruC6+YBknJkN7SsmHkHBDRcOw70yZo6kfs7Q7dC4HUJEXtxkRe0i1jKJde
Wk7erz3yZyS1jroxnM04DErNJ1iQimPva52XAWCOMljBelmESY1l7fKKbKzi1/ygrLjUq2wE/qIL
ozX/XD8wc/kh2DKY8B+IXfrpLuHpABY9jOq5rUDcSQQpEO37SN08GhuNl16StpQCKZQ4iLFFupEl
K5H36cvxmgGng8x95TAeJUZqk+KjIpeTKT4Va8jwdYg1uKwl3DvtuJ1LOORrzbgOfyvCQyTDqLSx
F1NSH6x98CGyC3WeuGKY2zLnmgR2JZTwdTuPxrRbBZK0Mlt/VzrGaJzw2+zmFJeIBPBg1ULU3C8B
p+AZsVMPBmJDEvRuUY2mYqYF4IgYx4Ur/IIMDaqar+plUSAdS1R5iabl5YEWdo119aF7wnt8/ql0
uAVmoFrSvla4NtpteDNgCUGLXtOBHl1/sRpjy4yWV5S3lLwg6OFVO7EpIBqohDV0dSCen5V+n8Y2
ojdKub46G31cKsvhJ2WwhQ54pymHqdcuaf9SCehGgvhngvyQwgvtp4AyXTdNIPFTVTFzinjfxjZV
QmKePvXjOCx7rh/gDybg5d0eJuyiocLnI4Fc/0xuzIdUWJz4etQEeRxSkcVzMkYAGIi95TeQFOqP
DGpyASKHz/w2VVTV8AE0LAJ8nNiGQ9YbOs731XKGlC6A28Vncua40fdo/A7L1PkQjde24c20X0re
WgdUXo7qisfgpQwtv+fR/8z9OW9mdD1Nlhhpogn5/KbfMqRlqpH48j0ot5hjnb8vjzy2ZF6mp3Vg
nwiwqR9TMARz6qYtwyaNySFGhvus8ib+iT478Co0nTNd7Ctvpg7lb5gDNhu+rDKxgfSQYiX+LDsc
i90btQceIxS0itVu0jJXR74Av6vEkMAhvaCwJXbx9Iv2z8lrkVbn+87pW5as17Qmi+3D/TyQTMGy
Qlbs5Vhm3QW7NEYPjoWJgGR5ZXvObhBA+QP/rtwlW3Dn1uI65TWIZU2vJiykI2rslm5PMHAGsxC5
KrsQvZFzQSQAJCWFvJG9gpgJNkvsw+gwjL8hxboL3cMTNm8e9vn+ps3W59NTO6lkc9bdx1yNjVHo
9D1pmSKYjCM3JgkuMSEkhGaHfJifyiH+e7/9BbafWFEDmI9++OetY9q32wHTfhdnMrJj4e0UJsow
B86C9RjwobKPG7CiLmnQPy4Eay3XoqScSYAgpWwxJD0m6e+TZ239QXE3CxoRpZi7UyrIxoacXJr0
Qg0eEiuz30tuwc38Xlrs5bE+SiiHuAH1E1uLYmWIwLRyecoMuxghBq8LHORW4+fIO7EO0vGTnJJI
ZmBYttmA3mdfkiR+sq3ZErjv6yTZlfRia43WS++lo6Js4vBHqkm1lXWwQEQZvahhcO9zeLfUu8ot
1p7IabZFDuSIdhe+LwnKpWZOgJAaxkiu3SXUHtlhaz0RXFNMccU7j5SPsrwBMCwPOqs7Todlwk6y
/UtotSKeojDmNmIbVTzWQ23Ywui6oCeppJYxUuXwO46kCPqsWk+0Tc5AS1j07hIHHqPzjwIVeTKv
X4nAwJxewWKLjHQKZavmubqsGkk+VDmeUiM/A8bzLHX6nvC2Og7Ze4A3fBmrbK+3v8BZHE5mR7I4
+RwtLs/z+IR82mjf7bTKBlI3uTbho9i0wVFsiwxu36J5rAeA7CyQY947CT2fdNw+LdtiERf2LMzl
r0V3yfZKZgADj7H9PRlOWAUjA3tC+LgVlA5D9skDoFAQ97kdd1BhwZZue8FibhezNS2pP0uqp/hg
8LLaLk6LUP3ezuO3kNMaDBTLQgES6pb57emAjum/2KEyopIoFNASWjQOOf819jvoykGp5AbXKo79
Dbulyiew9c+nXnQJBSfw6kXuOjUXqYXQIDeFpSv5bl0M7YfO9094TxuyhMivkPprSpHG7IVmduTG
K0x6UhgvZ5iEpEy+UCJSJAfxfFeGmXKISjTNY8EiRBTfjSc5k6hGHXwQQLuhxOatnfY5aNAkGAaV
PUQzeZO1/1l73jDC8oXojHQV3t2JFyi781xhcReu2djoRS0NzrR6XrHZ5z20G0rOFLDqggug1lMZ
++VCWfYDHiGPVN7CfbO3cGcm3wTIM6YkAjURm6D6bOkvMwu9IfzwcB9VBphjlSA5ajUiLuS8/ntc
pOhM4CyfxtBFHRNCvPqpatFG+FjB57VegrljpH/MeQqVbFCEE52XZQ7/10bYHcbVFSIXzWo0HSrS
UQn+QFFu1+zDzlNESiJ6tcweazlvYvoe5Lhg/v8VHTqlzIg3y0RPo2hqIkOYAGZdaVUv/kxcVK/J
9HS6z245tZF3SpW2iyXW31J/meyp8QyR3AIWNTGkfbCQHcpdD6+ZkX5R18kU/MxIT7fQ4g072Naz
9fMWWK8l2mG0rtt5aTquwNo2rcnf1+XAnNjN4eYbklXiVK9kuhoJGaEUR4/N3XliW9iMlUfJblSx
7WOP/Kg6NtAXjNrnozRX9DP8v7WfI1U9288smkzbfFFUtFu35Vog+w1MsVr4RQdTr2cZKqZ+q18c
RCLPHufCCvCN9sSQKh3L0KHfQ4/8HU1Vsc26SvntLXvv2O1psO22018Q0nIB8I9ZDioA2Y3FIi0e
+OE2n+TpwWbqZATgMcBwYsxHKxicQcmnIEmQAUtZKbmniUTZINiTfF7gnzpQelXL/dt8uMlrZ4R9
HpGCz0xb0Oq4lVBYmRqTtAbdwwZmRJvsyrw1wnNlnFYOPuTdabMRb9bajMVhrzQcJ+P58jUlLaSc
UziYnw4ZRU1TIEVAb6y53Nqqk9dJ9Nep0HnmnkEWzkFQx/1t2XS8KDxpAHrof6616TDcQYBEhP7y
ycVIt71gFsGf1BgJLf0j5oASS3sUyUsQBIoPCt1FPHKFVXvKFBT1zuTIPpE2oDqJKqtGId3SzLE7
b04XAv6sywgv0W1emMhlT2PEjDzgaOlWIpPd7SeMSQCv2Wgwmrs1U0GP7C1yXqdieLBxmG0TJruS
irLO0zUwK48XPgmsn3GZGWnDrlnWIuCePzGhEVHJRsZ7pci+MorvR8HoqIwRX6KHXL7eu75OymCQ
a4WEGDeBpxk+1d1yGOIsyEs0Vb8QnaeE6LEC1QZ4q0wqEqJm9/bGHwTcDcbFJi+tF336x0o3vleo
WLuWaUbIaFUvx71cc2QpqUUmamWqzlfyYobGECpCTensx9KrY9fp42Vld3sCfRTw67duFEziEWEE
9DXLRlWEYhVZP1xw5NxI5jW5sx1VlvOacwUcytnyNfLMfQC4jqOfJSUoC1220Aahkhja4nAVpIyI
nLhyhGArVXTgx7aQSPdeUQ/Jv6YQMEZ446IpKbdz30S8/nq+S8kD0BwNPO9BG/Rv1SuprZWeFTFM
iE2o3idwrytr9vamnv8TF+DrL1QJhMlAaIzr+eJJ8IW7w32B6uW32XzDdF4mZeHvlC/3O+ETRYOJ
eK4Dy+Y9O0LSTU97Qdaslc2LqXmmLya/3EKyoMTaRXtV2N++UQddWzif4EI9x11NKU3Qmx5ApMzC
F6o/4FunyhJS0X8lwbxcNcDgltYdzp7nHZnzYqYuENG/fXzRLXfIUD97Rv36dOvQxWz8qgnnuS6x
kELShYXqxRTIPaRPe1nIFT9A8gYWzexpKPsHD7nNrA48wG4plaVBFjAXSe2N8iaYMo6l2JBl3239
MzsfH+XF0dN5raMIo+XxrppV9aqtU/Pli82Y1yv8ASYlFeTGR+Pol9sEZBWITON5IVadhhGgPgiE
8ywhhoh6fupKYjToD5bnNXb8EJhkGqoTwZrXKv8AlzXP5S6TGL2/DSeb58jk0v3iwRPol+U5nwn0
6STDfZf17rMVHJKTpagG8kGxU/sOe9YVijkjiACCebGc8qkw5a+MsxnCH5ldCKVmYl576l+ut2wc
m+WHFDn20cjASZJiTppPi8euum3ZXvu6Pk/BWWs73TMIY+MUORCJx9umImaJ5NSZ+rH7zdYk6mLB
aMguyTQLGyhwQgQ/IQgLfPD271NVarKnuTMrvPHXj9biKVWeXmK/L4yxEZWg17wZGiBA7Wl4DZBi
zLRAQUM3r2LV19WzMje5unPB7bOuv3FcwXIc/lM8FB+M9k5bidzhY48218r28cYlVgUc31KSduR3
U8R7N1TnRWCpLHq/tGIhbDj2FwTYWFUdKYwK82iuYKl21kshszn803os6/SXcFbIXbTYZZbeV64u
HqRTZQxzq/6CYQlvP2JFcnWq6ZXiWwsz41MWT3eKgRngJEYuM9Ck6RtO+vk8xPMVqJd+YIv9jrtr
x5G2mpvcNX505CKnyevtBkPY0MUwY25neBpzsdNPjbgyyXcNw5q9cCqFgGiLhqXFMOrWcU4A3ntw
ATz5ymQMEK9+3Zz2lHKN05UQgLJZaD6d3WfEvQ9TgKNgHLpfAs/tOB2ZBUFsFWlwIZQ/19kLvL2d
1JLaL0ZR1zo8RYG8ghHOnMUJjL5VUmJ4MSZVwS854Hu6ohn+q+sX4NWYzZocIDmunpMi57xwbdtw
ccuY6yMbLUbYMQoLU3e8inJRDeh/w1pj9PXMErj0YM6aCOIg80oY+1rAuhIuK6TPhHjKCmodCjlr
h/1mWBGtJFwpOLhZYM8GpmmxifID9Vu9VA1w0/Y8Z1BpqIFRbDA6VbOVmICKRj/aFd9grBlbYHGn
JvoAL9yzTH3WtgISlbD7oee+hplgfaNu87jmF6228m/3GEGsEPY4BNQveuScZ4NAhwISQXSQ3DA+
HTQH78nQJx6VvW7rWX1yh7/luuMEuzu3TI2bt8I6GLIDBeXdIGyeFgwzzmNOrPSF4XdbxKdNMOY7
SQD8VIhiYFUvWIl/ZW6dnC2Y8OmZfxkDDMAeGun7VH/WfJWJ2G+t0guAUpLMv72Pf0KGMW22UJ2n
xf6XnKSenPbweis+Z+WSs3C/JMz8IOg81Ii2ojsO3KKgUISqzyPHEZh+vUBKcjgOzH3+AW5gkYIx
lHSiVu72Re2e5ICr/h0HzVxOwz/weFMYSJM4XxuTVpE3wuEvSmiYFjzhV1BrS5d8TzV0+uUJ5gIX
UHXixvBegTrlx2jSR6VVNAqAjPpzKlL+TytMMr6g9zLKqChinJKTkbpqVzmDEbBB3IxqKHP3imXh
gi6xefSfbUPu85gnHZ34f3UiECfrhDpD02ppnBnNJCFBA+ehQ1X9YR1FtXyUjcLko/f9Wr1sqO16
6EtnQLrfG73Jf+igV5bdkb0CYhWYRk6cSvYlnSsOVYO4X8+uCfj+QpdiF+HFiWRtEScOOfo5nBVO
l1RgMpLfR5StygrfEz+icz31uJYp9TxCNE9ITgSz5amJcqiFw4trUq4iJ6vqsIqxBGf5iJor9EgP
WSoggyq5I3dy+oNVenCRBfYs5IuitcF4BNnIzr62O8iqc+jVlByIJfc3Qv03gvxUDMVEVBAnpMTy
YmBRvWV/HoOCKon1RgoVL2w9qPPcpPBSq/fGyiOKEGY+NZcUm3PpH3Jm+h9tFVRDXEmYxoYrWstC
Ns8KZ+XYLCkcGqVqnu6K6XebxFsGtWDHgf2v5iV0wUCjESV3FQG5I3vzcOMniPhINapIYfyt8YUo
oI4Ki9AeLl6zt/O41bjvtg0mpKUyL2J3xpvEDmFJ9yHDOUfE4ifEICLzDOvgdmqW8p/DLrnbvUU4
H42yaAm2JOld1EYP17NB47cro4qfhJXc5Y5X8hXPxbV2jqXfxZ0KZCnUvfxQE/moD9QSDooBJKs1
6kNHpREr0gmtuG+eJZ+1Ojd90dvPMZMq2joug5yG9v/vqXzRfh1R1R7GrU3oMyMmvBJpwJyFPhhB
7IozNL9BkhUcy9zwVn9ziZPETgjvITRzj/SUB/f0/us6YNOQAjftuQe6AGNafcEitzBJYiVnYXUI
SC5N7dxn+hm5j4TIKTZgaI/ZyEsmIx8FyIfzmgJN+dbwQq8QbI3nZcxSGTwbvKAyJopJUnxMRXk+
OJEAG8oSgnrqH7/Bcq8juUo+bjm6V3vszfiNjJwGo1slq09hSef7GikclA5/+D3XRqkXimikjyHY
AD3YoRwmu0313T2gVDjOF2nbpEFjLoR6DuYaMF2MJ4uEcUCxCEyF3yCmPowBBZsB0rPRhkIJ4SAU
EgbaLM0PuitvUwldCctBad0EG8D7a0S3MhuBhtzB+PrY8u+/IepPx3FMSIQp4UUvaCZgiCJPhFYu
sO8RKZL9f27EBv1thVoJqZn7PzWiufEuxz3oeZVrXcjeXJegR+npWIzXpjGtmoXi7fnr6t3e3JL3
nlNJt6q6imtYPOL82YokAowN5pmXJXd1YFeL1L4I3LZMMPSQFD9Em21PNr2WPvngpXbE1+MqeA7+
VSmlyY0RFVAj6tZQgSMigT7aAz1J18bUi5DTl7mEZJzVqtTyCBYqHU7a2IoO9lC5Y4mvMVg6Xzl+
O3RGFJ/fAskbw/ClVudvbIKbT9rojsyV03vZG2wnzTGL0cuZOmwwvNkm+WBN0Pjwc6bJmo6g1ysD
aeh1T+3DaPj3hkdjawD5gRrREjSP/wSdgH2H+Pm2XR7h4xw8MLGeCcs4ly5iKX5JN2Sn9Kp3tR9G
M1KerpjnRj+9+lUpuyUynKAKMmcNbcQUMg1mwG8QKpmBu6RILC/71+Xk46rD58RFEtTTDAV7PeLu
qE4S8//i158LwhrCzqW8y3SigfmHLib2hk4jz4C7vyisH5/kb7S26/x67JBjX/U8tDFC1hG6hoBg
rLkpuoHKZwekoRic+boUbEtWDNCgS4AXyOKV5kg98HkfrxZzGYY7RoNdkQxnz1HpUXH839lIYRJW
Xh5cP8kCqiugCfYOMlBJnYXkeba8s9qVm5zX97Wc+9QerMqzD4CNftS4ogGWJFODTtAPJZiR4hk8
WxMEoRxAn/L6/oonrt+OdNcrPf55Fz9Ra7aQWgX9Ck7GrNx25xpSFAoE5Tw//hb6VOznIwxf2xjA
Cx6S1TBeNbWtCTxRUPfu49wUO+SEvFD8rF6fO/MGkmvqhmEIU1FPsZPjsCOzbH6wPCB2ATbr8JLd
PqDtPLd2MxqozmbKyzJZpMo+mXB2UlYFRh6joTttyMTyBOTY3u4nKdmznL7MV0dSjXPRFNzxssNJ
h7LqQg77RYKBNrZuFHXdRX6HxRxk2yDMF4rbXl2qrunVNEcf/hEqVGccwCYhMnKcQ8/umEC2dhCz
TN1DunmA5j163YL3B9ezUcdnPTvTqtHKc6WIK00jGIPRrFVPnPHhLCtnPUOxHzYchh0REYik43VF
ClMOY8poxBk/jbb9VK9YZT1w2fMIuOsk1zLrATxHv9NPHK4Yfhs0XnHlyTIe2GAYal7ROS+91YZM
LHTZlPt9Oj+VcMMthPtUNofO3PQ4MNhyvhDQgr3gWnBdv2drs6M++MVWAaTKXorU9HbzEPoYur1g
ILTATmv1MCZ+uC4mJg98CFh8XRFKOLUn65ushD/3nQQuaFzBh46QY06kTUlU0qDCcHzxPzmLOBY1
7dnFg00mHp3GAu3mwkN/XG9AzPg1FGlRxW5cbXloGeeOYiRN8un/aZvf94rZqMh0gINkf6VCcJRH
1gKC1x3CIxK6v5PkPi7WqTFTslvL/z+0sYA2Rd8AVSxV50JnGOBtICAC0hPjX/SWN4LolZiVosiq
Tb321CorxwSLiFlLmwDZb699gEZV2NO7yZ2nevd425dy46hCC73SQQE7snWNBTDJ2OW7uNbt/yXu
MQfn+OEGbv1lgdaOp3hjtdwR91ziZpaa87/N52dcKkGqva7UEll50I/2Yi8HqFx4Pl342xYe3f7b
qGjtDyu10fPBTs9dejWrRFGeswvGDhzIf2RkgbIv1yH909jx6RnRHWiJW6mRwzGXOQKn4nv5fGX5
6W+H37xo3wL6FfAUJfezs507CTbeaCLSMWCH+Qp4mBTmrVsBNzJzCsdMs+YC591g+R6GHZiSdP5x
MrB68XeAI74FNgHhptIP9DGmays7AbwNgJl3feM69T6kUvUKHYthus+ilMFrSdO8B8YV7cgfdP5h
TWqSHgmv33x83olDFkhoxm86SFpyDHPiQGf5bpvBfIYtegyFPhUt5EP0+pFqej581ItVK4C3P3Ax
hjQWatt/nbR/ViHq4q170YdMhlzWkxe7d9o6kpj2J79BQsesw2oBo+y5S7em/mVAisoYiq1SiafD
wWzwGHrEHXlOJ+I3od95oSf2xCzJoPX8FkyYsqeMv2t8ZX35ut/3BS/4viWhY6+QYtfgNGGvOmr1
PklfRO+sYYV8qqU591ur6Ha6ayeOzNSEJwXuXJyBGOTlG5ATDkbSJ3HZ4RP4AfKvF++NbEPl8y2l
V4VIkj/8DP0ppQmDDwfomFNWwJW3g0vtV1IoUYk6qbkEvek/kEgoYgrVupkulFk2+ja+XTrdygtH
B9mE4GfatakEqheRZSvShwgmD6uPTrtepdR0ZdSddrts338Qx+4o6VQsUQdxwxiXpY3/VMRZsR3r
7rw8yL1Hb3QRgJTGBgADmnB1rWdMb1W4WH617md+c2U6jUYiP8tkGweyJSkn6S4sR201QSk6lPIz
BYeAVnc4+jMawZ1zhvrmds78ik44Lf9/bQjTaJ/fX9aTD8bGMdtGc+0io/5BjebcJ2f/O03jVZ3B
uEn+/pH5Qd8j6Bq1mVRyv9FFUGcGP+pzRacIjrdlTuN2OlDCdxgkCdhbLM2lgY7S2SQ+yY+DB7LR
xCnUqydkO1ioVLn+CB3UuUm2WOM3rSjMWq7Ljp7jynrd9mbOK43TL4LOLF2KxFW2dmVWuUs91ktn
SDZRkvq9kVzk9U/yt5QHeaH2nsUDTewNE7NM/7CHr1lMD6xYBzhW2ZnmOM2LRBs6HiHM9EWN0wRz
0CFZqC5hFTk9H7zYYLfyTYxohsYlX9Wit8Dcf1/TIAFIOMqt0DiMd8Z8i8KvVKeU9J5D9sTJZ6IM
EsuUZdExxksaezeWDoq3zyBwQvG2E8FA7Vwbk+GpTrmgD/R1+EVEBGbqQsZddxyHlwqv3am1jH1i
9utkRN+2jbXX6BRDPhIMEMk7SbT42+XYlebSaWtwzdXnwdIxfi3vCloF/quMpfuXh7W6Awry6hXY
xb/eJ2J5nQW9MuHMAoRiHfcB1KwuWh1WRhgsBQ94i+eueQNyJ7AnH1XtGUGhl6NuzQwc39ws9kwP
VtzeJQlgccqQFWc+duEfsWv4GcI432gf7PYufFTmi1U4N4Xkj09rfDmVI0Ntd5CzAEDV7DW+8zLl
6wlswf5400ZZOIcvPymvts5CLc22V7Pu7VGgtEX7EVertIa0/uHhgRSjPzu00dNZkKG9JYXiAngD
J8iuqylXiQDEPndjF+N10objh3x/pX0LMCT71PELzY5NjeEgp1a8J15COiSInozDF0RYCbX1smCT
+CmX+2xNntNnu47EoK2LuMJhdfT61l96+GqgY9HzZfZ1Tr6V/b984eyOneHUg1JVtpA7vv7YnJOM
/bbtmMg2wexm+N6MEIjr+Gn+FmeBl55J/Jm++vP8da2sPw0Zp+do6bGVmQXo+59tno558wSyd1ae
sphK8QXNr+hp+qtLJkF/7G6LX8C8pIOfS/Voi4e8bwZFXZ8ZYyIkK0Dvok9ad5qk4llsNChoBKH3
5u6LBieqAaf9Hodfo9IDMPTPT+Qs7XakaZAdGE1KPzYDTG/VKzSj0goCbXAMtIDyNOvVlfOe7mvy
NjHrnTzR7C/n9QVbAm/2YfEW6DsZ9ewreglfcJOehNum2FVJ6rklmAY+W3K9gLLVqtPdajRKZdT7
jnHZuQr+mvSltLik8PtyktxPqX2p5ovtAucfi7GUglPWACcZhF0EpyaXHls63MU5aENIfP8aQiZb
/F7OpUUmXH7kaJfYSrN3quSHnZlg7qyJAC5idZ/Qm3IOt5aVxsV79gCs2lRwXENGItJ0rz0w5Okw
UaoU7cc/314q5XrLJ/HgzGGn0vb4D4j4c8zp4VSPtxT/OskcElQp+tmaO74xxivzlPFFLby3XVRl
G77tC5GeX79nhubOV1F36o/iq42EyV20DUVA4UbZYY1DZmMoEe9NrJGtjJ3mAU6ziawfF7nK4PXW
qY6ucszVth5wipy6JYhq4YUc1g4Z6ZU+ze7+7DmR9Gt21baaOeSyzaZBmJRfd66hNZzmqQVhy9Us
sSlPuYy0xX2clAatGocKjDG1vZfFSdLE3rIHDkie7RrpAsCB6lpG6MKkVXvjXvJWgX7DiAxPsFsN
FPId/7msJSiMUt929CXM/8iJYVGp47PXQ+SJ0V7XM9ocr9QQUWfxNAZyV2vqH600GE2FGbl/Yzby
QNDR3Cm/8iMGarUS4P2WHi7GDMfr4/vUHdgdfFVe7AziA2VohNt9hGvC61F6dRjpsdAvGw2s+EDK
rfQ7SR7IMRNUO+sCRdv8821j5rMvd8AUqCxcO5clvg4lXwH+NHXq2k8YmnL2V0sV2RLWpg3Lpqvr
XejbMUXFPeGeJ4vyMQ9XVb1ZvwXHKkRxKeAZWZSsb236P4mMC+1l/svVHrt4PBfVtgLoHeoEVEw5
Fu8/f8X+/X5y0djMaDXXPVpnQNMyseSQaqHbyo3NDaCSve6xz+5VQGclHvghlwxF0QItQJcvpmCS
9yKicjG1uEQKSFdPfUuoaIMFRhkh58MIU1rBhiUqEPtpgNyTCet/X2XED9hOjw/DsXXs71dqEHWB
t1M5o5oN29SbiWztBCgRQP0TRT+c43GEOXQ21lbXk6o3htJMm+Gzb7K2pr0ZRcHBZLCejZjmyrno
0xffDHqEgl7d5IqVvuGeRt6ZoML+UNJGfyEPkiGzy31SsDvmptLO0nzmznvsAHMzKcT61CdZlxTJ
yse1YHZO2CyiZbmT2MQhEWSIa5HGmYz36eCCVYcJo1VQS0bB56qjlecCCV/0gQUkE7MEERNmbjXB
xKio+KXMARcC5UmQmi5mVeTIFXW7qP8Cxof7gFwKL8dL+lDeOdn5MgluGCSZWnoDKP4/PgnNQEg6
2I44pRogLbaaNU76lbWxZbEo803on3rBpO2hq19hrt7ddsWsTtzPq3AFA5vb8InbzbwnBAsANmTW
sQ4IxTNvnVzSgX4h45AJZGut9os8Ae5lMzOK4oXiLkvtJmkOH1wnEFK7kmcPivDYIjUsJgJkWyHy
LU1YWpDT3v7GS7qvg82o4RF2WeAOkxUIMn81tajKBlN+LJsh++v/TjnpDULYU92rgFMteQcRjUCl
TLeop2rP//OcklYY8fu+nG7zv7XnDUnRHiApm4oThf27XXMld6DTOpj0YjF+3K3Y6oeqbQZMgdg0
GppW2znHyihMeNTX9sjtV2U4654UcX6scvAIR03J8RC8M/meK93UX5AkxwE8BjSFH663ctwrQYpX
fENbfaF9b0O+R6Aw/VXCUcURzhTjpiDGcVkhRXPdB+pECPI1dQDcZQSmDR813x+kyvCaKQ71ke1V
SREm6Wh80ycWnE+Arj35cdgcF7RAicr9PsZcZXkiv3A7U2oHYZz1Z61orJbsa8ZovQDUQUxtSiys
35zj8gyLt3m/EkqPKITFU+/mNB95IvsGT0SbwbSG/vQlyKDS171zVlPyH6gnDP8phRUTAIdUhHr1
y8T9UoC7t+Hl2Nam15F+vy/t85L9kBMgPYvi/OBs/gHL3oj9awKhX2gYEg/1rNlI4NqFzomOTsbj
ilTel1xVjYipmtRXA67rjwXv89PilsAkUeCX6gArohMfRlpPAiRMtzN3PGQbAl49hhthdLcv35rg
ChzMM5pGfIMBf+PVBBCxz5LCX6RtKy/Xl4ET7Yh/a+oaBEWe2Q5CcP2n3hULbaS+w2QvX7VnLhxe
P7TjDH3JR3IzuY+d9QH814gaZcJYQ3TDcHVa6A0WfzRbnujIKaAE8xWkD7CdI2ljpnmLypTU+Qzn
t+ZiYN3SUtn2Rgo5hNoGHUlXE7EaXKfBP5IAdqbB48zLbCsL/ye7b3zrZZ6gZhxlDvxvRpzkEaxh
PUrvD0zN2N6sVgZWMt4tVz9jxEE/VmTId910WrbSDG8eQILb4L0/JUlNOBURobTbRWxzIB6s4INA
qsC+pg3msjkCtv/iVpqW1uobF4YzEBV8GD8EWIh7D1BkavY4yEjCHeLN9ekoOYGYSavxiqkg2FHo
Sz4PIrTaZqpSYGneiOpteZvZwMjJYyLNsTmhVQKUDJhrrRuij1Z3K0mpuwJMXAQBtuVvmrC+6Kk9
6IQ9xrRWnZObLISV6B4+G1lmSTf2VQE6HbvlAk6m5nj+LBVSOtHoXVFJzU3tRd2ec7WZxTGzpoSP
DY6f5nDsI0D1o/wFzsLN2XtCi6nhp2Pl84Dhjrm6ibnrAPqjCW2Tla0hR4oAkwlp2sm7JHILxViF
Hid7OQ90YTVUWLpx5YFEedxOgUeICfsXmXhRgKM1KXrjftJvJkRtzLv08Wgkxjcb2dvekj/qFRr0
rbmAIs/04Qep1plDtY+fC7ap5l74QDS47x7uGBXX/XZ/F4zX2jP7B6YcRhTiL9G2lXxoEZl704ZN
ayuyLQS9lYTmvVIbUaAVT+Wf4YtWNhKPtKb6iUJmXHoyaDHM4yuMC4qM3EaK6+G+TTN8geyYaTKK
PcnsbbAskRBPv0YHcEDDSQCzvffgYLtGDo2gXwAVE4ILUu/jSBTe0ijMWiE/GMGcNTJTxeajIXj9
AdcTzZWZlIocGbTjnRwq0dymcLGRLuMeOs+hubhhbOas0jsNDiLJxMLQCXWdghIoy6Rl8xuutyP5
FF3vIXAqDXOGDqG6De/Kbc2iSPxQP6EtVJnZZe9GNVDue8GV0MS5FPR2xL+llz5oPvMWjPQpoqtW
E76oKeSf4I2YXfouVoUfZTVE1UWzUtVZP53/a85NXVL0SHnckmksUNhT0yYtCE/wOyKiaLjfzCGC
Ab9hYcRqqS3igfWFEBNCoziM4SLLkgm93KJs0gxasqWGKliMd+RbyeCvUmRFWJr+mXkR/IDnDz88
cYETF4paE7SpOJNTDmTEvV8GKjMuaGiemDivcj7vCB+9RkZKcVbuOHtgxD2bKfp2MZsN5WTvYZG4
/Y2qcBwVDNRgothDQXfc5x+V6qPKdkC4v3WnDsnawxUycY4osoj5nGZUNYjGvIRe89fbVOrvKfng
dnIVBCU8fLo1yOMA6OgjG9grJREr6ts/VpaIaoTH9dvyYnB3TkjVWGxY6NGmNHn9KEhtl6F9QAZS
jtdP9oSRHmkC0BM+KHJFsL4xkpIU1E8XBFss5T//+tt38oFqcTPEGSErHstJTLTJIXUanfhq5awq
CvmFrF21K2SR8ceqdeQ6Qlgjs/gkNOsNP86w6nPFnJe7rd2Ho8LpIOxI2ccWhSBFovL5jBm4mXeA
mn24r8G+515bDnf4Gcz/ZJC4kRWsMbhUdUNk6XvPUD2+XOtSVeCuhLgw2JEKQikk6NvarZ7EyQBr
TH5FtIcCf/YTp2MeTApL21Hjkwiye2olqskwDfKaglfuZlwm4LDsaHT4wRLtowrie4nT35B3CAQe
93mGN+ch2EZ/SI85fhhhlQOA6ZuNKqPsm3jOLeRMhwly7ERr4GUWK9QuK57adiOC+XfLh4K51nOY
6Uqg4eY+HYWuhJ1YRweQh0Zk50dqnvCQIKR3DtZOFfCmDcR9PuItII4Fq/royz9EUm7cN8wLJ1Mp
yMuXJSSsla1y09QZVNYwboy6vujGyY09wpLGD5mEfefUMphFGr01Pm73+qdGN6dW4LR7LAa/26wN
Vgd3dxHxyIjpgMU2tKflvLpTbCvllZ6vOmpxz71qYwK02tp6aa74QHUVPf0uBlk8gV4H7rCpZC38
DvwXPSsix0z2zuUEPFiunV551OrrY5/nPPYN51KMATuTaFap7/CiNkD9iu7/GeR8VgMwjFmc3fo9
rWOriPWiIA5qmcZsFoV0LubqBvle7jSLUS5jwKtn2njiTn9/ovxVSSVx4/9+Osl2GCTnbdSanvGK
1IatyosfRtBgvIMLwJP0E6Cgo8A//QajC1T9464GZn0P/URvrGm56KQfbXr5ImyQkHxNnsgLmPLn
42YzlSoonSZNUD6zjOEslEA8ACYiOMGbFVHWgvtn3u5w0oZ0MmE2V41gwvKz4ta32EfLIS32+Erj
6hocBLR0JeMoJPOvAH0aTwQilVkRncsYM58MrCwb5N7cqNmEGpkBNDewj1FuvekniLnEoSU+v9bs
PbcxWnfxTMBIrX+dL1LRiITqDnOSFoVKLuO5sr7W/470DishimfYBWk2MvxbWoBVAMjn7cR95n3B
bZGxhRJSGNy56j8bdcgneheYJgQqkfY8DV3sa6FbfPN61XwHRHZGJBiFKnA6zXS8uDqs0hBJ68ib
6EXOfE+eEa5BJifcGWZ32pb3qQ9SFL8yARxHKpuNyWyAMWAUMXw4Vqpjl5IqSBJa21FEHMdjEbOH
EbhqqJCYHgVQA13ZI3duMdeYud1hKu+cHgdc+JxcKXJ3Bid0smEtf7xhWZSjXQPFGBlwtdo1CmrN
VizaCr8gsdI4n1y9B5jTj9KaHrkZ1Hua05VgDSaKIgKm9kIv/qAFAj9UupSsWR4pEAlErQD2OKUK
ra5phlp+R5MSsl1j2fXeWtDJ+pNZW7oEAgQXZexjgmmNMzxT/6+rVkHg6L2F19PYOJWzsRut3WSb
rIoAql55YGDrb62Ia5j2D3CHnruIQ7El2JtXYFVG65cEXA8s4ReNhT6yb8e+VOTEKzNXxW61XecN
YrXQxebd0Q0WAn9jc9RDEpJpaX1J7jVTE+KEVEN6YVJXQjhaGEaCM+4QqWl/XmrpiM33bcOeJPVX
1CIoOZFI25twQMcKBgSZqBZvrj4AC+TAqXbl7o6lBEEB7a3e5FjfO/AgUkgelrwVvUQXNpQdgy+I
UXAusS73NydNXLEAroKQg/0VcFkwBZjFMMLbvaTy9YEIPqO8YVh+3KW30euKFgpDPnan5kycNiZn
RefNPEtVzmvGXs8WxTfcLY3xnk+cJ6IlPJLjgbLpdEd7AyCFq6DQ8Gcy8oKnv2YHaP/hDg+6x3yh
9uG7Pd95pRi6AbLm/u0dm7IribruB2oePOQfPHwBn3BxXYG9kIQVNWHRr+acMm6Wspo1gn9QSFkj
zOKk0/rZbKDUoA/8VjfnfeAeMiWOqRQSqGC2+qrDulZdTSZvABaspijsH9OaCn2SQaA+xpwv7NbF
vJ/AI+9pr1aRuql3AixA7DXRYWJ3C84ZCkBebHVmvfoqu24V9lPBRLMg8Mr3OvEHKnSdpfs5lnAm
+Got5IR7Fds6f4k0SJIDKHD3pjYrQv2XUylwgqs8+eBilIm0VxqooMvCYvGe2gYp4nj8LpB5Sb3T
4XArSNEp5AGY5dADNyqyVRmJsBdhGKXDirMwyxdtlyN6wqfei1/29XHq45pdKUpIEpuee57i4uOJ
4eBL5wvwMtvKNox09zzfdrKr+0DTCPdB8WfYt10fG+442X0nw3ECcT+NBkFYbkcSTVYpT3z8LARd
xI5Bp4QAcXHfZFdueQtLpy45zWOv02d82PFcPXpiVlDFxqOxTb1ylj/mcUv1PBM4tMrbPkR0O3oq
sw7XWDgQgL2WhQJeBRGWmNfCH0TT1NPBUm4jjUreFMUhQrF8EZQ4O7hWHaeBzPhZD2YVX++CaS6z
JTyZ9QW0Qv3AzgEt/UO7db/KesdqP5Aki1T8AcLUXvIQdjtngbDP1knV9zpD+B5+1ws3bagzWnkf
agU5oMejmElUxwEx3L+lwo2qTr7xcepFH7ss+815s3I0mnlrQy8bKE1tISN1TSE9hnhZa+CM+lCO
aIRSg6K+IqgpaLotn9TMM+Ngc5HPtrdV+QT5QE4R9rKIsu3RtN+Lyr7NYai9URhbwY3IyZgu9KoP
1Z9FqtVodYyN/cGzI7EVSqiAwTPtaI+f3Tx3Cb5mLQeZRrYs3s/1Awv02hQyqQblOPTKSFc8IIEY
hXV1JA10WdsPZB6bV469zSjRgy2vBAFw5b4tFRZ1SXhVR+CPW4aSq9wmctbUE7r0dRNicd8VZD/1
LwcLNlYDlLsblM7QZbu2HeGA9Iozs9Dxv+RCCyPLTjlkPXkIOAKY4Q0e1FjNUY1xZBNAWWphNsgW
TXQdU31K20KpP6ds++eTi50hycrREV2eris6M8R1l4qKzCHDzIlYmiHr2UQad6NxLY92+cHSwfKM
rSKRgPAeR1qhcAKPk3+Z1cOBkxbId1Pqt7WXLjx+imqO/IbvH+CDDLa/g6hUx7sjQSkxKp8eW0nS
Ne0Xw8fN0PpbHzB2aR2J26AL/0ya5nVS+/RDeYVaa8VhCgw/UdTeKEHCU6sAvjhr4bDOHF6x9MAN
yyXXGHpWkBmRMKpz1yadAhQtlHqI05VXVnJ1cUBTXIJq3wemH7HDtHzqGg/HAUN4LFCAep8+dyuS
iJVfabqtBYhYp+H2hqiXnhsD22riLjrWtR37YZ8sXtSD0mmAkhcVQewdDWoYkdk+0MI8Bi9knqyP
T++jpsRYGrTBghycQMOrisjgjIQ/YjatGO5zGgjwfTtM3R11N7i8CgX6cMBv/ISXEIR9q4odTSu6
FRkkvjb4w4UK3J4FhRgFVYMC4w9FBBIy5dDInjBIwZ1pAde1npejfF7ne/0pOOxi8mQjlirq48XV
fI7K35IsG/qMdWBkhMWorsgNqcQhQ0VjPi4vQ5n5pFuMu1L5LqC/rjov/AbDftud0iSgUTSHvrQ5
tFdqFQxftMIhTzmaX0boJwSAYL1fwv51hGV9XGnD9O0d0Bhh9V2fOy96QtslMOtR1YhapiaBykdB
XGsAMt9hYDWkBUZ+RiffXlNU9CHlQ/AGnIg3HUIcTah0Vj6Lp0PfI+x9OkYyGHM48/1SWW77ii9e
N/0IKqBTIYLLBaqzXHe+djrixiaVdXMYPYsxpJ/hLm2aN+5KogCu8OT8qJJnP+iJmRnvd2GTBrDf
oMzOG7FGa0GxyN8QRdGIe3jYgYV6m2MTBc2bP7IzECYLam5B4u9lGCdIhYPcYk+JI8AYUS/f1HJd
38RGp9ft2PZ1S0brM0/HCPvqKxK3Vrmi9dgwgieXBqub3p9kU+72Y98QcotXVDrSM7BNDT7vVtEq
cK2IwJsQKp79DQ6zv1Ap62avDYspC930k9OmbGGuAn/hePuVON/FHZdfb8a3rDQ/BUVG/tWwPfei
JK5AqvRl8P2abJu+Dok6RZuftlVhe36KlEWCl+670NiT8lj/Yv2l+620jCSli/uO5UlgPCBPb9jB
VlQrtjgFjuZitQ+9sX3002Yix62WXQiog0DgLce+3KN007AB6nEFGN7F97gNKhySgPOqBXFGK3mQ
9bzZWqYFviBtFuIr5pOTqMlaglXKv970BGHxoeKhHho7I6zdd8W797k7kkPwR7t5j3tbeE5MMn37
6FO/MS3K6e/Sq+Wc63qZ8sCH1UBV51KzNyNXGYlrrAAz9dlBx7dl5ifFMSqMR8+7zJxn01+tzYDp
5ELF1gQXT59Wo2VcJh1g4bYnVsoeR0RYT5TuJXuNxSCahSvmgY9uM0e6ZGP+lUidpGZY8STBQYG2
sF/ZDzOTt3MU/lHJvuKmLHOmb+TMMDzMz7sPRTChRFpl2/n1yGFesW2fVRrk1Gp08vHEOZcLOyb6
9S05ti4KXsJEBrmMlgtNpKaO36Os5JdLNAonfwcU3PKA5G/7Cue8a46oTNZ24SnBR/J465wlVCmh
IVw9uQ2ZuiH2u/z5+AMGtDNG/l1v0jQkNPVk0zBoMpk+/eHddDJluynyp+e908A4B3Zwzy7IaZLo
yn9GdC0KVZhbvmoGEoboxcyJN4Vr8zcgPFF6zQ3nhraDVgIPP62aCYtLHhgHoF2FjrRE8Mue57fd
z/mA6ymvhNgbew+4SRjslzAsDdpitcP9cf/fuB0Bu1WByrCyIQu6ZhfjlfyofYoEajz9vPWQyboY
vccBCTBFbRfwihVBUIbHGTiUhlYhfsC8EDfEkJGLfu69QeqPwX1cuXEwE29/hIJnnIjtV9r0fbH2
U0M0FyxEvXtY9Z96lKbUSvQSfT3MYz/tJREyq0U4P5ykAq6Fy2BOgAQi76jCuVH6ULd42rmsbiLK
YQbkin5LPAkoclaRAjEZbl0TktRPJoafsKCOAnoj3LA/MMH7Kny9LO6pBPkFHCl6g0wRifjwQ9Nd
GIroqaDtBZjL+2QjXhjHuCHbK5aHddTY6lO602NOkHUeqQkW8qHUjA1lersZPmD1sfFTSAh48V96
JpE4PDHDbv/YNUXOohaFrSWdAuGqrrMiXpcz1gNYUbJp0IPSa+CVLhYUdU/VuEZPOssfy1p1Dudb
/0lqIuu7m+ixoTeNqtdSidi62xPIVoUfGxfMKZFbt3TANmTk+0x4m0MEm07KzIi3dHxd6rlBS5m6
9mvbVr2w7iJOTeMy2YmPO1YoK3yPy/bvXK/MPtCFiEknvjE9sBLF2vG35P9oT2Qhrkx7ar4vsAnF
2d+1uEqyAJomA1VpT9XBkvH2CUI9JZgprDRz/CVo2SoVCChxJuh9n09RQYkDghKGQuYx3KkLz4SP
/lD0erLCrjonTu0SIutYq7GEPD8WZOAlN8p76L7QkyGZeg/Rzj2Eqt6LCv36BcABO1YUgU2F2GJL
0I3e23FCveMUADYazGDB6ogXMGIGDclKtby2hlvYAnkCnCXjoCzlq+bRtmncaTDMvKNF78hKIqsx
M02YrWRaQib5NIUbm70slPDfN+gUrAi4f6lEojsaJCWeQVPbXE3ovCs/RAIkUP4smV16ayYXSJix
2qX2hVcAJOx9HGkYXK9xYTKm6wkDzIp4Lbr8xXVBz/F+9m0oRKBwQChP+BLzdnizOtD745W22kSx
g32Ho+eLbH1zMX3uO786+Q9eitHqymS9Jn3Z/jzN976L+u7J+z0GdM89lYGFAodAFtjxYey7qrz8
d7oFK9ZDlwo40Kr/tcugQZWDgtnMaFYcHShq2yHp0CRbJpmrEj1GAxRcB/rg55LbwLbYh/n63ME4
TF4CBhl24qWSBXvKI52BYyQcrd8lFrDtclu8ambdHcbPcNzIu8UeEhnQ7uNwjFTsH1hdJMtDiwnw
MKnb+19tZGMcHuk2fJ7RYMzGGEwf656uRoOEJFlXSnjMV/CHKP0zWfzGqS8g7FEj/TbnIxDMQ7Jr
b5SJqguc0ofJJySqGApHGCqaLdmtv9ZysOkC/dBQxieubrUVSSBeJyfIXV3ZKIVyajUt4nDPaGsP
8K83hFf1LImtcIuSa8WX5GYtQCZRhCZyxxessbEezYXg6znL97lM6+jS4tNS9cyy0lI8xSn/rK6h
iaO7rRuQPkvk9GwYjGDsfpbsvQM6nxHKwgAb8vKr3fiYxHWgl+ll+0fBf+xtdZ5OBnwIhc5O8Z+G
ophByLPkv0a1MyvCrTIcvoxPraUZgLtT46oTCwhVHxSlkUa/WpEV1gR38lPbVds+a8Wb9ujc9oHm
Ssx4qU7zVvZBvKKvuZG3nsCnPVuhcvoUPSi7ZpN4x8foUihkpiHyTIcAZllILkkYgYFSJ7MoDnws
F405CgRRjqM6CJZ+GVQvhtUZKjUPL0Vf+OC7H+8HIfauYIxT/kWCPj8joma3hg73gwHS0DYtloio
Ox21c7eZ0p7uVqkTtCG5PWkXTEsyuZ7mVRG8AwFTfBiRMezVONOHUEhThPTUizuJC/HxxwSAL3+c
osUpqqBpyPHyP+aAoEfKBXlv/opDRFNH4Mk6ubjCpXjxSadfZgtOg8sZWJGwt64tQcxTZ4aF/Tqf
1WETmsekjCvzIlgdPmDof4KpulHjoWvhDPLkqsnkufGc67hccLUnrpFuyWM0vtIuyv53PV8Nd2PX
FHlsGZoEZ+Lu7SHd/1/3CR7u4b3Au+rCp27BNK4ESUwd8O57fLM+K22cO/Tzu4NsxSEsuzEuT2rs
mZDiWYIfQbc0KDxmYMjLJFg8sWfGd8ftkS1L/HtOss/Ga7nVOYQhM7nQeVE1GUtI0W+E7SFdsQ0U
OOw1DGegOidKuZjBrh8WZF0fOdB9pEnI73F5bNE4CsLpZlCsSLFa4uT5Kh2iRB1GJQDLFLLFlc7M
dQAfqcgBk2/CV7KtK2mKrg5e0dKU/pABzM4C5/inyTM7fHQIbjoz1WDIBasVZ8eKde2+uyuk1bJR
G9GrWV+qJe2+H50uLqS1JGcAxanAlnI4UBuRJUXvDS1QUY49V2Zawjs5aPSXWe5kEk73EPa+Y1NE
IhqWhucKsjJ9MWsSA3axVrIJWJbnfgvSz9r2YiU28CVwxKfDLbcjKG+z91WWSUVHDK07kjdaTNSG
Pmkxzyd58imPftQmCnxT1Q01wX9BebThJwFbjKtUqt57ulGvbn58c0m+LzZTTkoYzizq3USrK6bk
7wniuOP2faTco8GMe+15XAfTlPGbHCqtvR0gnU/Mj+dcQtnUGkvzcT5QlhpCkElZFO+heikKlJr5
N2LCmj2R0oZPP/dlCq4t21xeioYLt/IrfqS0/il8mWUhg2ez+G6dvU3+2NtyLzsJxUYCm/u9hQH5
jxH3HMbInFfqa5mQ7KDiHe4NHKW4SrxKgrozB6ifm7tuziskVuXBUnGZuLmPNZyrB8WaWppmaPzH
aC4CVRRM1RZwZWmAJ+pSuL/ulWRB6Cc2q8wly21ZH7uZ5pi14skqOrqhskJ4QRhzIVfvmdY/W5aZ
PFWPcwHycEx5GJLu8aJbmkp6Hcwf2ogbveta5UQsZREzvgzxznhAqZOM8w1/qqcVY6fG4Y4DKLII
BpbQKooXvEAQnNXgFYjamrtbr1v0yrTF1T+ufLpdm2GNrBXj8ExABHteEv/1sZzbWNO9O+1wALcu
C1D2218MhYEoXXlNH0oUMDbLmsxi3c1yNUS4GoEYpVKKwdY9XhK1oU0eIe30If3LV8sRxeIIPa5r
rYAm93FSqTPvGf/0Bik43GZVJFdy/KBWQ1HqrO5R7n4XDvPhJ13B9mTLdyoa3EK6V9L1aaJxRJPc
NbBY0pF9/XN8KHiUZdg9BtXxg2Mmvxpt1+tZiY/8zoYPlM2AbSqAFir6kiCEuhatlGRgpgCPdOyv
J5OGeErX/dviWtSNmiuq4YaW/KZuT3UPMBU/6PQtUeFzZBFImgjzpjNtvfoWEtZOKHAUn2lNukCE
Ovb/NZdicW94NP0SyTWS7IFA+xVT0gDWu6OKDXncd3jWCV9hhm3EFJ4bAnEKww7zylypRftuDdX9
ZRJ/i6babqIUSbcRT9a5Hgc1NY8OYOSMq1dYfNq5RmnYNdYJ/wsFidDq3X67/1mzLtiW7Gprg/o+
Kn3luC1AuaSQaJm+rvaMHZjAuEinGcuF/kCDJeUDvkMQDKe/mWCArGK/birzxmsZH0U6ruzQFbir
9Ol2wRgssmdnL+TMs4esHMY0VptH+PvDhsEYhpLWpbWAlHQ/j8C8Zelmz5QNxuWSNYGUjwjV9lV2
RzQuauOIPQrukhaNEy8cRhR9oBzK47IWz0wWXA77CZPndO1jmYjf0EgA+juTXgUMAItdRkLXzhgs
XOgGm4lXBRSQiXgH3MBKS6QejyE1ZFiK6iMnl/9xNX3IofoS14O+6FeHp/B2i9a7IdMM9Th+olGV
KGuzh+yyHfTFmWYMCMSnkMGiUletGPKF4tFmqWH66pyxCa9WtUIiCQb24evqVUhwcbnI5/u6P0YM
4JAnyegJMvRcG18HyWznDiYyTthAANwjDvbNKBFY+SovjBMX7MCSHKqxduURfsBFK7bhIlvjBn7x
Tl8MM3b6/hE6WpVL0vi/2YRcVKHfGIapO+RSnqGUZkGTrMyNeczuTPoyQVddO8ad3w2+euIKy7lz
XVkwfalbK+36sZ+c3bgf+rEq/FouZuGk+V74p8Vsl8gdhO0FTFaUtVhrz03fAbJajdQ2gxnNT6Mt
zj/NmkiZvct2fRa4+REAjavUc3IzcBfbtR27w6zXo/1UcO7saby7fvZP/qo3dy+/bmOVjNGqIK7d
bxlz4aQhlrn3U4tFKUcIn1NE6KAWeCnVOPrspRaJnO+g/tO+HS06iAGGIcfgsxdQwH2/osLMyC0m
Jb9MfEJNokuuL8O+voP7jar8Xna5PDZUjEAXoX2nDOhAExKLZ5APo/zI2+b6PEdRRvxt/pO5Ccoq
mHpouKUc3aOzVozOUUmWIkkJ3RaqwMjuAoHrsn7Lnw3ihlRooav73gtZlkqtiCZZBfSpILz2O9+C
6E50g8mxybUtbs7QtGDh1Q1ul5ByBsOC6Aw+5hRw32LNQ8dPPhjqpELy3oXS/5MFs3tFMt4qhk64
P3bCyEx6aVfu+esLFc4L/nGuvKhk5qqEts1PY+4iY8Tzc2KJUJcdXcW1RG/18l8kQzMpOngBCy5z
X9/nFFzHmMPS2lbl5MfMM/TyQDKS4SIReL3RwERMffkPFqv7VlNyGDX8BkN8mAkej3WDtGxpWlLQ
04RJrA0/ZoYm+nODzsACKtWNywi3ZLuH0DUKn2Jdf0fSICs2JhhA0Mpyxrg/2SLnCdEnRLEzV5B3
WENba29Gv03V7DYr7Cw2fe/JtwSw09J7J0yi9NWH/qOXwFL5N5PRhRwRPniq/IlUQyFl2UYw4kN/
Nl2vvXp+klA4GIP9xv/IxJLVJd3burcqAxCJ/FKSgG4DA8FVvJumyY+83PNCq2kDN00z606ZFjiD
OO34zzVCIdcVJNy6aAAXGAPq5ptbhIgSnvpzhCdJ8dX1tyM0Y4+3v+FW19tomiA2CDatxNIyV6dH
DKjS+GZi/Ayg7lgoP8IhdTCUsb9b4F+d0mbaWoEzy7KJpSRgpjUPsp+0ZYfZwKgw2nsNR7N04L5e
Lx/x5uaDTW/Gy7dMZRjMeeoX8RMXoiNP5qZVU8V8nKbh/+6qqFob9Uu6/iF15UzVMvrixqU0So9S
TkYdJrLsSAoSpL5UrFrac78YD5CXxPuCO1jqi4VMiNTFjlyZH6AzsAfkK9pAOqb0+ErM1ATJf6ou
jZupjNGy6oKaEmscQPsdyT1EF9lbzjuF+dvyatlC7DLano128JmUASOGFzrB8b+5cv0a66yoCWtT
/1IYjY979lDzwFklw0BJThJVIgzOVCQW9bj0ygQndkRjbEvddNzLm+F3+owq9wYubBv2qrVNElVu
fCjrTtsEbG+kEEbNVyunqeRxyqdcxw8CgDTqtnDPzZjPH0p7eBcbrLaswYlQqGw0kudYBKta2Rly
po7mu3Br35QO+pB8hAA5ou9D0Kiimu0oMLhSj1bTBP0Nnmji8DI3YeIPNGKrxZxKwZOpmZ56yLeJ
l93OdFsxAJQv872nn8ruxAJhIwQnBttxqnlSMMZKLhdLWAEj/xzcezT6yr5ML2xfh0nyZQxut83D
oHjEzdAdFUSRFRu0zchHrszvbip/eU0Nw5R++YRzPFp93PuiMHQlMJKZFgx6W6ZZoFGd0ZqAFST+
F3AY19jayGvkbsUIvdZN0TmTnpXUG3yblpuvg7TUciE1pEA6Kfo8j7ZcuqHL1ZSqCbqwJpHK28VT
Lh3E8RHTGswgq8l2/Y19TghuVtCcE8zROWMDDdThL8OkOq86qmACnjRDLJ7OIStgde7OL932mCxW
Qu5Osx4qMxd0pmvb93gw/nYpzlAxzzRb/kwLlrYkxxMDT9qq5NmyyDn4U48uQZ2S6TduEyumebmt
VlxkX642KQJ0R7MWZTAcggI+Go/4dmSFFQLGgnPFvyGQI3CygRuWODLMJR2bMyb0zNWZq5yWj+Y1
8Bk5aoZfadWeRzq5BxWXplazd3dp7/Xljv2on3ixhXA71Hw2lZw4pY/3wmy/TcpsQAELFH1R93zF
B1cL9jD4nDEH0qhXRz7TF6R3Y4JAplmoiCWOFszeZqUkdrT0wPYQhV3tXkhBS+2UT7LUBJPTCwRS
t/lmzeULHNyafIJLRkFL070IjyK1c9pLyWpb8QrJNseTIxDvA+RxEyHaSlAqj8YMYeOiaia7f2xf
+HEWrFo0ugj3nbl+CCjlYJMbVA5a3JNhdZE1DL/PiEmThwQLAdua73VdEFGEkIUJlqILJh+qTwbR
Sfrnz730yJGQiPXFAt3zcFtCPD5ZcSmC0UOn187koBHdEg7SPJxZChr8GYYCiMvv7UevONv0vcOZ
WXOwFuSgfF6l9JFdAHf1QjxS1cP+fUQ44W3vxBEHbFNpGW07C8UsvT0ROns1BtgQphHqw5SsDRtc
6jivFqKztFmuULOv4m8BrLiYJVF1Ql1DEOEXabF3ADD2AGrY7zW3ovEr28lT9i6iGJRxPR98PSLY
XhrGGbv8GUL+/Y7KIZZ/SALCq22tcG3adzMt+dCNA4Rds/8FFbnl00e6dxmbm11O7aalD57XjV6p
WER3JNe3WN1aamR6Xy9tNeF2+ssZRhO+8zJgklI2C6N1OhpAS7QoHTNjyVvE6cKYqKchRYE5wkjj
nWDyffKZ+TzDkCMmcKSLXUo4WflQE06K02wMiLyijuVfcTssv8YQPM0ji/StdiD9+9wAxBR5OgVB
sFHLh5IpeQAEbfxJrtSATCFasGctW3bmnsvllLIdL8FhrGnBJwPtAD/TEVcfw/EL1aCVUVD+z7uk
LA8bHP+1ueSQmAhHV6MDbSjA+62Zi7/3Q95Jg6pmQZ6QPTgNAQVvhRXu2C/kDcb5zHRx8XbSfplT
TOxbAHZv5ORgRayR8MNzeiJ2RbRA3B8CV1hJpdFDfmPGU2Vnl7SvQcIvjNDGCKd6VRb/tA4bU/dP
SyXW+VUHbk4A5T8YpUVi95VV1ynPpB3wvsaiWWAFggmmexl3DpbPwUO+d5Lu6dDQ9eIUhYjeUnOx
0hWnjtoE35wbyOHfDiMgi+j+UfsNAQcnC042EiyQa48lMh9lS0+u2bEzB8215Ow1EpGcN5j6UssX
FWFV06f9s3/4xztXOiG/9i6QSjBhuS5c30Y0YZrv5zY/FdHPd/7QvJc7wlErkVUvdJ21cB1OaK3Z
mzwdUIKsI+R6RNpmb1K2HeKYL3hxUMBE+nysJQI80QxUdbI8ZVKCJS3lbN8qgi/AzsJPm/aMLKf/
GpaaaDfmHM9imxC7Y6MvlSWNS9dlyx920G6wAN/5J8zJOJSMGcAF5rpH/mT7bDQtkpOkF+HkufGW
0FH186KJlo2p69QyKDjlv094WygP8SjKdTjOPEEkHSqnjXZPw//tvTni0b5KzesbE75UllRqFUtz
rcH1txwwbpvSIq+1CIx6RSe33Kqmx6QKnCNLm5XTzl8w2AtjNQqdeGZJq4oscBKIbqF7h4A/k1Tv
1fgrjB9WDoIlfW97He1ielTC58WLH/fOMpBrWmlO/m00wD4Guq6ZpCum91OSjYcKhERfPeFvpu3l
SgaxsNgeTMwP/YIHv8Fz2AbNugYplikao0oGiT+2G41K3EtONrW8Obfvj/HC2OJujbszZOUBnnWt
bgAd9iw1xdjJORUo9Z6/giJMiB+GY2IAJefj0Ip8pkZppuE8kRnfq+XgQDulugkxciSmSgXZsvJl
jleOaSZv92cJKmqSyIfmvCy9v7pf6NZfUTzzhwnVsWTtGuXkZ0+sxc86n+bzR23XlmtxSBwW0qtb
hnpBIIW0jgf8VCDFIsYW/k0szs28uB0Xyfk0mpmEyw9axNtPdLPUyRlveI45Ohlt2TRGIF/uMMNv
to+o8M3+i2EqZI8MXO46C381RhgtD4IZcC2i8kmiEPLPBRfzc3YGI2DBaUqUKihN3S4LZwqUj5je
qQdWolnxQ07cG21GY3xC/Toi+yrmOFmUAEQc/pghZucG7EkQE2KdgQlGYARO1kkPLwCyxW3WgX3S
cBUe85nJoRtJ5vbOWkhYsIsxfuGo0QquQj4Fb1wslqfFXihZYHMShSaLXCvSp5x7TSczf+DAC9mD
SH58UpXgZjQ8J4t5yVF7aeX1oHmvYzP7ADL6DIoImreTd8z6Izwfqac+r/SzIs4aum+p6IIlQfKG
XypVYIwyf9lzRgtn1MQ+92wp8WUV4WOHa+UioIDLryQlkCTl7rvxMmvH0fc6t9+l8ddszMp+RhQm
q7LnlMX11JBboa7EMwkgE4h0PXqKt17m5d7uRREjlM6VM0to6ODHIiJ9uvqQl+LcRBeXSJbK3tHG
N5y/94s5ks/E/WMF+10hqPW6Y8ApbYUkH+6HTgA+S7sYMIGywayWyo4bQ6TQSTY0pRIjNAj87Ljx
snyq1lVkALPyOqdpmbTxcgYzvY19FxMvBwis4fEZSVhOmKWNQd7uU8ONX5xu3VFDVqLD9ozqJU9X
VdAQJZKCMJ411NaOUwuJSk+MiqSy1RfhfJGEohhLaIMuMNWoGTG6vxN4N9i0R62E4Q0BajgHSQhO
mXSqarwDf6C3feoxuiovscJc0lLL0FSa9SJ75okld2kLiM15Q4/2GalsE6aIzJHbMyl2dIk93Qje
I9K8atWi1VgPCJemCXabWgYb2X8nBB/IIc1qsKG6wtHIbTJw1HDNTL/oMpDwceqqq5WApjFUR9c+
DQ3jUrYMkx8m90Z7Qqz1u/AAssW9Poasy9TMpuIkxPItYHuaozipF8osSvE4GTmHBKOj7yhoGDUt
3DFk1mPjr4Kfxyt0JF57Uqmug3/Lq6NVm6r6UeY3R0RfQkxBFGUztqa2Ox30h+PaU5G2B8GXz4M2
23mwBlkoi12oQu4H0EvJWsBPDuWTqaVaKa2X3BvX98aog1uJ6XAPwnqgffAa48HBtaV9aYfa3UJM
jtre5m5Lx/FIeCtfVRjwkgUEebvFz8muTQyLvwNPN2wvl1Oq9LvE0/UxypGjsSqdzIAivGeUI4LK
t1Hb1rjI8cvq7jQ3/N14PFE5+5hG8ZlxzntzaR8/DP0BS1GcEHHbkev7bNYU7fUNEUPTHqNPXCww
0W8OzjJFMqwPfe96kNyQTpbH15bcD7NBS+TbzPw/lSoYVLsV78ZPuXoTMxIFwlXmtjRlimfWz7MO
w5CScSAijqe2Hgv4HrUzFO69WAX2LDJfW3kslLvIB+CzdK3Lh73We6z1prO6yvhlSHuRztGR+003
hRj3pvLDE4+/gSaoG6ji8nMuAGQ9qLzvGrb9c/3Gd37DBF1T7QzJfdqL38vYSx4rvgaXMDC7l1II
J23hBKRMy4Y1tbAIdJHq4o/qvE3h5vjois+vi4F1CrTPNW/DDWEiFSScMvwFMCHRXUPnz/hzacaZ
m+1LPNsH+vyfZsk+pV1TMl7il9yDLsmTTdTb4B1vPicxJcwU2CczNeNKe5q/ZDKWPwDBJpPceXjP
g5kN7G3H4Q9syNGH+tRClovO7ENIaQmwimZCwwOQBOdJ8ze6g8SS/cT4l8ATMmhDYURokX6/n2BC
adxARHjKnscEoxYma1q0m34evzGGEjN0q6iJwT6Blk0JguDTZZCImwJeXz2TVYu0ntRYMmVQIBkW
d1WEb9Glb9KukfYlt8hsMzD9m7AfHmSC1qhYGdUe5H/nMLDEMnywMmbTRgH6/7bpZYpNwsqqaG/b
TqPyE7SGmwrfHwsvRD0heSFB8l6Thflt1+i3So5BQCLdvWgE1nTROssmy8NNdsmlGT7JAxebzg3n
1Me1odu1GowPLcng96QCohLAdwtjIwbWyQRDzcW9NDKn/aHMKXYN+z9fAuFvibJERr16zJwLs7jz
UOeTU+MuO0aMMJOzOJCJw74cPrpGtc/KCsxB9awJECtVLnJU7fUQcMBVjjFvZs/C7Eyzdb7JBwGy
+BbnELUBLLXtE4kZ/J0TABQ7VK8Iwx67oKVAyj0D801gTS8wzva1N074n9/Sjm0FeGXCXQqbimC1
z4+jo7KGRWnboxPwLVckLjDnuFANM+Tli3XHiBHOAMNYSnx+IN9GWsbYQfXaL7599Zvaqbz8EWBi
yQT4zKRJi8YhauFyNLLI4P10awEG/XwcoqTMrGxdavL0SmlPHVSa0oJb7uabV8/EX3ns4PAe+hiU
n2kgz8XUS2B0O6ewLWzjbsmH+Wl5Bhl02EI1qn+r4pYrlcbRrsrZrtWv2ZxXYz2de2E9wtmclXFP
aEbRDkalivx9XTPV+SEoyM2xC7Ezj4Ir6aeP1UaZQtN4EygF5svkBftY9hfLAhoe/sNsfNFR1lEe
+9bkzC7g0oKlf9qGbWG6H25nZmKSTd+T7xDrsJIhhEPrX9tki8goQi3ici/63YQfxStWiI0bjLQj
1IyS4abVUaJ2dlAxrq3250HkFpzQhWyi9xG7+NBPfHjp5Sjmr0DzNo7GOczbQTVsbIjIQ7xYMz4B
J21c8Y1REQgAzhplIWm/64WeXBY82LdO24osp8uyF3kxI3P1+dab2UxkU6aZIqc0AgXgNVEmdtIV
wPznvRcN+oxc9s6mAb4sT1iKS9A6HEvUBdytvCym/S+Ee0WdlweyYGosy8QSk4zfpjeikti0I405
w5L8RbhbIbhbKj/WFY1alnvjlSF/ZDythNP+a/AQuVKEmhRSIdoDkZ3XRi+EIshjVTezVG630qLL
w3zp4xmCiaThTqa7dpvuBX/Vq1QQF4hrvYOXcdMtBp1J8q23WtjkJwZA2jhoBC8wGBDas51np1Xw
gv9+FulKddKc1WaMZgQs8bGlf6L2fmN4UhyHvxR+v4ZIZaltSb8gdOVIDJahA6XJ32zbdKWVBhAG
2Rse0bl4tfVw2HP62FOYIr35e3YpvexLrwlZXOpT00HXFJ11H69dLD6DuORIypkup2+xbRcj/S8b
sIMeuFMrbN87LxgODblwe+BtjVt58Po0VudXClD2S2IvvVZjHubOoDmdOBEF8RDOHFZbq+Az4RmF
zazpCJdBSXCO6xocEd4f/GDmV0gQYBShjS1Ln6PdisuFrfZpAYjhfgwDb2yqh3o6PPLxoDK7afGa
24wMX4HZpMBG3cI3QS2vuPLCTPgoD9DZIjGVHCVWTO7tShMjM9jqNAwEPZMnoPWCUvMRqhNasTOx
/NSFfG0CdasGAoqCEw1ztQ1TxegNxVMuxWBZ62xy9pxDuYbgLaCtTC0y6AOJhKqP45fI27HD9Yzb
Xzh5HBnuyj80H8Xqk9flGQX6+0jb9jVV83M7a0eSZKUES1I8UZrTt9459HWcXf7nKeCU5sRHk9+2
vLOu637NNDOt3GUmdNWoOiGPVucEm+b33GUmhYve1+iKa1aBe8mpbB79tjuq3KievLbElhj//cBL
c/2ujfnLL5fMaCHR/p+7XmuRnUDIdAtvicNfd8MymdqjVlBtqf7P3E3Jq3cBn+hLAB9Z3TNyGhdw
8s/GcpQF71YrenL0y0yUWYKcuWybTL1O/g65GEsVcI7HTik3GbKRw5CYwAh0o2bWymAvu4xjMy1l
1EReWWcaSDFpu8NJpcSrBF6YXxIyOtkY5nbquNQeZTKOlGHLibtaIVd7Ps3Hrfd65CHFtG1j42s6
B8uO9WgJoX4P6OKEArt47AW/oCYd5lOlOzsf99kENLfqjlw4PmcHSzJslbepUOOOXc0Dc4GMrt5v
nYWV1zc0vpnvBdn5PxV/EN2DMQgKk/QVLmytUTCcrgLy+FTTa3hGbprMx1eBM8Hl2z9GcMAv2kdv
2tp8fZMXKqxsa2zRyv4FQTCw5nw28A5p0INR8aRC1CldsaWV/t9U0fq3Yib5Epu66kI1unKfDZnr
f/5+QxlK60JJU0IXLQ38fECmjmsPEfPEpVzQyPgrSQbX4JK7jhxPPLAhtmY1//tkxYvzqgX5NV8I
XRk1Y+CP6tR1JUhSJCp1aWxyZCSCiB7Q2CD/y27RCJFjVc2pSfnCgZRPV5q+dLC9rg4bnyvmbXN/
MVWTKjHyn1+lS0uk4LlYCBytwAE22A/PEyXiOVMalUtzMfMuxsE+JSRBZIfCFnk3tz17dDU0a68B
3GI4bBQTNaI8nDONhWhyU5SrWciwrD1j5Lfsg74/Cce4x5plTaOe9bQeThqbVX46ZQV6R/m/XqJX
CDdvc9g28JvLfyxdnPKD7Mrn5f4JNulA3N7IBcnNFYCnngFjXU+kPCW4j4KnZQKFTG3xUjdPf4UT
Jq6i52uhY2lO3KxPVdA3+4HMETAAcSScDMbcA7THCBRW/ITimViUc/n0Cf8OjJ9sVR9AvwshGcTq
2Q4bCxVf67Bx100J/WnE0iYqkxF/XOm1nN5vIj2ofEntD75/NpGz5JJaHxYgg5s5Ubyk/jZgLRVR
wbjhb4u8ZbOgiJUMznpy4O8pf+Muft1/kGfU3O+ENBO6vACgOgyZzlDG2eKLXoF/Rk2q2qxeepe/
TjIDSu0mmOMm+kXeN6ihvutuFcfuqs6jlyfqvy22AoqtyZ5xYX8b6sc06vExPK5VGh7GuGxnl973
qs6iz/yuSf8qWg1MAFZSGsqRFn6qn6rQoMvr3uONHinumwAoaCj1vaP2fisNQgwHKQmMABYujtt/
BRyz74d5yvAWqY5a/SblkR5t2niyFIsJzzwJmtD028upamdm4gRv5+SgS1eSmTPKPNRs0baReknz
DbMLSTP9e/vfSQkDY+tUZqJbGpUYyK72Mx/U2mFT7lMJOgHedbb2XIK8TclHEfLQIDRg1uiOnxWv
rSkEMX4OyTMK0LCbNuvIpIb7qn5QR3oEVItvIRAEI67ozxFNr9cKZAZpPOlwQKRY22kR9y4ICzr0
JFSyq636E/qN1sEQ6bo73VISiV2QYMs2tQQ/6bKOnVnXDRTyjqXg9fSxgMSKU5mkQgiAPV88zWfP
wqUBRe27+25PzClKMXjmGEBs3CuEBg4TF6JE6bEbJxmSqyFN+xImnzbAIxFaumOg+zqndCzJM/yW
jqPXjnAAW1f/43iKTfTUjc+HpRLx7xTNOQRcp7WeiaoRAQr+Ec5HuWdBwzK6QMyNQJqia1X2VVCq
BH1Z0p0VDi/qthnsWLrZLDsrjOQrLQu8KEf2CHujsQEuMr8Sa7bfn/CfILdhlCCFUXbML0ZpCRp3
UZidwiM5xmx6s3eEfOE3F7+mhAaCPJ5yoPisA9uDC8Gf0UsMctFacdmGLfwoxqhUpChBGjfiwid/
6WBGIFDlgwjYFJvXukuoPwx+S4RGrxBjuf4k76QHu0wmsSnz0yJGh+ywmzF3oqUnQ4OiMADKason
yGhF7oirhL/V0fPQUW9qODOMYbQr7Gnt+q1mPXtf/NeDryPVzkRWk+RBo9NnmyLo/DBbQYEvkdcE
qRRVc5LuY2K1aaCA7c97TiqhW+9x7ZGxEsxmdU7n4ZKOVUqjXxxl5sIWlf/LsRe3zGqMLV9iHqE4
ACNhho1c7oLkm1LpNfLCgRaA+sW2ySMgXXyFxd733KR5iifDUdc1/TIl/6oZQrr9/JaaeSdc/rvK
ZlFJgY5nED+kPScE9TX6dw9wyiz/EQLty+1CyRQGdT+lDRADKEzLR/Lo6tOQ3jLYmeIo7GWDGjdN
JA2PoZ56mwSLEHx1cMbD8RBRJjNCcDj9tT8YTkwreOfv4rdwIjCpkzESfbWCQTG51S2FEzbjOVOB
Y7U72TaFB8DAD2XRM+LwWlAXT0mLjtoi23ASpuTnDdG3sPyequ4H6m89B8gvFFE/Aw7lLCNcpqaD
zAJUvEP82kuD78GdRjTdMo/BOWI7fo35Y3wo+iyyR4pKw4J34YWSQPIZIjgISpycXz2JCLjNNETD
v8eSAyKoAjTQmAIrMfIg3hz2sJ19NgTKV3uFi06/rr0vxcPs7fqN/8PEp8dPO3Ub+LFXfTW1nus1
WqNrf1hcTUu3HAs1RHPb8Fok1uElTnDysCaWugxCkj/03tW7+TWYALxNMXpZtH12EYW2vA/xvi/C
bGrmPgI3h5hG/JWWEKerMx7oODkFTWncZZc1AILMkkmAmVDjAXWdvQmsm1eqlw2WZwprW9FQsiq9
Vqa0445UwOLxtv0sw7/FJ3YldH2bF36YyoIl8TuGWIqvEyUrszXp7IpyMHg5+pZ9kYVblCTpGqm5
XTQbiUUB1uiMMmBhQA1koB7w5++i4TAEiz5F1HdaKtmnKMDzJ2yhvHXR02/IflOswcNFu9bSYE+D
0hbqraKFLYY36CytyETfTwh/NWXJibhx3fbxJ40bmO/UIhPdENxZBKLZGWbNiUjxeAPdFAPxYEkO
jzFe+ELbvzCf2zUp7n5Zhi1FFJaNifj+G6SGaCSFL8DXsrNwvxjZ+V42/Zv7xl4zwbuR3mtcYc9Z
mQsS2JzP7LGL4yVo/9NBIZqFLwiUC4rxIfMK2xuLhAH9pGva9JWTYYzy2/LVU0kc/tDxnBTl8JHM
NZnBIWJiRQa73f59JKQS2PPudeLAKJ5Y5fPjzTwQv0szfwNQO2LRJIrYTmkYynbLLEU3ZqSdvYgC
A8lqck9TMhiki/QrHxffCeXVRcn9KnKjoUxBTQIJnHKOQtwBxeLxXH86DzuhIkLFr02Mr2za31Rg
0bkmSJ2ge31L/3JNVKursfMOyw+C4hJMoafAKcmoQCD9Vszvwec4oFhSZvXufQLDGsgU99xS8YKE
qYmFTxIehETCjcsGEmqJGBazufB7Rq3ok4724BVrB9lCMwrLqi6Lk4f2qL1y1o4FVrEtZQIdloNh
6N7LXYugWSl27IkBcFu8gbrEc08Q9AOUeu1dkY966Z18+Ezt0XF/Fp/KICQ7Bzj2rvkPgIV7ev4J
b+VMOnY672k0slTMzgO/vtf9kAe66IHzGE0cqr4h8P97rMkUfXAThh7sOP/rMKHi27fJ9vkFt/cY
7Z7SEnwqgM8a2bpp2gu3H26ipyZ15cBiqfGFP84PB0tsDI1ZQ8y7WGq8PIQl6wUCFuquLKnMNFr6
PMdOuG9+wxAZ/81D8va0nNTmLugygX311yOKTap40Wr6cjsuHaaKXNrALmdMNOcna+/TXg2R2enx
31ji8utcua5W3zfMcOuD72fIRGkro4xOGKCzXGptssW3sXizyuHmgjwjjM+pqBa4WYDBC3t3TT7y
kEmUUVVYbYGRWPZJfuGG/4CQfLnDddLQtalQYeaQWAZvhqTlf2+g3JEQvtHni48cDCEhp7mqllU4
LFKjR7pXPB4YhPM+qLNGL+zTmmEeCzy8l3VFIYt0JzfEWjeAXkv4/vHxaUTku81wa19d2al8OxTY
GR91zo1sEBKllGwxb4bNM6P8/7spg2aS5JdYvy1B19ft1E3bJqqIrdAk60h4kCDlvRq6o0Zt3+ZI
8FZb+dmmqsRL6TTA4dnY0nndqGUph6AadFaSxBDecRU1zcyvTXU3T4dc67VELnnHZdB8EqL1roIi
W9zz6nnHaOtD+W1XLQB4aPOLg/bSl3IBALG9okH08EWaVsmgV1U2iWmVLdBOWcmWGbIJNdNkp7u4
GpW2hXFL9eXxJ2iQCY+RYzk9QW4pWqVo50cbkrnearsTRM1FJaSSGokEgg2K+1GdMSMBa9fJ6EjL
LBHvpTRJ7wfgHkWlmnMFlVAVIbArRxW0XRNxNJy8IAa9mPA9ELoHkMHeMGUw5M8zvtMnQWytiaLU
gQDFWv0ePr4suClAiGsCBZCZclJmtOu9hpQNcrGkfQqfrfqLltu+RzBAtKO1vlJTEPQ15IX17QyC
pMTUPUAI1vi1BH5PzZKLsrqlHVoXGHhYycGrkYrsXaERP51vXdE4YVxk5fCTl9kAuV1IiuT7o4HG
tmjw/r75uckfnuM3x5Y6F71Xu3viXqyW7db0hcYEDYMhBmuM0q+3HU23tU4XGraobkccFxsEnZzI
Sov90s7oM6Iiq8oZJ0d609sdG0zYmvYAR12nPpJZ/05oCbCQZcHdGT/eJYOIqst/100SdnjMfw5V
LrHan2VWJmQ/fMQVDDbbNmqdGEtBvqATqWmVUACcYWYHrxVPmdFNTMMTSboQXKJC7u7rgcKNnKLq
v36WvdGV3r3AU16ef4+19D0i0271xv0W/IyRrC+NSsBGzN4s79GFK+5BlCPaJ9d+XoxOLM7YZorc
6yj59NWFUbKjilBHM/q/hg7YApQc0Unj6dt4e4urNR7N1nkGjv0Cri+mbe/jDfDylqNOJu6lMxMp
wUZ52GUoTepiuCFcyMwuFdBYxsXsEXTmIxw7lXl1X4SCr3xXO3czk+jLUWup6ikPva84DlQlWYtQ
hq6qRBv6sVNuAClf+Xa0cBcA/SadvdIW/yT7z0TrIBMhKSvsg7CESo0IMg89niEeBvUdHBbaf7gA
0HEVheXL4bGAQ18veKcB9Z1aLEaQ6npASmJYgIeJ3WkUVHejH21tC6DTxtr1m9AOTKOOlmeuNjT1
026whjQikoq8hjC6HaDdDKFMcC561ZgvnjmKjxCYLtmkvT6w3kid9Mf9PkVwXBRCFNjggPtaQrt/
mUKsqJ8aiyW52SKuRD7kpmcRmlxSbJVuUJumf14MqpFiNyewRsIZP+Hxej78F6UTeniFTdHNXOai
3azboR1VLeNqkOcsDbES7lWOi5Yz/eLKhmFcknaQtMlrLEDDtlAqVz7IU+C8jmoT4FQTSbKOi4yU
Ttl5Tr4QGB15suVY9aB7tIL41Cp18+oVJ9IqNMGvThZV9IBM+vfMZalf18O/h3iDwrZGDMe6jnZC
FhgcyPBJr69+oS2LKfhgHrhsbYQCZGCUh2kKUsk3Ec/AEUl3tNcbsVOwFum8ebqeoGWbSHDNC/ID
OZ+OBJ8ehC+to2Av6ZWee+iAROhGgJLv/95NU5kJWMXklLK0wi+7VAWUebgD3FEVbL9cGAGqSD5T
/Av3Nd+FVfh6cQTCBzy/orErCJgjDziZnWVASwd67F/srB864fTWGvm0HGEJGIkzbcnjRdrplshz
Kco5ak9k1Bgpl4yPsrZZ/GROYlXefwn719nBaQOq2ADsVky1tlbyHiEAtunO1s92+T6kllH1ZFxr
FbqHJrDPYDcjmUDKMmpuysaiYb0yb4EYaxoYQ/icm2dlckYvYC+qD4iHrrulSYWhxSa2Ku+e+ePH
EqR2N2Zr6gUT5TE5EBG2WY1LzdMcV0q+HRrVizg4KJqFopWKY4kYErIlpT4sL9roBsGH/I1yVXU6
HgGzx5uv6iy8FI88sQPGMU+Qn4c9fRp2CF2gqLreGFfuchqeTZe/TuUsq5hVyRi6k53sd9wnxGl0
wNVFQzFNSHnIXwuKWSBse6s8o0+wULfilEgulkBgF5axZxWJ8lup/l10vGCZaOWF6QiKoPI/0V7b
CSeL7IZhou4xv6LDyk/thYdjSRRCrufEaVrxREGy56EfnJ296bJLeQUjn209ozAC6D13gckBgfWX
vw5UB2KBZ42S0AeL94q+P1fa5jhrO8UlJVcO2tIm1ce5xZ6M60i6mBkEJn9l5wv6QvhqmJ7lN+WY
DA7sRZ0/K32J4fy0DSehMWBXB1SaiSEJ8ktNjix6JeTzwxQl2m+dmsNJ2KBlSNk7bSVoZjUXkV2c
/3dhs/onbHrv0broKe1QbsqNcvdRANpO8Sw97JRC6I/NZyz5Nahzo9nm0nVYAYQC7jVkj0LUOQzP
WTP7oTdRJIKK4SUY+yhRDn/AmsUq68EgKvOhpODhvVUDfDpUJrOgV8w6mFSvs70Y/UShL23sZqaM
muedz4492fH2mGW+3gh3gLOcDLDVDHoUCRO6L2BF/jNP1ciixGeYFn4l/6qH5B9uTcIwF0bzN05n
8GGuUtSat1VLN14ji5aAlJsscgtqFCCsqUuBIcYc8z4dgqBWtu5dai0NagluvG1izKv2KSP7eaZP
CyvwuXpJoHeySBmkRb7ha27cCHm9JZYou7mT9rKQBxtKkqVxYbKgTPu1259Tu6Ofp08fwSXnHDMM
xbmkzZqYbOWcC8fkS/MZA+8P3vf/hzyurvSmO1cmAoiVBg31Pgvtpg5VAoDmqxOvQZzXA/rPWcxd
VHMFzvtkAb8INBbvLncjb4KQOq119Bai8z6oG6sCDdfOJyHaYGePkT6E5A+PbjCuGwl02bYz46Bp
BegtAxUrdLIFGgtNbEFgdLK7bY40cfbxFmXB37yt4HPdSIHaIgrwYu0G6B8DS6e74GNslVFLRja8
hb8Z9wQibWfdA28rniMP91XV1vaVyrSUKX4FEBzogMKynl9YMFBMb4BNc4RTz6HtcP9S9SqalgdV
Nr+PySHfkXX6N1/1hQtb2kC45eSWH3nsvdv2+RDYKSYx5L1Nhd7TkwkkuDel/iotkTZfaC39Layf
2jei384gshFwYNjbtpEX6s4rrYTeUYWmAIS6CoSQdZIpSM3reUHJKi1I9249zx1p4fr/g2/6GHc1
wMrr1B4g6BY7RZlIOqQAJkIC1NoaWp9VdtoAVfCDDd3/o5UdMf+H3H+THMSlKQg+6jXR/R2AWkpK
RguGsUFg7G9wiJHSQ6nJEgQ12XrgJgn+T96X8vIesqryL4KSOgXuJbAQATvgjRVUb7trJZxLd237
r1sPf41R0FLvbUl9+wMe017fCPcNNlR7j7jMVcYP9AaBZRPCyoGOthYLt6P8ahsn2EKfPGKmmRq9
oS1kImNwQefQ504UMOvLd9FsVdZnGT6Lry6SwW3IRzFudczH0h9AhjsX+gyfAmIgOM4nZzDSsGRM
jmiJGv+D4RCl+lEF+Sq1/48E+wNcoZaMRUseVJtSb6idhQ1o7NDx9n6B06ygmW+W8JI/WibC3Sup
kwc0O151sRURy3+pPCRKlBlwlHH1iZC4ovSd+Dqk+mWS4KmHiTcBBfUMAcMeHzV0/VgYKhWSslIO
ZXdiqnLj0WtQF/3ZlVnPPFnnF8k6gLWgNJFxyOKCFV8A4qvuysi06iD8OzJ204H7BY5Y/KK9Ev6c
t9r/x62c9jDawfs3KRZAeQyl+hl0hT+lugBuwRlUaxuWboAI0nFVcNPYak04t3Fz6Clc0p6GPbst
RoWPjirMT6nLLPkO/9q1NTpkv95W2GAEFgBZlfok5cThUy63CK7UzG7XHfou54k6bGdvPu4/GrAv
oV1Q0dpnTL6Ig4b+87FPY9IpSqxBablNO1fkKCMbjSDc7UfX6b9Er8/CvQnJ47tNdLLSBhSyji6K
/5UWQV+OXd1YhfaHss/GTRN0FVe71SWA1fbvi6AClUh/p+tpFPq7iy1T5fS5rdQqxx7tvBPKy8ZW
tXBXUXQ8uK7PfgpAz9nyqxWG8D1WCtCdzyG7no32fYH8E0SvZ1HFeq2p5sSO52SIv0wtOq9H39Sa
IvDvKqWh8NIEd08zyqEsalyGoPPHR8jH/7Y+ReIohNDhEJ+17qPiPrxnGVlgjS5G9dHqo6YcEN7T
CbX8rbE5zF4+WubiNNSwSCMAiYFXmM6JUYWu7qDSg40ZOA8V3Sf22meo9sp9kk2NK3lLNun+Dt4O
khPinaQ8PvuIh91/5hinaM+w1IDs7wASMmNPvhGNDlOmNVeroTBC2bjKi5K1J65NCmqmIKW12zwf
1u73PTan0hrK8FC6KRYkPB8XnPjEMO3X27fNHrNJlCDJmBo6ydVYdj27MAEyhV8zljf322s1mZYw
EVU6unix/BV02H+EqA6Ox6MkQ+/mUGH2ZITvBRLo+tcOTwIWuo4z49G62JonxHB8t0Shdi1UNOHx
ijtwLBBRfr+QZkphglIdFMpf7QD0hZGvfRhvoU9Yl5B5RDh7aJ1u5/Pg3gJnf005XQqmI3Sih5r1
qvKA8E2ZDqs1HWRIcDqLJBSmvXXRZYtntW+hwnY+6HOgrecYTJ+Hdqx/P/kWICxKk/uAsJCMipzL
TkzonSIyDG6MVdD/ue6TrKVkYeL7mt6KPAfkghiPRf/HdyC8U6eit5zypVtAPDejE0jJv9/vONxc
mvEpQIOqFFzM+P/5y4z/miiLMMuCqXST66ng+T8tLzsTCOnB454H7PMHk7cKXf/oKf9ZoVBE33HB
B/lZGVf4kUVFIjIkMVU5VQNa3loNel+WJ/xn1kzeXgUlIy7dzs9ZWvIKHbqF8UQMStvXALRCFU8k
jstbYjnG6yipnjgOVULx0jAtIJ1m+jPsr7NEPKA4smSfadK44vVV1FPQJGELnQsX5WLTKD6jGh3t
GHKaKwsxFWb7DzP/ugQ7/3mn+cuXiipDnioUyXuuEfAvn/Jp8CWCvrgqzDRaPuREccf4kEoAC2uT
4Y6JkQvd4BprqWD9Sy9EaqkTWGCKDNWHE039qRfT19RPCZYg2mtN+kztGSj98AVmzFEs1zcTxhNJ
ZY4lPkdWkBilJnQivaRG9I2lbZIxy6e8Vre532C9JJ3fJPqum7NiEQE/qbbr7eprOGZ1yurEiuKY
cMp4/8h5V/WcCgXGQVjTwtS1or5CRQg9vvfV320xMJLZVEVeGl25pUP9xZGQMrdC2VFdrxTRcxzf
jTbsveZ7EVQutBDaBqDDW6gzEp1YOt3bQWSqrwtroGTExCYc+OUBDQeGb8N3A01T48SQs7BIoyYs
b+HDtkf+PQH1jYOx92+A2vsIlapmZxMmI0cMDGbXbRrqlXaLmG1t1JYb9Mugkaxvaku1JINMM21Z
2QaPqBrU70ZbytENdv4SlGewm6Dq5iLAzzkk4x8oFTsf3CHDYyAdgFCgCUBVVZEdXleTI4jf2GnH
yir7S2hmgi6gtWL0CjmzVH3BHLCCoSsIZd5QLy0Lj5NPpMgWXRmuYNKcWA+iVMSIjS5m68L7v70T
m6vXW5vT+x7520rjIC8JNxuAHnLJX736E99lHubGMTngOdagylZMMRF+BsBgmWZRT1XJuibGRvfg
lexcLFyOmVqvTvO5iogINWj34YwHEQreIyWD0W8ehtzysFUgZvIBmq9Ht0SX/rC7CcoJWhRoss9M
j5X9U8TQqIq9q4LlLrYqQHoy1rCo4G9um9cNeBIOwZB4ykaA2/i3W9gN5cJzNTcHADSiYqwf4jeg
hRNxhnLh+0jJf4ySm8xOQKzlweXxfilED6Q7bpBwj9AJzCbxc9MuJ4/GVllGmGMmockntfzsTJ1b
VTvv7FZ5rQ9nEsy1Of4EdqJ11lW8kfEYsYPPjlSS5oM06x/O4+W/h2+UaR5BdAzHFxoNvZJ5bRcf
7CvBKsTJ0ZodCNys7VFFJFkROXMSBYpxmWQkz7Vj+7lJG6+MNIjKC0CdW2pLwz//KQYbiUciQxki
Rib0l0PgEujt99NopwF+z+CQ8fjwDkh55IJbjaJTX6j/zOnSC7dt1AoFQlHE72H4rB54tGupm8D6
DmTEJUKtofpIqWPpGaDpdSYsi9sY1xjXpPos9Wzx+YeyJQ3JyTxZVx8S8qrtAd4x00ryHPbrZals
kMg351EOHEexD71VfowaCtNC44Z7KmqW2e0tN4qwdTLYulUrSqvw0agOeumQ5hE7cP8vc6oV4FVX
Nfdy+qkexofQbql+1XBukocZANlrrH49r1175nePUqq0/INlVvzItPXzpQdwHE9YuViZv/3EP0/1
UcLDS0seXzlS71MdzCZ+O+WKb/FJSjJOAYvmB8TNbvRzVK/pK+TSQsDEfpBvzbvvThYQxqPq3L9E
I4efU548SiMmhWt8qZfsNB08SaJJDwpfo8D8ic9R1gNlpcntDsltcyjUzYpr+FwhGVPuKniUFnXx
oguX2SATA4wjk5QlRwNOPNFISIJff/2xufVF+rejDg+MthcIhwIX4Ov+kfAsWmjGPOG2NKIX+i4x
j4202+18bZr7Oke3sU0HL2Ur6NamBCmYe7YQBkV7L/0rgqCBTIj0LVHAVS8O5mZC7dzl6WbXmBLm
M3KJ/JW1pfyC+FxHLyCkPMvglLh7oVIrsoEu1Pn+hUUosvkkgqsUxDyzdAJI0Rw7ZPgyAIGqiNE7
3M9l/TmQAQ771hLUSXoatz1kJiZ4Fq+N/Qck8XEvMmH0uMXSWn3oOFrO5owiAbDDKMdqmQRWqtuN
+86WVA3LQJE8Ss2Fhwn8VP90BFLtFz21oYjmXXa1FSssoY7+wrhiMmJRq/7yfk/6UBmgAi279Pwi
qWxtMgIcEstj7c/yNUtUhJeb1i9yn1BhZgnGnuLPZdJlC2w0uOSwCp/HyHHibqj0Gr0L7G32X+TD
/8xjZWsRI8M2u8r1rIIEA4rNzBxlF3pBv/GqKW1CqWptCHiT2CdLEySi5dSHJJEE6r9e3UQQDVM2
2BCNDzqXMQ0njmQCHeHtRKV5XVILfu1C1OdhuNxDWp5yMRDwz23pcvRaPsQ+Ki7eaeCyM1X8utMS
c1hsR3a3vdTxRz0xHAICK/n/+eUN6TFbXMak5Y4V3ICxADVMbkYHJA4+WsxtWAgUQ1DNRG52s7At
/sOyuTORD8mjZBNdBk2K9ei4EeNLKuYB4ZBctCPOHh3MBqpXxsx2mour06P4rItbsMKPleicIONS
FZq5pT6YZ5bWG9ng5VOzcjSbdC3W0C2Iu5Wyoe+REeTP9LpVjQS21tHustMioR+QGZLe9Mu3fBKC
179c94UAKDBKYDCcnd0uiYt+Oj7EAaVmEQMrC0rJIFaIB6bCqy5IoCtF+4IB9xb4TjsMoleZLftS
XtsqilLr+TzHNNq+j05YD93mdwdsGsUARbnsCBQ7+UfHsMSKRhoXxQBMF3vUh4sTrsCn8lZQ/p7X
74ib2vFUQb1PGIYkDZcm63RWb2nppPCfR9C+3of+kFSc+awMKi1I8UwCb7+Mbd7464369SU3bPFz
KPu9rPnJa+UvfvYJYy8IAOWdB1iVET8+y9KF7UcmPrqFeX7/FMra5w7Wzedi091kPhMRt3ciBUDp
YZeLVTJj/JXTXut4nP3M6zCyo+duHUbXwr/ZLqjSjdsBwYgWHVY0qSJ4pt5LmcY7kftDVHj0w9XI
KgmjDpaC3HGQRt5HhnWXGv3dfJDhdW7EGeRxNnN9jlewz3zJlUXSSb2ecmS8zzCU9Nd/sMZdp/er
IDCwCWGh+xyhHIPo2SugMxuD25TXqKJ6x1zATCqHw/9OtFclGiTC8vCBWiNP0+bllbhYXY3yuWKa
hjBNu3y7F/1BqIXAcTVTLkBVxIaaTKCXCCpD9Or724wpVyVJV5xhzoKNL021bhpcv81KMB8uHJYy
I3/lSLZoNjHChtHVD7oP45wBQ3FMS0zJ/eK0OBdk2w2WAuOb18jTfYHUJpdgJoO8+kA0xpe3buwD
TyYINA1UdbMIHRpUQHkh3EKZtsLc/nbwNT/yi9VSbIOPyKVwbd70GPmO+2xAwCREOGrOFgStp06r
aYgvv/bimTSxs0n6tVO6TzDKN5W9Sh91zbwEFCdN5kW1Xzc+8wS7a6crtaIRZ45DVgblWmh5CtPt
TvYBHLIqIMDk2LzDbEjYy/DjsadqgTiv3xHdAO74d8QoS304/Ti07tfu+6OsfaYUA0nqrVqcB3LM
2EoeVV5taJ0OD1wKwTj3E/+fWt2wKgXuaPP4AcckiYNWcyTvH5nkG8k6mybEQVJ9TvnmWDG22o5r
KbJ69LfrOmn5R+g6X2xler8p40Jm12vlGM219ky2j8kA+1LCWLmoFAb5h36BSDj0Mld58G7H1X3v
6FKvAYw2tCh6y3CRDqnkkL50juD6dQ9Nddx4fXJEwavOe/3mbGClWRPbdGP546Eck6sJAKqzVNW6
VEiMgwFT1h2hOxz4PopuPL+8cnSv6Qd0GgDgfMTlRSIX7gEMkRBnvf+24TT+hcLIckt2WNxlFffZ
Z+yWaAsRmJHA1wdoTSp9DTVld+cpXb2sH3c6/I0Lw7GSAi3i7avtZ+hudIjagDZo+Flqkuw2uYGG
5eem77dI8yM9m8QVYERatq9Lvx7yhZG+ndQXX7DJzCuLLgatneydz7jmrkbE5i7kVCURaKwlDLrH
m+oC8ZAkHhL1aoAgB72/7W1sWN5FrXrfBCUzXxKCX/l2T084FoVDeL/Ps8ZotlHWzD89LdNYzQ9k
p37QcmJprxkPEAlREmWCa03zIy9dPCM+c+S1jeposTgjH+LKVSyRsOim69bDPaVkpIhYH+F5Jyx+
ZRt+XKu2Pg3haewBUca44s8wbzOoT2CtNCFQXLRmWe+TP9CFjf0Uvo1qH3+qh4kEOuYF407oH7ag
4rLGIUUGrx1pNYoHMiesjOCQ6s90MzDeG4oWDjJCrg62HhC6mAq4RJwFB7Vs80I/w99YqlNgH0rv
hcObCj7NwGT4CLxp4YLe+Pw+0ySdeStZeQP3+q/YlAKMWtCCN5akcZgS4nRJXiLHrqUVrUu0lIDe
SUDt+qk3tg9yzPvNosTFJ6DDTY+KTFz2gz3tEtDgqRg8pbMRjPrhLzTjS8lsmK7NxL+ZeZqti9jV
ZehDyVTCPMliTH2GdzSqiZU+4zfno/I1N9RrvnpBrB2J/ZnpMm2bcyQoAHXJ87Vzt4w+ybPQVwc+
oWZxAk47lOP3ScobNrFsH7gVDGqjfa3DBe+MXrapfZSORXlLRogINivDUG4M1sdOpn72D8MAcUpD
jlFawLLvkbn0bgwUewURmErfiFxrvUPH+ibv7IPMcYJmuKrMNfML2Ll9lkeYy0zFiISLd48b3D/1
rtWhLZTuG6isPZSESH6QhWyuBJZvTz3J0kdysJ7AGDNOM2yCnbkyYboox+ZvGc+jSc4Eh+lk8JsD
8m4Z6jkMPWpmUZwl4BmHCDj/02uF8m4pR/Ai9f5yRxWtTTu6ccabfxew7o5yndj8hjEJM3t9BQVV
QQDu1hjmsuxk5mvp5Gp/TQhkmq2jYJFm7C47LeSbVMApkUW9ZBvvWvltTKkTHeCNbTl2FmmUusdv
gsUzc2uFOwFjHBnbJ8YGO5LYJAD7Da9Hf70Ko0dd1surKPdPPT8wixmTGxkfywAb1WlrcoNX0bzs
e1Zi0hUcgAA4AFhIZdLlBp521CxSj181sMRH2ZON1VvpO2xc5XjHMdS9f+pTd0ETB9o/yxKLAfCA
SL85yMSQXJYdPIFDYF3H9Sj0Gos+UoTrBVorK5C37GhjpGMbsh9Rf2kxtsTtbfROJa47LxFnFgxW
o4xDH0EnfUFq9M9Ma6WiMrKPYF8lsGtmXpHYLzIAuD9Zx992SfIOtZNZQDIrPg8xNIfRVIfWpr20
nC0lvCJoJv3FnLou/DBZL3qBT3vXZVFmnFshYCewDw3TK17XStWH+EvRT1SqJB44/zOCcGDWJDt/
IURYY1zBI29JaqJ7ZNWPkZOw9xsbhWLvyVH9wloL/1/ekwu41SO+un5J7cD2s/tYW/iWXevvpf09
lTsqLuq3vc8X0uP3JWym0l7ArpS77ZsC7Qrl42SdASGORqvwSG0sHrcOCit+ENxqRtasRGqNEdfH
mNz6wyMyjuz2sm1tIDdZMNYayk5xndzpznmdZaply8jNXHqDXeNT2D+UURzdKAjZDXgVjZ71REQg
f5KFCHci0FZpGA9nj5KBautXRVSCqmwgpEVcP0p0+tjOJF5cz1FFCm9uzjBrwUUYXzOtMvY7wq4K
84ja4JuPFyPezvLW+4+hLI7jWwWz4cb9+uCTI8+0rhFULcLL8PrIWgE3plOf4gkOLH+VCS3UTC5B
h0LmPupPvl1GcVqqRyr8WqLWzCkN7fSBPrmLM7NXGV+lV/ktGQhc8Gp+wE43LEI4RhlkzQR4WN7V
fqxP2PEbV0gn0qvCRa6wE8UTYLfCIKdeUlgzkw3ZPJ3zPKWMO7WDmXu1WNutYwVnUq1cx3m7j5mN
Z+6Dqu3Copm4/3/M4XzRo1TJEjDAdNGzqVB+F3tjCwwEcMQ4C5RCchdMNQ2SLlGmZ2Vy2j4q+Fmv
8VUrwiP+u37sOMmIAmP0Gw0swIsMJ1GFbkg10e3U1xnHrEro5BKvlrELOxiqm5OeX69pP4gNphoK
gdqpUwk8aYuDTbbgeMOHtYWPhgoJhQKHd3o00al/JNFLNnS1jPDB9XbzLaG62ZYvk4oWzuxIAD9h
MXynxaGUSOWyx4iJMzLnPpxH0vI0fx71a8BAAJogqpgugnBWtD4vxv3NaQnoLY//Ki8FGnb/Lfd+
8r1nI9zBEheaoC+vmyBgi8bw4tnC3WFBMZfrmA0IhcSzDCqirDxuEqNKOEGfIfS7xgP/o/MHvROG
O0ixl5pnUXR+CyinfSMkp5X5bB8PznJhOSLoHdd3G9igHVoRAYRArarn7dupCiD7uiSBCJwDLY55
GMQm1+g9tKcc4KTRyezfO1BPpSJabQ0zPQ0Lnu1cIwu2FcruI9+OzMhW7yDtEwLnZ/OxR7X69Mng
XHpjGdnVBVWvefskz9MJs8ioICFEINfnvpuhjhfU+LMaXvXkTOEmT70DtUMq08542gTlmS5pMlLt
ZKQ8zRTuv0kIcFEeHLSKME623TMY/JNR2C1sStsstxA2ixmPYnT96yj+xvKWD+OU/KgSoeow62lc
Xs5g2Hj+c+IoazTq+DrWomFrDUvVFV0Q7PMoEK7Yk27U6zqlXk2M9H51Wi5uZ8UkiW2lABcxaDgj
taMB7HkV3oN7T9bpthtbMR6KUfXsUV3It7z2ZK0AxLREF1lJa+VCZaSS9/fpLKzLNU7Su5h1jDaF
cB7nqlMpjpZT1bjRC8TSvtlHA3+cUwxyRI0kVBagYeo1J1oFCAe761MEBShNQPolgcYXg7W2dtR+
S0gphRm/d+Zq/fHCKfjUPnHXgChAvrQqhJ4bo6C4tTnI4w0DkTDV7LEJNHZkqHHU196XM1Yx+49K
Ozd2N8Pw/lNFCKufpEyQrLLz7fU43kkirEVaRcpvk04oaFxoIXwFRYuqpe5sE5dBWFmu3D4eDTw3
9u+tkLVVBxEt2nVvI2D4Cfzncx8M4974bLv9wVilPtJBBwD1yteQv45T0iGUs5knMqAZ9+udPyIw
wrU8CXb1o3osM/RRR+mRNu0U36/NsBDzrPpvyLOmCu3r5WFku+UzjSJYnxKEiLGkCmOyxBbXDnoP
B7kGsskstweVJENENkzCTAXBXyL1Y7Fyt/h8OhlHj2tW/7EMA90MND3z4kpx8h/USwqpqj8b6Brt
xaHH4yxi0M1Gp0tEAbMRPAxgnl2ewXy8nAbreoM4aRoRyObj8kaVs0q8ECPHQBpyi9HpEaJtRkg/
xXYaQVy8CatSzRiO06ihwj0eE/PLAVih4qavIocGLA0nfdLE2/JJIVIzplwkhwAHnSQ3Sn/fpJD+
qZwGc49pXuVThOGgunx2tWyRfsBq7pU+gXBc6Z0F0rpUaPDKx4gvSSPU70ua6HVjfi+g5rqw9mmd
K+rm6nFjPgvMjOnV6MI9KvAANVOXBdfPnncBhu3C6r3ON9vbM2VzWAzViHVeX52d5RlHFH7HEShq
5zjnk0tdtXBgarj0zOwJz2utOLeOp0gZMJHNxUuYZeioP1ZECcmS9gGDhNlCKQS7iGbdOvhhDS6N
lbqLijggV/pe4v2HSz6xskeqIXjRZuN35MW6hRxeSXewHh+/Icif8FJbQi9OSrfUCAk7Ie3oL9ZR
eemQmz2uAx3j+r/vrhq2gVlRjin6o2nsi1j8OrlvFECl03eBN4FzzT4G3sAaF40d1ST7aucSk+fp
g2CHjjv0eLLxXlhQnbtsM2Ihl6NB7xpKhRQrbBiALzJXS1+mZzgN8I6R+J5WidlEX7U96v2ftQ45
DDUTUbwUPgGttMszFAKWli9k0MByQQjv4AStMU9buVl7g18qyBPP+mK+GjlolQvDyTjRALCqhEr9
xM6kojYVP6DC8l/1Uq+6DivgaKvQSlsFKFop9fICxOAWkexSXLR+S+6DVgL0FCgcLTlB+It5lSz2
r7emFY1H0hAN2m0jrIITBvPjvszTAoLyJ1ZUvG4UB1GUFbdPFmmmlb1P4elyBZ+BuT7b/zGbsEOg
PagZx58tdHsPLv2RsJnrTZ39DJyZAN5TApBUdyYkh+cnRxeVDS1Ju5WocZURVMXtKPw/O8cY4FAk
JGdAJhMR2Y6wNIsb5wSppd+g4ZBOxKgIUZoXTh/P7/AukMuDW7cQTxoBZPd6yx13Eg0HpD7qYch4
SbuaY15Qi5bqp7srgi4Nbsl1IdIP22OzYCDs0d1LVf4RWITCmis8lm+i7jyS0W0EK9jFqXiXPUL5
XBPcnfA0ZvOv7/NEdV98qTpTbt50DxyyGoMYUYkE8fkYhSxpowbXsKvsGt4ppylj+tDzo4Rrzaf8
YIWXjhnSp0HfpQ9BofLnA5/AtpsnL7YWVlxrr5Zqf13mO/wDY6APVKrcMvVTXLooTvQhqZTdDgvm
bQrBTcTfSPGQg1yD8ku2ZHexiLaqLCXpof8PFmRhvcVxOZzUAbg/PQt31MH2Okuhgz9parNen7Je
fr++FWkJPvlqVIlK8P32QwIeGgSGXOjUjVqaIRYA4mlrsKi8OJRrbi4sUAZYXyQLA4mEvoEkCcDN
mvADTjjzAURuB9+EPSWReYMPCtJaw0FHW0/sgf8FLOv9KJK0vQWU+Vxbsc3AvUiBGAvPZYEcpPI+
KVhkZ/mlRARNNXMI3A7omKdCP7x3d1lHDjCA4xAmVPyaup2+UYzHlUhhxX4tOnuqtHz9bsB9JOcE
ujZuI0AyZ95MsK7WiSKJpN7vhT1wudDyjzzvk3RKY+0gObs0iXV+umanvnSHWnjIm6baLJTN9j9A
gEQ71zuTOcy578p4PtKo4JeVwBDuyBCmT5jfJvTgELE3fXWMtckI25euJHjhP+BF6bISPO3dIDip
LBhJ1cuN0+mEAk3Vz1f3Ge/8l42Cty6L7Ii+vOP3S3yvabjf7QqbJa/zxHi/KIyDuZ4McFVFyyuW
gF8beMrCDzvzvfwnXI2YCxe5Rpy2jBYrrVuihuxK1pFyUxexMEE2dousmjedgp4Hr9GmrDbIHQQM
26BozAIBL02I+MCLL9j552/M9Ym7q6KawBbGEMHp/t84RPIwqyCgD6hTvgwe7/Tbc5i3WAQvf4Vi
N8hKuYuXbAZ8CFnGK3HfLOQekZpIMYgEm42XUIqcDC7IydaDojSzv2njuuwx4XDFz3/KmCvwhjeM
Nir2j4BnTsqsuLv5L0KVoD4mXilnFaCskVEnbGagtOXjO0DHSf+KLIMGxJZKhEHTIoA8z2Ov4FN7
Mosedef4hQO1VHf/lUxQ114lVB0y1eF2P7B26vmhQC7oAafHHzoSo9o9MulSOykmndbrwlENrfiO
otp7JmklZWi99upQqm9kxn5gvpqcjlYfXX0G3iucEVkfnXiq/sfebsc3WcuyjAu1kwUsHKmiS9WR
ER+CQSRuFkBLtsjhrkFCtJ9Ups7lTRmaucEGAGSpyMHiXO8ZZY35dXo+WADdGRjOzIYUmxzld4Qx
VLhMwDKqi0nRUIwnwgYyM7eV61E7BHxfxJYt4ZT4GppqpxK4E9K1nM1oRezcyklaOgQU87/mw186
NN5lRbNT2swNjzKJblYZM0dynBUQoCnS8ZpQPQtXt6RuN1NKS0yNT+VaAkakkKH76JeqX+e/q1j5
wjxFU3dyLWbRQOVZalhsa3I8b8+w6htIwNHj4/eNb8fCZkVgkSI1nI070PFZq2nUSMTuu6Avb1/C
ikHLzzQouhSgF6DLp3lBv/r8EFPi84NeOJMpL4fRnMlp0myu2q5KAJr1IeYKU7j49wRmf/pY00WM
RHtMgMdWeklbMLo7II8Wa5JTAsl3+7QVQ4SfAskSf1lq3YWORZ00jNJkoFxkxwEUj0bVHLaAQgZa
5God/c4S9Ue+8xHC0KVnbXGXFOJPxcfkK+Jz3iGo6Fx6Dl6pRpIthQyQHtMKa7mRJwuCYJEYFTe/
0Gd7qTT/qOEu8qz/TV2AMcKZcw6IcWrgXALlvVlwQPe4dc/BcnLh5gM9XHHVOmt9IvjK1hBXzy9B
v/Pa2ipXNsN1O4fM+oOR0ML2ti8pPbjnv80c8nlJal/pbyI4CZlu+IQ+v4qcKXTfy24TgMP2gmta
GJJnO5fzd/OyomgBmGN5G7p0L+wWmpl9zetGrxk1vXxuwWCOjLW8ZXfDNmpdE1H6iov5ju8docSc
CyGOKsOgzPx7y847XLkJNzK+x1v8GwHU+0fRv5y55ZpmAnrn6ZWb3Y1BzitPmsUuYuOOqSmMm/i4
M73dew+8ERy6FZyb+PHlyEurl6Twfg+cXFu/zAK0/EPM3/+4+SYNZk98OqNx+aLZvjhFfUTvummq
TqGTJoRLmnyyDtpsM/ARf9BQQoh+hXg/LdAGZmhs3VX4M2pDFamOqVwHWCSada0FvplewVz0I4ve
k9lpWQz5q1QA3EJMSVbB6SPLdyahjxEtiSTsMuPWadFcDXDB7WcmPoUTLJLRiQcMY46SEvPmhpS/
ux1Z18GSK7G07MMpgPUctBMeyUvDavfEJ1cFgfNud3XhTpF3bFShmCupwW5LkO7EVY+i1jTOG6kD
xaSvY7OELVcWnP1T6T5W2yNIiUnSGzoMn3OU8mGNhf5tff++FDisO/S9SFIrJz2PEwSAMqkfGgyf
Ig9bOc8TUgTvCVfCd3jYHKKfoBQCVrFBjpp/JTuNJQbwICE4oPqLnjbo+deHqb66TAiahELHkybw
BPsHdeJYSWMkEPy3COdu1x6+YT9qqc0BYZ+wpMK41x52ZKRYdxsRM5TRk4F0c/4x6oOzARZfnzlx
i7fC5nEVuPrbMY4f1Yy26D12g2QVM2UIWU95Fb0/oqOit1JeyhoAlGMwP6qQAYviT5oA1JM8EYLt
G1/Tsi3LasP35WMf//9wg5hgVH2MsMZA/8gpPYc2KFK+W00Jh+nUY4SEQBzwxu03nsZg1wlTV+Sa
E+pRL9bserOluLJ24921NhwC247NVe355O+6xZV1jYytrnYLxvbBiHXu72taNXSBIrWZzZ1zHlNZ
SlNDm9LGn6cJrSEGZfdHZTKuy9XjxQddmZCRSMXKuYrRf9ZCQ7Cbvwgn4t6YdXUj6eGAp0EPx30B
fC/NFicvsOyydSovKN/KyPIqQXc39Sjq+E161G2R6Zd9J0/7Dx+xeGji9K1rMkGLJI6WS9VlG163
9wm7wxICopJthdRsUk4Ic5g0hXdNScWA2kEAabbO/HSxa+mkewUsg4sYM7lqW5UUDh9SqwaNi4DT
AL4H2phDf2kFCIMT3yLBiRclqFaQm4h8+A3uxSL+WEMlItCQ+oreHzKpSRjSuKs74rraNkic9B4Z
Gm6XP+RtIPhazev8w/8VXxLN+vqq4MhK6a7GVaFHrVj/XOfndToVK/lhEJhs9lQUd+JH8fdlpOco
2dqS4sCcFGSdLfZDUPEoIxJbsael3kqPMMzeKrYyWHavWjZ07yxRZP9E7lRWV9l5ffAEVTA9EJRG
v/W++2R0J/2RlHfWZygU/ZC0LcM8FUzKu/GXmGR5egvVBJqmODW2ex9yvUJfjSI1P8Fnac9ydkE6
HvSzbuDluhb+srAMh4hqlLE9uSRslxy2DO+/8qvhcar/ePX+tQI0S+r6rDR9tye8x3yN0zaFwyBs
cckmQsdD45ei/0eCj1ylWV4DXnllnwSkgWOmKI6CbxZOjAv99rT+xa2Dmnfz5e5f0V8qZi3BjSGN
S5Zkyp1TqbrueR93pMG++jECDJ78qPcwtjxbKMEb+VdtUGvYC+lMvddzB5js8UIJh7whO+KzgX0w
SRNkFYOGo6Dolq4F7+VcZ2ZF0gDRqqEBH63i2Au3NGnhuc/+X9zo0vqPxREvwfswaW6AXwWcBc98
a3fmCU6Xl3SD+5yNO4ShggJjtUWclpBpQOWFRzTvyQfCmyQTIk574oU4mnD/MsbC0iJs0j8YIs1i
smCzlzTQhsHE0ggpWmWUQ0s46DXKVa3Gb6r9gDJUdj+oZvdFZmCrtV75xHLPHwBQW4TqAHQc2VaR
6XlqO6p03/+9F0Im7DqzVVm9qtJNclXnpJ7mthCIp2WeHBGEq+GpTUMFyIFhLmxH+muwFZjY3hMg
CWeHiOf1Zhr+kdQTLFrqQCIETZSl3PYEf5EflpXnAXjvAKIL0BZ0N4oKArsLLw580CaWlqjrffyy
bp+DWxN+oFRyZnUiMNEcm3C3bORPjnli84+G96iTUsqmOaEx2IekqXwM0fo93RDHFjYbp1rTdV6T
H+5kxlQYsjcGXCap8ADpYvUxsSzAgNLLsxs2WL5d9m9AIj5lib5yHV1KIv69VyIKNIxuzhZ+SBoc
u1aEYmj/LZIavnas5oGuPvU4Jz2g2I8ZczBmQP5me4cV56h2UyE23zeYoDHGopw9oUC4XIX1oRkQ
J8xxkGxUFnpSCNklxz4dIdu1zkoZHj5b7zENU1y5oBVlmZu6h+VBkbv5jjkYWSbby1pN+393It7N
i8PQ9+pVKvxMAUbYDR2plhvoCjsqfE9IY8hLn99m/64m3uff6PhN97nlc7bSySKnoxhnXKLNwGkG
P5BD9c6nsJN1rtlsywZdQ4Cuf4i6K4SptqOWwOVi+ZdOUJJx4wGhIEso+B+6nuzN6fepRW2GvY5e
fyBWiBxt1MsQzRWQCxdMp2SwV3GAX1ccnv6IFQQhKrO47QcEGxh4ry33/VBCQXdsyv8qxCeiX4KG
1D+4qOnXg0Np82g0pRrchS/qz7dm/uW1EuX4cmqSru70Lsnse/jLrb+q0shdAjwyW8xTdVQwkHEo
dE83pzjU/VNiXqsjW34RyesTbkU6tkXzo3NUwwy++DJ7SYaq8+bXVw8GQQFgCCUww7pAAJ8RNpGW
IPc/PGYbrmmstgJWzAlJvC0UGhQNZI1r08FMd2vORCkoSXYH1YSfMm61xhWxeDKk2mOJuSP2bHD5
c0HoK9K2eRcSK7Pkl+qYCR4Q+gWxKHGKXqaGUZ+cZ4GjKCZEeHfegdcHzZTRB53W2zrK3c4kUPT/
8n1zIeRp5pY0qsnYaXQijn6oXfpcCTviEoXwludIMQyHNv7fEOLl6y8J0wCtEjiBT1J57cis6cE8
CfTw3QuO01lUAKd9TlOMHJNZ20Dx6JptNI3XuvIEkFlbF9iEl40rDR8dITh2sCPgKDhTon/ZOZc8
l1lN+QPVYpz+KAOgqErl1j2T7ADn4Nvjy9ztNNAWb7IaolPl9CnXkV3kGRpQUtKsnPNRha03ZZnr
gnXaEEdwm6ne63L0NJx4i5tBAyDlEwuvS3BPOkrxR8GTCKrIlhikXrCLPG7hiwe6IpaXHQdfloh+
QofCBISlhP1Tx/gqbyaf1v7pX2vswo+3zPdyAfwOSHs74ooV4nGiVi1LOYrQQdKYWRFP9BuJ0eu6
u8vJCPnglNfww4FrTE9Vxs2naAdjX+JnSFEGfyPF9EYhdt0tQDb1mdNWV4/zb3CHuHArb25ruzOu
AzlfYaA+GT6odjtHAENP0g7rd0opgzztXn+4deCjvKJ23/tQ2kzVSlNkgoUQkJCuz9lXP8ZXgs5U
h2dWW+pD7P3IzwNaxGy7QRY5+dVmG8JJ0AXpGpUZ223lDShC0EXL/kErauwTMApFvA5wQ36jxtEz
geSzcm79syEQIKP1Qab76mhkzfGVMha+8ZctVnZVO8nqD3oh2LosS1xQG+Q4ICcIWr33apCKynhD
X8YGcFn4dtPQdr8iTqv+EaFIvv9uBTOHmLLRAV8B8BynJCu9y8tGQvZLAjmdQldJwZu99bjC/zz6
49E31YuHFc4z+CHcf01KnT40my4ODYYm7/blpLFLYo4Sb2uaK3vCj31hEbx4MQIqlQC6YEknICOA
/BazvcNZIiyCF62NrUePxNSV+u1hsMhHPH9MFsNVriHSmHvjy0Y6APDtrfVPBteCQMoS0L5wRHg3
9bFe5mIU6CN8Kdmr3fVuHN+OZDKZUS66DU/67XnDD5ObifahViR+hnq8TJYO31lXRGR/JyILcfb5
tpbQas4Uwwjjln67EB683vMV0Vdbi7RODl9KziQigLjp+gxPbvXmTTr093Vl8PLutRlSZTbt1BhD
MVR1qAfM+yXPFpivW1ngxaiU4bt7JJUXeD9PkqzHwIg1vVABAtJc0JgAgT8sNl8C5fWFhU4HHyqZ
DkoXNbwMXAVZb4qJW7PaXZ/khmU26vdDO85qHFVWhkyWoK1DHByYyuMwlEU2xlnBprdqwQ6+DQ8F
/BIDIrNNFaDoLTLmyGgVac1SgTzdetfAYFxhmfq1FeHhaKWP66FEC4FQxfKv45s+//fxGkRYeL97
a6v/Cp56vd4kKX/W1N6vRCR9VqrJXlaxrX4AG4fRK3Zs3O2u+AmdGUKIR4zc2gzK5CfAE8fLIZb+
SiEoCnqrMoOuiqqhFhFNjsD1n3lxT3GjCQF0Fgy+ywxqOU6hVWJAtiGk79M4rmhoTnPoRKZdNvz7
GvZk4y73nKSiJxE0KfG6M6NXHkn67Vtn5a4DDLESMv+L2A1BFT4YoaPY9gDj3NRV7HpvJfgC8b19
dXrbiEGUG0WX6NSI6fk+yEVBoSLec64lldU0H9fpXC2mKIpW0YPZreJJ1SUJPrSvNocScV4Pne5b
V+BimqTgg9wg+AUsbu37Dosonr8LG9VGhOegm7lmcmFPFI2es8J/JmfnMqGmfTaaK8J7rjgsKm1f
iZV/GfxcVAMEEZee+qR26FFlQZQDXoNAgskakPle4c4v+wXVbYYE5M8fcGFypICd3x1KunSSAjfU
yXeH3WFJfuJSOjKowOVjUZqs9+glAUWAR3MN46hsou9w59qfqkoG0fDhWZ+Iqf8dV7uoiPDAULvi
sP5C43cKiVDShwHfQ5Nq2/htDMWex544E6d3MakXzcaP5uuSyBBxdqOiMmZrJuubktRS9yIDkVCP
qWr/MIOa1lQNlx90iCqfLLxoJt87t0Cd5k5gtisqJCDT2QBV2Cq8yNT9Slz93pPhtt89EjAs5k/B
R0Xey9MQM8gmke8VM2MBJSuwfFkzW/uRoL0NNU8dAC7mfchiMhpFhUoKh2PZ3kwYCq3hgfv9F78e
NnTa7z2H9UsY5TyDAcAHp5rphbdwcwZQohOOiP9V4u0cMXYQ6sG2W4p3L77Oxihumjvxrn2B/dTr
cUA5KxMSEgKvkhCDT6ERkw2mlm1DJqbEqxdIky+cB/BgLEl8UPg+m5cN+YwqVimAnQpVSwBFW1+z
ViktN69mOeZUtlhzXuU3cqx7RpbRAcIA7y01IPraGMVF2EO25m6hfkRUasDkzboGlPUzcpncdi3r
o7oTItvXaRKYzRqJYBxRDdP5LVowBw4xrV4G9WUq1W/KnlNlXEvaZb+j3zjxKAZsQWelhDuGClzq
hNKQE4SlO0zlfNYm0ktgqMDGiscCLK+/qnt7fi1R4+VpRBTh2QKUrXUYIJfqBId40nxXdFuswnuz
Ng3yEMu9ROEyl1v3u0e+J35qbUA/mJ3O5IyQ27NkroEQonLdUcFHQL++vhSqwo7BE0j9KXL6t7GQ
Sks92nsf8bG6m/t3nI0Bi1BiCTm9YzKp4EurXzuTUpgKhRd6yEZwYWqb83DBAUWpSyIJuzYLOGBi
Nm2IjgjM7lG7gM+X5r+lBrMv9NwfvpIStIn0Ykiaej0q6kacdKKcQquXwh6k7qlwrpuvxrYB9MU3
Fgyf7vZWLOkmeg8mUb1d0KZa1Dd5uNZZdGAxSW7ZgM9OwFO0F7kJlGDGfHxTAiDW3fnSUIlVYgcc
96HeXyayQWzonETpf4FzGrxHZT9F8UoTlvrRDrCra87JkodYa1szUoWEQ20JRjbJB/t98OxmoKF/
/nrGT9+YvPkB6/tgYm9a9PQlh5Qv2O5rUWCHB/1Tj8CUfmeteCi7AHbYBc7OZGgNsC1tVWeyeMAM
W/wNxrPKtFHIX0LGl0FsXilR2pJns4vauST2aULpBn/oHp3iQjSiC26MM4Zwy/r2Hv5jtu0vkWRc
lVWMGjLgN4Bckcz6raIlJd+WjlQ+lHlO17SvOqmKvn+dgYtd1wm26jyYMnFZ9GO+1OiZ0nFA64H7
4BQ8NaNXddPaX6sA2jLvcQKJVPjvozlc9/mdJSH7B+81iLpBZ9jWsrp7ln92uSp81t7XYlQV7GNP
SeiDp1+F4OMoAHFS4OfG4iFUfXJnlul6N0rsqXkydg0kWxkhbqxt6Qa6PM4C2t9u5Yw1C+S+kTBt
sVRjSEARCwRfyNDUKyrZCFUsuvus5ft/Ff0CDaUNBkT7omhl/mrRsoVUYBRQsOw+r+8alxxGtA3D
lFCc2TCdvqxc2a+15z+VnekTIRDgQ2CujUo/dho2nRBgr4/3RZX1aS3oNTB5aynCONFKO1SL/RXf
wIznNntVsH1MPxPEX7mr8zGduQ7qLgJp4+AUuQzkWIUYTsE57Y8ESAHtgQx/zc5fN0efzwXyGkm1
Pjc/c4nttNO81OcCaSIQLHcDWsa3od8aTbdiPbAdGi7Hszeu6vGC4WRIofQwoQQi8PhANCzijCaN
jE1FTVIwgst2VQaWw2BBn3Fy41yUFIp16rUdXFt4JKxYEYTxAxy+EWLAdNKNemSLZyzqLIrJ7nmz
Xeu7Zc00MWD9vihNTVL6ryJPZ1fpzsbZo0bi0iHmf4utca4q+nSlfi0ksVIdXXJhWURmOulEgjMz
pzXWNzUG7hh6rzwLA2yt2hsYtbY00glQ8gSS9odNrtZD2BQ+SkCTUvisQkIhZGCXIYYRdpKErU3B
v5wSLkQ8Rg1aFneeRo4TZ+cFTVJ8ouqOfljoVxASRzhGRMO4Lc0/Ut0xmY98lMJnescFFMVZKFTR
yj5zvyPzlwVN7KI4o52C0EVpyWPUtvlHqCaDV29XIVIHPaaQ6DK1VP4AC297HDVLROLXR1KHSClG
p+BDkVFhRCtDdXlKPDuSZ410KBuSUqZmhIngWs/e5ObSNnnPRaKp21ZWL6QoIQc9HH96mB9TxjGT
XVbz57iKhiFZd0Ooh0n4QF1D5kaf9CgqqQaRb0YwWxo4wU7Izwccm4zddF9forBdJZmiOwhrUReu
+WvjOFY7dKfB8xLr9YS0OBPCHUpRJaS4uIssSrq0j46pivrT40OChuQGsoTKWL/DlaxPUL6N8pkL
DgdkqHYbYBmxLhiDkBQuTwypG0Oj8s7/WDzOiq0JFHjc7fn/e0V+36EILJ+ElA6ji0ao0fY/tZQ+
3xQHeZnDMjQrtdSp83AP424RZqXT0qtE5NH12KrfFOcA3iDyGuLlEbsmsQOXr+AwNwX8QNNi2ZfC
/QrgxxCqIyJGPHeoR16QBB9fpkF0iqEtWfX9CWXRT/LCz1XVYXtH4AgTi3RO6NCRf24iq5etayRQ
zE4sU9GfkzXAJ1CmTz6osOQ6642z1ohyXdhpbniswOOOA0JH2Aks3EMCmTxwr1Y2lp32SVceDvJa
WhTYeEHtpA947xugtiQw+Fq5/ExqPihwqMdiTBLs63Klbe6iKrQn0KscbLjTHQmt1/JmOVysqyXR
yulAJABRDoT/6sFh45dRjiIB6qTXNigS0nESLnCkK9H2c5YhUliZevq8AwL+GWKWZhZp0qgVF1f4
xoLcB0IU6xJx5wYRAZX2RjJ2gdIprFp3qFl7IyMzBHbbbg8Nszc6F4qwRgNgSyk6tiJ1U1B2jQ/I
dhmRwiaPZ201X2TyR3Ma1VonPkElPIXEwoszhWqWrusVT0h1ubv7i6CZvhA8r5CRas31hVOFu7Lz
czXSpksI71T+8FUepCoRVxK1mfv7Q5Jqz+Gimd/tflCT/d3vOiBGTT/MZ0QWL5VTYX5/JjPPTFQD
AfqdpfzfcyghwPet22zouvEbOmiojapktQiduFqix2riTj0GsAOGibIQOB5OxSMVVO735Izzw0Sy
VNh4GEkLWpkUO4Awn8b4hRx8Dqe/OYqhNDQ/i7SNa9PXGdZGAhiilv5WSH0tI3ZaDKqiDDZiWO8n
ggLywax0XRSdvg37xKB7qtJLEh6kQ3JzxHmOVfSraFYunVDJT+hZ13qvLJ/H7gXndOS6jmFiIDwt
tTQCIL9G32HhXLIUFsWrc33ohscQ3Y+CJerSoT1FSaJAPtvqUg1bvex60LSEMzYktggbLrPO4TFe
XzKKhfmM11ADhF21PZzK/LrWWlyDLfvHXl6F+sUALrkVUg2c7BL7xcVZ/8Zaha8zsFliuo2+xj0k
+CT4yT7d+bH2J9iSZhlc7ys2OmvF8NsZ7QZM8MFgq9g1nJSGLRuWRuTqLsnbxRPt1za0wptBuII1
Mg7JHLYZwxjwk9DeZzNpC3aFdm4joELcX5zqvx5NVinyk+z+41K+4B89vOOT2NMCt8KYw7tUkUjj
SVPTEF1VZpVtU+M4WlC505TXVW005myH4L9Z2NDglbrOMOzjudW0CK5EnJG+zJnJmDx9fGrlo7fS
wbtXJsKJlvJ/0PR+bN//70hb25U4Kds3bbJ81ilFayxcPYOW7ecekxGxxcMh9yky5ysoEQpH6dEa
IpZkIvkSJop63yd98idwPvM+up3UAELh5Ed2lTCEMBpI7FRsfecIAOgPdozOEHpu3HRSNsrmSNRE
/aPK/5TJXgeJ6R8OJf8GQ6067WznB+Mt9YbTQ3ldvkwWKTrHudiqSBe0R3TNryrthZR1GMpN61vR
PeaGMmLZDdo7AfDGqTyJkaij7ZelPB9PkQEmgzRMJwjrITrSMW0FYsWdI0pKxxwLuF5hmKoJnFUI
i2FjYuv+/YoWNYaF2cemw5qM0Hk3PZ7kQ0y9Njb8kWoiLG3vJ2WQeA6VyVLY+siQ0+id4nmq8N+L
PiPInEJpJP/2pE3Nn6qtTE3KXtEvTLhHhN9UL04f8XV0vXWiF40GnNSEPpA/TfyjdOOwrAaXBJm8
3lcYY1cTWARe9H2OTh20McDekiUphGquL7Q9gf1OaNjtt7Hsk8aQmB02iRhqrw4oPsvhIliplosl
R9Z2El7kIMqtkSaeXLvhDkiInF2TCL7YSdlyq0Sj7g5b9lhGr8OBcLlYB2ETJuZwkOzy1lKjnoo2
YZaqbTLKbv/ahIM2/Qf74RqhTQt7iQE4ez9CMkj/q1PlA7InyPBAfUmi9zcAQv5ys/10bkhoxPIR
TXlVQfOSf6Y+YYgx0iu8uzYlmU3iEIz7ddLIUGpfIzTOJmG0ne1NzAS2FkOtNzybWP+7wJoQ+RZs
EjTvff94GiLOJ3kQTPhp5JSFRT+z+aJh/PA/ORsMQT9oxzGleEkK2SoWsvHDy2FMHefGnxqau22g
c9fcBfLsJlPHUoatsTwLq76U6PuEl4xlJ2mheoJqxjo+0ZeGOsDS+CT9m4N1lv+niw0X6c9zo/PR
4n3oVCEdj44timEe+YhjQ8TFEPRN4kqzcpnyJBNzV8UNAtlXvE+8LCHZGiSf5VsBuTH1ryjLIGkL
1H7HxP7N3/LDClHgmnaUepu6ELpwsVOBoSQddjSguARgbN4R2ogF4kq9k0u9q0fttgH21PHgXyH0
clAs087BcGIF3Z2AkiQbxjs5IntKxOJw8Ygcvcp6cWTtMWYscTWwpSLjiDyzaKAisolTw2xVJ83c
Qi1n2ibpS1DViwti2dBzZoS42HK5k8GbiG5A1p4bpgR6o+CY/sLtfDR3mqiT+JIoba5NgfYJ5cRF
FWKkk3XiDvH7GvY+a7HkrBSahWrVUZ44vN7sUKKjNdZxINCF0VJy4NB8RYUioXxkWAIVkQRY/Br5
xE76Z/1xFenERMFnf4HvaqW8ojRokLTlwA3UkXue9l+kjsrQbZ76eLe3NHVz3kAs0IpVafUJC8L8
2ohNWtvUtvkgLnmbDb6GC5PTNcg+WqVuj9eFWqvstFce+AmEpBrSyvuF+qUuVC2CJnCjml6cwP1q
6msvEf3TsZpZdPOX0kFzcer5rwWjC3mDR79Sq7TN/oo6Cut/y6ro1q68mjzNZVlU75OcVrzggfUw
dgkW3Qm2AHxgCk9wHSWEUl5K9Pu0utuTuUxl83Mdxt1XHHxENYsm7K3+6FiteUqNmZlZpUC6jTf2
4HFdT+kvhK1CDQSNtLQ0IUyuYKwKzBddzgwerLNEdbT14GywJ9JD+s8s9Y437wKGdPzNtAtwA5NO
5sTjC4EY2RVun+WTo7yZVC08FWlM+SlkYWyhUbz/JphFFv9moUcdG92O3mp+HzkB/FSszfJlAXDv
+BDh5uxvB0bljWwBDu7HqGF+nJmNdFK5nk7GxkqccXVCiQJTkhk7tDl+36NNyhP9O4u26zKgpdP/
nIQWyOCNuvKcGrQFgqBhc0VxdZUvCHawund7+saHYZ6cVIOQ+C5Sojnl9q1cGn9j0f5da5V5eIZq
qpw3aamelOFA/V8fCFTC4Ui3Cu1jJO/sePXOGZIfgUki4NWoc52L011phKxRfIUDnqf/2x0uFI+y
kpmDtslkhzNpEUy9/BUk4WQLuPc+Kr1CeNSvthOkNCvr+fs3/xymtlAr1+0+nKQhVNQLYDBFCsTs
5r0Ottc3hczhuYvhh423t3UCfGjiGwcu9L72txWIpO2nw7ZF+iwhGJTToeodHiKdqYUMt5dGTtha
5fBiZ2Z0X2QuHa+VxfXeekdJ096NP1lWyt8PND2Oz5Ubjzt4+aqWKt/vhxFUqYhKX9RoyCsH6b7R
K21FhbP7masKZGAxvt/vAgLQW0JmeaLqkxrfJEP3fSu3P+nPPVT2ygjdKjpzG8w3ffe2G+njq+4k
ROh2MoXJpZxEFkWk62FB0fV0zGrODM56v1GR0V3SZbFFCKfEDLdm53PQ9Sin1+tRmTrdT/1Pi6nU
5wNCLNLLA+HHEoolXHN77dClyadXYzy1r0a09bocbnRSdNlzgmKDGYzuvXa9WT1p0CktEbyr9PKS
fBNqzWLp+uNPAjz0k3Dxo2O6MEfENSQTNVXaZy/v7+HtH+WUTixy8zUzMf9KCrV8bgQE5sElj0C8
nwr82DARHagC35Siqqq/VKjPUUEHgwIPW3EduiXisDUmu74E/adfRbf/UbBmjATxpesqlVXMxFyl
IWvtV6cdf3YgBmdUk3DQQdrNk+3X5llh0NfNvvLtEpJ51biJDCs9xL97j4k3Y0poIiPrcyN5hkaC
kCgxYGAjjXiFGp75eb26KzHPXnLGTXSNqluZGqUh5g7GIlH9B7uH4SI8sD60qdHw0DJ0VYVSCHX6
wrB/TJEn66EaKcxJMTzTMyyBgy5ksyStp6o3tDmnHWmqToJkquZ/Gf1LsIuBIEV6gvxvuytFRnkO
7fIXbl9u/xCwXgWmbXxvHdH+yQac7A+39FGJrbH4WEQ6SMpEIQEsoBXQ9Gxa1fzb61X3tGt75gPU
kpDp3MC7Ax0tDJhvzkBx2FGczvJn+/QUpnTSBxsd0IeDSss7P0UW8XF0+cGXIPK0UeqU5ujGALK7
+BnlBjBv72dbPbBkKkUbSp6nSo3nQgFOFufIGk+UBtTSfCT7zT2G1y2zD+PgXskjnuMMlwkKFVGU
5aozUTrl4lwtUsUqbMfRo4GAa72Kztlx8XLe2OkxiA33b3fRh5cD7HxHDDlwpyEZgiZpR869yqSs
ezbuqSUVd/OF6l1I3wlYMulQPrXFssYwUlYj598ZCJNeFGyspCGVbe2WRxQxWihVkfIruezGvXnu
++no08TgGlHJfQuYOCdTLs1Nt9Xy9VIFasiVVfOE58LLPGbf/ne6t534SlUHzvq8/n8cyHoylMIm
r9P4uH2UiFKJaKlS3bvqABd7mDG/K46MM4qID4E/OJ9ksYP2I6A+K2qpFBvVb+Sdq8qHSgsp3z+o
fUuOLuo3c4o2RLPxcVyPfXzXy/T8Dum8pFa6bj5quN0aWS5vI1I9V5wHIYDvnc4K93TVCFLtGDDS
IKpWdJxhKZX2qL5eNYD80puek2F+NoaZagg0UpY6QOV7foPleaaPvzqWa/z6PRj5Rs7J34pupB7H
urwwue5fY7DTUjYQkfDhbj1Spa56P6YCho57zGXgzYyBicMIrpr4nYq0ux5d/IBrguTiyTuXKhZC
ek0Bp8zydr+g73k/RYaNlzl47pDxTBPH8x6WvAoaARkbwU1dUR2MUt+m5tRzMfnvXAHKkGsCjSrC
cV+gUoD7fcRNEPW7VsB322eYG7vNSb69mu9uQKBPlpoual7tGkhW4Ug4nT6Cc++UwW13GrukSd2q
Aw9UlP8QcV2VjKhcWzuz6zGGJ6WweHFOVgEUpIiIWIj4SxOBkoevk8sHmCOuk6Q1Xzusva2pP4t/
IvKJJhoPktndHXrz6o1KJD1aBZxzeEBtQnjZEzbRSoVQBdsSPKE0NAekycUx3kGRYu71paVf7Tgb
BATDPVIr7CTzJlMlpd1Sem0i8m67WUOzLaHB6n2D0fMfuWj+HdDCSNNGc24oQOOSwMTb+egtN+qC
lrDVDtcFK2OWyS8MwExvm0pvBFvsbCtyUIUhTm43MIb4wksqpQ8wrXkNSX7+Z7O034pkDnRF0xQH
YS0z+q0Vut+1VDkb1Xukn6NZ+1xRrHx/sJOgws5CAiJZellthq7WbC8g8m+PpkuLovQ1MU+jb6Pr
Jmot2/XF9WhxXyuZGwQalCiqoLfEoSk1q+gAcVdQJt0+6J/uCXVk8mxkHyKqG9t6gc+27i4fk/Fa
z3poujOkvKHZ7RDGiKLGxlx7EPOlI/2hwsN1l12aiSe28uGoxkG4JlaZcO3h/QRCpj4Ov21wd6J7
gnZjYmP60lLn0yrP9b7oVwJSi83XpPwcMXyb93S/fzpXjO67ORPRiRSboHZyuf5xfqPJOWKC6faC
rrbHLnqWuMKAaWVavhR3UoseYuZ+K2246Mz3c9A74C0wTHNEo0k8Fro0Y2Y/ws0wrvsX1H21NLVV
I6bvmdSupOdTWR7DP0Hxe2DB+vnBvEouAN/jthFG3J8rsfp+85+yL3kkJa565t+hgb4PzttpBCQW
T8BOZy3jCZAfLwr+QvAhm16UvCFG7gzoMstQ6lBBCEXFyn+d/ClXuueG8Mo/yScxOD96FQZJ9HTk
NFveKdyyBhDOv1hdAxJGlt/4rD2jJSmx2GvIxYhAVHYbaPjuIbRLgM+qA03zYGXTABdZfpUw0khU
wcycXoGEa+At0EZRB6/5umVMMCp3nQjDv+G38oOgWbew0hds+Odh9IfLWz6Ygp7NcP8e02iCxqK6
yJ7YzDS5uJqnZGeFy5e3DuIfzKySGPDuTeL7ivA/BCZiyiQxHa2G5ozAoCuSZkLkpPQE5hN5N4rx
pCTs39BmydGSqMI7YTr677pCOn+0tRsWQ26ew4zaT4C5boWFjd+YHtIA5rvkKlY6c+pVIfi9E77k
QcgEGYYEaHlNgZUG53sAARgmlgDo+f8oRHjeg8f72+AsGOrJQWwnMxeLlNMQgR2tUBx4zp/jd09u
FciGGXs41UCHyS6zs33ue1nrMTW5gSNmidXDv1dzeLc2haxpz7MoshFelxOtfmawG0Lw7z87xlPU
10XEScUfeHPlSAJBxu4rpwvz/qEOv1Quh2TUV7nhF8BMrCW6KL1nzZ3vnCnbU6Ju2/uS7n0sgyul
CIOXqqNO0UVEFrEUUg7WUDiwh1fzdj8Ra3jV2jHWm3tzbVHI/uwmi5wSLOWO8aP/iQEadATQekh5
I7rbkVc2YlsmS62BnuER3+RaWVA8baJUAfL03OiG2S5oFL3y0Ni9N+sQIyYVbEfoGrkGIfEAWMIb
AMJuQRzKdV6aDWrxe5jNcg+FfX6MAT/yt8rmFOYSGQo2xPiSj+z06gUleo75mpqJUFzBCZXvHO+B
eyR1ArL88rqQSzm7PnbF7Ftj0YjQF+apoQjHr9r5FTjYRgLBhVf3Brchj5vCOWYP8jgIqgpT5s7b
nV0Ousc1pTejGA/p/vRcB0yCXae5nnaPXk4p25CoUE08sFdLAwVsoP2N0jBDQ9l5eCGbvC65Hj0r
LArXjLl8s1CjPObeLc7w9WJBkPRXSRX4FoNkbfERv0PRLPDIIagYhmjZecyakT18GcADwoMrAi+g
pxC9jiJfKnzDUyVmL41h624LYwqlnuIWnbeR05Z6MpVwpUuScoo52RjUF34w2h+IGgmccX2pYdts
QWJZHkvHiyP6f5BVaY/x2MkK/K19seOx462sUf896Q55W3k+IsFEAJwqL7MBh6GjcKQ8GFRVDbR2
CkBDgR3ca+zdRgqSua1XJ9xK08U/Tl5ZzHRo6Tky5mWUJINCIv+Cs1gpw3/tEbpNdwePKYyNTQLE
TVQayPFvAcBMUvaP4kRWmmlwTXIAkczjysRM7ZkbHlc4Hx8jEpP13pu1Vy4AqWaF3oGgWqkHwEbI
iEzXBfXo2byY8udFtMf1KVImpu/FFopwkTQIYdFykqS/jxXi6Ots7QmjlNO+C7lx9BJRds+3C/HU
HXWHkT96SxJBh0vFbiAz9JuHzQSQWdUs5lHX9oNC8jmC77dl933zwZyOHEAgO1WhaXemfmnixnie
Pz3A1H00cLyF2f/CTBXhTVSL9aBAzERhhCgAZhNNBJydECMSxukY9rVs9IWbX0OAi/D+1Qgu8C2O
4pKWFtuZDgsUpwMJN0Xh3E/sXM00zn81jnMHiP9BdTgwOf97j7Ct31FwrAVejVW6CYetSVnVcKXV
pff6p94I+z8sD/aKeX+avBuZ6RKz0JCi/FYMurRQfqvj8ucSjtliEyYQnM1sHjibWbpEqg4VrU/b
2bu9465uVAtW8nCyvFm9axXWKF0WMk8ren0EaYqz63iOZPDHgytOIw7jWAEsUVkXUUyjz6H1qdUW
X8ZTBlHbBfRP4vq0n3ryIdM2GUBr028WcDWXe3K0lolHi7C6Zin47umaYFtbnkNy7/deGRMkCYDo
swkCEUkfCww3v+ZXVq6T0PnWPKy0GzydwQhBorjwEY9/7f7pD4MKQiZyRAONihAaX+JFwxUhkhP0
vFJI5gDJkCJa77wixdCNeBsaDHalicMO0XDeWR3P3ZyBSBkhFUMMA37vy4XKt5y5/R1NK9DOJQue
zYrkfOp12UUfYO7A3/xCjZHOolXeTMyE+vyrVlrQ1e5jyrOWSe+X/dr+2jG0AUvDdCMAqiH9fTN2
Hz1QSTef50ScD7+JSDlyEsM741Y3P82gblNlbwH6xH2aE5y9nrsFh206dhgDqOf6tvTAnCFs/4l+
LiAKJzqBeew4uf32yBlg3nfU2voeI65RIPeCbVkrNJWDhaWirOrzbmpvrhVgoEVguxYQFOdC5W3u
NcqnbcXorzAa33gq+IO2QWV/y9vpud0lLOAaQ0/5Q8AjuQa3yzu+VwdKfsNB7w18VrToSDRRzwoX
nUrQHZwCOWRwxDTiHv5iezcYgoks5ZqsPWz4J+txVYXgGDPFf2OLFbWRRsdyDwNdPLcbc7P4S30x
0LZ7hWT5ePF4ctz1wnzwrb5Rpq88QUiKJBKz9zQt6a4ibK8kR5n3J+fQ4bKV/QBXDqu8TGFU8yjh
mGycuUvYHkO4W6/gBbfVxAzKe1joNx6uWcZSelPnQDIlmbyb3xJHI7U7QPyCcL1dyoaG21ye/Hsb
w5wZtWXYbUntDzdTIwez6fDl/F8BEN8ihm+esGn4ALPA0iFFuc31y7FPkgd+/iw+zq1tEWxeUVv3
aaen0HJcqLx0R6pgnbU3f39znpSdPDqFKRd2r+uygpyB9aLmcW+iGImm8ApEcWNPbyxisWsTK2s/
hrhM2nWmCo0q9tPJX5rZTbHBjl3Wm/W0KlawCGJDBPfd2JOTh7cSb1q+x/XzqrstIoVoFQ5otiNi
/llml3qNiwiDpJOdFYAvG7o3EEQS3+UYphm50K2aKeiPKWmCNYL/bQq0jafpd8RVC+IPJ3dbBpjc
GXhOhDqYen9bwet9LYXO8Fn4nFFdb/CAOEwkuPKdmQd59C2Qh36bCiPRc/p35jor68kjZ7mg09cS
YOm8CaQP1wTdLav5iOPHBxhIWyg31TBOs29bmM0WL8x3SakY5rKACABZLGs9sIqtfzP7uc5j8j/c
zuuvcvCy7B4C6aaCA/hGxBB99xArG14eKEWYYTtuz4QBCrX0+OQzgTN7zBKMt59G9sOwxQHgs7Oo
mkv9coTNY0SIIcNAal2j3+H1Ddx1XwhS2wIsUX48bku7imiB6Sw1icb3Eon0Pfx5EtKkna4OY1mm
HdQ4Z0G1Y9e3X5GK6bFFYV7TpJY2YpxbUJDYrF/K7SzYav80vpDQToZsYa2IL59WCewOgkw4k7+K
MT/T5QQJMY1kI59hXiFN/WFtGpEbjGjrROTGt+1WHAdk/4IfI4udl9qccv73K7w2q17DDp+nV8Ev
55BWPhYxSlE0WIeSkdaq1Xxksuaz7Xsp8DiSCc6BDQWmxGIVOE/AqlFySKXU37VCIFyUinRXnlgN
t6EIcntEuPx1arJtZmhngQE0jQ5+R+VYh+eZWJnO5vNgNz/0WYRABhAp4WBhZ5UexUMzoYHPjx59
p+7ZFVvkVrlUS3RGJQJDLnqaTkE38qizk2xjVvMj+hjRcHPDRmr98u11hY29z+cblnXZiJ+hPZbi
cN1g+8U/6B/FGIqX/IyEr+XYyoRIYDfQlBPF2uzJSeyTdBquWNGmnGUWZgSHeW3qsVBgS/7d2ein
hamgth/yUh+3FUqyQQbuFGsLnVva+/V/Z7D/8EexpoB9ZTccAN0DvOQW+sZDk8vjWTxJjrnghQ9g
OFzApqOa5TLHX0GZWzP1a6A8En/ErAiJcIDhdjVYCOqkW4JpW48hgF2ErP5YW39NXEhTuBlK3NDS
eF9pKZPxFTPku+aDdVkwZu+anw+Duel5hnbhuzmiivCtkhB3RNQSYIJSXbkIn1eTHclRtIgO+uDg
ihgF/BtHb22lOwMshPgG0tAJvxVJGSnNGIWYMfhnV7yMMR1yQs5DiX3gOZBoCAG24H+RevnK667i
JhrvVxERvlBJfam/LVcyqvYyzsOkvYT7xpPRcctPe1yeplYCoCq+PKTT4ti6HRmXbK02O3S8CFIl
IA1liKVcDStsFY+RfQ5KzABr9b90jsblN5Y/dCQkcBf6Hz78wQCAug3VtWLQuNGWKSJH1jkMLLYN
/X8cJ8TgL/22xkduaePunpXmUxhbsyFE5CgCUA39KnVuO2dxw7RHkOoR2Lsa7jQYy/cCE6z76TdT
y3S1Hp08wCANlIa6PJoJX+fLFeXKqGpWlo9Ry14L7CKeH2Xt5n34UyQ9Yrf+xeKovONGd1P5VKti
BTOx4k+qtPttZxP3J2ATEoZiGNe3xEUg7rDDdQ+JPQvaXjX00BNyC1djPBgDFKAduQvyDmdaOMC7
8GZSzX/HiXWNqfZs4zGDHZ1dx8PXd1310vvy2cXxncZnL2xi8j+X1JjTe3C5qn1adDK/hPRFaeL3
ASpeeB8Ocor3B/WpwVITcZ2sBaEnkzaHp8C/2do73ItujFLGmt+VBtPa0HB1K2L6t6GxWE2uX4bT
xya+tjsD9SgcHkf519HDVlq9RsXLtn653Q2i19Zuu8iynAv35ZOM+Dtj37rjNpGg8YJT7+fGR0a6
6yUz/Y2ngFnZhj4q3g+lfzIoyolX1ZnGjP5uMnI16ZGJah5OkpwRvAMI3bV/tAj1hwRVTe5mmydF
0KdmBiJ7+OLXJlbRJF+ysT/I5YzghV4soInBBbcKCNMwaoamTQ8WVvdb+wX7ZLHAUhA5TYEgmWAG
ml4uwSNN+1SbfpaAQN0bK4GITUvEqWYRH0rYwQ11QAjj3/BaHGlYhnI4a0LMxsNSDzKKKfD5SSXq
tH3fpP6sGFb/wExgsImV9+MdmjYWa8dZOXSxMQiptZlGSFlmGmse+Vrbf3NPiL91QmW7K+QIIycB
eF6shyBxlIn0mFyTDxTv/a6e/HVqvRxSgAQ0vdc8zgSr4pFNwtKARUbH8Oc4eYKb14Cpra6KBOsA
xd/Sju5pfpN2RIaiZlVf1jA7r/Ek5o8ErSgqdJHxyf5qNTwpu2dwGvLQe4LAi5KhE6NuLnDT0drQ
0HWuYt3/Fzrw96NWoIRW9MG2jNKqzGgmDvMsnfUqQfrBPL2PtJyYFChzuoVO5GokdKvl6n2AoGlQ
B5t80hkNorY7g0fe8DLv6l+L0H8cfv9tMOULKZ/yOK02UpMhg24LOJKOkOqCrhOiU2R8uJwXc9Fx
1/o2nGBwZYj92OYL4jqFc4QkC02OoaVnqWCs8wNWmd1OLuj030aksWYmL3aYgrlHE7AGGwoWB73D
GidaWhI4KXuotBG+8dtegi3O4XEv8o6Mx4WTohNngX7BuIAGpi+y5mk9e52MZjSCv/wSgbrg4IS3
jSSPrgiwtIM1cz0xG3lfZTvD0ajP+8Ib2uPaRz81iSY915wAxV+mveuSIRd76ZtEVk8HAkVTMSYx
n05hMZBzsFgIYTASzQYewrUhyP5crWdau3sJTGtdPNeYMosmd9vsD4es2sr8c7djEoG5uwtnxhW1
oMIKSVag/ot9TxUrOaImtpva7KoXyT1uIzTmmsGI8dOdmPmPjzm0wAZz4mcbP2n4iGgLaeP2w+VS
tYlYvrNUjZWZLj9uzve6glDZDkXZKEQ73efrlRr9T1FukP1HrdA+qWW3NbwXX4lulFvYHvXS+NMU
jS0tOGlPQpHWnDqahnIZoaz8XhFshmFzs1MzOzaUr/weKqhmGCez7cSh1OpQ+EzHJLk63/0G9U4w
C5A2HA9GWNnZBPp3B0iIvP8CfsglkNdc211xcPfbwHsPZPIXn2J8VzfVj+KFi2OVwW0mMIWWdFdV
PkVqo1CLebtsINYm3M0urkNMXZTmIGYpLQyINwITMM0sg4mqTn6n/GfmyE9p0oVj+Yij5e98J9pz
R0h6vwzJkooCW+NlJf7Jy6YDhbCUgVQ9Rr/X50jW0jrKq/yv8/gG1DRDrVubN0gVi34vAxoolCN0
5mG/SgesQSdA54dX8N3+PANMwrHISYp9sBTh7upiJtv8YzL1VpM10rhDFu6QfKwtIM1JX5Zq7IRV
HWwK9EKOMC7141nsGiiR4jsCmK4VgdvQCZx5VI6g8fHChBpnrlQp0HwS4mt4H2OkxVZ1yFKpojkv
+VV0x1Jj55qz+3tMCX+bTAXZi5fA873vy9Yrpas30HDTswUl/kSqANvFy70YXGdbqaNYGDFXvxak
iFir88m8Rx1ksFFLGWxR9/nFFdi1nmDTRZ/8W2SBNFDFT8xDUlG35lW1pv5ra1g2L2KmAHBeX8VJ
HRtcIQm/BLn6xzcQ/USJpXu2zsY0ba8fqTZd578oJaByUyqlJn9SsIUPg/BHEMJmVTLw++G1zpWL
f9I+hlNAdrF/BZZynvq8uueEiz8iaaxACQnXMF40Wv33NG2d76mBAgl06yMRUqmmF/auXCZKZqaN
wjUVg7kbV1T6kqu8I89/NKYHRpOueVn/r2zrx3CnuOizsszRizYn9rSV23qeHzolfI/MS/OfTxm1
SPCMDoDR6zHyPwfW6Njbp7oituy0HVCPREMG7gR8/rQbPt2w6jzM94BehfKVCU9TbCkWhX2rbC1o
cR3LcB5Ib547jmcPf4tt1tD1hmVvzyQl6mM+o0CDC4yTaRvExcp8qF8pM7TQ011hNtR1XjbnDm7M
QxjW4hpv6Mxa5HR1w5w1WGG/g5V4ECOUfMUqErn6WUp34SVvtOnnjMTrDRD0gyImwraK1pAtVmOh
RBG32jQxuqUBJlHEf4yckdWh5ZgwDVUeXmFJqd6cbaM1JTBJeJP9LY5hF0EMhWtvKmx0dd396b2e
KcUW7JOzK4JJroJgTY6frS0F4VeK49njgoE39AWQMmmbl6sw5PgxZIUCJ5lvavh9OG94nEEIwv99
xTym8C+Lxb0L3XkMPbImNXCs8bttm5q8DegC1nzfOIO3/Tt3lLqJqo88H1WnztiJPZUsk+IdTcZy
h9dBeSsLFVfspDbDxoef3+WLZ+xXYnNlwcmec4XSRzqA/NUqqtgmLFlCKvzz/Fe5g4xzynv9HgZf
BPMOiO+yJnzlAjTrWTr6zNyFWAxNp9IhlnjBcWwV4ca+EiCJqcpF6EFafAdz3H+/MrBAUg+xnzQv
lE4Q4Zpqcmi8233D91M0R3Widt3o7ysb0/1SLGxymnKFxTqtozW8EceG7yy//0PZ6FABqcw/QccH
u1XTDcg6Fn/yzvfqLdbn2lDjexR/BTAOgDIJX0/M1XbG3XNedXwsEHS1SB+CxOjk88PNQIaWIM8H
K2/8dC9PibQ5+jbaPoP9JlTbD70MATsp/TplvJOOI/Us8tMGlED/+79tVp/v7SASJC8V0Em/CFHG
29fsXgIiJFj+vYoECJNjaFEPo3wM4wm3i16OxUSiDuaqOAnyaGrMR0myK43fD6fR6qmQM8zMwQJq
xajhCmgH7AST5ubnbRgcKb4JBJaUnG8SfOJBqEVAF6UfjCKNqoDC832Or2y4BJMLFwa1e/b/6386
8iBftGuwOTQm7TtV02tDZuXW/09S39A4HksKRaalLkzGVNAPv6J7jhkPFRdLRV/XaTPmmFy1Vbz2
JyMapmfC71QoS7ty1g1iolJ4/vzP54W95XRGo16ANlusRD6BaOwtXlCJ6jykmc68qFB/PIBTf+q3
ezIgXmCkXthPrRruqTKFx6aCI94PZqKnkXlOlanUZCn1XMnuVJM8vUCDuluLUJUgjPY7/8hNh99j
jyqx/Qu7/SqY+BB/wP73uKFdWGKgWUYxBx2TO5/zU2cCLGNhu2H8vfev8btxZnrMo5//VXHvFr/X
dj5gm/ImlQyXf2oeZ/vTUTzdHZFGY3cdRlawKAbON8QnOYYL7ys10yZ5CorU7lUI0Akl4auCosAa
v1rg3ye2giuhinhl64JVqEq7PIczD5M1XTBc8Ess+EtQF5x9WLj7O2VsOTBoa8wM7uU/oWsXJCK+
lSCSa62afl4QfONFszQXH72GRN692cjh0vDtbUWVsRxOq8StxzX+EHa84kQ6ROG2ghy968PtspUm
uZBhOW7dprdmNKp3RA2e519m1BBbTMnWfP59zhQik6gECeAu8hb23Es5gFCFqa5et+/XpNMz0K7i
9Tyy3Xb9mBQhJGpk/pyFsFGF0JMWdu2KA3GSHggnH1/HqCJnmlCF0OreuMK/k6JYejK0fX4yjJz8
pkLi4P9LzXYtJv9Fy+35Pn2CAM3FaMNJD9unKpNwbUKsm1Y9pCLW1XhfhZwDid9/jICyG2l8Czsr
/+dNO360qZ//rYupi3CNfk2MHMY5F0xfVNn6Qsdxd18rB4F3138zuHzTbEjRJT7ptdFLRbshHZr7
Y/dP0QyD6cqZsKsVaoUn4nzpUmEPHyfPhJUjbnH38J6iFEt/sLrfltDfbVl1QGPCk+pf4PvVADEj
lyG6Zrfop2w3u4XqrdHbZR1o55WZv8uzyBT29J6KAyz9a/BQHvghdLM9m2zEJyFDn/+euKLvotBv
di4pmDI0chGR7zsE7LqCDDW5IA1mg2sW5QthaHN4wCRJ9ZmXrQ0ToS9kNjc1hhX3pUtvlV7d0EWS
8rsQk3UDecq+ZDHQCLKmLi+BDcocWVsT4+yUiLfrrnsoTgfbHvsp3OffzS+GMrSo8Sbg0/7AaWkL
K/SRRPfY/TN58BGoS7c2tbNWWmsQkCvzIUkgbDjiG3PvmjTbxFHM3ct1N+68s8hWW1IezdhUddPo
b1ufaAdSUl9DO90SOfH08z0TsbJe7XaA6qpGJXKy+dARlLf6AHkyMlNPwKZzmG1YBO05u5X41jNu
AX7G/frc8RDu8kuaN6Ww+O3VYCkifTRalwFNx3W6YGzYhdmKBpwdPANXSWvCXa4PL4i7Ci4wfHlW
dZqIImRbFkfzHb/KxmMuk9kj8CS5SB4vOATapeUYss6QdK+RSIrDHGDrWs5Bvs24JRBFp8suMp6L
/1CVIwnsUedWYXw67cSgGUuwU4nYuSZoBX1xPLpYrE9tB52ENdcAzdAxyBZSGiRkYBSuWdx7o7WB
rBHNkVM+o6s5IVPnqK2goF5ot0Adnwf84OK3GKDosTfgAXJPvpGX/qZiYrPyI+pQ00+QD5xVB36n
28eiOVbm5pB6QQW38ddaLIEA8XIDOSQIx81pOYeI3BturrK/6jQhMSFoEz06wjaHh+EGHZWRpyw/
e4MgVBB0AzFPrfK0whqdwgVASbsS1543Cr9pyk6EXyNE68PiKUsSagC0F1k5Iwu6L//rdHDbxgeQ
fpUhhQiapJ4ncstRMlwdkWtz0l0IxI138a7Z7Z9MRNWCG7X8oP9sm365jriDkSUTa2BjM+MtWeTL
o8Mp5YKoRUfBEpbYY1chv6PR9LPRgST3wi9u0rnRPU0rUmZVQiGGUAAE2ytlOtKh9ofPC0s69SUf
+GI+siW2UyOMbvxYtDjS1rGoZrXHv5n37xA7WwnmH5+Hc4WD3d4+8EaVxMU7AeR1+0f4e26dTipb
rH9UGwPXZS8/k6nS20He6dZFc03P5J1RaIXeMNZF+cnvPxg4hPW0OQyC7g4+H63zHf5Q7rriwKqW
nSKfwDxUV0Xfhytkq0jdBCP5NvP0oPuKyR9zKTivBenFdcTRNDrKSFKB3KdcdbPNeVnzgdjIi7Uf
mF/KzFxOCUefuknNj1pJbbPw6ZxROEya3m/+njgYJ1VoK8Dwyaia+lo9uB9M7LLNlCJ0pVccj7Lp
3tauqpfxj55Q7axRVgyh9PkyMumwAMWRwohCqOAfokZCf3cM1oQAk6A0k9yc8B1SJV4WK+nqIYtb
Ab0oAOyLTRMWTEAqlgqeNC8yXAmqtQO4exYNBW9VoLDq9ttHsP9h6tC/Q1sVd6DQLjmXNmSmVZZ1
tMnkAWMiN4SP12yStFTbHIsAdyCOrVrBgxRkPf1XAvmlHOWr4Fi8xZqsd5RdEphxkY21lj69sxXb
X60XFQhZj94zePdyWszZSstLIv5Jd4ZGgojkR7/rJy2DOK6287sPlfKMiCm9r0mJHcLxY27rPIdv
F8zGhF882lQSEXspe1AEIHzb/0N3ui/kM+JshOvym3L2+a6owcL1G2YRMm+Fd1wKY4pRclptO9vE
nmXUHq7NIkyyNIJqgZzCP5FLrhmcdn6+yGraiZr5Haz7BtgBoU7peBqEnV3MJvgpChAAMc1bJ2CC
5cEAGjENwwL67pmBMt30KLqp7LJ4Pewo01jxDt/Sqd5YATf9RuZPLAf2iduEfth4rot7S+GAFmV6
QB5etjv6c3lEe0m53S5KCvUyzOD1pT3CmwV15wjxF57JSe/hgM4ew13x+CI+AgYUQaar5SdsheId
GGxWE+96P6xDPR4HF4dLRdLzXbI9LHMl7dYkzYZlyhDwvKv3uVUgPLnxF3iegD171aRwDBO5BrKr
5z5zah6ztf3pp2nUiFcCmcjnz6To6IMi+zdg1815GQfvInCIVBXrqWdzm6qNjwcbAHhh+tgL3Jku
CMqlG9/xgLJrX/cXt8Gxx4ByOe3HC8u9T7x27mi8hA9BJkCo0555dU5X07AGC4mgFdxRDIlVv3cw
SxTfgJfcrMTqKtfvj2yJ/+B9/3RGbpLVmP8ZwWy70D/dWDb0mQXwGS9XT7T46pl/X4NARJQYzdb9
eiHVpkadxlgzBHAUvGrhhxVTrJENZkzO/qppOg0km285UNpKbIDAITGagz6E49P7G61cEYDrroFE
KuUIxlrReYdejZIVV5tbkhNR0TPWd1cFlnv8WJMKHLIl7vOBsJn1MVvANxrLI2PLH+jb2+rVXjNG
hZw0szO7qw9Q8u/IJnOrJMs/hfdBoFbeJqZtZJzargGwodpa9U6LwoVczBmejDnX38EJUC4riL7k
K6tLSALarGxMsj9c4M8V3wgGgW/5YSlcXsbKtqc0+agGG1Caz3kCl7zMmtfPEPXKG7NLxmCQfly9
hYiJc+lb9QbqgKq1YWj82CZsvL4qAanYkm5Qg5NN4pplA99bqU2Zr5cFUs6iLYQYACEk7CUFsUTL
6D/aQA1MgkxxEFRoAJf9G3QanDKb/KiggZqaNypVyMh3oz7LoBlnvdoxoA32X3Jt4hThXeQIGSI4
eZRjSB2AgYBaYXccySOflTGwLuLA2Q8WuA22GWaa4VBMbKZCDqt+L5x07e9mmxqH4XrKerR3OiXW
4ITlHcs25ZMHVrNCYMK1led/opfAu9a7JfSck5EkfqBnnxWKg7xaP96TIJivr0ER1Db04wiusGpF
PxmIDwBfNvQZA+d2UeHL4NTU8q0MVdQFdakDnLyZxKJ47tMYxV5LYQMq2LiD3nlUHWt57V+1YDnv
3O3j3Kd0ArLtSLY+Pzb1kiYtVXhqZx66RB1Dj0qnyvN03sixN3J9Pw0jViN/mse1YKzpIBptSSgV
DdDI7kBdxxcMXUc/LmzCeeggvyzKt42pIorZpSOIOWmAWsWhrBIAFQXM47y5q1iqxB/vmvdOkMhd
Ib0GgnfAcstGLDf078DxriUqjS6+o6W1MX+OsusauKr+Flqg3JwqjRRDaftWN/pRhOJVbrspTlTK
SkWjglaOXdWgB/qvxrunDVgmyI+fSQn2tsjcEgPcLVDVG1/baP9uZciMCSTI6e6MX/3IPFXrTIdI
UU6iB8w/mByF6EbWNYnksEzoqwF0O44+dN9Mr/ZKU0f561jTEULlum/cd0aeK/PTp/+UztLC0IJL
G1QPKUUJ+Iow5l/CFEtPjkGJq07/BmmH7bIhw7kBFSthyCyqEpbIsCz8g8Wfhatg5VHKI/J9YIXQ
ZfdjKY/OuekZjB/ooEgFKhdgCwm7p+B+vhJz72VGnUyIaYS6KqdaqC1qf5Xkn1JQfLjhbwJvMi4N
k1MJFpmgnaXSWAGdRtjtmdpLEY3WOLX4jWjoOec0c69YUxms9R7p3v628CPH9cABGmSInelHgbtu
ZEP7mn5crglMdyT0wO6VefzR3vhRsLx0fEII61oazfqOq+3hiZdcj7GJf5F8/lPyqzc06FvxCXTy
ooNfxmG3WU54+y0qUhShNxh/UyhPGp1TL0lbAeukLdD03/VAXxo62+poOsha4J8I+T+w4IlIhFGS
uTo41x4MzO7ORprGrBWRg/5vLEewY0WfKbJp4g9US3CcdW8lXerdoJNjWnEJjP7dChpvi1YD34P4
lHx03WEoDwv9nxnKpn/ZUTY1gK9uk3lPPWBTi1vyN5Addu4jKA1jxUq2bypqLJ928Y9xYm1+XVBI
DfPhtEmOGkMCmc6vvCPOKiWZmmd8sfGuVGygszvGV5OINJMhXp4rQILVHxkN3DdDpSbyBCE7BS63
AIZweJLCDZDqXkxZBzQxQAYzzIyVC8A4aBCMHtMbyB8IRxN7GFPGH3n2LEn8cA7khQM9MPLsUnRz
9bMVAp7lLyQH2lbUwsfgz2BX4guaTtfgbkLg7FEeS6ax4aw9RB4yn+WuJcDtuTVjTLyqADPPgcKB
80C9Vb4BxN9b5Jx8dCt5akHw6TKeHzXrBjSGZUJPZUtvvoGG+1Lha+1Cl3W2ExpGwKGNkOmylpA3
jtnKfNEd4ZuHD5rhUmAuuq8ABFSpouCQuYNTXAd3jZ4HeyvaYDc6kA4+vESYsutI/T4vL1qM+Qla
Gy94ynee92lDrA+4qL57DWR9U+ZF6ZvpWPxpIxrZmBTCs8pGzls/8MYvMAJ7IcN7ZMSJhzuvyBgV
mWx1vVqesdDdx2OTRWtohzsjGAJQhSJT+pktgKCocgmDSKjq1bDg2KAOtzTcdYGEYQe6rNfjhflZ
EeO8T4dPfCujozO7p0Q/auSWcJ4mrpQ3KcxlYD0fd8291/3fpuEWmYdvFe4guEMlFbKyeD025zPx
ypmpZ9i0wtSPNPlUAqxSqdJG/qJLgbiGBP0FYY0F76aqZPekSqNKpLjjYb5iXvk5DeDJ75aDSEgP
yGuUPnEtX3uY/RmLF66VRIYLradNwwXuMM3u1E8CqZcJ3uqsFmO0btZBe2ayqq634BlX2kAdVar6
g7C/AMx9mv6cJyJkNKOcMw9M7tQpAJAtLze8VrQFG762W54EDgTQ8lK1FJiQPEkjg7jllQuETS8W
kA2dHdu1tCAqAHiMja+sGdwH6d0MQKg5a1z2EQ6LNBTE5oNhXVPnMdN9j69sOuFOaKqC9/Q0boeE
4NDeb6eXKUPLi1k+rmGDnQL2bAJ9ANMlKZ+reubNXqpqH66Xh2HonvvfVqqAL32w7LMV3pu1ZQ8K
xvBDj9MkSNgmt7y7C35PLD+GPUvGjq0Z5hxY4tpEDYCsIndM+9Pe07otFPXQopeqFFSe9mLJYjYq
6I/DT3Pf0SM4vHfCl/xstYy/r2DsVV/pmNF4tyvzcRoClml8Cp8PMJvibXyiZZn34ZDSYg9V/P1o
nG5S3IarJHlnX3Hl+ISxkfo8enn72LV1uNzgYe+Q3dFuudiBtiVaPI7toz2y+JgnAWsj3SRNlQb6
SFr6310BXVZ0uDVUErIWoCzuictlPkK0I7aByUYowVjoL5ZMGz5AUlATbI6CZGe58eX18bZN15SC
fT6njYNaC7qgvi+cnYdP5MP2rujZ/EsKHrFNsrtYPrevJ+7hUSNZznh/VUyMrKjjT5J2cD0iJAgK
IU57PoIX1kR3dlI3uyN+K4BV2k0+WsMYnTvYTfH731ADIr2aXdGY0CrB5y7NJWP3ZVZ+t5lHvcQj
O/WY89oBt1+kKYL+/eu/5VZuHsvwlbxK1HsZU+bHSVUImY5HeqSjGeFNhAI2fg0Nw/c44esNMjHz
J58/EV+WjmiGqZKbtSDt+MjOSvK0bgIQX3sak3fdjh/aEvQEUGSuQz1mo8bllaebRKnbY5Tsl2g/
h9PwpxABwelaSRMeSRN9TgZQ/hZK6fptN2lTQoWggyOL5YRX4ip38aoXZIBTnr94Qseb+oGxb1Fy
BiNLlmJkm3hMpka2J/+Gs+RDG8elO3kWsN4OP/6gIVXvlC/g9c77ssITB90BhSBC8g1i26LRoYH9
D/o1D798pQN8j43gVZp5PiGbDNYEAIwV7r5zQV4/CGAbfMnxsD8nnTGhpRPrnYxCG7aY+5P2OZm9
8ic/43ymF7uN/VpqwkWUesN7EWc83GNXo3Dbhk2B7+7DkJA9WxnOJvVy7LPXfyITwlVvOag8Y34f
pPcEYP2eJOQC9XYzYARYa1q0G5PNqhKoFJ1mRmzONGMK/B7OoZfswEIZm2i5IeWZ3jZiLjNUzeHz
4LmNLpwGnu+DPoBJoUGbgU7sduUVdScNWVGuaP9SEO3hwvHCBaNKw6PdBt8o0Ne+Iv+4vPkF1YiK
uvWuWEsMhd0mlQNZFTbu+pZFqRBUQKgtlxcPz5QUxIufzKqnN5hQB0um7lS7Zp0oQsvbQ6nONTQ2
6WnZm3g2U4SkKOKJXuoTw5QrrS5XKnj8yMgbVYnwd+L/p6eq0tr2wiQ9HQBwFFfJRwqtfG9rBsHN
wuKKgCIz82LRLD9PW4JXW6eV1EE2IQuaH/Wp99yzjSIdf5ELBn5LqKIr7S87G1MLRNHdpYHoGI7B
V3AgbVGVdNZ6c4X3BqvnBhaVrO4XGqQpYKQDuqOn2P4SSywt4ZD9SYJ7botTExGLnvV51x7QF97R
QZkoO8ClBmWjCtiLNddGF+b1VIDFc3oc6nXH7qP4guefWRPGupWZroHxj5mK2uOdFerPR4/O+tlF
d7gUjF0Zqp+G0yHoW5gemnw4BuU7SkcvfRO4GQD2py89WZZEqmy5CqSqE2aJTu9huKLcUA8JXYtd
yr8fWr1fTBc/FJY49eCY7GcK3AoASVA9f+PNmx2/pT7CdoWFm01EQmWhIBj4LmbqB9q/sSTslpX9
IciyAfIT9LS8DgxCoG6cyYsvbl9VazU1jhZjMi0ihaavf70IzCJnqBJh0ZRg2ng8Pi6Ouw/j6LdF
7zqtDxiclzJ1UB/jvQquitWHtGZUDNuSZtNgvwbeoHigRZBQLpi5xcWrT2l4SKcs/tekfXH2oy2V
Je+Bf/YCL+mV0wIFj/3ZvYgxJRc8wKtGGF7lwhRUbsUGf0SZixQCg/inRFTz2wjbKNnIKJg2TPLW
TIXFoB4BBzkp2tBJO4qKdHprezwnfU7sTo4mrdwz75NzmuPlNTS/CtWSL50JW2u1LvxiiEJWe0eT
kxlkUQEZVfDSLvTkJUDGJk8GrIR0XgI7jXgkFwPdj8Qfh2V/2MZCHHZ1NBo/hNmiVgZaqQi0g0Yt
OXolt//XTds7LztaUVJaeXSLM1Cib/VQ/sfPphREMSZgzg+D2O9OuG3K+2h348GPZWGR4kh+xVE2
TliiaYXsPVHFgltHL8QNFgys8Ax26yb3NMnqqgZZUsIT9BJ3AG3PAnCcK9qvwErf8kEj4aPgerjA
oPSeIV0CMMu40MDCOpT4pmbPnfBPZs6JmuZ6V3F+nUaiIz0lRKXNzhM+BI7O9x3gsXUj/YGMqjUQ
6PtRbiHrvv5MzyIPXovw5BP18W0ykVofdGvDD6WxAmquo+y7i4TGMvANxOWvq+ZfGL7UxWoY+HEx
nzq4/J+EPSt5JwoT3HipLU4zVa3Y4oWqQLqoW2CiSAh75wtkIvja/5XdL+CUE3CvzXdnDhfmbCAb
Y5txUVATscIHiy7I2FlMrgs+uEhyBVcfn8U6iP6B5F1a+b+388SYcUC9Zk6sWg1/RP54t9A3Iti7
cdbTauGPvORWAho6TsxIihFCmUrADVjhQvyrmYaDAXl/Sqg4PDVQCAF/S5T/74QwiUbyDdNQnpiF
AIuBcxk+57yGBZaNyXhajTNTK2S4tWT/+kQ9f+V6z1wT9nTBTtQQ3F92kzGv9NyT3DDi5/heVJON
15Px5EezgbQIcq9imj9qG7oaTY73dB0ASRhLQZ8Hl0WDjXUgYntcMl/yg54C5oxhUIXVPuq2abbk
sXcS5reFsFQ2WPOylgbbcBfdJkwfkHBv006m+gUKdDJWJCJROb6AMWXYfCkyxzpy7Aug2LqVtdid
qgNCnUC/Ie8NCoiZ3CaVjZ69G6wNOTWRKBSr0jdCOe62ryl1kux6gDXYMLFHit+I20quER7jwiIu
JvBsp7uCWIBA2UOmYTkTRT4EzZGw0yMW9HDtwKLDsllmWnHaEZmr+JymOLty3YHovmHLjRoJLJcF
wGr0iv/cMlG9Jsp/IloxderjOaTKy5V3B4Bf0qxfLUv17+BaD8AoKKr38rUL4d9Tqsv97MRFkSy8
rOqRmjznM+pwJJVLChTED+I9HkBUsAT8t8lREQylBM9g7wXBcsNKhw+QELtoTDz2b5U9mDrQd+Ru
o+CXTVdEw17QeaAIjUa3JLe3c0XV5S3EIjRYKXNc7yTM5B1NrIxnq7OcE9Xc9gitZmlgO1eRMu6b
nx99PxsI8kjyyF4PeLPx1tWnshLs7iSY9zruiYMiE2XC8eeQT66gvCAVKGTkMMDLT6irO4Faztva
jQqvoOdQyWmhczZBUYrvkNzAm1DidLiRu6vcY4mFBUWuwC7M4MbKaL9gy/lKgBdPRJhTXLccrx1c
4KXrBm57JEIWF0FR7I3xHN+wVQeTXjcJYU/C7vHKXBnTNWg/xBNB1OZtvWUY/6vU2kxFzMeydBjv
1uZyTxHENQ5G3FTFrl8c5Kxzu7QUv90jfB1jJpTvNIVnog3vLTjXnjdTj16Tmib2EIXO6BUMd5nD
gkFErqeYghfaq7dixBsRklnSrt6dciKoeWT5nOmcN2nMORikT08moVWplscvAEZxFW1H2WW4Us6+
WVgj26QzUe4uvEfz+fyp30JhTXWiDRyJby+Nu+Zw0GnfgiQD7D2NSPSDAtbSGvdP8mTOg6hyDOTQ
ZWn70XXzqvgbGLAXtRRokft8j7oJD3VBlvFbG7PzJQZ561c23W0uD0qlL1S3TQQ3KEktBNMmHrYO
n+fCTPZ2c1bRqXvwvqyS3+QB7tE9bKaJpuLAXko24Mqke00ivlnTJZirVMcYp9r5kuZwkIZ55q2M
d6FbnZtUeCg4jfYHuPujnHHdWvk/ngjtU3lWsVRDu8rRNMJlSuMaNBe473qktxab0NTVX9EStiHo
z9b4lCVREg8njHfF2/78uX7xziCblGAJVnEcfblwZdBk8Jeob2hoNcPPNKrmlh8KPucOZfF6sY4d
0f1/eJ0XK9Uz8caJWg4ZdlW3cIaRe+22wC5U2enLmRk2vY9NyA8qtuxMVupyeTR/ezR4ekdMkzg1
FNCDFrmQgmJ5eSQKhYKsKXBV0zpqS1SeM4woChMR4Uktn7uzhTt9v07ERGihhDe1J6LAYWXsTzM+
RbGckWa4WhihMAlN66eZN5MIttT07gQS4b8B0cnmB+DYsBc1IJegF9v1D2yEebMKcZ8xnJM+roCo
qpXATYfnCMC/OuEpv/4GOPRvy9vvu7prRekfz+o7Nx1ONZDOHmrc01gJ4Mc8G1JZ8/FqTqfQu6ux
P+9mFdx1Yip6ZcP6KgvyNvRxOOgNvK77qQBw76oloiLdk9nL91JZMeeWKgFpN2LFtmw3hrmyE242
MScxMmFNzw3OokxIXNXciwClgdiuFDazKs3I2de8jY3g58bYQKEvMYqk/Od4dz3OwdI6qAm5Rayq
BJCyY3Mt4n2VEZrzEeKCy962gHF/8mXShiC4MSqbZHQgIaO+8t4B6TA4zlH6g1H0SdIsWaPWaAxs
sIB1pWLPSLBKOvMKdDvYYBPILfFcIiSlm/D+mRi9Lbix9ll/Da+VxK3SnhCZCnj+ZMAuXlTC5jGe
XOVvXRyYI0aUTsvJpcpaYbTjUN1R9cVT2C3Ff9fUaAw2xlrplQutwVHBmW18SueVpb4fFXk2tsKj
tjZwoMM3aO07Io/CUTDMaq4E6O+D9fqAWmJtmM4JEtna1QSuUmBazIK7/IF1b1jIY66AM1xVaoe3
3A2lIdvHJcrA2NYPXmV8xCo9DWZjQkmSew37tYyCVincpdzsLQl833mFktNCIglAZRsYb3g2uF6Q
kocrR6T3IFrf0ADU+cn+A1i4woClbY/W88S3q7r3Auz4slyGdgsjdVtRdVRAvISF+D1vX8ayEZgX
iVelSMX3ZoaXEkFEuwxwdBI4jhWomO7tlY3MrLtcp46+0Ks2n3VI9gvjcGo1MWzfuNmnRuV7kGp5
MDMtAMPIL3Mq3mOmYq6/pQ2VwYCGHI+wu0WfXXPT40BqvrK2FtmrypjksvT9ibgETDrANjJkMzS+
ssw1uma/l5rsBQIigG/cvjD2teHiiaAlMxQ0ErFcEnb9JLlsDgO+weu3bp9VOsohUVbylHjfsa8h
raY3t/yy5iGuwERn8TjLAdPI+2fyFT4/P6hlR6a9kz6Sa3TUX2o+IMfC0jbpkOD9T9SO1flejL0+
rD1NADgAx2Lqw6yc3XI7rK9iOXOA91yLZgAipNxZMOBTcHWMOyn90/p2mthIHo3+jJRF4ycCkdBN
J7KJiyCy4FP9wS4QynpAx3LSN77VNyEBL68bFDgqH9Q2UOa2T4iGuD0GPLtSy3Hjsh+F1ggpsFr2
2d3nOut1SKvYecyZPnPACl2T/IxxTTg8baGNzF11TM9N7qC1sbdnUZEx7UD02l3t7KKCCFJvYNi+
pn5tsnbvJbkprivtp/R1yzvEkBGYbOIOZiA2UIMm1pw64f3524PpIn2UzwX/ZVBZZF6HBdscw8Ut
8OAQ6AgMtZl2p14cBdFouFESNueA20OXe0bnLUf1PryP/w0kz5rSyrB0MvsHqxkApeAOAwG6/x+G
NWacn3F5PZkcHe/eov0yYIcmI7yaH2R5HqF2unOBR0DhaA7hKO/T9D3vPjFU9wKOYcOOL1xQBOxw
eZbtBziYy8rh2vLuDtJARAEJ6c6+YoPBOrL9S6pNXUuAc1aWdMeoT8LcasxzcswGDB8gT1TyBZ28
F/VTEVmdbk9iU3c7CyVIT9nvMcasm2t5avrp8YdPJ/2qYm3B4oAdLd2akOIA8ta6i1Xo0XLPAiUW
C17VUig2igvaoMFX1iu7YRjepTr2MBntfAIy3icJtJaV1D6rch41BVuQKlxnLkEipvkkpStd2ehR
qJaDTOh5TSxL5/dY68kr0m7f07mVCQ0P2ARIWnE80aDrkuf0cCeeeDQtuwJ98BDOjZ1Awf+rlfo+
HGjMbrogm1F88+8YhkkhP3xEKl/ST1yQHP9qPU20hgdAxhdBf+ESRPLVEso6qUslG9KuZVXHkmkM
zhblE0kn7AVCdLm5fd18Y/ovNL0MWbpf1MDp4E4cxoQIbIGx1YTBc3OtL8doeeIzcNt5X5tPRN03
omfcpcuUdHsz5CI+W22OV8BVPur0B6+Svj+mUBRUhCRTb4IJX3SIPT7VS0KRuOfTVmyKiL25J8Xd
AvTIRL0TNCNOzIe4KAGcO4TujxHz8pMo+oL8F/vwarQlOuk/zbmApn1hIcKWYolT5URFDh/X6kWA
d4yFupOqjou4dszaDxdafpXmpJQeGbz63+U6W5vcYJvagbr1YrAXW9SBl7tyE7B4RAbSaOFhOzvQ
UzYFH/Fqz+ETYX7U0vev52pPtyvOXv5xWbs+62g9ruVhKhQM+Lloc+3TRsYZ3IfoDgqwYSWw/RpV
p61l+bq7xDialQxd16U5iqJNe01Nl0dD4Dx/fLovRDLKiO7ONVHmh/S4lmdEeLrFf+y+KLntz0Yn
KGmsjJn5CfIbEmdG38r5GB9vDxOcw7OpnCaUatncn14pYZiQ6+cJx55qpxVRDzpsxsgRPQ6Rbxis
8fkyWdjG++yrCFxzWmb+dtecNhOj2x+K2ubrYGbyzp3MqT8keiioF8O/GuTvBZZS4RJNnKICATIv
Qd8o45osd2GOrc0B/JGz37aHvjvsCz3jY43nt1Jrf/2hrXv831RrcXKyoFJZvBcCU92vfJunE/Qy
mlKQXy4Oy2EANjmGqIMOq/kinNk5ifLVZVs3xc9rA8OJTcBJFxbGTVr+jYlwORQ8fDRS64ckcSRE
jPFq3SFMvOydDg4kWmi5sjRZZjGlKzluAExM54XpP4rwz2/Utn8kndXwaXCE5PQO67CWa4n872yt
N8RVxOK4/Ns32mI22RPhSG1COaUzAXmIHhbHMMt0HD6WrGBAMD/tFKUQLnXpfVinamS4nloDk7qa
9t46oMtp6ianSGDRlBaU34vzOPlM2K359xjnV9Lp+yONbZUL9/MW9G/jAOwU90Ji26CUP9UW8CVx
OIeiL84wDwNyTFUMYjg5lsijJS6CVYASbgShOGMbpAmw2QwmAdX8IUXdH4dvogofZteqtAB22nu4
uNySOm5MYGS7wJoyujAWLV/sq1Gj1ykdb59A+pZkhKGyQE+PUUmiXlRn/R2lAb9+vK8+v3/rlGSp
CCtoRh3l7Ksbxgubf/JwtTzqFDH53ecHe6i4+6iqxkOxA7/KO8ldCf+nKoI4rQHI0dsuUwK+14Jj
iWcC61beNDh9steWEbVc7j+qHJ+LjeVDEu1yl7P5BC3Fho+ogSLHPSo2Z1zfppTxF3oFu4kugxS8
ylFHgnRWfJgKsHRPLPj02LK+HbgLX3F2P5h8meTTfnURuLbpCPUsJFKEPrbsZISxlnknkHHHukIo
zI1AEzKx8eHWsbgClT4dDH6eHjPjUfVXn2V2e6Mj3raJ2EUcN8vs8BgboVpJhdZJS8oUdcbqm+RL
UJhV6SjdnbkIZXhrLBaG8kt4dkLdHAKzvVb6LgO0gNWGDfcWgj0Tb84xXqLcZzbASRa5FGHa62I7
+ivHSbS1JeZVtEOb2pPvLv9M7E5ZqFjy4yZB7waemrtKBsEKgeRJRjWhG1MQO6urgRXVjOzi+eTi
qNDUvtq81ll5SsuvFZTTW970EBl26t9HSJC56KXOJLkLZUzePIIldE7cr2xHi/xMZT+kqLhrSdwO
lj8aPY9MRqhsdC3IZum/0pdCsKBjs2yIdjApPN4r5leefw7+FAspJz9KfRPm/oXv6uNSdV9O1k1V
1Pm9YHglitwLOVZAqQbrLvkjOLy+e4nLUyf+0F3/FVq9FEllLH2zN9ty7HpBpb8e1DqXmWYFtbZs
1x5wSSTy4pguaKNXSAovBKuRvGz+7IDWqP/YhHhGiaRd32he/fvRAhsK+J0RULv4BRuWP2BHEeuV
/Sq9TBf779tAPm1jWuI/pVk+uaauekfHDtQEvBCScNm6cS+zrTXNfxKlwxPUVM7OKrs4aZXvzkhb
998WAqE5WIoaTkIpsmiYCbZRyc67OR6b8Xfjl1HQS7EhQsHufnyfOkEgmuvuuT5M4VbHNyMIrxBW
Mfzc+yWU5sSMzII8I/pVW4LMfsPzqECoDjgwr7sMZQP185mYNb4ZEfjuRETD3TiEv4kqp0bzIDkn
+mgTlw0UJTbSmlK/m3ldjTi0tRETkSuyAHH+TPP4SJmT9EvXehuqW203PZ3aQiQZxGr5sJMtUjuD
6dJOVxdSamUFDWGc7tW/y/NSN8TzEeZ9CUSn6TVDj+nxykYmEN7CEC9TIfOeevMZQAirm5s5OflA
NNYwclXqMDrDIMUIZB7WXMEucsfPnA9+C2rcjcOMIBkvB1ba5ih2lwq1g8GHE4d6dlkGPA5tECoG
pgUYgRQI3g7ehxA5218ySLZkwLINQCB4NYS0uKrqicoEr9aL2sAXLaq9gLYvs0d+YnEg7RbZYY2g
mW4WL5DwsjvD4coXktPr92FqLhSiYWulmsC6AjpptpuUtORkKozEYT/URhp5MQm+RkekCiTJmQ+V
LoXXG6w3z5x+4Ywj3yMBY1ZlE6wVRU/vXWKkBJKBk2tnMjc+gpzoEDC8ZN/qVGsb8Eb8y82qK22N
l0uydUH1BcBoJ4JaPUw8XcFo1YvuZUUvhNfId6oB2jShaGd4kIyjvNKPTzABmMIcgkPIcqL3/EIn
s9S5xzkaqeR/vNfj0+s8PP4YPkEuAwNDSvnhXkCLmTId/Qg7ROSDK5eq4ryhtlfKE38X6gD9kS8A
3eF8zu1bhTRw1Kc4cdyALwSDcB6Yw7Wj+hT5mXNXjPiwt7v1t4i7aIDfwM8LFl/G6nefMmLdCoKJ
x28k9pnm5IrC1mChc2b5BR36vwVzMcAHRSfrU/ZsUviOpk2UUdXzoBD9kxPVWh0Y8KC1Q03VDpMP
+kA6GDtGaN19ZhBZ27xZd3hcjgxYTsLEvUbC4IlrSHTh16PV/d76N0tm/OwK+xlTVg3J93bSCsn5
lvq2OYJGB+aZ7snrzYCc60FOPLDRawUm52T/nx4ENsFbpvNp8AAzGST7hqjkFREYCelJJNXIctQs
1tnkx1qnp9OSHIbdBeBLnq6guWPzNYBMVIkBaSpeQ2N+2usVJQ90hpruyqXlcqfas+5YAOYVwaDW
hgfGdPkYH+l2T5e07AlVOHEvXmpHLgDi0vwsnWKSdbp4uLwecWUrYM3PyHR3t4IQkBA71qNF19w4
E+C+5CP4Q/l3vCCCt8juX8uhygxEUkLlPNy4Wp22Ivgp8BvyHE9IclksSMyuVra01878pV8UIIxp
Djh8Fj+uO9S+J0SCBQ2u1k39EJ6FzN0cTreHllVePRMPf4I6cuu1B2eNC0krjbO8TPU1306NFTdw
qDwxy8b9wbWRwzo5IaCVbMbXz1NMXAkk9frHsFADm5XhEQ4r8pk9dJJX2nlZ0DQUD/IqUtTlNc/j
VxXsbkpbegdrfgljgXSqKBXe92o8kRoKNxgavVheaQdmwhAlzSLkInCXdVgaYDEpwj7/xtYuw8m8
AUeABYzTv5WJNw3BaR7UxL8q6HWqsu0MxJIiLAhESNhRM9W3bjvwCM3hYjG3wvfgpVwMHmfzYxY8
80SieFy/pijt89RTR/TaQK61wx2Tm8ZwzNoUDS27ig7WgatrMX7eLvY7N16gmtTG9E2aI+lDRytf
kjAbkzmFrny/WSHCielmbsYQuk8BCRSEQBjMj42I6a3k798N6RiNU3KxaAVR0BkQS76kCEk8N0GN
tdXVBth6pg6CztAKa0z1TT3AxEPFsrv+vYCS5DLOlLZCDe5ZF9RH4lE9b3ThqlHIcQFTxQ9ZUd/V
EdR/Kndx+8zJFHu/cIGX0ILNNjl+pzxQgrk7GsHHnmOS9mHOzN6KR1eCgA3qx5cYxABTisTGpWj1
NTkFA3nezZ78PhCBPGcrKUMjd6XXbszeXFlGKysfCudk2rKuFEWOtLcZHniKtu1MfZG1ThTMgiok
S7lWk73bOyPmefoiEaMIrbhmdil5zsw+zfAniqV4hVYrpfct9r3APfPlN9D433Rwh9BaMz/vfEIM
Rv5+ZAT1Jqg+RHHbvwjBLcuFMrMneUUFx8qMcCTGBeXBOod4vw59JdPKEWuGt1gH+D1g3R7Vyn+K
Q3R9lDBEuaboq7Jz7rJ8vahkNXPZH27o8vHDPB3+P0ylnbJ42cZPBedgWhMs8LjlyHD0Vl3fnMJV
rvES9ztoVZrNtWGq5qUwQrP5dRYp4HLLaW6uRMoL7bXPUszvpzYR02h/u64BV/E6yXWTPl3J+iy7
upmWL4y2IHvO96mJJVNX4JWxGccr97ewddEq66g6wUWKrqYfYntTQ2g+66wpXYFrK4TEJaMWVDCd
GzbTqv4VkO1c8uj07XZ0iw5TZnwkrm67h/MJDGVmdQFaayM1lCEpiRYTIKdE1DKdWuwKL4kj3qbd
MIdNbgL7zV1LEnjht9l5LiWMBOLeDIcVHGlDM2baUWd2ua5//8ukgWx9hyNutJNPOb5PofbLr7Yy
EHuAY9pKxpmYdCKztv45yHcrww3Bo8F14udJw0QNDpxd3PcdHxCGOWUlQ3xyNNy1NB16+X3+QJFS
Yc75KK1GsB8sNtT0uccwPoT3mPPdL6JZDlxWuu+TJwrzUlpVRGxOHFiW5cSVsrJ5X+xU4zgxZh2F
r1BdOmj/Ok2/Rr4lvbqEK0eRvWYvyanyed8ghVh2jl/C4Q8EiJPadoOSBQlhuYD10IwvyexT82HQ
Z4wrc9SWJUimW5HP1nEfWAGHuaHRazwXAI2dNoVLNSLQNcmCVKOPxskVUpgjRBwaLfhjNPG02DhK
OQeiOIsO2LUXzjOsUiTkqIY0OUy6pmQ29c0+sHaDRtbEhN0VtuHinyEy9eoztR17RTSnkZWHCkPK
OVqmJtH1W8VSFjqNrv+x+2J5QH1A2nN4JjIQEC5tJZ7jBvHXEkFRGjQ0lciBhYuljvlYInERHpvv
gm235alBlM8dqECIhM+FwlTenvuipzwX8B03wc86GaFKd42AaZsILeXWAdaCK0Tdg8BLGASKeLy/
qSRH80Qpr9vlyr+ncg0IgjbvuYaowgPlpn/BqxezS6YUhdCzIXAC87Em+ijDmghTld0DCO2bWxii
hx4UIgwWHIREx8vuwiPSrs1hdnBVn7bC2gv0uV2FW0WxrcRNsoQO/g19VTzxTm0mQpvPZXF8h+Iv
XVievgChiacDhmec+rSYvejQIgLjKEBGgnGaxGw0qbn40hTP0Fffx6TcVD8AujNuXrmLAa8/yA0F
TF8Z+i346SyUmehTWkE2LKDRvSkFIDrWkbV/H+l5Ll4cP2cQPfwqW4arvdHQBhTK/d1FKH42VVJR
WfxgbYJzKY2yZCzboPXxKqcRBn0o8iaGElgdGSvmoe9iJHZhb89/2Lc+qzvhf6nFtUnemVm9hUrX
BpN9vRWWnR+U5dSacMW1xNFxwf8Jsuee2DWUtXI0Rcsv/Xs7xW97RgOU8YPvSLkN5Ul7fBYfNrtS
QpVxUmMy0waPH2zx5lBBSSdYuYmWuxZL8ftvLRKmmDrftwjz8ixgj4rQOUdUAUE0wAHL7jOkFTfc
ufJWvxE+Di2YBvN1Zz4BhJADvpw5efi2bbTbBD2Ah/kT7huWGlE960OPr8vDtoSWi/2lppLbD3+X
pfEDizPYHWueM/8aXyWWODYN/0WBKm3ksGek3nWiRGaKEes7mwsDBpI2S3ah0hfQVRV4sZ6FNhAa
mwxRNuhDb7pALdQY4HfpSLFtk+L4N92laoOx6XFwEld8AFmZX570ZWGIu3TtT02Xfc+q6fKa0evl
o3BGcLvf6LNIG9tVQUrM/cMYDGt0tS1c3374xrYF3u0Zxwh/E+ZW5XkLjYvj22D2HbGp4yELuePf
tjS/R8DJzHBzrY36cwC0Zyq+WwENxTHg/4+Y2dWSYT4rXWXFUyIKLZKKfVs3ZYChIeiCTFdF9McY
0dJ8WP7tQ2wz4DqBz+Z2mvAYTNJMkjxKqruHcUbfooFI3R3JiL+yKVF/f8R61glNrOn3etI4APO1
RhU0688BfKSoyhWUkWK5atyYBzY7AZaEg6JeQweJZVI2fO9gpD/1fMZ9AgC5BnsI5y5iQdYpyfbW
agQ2WEuTi8n9pjvwYu6RCRHLY5LtuW8JA9OymqNit49K1FvTfaR9wlP18fXln7E6hRHPd8ExvF86
hQJtgrX+WU8LEsHna2E3HXAqAcUNDi1SYHHFcP3R2dRhxBOBHx+XsKlKRaTd+x8Qh+a3Uf4BGteI
5QnISzZEXsldPJ0HUr9gkm8fYtbdF5Xl9n8hDrkb2iW9s07j1sFNhOy5M+gHe5SCrL/4HpwJqreM
3w+cJK8utpBFhjcXpb7tHsGD7QHcMuQNtCZoYa1a9ZY818ufdibdvcIRe9Kqkwd6oky8AjLdqXZJ
9oQdzFM8cXvM/uUOxLhNvYoTZxh0KxtVcjbJeEjVLOjCAX3PgZQ+Zaah5qF5q5+fl8UcemF+OgOQ
i6U5alocQlRwXMtb1d2uCXUtdb48ZkC/QbA+hOlRSNnFE/0W+JWFrI2800x3vV3XgUoNhjT6oVoa
VnOqRwpVNZxh2syg27WetU7sa4wqnFkncbVnyo4Ch5rsLHNoDjyJeSplxHf2gfgbh96iBn3OhG3B
r8IIzn1i+n8dVt8y1VdgHya3EudTbEIlcQnGz7doEOwdqLGU2ui7e64f6X0o3US4hyCG205Pom4c
S77THPldG/dR2MZdTjnDpDkrNMyh0Stz9fHzGGNSDc30toEu0SoK1BSTevn/4V8/D26xvVajfK8m
JR2yGN2rUIbsXAsQJVCmE4imFXtNJ7LAGIhEwyRY9kFRAHIRoA+zZxBDENEoahJ6Q1V0ACdYfkis
9azuk38nSPRbSkJk2jzheMjmyIXUv/OgZXQghk+SgrcUs96K1BTrqqNvH8Rf8qJXN43GdFVarXC7
PDgVX32iVDrkJcDTfCiLk7X9y9ps63Vdd0+gCJKvt/LP3h/b76tANpMY+5W2O9waotrpxikfzkHk
CvtpD6NXNh8Mjjerh1udVmpPv+nYsmMu4UcgvS1zQ3ZRomRNPONAmkLJcr4j70+VNH65FakeLM3U
v+CSBJtOzo2xP2/MaDzHP+n1PqFiwFdBJYnj8IKQzRy0TCPES8hL5BGczU8Lz/kHYvA4wzrF/Ux3
S1fng90SSb/W9J3EbipiXgswm7PR3B/een97lgGM6tp7NIM0azA1yfFU7yp79heVDo789EY+JOl4
LX5pdsdOCxSESWfRJ9PzGR8TYDMqZCmeSy61kbEFzh1XkuIp3YHEsIzubzogweBvBuqFEu/hucH+
gb4QH6PkjNt3/eQl0Jd5PtMtYKRzeor/0U0G4zzVc2xpJdAytzveayzpd/AvNIcxzDnUevRJGtok
4RBjf693EeM9Qpsr2Oxa/S1YpuwSqRIY53TnnEg8iMFdkFypA1mmJN0VsY6TnVW3Ia4H9jIS5C8V
2VzepExQu+I8EQqRXW2FTW+9cX7GKeQOe8/z/YF0n0Kp8bzfJTsBO0rlcdiHTbOx3BYFQdeSTPQv
EnUE5uEw+JSTUx3MdHZ6ESuIWb1J6uUM03XGc2UBcdGt/h94iBubvhzHj4OeXf/cE8/KYCBhnlFo
mlYnZragsFXPd9vVWIVhQNlxZZsTZLX332UYz6SeBcgyBQGV7RtAbDutBANEv9BDY2s0tnkj6v9S
BeTJL9XaD6FzG+qoS0sfddvlGIaZaDGQtnIfR5byJMmZ39lo/sp/oXT+SExKY/LS2cOzIZuvYb7v
lEClCgYLk72rMc+KtlMsL3908rJphsjcWliY0O4y3fHxn1e8+wdkq1akqOOydb4pHdapRWkjRdyt
gx9vN0kBC8hvrFZ/Ou+aYqba3rq1lsz7/YyXXH0msOWxdyXzKdUJAwbQo8/KP9ChaBhSQ5GJmbmQ
bKH8QbCtIE3RBVjyCQKIdTSesQdm13+xIcQ70w0SXD15/QEwqPeRZXBttTPVwzO7IwOjyqYf6LKv
xcnBIEqvEJELk9Opi14nrfgvua8Lnn3OIynPQy8GVEmmDvI9u88GUI6/gjiKm4myOh8l/is622Xz
rj51HyCWKKB/LP2fVSk9hqe+vsL90t12e610qqZ5ApX0H7JChVNAGzrBofSOy8Vh668+73kFoDyj
vx3DjwiJfCDnDbvgq/AgKowLiYlREJ4YicGBNgof/62I+lnLIjB8J7cHXYaiYYkA8K+RQcpcm552
kWKrw7TlZCClHkUGROS5VK0m+7Cm0AK5SifdCH6vqK58bDjumquBO+fsJWlmnj5QPrq/tQ/IHpCf
WQbkmVEdMg4ozBwVlNI61KuZ22XSLIprvN/RBtVmo8crzyKaPNjIuk90PKLPYOIUmqIx6FjlJS5z
8Q0khPfO2z/IJTvWawUmp/aoDYVhMAVb2qXXb/f6Kk516E07CSGNlfBNB/dVdX6I9mspgK9fHS+J
LmPcxggm7CByDz1kFTpQolnHLxktm1jk485kFCZnX6s4d5dhJ9SeeS1mhAM3fZlD1ld0tBtnhcDw
3YbzcxWY9iDRUtYaTkTkPqFWfVPiuvBWV0RRyUrFREB50dRcjwkGd1396GqFuJwe3dSjE53k82Vl
yuUxdw5KymwrqKdT3wLSAIKC0kvJtuMslvNyNZeO/SWVXYyaBDtJgWk0PMqBSV5ScxlRlclAJqrN
69b+LMFCQTrCwXic3ghfnLLD8V5dhzpvEPQ6q2qDRpT4mAk9n49VTMhCmXyBOomhvk8Ssb+VbcBS
CsHQJYJN14XIx6fgawylv0Jxzo0L7gtDzTLeOwzUSdnpcGPbv1egEc5PRhwLDI3jSyFuKhpPzQm+
VwSqAsztuXo8/YWSK9JpwKLuF7Pcd23Bo+wA5ldUO1bC3+/B8LvlgPObc+8HVKrhlMepUTr2VkmL
DzVgd2iqTPFoPj54HQPH1zT4Rs++hOfg3UVSFgCGL/gMw2XrNqfacbFH4KKiYBPngRe3wZzUejlS
2iC82t5aMOrf5jg9tm4dlKxhnsCe4k2Xifs/0aeo726Sds+6lXOimsbBFUwr+jQMzh1+zB4a/CNZ
2kYph6YW83VYRZ4P9cZGOgpy/yb5G48sTWApmPWi05jgwOVlfAdl4y05lt1qVjU7orYxr+1HzoOo
BkZmmktPkYngwIUZYoRYDkcYsybgx/wZC1R8cWZBA8kIVmcy4pnV4A1xHhZRAGmi7YsugVGCpi8m
E3qU5yK4eVxba8L212h5P+gG6h4e4j6FclM9P4aIB6aQDRwm1pyySx5HOKgMcUF74TEIu5Ui/8z0
JIvP+HdO+WQalFc9fOrsdMw7UXMQplI6vS4XTm/QPgifJs4JFOchMBhJVtF0UoQU+dWpWccqiPqS
mpnEEcLYYWngkodCmZzClbEyKeRIW/dz1Bp/aaftkF25XA+TwGpU6JenD7KgjIez7r4YSrNJ3jZ6
qWAj19GQ7G3QtV+wIJK49S6fsWlcrLiRDHhNLk+lyo7d9+D7eSebWdFOSD0ABqSQstXGQgd/ohQQ
snje5wrsmLcVZ0LP9+Fj4YenA0kyAeCNaxMjm2zHv53ZIu4A/0hj1/k4iOIB3mGLuO2SjjbiFxAA
IK57ktKe6C3VmqPthrGd53t4S3tvhMXqWxRPU+aIBSfhVqr5TwTwMwxh4YAHd9jEp/XkYQ5mKd08
UPcYr7RrfHHqy49vbPiwXN+hOuZasUPkNWBwTyLWlOhIb6Gz+7oEZqOflCVtuIgY9xuxTyuJiBmR
lJva1YpeKmAelH+GRqVHBR6R41LjIIyfIF5EDxvA54DT79c83gJbavPl7pk0gsnoJAELxrUsP1L/
3mYl3HhVvC3c7yNC4lh6JusMoc1VHqE6NDIZsjPR0DgExQC5izULrBv7ABqXk3ziGskMB9J8WqGU
bI4tNEok37T0QI2W4+g/ZNavbh8gzk2pLyTM3kdKtIXtZN1hMXSBEVZ4Z3KSViRC5ahMdjJLp8Hy
hYBANb/Rp0TKozTQiGUrTRz4bP8aXYti4c+6lMAK2HgH8QOToFzpO+XcG8B/tRkuKWRmn/RZlN+Z
qyO8oEQEzEFwhzzGXUOoLL1SyRpaPgusvOQdwX7wPlmj4u6gJsCc0yCut23yUQHcpHPGL0NDiKAR
g+8J4104gMwrX/02Fbf0a2fvll7Hzm7/EXqSeMpsTH9IfPqP3fIqlY0KBIhO4gWDIbWQSdeN1FTx
qAMRuPmJ1DMFfYCdEIjvN6ZckKVb1Fss2PiXlG6sBzKBx80RHRThq5TXe3KceDT91WNSImbCsKJ5
DLcaq+XZNbxukXnhNaJlwPpCf+SFzoB84bBghanE0D4lodzMvFBC5UpnH4Z4SdVln0fQ/IeOhX0r
URgDoyjEyT14IDlfwztvNJ+Rwc16hgtOf1dSvIny/uoNl/JprM1AVHdqFvg3aZhT+frSJB8KrjH4
veANIJHhcrimw9zrMcot5+TcZ0fibSz268b1ThYkEQdrChhGuoJK4ZXB4qsR4JLT1WXCwFbo279g
naW6+e4uloLK26L2b5A8Z58OIf866784S3Ywya+8BeDeKQiGpKpOkm2gofFGwILeq4ftadxlz39L
Pe0+RFN0I/5GEtpAwyvT1kRfo31HkPCHvUe38nw1l+0ri/qwGMk5G1liLMZu/yj4b9f/Pj/CiuWu
7MgVbAak3CN7qIXrXy+jaEssmgfXk/+7/7vQJ5aS0ZwewZm1rDYEe0ybAP9dkh/U8ktKvr9aQpD+
2FvF6aODNKQK8GowVjh9wMGfCO4zOcz8EKOyCwmoNFR8kBaOhDg0sd43eEiqJNCtCfHgwpFAR0Aq
/SyAYsDQpxd2mYPtiuVFyik8vdiaUBY1lsXuOSCbYuCe8tUXDUGAACr6/OlhDmuga7WdV1GmFQUS
NRKhZw7IqgDFFQZ9X1Diio9ZA5i6BD8Bvh5FI/MHMnE51CtBowUI79zSP8Sa0f7PD4RajzJsTrgX
NZZbZImdGsF24a0gw/fchHHRMA/kn/4rHv6wLPfkYVAqUpH8virivWVED2/fVpzJ0vggEpLnidLW
xb4pkqBtc3zozM66hRX0pvcdgoAw3m0e2g5Ao0sXXBYxXmvdAPuv99hmoS/102MEonOao2h9XX1v
fHY31JAyIkMQh/0/W7KhMdE0H818oyis0WHbPVCdOCbr9tGFi9SIoDeTQI4mGcThJU9XSrs8zWXB
57+TAhH0olUla5jTEOQMNgxCib7lI6YhNtgR4fQZAggoLsmiEHWhpBy2FXDdj0VRC6Fn+VmYsMyZ
hKrwp7EpN9AO9krqQA7Kcx3opoGj4GwrX/YFb+MrRQb4yhMG9iE/2b+0blk6b5Amp8nC3DGQVOg1
L68fXPiPtF2auPHcJNv6uoH3br2Skq6aUg0V0IrDY0SrM33+9KfMklEf0xWbv8iZirKEZulziwfK
ciqPk9AM8iM9hN06EBIQSPDJYy2yqyjTu/HT5VU7EvXNV9RTP7pG3YHCd4vmAcNM23Gn4ZgFfp6n
S+nsBRDXJTqzlk/X5L1O5aNu2qoeYmt3Co1cXFsF8M8+Yb+lRvDur8aM12gqT4ha0xWFZsLDQyQh
jkJtHaXhZrN+02dgYHmh6XPYPhWcsQvsq4iDrhlzDgmI5ZPTcXcafduRZkzUglzEBfz5ETLzrPva
rVNMsPrBcFZ7f3XMeDi5QovczW9kZ2HuT+V0ASuwjnLNga9Wlz57GYXaE4XIb2GaNA/9OaI302zi
9/5/wciqghtXMlTUXmiZ9Hm/PFiUzXVaW0xlMNqRvEr+QYrm1rlBDc5HXbE/ncOyjt9ETiQj7no5
ThLBKqBH88oxYud1aHLhCeghW5ZGCHGzmgLqMu0nRGcniqyIv6IU1UrgE2H2m/eb094M6O2s0tzI
yIrX5slDbVsP7VAoie0/WzGCfYAhxb7cyrv4u/yGbVwXaotUk0o0tt0bMAIWFfSYsK0GENS4gx3y
ApQZU3mHPTiUx7ldN39vYqWGj63TAvYwJNmK/Xn8qHaya+I+WTjNt9kCf0pfmQETJazSJWdpGgsu
wnrKIZsCdxOXzQ4rxBD+bE1QTU91/ojuiVPF/O1ubmONlZC+THOgsYqTOKow9pKRrAl6/Wos/1r+
96WIElFMAYNzNtqClnEZk1hroVpCXfni7u2umYUnRXujBN1wmUJNU2wmBnK+mWzGyHBi5QCMMN0z
+pp+BbSi8LRBSbMtzmsx9vqh0uHOa/+xrc1dkvz2p7n/zSdqxsreITWwBVtyBTJqtfuU27V55YhW
WY9ail/FU37OC+JiiWUeUPP+dujH1tc1a86GG5SbrVDZXqGzryD5B6Na2PQMGAdxjSmVd/iWeBp6
LuXjWADPI2rcPC5+zVyoCzPbS9oxSWMPbEq9klHPXb1iImO5uXYrEdkLePYVl2CI2x9QGCnNFDrZ
mB+CAN4U6tBtKJsxuPmQEufzHSVmRUM8iL5TJBgcwGezqYZwRcZb6AVJ5X9IATDmTyPoNdM5nuU3
pESAkQCCUuJKZBCtTlj/A34YKAwbnSh/oXho7G67loX7w3TaJnemR0NBIVWErF3a3j3leqUF4MVh
2kT21IXZW9JcTr31i5gZ5pdal6+tJF/qVee6w+Biwlo53lWJSOlwPU2eJXIO6Qen3oJxeaQGqevb
/D66/yPgyuDbsMijU2wLCt2WhkfzplhDBJFii/wzhiKZb+s+L8RQH8xF9apw/Xle+EerkA7QPH1C
P9UVzIn8xN90eYQFszBNQdU/ssFadjxZQEtJCXhECNBriOdhabyDNxJz35P4xEIsD3ZHgExwC9lk
L7chWur99ZMvpKF9aToHoSFPJ0UActqH9OUhXAloxJm4ZhpuempcFKsaTc7tfeKxByRGX4IQ8I3T
hK5+OSsD5l+DMOLyn/hGME7o4RWrhPGPtWgc9mOpofk0pX6qErHniDKvp/nJFJXpNps3m4ZjnSrj
Ai2Pp0S95PXNaluWgEuHvNjPzl9MWCUCriBaryTRT5wtnpPlGS0bqtvhRfAEjoPqcZ8/0uf3rmJz
CsvgnKz3qbaRGa4sKLi8fvNxkr5b6uStUNu52OPvIp7JOXc3q4Jt/+6WpQfxWU3MDj3Q9kx/1Lcq
bly4abZRSkK3/P/huM3PvBKSyVgd2IpxSblAFbaPPyeCe/rg/gpsL7L53AoyFpjWQe7dh3/5cjyI
cXgv1F9juGETO4KX6BYGYKeQmlkVKQ22LiltypLSFZcC9mzThQtBS1bAJ3dDWuRu2xUSZnuPr4c8
8jNTGBOKOMIgBrzAKyh3hGhL3czn3d67Fq9U0Z1iBOfn88qTajSoCOzyg10OHd5erzNXCMXqFtvc
K984XlP6TRoDc4RtrmcNEBCmME+sWBYdNLrVbHAHtMf5Pcaq9o2vAjG2zi3BlmPsoIrIp3C5VDqa
fM2FQ2z5EcO9B1r86rmIyLt9VeG3nXLkE2PTZgBpVPjl1U+1J251QksTgp6rn5gc3hyTFdRPgtZT
w2GUQmg22QdIZYseJok+g/LPZ6wGF93FQu9PS3kMtpuwM59kTa+jUvz86EJUaTaBNotZ8RsRkaix
0th+WWfxHE4zzVMF3Ru65JdhQyXamMrdUVYLoL/zukUI6ym7Vypo6IpjPUQiDCMg8bUT3sJvzMW+
EbOjp3HVKlE/p6CGRD9fqmmcP9hev1Ipd5legOoF/HM+SAEoFm+q24Um7omhsubmgZDs0rrNXbeO
zQzsYT4cGPCBhsrvOc91huV2mlTN7HH0D+wK3FZNDb2KqryIUzlZPYRwffxW8Pu8NN1+GFVqkn1M
5gHuxZPHsCcb2Tdgw060AbCp9sbxhHXUt8UvJjvbYJc5STCor6OPj0bqyKIJYiL8JPwNp8oh6n+G
i7sLR03c+wiWlf2dazWPJjIu+rxAGtEW+SUXMmqPW9HuU23sW8v33udy86hQh8juyb5gGDMrVCbv
zBvR1cfL0Dxrw0q9Lm8gJieOk1aKwwHwAD9W7up6na02CryqgACwSyPQyG9NYpRbXz+TKWSxUFzs
WAa45WDFDrHMxW4fSqoxks81Gb6QGPA4OwtIR3vdKLil9Fb1rB449PrYRietwkg5SAwt6TN4QoAn
JSNhDlYs0GC6ytJPlg0qUF1js7HR4lXARJSvbkmojkBkHTyyU62QYWoPunkw/acpxNapIW/kIyD9
bm5PfZ25nSTePA0Dpe+Oi33G0u/Eiz9Sax+ua49Lf19WFME7y5zkgazgKMQ7bapGcMlCfKobJTgP
7TciHWa86BuZ9kf5FF+XUg7h19oRCMcy1U3I9Rgv8L4cfVTvOKriRriM55bDJ48JfX7PJBicXyCW
FUiq5Qyh4EdkZvmb+HoVNlApUf9xawaaumvzWlHPDXdDLD9axBlwqGKCl4/b10Q9CiXN5kuwrbeg
QjqfBWGGoIX3u7TCDMquoxwtinPgKp32zjjt1jWwskfdT13baXS33EmBQhCRxQApk/BFNWwzgKlo
NTW0I/Sd67PrVQjSjJwWu/unkyM/J/kORmIPtEpMGE1oJ/X7uXPabM/ngEmP7Kyt6KtyadQnEdxY
5GI6upphoFsWDrDiB47hhV2vHh/iWvFxMkeGf7EVj9hZD7fAmUIoqgTOXq/pk1C7qUFe35mm6LCw
1edJpTYajA9X33kMHNU0b3sKg2V1viASlCGSw+9V7edwbUbVe8svoE15kSYwrxxYkC6k+8zmtbi7
62rcKKWBAqJocSbNV+2N2oN4CUvrVGJkdHZnn+E7qEoQtjqZZd5ILw3VGubShO1THlINLcoBxQIz
8nJc0ebo11wTCGKg4rzDho1MHnWvr9CRx4st7+k5Ot8G3F6OpxgeTnJQltEi7OdldtpUT8nF9EcJ
yq/9TMvKRqWTMsfu/OlU0uVGQK8XhFdvgAuZmC58gDPkhmmHkCKbNCUr2X9ffQNdI2ulG3KVdj2u
qEEwz7YqrDabLWieaORsmac/ppoZWaBisKiitCVApnCwe+hthCbaWic2D/iDXPS9QlGJm0T0VrgJ
24kov1Df5hfi8oNCvhoPZ/4o5xtlTj1NNhfkOS4NGPTGwgsSRgBTTcfOSMsTwnqWHQv23msyJD9r
vIlKtO8WSVSn+o8wXrIo8d6ULG+AFFvuvNaiv/7OhC2muSJwn5yjudDkGedDdl5JIH1+ZkmsYiVZ
gxW2ONBc1R63mfyt92C2WHmBq1IDXco0MdLK2P1SxZc2+mXpgwv9mjKVkgVpqjPg3TrB9FbyoRws
XSagIsTofbPLJRdKdg/ZQY62qgVM+BfC4C31HztI7nv8VfxKsAvd7FdJ/ktiOen3OmOzdJtdc6ZP
h652JD0QN2P0/VvBDvKaV8DjHEYUOjLM6VzrMKqt+YeWg261G5QuQ2nW0QeZ+aNAYgeWprmeiz/M
Rxq8NHnb5g+ixfcH9wjfS8HAwy7RSHkRu0MJDoybSVXPk3OfqNZRYCs4pRGu9K1YsVOIa2fD89BG
FPZKv55rLgWi5CAVhK+O6eUM1MSheazsj85Tcxm7KpMVptMsVe7rl1i4h+O7AiME31TXDGVXyf5T
7DJAG0bgSpOBfT2H1X3ov+RmM8lOCRI4UkkAS3vmkgLNR0wssbVehPCAo6M0CXe/2atWFlkHIwgM
S0iOaGPIz58HMGW8tdNLFQTTPPlrGzrNwYbJt183udDA7K8ni1/3f6R8zOjfqpyp+kycskH5nkD9
YymSpbswwsBaIF+MtzrxrMmlbeSx2g7R82JpOyqczwj4yxRC2NNYvK0YOGdv8W0YJ/PYXiQP1aSs
3G5snFdqDP3SGHcQvfRtggX3ziGgIkLobTyYdh6Rfyhm3S4ObxENW+XGf4qNp436Nr7WjpqpZ2YJ
dzdwIrasn0TyNuOQe1izs8EjsLIcRjoDhJEtmpkBO4hPDVAURaJV5dG6g6uZcrxDH9efwK0HBsnU
zPPTLqvjA4BWgqrhV9/23jZIGalK6MI86jjT088iQD+/qATry6PmF/CuF5t5TA40XpO9OnjdiMZ+
98UYHY+ejnK7Hitz+U8fJJ0BXZfKdGE/KO9rx8UWwK3ygrdnUiI8ncvT5z5pjkerEQwJhHgSbyDt
YuvI0hR5vZKSDMhRj9ZOT6QGknIVAC5RO3iY9kBmATlBDLYzCjL/1WuKfcE6m3DBqX7WZ76m73ph
3K4c/SumsISXKzSAi/FZC5S0LuNgswbh3PROAjFg41FU7xYmC7v2k/0xToHfPWZYvSMYf4I1ws9r
8KF6jktwRmz9PkcA4BQMqfqtLd7+f8t/PW+P/KGUnYaMOrfMQlHtD33gft0a2j71l0Qf1Tp48cyS
iITUS0sxAcRy6BYFRRn7UzqyPlDp+UDQ1b30M4Z3woY6gULiUETr4Fi4QMjR4ulREvZ2IfVgBxdL
9n/f2VcZmKkCMJMCNx+qBWpyjyHQUqIUbGo3lJMFwVN0xDekIaubWUZ37KPoEivOrXQTJXsVh3Uy
JkEGOHP4vg/jsZxkYVBtAdW2ikwVAhs83403weyXPz084WbVaQbz+XqMCPY9r+xmBhRWyZDBwIun
lJTjGHM2YP3vc6iY6+O3Dweu9hJGIqSKt/4j4/yoKlBAp1HX8bo+CmFEU1b440hazm2J8L8D56ID
yb2fd8E511MJRkaiIuLLcBfKVb80FcDKo+6nZ9EIQjVgK4VLQgItiSt8ag12xmJe2LN+YoQkPgcT
qxf8tDt2eDfz4ApmZki1/4z29W1FCILdcRXJFvBVkzqC9dK/i3s6k2miqYyW5Aw101tlMenVY9Gz
Eri5wpSDUGnzyasMU4MM4782muQ0QwKPDD2LI8r8Ukfz6I8PlokCBmCjyMqSVkLVQUiDytDKXc/b
+MeSd0HUVWxg0WISEoG6oN3XhccqhoSPdPwx7McmGlpDJ39i2pzt5q+kYhlf3f/gv/j6GpdwRjss
eY1gZkTwPBQ7PSaaQHBr7AGWPH+qQqIu12LMhpHde4XpRVk6JPw+B7QSruzARGn2hhQkH7kTB4G5
d3md/iEuovU/3VTmHVZMddq0bVngo8zr/0m0A/3dYGOxEH12iuUUnAlDXtr5kMcXGRdna4fgHHn4
TqY5Ru53EMve8LUGo6ss1jfUFFEe4rWsKE6Z8ibguPUfXiAaaNKcwMfo/nVp50D7G/ugR6/SOAuM
6RzgZuHqoaRjRSlvSxa9TBqNl1QrLwtJEr7VpXGYRWTvhsDK3tqLa4ILw4u3sboVF8iIzZwVscrc
zsgLYNG8ivJtAIpV6ONZ09w37QKRXbt/b9PNUKHPwAapW6e/2yXAxQe+T0NFScEPRrWs+XWIgoDV
ID9OOILnkyK7cvuS8E43ebBiF0lrTjuZaxC9d+r3PxnB8a7SUIUPe3nvhbClV7/jz36vKXu7Tzi1
cf+hS//9/UPzx23J+UWicaT4gUiEoznSAhLxbmxW2Eo4RCDB9gvBuxURNn3EWI5F42POfwn80f+f
WRHyqM7gZNI1yKUwO2jnzyLIy4yOKre0mODs5h3sR8m4Vnca7O+mFTnCxO5OO5qXmgMq4ry/R9KY
eFQLfLv492O0Mie5B0Xpj4Fjp0zY05uyYqcQoJUpQG0xO922sRUbaGUl3wwyvGLJv+FcogtP7dLr
dBzqjd0xVW9+9Nd2unNYwtIGvrMBM5+qMRFH4t/M3pyyW/8tJGEuCB/fEp8PVQprr/mS8SYlDiu6
mzR1mfIMudEB0rKAKhE3Fmc+bcmhEioxJFtHjI9f68stLKnmvaw4XdBC9vI95U+qeQsLuuhHJRSW
+nxvhoHvudG7cTdBbfpGIjOMTzdGBi2V27l5vELUHVsrOtRfxpyImZh6JCbCcMyfo8kvDRB5PdTq
xy9glA9FjOedtV8/D8B4XJNdaO6c6k2ftnbAK2dND8XseWC1SCTpPqgAD+SUP9xSORk1mBTVWwuS
hWqO4RRmorkRZo+/DnL9jh4H0PojrIBKDaWBVT6iYHeQnmvBazrwqxfs/UQODfXpZYwYOnv89NAC
3KUJISlV4XZdXB6KySghhfR7PIPc+leasrlcDEV4kMn68A8FkPrx5PONoAUWx/C/Vh7DBQkOoe4r
kjwDuwwWxZ1Do+dLAuEDx3U4hMCCgyVNjfT1So8qiIKyZml3XciXiQwmUgzWKVZYaBFl6GDpHzPI
rRCrrEQk7A0Dr5LRryVOiOvSqTr5FQX09JKmZ7W3r90NDMJZ7xf+tP0oM19FP0eFeUi7+4S7dOQD
2Svi72zvecwCG8Nc8v7qk9Lt+D2aP4Ky3kp8JEqF/5Hx/8RKfhYNGDHZCmFsKAjUxdkNN71Hhufe
NZmmOjCXbfAEJcK8tm0SWD64oMakqNkxEVCLQkA/pYo6rL7oj9O6pX59wy5hg7fExMV4614p7aop
zPjFrKIymJJv26q3f0WFIy5SKA/1vL7rw0CpFpeAn508B2mV4OElcsdVMzEEJujxSoJ/H1Rs9Jy9
Iixg6ilnSyISs1dUwsJoWjYeneAGqaJtM7cCFIKSmiZED9qYsX2XqSdHqg4Ah5vsyvfQ94gpZ7Sv
whpU61MgC2kuZDe8XGzInOHskEezsGaPDX0qjjKcBAPv6WdNvTCFZMcI4MGV3QjC6Ru56CA8zOwl
sb4KF3HIPsMG0zsxnSrLLFFQA7muFj32+0jLAW9yxQAXaoULtKeY1B9aarRVtkgy4ljNq2CoMlav
uZEl1sGa3iWC6nNPg3YqvvE8ZxuKK1netwa27ReffZ5nkVOEoM2WYsD47IOrNYgntYH5dJAhM59V
NLWjkV5Por6jds/510Samfk6niaTQP22m1ylLYXErLI+X2hu9BSBfmUTmYa/wOLtgBkp6Vzf+ffd
0bh5fVw5HB2OXgAt8m73J6euQkIng5CQm319Cw942QO8oRSBYjQEdiuO613ssq1sD3z/QqvLCqky
Vyu/fPCaPMudSxz/oM6FVaSCMuyO8Hi8/Zcs758PQqBqb3pe1vhsAA5j/sDpOwI5g9kIROe6DiOP
qDgoRJDzGKkNNxkfNcyXLEP5eUILcvQk2q7N4e9n4NLgsQhR8CIhEGmWj0d+Cif0gNRcYWenfdai
BqZryYuaSLIUL0wvCd0+7iYzlPvWAyn8hAWsgxYJNT6GIr2qBt8IXPDEfQ5VnrKYqFnvwr6EG5qB
bv1rFmDEDWpuKJryy0hU+li6UcWaSxcpUTdRZipVB3AnU0IrHm5qjM2Z77Wkr96u2Y49HAadX+Ql
q420/C8q0IGIma+AzAyyzkN7OSr1h0wLJ3kbkNK/reL5gl0JbR7z8DQVynXYrbKR5K498nmLMDhs
ydGrwls9unTKJTc9iAoUnf55R7FxsHOPlDkbTOo2xfpFVmcTVuSSnRKmtpg/4beUNSgUgKlzqnJA
PjR2oBEMPaCUZUPRYSCEGXFaRzfT/13O/lMUowAHmud4LBRZy4tRJSSoLQb0ol/mBJ6wnSMqeGAG
MN72LOEaVtmfkydDp4awkDFKj2fXI3yB1woetqNCVYq6fwMtKJDYQ0zvVAO68K8HxQqdn6w5OXN6
FF8SpDchq9KdjyHfMMrz/pR9Y0Q9/bqDAdyfB+YZyKIWTj1c9fYbsLJOd1cd/1Lyj0uGpAu2744Q
vOqiO/ZOrfWqfNu6jfUrHEtN6uODTU2PhUZc2Uxu4g61VbSwiA9kOsqi7ubXg3c1dcv2D5tPJj8H
HeLBMfil12BL8rDl4AVkeFX0Nohk5qMkDGLY8SesreThTm3U1XQqRRAQl0Q02Ppf96j2HSk/dDk2
AtKQ/L1NlvflKvsJpBYmJnEQ46P3DU/m1VZnIz41P6mKFWnkAnYsNHJ3BsPP3rDqJQdHvyEx7ny/
ERezLXOhmM3glGKLuxT6BVJmtlXw2A/pCjcboLS3AKGwp6p6VmTlKk6gMeMyXmSQeYM9+7jBhC6y
2wtbDSPO4L/dYXsZGIC4Ocd4vl5HzWDBCOIO5iPL1fWpqibNm63f1zH4+/p3nz8yrx26fKJ5yKtG
iJJhSci32J5BPoQ4+iK/ZwyP2ipHfyJcZAjgVtUkJF725ghfhB9OE0iwv3/iv2hjgaQNtrptD0zn
fLL3AKJYnfylMUSXx/lAXnrtoE/mY3eyV+eUA5G/YswvD3BIpW9z9STI87usIEjXn3SAl4mwkZTX
/g3eDkwEx3Ss4yWEkfFubjUTkQ9ZCF0mg1hCz+VU/4Z++444nTSN0P2FE2Al09R/wHM3vuCOw+Tf
qJkQ8Pj9uSglS2E4P4KkgIaxDj95tJHZAhbKFobQmudLWkL/rQqer6uBaubLIVW+ww8Dz2xuBxta
luyAXnxtdIJ9llA7kq7FnYtLBUq5AWNFBWKxPy0gC9c1HxkZ1yvbQ7yiiK+MnSzHtqUI77yyAL4z
V4NK6kB4yVZLDEJHR2sXP9X1DAaIA3XDBrJU+VWUnd4Owq8RVpwAc/DK26hUIhfHq1XvlFQxbXdJ
EgRGJ5Hxe9oShkphMH5psIbC+rV2PJ485QUrM8f5DLrBQVNokWKUUnZpNQ1cubjFQv8b/0to4MF+
hMgM+Fu8MGuYf01uLItNXgTk04BV45xLdFpf4W29znCoGcuANUkw0u/YrfSaN3xDGTDX+idsDYLT
E3QNw/7STHtcVu1J+v7iDcpoyJ+4NLf9gdOWVRmPBjCGW4UKEOm8Adm8OXO1pyQqUpqKw1MfonGN
bnNLTF+jogYiHpb9kAtreGdXSL4sAYPLOVqZC+wD8q/oIFmiCSu73KhfA3mTXqtXcqjgimxReLg/
wsm59fuTtc+/vrpRXyxGnt8/XBbKBrshCRyUcYWzwctE/THymlEPnNsTBolJ1GAa0ptjajf/spGa
EUaIzvOYAHWz2Wwe9mpIRZkQNEfhWVsvlEJSQPIccaS5Kh550395OTFTGxF4dXTkn29BQmhnqHM4
Jwp0qSs1S7hLiDfsfH9vqOyCvjmt71r3hWP6zSsfzi+CnxYK4e9XZ2F5eUopTy0CBNlCBlpEfE1Z
Y4m/qao86BxOfWh4NDsZiT9f6LNLDgo53cL6wxk2gE072nbadscdXWu/F3i6DVaJcPqIP+g6IuYw
xpemA5LUY5gSNOK+83daJDeiGoimkKdc1RgtmdvffIcoEl0jHib+BaChkr0va9EfAGRzilLLsTEy
EuzBUNhlVl/Tv/EdfZQUKEO6SGOtWs7B2DoXQm5gCwV07D4E6OXtxUfmYCoMpKmvxCCEkTHGuNrP
rhlTiEHj0GrK0UgTIhC6ekZGIYQ5fRcalh6UkEVT8wYSDAHn+lZspnS9tZm7eWmboxh0qX8cTPp/
peCgJYZXhV5SqEIUzc+ETDRFxvPlpjjrHG/fKwYHMAKvpAK45RWZ8Zwj6djdSc6qBGgs7HRkkvtQ
XR0kfcfeWgqAxrRrpfIS81T5Fs4CZFaovZWCDpDY3KHnv2ob2sgOAHRVzEop4wToJFk8DtayVR3j
DeVprFsfJ+7Omi8OLjUGuNDx0o9pvaQ62Vn7R34bJdzYDGbFL0oZo5bEmGyZyKMTPqsM0zLh0TrD
otCHIUwUvAgvOCP8cEeghcscL8m8EMV/ckoB64iM3SUzcQm45VpuCKv7ihrFtlwDUja1JGqJY/QA
ULLmOtW/aFMYxT7X4OvV46pIuF9xI5psaS7tVyTAt/XIVS1JUMF2z34chBJrWMKXILjxnYUAx5WT
Cw48yJHbI0qbFftiNDXpcjXg1e+BALZyswiuhWsHpm0b5AlNZySRZRG8rtTcdNL8df1Hj9XWRMws
c9wLTaUyewZazTUNJr3ej0NNbAZZrluswQ6TqZ6L8JhYNfwXTe2hgXioFKPgppWKV4otfImBSTWQ
9oMz/WUVFMBnZDyaLQj7blITnm+kaAJQtylF6Em+I+/hTqk68BibdqlcvC/WSGqQj7bBrsAYVzqk
uoWweWmWla+jpmd4dCpm7Kp8RAo2+23Kr3coq7OmTlTuGUD++UBvkhC3/7S+XvOwC+RoqLXlyqp9
pGexQdyrPTLRGmAXabgWNlb7VQtbJZ6hWrJUw6NSVl2e+Imc9+7k/8gk8fdNMAnpIxDNNHIcr6Fq
SNstFg2sf5FtXUO5VgazJh8UZQO/or6Ppdx5Yvc301o0yY9HfjmW2mBQeQbKfRlyl8HBgGgUjGFl
5IanP7eR0ftt7wXZd8ym187PUOGTs4rURTMH4JoumYRAuCR/HfXkMI0HNv4R4gfwq3EyX3qwdNgr
WFy3PqUYd64snBV8kraxpZ7eK5ZQPOEpT0SaeKAJ7/qVj8mwmyiq4ci/YEIQZWtfXbPU1w9x7gja
+wL+Xwtg7FvkgjGyLpnbs+6fqYagamFO/swhFZoEYkX9nibNocOWw/YmBTuxNGvDwdQHUXBHw3Px
rJZPAokkTqBT50uSsMvW/FaXCUYDqXRroAeNvnLZ57Bb0CvJLnWnuUhVD4/vVA+JdzQnAu5kGcHu
KF0MuRYbQoWSTYpQzk7755gr+syonSjxBTortFc1dPAqYDmQ5HxJM9Ou6VzXUdKKJZYtIIxqN0Qf
qPNFPvunV8RztKm3URYS8ic0MS4gPzslEM/s6VzGkQ6GabSnVUXRG3u5rhZ4UldOMkFxQ8X9NJM2
L8UyyA5s9iL9rnbhbHEyBh/0wZCzhj2JmCF6E0Q5T9iqzC/F7XA1I9j52tiHNZGAPOeJvoIVzFoh
MmK46PdRstFD8AHQFuM+hE3JzlqOgQoMH//VFTa7Op/mRehV/QkA658s0l7IhMwyEy4imFO1A6XI
yAGR81o8/VugSpLeZhC5m6nKSYwBfNE72qe18VuxBi9gr0POCtr0djiE41IKPn46mIYjYssmfJ92
idykLYSGnIaJCNJSFrIzuts9PQ3CqP+vpbiRWuJFR6xnmmCeJfawzwVPY43+FGQBu765D3fmWLcw
+fzrrPGK5HalVma6LB88pOw+93uMWzF7U755Z3/PS5FvKZpVWE1J8bR0CjxXTRGlIZYRaoVBm9bO
8UP5zxBTgKO6NBvigbUpd5CGYirFJr3hC1/qMJ8e1Fd79Okr+0BqkkWPceqmFrpV0Jf31GmxlSrU
POqt+NKvnIZ0eRFZs3t0vTjbpQpLL3ZunMuCSLEbmoba3/VDAW1i4WJR4GVYDoWQihuAIk7wC31a
/dNZ49vJHldS/FLvUJ+0nRgbnYlpyFJUGdHkMg8TkjbqHZlOeclDcZevrCYDpVtE/kpwml+6G9zT
pUvskPRCFFY5+mY2P03MdarQUwvn7XMKB/T89cHvkEDQ2SOQqfobu0fQwKaYjp6WZ4EtWSkOPGwk
n5cMv+qB/eZOnavI8qbwXjrDLRv+2GjtFWPqiCaGc+SmHl98kxiat4dl0Y4YDDEj3GMz+5GLMH3z
jGoYGLUO3Pzz81pG58u3xJ1junKYBQXliXgeo0slzgn74pFhzRNPXZl/JjwKkuKymMPt43/uzI8p
rN4pZXU5ApYlGjjo0ocsi0UzWQL5yy4Q0o43V/NDmGEcpWGPDGiBUMPT2r0SAZh7zbuyjb3kOi58
WkaFqYmH2nWMEwQM3DZUB2BRy86DTnHLbGZdFR7Jq+GWbnDv0+7S2J7LfOdoI+BMUnCvV44s1OKz
Nkn2u59k00bN5VLQAyi4l7G01d9VDx/ZssuS+xMvPtG1RQoGx6q0pFdHcSen7qGiqRL6r5Vp5KNA
8hmKqa8dPK8SqT1lYFMZYW2AvnAg9MiJyhg2FPk2se6ktWJNpcy1DKQLieItuip8iU1vzueC8gv+
UD6jQ+1wXmeAGKKAZ2Ex/ep2jjIyZtP4tq8efJJi9WI8XBwKlgDSwMNvG/aZJ3P8cYPx0NnSi4a2
0HAqAG2vst99yo1wap8cWFTNuJltonxHTyAhltiD2u2tvQGVbr4jMB9Urxs8DNDN7O4vgoJkNMuU
LjY7VLpfnJv34iV+3JLPXeESGLGps9CEKxST3gy52Cj5LPvi8TIRd4jlHNmqUZmWUaHAIjZQCjxw
uIZPU5sC1zDB/Q/5EP9HfQokjCQs9F0awRKc59AXrRwpRuvwxmvCKZjMb5e81a5JDa+0cb+J3xW5
W4H6EzlSCJEiBM1ggmd3g+uPgYFRQ3PpcWU6mbSMAN7K3AcPcZQzV5QyPBdD4Q4q2JcPgiYEzy39
zaK6Hemn73Y1xd6zIPxSLqtN476u+s5coB0Q3DRPPHmCbAcnTX53fvFOj2SLeFR+amBVoJ7FZZKF
G9274whRoG5q9DHtsOK4FAr7bwngwo1gmwd3Un58w0AOnKebmmuQVnyKuHciatpfO1tddO1m+UpL
Gb6WxicU0JZjLTVM2PTfr/gfwsl8waLwD6i4x/s+dfsHTrakH0jEx5DlS0txwVUUjzqUxhL6Xekm
SIsqzHLWPZEe4hGKpkwfswTEiixF/lxGPvGerW/sQq0U6/uIxOUV4VHYfFNPfkWd8LecrqvA9pef
dJq06fCjQrBig5d914NRKKvNLXci1q+Shef2td745aanD1RZV5gc3pUM7Y9AetvV6zD6IF52QKw9
war9nmuC+4l3QjTZi3oi5PdtgBWcqK4zEd5aYsQQ75GsJwoCeiWRw8up8r3HO7AfR378fg+c2n+w
vvFfvpdYdiIocoeg4Ml6s2wxNuxYp3UDkeTGI3INPSzVCPtcBxVASZWQ3HmFoaet5NSdxrGqXV7v
kr3ZloBY8PD0WcWmw9aPppsHFb2q0ook/ZzeKH5+cE4xpYfDdBlmCHuA3ArBavg0GYGSTT7IG2i0
OCR8CEnJIAAdGnZjLZgtLt2k8kSL1LYA8Zix+D/kNyM6ayVyV86xxFM2Np7ODvNhFD/chU7yvWUN
Vb0iQXz8BRhfHqqeHOQyxm/Z1i5LXe3ASln9T7WLOdPJ2LUuGl9EDnnccm6vGdvrcTGO+k6iQBrR
T2pWWbo+C1T4YClm2CCS7LcSpvjTOfYXP9N3MzX+ptUwQ4gyKzeVxrCP76rn8qCsRPK7L7Gjk8T3
v5MaoT0GzJzljiibwxsmjl3gwmh1NihBTPf4imSJNCyExb8bs/wFI4Uq2Uw7xn2Z8KywFGhjwFdM
BsD34wsT5bvksnnmAMfe9HH6PO9Xk6OWEc6rc+qf/qOtvWdsh6Nb/HzF/E29q0MsSbXdBxZUKosG
VVf093lv0XA625jKUkz3KVmr+uq9ybNDQZAZafazqmzFSJNBtlvuqoU3RBpmJArokmckbljK8LeO
EgQMazynbJ4ZdQXQbHazpeZ9wP5ZmxUSBJteL0XRhqoVLej+DN2j/ZBlVDJxau1upZ9ZqFePNaDH
aJaUH3JNiosGVxcwcoyG4EPgDQS9rYzvdw4FNC3K9ifKYpxLwlojwHnGsyKamXByAUgepfxc/tbN
DUVkubxYvMxlGJbh241TUpfwyYQ1JWgv+35OOzNjIOUYRRiCm5GcHXTuHzwIIC8ZOazLoU5Twhrs
mYo8Re2p35GId17xv6Gp6Xzx3TiT9PgziCVcKWrlYclO10NMMipUG3Y/fxY2d3M8z1qkgzh2kimL
AMvqORcdXgiBPcSwUcws94lPWfcgRKXWKEkwS5h4h4OEXWrNRRGqoLufRt6lUsskdwskRdKzEIh9
HYfWHHQCU/HFKyjMhCAwggWXNy26zanpCI2hd7AN4+4koY2dCyaG/q4sS1zJCv1X0jeNcUcvPB9Z
r4P3xfq2reQb4Ng3VWLCvNm+O2htJGXGwzGd9XPDC12Y1Yhle+bGXLcv6gy/8cvOPc0Tm09fF7y9
JNL1NmKykgsmu5IBU3vEh/DVgXJY5eMMO4ACqL3oK2wOPiBVWqr/aeD17mXcJyHCWzyzXk6XkYs+
ZMetEjx/ehlBbYf5juNDjZAVEf6Y1jCAPDLtRiv6uSBtNn3BnLo79l4Mt283PpqJDW8fdYU578wL
JKs+iBmgKlMXmUIisdh2XWdwRGH0B0oCbNNZJlt7s5ApdeKLlUregf2sNmof0jynpKaaJiqS3UUl
WTfxLbjvoyL6zfrVFSYKA2W4DrgWQu45fNfFQ0KLiwuo5eeINpp2ekqngCwD/xf/xUuTavJ7Jra9
fFYWCF6zz74wyV1UafvvlzPVTK8cK+fS189y1VBsLPqBpncQaRR6ldfXv9UZj4PcH/wX4FBx5fIp
6JjGRD4d+SUelZ9YVFuI5Sa5fD1LNH8eZPwk3BYIrNhGmyaade1Qbl3FCcxU8UO9q2EF4PRBkIQE
IDbkeKNnxUkXdrRLzsl3oyBJj6u+iAQfmFsHO5aymaNgdIeTWIUAyMVYUFk1nzLGtB1OTJydR6Kw
ixU0SJTBUDzvCx2bFzDFL+kiqJlctEqKAxxXTZ1UFcEajerMaEYrjnLxBQo4GCzfqkDBZR1eQQDp
BzjOsx9+BpL1XZqKW4GqTv2LZWQoFfWdpM7FuN7Z6fSEsUxhvVeWj7hfNSTZE0EvJJzKFuupvg9U
1V0nmw3trUdHzNO2wmqg8nAHSzRKbOGOWHOm3664/KVBew2XSuCyMq/aYmIj1DWBRcsSb3c1cJYI
QyKmxPTeRjdmnA9Xu02bX2sBl+ohOGts9wcQzCiEb0P/jzE0pnltl1fCRvXFmIEg2NKSaYNWpTJj
p6QHxfwIs01regO49Q5cM6eC+7xex82U8DhVw9PAPSwkKFL1s+kFUWq1xpEuJG2/eXQx0vLJzF4C
mpUX5cjFrh0Qr0F/RxU3NljiWKE/lvBMOo+3Xo888KhVrwJfWumkyMk5M6s9TQ5TKd2NP1zsA8nN
0TNqED/e8DdEH/XZiSnX0l8xy9jqfbnNs0mHMnPv1x9aY7eubDjYn6dsZ5C2Nuzqa10SA5FJqG82
3+llkVPnxoQTatBhBe8I0SdizhIx2AmJEkYaY8scArCDvn+Rm/8sCbOuLV6dQuYcTuR71T/pgZlP
/BIrptm/Co15YbfyA6lwGROQHYbT2+NUunpM5phQpvl5efdIvetosAJkT68tJeyHbqziDzYwtfl6
3rXN+wAjcHeJz2aG4FWrr1bjXD64iQgY0elhVw1EA5u1xWtab094OpZ/1EH56M5IxZeqJktlg+So
+DkD75S+N6HahYrGkQUEO2XIc2S9GMCWXDeqdXZuC7Kwajtbc6UUlHfiljZVXxUNIaBICQWT3Z3M
LDaXiYUv0QmgKIyJgRgH27Wg0qIGEUd8knyfSDXotlr45K2ZyJRbO7cLoQXiR9nCv7cMVTHnlY4g
off9YIgS1Qc6nceFd46pY59o4cITVv7L9qLShqfrqwlQYkD11AzQWaqe/Cco2jNTz8eeZTNMo+tU
6WF+3PZVnJb8piAZDSzo96cUw6yd5sb0GHI6mSNCqEQZnqXs/DcvSZCWC9itebuaRPTjooOQ+6/P
0t5NGsTW729xUPTeaQCMDJa+mr3m8R+AsRI7TC7ahB46cnIR/xQsGxZaZdyiVUmcNVD3nxclXJFB
mbAkETDDxyGqKqQfXQQkUsRBL8kYyrRtKeI+q1kJ3mSU8oQ3D9kayAQ4kM0P9TJdllzyiwZego+Q
e1ttedlZ4cEbjW1laIyq2/Xfxi6IyW0Mi2OtdYeoSi0rXcETJYWxbbT0vnd7FZwskJby/Vqfj0y4
RbShjtW/CvYLMbGzaQRRNhXxHyen6j8yuYSkzewh+3GOPk/qtzyiAXaGhBFk+tXg+ZzmsjD5wvgk
G/yIZUckVJQwPkWVU1obW2/cv2BhTGac6Vbgfm/Z8ZXaWJwo0fheOO7owHyl2AbfzT5WoHglljhK
lS39vF8Krgtn/Qeu4eEGVSXXOeR4a4TsaA8JIa711lGcY42ggBdSpmybXLOT/S9AcZti/9dUSlzF
Yilo2km6nkR2z7CW2NMd9EqaBDFqJNAZpqzvC2CSFOHNc6yy6iGDF6nNsYnByFFd1iWEZecFcTZG
Jd6oeSjNFdxbQniYmUwRPzMgdT6yMGD2XysrlO2C/3KHyhO/g4lTYvIe9uvryt9BEVvpxSRI3GOM
cBQexOi2kEiGP3DKuRVxgtadKpnpJlOWXtsJiQjUGaVIiENvfqw0CplUJ5Khauc9sClQ10Ftg/mW
TGHKwyt9cxX6bTqCZdsO4JONB+itf0/pi1YBp1Z3JvMOb7J7TSmP1zuBUAt46WtyTRcRxyiG4RrU
pIwIOOcXTy9A+6/llwoDl7BEJY/UEI5m+VyG5qdU9i2LZ5TyKz8JQONFYqbU7XfBylYuOGY/Fd71
NYLPdFq09jVH+QmzS8WQhbrTbl8SNF7Lol4RO2JMtGq7bwq66E26U4xF1zv3ihCzxRzLCiGlX/us
5aFI9RcUPso6zwa/zbkE4RqORDRpFqPLtcjI5t3YMWYSoLtBr57B98XQGFXMuOFY9h9XHKl7cvpY
H2dW/+GAHzVGNPaAihYoT8jzCYJWm2mAZRp5xvgodpQl0nhpRFDjCaFU+yde2eaXw/0G7xsUOIXs
mgTa2XQOj510BDjI3cTQp/CgCNsXwPm7lIcDXgxhYSI/GmkD7xLj0SkDlPkmMFvEb1n6eflrMftD
w5017KZpyZOZHEuebXdIav3m9iACRtp6d8QoghBZZ2y7pTEVpDb873SXnSVII02HqAw4sKobMSzJ
FRXKRcIPad/T1ANcLvwwJKZoMP+1R+uXdm8NFJszR0zYMyIPkr6cxfqf3c0deCdC20vVFZ/sk22A
rGbIeUOMR0suMdamdJDG5X6HjjNKNc9oHJVgEa45rsqZD6f1no8akpCxfrp64DLz/iIxVW9tIJXG
ZHu27EZJdgqDMYzqRo7V92/IUmp+n591jKZ9Fl9ThExpl+ZV+ha0osjNLosRjBVJVuLt/DDKyf9P
baIMEZAZsReUIfBCYxc4UmuOTno9seHjRPURhru3WigYWSXDvSAoeR1Mz3Hu10Tr9wvgKmJhKxBn
0XFEVQvVchuwqsW+PZGhaxRpoJYJaTqKLZpLqHSYcoCBQ7x+STz5+UJovt4Hyj4q5RYalMdUl4xH
GJKI887zelDaRdHwUHO6lYofMJ7XdZr6XytSlRCl1V7KcnBxPaqpFCawLu8nx6ScDu+ZsCTzDZA/
uTkJTx3IqVJ9k3ItaT1BPv82yDGkdrRJCnV8TCMiXn7FC7kVYNaBwnVnQ8ysZITKJg+qeIkcP4ap
D+hxwp2G6bozqoYntDX9jq+00l9rLd/hTEJBnrTxlo6FZAwGptqUAurrccATdLz6oeGMW8kRLL08
1eopD+HHUouI18fnOMwu7StWON+U7dpjj/5EUiJwe1nmuimPv4AEL4iHasObSmaJOqyoMXLqOAi9
w64lkcfLuL3SMA7w2EMORcdGEQVvstxt9/BqKSCcr4IzslPrn3wSQ5E0MFpZBLj7ARIZfm0iLDge
2wBdAcGFqbYjVPNLyfphZbUjr2rFy+LUMgjrSVQscsr28BpCnbx4Y3i7ISJPC3B4lnpVNDa7Xd0d
iwberCMjmbsar3cZhPTNm7T6r6qrwaqmR2yCuW4n/xF05V8E7AH8SJtxOaROL/TRkhODDY2fYrDv
8LwEAN1nYTIgSJlc8FPebqsrHy78krhSfAqUnjRUqapGTeypJ5QLNZI0lj8vjev+enSC/nZCQS4o
eQn2VN7KVwCHP/RqTJk5/qrSK5qCytH94PEUNGVoAq0PDBmt80uQHpGjW2CNFD7w0eAwaz1oIh+J
V7kg5osmlaTQP+XSPF3BE/e7E2DoQYHlW3EbRNZpDRTnOWhrdEKVjMn7pLVyqSQazlrVod+F5mhv
yh54qtQuPuX58AKOIOVQqq4ZUSidiwErDQnwfchJLAVpFKoa6a3LXSWtkXlmIdUXCNG4nxIHM4Fa
FX0JHwd60CwXTy/oC0Z4zANR1sPe8QwPnbiIB25QFw2Hn0iwiDVLnaePZWoCUs190JdesbuZWvhQ
+kbijMTSoTB1+c1SkRFI6VXgq3vDcvv0WJCAepLgGem+cOq6b2bA64aQqgt5tBkhl09u9fJdHYMF
gKpM5T8vhl3l6r7FTLsKsGa3Gs8CCHndiefmpY1b94VY0SAbigtlxhozqod5rPXMhYhD1DAZnJlx
nmloobtADQ/ka0YBMfADVswM/if6BcRkNet8t8lzw8DLwX3+UCdeTZQLSy9SSmpZcU2CAWo/Sh5b
okUj+jTdQxlgeQZOf34F5/VePOqvE9xiTV3HgAZ4hNRnA/7i07ueCKQ0jZhQSjwSsi2c3ghIFXEP
yHgh83LnTMPpOE1vCnsqvpE/ARATCjtU47mxF0LsD7049YayjkuQ8jbp1m3VecBUklBT6C3pHOud
xsI8YjPHHBlEI53A1zmJKo9u96lMa94kwK67rVyHdcyBaGGjZCSkJoTvc4NJiCiMELhsTxbxgAWQ
JsUq3f/weqVLTaeHa782mdIYyZe75W6ns6xMJQUdvYh5DgSC4SYO1A6AFhgVrgWHKE5qlXt2gaKx
6Xf1zYhTGjA2grbx0LVTcvMtq4+JPXgaTiYufAtOflP+l/5/UB64r9QgmHa9b84scsrEzNOUqkk0
ktMixoneN4rxEYR1iiaX+x/+VuvsMWMuNqeFieWzxHVyvfBl/maJ7pw5LxgwRfgmrO2SEid4pvBy
gA27gvHw3mhHkR9C1Ou8UGSnaH9e/Lu9YB/EDbv3f0YhkuSpZXyuCcX2i6D76Iwx0MXDrN1MeHrH
IGqm5WdKLO3aGeQ3OdikuRdiVLYsUkMDEnzc1TV2sca0l7ZukDzP3Vaw/IwYL/Jvgh2qGRYYfsBh
VpCLjZDUv9owzlhzmNKbKyJb3PSZ69VlB6MgBucxPqJy7P0plA1CpQx5vwLdFZP+qdTeSNltW5rc
YtP4ehfJxPEDbKCGIh0JeaunT/DSGKhRKGfqQydB5Hl7k6NYocERwan9+lzQAwch/zviYWJbW7aR
2uK8xrzykMNONUVZK01nsi32pokqShX3gKnvLclbixPCnAOe2dTFciP/uN1+AGrLjP7URrSae7Oj
srP0v0tuvE0LWt1ZzDCaNagMvPA7STHlIkNTz6xefFpgNyQ0Jt3iqeEMHGht9Ep9qvmmLUOef/q/
/3XYYrj2Xp1bE7FzT7Z04O3M1F3/3wB/9cWjy6mwR6Xj2AJb2RFelF+4PXS9XTrI5qGBmSTWuGsD
10y7z+tKWQeitbjMXGLzTtMF5/k+aUmAifGgjNGNKaw92zAxJ2c+gjTWHTOE8M+wEximdK2C4gMm
JRGGEFerRCb6YCSb/Rf6FnIBExK005nsof8p52/dM/UCzSxKKUB34uZBC58PzhGhmvc8clcDcstk
Wv7mDKXV15ezzqYIHBwQSkFirYpGVIq1o8mjU+eDbZLaxFigWsrMruu/jTLV9qA2EqKvbasMQ4e6
zy7DfFUbXcWsaujAj03npEYhWq5HyYWDzFyCvEeMCGVqW861xtlAW1QlADXoo45S2e4NSKPafopy
FxLnUOiEL+QPH6yDaDgNY+jHAot92pL+C8hGIYcOjm3rZeJVqe3F8sn+/Dl9ucq+WiYNkxfq3iO9
b7goXpkdfTkz2PsxJiB28EcoYMB/90qbAUlntidQiSqvpcAJMZ9fJ7mPz7kbAL5ph3DUXio1dpV/
gCztyDehvx/o72aIB2LVwytE/Osz9j7N/CWLdFcO2P8vBrcSlqRDPQnF8hYhfnhh/fLkKELeWpB0
dJqUObB8gTJkwzH1/4U+YVwsBGM8MKLqBLvThCIM1HIP07Dtcp3InvPo2k/ct0WJ8zZxe7mSlcZX
0URdh7zlwr9uKsEyUHwSU+wD2PnQvSrg9gezCp/KwbAwStx7cltNO7g8lpPY8biMOYtyhqYFHFYz
DuHeKiohl/UfFujuUeIEDeHQ3G5cnXqkdEL5Ym38vn+9TWKxiFc5lYu5HVNL4r0/k/aUZXBf07CA
ladDXIuCFs++Hx0ezxE12rwxXXN4s5RZ8FRBfeuc9VVb6p+Q8aAuKkwxJ9vLIIFwEF1pim+PKui+
cI5Kmokrt9birMQoFjWpr8W55zPrCs1o+k2wDgeK3gkLojLVYpf6v9eWJvVHTsCkZoenHQpEoDHt
uSPY3aTMcDGg3YLQKbkjQqbmMPFqS8a9lqI8GSYZ7lKpB1VbOURB+jpXUJ73VC3iXB6ZCopFSZ5O
L+pDjzQTwDQ7AzTI4820fviNL+I4dsF+7IGwKiXdJc+vNHPkv0m1KZHFLMRgO8GrW+OybHLvroIa
X7seP1AY0x+EzYz3UZeCE182L4MALhD7PQCkntuar2KX2DQY/mNanfdb483X1GPM6JJJdy35tqsX
nvZz0mD1P1yKGdozAYviD4+inXENHMxSTELHHxktOUac5+GC0ZQsSdAasgSlJTYt7HqS+57cciVy
GGXFbmj8hBi/Z1a9wdS0t+zPd6L5TtoaWdcRVzKyzhkTSxDW6FaN6zScTCTgNc9hlJ3gNGLTg5Tk
B5p9t6rTOYeBjsRZC2y+YE/JjcflNFZn59g3Xzke69GjWBm0ahalVmc1GeS2jcUQqYvfwWlitHad
UMFz7CJ81kQWG7eDaopgqcqZ/EWaK19uVppkeHpR2liYnSJzQBRZHbcuUYxyrS86QW8vHyFT9bU9
0OLRSZI9TmcqRUO5HhN+8BqQOslryDAHKFwF0AxtUZlngl4gD0mtABVHpJb9Bj61T2xKfGEDgUof
Am243nKDCikx+Lk9QriOUhcOYLW4LIPyn3TFa5zwGYDQqn4VFC/NlqU8ogizotqf23vkSc6EZLTq
IfoxT3xakE1t7IM8WQXi5LMEPbSDWPUoERoKezDGslf5A9nrN0qz4cS5g3yUdiP06dW9xJsE4h5o
JCZb+TCvsjyKD2lWSf27JKp7XAKVZgGEO+vhk+mSOCmPndrJSg9SK6uWREdnI/GnRr6KudW7esDm
YK0ynYdNILHqAg17v3VfoCmND7uc1IRhOJNLs91MqHjRtkihUsBJW2gciBdodKqBQ/eumt6R6fgK
d01dCKQZCgWydY20yvAKu+QJm0H3rCK61OgxW6MG2hmV28Un+F36WMpnXKFeyqrqNfsX9xZG45QW
HLOb33dok8kl1r++Qs7dapLBPHeb+lDe0aQ1RPdkdhf+wbGcO603WlmRUBpRW9cvFgR1SKJQ33AQ
GcobpIXtT5RrJ0Be1GIlk9ArkCW9BD1jkYUz3zOqzAvSNfKisCPfqTELzrjgGGAeoMhM+qI691r9
No/JD8AeEvruucS6QmPG42wbs20cYh5ti2UaLjYTOZLN68b53GdxVCe3t7Z/9kJxq7dRbIx/4fT/
IanRcgCy6Q012dSHgOZo1ghKwL6uFaZYhyr7vl5yZ1yuvcyG72ilCJ7O1jf3YuJennFH/c2rJ8xO
bsY6aBPE31tzkQ0A03Lj/K7PmJRoCvZDl8zWMnjGyXaMcrpgWsEArUp/LrnP24Js24vG6ze5oXOi
/ldB7RpmaXJuyKd2MpDrz1sYA9cm43LZ0E75cUfwsBJnSAYtCn0VvZ2i2pDhipTuyqzLG1ntpY0n
NgdGMnPdW7x8mkg5fQRjB0rZU7Uy/b0sZhRw0MbEEmEunUFVxvAY0RyjEoEoM0qBYbYXa/VS6ExN
ZT87Cryl2RXEvQmM7GtzleWAM7GzcGs40jpAP6WoQnCTKGV4JtHofSkj1HPlHPZfBjE+/DfaR+nD
F/L3d0xs8Y99yFch5EZ3P8PmE+YaK3hXxOk1NLS/kqi7tE5KkplRCLz5sRmTsYlQzFt4/ZPB1ARK
qTi9/x2BtoKEzQO7FTp6OXwlOlf2PybULNF25gwksQu0ZeyWjqVGf80uw/K1qx3qSw8lT1XZ8/cz
OQefprebru/Yqui/PsffUEgZ/nxA02JXCnk7dKZ8FFTyU3Ud+pmWbkDRHzokNV10rmIrvzpDGYfG
JVGpYa8WD7S30LvGZxnjWbd3xpaqG0C2Ub6BI//FCVrmAE0Cezi9UhXZAjeqrClqEZF+ogynzIZi
/acqY+SaiVPblECArxJqo6Q7pgUTjlZWTuRErlqP6nTzGQJRfmvKv4QRv5c4o2YsK2WL2MgmRZzI
vx7rRAdC8nKWNlsRy1bWduOUVpyi94A2jqNzTza5ioa0FyU/qorOdZoxtNVo53zcHKZITb3Gkclo
3L3M3Wgm89ILIPVHSxMJtZHhNnc0QSCEqLKiRb2iUJX3bqIksGFfzQKK0yZrU17iWPKQO5geRU/A
kzrVu16CwMwsbqrADUJUCXspmYa8DlSzwBvBunowS8cEs9F7Rb+lGsONQ2G9MHjRxOTe5ON/Trse
+Q9NnzBEpPw33jM7afNpemncpzpN37RcHQ8iVPlkAysHCPUoQ4XDrm1RwUnoSkH39pJdKGK7/Qi1
v6zASBAQQVJ4xdGsb37pRU8zm6rLSffNSweDZ6VQU2FAU0W4wmkxlw2uN5Z2QlusybiitasP82du
AkwTkAkkKaf4kxrXAjoTGWWbKHwNtnAqFqZ5Ts/dxBdqGMkWjfRQuYoWncOddFY5AGlGvEQ/8A7E
o8Pt17SYXyMK7sDzME+sQzPg79UoLEtyEtHlYK2FrIqnse+bBQg63XxZBao2Ktg2HtJQ+mzmHnUW
wz9OWJng+yNN0x+VeuSajeExNEq5px+HWR86qBAi14H/SN3ETBWlLjDofxfQhTu23jpUU1tUPIhf
lqe8NRI+Lq0N2Xxtqp4K4UcQYMm9ZNGXVnSLJZJ5mX4T/JLO1rZBgm+MBafH7n/mwUMYhsoddZBN
ytiMUHaVPZHE0NL4uFjIXFWwGsnGhTnTr9jiaVyEZ6op/MKt6kjG59A6k2e0QJ+w66sFPIFUvX8e
Yn7hZCiOSW+gD5kjzA/ArwJnTiMU1mlV4M4Zup9bkk6OyDME10BIXOh1gwW1l4IojLQekE4yikyq
GThBUjnTv0gmldVX4QWK8x+3/QQgpFAILX/qIPlogH0ijzIo71ZLAuQ1ZEDffVTlQLYX9M00HN7x
Y17tqhc+LXgO/2f9/kG9c75Rpb9Odq9QTHkDkieGua/ckBaw1ddR4HwUR6vG19666BJYVCfdH25g
m57XJcbQ0DrvhW/rDyKNmKycXSfZy0EmzKepHHQjriAuBcYVdD24Vd0dlyZgGQeNPOejNTRkoA7P
KEbQ8/RgNPbqLClY7xLn5kXlIZThgZ0nhPdb3lek2pSfWDT76+bSx5+m94bMQ0aZv1yroAhakJyH
nWNezbxVS0XZCyK0JTeyz9kvVOLkqIEGlRta3SMOwjmAJcC110pHJyWqnOG/OLSi7wz/NvThnWlF
EqaXL8O7VI9AZjpU4PY2jszmi9Www0N7IfFr66rumw6L/BxKiw1SY7ECd8ZeephjbK6zDf4SJr2n
2F67/qllsUaXGUzlbt5ycAIr6IKPzJf6JWesFlFeypGNMy4X7vMylpiss79p8DZsIgOkOl1i7unR
KWyblHJ6PlowN8PSDRydemXyc9P1Yvh9HrdXKOkAf5esh6oYG7jKt0gXyD/nAn4xRXyF27wFjbYW
oao4M0cZdMFxF4D38/8Uz6g0LtqRR7AKnEqyjvLLcGQDH0S0MhhJhB9BAyGODo03rvTJZ8DSwy1z
ds+t39hV8F3DHWV75LDh/j4wTG9LfA0shodjlqqkyWUueuWbrYyiB7cWgroISxR+KX5LHX16SUl/
sjSybmEWgzNnFDvW4raG32H7ftQTYtbYfrNuG7niz+eQ5PnxiXkY5WBzNteS4DeZ5T5dakeWUHxq
jufGfDmsQoK6cgQf0VASlh+UycrgliW4xGecSoew7vzRChb0X400beCcen+1reQzTre2qQPJ656o
0EWso6hQ7GaXrgBz9g85k6imLoTnduaaScQESIb1bndvBvkpoNDrixwHauFUJffPWZ4WV+wkdrrC
A34aSzDqtB0jEK5AQBP5ZIcFor6N606kKc9wSvQuK1H1tvJE4Ks0Kc9RGXoUJDIbIn2fhrRlMIwH
eSxCFrJSAzlTEWd7tBcQN1zLFhJj3buH9wIB5lUwvYatmGkj2FnSTnh1NH0K1zR6fcB+ttktj5Qn
mGh7Yx5f8cB3BR219/kaTPbwkMku+mZi44sSpkfPAPz5abEEVniz8FILTwmvEQMndJBx5dzEPh3A
P98MTaHbgPx4mzxPOLigFlI2XZ+FwgPOyniKkipgtolrR3ex7iqUXEqw2xP5tA2CdfmMCqmmBUST
EPlgN6PyZ0SkZpmWEuezjs1l4145OD9NPcWFIpoeo5TXlWqAC5YTpsYnwqP6cLnuQ5wj2JbLSud9
zmr0RsJygST0Nii80RmGEdiXSUOZnfS6N1siADIJjl3hyDYNQ4n332mkKKsLSLbd00SVPQPNhULi
FZrfPmTlozE95JGl3RZO+i1E3FBb9dYc10+h18P48uGEJC8AzQE93IJFw+pW9iDfqdRGf5Pvz+JY
RGHYkk0cwz4ViEBAuUL1bSEZQazRwtu0EEOyd8x84apVjCSmIkjM59Vz8bGS+j7rTCMjwCQ8Grsv
piqdp00uTZFlOwsJsi2pb2q0X0BoKp3JGD/8igU3CfbUEdVanQYj2vLfl2oM5V5MGlBU/u6tmU66
HAbCkj5ocWik/YUaOQIAcR6vsLx9IhQMeAftgLs+Ap6GlvzQo7CgCUD2D0SFOKJhxkex102yf7he
mfJp/PBdxjAGnUtL7Xo+aZm1iQmyAnFbl7aOyxpfqg2cNDBtOiC2gR8KONEzsvUflO8XYhSOva6J
cepDi9uTt7MjrE3B4On06GoSJ/xh1UTDWRmpOLz+BbeWaUMYhgNx4dg7jev/FHdlx1ppRLn26e2f
v+ujZJE4StdZ5uMxlNpP7B6GgHT6LNR2066kxwX+TrBL8L4iq65tMpPxYPDQ1Gw20nvfP9E9LTdD
iPqOwwqbsj+Wn8GTwUe/esHfBgLu4XOrQBWaHsiawee/itykL6vpWqh85tzRwxFby3ERGLIsIiWm
gK5xktRLP7VKsSN9se9xNq9m6oItrz3WnezvpJPdbSayHANk6co9S9LMB6aqf18iToY+Hy3tSBR5
vNz4Jhh5hgx4Rwlv9FGC4l5RJm4XBe0zEpQLuWURAy3EwdiCd3zV/PkjQwkj3mRx6Epx9IcvFkDo
FLwgyqfYZpxdwUvk7IaP5RKycLnQcT4yGRIceut2dw83foBMY2tsUgZ79vC4bXdnbQ8RH5Oxealz
KoBHVmyEWizbI6++Xu15dQGELGaJCdXW/Jnwjztuj56D1m8I2qAlfcBHizrYJ45yjzIGVpSPWLCm
qWClnBcoEoQ3UwR5AOCPbJQOYXbQcsoEbJa+emQ/E8DJFw0dWRQJB9FV957sG+75D0cExSF7Tezs
10gHlE9rCb1I2ZEM+K3FnuPTlafoabGk2vxhKDZIvqvchrcFhp7H1t21QClmvyA2OFFy9JzLhTWR
7x/ZPXBhzq/TI9mj1n+OMVeF+avthCcLpsuS8J+c6/oOozHx3/LQr7PcM/0GVPqjdvR6AZMkZI84
DG7Inbz7dDrN4bc9gGYshitUoANep+3YFWRQyJ/4JaoIbvUu0XbQeku7UQwKruo8T6dN+WSmUSNO
7vFwopgG7dsCTgz8Rzh9UpeNd3NCWGGRxV5ZUwYKkal5b4P9u2XTULgXIeqn02cfDWZNublRshOY
EoK3u21THgUYXUUSzS43ZkXCHiM3bT8/oxdkJxIQdhOVV87G4RhY0mlKAhVClbybQ+JhLhLQBeSX
AI8vZHI2qo51DnjZSFsY7CUIoGrgZ/7X/PuVVGCg+ssdWRMKsvMBucfzweti/jfV3/YO9dhQuUMa
wEBUeynh0ueaHkCpcIlfAbDSi+p1LS0UKzauoSvxljlgWFL4Q0yu+RCWFak69yejkGq4Ah6MaX4q
FphrO1XXSDL8vd6+QJalFdOl+gk7+Ixd5BRmPz4hYwDZMvKezrNnwvrWokWqf09HMDQGC21RAoPA
7fBvqz6WMPT3gI6/SFSE6UI0IUjXWCp6a7+BJKpKjPNWCjHZ3zIOBmwGZPEyfx7SzNSAE50cpMcO
17RngVB73saEDRH6UUWLr5vjU/GKgq8PN4BGjEb0cphmvSn+1f+MyYIxYF+Smi8c2dDT5UftZATr
oNUuqACvGrixgVi8mUQDirHeOgVtZGZW//qM34eZtUg2TBHzgWYJnTcoXwgU7Q1dkQEN9riYKCuj
hJZxEvbeIdXZCC/dszr6n8ZvnLhOHqb3jP/116eV27zGDdAcdgenlfUagwHksXaW3ugAtx4iuv8M
U82GA11Qm174ze7TA42rqqUxzHCVuf/NSFLVmFkpJZU4404f3ZZAwBGJ3hlLsSx0HPsK68iFITa7
P1e/p0BTtfTxAnRvkEXtdK0KZUI8Gt+Oo1mt4NWj3+tJsOo9MhpP31uVw0foqRnEFAi3H4/qwXH3
76aiRLTdfXj+VE7estMCO1oQCkNjjwNy6JYXJtsjkrr8xzPp+YOzfDiqCE+Q/FnsjOtrtzTTWSVy
plrKmcCw7K46nc1je4e1WETTxhIC3IKNjOnJWV1EZyh7evb9hLY3n+6Cwt3OmhWmsfkXPLIRYa20
swrEfaM50nw5eNkPfNRea3+aZ/UeqIfLe3E2nI9i+chD+k76J+dxXKWdV2q6kJ8zfxemBy06ra5T
NdcN1QXBYUB4nuy34vajpsaR3cuLRit7gzHOPc5SrBEN9moZTUIMeWvD5SgeQ/DCFIL6XNExQr2L
OJDrq4w9KRGHVuP+hqPEsVue4CwPJzYxCvQEJ3A6im4utparR5Lonux4xt1KFQsQaGKtv0umcUUj
wDDld756emQmH72YZISt/qKeMMEwE1Y6U6vidCjfvYMJhaLHY5AfB9OxQc3TMjPGz3ESD5IF6+D4
mXPfB8GMBCDrrBjdIciLKzj/pXBol7QQJEEVzdHhGhCuS9E7UrBubOM7I6EDG3BXy44TeJR6Dm2o
RU0fDMye7iuO+gImd5u2Sw/TcFEuKoKPZvU43Rmj0/ICFVZqF60tnm3tLFU6ZNu319fzYELtiu0v
DqvM2U1Iit3qdrpisChi7EkUcVcW50bEOG1Qmvyi7YU0naf1Fk948S9ZU+0A6WyqyVs6E6tZmG+N
6OqYHweYE5DwEzWs4DHpMDF0vb1iUJHiIsxYjtUhD/1K0Nhm6lnMr9CHpXX8CmIj9IkqDrO77qlp
dQNhnSVHJZhPZ8mBhpRf5NqL2081j/3UZNTX8KWLx2v9fu3kp1oFvGFKZ3kOa/xiYZ2m6pyE636q
Y8JCU/UUVGJkNph9pphya3ozCxhoLu/wWthzDP1Su1d9IvNA6y4kjFsE2/9z/uhN+QHf2J5SbA+2
nLVVuX5srMXmsZzq1oaJHOLBhHUEaO9dnZr5G/8bcp7QNFMRj2CDcAMiQSnkQ4kbAX0rIPSG7y0b
7hzF8M+NG+wMeyIYbK7QBm8GbIJfhxkhI1wXH1DDtM+wnoEdG+ONTjMYM7KIaigmcnlKNGzcEHH2
1BgDXQd6tTG2zYebAYom6xzS/qmflAzivtO6uqJqSjVp5Igyjmuh48qtZUH1HZKE9uk+gIyKdmy1
L8oTWkbS7ee6PEgAHM9ewa/i373BrlRj4fvCvs/djwRE5F2HdjtruOdWCJo5wNFB3xJEjMPrOHEH
ob3YdOUHrnsNegnKc5Y9NviG39vIZvJnl6eLxVTtCKOxIXAASOyyo0BL7ikd4N3clW+Wm8QosQQi
hDOcTvXCp+NKANADxvCt9x9O3EZffcTj4q70D7fKNEdf9PY68zqTr4b6xjz7Ss9wllmMZtw/ip4v
xyYjFp2Oy1n0p/mxbGdaxNgK5IEu307bq0hmlR918+rhaYVre8aI/p4p4QwQAvCao6XZVIE93VRQ
HJW2gzK34XpZV98n4MEjHVwmMPzwbdF3TPfT1nwdhlBe1FN6hEUZXb3R3oavB3TwgHLPnS3mw7Od
KgGIgOZWJPucSPolafgAIlm0v9eXPs+IhEsmJbw0xWlHG07ijNLZdkc9HXYqU9ET5fA8Pp/M2YpW
t7V+WYaVt+Hf3xOxwmL3SqPBqxqUJhnVYY6eAldBQX+whE5PIlc4a6QLbP+B5eEby4kA0Wag7q04
b77kgaxw268jgcTZw5P7mo468wS9UJ30ijZl21NPUiuDZz2zFtyruVeGv7exgMWY/Y0QaS9KZ40+
KgRBD3hLBAScCL69y42w6vjnaLBjUzpCwd5fdaL3cWurrLBkwtBpLZCp6L70A65umvlGlZZIas6X
WE+7/HmUyn2x3kUpbqQ8C+18/2gGynS8vuC4DxiZNiCLCj0EFAhyMEYzjAHPPs1q/OuYc+HRqv1U
PhNpWGp0vOTBfsH5SxXcOicd+f8KfZksjDtQqJVQtgJSM/kruAS4WGKcqbs2Vcfy0bMzltSGynPq
YTmwNiBevGXzDtBV1N8n21NRX+u9LacuKRl/RPV5q3I217XQFuu/wYqcIug9YdvCCOdVoIhFmyJL
puTBqW/8zr3P0zsgULqiGj53sWMu6xGz2ErCp6htyxCom4G+0qXwdRIzuwMKqTav9xkj3SOVfl0L
epjLpbQfT2P2aeAUCwdsaLshjSNKqZtaDO3sJZ7C88yQ3varicujYRA+q5Ja6We9qUj02QsKg+jR
7Ybqa8xHNgUIRAXJfulmttsOd3PEN7HM1Kj3Jwk7nbNlIbbfk1xINHPspj/T8cnOm8qthRdWPAgq
zA8Jog3kuMojATG6JcNu5cIN4h1inOloiUdB7BH1uCBIdlSz+O5h//Sy5xZ4JpAam3uGLs2nw7Ds
jvUMfpvtoVbEPDuJohfvl94Ybeb5JB2Edn4JdAGwFxjI/pgm06o2z08/cx9PIMqlFNV2eOTrklJU
ewLhq3UETHCydmitU2bHK3BeCa8BsPa+yaAQzTnp7yiUI7koq2oq90QDuH8/X2wq0z3UARKfJiRO
aFKsYcCXC32iaRvFmCmBOP0YGezndzQjyCkFk+1ct0D5PrxkRko/2GFTpJfFqRoKOkJBkuXDVRhe
BRZdFJZ36q8esFn2WsPpqdpoQa6kXAIhGhkqIatq722F02Kw+PBNlydoKvO/a9qOMjnCkU+S79Uc
2pkTT2Y2TypiAofnsCyK7Vvon7rKHYox8bFyl3RAPlXR6UlGYapi/YQcvNgPpFFcLTaWzbwhLWpW
O3UCj0lbBEW5U2p84KcirOKTT0J8YoFCEZiulqZQ90zEoxmJffhp6EXZzljJ+SZm6il1VsYUGDi4
/VHd2bijPGyDsaPPcZBoDSQarn73AdXAwEK1sW1q/3NQ1fSOqGgBQajQ3g8dx0qZ7dV8N61csIxY
fawE8/3hmcQx8aklmXkI4V+WOyTT841A6bKQyCnqeB6xl6dHGYN1916wb9B4bR3QXgehVbOFAzUM
Vw9b96zTwrnHBDBe8rsbePr4L/dZMihIU+nRhLTNQVgTuM7AJXedhAE3fI5isVz6mNNs97GPfhxp
LCj70POHWqFu3ybBdOD5dsDT9BlZQgTWRiCm2phNHKhEcAEFJOhVYQYSl4HMZfW7r/B1Zs/2sxPB
g+8LyJzYUk6nlwS4rQqOkmsT1KkNS9DGObpNMPtTF4YWCjQDT3Saz6nHmu77lx6fRSUt9l+xgNHM
NDDvBtsbnuY7Er51nfTg0DltmJ4c22ACezcH13FgN+CSXzPIglbbXvsoHOuHZ6Ihq7FfzJZt19cN
SQKzB4BZr7EGdUsfD/EkZmIDnniz7sapwZ85i1KXwQIiXmYDvjqvaot5P5/+rl839UzoLJox3vFh
R2ZnAns/io+oi4wO5Ibzp3ubHV2klfLRAu3sd/iHqaW9GEGN2tqWz2vNXSs9Z9w68LFzfsEHPyPQ
e9v0+UifYNUjdLEmsSW/QIp6o1/yosnMPROXRtVMhq5N0PQUKJPbW6oqpz/ZdWTnHSow3l9jmJ/0
0iQcuv960SkDSQmSkSoKN+xBpKYfiGELmKd6bgAhKh6bag9BMqaRV/75+wSPgQT1Cs7EpZTeUw8o
UGvUtvohmadnaGVXgs1hCI0eAgFLjYXrGerpUK2egnPb5Dx1XmRPWLZSnna7z8PJ+Uq+sGgwKpaG
Q4CQOK8tn1wybJXtKULq2M+9Dz7yLeK5KT8Lt0TnQnTCpRn2KJPpGC4hDqYj8HXvDE3FV4OgRA0y
TIvEr+36/pBTL+XTnyxs+aFJXkr5gTv+vNMR0T6FfE62RECqQrupzzsHY8WBzd8bGmdxfK10DtYk
zIiEgRlXuKisJVl71iLOl0vdnmQ7Sbq7OPt4f+QWAk2ECyOwYGbDVqGsjkpeT+YPjmfJIdgIFJMh
k6nFUfym+lWBoeum7ioLwnoNCqeBIbP+2ZhTWGLMe/aJvRTYEOxypUC3KeBjPCK3abaD11EdMJf2
k8RZjH+KQ3HMSRxt5IR0gdzqbVypS+M9BlWJYFLTs/qNXKZvI+op08cqBhLFptpLHoqhL6V9oGN2
ZmgoLMCWPAsh/Je1W3RGDSZeQMhYsGfXDW4+R8sDuO+YG7r5+QnhxSHLW6UjeNHcWRr/jwamgsX0
jPQ/mSpjn8rHatHDECujXonILiWLHxq0C+EInO2TZWaqjWp+LwPgw2zJnDRIEqQh2gl4SvzHxrPp
3qU9euOg+8IFJjT1r8OU1Oa3NY7ggs/0YeRkGUGA0LDXBhSbTG9gvYvJjy7ev4oVAnfcTOk00Aqp
MvcyNxRlhrRqGdCGj+bPQY8F4prfs5bGWfIbedPklsQO7GSTyJOlgoBOHO5oqtwpZCYzqwSHL7x+
zcPZ6iTR6oWFjrM75BG7DHtVWRmY4HF+wV0qqPf5iURZR5kpkl7asqkynb3isBDlUwjHyva//zBS
BrEStmHtXDW9NTKdPdIMl0j6EM3GRc2aBWjUXN2blkxQ+WtWwqQoY8C5c6Stj0ZWI5aMOUv1CUO1
DCIOV2QDRQ1747XuBhSL4FS8GfKFQqNLrpXtyPGeCj/h0YftljEeyDkx7iG59+fiO8K94NCkqXZ7
Lq5nClFxOxxShnBIXqZ68EFvtktlFKL4yC7gt+Rtn6Xi5xOxSPzvQ3k3jQiBYkBzl/oqY+RlSQmB
/xiCNohJM1BIMuc52lQvq/PtPZuillqQelLzv6Xud+UgK3QBdnTcwP19T7/JWivig0ZTD9HmRqXv
kKVKWArczxmdtogtuJ3NCCnxXprZUas/Kp6KWpMVIf2/7SFQvra6BCW6feWpBIEskuspKn0dRWsc
KZ0WIg7qrATxjVELWLrxPzMzCtU91Fr0fqX9a4/OPwJQV9NnjPZhhXAzXiIxj88OWk202FcTn9O0
h7dJh+zYJYeTs+CJGxuHX0/9Ha3m8Z2THOw2fGkF9u7u1U/7LCUztMVsIMTReCoppUK6pNbx1gir
PfbmhVT5WPpZxWuNp4Jpq11dgGPOfeTCptw+fK7nBBoAql4oRpbZqdAjvo56/0L0gD4NPk8/u1QN
VIOQsQjwFQOQZU/+C2ZOw1AZerVCkqHLbjV0E/q9RKbgJae+WAHfZvxySnApszip32kEL4GBIa0l
mHqrYaduzO0DSJRValVz3E3TDjuOuDENxju5nZdmn4wWtLLiUdCEg/cb1liKkljIcxvPItOvRZAO
CdDp94C353j1iCdM/Yoc0QQtMwGMRadtJOHdWyW1rQB5n5SyMnlWw8s0yTULQ6YjadU1id2Dqc+P
xcPPFGVfdCA8JtMuXU75YM3ZxK6B+8PHDoIqOWR/T9kqNzRL3fLm/aBjlW013pAtugYq+vLKk6cH
5GiOdUv22sNidTHLYRRef0saQBENZj5ClZKMYUIwl0oJ7wrmfhqxCd1zTJsbx19N9bnkTflDeq5X
rmEPStHtAqZf+TUnesgRoWtYnvT1dPysFqFXrjjXZgffUQ07NRnnqOdfht4+MS/YfTvBqZOyX7QM
z4NcbE4Fa5EE5Xs5YCfzlXD+nT33ewLG3yyH4kOOxnQiJtG6mxekXO7zKF6Yz0yJXv8bNtFGO41i
2J8HqPuLfJ6dVYUPT6KOzna3otDvIWd+rzO7CEw6u7KPpXFEoZRAIPIhZxm/pEw5bI2SgON1D7JZ
f93102iev+jR8TM4cMISS6962ZrsJ20WX/pIdP2JVB93gKwL1f1+6fB4fOGfccIK1NMNShPSVKXg
weIsXAgs5cBOylL7SwKQnoWf6AabCY6u73Md9vDhFBPANpVjULsHfzchNnkjkZHEckQ90JPOp785
oU6cnke/ycOnx9qXGD54AzEygKyGOwy1U2vYzPeMc8hJDgdzg8o6s2YJhs2Z9jz3MmbiFI6I5PIA
EcG9KAE8o0TPld00Lm3FDsVzUKbza6Fh6FZpGbyaTwDQ76o/JILFNxtvRuzv7w4Lisi1F0qgSSS1
F6OgnogvT9tw7C4kII4uUfctr0arSxcPApMDAK+vlA1TJx8Rh54o00U7t4SQb1o6hdWQ1rPg7hiI
3vIT7EeOG5oJ7+f1x40bPdhqRKnmVJVRvDARL85Zs+8G+BsR1YXimr3bSwdqRr96KJI3MtX5U/8o
ZFpTVbHlIqV5WZnyFpYod058eCz7JDf7yT5N6secbX9aP3G/3FnaB/OAmrX6vi1YfNGW05/8CNYe
gGacL+gnuM/4IXf2LZKpoybei1n+W//Vvo1xC0ZanjChK3gfMjY9G9BRqg9q0eaNy9rIzYI9yw6j
w2VtRyrK7kkP80qrL9tpZLAJ2H3Ojv8/fY2quRuwPMz1E9P6fZlPZ6bQJI0jqCsQz29BnBEA3vGa
HN1YhkTlZgMlCT2oGnsqYIlOy/sLnbhcKax8xHxEGoYsO7OEWPijOmAAqm2FieVS5WspzQbHEwKb
9VF1hPfIk+AgdS3EYlxTncPo5p371VijNW0Rsxc2bB2H6JQP0G1w2ippreE7RxdPdObgsBTXvZe6
ZzBjhhI2nWUDBdJ0dbNboVUV/27v/9OJRY8nsmOXoUA5gkFYGhj1pxC5/DjyTtLbCs8PH/KkxGDe
XJ33KC/sQgReSi6zvYET/cr91ANEsfX454JUWGACY5UppxTStsqH6WwyzP7wr0ehl7Ss4hbLf6nt
gPAS/NzWnQrdzVVGIQk7UjG3a33TpT06SRfR+5nII++UMCbhuWfPuYSAf9ywqFRWnyDwaVUGhAyt
wLRk2giUH6yHODq2UPWoXVnHScHHi9PboL5dpj4xaiZH3rq01BOLb1HPzvOkoiDDqIUk4IMOy0jT
MaymIEx6fjyxXAklRb2oXN02P/tnkJvZcGN2U5M8d0JEQH59WEcHKW2gWyAo51YrVFF4CQnNE+gW
BDqdcYgCv4jdwRPy0e6RM9UxeeLZ/GzChmwci1ByAkncE6GdMLx3/fVMn2tFPxKZ6SDrAanmPyqH
jJhWwLnEhcT5ueJSDfxBPPLdbbAla6g51qNoDP06dps09bbLO9WM5/xSltQUD73CJroxbLlrPote
CbGGMVBlzTGOIYrj7zxjHUWdF1WXJMaojz43K6B68ZnQJy0qkpUg4+GF4MTogsnp+KSUhNi3P/bm
wO3VBjbikn1Uz7PXSM77oDK5c60FSr3c0dsmHSB96NmaZpI+t/KaaoF7Uow/Z/c+LWkMyobHzS1y
ok6wTWjMxg+DungGr8JJSb9Kjt6pqcNEdj6w+bAA1x0Z9XXCCv4qkmlzIOVo5uPRIqbaRHmhfE3u
dicdymnU0INBl2w/BiPeUbIKdan90Y78VUUTg6arFl9d+O0GcGjPMm3ablD2vWJ5uuslEj+r3cTG
9uvL46/PtqUqt7YYxM/QBAwPi3vqzty/6PFLw/9wMIwosHvmkslWiZOr1SnAckOAIdrMRR5TyOyt
RrRJa/YSWr0PAxrtn3EZJOiucat/ChtmnTMCI5HVK9wc7eU2bX6XD8acKTm+SWELLTHg9wFK+EHG
ja5ndHFSRmEA461lJ5jamtPP5+suQ05XuPGN2++ZOFk9Mu49nPD4PHQQGZ2/CSaRGf61Gs796WzD
PsaCuqD2rMTE/REyGYs9Ygd8OCeR7nEKfLKHzLHgwj66OXKr/h7e9XxNQ1wajkj9r5GlT5FhyeRk
tMEjUUTtyisTfmlm6CZP7MZKJP5UnDxDQ086dsHYO7r/03MgtvvuhU3TrufJ6mwhbMQIJxByF5mw
BnJVeUopxu1OfXp+KKbUnTVJ9Cr4gIDTS4k5CHWh11tkqbbVX5xiPLl3bp3feEXBubopm+7i+x6E
iJVQ48nI6a8O11nh1Ajh0mlpleojDfl7JkAQdoiAochywPrKC7BAzYfdSoPkRGtG8haHk2J3NbOq
dehmaCzLMkrcFIgjm0OCB2FMMYiFTgSKprNStoG7xFJqD3vL7F7r0NxsOU0zGRqKgtBtyHSRfTPS
tdqbhYea57rYeHS6IBkO0ojM8EPB7kLVdYeT3vsHKEd+x4xobhfOmahO/ma1JpgQm2pArGWgwhBf
2+FL0umy5S2q1junWM6h3+w6C1QUqKpO/hTbQbw2YaQmVwfS3Q2MRociWPnrL3fkgc5x5HA/2nvn
HysJuNl91BuY4PYG+4k4a4ONTS88nSKMaOi0dAZqmLLi3inoI5s6YE/VaA9GcHiANHziviHnlEFD
OhHgst7ujvBiM41r5/RqwTw8H8vIziNKWAp0fAOcX83YAc40rRciHZcOk7Ts9avdVSVhYSOJB31m
HAw8qWIk//wjXq/22DEaYRtyOF7X+l59RQBvcJD4b1BigNF/SWHUzQLdqX+f8HY2s2D/F9jMeKsq
YVyrjEglgjb1selguQP/kprni5TY7kaIsu8W5OAf0MiJ3uz7HYtOC9+2dd1pEPtALM5kgJ9ex8zJ
OWGK+5h3zvCniJrhi+Pfz1QQVvS8O5GddVl1n4Hk6vhZA4S/lxDThF3/7AzTgGkiRK23dwFJUqfv
4EsCEbZvNwfFFaMW3eGy1QWbIYoRtaVorlSGYT98EWzxc9z//ALecRd0sUo403lDXYD5BiCA4+LL
YEj1tW8na3xkPgHNGk1ACKT3A+8p9Rr9o8gX4Ac60D3tCBnBxzcM9Q2T1EXro/IuBHV3ObLonp4r
RlZjC6R4+BBBJ2XSGUw9+KMGo83IaZbLAI3wnTOHlt/qQb0n7vqKlpsrdNbK64f7dB/zQD2K8ora
cS/DMYCm4fQQWXB16WdO8ilrQT6Wv2jOVNKLPhvd8xPsC9lM5nRvRa2bxHZfi/LQHmjc4aAzVHrc
pa3i3QJUvlDOWv/UAFvyX3gqvfxlal3HFEvlC56yEFFXsUlbTcP6uVdlUJzd2DfNoo+iXPXxsJNS
ZnXOScsruGqgpZQNC9mD6sCORTVL4Zsyt5FezmS1ek0jqtIL++0MNvcQJEOCfHxJR44M1DLv6Spz
mSN9qBb+4y+vuQ6EF47OC0qscsoQDV2rXUfUo7NZuvvlBmwJWtw3enGEjGs4UFBlBLnmsoGF9S2o
ElVZdObiHNOhOqVEA2+dG0jKHKxrvXSuAKsmaZPUD59JeJasIi0ZCqCCEJ/GKZEQRnamE9TOgi1v
Xjarif/DO0LIqdh5pC2V8jWNB4Ip/5wIVUdwtR/Ydcx9lgwyC2ZkJymKQ8kBmolCaNMy2hqO3H0B
7gDWnz9upBpcw/eb+NdkU4CRXq0JlhiBXdhurhEO9YN3cjl3x0HrpH6R9Vh9uCW9fCv8BNQsK/HQ
MgzyTiVVj9DrJ8ckKAC4KtLNi7G2jERzCiU5orkfSyOpY2r/0m/OdtMY9ekGZcqTwCABgm+S4Cn2
pmmX9Msrkc8R42r45SoeI6wbKbP/32PFoWoW0PUG7moRA5BukAAxlkMYTV9ZUsfJUeNLhlN+JREz
Rttb/l5jc8qalETERzzyIBHOCx0o4Qxp68wOfWFHdNnt7y5TDF18rt2ttGqBYz/Jj72OgUm9Zk0S
4uGv5Egd4TowOlC4CTZEON5yVvE7EK0J/tv1nUSkoC9NHqK5gwkOo9ewUh1WsU6AaswfqDdjPKZd
jyjEAH5/OOLDW54tz5EG+hqpqWyTBbVTLZNwnA+wi2f+j1OemojlyVSOHy1TnN0RQD5J72UwfIJ2
jCz4Ffw11/c6mvg47LPywxzmV/7V6NNqrpUwebZ8EvULjZ6/oHZgqz1YugDxmqPa+wARfshixoDF
bZ/XEJwb6xP6fj6Vkjt51U5CkSoBEpZC43QqlTSXEfHjBUDhWAdLwNugX5dY7hL1nqhcH1JOggtC
u2rUbiOvzG46ifktPXtLgiNimY1ASumPcI5x1M5KS0VJtFxxzorO1m5DofZ14IP+fw3JnFO8C/3S
L4VMFbHIISS/GUeiyMvXzXJzEyvEDZAk2qXFZS95/Xz1A5UzEQAojMOm3By2F11bmsbLcihro/XL
lVjxh28/IwVhXUEMTLQJS22UAEGcHEBmFUJjolpg/ki4N4VoXzvYV3HnuZR+PssZs0OGyKkEACyh
EGES4TGrllKoWyxdXqca08KzH2P+B9XT8HebTHcJRWiqnDzCSpIBWejK2ILmTOA7VnSSjWz97MJd
GDEHw8IRp3Cc0Uy/JJDrQnbEIxuIhf0wlgLVhSqLwtBkKWgZqWiaCA/TdbtKtOfypoJLo8Gtjfuz
xyFBGhfZJx/HsTEfS23dkHNwcfY0gN/O2N4JjvpdAmH4tlkigmRNh1YR67ueCzJ+w5OAf9GVb/rn
M8DgDGwCvOgCFfebKPlik/LYjTGLdVBO7fFsc+SnZPw7+PyyLqERwxCsBKztXsAt7GoisfKToQ5P
jT2CfyFKMCLa1QfrOPf/kflYHmctDLRnepjTxPg2xjQMuYXRip500yfz8l9IfjRi0IIwwl2CZf68
AXblqsm+Dlj7PZy4Tefkbcefh1ZrykSAzbIHRA3iVVT+chzuD8bVV5UwoalrpGgr5e7Tm2A2CEt1
atfMplnm0OxKWchKBubVvt/SliT59WY2It93SrKnJiAQzULte01AOLM7R0jUti0K1X0UVOWmDv17
FTEnuM0+9HINia2x8aUFXMpNtrImfdNDdiwMBiY1thQz9NQod4XD56VJcLzwS5xWPlY+/SCbNKpB
QnXrXwUEaGUZD4G/hY8keyX+oSTvQWJc89QXWXESpjF8eJn7TvHDUzRzNmmFOFhKeCdJkO+LFzg1
G1zowR8kkM9/gIaj/QAOy+EcU+STmpsYvPVWBL22L//4lX1Wk3AJ5j1fFrkJo5pe6QHouClI8CqJ
pS2pPkjmQqyThwuN1sxji9uRPig6TwAdgXyaDBcpAeNzQ33HeybN7rHiqQNJdJ7UV9Svp2y1MEp6
6OlYDCS2T4oWbQtApUEurlHntODbAzOsZDxOfdAKEYuEIB2B8Y4w6Bp2mTV25wsIBoAwcHfoI0Tv
L1VPM9Sdnh6hdFgqngfTUGhmhHtpI9aiE1VctlgVUA3NgiVqfamABy3YTKjAyW2Q9YEjoA3Hg4mq
RMjqrf3QaWz5uDCPqjG2FyHlvzo+lHTeHO8ma9WyVMs3tJr4C1cNsXbG370/jGAp5O8wLg5R/Ago
rV+BvfLCU15qlIVjRkl8JcCaau04aMvLi2Q07NHzpKPXocvjr8PvbkFpvDI2Cn2lsrHGQrVBcg/7
537yQft7qhRTjE7ioqtItmt/A83M/nrFY+bseOXXcBmfbKXkcBNXvptYujR2TCaGy12URIZRxCSA
aTXF8Gu1K1VxQPUKrtGRdqJWT5yULhdLT3+rJk47E39FPVXlNgPbK7DYDP4hbMtI/YxHt8lA9H0d
pXtkXdZBp6vjSBN2oZBA01x2sgKzH2xB0Cg3X72TsxhDV2CPuMNZTWU7maFhbqw3wtd8MhE8ayRm
Np7mALprgxawsc4XJemC+hoFEjZ+x9NNG2Vv3ibLI1dDFG8REbwJGlTwAYf0U8sZ923xcZjECtsO
7WxFKTPBBPmecj6HbjdDCBu7Bqy9naq4K+Exa7pZKleiLaiSucgSXXc+XSOO0Z2BQa3qfK4DiVah
5JiBZxTjW4FU/sRZ3/aDILJWQLsA6ebgJLxbd7VsagsX2mgXbkqbbjBR6q9+eYCj8GwKtNtkQQgi
PMw8jyoNSyVEeKO/RzKO6tTdW8hDn+1spZGhXvjNoRe0Ndv5sW/l/rUVYTz2Nm9gRpfSnXwu+SqM
cDaKZGW8qu/95XuNNHkQu3umwre51y7rGvbKFmeYMN3HGBYOuK6uO84VQY+vAfdh/ELQrpTylZim
abVi7YiGlWU3ctNS5ZlPIARGMl8s+mQA4BX8CGyl8jBKLSV77p1/5gJszwCglg6qnlbNgfMpm5A0
tBj5r66WBVVI4Nrxg+7dcGtKGCJPTkPD46ohZ2SyjiDCROiKyMKYT92IaFCgoPqlZ+i46HFyVzeL
zeROKe9ZRVXTWorUN3NdlrVM8BePfi9IJ9OPPH7EKKPrHOn95R/+rZ0xynXuu6CoqCDdjVUppxiu
l8leueJJ+rXs3BAFffDCsHEke/Tzta6d0eJnhY9f9Skq4xzoNwze6ON+JBQJ8yizKXCYPIXgIqxs
yTg0q18xa6OKW4Ue7kliQo5WHWx/iAEVc4sbBXhZ+0VWc+BkGUSL9+N33vGRnXVIFpKLpHOAfaOA
GGmoLLwVs3/vxZkVUMeRYktd+6JKkUan/TxWI977DFTtTLqYLX49m0ElTL+frnkWVm8cUqdcGxat
zQhjaPaYzivPjVnd+87iD3Leiua7cijBaCAQcLttPP39VQQcIJ7MUYbqnhApajg0/OXRGjiv8xYw
YXRuyTEdHVjrmyxnn/1sFsAko3eJmuOwsrI8cDZU/mEEh2GZiLEI+DdAqTLdxCJupk4aeAj/t3pN
j34d4dopE9TFqAelgByGFJYlw6o7EoAuFdED8Lhslz6Ix0uTDE60mKA8gJL6wsUNwYJZtMq61xWA
7BD+n6MBfgc02q9Np/b4ibgRRxIDWlOMd8Ak2G6wXaamPuD08cGdG5rHfryMeyW1S88dVHexF/HU
tbGzB+/DTtViIS97Ygm2nS3Rbnmf1WMquK8TUVJKTv+EEqPE0BsnrT11IY4GteR+uDjTm7qqc9iR
+PNoABJ9zjAOh3Rd6yNUWmeYXBhD4uPjuRWnjQ+K1H/XTq22aMIumE/88gDxWq+RgqbwBJDA5AWS
JPxJegseO7P2aQRIwY5w9iE6RH4Fh8CjmODVOcVyQg3EuEZLsIiLxH6X9sqgtfL6MWtflDuUOxBN
02AgbIfK2gJziDP8+w0SneCtTF8i05LUEPIKN3fCTtEPtZaYeApTFyHW7wGomMjtM/3UI6+N6vDl
PcPNZCPO6zn2jHIhyQKq+1P6Be1+6q9wDj4oUbXj2cR5/Bz2PvKdwPosWzBGeJ17r4z0fIHRPhFe
iJYH6G3Ef7KMeBw3/W7Rb9VjISNs9NX6d0manfJ2a+ErLWJc5m3A96Bgeux9cEEGkAIFANycV3cf
ig3Y80MtScevvgiGLPnLb1C87SrDCzdzRQC+s3HixoiGXIHwriIenN9JCW9SOy+yGCDz2BDDALgg
Q19Kwy2HDomOptkr1rgEDK3f1fTLVa6iFJSPL73TzTMliU+MjWSPwGW3cN/Jz5vYdUk5D36BCd6c
PF8kLSTjlukVEPbaoW6aYym7cC6APvQT5Uo6B2zXqXWOI1a12HpSGjqOr6GSXDddq8+kJpHZfnRQ
SEIF0Ub1ieF3DtE81qFLhhNtpg2kN46lIpFvQl2vaz+IyO1jPMVvnJRqXllqwmhjs6kx09VCpsbo
HLxegb3jnJmXkkjtHozhoU97qIf4mUjDqs3k0RCzQIFftY47SqaKx5/+O939eRB4zDjJ3VNc9mf9
PbrNyw01r/31Rj8O3fhQ61Jmi47AbqrEs125h05P0ouBl8V4RSSR444iMSVkA1s4j5AWMilOn4O7
21cbyYB1CmfZCRA62XlkcgCH3i6rueQIz5PfOou0WFU+GC7cwk/sIo4IDTaHAWRfklGQDrw77tLh
C2dTvA9Fz20CHw4gqEtfTfSO6gD+RXV0fpXHqmTEjr+1930i+Zb5/+b9rMNUqq1GBJLQJgadegO9
ZQp3180+779zp+422tvIKpqQTI6/QJoznx9ZURQyad+OtKqIxo1VdCqkSYZEue5mNvavbzy9htyL
NBla0+ImzKPL4Se6qZhdce6KCeuXQPUla4WrJqbEsxv66jrMrH14TRl3oTm4qkBc5TqV5sGpm9hn
uEyCQLhkhirYghDfSsLh6WkR7GONF6GHqPlNx9AZo56EK6Frsr5nOQDaUb5pMd9x4S49mhzwam8b
2AGnlQL/Ib8td9fLE0tb3pCbdOtM/uCBMdYzFRxASVPPVorGlts513Wu5SAh2EztGsEAOWHXIS5g
b302+UdUzkaS09qrx3fmwnV1ERWm2gcvOMr0+N6FiaMI83fWGBwsV7Q34vVWUCB5bK47N9ubP8Aq
Pko7HZCsRmM+b2mEcpJX4ldEkqrR3yTCsh715dmZaRy/Hcp1u/9g86tkwrh0ysVhuPf0GMWuRXBR
7mLLDFo0W/cymmgLFHIaCGYACReKZYJnaHs2HHaaWKtNfn/4lnXGThFJ0bNH6exqv1iKdjGQEW0M
xABWntTHF0FLu3K7jFHA7qAT37/dpOZCMXeuyz36WlcLNE6Z1ca1onBnBy2FB0S2PuaaInvEC/p8
Ty6X+zJzCu68gQLDmZ4V1b5+yj7AcRuNZq1VnTTF2k8VMflf2gG44pVZCDYEn8PN72H4jOrvSTWR
9P1skJMjwOt+gTM5ETvK+AJcwgJnwvU5jAJAkEe2P+5LKmtQCwUnl9zFdLiG8TTDyIUrE9cqkve8
v4NWI/jgUlVQZHzlsVNV6KEd8ToUYJwi6+4w5W6TQziidEN4NTsscTtIQR8kHJQGEBc9KZ7FJldR
AvHHLsCCm2/XKbFFwrMJabnup87XgOWz76DFp1HDi8hYA1nnU7JbRmggUoJsCpjUX8EsZWJq4oS2
B8+hbNPDfjcSoTolPanenZ0oug+vptjkjvfy4caz1lZJIPirHfz1lf2SIYcHJKVrVr61RDE+TEs6
tA2mnKv9ni2/HFcMYDWE/VZvhYL4813npSu9Tq7FytJTaxM69U79hvwG5e4a4uJophA7gguaVybA
BdjsiYtsbXIOiaZ3YL7rqQoU5iY8Li4w+ZLOejLX0VkyWzT8tIP63v4CB9gywUH5DZg55nlA6QsN
21LL7ol2P4QZxJcVKek/SpeDvHlLFRnFiyyAljrhdu2IvJE1Ej3xHB0/rSEGfeRosiue9DVFDsjn
ZcRyQG5JEZNA0gbsJJiHqNDwgOGORdkAIiDDtv8ptYpAhhunc63zw1cNgitM1xiW6eAiT7I5c4N5
UpMm4Ms9dFT95fOGykzxff4yjqphTGU9ZWV4uRhnBZvRTHwTBu/z8vd4fzzJbr6idU5qSuLIrgFB
uoHlIrg6A8NOAmJMtcrt4kvtVUvbNCgaZuSQYdgUjVlSyYTavoXqC3d9Eh//NarUMGGyrPh4mWtg
Gxg7snx9V34SVIs4ia9buExT/IBC4U6Ib0ajvgOTS2mTFyHmMaMKeNylAiYe94w+/8GT/dfGNyk6
NPzeQrMH/ptsg+sG30NckeOKz6w+62rdb45VH3gXJVfg5b1AGBnw7NcAxmMBiKK/6yRNp79wQiKg
BCOG6MZiiH1UdYD7NobbTn/S3c5zYla/1qKReHXSSpmgTQpMck99rsN3fnLV2TDWWa9fh71eqHGS
KhOjfX7Sn6G6BsEXvRtMLsXi2sJGVcTcQ3TrMAhBxmntU/A6Y+1VfX9yc3yKk+vEXtq50kLFavwR
tsao4JT/kDLTik8rBtkIwtP47XRprfYM8/SAbCTXMTS/1DomTcLSpTzj275h9MTUDtKTmqWQQrlX
Z61px+FH+O2f55w6O+mf1OPdaTcmxh2NHodPyLZW7NU2a4/FDL0aj2rfndh9dHG/S6LR+ApCXAa+
d3bc36k7GoNkdctx/22iCP/5dkQYrcvedv5a4sYt9NSD9svk3W63OIote/mP3Mm2zihjIoyvpP/b
ceeQp+u7S/uV4MuUfxhio2u7Zwd6PLLJptq8JUPpLFzeY7CDmhzl/QrFiBpI5pX6eJ1zyR0GFUBH
CO+a7UYuYLEl/Q7mt7z/BVgRUSDN2rxoEdAUAZ+ag6LABHnyYMDdtRjDXT/SMrb3Ok5eKVdAf9nw
BhdTF80NM1xrTUZg37UyxiGd2tso5YhLuiKTxrUz7lNFLflQ9Bi/mrFab5X8vRE3+TpgMecQLfIl
W2xK9BM2/TPOiwlhnsaJQNP2IwWh/Dths5tGRk+LDepq5Jb8WBzJKNncMZE1nFGmN6J3I4P80P3b
n7o+LOJVb4ndzIcEPgQ7fzfAG4QtwdCgAOoOeXhSncDn739dFxaeEBysKDsIRDC11oN6l/A8snie
KDn0QgBolF4m7Z73Z9UZHzlY1tCiWt/fIps6pUKcoGxAzkD4FJtXsH7YnWoAXvHV4lJNHuHQ4cTi
xwzRTTz1sY6xrZx6Qrc2yr1wd+79yqKQzmwVw5fbjIwTpDT/Tm3lKyyqrBe1boK9BvHBu3C0H/96
TZ5FkYMWxAdIoqPYTKI+YQpE7iAUKG9NffCUw99azfVvztLyQ4jTxmBwOI9utT2IeMkj7xyJDDCy
J/tXeThTahTjuZ8Jjd0uAWiko/hKqVBLLnKS+6MjH7mZXk1LWxAarRYvTd3dgPEkPpqAfgStz1B6
1s4bpJTrwfDgbbd+OIsl/9+p8cQPL6HZE4LFwOKdcWTRTNrxd9uuq/j+rtFGVV+stvPSWuTcE7qZ
O9sJXDG/gSPr8MJ+IiAvv71+/NSiX9sORjUE6lup5YWU1Tu+ZGuQTBr3tY+PRo0HyR1+n5sTjQz1
ccWWd2FvBHfyEGKXcgIx8NoCz2hi3YJp8+2JpZ6gb8hdhuDAssGaavw+qHhylvbLG/wE6TuqljWK
L8dLJltL1aDRCS4Wvec+LOr/mtVkA1BdVRLhv8rWZh6RY6o1VeXzD0npOK1tiG9j1nik5c5k4hzP
7FOUFnO1XbxsQGvPUohPiii8Ooxwwkfu7ncUKXj6itI9nKtGbss9M1lXfmUPNa4JpM77fTWTfpkm
0kT03Na5b7C9Z3J8PHceNDIAvPMnhty3YendzPagC6lcOm36XvmKzdnFneTMnQocLQYu+3ClTcLT
KVM3HTJ6p3zuXbWusfzW6SfprWLnVm4IsvCa6BgCMfLtQEJ1Kp2tnOZwQgiK9ZFDjJcD0Arf8B6n
x/Snwmd9fosde41MrRXai+4Tep9d8lf/wG0sf+PdRntJ9hySS+WSTL73XdU8maKjKlv7EdgBiwzB
le6yBEJxLU71LtYHnfvp09nCIQEPTB6RaFoZGXNSNzAGy3whVzY+FeDJejirZtPkm2mR9E7irI7g
gRO4ZynYpjTr8zFpVXVmxMm2Wrj/4F92/9Tqb0wL6okTLE1OauKoJw0nCloVoqyh5hj1TgES2Kol
blux4os4hfY2QE39n+l5gDyWwCZEPhTTZ5kxv/pijK0zupXO9mXEC9scE/Ixeq5kH3eHXqhdrAd4
w2H4h24E0Z0bLUA1Ar/W+cTORmTUu184WUH/6jB1o+6RXl/1JTAH8kgbljwAGs8gU6CiSH6Qamgm
wwxG/tdbX1fZ9yqQc9uzwv1Y9n+VX0/8ekz9eiKcZOroiOnp/LwWS63SgPBpaQJyN4fJruxNHor9
LFcRjZTmQ5HEikndaFIKZuM9Pd91VNMmM7hBVirt3+216zbbLifY4fxB7/p7WTBaJkivJWnGH4AY
+EG1SNGKTQStwpKMmvTT7Qm9+wT2e+mjlwiqWaG+Hdw/OL9SMzHAKGglfdTdOtGHs43jifdKoiiZ
5ujTYx1zDw8JZ6KCqsQoyd00KpuZZ4vMPATgHzCrlChtHkTH+aAnzuuca3dSMfsuceXM4iElF/fG
+qO23d6N7L4jK03wG2AbcRkUoWOD13m5VJj7870Xxq54CBINAa2BLELyPGuxO0JmG18EZ3z3so6D
jxZ0azpG9zRSFEVOPgTlJRN8J3rSkc3VExSz+ykON4HRn8mLVvCm+igI/DiU5Fdyu/aJQGfPa/C6
h7SKIcbzOnVTayP66x7khMzLI6BAlMn8z0Ek1k/kEwUFrYsl7hz5kvAeJ2RZ2pa1qsH4m0j819Ma
zkE7c1HLw4sB+7QA5yrie6W/sOOQGDsXB3UjQ3rtkSWCAMVnYWYmagSQAo9GmmWpRwZmoUCgeRqO
UuezYTsPZ4QjmYyp9+VBxXIcJi7WJj9eRBwFOM3Cms6wE9vBloePejfFKQ9G22mYrHacEQ4PntZF
dEdZEV52bnJ1VNWfzJD2gV3WNcQUo8NPSavUhS/GqZlvULkU/bAh3I1tUvn/9Dx0t2xh9cAq46aP
QMxhax4c7fCTW9MUeszkwnhTk5UVQ9QPMMGocrT8TPfxlvUk8rBd+vso3GEejbBmxmN2n3iigam2
uX2M3RgXm/dkCt4F9f3b1cYhr/uIkbMz9U+J7+2gelKKMEq+/CKuul/UGoJPzffeIHf+lSh3Dzdt
DHn3Dxz3tw/CuElEgA32SwmRjhqkV1xQCRIMBAVIn39P5IbR+RCMfZ1qC5YCXQiKfskvd4Q1QtEh
tIhSaK8JkGn1oE8H76RI1F2ZbfFnnzV7WvW/VQ6ikzwTygZ4pV2IpZqDwKWpQeSyPTYHpUHsdiI3
jHoRjFbhdLMPaoIiXqrF9IZw9MvMUTGs6P0tO9NJNY8lbMhG6ABxn79RWQXZeN7wfzOMV6TFvtl1
Y4DHb22Hrs6vdM/Jhhbm+b+OgZJ/2IEm2YMZ0y7pRrAXh5YoxaoyNCvMApE09v+/POM+1mzqJDdB
B6MgK8Rh+5FJnrYk83lEzsdDnj3+Gh5YBxiCuPtuy2QQjNj2sKXFXDIkBqnIQNrtQoLqzABAw49N
ewzEyN9H8HLtxLFHLc1eDgE/VDqw1R3DmHdDkW0INM0ciy4fUEdQgRR2txgxe5AtaV3lns7Cm0tn
DTh+cWyY72E7dSuvsffGz5iL0zG9Jd0n4OEDaektTOgA7D/aMVbhVfTuWdBenln7k2OqSEkT+4jx
K5YkEsynX0GkkdXV/++vf54NTj0cgFhxhcLbGaSMUYAXPUheifX6IAu/dqvCzra5Ei5x85ipGgel
WRCCWs6MJ2niWPaUPtu/R3IxPdm72Vd32il2ENPusm3tMdH390+nlX7oCyqZPLRXMgR7x/b6JmKn
VsOG5+32bAftHsNRFCQi8HBNim1n5u/CfeeDAw3wGnsxcwYefUE8UUt958MiQxehj+frb/QuWpDh
zRRZF3d1+pIXkSovH66EnhIhmGxzDvTPtpo4mJlfAc1FVvh/zkVHqqUl+Fu9krGTlKEMB7V3qyGy
zI5AilyKlzS7amlL78EmwUFfmU/aPFv1tsceNeyb6dgS+NJALHfL6XUCEgl5fSjyLTduoP/Hu9fO
QtFTXbl/exX3ordQ4DEkgvTMggF9Eydt9TDm5aPqU1TYurHdKpfN1QhOCj49KPBALW97/+FD8V8Y
B28qqr0JQQMJMkID3fA72CrpNrASH0PzkRUGNE2/VnkhbvW4yAmpHLydMII2XOCTa/3IFgUDeiDj
6Ld5Kt3/3jznnwEhyAlTlWZXwYqqzMrk6gSCh1aiRGn0dGOmD62K9hBqTQisnJmvC1P2IWWEmJ6u
ZiBV3Z8Xea6vn0PjQF0s9jiRoTYBwWZ8fXMOKbnhfp5dpW0woPq8SRAj1BsVeKYl1g+3N+8c7+dx
ooHhsEmdcjPsyozQ3yCa+Kl8q2BqqyQIB2mKhocQa9VH92ASfdBj6Tev0ZyRm9OexXbMWIv3NDfW
QxuV5HsLEAKq9V+UqOOOINc/Yq5CqTdLxa1eZCocv5J+3VPptxPtd/r2g2Sx7jex+55weN8yeHWj
lVCphPQoyb1gWSLck/FvT6WUoF23N4lI6DxOsTd1yhVEZpQca9yHS/0Lqu+DrRE4KX86fCZGYCgY
8a309wfViV+f35feMh5MnU6+viYosdg8o3QmAfbPmJAG0we/4sVuCpwzjbdjfKknAFT4+FhkHobJ
URcF40xTWMPCaJsjlzr2/G9mPYrX0J/MWEgL245SkwMFXPPhyCzJtZWPGh1djRk7uwH3ZbcF1joH
pPc17HPGpjGSeUwisSZqBSkYY/5IcmpocK861WXYYtUf6l7mqztoyJXl2GF1IHfQakPlUA4iQufy
yYTbDPzL6kGUips32GBKYKG8UoMetkcRdKm4XPWdRBQSYG+84tCFEXrXfJvNCFiVmtV42Mylb5Qm
r+ZgbIXFyldOzXtzdzXxXf6Ex8qtLuzPVXO6iiHqSkxfYFQBXV57MIEDGODuZ+UA0ruLJuEOSckh
Gx3U05/7pe/xSbuftneN7C6iHBFIDagS8lfu8pmX2ayS2YGHF2JGuo0gMQU8T35V3Dy4U9jAh1M5
gpd8YJ+tUGf/yGDtXeK+TMJbPeJRpsrwLmOz4Ap+7PZPy32i+1xShD/FsV0elMPgGpsnRObgZeQa
9rpRqPnKsOPBWZP9iydnID/RpXPnNHHGUvaONBxWwwmZ9NCfsp3/5vY7Am9Jt0nizUp37tjG5rC0
Kl0OuJvH+vtXiuqPvjYvcxZ8v3uVFwgLAh6+aJm1BArcMiGt64D5i33vx19/QZOJimEjo8YkO9Ao
oCpmZURcSExKn6QTUsrve7SBMWFVUQ5dYxtkV8d/wB6BCcezJ6I2R/gvUJpyuIFCh0Vi99q2RBCv
QIVzxgvdu947Nga/t0UbZK0p+JXqP2t9+/3KQvds6eg3x7mMU+xeoDauS5lT3SyvLxWIh5cAt+5F
ote1xj1zWNmTwqNO7x2KpDUw3oTxDnvztORbw9DIHvosjMRT8HSixbOGQVR/Bs6+CizRqJt4gMTX
25lDePNB5Q6J188B0mifVIAkoT/6LQOEgqIQa2l9Kxj6IXVG3wMRCJehNP9fbIBCmQ56MSiOpvPe
tdDeZf0yQ1asqiDFPnwDRbIG0QJYF8gJQ+v+wXEyiDKQYxu0YLydB1pZzo1i4Qw81cqQcxLO58y0
k2M1uUQ0ndZFECzvOfVKv3hV2Tc1mlc8xi5R7Py6Fecy66izp8yXjp19Oowswqv5TEqZNwnNxApX
4aFY/M55nzN3nbjEG8ZWIPTVUOhlyQzGKIpTHfUs0unnCm6RStZvLqtGdqBiYS+htVbiyU1lDFFZ
eihqHiODjuIMlF32I+O4Jejq8i5d7l3FAV821V8qpB8p8akAF5r/bIhx6YYG0fPwE+Jnrigwb79X
rBKz/2GfdRbkzu4ZBnyttLVi9oeL1Qof812vIeCJQE01W1uEKJqUKYgjo1FQYiw8GQyIM/4ca3jw
1Uh7iE9I+qwzLQ6A5Lnlk3DNrsjr2A/DVl6GC0qp7t3vForN97bsQ1qI+P89MZUBOBqnu+Be29hE
tvySb6dmUvK/6qpHnhH070a/3D0I3En6A8WcWidhVXFkw7wB2K991vx12ZznZbqPzp0lURgAFM9X
JGnw0zi+h6wWgevP/Oop0DjVhua07pHhSUBoXS37ws4oXcQoA2urC8EUD/n7Xtgh/lzYy6zCJwcb
/6B2ipqj7T6O+wqT3oZB15uQu3PNTdHiulfRSNEbvsxQL8t9EvUIW7FLwkQtl9ylWp0u4hmNJ9NH
mPGvuRkdtKrdp2R/Gzbnuhvixx68MRfFkBmDwcmeBYWVC3Ukfbbg51z16vq/ihlCng8etrSeqd+Y
CqCPmGTnlTOJ85iRXccvyQLKaC6YS1S19fbJMmPpf+yI1wSVHYjQJKtpbcL34tJyVGzlDXwUY3Xc
RtKR6q7Pmsea2BIBb7A+31j8RoxD991/cMGpISbNUg4k+sPzd2zRylZKTd4imhjlE7gryM0oGaS6
A1b6cvha4oHBY9TcGfM6PpkCiyBXg5WmsgJ7WhJIRlt+z+heFv0Kzgi2T0WIOnhPt0mrMcTuamBa
3TAx4Z9XA6dFpAyAThDWzHfQyC6fpanvVmf+/0gXx7VDZ/OGiz+9t9yaCuzIMY802gVw2/JeW+V3
QpYgP2ojI/iqhqksDUhGg97l+R+VBV6E1RTN+aJZIW69Zf/fNznht5LCluAS5RGnOKjpyp9wqpkR
D2vgbcTvuF2uYyV57ZEKqKpZZG/9vrreciwurrvvM77A6srbC/m0msyhN5Cv4IozwFlJ4//CAL0t
DGk8yqrrxqZYv2xIF7K5vYCNj1cpXg6Oe6GAyv1rmFkyzBXPzewYh2rHxX1mV1GuVsFqYBNNAwrr
c4JMOMEjm+YKUx0qO48D1sVh1IuC2sO+TMQNdHl2kje5vlfjgwHg/tcjklxEMpxAIZneRy4sIFol
VnXD7qd2GUyUrXp9//gb9RZ+fsTBnXZ64DMEiwBAkMId1xwFa2AlwOfyqkHJqLYm9d1ZqKxOJvnn
8hQyHLKsBlEEOTSnSuZPO1sBduIyFyisjgZZrBa7clYaGxQz6Ea1xatzTdHasHMvDkwyqpZR8xUs
HV5AiKsvNM62YKmZZ677ZsGZNC8u056BFIAOAl9AayXXzp1IRqEvc5/g13kpU9aveVE0uqFjvfyA
eqN9N5G0ZSHzaHVklA19c1icRapp1sPdACYrnU/eri+gjsfLVWJTqsUigTTbzU1NN3WUq0dISVCO
dTVFmwmq+QERDIMpduWOkVRkf/AYH6Gr8wYBwO0HNoOS1lWhdqUGidzO6uvd84mCdq/oCPBL8O3R
J2BpZgqE+D2X677H21yV5qeHwPbQfA+c2LVrLYKrSYEpSasOAEyHEO6hwip7LprFxmYLaIOp4w4P
qGvl+zhKYGuJq0GbH9xPT+Ntnz7IaO0uOfu2x7gVB3PT7q1Tst+geSqThVh8JiT3mn8rF+YaoS6Z
czXoQe5XeHAkLTk/cCX4DSYdl76EmW5IE6wb1cA9JzsQsrsYQFvL8iGDnXpyBIFUEM36JmtKuz1G
BVf+HHU9Q/sW3JC8KndGrCm7sWt4yV6GHUkeTZ07u3BtrdHVGfOjOcZ+88po8KXlnIVIGzOVs9+p
VszlNiJaSQtIvuWoVxYnUeouDEh6HGBnC/jSntTbdd7GObMmVGsnFsR3BSlc/J+P0dm2ECk7zMg7
4LF7IcTt1Pj30duRDGA1eqmiPrva05Cc5/SiUEEvGzij5ftypdLhQX28VjvhOJ/sS0XLuFMqsYvz
qv/NwwmT5GRYY4rI5ZrsC2kwT9Bne7kxYKUYi80D8kKPMMi09asEPGE5P5k/dKctLN5TeBS0sUL+
gRvNzwgAcfFvvJb0TQ9H3ltdz5qJ3uznBmggjcfAVeU8yH/M8SzsRzEpOuKT6q4GpY1GMMjH6AdX
P5gASgbQP1U/yLnCphnD/ZEXlbUPzmQhr2mN6Ut/MhfO+rcvuvh60Goyr818wMsOmx2ERpGvoGGM
JjOcaYWoV5mteisiSqJgGQU3pjJzjGV0XU5O6Cwg7hyhxu5CkH/JdEAIZvRFLtzl82PVIghbgHUM
LgRGs+IGWM91MUwqChQ7cRdcNCQ5RkibBIpbSSGATEHnxFYJWIo0hJ6STzHhTCXDZgzL3h+YgESg
JfSyi/v1VZI35Io6BC5sbppLJ60JNzyi6OUGXUmCWeRrrK8XEmKjQCa+A+6hpr0uf7FqNls9MvzI
QPi6gaS1DaIhBlhaufY7XhUAKf1dINTFF3mjJwDtWdrzo1IfvY5aw7KORU2pEnMpCi3lNJHFOV6x
nx173pkBycOf7wJz0j8JEdL4fT1h70MokNQaQxbt2IvP8GLBX6U9IfGKx7um37T1saw5Ctu9bH4q
h3BGFE9wujvbjc3/EFA0tE0PyJl0F9OlgbBjs0NiaPGe/qr52XEABY5fMh6cmksPC2deqL9LtBaR
tZZnTg8I374m/RE8lDEZ5L5MZRmb3TeYRAeaZNOKztObDvWhPJu97A4p3+dm+sb4rNSoWKMR4VQX
zwMsNXQkTqUJfo6glqdWMZdvzGfMEz71O4r1PCbkZCEl/oUSIyNhPAxkLaT8imXz5+pwbiZvy8YV
F9eIB2tjm19wJXEw+02g7ADNlgwkEcRvGhhVBf1f62Q34v98xyoNfrrug3565NIXgXQvqOhiEn9m
omOLwpFjqWh4KB92ztZaTqcBOn1D0lQc9uvH7osDW3/xYNg3RCxoEZlKZoT8mBSj8DyaWQ5VH6pH
7b5QJnPMsCY6S3j7nhRFJJkwVnAyEZuLfmpqBja+db7GKMyV3Z7mfCkyLg3ri9Zk/828gysNu+sm
Yzb4FYt0JwST9gMYlxcoCINhJn4OrgHQ1SODtSe3k5g1HLoO804d3X3MKQt1H+fiPE1DN/ge2NET
3e4KiJ6ppwW051GaeoS6fNRq0K8jtiXObzWVGyL3HbtbqcE029pzFi1yEaFL+hTNk92KG1ZwnY22
V2apVWVx9gVjA01myg10IJt3FPfgRwMeNwy6vaJ63GZ+E0qSYq0HgoKKP2EsGRoB/I8y1LdfJ/DC
eJKOGcehL/F9uKC0B0pThSwvHftBvspELjRBKsQmWjHLSqpX0ybqU4mEigL4UApthBm3fHhP47oU
DDCBP16p82hEgeQVljMJUdvdjn+aeikLor6aUCuYdEtA9KPpQv7RTpWuFyRlZyYbVqQUm1RoC64B
AggctCZy6n1LeBg6GQAir/8yRQyLDdCgeOrNdsNBxC0tbzw4iNWOLeyLLLHWp23M9CPUMSRIcgcx
j+B+gU5SdFQ0RLBP6m7kyScD4FJzak7CVvl7pjmJjoVAj2rHZz7vjjjoZNpTZhuVCogEeZ6uZ2rl
eN6nWCrbn464wdzIp4TvZ697aGsC8XKb4QVwJYSe+fTGUMxc0oLSH/E9G7c+aZjkxozxJw7fo904
KoBEvYrBX8BCX3CIKE2JzI9vjOQPuTIKJqZWiwsmQ/8pmlxMh7jXaH0Tj8oIEm5Th9SY3wgIhXtk
XrAlChKnVWXGXQH1RdEDFOjNEY4jA+pPgTr9mow9D2MykHIWvZYl9i6V0Mu85Qcb49nq3phtWsgP
nf8d3BpUJH+m99uHZhuCOSU/Ur8OESAOMVeQVIZRczlxLh4cyy8Ez1u3jKMduelNKhAlOytah7EP
tDn9RWDZId+uF94YrhzQ5WEAWYTnr17RW9D0wmv0FIN1JGmWfOuTY7uVtesFCpFqnA7zyYEPBjAM
KEw6CGCmRnFrLbBlRE4dcSlBIpDWvibc7UgJw1kwm7pxgjzG6jtAwjNLyUgnWQF0IewLOO+zSg/W
9t8N4b+qyj0RcqbNHk5h9M6wH3ijbCt4ZX4WM0SXFcn7SrbyNL1I5jf0sjHjCCEiapJ+iAAqAunv
zPjns4jbh10iiUpvyIixUu07ny98GNxm8Ut2vjt4Ix3KgLiWjfqsVthA1nbW8D2ikJ6PZuFi+6Ps
a2JYg8M3/18kumCZnoojzibuAuZIHfZyVztzJ4fruI+E2xk69Tngml1QA/gOOaIyNcRQD1xsBAi6
oiGbPEX2d4nnfdgBwl14pnCXYeLAbHo80x0G+DBMTwluHzp92YHUW59iEv37AUZPAh1G5ooGK1UE
WSjGN4nAfU9Cft9cZWDIMs7mISnzcJ44tNY9o232bHpHB6iJgMqi+G32+KXCLykaLPOvysXJNooh
XrHvOVeSAeU0+KiCu/j4o1lh7mfrmfazjIH3P9M1dd/LWtkF+em+5IHADOvICCniTirz6QqAlbbn
S6Rbqj7flJdPZmpYIzi2VkM/qyeg95Hfhm8luLtph2i7RMmG2NGhyoXgQkkRBzLU6zkTYzu6aaW4
hv1VxMT+rmHok4uxWdQZ2/o/2uNzTidkImUxPalZjNJHaM3OqEtFRwHMcrV88zAInjy/oOnIqP6T
/0w6BxmluyzQumt+mXKEuHMm4Vy2xeU9JGhK0lnLjPiW4S15AjHH8I3kRBin31d40VXrTa2TYDNX
BASNoupzz1uIip0gq91vvYWkgbmuk16OxVDcO//Da/4CN+UXuRUdWzycJRyBQCLeLb7elr4EPusI
PUI3dUEmWrxsRMV98D2gphdko/jF/ueyouY27XI0/NwL8xug1orwV25iPZ8oelgDuYGcJubju+M9
ZdHgt8KZYhDdRuaqg9gx8/X+Re5uB0sX8cEjB+nChe16lSrPtrtFnyEn80LygeWBqAxwZZR7Qvrj
wZKBkI1JWV4qtMgATg/qwL7k0ElgOFw3NokYd9ufiaP18vgjIVX2vqbnGfp8scq9Syk9bv6/m1rM
6cUI58xzhs6lVrKfn5MLZwQzZgeLPDz1B8vco1X1V92lLpdekiir6e35nqXHpzUVljvWbBalbMHW
ro5272qpcI0Ydycn7fX1A32kYSaevW04Nxybj5zeaDP3NNW9LTqe+NbbTVM4FdvtOsvBqBTGIZAK
ebeEBXbfwDIFnaLxc8kbdHvlN7wusQ/lWr34IsavigzWus7BLpyT5CN4B87j/eB5nMvpdEYLECIM
iI7gm4cCxEJQ6MhwmRG5D+hc53BaGF5IiyQU/TvrfBTgYPi8DWXpPADX0C/LBzIG0fevFjEx24Th
wwZjEAwvRyMrheVfpAOaT5wVYHd25uu03KPfOnI6OzyeSA/0Z5wIdwa6gk52nzlNyqwAab8Jfog2
Hkw4qXE7aNBdus7xvR0CVDY5RsOxCImB6zNKd1HWfB4qN2DcPtbMfIwQSZfBKymMi6d1Ru0kw0RL
R5G6eaZMVRWjYqc+EY53SrCD/hD0Cqx62PPQFc0ve6Tg68GKqW5c4NstTrkC/06YBWwP/OYvppka
V7gP/ysQW+BWRuAW7xGdUWgOVIxFE1VJC8fOSvVwwA5ii4uW35Qf3n4ZfXYFapWVeod8siMNZfNm
dknTx+zrsVli2WUrbvZHY/NLLohxt78NUEAEX5Rpa62jdzfc5+SEtnO+k5SFuSyEeA2cjbo3HrwT
3Mr0HYF95bqeImmgqbN1S5rcX52SrL7LsRTbt+hq98n2lVHJomTOwQnnBIa/2A+RndLZ/YZfCASp
67xkAelv/+MAI600ynXcKx7w/6OQWWHVI02PqwF8Cq+ruqST8ClDqxHazA/dP2sosC/9zHzjypKm
8oLtrS3K6cJLCGHe3LLIIk3fa9FZfPQuTzloLJ6XGVnJQptgIPzw4hcnvYc0lwUq5v72HTjvXoiD
+QL6j+8yzyAMlaZlckr313G57oLvYFCyaZFGcVnPkvizqFYzqyuL7J39Ye5/b/ALfYlnNs8Q6Pv+
TdIre4sLF4ahL0uKSlnv3BYsUZZnqi73RSuwBWAsPoGu4aahIWIm4dvRDjaDe9QuFA991U9f29br
mLv9QbwrxJ8quv3dg3XwShBEAHZI/454G/9xaz3MZf+DZP86VRGlvBqjuh7lOH9pam+zUXgqFXlT
3e5fugPxHw8UlpPjqcjrLJRpEie8zGpsktiyDUx543Xo/gmr5LhPIB6Siqf822bbkUjDQNbTFWea
7+3h60EwALXuBXBRR+4eCYfyp/aiD7NZR7uuoMk5sy+aDOfhl2hJ0gZKsq+deghgpGKU8HZeUPOt
riMB5lxufEWm2gY0+aetbuvaX/KNdj759K76BznqTJG82W9NgTtQYkm4/66hbozsBlo3xVTdQ3LE
7kpOrxcmKKwosmzrNCIjVnTzvaCPkerJmVo+kfmafPTKkadPF8q66WLbB3wKLylzYaVPnCL8rMv/
/st6dUqynsol9dMKMwEBmcD0++X+dI2K3Bwy+y+w/NgeR9kXPBUVXUQ2kwNo0EzV2VqXkaftVytZ
gQiRqdzhixJV1X/IDZmeVhPRx7MzqSH+NYeaI2jL5cGQg86TpsPpj4ONnJkp+KvoOC8pGvIXq5Zu
/MppgcCJwxYe1qSfoQXyVOdWgv+nfVOxzD4ifOvTw6ReMcXB/6Qyp7XeDJjZ60drVfgvWlCP2y+Y
v1YMlGrzZ391+4PRYtAAueZtg4/+3w83B4zVY9As+c3Ej28u3bxEOOnPR1gulJ0/MGgvkx+3+Khh
9a7jRTP/pZbyNplHGi1pUNjvK6Ip3SRqM/dyNmWJ7m7JtYZdUlWIWOqL8MqpaKgwVtV5OOzYgjcN
DbOLSBozU+jbviES2oXojydw/V2/cQ5Yc+0+6FMsKUxPrq1XEH3MkbqUr50hOup4TuPsPdkxjwh7
Dtg4gEmDDSTMtV5JWyU1ntodk95n5miXTOjqZnww/BFMMoNyn5OcBBz1/RypGxTvILG0AFakaAjD
4uyxf/GluUPtV5dsmspQpMzHWNvx0IvRHPiXSoOzhoF75fMxntgB0iVCF/r5+XGs100lMMPsyaZ1
IENAvs89msUtEME6V0tDh5r1zeAb5RLOFSHG2zBWSYTEI50a401KXU27xk467F2QAT9u/RK2+Gt+
V4LQVo0mU6V0U61wxXMBhYnyfeiA44bma776goR8QU/qmjXOSAxW7oRyAV9DuIcIOYby3VRlFcMr
syZey5ehWHYSWGxds92SqvjOh8pBxZ6uW4nJlMOHG8WsneBWUH3xza40Kuqf06fAyed3wugrETZj
DNpmIG75IJ7ODueiIzQZ4oXEhtLovO8Y8W2opJ4dkXbXtRGxZ3xDSa29kH11Ya75uvK2xcUSziqs
hKLq+DvNKMbBSlf5XGe8vmgCnZ9p0ZrNdM3NDaHjzJMzLHnhLTaTLB/SaN2JNahBI9xj2mDLS2Fb
qwwD8e3KoexZZaOJUIQEREYT8ZT5z3xGrKZZQoAYLmUGoI5k+BtIm2thcEm0MUhCPYFZ0GHLK1QX
4932kJDgcuJd2jbT62JGkAyM3KvuI1z3dQtKImfNZ9T35uCbC2xeeFQ61nCp2f6FVjq24A9ryYsB
W3VHNjthNWpB4dfrTT0Xxd+DSlYxBK84Vj7GskInJC8wXzFF+Uyj5ojM1Bq5q0Mlmd1kzh8LDYcP
UwOJRMHuUEU0W7RspJ+PynH8sDhxknjcJszQvIt/JwN9bJUnentsaZjbQsHtgGmU29YgWjQo37jt
wyDIQtYZPi04OQBAU0PQ8eWXAfK1HwBaVS9H8rgK9M4FbxqgWgVW6xWPeFoXnXehaHs6yeiI4Fo7
6MjGeSbzoIZZ0WzvqNBwHFAuUkrg+l01MH/U/X4v0mfWwonnxk3bkweiaHEOG/2NszLzC/drbHxc
d7qkfhjyzQ+F1spBt2ThyG+wcBDDSznrj6AV/EoIYKJFAYBxIsYXaIvJxEpqPiAURD2nXSzM61nL
YrPLk2KWiUTH5W8ZETaxnVlVOnEGbKm6c6hX+izEBbxXkoGP//h0jyBerHS+GOVC8C4tWVT+SLkL
ZwxQFS1kcMnyo+U8/izlyBDl57l6gP1kcE87FvvGZ6v2ZTY6FgIdGPThtLAnCsLa6qUG0L6jP/h5
9ciTgnWW4PUgExJ8NXN/afD9tvGntzXtTjAglA0vBtigfw6fIhp/jcm8+LdZC1q3Ux4/imnz+/Ye
MtDkd7vlymdA9Gz9pddhHmuyQOZeWQkZDnSFs6q0She9x00G8XEQT/5utuTC7Yewkbvh90tbKg5h
JHyjwwjQNZC1insTitWdrYA0if/HMZ9vAJExAHrWAkSu4gQEExg6HS/bGuJCIIud4OJJGPzUFaUE
oyikiePGsiXJt4QA9TFB7pOtZn4cvBw+49yH5OytFQ/11yKqDi1sihFV3UWnxKH63uPubG+Tz+4e
cfNNsg7IlqEJNEevm+o72CJRGM6tuVm7oxo3uXp+x2xixffDCrpmX/jfNeUiCu84hNgVeEoPfc6v
lyHhydBT13jEAGfbPQF4p8e9dWy1rFMaW7+dywkHeHGctQzU4Krylb5cd6F9Lum2GLtlfxEGByQT
MlFNZ9fJk+ECEEyPdFagFKwhFrrR2BZeBiWJGOSDLA2f+d2+trnXwPSIWN/GlZWnTmquPXoPUdVZ
uSTM7W0kSu/6TuxH431ot8MRlPQbDmbf23+mW1AR40hrC3rudmxi5qhabwQYgEuL07TkCED5p+qK
GeOur8tdeAYRnzQ/FwIRpqfVqEslZRKr0+G5MFDst12y29ACZ9SrDq4TTTt4TAOGhxAAwfqRXVx2
BKj+0ifOsE5eCcs4eT5THFSrAYGUQliAYf3VMCh+fv1HipYEqBsLTz6FxL4LwPXD8fwRiGgTzLlQ
q1xeE30BCX/mii7azoQhKZZoC0GW1ec3zlXulGoZ+ujJ1YqIpaAoI610QWbE3JmWP7eT+d+7QM9W
fT3JC0z3vu/7qbTMcplabCMwVjLtXD+A9aUT3tsDZMGh5IMmocRt7OMTchKFYqol44thDjM5NfAc
+bFQNiRmUCk4dcUPBb5X034+I5YZ/6ctYePQjZlLyw267E0MfD5lS+ufTrOz9sfp4fVIYEYQKxzx
PLaOrcLRm3//pxJCn8TyTfPj2pEAm3XE6XQY/Kd4y/Fi/f4JvMrXFVKqKme2mX/ck8FbnEFvHqT3
sHsQMfudD8DcDuey4l7NiiNLDIULSRhLKZSYIUzPoaiEnaySwVPPgoUea3sNn6l+c4g1BsLCg5Sv
1ls38mZ7jgWSSIAJS6jJFKhaDYo5Vq5mDg8onUi3CELdKGPKdvphafiBAlwH50R/ezQmCriDcljZ
EJ5hlTzLEZH3ns9yL4FQlWaeXq5IEXHdis98H8pDP++4VqddrhNgjqpLpXxLfA885tqnF6ed2zv1
TQiuiV1gZP0cHWvmYxiwmGItKx2GY96MG7Wwos74l5VDrEMArXebHa56WnkMDuweHGW+Tk5tJkXz
H2yNDLVqLuzaxfBNVFehEMo55iRUAb34GUiF3dDJWgEBnOqBrDUdmmv4XtH8oiAn2KHDm4jKE33M
JpXPIvVwgOTRXTL/mO8nbKzkBPskdGbtdsaWTIY9GUgRouxB2m7sbRIFz2/wRWCk+Bs7WKabW+CE
g1m0fx3mUq98xlrzV5ZZZ0cMJbDhUdDRIp+bkMBBXG2iTp4/G8btnPhZ/fjKXKNR1dQXxEy77GBt
PwQyXw+xMhPL/44LZfEky8vt91E133e93+ATdfMn0uUQEFakE9DPOKqRYNHGw0GEThZUDC/BFYIk
K5zmFjBYY3tfcZT1PCXeD2OSKCx2c+TN9r05PTHBQMpUrEULWSHiIKumrSfmqtWFEuOKe2vGa+Um
Sr7D1knDMEp98rishEYawJxEIbUtK29u4EgDYOc4ozNrWBV01a7zMUp9PMiKg9TXNAsk0PSMa3vh
gh4x18ln4L6aq4rua8QbCY/IDPePguE1+wV6M3/v5srg/rVMYfpq8T6ScyXebK/+U59CaY1A7l09
+ngnNrYmEl55QWzmJ5IcuJYdWb/1jGA6GzbeGw+sRtM7OFTfBI15aD54cFkZlJ+KvcaZLA6S9v2p
sMOD+BdxkEy4e7vcz3UZDwCyu/N426fNmdju0llTVHwDozBIUrJ2JfJd/svZ9HoNeT9M0FM+BC11
25kZwqIGPbcO4pBTzjyzYd+MXzojs5YNMbhhpxk+s6/XIRHnVhjuobYvfos2y46IC9z9in8EnQmj
oI++fr9d8KD6se5/RgBRHFUT374gqAp+DCUZHCliban7OXIBICibMzTjnPS2dgWSrtg1ua5z+d+W
mov0yYd4L28T0AB6lA4OW0isNg1tT5Tx02k+9ysEW/NZTxi9Vx3xFwDuS+eOw5Mnr7yCH+PKLO8h
kNcZzdetPrY2J5izSCNSa1Sd07sboJ7cwjDLBjFze1fIMBCu8nDp3wkDt3gczzZ9RAmmU1imqqe5
7upm4f+pnCKY0Cjm1VZ0xe0mwLacd1qYSvggb+5ZjGkaFFh8Sp9/wJo3Hw3O/qyRfJGoUuyB44xN
Gfy89blEMxxxvCHazsbmknLeEz1Q5TfgtP3knkBclmbTKH7MugAOlXn+/5QAMsfHjZxXhgaPuFnW
gnFSGQkmgGvxBBgeeYj+NaK+LRKEeAtPuXZYA/0IorspcUgPBXCgZb8pCzLKqXn3GfQn4qZap9QC
iI3+rIiIH5iZfOeG5BQqcxmbMbLtcfzpLHdW6YLqlk+/olGupZcOy3UuIDI6ltZRdMukv0dqn46Y
QtnWcyvgKgVbwLj68+skwsDEHCdU9CBAk23rD087S2TZ/Lfw6wCGJsNpJlbOyo5dcDWuwYLOElmi
oedOjJB9najPAQLPZRIJP7lcr54yxJYcAfSeSlrbw4EAS6mcye/ctq1teZ2e+DDXihJbuN+9TE5Y
oRYN4LIPHzpvwAM4Tgci8uyT2sAlGluODJk11VX2q76SQqKEgML6W4ptesNc/593w9b/OEUVgm9d
SXYDz2XgHq/Vw7hM14VmclZ/8MpXOdOfkYLfI1/w5IvIGCXuQnLgpBPVPGsphpf10kK9jmmzS3Qi
ShRXbgrT4KQfjnKNtynV4yAEO2djc98hQtKUumXJ3oQhoRdX0V+OqhZzLssNtxH6igC243gDLgCS
42OSyUgsfZzmIbMtBuMAZaq+LvoP+OLMYpDYvZuSAUbEfGgXUdY8fxDL47+QO+aBEeKgloXC1qgI
thX2Khmb1BJyluu2tvpqxTYkN12Rc4RZ5lLQJQUqsMh9w+oFkSVzZuEP1EWDsoxTyGjbqeQ7ibeq
FIAwyWKb3i8QwmU11+b8bEAdzlfUX2ALT+OWBgyB3GhtBLDamkfoCQdcSoqIdbEmvAMycJPrJEwi
pHb5ri5ayYNi8Vto0ZwTOqnT5jejziQIGM23cXOgpWnWnTdpgVBc3Zf/jUy0qgTEZNHou9YpVEs9
3Cg3lymqBiyoLHtDnFamSQAPvBKO5J5jnDxMghK30B3yrs5T/iN0PJMjGxY276Y8jEGgGk235Rwp
Tb9A4ZoILLzOSzCIu/KZhhiHw0C2ijx2IYw8+mvZG7DKhFtDrMtdNIkyPTPL1jm0Gk/EwGBK4H0B
PrIvn8CYYxjtAPyGL6JDaLpZtNCjWsJB8ckbMe3b56y0+mSG/SNRTcZsPjXZeVG3mK/wukEON5po
d/0jA/vu0is8G/KcJSb6sp6MtZM9iLyibYcjOj/5Dcf6lV5nrOUJXknQbJZdXtCXAbAQekGwTvRQ
M40rPGoH1TT44Cmy0rtPbjzE77hCrziEjD1sOj2IXDxx7XH9P8ciNdoiOKkCh5GLB+uQ8/AqGR5r
EUvLUcU475Hpl5IFjRHAam1Mp6cmzGEoX7iKcEys8KpYP+ZJEIl9onkRyroQRJ/B5oogW/yNMQNO
0Ukd63Z9makVS7kViYSbpFgY+33SiPoo4zyte6V1E7A82+01SHI3nBGg549pJOjrFB8Ww0lHXtzY
l2ZIPDwJa5qDpkfPkyv1G5ry4dsOmNOS4e8eobMO7NPefN318HW/bG/jUSxhj8nanWEOAqDFmvRV
pZFg916o8Iv+gj3OI0+4j4UQMd7q6LZRJtMwZF4Ts+qxI2HNJwqXhtPSf4rRzydBrzRXI56e14MK
lngpNeO4GYoVHHAH3mmfuSZV2Ut0x0jO9o7jtS/D+KLi2934wWgDNHqs8lXRO3XnBas444s1SNZz
/TAYcg4yB8YW08VeenR8xTh8LZlmCv38oErp1F2dB6mOawWflirSKa5bZ+vaKJmjpMM9fB2ooVyz
NnvkxJbF+lMpTR9Lv+NgP0O8SAeHYab4orH/yXrU5Ws/1Unoom4X3hLiZSkn2k2ZwMrMcwNXDkLi
Ckzru8ZAOFVSyiKHHhri3J+ZdI7twgDQSrw+Kf9i3FkJXa2B90EbJQL6TiR75AKFNmNzUcypxpsQ
poX7NLDTw9G7Jm3zIlYIpZjPDDY14EgWeNNjhHk4GSS/fFxu1W9FeiTn9HcktlEm5mQyz08ex0Kf
/FdGzw5/idztVnafBWiWgyOeUxeBXqFm+i2OQnQQt9jn8iAxBl8O+wkvWUXBVR6eo/ln7JrJe18j
u3LId6IE47PGEBXqHkL+FMGW15r8lwsIz3pwBofGXUdBvLT4F0w91Gmkp1wSukgCyO6XZMi7Ta08
ClP+fIL/df7SMgJv+76mRrI3WvRAnys/YAny2ejE+BZKnDb5ARpvti1YMn93DfuJAb98hUeaaIb6
usrwuecFuLMGCuDRGi9xy6qRSapTuBsHZgpPVwx6AZHPkH8OzfiolDRDSaIy9Bzs2ViU56IbQjjo
KhbWv49dYOF9KwBHVi3az88FT7S3F5W07OF+SmC32lt+wAD/KgBJXTML9CHgQqYhd9c2OGbA1VRb
QjirFhuGwWHsazquTBxr7Y1ZwsjhWqTv6du2DBXgBIgNEJGiaIhQuK9aw/x70lu7f2HzAavVVsI9
s8DjMIU7NQrydS2xXwlv3YHygz/52GPTebb1NoCoX+8HZi4XNaVY0M6JgTcUbMoCvw1/4IqM9fAu
p8f4dlVJIZAPFB75i6e+2sr//71dI0ssr58UhrRqfkNohEaz6eia4EGOAearImvOl6oeQmUWP8Bx
Ldb4OlqBXOqbY+oYTqKyOgOpKua7Zk3bapPlolTcsOI2BoI4GDFdlZaH66CR9n+K/kLHHvo6X67Y
l+q7tD/cRcHgOLMB88VEQtR2gTQvvXqK5z1eOm4EC2XrAi6elahgHQbQ+gSE+ouVGtQoO1fCkjLG
BnWZsSSccZg5h9C2F83Uu3d2zoO/JcfxeMfOGGlBbhEp86io3Cw5WA9zfXrf/yqz1ZDP/W0Q+cjF
NyfB5y+zMamqNLumIY7VeVNE5L0Zjcda0bF6YK1zFqw5wjWUg8g5UXnsxIKir5no2geVh6L8Delv
S52ZZsXFWdNIuRit6I4xfBxjrxgt9JqQcZkeDGKQOhEc6XEFW3qurVjd38EK2gs+QQLeWpIsPUnZ
WMGQVLWn5pTxmzOI8WdAkFIE52qagRJaL8omqqy3YmlPuOUcy7doXg7vKuA63ferh/+BB9rqoKme
BRl70q5e5f7AuVO6jbzW2bQA/918S1iUS3aoBW1Np4Yx1CrAYy1CS3W2UetO/eHw2qY3ypJyL8JP
KJfmeXNlAJwbAFQ6szZbEyLuq/kFaFQ/is+yiHRW3Bw97+mAhuclTxClTwtRBEUCgVAC0Tsry1Ra
rZfNcJaFS2lp0ImyXvrX4f1Auv4KBSHl+nO/CSdkZaPJvAc1c1y4CANWE9QeOpdxO15BHJj/yQGI
tTCs0LWEa3r2K8aT8DwoNUZhf02M7n4mcZp0nuS81ZObIQTqB7rQswxDmEyfw3Bh/D9ZUaWGDfmT
4T/oXPvJW1M1360TTJ76AirrwxX9LxHNNzbimWMZZ/BzLUNk/AEPW7ipPokuVomTwUyDa23jgYxy
1NnaviJ0cUufHn3h/jquEwqjPfxZTVNlgPwyZDTHrLmIPWkcdE/OnenR2w/c0nSXV3jCgiZiYgpY
ZnzHPw54NaWfCGrBeAh61yiET6W/4uU5tn9Lj5bBjmSvgxEZa5VuIJtonrurtWlhVKp1en71+aDw
s9DN8M2aywklz0KAnQRkh9IZtUcI6ednccMQDtlEpE3JN4KrB6xalkVABvm6imrV2K4EosSvubiB
HG9mnrORwEMD16lGfbr2DUyRrrYeyzE/mdSzyI+2VFUalpw6Mq6YHAFQsasJCJjFSjvLqAu0lKfp
UduGkIpS4HilbHffrj994Y90XpvLIAu/Do0mCeK/M0aHMKlijWFY5XRinhqi8Eobq64aJvMn0KzS
3WtlhPC89aKtB7BUTg1YHUgTfDUfaz6jYzN7nBSz1j/aWnlWRIB78uti1jjgjb2I2O/ih/S1yRfS
h8VWBMMGb/WHUbI9Yck3b163pwKXfsbQcOmVA2R434luaoPj2/U6ZtoJfIz7SmtUlRq8Fz9GI3QP
69rD+xOn6AchCsGgEWd06gLBVeap9voh48reut7hgXUY9NVmCNcng4akEC/WH/H6UPZismUYG4yc
IV3jyhx9RaUEof/KzbBIb+qzWyNQyrQvxouuZWWeUZfVr8J/JDvYRzjdA9ib6ZwOh0dpcU7JaZj1
wr8r5Gazl81Rnjb67G837j72S/4Wal4qHEbHWDAQ6uxloIMTp2jIZxSoiqCgPVF1EDxlt0C7GNU8
Hv7WdK1NAp6aj1ttmW66/EP1TXGGOA083pIlNYUnWNtSHdNig/wAbJF8QnD9hoyfZT2UkqkqGgoL
/4upU2K2sc6PIfixKu1NwZBLZVjmecqxYDw3p5C5CHOo5J6BoKpFnpYIqKwyK9xOoT61m72tDxa3
Io+GGdexybWNdHsW9aQXGLbQtxOdCq/cfpLqAE+tWvMwo9+oL4Zo311EGQXF+pcQ+IJVOkWxSZiZ
2lluEREdKRhMDN5rnVPUFaKAKjENEDarDIFu3Wn5kwUD5rqS+PX7neenWWbnMVlCX1Sr50kxrxDU
vpXn8mdpWMgRdPjokNIPRcdlmaPNlnoVPtHJFg9ed3sxclgnUasqbPl3VAQg/8zgsU/V1hqUuEB9
9NdDqUqQbmmuJIO8JoB2afKz4hZ7exRv1QTh9krvyZnEkg3yyZ+g3DRMOxOSqvjMws+aru1au5Ur
sxCvRHpQEjWxpVjRuUBIaBXog7LmYxUl5EvJzyeJuzWZLdJofYEssw5FiHevBe9vFAFmMQI4/CTR
ZN2pjruByksw2zXX/2EzvAuOgAB/W1Sh4aHpRiWKxbAZgekKNudqTADoODBKDPQq8LWMPaaZkGIu
790e8AmyvFLi8+jC0PI+ZMmJ2IBHF9+ghr7VnmeMmwTTU5qLXLGJJ2KBckLNXO3gn3L1ZWWmsNmm
cyKlPfeLdveEQW9/c6NSoBkophQ+MCSfNjxjlRUQMB6ffoy+aj0x51IXBwKVRtwYuCVdJ+76r5vF
rebEG6Am+vJspOhnzBfYVWj972f+8EAFR7E+QRkZ2cvStvnaKvHtqcXnkXEgmxVf8sYbFoA8oW/b
srTX4IBEeBWBjB96fOAAxkRGQm1atjQ5l27JF0XTguqhR8O2vdwBPwuqukjUUcAGpfP0Pb87ByT/
v9X4JoFdXJceC9gJAGgVs+Lc1syzjlKxtB0vKxQDANMFAaVIK105Slgwlugt/wfYwGhO+aYsI879
jsfB9fG3O51i2ggLvGiQgbH+ccU+CPrEB0Pw1R3P2r433iFL8r7CDtwge88lm6cv4Hevo17SrgN7
xrbegRyfu+TKZYVkvkikH3o9mVvDLsXYhRcZzzkaNrrXEeRFACMPekAXYK6J1IPx6aEoJvbr7Q+a
r3sb9+4Cve2veqF1vFBQtH+bwExmR9WXyiIDrArmLQRXSFp7g4mCwfXhalEFeMDXqf32Fs0SJLL4
v4mM4GuI61l8bkgpCeuY7eYIxAfaAAplNyWRVzwefC/XavVPSqzfeCEqxnsb7PHZSr+UDQ65p8j5
fVFF1eVzLNS2YBlZhM+vDqOW41OE00MBF+57eDm3OKSqnWqwhULdf9I9XgGl1d9/J40lQImsf6NC
FZm7aSKs2aX+fY4uA7hhnbZKov2lPCo7LKdjH0sMEShd2DMCBO7FH5dV2gaLXMQpVbi527CEp1bt
VGjeS+v/dafo4fQzPjai7h/LH9mWjT6/c3+NNu9tMEX21XIhEdRLEFP7ry6ww8Nk0mkhIL8mcYCc
BMM/ECkDv0ssVIhN3yMHbDH0rj6P7+OT6yiYmQCBRpk/F2g6MMIeIK6w/mwgXkJKVApn1wdm6Ng5
zJg7wp6D7K/EP9YRgAEiLxsfiSTSm0Zmr3CKpF+3w+7LSMNO5yBBHdBlv1NrPu+PbxpanU3kPOgF
EIOz6lI7BABBuCpmekft96pZXgzifZWUUyzgQ0RHotAuUnzw/qMfVdjtk0oxBKbZPFLDIm8AnWES
rQ8WZhZKiD60vtUgQu+EMWwock9mH0Xu/vRxGuwb+M305KCQfG4TJ5gzf8/9iqu9STVrY9nhf7zs
apculL3rX/p4MXuQ30XX40ZtoBplgyr/01MhvWPkURT4ICOpxJZqgMpXUt2nAKcwUYLcXO3HGZDM
QaIysydERSOOCUNQ6WH/MokwZXToS4awp7F0ZhGWIvRkWHPowOT6wvv9L2/rgjkv04lmVNMr2hkn
GPVk/wEdcPdiaYkZgnlW5PbAG7feyCNx+c9yKQCHVbVvqRc3VjpUY7DDGJ774zBud1hpzzB3sNB1
k2kpi6g+c5nEtPkFiNifapMLSFE7RRhofh+B2lU3vGF29iMFjjJphRSGvaiECtC8WqG9TCF0hkSR
kTu/UwNDJZrGUufnRWQQ3nDRNQcOQTYfCsIZqpIb+yUfYAnSPZhW2Y44lGNYNhLk2/Z1HaEh+uVM
Q/0JrVgC19dvL49KaF5YcJra8Fya7MwRkj0GrHZphAUeK40IKc0j/Ly0BYfXya2NFazfqVEe7hYW
dpSMzCuUy3X0QMg2T/TWeFxVa6m1H0RubBZvWVv4daElUn7l2xsKPbujima+MtqGTBtNZ7Xf6CMF
PEo7WgEEK0ctHR7t47yTP/VjSFK8Mlv8epAF5RKAUPWnS4+wlIzpz3XBZcJUFT6DcoDXMkx57cF6
aInOtU2dWaWTznOl/GvtirJmUvA1mTXtS0nvRHF6ArcrnXV+XWxusYHbify/efMVFMsbwIa2KP+E
MW+YZdzq9Y20ENMjHPb+yQQZcXCxgyzL/SvWxOdc7u0glseg1K/WauKCZLU8xH2UO20BeZy+gQCe
WiUAl2ZbVUEgaJiiQ39tKmojZJ1tzlEqjVxVPxj4XmENw5p2ESvm3mBH2czIdi45uf/jGirZEsim
TVGy/fzlwC+lwqaL887cSDSTQKr4eZIpCS9DHPELPzFalJ4ZBWpKUlo85TSPLGJESH0D4THWrIkj
k1ppUJEj15e7ZP2NhbA6gDBzKdJ3vUb+D4tDSNwPC1OYb3fp/RcK9LVG7wsg4fZIiYJhc6bRfiik
SKSSPXn1EWrfChj4MZPI/7tAMdrWQb/ZVGf5ud/55O9IJUudDc0w5s20CfPboT1xiHTXEjow0iMR
e/iaY/pa7+Sh83UAHaKZ+WjFPKRrSZuZ0Jcsw6p/oIe7n3KMhhl8PkPRMJLjahSwzr9/98VuwK7o
KWo6Qg8vgT+ZIyJq9L9ONbqNGwa/rHaePePeLNptcahNcndzggZHWo59VAsCKgkxDo/zI3dDp049
y9kqOTCr3aRJ1AwKaeCfcVzEHp6fLZPA7aeADBvJu2QrHFVujwUhjas6fRgT0rlHfXstnb3pLCyn
2JzhGwTqB/BnW/PLauG9NSVXQVs4/r2BnmyhA5AiqpDaZlKgBDXI2TABwY2/RX/erVU/hHkKUdmH
UlmimEIsYGBBkEKBwlMu8eiyoTHkwF6Z4eEmxIQLSCfBoLRIMjwtzVrtN3C+SgwYeXNEe1CaQini
5GOn/7Nj2CgnQ1TigwB5JMpkCQpQhtLoTWEyxdIgLrNSu1Gyp28Opu9H7hfkQ7RZHIt3l2qWHfPo
Zrf1EcpMOMDHddn0FSYskdWgxPgomkqcAMMx/sG2z2DB1jzZBKtOiUCUJOQIj+ZPSUGM/r6jG0/H
B9UtwVLfuNu43N00NBIV/YXd9uvDzCTH4Yoy8a15Ev5zKN3pmq95yutpo3AWhZvMKI2mZDKm8Y7b
y/Ngg7EsGqvMgyyPA+SbQHIlQXAXeg78zqxpSsUB0E6OFxYmbHPNb1EYwh5QIp+l1sTUP1mOA51Z
dH6RcYw82pmU2qPoI0lflQqSCGSohTz4YvnGZPTy1hSrwDNh4DgnmDtGZnABOKgFMKgIFIRYccGg
g2R79jvCm6aSpCFbLNp4QD42Cw7bxwG5vx9ojIfU8JcRAXxYk8A2+/++uxqhTJL/HQT3ANOF0q2k
zQl+TEO9aTFj45qjf2CDOxczYH3oj2AGfDKtyVu6O59Krowv+kw0v7aM4V8/Xm9wT4QQFsQhe7MC
cJdmpBFzxQS3DtAPFn7yBTn/xwXwTWHT/oEJr5b8KTft2SKfVpBoXBd1aFoAmDyA/1QUZl5+DPSS
ebc9qXwQfccl7eloifKwVvEShmK5W6l7ejr4P6yTg/ZSpU/nudFuCw418St4QFWp2W3BPZ+s2TRw
oHHy4wcDOjeJ6hs/iv0YrfvO7n8QaOJIBbgWyB0hd7ptqSzxcqL+H9cORo+efEdcyrItj83iFJkY
7O5cJDgMM3AUITCpg0CnTrR8x3YCEC31ajpLfyOPR7nZLMw5ldiLtVHmxw47nhXIcU7QTpRo7Lmt
ZEiHrZYOxd1X27TbuITteECunQw3+d1woDtkooOXJC+Y8nhAIQcyS5MIEps0FMGuSYNWCIW/Cnt+
M7R/o/rhP1VGdV0ZXS6CKe1zRVYEMfAlgo5AKbH7Tw2mqpA60UT2hvf1zyWXPGG2qzmXqSoNzRSH
qCaPY7SNVi2FO5SKm/WCLh1dcMMnOpI2j4nbfD97tnu5dZjruJC+IJ0xGtuUFNTpI2RQwNRwsNNM
9KR5CQ2bstXReA/Qjq9BKeWpTe6gBplETzpWg3LGZbazUAMzYBmek8XL/ueOB87/g0T4oeZEu1Dz
GW03YR39FaFmvsG/9EsN9NbkETnGUEhsEW6h19FQRmwJtki4xnIB5XlADrVRyrN7xSTlpCtbHDq1
RSHqosBCxV4AOGOzYeTL4xsyYR19Tj9Aq+o5cdrFNwbp3pI4U+WM2BubNGDE1Hf/uEe2mNoHEmow
LePLxMZRV2tJt13oK5TVANFTLWRL8yh0ooOjyIdOdbbg67BRMz+OZ8QkMl+VusxTe5P5Gyn3tWWU
tzN///HoEcUrAtKfUMMH9EkqSz6AJcdrQ1zYzfomXRqWG6F/zgfCr1xRXkR5YDkAXOcVYfba9Zp8
6cNUQTD8O8JRsrltwY250rVBmrxjoTBEdnpPPvZBHtoT5Ws5wsDG13OfSP51Z2pkPcf/RyEJZARe
p7wL/97UHRFg2N8Vt2pw9qtMrsZicpUGdr9FuUSEP4ugth0lTTucuP90Zpn5YjZ6M/QiymYlYqwV
4rJQA1HQ6TqecrFHDWjW21wUdUeZxD0I7iAH5JbjNW0hNFxRnOXf1sQod6IKsdBXBf886wWdxQvk
yzc0gZPHTG6spPuZApC9kN0vhDljbrqF9gtRYNh6082Oowd96nII5HT9hDz2zHv56Gqanz6dfGlC
/ruIWMVX1RB3hkvQn4PAR6dBqVREQwQbPsIpkRsWREre1bbUEjzhcDbfqeUkWAzltSe9zbfjH0sk
YyZNRbdaEQW4+czYbepreeMMZ+23u60F8YOXKzb3NSDqj9k1KihyB4to6s6jmcVRcStEtmELO/Bn
S1jIUkEhTFvwW6wxds1gUAQEZyNNrw5Hf7iXYlvQjVxloQPl++QVLsdAnAafw1b+XU/Li368A98Z
LSK0RCcMLv6tv65JKW7lZP61Uo1h2/YmIX09vm4t8LsHdxUiey2qf7DbtqajOv1r+9EXbXepi81U
Z9E5gZlka0MddBtMefGsF/Udvn1mVXPe7F1UMLAhNPfJOHG6Ax/cHkpWSlkcqYtNfPWQDULi41QF
yEIjwSj+WNUc5W2TLirhQ/ng4Qq/STCqKpiBJ1lhDnKqjoB021RrhcId5956BCOLYlmHANnLMfck
Cz2V3C2wCaQb0eV4qdnH/Dd9HgKZb+Ot+yMBRl+lutQuEABr4kV5VQYX8f3VjKt2VVKGQa15EFAS
Kt/ecKXt7AZ3H4jWVxlMMgn+vAhYBdmnFM/ztgBLcXfqjJcdTIxLgHg2Av4gUJvvvmyMaUnlMNfV
hW695EuTqZXhkh5Etx9jt2Ymx5db/+DY/MM9oHnLLRKDJzZf6QDjnbrJn/VgXxszWJj8GqJ3XYK/
BZLzgEWAv6MmxYu6sEKOZjuF5Oi/bKGK6CNVcELOdp4+InoOwLdfRaPymz1hts76PPh4arrIgW0t
7ONJi5WmxVell2XiG+9ZHToOhtkoQE+Pf/pW12IY1shiDtyarpoNepPcuxWcwmroqvF5AHjb70A8
WpGEwRioC4V7QP8SjrTAL8f9l/k0jy5YEObAux0kGy2bMNtyvfkQioqywLpoSPw8YOtsdmx45ypL
AeVOoc2OhP3rEsSqKoq1jhd4H0lzrrCbiSxmXHy/GgRSQxrUFg2DDbGIdtuGuMy/UKQK0hjoGB7p
cUV1bdA1on5RClroO9q08ZScdz4KZK7zBfxiYDZ88cPJDSDLA46jBFkviS1cfGe3qvNV9ut+E971
R4w4YN0KuMCvYzZWoYhhjBw7ZaC3mozw5MONUXaU672IXVW2q8Zvt49YXRfEJA6mEFgJpKdM9Z4L
OY13usAp7jFAHbg71Pi/V3ZF/Enem3Rwo80PP+nKZaGdjZ3qWG248gt8AAJvjEjf4dmoMfs6Z2vQ
+CYxeip2leOMn/un8lCpizWZqFHrFm/bRrJrMPJRkD7wcMmZsIBQsgTX6TYuvAvXucgSc4syK8qs
1mqcVc+5vKbJtsmRulfkooq/rgo+6Pne/iOWAdIauJk8V+yBxDR6hwZ3CoXeRYtlCwPh1KFPUjDM
XDWaISAfZpNkql2nNCZrXjs4Qx18FXSMD1BuwGiWZWq0IxJgbG6UZfgfv0Tg4B2jU7Tw23qQ3AtB
1ZP+xRZrXA4I/ZphUVd0xeHMtVsK2EuyN6NLn0mPMkyomtL6Rp4bvYDJZyHyAA+H5ZzM5ldmXhMS
IRARgTJtqxtg+utTfnTvIgKrPAwEtlAQmQLqyZTTdxfjdUeSbA8j68Hu4xyK2Ap8akxYYAcQWfuR
hsmWtuPBQYb9C+pERsxFwVQ//dbBqmRJK/sdBk8vRkxyyWn63lYw9AuRR/CuRinogglCNfye9gU/
itPNvQlcQNx2K3D3CoYsDC74lTXtZ9sXhqSiV+UxvE8qQFVlZn1waNwB0imoto7gt/Abcn3O/hc7
faLw4i5/1sv8zb4joF3C1ztlOv9weppxKZPzSoWSCjFs+iQyuGbaEKx5T/0ePpekAERW+LcI/Ngi
smvNBiY8MuWH6Pu+rYWfRbHr33O7H2JmcIaqsftUo7ze2Pi3I7PfLuYH90NVOE8/QwbnaVDVP+Sl
gWWT9hjP7XaaO2R+3XLNATtduuMB2Zxr6D2lnwvwhK+JyebWTZYqRC7q9958FMEKBKh11FTiDzja
DQ2Q++2ROj2F9CAgKGmHKYFOKY6JPdle6OR/q0390ZSgiinIrDdph2/KNB2Z2k9VShVcW0cFBpj+
/lOVPMY+saE+p3XZiU6CMNMdYX4DSPWvmIBCbEuILNebokdxKDktiSWgDNATpZBT+UN3EsN+q1SV
Pp7tbbLZpxY8Kea9qDgUi0fUypv59lvoeExNdg87S8fLwqzX3wbquIPMV8b/c2Oujs9wY5gqRTpW
77F5AuZJT7kj3+UNsPfln4Ex4ljHfguXjjn7c+6OiJJNAZ/gfWNgMn5lOtEtblbZg7BkuS1u/NJo
cgZmJRJX0K4g4qFWNBjmhfczFDin/+ffUQDRSB9o7rZNG7s6iD2aX/PmoPwhx7IhOaamX1YgEinQ
zouQmu6pAxkGnrHQoxzHUkZ86KsO7IdiyWdoW2ucm8lPPJT7j+Rc7Xwktmh/GNUCmPLrrWOyhIUi
4KSuZw305wBZDaHKuch26bWZpwRIBLFE1m7RkJhJRtMPe9vgAjmWTBJJ14mAtO2WLSscvgnn6nBu
3gbtX34cVzrdn7ZgvISUF4B6wruuS0hmquMueiZcWrr2xOU6bgAeguzZY9JxyCTx0hS2po86pMOT
LwR0w4takzDL+DMJvKTR4UQC/g+7UdOeUH0LJ4HYTue6Akb4IzEvslLxLuGW21ypPlSdw24SCxsg
Gr0uqLYPeIEQpf6UfSpiLR4xmGgwm26YuQVDgGDZH4XbWEtJyEQcpKwzHTuZMChvczDyS8vY/Nys
6vcYVBFgnCaZoK+4QSCENjIqNK/2ov2CAnySZzLttkaf/sgFVoiCDETN4eWnvaEllWVwkXd9gOm6
GDE3uoXUvl2nAF9ovw94urHHzW/1VeB/GFE/3a5ta0g6lrEBf0sqnGNicnygK0SfKAjdrn8XFWtA
tgxgfa4KTPWTxKSKNuNLwkgx3ax9HCvRJlmm4OQOBtpm2aQlrKWbzYtxlc3JRx7fegylhPiGcXCl
Xuy1krJY/FZIgLoepYf+FCtFBMC24lCmHbVNsQcQkLLSNQmthtxHSCI682QgVUy/WAANoZCG0LMt
j75sqC2tzmeloX+nf75DQ5vrnurfGw5Ky+lFsg19KPJXCJBnOvhpu9fqW7Uyi0wC3X+o6Uk1kTLt
fwZ09IqyDRAc+mSEG2MMWgHLdbwu34fTsAX0DswX6vMVHx7MPsqatCkAGQ+td3d/jd43W9LejTOt
GjXmJCUa8IfzLewPyej2ZMCfoCpNdmMTK85j32kathpsy6Aw7ghSz1tgvyVj4TQPmqEHJe6ctD3i
PW7mQ78IuQlD9CzFWPXKXpHtPE0/flnagpxJYIUw2qUdmZSMc2QSl6uhpK2rrhG3vnFqakiL97Ba
OmnIZPRvwtenRSVGjtF6R0b5geWyuHrvx2zHXpVK8/ejPMNOMU+jsVpMh1BQYbHGNYBUjK0OqdFD
kaKtg2MhLl/vqkjiLT+w3/RYGjanbTZfHaLONxJfiNFEJwo3zp13g7E0Y6+CeilIeUsDNH53qDUB
bFrwl4DcQIOWKU/RZEnvMGG5kNM32g3yKLaAmxIvp125Af8YcWj6A2mBjtsBZ93YpsVfwYXSmSEj
jCrzWUNiH1ATkPZeuFlAojqoL8d7kWBopZGGzyl2F1UIDy2d0JglRD2xL2DB8TPYcPtoDnDDbAP/
2A1wHpftRTgp/ra+8UcHuLooRaLr80o/BMhgE+tStunNrecjhQ62EAelb8z+GEKC1qe4c8SU5uth
4ZURewxBJefxe2lYKJ8CwDGWImtOFJpnxli5QTQmuF2vf7+IQDYCwG8lW1imxoKLYhnyiNzRrXg1
Qfj+yZGl4U91ewGWdyHLU7bLC+TJFOHvMmOM6tl23/W7PCxzlsQ0ONIi8N1ev7vbynXuHjt03357
Mwkh7HCIgGks0n28YrVWk6vBQ7Zv+u4yfYpY0e4PVuKuA7mCK/zBwz6Z9P/CwpjV6fWvecMGqGKr
yvrPL/pxWQBAKxE5oL5SouYX06bEulhE1ez7YSJuCeT8zwk+DgvHS2fskpMhODPgDXQudI/wPFQx
EhRP1rFXiuphh3eEFvAA0XU3nWsH2MHkZDOP055Y8hDAb16MdNzcsQ6tg/1SWslzaIekSxNzShEv
PpI3cJk9BxusWtuRbt4xi6WQBWwBlbSXc31WEz6iqgAv8Ogw/FO8ageOOj82DwrDit0tr/7bBDHQ
HSqleDRrc57WkscXEjWtXFqib+gtjp7aIWWfJY7gbhPtisCkZJUaZ7zCETKun2+D6ZSnZif1oDk9
dXyCvyTXn2zm4HI4sSvkvM+Z3G47Ueus03HQ+A0RFlNx7ltQyX1eiJ/FL9WqjcX7XZ5736oMZjs9
dsOu/yvcz3upEPlbygG6C5gbq8pvGfJ+LwmqG6tQBtzt3W/Vm5xYon8FC4QTKTWMNxSDhJGP8tcg
hV20HAxed9ZzSxdw1Gw3AwOZpzf0d+IGLfPRiy3srH4w9TMFjRVuBSNrs1y0xWp9E1kGFYQcQ3Ua
P4aGkubHP8+uYpTPTA5w4gflTBRl7XsYbtj+qPbG0CK51OMwkXE7EMrbNQhCFaOoZ7FoV/B+cLH4
3f2ZPETSdrcTEooXKnw8JM6V9SHh3dA8JixiuR4IsKqdG5SLKGUIMwkTzD0BVNL3uQmtkgPAaOR9
xdHBLAXF+lVtc2pybz/AoiJotLpzAMWOX9Tsz+JTaDTfRC2L0BMu7ocTuVuaJHHD04LMHJMad0PB
9x8ACpegu+mjSM+2vMaJUwl6q3zwBqg14cDEYOIrwsLdjzMsAsYTBjxOkmnDm0D3ypkXcYIqrv/k
12rQ36iEhiu5rurOotftOHtHuUH0/IAqdQPYGC5OK3pZzi44c0YWkY3PyPzZ+fGhiMcQeQNu/XE5
RKwrZXnqm9v6YIuDuuxPfjXG0anRTnZIMNT0tZFp0eaym1LYCTFySfRbe0rn1+LTXw8gtf+0rhiI
x0k3C0o7Hq4GEo3VSg6OxmGmIhY0XUDb/u4QbKJWaSb+vsYX6NZxhLNGEvnzifWkyaJHGrNnieJc
26b8a5suNbvVJiWUL2HQDQUnZTb/V1h6Lk/799SqxsIO2nG/h292FxuGjoA7sUvFc77Q6jKHcSLR
1aqblkO76fuAWgHbYpV76Ql3yNIfSbLALp8mIQ1lgqxKVMHLRcyb8/6995p7yuKwOzOShqHK8x87
96heOpKE0r+SgIRPFjlralZ4ap8Vipkbq64EQKMyEK/f4/FjUm5zBKWmyMlgYuJhHnLGFAY1mp+Q
tmUWB49zfXK+4rmmgtn2zH9CDPFC8LSH43pXRB+aCzy80yH6UcEoksvo5ayyqdycvuiUCx2zmq7/
qbrpEnZxAr7orqMwymmOqLrKIVfah3j1eQhfJV71QNRZcOhBaj/XzoeE4Qqxqrkyr5kUltSTDy+D
YKyJ9zyONrQbPsyuydiBvPJqnjWoUCCQVBQscOoGtxd2NayUqdjiVRJqyUmz7j4qN3iG4FGltyWb
vC4VZID4cJ94zBYD4J6BunxscwAbzSExwPvxXqKY4CK5YGB4xj1foTbj0Ps3WtEX01OEKH1KQbkz
AN4UwtcgcTQFU9iKfZh37o/niihuVrflv5Zx8gLlPCqG2vNbBOa/pVr4n1tbhSZZLzm9MH805nc9
qVv2uqzpTfRc9fHeoNA7eIrmMBWbFLJanMBHLqRLU4k8uYhceaRDXxgKf0W/FWr7sFHCOlBasJXj
zq2i6X6R7gypeoVNrFeCZlMRfl9cQEFEIegiznTpHBMaI7ActtwGtKp2X5yAmaT78dqUtlm4hm06
wcYjIfS6R2U+HzSvvGu5xfcVLR7V5FCbPjImuGoPmbpxAx8i3zB32RoQ7D9cgB73GWMLQvjxCabe
ytjLaFEkk2LA57awowL2jkJuToz55WhothtVDV1Y3INO/mXf5SmB6rOgVTcHqav0zU4ed2+GpH28
GgrTHp+lywC0YTM0jYvBbjWe0DknqtSx2jVe1gSJ6rLHOSyi4380zL4CbvbW6Wib15vNbFiQn555
ipZPohJKeJ+H5Db5WPQRqlNdlqry1TFXQFkCeYLJ9H5MLfLW5xABoD3HYQO2tklVCsTdltHeA4xK
3AB6DPdxSRigmOmuF/aSbuqIF4gV5isqQshB/+PtjUY9Z/jKe1eY2lzGa9jtC8wCRUWhQx4/zcAn
8T+XC3zI8uUp/KbbfXWQwAtKEm3ANrtOMt0RkcGbJ9HcHbkpWAi+FlFFiA34KqRqpQ7rQMryOVWK
4DJ56jN/Ab8bY5v5qwGfEqT7+9DFlYftG7GSrniH3aqH8pAl0oE/FjmbLgPygrUlwNr2Di81aCnU
P6M440558qkJvyWjzyuVhkj46aj4q25Dgfmqr5BI8g4qs3TfVI1IHRY7jKR8D1sVh1a1o9lWGvdm
+og6ewZnt2mrkd022/a/bjQxy6FYW/fZa1O0pLcP6vClGo6tP+QNuJfJDhqk880MzUKDV6lM/zGA
BzIg+oVL+Z+0/u6xACWiZl1y+a6sOJafxLlLF3pt1u1AiucjpdhxLDIRZ1uWLs2iH2OO33x31jMa
2w9ctvBXFz1PHHTSLJDheXYRIBBYYG5cyWEBtB40+IwwKxx9iqe8vL5JXMVDfwmK3rK9Wv048Syo
qnVkzuLMKkUWYy4rnua+EAvEtlhrksoegVQLG2ohXi47ItFcpZRHi+eL3I9hx+ph5y24PKS6WyLd
/z88WNJVvSPnKxd9fNcE2qSmAYi+YnBX4S3pMSuJ7jWz8FHURkgC1kOXi+/d8/Kxauo0hIdBHQCZ
OlIdIfE1LM/SfyRU9eDQ1bWl+VYboVKtlOZLA9vr2PgKeFunYqgwtjaKh+wh1h0Tl10fgiesiI+q
oPA72CNbEWd3NS5BRskZCD33akkfE5KomCL2Vrd47sE7jLJ47PaLVSKNhtJPr/60YGfcTosZBjKf
fVPIA7fOwXdb/Zlnwuo2hQyfDiRcNo28i60us92+VjQ94vC1msANyHicNk0TTnh9yBMCc9TnkFfJ
AvS8zK809btfwG2nUXEb7ccViGxMIz0KbyBtFLRIsMgnqJA1k4dFy3hmSa7A7CsAmH46WZ+1YqBF
0VjbJhhHMDVnNE/eztgmTW7NxVGvx67PNldVn7TPXgjvpcu+zaiFZhKeXJXwYsAVeOo5yan3G6GP
QOXX5wVr+KrhTdfL1HsXCHY+dKV4mjm8p/Egwms0bznYppOUtGaG0s5WYtUsn7QTX/uBVaLOLad/
NND455+pR9IFUUSo8ZNftH2xVta+bbD1ooc8PPnGGD9W79CUsW9EWLcTN+dwv9G4Bof4bxOhDnLq
aw2se/m4FjDGXIJaFxBBHfUo9PKdqrfTjCIVXp23nrw1He/5eJGZNwaXmS4/1Ftne4BRpH+bj8gU
XEmOJsbNMOKqS1vkxfD6g2RzWAm7NuI6aVYiAnF5jiEt6mzKYKWSco/B7tp4n+SwyrBlpKyWie7L
tgyoGWfol5eTn/RXtyW95rtksE8sxLUqk7eWzZV2Td6sWSQaj8YfNoxba8IhbLzX2haBA25AePqh
OQbkXhU1gx4vkZ55da0XVbhgD1ys0HC2Fnj8qcdMQz9dOldXgWKf4Fq9rQNHXM9FS3m9OoKEVyqL
ageEEhmLXCJMyNAHGtz2FvEyBIcxQE5MWyef4G5tR/9uSp5yAEcQ/xT3Rp6K/W5VloHKKOPK9Z08
8S1zPYhFVyXrK5UaDO1w5iP8WU7BP0GT1uP2s2K2g18anXetREpctP8/9RMhNwA0t2grt/deSFnY
c4/f1NzbdVF1vGBxVpnVFxQKLafkj6BK5SvhQ0itaQVCItnUfHRgS03YT/mCh4WiTuP0Imh35COc
H2sJ5DAMPhLU1LyT+Mb21ObmDUBUEqJ5tx1XkaNAOlWBFll64ttgcn1VjPPN5vQDvOZ60aDxI8WD
cYwcwxRHpqVuJ/8uFWmyK23G17+IzGxgCKqD0io0z02uVtmKvf2m1+CH8/Cxdsxft16BmY+Izn5d
f+pqcECvIm7gjrlizFBKHlJ3GNUxfVFx3O1MnLKFAUV6ya6pU9KvIMOga8f+Or3HhhnVasJv1gNK
+hiNI4OHhkLmEXm9NmeDOQseg5lKQkOmCCsCHX3+kbDZAtui1swh/RLRB6g9urxSmWWd7ype1C8m
hzF5R3kpf078cLmQTrMMJj/UcIKE3quUGGZ7E+fBkJQ/8OUYv+vd0u/OvGq/ZEnb+OpIw29vKsqi
C/x71we2xcBCLzolN7smnnGME3aUitXDtFOd5Cr+TSv8baogAS+/bugqb8tb3tVL8PPxt26ZZFM9
qxiNpZcDJBbJdjjXLHnvc96V+0EZBjUyN42GLU0mYiYevs4yj4BuW0NbvqEyHKzPZ+QprxhFxHVe
+TMTreuLcbbv5xGMDWG86IweXCtaV3MjQROldqURl52gtEY1r4Qcb1kmRYsPIV0dgOMW2DFoYs5U
HAMYPRSLvlJDtDITP7dzuNqm3KLdQSZ8K2SQbC43Jr0s19xqh5k6dSeCUwTj9r00nV2pZHt/TNRK
pycCgUPSaKHfXAeSEq9tE470ZIwqECmAdYUSI+QWI7V8/FKtaIAQPpppDghZsqoCy9CYxf70s8M9
tAGHD9enx9RSJgaGLhJyTqXE9lZj7mwaH+ak5qBxgfUND06g54o+/Sd9L/rcChm9NiWh/i6BvwcL
sJsGjOJbkI8k48SMElPVpcU9qWbc+gkpatGNg6VTedQnk8ssBz8hMO06P95HvnEvC3nYFgyezknX
qoYbZY20U5YxFhzjfNcIUcPwxWOpIW/sHUB7VY3qWl1qe8U6DME17IXUORFNQz7nebc8AvnmVzZd
+/0DYbTcCZYGiiom1j52rdzv5SBcMiRUtqVQjnd5PzYREf8G6ZBaGdTwxIoiHPChpttqgSUqX7KG
T6h3y1LwrUxpAX74M+/GCxJIHsZ5AL9BkdM0ON9GTCANLA+id35ENzwU2lUpjpmLGX4CFCKMNpbp
KVF12+UYs+KjhR8XMHbI+enGUZkzpaV5wO6pm4L731LX4UDS1co/JRvT3rx59jl37ssUZ1tysKHB
GsUG2+oZs/2VHk8u+j8ZTF1YUhU10YER5DzkriDA/afbs0QSKbSpdXFsk8Ulj+mHbPKW2Xu4w8hs
BXaniNBulzhNzW9mhD+sg6cfq6QkkYzbCyfdUzyuTh3dYZS3Qwle83Zdigxw033YBnF5a1IpDPoa
Se0Y1k+ItUsg2rzjRgNUP83NMvodPlb+Kt210ljCkGuhGCTBmTLd1Ze7q+m+e2Q36UnSxVORCIdR
dp9kcNFVIiUSrEV3U3FLqp3d8ix/lQ1xmGLkoKADUjtgEXLe+GPoDp1883GsRYrjtP7J+YxLKuaW
AeDf1bmpqIW8OXn8mrIFrGLqMvylgx14Iq6H3pvmz0K01+9B6D5A1akiHPhZO/ZcA9owRa1im0SS
SXTXlRk1IpxYTn/lnGdRAx9qYv2JZCBK2Hhod9O26AJIBUf9Cwm9wTAEfcoYiDC5dnxDJDfWGso0
BWS9Sufy6X5DXpTYNe2gGJgrnKfVdwMmnHdjqunwTcuwVtmPcGejJ30UuLEoq8aznje72PGQZMRK
ZAC+ZJ5QQyPB3MiACXOhR5dP6CpznlWPTsxASShtFJ+ICNrGVyTQGhNrSnU7wfFo/pA7BLldOZcx
m4wAScSZYhY5VKj5y3FEJSqwqiqfcksB7tB5TujH5ISq/oG4JolUyIi3OTTYc0SBMvKlmSOjEADI
4fMFRmD6uezJweKWt/7XfNh7kPphj2ADFd1qBUkkS7L/VDpdb4ud44IfxPXBig+Xx/Bq2U7gJO8n
0asSHfpIvHNul9yEWzrcisJ9a9xgntQWS3PdZdJTSI79KLKSg4CUuRnDzrN1zPZKkFPfGAn1GFDz
1LkHYQsUQYyk1pGkgyIEDTgxkaFUaCnCL/TzI0mIFfOF3Yay6nkoRMOXSw+U+XW+q2dwK88IMLI4
+Eaw72nk4WVglmTjIQ9OuByKitdWUmLk8YuonZsOlBwfat9HCAan/X0SzdVPQBoi41ZaTCFzPoj0
YC9Olr3Yp3zr0/VEqDQ9dCP7eLPjwX/howG1SYkAncApiAJjeMWlGMfHxIUUNly2leNeA+cLGhTX
n+GvM8IC9oVeHdHrF3cGu8uiFsCUzXYzDF9Es/Ya+8pEEEmoMehuSWeQSwCVoZ76inpiAcLvV0Ij
JcKGBWq33cbVHQBKoqPS3LeuBPzhAUXfTFnh+Ihy/aUpS4f5im37vrge8vboANuVAGRXYaIWPkO5
B6pJxKRejnfKST34ctj2JZZDf3vByQOfVaUF56beAM8IxPU87LK+hzsFP+1IdzZkPL1+A4en0USu
gOkClGumUIcTOMhyZWzLKPfhHBC6jtetoO7SLYq6N4MegwPOkpjLEWiZ/n+B418CKKd97ZoN56Lx
eJ+APTMzR7C9UphkM727uLv6TRT1JtwoteB70nsYr9WwRuVSeTRsdMq8Ogx5mlQbgN6h8z4Te1ZQ
vaanpJYphncLpNNO7vqiLT+Coj5dbcNU915ti6cPL3+aFM70vvz4dDEiSduG+rOLje/RsJg7j/Q8
BxFMH/BSISzkEAgTaPlyJNrmBEUYhFPyQcJDFtbplD7fyjyoA9f7B30NLNLNSivlVV5cCUzBDAUo
ImQ93ca03LoBFUy8FCSclfyC2VDV4gDrnFPfdRYmev0JC0EwZCZGzV2ytM+SNtJywN7XWw2tPOLb
05sAoza1jTUc15MNWAOXbNq2qmK9VtgXfXCIa2+aAaQUQ1pwBXI35aZ3eVTebd/N3vBvCzIgbUUa
JpVKW2Ca+iqbDipkQrbVInynGlQGgUM5PM91Mz2B/Fr52FLhK/q+5bTb3I7nhO3BGYN0J5SuqXjH
wZZ1bAEsazFslwO+frxmyUeCXWfiNxz9WxukadExd2pAqoxwRd7HaM9DNf1ahcrBXX9273wk0k33
FO8wfckhsFl5vfVeeblfQXyseKP+x/bpibcT1hmKGSaDJs9JMZzG52m4Wnq+18sBNoWhhc5mcDi+
L1dSzoVcX07LrrucH0hPnPSlxnbf+izlwYGUY1iYnRba7+iMy1HiRm5OvCehnTdryCEt5G5b34Rq
XhJAWoWv18oqipTGuAsdcyd2AmJYO/lPHcjFrlI4n5Cq1ZoifokHV3IbXfJgPzSlOmRN5fqNWcDU
4xb7uhWrjWoL3Hgg2blKfIKGtNJISnWFRceEnTBMNzBEb8Q7gTc5DlryzsTLVyxxTViE4aGZX7H8
nDAFOVj8wQD9TrsBizyyrnQSDPfftrbaC2Lb0UnPTXwtBOIKEGb/6X1iOgk3Xd9QF69Ud7nS+sVA
mo551YSf5WXlJzOfUNjnnbSqs3WEG7FV+Fu3Q/k3P2ttM4MXtOba0sVq2jNa72+WwS3wu4iAazTt
OEXMUqjpkyLc+2KmF08Go2gYeTexfDFzJ+RxVwsptM1XPT3ZLotrgOwdcTkePiIauopucq7MOAFe
TSW2g5aGvkTsoR6ntDtwMUEmz1gnPc5rLtvO5xNTO7O7kZNiwe3dbOjnBmDjmMSsElGWYMGkprxy
nPSLtrJ2UTWrR2wrsg78uSGGR+W75IKg71G2Vfa/QEHQdmWeMbtdoUUz3e4MCINsjzzhJe9nxke9
jpUG45/AgnmM6AMYXsbod+OCD+QO1VWJxczvpNltVDXeD6QMz6y+C8h+uM9bM4qXtzHMrLK1BuXb
sXUKTiRkyF3cMmVGnw39KQTdmmBJE82ftlJdkeuNzEeg+M+H3dehZqNSg7QO8QnptkS9W6AsqFEk
YaAGpXh7X5xgYfFD9noDUesHcAmdXvz5MmOQVgwKzEiDCXqpY67sRrQZk83OGB8ksGWwHnYLwAtY
v7QS5XNALw7Q0CeIdcsueNr2lDHU8p0u4PxY2r4oAIQbJhlV8Nyab7tloK7xdI2NvIEAfArG1mle
JwO6nm+bTmYa3P7VdGuOGOJNiKh6eC7VtM/J8el2e4k26rd5ica+H9pBmUW2uszY6PKFFcKauT57
yi+kGC1L9D+XD5vxaW9Viwm81MNWiYJUT5meB1W0JU+mMI2WrDKnN5p491aadNOjz/nOkfewtJdF
B1YMp2Y1msU2jxIe7jL8NjzSr/zN7ggMCBDewoZqXSd6MR1RIb9pwaRKt9QlKmzr3JCb24NCOrUq
+Le2L7iP3PKyIioy1XsWGWdyVhBz2AbE2+iACACn1ROayRYdoThJHE55FXnlmVy8spuSccmS7agh
J1YZGyZ/JDsgTfxjYkEgiJtpYyrqZrFcVqqmF2iD00yU4PpJ0mb8CRl1zHa5nGsv1ko4bZdSkaE6
Z4zvg5J/p9tu+NrW1wkfgYIWYjV/Pwb2tGjxM0d8CrlSQqbb707VsL4Go0CxAPsoj+JkIyWgcaqY
cRKEthucjs7hhhkDn/7d1J4//t2Y3lJ0LgMTWU1dZ2ONwgWYZYUr5Cm0ltjluWVB1kKhEH4F8+7n
6u+obzVXsJY0p5oltTLexYhY7qe9UqCeeY0BeXdJQ5+yMRZgLNAuQ3viJPGMU3z2OdrzAhlaKs2s
t8b0tAxcxFEJRG0Vrsyn9r387rS8VR2rLW0/YvwwDlDnmmwUl02VEV38nA2ctFm8fYPED2olSA5e
Ks76hAORFCoYT1ft+IH1NADQ7RxaXTSZhSF+bj7uIA2pfVfpNQD+BzrGzZPl2oUMvS+/bakvnOeb
tlEJNI+jGJAeygiVLDdRDtOkQhLGVVDvv6Al1lYWZUM7zfOV210Pm6aDiRAtgS444HMfa5PZIhwz
RbAfjEXq5wwPQ13uOjGXPUZCjTKRXH9ZSCRYpH5KJAyJRST39hdAVyjB6GhdNFtzGtBszKlNGxtn
OJCUNY6BYMWgtBRuq+Jyi9BrS6gbVpRS0ghLD1H6+9g7XIuAIih3skAutSXhbzfomjlwYrgQoEtI
tJbIK7gc7Yf/DytKOa+REl7cPgLuff0DFthU3IP+XqXFI7FWcugWLI/q93HrPR/MMVa8/mSGcu91
JBNM2/wBaW5INEqUzrSQFkD/Y3TbOUAZhCF4oR2wyrWgjQJhCNUmov81FhowOwktYCeW6bGdkHVW
oMWw+bMHKnWKdJBldVOs0OoYZUqARJ8l5WwvUETplJc+jyxIwEVJ+1cpo+kVRVZ52ccpjimiPa3M
C71A7Ea0Uo7QycCMv7XCOSqYSntVrZilQhCRfRUcs7XfZOrtgEVchgcLvpB9gfY6i4XrBB3qoyzH
+i9+kUiu0m0fVgNTbdrYAg1UI957SxuWUO8xFiyecLjtFYbmo+oDZH6pd784eSohM8d0tKMGv6K+
iUTl5gtIaDuFJqovHSmlqbJ7/SKjzxOFbdsdxOopVTkYcvCfvyKpYWDfcOujM/K4anD3L2Tb19UU
fYsvdDAmlzEfrIgOT9QoaEBf/Ub2qiYs8JsTIhoGUFyleoF8mq8LBVs8PGgqNovrMJS3kzO5t2ik
4AxBSOYQMXibNyMeOZgQkhVRqEd20+i1RQdpxOLUfdZKOflQDpfdO7ihlLQya5/lkQyK8nWBApZJ
F0/bnzzcG8g1zqbq6SRXkrVML/3dytBr2L3ON5YfWvwxg9LvyFeSbC+rJsMECT962kPItvptK5Pc
smLQBfMcC3XhhJI+HdHZTS1qQkKG6ztRyfxERqIULKKtJKCVKkALjOjXWRj3oaPAZBhevXhAbWFY
zIpWUlAzszKR1F7FdVISCpBnQBRIGNs2KukmOSHGpua8fDyYbL+pKd2LmHSijkq2jSjsJs9do6i7
/mDYu536Q2+gyBSPH6GZBRdJ/M56IdFnHNaff/Z3YZtE8NHQLxILmqKy4oluw4sFz6DTuoE3psTJ
6NAeZxUFfF+Wv08bPKd8/JZMFLqqorudr/DuB/nFyq7STKh+HfmIBWJoIxL2Ik25NNvb/RPV9Vu3
mvu4p4Bue23YMIbroQRbDz1Hziw+hT2AXdjYwmfd3T52c/977IlarQuM6hGHJdct1BWoHsdbgOkq
zji4q1xF83VT4OStp+qFynrvqhRk3mzDuwjZlk6WW3Xle+F0Pn42EHNP7kk3eKTPlynOtxSBeKoT
eFnuiZ5Z1/9IL3N8tIvNEq94RJr7Q4h0Wv+/EgH+1WEaZ3Ah31R/I1u4VZi+jc4L53vAzZAHorbI
4VTW9ybmvEVUp+fDicIWqgoS2FbeHF6PqdtkRDwWc9gtqFNatB2OmBKTUCx01RzmXQDT/KtHjgSy
V17AGfj3BrshMUJgo/MyznqnxmLG/ie6OjQpNhwxTVLihAFSFNV6be5zEehGb9doZ++42bU43Go+
+2wVW+KNgGZVmoKJznJWC2kiYH3cNnjfkNxvZw77A/zBd/1SL5tLfxglvZqZhneNSuZOne0RIzQ8
8wdq0GmqmGGPWEef/mn7feoQEUbAlZP/TknhqSfumOydac5MTy+PIC+z2GYFAaDrblanlwUQ4bdi
q009E6bI43r4SZdtMUF6R0pLluJAQzb8VjXtXj09mol+jaBiIRco3YI7phdTx+ONF8TnmLVlXTXs
V85um3+GVOJ9SDslr9KLe8D0j4/y3YX7Z307VC5JXZk5571N3ZNiW7L+i+at6stSuU+1A4V98lNL
5mMelCtNT3D56kCjQhiN19LonfN5UDgg0o7u/bJgGQpig0GTd6LnSUM5UABoHoPYjjJV1Y3HZKSs
aVahziP0mTOFhj0I/QovRxvUbXoqDcMa06Sa1Jz1MrsrLypSa52bzmFZd7+96qwiRT3zrJX8RGbM
ii0VNx20AOOU2pmuveCGnCpqLvz3i73TkDapnpjYdVN7VT3c78OoSLqeH/TWvovRi+umcqKxKDFk
LyuuZp86QPTFy7EbCeBF6gVQNJkm5jPlnsPqP6Sj/dY6n/CmvDFlVk1nXsTNyHY/gkesvzqx+MP5
39zW3h5ap6z8QwwiIO1mKs6hNoIYwuSM4Geyoknav4LDneDI7hT3hFX5YS0FerYzaArvOu1CwISE
I3HoYkijobzY87+idNUtowcF9rXy46HvonecY9rLRiuKpTIYXX4lqYAaTnhDVJ+rnhaHzXa7oR95
u1R4rkr78joU5nh5ZbuPNcm34u/j9AXqMHwmGI07qB/bsF1I3QwNW7n1IbT4LTbYaW/8tdbjjhQh
9Mv+GxNUcTWPm5EXZG27eIJ4TjnVXBF+RANMma9PnjmZR2F7+L9hMUUAMd4rXPk/FZW9SFFfdWOP
4gGLgTqv5190WhNZpI9bh5OtRBpa15gZfQDfDHjoZE1YhqEv2+3n4isaxSP+11Wpqvb549TsLn4V
ZSsZ56sz1NzoksAgLvdNEPHdbbJgO+eRKRoDwg46nN5FmFexsfOj5AukypaywwhWHieip856I9Z6
9Ku2/6aPEWxqbvczLVxeGYlVdvpIk8txbPL9cGt5Q725lblTp6HXLMWzcuyHueGtdxi2vwYmecxG
k8ibx+GownnAge0R6IJGZY4C15TY1Jybd5PFdAkp0AIgc1HyDSJlOnAXbn5AOL1q6u35P7YPhL8H
SMVXZ+3/EkuwdllpToX42oKF5oydkaYQsvnyI/Pjn9UK5jHvmxgTRM0e9HhbMebXpphG6NmbvXdz
2eodWoZozY9l7kJ2LcrnBw8jST+xjwKJpIHYuf+H7mrQo3A1Gqb/++D06GDOZxHplzExaWQkhbP2
cf1c+UkM0Sg+vOf3t6PknzQmu+uJwce38IipGMmuSOlgebtP1eRIB9tyJNg7PXyCFhrxAzushsWC
NprAquajUA0i58oXHL2ITcRJbTA7YP68tBaL7WFW8n02p+clnZUVYCxpBUJtPMDZwZ3T4dBBN+Ve
MCFA3UFCOa6CHyYohvJ41osUwEj90XHlWMfnjxC10CtmOiNjkooitHcERHxJWTrg/PEqUz+RbHOu
kq3NQ1Ky5ZHUxf79qkWRDreONQhw/aA9QvsBvyllnD3WrM4qhRTQL/1jETYKhdGh1C14U5wzExYd
FdjmLGiddhYbIC142V/UtNUafYgZZVZ4zwheLOlCGJYec3o+8gBAr5HgXSfBJE+sn040BDx+586g
pvcaC/gVxNGJn/cjGDgbwyGO3cVkubxfgtuSyZ8ZudUn1zEpoRdIivZxyjocoQfQKf+HQZAe8JiS
abRfoLEbqfR1ZgLZR5m6j1/KHhRFasaYpyzdb8N7ge+/ijWZQUk2eN7iHsU/OJjs6/3B04szIj3/
hgJ5tlsb9X+9pUzXW2OfQdgvhaNqHSh/CoeidTIdnN4zxRrfZsqYosAaqJXzj56eaKYXLGcOzAdR
8owFwdVAtqietXqL3G1EBtN9trgNk1boYD0Q8G5r/PCzEcE7sz1aqls3eJAB7OqAesOitHy5KQSG
60UuJ0n89aRl9dI0oA/8ZlGVyjlQ5ZOF80znb6KOIbO9BCWfigGw7kVx13jEoziLI8IdvC21cb1U
Zq3DEeeJ6ozolLrvVM7D4N8Ynwl+XpVNSmcTMPNrKmnM2+nMzJCS4blbJaRoS92dfVLq1fkta6q7
lQhsOVubM5VjAIUJr+sJcAqTdHw0Xe0lyHN55JMxKOo8ORDf/8xfkjM1OWK5vS/0VAaAppTQzfO8
/4VxxLu7xoc1gFWi+gSf7/HAD9jaWOq5wkooiOUhwbxtqRxA2CJkM7Owjzft2LkiGX7AcN0sqxHZ
3eERoA5bliU9K3HsrzQd5B+lUGJBjRR099R1W9dUp+UNx76tKM94qaNpJ/x1zGOEGzubMrivHZ29
+HeWB9xoMXd7XF9aTWOEXSQPGo33a+rtV2i2j31WVJXRi4O6mLz4sVBHhX4O/AAz3pUUiDm2YrRA
EAvcUT7dtZFWjf8ZxLguj3jK7ONqI83X4z7hw0JXBAHw8+lVBpvRG+DhbjHUv4O1XFxd5sSydx7t
5u8AjSBPavJ6a57hRYkyCyDlMMDq9XoFjdZfyq+WizJmEg4KqZ7ve55F9b96WqKuDeaGpZBAAqGl
1OA17NjeO565QlksKEGSZKPahmc5F/JaaIGGwxZSMu7nG6jMFXxFf4dcJfBOC4LXqXtP6nVIpVd5
ckc5YAOU6wsObC8RDY9MlvyUShTZKJJ7+BrcUGDFGX1eS9+7MY3aKfpdBsVazpKhEQ/f3GJ6McSI
/eEhrxb+gKNKTiyCRL/KugxbltwIOytdr3DofBnQU0Ct9jpiO2QQ0MvQdxVxI3Hue3EEVOKxLlGH
hRP4eSac6oEJZ1PbKhc8OveSMc5dKz12sXPpiscBMIr3Z4Lf5KPvDCxZwRjr5PV6DGNwyaz7RCYV
QJjbRcuPoIYiVvpkAIx+vnzaZy0Yvbm6x6KnlK5sKGIcOkeWyBYrJgY96bv3zCpyZcv/4OTxV6G1
PJFwBd0Nib4JglcZJ+SH53btQCG784obmrhs2DufBZhmsM3AwDrh+vkt/UCsiI+LMuXc12ccgB04
3oqTRCVJhNtG/+11to/W1sJLezfsrBCCpEadQ/nF3ZFRltYK/Ia9Bj5m4+aiKiSYGMKveZOefTYL
ObatKmFtX9CCAw1e6Fng42ShTWI0+g1eoSxKmgn5iJJyZDbepTOx9ChGCZEFcOzugKEw7k0xzYJF
ksYK6/PBxgfRoMSuMU7Xrju5njokWg5cwIygfAs7JC8zXFebdNsd8u9KptAQQCVMQO2FdZAxMKj8
J3jwSptKL/AqBFrFlxY5pIJGyDrmcubeWeRXt8Ph7fbatBOCm5LYEgns+5P+8gZmvcpoAP77ZMWq
mQC3JScp+Qk0a6xLetLuOsAEF7ER+JVKOa0Vtt1RlRoAW6STf15QY3oe5Q94jBADmXF801xjqkiP
UAbLM0qTOF/J7fwajylINN9zC5O/1p9YUJsUot3EjKOr6yePUEVDXbNm0/Ma9rQdEOu7ck69SoCo
kAevJSDBhQm6bvMVUUGvCLW+8hwtTVPlMETehdYsWz4hHimIC3UnpoyBQguTc8G+r785aF6/FIGn
nwt1rgFPi8Ry6pCJN8+427lu3uAj1Fe0ddUDdEixadDQudguWBOBvtJNfS6PwaemkFL0x3HYneap
ydvyZ75lqIBrwLWwa2HwMndH9VG8UGrZ6rCf/yLZ1zCBaUi1Nt9BWGfm8OYZmh6NrKbKDLzCu7+z
1dGZEcTJqQeNPlsXLc+ggckfeKtcWAGIYU/BfqLBC+eEvKQzIX4M3Xo41nHQxSK/mxFMXOuUiEPg
ssf1nDszXyAk10QYkElxkmo6T4DwqnX+Mz4jRomBMYsloXHuDpuWX5+Q4mL6NHC/fdWXH1D3prXn
313+E/0iT3hxTibmI5S1Jv/brhhxjMp52O22S3DGQwKPKnM4cNv/2SKuCIlfxsANK8HTVY83atdO
8NZbzuzthHnVnEceAJ/kw2UYQsPMJDI07uKZL7d7kFZwPBZUiyih1QD0VRNzSxAa8ZT+JZ1rVg1g
BsoCOTXWiPX/+3u4tXj0mOtnxG8rjsxev5FgdYCHeAXMOAoX/K14lXWvtPKo4jADpX03dU0ZnICP
nTxCwi0+mSa+wFIJXfWcw/2VAERmsgRpJCGqc53BEDb2+HxuYRcCM7UcHDhuNx374VZuvUT9JOzp
fQiYBRaaUwzSZ2ShAkmNoGpsXPz0llepSBpxa36o+ag1EIZgmU8HN2i7WAb/xmSQmiTP3yeO0bCu
oY9mIACo0ywDX2SboVCni5fPBL1aQtWhjl4F3U6b4pzDGq652T6/v5bYlNEpm58Qv6Bxsl4vhA7J
Ub7iBsUlVX0b/mzOqsD809DiexmG+jYkrpC0wbKNC80frZiH/raehIrc75YBGmPSSFh7Y21prgZA
z+ja3lIJ9Bfsuk0sTKibB9aKLEhF7v4Z29SO53MYY4MpsXRcGSiXAtSoTVruO0S5dVlCwQ5Kb5kr
FLmuQ1cu5i62fe8mQgpuay5CKFzh0OuKqrw0Nhb6SlSsYppaCY8d+KUIrlO2nFfoURWw55IkKnNa
wdhKMbtQzlo/OEE9t6YiD+0U9hlZtz9kHxN2edY4VPbE7XFSCIDA+jRKawh1YcKfR6JqXPfKAOTF
Vpg5TCX93Yz2JZpz4PGX0AXczBRoMMzX5hPKIPHOua+wdS4wwgy4iODUWjfzbHE5NfTp+KoQG/k4
fFUt7IGb0fNdptm4EDVkPzJZvHRazT7Zyj3CidwtfKUyu4+B3rq8PNHYldb8UDhzuj/70izhOfMh
QnczriR1y8xn9G2MshR3XUiF3eP4z6NlXi6WXclnLgt7XRYIZqxzGZth9k9NEMJOc7JqHOpkIrzG
GIKB4KDsWgIQErhzv+r0KLKSMw6X6DVkYZ7BvJQxWVX/Bud5aql/1k/Uf7XQDKcdOxXXV2hnPbMJ
JGKInbHv7dQ938rg0e5uCZY0ksGBeH8MSH24pvr7TNqIz/kmvjqr5NbKpajjTW8+pqHldipNK1OI
xmkh57wtAn/M8qulJS1lqL7T+3GscxtIEOgMm3LiGNqPMgWch9QrGH+x/gGHBMtxZmyJNixo7sSH
1K6ChJxarNYSm8zBcsae3GHcP3H6dzYC1Ok2S2jgkasaAa1zZeIVgf4XCqEwhF1/yESRwB+s6XMG
r+DPUcN2ui85030DKGxT//6jdMINENULCfNXzlwZDcPpWZRtOcehMCIsAoOI0wrzZmetgC/H+Im5
7nmGg5DBEyWm7B6M9+OSNDWDATViPvFuapNEh1kYiKy9fYkG8avxWrxpIL/E7bT5twQ39VwtY5u/
8QzeVdw0aKvYPLMWibk9D6iCliocrhVFceO3c/GQcYgXpxZTJZH1NUHnrx4Kt1jFupaDaZazRXJJ
47BNIkmtD1Lna5HRWC4+qJAUpFif81Z4X/fJ5l+CEl1vmqBHmYwQY/MOazgV+Cw7mLDY/xnI2vUV
PYPDx+GsTEuTU7RqNIHE4Kpz7E4RGEMIbHMeuji5Tzfq4TXzDqxwAI1MdUYTQPpq8yCmds7BuxeB
DWtOZ117v+6MRwntxL/D8+FYd5fe6I53b2vStKZvf4Z5zFej68Hjkt5zva5z9Hgen9/WpwSTqnbh
ohVFtlh/0Uoy6ZcXqJOl74qE7JHBz9+5usMTh1Zcb5Q32d29vxOAYS5nvahr0252nrWMn4xbuf8t
rP86FCdFODoApoNcJVmNFhoj39U9k0ddLa0mzfgkCxAn4ZSVmXoolFf2y+Nlzxlvxy/sJR4mZnTz
DVv2hToUujkWecCKhIdo6ZQeDdF5r4NsRAHzwDGri0P0ubqgGSwE6e5TSZfHl+WM4uCSTWlRvlYU
G1qt6NFyinGh7W11UvEbAKYPRU62Ak6BNEncdPIZ8fEDUlqt+jxa4WzBm2a9Gr+WqmdtCGlZZlOe
vZkiLiKc/2FC1qQb7G8+G0Q/wr3tT/scLDYhIwUbxMYeGWanVCST2gqET+JoUeGk4uj6Xi2i6tGY
HQ2CDO/Ra2WojjiT2pZieblCFkICwCfeAVv/QuN3SWaWRR4Lw9o5oNdW2bsmPG2OTaN0p/ruUzyb
Pdfh3ewaDpu4H4W56Afkyl5Dnd28tdWqKv+GO5l5X0P8NK9gARz6kTvm1y3fR3wTYm1avEEmpnCn
W3QTxGLVWU8d8WK+X/1obKKvOIR24Iulz64C3pkHlkPpb09LkPONVSnBJFbYR/N3K2fLfJNZsqcC
CoxjZTeY88rR9NCsc6CLSiMhIV7bwNAFrdswJeM3pB5zFEmvstepAoJwLU9lRasvpJcAhD4cNIEc
/ryziLHA21qrA+mICqhBUrXRcfllhAHW9y9eKqEu5whCHUuuxK7d+0783S4AhexMPxBQDBVenitL
HjLyfn7KExGSpdrwLJsgFrVerJRze+0WKkkIhgrM2gB+ZFypevD43/2Mlh3GboFpckBHYVV65A2j
A1bNXyp+tjavLYfeYEgfDuZau+TXxKrU/sb9yMaisqljDmtjW0vThaHM//IdUgUKQD5HdSHgc16l
+qCweErggYbiz6cuipPHN7GUro9kCjXfAXR1LtvO6feJR7/MTl1VMXSBo824JUQ+JyxGAwYneuhX
47aEauNHH4ywEdcqLSZCN0uqsniumnPWq7JyGy9xRu7h7xSV6m3Up07fKi7/6HdlsL3sUBvHoDE2
8wcwa2T3VkoYHOrtl2rLGbQxY5xafcw/77SwoakQdx6SxU8/5N+GJPOjqDpdi7qAFSC0tYjXCzh6
jMb7G57MU6xcmW+s6ZA2af0h11hI92YgBLRMTlVjHQPgFxcE1PuM1aMEa78k3x999YJGyaE1H2KV
b6zFiiG8XRf/uDM2TXQZP5Bq+783KWRdgg1HVALv4wd/MOKPSCOmCzWVJQcFI6lV4TA60z/TYu5q
ptdW3gSYQL8BMpWY0C/ILvP1iuullXUJ1/4aDgmSZBOUQg9DhaY5QOxMJMSB/F9hbH1feyoNZ0VH
YbZK3z1O071PG/sms721QO5EfPG9KNe4MYGQ1p+dzvFYOPVMrVA2WOUl+BCBGZunnfq2CAlDJf5G
dPc13woSIIWpljPTCvJgQCUYuRC/B3E3xu6sk8vVZUefmJL3mSrwlUY6yiBZ93folH6gLkxDjUZ0
d6GzEbkNU/fju3i3WRmxx+Ypx1D60ehjmBgPzo3iRbTw7SP2FjZZno+LOuW5hlljPCiCyv+e98Kz
ZPcn9rBCsDAMSiagc3vUSHtaTN4CJVSqnogqlsw3ComOxt+OoCPXEwZzzaOvqTR65O3Qfjm7gX99
B+CQYjEiiaAtuXCIv4XIZhBADHVDeQJmBdsmQBpkmH9LSPfkGspxTO/4WuNwyCGZqEhrTU+G+VB8
dbLKBnM7Daf+tEmgAxDO35rF4WZLNK8nwDro8xhEDVYhGxLqjXgK8Mfgs8tpSB5G3gDKe2Uvm6BS
WPMQa2wiGNjn3EaudfgR9mm62KWx25hfRHmAk5xr9Sp/QXwMQR66INUm0/yvFIL2DhypscNcF6CO
muikdmiM8du0ZmXdDgtY936rtCVjsJf5lTG1UUh2Fk5mIIUiTvizSu4B1HZaLs7vaLEhMe3/YC9b
+E1e9eKswxl6um5sJg1DflSk33Wuz0ZA1EL+NUj468jcgRjXZBIA2lT9F9kuQsC4QvII2RGdJQOV
nGIJWnNbvTBD7nlFDcexlVVJHKGvWBIRgiQYyK7mGj2ib/8zX+ZBeScDq/n6JlIkByDm8drYSVEW
xpGwrDfXYT+h6wIfwJy416EZZaaRvgHTnuS8cOEVdZO8VyTdBeksv9q/zVk1g62ViTx70YgYLH7j
TR4Mba6CfEK/X0jq//M3KxtI0SpyjmgEPrmvc7hJkposEpgE4HSq4gcIlTTMF8wsHovwMTh9R4Tl
EdxGAzyGvaxKgqBkxM5y0eWIizxiANEf6O//BcSnQnli/LWvrNcMVVU+79/WqXjMmYay5/GkdtQN
MuWlENsN0piD2FNa2tDnZmqZX7BcqN4HbV8VU69G5X7XSbZUwGoZb9iE8s1904HV2fx++AajC8X1
L0f2j1ivOXldzasZE46UsHUWg8RjQMIGQWx2+qI4DBuHaevmIW1OYeLMsH6P7H7iZeNnwEY60ouY
76ngDywpG8Jyhupe0iTGDt8wvU3DBVYqI8JFIKNXpyJXt6WPkxRDrW4FMKkLGOnse2Vz+aGEarm8
nFcdBcStj/V9PNIqePiGtHjMG4dy+p7lL8ankF5prp71s+ijXRP4Mxn4TgBVTeYPQypwNVgAzq+n
1dBfP79Vlrj2P9f/4qzSFNI/xZdXqSarw9akpaKNgJkn+YsEGRaRuTgRzr4Kz+s7kOM10QALYQaB
QioYCF6FcDCJ/vzNb0sgTgd52U74HEqulRvu4VooPzPD3swpXShHvnfQiCJUeyKHY4ucN2wD64vF
N4m3GMKNsncj45M5v8LzCvF0LqR9ARAWltTaXVWlk4OpFagtXBr0F/hxuACBcd7iV1MfAKR5p+K9
XOtJTSbwr539c2USa+D/6PH3yMMT3Vbmf0Jn2vloNqle+3rPy2JqkQnDb+6x1unh9uPYZPaP/SXe
EptysUBDsJ0jCIPT7bhhVmmPtT3vK/rIXxmBTYaRzFLnWS4da8+WrDmbfOvg/0Q0cQdarMhaz2LV
wS9+C57X+rnXBrlRyW5gTDsON9ug64XhQQRhMDgh1PFsFxvwRINxi5LTgbbpa/VyfVPPtJFD0+24
sBDA2HcNAZvOLshxMJpk0PyEbqBjKZwrHVqglUT26DWyyicTDG/BXU/tb7v0mTTX1zgt7JSuDfnb
WfDcWG6+QFP3x/yPa7LgcB/mliA8RWBbW18Yn9R8EvIw4ps2TnIpuqofsAm2bAi8Yhua0Oz0S/g7
9iZKUPozGgEJzJoopvgFN3INcKaVbHg1jKE9xcqwN+J0HYijas4TSR4ZNzFdAwh3fsjUsZi4Dql0
eGr7dn4tS+rGzizxJRrIm+R0Pqc8pHABLIWuOeikjJB9jhBmfZR7xuROcW8BRIxBUlyHkUlEc4Gk
yOVdeK/44aVRzuGEVyThaTna3Ge8knz039cGKcZQK3ExjNeUnOjWnyOB84D7p/Vdsd1uTda8NnZ/
pGGGyl96hUorEyCnMStsxSwWTopRCq/CRRdg7/BZjyHqHmOWBk1KsPUanTVaCw7XhuYLuWBfkjWS
kXDVfaysaKkpG8oShOdDenV/6/ObncdxQDUvaX0kiM1LaCtGhny/qPwlWoW2Jr25AY8bzu9mBEfa
xmqfv97aVZCT9gzyVBvpnFAnrF591qfvajhkSnAbRYVFFfKiX7Ymal0tM7CMZ74lcF1mTiZJXXKA
MKhzJUh8Z5eKtoZxu9qRHdHN9nEauSPORpX5gLKafMt/xfmXZvu7bWquc9x8bifn5ZNG/Z0Q3JNT
lg4sKcRMT/8C/atDge3po1yrqADhdTrFH03iAWC8sTsvhGHk3uWb7RXEwsHJyBDPpF6UTXxOEpdJ
KCgPVt5EWWgu2MGfJiB0fH3o96O9UXuQicFwyWPT+duH+LxDgPehlaYi0h/WuINHqS5rzgT8g0Nh
GVQJZ78HTaFI54IpjJtYNARJ11jhUOIR4o6hmUywmNhH7j4PGuQTS1FzBH46KZ1LvDtsB9NcO8na
juPAGtl2mHVG7xlM3PYdpUaqx4OGdqWsgSXA2wH1cYigBKCNCDDEeErbAUwgyL+qt9rOZujhs+t0
+EdmuQ6giBiUAK+YbOvUWCNKIgpPVknEMfx6PeyEPh3l1FncmgawVaQgsRSF3BUp+N5Ktc4G9KPr
SgZRAa+WFMxx0BhGASjdenYwSinIUYlsye0Kg4g1eBv4u5+EKsC3k7z34Z645u4nhtpvcQ+BBH3w
7ftamTeKho9GepsWzRatmRN67R2/e1LB9Dx8NSh8rw25eRnMA5C8TRzeponrqRM3ZHLCNfkL8RqH
P1A/YVgKBjurbyJII1lOXEGwXWXfS8pmDbvNEJzWqY7CXlreVs6UxPehSiufVjvPQJwPcNH6K8Lr
Mpi5dOyQ6IOZ7iBbzoLJmemNsIpLbbxv7U0+srXb3WN+niBJPA+NXVs4XYy9EnfI0I3P4PjOW2dN
AqEvd1WtorySG9gNc64ZHV1tGc72ezN9n5S0vmjVnYwR5Pxnxh3rKWpmHVuIadSrhpgRjrKqvn3m
PsA9qKcX36I/kThKZm5zmUREOjxuq/GKIN9KN9btfpdZuN8fQjGiOkzlUL6rjiG9AXA6EU3rl/gb
zzDRJxcGG3Hiwyr5mRPF8PIEEVP5mi2SbLgpjkselnsVLUfsTTlcvEwuuTkMdC7AQtMdXNvGVN7V
q3Un+dnCjsVLfdXpeUsK6Dp8PfVuzAop2qH3TMtvFfFN+oyHQSQaFrISAbabnOPiisYNF6HTr3Aj
LSA2+GfLl5EJvV2v/I0GWx5Md0o/BY1au9OwxTm7drrf2cOLR6JzMVYpa9wb8nH6mOV/6jIji2Zd
ZQwB7N+HuA08h1YrNHUJuB5AjXTh0fqUHsSlzx5pq9JvDs/kwSc/eSMaUV3ypO/PugjocgswSC3B
4lh0cEzDUkWXXMb5rgZRis4sMDs1KKwDi7NrdZSK4IWTMFXRKolir/SxcQTLxjZXGPE7lXxwaG9v
uaBfT6m0BQmXWcXrg94x6KvFIa7kZARovoAuTOv68PphRkdsRxDCy6gS4ux5IwRLmVCwAHb3IPX1
U56/A+W+kp1r8NyjZ2zMTuglkfqLZgIw7TqKYm8BnRKBWSmI/5qlo2wvxZ5AesKqBNUdOj8jrHQc
yAvsIVb25F9z0NOp2lUS90bxhnocyQBkuDDujL6djgsBw+gGoKBcvZ+P5dgHF2J+snIPkSUCGwsV
gudaJoHaIqDsVdNB8BNer0R/Cyj8Ga48y8aQnDJMD3aWa2EoAXqGVn2T7uFbldpHXPAz3EDqnIp4
1sxUBFXgw3cSWicbA8J5efcL8k643gr2NQPAzxoZYK3RGAvDKeQfQ9piKrtnjNNbOxhoe8/qlUhG
fzqneDqf5sMQLN2ciAepUZHwNIEPAQB2FRsNyPF27clpMiGzzXlSf+eDJ626fg4YHutbAYRfl5rv
9YdDpzK8h9KQvI5mLBBPKaRmCaxcyJMxHQvBCnZ6dTqdv+yi5wNSQpLNOJIJ04PeLFmDPPQrOU/M
Y9v+lGAYLRQODv1Q/MPJQOgxhEXJtil9Ku8B6fBgutMwxlCfSpRfP5KbEl+4Kn77WR72I8KXPfJj
Oynhc+Td6jFN4p3xEkHG9A1qSBfUf2faaTzFVHS8PTcfttTRpiIFWpe1uJnaX09/Ud9cDcMcptiL
EDqRkpmjAyS4dAv9AJ5bI3F5kZX8fI+DWhDQIia9Vz3+1uBkqdoZswQ0mD5pb5r7Lfn6nIsLRhCD
+ATybnQOoDKCK4QpXlJZZZNxq/5+xdZx5d+bRh36m3G4RgigbFezvEPZV/QCZ6M37U3N9PIXU+tU
iFa/jNBev4cqxNkKUGUtFE388OrHgEKvgFASakgA6m6BqPdulcFycdAPH8JVpEGxTcb5iyZFTfFr
X1yi3O069AtkEwf2PEWdfRM8U/9Rg4T4cC0c4rJ4lvXDvJqBcXfPifqnDmy6jJ4WUNOOqvvBK5AP
36Y+yNTMUQC5y50N1fI5pQ6jTGCe730leI4OlzFpoU/YVzNnd9QbqYt+ovxciS6MYUgZTSyMX5m7
b209dFuhq3JkP/6nV3Mne7p5rsYsxqIsa2mpXsAuwI3Tm6HI9tAqkRBpm8lHtyzXyESOLDFcvvvC
mJJmCjvAzHYT0Oa3P8rV280byiVuvCatt0uPUOnQIFh6fHDQswwX4tXomIGRRCoKNqpSqKKsL8T5
KsxEQiTIqUU/gO1r3znCvSZG2i7VuC+0D0CmCgjfTTh6Iun3bd/6FCNA8sfQVEu/7HK3g0Albq8o
9Kwimz6iJ0hQvlssnuMfvsCN/TMVO6GsweQZn4IzV3XFLa1sBo7Td6Np7x3KtRJKL9DAkiRaIzT1
W/vJDyfv/vJuosNUQP6F1zJespYJj6RYuR1wlLrzbRwnlNzALHotpEJAUpZLDxzW0vu3daKwklvk
btzeR9cR2CVtQ94/RVtRAr/R4zDqXQQfDX8ePgMLR/QyhxhE9rwkZ09qn3CKx1OhYLsSHcCbPHeC
alBBOObZFNoJtxMCSSV36dK4J2DJiWVjVNheBZ4IVtDBeMUvUB851kf/rD8diI3Ya9XT72C5pQ4r
LdHWQiQov1PoV4wP5Bg+6SPv8+kzF069MYXOoXoPFooDUfWbL9c/AwnOe9Q1e9pn2Mwm64Fcg2dY
iHTqEbKWUl/TcwfTQgxf1w+0PhwiP9/MxLrxRD4bu9u9h3AE0Hut9E3KwFZZsE8RPwqjo8clE60Q
0fdD1pUF0vghssu1xOyeGRcCDyM67Eb1THHo1qYYdQAVvvFZ6gouR1Cahv8DhKaUWStUjqVMbQOJ
kN+ZOc1zHy6pfot7p79JgVy5eP2fwzONqOrBLfQ+HzlP/aFi9i0kBM/qL8AkLxZ3Xg+GHuL9GLAW
gGCH+WS9YpzelXmaPnGiKHiqMbq9eGZpn0yuehC99N159pDVqHBTZNF0zxRw+2WoXR+GW/AntNrJ
Jt3F4uHTEDAtWK5CjHQpjr/9tLYVN39jfkYNtkPqES+antcH5HYMmIY4cye0DzMm/gQNIaWKEdsB
Tf0rA7N0oMeSELw/dhauifkNy8TaQN/ezpETCqMeh+ONwUIJ7LuU2Eu9EApTOPglcfDniSHfZZ45
iA8RAYCOGoEbrEZEJEO6ul5laLjWbZPLxisScA2LeU0FBURARTVGjhTFQdx/+EVz5drnEppBTnQG
hqfVrzJCCMMUwhLSQLW2/Tr3HLieh8SX7QsvvNz82cf+i/VH/u8RD42icOWDmQlVJsKCBQr1A4Dy
p//zuuz7GjUh5XEzOLzHlp/2xwDjDz+ckHJufccAjfHAHO73zZ463+1qoanjbwE6PcdX1vxKtlj+
IFD/ijzUYb+Cm57PImBpbQNHxp5i4tFsvkofSrwehJLXk4IYYQ9ny8bwYB2m3VcxVY92l4pHWlZg
Fee97zOen7SROKiKZGeDF0vkrxwNKpHLieDkJjlS5fehIDDzHMb08Mc5E59uvh/Tg1nRlxrDzf7o
fi+XyW9tO3z8GMC0L+KYcOiJfRb1QHA+Tn/cqBo+CSqAVe+BXMbhISCw9rw7yAE1nlCljayubpwn
fwitGqVPs+CKpp5tGO6RYJOyrLLbs9nLoqnoKJM93mefwpLA1Hp+kKLd4rGAcPiLcxJG80r6GSlN
m1qJK6GF3xf9o6m7cq4IwKHZ8TrQRMHco4W6ktyXWQ878lnNe/gzriDciJhKTwR/3xrKQ0Cx6czH
2sFHNDLAY0XxqJpjCjAe9b7i7Ym/KIgNq8af/FYXMaTzIJekpKMqaRjRrFOYgwzx1LXZ/48Qns/K
M0CrdXI1nFrbjwcIiOCvVoLS1b2xj6/BIQijeaJjA0+V8WaWJ/3wKjJRuwzFh/OzLKDb9FzV68O5
CROUfF7sLhI7XG4m8uD5UmYEYektESYkf8g4wNb8eJUx0MZYSbHnHhZJOF9Ao6Wrh4lTXPuaWDjA
Z2uLu/duhEKH7mUrWXf+/hztcmEvgWgFfOYRRsmka2Qxc9kAhB+ZN0jF4wvVsPetpqVU2El7MsH9
LkJFbUZmIvxERsYcd+hkewYXE+MtJ44o9GPJTGT3u80jwVvrkzlgjq0CX+OyeLYWYzaihl8oxVkU
iHwxkOYtfhzjegShXuUYx9HUrmRwz2iWA4RBYpCzcRzZm/N743lsp30IRhY5AtxYlJgx4yBhqrbm
J+k8TidmhGgpVmSzArk4efFGjk9VVVY+DLLZGaL7ingFdODBgHuYG0M6KdvAIThRHuVn6ckAVive
Zg8KjCRMv664vWghXZwzC0S5TeZVLGVq4iXP5sLJnhQ/FslJ9SdmythZj/D9OwH31dWH4nmMCLeZ
9HT6+YRS/3RShq8GvDkKL/vyDY5zhBVJUftN18/0nusRzIQ7vrxaKOgDsxPq2mm2K5Y47w2NOQF2
S0f+4fS8kRLttF6dwIn94MzrMxpXymezzBbs6hoSz7r44HKE9pksF+1nuOLQaYBaJ8aBLgG4oeDK
B/ivd2F5cXd7OCkPQrDkihIWtJUpMVzg4EPnsCNxbUux4gZTIaoIJUGI9j/W1SlaVZRwsu/oZZyB
CB4pIHxvp4QglVnitKaMbBeEgGMsnEljq7aOrl5Qz0xMZ17m7XTxXN+dSPmq8Nn0IFUsEXfxQi35
rs8RlV0rsXQOykJUBadnhmh3pPC4df0FOfbQYwfzOi1xQVUWhOdzw2VtjW0o1sD3q7p4tyzmjEbI
A5u0/N0epqAqcA2U0oZtz0noX5RJp629Lklder5pgytrV0Fyg7buNKoBf/PxV7Vj0pa3I6tgrBR2
kobsQRn0Tl42TXVp5b9EtA2TfvFqKsTxMLucnvVCe+lLXoCnSIy+3c9LVLIdVARC4YM6ZkHxkhKr
D5qDc7WxiAO88lXgtVUGS6W5JWVL/paW8jrA1g5RtJHHeZOZu0Y1BI4ysQ5JNJgnIGWs6lkVwsfI
uUFhmVRseBgB7f9KJdmORrW3LOY/4adXf1+LRa55wjoZOvct1koYKJ+DQh0gdIxXkwzlg3kPZ2Mn
8h7ywejcpmOK1TaMad6blJgSYLAlzh/C2mOP7kduFekpYUrvMPiH+OLqTzontQRYyt61jyd+u2tS
xxCnW+81K3TjAEQDFdmRGx0f/BogaQsieKAysgtTsQrSFu7TN8+Y8ah+cC0cW+LQgozy5uFzyR28
Ro7Y9PJvqlSpmalrETtEk8wexFHnfFWnngLfsSKczRFBslvo8JQY36QbaEyKEiigh5sIoLcmuYEC
UpnYclRfWMpIBRoNCIlEcM0GGYb92pf46dkkKTqolsxcX4DXybwL3oATC5Bnx2qMDi2IuS+rw7Qk
awS12236yH1kU1plNpmj1wZCRjqu/tkkOTmGcE96Liub6telKs8s0ZL6Gsl1jPQNlt8EK41WGyS5
S6EI1pm0ZclomHLiBEtQr3S7sFaB98YIR6h2FuK3y2JA7TCjfW/C4oB6+l6dBOxh3l70Tipo8nWo
fodFo9LLralfx+/xiiy6eRzZ1k6AqIyjhDNDS6rSWS0O/lQ90GKQfbT7jK+bD5rzQDg5ItNn2rFx
9EIUeOAT5KsCpOavB5yJBQ3elkXn5exoVTBZy76Iy28iI6a4YDXb9SrL22CSr9in3lPF5TispbYV
9jRwIyL4J1dQOM9hPHeS+PG8nQF8UAIl4M3/QrDxY6RClXyRomsm2qzQ2dVtpSkf33Q32gdqUE3s
3Z3W7jaWqQ1yUVyzITRhfHTe5PCJ5A61nqa7swoERbbpy0PEn4m0FFdvKQSoKjp/pmeZ9oFkyPY7
Q595hZFAspAlRJ+dglhx4/7n0yl8wQ0zgO1SqvfFozpcfGRFhqn9QhrHDI077Gho16xUVuaT2HBP
fqXNFPOTaPZOsBC46K33NdXVd/1u7W6KZLNgcGIxUlAvsWr5SDizqqGz1DyPClfNucMWVrCGACim
w3WrufHBm30mt/F7ACynuqr/QTdoQXh4zreDUfK8qACwoIXFGinfWj3w4PxNXFGGx2jogu/AdjbQ
TSDyzbuCPh8MZ/TOKt4WolKc1ZYOUFN9kPLc2g/rjxtyGHrwVs/xKZwkIZDYLfwtMYEOsii7DDmg
JxXbmtaSeNj0pC4ZFc9nJF+7LrsjGx3ClT58x2/90PyXshJbBxJN0Me3u9H8OtXySPgrBtGCNm0M
sEZ37EbOpOUxc8kz160S5tev+m7Svbnva9e/l0flszTJxINreIYuNjfnZtPRckUtBbCvi+fUc4Ej
5E1KTdm5grKQF9FxShe3dCF1QRLQZQ5V0o9oLgKLNUNCqsowoPsInzwG6c04pd2B94KkYeZR9aPJ
uKos2qLy4IzIF3NOQDP+/2H3r21VTaA+r4zWsPERn7mkgSKnXUqAaA6lao7eGAIr85a7y+fU8e8e
d3moN4urc7uSnojyUym9LdeP7Oqee4SOD/0+0Yxs6ITDy0gNho9WI0aOjMh77y3DmoMHxjt5WJRm
AYbjSZHAbaTLic+DEvJnCwnpe6GWtKuBNEJHrwMZjYZOp0hfI1iNRH1ZDlC7o8RhNkd68yUwwzXh
GAr21HyiKz7dZdmzUihK6dPHCz9opgFzw0aD19ekOmPQyh9jDoOY01zsTSFHqHl93FCyIY6nxa4U
B1fyxwh/hQ5Si77MfB+w1GVNJ0A9xq01rv3TLMHcv8pvooyFds+AOw/JfxUr2Vyqyo4KZDwI+lLF
6uHqm4tz1Fk9tg/BA7td/8H8+VoqIWVX8ksbQqEwCjweqEdTJ7/GaNB5/mlKu+as22Yfu4XjGG8i
x49Xd+L8f2mUkgbNxMrKUS4bffOPCSgTb7iDvuUSm9ofONPzTEnpSKbORu2K9UzWedDD7Uf8uLS3
eh96VcHP0dYg1WvDZV4w+Pj17npwEGkUl+JnqwgL2ZKTV7S6j8Qbnm3gXEIqhScFvnqHMuDAaXMG
dbUjgnq33jL5c/xDl+PjUKesImrKcVqs5dE2llfAvSn0bbalqn3gV64P2TaSVS85vt9EDmVLsu25
kEqaCpXfwUjS85ACzdX2sdEBGtUSMpfmD3Ltv+3Q8i+8ikJ0hXoH4C4kiWhU9FLwW8XDcZupOURh
AxRugf3chIl4u4+Yojab3xhWo92UjxZGEoE67A7NkMr3wtf1SvPTA60YfYObZ9pCGOSx0vcD23Zi
nkBQ+AHc+NaQLuyVpISWkdQVI+plR1dzCaNHFUrVSrkeneE4oqw84YnxTW8i0bMnSH/kVMcPiJSD
cqpYGkKqp4WAEpyBBub0lH55n8Un8GmmrpgVi/0xifgwp7VUgZcYHD/DrP9JzhSpjso60TvxWvzw
3jXv++8PTV6JgeDiubibtKvsotU0iwpfjKlvo4J291v201fe+odtWVB2gOjOHFqAk4wKuJkQLpKE
qtp4KIx7WD8sWho9ZuAyZcZsYdipYupFiSrQtu627ZiAh1zLasu5HV6jxJAqO2GFoB79kaLqz6bw
dy/ik6sHTw91CZowDWX6okdWYYfkZ+lOAmRRMdepMdSaqDJQ+MbQ8sIOo+gzY0SgkWiNS4eQAnjK
6gd2S/zbuFCNg/e0VY4io0Tc29sEfktcP7NQQZNO7Rf9ek5kH23mubE779PeAWZEG8l3qKkL71dO
xiRHtprGn+nnj57iN/NlAQUdxmORQuxJLgAzkWGmNPiVmsV4UwSvNOVEja0pVoYAec7pa1jfWEsJ
JkK9ByXrQR4vtf6Vaf1eLm4fsYuSOLvkGKsiRwvCrUsZRTGj9HDXX2alghw7LjiKLzkNAfHD2Eps
Qj/ym9sULfOkLB8ZtZKGAttu23cLmYvJDG77JYhy2rB7Buljs/UgnUbSs7i/GbqhH69tBp+33Z5x
9HqwNQG+mOsHfTm22uJ9wE+zv8zEua45Sq/sErB2FjJMPN64PZ9u0Jy8rOripYq2hka9n2SWlFas
1UTzxkNVtYDOgGIqae+v+AMs5rN1r9oaMZkW+kTOKDQLCN8tYvOSsOGZXhi2EjjYWc3DrsN8kiKV
0OkcndZSjuLiZk8aMx+SdHLfbwEzPskW4NpyRoA0ITVAARY1VKfI5q271Jb0TkRCKVNymU+kvV/q
wQhuYNlRZTfnrru0HbrFJ8bJP6f0+d5Vwgd1zuVTVJV0zyBPXycNnt3VALGho+7/9tsa2IVFy3JM
lIPctKIifI/+2JQuRNJ7gpNvGWXZQ80ci4igqROE0YI1GotjBoI3WTyI+nkp3PYFeJIb8pxfzDj+
dNGz9D7ENcpUQ9X9zIT8uhRmFqQ1o/f5Xatpa4p0rXUlCWzd+7jpimexNtVHrrZCgiNsvz5N/VIG
izWEIzS/nHz7RB9SyVUOHKZrR9C3dz/Eo+cFjIwE4QkfiQFv9YsCdw0YZVSEU+Gmj+Iz3WNjd9Oc
Sob3UUFGOlgFQwNA4rhH92J8p3Dl9iA0Ban9JPbpwf4efP1sI4HF5zLm7pgE0wh84q1O/oRHTmxU
LjW11ALmuG+wITHbPkJgN0sCHKv0ASKw9IHNWnz0gxCPmqEJak3PIGprp0HXQShYWJIC5JjhyPbe
XmaQwbumGKf7KNLX5xIG2RYW9yanAgUXYfv4HhueDWtg7Es1PpMFlPc+PLjONiE7VlKF2wAmH1Bq
WWNY7791Oh5FYvFC3squUg0Adp8JxpyXGHq4Hr8yZrzqt1/JtYHioN2QrdrZHmcyRGFLh0xzFCf+
CLdX1e/SGARXiDRf5j0xd9KrXPkoPKWR/2lkOxZSlVr6acy8NeTY7aecbKx3fIW8VrMyj94iyL9/
gcUfiumJa/VM+5l10p52dIlnPz9/EljwwV6zKm7yPQs//Rme5VGEZksIzOn1Kz3Fjpsf8GAD3Qtg
+Y2J3VaysvJN5pie1PxSr5hYlSOHidwL2ZFrg/9AA2ma7AW+dej3o8FCCRyjHD1qO6OtheOmMamV
Fp43qBBKoT4z8RS3sJEmR+/AFMJvtPxjzmfOr6fIheKZhNvmQ87Dc0OX4Z/aeLWxKjgZwqwhbZUb
t3+72JVxP+V3xKSKhy5NGribrk6J+eBAfsUpApAcszSHJeJtZfO1rjiPQh8q1cY9HfWsWflLwhBN
e0Ui8OIDIDqibCP5eBGOqhdsNnHcj/6AEhJ9KSntHACmMw00YFSfxT29qorAczdtmzW5npnRCqte
3DOvGjX75y8/CTtiC/F12XZPpZ/fxgueUZHKCfgOS/Tx6jlMtzad9ila+nRjNELO8aEL2lOhs1B7
z0oX/2q0avLNxvkvHpXTWj0yr3rB1EgLRdb18W3+isLDD8KyrVF5vrayjgR0VmnepiAkBSHddG6C
0nOGqS1XoPnM3oa9F7a9zv+XT4IjuABP8ot+wBrvQOeFbx4SSsf7RXLAzQyTyiuJAS4D0plQA1yc
I61koTrLZiPjq28vUDugWtIMMq5qxFl67m0RnT7adGeEo70N5fHOfMt4yia8vIKcXLIlb/anUgSg
8gDhc6EurZiPDIKEOtNJ5SHPSEJHQiUrcGUXPrpeF+rY2Y4OUaaA8Xp53SuGqfD8wpLMGZGb97fG
jT3gChlLACAnHndj5Zlm93XWC1/bG2Y8XIOhk56Ai5n6CmSpK8mEwv7hV9owgLUuNAhe2V0SMFym
ZUNyhb+S0WDWxMvqFweRu6taauX/wGDuPS19JD6rV3y3ImVLoK4G0WNRBBA1LRPYz1WubIgXHUiF
QRWG1ygEwpdK/lUgaQdI/LcgwZZOhc4W22DKKBlYlt5p470ch5aakBjryL9peoUdRnv6UjAxHTq0
mzW9kvZ6IL+G7Po4mvQizJYN37SPwIBeHt8R86nGAD6XUG+Y/VE4Um6qwwD6E9m425luMzQSxyL3
+vfLjUd6TZ0uThfkbewsUY5ZRcIdd3ZqnnuzlMVNW/IoOqRSz8+QMQ9QZVO2OWGfD330A4xPU2dO
/CUukVFizqvI59amxwf+LxqjGBnaRSG0FJ7hrXOPZR56icg9IbZl7UV3Xy7TnXNJXvhR4DGCrQr1
UQq/6OyiOqPQRdeKZJNWhkG7JeYaoN+exCnDe9W0FFoQhYLkebSJ+8LxcPq/EDQPuV517cV04du3
Nrm0AHXcUFmqmTt9qAc265Qz9AGDzeIbMcwthyp5zzxVKBvislIx4t2S3fSNNxU5vboXSC7k4phm
Vo6L9InwF40DizbLAOjYCiDjqskiSF6OrjLCP72ne4AYyOuf78WtH5UDn6GKuD8LlwA0iqPbRG1q
nuzXxqJcgAKe2bMVfwSB1C+/c3tXFu4jJ12vQgXoyrQIHNxYdt13Ma+AREcLA6apCEfcRB8yTNqd
DoaGvBlc/u28W6Jd0m/HG/bMdo5uziIf2V2KR3oRay1ZiJt8TFVP5d0bKrLckueD7YE2ddI0mMwI
+dU6k/ob5qRUrfbTO/EyjSj2bzlEV7LOL26AiY3hhlyTtoqHv6mglf+fx8LfKPrZtwUsYfbamSgI
eCwsk5X7cO3itDlpkweKDaziktwsZ+LIT1f/7Y17GEsQeDSihEwkEFBOZ7xAcmv3Tsg0GbtIRfNm
rOke/a+Iwtxb20rfNDZmdW+XlLVstkSOb79g6mPKfCEX7ZnR7pf0zIpK3ZT9edkcIz0MVIOgBUMw
F7Ys1avsVgqVqv/6p1wa/8asObI8uF3N87gmaIKsu7Cw4kikABnnXVrMbNNC38/a01aulsjQ06Ml
rakDLbu9EF3Vui2j+SM/Y9F0JHPZnf4J1Sq/zQUhZ7wOG6LeCTY4Kq47QyvOkvxG5zrPsuTI0IAh
Y/Hkm8lrmQ7PO0vAWDOuC+TleIVeIEnX0sOT5MWohIb5W0qoHVC7m+RZl9xtOx/X4GsQ4x9oNBqn
kYglSawdVJSz12Qp58WkKgJy1ojarYufNmwbMkVSVC6BEEAEKKhBazxKjYrq1Izph0JsGM4bVS7V
NlfoDwiJLEVUaLP8JLk8Cqz5wEqMDeTA+uFNNVSrwSGJLq93Mz+qJSy7GXuF7W1JDc2Y0Zoa/PGa
3A1sXYLlHg327xalNRCgasn13dHtO6K8yXOv3EgvqIvA92jvyJ1uYw8DLvNcmKFgMqD80FjmfI54
zkQ8bRNaxCswerI7w3ngAWQD/dsPcm3tJGKtSbj3G+7fP3bd2ia3s8/6H1+lYiXKmCLx0pFA58iF
o65EG9rmXbna6orpTXAqqHKAzvz1rtOORT8H6SnOQapAIvFCJug+tm5/5USlupECifXcQhGWZlMc
NjncXfrYAKuyy3f7g37uIIFIkCcuqLIFlbK75CkLE0L3CV7xnyklf65YWtJN3GyFwfjeKe1X4Rug
W4jpbKWHj7QCtKfyLmXfSuwAY/KHxY0YZf88YJS6gypj9rv/rpf2e6omRPI3ekrXHV558+Gs5dae
Wdwkf7zCgHsKAPVIsiyP+33r64t6GM3jzF038365lF+FU7pu4J79/IY8EuyGjz79NHAzquVSwaw+
JoRb7BlVnuL514GcohAOiWbW+y23vKE4VDqAl/BGbcnwf/bhl/kvGBDrOFaQtCs9luSzCM1bxTtj
LzI3sQXed1T4/F6+ObALt4YKM6c6Hc/039eHJl+Rmhdqt6hDxekCfJZCaGUF77awi0QEei3GlHiH
ozJ+blapaRldO3zMstGkuDJUdNJlkPU1/+elkBjU8bxJrJW5LrEMTNRjRn0usg0UU9Lh2sW7DCGw
xdvBHblI0BSEHhoT05pIqbtcwJBrRWHI4lJ4xmn0YKcoCipah6GVGf8D2y6kQYyA3J7e5s+7EQs8
30U1CAvzZ9li0hb2m31uLllcsqwgAkV9ssfiSX51xbBA4tqWXeTjSk8Oy+RfPb1z+jnooAForVhY
OCKmXCay5xKd+l5C21zLfXqoEMs8HWV6Z6rLWSXLF0nTywD04aCueIVJp6s0/UFk3t/oCk6Wp7Kv
7lWB5KyeY2KDuUH2oqK5cQqQltyq58MbTsOhBn9ir6X9XoJi17+KVSr7XHhp+BKX/wuzJDfmtkVg
q6puNusUl6r3C3dzRcOFIRhZqft1yV4BEWSzo+ZuiEhUi3r4p5Z2bZ/MsmPEGR6fYQtfvktD1oBO
co+2YEx0A6gJ3K49/pHtHTfBC+4/yjZPOc8VCi9q+HX2TVLqF3FRAjI3O/mnbw8Lz1HR8fYTZCSV
1GTGx7j2dl2SVgUgoSP5qfk5m5gdnwAkXq3Wujj3K98ll9eCs+ir369hRHX9S/UuEF8Gkg2whmq7
Ryws+3NkL1VfcIwk5f0/mAgWXbF+a/ib3SK1iFDvjIfI0+ejXNw3DlcSfPwA/is0jwRLELMbdYWo
vkAlTUGYLqvoxl2XHFQEPvrouPrfuldtSWOhe8GpYveDqQav1fVAgc+ckOXs10ZKf86iXhTPeB8g
Fgd2CVKsQnsdgu7C+OQE1YY3GhJ01kh6mepZvt4XJ4wAnvPqng9OQjjhiErxk6Y1CESJlyx1x8p4
+eTYlVdxSgi2mkYFrt2LIX4LUoOUHTmkpEThzxe7FGsY+xcq0YI8YNG4D+y/8otAv11jqQWBjmtM
EMCq8RPQypUazBADdp9/OPQvy5WLoFyX3mDtEuFOodXHhFKx1MEeeMqYhkHorsGrbQ+FOOvPry/m
VE7QRECWZkQb2xNht6WS4QHkotS+td1cgD6avnbz5yPilf8NWoQI5MjSw3CcYsyF6UuWT1cToTjL
nqDLEAcFRaVZvCou/+0Je5iiXxas4D1UNPh6UoH2C5vfL6v6M4CCcPbbPR2xypbQUr4bGDv81hC+
J0Qp4vFgNDWuw2OFDwzZbDfUZD0OyDf4Sjk7IwhzICgmFlypANP/B3EvBg/z0Cp29JvSGMSD8n+c
TIMvrHyEoynz8kiHCHXuiAEizF8fcAC4vTtZAu+nXUkfWxG4nBsTmkqPtRpXQV6Mi3wjjS+SK4Pu
r9j4tkUcBiKP+0Boc58qKTxSztob1wtACWPRuDTq0iAsCBuu6aoQnPjG7Xakk1ZGNUAZS1pFoa0U
LMhWy3BNrHYRtEDrR7EnnxNI/SzToD55m+UUyLP3YAlvcPz7TxXMz9LZ6Cb2Dn3iCgHyA8CI02Hs
f05FGSJj6/uaiWjmklYvDW55cpuCAtsB7c9JQiVA1Ex0E63WWa/fsAmul+S7wLS5F2vNU4MqcHZx
AIa00qemDiWgyEM3oWVyfi7r5mTpVh9iHQU286E96cYWKK67KNw1znjJLTou626MSY5iKxba3csJ
mPDZv5MGzSHQYX05NNAKqrW4lOXZzDKfhwuBz+a3eYBxE/M4AihyXJDIs9L9HqpmbAWcohbcksfl
BoOZ/AKApY84TIYEPHVTTLLpKSdnUb9VIGRRjhSBWhvDCbCb9o5BpO2CmewsaFlaWGoqBJVVWY+8
gLVUCC66CtYkid2quDAoLio8HmvSHvLSv2ch5nulc2PptZJAm+NHohM+2zFZ3zEmw/+vBqjybcwx
w9uJV/foqhGeP9u6x3OiuzM6WIvFKuxG0oL482tHHNKdMt4mB5FoydwdHtyBkjPxa1dGrB5Y1YFk
eVX5vo/UF8ynMQYq5E5DjLjCtcR1pcDPmVc+aslej3U3Uv3wJfrHNK8EZsGBnMLGJg/M3hNqVJcP
OGTJderrd5fLbd4L8fGI4fNBGcdC/dno9ssU/WyDFlhFjz8dqA6TuPsMqGbnT3k89aPbgAVs/yhB
og2tCZqQg5/y/5TlqBDgpjkPae4/9qD2l7O1y5fZVg96e/LdKgvoLn0lMmZoQUymXu4fYO11ms6+
sVtoL/JYaGJf8JLENXC9PuUI/CApqyYzYjg4egwyymGEW1naQCXRa7elDhuZG7AjlYQB0I4we8J9
2uhzRhvbHjt99ljdVSpth15PAYgJAez55tVffqb71x3pMytlwur04oiTUnwoJfHBYO4aatfPomBg
MZ7C2VkuiMcZW2eISRXrUn4ZJMW4cuCT42OVEzrLOrZ9xRuvIMO6RwOgx2hEVZ1SdiNrOzb7kIok
o4dOzp9GVH3IYYFvynkt1+8gS8AZTlw7dNt3bjA9qd5FL9QEV9uP1WmDh+XSUkq14f3Ca8YdjNa0
NxHZsWCPwMKm6qgpt79142R++Akmdarfrew6hgFa5KPmJEdzHO8SiJJaOruP3oQVI7s6m0WUBE+I
RKx9p2q6pgfkt6BzqEyCNveVtJW2zCRlzABrohYr6m0Nu1kZv3E5O8DPsKg0MY0h2YKJiTKd9YqS
CfIIJTZlYRrB4Uk1qFy7EUEG579TSFWcHtnx/gVHS7H1hH5IlSHHcCE4ck12dkmcG7QeAhO6SMfm
r1d4A1VuXkNfRUFKX2nHr7g7mpH+0rD8EOnmdu0htpXgz4DRX39Wh2YNF3CGQrCFnBA7QuC7YiPI
VnappMB82cLRFtOEeh3W6QIfifaDHl1s6ip1nBiRjyIJhu9+o5FLKsI2XVAeLzQ3PlL+XB7XleVF
SKyG9kJe+0tbmjPHdCcASXQ9pF6u2HC3wIDcrV+sfajlOEehJyhwPHfVX+a6yopdiIDYmC5iYCLA
ZYxrCGVHvceZdSSqpgoCuONYyqxKwrFs5YNoEeURurpKGf/fAG75gp4zF5rTKqD9OmF5xxVUQQWt
nIItmbtInrrkHdbNJR3vF3SPVZcFH2mAMIR0nZjMwDNo4B8cy5gXF57gGq1p9RPk0KnCLxWn4QKD
5kGwyQ0h8sT5+Tla1xfXHippc6gSCvJwMap5pK2JZdejbYhnDjpQEAJaHehTHlzVoKXujcI7zvQp
D3VKdL5PKj5Q3HATgJV5SzF72g2HWANGeegUpassCFGrgXXGJ0OUrmtrGX50jXTm8a007/T+WZL/
olCufd+EyqVWthRcbPI7Dga3QPJLBuAmN6UUDWoVJIc+h/HuDAW4b6FB66Hs9/F75+m9zJw8l3/V
DjQC3PtPAC2IEy4X+BOEp8pxDpvI7m94+tTFp1b04X2Mqv6xqbzwDfwaHCMrZeno7XjN02QJchJK
y0gzz1cwCgR9CsHZylwqGeT2Z3gOBdaRypcxksad2wBivtp/QiYpJNuPGqI07igmH0y7rgbv0JC5
TZ9fl3FVni5LPTBU/8dNlpuMW8P2drhZoz+ZihjARKTO8MWDYwlbheDNMwvbAEPHxrxRBaPfBhMf
ZE+nqCIuIWgpHCnlVsvjPEQ9l2QfHlux9gRRtvt5gvQrjkiWa9rZlUUbvNpKIUMzVBdYqP3+/Hx5
K4hjLQbIDHHT9qNBh8x5g6XdZhPetKHYIdgImxAco/76t6nhabsIPmwvVnNqLn3Cu/ZdCvBLKkV3
r4Twfi/YQr9vQrQKTQX1ZY5AUJPcgsSA5E3qdvn3M1u+6phXtUgM+O2/Z/sWfFfmHnenaANI5AVM
mNmVhcWdoJ5O+Bv66XAnjNbi/a2Mx5msSQ2j961Bt+kUZUzHt359vxtHcBU5J7egXXY60Ct5pk5Y
gbOPpFyzmDpyIZTRTwfCUPJLo2BWwhzkCCcwmzk/uyJYxBav20M9m/Dy9TaTxPEUOxfd7Nc0sC70
xvDG9ge19aC98ufeZljqC2WP/4d2emkCW3pRgkA67uPVRq+fE353Xau5jGfalQWCO2QUC1JHcWM8
ql6TGO/gIgfRicDKXKDv5efQPGv0/A7qN4Kal9ohqq/V7F6Wdxh871wsBLD8bnmu7c5Q6XInyava
1AMehIlpPGPn6Lld35NsUJDRh2Strp+GP9tHWoLg/nGwNo/xEnEuPkxhosSGPj+7P2g9/wChGq/I
jI9kyqXaXfbmG52aqvFhGOFC6feG/9zqU8uTV7WU2lN6zJm/xcxcqv/eoEL7UlEBb+k5ZHwskA2l
cY1reUZPcJ3HF8hEAoUvc2OYZs9kyC9bq2uQrF4j2OjpbhaExJeFDokmDkJ5xDPKJWwyeAFcwX8M
Ei22Os0kMRRe/suDQSBvy9J0CiyICppySY/AF1M2Bg+V+jorLCZhqR6n8C4ZSBFuO9ei8iUd1cJX
V/ygSJvumChlU0WJZrr6eTMBNUR88ZDHOKa0pAGkGKqiMcQi2H5NScMsJ25MYHDbF/nVOkMLmi75
HUj37QHjX9xr6HYc6pf6dHuB6y8+xMbwxNDT/oRL+W5c/6lilR0/4tI9YSkanhNoXFkdPZcVeN1F
q8jNNfoxcUSux0Xd4gY/GAJ5SLL1A54kQYvJ42HwslQk1owNezNoInp8/Eb9xHgRzfKCsc2rvUM5
J8UI4JaXmDodhgIeo7NDuJmPDFBvI3bCXZq/K3hguksLjGS17mU5TqoMxUx3AbeXULj0DThfVUar
JkpdT2DFtKPh7A48XZ+awWP90UjAShqi33Nj1pwayaw/sC9YwCm/PU1uAa/I02SgEsbbEnTD5T5j
js0RbupQ41FEqMOf09ms5uLqr2j2sfmLVTBLZAtdwXt9CKOUfZAFyeGuxVs80kdRpatugKsoN02n
eeFT9Us8PAHb/KMGgv0luOEZyBU3Qhd5kRmqyKYDS8YgE4JBUEDr+WKQY8ssqKKUTHBhsI3glN7+
m2vunKfEjE7CFwbnlHZfDhDj0TohzblhIb8v39HIN/DHRTokhGiqVx7ocbmCFjNitZ8pYiSDlkbA
L6HXd4qTTKkyrQPF1y9YYMYnh/mi5dnYvAKEiLDG5OFmS1gT42Cw3w5dfEbrR0Ms2w7MFM3XzCjc
dIyLymfn5fhwJJo/hpKFCJWdMx6ANj/WK1wjd5Lv8RyHZylH2jD35P84x95VDB442ED6grrZaWoH
LXwuNcoTKOtUbJGyx4SXV8vR/nKIiloR43ncwZfo/Jm6w7Nuj8UaiErSXisnZ7D05v7lFadBFIdN
7lrC89v+/DLDBTzBr2nR9KSUSFBX6TdCwMEl5kKNduaMY+3JGjqPr2mkZbWpVgSH4Q+esgiRRwMQ
CaQ3WRsayKovbwTnELODYSVckWo1DnIsUPcXmgyTEc9CvDdlYlk1nJPAXqGgtKwxAu1kZ3dR/v0M
dm17CE03y0b8dw5Ulwb+i/+EncxcueMKVDsQkrE5eKa7ZlK3TK5+JvAU6OEl3VTbwmuyUvt/kWbN
Q5Zb/iJWqweg+2NkTTwNJhkhqjvKLuOr0aXtwpZD9Urur8Fp+celcUuYXxU1EZOUayn5s8mjUf1f
ps0ImrFcR4tm2NTnghIBdkltmo01zyP/WzlKoprpMK1VD516pOIl+28AvPvcB83IqcazRtbNcAHD
4UTydI7/Fi0tv34esYcrHY8wsxWCoxnHSifM11sUfBvAAWvzByABI+zBgeCxtwIs/IDO9FIA54gp
cmgvS/ayXpUe1p3zrprbSooJj3eUb8y9nmIve++DcMCDjAxlRD+3R9K7z5F749k2UJ7Isl6CVS+/
fIamrEkA9eGAxiAQmYgI9zkchd8GllyUHAm4v/CuE+RmnQ2ZnSjqY7gniuEQ5FVoCuSILvEDEwf6
afNsQzjl4pK84y6oV/FMWo/jdss8dXaozT9jlIjUdibud9xOwZIa4gVgsY5yj92P1glQ8fGBQMpO
wsQUotji+HpDuDTJEEeOyVxscKY3pBXn7j+C1Fh8xHTP8D2Fa0lFHO6s6WbIl3f5PRhRgMmEHo4V
I2Ql/gPa3dlCAlqaQwlJZXGxyrcaNm1hM4XAgh9OCBnxvFl8iE8fm0hoZG5IyM0aDcLYIAjjx1qE
WQra+zJEi+ow+vp23sJ866BtOV65ZQdX5cIJxjeD1hHqzmrDwUD0IrYB3o554t9/DkqdpEKfmPye
48nq291JgFby/Y6Dh1od4KnWSvpkHNqvJe2IJqHNHf9Is0HlwzOmyIh4u/5lkDVv9qSWMTSEHMgA
KaYCfvvObByKAbts6iRov6EKJlnhwL9g0aU/XCEDPDRdtfdorc9Ohzc95luJgO5FrSwe9kfCaUwL
OGQBc4bzkgA8Nfqv5Xv3T7U9Kg7VZKukrT35Es4cs4KiGH7oW4d7hfncgQOawpybTc5GpiUwQ3Bq
MTmC+Fh4GVJahOZAwwFqOgrTHSbb0HHGl4jb9VB2mvQeQf5Z4ksacalHlaNMzz0BHCzR4+8Z7g1Z
9kqvyGztfjcRx+/wD5vcEKm3vU/FH2EJ18Q2h3gy29ZzVqsGkN4PO+E9eTEP/SvlU0m9mrB/tSRD
UrqhWqlPEkn4IE07ngJs9VPlypOWtPFqxR6szys0ec8KWVNT0FVXipk6hbL0Ax78TsusyOCv+Ae9
DnRP30AyjWbv0+HvxuOIE4Pj+4L1tWsZuc4OJWHX1qwx9hJSXH54M9BMVEKN7/6aGVpYqih+UNP6
DrHk86/Eldo10ld5o7VJRKCqSZJ9ZzYji5AaON+vZbUmeaoTDg4qf1qzM1WB0vK4epCS9woeuc1l
iVDWERebzJlveJ2f45rF3AulJkCtVPaDY9ykTFX5Yv2G7TH9J70Ay31yT4crZuFHNdC8O9DTk9+c
VuLIDjpJwqHhycwa97J5kp7pG5fsZBBPlVZd0Kq/wTSAEvsj8bi70Wdc7y4e6+2Zkf7Ptuxw8hZh
kXcbkMM6gY8wGC0/2A0pedOZX/Hs1sIbzwbWJE0rcYPQvDY7Tgzgxdk27f8jV4pHy5C0RgHL911k
jov8eDal9ru/mlvO2yqrFtqoEqIT8ePNcfLHnXJTGwg2amUnpIl/P97sEtzdD209MPywvJNDcGdz
TzvrKi6PDNUri2HSdMJbN6u9XlyRwSriIN7scaeUz85J6RiROrcKlsk8A9Fs0YMcHSNk3Y9s39kw
Ii0r1v/YjJ5kFFguzzx3JpGEbtskwl+w27sspNfYUVQfnlqSZogJHCtRbIj0s8pxPaeRKMUafbed
Evv9RsA3naUVONMDgHu0yu/RIR38LTFto951pNwkiUzVme8u0IDOoHUNzQPPIl/K8tiRMQm9mGA6
hpv2r7INt0Hb41DmVDYo7FCDcPijbdTUXtUXduTuP3BHBErLhO6HMDwqIXoUYpIzDfZGKHQf5/HD
DGOK7oKq+UjVkxae8lDYhi4PORUbCQVE4/xMnO6Kx9k99QrXtRrDKSzdQhVX9wU7HzYysmR5/At4
vAIDZpE2h68p9XvthpCOXBYA2DSSCZgIRwjo4JfsITYGFLXKWMAIudWK5BHI3OO1VgfNnXGMERHX
6d8at/KnIcuUDDydHNFMHN4yk2Z1pxcltV+jVd6WtNtfQcolqLVKWAbWeSaq8BzYn3mUM19SKzRb
qd14AZBAbezeuITnV0gN/j5fm8jRkuFQDB5llpFe8HdQ5F2vdQ44PFbKiLShYm6V8WDZdiYjaF2Q
DGStjCu89y5D9Um2KWPfx5bzJLiOHdxHV8jk3fb/Q2sdONUhL/vA0Apq27uJE6X+06CjO/OBBjrc
NqqLSpgs4ejoJJB0L78oSyAX2iTBZPeG3RxeYm0wh4xxsl0CqoKAWdWBsTrEcIqRhqBFEnIDrK2X
1/IkCA0hSsiKtTyq0aa4fAz9JU3RmYLZ6eILiRqhnB4oHVajFCFwKo6eCTNSgeblLq3YWGIk2KC0
5tSsq3M8I9JrLhC/05RvNRUwAPs2KHlPgPuy45Cf6qwG8qcCb5m8oV3EgKmVppqSaQ6Ony1/zOTs
lfvz/NCKY7hia5TuzAzbjctKvkC6/TVgDooGoTGw1gX2GIVikPn2fhh+f+K+bQZT9Wi4qwm+fZc5
6acBpYoGd5c7YUjexmFXDaOjIC7FtYgc4P/LKSeMcS8kMg9LVs5WAkeXmcKWa5aGqR9GFLHRWdJz
k3FvVom+Q6X1c/D80R6cICoxZ+wSf6hGkSqK+Qq2Aop48ko1IIz9mJS2p7WY16KzniOfrTCzljZ8
g7NJqn+hcdbGYRNKAlb1tdrs/zXca5gJSskiMTFY1xKjmKe7xMMafqNS9mqOe87qVIqj9q8sj2Np
Ptfe6tYBIBRWU0D2FCm3KXUGslGnbjSJOsIR9LHEukXyj/KS1kC+tbhHvlfFx2m+jYuo6y3rdRny
0eO7b6AoIRWmnPZKfYxQwWyQCrUqr4aWe/EGGEBqMgvlWQ622wy90ccqYZzw+MbJu2Z0z/9yhgX+
wWfdZ/BFMo7EDmpCxZSaBg5ydaQWR0eNIZ38CQDMUik9WwQhI3tm2ly4iy+pRp6QzXNpoHcrn5/i
E9UU+yi3euxh+Yt2ddOujsGvGPLtM+tg5gteYMWoytOZH+uVfgLWlfxC7QpuFYy7PNDFKs7Sw4pu
EztDps9EXnrk4IvEGKtXf3Ux6ypCsxahGWd0cSFWD+pz0Knt+3X1eJVX92g+q0Q/eFC2g8TA+8iP
5OWBz6xjMhFVVhG3UYOeYp22oQcLTZEK+TqUunzYZAo5N+8F38GxTsN2dO4osp1j4asqwMNMB37A
HVhhMcJH4o+W8GePA5Q/YLe69B+FMn/F205UAZ8OJhWRf9Ef47k7BF0ZG/lWJ+5PquV15Do0k68d
IdrAWZDtO7alVmysLNcgRGMPtEgBSTd124nyPij7Fn2kw5zoA6cS8ld9SwdhQU55gccnuEShvolU
dM008NaH+I0PRD3pqthd8ofQU0qGwv6sumj4OGp3O2/V45S12KH8HhgGmyQjc5hxoHGwlvyW1cP7
RTaj1EGRGStP2SbTuSK+T6CKzjc2dR23tVBPnssrhWRm7bD5OBm6IgR9E0NlaQsm4n91ApkO9tZW
BfVT4eZ8nB/H87lN/KsrlxR3IlRQRmczeJu9CFzOKMV87Q0tDgKUIDNIqwjqfi3ZNfM4cho+M1yl
jLv/79ukajg+DEGDi2A2iXjdd9nj4c5TYpf4k+Qi80dmebOkVkKHjTxXX4LXMUTna0sPPcKUVJZh
FZ+KJVPeqw7ejHHSKcESdTvWkirfgc8gzgFVzFsLqxnYxRVU5CcqK25L3uWN380gMf/dpMEY3H2E
t1GK2+X98xEFj7uinmtcvATH3+eIL/GPEKX9lazuUUviu6O711pH1de+B0WhshuvOsGX3zN57mQz
rVQZrYDg1/jG4z+gRyLI39Zu9zXYoMxCmXu9bWDcgTKP6GQXFmpJfQGxu9ZoA0JynumoB59UZaRh
KogOOHPPEHzxD4Zf+jqZydkkjl+i6M5Ad817QR1yeJNhATVSrNqlszgcozKuUHN7n6RRZVZhhxHf
bUFxReJbN7yE6+Aj6KJ51yFRz8t0/P5yErGuHkPw2wklBQ+fSukPKwEVZu6CD2fUxBaVZvsniJbb
2oSXu3hfq2EtlHROUx0mmCQhorMZ+dscAlmHQqWeBQ6XlNgmEKNrKpcZLiETmT2lLMTPQLWC4+su
2rCOpx5xhX2i1GgpqdgAC99dcuTwFaRvCRCp3SxuwIQRtJeJ1+qB1TSZ/1OusabZRhBnkZyCdwQK
00TJJWGPGEy54Q7cN/h1IXWG5Pu5u8Md5yP1qZUCUUXORf1I03/DL+X8empGqQubZTYllOvx9Wav
6L0xTeKiOJ5W1+74jrzjdAYBfSXZUkQtAJfsP13JpAQ37DpC5A9Lt+JKZ89/5H7WBusRjBkvEyAG
bScVa0CP8+MLD6rN/FgjQQcDTq3UqX10Rfleen6kfYACMesKvptITmLiMC431887UF+fNjLwOKz/
s4sTsCZISqVWKTEX6M9WckDSWh3JOLwQOalg8pmUjyLN0yPRR6PXvIihjAAlUvPN1/qA7xCiFHhh
ByqBar78VSAlCECZoiFnJd5pzYrr/0mxBocu+ccMsmCR7sew+JsXGpxJNY/UqhVf21zOcDfJJJym
ldKs832W8+L4+R5fiU19hR2cSREvT9rJkhtkf/ub4wAmghf5Gf3popidICpGMypMH6Pw4iHBX0nf
pCGhS/QhcXIAX4+RF4/wM1aWSrlbX4QDqSu6TeZl9TBeb0rvLskNEou/pdOuLIcEqwS6tSpAcr9K
On8b70q1O0VVHSdfKT/lwFK5b9lc/Ey01CXmCFnTTHhAfd03nrHk6XGxPCXzF/8c6H0O4wL3axmr
rEXsh9Ys+6ilXw+QimtNylbZ6lZ1qFKOm8iTEMc8nB0iSnd1OJsLhmdqlOAsVmuH8EuoP3r9DBda
lX2y5GvkLPqd26JS8Sdxgd970ahEMsDAWGodXvDrJtrfdDqMzGe1qB6rnnVRe6zd4OYd+NVQSs88
PU8Gy6NkcL0QBMxYcEuUeyfbYavualmMOqij5WixBmkhmEmAP+62LtzS8DPTa2d0xHAG990GW/Nq
twctdrXfzeFR6d4pYHpl+Wv6mccc3pz9AlAfoRbGIvi7994DeN4wsFFzbPNBnIs3DYZPLcZlE4Vs
+svkRwF98RxVi3K4nl0fQS5c3Ufnz7C0SMj/5UcKbNQdytbBQNhwSyqrOvMJuW2Xkefgt3QM9vJs
o4ycHLfMNH3TYNNpeb8mtPMARXmau1Y1gqtHfLRHZv8T9JoJjk8WsgTOplAMEJ8/TZLkIODrRwcm
vqkfdepdl81r7PH+5Munw4X4BYjZQ6ZxRuSI9ZyWuIq4ywmwDgydK2NLbdjRIHbgWtTvKL6RX3Z5
9SFEqfaLTmxz4faaVwOQgy+BWO6YI5iewZ0K+O9sc0WmvU7kMGWVTfv2JH9F6rChthS65iL7mxtL
QVB6ouKhIeZgbeWpDzihZpU1dbQ5bFjJmS6zE0ZQVC0WcE14EOSKdo0BDFrP9r1JT2vhblajFSPb
ErPioen2t6OCIqsnNQnQhlDzI5NKFfnjgovZJ22eYQd1Zq8PnzhbC87vZ7rRUTaoxHj8WYAiIZB0
uzZjsM+MYUtBZKQqJa+/ktr1SpJ6GhH9xEgxlK9sGy7hBj7BzRQiwun52Rn75gdW1z7uuiaczb5x
54IgptCtVBSL3r47nsvbD4c7DePtrD3ACKg+xtt9DG7TSnvyehMPW2+SpMelNetPNsGQHHASE7n1
EXk1RaxuMJ2/hX9/X9IDE+y4sueKBE9FgCarlFdgzg4pwWfgppVu/8LKximKNYBKhS9V+npCQK6R
OQZFNlCEjAvB8FVx+s+FqsaJM1PKwmRAoZyDRce8XwcAgNKzpxDJGZ0qXGiB2LgpLzZXEs5g/y1E
BhgTf6zNEwYOY4JkLZmlLudLkiejMxkc1E6hLQdCUnuGOfzv6dkvkGY5O7qQLBKUMabTMXq9dOb/
yG7vEdu5aFpkfkAg8kGYdQFaCIbVHKXeX6J6Qc4vwvpRXX6Alv4ZkxrV+qr2wTVCR9X8vW/YEBf8
kQdVvY2/3zU+PvmCUrbuBQGabAYxYobo+Gl0GfROVBqtIaB5hSya/Pee5gotZTNYtcDQkWoVdjnK
/zg5gqhZmEY8WTggMxEkQFThEXdEJ7I9oAMtUB6eGVtgv7tVJ6AAkzTB/OeZ9m8ZDhmETKRzXvs2
mzmZhSDCBPBucFUnBv8mU5XWjVj6Y2kcxpPFd6dxewS1HfSiBAk+YlQMXtl1BT/a0HMyQiJ5FkTl
8BM9PDUny+vIDZMNwUWEd2ajXge8Yi0+ziaF55fdoUp9ySurWuwUFvStXWbo5V/nFQdQ/pXIGg88
Z7JklMuQo/g/ywslLgvpbZ0Dp5pi1AR3sy2K3wLumwjdpZOGhjR1PfnABhmpypwtnM7U3XbYMfsG
/I5WSU4i4KsOyy3ZEX0Ohg9OhFAbFgSttXmtzKLsHttAvp/NeqepxfsL2/sXaHgjDVsWYKOG7YYR
/E7drw8vll8Ln0M4MmAkRB/JFpidtF5lW6LSMD3C197ApN1JBKVNJ8GWwJsCWDid2CN6uFeMKud1
u9P5Gbyjbs2C1ad9kVY0MxuLt2AqMXwQqsdFGRRF2ZGU9nvnLp3LOYaNWE3ap+3U11yLkgBYZ3lf
8Fhm/mAHbR/MJ2D6A1uQ6qnUEqwmthetuT4Sq79zsc5VyUcjmi+9PswkTh6Qn5/KzNggQQtMAGPP
TpeIIzn9vrsi77Ogg60zxDRejJjo/cmeC2xYKFWYMQ2zDaQLE5+X0WOES5HY74YEKmt3ekFT0vKr
0knWLQof7rIYERSo7Sn6oXPDsKd055REgvDMinKCL0pQlnH+KEbhEGVBwnon0+WU4Az8Ye1M0I4y
HL0KjHyLZdSz61qRh0phfcccPKWe7el8xBxkXrSIQrBIa0SL6fCaaJs/PIuaNGq1I+yVGHOoMZxZ
bZ7W7iclChZkCFRq7y/5fRQnu6rVJ7xaOMCwpW2MwhFCY108ru65OMye0P2yhs5+UHWWuk/rJJ1u
opZnMVsxycG5qYzpH0GcWa7L0ffPRKUgA/KshjbV10K6n6XsVoljVmrEn0CEIRnudHSIWIK+Xjdb
VrXSDKhPdFCCdkhsXchntVv+ynLancW2aC5GDaMaBBN3nX+kPHKbmUfl5uO54JVu2DLkwKoSouQx
rym9eKdVnEvAKWXF5GNcT8XJKLXvMD16IZZBZQ0rV+HFgaKNmfzXdbUykfKJVq6wXxYtZW61WY6Y
uPzGZgDitNJ8cVI3FHyIvHD1Kn9dbyFtYeFKRGKlKDmv6WENkBVwoSnfbWRf4LZImDjAG7m1kst5
Wwf3wPdXfE2IONL8jUdN/HLJLuG+ExBIyC9uKwE/PzZl+yQKi8yUvSwdzuuYCn/cYce8E5VmUyMF
h5eP5U3RgOU2xxsARY3b0Ci53Ywy44JiYxmlW3OhM7j6mNUiJV0HaeLdDpGwf8sHDlXiuqRGs2tI
XBRySultuKU3xeaAnCJoQhjA2ICQsYtsQgw3zqyvunPa03yvKrnHHlGPLwxN9RCXh50RcBkp18bn
mp2tBWoch8j17smxnHlXxkQJJHf6fNC9GjOSxTPOp/T2x+iUbqzSUuTCf9EDF0US1IJ0YxSk26d5
pQONh62PjFpNAVn+xYdR7iB5R8ZnwL+owDblh96Sfww5YcjQyGIPTFP1FK7MLvMCWsv5bQlQMjmk
Iga/Gbdbxq15sO6SF5dFTq0Y8DVTUmH4kKL+7kFdgvm98c53t4FUtQaa8NvTs3M1+NTeWAhw93xk
7g3CzXABCEnamSFdDPGVSOmnyOGtiCNKecdyDEe9IcY0kV3ORLYIM+joFY1ZPYYqSRkkoH/5YalH
WbTi0Afamt5CAeR49dyCucdZnGdb8OcoASwfT+6FndYXoN901AzwP2aADKY7JMo2qkdBkUW1qeVK
s+2JG+bFTm/AECaqnwE3hUgQqOpyKndzhquplVNczNmkzu+JiaUO/0j9ulmC8MVSXWPppLaiQCKa
BB576g1xXR8V8Js/gm9/dxikbXJ0kP0sMZ5Y8WC3nUh445V5+ehq/9puWvTvmzDDQvvgg2MwrpdV
3+zPoeoIxpnDNnEAKJyaZQ/fu/dhlxNqrZ5NSRRexekMOzYo+KNR9GIkukMEyJKYeCMil9dSpgHs
tRHVhwYU9btkN7tD0JyNb5Y6cT6t60cCtrcBWX8YYR8cdR8n5LDyrTtgS2qtKlqZjvocBzVIx1YR
k0Rj/yUQeyUCqHf9Kl4kBm/LxNnB1b7ulcCVyI1PCgp/v9JVZJ8gNWh4fl5p8Dt3OU/GYU9XB8W+
rTXD70L+c5XqCFLZO4vsxdwYKTQYDdV/kVYVIyNyFEjejZbHwJo06MTqDG75iUw4hVtmtEoWVr0E
9+3FwAFKa65MGw4AboZe5H25chqLl4P2UGb1GHqwPFtpRc5CSJy5U1fmgqBWLar6547+u1tySbzr
5rm1uIfMYNr9ihx4YVNbXez81a5n7EDt4qQDMdAlp8cQD2dZWlNH25jF7u4MMAGGgQfpncIt9Vlu
vmyImWtRvuahxugMT4aMvooxFGryFkhfZIVn5GgvWs0qUikCjLD7FhtRs9kVzBReTfgIneRIY48U
0+wKNypvYQ2bdof4EE3+ZsTd0rQEd85C3CwGeuMQPsyrVHqDpwIQLglafq8J8FuIRzWNGEu4VciL
baltFzQEEUK06oYQefNDdQdde8Zjqi1nxuG5Ksz4x2rufSARMR5HTnR8gYDRuT5UHY6bYTo3igOd
5IfAKS+CrnzfgkNl5w9Y2W9vFxuxoPKKn9NRz6oh9jESw/KbUFRzVH64DXQNr2hpIn7zfHpcjhT+
b1BtlQ2P1VxG5TGSehXvfnHWMcWZN9V65Es1h9KWGpGV3n4mCnCchuzHF43ELQVqGr/p/VMOt1EC
N8lFcd87ucCgjMhO71Yw3/aIlbU8emcrKUkws6RlxP1v5KgatYfaj9CQ5XbptT0WkVcZZHXj7r8n
pd5EMmVl34nHxa1DyRe5QVRLTp2WwjLKuITdBt9bRAbusLOMMqrTmKJ2QhcOR5ISCePDKqYA3m2L
Kurj2a44e5+WTn7nBEkPdWJx70bb8UydtwgfracMlY5m7YSy9kBD0j3Qzxh13LH4Lqisq4kBJrMQ
fHuJquuM4h4esInP7bfalQUoFzAW4D8AXXLVWO+BVYWpxqEf654q7K9kveTGvdNkUi4TGVUnD9SM
8UGEBwzBF6Xj2GhFPmLjgSDw3fG9EMO8rAtNWqRoAkPuRZzhTznkWzGHU4APeUaBH4oFSQIfJTlN
PH9mehbrOzBECMJwQQ/AYCDDwaeLALLEf53s7NRoyETI50MDYNQCF9EahlxdvRxLOsCmyPNGTxQo
B5+56e5K7b1o+po7OZz5hYte3JR7O6TJqQynmk4qcTUKqIu84+YOVcazLZkv3FG0bL0mhM+D2pzS
i3XgOgfMZe9cBj0uZCAc4t1pS6LQwj6iePeXwkmCNAFiHVu/NHoC+R4MTOg6g7qxWDpMJR4/CjME
YmGKR0CRsRxoJvjrG+cLCvs6KYizzqeUZfRdeax5aYnxXyneuEMclIugJZUf5cn7E6nBqHbxq4PT
BFdo+b1pqvkjOdaw4TLvsWBT1gCcng6TxLpQJ9fkJptGxCz2e1aUdPSpkxN1ZTwppD2nq1g6T5s+
nXXH687QdvNJqlTYg5M/MffTe7K0+UQtiMcVp7+ie7I0vEt490EZCjVj4uR0vbjrgiP3c1K673Oo
QhTnrLxAIwC10YJDmNuOCRAhqPonZJQED46BAEM5+4Ncgv1SnxuBIdLSoFklH3DLuFngWlB3cmTG
X7R+CQZR20u1WiZJwr+Vl1V607AdkwjdF3ArbbXtEJb/rKx+mkF+sFEu0sSTJFhsXW4a5aHEjKTd
m7z2Ad4+1HlpdT7y5djWe4+pj0cn9LhRa0C+TAI9UfCPhWqn1iFVZXli/EEuMndXV6QaYYjyHkmi
uR8NUYechAihqLviXnIthAXD470ad1/nx+WBZdgO5P+oPUdEHEB73wvSE6Ui2/ga7/BFvaI0SjRc
23qUsc8iPfjXKMOZlaDi+TJhvlh5iDeLZcm4ws2JCztaMetbwKBWaMf+Ceci7lvyTLwFCUbuNO5y
P0wkwMHh/TTX60h/+n+TH7dmfTEJOQGxV69k6WMB6tVecV4dLuQKz/FxxwvaMHxlVrNU8qfQfZ/P
ob2T9OZc4rD2JkbIZQpEdjj9kQVJBMnA+q+AdTAt3uwyLMMc0HSBeyRf/fXgSDaZfH0/PY+2PZZ1
trS+MlLpPc1INh11m8wPSiyHLo0TaTYF+5dCIlCWQEWJ61HvFfHUE61mmExHf+xXDkkhrVopT/Md
icEzUkYclln6+AP9tUNjwcx8Azzbbvs1VvPql+hGif7SGE02iJBZ3dMzip7BWxukFuoWrJRPSANE
alk6YTiuazkqqEtS+DY93B6wMTz9cyfCG18bt+ti47p8SkoP2RGLtog3K1clOeOvk8Yo3B99V/c5
kOvJHGxFv+xA0ckyemjiVS/yYkCXg8YgRB/FobtL5mKX+R8KSeU+lwdNuQPk5BqYaTU5CZaD+XE0
Gq3P1IRZRp0QE31XH73jUTqoYZux438IhfK0anCszFUxn/pcHiL9rflr/Lo8LKwqPAyf3CYcC+K2
Oi2QBgM5f5Iuo3gcPK8r6VyNXtBklLLHegc6jMrl0K/KPAf8JFaLH4MRPmSpgJY6WDZThhLb8BkV
6a6err9RM1XOKmM4ieLPmTGJMmrap0MIHXCjEb00KhrJQJrzf5lSo9zCh5hzGhEgjGaS0wQGhBOV
lxLEH7pkB2Haj8YFlS5ZToUnNSdJroZDk97qPxHefHnNiA6KNSs57bgioGZZZqU15+lFmRRE+Jq4
eH7JTsDZjIdET21brhoTUXFbUGcFHjkWQVC0p8XxpwM6EoYU5ApuSOxu6wfCe5HcGOP3l0k36u5g
xu3FflCKLIQVypKQHK1XYKIMnl7SAN7iBADm3WPfcWIGFadZNWPixCsKd3KGHSisxT07qMqZASMh
S9nu4y1yT1C48EgDricu9y/XG7yco29yXuQp5rcHUO9e8KhEuPvvYdMmPBE9UXDs/duLbkcga5r1
/H9mfKtyqzqRjwLlPwwUs1n8nAp7rh9wv2HMLI8Co32HJaNwgwpAmRpp6LXIxtvgAmD/AL27EEhM
dQfuMG8FpteWgUM5W/m6QErXa1fC5AmKMOs+AqsWN0DQnVCeXj91tLF1TQbEb4KRgG5YoWYZ6iu4
UlZR3rcjYbZgI0CgXAMncwT0+28iCYuhPUS51lqERWa6wqF7UeXnxhG3m5C7FoUiJZB8Oz0ePAHo
knfUvBerC9h/msqXPCwP3u7pu/hHejg+k9iyuKQ3RH6WWfAouO8qDsi8MrnfB13C85qVH8XknE3Y
Mcc1z0NzekKqVfuCRM/HKqAenbGaQQBMD2S3dPOM9z2fGAbu4pK8HIuWRM07/BPZ/b9ZrvHB41xI
lwG3nvzqCLBxLYIKP5uV7Ys/KQWoHTvCfW9l7a/3lhYaQG6dfoMQA4jvQ5wRhwjdLT8F7q60BGBp
NNJ3LWCFwZXHcyq39gL/F2AIPf0Pi5bRHz4zfxf7SAUR8jQo1J9/1HVGt3wMpTT3ak1/HgskzV9g
RXcxTAOBE7x+/k/TvXyxe615XKDWOQw10zWqMMiLh4hxU+uJsarHUxHTyjh7f8kOIwW+zPt/Qfje
ypPHLLL0svt8GPrEQB1DQIrBx7H0gsCjtwE3O1xvp20MJcAB14FEpll40ynqCHL2s2fIotaaDVJQ
RZW8Ujd1lrZXIZrKeWySeLJRboDEYC3gZZR3dc0oKsjvR8BEC1wjeqNVFWEnXl2Mp0ylmDT0eJEj
gB/nri2WshLbG43N9L58ol0aCtbNVmaWW5yQllwPNdQO6840bWaOzgAT2Ln9EyZLIALLxCZl9AUu
xkQjlJIC3sBe8tucg0S1yCqiSKsrhOOkNlvnfVAMabDWJcD5fHda891fdn8jQKARH50nBulrUBre
At2xZi/hLNgKsd77v01g+Ns1b+rfceTpzCnVp3RpkRoejESgHE3Sb1wAaF2AkBbS19//diW/W5dT
qkDUK1reUGdbs5ProXyrwo0tOSz+XTmJvYcVTBTd/fOGnpkuWV0tUzTv/PBx+1q6OuGhrW0C8aoV
8NIjyC+TLH+03wV7lbS467RL8xQdgfubdp9jIJPFtsfPyao8JVgU2bW017rZCqMuYfEmp4jwG5sB
SnuwwQ88TpeyjE+sKLXBUCEt66H76e6dIgsxrlKdLV7Q4WuUlufhHpcTPW6SuAi/XLd6knEdwnFN
Jyqyui1fVj1S7qFQGu+uXUYnkOLkVP+ClO4sts1N3VNkVUssBnNBP35pWKN/cqNRJxe2XOaAeRK5
mdYFTN2JUllBoEwdU7UW9PqYCNfI4Ee6+teTdac9CkQ/L9Tt1vfPuQ2KYZfP0TsR32LmgvIVGAUa
O0n4UGqsZTucsqS4WfkNmkQeet1nNQ7JN/PYPeQoMPgrckNE6VfQOB6sKHcY+T/7vBaHsms06k7K
rUOZGvGRSK/LY9aqSSXD00sWRYTpGiKdDM8S892s3KBjMbIpD8xY/hPyr1uNuRcWkjn3DMsrpTcZ
f4c6BXLnj4AD0mGcR04fMfSFR56xzOZtmj5+Rb5sbLEPRbwCTmHRxw30ulfdR+cNBdiJp74qBmvP
YL3HZQF25AuSC/gQLYLLct5hnZdYjXTZBGi+mxDhpcqr3YJ2VmNbGoBHHXaup4a0AYq3euoawrJx
iMedcYpoM3QKvrM6GaaDbSRWg9C37cNGEAfsV5jyGs+Y1eIhRZQPViPOIRUPPWn9G+YycnlBbO49
eep4u+aUNBRbDidkNgQDhu/4Vtu47G56oNib4L1qwCQIJb3JiP81WATXgkeZrqBaChGLwJVIjsZM
fyZ+F4ggcrEbWBZKIix2kYxKrQurSlV8VRk1nJKYzWzXP4ulg/VJDn/dqzXh8c2II3CTIHgJ4lTH
2AXlHcQD2ers4okJP56z0x9siYTFTVTL5Dutug1G0994J2M2wNjWW9qL/tQUnuawE5HYXdgni7Pa
GM4+mX5slA7veAPPPyPc2XV1DgbzM9eOhjs+hR+WP0aBgirXjfE4sChmpsj2beqr/cZHqbrx1jlH
D5959X48yn5ffsqQCCEtRpt0dEvhJauHejJOC0NSNT4qIrPAZDIBNfk6L25R63xYf/L6VHng8zBk
JCFG7vXtKdNF9Y197IUdrLIkHru/XbGM/B310bTkuPGTFA2aldfbUjK9xCpuEzQFqwWtKjBmEmet
siGjKRMsjNQPx+YUlQQYthy3cbU80G8G2KuyU50sGH/CzYaZux4lFW6MNfoyndKphafrqItuBMEv
X69uOihAlHIS/gz5A94/NrFCKnvKSns75/B9Ea83OyD9RTX1aDZIaRWx4pCpt5E28o+BKHl3Peb6
eBwMnVXaAZlj5CdLNT+ho42jKlDF+ts+X/uC53BpdCXfVXUz5T4MrJlg9boWQF4dtH/UrRJvW8Wd
Ejl7FkzGVR+XRPnkd+OqfAijXvp86yx6TFxIRS8gxSvCPapDMK58L3dZRFqpCI2bUNMgPIQCDmSZ
oOP89IUCp/Zo/Ynmiy1rD/Nq0kbIh+8ufgZ0RcST8kkIDJik0kR7WfRxFmSnghzAkpIkzbJ+OidS
wMyz6jw8pfXtm2VR7aBWThsf6ZE9L2e+oL0x1YplC92xNBtgMJqh82WKTkl0Wvp3grpewtQ0hOMe
jhBihu/vCtOX7A4gu/LFpJbe2psvTaRZ0+09gUVxdSjFsovxT6oSnfFEl8n09zdlMgontyo6k+30
rzLTFP9L7HapwKgjCgVELni+rtxbgs96GqmGTwD01Nvc+X2kKu1cLvua9DQkvrf9YktBVVYijGhm
1XsTTvF1IXcweMnMQqN5hkphkIH3tvegH4J0w7Eq7qW82q7wRv7UUWn+onf4TDP6INu1Vn7uiBCd
wL1nfInOTbjyVjqqOgABaKGA3k0Cl7lmWR8h+LLtlYgUP46Lji0IOqi4eMzZVqmwIl3bZ5tk+9jr
dF8x6HKX6a53wLYq5/eZeIpIITzlWtbbmu2cfpFzVTtiobFRpYNoHHiQOry46/yl1kSeAQ26DZBn
6gsJLQ8Pq6AkXfCQa8MC1bXZAVtRZ1gK2PIZWtfBAglsi1A2TOlULiSOA2ZOzZ3YSF2Aq+uJ4yNj
AwrfTogLh+4vmG4+5KTiytbpWLNn6m2e5OjjLIl6u2StDY5Er3/tA9xoJJGi/Rvr4/iYD6P3CslR
IpuldruC4ly23CRBuru3MI0SnlmKJIn2TSOds89hFmBjjvPk/HhuKWwjSw2oJ6M/8VLMcfP3okPe
aauzo8pY7d0jroqHlpnjtHVoSWQH4vACzbd93dSfVNy2+h+uBDWUKHYQ/9JahkLZwkwxKcDAyxTI
q/4PLg/+3BpY12F+NXfRQNlm6a+CpbWc7sE4pdwdz3N4CHC796qV8dTZvQaZ9KTvq4QSb57UxhQB
IO8zyf6H+fZvf9Ra2gcHrAhhB+6Tnke/ET1DCLQ1jerjvnDTXtvLsAGwwKVxKWs2bibjOo75I6hm
j3VX5jpU4ZO4enqmcIHDTDFgBmzZoFYCqT7bTtP1G1iDrSlMLEJYjqzigGRwIEQvQ17DB84Mv2Vo
fzWs7eXk1kz9XPA/BjdAo6Zt54Vaw1hPQ5znTHwvJHtIYYiP9NMSJbnjUM+r3FPRPW3OH2Rp0Tzp
tKiCk8OHyhCAlgCp2f8groQoHir1bn3yZbsOHCC6pERje+RbFFgLcQKgvpQo75rQpfUqh8ddzQGR
cBYVOQM2gyTECGfRktbzrboQkU8sgmvbOHof1YSjp7/rQIV6JEzsYWWG0w77eyzApHHX4hDgWg8n
d8TEnll+qiXA8K5YSw9q27jBCG6Z6JuNr8DV2Pby1DG0s318Gr27Q9q0pEvGKMT9xVcQefblRTEh
nwVODUpb8hbuHmf68GuagG6T4SAdiVYnsvrN8DHq9WUEg08b0T48eAfNj+n2g7Xp0gNxe+JjGO7o
6xo52jQ2SMTc5zdFssHsmqWpI4Ka4qI+1RXFcVFl8CBCAmFCROEzgLURgo7A6aS+H3YVdEHRw0JR
ZAp216ErFjb0IznNnG7Oz2KvD3nC9Lhi3ABg0qdg4BTTL6rcXYsurcmfq+jwJPNbW/G605lSU+qr
RrFkOSjxlRxYaF2451T7CxtUcCTk9hwjv9BXCP9VjT++3ouBq6jkW1izrGKALl0un4pz3MLBIMhc
2MMMdP/ewHpWvQyWC8Ykt7ZgUq/5mFBaH9X+2RT3J/Cum31LXyKs3x4K8VPHUFhaK1+f21PbGtDq
22H27w3N3eW3TJnN13cIllQtTO/oTiDfLddzetJjLS9T4L6nf33BmjSXzsKPPDdKm8lL4kq7pFpI
5L8BNNegFR9eqUscq22VoCu10eJFzZbUJXsJTbLto2qNBSybT5mU9f3QxxvX1RrVToxCfgY0r452
9JA8RRI6/Eui4pjSUgBDWXLNMs/Pu7ThTmmI9zYb2bGDZSgvVrl5ZICqd0Vhh+80X1XP9Km8KLVV
ZHFijWFE3S/6jTtiUHwurX9s8dvhm9O8IeE5WiHv21HkeLxj/hYr7GbGqOnJpdHCsZnhDe1oyvPx
vSOXc3yAyHo+MIPg4JEGxWF9j36KSItKFpZ1wqQ7zmm+w8B17tFP7RGoI/ne10LuB9VZOCofu62W
vp0IhzZDi5sx+s0Uxj9HwMDFiOSwnymE4LFzuWBQDEkWZ0oO/h/sQNjPW1AyZ389Cix0yWkHTGd3
OEMYHsvWNsll84Iobg83YHE5e3ia1q6B91JEUC9WqTCT8QXn3vFnovAMQu7Mua3xCIuugXrvnxor
1+6f6kSuTmE5hkvsbEtxA0vW/op/+h7OMH9fgnB6QN7BlcaRK6yPNelB8OT/WqSs/TxZltq8gPrp
Nmu1r6HQfzwn1UepWqgBDVmNjMeoLnKd5CbDzH6qiDlAiSI4D6bnzAPho0AffI+nBKEvFSeCwj41
ElOxzerWDkqX6H6isCQI/LwAQBIMj86kilDwOXorKeLA5ZBwwgxja/cD5oaGjl1Sab3qPAxsWdH6
F6Xp5AD0g4yJt7CkaVuXsMSuxVkG6d3+WqSM9OFXC+beVTBPsj77s6CSoPwnsHrTd2R8YUUV5BqE
VoebnEp8O026ezflMWieFGqhSGsMQcxObeugPqKkZn5OaVaQeBktUX3CEKCMbKn8tycOYjXGSt6K
5Mc5mhd//1DkLFoFsYZ35SrANT/ee84CaQ0lzMA33JiVmEXescxYgJEIoVrRvh5OeX4SabQ7e20b
G64xYcOkyNLm+d14Rm0jcvqq1NL+R/k5mt0DoZx2sL343zCYcA089GuIatk2esmL9+o2z+MgtOl2
ydRLBoahf6stRifKuGHpTjDrtTnX0bgeBUffBt9GgRqJ9CHYgDfTmW1NOHefuv4XrzXZHNQUitTg
flQkihPOV+DvBCVF/tSMnE65Ecf923CZZkkA2y2k1FPlI8pWVIYrHm1RTb0AQjd7HlmWawTq0fSp
8Qk6Urgzforn+f57ypmkMtTz9q237Ifndaixay7XvF0fzqnB1R1mtmtPLqK+oR8Y3J8R07GI9lTt
b82LBI7ZQiVjt0SCOIaoYoqPLBsb9BLtcXKMSZTrtBDbcX/Np57xDRwo/huT/s8oMiEIWpPkl+un
K6L9DTARXqv1Zs1z8dnxAdWc+XkYhMYAmrcmS7VtL8uGwdhWAcox4nMfFDQBSNMLiobzVZQ/esaU
q1yIN45VxBJYZSS2USwoeq9Y4syMDJwyCNOFCJKAFSTZ5qR8GwHQ0ckMW6itEsdeWhbxXl0Wje2U
RqlTFCziPcGfxkfifA1u4SakPOccQZdDzDX1jHLkSUuWyZCsJNp1BTpw+IzyDqWTahd34Kdj7QI3
WWvMsJtv5iOOiQR6myp/TyjItHv9gVC9eUU5Hd22/tmSpluaVxIlXkWlUyzY82P6q6zMgAXI74Nn
fGoc0mzEXbEyIY847gIU6bKFHXwbAFBw67783kb2Onvh+Joa2pyhL5bES2eMRtyZuA9+1AA7ztdw
A1zE6qvaiIzRFEFVPkW+RutuvEXKvjfK13lYjp+zQHTyTH8o7Yu4sGRCFq8Pd4ZwgK0Hk68fWAAw
Jwn2tYGh49PsmSLiJVGYB9CZNUCrvvUsqCYhaCG4Wq0hUlFAOoiCyVF3RTT0ZuYLxiKFrcpOqz4R
PfmvHIBYMGnRNcFbEl7tRVf9FsJ4Yt8RMp9L5oiMB5D6tZ7JlV3P7tC0ygAvBtXWnMcmVOBWnhbg
PlykJ9vXkMs400o5wkoM3Z35LDoJAQPG2c/QWv0twK+VEA2TJnTjUa6H+G0fEJBwx7t5W6Fs35OE
Wmz6rihipKQ4axwyBcnbsZ7JPLmb6AXxwUW9f0w/kYsq8hosXIMh3v3X0/R0fIRsvGYWDxoZo7v7
/oeNLY6uzGITpxSu08EL+MaEOG4Dw+P0HrSFRuSoxR+4Taz74Nk7m1POIlweOQbKLiFNVH7YG0aM
6UW4GNmtTQZLYQUmRc7vsqk0TPt7fWTdD26FLz+tgSAK6w04dwPhc4GvDQT0wCGxe3/Ne65ryuW0
9VrcebrEVzu4G1BYPUHS+Se13rLvJ/XUgCTsP1pz3kYgnZ/l9nUbcNrM+Vjq6sJpf/MpFv5hNiA4
klgSJUO3X7Jz3YS1mH/0dL0uqElC0HISL5Dy3PEbARWNGAqqTXDUY1zkTavtZXqQIooHLmws/FMe
YuTT1RGhXe40woyG0G99+KomUpi0GAYfG4oftVAIwMgIOgj/lph8WLh1QFJGDmcU3opktirVTHIv
aC+naTkS36QC/eMzXeUZoglEGdPBhKhhvkvz2msQycy9dacHlebOGQxVho7DEZFPXvpAzimfqNvx
aEzfeC/mBp0UBEcTGK5vjXkAqVzFlXNXdLvgcb5SuII4MNhA6mVCOYcKSGbMINSbuIxAefStX5vR
UxNOni+kUfsycKpeOsTJhIhaQUofm+rHo22rub/kOv6JpWsoLMQcSWG3zIGHkOAL+uM9sMYVEdHo
hg8hXOO7qO4FruPWUHk5yfIIHMUfK4XaBnxjuQrHzAUmv/QBDQVkxA9bEcVxyXMo3zmXz2AfW+9C
S5kNkr81DG6J7nPlJBU1jINoOC7armTLn0qJ+ey1OruBU+hEQZojrZ/LKVaVf3Z9xRnd5AilU+s3
/1xTZLVH2bXvCFfewyscYBn0fzr/D+4q1ih9GrPjod2Tj+hR8uHA8sAFRvdvbW1nVKXAMyIIZPyt
m40IbSe25c3cVHtB3NE2JloJ/mZTRiOoW4wAMi4B48pgpnQo3IBldXwAB7KWKXNBumYm0x/ekdu/
B2dMCRf2sonQsOp2D2HWUc5v/jynS8465kTC+OH2gyY9UG/wJ2frfjoLsDXw0246fcmEsydHkyW9
jB+D6B60Gkm25880Vb795IpNt2H7s1akH+Gxn0fvEn7W9rjFRfzKAM19QDMOcKEL2BUtOD2GW6xu
EWDYgA/fzLTEphQhZq6fofDs+6B7/d/lzArXj8CeecjmAlNwxyidKE94RCAyptCZ1x2MrU/hyeHE
61kQum9yyNZbgpDUvHUCwKqjDg3XaE9j3B34wN1jbgiWX2osKVbdUkWeLKsCcYMqZsRGrdSkcF/6
GJo/wKmK8hidcCubkj954PN4Fw3PYipZW3sqTXmgOC2aGJ95ffg7Rp5WrwNw33QH6jfuj0VE57gx
mdfmZfjsufn7kG3zoilXz5KvWSp2Ddrd7g+b7AkjJmCAVjGYncWG48/EmYYDtV0Tk0aQp2Efa3eA
YmChaSmghvaVsa/k5FMyORlTHULjdkZmWBu3ouRWWNNp5PT4DCJeDFBJbeMfaWfq+EkNMb/jA9J+
mEn26yqMlQ/8PHNB8I5lWlGMwj6NFJJgiNChhJtfTQaiYdqdYEKP/RT4BmDZZ1H38WCZg38e2tP/
Soodn5T+uqYabmE1poHQfbTL7RDCwmgCFqZRvoDSPv4Y0xvSCxZbYGlPKDYN3E7RoFqUA97AdjdT
bUmPs3CIW/Q4QBPkG4rf7Er2T+Ex0jp9CJneBkoXSUyq89rDM3gsTzrIWVRjZn6FfxmmHVdQrNeG
6t4AcF35AfssbeopmSgcAIns8FAHmmirqMzBZdXntx17q7Ngp4FxWxQdNoDF1wnd865V6E1hxImU
xljapbSYi2IVdcSytreNUlrdPcx3ldshIPyo2w7mMy+OQAylUKu9s8L7hmxexg9/EOWfe+F+HO2A
G9x1bkLfiyiotxqOeQLYQ+/VQbVcSDmNyHy624kRVRAjJa3+x4whOKDCvd72/HmNX3o2SP3YaBAp
JdV0SjqQwHST4dMJZI1eW7a1qplXY6+BLFL8s9eCmXZmAvVAaa3DdrMtjSGfS5FxfwfyrHr4/BiY
3qGF0hv+gsFBNKb0srlbeSIXQ4sNkvHHzvF2SaaqL3uivKA0dMLjEwvxqwMxpSNjITBpUK9IXC29
c21KyikbO85wAXG0rm1M30yvV8AZqI4mVIBxVz5ysc0nbJRX1lQva7CFaqMDjcFG5uW7s1K5gAYW
7knSeFBMGeK29QpbM8O0C0hyHhEtrpuBqqLDVIuA0Q5/UlSBlUw3GK6LVkb1eG/n+Wcp5xywgBrs
EBUt8Fm30G4DKtMYCwqMx9xIWWAWDZtXjocq2pFmvEySqDjDErmjALeY9ltdEYnOpL28GVbeuxGN
3pA2qGHcF64nVngABUP/xWnNckbzoAXqTjWHEXJA9Owq961qGWvBv7V5CN+7iSbRU/XS3SOWmloc
mtRTAirKVaAPgifdvP7jI4FC6ckwHl4XKpuy0lgzehFuMdhSHd/4S9ZEE13c/TVZ+n4HHG0tZP/x
RgUZzlIdt/ItR6/RDRW+6k9EfMmZh8MHLi20T0KARQ//uCcXTkcBPrkHeouQQqnBaO1OgYaW98QF
XnMiudzLkqdFlLjkAQ7nE2rbFG9huJEj4GUG6iw56UaCEWsCqXNdlBgJ8LdCyDr1vkY1Izralt3M
NlhlNO88krXgN9FpA8KPjCLNumpCkeTj2LlrkeKlnMVaSDS4oWKbKtkYVGYW/Rj952i4dPHv6kCd
nSkM30CZJh4UBoRqDo1eeMoX24wcFuEZaKw2c8sMEvN9id6IEsqL9ep6jUiIZO55ejKCUXpByVGx
wTqE/kJ62D8wYb4+2L47HYgGA1/4TH3SSgo8R4Isd5C2Aw7kTj4277nLIM9OL3MgY6KBecpuuW79
xMzYggIJQKItRsHTdaWCv/syJTSttZPt6jEC3vNwJ8IbcpdB4hhy24p4z5nXmh+/5b/bGk/WQHKA
k/mfIKg5Vg2zatFFtrofvIzP2+2wF2bNYETkFaYAjttSgSH1vT10TYhCLW+NTv+47D8teQpTe3LH
/cu9e/5yoMFB+70ZntSBterGDlyK2OTodB7M/wzRq3ZfbenxbqriZpLn8MXlhPetdH+DFGBtYLtm
oZ7ZXEQ1vD5sK785WH1aAgseuQCTgD/fJ8cvgXbasMLUSHnuCU3qnKZZpw4AeI9x1c+9bnFaXvOY
sjRgGzfYVjoNhpDBeNeW1JoI9BcGZpRgo8PZn68l+EcOorrCh7dVo8lU27uljOvP/mRbnVtPbuUQ
1plmspZqkTMxVoGuSJQINXO2uC7ewXVzwN+egxZ8Sat/gS7STeZ9w99GcXWnIzYUQ7VuCIcibdi9
KP1N6xoUt5lz3wCBF+xuk1hfDOGDpkfX+l/f1S+pufhqy8+9wFNguAJzTUtQgoi0Ga9L+85bwsEB
URbqyIq77x8+poKLTjccKT4wfu4q75jdHKEJy7ap8XnOWVkXumTbaB0sWmkYR6uQ5RNPNe7g0pLP
z6ShnJnNKv8mlWsq9+dDz3ii5vfY/58gnR8QSv+klzvTNDU8FLBksr54ftOAfEjKluxZ6nUKtZ9C
3OSQCg/OKTz0OLIsCvuxtu72gbnP7Tg2zXuoS27XdnaoS8WTxOG6EdMqshXa+kQ9yKh62Rs8m1FV
6EIua9CMc4Ht31s/KhXAfYemgUwS1laulTJY+r5wYg8tCkaIgyTKeod8KorczWpKAp/gyIp9EJcO
Zjyb8hlLpRcEGKgrsv3XOoeGfrjBSMT+kJkehWgrudng730BPTqOmDyRFK85eD9H0i0/czyi4ABm
IpzSY8ECSWOc4xMKXfWtPoLIRsNwNeBuX7VuIG4HH026rdvmZknfLRMaWnbhcDl1qMry4SdNw4vr
vVqUgb1R+su9Rb4gO00sktd8vDELwFosbz6Qfey/qe5KS5+0J5yEp0TYXME+T731OpsvRd1/yW2I
o1hQtq69+RyVHaUEWsFm4PLdWYFg7qiez/EOFTE9QevB0pAVLAD/Qe7lwxEM4H8az6c6LB34Nh2h
4k/SiOW1R938asrZC2RxwKtSLOT5+ROTSm+R5rj1N7frDOQeDsDnNSY3jP27/1Y4vSQkhmbeOEiI
OSdpUltZhPPzKc+or4udXgFHfbBy6L5FJO27WengLSajjhURc13BAhL0pOdEFB22ztIHpSbPTQWZ
HM8iRzvV/Hed4l3Eex+WKZeuaCrTYff4Mjt6qgZftK054JLUxjUEn/ox0/UArifzqk97pK6P7JsC
n2jvq0+oHLqwOsX5kaBfga4nNTZV7GwJJowFcFtb6CHBuQHTCNx6fcfxJfzi/641mu4iQaDQxloT
mmkuDB57SlApd/ez7Ydn9hZJOHB0io1ukz7eZoMypDQCg99KxNDljIym85maGWYMtVp1qSi8/IpV
9g6z5yPBUnh7dA/WIrTknhld1hVr2+Y4NFM2iNDYr8j14ECXavRF86KhA6hPkMdDxUoPaYCqYdlA
jkp2h2ZqXFREVl7azxoUB5rJ52Te31RtnuEBPhlBHDHxI9foKnBGAC1zJOCPVbSRgCvGoAMMZ0kh
tX8k5AKnJ3HNgJgiXS9AoC9bjwAE4ZJCAlKECZRDLB0nXPMF4cvgpqY+8QOKbXCoVh+p6wQ9jdd9
sszICM2xm57+tloC43GCg5dj2vWRsMXISI8+j5eSNUn/veWByc/BoXROkvA7Fi5UcjRSSE7zCdm4
2oasEYJhQJ5fWgyOCrQSOQaPGo9BaGUUSbD18kjKOQQLrDdP8PHC8dMJc29aHCqhKuakuQ6d1e/b
PXsG1anq8zflaQ3YOCYRxxFJm24kFKJSKwT8OwRexkURQhLDravLXyxHaGbvLSkqWGTe6VOBiFlF
2pUncaDsyOzxopYIhwuAH4J0OsWMhKF8La2nNIoAlIClA9xkGPR298majQm2+O3HwvZYMZ/6hOKY
d5BkMOAFl6E0aAKWRodvUTJhEHxG9mvR/ICy0YkE1vYXb4R+Ss9xk+W9aX3K24Eaw1mMaQXOmzKF
pfs5LW5FtoBO03gxtZ956hkclVeE0VlLspBOVyUZZ3Uv+CDmSoiOZbwJQ8QwqZyGsOSGj9qc34nm
yUECg+4TMXqzcK9DdL3k5QwJytuMxE+shfE781MVoqoaeW0tNw0MUPPDYBBn+TSS3nHnA3dcMWA/
qTKjWfVyvRBdJ75LyMfhO5g1ghjea1LdtXmThweatjLHWOa6qBJ9Dw78Gzqj8hKjEyGBFl50NC4v
bykqL8QuG/aZZhTgu8FGEdBl0XQFhVEaTok1yHxaR18DhgYcoPLSBmY6Q4tyNxFRS/uk0CkSJ3TS
VEBaWPJrTk3+RDO/u0mUCTUgtIjX6eG1KHWQx6DB22KTyZdk3sTpc7l77F8/vRgzUvOfk6yew2QK
6ci0DvorvlNk/8FgmalMF5lVedkiS+hfQ/JUBAySbzaZzq9H23xoKjv9I/l5Rpv7AEPse/ojViNd
BdJPdAl9hOkCPUMxopB4XEPM6Ci411R1WqO9QazesPG8MEkeLTYH/6AJj+En9qUOqUyoaHs/6HAk
BR4gQZPGaqlWZr2oGZlFK+HxClbUgKe6lCkVakIXmVb7AONknIOpv4MuBxtMw6mCk+WOzwvHE9YH
3Onyfx5DRJz6jK08mYAILLu8aEnMWqN/gXO2Y6MspsurlAqwLA2BjtQ37e9MFPonUhYVs2kTnSkr
sP9e1s4fgamauMe2dDpJrfIzSjxzGjoI3nPfzDYAuNVX/oa+dnPkykMvNDRH2jajni+mhASG2SL4
sx8PZA7iWGtQELlhn1j8ZBijIg646SDflFHsFu02hpnwHh7LxId+wc9VkHsvT+wjBMUgu78WEzdl
QVEL98u1tx7AkVFVgf1iQnvOOU+nshKukmCh9ZULyNhqQ1yG2TPJre4IlC8xOnLoWdj3O4II0EjA
LBso/chaY21F1Ska9wp8AyxIwnlZ/+XKExR0+kxN7Z/b4ixLhpvLqMBJx3rDrADyH8wSo/nzMN+f
P8veayEsiKNuW2W41kPrVA5Y5adOoN0WPxSn9z480gGHsR7RU/E9lMbn39EtqItk5qVJ2ocEqffC
ejPK23S0vMliR5JzfnYF8LP0ERfWneyHtKloj5KRWGa8XKae4ZeKkrVi0khkGs3zbLFHOwrgVKQg
6kp3oaOjaOWPdhxCw6aeWtT3uejoi7pPYZKelr4WDncyRI7YUA5mBOI8frgaIYgen9XIK4eNWNcq
bJDJ0hKXBxvujKiJVB0UmT/3D44YLKkRy3Cf+8+glVPJNa5YN0VgpyXHnqtAavQ7mTQnsp/5ZI+T
ghJqIpR5QpghHhF8S7m7DNiOVeryUyWZUSVmpu7uuaRFj2CTj9RcG02Hijv7gqoeTj9MiWMyqck+
KBUUw+XY/onwC02N+MHBWrgN8WyKb3NDfSPsr0Zq7Veyf+DXaXuN7SJBq9XDnZ2R8wfphtsXDgXH
p0HXhcfalXREptQzCZ9ubv3Dvx8peb1fs+LXhqPQ4F8JFFVui7zXhXx93SX2j/IkxZ1Uh72hqF5K
ZqJOzp4CgLtsV+uYWV0J5K4RhTi/bfITHZqjJycqmGRtjk5Gec9FJupYV48FV7SALxB5P+Jg9mm6
5a9783Zo7+BfA3sk7HwaSzloo7ULZW334HyV+AvCAUTntPLst/eOlpzf4ce8TQ/G5Yn7Mm4yHimQ
3nUALqGDKu/yrWlhdxVWqjjkq5uY/tvQ+4DmQ4zFTKBWDGt1CxYX3VMjjysg/r26KbXWM0nq2rKE
CPBGPEbsVM82OHxTGwoXDyQPINwIM9ZVyKdW29vvg4tX6pR/Kwljhu3sftgx6ooXZKc0VdmyRlQQ
HNTqYIz7B7ubsdbBAHvnGV656HOicwkhZoQpmHzE1zLVTABnjRhlYql6kJvl1DzvEOBkb3EquQNJ
FZzvCqfmGVP2BMxoIjaS5f7Bx0ozrcfW+SmUIKMpt9iZlquaK3EXgLGeiG0lEQUH0IhT/3K8ffQu
e3GtMd7BGOazdk6bKRC7yO6+4OjGSDosEAQ7pFOMIwaGS7Ws3XeXSFz5Ei/XqnegAQlnuEIg6NSp
4F89RwbwngWqTFkYGjHNiuqlvYXBXumjslKqJaazBmFJbfqkaXyuuNc+Guq32Kr3zj6iZvptDN20
+5YSGKkM/ad6dof6cORyX4RMIzq5LiX+UVZQa6Vo702aEDE7NokbNQKTV4I/QgG9yfB52jYcSJkZ
ZUnwMKy6FdsbXf9FUaRc3uZAcgKvxtNGgSJKRkgEdsvvJMGRr3uXnZI2k79CBLGU9Wf4LE1Hhg5Y
V4uMMso47u6Bs7FwuZDGjZnJeXSjkj9fc2nNAq38NY9SxnO6JPaxfbXKY5ndHTvdagvnxyF/Osoi
2WbmkFO9dDsZ6+roXtoo6yAq4FzGaxCIHXfBA+6p/aZP8tAwMbRjts9G6iV9M0HwqZVInznZv/wO
L9CpheBLkoiAj00jFegXoAUFgxzGzLcveitGDpiSmbaNb7vARvFyjSrzEYhCcv1zCtEzza5++O/v
0H8Oats7K1qBKFlhuf+VdCcrIsMbac+atXjZI6QRYe58dH1eIny8zs5zGqCqlKhds8UokG38LwXY
Ol3v20Kjn+OaqkAKQhE8nJ3O2jHw9msJhqwUPFSwF2uy/erVbZpfw1wnlYePffljh92bwgwSsiT5
B/EEfsgCAFixsvylMQVp8SvTYuj+gP7oI6cpaVChYvrBOys0S7YQYSty3Sj+bAmV2Ye6NKB3JHtA
dLjjZw9VEoAErMjBInHTBIpSeJoESFlPibclU5WGcpsdSrYEEW7eiz7HEUkev2GfsfYYhRVNK2d3
/Q5p8/HJMnL2SwpqpM/79blDt37Yd6NUocxnlLwaKbZ4MLfD4JwaUkj2jkL1vF6SP2DQsejOfLRB
Qamqiwgz8IgH+ZyZ3qqXPkuJaH+w6hV8T03BDXTFshhPc3yUfpR489vqCBjevsVQBphjdWpEplSQ
odQluJEqmTHI0b7NDB5e/RonQsezpZTjCKd4KQW2zxQuVroCB0A29xHXvUVKOrRg0X5pQyZqUNjN
fSqsVsND+qZ2yK8uxg+sjmNCMQwEKOTmzP0hY78v53JUkosFXAnLyG+OMzFhywMnb9CAZ/uSPFOi
yig+5zcEzOApaHG3KF+IBFHCgdFc36srcJAF4t+0cw0PXnqeUx/N1Ve0LK8wfmsOVddrxeTeck6e
XO9rZJZrb8IHLu8JvqkhpulO/7feQpx1SAKuXb2VqY7Uv1fMpsge29o6tx9znnON9Hofc2NQFOkx
/G6jVpOB7ZG8bK5CgVQx3QrZxhe92J03xOsjsQeQhN39AfhZQ//O2klMd4EF/0QPwg+WvpFIZE+r
sGwoEXoz5bX2qmHcTGv3PJA1z6W4vyHVtApSx3PX6QaxDLnjLfHQNiY0jKSVLNbTHfKEyGzR32NZ
jmKuFpa79GSFxn+IV0E4JxB59/7rmjoO5Ge1AUOzKBmNKMEGNlhHpBTWLwKW+ptAKz3jCcQgmG/d
KVuVJ0nGu7yUWnTgoOJ98jsqduKptIvWZ1xJYcLGuOO3rjuFeq0+g85wImYJqY2wHzJqBijNXfRp
E4J9inXAt9P2Y7ktg8ZYGY9p3v93SN5l8ba2yeC6Wnx85LZS+7p/5PQCTPP5eG256VPoV3U32z7s
ZnkKDJfk3MOC+f1/vwKUFlsGGo/9yj+dF5fr4s/29GC6tHvg1a7xqhJCgftGhsYWMOCrehigX0bl
s21cPQe7eFXX2l+5boAvMFP0XQpAGBnR616/fljLxHJrLDunzBuXNX3t/4d+fYo9hmid9+VYpaMa
C4K+1rKlNOIqncHoaQc/4fr3pzgAQXHHh4VxIdcRBS6cVtHhmrh/VHF4a65oMAvYGsGxsiFDPCV6
eyr0VEWBkyQRqJTern55v1LL7RCGaur56zA6yDOr9wbD8q/e8k3dyYeI3nFCrY95CVTd8ihL6U6E
3GjZUArjUKvr7Sv1X2l+mXelteKflG19/YrWRgjXstR7opoi9AIcwY/M0yM1AWosSqJaHp+qJ4eb
UFYRiVVJMtG+drNFI/FRwn5UNMdn6HCJul6CayvGe6F/Z8laY5g/CTh8Iw0fH8AQXlyP/XD9u4vy
ScZM0PIyST/R7jropWdwfxW2vtPWrzn+9iiEEtoE5AfLK8JauEgmV1Bx7wa7hZD+ZeVqURBMq/0F
s3LNvnDtOmt5+tR1Xss1djOPO29Mj1/va774JjU5sE417tB0Smz3fRca+ZIM22ZAY8JnwuTYoOw6
DL/PBSZjuvXuuHO1HCDo+BoWUKA/PRsN4dm/hxcbQ1PEb6QdiUEZ/QfHNtHizQxPyKycfLLxD5Nu
cO163xh3gzmMH5aDHBqoyoxLxZD84dcH6ylMN9TZPO2ShJMcpa+BoRqX3Edi8FqzOY3rJSd2I0tD
CEZNXGxUMrpbTcviIeEiwWWBuFCFePe7pCp/nJw5Lo67S62IWh5IOWfK0iIdQeySqK5V5WJNzrgC
A/4ZBzoD95CyDAAGb2xwpMCYxOPE3vklKskS4HfElRqdbyPhVoy4Nlqs8XhN8evGQb+EBjYpt77f
3H3UNEpv2whvA/9A7R7HqkFNkf4S+7mcjfLZ6+asyyU19cbuD/ICQyqojrYdFejs1X2TZh69T5z7
wrTHsQFMf58lEQm9Vg8bTJS2mgMG8u4sCgMQpH3vA9VgjdBUJrjpqXMtBj6fEr8KRrif7YXW2M3F
wUIpFDerXDA1f2KsfZtd2ssBxV+DUt0v2xjfYBPHH6q1dL3eB2UlXF829F0BjMtxOK1w6xXqtsbM
DaO9ULNBZg3LXgL19fnY4nV9eqMSh0+alCI1nMkPr8y0Jq3xA7e+wJdbsMhMuOWFzKtPUACA5SdH
MvPOio7MoDeXhrTbaXjdWTFj/8ZIlodMgwtJn3pBnaV9d8mR7ax7VHSHHbuEaXbMTUiMevKZHTcO
FHCmLz3BtZCRW8lTXCDxf/p6U1Yq5pjw6u+v+mDqV4XzwwqPnegnA+xsU5RwzxO+oEU5dSMbpU94
I7oEgZUcaDa/thfTMriboX290yfVTiqh3iH5RL7kLok83z21Qyg1BvWWoU9iyBeBGzgMqSOtSEuL
GwOajiQxfLd0o+wWFwrPMw8LHj9s6VF/+fMA8Of4xDHmPzkupyobQ9EX5ipo6a1UTRjb6AjwcyYA
OOjSV934PuUlDozYFU3IdzUViyBOjhOHQIs/AJOAoD0WHQ1jMOxKWfbFr9JK6CToDO294vDjgQp/
cAK1vLo8414BK8lCPmPT7X0tUHsePMJkdxVSCV2M4++19FBcu742HKYVRqx3j2kkR98Oncz8nPrp
woPqfmHAZUN/oaKlvzq0pUWRG5EbIVg+kLHJKP6Shwp3tHyzkaHvXDpfxRBGNzXlAg+ZIdx6x9Gk
ZDOeLVlYWjw6RiDAmWA9ZafAEXdzrXlJNBOAMcyQV7GCFRALLEoal493rULOnsqcmTXrMZY2VlrB
xT7LDsFdKe3jLc8BLkcxZ5emPDOLBjZTld0XA9YL55r63mPy4qnhVOEeo68W3fFOvN0xWcwYjUn9
5tG+uPd/g5+ao1lUu29yxtLIeAY8UrZW5goC0/V43or8Sz7Mc50KQYdOFkLGxDe+/ciOjwo1YT8j
MIocFCf601c4Mh54RJThIKEU9QaQSB+dkMQn9ROgsUYqzzKhODEK9qLCip7fEw54+mulvFPzd9lc
b1yp9BRt6XjgpgIvCAUPFIxXHhuWAjHFjhramfv+K0qFMxUbMu5PSNWdASVm+gj37wHgdkc3sqTd
gFx9zJ4wJ2ohPnO4efvXnkqj5dDcJv/Fi3o1do6COCFBXPn0hUoyhBtUwj3YQhurB1zovgyhk/R4
Kn+/TSYHAO158pp1se0PMndVt0SCAJ/U8UjKgrZDXHXC/rNtUbVozqvRwOQvGEVr3t3tr1i6NimN
VWGBn3D6ptQoeP2ouT4zrXjAQFoobxywFgccSXmZ/hD5ri7uPO5mZa09Q0+L8UopAagigvnCRbHG
FTw47AaLYgcFj/vPmJL+AmksGRkvWHV87r/MyfNljmPvjljcIOXvdfypmP0jtxTiU3nMqEK8Cx2g
8WUrZNuH8H2pBbh4y7y3OaZGkoLpDXwlzlgd0ZEGeVFXtreVVo+nP/N5UoUElx7jqfqRPSaEDu0l
VlWQFCua5e+rEqixCC+Gl+ADt9eD6k6TciD3R11H3LfZTIzKWx2srSU+0vwMiF2iUbIioYULBsWo
jUI4T4x+WeHIpLX0VS//aWeFEVMC/e3qGNDgYphPMGvLDftmipifikQDfyB2KTyAc9IK0XAe9cPS
X3OcxYcC9pLADr1/JIBYk7GAoXH9n656uBl/hxdfXY+4fxunarEJ/I0aoY5CZYRf6NNFUjlLdLqS
/TZVbu5w9ab588HJmV4jVkBID2a9MSDzfFeSkpVq2zSxgFq0tZyiPwtnKRqVnacpbb209PrNg/VT
t4KWbn1CL2vtaj9T6uyQbIZ8KSA2DfKcwMD5JfYMM5p+m6XSdX3pi3vp4h+bD9r592MYbucklrUQ
JOu3bmK9H95UMPcBLBPA012xkK1zh0yXc0TbOMtQ5ADBfFjAftxfhUbv0fMk8ixlqoiBufNSOMvt
CktY+d8rd3XBrUHFY81EOZgrSU233w9jV6619VQ8aAPtBDwu6lM//DTcohZSsvV0VhqdFXlbgABx
Qn6anhuDJL99RRBnEXQjleP/eXgYqBJgDnRD1rHmgIBu3M/BdC4NwSfQLDa5SRL7kvkScltHLlyZ
RlbiUJsAR8x1bRAA9XiIuVIDhVvbvPDlg4bCD6PPBi2rwD6/AeOjmH6oJH2Z36uERW6xLUOHfWw1
HezDv4lH0rNTJx2tfrdnJ52IRS3uveFuj1VO5DoD5vInoBNMrYSIkqEtMghW04wFU7RWjFfkDqPA
GSIpkSluK8nQtuideSSG6UJ4jVUO/rOURtj8O//0nP+I2Cl94xoC7W4U13MM5+GE5RH0cDDONK38
XJYIC6lJXL2RPQAFq9xxvnm+TsL6Y63qGHsH6y/izb0lgRWhJtpjuuswih8rPf0OWBFUYaX6nNVH
0NLf/4IWTS4nllFq4b488GIWrX3rJ47MGomM1VVOSH38YEBbfFgDLn1bKtamB9pCLy5njUtkm+3L
oQjXffMUNXBHotkrYncDvhAZ1n1guUExu1cV3Yug1rT2iXyQWxxCeE4Mc77YLD78/Slb2GEaDVRt
xebksUyvoEH4+DkL1Cpq/vCMszg3/6ImzzZ7xqFLcWg2OgVfLKnL3BbfcMbCCfSB1vUGG0/NkyBV
Y1d4GtxTT3GJ87EenP/EPOXoU0hxCKcaAVEU2qpZmi+eLD+VMX7rPlEg2va6+0fE5jgrgN1pPOCj
bJvZrBgD8lrbN8BMXDu3ml5uh0KaHRRZkS3eM+X/1jO1vdtJLmN4BSsfMRry5xCIkSVHZIqqdXSF
YAli6OA8YWQG9Fl7TqhsRJtrjirJJ1UX9S5cNpLM22GIw9R3ed8p+6F/CTpMAlBwsvsGb91IX1Ys
inNtNJWEJ2RzJX+D4xgHcwikO45qKwG/yDXI5fGxU87jheh41CxjKnZtR5yeo8xOnzvSIroODPY6
grKXT6A3Zhn+t7F9UKruPHc0j6vY89ye8o5HNJ6tNhsw+U5Ns3YnEs8SId9ASgkD6AgVJFJTGHqL
A8B2GI6zwMFHIakIzuC+P/3ZcOBDTUcoRcIE29ceIKT2wTF8Ey9Z4Lcuqq5WMZ3bimuEnPoP00xL
+VP1juGeo/R8i60OZZje7HAmuNGmmufeeunOn+uhU053RZlSeMd5MMrKU4ghwEYkk/7QQRXNk1y2
fwGCWQ72AvCT4LklisNpwWPN8c/N6wHHyHZCUzBq3N3YUZCwpW04iTORDFotGBC4kT8zz/zr/zPo
qT2esSS+xZvaZ8HI0ATJr+4uyf43PeZcFR84xNLRwhsaqNeURJF+Xp53WxjmqbNMqGG7MoD2a0Hz
SV6Gi0dx2jyP2+suv12n2edDCnjcC3eqS30AoPlyIZwyX897QCnxQ79qQUzyj86Vhiee2bJn/4rX
KR0ThyUoGq4WUrhKzj53rjZ89GU5ahmMwzktFKYH13ckNUWySFV3YyMbikSiyX43mG14Eg+WY8PO
uzqZiJDSfGnR616VAnq8JOKCwov+NRTSuBKl6y2zFaUgnPI7jGRUi8GQhXmFspjtUTFwWw+BJrwY
R7eIsW0tK1QbdHm0ZnwQDt5yRZldt8bZ9Fr3k09y1no0DbNXN2s6nu/M3TDn67Zf1T2lWliDaeWl
rBNRmGGdqE6PXMCzivEW/NB2ohqFz84s/mHhDo2iwAAvwNZAgc6f90ZBJijL3VBlfVE9A1qq+Avb
d0vX2YYWCyaXmJxzGl3Fqiv55bs8dRFWsvY5rhPUcm7dbYYpNzbCE3zr620/LVa9keAx8dms8IHl
cDqUEkwv84j7g1xBIRVU98YeEgghgka/fpWa/vyMdmlvKvpuZhLd8EQrl4Y5RqVzogd1HL34dzFS
S8eHuuwv3XD46+ILGkWJ1h8QBItFu6fm0jndVnGqM4wEKnmcOD3dLX4zlNRWM2iINEoBoPR40w3A
Jwf4YLDAhaccRbuPGH2Vq5LewgN77n5y/3eJiX0tp+xtKyxLYR05AchI1xq+QaGqiUgKyGJz5tPv
SAHKXzPoTcrw1YpSvaO3UbSKKKDzYMPRz7pD9S/KApTsgYOIAOnaXFeRgxEMVQIjCGPNgw27nE7u
Md7r6gnvB0p5jP6IR8XvG0RlmpYD1D1aikacjSb3PrZr9UC+dJxLWIQffyFRl48iO8zbpLMP4Kde
3MV2T9JCe7givoDlyVstZud82x2BMM1UeyO/9fg22v0EcZ315y25O5FDJ7jOuKP6tOE66B1yQjAx
DgyZ9I+3p2U8+hF/3y8YoLCKE+gIMhMc1Ju+QRNaSq4zlf3mlJNcU/hhU3T2DWKfDY2/sVyLD9Pj
dSFhgLFksMMVvh590VZF4VsavPIidlUrTt/meqob/ULjpxb24yaVzb/AL84bikkKC0lG/dAzkMCT
hpUfzWqP3B2FjRG1OWMYHDtfprUuv8ESW5882VERQWRUNZhc0Nc6gbGBi7O889VBv4I+bl2S+mMx
WwCSu9FjMrrpLnMR9qdWZhPOHRwjnsMwudfs2SIXyHdc144QK6bw2Ec1pmpnbT96AYBRyxsCqi1v
f0yjrd4VMy/A5ibMPY+Ab63PzbGOaPA5qp00w1QD8oGnswncLiJQcRJpXY0BIYNx2WYWvYvi+C4z
OdEAku/pbwLJKGbamjhNKGN6Gd2hPKo+aDRbWl4A42VU9ekeZsV9mrMRfzlihuUfMZfCZVNXkTfI
Upw4DU30ME94qxn7xqxfuVegcVLFJ1Y/8AUmJhsg0nK8dTm0DNGjlVbau4m14PFylZohSgD/hila
/EC6jwZKpoCm2U+EorjWQP8iHw9ZM8tHdSk0GGk4cTwiaxMhImYMpxxPzpqswUv48p6NwbqOVyhs
/3z7KRzAvDS98VKkb2SGBTTs+qbMTwZ2zkZ1TXbchgBa/aXKz88lFqejYLMxuG97JoLaOqxRoR68
xGQY2sNzFM6lXapW0/3Ov1a8lCwHgvxIIQE4PwLQDMx8lLAywWTsWgliXcdb89V72ZLI8kS517h+
9jNAKeNMyjnZmQfxcrJ6/jzPFQOQ1MkKVSn3E3Sy3UizMOjLQyy4rgs4QY80cjmPhaBokOuvS6OI
y+jA9fqeSrfKh2m7bTBTgdBxoAPuU5aUxLZ3Mstko4Y/y4xkr+vTcpNs1f5j/3UYHcCAmVOP4+KH
ibOGorlus0WOxAEz4KHjugpzc4YP0gbZExAdVdpF5Qw+AMSuJDokrE2dv2+0Nz/qy8lMuJYLuVnC
Q18Hhz/yPcXjB0S/xtXdFlWuyJ+BQ9CZWModCgazUBa+LKp3AYtoWdlCM9uyctV8Ibpt7bWLY8gM
+JBqKj9PUBnB+VtKcvY3kf7FXQEZpwT7oAxu9COVtOlFUY/jpCM4YTeZGKKYZhRxS/1jz2kc3osW
DAlrmvv+0uAKNugGyCWc4DO0bdsK+zb1EEvnCDz6yAMhtabKySu05xKZLN/b+7yYeJUnCndQeWRJ
k1AMoLh/KoMuZLwjDfmMONmx7NwgoamXQeysKBVF1ze4Y69K/Oltf7Jvm/oDOxnfolL/1TKRdED8
Suj0Vxtxlx0AUjkV1OSqRdFuBsUYQig1Ew/TkmygFV0NtCHtny0yzsWrQhWnB3fxwNU+XhAm1+Mz
8o3qMSJc2Q2N1MCVaPDNTQUlGFMEY95rsRvNcHQKr8BXlsIYAcxdXdg/5Pzd1PXPqxe2YomyZA2L
daivJWosbHwa5ZZ4oUtKgmcF6TW/12HOmTpj8pWq6uRsTokQB436E3/KUZigIrGpS4a6/o9GGPrM
NY0f5mTfrmQUD3NTBzY3TXzwwDUsKN7SPsxL4m5dPWMOFwX4YPOKkj52ImeV6ntUC4G91Z5HTlF9
o/Hbjel/tkT3xIo+vqJsyx7MvjKXeCOtlBPUV81h8OH89D/UVC8PWSd16suAddr0OrI/dE+J084D
EaxLMjzTY0c9vihplN6cEtftUVomTsOuZwDyLZrrcsIPlh5vAN5bTXcWitLy05Am77rAJobXuU30
7GMwVKcabD44nORNbTsXjgBtrFoeOfSf5ASf3Wq/bgVSzfQkHlBE8i8KwwxThoVEieFefc/bDVv3
TSlskPRsCjs3xxT9FCml9acDZ7/LHdVZtEUq5A5H9OYALEpT05HGE6p0dCenvVQdgTWXFNxMfIfz
J/+xZZSIqFsbI/B+Z6WiAJEaX6pu+6BtWgBZRrtHxKf4fcD3wLKRuY8OL2Mdsub8p4seI5LMpD3L
gLZZCvd22NmY6//9Uu5l+3XN9fOerFYIfmdcZYanr0qE9p14Dfg9NbJQcaSMRl/tV8Ug8TOM7wfq
57cBWp6eZdPRbO3ZzzVk8oC8l1+J2EOs6qm4eX5EKpb8ll/J4wqrMYLLpVBOZBa38WqeWiwyJv/P
y1ed2ljnVVxwN2VUYl3COZkdjBNWVUa4M6WCJYoJWypcdcIoGrJ6MNiHEINTsGqAENWfQ6ARI3q8
LfVu7UIZ4CjuzxRNkPNBYfnm2RLi94C8vuO5wU3eQkmZKhk4MvMb4zB+qwfwBFcPCEKljAzYxGp8
vHXvzCWNlDpf4D8o2QpbKosz3xxldE56zE6u2Qtzj+FhZK4hJBBMbbqJrntQ7oo8zYV2e4xlSRdN
fwrU2u8ix51u3MMohWJ2NYPaC7gjlIeL5DxyskdUYZs6gMclY7Lp6dS9Av9lBzCW58j+Z2ZFJ25d
iOO3CRovIvAbTfgObf6c08cT4wemVC0RqQT+NTEG2Yst86F57LnvodZgdGscdKfC3O0r9stzqNhe
JRVs6p7uw+kgwnBGA6rBEnwebmmEfOS0haKYy74O4d+VE3xKtdHJ+3MaG7aqt1ojSEr4hQ4GCeT4
kwfRK+AAZVTzP47O2Vr+sx2y+ERuzST4H7RZ520Nn49sbg3+Eg0KuKwXxagpYG5gxAOENTQ43WQc
9//sB96npS502PAcRmsHjy1ZXr2CggioXLkr5KuHuFPlq+yWALqZcNuVKzGpKGgT33VVi3oiR4yP
DyNvfUFiXZuyg8Wc+m+M5ueFf7On8uAQMC6QycXeF0H3lH0rtyYBxDShWvN4IEf4Uz0/RA3isAmL
UZStKwX72cRGOtz+og+PUGcXUE5Fx17drZ9uDsffFzydkcXIFu9vWxbjq/WAIYrZ0YPD9+1b2lPB
7nSr7oPmobuCVT50NX8D12aU5Ts+YqJDNc/oDn0Rd0REYsQW/B6P7K26gLA/IuG1HXq+pL/h5FM8
dRq+N5LtmP5vuYbYgwYjUl/iA4zxoswdse040XkJFLrM7c3MOz3EY04uK1acf59iNdfX3xNTkcUA
tkwyaDlGqsaZ0o9MnohlrXjbjY9T2CfeGedArcVRG65kV93QxY4XXvNTQzOffjJtJVFOtZIALXuj
dXD8a5cp9mijHmWihYLPOd3XnTa3QP5bchmmFNQeUHtkhNUT7/ztvNddlhM8A7Xhz/HVIRACEqXQ
myu7b1hrlZ9+mNl2//hZYzv5DmNLrE0pEslYocQXEOL5EPHXkFvPoW/kB5ZRfnvd6fxoOdwtVrxE
BUqJ3uE4yjYugCyLoz5yyBECRyrINYce7PHm6XfjlR4rPm5JSHzEQZKF3uHGrShFAC0+2PA9P1eu
61hKAZfqhzSWUedh5FUPKuApo6RkgMAsOtjd3TwgRuaAi8xABq1wyy9pDXhxW+fia6w3qmQG2KQ6
tZc/kzIr0enEJsHNa5wereFZHPBlUgNkEzvKRmPpeVnQTj1hcQ0gqQWKygNyyYw8hMOfpJJF2asp
BQ/iSKZjVo1yHZrMgEPzTgUwdkAdmXpHGQ9adypd2IsBsGn5J6N/mLnNsOPSr2caP7yDX5jPDLsr
Kf034K7fExxo9O6bKAR5jdrK/LbjPTLbrRp2xuBj/aPutat48YAFMauX42PmhNr9XFqe5JRoY24D
XdmxVjaRdk+0vL3SO551YXGNBtQHnz/sn6KO+wZyBcvFGJI3mMN7nlGUcnVT5wgRlrgCIoeALAOc
TcwcoIOmKRZitPlFUrFxqi19yDwoarzEgIDw83wvcEbIeyBjTG6PhicIjaeH0h2J1JunPnHECCg8
W029o4oi+oG6/j8Sakhz3GiF9vdupPxWpWPIBnDvVhJjgu44jD6GeNo8qfc7lsvIombAIkIiaw9M
EKE6rNTSQLqqIsLd5L931dG38Mq3vqVmbuDFEVOuZTH4CYxgD+8Zv62347GQlWe/x28gFTuq3Xkg
CaBM1/Pa/pKT+rpXwoFTqaVBzuFBi39+1h2a2b6WrucC3X5jy0xiz7qVhRutb3jo5r7y0z6Nv9CG
U51QEzCZ9TNUx2Yl7rIMpOfQNctGMIeVFg64qUWWmwywWc4VjN69f0njeknh571v4cfTDqanvjzo
rOUPb7GNVosiAkplicUxFypZ4lqU6+X+A3rA5A+grmhXFo02n0TqA075MuVEAINHeDFUMyVW4qIB
kGvZ+G27HNPqSZiKcmtn8A2zrJjA+L/ow4Y7m72BjvR3cMHun4clQ6PEGRdkxmXVG64mawTgFm4l
4J4js6s4BniPs4h4ju4k2mZlfBCp/ppDL9+RFQa683lriVCtecXW37h0hg1t7A00ei4FSlYJBuzK
Jm9f0Sqc9iQW9YccdL9d+yXzIqZjW+BFk4Cj4i8bJFaebFdp8oxjmOmI/fxjw+8mA9tx8FSY7aXr
0etK2szryv4JAILxAr+4VZhN0QIRYL8gMqLDvsa29ZuIFXqJQ1Ul/X0vCw2zTE7pCcUAuFoLkKho
VQQ6+A/+22J95nMWUSFV5vl38XgKxqEb0j89p1fpai8Fz0FCq0kHJAPIVb/Ip80ErsdyEfvAl7Gg
a75/KD6QAADtjjluHLbIM0Sh5KR9cfxGR9i9uWhSbOotcOprr0+O8OMFyo5qw+Hj0BuvUhhpLejA
T03jyOm6zgT0iBYb0aLBuamb6hs0m7ajtGsVvJR9+OtdU4rIn2dw7YWmpLepB1QMQ340R6Dqv79S
fDXLXpR2Q5stiFZRJC/W3o5mxYwAlfmlkj1xSiNHcf1qthT/0TT+620ElatqGB7Q8W6Jal6pGyEh
LGE7QkHVdNJGz4Ks2HKtRYQyBJAfYp2fWZzgQZBk/YNaBajGF6G0fWWb0aJ0Zt56qbKm/xfHx2an
0KJj0T4EzyHgZnrNN5mH46arjY+N+ei5dmTlOk5QKV8fbjvEnObCo31sAUY36CF4KGDqcEkBM0WO
LuSlfiehGLQQXsoyayiDGUwvEXA6ux68st7V3vO1SZ6FDGm7ycVY+5XTWQzlBp1KcVHNtjValfd3
3VYS0O92YjvcYm/awt+wWM4av0Msi0SHi4cN105jCXGDiS7z5wd8tf9B5dxnhZwXkiFWiSx9N7wU
4xu+QQLp3Km/Rmc6pUGgh7iJwkQXgO8B+VBl+nohh1pLlWrjMy+NZBfHLAKmGS3Z37UPRv3A3t7w
8Y44LlBJxPthCzanqryr8T/n2UmbNobJP3sMox0VvDo/gHmb0J6oIReXXTtrSpJfoLK4V8CdDbFO
54nsanZOVI0vczBREFOmtY2xNKjD760q5eAWfn1GlOv3qOeiws60uAdpGNS5L6NVOGcBVKsgsPPc
RWcD8JbhNfHNcsGoXW66bfyZl5h+rNjXflaaQEWtLmRjr1OJwytp8DMSc6uQklAM2FaZvuSTkHpP
wWbeA8vJD4sCv2StafxBQRYF9S2u1Germ7SKV1C4MNnLW58LqA95RXPxhbYou7P5b+H1KpAW+DpP
myshBZnChaVzHrsMXw8HRg2eW6Svn0XIa/36X/b6ticS5vyK1t45cwmt+9YCuGf4IIjEJZlXM8sS
npqCFtmUii2g7+aWr9NIEHDCMaoiKwDCVMjgMlC73D30Vc7+4H4fLu879uu4NukESoLywnMB6qGI
KEaR3ljGc9MbiDQofX/ra9nuIOFgP0gyUzXiFUlkD7XuMpSsY9ewwfbeYhijOcjcmXgmslY93fL8
RMGlaYATZyy33cbQPLSTCV2EqcjOhU0CDLy3ZLFNSVrHL8x0FM4byldm/fUFAUtzvbVfme7HSo2h
9kWNTnGXgO/Xvn3c2h6AaVQHG1oS7a9dC6h3sRnEWAKgjvxKzlRJSnBgabn+5x/9gxraRcUbwkB5
DcpQYcoiRUe6tU/Cp/eHqtX1NEVLeEJQ2MnfqfZP6upXOIe2fi/FjgT0SlETAUuH6xdmFFTzbc1/
CRdBx7TjWGsXi6KWucwlPsASdWr8MNfppRgY1CTsnFehOzmBrTgd6RY/aLx8UNcbE5GIwgiB1ZS0
vhnRY8rjwXx00zAXDrH5arfOYZFt2ZZ3LWWhsaMPexzqUdxE2bChNKyQ30KVuIsJFiH2nAmEJ0Cy
UcqmNdna/LU2wia+jAukuacsfFRdQxS63n4cd9ibM19eUrXaD4AV85Qv5wjioFBKGshw2bQQlQ5B
2rRTIg5AJyZfVwWSYlmnyA9nIIQeCyRsvil4SAatUklL3ihSYBJ+SJ1Jm6ubWUukuJL1KfPYwwni
jHmLKYZXHeOZlIBz14X2VHnKCpjJ3R3NYTrW3iMxf53dQMYr5EfZ80V68zgBKChca5DhCFaXBkY/
J7hLDxk8DiulQqdKILLI1ifZLYQGIyP4mDc0Y1JuG9ETbpHvxvkS/yAYWOtOmEfk64I2f65KixRv
5v6hfcWleSjZCfr3x/vOAZqdImy3hcNtXjIKAjAypCegrja76ZtKwGVGmBRBdqtXlhl8dRuZ7XUd
SWKoYD5fLNvaJjOMVKAUXMaF+XzB4mEjCW4hNGHJToeafIqAAzndBsZCBxqZaM0lKi54nfmMY65x
gzCSwXTe4L/5pnl4EYgAuDJIaKBHm/5P6tou4EqjN/+yALLwtyFpi1Xz4ywKg25l6k/K7HrOSBJm
zh9CCYrVBJd5Z5+PuCESV+tiEVbctlcNR44CrWuJueSKpvBmBsj9XKrXMUq/i/HKHZNyssRdlKMl
TC3IHKJ9s9DTfQKHiiOEyJTD6zZkqn4ManH1TwKXSx8FHPYZgFIadbFH86SyfI40cKaTDT/Gcu3n
6xS5OtEOy+vqZr/5lB/77BNXH4RJXrlBrt677GE+I02yusbdSriAp8BQ2WkhxNL5VjdavlaowjoA
EWw1a7AgKt+FLxo7aUTgdD2xFddMcookam2c6FzoTHOqBkjRzxre/sItUqP61IwAroWj7fgnEs3r
dV4W6UQoUxPrUdm2kNEzsy/L2QI/z/jsUlZjOuxd4m2uqv+KnsHnNQOCSinXvdihDszy0PQQdcMZ
7g+ldQO8TMbcOl8rkMsnjyHoWOFXkrl+OErM6MKi0NYXPM5v7f+UZKmWFX8JQODJFO3rUtMavTV2
+b9oshVv2zbGSvS0N8hiTHd/gqDKpxv17VFFKGgFHFlBpD85Rq3bxR6F4ei8S+I/YbCsMsnVRJ/h
BslCVlFx1SizZbI5PHEW3yr62bIrN1WTTY35acA8wNErx8f1U+ZkW6cE20pOW56OngrfXFt/qgkm
gRb8sh9abg9xwHvDy8g1kHWZvqCup65MwAYeZWnsEP7SyFvBmKqrq+Jd/XuJR5+cWRIG62KIpalG
2LnDRnShnWjjwjMDhznyhld+4TaarlQlbE4X8qNmkpnY5OphX9XwArzoC6Q0PUqgsnc1D9WuMRXL
UDXr6ltgm3gQr1gtVxvXrgOnUJKaMF2ytSxb0/GtEHNcPwosPn6lsiET8ZBY5obRxOpbWrE6sFuy
Ob+cXHJWJ78xSzvd+ha5sPpwkge4os/QVmFGUxPpfqMLVj0IHm5WRNt/dHfJQ949ObRVsinztATJ
8p+rqcB3r1J84E3KsKKDc+yf3kG28mx73Z4BYeDe++xjMbpGi1RxsdNwH8XAKiyvgjjqXthTO2hK
EIZTrCjgxWmMYUIQ+ya5TOHa5QATos4IO29ewYWKV5csDYy9wLiuxjAMOkZ0DdloNpgpaDIX9kXF
1K4Ocw6RcVu58xlK9zub7D5z0/wUkuw+c9E6Cv3GUumbgyCp2JbEoJG0fLtgVsWS37TPodXwMRee
6YCXQUbd+vI8UntSS9ygr4x/nyILoA65/mAK3VeXB/lrBVBpIpnJWK+jBNuVFQ6f58l7UT+Wxs4a
U5w9wlHdFuowytde6cbzIVBWiRGm6PWN5E0yIxp93E/iS5Yf4W+UABzQbWLwFNPadcKRLhB7fv5z
Z6fsX0oK27QY0rCyVhGHxQI2F7oLFJNWrRKlL8gx+xyC1CE+lDNJJywn9pHI+CQ1N9YlZg1kASWb
aPC09YlQjJ4Z5/S8km7ctd8kwyc3J9zoUvtsIfN18EbCVZNXDR4SDG5p3p0WtEoNKt0LWfwOTwbB
PZ/6Wf8nR6YWDkZq6NdxMddHS/ry/5f8H382B632p4HFVn9KbX6dLtdHj5+EHbw1+tinzz7RkBlc
IBfDy7upPi8voicn7g6RHg1yKN+b+hDm6m1qHitZ6c/zHdiYaG21kcJwe2Nb5ZLEvmJKPmCG0jkx
LqIfAsl4Tir6OuvNw2WSdRRoK7lcHsv3RpSPDdS8V+4hxLT6zbwbphbxMTWlHvqf9fujqPIaqbsy
QtTjh+WTunKLgKqjAmAASNlIS+gqnI0dog4aZJJkfZXUFC7py/BEJWt/HeHpJE3sIGzdnpi5x+Wl
z6rdUMBFmyzuG22Pde1zvR41+xDw6DxOsia11zRAUXLlxkELQ4Zsa2+xMKonnBPuAD21uLpDhQ9T
/HqoijOdDxxewmoO/TILr5ay245MA3o0gTY9YI/gRzmfHZpDrpGmvu5cbVodkpcrvuL8Lx6uJHb2
CVzAruqGgmcBgUWYvrd5UhB70b0riEu/rZ8pL4/uunHDsH4nzCWykgOSW5culkPgMSu29V2RZ3la
f0XmWia7QDmz8HbWuPg8sBZ9uQxYK6iL359CD+Jql+CtZNio9LD2qiBsEex+4w4oBygIpLzD7/5u
2StDqT0cqr30MVMvLD4AmFHIDiUoUQyYnGcuj3yB/Co17wP5N6P3ThD113KesPudPcB7p/b/RpNH
OzwIyOw1FhS3LcwJTOnMdW9C6ujnjn4lHL0moVayw99JqpZk8poo2oKgv08ELD0Gk1y/CK7Jp7Ts
hozM5mUc8IUcEYo8NcMGRBGm5tPHuktywugDxZC20ueDLQZ4hIe20kk3Wspe2oM3xzGU83E+khpd
SDIi5JAvQfFT7xxUoXGbvOjF/TasOe4XxMc0v2bEYs1WZTuV96fhkUkALgZJpyAdb45zdSsVqjM/
Q4/EiuEeOmFhkcouXbhtyYq+P+DD1/ARHuMLKo3Te53X6Gk5QLwh819NDJn+d4B2XqA5oo+23Wyw
K5Xe7tG5ztvjCJC53UR3CiOVrjTWaBrKaqt4nO+f1yR6TDO0Ejnx0DcKnpmf0887cmmoMB808tEF
wlXkYCjgSVtmvtXAxkF5BDMcZOe8fEUW3puH/C5Fgxaw8aCjkZJUD71Xs3TiFKMHtQSoI5LnPd/0
M4brjp++jU+D1p0u4sUL44sG8ZpGAEQEzlE0oUlumZzD4BJ5yyagImpj4fZhstjMnCayTGz5fkDG
hIJz1jHxHbJU7CuZ6OA4jNXRP7r6u0JRSqw1Gc+Vcf7kx9D9NgyBPnZV7pz1BI01f3n1qISxuRWJ
VEzIG4Kap+6dPnWIQ9hM1cQgNQNoBJAG0exkuEBrOm4JOrDRLB0vUA0sYsWfTAbe7dI7PZ+Do5aB
OdW6sVsBSoEXh4w7/K5YVtI/4NTTQazfsi2V6jrUZm8Sa+ok0h9dc5ew/4PBGCi2kTUIooN4pTZW
xM7YgzSQ92avVcq5BI77iOZ0s89Lb8Lnt52468/ouh1xkpYFX4hUzKm3YScD4h++cxNZF2gfsQDB
/9LqyBngNwuNN/1n4HBiDecbtLnyba1Rljt4R1ciK/uYOn2IDFB29x22UV5crHqohgZ0RBT0md3p
gU9U2ANd3oAZEIxLo1A4FJM5hPpoeDIHcdEDm2Ep9UvnLmm648y5c0R8BZsf6AfmAfn4/ZkqbkfQ
4ewyYgj9Zf4NcTPMBRQATJtKPPrlQpbaQW2TsUCAHQeQRzaNfi4w/CMGum3qMwVQUFFSONMHbMnU
RJ2yy2tWtNrObvRINZwR+g1HGusx94Ey3fFtW/6dsI0hWArh7V6iDH6kyhwFdSGXWYkmLEQrDNC/
SejPyrqmPtCvo6NZHfexbWq7szSDcnrHlN2g2nXpiW6KUS7GasE0MhxQseN20AlIWa1EIa4qsxg/
9vB+pNcqOSPGhkgrfUOGG3lJeI9Dg2TuT1ys8OgW28I6RuJMb0SLNkT0k30qeDnmJk9SZoG6BQYi
wkD7BnX5fJiVpr6GYHzAOFerIDRjBi8bRT4NI5KsnUSs+waXbqCTNYS7j0+zg0kk+SsebiyeRh90
QwJTvu2oAKyop9E+gpfa68VC23UdygyLE6bCo8HUofAuME9ubtoPGqaEpe0w0s7q5vMxIXqw7NzV
nODtQAALzdpWlbF5kgYSB+qWk67StmjM9caItgiZV/WNzf0tH0FtLGDHctzVzzmhzBTg/o+VRQfs
DAIiVh6GHZwcm/jYMSX7KV2D4X9T8HFh3EeERnBG7pD3bGaezwwXptALB4xkZliPs/P11Aoat48p
0OZESCqPgqFaKxBPme3VJhAbvwpAtdUB9ckZ6aZ6L9NLo54jMhAXfq6hWA+V3mYt3PSJGPAyGTAn
5BKU6JHtDsjvHHFhYoZO46rz+QCA6EH6b8jo20ZTVJghHGKDkKW17p6v3OueBQiHJIz0eHyhP5hD
g7RfZOi2UMRn8lWs7db0xVL3Y+FQq+xEnYh3kJ0SMgTsediU0gZoArxW4HVbDxzDLyJBj8THhJzB
CEw+3WgLl2yG4bUBlK6J/SZ+qoRPpwj3Ka8Aq9bc6Sz5y0drBSPa+yPN0R2xHsRJ68UjD0EXNFB7
l0eVjciznYuCgw+cc6jGNOcvn2lXNrlLxO/k5UIOPyGYYxvRvHOnYK0XmA8y9QKxvovyCvifPfWW
zIMjghr5CEndoFVFGumC6qpyvUhsxPzQ/dI1AGhMmGRV1+mOmEXjqD5Sy+Dv6ypurvdJ8r4NSYM9
LhgwSGbwm/v7u3O6pbLDnpHL76aqwGY7bTQDzZl2xrwGwBr/MNpW/5cRsTQ9jzytLAfmrfPWVCQl
H4z3PAt/FvY4iC/Ky9ysN5hqrJmpZRuoQC4mJQ7X5qeAhjvxM+fsjEeVgbNhH0f4da0AdYUgOKYp
H1IvT2FyxwhL7jnZzdJHgx4QBq52bemnumFIqEm3U10at5banNqeGUiNPs4e4KTkWYyDjwAw/xvM
l3ghlfyjIz/ruOD3jXDxT0cIEN7EUhlAsoWR4AuhQxIrhlY9RZbo5BVN8LhEy02QqPC1NQ/mabqI
lkiISvh765AUkcMGMOo1KAUPIOp/6IxgUaGSSXMtIMXwpwYaY+zpVDmGGWaH8CfK60oKTbkGwvfT
fqVDZgYW+lHNfZYllgv5vWb/05zApz/j4Sqyljplin49SCHKGRvtqaPoHQ3JBUCEM5VJ79U21/F3
kiQoW4bENs+ZAkSk/Zz8Kp9r3zWfPGeNhPA1x1TQbwAt1LkdfSU8ygIuZpHYDtYMzCEViecLeJwW
6zvtprhFzbM2kR0P7wdPE8nZF7UU5+/Qe8rmJZ7kFiALbw68Kqq6/pGwWlEw0vdJg3uEs1L0wqMC
TE3LtHXlDttCRXP7A06mMAioKwGidWAeTrfhUG0sqLxZCEFMyEkuLstNfpGa3JxtVeNyZTCuIeHh
24uDlTINr79jxHl5nYHYYtvCfKHID4+IosDrnuEyyUnPBLE2JVC8AtBCnMvN0Bin3RqPS3mPSFpB
WLcMHNuIAwcKs/rq9V+90lBquRe5JVcCAQmlgPu86aFCJjwGbwLoDJtRccQoejIZjD35td8tF4ah
f8wBeJdp+FkEefJ5CHbEmp/jykDSfMCIQhDDm6ev0j5kogGAgdx/qrqmDwol+YifJNsPzuLnJoVu
pVhS3sdjpmr5cH/HBv/TDP7qwxglA+yiHYjGRi8WTlVxHY5YENBKeCFLbAHOBas7yrsWo+46ogCJ
8suM7D8vNwfoACTgW7fiEsmCa3u5sb/+CZLw7JlBZPUJ/iCJmP3Y9KE/efcgbv4TCSL/f0Skgzvt
KBgIJKoCuWQmcvWG78D6rIAa91wVpCYla5ekdUiZbXsP8S/v4n1MvIUegdBqxIJKFeBmzZO96V6h
hXAMdDcTtZ1Nh7NrAyHmfLNs+5P2t8xW9jP9bMkDfMAmdLNMVLfV5vZM13eyMGdpKTB8iwjK8bK3
KyW48LE1Qu+m7nfkKhu7O8LJBX+rESaUGsxd04Qox5CxWCQmLSQhaBDaXAf3vaKdHQnuL88j3+Ro
pC8G6u0qG4y6NgC+q0Wsra0szBW9Xc95yUONwimppD3su4I8irZSz7Qr7ybhBtd11pNX0Qfj0ji9
zG7S9qkhCiCvViGkMGASZPvsDU1MU9gT8KuR/UQc6ZfqkPxS2xNSW2O4m8Wy+m7ijqENhNqoYicb
vyj14d3B07aXjjS8ncw8utRWRsHpBtJcWVWhjT0Fjw0EbG0XQfWVHydY+KBhaEIpXatohb9xtO8R
tr0l3pe84G1dQNUrUODmawcUMQ080SRTZKWU6woJg/jKqKkQwh42WNaElkHl7z98WE3bZVMJkRhg
2D/VrshPQCLVQ1fsRFe4k+E181QbB14HHLfPgmHOZVoCgdrhQ/67T3ozIWyC+3CJeFrbK/AvEl0p
zGMVxUNDt+eYEAoiXDPMSjyBGLnOu6TYxcYqcqftjv6omr48//dZX9LKpN/ZixlgyRQylB/7gAgG
baynynTlblqHBENuSHkDv6E45OOo3V9ShIXuw62wnWbwk+00e7/P3KOwcifKd4AWVtNLT6jIlXt5
PAzTzW7ekmj541MhqOgTJ3v0Q7A9//gLfwetvIFndxdAfdp87dlILUy36q1jt21Wn6zh872dbMU5
N1lt2mbxGx0qdW7OkH5rghbi5fdGdIuRD/JgBl8iwcGSTbFMR79t3AnTPThObw9CY7Ti3C7/MjDI
h2wT5C4BE9q9+7lW7IgijtF2yxcMm+CbRnTSIt7027RoJghsh79i2E56bpVOCqqWMFiGBNftm94n
+pSNhkNdeyMdfDhNpu90DC6ce9sVvVSkh/NsUawBXOE3LI8DG6eE6JdJ4e1y3x4Ai7whjpvCIvoK
a/EaUvm6GqrlK+WwLFNtsoOb7TyF037xQ7HTzww1H6I3Ya0oxdcHtw7ey8SbYG63/fvjDvb/V3NN
RF0p30V+7YerSy7ID+zJ0P1HFhO1TjYK5dFpMema2Vxkvo67L6zA9jTbCbJLReXfDNTn7BrtW3ni
o1drq8Hcxd0PiJi6I4RSVJEepv3l/u2ovrbWXCybhSVUIIPe5/KGhHhfhr0OAX6a9UJQYgBbD+i2
g0p1R4wAEJUPm8Nsw9ZPHdKDEil9BGDPUrkLZhQEi/cyukCLlWnBQ+NMr+/R4phi+9+qcsxFlP9V
G29pzsQ7i+Cc65IaC/mcnmrv6yPR5CH863ugmPaz0JO7zAGwcE3GUUyd3sCjYZ5uW72YIduny+qx
x3V5MMyV4AtwjmN0G/mBabiEGB7vBeEDHJiFeECBYoKNbCuhkhREXxrCyPmrtabx1lxDv2O6/Rr+
VfEcaeHG4REMgsMvL8tBN8FGIgkITUwVuZ1o23xuubaiu5Znt4yExjfoShbuqv5uD45mtou5YMeH
2/0CmxUTl/cyB66GHAcX1fhUpr5qPDx4YTa59iernPmIW2speFURwHzH2NInrjDvAABAU+A4jeyA
bxNa921YlDh2j4rN+26MmlDDlpa9Rhy1pTMAZjKbzPGv1ll57byH8zNH3/co+JAcYIJNgecj2ItW
USUuxTcTHxFWrOBWuw20eYCBSZ+QC0+Clq3Av/2bFgKUDI4VuDu4x61v+LDMVvdw2qzJ83Ctwn3f
ALiEuvhUK5Oi/eHEuCYEJf0TMFp6tvydj0l1gMJRz25rFM8JHk+21ZTUAtqhSsO14AVEbroIYAwh
+oHMpx8GnTUjgPkVHfuypUHR6bYPmP2lgjlt9gfDAOkpnqSLwKj1sI09tFe6QGlRxG0jLGbvzdbD
nIGuPCpETEDOJW+ejYBS39c8tD36w4WYbuF/UdGXRhQQ1JnJ1y8AG//HeIpcqm23BuyitvERFsCV
Yb/unAwJ2h4R+vcfYNWr1u7V+yR949Q3EY0cF9oOyU9TtddwBpGU0NJJB3B5bIJARrNjCUfZrGxH
6E5RISAxaMLoFiborkbF5oeKtLUMWV4eDKhBeDe/CzvTR7nAbnKn6ShqPgChKCTd5Egqzo6ICQiR
+CU8sqmClVmX8NMa5wvhiTKEeGmMXA2QlU6zK8P9+oLVeRrzcPfOp6VYzwgySS9mac5YWm9kS4PD
Ghk2M1z2TEmS1j37xIms/M3uTNbhDK8kjpZBIUA/0Zcdi/5PbmKMwDcXoz9jrAe3Yp9c8Uo9HgKN
3JA6TXSVnxoBt8ho4mUwB4cHuFcGtSEEO1LvUb0AhjLnVkQcOTjub52aoKyHQq5QtI9KE7dOzIJ2
YtpV9Nho7jPFj7Rhe1mEeo9V5KKBvKXmTF04yFST3UT9l4p0wLftfnsgl3LKrqP1GyDhk3gLqamM
glbbhuDlAPYU//FM6/WuU5BqFKywlvYIOQZrk6mV/HsHrcQkBAjU/w32xK+bN/2M7SFiyPAwLtq6
M8wmAc6Qqg9zyklyHVY0izyTljlfvr2LWavTAku0vUF2cvbWoniwoZNk05rtOffNjgpUOgIOW21p
0oOKs+yAs/jID0aKBjMG6kss0BAYS29+Ppkbm0WHDqNwvT4mhJc/kVZnDJJpVzdd6KQeD9tHLQNS
6wfBA5+nARzEu0oZZKHicOpNFXHsmC6BRPjw2hjupZU01nwqJHoFuQTzcSEy3QyH5az3nHud5M8w
PykwtwCE2e6eo8ZvXSERHFrYLy2Cv9iXZz3bGSN82wIyS97M5SQJDONHeSrW1njdPvpjA8Dto9LE
g95IbcbdPb98UVpWXOe4r6qbYBJmHXbfND8nEyvgZqiwBdxyyUp9sq2qxZ7M0ZO/5QhnY84zEBsL
OcSuATV8geeAZf3wqIEwyPwDuiVCy1Zl2/BroHhDgQ6IJgWwc6u6vEovcGzj61trdAuVSeSQatKB
X/XckXHPdnUGlWlbYoYwj6mzC5AmdaDUXXbTtPj4ZiLJY5H/d/YrI84nD23xVRyvAO9nlPCFQL/0
atv5kpNZw+eJMVFFqAoIJryozQGw56ag4z/arkXVIMG4Kpum01ygybx496MylH/BkcLMoyR21BzN
nxjDB8Vgreq1xkaERoxqHeD0ss2sIEMf4QB3tPqo+ajXUYLWRBMWrP1xdi/Fwuwx/AVrz2AxwWcy
q05Qm7fWy4Qv8O1l1sjYd09X+Dw+w7+yX0wnu9TEJvGOBn88wnG2T9YxNVF5u7hj7bKVKjqi4oNd
bgk48ERg2+0nP0s0ah1T/6WG8Jt9aVbqfSbcZaLD+TYi2YeAcJPmQAI1c7BpbsSlLsBw7U0GQQcb
ZwY5LhVhpgGJgWbaBFU7IJC3T1qco+JYLvUrKDuS48BIQIP7V6U5a/e1dbf9oyDuxrkQzLmsbesT
lF7Ob7kLrRlmPNOcTC3I99OUyhbqzuMELRgeqD7esdHsNCiGEkGSHy41Sev+GqYSb1vBPN4z6Oiq
G5SMxNYva1ADKgMJLkUvxfF1l1FJdObx013SE9KXlElF+DpjYMWm/JeSjxCRlFRJMay1zuWIxHpc
EitR7+Rf0l7pVZgyQg36eu1utGiMXHXMRCRDMFeGro6XDVATf5fthVZGO34j3ISTVX9WInebL7wm
0VvghKLpoHMPGvrxHJZMp/nDmmVIzzwRlkI3a/iZwJdbkoRQ0HHOT330E2owrze0ari08kY/bvjM
TuQyPIQHSKw9BMhms2hHxAaUgxRzZkMu0EcAHB+0hDS3b53RPaCkMIh8sbTU3V2ipMh94RCi6umH
Ju1UfUSiu5MVqGfz7FwNYuVgwk4AAPsvmG8dJAS2QL6Z/+PXGssKAYXiypYsjoZgxBZC9Jq1g6qR
JiCOslLYUXSWrXYL0VFHr+g7Y3tEK2wbq9IqD8KYCnclQuywnJltEqKHA2bwaJ3zGP7BBFvX22Ow
X7IPprjEeswGtWvYXiXLSQbgpzbbTrp6UTQRzFP03wDMClSvCccd5hhn3pTCBh8r3HvSAzE+mG5p
NgJCR5Q9+fw70Hjx5/qW4SyS+NxDYKU/7lbe9UAANyi53oX4VFo9fpEl8G0wuh91O+joKCbKLsci
/fVWy2o6JuiJ3IILdteSVda1Itc10ABjpfvmdxy7B16A9ZUpdDeL5/aguGAFpWxVWAKaj++ekrvW
FbTWC8SkJyhoITyN5Vzg5Kyx/rc7i4XzLlQ7oAqFY6cSrSTMmJ6Ur8tlH9Vj5Ig9KsqdXFTLWlVc
4ROYUlfdvi+STqJaNkWyz2YL+chsMP1/BG/w0KeeilbLWvhwJLMlKQbiqK7dmeiEom22n/2gmzec
xufkOxt9JJxeC3ix/MZw5actpMl3nnsHI89NvX10SavcrXCnYmvPqVFjtLdn0Z5CQwtIUw74cCVT
WiTtXgUjIROcJLTziVnxKL2iPNnCURHjk4B8n/JsdoY/620qeeezj9lAnC30nPp4wbuGjCyJwetD
ZaKTm5hnOAolymUqonhyaruWyVBy+XrLn41IBIEkvB78BbugQJitx5dtcOlgjFewn6JQtdHwAJDD
MFg8+36NE1iQO+6NS0+83vYoYezx/ust7mwvjitwBhel57y+Zs6gD0ffGPk7wTr/0P7BeLCoFRVc
3mc3sZH24t99PbL6vjYQq1grH66UQvi5UEtOdYcIx6M5a6DmrAqTyl0ybw8OH6pclwlgku8aIu0S
7i96R0MdpDUfH5VWem7tWmhuVANFlAp0QIVYpatJCZ0WJ7+ruWRRd686/LuG3FCJGZRC72dEys+x
DGrLIoqOIaJZuiN048LbL29I/VPsK0oppmXhwEVPpBD0VirOEgKodP7Bz5+kyJrncmFVEMJYW/Mv
NFp82M0vjtvf6HuNj6gzoSkUubYUSRsLLErqMcHYZ0riVbz9rcSf8F4YuU6lKgyTfnDgt3fq7du3
lwEvCXSuQWYax/gp+KE3aywiAlSHSO8WRprzlG+REiBZo8dziUCa+9tc9P1wXFN8g6rO/cujZTAf
3bQo8q8xKd75MCkSf8pbS4ya/yvtqlwBkbCU9TNi8h0Kn73Wlui7sbk5JKnxS1bFqSo7uKxZgZNl
JXsvX28B7KRwq3gXX9zJ9ckN+fMFGtxcWiyaqGHtpBz0zaG+O6feY8A0BwITkJYerX2PQYCEs7xk
iYUygQuus+kWo7q98JLOAqS82jNlJKPkAPy4jvlzadmObcMIKXyV5BsZ4pxIYhSz1Az4CAXlFBwq
LFM+vUXYHRYAHxuLoesuL6uSK5j7gHXPXdifS2HZri24raBgVLbNgkH1h5YGHqYJG3R58G6qeqIA
RVu7uxZewKY/efqL1r4vGB/N1oL8Zput9ZDVBNfcFzV1X7L/UbCYmUvlle6AFVT57cGGiLEnaC/r
FEdLPviP8kURKlLidAZ9xftq898gsq85EPq0YsflhL+IzAd6N5zUhNMhG9XDwM9aBR6tCwJfuuET
F5G4aMZXiyHDgrpouUSpOxJYGQAfdMXcJCzUHMbM49p8EUUWnLjACRX2VdFXskVnBChVDJgaWWj+
w0LdMVcv5CrrAzHt611UVda8W2I5RZqgRHPlUiYJweRWj2WN48KVtXqELegzKt+biZA34js+aRvr
xzdaHdIoNASnLLeG4+ctiGGu05S6g/jnMofq9iC9kEktEADt0gFSqIU6ZGUPWYQkC+5pCVpuOCUW
Q0LnshxqaMy8i4EHtkYQfjaaL8bD2IjlIAj8J4Wl0cJW2Eyf5xXXNcr/O+Zb5or/PeNUojYR/8sX
bs00e01dhHyY/lEWeOu7bLwiQJL7U36y993Nhy8eO9Lxz9JIKTTlN4IFL5883A4meRtSml9r9A9Q
dwqsVdMC/SM+baQLgLW7HZx6Z0gp/Lf54pyaV7ZQ/3UGa5ObUXGh2Bf2QrE91NtBNxVA+TMCUNIi
ouQcvqor87hCqPTzB2LR4/OcHdqigl9q14emwhX5ocRDA1pa7dQHacEGEUPVBjsvHrhOkXBShFgY
cOENai9stHPb/fFcIJ8uP5fR0QkwW7/1pkLs9Su5ejBgOsikpygAWTHRwtyd6ddhSg/AwhAyfyct
YJQsm08sXLE4VOJevex2x3kv0AvSQzrw4MkZ5MR8bskBwv2qMRP0bOdy9RUnodQKw1EqBs1Rfj5N
JKBQ3JKlDdmIfyzWSO51T2b8Eloy5pqocEU+YfP2Ez8vMFoy1budUj/T9cDspxY4qhwtVh3lLtLu
0RyY0yjY0SasNH4p1+sEAyA5vBA5WuRjwfSy0c0vAKcsE5dIinBTF20Wu/OOyiczCaEiwJOM76Vd
K6nGOnwSTWh+71mJIXUzRJ1/FD3Gc+5Zw7sZENqSVN4d20zaeNTepqUeqMQqHoRgr4pjQWbCEXhH
dkEUK3rRz83LMn7HZ4WPuvpUi4ZxD11d0hVEIISdoVjTiYALd0VF4G/IG5ejT0FubfEbT3KkpUyN
adeP1EiBbcz9oJ0F2t0XtMTLa2+mKrNT1zj1bcRpQ8rejyoMuBC/MhYprzchAAuJyWm10UH4t1C3
m5/sYcBqpOhiFhPMhnMzkd7fX1Ng5prlV672dxAp9K4tToH9zUyjJE0XvuGp33U/MbM6G96v05OY
fp+6Cb5GXk3jeYKnCCKdYM7/T+bkHUa31fYUab+C9FeOJt343MBjb3bWVgIvFTIke1R29NiGUJO6
ILvibdVEnzgGQVLUnk27ZSHh3n4VWKGNIqW6qT3akkoYSjk/pQncgy2Mcw5+9/fQvHYAkWCOuo4p
uDJVybZ/crsZD82MEdtPQPJbeFtXvATsYTmAyDT5Y+HY77cJLpFMdFLVAFCBmzfdwJS3LHtnqLFy
xY3WcezDo06HPT/lk3mv+XUGvyGkxPJe0SD++zAP/HRR28tYxBgmurFC6xnDc+UKmVftiFeGeldJ
jsRbQdW66tx/71O5QosZfpL9b95/tf3tIspAHdsbz0V+0Tezc+nc8J2KAbAZR0BedQTZ0Ir6eR9N
szk5W6sf3lnlhWhTTc7g4KeNTIMbggVBUcvSyeug5nwcjKyarAN3/4cAOAlHsUKfQGSmFpjk1oda
n6NxuooxQKjkGTP5a0pc5mhNHB4F4FCs5j+FBC0OKjRAOV0Y9dRM/Yw7DFRYkFW1lRvxnjzvn/zb
VatxXf7j3KStY31QZ0iNBv/4uT2oJ7UI3LonR9XsDtetM7mWdWrWmsDLGn6+2qvuMat76kNS51dk
GoMxEu0Hy7UrXeswJgusHULQc4k+Um43JxNLZOub5UD+rbiVmhC/aBfXnkqHpMPVRqSxxvnPvzPO
CkIXVMWjU+5B/ftSK9HUQoVHC/xBke4XJ0v41SGYJip5NED2XNpnIO3u4cjoEDF4PYpIBTyLBDd6
CTETr2cAJTmhzB0hH/IAmmW36co1+WjwgKSpS+GK7E1XS9un35lPMb+bfvGR5l5HqgFseIuX48ZE
yfmTMkP5TjcxWfKLqFoZ/aKA0X84HGNws11Ll1xtVCewmbliA+d6oSZ1PPPU2/uesdr+QzDaqtia
beo8whPdMli3DYymXf3dCC2cmwO1cnn8Ihgi8CXM4MlMdl/K9mfIR44g47ms1fcdBqozkWdITzqb
okQr9luCevnD+Mrxre2xni+h/NmPdr1xman4u0QdFIdYp/ftDqLNc1tDcS+BBvNutimOcueSu5qa
EFsDxkiVnqqPs19exuwVjJMM2xVaJ8YZj8QbisoNsBzEVhKAVnjzMsbT2mqbJUqMTeDRWExjCmXS
JqaHRtVs8cEiMLqFB9JNxOU2xAbgD9av/fqH+RiGtlX5VpZ0KED9fcaPnQpz3wRqVd4IE7V+bYXu
df9XxGWLry59croT/Tukh/xsDy+Mu8S3oQaiBz7a4pW7ekosZAxUHiexLUDZo3LW2PpB1UZl2jDI
XgbWtKHj8e8xLRlMF4ZdYeuHs6MoU8PToY7zs6kSUQSHEAhy5fEDzyS6fNIk4GaO1WgBjQQM24LL
shKCDhUnYbjNwNZtSDZfWUoSt6PopiBIkhU8NISVoeLnQokoYeRRAJZHWJ59Ev2iyp8NccpzEHUL
ZWjq5I52KpMUUPeWHf9v1HbbmuPBiu3PqYhY9tIAC13OQckAoB3EfEK1YWIeyiygCLst8S1yzGVo
+LKBX82UoD2Vg+6QacplD60nAM64OHT+GupFAw++SMaMEuHUrecmmav53WV4cWUKKwAx5fz0ZU27
TKDW4uP28WxMBFO7HAxR/g6SqsBbZDlA7g7Ih9t3hefPZ+LEu/OYUGqafMmMceP157aKct/Rn/K3
Q3Nos6vp1zXRacwF0s7L/lCDbTHWcOZm8Te6Xo5qtfklLOub011DsojAvK+hbLYuoN8xHFiXg06k
NZRNfBtCDS41uABVHogT4R/YrcPX6h1VofXdUyg3Vlut3GMzwAStA0NSjdvtXJZ3FkucCcm8KeOU
z1SFb9en7ybUobSDuQNnhRCkf05EwtYzYV2Nc1oAJm7IMaDBjp9c2BxwidhQP2oZHLVennh6O+LN
hzW+Jvimlq3lA4BZTHad1JFEEGuN2HIeeEq0BE5FMustJegp/eeqM7ZpC3POlQVsASFzGvVx8kZP
ht1VRhXLXpykjjh1NvIIk7GoUStnP5Jz5s7os7trqoh52aBVdJTD9LGQgQAj8VU/akdHw/faNZKl
p+s5Cc9/9AnEq1ZcICpt5Cj57Hz/To67kP0/zZnR/A5SXJZ9QEhYhItF310IGrhyFF4NmeBh8/91
h1P3cNuuwty/GHfSOg7trsqo13QW/rojJSj6/xB+/TsmU1H6t2xFSQQR/P5fDiMMLyCpUOSBXjmG
/ZDpQ8SMOCbeEqkxjOaG8ru1iZtDWi0mXScMXXyvOrR194gGZU2mG2slJGUN4uImIRlK/9BgC/0D
IvEwmcxjis0u+3rEAOro/A/U+b0PrEZ0A4VLkblI2Ilz0OcC6nnISHeKf2RC4hUFfBFzg9KvXoK9
LnU5WH3kvT59bVS4zzrj4u58v5fdbNPbXs5EO1rCPccsmE9vcgbi8Jv+qsoH+MApumM3KjTfLesv
qzSLwS1r+cJE/K9fnC4f1RlrtrEYlh/OvKofn4094eWUjwcU2RcXnLlSp+4z47z9po7wxaDExzuP
Mxn7qApEIyO+7bvZLlGo6PGnvr+V5UbCwALiChw9EzF/1GJ93sX/uvvWd36dqTlMzRocznfN6oYf
EAm4h116IY6ZaWTc9lkp4VHTJIDXRPWECzLf19dGPmBb8neB5gfT/t2gKFjNrvRLODtVBW62j8v7
fk+sp+OHwvsDoRVQhFMd4PQYnGcL6dfRYeisyCaOJ0PKJpAsQuK0DxBq/wtDQWXqtYmHE0JYbS1u
/oO2M5FFt6qGXmkZCxXA7Hg43crul4tb9siy7lS645oap5FCUxzpQoa3/lh1i2SmFmaNkqScuUGy
+ZfIKqqZj/eJZ+ebdL89N3TqCtZ/CNb6OAlmGjXoVimcqrkuUTDfTORsmBS/hyx+mJpd2SnYyxzW
eMegGvuP+BmUFonfzO5TyEK+HXsZoUCzdIKQX0BGYN7UQp7CDb0VEfUkUSIFPeECZsMDV4F14BNb
04gXOJbdFa19Q4WspFsq6JtCGdPMBPm3C6/zissbJyMpv5HepKhV1qJsdHPdS3sJAKBVa0aREEcm
cjK7g0YnLpvSDxHjKWRDDRP04EBkZs4ZcnXUXBlKAp05/finRUKCCdXgEKnWLDvFfajDgJdX1KHi
JusrKUFdBI/kQOgo2CySKQ6Me9UbcdIAJbnZS9ZPkGvDCC6P0/pwlbb8bnLz27b3lKdzleoT6mcf
E3QH2tDr4zPvRb/p1kIeYu6TTsTIKszS6AqQwSXy3mpKucYjl2uCqSViMaLOo8PM+8QowYuCWCXu
aIPvV7tf7C1zo/DK551tY9nuM880jkDesYBzp6D67QnKeT13vH9TdLngPHvME8CaVGvl4wy3Re7d
W0Z79fzg0SfxQ9hI30veXsfMV0JSu9U0NdzJwVJvVIhgeww8fMj5YVS28sIcR8m+s1LR0MFoVYhW
04sh3+RCdQc430c1BVuyt7C+mXGy/3Ykp11RZOwnYr8a1P1hrLIrVrS5KWLy5ir4U8cPpmZWuyXy
pkiym+NnHbmxP7NkgC9Tw+0AGC79BljUbopSy8iB4vlpqKrjc3lJWhxDD7g9etY+wedJNmYP8HCV
r/Vf/w+t2C1N9aI3KMAf1hRDManig3WA1lbtoSsQJnn1TB7ctpEWCqiY7VMZtAEU2/X0oNH5k+Pk
bWejw4dRp3PHWg4IAPjgcUnLzztNUI33Ys6Krq1POxWa3eM7+mlpWq06q3IcVNZCS/otTM4xMS27
pI9oWro+thEnqASVJ5KVqpUiOYsiu7CgfREZwOuNZQj4dJC2HsOKoxhtsy9/xjaHjd8aJ/EHgDwo
jlSf8Av9IOr7FNkyqzXeuQD7TkJor4MfxibWYwF79H1i7nSNyAQNKIhzonmporHFOUYWlAstUuMV
KsFwTcCrkhnnnqzNm7rJpGlOVMoaOUl5Ryt9K/89xXoWBgQsk563vF8wgufPtL+2aJELy6IXOsuc
EetXd5cqBwvGrAu1CfpD/7HURZ0ZcRhM0M5PbjlfcCfU3MbTtHB7tNs6jTEFWfkL1KH/ZtsleSdA
o8kVkf5ZgG4Zyn9ujgm4ROsLniP8TRFEw0smVdicJa/1x6+6FnFa/U9vfCrcZhZx51qddbgjyzQt
yqVkyVXBkMefxUJuIMTiftIntbYoRpl5snIzuMXza7g07i9I+pK1pXUbvgB6/Vm1969R3LS7r6YX
RN2VcMdNTFJ/WpdvYiUXfVvBrH3rUFsmARr+OMmQkonl/i9SSiDrWH62cmBj34e76ar+ys2FB70V
x2J5El4y9sP7VbwO1yoNs0cPdYaO9aX9pgSVaeO0+K8TBz58QxLhNpouU3nwxEDPB5L++BId4mcx
zFG2C5AfHjWCGa4/73KYveTmoIVRMd3t8MuSq+ewZtextRcNs71ZTonTsbK9XBdX/CiGS8cbL6iZ
zdMi3KLBjnr7XzT5os6Oh+ouxkFrcGwr14s5jX1kkz5gRawKDVzfOFbBK8N3es6ZQHHQIY3zRTcx
bSu6hK+bH0sa6eXS2tqNXDptYTOaAJM51Ip7G8bZyEDng6PP8YCgqpMcjPqo+gZ1Ttfe6rUq68Ol
BhVL0E4c3F/1gAkkEpW3jjSJyXLE1lLadwOGlbPCVO2ae/8wq9LCSct7nIOiSWCrmnIJSff1LGyb
t3rWj3QbSnihyG892PGW1hVG9Mni4dhCFpgZw9f++AVgxu9+zmrvdVoqckTmFJeQgLCBPjqfsQH+
G+r0VAidSSPFF07SM2qdrAOdTGFTgFr1NXDWYXSP7PVILGZ2leSKn0tpY+84L7MuFKbuMFt3jBx7
pwtpkLcU2vXL1BVfIHXAweHkMogX493UMf18f+dHuIu8/+0TggCBZgV7B0o3EcwE+KoCth6g7H/j
bRGzTUM/ObVk2F7WTD7iBdngyyCeh+BbvUMWjK5zwJyL8wXxYILLIt0WPwx0FhsAIirX/vF7ApkA
Cf2Wa2BfOHLPN41+3AilhUmW7BJ+RKnT/gOajyR0VGoN3U4H/4ccXfXTWWCww2QyOG05OrKkxHt6
S8BILqwG8CJAcQhS7s8TE4C+vd4GKSZy3dLYYdWWz15HS8dyye79TmsBb/bivP077iCiGg2lHn7r
toJlzJ7b6fw+vVOHyvzTX/abHXRZUX16ql8Y/+thzPr6k0vyTWlIpHj+sf0Z4Lcd6HRt39u23zPl
9jqMzUDjokg6Dqq1We3ambfw+QtcXpahhgPr9tyByTCbqLmp5GDWWxP0RCJBPXaZf2iHcJhhr4ET
K0SRM7WMUUfU469UqhMRY5BmaTS26eLChVr4y5R1kajqY6YiO2OlTOZe0qtUlUcPCidNGWNeoAiM
i+sp3l/U8JL7Ei++CmA5J4FgrRVhpw3lxkQy02k7KxHQeD0WwVmHTwRUkVR3Ta++UnYhdHsnAUlb
+VnRknaSgJuze/p9DX/Y/9+0u6grOaMtpOhLGh1LPgMAEZ/+uy+QjNKRhCIs3bXZuPRGq+zaXOyj
PxTRPTtyZQQ89ADp8A2FO468bBlwtFOIVpEryFk1eSluL0c2MST7PnEzGMQJ7jYCB88tJDe1zvO5
Sty56+zY5Hw5b8EBq+dGfyw2ukPBzLz5Lpo5TC1PibQspz+Tf1bfIB20RpBTsxz8pcgWJ59OXnSz
jihkcoJ6UBNSl4/rVR8ruRbLPiR3AV+LoKvVxT3vkV39jHv4sQlz5cbg3Y6LfROir+BgMC444lPX
ckKcf5J9R3SOcW/OlEhNDU+ajT+NJyKxU3Sm9stNy3mrl2XnWgvU0ZA3O9nJVXaHFPO4fWpcYuDW
N9djckQeLPUNDYi8g26j/jmCYLchNkWiTLNqgKrrIokhD2IlhOdG6iezDm/lmhbBghns1yifpjKk
PHZBSaKf2O+7pTGYU0Oy8eOppPl14NhxvoXB+7neEZ9HtsTcPGNVS5LrxGvAYhXMXLEFtv9EVcrs
qIWhD+AJza0tjgY80tdnNXZj8+DocT6j90a2eCgURNF/hrQn8NHCjayacRVxVbgp0MzqIN7HRIpi
yS5o/MkEtsvZms1xdeFtcIujFdCs+AX47jVup3PQEpAxlcz6L242WPpkDTMtVFHZC/tM9s/MvYOa
y8Dlkj38ueLV+Zgi/Pn+1ZjVdRP2kn6pPILILePmBGTfXO/fFSy3hgzXZ8rTzFI/AiTkcwCw8lqL
D7HBkqlrVZ1HUhaqLlzchpRcPCo+s6AvPwNfk+ZfqAah6EXX24kwfGyOqrypucfOmguCbyTSKE0d
SMST3Sn9xFvHWTVNsfejEc4xkAf1vA74V4G79blxEADBQxYpzQSiM2ojCY/BgO11YG+hrFON3uN4
3j1MjPlPP2FSr5bnA6+eeESFesu4bfaBk7njLOYq+wc4U+Qj6oxmVJFcaRkfXcp0V8DsRvBaIMmv
HKiI9OivmH1V0rQ//MW87uq7kCcNwbb7VOXga0kgAYBCE2h5WUo20eCUW5SG8xGRiCj/Lg+B40iV
5c09bhYlAlhb3AHh9kPHs9+kqM3F4Ei+pzxgO+NmGTalZ9OS70lfUeTbckK3WeiTldVK1UgCtXSf
3kPaS3f31dCDWsMIWNBqHG2j6mfF9eAtuuGoJvOwEGJj+IeyLlv2U9pVSAJrBGlIwEmV5C9wOLb8
IT+bPKoJxpBtrmDnGrCVAkm28BzgUQPKUDuRhNpLhXUFZPMIZaqtve7uW3Emx0BKpWmFcw9yU/Q9
gw4fD0pnGactc+ifgjTOj0l1tmxgObFglHm4XsHBKJNeY2HobJ+hRu7ch27+athiKPAFBZWZneAM
8LNN4feSNLZSQWn1S8w5R66Yrsx7HR3qNpj8PWROyl/Sp5+9P1itduRnC2JoI0Ud5cqrjfDucp9G
Uzu4OZcipLIX+ThJNBiYiqo6kvhThNAf49z1qIvaUDJR6u7sk7MW6hM3QIsFvUDsyrSNPWhbGFXe
/HEaPhqPaZVRkQOZv3TCFOYALt+eKC4J1lQLqbxteM+9H7JPXgU4h83udWZinzXIZbgmlnn+0tEu
fNxD/VUkPLEADVfw1GTD7lk8lEr3kPGeYl2UTCdSHCqKDEfXkVIkrqBL020q3rDIohF0kQClboS6
gwMjywaxYacPp4o6AC4U4WhWS3GdF5AUKszlonMO9WG2ZQU5Lz0A2vgKU8Lq+hmVE2sQpEjcbD/f
32j4ANnXVytCqd7BPJ7sB0HsycmcRgfkeuWAxw83dE4ufSxnLS8aXfKYM3yt0rHInK/luC6dxVAH
sVlkibiPrDRdTzIOtXZ4sEie5C1qKkbUlps55VsiYtyAgemmHYbEgpwDV/VlYJAo9+SyaoZZuMGe
PikSlD22RvZoqgbCVg1vl1ooa0Frv7jmME0i6Cakqar1K2mwg5oAee7oFCrKskbb74dTQ44IEGBB
e/J67Rk1K5NxjlwZ6juj21qsiTjWHdrlUKMNtitAr9hemEvRzzC8i/t8QWFM3aaY4EEMeJlpzgsY
RgDq7Ckm11gpyqW0di4XVLmG/ldD9kOqxzw21sVehPFAdtQubBtRbbWx7PKzZtuBhKAA3KDfzh5+
yJQQ0q4STN75j4qgkSlJcM6/jRhiFIpSm42XFxF3Pdw2Gtgh0Gtzs3xgM1AiSwL9+SxXyZUsioB4
Pl+/oEkF4IOxtcwUsTFRVzFjw/LQpCG0CA75tQ3tGLrNE8XrSs5bUoYV7bv3XCgBw5Inv7Zzpcbs
6dAzunnGJ/Lgj4ygYEk59uWHuubbtM630i1lURzRY/vo1ZzGAoIrzMa7BAP4Fv+rhPGYb+fkMnjl
4uJHXlAUhCxZ1ZqeXiRvkDS3njwo2dHFs0wsjXyyJ4xsMoW1sJh5KY6RzdSYqEooyFV45nvdQjBW
HfE9aAHsLnl1a+Jpehh2KBoreIU5bMNkSjUacDXXNPpwChXsaoRm+saY2urv1TEkZO1pCr4t4oP8
n22O9DEEfQ9ly5RWYdfNdj9wlxCg3gb16rmWJEUh1ICwKrmA+lJhvh6WLK4SlQ7oMoRXAFamupbO
CkViMdYUKJjPjscJFZ1Ful5eFiHQM5p2a7dWkdk53VMOC0ib4AZmC4ZS9ymdH29iqZQjdV2+MV2v
jMdpli0NqRvzOqeAAbarE/MUUjRfd1LUrvkeon5bvLy0fCUrEmuBT2iRxaM9m9mXvZGMI+OEA9SN
W+6PC0kGdPeIcDhtA7Or8k4lkZFeeOUYDO+snEW+zabyVttANKmdPpDoRyP6ec0Knnq2fVSY2NyE
kzdpq6fd9WoU0Et87bKNfQ2ykjvWB/oaweriFQvRBITxom3/ssI5yxJsI27yfwXiFCco+eThFVFM
XQBHJO51z247wKmImkjLoZbKH0zPTYyQXyGH595QPx5GvM3VAJTVF4gBsQ3G88VSpXRY+xLvHn0s
9Qd9ZWneFdsekvREZqBWWXcRiK3DEgyVk2VkWAlhDm+n21Rc01XmGMgmL2l66mjFmoApiiMjd88T
FJb9wEHHfaw4WbTjiCXrZPnMpbogeeN+JuHPexjRR25G0Zlenk3lYOu9uzueYZD/8BsglYZUQoF3
b8bhAWKDd8tvYd3zeq/o61FFG0J3/thHCDzntof7UrndPFWXsj47QAzgzuk1F8YkSTOyD9xHUcCs
yqaarZ3bnNephVUo7b/400umjxl9Svyko9P81KI1sfU42AoAPhE9ckLJnEboLwbzdMt2CQCy3Qsc
FJ9t+nUyXlRIA/0d293BMC/ABGP36wcepHpHMut9do8XtuwuK2NTTPZdh9+1/U+AJXNNr9abwCIk
ebmyo++inetptuepLTDKvmk+EnpkcgA9j0pR2yPJxypY9PUH455CZhIIQcYPRcOt0NfwkIOl0qdM
2i1q3m3m0b1GbA+F+sT1emUwDdZ2bCJn5uAoASyHMFA6LBdiWQv5i7D+rnQizRccfWXGU9OKzsHV
uTlJl3nk9fqu4p+cf8k/cpdqKQ5JHXLBrlFXSVV1fMFmclJhIFZmSAsJXlCf9ItnbWXCQtyR9EVe
+Og/Fp9VOJQ1zv5DeKXUcBCyTy80tl63oOw/M6LA/e2E61PxWHbPSS5Vj6tei9dlT7CElrlaQlfk
ta2e45VfJcFGKtlvF3JJZh60U0Xaiccgpqyf5brIli1DllB1z1hbK5Dupy5gvxeThrt6MpE8gISs
41go7rvhMhZWgdZ+ErwCijXHM6/Ym0Xz2B4Z92U4G4EBpMpE/xe47SuHlDqTmMd9tG14L0ofNTQB
kbcvrAu65B9+gR5rCZlWB+23ZaEjAm9Lgkms222E+5ehWzU2RYx/eGswc4h7nIFpMSfwA9cWSnzJ
Yq7ElrrHGE4WLkNNVci6jQT9ZjKhykXv9245EfWoBBwoLmtNeIZcCZAgUbyKZqyipsLJeiam8gc1
sCe0AkAdrDCt69jQ0HLrn+1kF4FT2JIRhoGQPL6iXbYQKQMsBaRnoWL5MUBKOIkrVIkkpFrJ5FI0
5HF155YFQGsVxVAuc8qSGWD6XygqcOo4ST4+VKlL4OWSNic3SfP56SFSTIS8HBze0mZtmyTc1rDc
EBmg1a784kYT3ntwdi45QV3f7LDTilYPXlj7JzI9ZNsbAeCacsoOlCG+bS5DKa6ZNO+V+1YoipVw
y7RyCoNjAjDbcvAlvaF1y2o8KjWi3IIX/5lUBvsontfRRmTu8VBykXldLrlAmAk8ZEx2DxwerviU
+KnF1sMH8Q+NQojVnc/L3z55U1oPy9DRCAgHOm5JUjSQiUinanq4S9rLc1VcuCQLgqIN1pnG2QI/
y9zcokMlk8y1Zk7KoI6zP0idc3OmEgAijX8PPOUiauW94fhB8Ek4gZgcMAUmDZX+26stN5Sq2AYm
vekI7G9htFhQIDQfFPOIGowo2p//+dTIR50SZegnyPYqjT+fbNDPP/qa8dnxX+8rx3lAL+ZeRRBy
jjaz/cNtgYzu0bgOP4NBlxSM6dQV8n2uKKxntixIRJ/oJ9HU5w/MS7zSMwdsI/004r0z8EtRlnt6
xeqYmJLpaEbG+jphTPehPNTVnoPSKxaACIKel0VYU8h/+fA6ui7mu7yi1k2QmRVWNaKFaRzWnqFf
N2WnEv8l81rtRyviWX2/7uoRMmrctok00mTUZ/3h2QKrXZBRRf3KczBZkIZRntNywLe6ReXOf32D
BjSakNUweb8ImwHbUXFQe6CGtQ5HHzCSux45dm/AXLVjCMQYNEaaLWF6sstHoINjYq3cPnhelF/x
SKXUi1TeacT+tIWzf9T5kmUoMI1YablM3FmGs1jtcOpKT+5UCeFD5Fm59mVPWUdLnFUFS3NRYNXu
4TGPIjfBXK+xc9/6WvhOFOOryk3FrYNOve/Wb5cLg7OQLX8457Df/jTumwBxtSJWKSStJwSCk+XL
wdVGXw1m28Jb/Ya5KUU7cE8bRLsI0l45xHKIA9L8UIPuZ957mfLDV96noSF7/LY7KpKT5mfD5gn2
+vmXBUiNJDqnJM6+zgl4fJTHHpyV8CUx8bIo3aEDb+dKuwRjZx1jzWcN+yUPpeDxSu3CEArKAYfI
0WI13Jr1FBvG50Zb/sKjF+Ulm77uYE34tfciC9IVIh5qdIUyINx6qVq1ZrRVjrsr2oBCUIwRXPlD
7iD9XESkpm8aJuDESBzZsCkb45UamwrRTU6pJTg/J2gk75yx7nS3fluSaSeyt6uqUwvf6TO0E+x5
qvrOSwchhXiUbEciooZiMXlr8VjkJ/f/qduqTbmNxizVb8PQqzLyNEKkAV1+HXGu8SjLRHSK3QaH
AAcalxk3NenIRhvxaat5xdsvrJ8y/fNTJY4CNedmDKFr010lYXm4V4bagDGdUdVOuujp+iSIjTEs
VzCHqmcHPWFrD4tCHIEzXWGp4G+FYNZWVtwdjqci2hXSinx0hIqMRO+TJtCXPfaWAGMKdEc4tFCb
S13naIWZ4KhbZGuPxaw00kSWzw5KC15OMfZNtIXT4mVTP4plNtjhXQ54KoqlMmG+pgmujCFhHnt9
IknchD3CgNrOrrFk91aLMXNwuZ3q64D5adv35duYST6fB7fyGdx92l86CDP8hD76ylw7vEW+qina
oO8rduRw77PaOOMQlQOAES4GQW+XSqlwu0NiBcSgzhgSaiuwQSnK4uX8zF48Eg91W1VfC0UpP52U
jYyZWgdIslUjlOg2Q3ByvE481HBitIQqj/ilsVLWRczU8ys73KDVzkFWjU/LojS9tDqm2msLZFoO
QNliKfXie0vc54gTgECphlUz7s2RVtkaG9aKI390Ln9FvZ2Ud/FdsOSIoePn7Fp62IG8+HFeEUmk
9zP6N/63s8pwUunJt8tzfkaezlonHILVay/P4s57aMq8Wb/POSm0UZ2YcGsFbge3Ak88MX2bv0fT
m1Bv62kYDIEuQvPVpJXCmZX+WAb5Yn8DXLChQTJ6iAKC/Df7EPB5rHBkPAFnblcA2Wmc/tq0dqz5
D0mV7Mt4ehFD8K62Lgoj+QLUn/Zo44fL2OY3d3LMQh9XFOOeQTFYVELBV4LuCykraMly1X2PG7YF
sPlr5NtmnSp0AbZT76o941+VCiPfS36rCOgXi9nIoCtA8AH7qM6acArfvZ8VtqNzrfEwvAIH4LRC
Zf/0JwO8gYzsIqEXznY6P1UVotBQBjfmRC6xQ5jMIC1x+wb68L8PEFSCoooZBxUiUfz3338Pj3uv
KLXCYgu3yVqTsbk4bkiM25EfnHkQeGhziLijrpIFoLFwnPocMovKzFfSDfZXUDetZslb3hJwWRsw
m7hXRKHJSF+y5iLz5L+GkBGsTaJVxbLEcUy0ddHydpb/Vw4yZHKw8z0tybpxMa08cSsPiKOJxtrR
asWrF+Nm7PCY9vDyTFPtzx9pQzmG6nzayIMW3FTrYkfE+eVwQIANgxGzM9JzI4IO4/o3Op4JSYmO
Wd8j72bVSWRIlbo0ORMxYTWSg799ljbqq3yPFMbu0W08O+Nj7A9wcq9CQygDIh2hDCSA6gV8W4QY
0CNMW2xRJAeTXiYthECCvu0gBi6PF3Ij7XdxU1aHnP9V5EDTl9LCcEnMPy87GFm3a8k7eKewMJOp
yJb2j9ilXjgU+HhzfXn+sPbZCas1W89h0cRBkh+j8v8Z/WalLTzIAYK22CPAHyfkrSU8FuphhTux
CiHjWzd1G5EWwV1AJmDyI05ay11KAOhJLy/Xq5plDpRrc8puZVJYDTcwNpFkUe7LJ3ksO+cHkCon
Y29jqqiE7BB0+2oLGf1CjPxxNDA3gXfMeYrWCFoI2q0VlmDJsJ42+a0t9SmeFlfVAm0Pd8FN4t0U
onw9nD1k1P1vLbj3Cy3dl4HRwsYDPgvAZfNfNY4kqSYpW7empNIzwQX9GHdC9hOOzVbkfE6TNND0
t76t6wagdAII6qT/QZ/qEfLCpKIfwWvFy7CtXmqWAsHO+ptgDsoJM2RGJTSkOffroQ+g0oftiiyO
uRAv+azpWDn1XG51CF0b+1a0+6Oi8HOWGBzVfeezR+n1PLofhCsa5xJzkgc188hx0Ojb2Y2ZaJNN
eXeTtf0JAtdqqnqedKbPDrdVy35jaVNtwuqvDqm1+O64u64acEuzn0IOWqStYlhKUNYzD3e/3C4r
W5gNrbD3jtGeHvCOYx5q6iclYknhnRLh58orr73j3MgysdWhZWuvcHA2KYtBmVzIYw0ARIeIzJ22
U1/CRME2/gHNm++NZVooJdmGAlnniPUNOy4oZW0ROCFI8dFlXltlNgiAV6GqsKbU5uefWGlKBoc0
iYgh69EAWueMNK9qzSIqZ3OxExE+K/74HQ04X4DjqYypwknp9W8p9ZQMMp0MW/cHsLeod4qH1hOk
ZBuHFI91CHvOOnSDOIvf54mlOl+w8xrJ7o749Xq0zEZKnklQZi1EMZTGmkvtXEFL8VghMR7RxBBG
QzVzZKIAgaIUcHPIp91req+gLwnrm/xqpIN390Gm8yGutvE8BTVA3IxNtffop76GfAq2rE+trG5O
aIX9Ld79EESpImkTkklEeRt+/Xh/G4dnoZsmsbYojnb/YpCO2H+f/XMUWx01O7woFPkEp3QHCkW3
ua0a8Yx2Tn2jHgjC5cDyGz1w5/dG9b/TXNsq9zlkQ6dCPpoi6pG9+w+Mtn122btBEt7oPEXf9UDE
PjY5+ZTx1eMGfb6LITP1wue5H9et7tn6289zU1WI/YGXbiZHfj6NaPKiFf7b/wIejmaKp7pvdv4Z
OOIHJQSZguTCbzFamc6CUFU9YfskudK8SsqXv10eUkjaulCJHBKhq2ekslF2Gc9EO8g5MJLzch+N
gyoy42cn84XcQnk4xm6anFr7MKv/anUNbwVaqRU+XGkC1lVW/lc5AspN0ZT2fcHeEgnGLO34tZpA
BGRmXjo5njAPzoJvMgfA9ro/s+U7lEttMB/7BikVoJJ1v59xvtFDc8pRMMJf6Tk0Mmf5dmJSgmz1
E3q6Cp+A6I3rpVpftBlHG7Y1Om27tspCGnZjC6UWwoPyW6JbM4eVYa0npWm6B3ZIIcgBvL2PXzyl
31PEiubOfnUk0nyjlzH7t3hDkBeG2PU7SEOQWdxlhRoCFcCTpaWJpURjJwpLrKJ9EUjZk0QyqVQZ
xw8NaUHxFgZks9drT4MT4QjofqugeT7X8aaWNgu1LsCiuW81Cprv0HsLA5DCdYE4zixjuAaieugc
kLpsuTOMLT5gLsf0zPdCrbFfAg9/9WpQatm1jTtTtNwsHXzTmUQQ28A8fpQlTPaCYigL+ZK+OkZc
1d93GklRRauq9WH6wZtdDwYMiCwuaPkRwjJz/ujKlEd0D2WsrTRdzw8Vt61TocpX/xayAdLTrarP
pWAEaS/EdNvVJfP8J7vfSILqfRrbffLQOeUaCQLoYoA/KB8w153NOSirzHn58q4DXZbWO3QHWGrx
qhmS9UWo5Q1EfSDPr5Gi0mkxxA5MvDTm09Rqt4onHkEBOJ2ff0ZXmPUqMHeaul/o8NSK9n/yCKt9
h6pmZZyyUiMJn3Fcz4c9cb2nAMeLOo9HQER8wewZL0juFzfdgFTTJ6h7bNXS0JNk9iK4QBEtfu+b
GYVsTRnUogW3GyfWWhrnjLQkQkr+Dl3NoSFDjk73vpdNpqfFp0pLlNzLW3eJ9uD1sfnVpmucYd19
/3f7di5rvao85F7Ht9+PKhvgmOh05MLyOQ/e04p8X62XuEg/ASdLC3EUbjPz1aMUIF7hX6MJQNDy
SbHht1yohaFbW2jyyD17PUrY7xRWDgofrxuk21aIPCNGKCdisKEqf8cxzS+FhCH49U7OHDvjX5DS
x3B30p8wxkkpKAtCrCvJ2jd3E3fA/cUdlvaC5ukrKZBqbRHG+0Aniul3m6ikJczXs5v6/wEaJOE2
qBJohfmrIJfnevx65vX8F++vCVeDHwwLH1XAu0BRK8Mo/n319K3NpCqxDJMfLisx4uRxct5ZWyLk
wzobr2MuTvmKsst15rWWD2T6O6Oe7bcWFpGjYMj+Y9D+zwiqdutXOOlIIkp2cR2qcOj4qUrtsW1j
CVCiNQRvoPIlQCoMeEC0T1NsHki0Na6hMz1yWH001v55FJjfrdNx9jQfcBi5pm9kdxPgqQyIhOhh
gr/fd8Ap2N0+cfDVZbQw/jYgK07oPL7TzsH5NSmBqTSMLq2X9r8jPEpRLNgdfSnKftGXXNPopwbz
Wa9ZsyehxW7hSICfBMPli8ddJaxx7SFAYUwC/zDP3rXfcio3B1QSYE3qWNOBOfEzWbAACJSv1rqn
MSfx1akGhGdXEFjTB23CX4Ak6wUsX7annYFu3VLLOzDnIgutQgqw9JtKGBnnZ92jzhe+HkGTsKk/
7Rfv6AjJYhAKYiPw3hnbzJXl9bC/4rK2UKWxHxiVAsAjC6rCVOzsXgOYIH1SBqtt08qsSLvR/MWQ
hj6z/qrmTmX7BT9TJ/shfHZrnz2HE0v+eNH+IxrPeNEboDwBaLZB1RzByKRmsR7+ObtXhAvp7yeQ
SrFuFqkeVTDS/p5KWHgl92pzeER4ErdMMo0RkHrradGUY2dty1vK/rkSY25/zA+tW4BzOkUxGzvW
RsdaeWK3SUOZGtVO3BFiGyaQl8LIvLB5X+DtOdKrj5LaGf8huFwt2rwQm07DiBhP5T4IpO/AHyUF
qYMd/0XcJp8rRSAxDSm/UgNXeAqEEgFMC/c2RWqCZB7P0PgybHy8SC3GLdUmdbiIDKJNvY+26O3U
AhkMpqr6770dHTbGvE3A3PgCIqvRjvtqPnviHNk4adNplknXc+dL94eFsVJW8Y3EVH7jcdpLqV1C
/uC8oSyK1iOMuo1Dw8tWjutdTaStAt7zzQ3G7KNDGt4UxIv/romrSdypUjAnZtObkYPaON/Lq5yq
4ihK/OwmX9kuuz3XUDFE1j/ydubJxLhRDk8L443pL7ixNpEnBprdInPpWqtOXLMsVZWXdCf+w+7i
FuVqJSUh2EmR7A4XaO4ZM+ot9B4qrJJHwLVidPzfNoc03V+DLXrKAF1j1sybEtm/5NZLRPSD0DOC
n9NBFnydKLHefPLVLJ9M2+qdZr51VejmR+AJkPFNfPlRKWFMEBstTTlYXDWESsxg+9HALrFlHUmS
en/stZkkny/6Eq1nETvfIj/F1EEkSE5n62vXwEdUXH1KYrs+qRoeQ/fVyoFVB+DSrZbnA8IvgX0Y
2/rxJyShtXcTeRI9XoS+lipkV+ptg5Ij3cLp1cgurqFO7ZavLgw+cRp/ptd30Ld2JLGAdbw86U2D
QjrroBsWUxza1JleqJjily3l9Bs5SJPZJAEUe6YtCprjsM+87MYzx2FpOkG1cuJGemFZsMVZAvOw
0n+KDJIGj+yP/MDSEpcM5Pmkf0PrnOiH0ek5izZ2/lUCxdMbVgykf3Tuor6c8BA6v42l7BGj1Plq
vBbMCh43MjSWhy0HNp5mQzuxHY8nZ6a5iJa25RKkfFbFpJRwxRpUJ8vUc4qgxAl7lfNiKxvCmbI+
XLuxTT3Gp+lk89PiYYJUZ/prSpim7UfbaUDyV4iFImmgWc+nBMFUqKerxyYFTV2lsRXLJasfW85Z
Ndzlz6os2WGtvpFnPcGj5KpPiqvrtniKrAOEyMkV34vYUAaBfSq2/6/NbjeEffM8uBo7T5wlZxZC
gpfci9w4SKAZ5tvJu73WvJnhKzRXWw+SnXMvOicY28+hfH0N2+ZQQTfKtwXSh8eHpMXrgeqF39/D
4DEZCOh0wJ0a4INK0RU3bwNCZA3EEUCbhFP5Pcyxf1X9Ez0gl3OWrk3zB2l4Fviv6a+1Ibo35U8f
S/k0tf1lEUgRRPZEWaAzyeiOfjiKEtVD9JP5ICviVYS9U3j4haBxsLlv+Fp38DnO3xXHcx0i0wyQ
OT6eur9B6wU+cOWp51NXfBJA5ddpCQcQLHiBrRh2TjUVZ4iI+AQPZEEaHJH/FNknMtlSWYAhBNHb
FKgQcFXiMGD+C74nSpYndO24HEyFdZJ6qT6FscaXcndotJy+5mJmmVE6itX8x075wG9BkPjGphdc
kcOuSNEpjnnq/eoIIHFXFAjCe3SeZ+4wr+qpdl7w/ujbKvEOXQe7JrxqJ9kyoZU0OqKiPBOJVzKS
3yV4d16IteJeyFdjrA3PNaV9MBs0Av0HmoRwm7NmSR+cqCtpTYRZ8HSMyxzVyRo+B5Edd6t7nTsx
s7YLTPjQAtLo+iV0Lh2NCWTENgA5NNhK9CriiXCisih48lxwNJuVrqKRNS6XNidJUL1iR19rxASx
PLCHuuftWC5VBRTyAWAuL2L+NDo3n3yfbJP0YvDDokYkGA6RlZ63Vr3DxRExewkotKG1kujyTU/d
Dwvq9oft67Gjnoh3yO5PL5vOhyTXUhmadULSXxoseVLRwSDNde6rUm0JVMEjQNmORKZjbOtGS2/T
R9WAzRnmB4dYedlnRjE23/4obNUHcXJq4CELxUKmYt3ml6Zv1FEkXzecFHN7rkGPbh6lQDjOUpVP
lqT6n1gbcqqhkBJ5z1aMTC52mFTdVUspngQgPkh4eomW8DR3c22VE0CP3s4bUqUeBOU4TsDcyIOm
awv81koVIQCwsHMV09rhXjDsVs6zvYe5glGtN0IhJDG+/OSjOrrd05c2Q8KpCwdzOCu/OxkmBSXF
ujBZZhU6/q1bCvi7dK5kL+psBKDX6iFIlTB7dAKYmpJ2lyZAWGTDzSGcOBfAbdiEA04QqWAQl0P/
BIh1FlBdTmILxsW0hqBS0JY0ATurSnpdnZWz2ar/Kh64k9bR166k5KWEJInK5OVbV+SeZ81Mfhoa
8t6aYXOlHaVjpIcXtJVii6GVz7Acd+fU6qwvX4zpMd9GKXvo+KH/lzH/dx1qdL+UXPjTVBkfUUeC
CmG77wIDJXQZyi4pNHT+1kwfHvGpRdo83TQTeLdIprKo5TAslyv4i8LB4gR3ZURic0X+qkwYltmO
wyMSR/06e3tFT3H9t1zXATR9qR8CTng2s5+5pczLogfrguTrwdHM0qOqtiMdf0636ZkkMUi+02if
HeT4CjZeAMSPw8vVEnpn2ArisB1Wg2j1RnJ1ikRvDW4+jWtSYuBNiChz9xYYQO4kuZfuS8jHEpCG
ub5P//XEdZunLKZl2MQsY5NKuaelnuImmKbFftrvwOQP017PonNfMcOt2IbTHmD+x4kSwb2pdONr
pPlxRvEmaFwistq0rzj1o7SzzzRmow+WZc6YnST/9mpmbj/6FZDi/jIaxodyD2CuUwKsu/ftzNz5
nj5O8yodk1KYN6EnfrM+cDL6vTA0dsRFqpyEdkU6DW1UOTOPWoWNJg3Kqh+UJKxLmgokU+dai5kH
JYXY47QHPUkvq7/mNIeLti+6ByHCX/lHGiyD2dboxj24xhLJnU89VPkHQEZLtJlkvGxhSHAOrZZZ
RxumCntpmXLghsGvnifU2EZjeIyhg5C5A3p3lmxdSbE1oJR7RTVkHgWW82RPG+x45EmTwF5Ai3uc
vkn3wgkT0fFaveY7Kvx3e+My1ySCJyhD1jgS1gH1MrR4OoNSccUhMQ+unP2W8cwZIz5KWWtgR6ZX
/oSW11Cm4NM25gR6NlqM3z7qz/Krs8cGQe/5q8hdPKeAf9OuT6L+sZhInlraZ/txZXw6IU0FA09H
VqAmE8vlH3TmgWjWPs8UIbsMIjHOWzFMQsOrDwoJfyKq7+k5SsrnAVqOpi5Lk71rL2YpA7bbP4IZ
PH04RZTcY3XqpahUrCUXt/io8NKFDFCV1HnxsYURT4fI6QEeGVOwC7IM7uPj6ZoGPY3slQlJp3ee
IygJ3/5MBwcgrkFU9cq6apb4DaloZwxuveetRqCHgiAZaGyt+m+rIaiFIjIz6Rc6Kt5AxL+UiR9F
d04H0zTQLxZWXm2NSvyRNNivNRwDARn29MKMM8I28BNB1p5xOs1oj4r3dY4XqPPpWHaN0TXqaN6Z
s2OUa6XUS2wTQGlZxLq8fuDOr6qzsUUGevAtONO/l90sdN8OOZGH5Fp6PyGn2X8KGq/ado+m7rTc
LO0HPB4a93DvFYSlvmMskEwrnGOBQ1NXihMoRm3DbNpS8rLlzXncGgSE7y0ITZCOIcvU7z6fJwxW
uyHCzs8lCPXAoNY3dLxNjqM9s0myTt+sUXC7hRSEZcEcKgjaHjWTtRtO3KYkymKknZYZM3z6Vh+/
e8ROGWFrF9crjdG+8ScKDL7cJX5xEz2SY6k6h6u+/0WqDftHQNojBQAfqh23OTU2VrGwxGO3oetm
L2xb6BxZ+rOjYPGeejux8x3Kk4ZJunwhjR5EFr2s5HC05YfToq8eSNqm666g/DdJgQ0endtD2Zdr
bIxewvtbgXAvNXdKFMzoPhKBMmjMHM4iaPu+4f+fhU+2rehAKY0WMql5+T91+1xf0ftkjmhLp4Dq
7F7AnKX7dw0Awrdmt9gkJQtxM3RnDQJpa/zG+AkkXMGfP3DI2tbeHimUG/RzMeoJQXIxqCgKzmiv
6yaVoKwN+DDrUJt0+0WZCAIe+FCPUh1TKtis4lFmHiBt/C0AAQsP9L0e9n8xNkTnIl7cZIE6Q7OB
Eh91lPOtuQiGfxs3vueoJ4sH45V5cXY+9O+ED8PPUxT/NAMaQL1ptIjcHj0CSwk/nIypOuTjK2IK
bJQOM+liT6VLwMWGkBdbajQjYopAwRPzc2gFmPiYest+fHgPNy32isnmB8r9x/AqUbi1O/QVmPm2
u0+iH9rvaCqmitE3pegYQ5hHcN3SddAsgcFuoMP7VMHQQSKE5f8mHUut9KJRFdu8mkCpKAdmja3L
qGYVtAMvt0/KlzcC+ogt5Rj0jNIK2k/I2zzhV5NMFV48OCiZMxdwDB3T5u2Jzqpi5jSfQ8HCx8rZ
lEUdV9EuelmgeQ1fILMAVc4MP0MQNFyc9jITBwSwSG+7fwuaWOW/tuhDZ8shN4Ikr/Z2KoOMNmYu
kZgh9PtFPEiZTPYtsGct3TIzD8b3UXBZ5TrK1QKN8+2K8nvMS1Fyf9p5KCijvMfET3dxhmwjG+XK
tSv2Yclvxr97FSuqjma+lR76jclc8EZ4REL8MVdwkKYOtqYCHcL79AuuJb8SqRylFCrXwyYBH5r8
cjsZMUpYI4j0JZOh0SxgH4hfC9xOQNnGLvf0lCNtqSLnC0NnsXLgqJ/C+tu0TfnCNpes69sW1PKN
TGh3pL35XzGkbNTqcaRFM21HlEQkiOwTLaVuyApA7Av/uQVKONa45b4uNHZ6Ca3PmrvKIIDHwO9a
HiuoJm9sYFQ6CnFSTlsVfwU52RLKerRwvC8CSkG57nLJGeZSSRRSvXjcJLzzVzLyTIt4GZV41mTl
VKc90aOinrV8zLLE8aeMW4cFqk9lAXp1KoHaLl9fjDzVIcBUWlSvs0OjzyUv5yPgXufFNUryX9gO
dblOvYHePV4bOmklUB6ZFKlTo9h5ZRmi4/pjK7fvKv4p07XhiVrA8qFBOMSfRmzBXfLUMwtLH0hd
aA6XLt2+CzhLryjd/HVYuV7dwCqTc0xCVQpcnX8SEQweLMs5WtuMHzfqG/Eug3K8tIM6S4OWuEcI
oR+62eg/7CsJYw63EqrQxZUfnzQZWS968IsPLjjVqX/SB43MQFGPofkC7LMh8CjK/yR09xJdn1e4
bA5Wvbtetmee7UfZuw/Qlsg72kBUMqeFcM1FMYtZApImqOaR5A3gVmog1bhwSAsCu4qZO8OHP5Xu
P6CeshGAsYNs18hzIXQX+6qq5mr6WwoKieT34yTJptHSVaKqfogvLHj/jqAFHjUsR50PFSlLehCF
Qf0KOLFVvJX4w/F0SxWNHWaaRgTiwUDsB9Q1ogpkBOzp0cQT+s6hKrJW5TvNLUG7+YX6Qd/u5F1U
o3pfXeSpa6M+6237duAnNGwpHif/r5Gz6JveDtxuX0zP66+EJZfZBIh4KRT7jawUe+So7j/dY+Lg
2dOiuoBENmgO5aKkf4PejQ9OXO68eOhAEpWpGZADW2OGebln83l+G9d6qhD9Re1GOV8Du6S1C0pD
zoRnZTkPCggIhVqABE6qnfIrN8HRzI8BkX4AxzxtZRjAsi9k0Jkf7s1gvU6ib+dvq2PakTQCIM99
si+wWL2/gq+OX2J8UtMoaw85O6xJOM6py440KTiYmiqV1EHiB6fAPH/EW1mOA7qDQL59uc9t0KKG
I9ZG+UZy0MOcwcTcZDd7NpYssJBY/JTJBC3mF4ZYyUa8fVCP4DSe6KzXy9qIcd80CLuFgIYgyxf4
vLHdNAxsWJpAs/kE4GMwm07L7vOY9kjDbB1a+g19umLFEdiEzyXDm6GxQ6EVmuQxOsRP9vE8k7++
d9LWAJzP8EwX8LgZtINRlxnAoDj4DLvhYhcPpfbCanG3XS+HaQ9CQ5xO5FArmNLC/fD1JypQWIP+
QymkQhscB8rNTqnK7uFhkOOqlPK1wiIns3nhvz6NVCrkIY3vgeukHcbKTiCeFFHMvyOPvdq2XHLN
xp37WVKNhNEp4LrOvLlmOnI6eT+x7Ax64ah4v+KE/WeBEYpaKPrdop828Aa4HJy6yl2M5fxuTNGu
ibvo45ze8qg6uVxcqBCnGjgAJgponYcg56zk4YPhBekVkHKYkiYqG3zTwDDHrJH2w+D9VshqGeWy
5BPui6an0Xw8xBUSjjptLp5dS9SmwzK0k9WUXHFetmyOJb31mQjyJkWSWc80YGRaZ0XmpJmQxITI
Y827YfAZ90v5wpXF/62UPlpIkeDs9hoDB4HmQ1QIQgRSql8jPgl/9tI1095tSNoXwITZ7zn4A00x
foFDPfkpRtgcOEn5h5GC9qPsm0s6UtpSkb0WeuNPjQp7wTyTXi1Sm32nRuCjO/93MJKr1ETswDdd
B/xO0HJ6BSinwpgvDJY+l5NvsobvF13bL+w+F9L5c0NT5spKw9d8Rk/IPk5XgQOowI0/IBs4PaUB
QuogjNtQ0lA6ifucOS+orNZjm7tZzVolGFZNAd+B70495mKLhLSFDcAhDP0gcUNh8bSR2mODPqDt
DZpmMY1fFim/iHKRrX2gCy8CPiqVtbAqQhMwJ9l3v9EpoesuQJqNA9V0ctDxssOoDisRq0EJ9P6h
Eq6jcslKY1v5j+CV07Secum+sSOupZWWHSVcRle28M9SVX8Hwtwf1qLHp3MGhFiIQ7y4/2IPucCO
gPY1VQsaySH+cux5WyYlMsh6hS/hI9saciAwKnHK8j8ic9iZ6O1wzrYRPsA0d11OidcWe7W9k41x
Y0u5ZTbZI2Hq+kKNDwFQMMPq/YNqSMKR73s43K1yvU0l8c4NUovRlkXkB/a/J7p5P9JeDgT9W2f4
bjxY/Agtc55INZzvjpGY8o5xjDpw9Y0uTLfsDtEzwV68g8uYsrUjEDQbyUH4IDXNl8EUSX1/k9V/
fsZzPpYywl8/S1kO+QdATM6SGTQzWyeBSR4RQc2sZkGy2K1WFhCZDVclPIj8qrA3hTmtgOo0ztla
g2v01usu3cyHzwRDO+F/rDqGbgFC31tf63f05MZguIQwlRWIRJd1RqCZM6KXGWLUOMShqC7fW0dd
eD6L7RSNKamVZ1NtaOUOlMCs2QctjsMz8MoK75ZAXbPKMxXqQx4XStNMINKAw7VxW3jqZmuokkrh
6yHp/VGAX6xU9XxgUCnhEzWOdl6N6oJKnSlOG2SWRVAvF1SschpPSqE7IbbeodC+t9IVwz1iybJu
jCutAHUlrGozQDnqbzSJVInNoAnlJxWtP/bxMyPczss7rl/8cdbKtl0zr8EGCwRg7immzfKGkZZz
YwtloDVM7cSt19menV2J+doKPdZijE+oRf/4y9tghv7KCgqqE5Khr9/n+91sFj0mIjAGUfVzX0wO
giAhvlYDQt1bnlRmq5SAhlvQsWmo5o19pc6dUA/zW2S4rx97q1Vt/b+5lvsbbeaVgEzD44r/p/zR
TYUuxuM5YicCZC25TAt1N7tj91BerU00GHyVQ8quvs/Ib5GpxaGNLzz64qbzVJjdGwCztpegG1rr
GhpksLwJbw1nZ9FaKeP73rMhgn2eTuZTfF+mBEROrWD5JNi3jabuARfKGnmwvlhZtLWjFBBq7czC
qbGUmXdF8WPDUzl6tYGOgwAdmNqWp0DzMAc+Pvm+gVgC0WwI1Upnf6TgHukGi79c5sLnkKsao0B7
NDrcXmNqtLNNVB9p1EhyZvJkld5Ghjc0nJCkRqmhp2Adt2iDCTmeLbFwgyF2epDsxBMAOAdcNEVS
LQYjwlrXeeYfGKgnNUd/8/P7pHJYDduFl33zfXR6L21iowRLABBuw71wcCgyopu8lTmhTN85NSxA
EklEpXvLlCVCR2G2Ovoyd9IRH2Yaq9a/soKMwdo1A6hpQu2BTdciGIhxs32f8EAQwAirdM3ZehMR
ZPiYb+AKMK3Gi55rPY/IqOjfz+w2gButkOGyPx0e4bh3a0W+yKigJKBWEBlNQEkYFRF1SDRqN5rf
6/InN7IGKbqZjm1/tNZQ379nyg1OYug75iLxx07F8y6RRNBo49ZDueEUaNE4a2vCd5oPJWx17GDX
JcDzDHFc2r6TNfA8O+nLBwA0hDMkqcV1DxXMUblf8Vy4sPjf+w0qgd9kSACZp+qIE7dgF/Md8kWn
QEJBBivZH741LAmckalGbQ6N1AVaBc8DYaWqSfh2kjaK3qjcB52QXeENEMTH5gKviua/nPcUarY+
1D6GadjVaLqWTSKmly/jNpWWRXx1GK4Uae42TYJkjpueiZWpcuVWbjGnrDmd7mMNPN8hW4hvB3ea
z2kG18fX1eesQjAdqGS0nDv8fxEfcyNe90DZFbhG2yutLcoibzeioumGtyx8n4qTC0q79mU+0Eis
98v2PbFeG5SmHwehykSwYqeJAfzj8DI9mZwmdgljFezLNFS+K2rSLUnRHqf/5biOmyt0tRye584Q
RQvwSuMN1lEXoa+NrnZZC41Uxae2urOho9PGR3ymxJw5s/pjX8tXrNlZJXfEgKB2kvzMKdTP22w+
0xwlYfQoCK0IVRSSOI5eitQz2lTyH21ZDKLsldXL8dtcdSjnK+FUFFNehLDRYe0RMdD7ZGFBrRxd
XekO9lukzEaEAYifzhBcHMCCd2s+Dobf7bFfRMpDO8SRinXR9C7dx/BKxKPrCCWdSSD8cJLoidnd
iHkcVEHYorjXM4lDxd3ypGT93hOBPcCwpfuO16fFbHdRyqkuoJPfvzoYu5PSnoRpwQbYtK3TGa+l
6T5OaVJTujD9om/Ug1DC3I9WNp5pF9EK2tNl/lAmo/2Xcj8G/ysuFYHa70yA5OIJ+yZ5QfZNCMsu
mWz+cy7LHAkesITtSIUWHpVMaUeiyJVj4y8y5e6+RO7R+omqxQp6m7vkXWl5OSGTgR28xRt11nhh
Hfg8UXvqUdl/Do5w3o2K6Q09C6Scb95qJtmEkLHpS65oY+auf678xix9RrDuNtkKLqiNAY6snb8w
IDq3u/Hl4xlrsKqv8ft5jWkh0FvNENJazrse9dVx9AhymYDETUefcQrB/IcqutjB7vw3+O8/zUQq
0POySGbtq70IJOlw6eVcPqbxNsPhm8qaA6cEW40bRsvWC4JRehLNBO8gUpYa80Su4T6OeV9A4BWK
TASx5eP5RI+jHpefAztcXW6V45Ana4gSD1OlvtdfuJZDODHZQGxJq2Sw61bxy2C+uby8tDNNuhnj
ztqD+/NodK0zJccsBB14e49FE53NKPbaQMmjo/EFcuPWZkyAnkuDg6vIldCmYy7BX9FLJVZCavec
MCxpz1Mu7pQX16OFY4nosG/9BPdmOg4jCrETNKs1Q8R3x55gq6nuzlOIByUlxubqqjAfHgdc9R4W
DAjGh7F/QbI0rGwmU/KWOSukhrMKDV7oXsqm40WUnTt9WagnQT43M3H/GJJYm6BIh8rK/PywtiT9
JrYi0ljjG/+lo4iisMA82Ffa+fH3b63cfqjCjFyo1zTYiqhMcOCit6Fm60cGRgT6atJmw7/xfG9u
SqpuGjz3rUnZO9YqdYg1SAs6829Gz2+XuZMoAIQ7zBCSjnnCtcxn3h6As330jQAIpedn4t3XOoqu
zSoC/Aj/hekc7oEIWdWz8IRUXMnZ6OLIEMtEGAu7WCrzM0ggq0JKagfM6EMLiBsFjN9ZcI3Q27Mx
nXTIaY5xwhycLfw76DTZnzf7+g+41YJFEHpWB2kZ3h5Bp/SfkDquKN1k/0Uin8xTM3IdVzZ3PNWG
B4U01C2Y4bXF73BzOSY9r3VFsSEkiHjdHL8VumUj5sTaiylPLEbUvXbvFLg7lohkmTmKXXfEUZnr
q5cBI2mFEQqTrR/v5Xw3n7kjeeWo2apNWcr1/7Y2UBrfJYcXDJviIlI4rGsZQcnXeDEhqjEklkma
q6ErqNYn13bakHxqTgkwhuVs5PLn2PcMM+Tjpoo7XcNfbZjVMl8il1bKjVUETWOoVIYF7BGdduqx
cMQ2Ubzlj/yVlu7y5BOWv5FC3JpTwrOm/m/XbWWgrg3EOReHy3kZ5Lc9E7ZxE0j4sLljwtA/pZRI
NsbA0qIHaVWjLqtIb3C7u65Dm2doFrVn/NIun7WAk8oF4zpJoL2Lw1iucAMLyjb4WBFymvlOAVLh
vMAiIsxEznAZWyWOrIn6RIKlV/nE5JeYhsNgm2+QGn/8qvuqvyRUCrar39vkWG7Zqhm7jiPxAb7p
Db9Zwxpib4X2jPPqAXHdQO3ZrTof7eqy7Gr2EqhRBAzXdnG8KiukPcMXWI40Rwh66L+jo/6JOi2R
8TCYPDYfpEwKolQ5HCqU/71yKmQWOqlp4TgLvSDlEU4jNgdG6argIRhotyXJsXBJMBek/Ey86YSi
HdnkQ3rHiYLMeJLQYUCgQXuporv+nuSjFHcgyvDT6UboMZXN6LZnDMtdFjZ0a0jf+yVM26ROGnAf
uO2M/pFbPHDtoE2dEj/0P9LpWACjKWN+HqzyYgcNe0501ZvtMDZIE4EIVUQjSfTKldllGdk78GvN
hHC4sY07z8eabBsPNgrNlkHBBdOjcuPg23E2QhYaCDICw/Ro8edbtjK0dlVW/SptkL2FuUlBuADU
qCjrz05yCUrV4i7Khm1wHImqW5eAl93qhSScGc76zJsko3TAm1n7MUZcQAq/etIhyitW512AXs3j
abvvn2OMvY2JMoN7S42sWLQ/4cwpsl8vsMVfnWS4IE+3XVRK4c+Bp/Mep631OtpaS6VSnKpSKMUb
dPNCEVAy/ozzh1M1i5D7iCMaHKwXuAFKt7sVqnrL/ZWbMMAI0GQ2EHQc8GoZ31hh3Sgx8PMFC8lz
vr2deCnCNOHEh8QFUmwG5X+Fsk1ucKqVs4EzwHoFmwyUa2ti0yTz5oLgIZUmR1noejIxkSL8ZFOh
OmrkmavYb9ScjvEhVnsZtvLrgyQe8mC1k2ZIUgcPEHm4RVl13zZDI+O5BnKJ25nuda5EuPUbwQf1
nHX54gbI9zApf9yaRm4YivlBbKJjeXxUbWJR8mDeGeEkPK7tPpFHM7Xwi6Ixfah+2IWAZj1a/rjN
b9/7tM5Eoo0SC/nyPSd01N3FtIM9MRXMRZybDXwjOS9lAphfv88o7SjG92x4tG6SwtBRxBhOBurb
25QRMncXqooAaBfxfd4Bn/22xgdQ+sKf+9nHERaG9gND02FaafNWDwi54/Kr8a8nHtv1+Zjlp0+u
Vq6OVhSYUcdODHCouYTpSLfYY0gndsa/90+enlFeCTOeWltf2B2whDN/zT8zIanMH03gAXqzSs7y
/nPY5KzJbwoj/2lg8i2fCRgBxTEmmnN2TP0ypb3Xria680HhHTE7cFnvgo4DOi0hQPxNyIFrq3NM
CRRE3oR8dY0wpz8lH66lIkKInOLMywsYHnUKOaanp+f1ICotjtcpW5oiuiIGnoyDuxzj4qdze7RC
+bHZVVAK22iD2vDwOG3TAI3H7wHyjVbnys9IkcUL1qy3TW9a5APpzgc+U5Wk8t0vKWzs5eGLyAiW
FTYQrpkr7dwr9hGM+sR2SdqhCSusgggnPpwzb6HWyiF1G6JNv9bwxdQBKOU1xjBIa3lKqhidjEak
L7UJG70aY3j0B3uB/AQEv7zcWMCs5Uuo6Js12qTkDJ1zZRwPIwP55AH5OQ9Q0i+M1XyiOOFW+eBC
wLatidJGZoetYSH2J4NpCGFUhu1quQXq456oc+6SbZAJbJFJORPpdtwjEoBZWPIcBwJuGZ+/pgm0
vVha5NlLECce2C8vVlVK++IRq4+rRe5LFdFrIJNriEqMXq7e6eK4lVlcg8ISAR/Wkp4MXvri+r6z
obn+HYPeYGL+xQ8a8Qph525QghN3gIncvVk8vWgRtxS2La/8B+pxbQMIfaY7YsShs4wlw/aRMCA/
SApcOT/Q8XxwkHgEg6zwQ2WT/SdYb/RyueMZttGY5xm0pgSWGPaOIVn3Jrzo3+tIW1dM3vvsG7ZG
TuKi4Q/rO565qY5M3XPM7bnq7iIUDfvySbbIIQLp0qF71YhJmPDvszYtfKHO0FEfKy/dAiV/SDdh
gtFkHS1SRUfm+mYeK64PJ1mUVeM0dZzrDi9xA+RNSF9Rw46gO+LwDOUMbQKfYMC1sgmfuJdRJZcv
z7KkdWRjBh4xz4XIuy0J8+gaddFZe69pzmWwIGpId7xRIezvGONZdHZ3uAxCftVB8TPAJA69TZVV
X5HwdRPVS17++CVmDRe1ZsZwbhRLbMk3Ivg8h9uKC/tEDxg9fKknVMcN8aHEVa5AtEjtzliGUgw9
x1H1VD9RkicTz2uXfwOkS0D6A15CPqmwqAPHvRi0whnRFzT4C3c7ZJpVQGr8dOsxAmDDj0eM98mO
d+b6Bcw8N7utPFcBwNHFY5vRgBo+V2G/6O304slAvtC9ZxLk8p4Ij0gDbjwAoNa+mGLpwLsT/wKd
/ZMjCw0Kr9pfM/oooOGK0W8MHS82d9Ih99KQwjd+0wTfdj8IaiElDjRzMk0z5LTtLGfBBvzFeqVO
la53qbttdx/OQcVJQGEvw0oL+RtkalStBez0FsGH/agAiErftCwIO6v93/27xXPCqqJzbjbN+kE7
SR8tQzIBnSG9wnQzNATBiRsmiIQr5N1FIZ65BRN4JCDwptQTSfjYBGmjaPsMOYjtTu3H4Yc/5mHU
SafGcSK41b3AfjyR76DiIHRZ2V1ap8tUPtBc9IhX5/A4mSbaFweN1zvoycgyDngIUlC/YtlcOfWT
CTBiTfQxV2YwL08s+INRMI7lZS+y9SnBthnnUy9fFfDoeY6jsIlq/RAzTOwSWoYjza4CxHsDIP1z
9BJC59uavG2FZORd7jHhI1KUgVL0HqiqKN3s2D21/bnmNZRdKZPiU7pdbuh4knn9BwrPBOTJ02vs
aIHzC5qq/6ii1Kme5vymgVUPYhdEQfI8xEM8LxkkgEr3bybaugMCmHuUN46kD+ErVtRGM5SSkq8+
BqWkL4n+wbIkozCK61prCmevNXQbCX+lxuo0gP0ulHoSUmIXBOri9GjPeY8euobzbeJ8Pm6yEs7v
Kb9KGZ7dvqghYLHFYg/NP4B+RCFvGgjff3Bx6QPl9vqJx2tX2KJx46Vf4498NR7VNFYHQbmDGQqS
wjBgc2tcxqw10ZUmCPxer6RIxs768EKw4ZdJa/+awHrfnX3E6uTM/CVRyZ0dOuBkeL+u26FP+zBa
nXHXHY3AlcLSBoFFgymUgc05FSuounz3XMJ1AxN6gm6cfsHLJvvgw1U7tryflF0djcJWZz1c7grA
4ccJQU7f5yTqS2s6kNCA3oKMIaTk5+Su5OnSFHajrazcDuw0I0BlOjDw6O9HdjCosBnC5CbDnJrb
Azo9+XP+N9Qe18ErEO5GpMK1NLr9JPUQ7pUmzbaEOGzDIPQ5o3ItHnUWu0Nw8lXMyRybDf/feYKy
aefD8YRjAUmRbrEkBLHOfE96jKIfT4im82tXccLYy0XdmLHooL1hq+MRg4mCzk8thXj0qiF6zLlN
rOQ8DADbnvlZ20ICvl1Z4rs4GPnrt+dbOaP4sr/IXVGPrGsjPv6qV0FU7j5tedMZLaaCXpOiiZki
+7MqN+1iHrICmz+44G/1MUg+5tdFIVHnpG9C5hqayrO4vC/ZqyqmOlyUMOLGNrbdoWihOKCL4pOU
AZlCsP/HFEQuQf6DSy/nPySBC3/SYjlJreAJYQgvOvgu/gTQElDT6qPT/X2/c1+Ku0lu8LkmpWM8
YzHGjkc6NkNehz6G0l81MrwI3j4oKxjaKTilYh+PfV7IpzBcQJFDOR5xDlAO0XhaqRn8UK1Xad77
I1GPMo4zHFmybjQ0qcl7pM5wB8Kda2k0q6NhY+vVcB71aSllfY3i1NIcGwuYcu46/ikvZRhRljva
yH7m9mMNTPeyUig/yUOE1vY4O7DGv3KPJUtwCwFZeuvEcRs/58oBvs1ncd+Dm7nqLIpS6Cuz/SNm
IPAS8hFAJU41fVejPnuEfC01imMPtsXqc8t4yV0e06FjXcWBdQuCgEAx6lnUW23P7ZZAgSB6FP+L
8Ar091DHekiyNozhSEcoVofPNBWWl8fSxrH9DrdafsEv5qTylU3OowaVRFqX9vSzHL8dE8q+pAoR
hBid+BIBuz3SfPaqcVE5vv8jHOQCnc6PSAznfTJFTBseEqk50Dz7MnCayvf2Ta84MprbPfuU6xI5
ylj6DI/1GXmXXApWa7BaM+gbI6I/BQJaXr/agsod2PGEmVCBwGxFJFYaLrphZ1hewhFYXI4yBdJU
reCFuhjYChZkhsDClmp0EiAGh0xbFzkSPyF3/w3lIN80SFOYPjOtMyCGw4falr8byWlx9D84s4RH
lV0KSDIFnnz9AwDb4P3o0V8HEuK0Mw5rfqIhZnc72X5DQfaOWZwyvoHYvr0nYgnoGCS2xQ9ylxDL
3O+2OXZooEqbpTi2CcW9oy3eUuAxCxuF8I1iYNB+RRlKYNmQH9UEk6ObDAOYvjjrudkY8y4UQXvT
cBlkGr+wyeb5tsfPwt/wmewzN0YHyvGCZtcPuqvZmgA7ZdDRM3bHst50b1vqJXUibRV73bammeKA
rGlSbqRcr/Jj+ZL/UAlUsKNqNkdtfqCuYKqdQmwdyWr/FT1B2IP+eXgq1HSsTDCqSpZOlp+6De0/
OLaHXXUX4x5IAPCBT3MlQrtZM0zYVCq5VrD2eQgr4iq8IfVwNXVL2pjCm0h+ioZkZloB6CESU5qS
yZ0FmgixJOx903M2XALNopmqiOEKpLNvJXhJ7HqBFCq/pW5nRLFOg5IM1oX3AAQ7iAMrm11+tBih
Qpyq+Gm/l34dsqqbIWFQjvpRM1n9HxixaJW7W14Mjr1xZBZoRdo6kpgPTZL/qsS3/msPdGGFsXKm
JcgQs7pSElp0KPzs02LABG5bH76gNrRoJpFejzzBtRVnh8Fa5XQED2gMnRE68vvImDiLBgH2OVmv
z2EcQrKj1+uTNAK5TXrVo/+zakj5M1otZ/L7yA5/PVDoRRseJy5w53+kRWEV/5k8RphWQqnPLB7g
UX38FBVTUROR1EzsfqjwbZpJvfpC2oqk/2TBG1QQUBoKAMfRtQxxSW9wwSSJS39T7bzmAwV4lmB9
2F5UZmTCGbAzMvZwgWGUcjd2nbMxuW1EEPggOHuFoWjEwoZnD2gqaqWe5NuCbWGEkOngpuXsCwRt
qO7YgaGk9+3D8p/7IS7FMN0JdB+ObCKmkM3vlz6EKZwxcvGmWsVVizyTfc5HQITgWMOHXlWS5QHA
nDuKG6uDAwyaZPpa+KGiaCcj4gQTXdQG6rdJSiN1a67DboTytnYrm786Oxq8HBqQHJvIZAtAFsMY
nig9TRgkbQrr+CLYX+mhHPlRxJyY4NWAU7sEcsWUmGORd8cZQMCFNN43rmE3mRTIeBuBVeGce6bV
MLzeO107CBVo2H4RfhKu5YRPV05oPNRLb0eqs9bCu4xtpx6VzWZfWTq3CcdJ1q8BfWmB0Jzt9YFt
bigMFHOtjbkfoXNNgDjdpM0L4+U+G/+dz65dgvH/fbOkkwOrje+DqgXLg89KfHhOC2yqM1Mu0FM+
195Fxt9i4pBGnnBGwME6P1RcY2K2rmofRdlSTJCPz+xOUMVUSK4a2D4OI7V7HVNUtPIPixLpx5K8
GxReGZcD2gdAskTRM8vqboIsdvfmnRC/610zCOvRCIeLAyUW0NMF2y7np2QvUkVLxHrxNhP44Msv
9qWlOYNoB+OOe66G6HCPCMuz5kWNP08x6w59wquIF9QCZkqF0Qis9ljTgfyi1Xj+lCNK9ZSqSv0p
XcjHyzgp2xDl3u8jPEk5YXrzA9F/LRE4PIS0xJh4qJwd2VBtKwrJi+7Ppd/FSaAFKQ2WYs+qsUZN
y+gIz3ED6UHcbo+jBPSSD9cNsTfFuVZeo5CG6570f4fS0oj5aeEZXX3PRP3/FvMnEq9J2GUfqYOZ
ZUo3pyoowxNW/DEI9f7cbutrqIN6gcjg+iXVvZp6Oatg8Q75VqS0UT1qv79EnnFfu1vRL+P9S6F7
mxYzME7ru46w9Av5xKW5zA0T+g9ccj7GAvzzDksjmE9JZKY+JVoDBqUfDCqN93TnpKq9nrdI4bxF
pGzyy9fuI42a5LC3jpb9VVEnowivXYxSX2ltFKsijftxIMaLlQQhxVGpS+nbfZu8xbpITesDz/3d
NmErU2aWyp4YB5k3GloHfZ0AIsOT8xihfgmf/8clcr6u4oblN+ZA+iZqgqEVM0kNS62O0zuKQUMh
LPecB4wVWGtR94/UKx/SfnEUCyTVbmqc1BHNXMWbOO18i5A+dr9KOSxV40RGlKyzWbKTv6Tqm8wM
KhCaf+rN5k3gjpcbue+stMjnazjXGgRtX2sU3DVyMteuRJ3dEy/WnhBZobgN3aLTlSqeWDtSVa1b
3piH3qEOXivkkKWM4cBkZfvRei+Hp+gGrI0g2pMdZ5kCjt7MileutRUqvbIY9d0QIg7/mGNL55+3
H9Oam5vwinMAa8AqP6t5nyZ2Sji+vJOrzsZFYAiexgiqJR3XauAA+Svu/rHGrYj8o0fCkstdGzd2
DEe1o/RQOtiHsbanbuK40qZfeFwqjaHBpNlhG6QIvLTFkxlzFInvoAoDSuu8PAEGWzV+CQHufWlx
MqRRjRBZXHd8+XnMOQSGLqasnDwwtPe1DRHauiEJupw/GzsloJ9jcTY5N/45HARMutkhz5j6fiFo
vHeZHvkQEfkpBK1nzm/xh7y3E74Z460AufvHhANeUL8U4LhHW98z5B7OPDR/I6HWj3yBj8pBTDuS
/DZL9Fhs7DOUZbvNEHxE9k+khZl+0BQeiMGBIite8hTJk76dqpD3MkqeR14MR6+UtUw5q+JuwgsL
K5EaLEmhiiXTu9t3IpYLHkdzpjJMC1whmN7VGW0iMEnWIMo2OJ5zMPgtUGEg3pzJurCcBnmiJVP/
ub3wCGw3Ba534/Ije2uVP/Tg9f+AnQs3i0KfRYNk30kNZjEAZ6bSzbfyfvLrFYLUtokSvutmD1T6
z1RJpAriNBUtmExWW+rj4GQqz98I5H5VfO/gaeA2jLquZMadw1OvmtVhblnq9JOHJfP4MTwR0I+S
nYEWTiRl7CYM7GXVJucQ9F8Ain+t6CRligushZrg7VqYiTWqUq7FNG9XxhNQCeoLHbyY/CUxZ6xI
mIPh+ySGswhwRhCGC+CvuUp5UWTvMk3jOnlIur1F2t2uPy6x0BcIkydA5apLNyDn27CD0TvPFA1r
Vu/xt/rnQnYaJc/7pB7bmdjUGxIC5JItPDH1O9oVRkfrtHz/ljm3gnX3qrzjsNQIg7ohVcaB/seJ
RrfhepXa94iDDSP/lEKKM8SthnlUn2b7cXXiE5Dv4+y0uCLDnPN4KK1jM+4yDOuABMrzEWGScIII
MEs+0P7cBYiESeXQ+eoSmurqDVx9FXSzoOIOkejsVUBWnRp0rzviC1OEkINDWC+eX8w236uOuAaj
IJX08qHXuRHcJ2W2TyDArscssuPFk9uxhWCefNUnreEh9wVRoGWRsyC0AVYpeWy4LU+Xjrqruch1
xUaGa2qYhP3oqaHCWUQbPP0baPQ77ukupzdO+4fQ/kL+Ot7z7oDH3Tn+3qdpPexk4Eulp0+O3QoY
oAMZWikyCFs3WL4FZ+O09FtpVSTTW+C+HOxyA01R0xTe+KLhoadJnWmHtZoXfxGcnvImPot1/2b5
bWIvzYI/Q3Q88kEW50cAbmsRHvrtO6KsxSJEOS54F7dJk+JRLopDPA1K32d9Wg0n5aTnCTRsHJst
ApmYPJM24DbOX3HYtp7u8M7dskIZWWFyU5KQv1/8MYpxIgh+6vrGFF/Dl2s74jQW/3xycEiKv4Am
nCTC3LH6XPfw1gBoTo4iKKX4H5uz6b9RYVysH6iVUkh+dpKORcHn/r82MM9ve6Xw2JA2SZm7C5od
HBDfkvreyc6RL8MSKuW8oBmfVUhGT9gtQUN/E949vPj9O0ysCwI7ZsUAAqZ6ApWmtnuGMX+vxluh
sd+1Qb8jouqHLF5GHGo1fnAHBiQtjnqHGtwbgEpIsTgvJJYS1cjkBW0gxfR/QyQTaX2mHKI4PWVq
K1syoRA1Gv1j0cxfSSWvsPCsPv8tCPeWzu4pWaSC2pseOZCj8Dckk1Sxt5jSiSxUhJZv0J2XQ0MQ
8OXqVrJvYpBtE17bV7awj1ezXJ5tiwCHKow0QqyD5gMFyoxFFR/6AyhGEteZrzQn8pltttR8ZVoV
3asVh1deB8ry6OFypT0l9XvgzbcYbd1qTTsYF+eKtCQTGhwgv9eSWijOs2JaDiIid6LJ91JSc57M
Rkb4exKOr8prKdY2Me4vw6ZFlceXCuTUJMEMdp5LDWbi0a567VnZdFLDTvJ3IKOSaHLo1vC8ujWP
2sU9hBj2Si581/5z2NNR/Q7t1DnFspY0cfDY+ExhqK2VbzkzeVmIq9XQijQhEPJiRZ0g5AKckApN
QDyNK8ATkxPuwmXemhG13sg+IgbKxPql9vyGfMmBGoZ06v52o2O5K3hVLZC+z/eRdffeau00JC4x
533M+pe4UHvo6zPHhNrV0l/qxo1kmt2Q+EzJxbe/HyWeFuKNx3St22dhCv28ONK/vgcXSTbUTo0B
V3JvDnJip0zgJHfWdgPZubRBl5aSPjrsFjObnUoi0ogUUs8KKxFvJ6v440M5sYoNI/iNBKNtabrh
Tr46o3S8Ae9tK/vNfYWvbSy5DFAGVOhJEfx83RnwuHqDeDvgQpH0MkqmlLgQcAJd3eCX2Ur/IRhs
pWy/UqoVB7G/S11huhl71aBO7/JDDplanrB1hiy0UKEXD8DOGx6trN6G+iqmu72rqyp+YdKKIvCh
0sYKPvBrn5+MUvXePg0meZ8o5VWhd6ma2WgJqoZfLes/P8X2y0bjpCv+OuJmZ7bLLq21xCmGlT2N
W/cuegUMk8JcayBYoCHpNWxGm+3UT0AxPhFBE/pOs2qwYZ1Gs0+QpXy2cbAW1cZpGAOUjUij/Ww+
Fi3PD8PDOMD2W0MppbLUW5tZkYdN0id9BsVvyZdIgwq0E+0X3nx8FdynRju6Nlb/1uN/8TS/vagg
u53cVN56tjo0W0uUurQngLvodnLGstTs/oBxZI2dsNPbVQmIX3t8H/1/KbzB+KWS7k8e/he3ieAR
RxLZcm7hARKrYL/R8I368SWxpJbc/blWVHPawanLRnonW3CSzBHV52BSvUX4GVdc4f5D190/zy4s
ML7naQc8SXUga7prK6B+7Tsm5Np/IUj9HHfZdlDYoa/FyERBGIlqLPPz3ZQ9ZesoALgB5MpCPbF5
eShT2cuosZiM2MedQAl4U9+QxNVftScMEaixPiujN3csTV7dGpWQzfaGRemcvhfBCbjsbTWnquXu
1X0HVRrdCsOfyLVpdedgUzkj/8/4An4CeqAM44lgyxhCo3ZveyF+0lmJyrMr3Mwd5JkYzZ5YIKjB
BCzXMl1+ZhvyPPiR5I1Kfo3j0ah8WQyrMlytMtnI7TjvPX0QC7gcjMA6FgsOZRra2PsUBP/xxyGJ
siHfKSWBzF60SZt0miZhtNPtwmitlGqB7MR/ZNE9DMRC1dkvG43MrUOpNXo9ebHgqleHltmwkw7o
OfKQHuoqKkaIp9hwwrzM/fk1ekbyZvL8JfC7IVVHy/IYaJNsPm5OBgDb7LUJoX53lMHMVJ5sqrrd
zGqXyuqN+o3xNU2n5GjxXYKSWK9+qw3ARuC+2cKkYF+Y7i0Z1WqafkTs3nt9l3HUrkk5DBqd4+yU
U80qnaa0V5nTjK63wvEeEnoHSgP+jTmdtlLEasZZgK67vGmG9etaV7W91hb+bPxSFcf/9vHAEbcO
OVI58itsGRcT53rOqhXxj2H3VlRHUa+owdj5rqVFtq+hvxj8riEAMmekWZjgevTPi/6hsslV8q1W
KxIkj32qnfU3d2viI/SbRotpfUpyKAOVY1YllzQwZVkETXp3Il/2wK1776eu7maDt+tp47eA2w08
FhHZFurrYnwZYmLsv2oq+xuEQ+14hIZQXRZJKf0iCEcH4bq71HM3AdtcxFnIiihy0OXcKKhz1SdD
Vn6XA26nUEp0YR/SC99K5f7tjaeac7zGFRrUhLhFL//t02ixJc6ZRzb2yleV3GlrxaUHmjXnUeZX
oaU+lAv9WI6wkaDEXSvn95A/u2CsthlvZ/Ms3IYyVmg0oFTHQ+Dq8ss7p241I8PgvYfCfVc5lkQT
0W/Jj3RaTdW50BeDbZkrns9JDWN2FYnnBdbmWNsENttUXjAJeGJVEgLmVqVPwdbFDYQx9RJctBxF
6uaf6i8ZI9m/cB07uKloBXWThkvjJt0paptCTZGKSX8GtTdqGg0QlBBo/nVGAXXA7yMZOvrf20Id
iWCfdQSGA1ML/+k5FWyEDTJaHtvbcpYvmzIPWVDMrkYAIf2OL0G6I/SyDjJkZ/fb/Exoxu+f4GKZ
NqbZM3nkjUuXH9MiTWY179d04Ovf8hf1PGLPiJTdkHAZrN5XclUwrrFxiizbulGpCtmHDYRAPr24
YkLLKuTLFbC/hdb+y+Xn2ERxZsGmMWPfIUsx5WxZCzY+jKiMv/heNBzotZZmjUfhTz7ZEbVJenz5
UtMesgmf4njaqCB4h7JxjSmyBus0GKY/ZK4qYRTjEh4gj3tkiE4VguGp351rqf7iC+lC+OvCoiuS
JoiboPpMBNhCxMxwg3D0P2ymp6hVZpQ2jI8d+abeDNnkGNm+FaQcU5mMPBTci4NSq3YTSamJsWSF
qrgeHXyfcgkitnR294JfIzmG7S52/Bx7K5MigAGXp7Iq98U8rm0+ieFKSdluMocOZXmaGg37ubfP
U9tD/mT3/VT/G9jy2MTbHFL+m7bbw2y/IQr3hyp8+XjO4SdcOATVyP2aiY6gkoP/Us0C41ycoD6T
Hyac/fqIgtDlsO1SFelXVl8zr9CikoUwz0Ni7VSwGGv1Z8Ran0dSGp5eNjNwW7nrz4smo4ohujf6
L0JhcHUqF6sJSeWYnmH5zEf83BjnALpkixCckH4NU0X0tt7LEOwDIW/G0fhY2DMvFyVp7ziT6yJm
9KRZMMQ3kbA4zWvdEJfiiUt+KL+SA7VjxL0REsaDFYJaHLnibYDXFq9vnN/L5qhuZuumgBl6t+cM
GJotiD9/W7E6bUdhyWT0Snjy87kUrjmQfVPfC/ptXLMlGDbwNHPDPzsxHEyoQjO8M9kbofFf0yVO
FvHrlJ7Em33dYaRXbLau1EHa99mr3aBNzbJldpH5a0YnR2EfcbvgGTaED61qtP1FAbVPIqExHwcw
fDgU64vx0tgC7Kt30Jmhciy921pS3YYQBBZ7s23uaN77rexsfT5dqWLhNFdkzZu1a2P+hqWCE2iI
MhwMbLXdAq2mnfGXcYt+1Unawp3fgA/zMyK3XzswXXAB0991y/oJpYNWNxCERSjMCj3HiusWSoW7
9nkCU1MkKvektDNC8eiOmLBJtZyDTR7vd7Ovd7PNCrki7EpXG+HFERHqRu6pq0QasyshgKLuzS6K
Z0qNY53vLUvR+fE3ocG82ZJESCCwHEnXY//j7oP7n1Nuu5unePZKUICmrx+9JiqOpYAr9iJuS8yc
rKhoePEMxO4jm9EBCGFXrfsKoeNsjQlaDGaPaymkK3lV4EXzzlazRcjf+lYe/cceM/QNv7V6ZBpM
NZINDtQcLhZMDuwr31rtBXXgna+k1m3zCeIwmT5Li61Cst82vsv6HCvsn6pCj10nsCyXgJg0pD0F
7M4lyWVlYUJ0aCTT72qJgO6bMr4JPKCSromLD+k9KK/pfUMIoLkHO/YHopu+KkiXlNaPk4T7kyVY
dPzqfwOHwqE4Em3UD1nXOMNMCSG1gIATewtxxdeBjGuwolTNSpiET+tC3K/9w4xDf7zv+ZRF9SXH
Ur+AjP6KfzbbcG60XE/ibVNg//fde9SoQCky5+pyZidHEt8AJfaq+ZIwID6B9A5dDxME/B1mUz7H
SCYcAo87g+v6X4nS/7gZz7iqgMiBx4KM3SYSSW59Kl+INXJfXQu2wBogHaBYvvONViHbbfQ+Ze4t
Kn7CnAqR5BlV9gwVXk3jF7g7xyj1YAADXUiIPrtTAAWdu6ZgmfNTl3agqHs55MgByHFQNRKl7eZS
JFPOZNVTrI0MnkbFxFshQEAC/BdEer4PtD7H5gTrcbErGdPDqx1LEnAv4bOU2PVS7GtMSGAIr2kx
xDXptgAk53FQEPImy4vE0B0ShuM78bGQpfigcd/EEVQFdJTDS+XPq4C7f9J0JJHBjolm+nmb64FW
L0bdeLr169h9J9p4VWvE5ZnKPyOx+7crYDhgDaMbCFIvot63iKkgWv8JwFZsH/cCRp3FVFLjhzT1
9XU+ZbGCTjUeJs0wL+2y7AFplokhCr7fpqIJfSMO9+ahGHnoH5JxPvqFDsdbTJGd2OK8wA4V+eAG
o0VZYSVizIDC1C5SZlrS1OEBvofeFraDvr98JMhx4cLYriF9/gqngSC1llwRMBlrSa1LcuiYf8O7
8xOx7vVgjfZ9nY79TZcs2zeybuFQSSL3zEHFAssuSmaSHCz/UCSgc0lVeckEUxP2TeIhG1J3Ni6N
8r6kZhSYXjjFlMbrG/Y86idfS+0dN0tgMGeECK5CDtDOLRHTc9qLWkWHrzxdTVhUBc92pCdh1TRC
0IYRa4xGBiOR9WlofCPFGjCI8is/9mEeyBGFJ/5+E7VYExhkl1folnadDyoGcPQXENWr8NOmmMHO
y83N7yF0nsRMORtAugx0N/Rtyev1eKkRfLYsqiFHqH1dzXyuIIKqYKRnEeJKDlrdZGnsDV67Nbk6
mBTouopKlbK754iyekfdNS9JEdkH0rleaOwxgXDRh3b5Ge+uUiLhHp0ZPbtSLhD7Q7KZzsNvxBEW
oB9PGQuf7xSLazHjkJQ0TedKo4V0auWLeKzCevbqBKMbDmqZHpzFXeY0vje6UPEFikmzAQKrDf3B
jAWK9TJCcn+PjSqEcq41kJGC+RUe6ay4DPGcgkH2rz8Di5ZdnnrrwP2pmsrX2+cANwKDj5+3vyH1
ftAOk1TYa4nlXsJFvMFFhZCHGEOrXN3ceBnk8YfHYVctCdkJJeoCUXg/N06ayHlzdaHaqCcLAoYi
f82JAwql5fNphItpPrDxct375uIS+2pzaYY+f1IVw8vpJ7j0Gja3QDMR+hBzFNJJOy1DaSewAUWP
trYhtLM8y++hPK5sr/NWbzjgxba9TIv0v90BRT+3pAegHaz1ny2r9wACSiYGtI7vJ6s6FRJZpPAN
yfV8ZRIl0V9q35yXXb2kLGIgMGJlInc0HFm2BQR3rCWNy34mtLNuB+OtWv3tjhkUqOUvxx8amssc
wh64X6O4qE8QgMZMLcJmqIomkGXo4WNWoy8muXP7Q+dyZxsX1EbNsXMr59UCeacMkCCr6dHdRt06
M2je3cxXELxa8UiRG9vKQLBvfHfGf8IlyMajGun2NUAmGtgYjXxML5bttiBTYHllHWKGywMHDzpJ
182WcOD1XZ8s38LBYcV0DiQGi5PkG2us21KeBNArr4AC3OVDWmeXvUIrcUOmJMIVylMaVskIRXqh
d/7+I7Nj7w3v5YFjXLVArjJrs5PqNUVwp9owq1bYV4T+gWsxb5TNkiDRBLvNK+OM4vUmbdGEOUkn
3m6/rpzOlqe/fC8uTTCrFpoRYcLk+TjUeQy0IIR1y8rWIJ9OwsHz43O67gmn2kaWmYGBORvBkUL/
IKJ9J3r0fj9lX5tAGf1Zm/l1HoydN//XKblqoA0Blamm5Xy+Yh4e1oJJjA14KkEU1mlreOy0Cj6G
XnMP5GLVio9k+agAsoU7E8AjodRe7aEVzePTSlRZzGFmgpag5LWiwS55PQUElOhCmuPVXk5kHTrY
Gn13HV5JeFObkwTyKiuNnw1ilOdPVOH7q4UoMxswZKY8ZvO3wRRdIgHFUwXjpl4WrqyOiafy9++u
xpDog0tt0+t3+0jAOfR6kj3aN1PrWZZJZiWVIED0dOIu3yR5SF09S14hNc8mW49A+1egj8BQG9C1
YfBmhFG6Tx3TIGcu5bhqXJS8nq6fTE7hSQDLtlaAXCLk+FMdMa4yO1dTEjPsGGJHJsivNIptbuBh
aorEjPTsFVXhLEkjRSTl06agZKFKwo8xMqn0Q9C3lX9yMutzepgCTfOEmZAI1XJLD0Z1kKcwJgxP
xo6Lk1c9YzyTXuGlNGFB9PYWnDnvvqIsYJfW+CBNm+QCqJlTfCBkKfBPZYlbshO4ta/+ZBMqtS0o
ZXxNUVgzaAozIo63aaQhOrDbR1sF1nDLKKap1MWkn2EQPnsr2cf6A5/+IgevmSW+dRQGEw8DwLjN
wZgp0H9AGr7dS05WQi0KERijKb0Oi6b5ekAczHiFVkjz3l9YqbDXnwntwPrmzButX8NyG314qVop
8YIqvWI7/Zemgkuqjk6GX4QNA5ntj6P8QoOGZ91gsKzqiMOlzLAHbZZgYefELJX62hNBMwcjdO6H
g3BbfQBaKYo2Xjg6O+6f8R1NGeypeXRaze3iLmw392HyoylYyWu1DpQWJCdiumP0UypcZI9xIk+j
7K8woHLmPjDMPieh+CUR46YHw+ofaWm6sJAqCQDPuOY4sjgjVxgRDiandju4eY9YajKre2bslDpJ
HKb2mQWpOdfLx6TmKMztJTRkoeplcratr7OPkh2W56FIWiiAbw3tgLUCmt/afrVRk2SQ6H7hKU0s
OdcDVgptHP/nqBwCPRs81HEVPHe5CxDVFPhpUOr0EB2CctLfTCPI4WwH571BkARpZGJbi/EptEDo
SbJ60cDcV1sbMahgs+4HZehkx9cQIex9QFckBmzJ1RziQ8Ja70FBXI0pVGI3xVsFHftdh1RGKrfm
sKEWvvHtra4DmundQp6Id8ZtS3QS5HEwp2PT798Ef+CHfB2mfYExMijcFiYTyRGbIxK7BSNNxB/o
xrW6qbJKg/oPpcrqJfwpzyv7LqLdM8GpIvBdZYED0ohTnWnuS8+x5WN/e7sZ+/ehFbwglyPGATEm
Rsi1ZvdynRfxO4Nwwf4LPpwftKxDQSWNvODPG403BRYntnosef56QiYtXLY/Z744tbCxCscX3cip
K5Hd3hp9TIFLrvbfQ7ZUNxJPaaIlohqrqCT72wEKA+N5PJqo+ncO2buONqlj73SCzWRSbz8O38Gj
kH4sydlSNIbcCBfhdDOxSFZw+HdgwJ2EGAC4pd4RP93EmfRvjjZ+j6ZLKne1P0r2aOhsQV4zPk4x
3AyNMAef3o6Sx0JmS8d6mS6DLv0Dsdks7tAOcdEef8LwylVwwN54M93zUjESwMRpYAEWIuO/Llri
QX0IIvklRg5xuwr+K23Haxwd5SpnfckJ4a5O4powId46lgnyYgRiszcJl65iBRTkxGfeB6DO+GbT
+sbgTqryvLlPVugwF1gUdZPSf1dTz5IzCl59heKkjbZUEtiUm7rIjnfpZb8Pwuk57d4RC3pgIStT
61aaQ2APorWfzytJC11LpIF2jP9fm63r34Cl7ypYHJI6mqBDnKMcmbKtTwGBZQhj/PwiK1jXC8Mq
kNAP2SP2R6YKdd5jVia4uPfoaO6sMIJjXoF4g9XABJOlvWAj4tuNszuDGeuww+4aSjMj6F25kMB3
Sfs+kbnEgtY+W9QbB0IvOuMqaiwBGCqsTK40rtlucCeb9eftNDUthU91CRpFiezfX1Y6agVPMqCc
HbC78HC6TO5ckRKK5WJNhTSmXIrURRwv0aVyYfNi14vNyD/7Je32vWbOXcjWuO93TUyZYAJJEWGr
RHVHJJ2/VtHhTngb0zFGWF2EkJQfvCZLCOZP7J9VhRxePlPNOdqWuD5nAWJj0we3NvhOg5mi7Kaa
Nq/1P5D+ik+QB1wMwf3FzT085Q+ofGVV8urLrttiLlbDNhH3WB8j4QQltAA1dvaC4sZXLVoNrtO5
iFPo3hdM1fCMCepBwysXqiym4RzI5OmGJTDVQAmqLnIpaMJJpi81EtBw8Jo44TSj/uW7hLvLpXq5
Om2vljb7BSM0gS6sQybpj/Ddy2DczNHicgdiNisRvtvzCAnz+u/mo2yBOBi5LEvICG2PGjWrek5c
NZZBfpG2uS+MywE+T/QhXiDVg9Gq0NOk0H5ZrG+vL0kF84pet37QOJQ2cg5AMskvpNHWmcrLAPBC
ZUSxewlqYe4a9wAUBiij27fr3P42C2k4ImooZKx8vxMTxK5mVUmVUN9THMPCdnxRB+dlVubyozQT
duldqUnJGNw/nncIO3fVvxeupc0Ym1qOh6282ikGA5ODMy7cgIOBq7u/o7P59KGyCSM3QNO4ueol
pVPVyMdcxCehrgQX8XBU5/8dTzPdkOmr+K9NH9017NZ3WjEhMYqpIk/uOkU1WFqd50yYEOI3H792
ib0uNgE4lBSpAh+Ai8HjH36gfxnWiaruIV41p94WzQgxSCa9p21FavAGPlSzrp1Dtn1pSApvLAy8
S4NDXpEOrjoAtzzXIFnWtpva2+je3oxOg4FJfTT+fSmdTX25g5sfrNvyfvGUzWRAMv0+c/WvIMpM
1c1d9iBB/trtyw+U0/G6IwGrfSOpanA/necuEE5BJ1/RtyH0qHSdhz4cDauoTBEahq7nsV60rRlc
bdC45KZP5njh6GP0WlRgTnJVYnI23HzKQ6HvResEBbN3YgRtQ48NoBbQjQsy+ptU+CyPvIRCt0i/
8YOJeJGMWDABjNlwF5+80jNRuTfSyzn9hnfbSE8jXeZI+yNhdvRYTdytELa/CScJzJQDc48EbcXK
zsGUeohz/2wq9tNoMPFPLyaCR/xpRWLxZqNmIhoUjWmEcRD7eB33KrjiYguDdKlGu4mKbyTOVlqf
mS3SymfzJUoOEjaYm+QawE0/fIdgrq7b7QeUjJaWwYKX9bqUX0NabPlu+uegS0vnYdJLItfH3N3d
TuzY/Z3/UH6qUbwI7FjY/DPE/+bPr2pfnVrfA3JyIAOachByOQeGWj0JMa+WHDbRL3g7w7Fw9x25
LkZcyTetHc+g+VO08enup20Gnt/BGmvdCWmuk4PV9x14QHvtp2fF0zI3dC3dCcO9InXJdC9dX4zI
rVRCPdz8IIiYriYFyIpGKZYECUeL4glUXd25KReCrLI7VQGZKy0SgX3wJvTeM/F220H0d1uSq2qD
BCkLFL1ev8OQNN9fkORy6TvmJavIYvrQ6Jfne3ngTcf22SDXZcY9kvQhhyKHTbQJWol0GcEGW+SU
iI96CHv7YfFAVZ18rcAuV7ePZ1JEYFolh42K5ht5CJZdPQnsgPzQz/SNobdYjDbbpBvk5uECFk6a
LRNA6ZuJLpAGp4wfiX8rOaAk9uqx7jbl5FfBUnvIygGXKAqOHz1bZFBcMgHYGZzgvnq3HRKOd5jx
08DYs/bYQ805LJR++xhkuz0oj3mpv6sSU3kHgPLpPbIfTM0QDG6vLa8h0PAP9tJommaX9qL0Q4so
zPL9WF0v3Je+g3jOxs7ph5yI4qtpq4GiTjzafcjaykFgFX1BFD1nqSKw5Taje83rmRJ0XPam8i5k
iZZy7nNOFsVi2sa5SdaUbp0KaATUw2XMpiZqVWD4RsgGIkPCAClUaXHZS6B7lRMumhN8EP89Ap1F
BRQt7bIXM7SuritWLL9cXWg0smfM78kB5a9r/ZA5Mp1Ehatq1MfX3ayzzQG/2RAkwPPg7pgdhMPm
n3o+1zqaZ2f+0Ubt9Cpi0yg2Beiyp4UteMehsnRCOFrLq0pKCvAw2hLksABjybk9Vcv/cAFw04q+
YXjlpbYkvI3U90Huc3AcERfcGpm7+32o1V6osn7Qo4Gb9Mv/rXK2Ue+omSKflYqorIsIxd8nuUH7
d4CMoeMHacg72OM3BZELzniMKf7KuW0D5AxI0N4YJRBSBd/KahE8OzhVm5AbVPjrCQYs+9FhwV5w
eRvDmOJpstGA+YZJp5FyTAIKAGssSvOEQWn3FKhQZu+QQKg0iDviaX6/iYA624diA+ZOqBFyaCT5
VHcmtwlkw1VgSc+QbgJ9W+8g4r9d+HQ7Xel7t6by8wa+S+3AaxWNCdmuuos2zvvYJBnBYaWTuS66
iQeali/mIN3PffM1SSK2znycWXqiFvmVpJS746EbodoBJGZesaRVit1PS0oKRRQo3JrJTog0aF/n
8iu1SNlKEilHhBj+xLQlNumPGzC6ZIRMzekoOCnqXfZtpsunzRRTLnnE+U1ycBTNstnlLWNS/Ig5
p/S0J7sJ4e8ekDJiVJu16IlDNHmMCtSuHO5tYhwI1H3F1d5bFGvjuCvvRt7pRO4Lgj1emA//gQsB
UD7+qQDpWxWwS45SpZwcpU4MP0BPrbrO3LcReFYqIfOMMwCXEX9ZxHHZcPppNGWUIgMDAcjwOZmP
Ffk+oc+PKu5IaAsWlL0xTHRLmUTlCYIbMlJKVGKL386wZjevd69t4orqDPbWXnylrlbve3Uu0zkQ
D3h2Pfu+lo4aQBoMAyoX/lnHV5yTTI/epD8GvYU5M+VjCycnDCr61wQen9H5Y/mgKQ6zjyILdEI7
Xj/0++6tq+w22h3dRGs172Gsh4hQcUVy0paaQWFakY26F57GM/15xG/D7ilMd8Qm16NRUq0cESuE
b0HFuAV6Pq2mtapAuNVTReuvXpmyWKxSLT9ygSfxbZzVSZ22dc9bwcgTcvUF0+USo6GGSTt6sFoR
IYWmYD/Gv0G99Hj8DZ6nhf5mYmAMdYM0Rvz1MfUyLkeknF4KmaEHXkCl3x+zT9Nm5lPFHZI+gwPI
0fxkMGMZquS76aoXWrOrvJsNW+tibUgahefcsddDlWUJoQl3VnXp+4jvnWKr1N9/dxJTcOAmQe5O
AUWamx2WYwGwRgYYkvlMTbVZW0YFhGeL53wC92JUibQzSMQ5pGJIvWOPyT8+jz2MoGY11cUpvbkJ
1zJfeYmW2lNfiDpkNB46T4zEZXoU3L+zM+ZYOHuVutqZY9/9XrNSjNoEuT3EYS6V/kLdOZQFJVjA
KFSDal7Yt7T0ww0ozsJG8rW5/gN8YQ6xP1xh4WJIPDSK1SILssz2QkJ2mmaP1VGDIHbIdm3aR8IM
qhBHN/n2iDHv9acRCAJlZleAh1ZOPEBbvbuI40l/0ddGzjCecPrX10pfUgmiXmfj8MZDnjgam7mv
Nr+KW0jfLD4QFsrQtjUOOeNe1T7eF2ML9XMRJ5bh5FSdUXi5GoDs8q6NihIPEFAHd4Tkkj5XeQeT
qQkJ/K8kh8dNFYvj77VrluRQAcxBax2PrhgovCUUdDpQdqJbJJtIdSnqNbaqY5xHMHGFvVmPH02x
BxZKOAU9s8CohH16cgjPIs6ctvyhposSmgHHtGcimdigz0Rl60WKiauvvDLKgPID1wUcKWwbi4Y7
b9VzU68DTaouZjpeHbVBr4pYVKQiu7AMFFD3XdoSixcZ1tsu0M11OAFmY/UgQY32cX8SyX90TCCw
ZMHQi3nFwtk3hpd86haIgzocmFokTROTLfI9sdTd2e9m35JRt2W56lWtDTX61+d84GAVUwrWYdBR
6xKfjXddsmsfJtwkGst3R1Ap9Bi0Whj449Yse4kxBUDG+iuz/cWh8o1CoZCJVFUx1m3J18+1z8VN
R6TczzqJyJ9psfzF4SqAk6L1Pq4Sqhids0IXVGN6Ie+vmc7vGMmZQWY1hN4HkTRJTLnRMdJHCykG
uYP3NUSdknY9g7vvZtNrkwiad56nhQ1vCIoh1R+uT9yqeMvXB0shwHnRvuC2klPWTs8Q3BXwSwUS
r1DrqH6SRTW9LJwSPWwDl3Pn9DLj3yCKKcAlkCXUJ4Dpm35v0CgAMW+KqZJ/aDKg8MSZIayDd+qx
WeMnnOTe7xZ0Lbih7x2cPxb4zsw2BKXhYjDqTHQZ2565QwAofqpqt/qNwhKde6siMHa92eZVxATx
bTq06+7v7/6VcGia2HnSdU8L1kgjfNzLitZ53Q20NOUue6Yx0EcG2t/QAWE/1pGG7PRO3hVYcGmJ
I0CW6iHN0ubZP8dzXDEzkOCN6pezmKECUEjtiuQ9p+rQE7giV6Q1+YMvcuXGTl825Kdl/GYakraM
vbcdnKpbCwy2Cj/H/pAlNHfo/IaKwtkfvu6bkpqpYzTnC4mXOokEdC0t7AYCaW4j8O99V6Z8XcDs
OQeyHz4CI1XxE5RIrVLDvuetck529AKkHSe15sTIYwhjf5cAL+rIE+h/LcLZZDHfM8XKdbVJ3pEh
Q1hf1fX2SctuUkYxqeays5ae2jr6wR71egEQPd9CtEK/W3z9M2urZ4qI9704ht3OFrFl4MXt+QNN
GsUZkvT6zBxdgs+uxNhhVUY4vPD86vERIHRZEMNz2XSWu6WfQfRuFGj+iIJYANsbqfAliG3H03bh
/L16sNss469ccfhrslcJ/cKoX2RkNeMz8VFzytwdBQabDPJ612nZz+4UvvZA3+z0o5oXwSk+yUlY
nYF7vTNsu8KvZioQQw9+e88xFh3yYm9orsZ3KpGqzmTo6Kq8RvS6ediQIosBEtnd5r1FX1e7e2ii
YzyIS9d0r0Fxb3tlLnp9QmHJZjfEEHlewqfntSPYygolv/e7kXtBo97spobH+VNuAcJIEIt6Iqi+
xloUp36rF8/TyLDcDftSt7D4Cuebz518YKHWKdVX7dmCYWA8KKJiUUdqNxpjblmU5CWqnXWYG95K
9R5ttf6OYpOpBVjv+WtSziEvlfwiz6u358qxXswjEA19E51CDBnOzUgzeeBbL9ns4MeuyitHaaEy
i0Z1tTkw6GMicvnFL/1/4FYnm3zLctyy6PU09BDSzMOkLs/rlmbfzdJUb81sfPYJw6cHBggutk6v
M8Z/CxsE2x5PwxfX5EVXgnjT02X1dgWWy2LVLDXQsYznxG2eqdtqQAtXoCKnOtsPwnYrPf5ppMBw
h7SAT4p40TUhamvxGXdfNefXXRHDwkb1pd0Kcc5XbCdBBErmjHue6yE1NHg6QVB7fRTC3Dponwga
imR3ntPQWjOD15Yno4HaE+qccRIps2us53dZ5C9PtVol4Wt0ORg8uT2dYzP3IDQYlANgauwhppjy
/9ve+bXp6NK36z5SNk8BS69Cuk8eqjCq67eX6wxrFEexT/9thUXXx5ZvK3q22YVHR+23KxP5FiS4
3R+UaXtde9WWudzPWZ/L7qpuZ3CziT5AB2vjp0+ykkJtk39Aj26HTeEUZKG7JOKuUuiLMP6z3l0p
o7M2Cezj2pNahZYPzEyYyk79lTRMCXed+P0grfNX5rXTNxjGj9mSJNddXlTpzn5aFKnb+K4Kq8ru
+uJepvCh+kZnrkmOuz9HCbP78sg2fueNkoEKlpKDUF82TqNf/VDoT6v1D4saOJDx2oEHgXQEWzDy
tMO/51KaObhxnUlzMVROzA7xa27IFN5R8fPCdD+/gDtZyuQrAiOwW1vrdZgGn2xyPCW2rKdVwRj7
wU1MQpGYE9L/vo+coez3GMUSbOvOdHALpEUSHoo2SxAW05aWh3BJsuGJdE2Jyh0s6Qj+1uqMLaWa
4euqXDtLs8EzKctqZABUegraZJ4o/ZsptE5Lm7bCcQoKfw/QE1u/ARItCZ8fCiMmWMrAKjLKvEp2
MOSQmCt34IaJv7K9nLgc3aztXb5erNY+bezcFCjp8Iew4UTKvKEhrfEswzMWsJulru1eeP0Gmx8h
Y9moqjybsr+mht4YNCT3TE8oadBiIt3orWAI4FZ2jnU9C8LVuXpsuEELUYC1WytAggGWHzJB4ybE
3nkA36R1vxys4AAs5aXNlVW5C5BcLviNKz8UjugEcYyYNM55JpDrokzySzEt66uR9MB36N6z9bUn
lWHOfNubwGLaoMK8oU2zwnP2vwym26sQrBugjkfISmJpDNp1/hNWRaEF1OZ9QgjzwnKOMkNOSjnu
WSY86HM3zAMFGRvsPPlOQK7cpPzw4iOXldQ/23w1ikmrJ9DQn+Xhj4TxeFqnMOlWRpsjRWG01IGS
fD7FBK+hb72gYcXj3lue0aXgkLmc43m3Y/A2laJMi1I6xPAJcS4OrsUB/lgmqI9gK6k3F8iw/L8K
QVzy5ZZGLOYFVAw1tyWxBKgtBagWTpWuxNrbFB+nuIQ9Rk0DSGIJ3pPYsk6oU2mb4HMD6DwM+rRT
iKbaMk6Lfv0/Yg/tXwmEmgWvNv/Vo4pgWJS6tELMiDRlHSjU5Oe9y7AAGy21vDlBoqOvGwIJKkO5
316jUEaqY6y0/ukomFXWS7T/8PoDrK0JbnUX2lAYRG1IGgbM32s4KO5q1uMAcSVPxaRs+RUSSanO
Hevzj+G49c6vvFEVshPM0Z0jB+mjqkAWYSk6IPnFztXZQMDKt5Z10BH5lZ2rhp9rPBmuO6XC9BfT
CGjARQ20ZGKy4PoDsZw1l/+V70PrUcFge0vd3+z8ar2fuC7QyDT7kARHArlMWEgSHpyrr06aMn0y
2KdR5jAJG1pIWCStGCMgEuLjJBBSeP74q7nZ7CM30++3ARpP2mmWzY38HHGedCS/R+gd73WzWUbS
IQXJweRR1JIUxKTgdmxUhemdCkch6Pn4wiP89GXTIhoyz32pmbOkw1d9zDJXEtTzJgQZp7HzAbI2
srAV3QHbKRsW4sMd5ffVbVEngJnWzH87CCIDT1xQaPLb8+cn9mSdhXas9ptvqPj+ly+p9oKEs6Rl
IADjRYy0SHfpl/U0Uvwla7j+1vONj8BfYyx4/99U/+NVgm/jXf9bmYMJ5LEIQ+i5stQFi36j5dnB
QZLTX+cugNbdhW3QsSC5X7ht99cvuiuwOtDssag2k13bH19pBd6djJpQ9Rhafp2ZG+DDtKFpbwr8
c6UVsZvPG9lROZIy67JtPwT7rQqfL19oWmZIsEfVE2hxHTm6bQaJ3JwoTdgA+upiveQMjmcp2U5i
8thBTMtkeRjV37neAqnWeBJuAqpBf91r3r/UYM0l1pS1q1v7pJfFLTTMPt2Hx4aDbETkjNd2/EMb
glAFKer/P65DrFNWwXq7xI5BVnv5y7jV24z86au+r86ZU7JuXTvJ9R/oOzhrTw66po7IBAC221zY
/Z82zVxE655YBh1OA/0PzjxeHBhVj1i+VvlHt2iKjLvBCex+TDVum9MznnzERk2lvAoEt1caswzx
zo2lsljuOYDLoL5HvBLsOTqc0I0EiC3iI5R8KDljIDd2YyntVd5ovBso+3yHnWYxAk7oOL/wjy8V
TBtMz34IDITVbL/rAa5HJWjwNiHoaoiSGxE8rvbCGdTY1MX+5195K9gYWYoEeIEfaNE/xtSWQsQ6
fxPMdtrQuNuAL6Li+fEZKJP0yC/CSHBy1Gcsv7xiHricAF1RQUC+5KHWz7356utV64U48+/en7kG
+oqAspyvbJkgkuuNi1EJLF2SEKcKvB6ZA1l8nFQJgnddCKYjvk/1JFDg4uoGA5Jv2b+4iEn85dG2
qUlmj1To2q/rczXKmgt0kpdkVTpinCYtoy9sEYLOJdohnG46XdebW8+gt+jQu+P8/SMWQBUl8Quo
fw7tp4mOOfTmT+/5uZTpFXw/cjGpnp33u55X5BbdnOLFGAopM22gEkNrU4LYUkSbuMFM6bTJA8B6
608S1sSOwPHjwP42HiclMSEFzPyem5MAN3HcayO/jCQ+sl1pdAKjoCfVTCKwis+E8Mhh4jUR9Sv6
7t8MdJsS2Dgnot9auTuwcHDLRNb9l0QLJy2HHwQGhw3rsawEVV4IWyN/xZEz6sSfHmVDlKOoP6oS
iNW4UzaHVRJfUYdUx4KAMxIbJZba7wDc38nvDZxsrLa8T/JP+LkymbCCxbYACPTGZH2xRjG9FTJ5
8KVfdwCOlntNzURe0U6XihlTQzorMS+iZJ6Gu2OjGeLPugwyAXuByGQLG7+9TUVhQerQkUVESe/l
Z16RSjP3i3jmfm/zwECqw3X5StBMfq75Jr45aO7x2lZY6WGMJON86aBNMPX+sXXqa5qaTJoYJO/m
eaHGGFft6LoRtHeYs27JKZ6GTt/0BP3Y9zRLudvhqrABAJL2hhc8HQ4Y3YOrwEOpRa7doBvmZ82d
BfU9z+FT4f7CuWQlyIYTmoBK7sFeqM0fXwdOg7U5Ed2resXuJaOsGy4ZEOv0WfPRpCsVA/bNn7jb
GxNEE/OHxyBjAtJJIpz2i0Eztw1fpKnxQZdFT9Udg1xZAPkrmk5gpHtHso/+2tA86EhNIQXAJjh7
CGrkjoSo5Ij6i+EpAz8/BE5NB555+xkUELiiT47G2wfaJt4wwkgdBEAb/mTUupdlHCY/AGUwimal
4HigRovmjwWnKmb1Cc6wOPkEGgoUrXRAjS/nJB2/rn2u/4qQwRg1Qeivukf89Dck++sujflnInMW
wEazqYQ0hz6QOpEUF6tgt7rrwKJ9SrPjJuDAFCZvJmMGQmyo8j62lJwQJyOvwM87agwnfT/KzTW1
meAVyBUCqtc7u9lqSjuoP8XjvAMW3uHAgJ/LkOyf4rw+oGg3y2PT6PmMKKoCcwwwdHzciSdoVXiv
3xlfvbCT0Ws5ycisUvfkB3K+xkK2xaZ9F+JjO73Awz7+6StxEogaLG6dEKhrGazhrU1FvmbWjYUF
Y1KcRzKKoJUTaJqRP6RsDjoELZj1YYlQRAEwfWm3ECBygugxVP8pPYu8yKj2N2sCw62HcCRiQGlz
yXHVQvNsE2J2wTE9LoDZIej0GOsPMaTdT4jhGm8us/fV6Gyf7E2jR+IFJaBuwrjgfFBbMMj+ZuvL
mb3KbsmyPdVCKXu0qTq9jLZo9VJgqhKurO1veObyNA8OFz6qlPUo2lSH2dk5UeAIyafKk8kyoNpn
D0/qkh7lC/BfYWESJH/BNOMJnTswESIYeDmfcu+yv0mFZuGuP6LJF7jPycOW7taB8rOezEXQFxni
LH8PPOWlkTluvTEmoLWes0JhtQ+uRFxFVoF8y4yykUsbqPNWPQD2kNr+bCxdUyPMMR3dP9W3ksmD
R3h3ub5uLO95vzFEW2LmTlhuFZNKLxAdlMZPo8a+YeB9WZFrMvddG8WWIXoivr1JkW8B/GZewfa0
oQZ0AlN/TQUkuQSzeueweVW2s/S6V13iGN7H12ASTWayIRM/6bS32xuwI6oeS3reMPnqXWF6ebwW
5GZS0gdIXhMGJ2fVzqn7cPGUbf0mVFRVUEHbnLCEQhQFd3qEeRrSTrZK/r2v0nq4dGzxYlHCAifz
/De30aYgsUnWYpmC5ElOazuqWgAzc4Efih6FKLW27y4p5GPO7BFztFsOQV3RiLbNEhvNiEgpyoKd
i1TIN8brRxf1AhuF6YL45UBXID1c6vAk3rWL/u+tjVF72yHmwDtnOCpB6HWzrd6G3tapM7mk9yo1
3aiAGggjbrClsrgJMVo2d87TDHO83gTaFfLdKC/C9yg1IX3Jf53jwGCjJ5e4OZZ65ce67offgMLT
2JbFE0/eojYABOWC6aWtwLCaJ9GEio9MQAChPW4fYuHKndN2ANGwPnkH2M+iAY2BzS5RfwntrfH+
c+69L7AbKV+5aNfuWKuxCc0vU+yCz2zFuPsBavKKf7HB3qsxcuyn5N8S1SUphVSyVdek1ttAIEAE
q4YYs/LA1oXpe7nu9DOMVkgdoCQzhCk6KquDXkCyg5uZOg1tC7eS/FAi7ZO8W1n4nCb/+nybLEy2
qpsfIWBcr21v6FN8UUjvDdMOWJle4/4uH/iA2PUH4DDaLvhBrntk8w+5ZnLxKhdEv/fiygOSaox+
FgDv3CXMSPqP/eaYmb4sRAOYg56h6o4J/XN/HUcmUvaquJ/ahi8nKS5JZsNjCtSXn3SaeDbp7qsf
3R/MDtLZYWRRQPB7yS27sAy1j3GES4pHlbRIXA4LAHUKgCisvyyTXBPdB5DSTjOu3qK87IBjFtuZ
ZC/Xghq/kDIes66w+rInHxq/XNb2p/yp2hQK3c3kw9ELK3/hVDYJkcpHW09BAdaJ8Cd8aiUnxaxp
CKy/J8kkJY904BSLj05g2bfdU11Ckbvyd4xpXp+ETVvdAo0RK9QhyGAYKEQpPGfmTHjdIY2Ke89r
NwSUtWiT4ePw0c6q+1XjjFJYOw11o1sNTJnH9VVcezj4f4oGlmbIFlxNFl7/Gi2JQJCHZOY1ZjL1
x+KgR+po4Y8MDOvwbbMUuVHzgDyGiUyBZFljq2b2e/jqdG6XTz8lKg4mzqd5oSqInfjF8T06B/Jt
bcZK1yQg0VI08dR9SbE7j2ZXcLqoDxoTpLg4bjFX9zmMf6aPIhZtcTJ/aOpd4ouBQU0e0Kjn31Jx
W+6KOXHBM0VYd8F6sMnFQsJBs0G0F+Qo7Bhi9LQe4CkfOBWsZK6Zbphhf0AMllzYiO7sGumY/gJZ
kL4X+Y9ip9TGHBhZwszoUYGQ9pjXlyIfpOnnTRVshAC+8gFUc1aZs7VzNtCcMWZ/9BBlq8SX7blZ
zEYeZvID5tv8qtKtufcz6cQeZ8H8TVJ40wmIePVGZyc8PJMMMsScd2QCDvacK76jYreQaEwVMW5u
vo5aqKyhRuMoGPfpEpIoAszHDKXGK4i/8gd4/nmV/ByAWcFDryH360KLF2yUEVa9+W0MBs0XZ1E3
2W/9ZRPgSE8hm87L0J8BRQBaEUJvH0NCcCH5F2lww9wWvKkjbmv+Bka3QJVeTIOP+eHGah1BQP90
NhksD957Xz64cflmv31H/skHrA/CH4MH9FMARDHncTslK9cB+syYNQ9vvcweo37+IEkpAe9wE59/
JBG5jvq2QoNHWX5QljrVuLp6ZjgXwVtX16NGFl5kZYNb+VlHndQLe/1rmHr+sCRJXqdoCvrJz5KN
giwhE8vlp2OBg0IEOS1G8XzJHvFlSohPMMAGAX6+wtpGE/bCVS5khnuxVhMmQcT1tf9juKX5rvhi
PP+95D8+/Pac7wMJKgl2PBiCuP3469ndlcK3zLc0o05rHlzLiNPhrgp1/+q9+T9AB4mXnF8RHgje
+J8rWzdSNJwWlSh19WlDdovuLsMoHiPb9PA+5hXoXAlUckrckF8Kav2etKfLvxMFGohjhVJJ/PU6
abNrzewmNgTno5bTVUF/zrSMucTdVGvA3uARqJTNLc7kg/al12MdDCW/ikKGWmVvQbrZTbHLvmOl
1RQkRXHbs1lFqu/wPN2LWa7eahb1Nqpw6pt+cS5oBSqINWdinsf616nLsz/T9a8bVuZ5enrkzh3M
9PU+ouBQqEIed32Kc4Dd7DQ00p2LppHVCfAEdOmK+aLNAr05H1qZEdUG6NlMAI0kiDZ+Qit8Hlfx
t6XDVKUSEtgH/38UgNB7hSBNSWYMRdeUtmSArhtuGabC7yDIEJKbBcjbYMGJAtChTD409WWZP6z6
8uE2kYgOMwSaofqh455vYb7AQyax9td/VOcrFKEZmfSDA+io1bM9aFn1UkTzY6pK4pQONc3VRdJE
ro3yhS1+EC7+EPOX4Q0g9DXSnFWI16ePB8HOXpk9il4jk62PHWE2BKGrSsVKQTxQCFf/iFjeoMmZ
q192Nr3T10n0tXOTAbu4FvURTk9mohyfKM5XTfZq1rZhDDZ4FPoUH5b+99mEd5VJ5CktWIrajGh6
boWVFjQ508jMYvjis4KUvVTb2eY4vBzfm07ytyFKSScLzh1tbQ0+oru+vY+NOq/BCU9r6X/UgCpN
q2UQbUGMi99L9pdUG4RyU+cHqFhJtOTF/a18t1WdNcVk0w3icXHO9TPeKZpsdjhxTw9adam1D1H0
xu76VfAnlNLc3qFZPPeJ1HgpiVnLgmDXTagme0QhOwxG7RF6Y/s8U54xPvRJXVNd+fYravRNW0iw
rwcGeB5lUNLIULNGfWq46/MXFJoRDPK2M13UsX5F2au6lgZkVQ2qZhF+P42+krgTV7AsBCFjP5wk
ta0UT9ufxd8iFWx9Bk5CzYI51xf9UKG1XbpH9IDNp19UMe6OwdK+1IVWEx9aijAZ7uLuAYNsDYWW
2qkNeILluvAvv0/UqIx78fFLaRw+vvTPsWAdS/sg91cNipCe5Kxg0qXd+VJgN5Nvj4Of3jNZeILQ
erH3no/VlpXNF8559OSpeK/CpVy9md1q+sORJDOrvTOggVMxcABUnY7E5nIPhwKd+0aWChkrRHJD
inaKXuJKS0SJ2xIXl7CpxxI2t7zKNIwEetQ/KlWyUkWoVNkU7QhtJHsr4BZvELa+LHGoMhJtfn60
4VRGDVHLtSJ3uZGsxgCAmPJgAuik88YR3GXHWslQBNSRIxZD4qeraCnpAmg7Lj6d5Kmk3tIWiFny
/q4sjoQKn8hQuMc9waIfNYQdCZXE18xhVXlZLIP3w/ZnLldAscgxWpeeNfQrLRWm307gswp8INFu
gJ843FpSeDQAbh53MsqLKDpSyNu1lJoMfjBJwtxXuRmNOXvU5aoKAq/YxY6KOCs4nBVhpZiWDrx/
FUlQ7gFkYTLBuwbbfCGhvjtcE6IzAWrPumwQm6rryO/DqITCoJdt6ZQH92fXx17VASrs5Qhf5Pfa
NTxfqt8TzW+7771I+N2hLjZZW+MkTj4bCHWDOkG6j4qnf/oXg//ddZ5QjcaBax3UsZdYs26+I+ko
6Dbka2LzmQTPoHRlT63zsDWjrC74Q65R+w+Du9iXUiIlXf2yJVtWeK+vAHm/aesUWyV8CVKhLmZX
FwkuMEd6zkWcm7kD+XNnzUMkS70yLCeLwptrU1FYs33Ck9W4uuyIR6P523Qbrq3Fc2lW3yyvaHQ4
ua5Q+N/Da0OlXs/nIav6vT/aE2VxEGvvRENvo7pX9NRe7FeeYm168+WvQrjrPiTxTnriBQh8dD0d
xOUuIXIP4yu1W1t79cd54k8OUTS3+vLMB54aVb7H8Jf0ispd5BacxlNGC2d8UuEJiF9ldd3oQxiK
ZOibzMUg3ZSIMy+Ba+uf0mcFowLKIAJUjXm74fn6LxceOL3M6ZchPGq583zErLm3j0hoHQdDaRto
3uOYPZVIC0DPXPTbDaP4KiqBjK2breF+X+LANwx13NLIzajQ3p0LUpCBsq+MuqlVlrA1y8FCG/U9
SN9vJ3SNJf1SJZVzQ9I7seZtKSTRF8MVq5tYrW5NeEHPBLYvg+3L5ve/cOiU3zEFfnI7IulKIMjw
usUYNGda3lizwesN5q/TjSWafp6u1goZugld4hmjvljEFAmK+AA7k9NDOa/FYObWA1htILwwARQg
q0dWB38eRtRLtKmJ37xT0pUxeARfRGlEo5Isxo0P5AyFjjFK/6N5iYBE/Q1EC0iICrpvfM+L/5TT
2/GvqLfZv1u5dEAkGruPYvocDfKd8DAMCOxEqrpXdXDOzZTDqZXPEFuf6MlJScttdlGqlVoQcXb+
nP9R+Jof2fLynRubp59D4iyXxOWqryLUFtToKkeXDO1Rvk/zqHr/Qed+f044nnW7w0LJaQ/EqaSn
xalp/f4pIwPw7f6Az7Yy1y6gbuOjLglUmvKIKirM0sVHo2OoNx+rs5rX1w+GZb9/gl6mOne7i3gi
HXUWYftTqFGP6dea2tJ2GddKwn3GNumMQf34R96bWdr20lc/0gw5c6k+76hjtoSUo7Xp71msIPRd
5CmXVvKrtXGvh+PZblvvhC7NEan7zk2YuHh8NZ5Zd1kpvpKA9yDvOzvYKKZ4a/i9V0/qe0uenXKg
8w+KVcw40xFDajReYrgBO1EfnSsiQG81HvLeFGd3U01bHe1W/ERM1xFSPLQcnuZpITTj4SBdhxaw
wjwHCCGza5Cr0lQWHXaf7+IjtsyKXAL1Tlf8I8NjWH9toPgoyP1F/edIEBzjCJe9NW03V3SOD6Ns
1FpSwIBtiGj+CntVNYeqoXTiqffIPIBNLyFzbhJO/N22+QQLTOoV+mI4LBms5O61BQhjWN4+sjNs
8ShKQVvA7IBI8qtgN7zp82XNohwK6yRix5Iode1cucGxJz7GD3lduk8FhbupV0Cy1T4tNx2rb7FX
uZaJ7lZQxpJF4S4OTp1d5YDzfFSyVlA+OI+AXzX3CPW10ZgV6HSIIazWHZIc7P00556sRdI1Aqp+
CqFUcCnWZTxHf0MFFrtMM63O5RSKCxIcU0Yj3UGnEHzPpD2gJo4SwNZb/Kpzk7qugU6RtG6Oa6Ze
UlfKFrUqPALWAfTCRMlw0Lt2mzaRRn/DDsp9pVMwfjJDXlUlro7SeQTGPlB8vY3OH9+hS6Rn4jZV
Flohmt8FuGrYVOeCMjekmQX6tQewqvbfuJRbm7YzFR+s90WX5FjYGwGPRONaEPpLJk1YqVMNkEfG
Aa0jzN1Hjl4BiyxCW2SAmCdfkUiraLZ5jkxyFTDe6cjTdOyuykDQwvgkYCEQ0FZoyobgDtqvgwEu
9hhCOapbW/AhCVIclEpx/bObBCGIyK5KQeJqm+qCZADGmAPoYSIZmUsExqlaT/S/U2UhZZH29pEJ
K6NFAmAMfTC8K5B22ALtyY+mdcKJsxe0ngj4VpOpUM7uO9AoU2qx9WQ4KFzNge6t/2RVePU1xKVh
6HX+uzpLI8nd7CQejWN7ePruOtfvXmHMxtsHe+umEyWTKhqqTnWhEkkUJg4gyFM8ylW6q4Aa7o2M
UpUiElKVAmT7xMgCrMLKCfc6ZrvA+Qj52JPGBrop8+4/RRwlKea7sAadrlEI9dsGAaSWIjtP16r5
AyhEfMeXnwWU8tmbJf4WuTZWUb1YGIi/10vj1w8CtZZjeoI018O9TW9EjbxTsNz4tHRPHoz2ewpH
7Jl2dfxonejCKzVpApYgybhx/7PrT50HbAP+vtImTa54IAZWnEfNRaWM4fHHus3JDEuSas/p5nYN
Kp+iMuCrU7xM+1mpKAbTzfcYDTVnCebgCTMZJqv/Eo5OVWfJTkF1ZQiqK6lbS+zJIHhOwbWvEDtY
+LqiZlf+78ePDsSXBK4c7DdcBmpucO079lduumKlstmRicl+SM/0Yna3VvxZXyQkqq5ULliIqn+q
HUSl/1myJ9hempbkdCebvg2JFtnO0nGBdFh6gx9ghMHnwanWE7C0+Lf8dykGdWNQgRWPdZC/dSfo
4brwmeGH8R8hpgI7HRjGOrb5F8J1OAEYZg00jcp0J2Ll1cJ1TUsVfAgxEtSTSY08AoknDiRuVah/
Iylj4+gavlk4VmhqBKZw9DHJCjemC+MNeCeCgbFPPB4kVezyJJ7Zjoyyr7T+U9e1yJt1arh87L/Q
0bVi18lHXDhuKnPuSNHwJa7vXMlbuql8uyk0RQJtP2BFryaku4wSM91Zqt2yfichj5jsr4qc46/S
vkmk40H7LDojakz/2MNdfnWXp5zARZJDTfPtDJHk1oQU99S42GF1naTVBARU12bspzSAbzUxevVy
PMulxUQzcqWGrmg2AccUtGXgO3jgmZb/vWcvh8UWHbCGgvoi7eiSn100gYvNE6P4vrTIgCBtD3li
krOYazBMBz1LoWP3z24by1k0aj92XA3vpk+M5G43XwjLqHSrU22nfJwuLwS/HqbOqZp6wevcelLQ
Qy2eHGyoG033NIVIrEpNv/NepIDVWdfJHxgJR9hiGGt8M6OZdPAkdjoKeODTOcf6oDpc+smH+aNx
pgeIN1me+NQEqgosrzx8zaFeermopAsriFhhwitvp2lemXD3YCI3IKSmTGZMgJoTCb4xTkhkCyz8
UdwQYk3nlatpyW4Ay6is1O/Y1Mtm2PYGwbsaimb19CjUWc8vx3hoB/XNllYaAHLP1tasp8C4KsFc
s+kJ0/zLSsSMIVheU+9OO9wv8prOZOKeNmBRAR3RJRG65wHkRDCl2AFO7S/1+VY/wdLcwOPueZQr
Q8lZbSMSp7SqH8dM+dFQ0g/yMyBNQUDh/fcwDrctF8e7hhw30i+Q3lREyICioECEAK9WNndZJ5os
CGbvNzzW3i7L0wOcOtxllCLvlA9yw68zo/WHPMItIvAqdrDC4aJO9sJjW4yhk3vfnQQCLsISIlGB
wxOzCfQteLTeGxbgpajNcmwcUtFUiG4e6UAFSZE1XtGEfgnvpAYMZH8e7xPITCfWYDxyqDftkYrD
B6ob3CJR0KiNJ0Ec3IgAIZmnlgUWaqz3tzNaOcRCP8R3j0thxahsH9qENNJP+R1EYHVyD8MLrsbt
Gfan4ivMz9SOIl7PdZ8ukpehRj7we9oNYwc0CgLGVlwh00AbhokqFFNJEmOyk1hCwujmzCF3Tpxs
+nTtJ9jBvUtX7CxUQgXp096vqVtuRlsR/BrpnV01pwmGgyXTfgUMbWO21j/KAJrz1BG6sWayT61O
OugGjvJ3l2aj/msiMwX62HhzY1BTQngW1flgTLNo7pWs8X5gEXKOcaey7eH9b78tAr6hy7SJAibz
4ocEDKBSnXFWUe1Kvtnqb0/X4BZBNdgfDdX3XnA8VyLnzQWWXk1NcBoHWK+O1+kytERqWG+/6Cqp
BFmsSkaCtlRwq8IzZyTvMQ5m40PYOIGK75G8kyvf/g9OLXRQW/2E9j8tmSWoS6qDhJiD/lbmsTg4
RIlUlSCb6rgic0CU/xPQbPokTCCKpJ252PpiKh+7nptk/KxewDjfLXdUk7uwHObfr/efZY039Zrr
rget7o7D8pKZ5+GzB1qzrvJKyfTsjju0N80zNmUSGS1FDJBKjbSyJWjArhMTKWQHxosMmGXCI3nJ
ooDaNYNPSUBIOy8g/tAyojVG68MQs0zYUFLIgPeOLhlXiSDs5TUQ/8DA4qGgs7UdhhlQnKzxA65X
yjXZfFgla3znnuH+MhH+IoNFlpo3Ky48jlvD+hzUgLo3BaUdwuy2lM0o+T8vRlqAuXREaYpid5o5
GvEgVSeIzwN37wvAjuaVA4fQZ1rIipUw/dbrFnrmzAFBDTZs9tAozqAzxYePdNPXSRnwU8oabLJp
eJGAYkiOUFQpo8zDvsLzJFb4ZnPoDP6mfiM3L5rJ75hfrHEDLMaUMznjMNXQut0k5Lhmt4hH5di6
c9oPIDQ/efZt7dqFKLZwS0lu3mnZu9JMFYVE5veVXZeDlfeJmgwdeM1hOh1usLctncjF883g0OgY
YNDXYIboL1TkF8cmmG9HKSQoH/C897El3x/bqSpeZeBS9uq+2U+sFqCTYTngKjfbQ+6B8HPT1B9H
uBQi0Oaa/B26z8c4JswbV4G1TtRRaktY2xrZhc5zqR4AZCxFObOeAhlBaTWA3VO8VjqcEMahazz9
0ZkshHzWAaXqB8EB1L1DkRc2DtWSD4lPB3Utzc2Xat5qMCH00oT6OKIZ1d9qmg3eZlG1dslPUgGI
Skr08B/l1NRSE7htS+vyWwo5RZoaR2C/woEtrAyH2OrEkr4AyIi8hYokF98IkLTDbH4KLYOVDA8V
z0yEE1Ujx5yjdNKjJSc246wfoE16XCPVd/sE0PdL0DN5arQ8CfSpEHHTORppSFrN32hOjhg3R+mR
BJiTqMHyheKOrnLfIc70LOGS1vDhCz37VDFlOYsoSVPR3V+5ntozhayZeyMeJGQrbrcLpohVFtcJ
mCOpCSnnKO7vaaIl7tZguhNha72yk14rGZMGI8EUDYx622hEFEO6Mz4S4CkEVhEqx73B7oj3CoQb
6hMT92IoPILMWNT0YqDkCmxwg4oumHjwRTLCI1fp1XHpKbknf9oMC0iH6kIunl0tOLNnUXs4x6BU
QzvpolRiClbNaw3caS60GY1C12cjyG9UYr3XT7XpaE673n5G3AK/wlHcJkyk/YFZ5Y+YSuAtOMBa
b0BVFCGpGKxnazpqqHni2xclcJRJl9DxNKhJsy5OgJwxUXzn4fAJzM8AsFNGn/Qmwr1sSs9Z+jzv
vo7MXyBXQjfbs5RNokrOjvxzmVGklYfXcRrBtZmBWaSzZGzWYRbnIDphQXNKsRC6+YGr8j2jDi1O
9Stz2RMhx1ieM14qdbqYmwssWiFW1EJFljEG8Zw26wgIvVH0gCyzdshP1g4L1pI+/IStNXWaoysb
y54QOHjV7UH9B8/S727u3eJjN+DsPUVPpBSnbuFjU6Ofl64XVkEmERv+W9vFsl4D4xYy5IdtpQRG
qKnIH5EbqYuUzktcMSe6RWmvKC9b7Tb6ELvDshoCCebx7Bx6fCFLO6gBoQNShd6k7rmb86O6caCM
UFpSiZOVR5Nb/4r/SMJDtXIEWGLN/7/v/m3tGeNvMJ0u40rpz0Fo6h1/nvsSXTqnFVnt+2kOi+Kz
vIBKe6Fxaki2naH1LCQzh2tn9CJfxddMsFfEa0ThVTd1zaoVEnYlsRtdlZpUVJD0GypHERg1Jynq
Xcw12k090Km32KyVD7icmf8Px9ldPyB0hRyqAG+9FJzq2HwhIj5J9rXEMgf+wCmSm2YX5acEDMKB
jITNLamIXENBT4TctjwW94MoMj7L19EObYbq1YQDbpFwizr07sa/ePnf+waK0nRtKV0siLsWTG29
wM47X7Kx1ETQCPlcLnurR2mGOJPFWc9l7Chjst27EfnS8ZuaWmPWuNJrBIzgXtHD7kwas2Cl0Nrt
+ShuV2/v/KbEV+omJrbhyfJqx7qPtflmhNoLuFC8VFmnxHc/lZLbLhd+ZppaQNiWvkXFOEE9xf7i
kUsSLcNWWal8kqYRGCO5Iaadfs3Bi9GrsjvWzZWP653wB2gu4nHVZMqneqzHf040IQwlA6a53IEd
dbKgTF0z1+SpiqqpPJ7BfECP4ymmpP3vtJZpchmjYv9yGV1kR0A0ihT31BPjPphhnre1hWJ/lz9K
ER6IKlBl6Gc1musUfgg0QY/UOj6GQawPfS8IPkIMyXWOc7U9KgJZ9fYdCQtFp+aZEG3TjBdqgue3
BtKzrADMC2S7qn+JpwDSgA+etS626TnbbR6FqZfpEReNRHNjgOf8fvkPZGjqlrAnkmVRMHdlksBW
imXNxknozYXKI2KJhK2JZp2UEmUYVsNfvZW1hKVy2w6qHytAD4oVl9+wtdyCDuvZZPw1ziSub4ju
zq3Qf4GH3NZL3Voik6QFpC67BGLD4eCUfTQvj0UT6oDCSAQlH27wLguXi8mxCkoGsM8p0BY1Ggmf
x5zU4m8d3KGSneovjlZeyoWrx02OKhkBA8buFg5pTdXF9JyzV58rHSXl02NxmtYTZNZZWNQ2AFTH
vjUeMnJzDkDC9pAWapoRDpwG1+PN1ynblcicsmSbJLLQmNEgO4AvO4Hj+AxzUFC+KiBAMQI7SoSk
OJkDFIJVFybE0cEoO9cfR/5LsP44/GvWT8Xd9zo+BVMpuPY7tj9rpPRJ1+iRKXEaidBdKt5J7IqU
nZElOHGT6gYPELyvdLhJhQcUugb6GfzeYXyAfi4ZS5HEEFeeiDGX7gqBj34a5QldNSQsi4K54vRa
PGX+LnxZy/jrlVkLMBmtNCfzlJLA/kkxs5hqz/NHYbw0PU4wWEvSG0h+5kSQg9oyDbPZ+fr/Uk27
xU4ZkTPLX0wyk1bc9R5OMWeqI6KO8+LcV0PwHoPMGAuPUYuXoYaLp32uNNOSPcJz8jZnPnHqUL0b
e6U4R1aB4IbMZiwNNrvL7OV0wSCwtOasoUf+vv+Op8dAqnP+E76fHW1oUUQxqm3wV2wlBZjrFFvt
5DCuf+WEB2HIyQ/kxOka0SHcbW4VmjqEmxkzo0fqFScMaxdUPgquiX4CXzeIiII7ZQdakBdU7Uwa
cnehljOTJhuy2GbRiSNQd4cH3nioIfKL7bd+CKobhwCFEM1PF0ErNQimFvlTxn/+F6/HDIbMb8zw
4ed4c4n9enUazLFH33/29b86xf08Jlzf5HVbaVHofI4XTnaZSVOoRWZ8bP/5h3VtV/eHdzOmAFoF
ZdWG63krtEiUPyjujBhZKIye9eKVGzXMc8gt2reH+44VwydIs6pthaO0/QeBe7u8TDMYK0TgwIbJ
U1mb0ruaNKHbvqO5dslpbORdAW0DoNpDwoxwnxQpJ3lTvoxB+Us9FZPWvZP5n2enn8ykg8gnO3Mh
cyjGWdBkh4zN3GT0khEGEgzCe5v3PjdZ47rqnEdY5GxdOuyYkyJlxyrzbjLZ+wbcjoh6x/PR0TFw
2+wltvJzG9y0oGazxsZmbjc8hYZQDIXgDWPHSHl3c76l1UftB2l4LVujMnSifUp4CYsvE5dabvec
CiKT0u83piPBfZA5a4fD/9akbjVNnlfM00FIfqc/A2k6JSIwyUUA/YHvBefIHf8WmOG0aoW7AdP6
i0W6faGlHeANFHgNEJPdSMUJdSVRh5kRf9SWdasaGHCC9xL07Rh4urawVOr4FMgJIwSXjiilIfIA
RE1dNVsg7+8QnMosBR9WGWqkV26lfAhAMqtJ1naE5wPFM2TA3/I+EYQ//vVQ0+d6yKerJFpsoWbe
1wm9LcGjjV/qXqKZEtO97LdEBTBaKNyctWiSoOyLI37LexP1B+d+BJmmrlDbUlKyufbm4okRcAX8
jgW8GG2K9LlbdHROxCc0pG8bmFXulLtE09coscQ1ZdRthwg1+RGl6JVOhTIbrXOG+Y84sAbidss5
OodK9RmgwuCUip/iqnLWa3D65ndTn5m4qCUh2mD6WKTJihJ3gRzHs4Kk//0a2TuA0mgXulJ910zD
4JbDbNAaInadoLeMJzBo6/paONDz9p1ffA0y6sygkzFUfWVQ+MKs74gRqfZKIYd1xYHUXl1Q8O36
CELj3lEehlbnXRTuFQ+bwBhX1ZJ3O3Hgh7xgZi3lKZMGRPokLclNuCN1GIcYnbpUmF9rdhx87pxf
iAzfGIwFeK7mueC8s5af4yw5ybCV0LUGPVyQsAoUi52+HoK0gUK2dBDw3AWJ1XhJmef0e5CoxJlh
hVDi9ydtSkUoaKl9svEADTW3zmsRiOxgiltEXAO4LvfcAYwpHtjJDr00Y6804V9E/T05R3k56+t1
qUUQS5iDTuVKkWIb6Jru7jhcw6YtDnPpwttYda08Stv5bDGfrljE/p30GULBh+2FticjF/q/DbRU
f3724C16rmwc3QQKdXv9AkXAmGCS+LpMBW81UnTiQsKNLVKMkgGAq4UnwR9YYJqf7/5HYHaSwRaT
4uqhG7HrREv2omRDHpz6Kh0/baPcPc5pdUBf+tHf9BH3Eh2/ANB9DLoc1/lE4pljVBGlcpR6UJzK
TeCrOo69SLbs46sCUfDby63UNpX9kds+OHO2crX+5x9AwlRdPL+EtEksOr3+My+bdR43aOSsNHzb
LfNKLorP5DR+xZxe7Lwr9dixGX6Hv19N8CfNo4GRb5H8EOOOKcycdHjxRnZ+XjghyOJcP89eRIJ/
duEJx/DOeQM3tPnvgTfHfqtCh405yHixOSbZyHCkUIWYsSdJ+vUzyKczc+Yg8nM/9D8MCo3ujkAf
yZdrTwfulK1zQfK3b2QDmxcs27b8S3v+zSJNiaswWxp/a7UPdXqY7Th+4ZB0OmEQmAGN+SSlzrnW
f13SpctksURQuRwkqu6R8eumDFC47W83/OycGU2KgLYqM86LoAZaqoGtf8MNuOjneT3eV+kgQmIq
U83P6rZYHFqACwZoSej3fg4MJeq4R52eAxSRqkdO4O7RvtKT0JHA5CEde8SUSkKSU4OcpzmiaXPs
04v2+MhW30DKy0fVVYi/nr9lD1dmLMLNi6ayKYowzg2q9LHNyjyCUiEvf0YjD5xlil6FCqS1nkft
E/MYZhyjVMfNF/oOZMPzCcWjrIj6LaGpVI015zttIuV8VwVD4qNKnGvYJ1geRECeUsbADGVp1PqT
7JJok94g+UxjwWZq+9pKeKoiwtMH4hFdsV/x1xYl0r3JfKrQYoOEretOIxCDq1QhOGcu3SDcFhkB
Kh/rq/UhYDWwhv3DdZn6+iV8dFTrqNu0XmZOV3e+n1BKxbRflejEfxrEAVkOSapW8CVRrxp3p64l
scs47oDBhHEzZKwd2u8ZeR+MYSlG/2xK2qsULygbiFPUxq2YYeLcZ0XMui3KS/W6UosbwACVtAIl
g2TCQ6mvGTJDd/9zOo6FIDsNzBtCjmNTNsJbqjGZxlctt5xGNEWdqXrb2jGrCUuQlwC/jY/gAVum
jfbBT3PVRuE+Cai+Tj7/hFP+QQ6V4ylUgc+ya+5pVoLID59+Ls2KRh/zUfDbGbv090TMEMhu6sGU
T66sYCZxjq+tZ16GnCO8fKVnzylUyxACCUDiVsa/iLQsRh9qzqonJanVK0Az4D160frJNBVgiTkA
OQdGA18nxE7vtFltKiez9ryt1Qr5aeUAD7juPiP/6HfYgFQoIrMm71EC8SlcE5GfS1nhqvKN/cMM
p8AgaZNT0uSb88oG0q+cjxsLIEnJ352perkqb893JczHKi8Fk1l+Zgoq8f7h9v+73q90yABFE98o
GFASr2b9T+Zq6qLLwmNMe+RHhSKtN4N8pHdZMoAV14HXkz6qGf/mTNVmZM42Urb+bUoFspga7vSA
EKK3yOBP1p//EEdD2dsHaNyrn/5vNowzHZuUOtOhkEI0aDfnNE1SNBug+xtrMWNzwiGZ4hTul+Pb
r5oF0W4cyboI3E8VlOdLV9Qpd2mEvtgm6msbYbUgYz2EdNXF8Eh3wSg68bU5JIzu0oJvva1MA95D
lGNNWEpca/pCvOZh4ildnwaDCB+zpjdFFZBTVCULTcVPmRb89ZxrwZFJ4pJ44HyD0z369XZUZMQ6
VGf0sQ96zUYQR+qrcPiE+1Ulm91Si5W2n7AzkD7yYEyMYVBtGdmhwAyPlfxKmA4iZz1qv6U9NIbb
Q0F20uKWzqsDvCZukj7a+RNpU/HBd4cqUR+zhBDtcwXONwPMQ3CgRJiTE+0eHdwDhxE15F5BomN0
6xoKlDRksj81Mk8MhF657ANDiSkiKp8F7dPZbBW4i2lkOWOs1lDbHL05wRXXuDmLQJX6xt1aWv08
b4es4rwqD7JW1ruNGHs73TPUaCLp7WLCiDfCdUk4UHOpEgnZqs1ZX2gl8lY8MBPpcH8MCYu8n3fn
AtaiJ80B51xIwaO2qcIzK0GkMq4J2Km2pH0HWtY/3lEl7WttJRupTmKNdvFFwwlM6wQwA/gQCqAF
eCazuQLcvPuUnJqOY5+m08m1ciiQ/ywgZfVZDiEKVshiM50KQ5CZSHcL8mMaJfZ/aDqL7ViGPmfB
XcHHYdKQwGd6fTbxjRRINYOv62Qzyt2fO/3EEN2WHtFBKyvOhpITPnYj2b367D1G5gXO+LnKql9G
zt1puopHnaIZLXW15n+Cl7CCodR0M/WRWAnzWXB7Cln/PA4ta7OAoYOjnGTFpcm3mlxdxc2AXBNQ
yYCF+y23B38VLF04lAMalNL0DKn8IDnBDuRtiM5vt5jHWIPwOfMcb+ZHgMJ3+87pF+qKNrHqcvpm
q1lK2FBDmg/IiT2WNsiwjqBaCLHppxEH/8CvcEDFZVULK0NxhSFJT5AJEEklUTn8bT2B7X5sKn2G
PI8ZMnJalmVN4XYI0zMAveRfFQ5r5GXe4UfQnByBvQnTnLVUIZ/oAFEUbNOqQ1HqNxtInUqmaxGx
qKAHI3FiW0xEDTFJz32FQvnoH/Qfc1CXjfqF6YFkmJxPdiNmJBXTsXLZAnUDmEPqebt8AhGkBZNY
FuJwk31fFrPWs7V0/LETQR6iFkzdpkBJ0nDRNXjHcLrc5BT0Waf0l8/2samAxEc7b2jX/3J/Coil
2kpV4CxbS7R976QBO7NPM7RlrunGyAw3FgiY/aTmJxG1/3JbRET8sp3y/EAWZo43lbp16VP1QUv7
1dIm3C9uTJ8txECuedKmIPYF+XWv+VwzQ/4BytBuQ6B4WjdXaX+srjJ1E0K3RAOq3LPcN6oOr+bL
LtKmpovY84ADnDRD/TgehG5Z4FuOO3mQnuplT7BaE+Ox4wI2ym5aGJsW38xoiLpz0aMDbaiN5PdQ
qHfRYIbvCHE+Qdbr8HV6YlIIQDaKBRVRLTNRmBhcGZzEF2plwdeoPT0/m+I4X60rXddoXUr18H0b
vyWGGbnIvRzWoY4YqjFjltje62a3JcFw4ke7JkuAs8+HYn9KvDcKIqcMnwj0XOdp726V6soDN1r3
uuGEEvMCgeVyjWqPKcB8+i6QThmV5fXsMf2UDsA4RMhlIsCfq1UIhRUryghV67wnoB7Mo2WYgt+8
NdpTGpkcmGxhk5Ye9ct5Jeb+Kt7xHsIzY8WOS4YKp2zVU/1kFgM/Pn4Ii2tw9imVW2mtW/VF7BT5
nQjignOHrZV2S/tck28Ac+uBMmGI77UnppEFuA7lWrDGJc6VZxZhoNX3WtT/KOnFbDm06VcXwqvD
JoX0GJsj/zwcViWT6G99p7jLkinbF1mR0C2vpEpXjR4Lg/KCnDL1gO/UB4lqHuZf6110u/wZhKQR
j5XW+DHEU8GsLkLLbeVk5vFjetrIrUCW7Ge7ynovoAE+a0dn+JT4D6vXtDCnTol8g63SMjqKnmg+
CIsn4OKPLcrA7DyUB41jxmoaqQFVmjZnpdm3RwDjF0tR2alljD89/qpbUA1yld9zKmnSsqsHcXud
mS3+iwtfaVdpQriRVKkY6fOE+uSis+VGq4So1SmNs+TTN0IIXk0XjbVmSeGPx4eGaMYG57nJ6Zuj
MMaFVL/V3SNWqyqL4dfZ/a3IKPhgLnHvb4zpQSBrEdMPfVIoC733kVWzAjhAWVFn6AjQYixSPm26
QqAPeGKgNEeCYHONp2TvLJ+o4xCDYZxcuayVyvhShZKkayonJ8PPaBeBam1vJP6JaK+Or2Ah3bC2
GZrxhGBgKqbxfZ/9Oq91RxIYc5lKJNOZ1V9CzxZsDzh2yHaeMNp+M8Da7L+PfSt+Mn4oP9/42aQG
hPRp2IY1ltqBhWaxhNPU51o79rJcIq8U1VUhzx61OqemYrckAymtVS2ydyOrp8Q1VgPSJlvmIY/b
aGmNkMfTyPzYqoycHArzw2VwYnHl0f8y2RmDMIpgsGJAPqy7OXinkLSAqkUCWSPCDHr+I8gm1R8J
KUYr+zfmARjNPm9/41LyBVqjtrepaFXeIZQcx7lE8Qn9+Rg/nUL2JM6AJb08GifM4uGxewAcbKfU
3Os7iQdimrm4MATmaGzLmpZM3VcT32ynlB6UVszwuJmxmdUqnM2MCFSO8/m8UbiHiVxozTpEp0R0
+t2kS43SevQEYTKQvcYWtgAhVb6w9nnu/NomrfPlDRiNcYEZFYOpGCvJRiR0wSIyDrDmPgxnW/w7
w3t6mBHghdfedivkgh/epy6cIxNjpNB2JhzazOhkVmv1gTvqBw42jDmS1AK0x7DQoMyDkN3Xg6jy
ElOyJDtmo4Wf53kwKEHwh7oua3A1Hk2sFEs3hEmdMM+5hK/+7BDLZkCZqHOG529FVQbp/I+r93hR
cbxC8j82Dqjye8mc8Y6G2XijLWCuv0glrrDGKvY27rLtoaVbMxJ8NWyeqprxD18Nn1j/h1zrKLYY
3Xx5vI/OKfBEiFehFJiO9alrYsDnKCyBPUY16+aIg/wJN0lbBDFDz9nHDxPWJkhoGNHSRsHZvJ7f
GbdTFiIOpdwK2MvtpKddOk38QvV0VAqa8Eyqeb+tFP/w3rpbcc9zRCzCeoX6ygwyp7URhTPzfe5x
oC2ZLJAyhDWaQDP5z7yDm33IDXvU7r50RfyxYM3BRSrirhTK+FXFUSbj8T3/F8MkwDrkcwVTkqA5
5HhTDcz3xevAlJkHK9pgQ9u5ogb0TqgRKklYHKwgmUCpzmZi9s5RAnz0+IKJZkPqGuGx+NSbeJKr
U1HKwvC9OYx+1sRE09Os8TrisHsoK3SLu5Kd5GkphQMecVkq9lbibr3IKIIHrvnsYPrfd5LII2UD
iIRNhEYSbeOfHl7rfBc8mkZNt1NedMmzFkg7lJpS1ZSSyTPitdN/clJgRdHzo1md4WDUZNHqJhCX
YQlFc8tNVGGze+MBKXj5gp2oCCYqus72uMvlrydw3OeaXM0cTfejDaq6uEB3vGkAYW9GyYMLgJpd
IeqK+vV2SwNIrtgbcN88dR6wk1n3BLnxUgGEqEFGFNIcq6m8SrItnIzytsanNVD87xNpczaHCNi2
iSWtD+XdyBOOWzsD2pRivVV0f5tA0VBOQdEfnkn2PFH7ISeLTKhbwKJ3EM64fr1VPekDmy1JebTs
xnLEtPXzv7DnBx1bSrZgTWY4gua1CbTtkNuWEBuombpw+9M9MvmFLHsOEsMLoZG351ixQOQUku42
N/TTlf6OoVlv0iYPby+adclDQ28q/GNmYOPrbzrLNiSUO66tIh/S2ucoxa9MWbAldxiKiJBOOhgc
TQNN7v8ktpTvC28J++UrOsEua4aU92JXoJVDLtveb8FuI+7b8oomjoEfpb00h7SRenXlyWTOXpGN
P8fRaAQpO1lpbcLIhL97kSN+B62kXjeSmhLBL4KR2NXrMQHOE0ZHNxjP0suUkVLqf+k4E8GScV10
P7DjreRMSZ4sO466+iOn62tFJ+XYCsLwM0IJLIyH/fTn0Vl4RKsx4/LqTzqtSPjpC/la86jNt26Y
7B8iSV0dOSBk0qNavU4j02kGq7JJ/FJxDBMuzDF9djInPMfXB6iV0rv9HMeDSznX5f/sfKUIIdbm
3UcYJe7ugy8MDCSZ2TR2q9BmcGFUfT3Gt/u6BlF7A8Jxmeh2A0Dy0QLvJByy1q2Ot+xJlL8e/Vdq
H5TGN8cXKE1p8xiTuC2Ic1YIsgw0II+yVtVWBWUeOBhwP+o5w82/ZDOWf5wKh519dnRBG8Qf9beQ
kLE0ZD3rcG5bS/1G/UZzAsh74mdw1yClUg3WNGYVu2en1dxO2mjH7BqU+ymJbzBjsHr8XYakVYew
lfD2SGU6h8BTDdQ8g7bCZwL+Lywpl0+2eRhD5lydyj6lJIMCua9GySbzk1EdYZqWYPIUNBQ8PoeZ
/AX+hzfBnyI2FeAiZ+HklzvmfL6Y9wLgKaHs1YtS+OxY96KhBfzmE/Hu6LUUL17NJxR3RimFY5w6
pDAARhRziT+eJuo+sMv4lmkhcd6vCZWCAImBce4k+afEVe0U73vxL2gSQXdljO7wzofepSvlA8Vq
wjCFmLPvkmVnB03g1e+wG4Gn4SpmIoJ9eg1Zo8xvhjGOCLMatM3MmFm14LlUbPxTdClLszz50pOs
FwvwndVkv4TkLmym9K2vsxhJvMnBmZyvhqkOr3HOcQf6HzMcS5AH6L36Ia5SI4+gFLSNKyzFdJQD
RHudXw0rbJ3vrrdESkIQ0pRqpX6xUnRLxCUm7iU2lAJHWYCjmyQ7KqV01c93UPlLD0w6xY1gxiWW
B0KLZ3/jXKmtPaHlIcN7uprirvlfMZO3yq5VGPqesgUqL07oRFqlIB0GMIvRjL6RgyjoAh27M1WY
tnkTajBbA8FUYzAPTv8MT7snwmh28gaB8Hoil8o9t0LN4xI3E8TI2A4W818k+hWNMlJ3EhYgke3W
ATX7/osAvvz551nTWmBDgwI2QdJsYPPR3oJPToie6e+ral00TbUiA/5nK1om36i1Uy3uX1ZBafN6
fyBxXx4/YVjldMoUqpaMMG99HPLCFGkbxXWveYtxeqwby08ftSrcVEKE6BE8pThfh5ucnKOHMec0
nCcjUY7VHvp5SUgtgcwsrLvlcncqnT/G5uh7nY8RZz85GgU/7t+sBclhRYQ8FWSTLba8wo2RGvOR
I1Vt4VyB9zmhc1bQtVuK9Xrn2H33V2AH8/hci6qJkIePPmvSSyA23ShzX26DGy17ci2beFHJhIYT
P/k3JgL4XHUby5bzvmRn/ax5LQWCW/0hnwszYeUPaclgP5u2ZlBLQLh61IE/tcCwFGH6wVUa9gNp
VtCZ1AuqJOv7koQ10dxv9lArC3G1axfXfItM2MoqhsuOMwjtuxhMkw0H8eqRS1gblLBEWsa16CYs
KwhabcHzYkPoZR+N8mhbUfm85ekeU2tsRcNu+XM1JdoV9IiqJr92GZcYPlyjJ9xKkiIaD3nDWmRJ
FHrLzbORX+yFEbOQGRM5XbDXZP3VokRS9aNYvJiNW7yxUQxWHNmGDgaMNSYJlj8MMo7xEvhwMJ2s
m54lZKPDqgdF/WIe8Na4xw6RT8u9X8SCvwizv4A8KnURywYugESAJxyE6RQK1rfJGxNUL+Bnq3ML
JOtlIbj6Iz4HMi4M7L7Q1yP/DCL4+VYWD57qrdH/gX4tyloZ+XFfHsQxY/InaJD9KkGCFbrmLP0B
CAA+NGbAnmLGF6LaLGWg35bbKJwssKYAYGXnNEEtWRdi1EFvGlpPM89Or5qf+uOv3mK0JwZaPCn1
zxzTneiCLzJn8Kh3ydBPOyGCaPuJDpS4sapEsTDFu7yxmgBgeY3TkhC8bRQl0xFIFFmZkNSS8lCt
iKfZuV/K6zmkVqQmlDtEEe/9/KGzdZ/7oo0Q7TFHEHCB3+/uctv5bEtdBOpkluJlAV0hNODwnCUr
O/JCFouSb8BYq8wIdDPBBXHmCNmCZeDe2QBAzSocdPxX13oQ4Eqc0LgyeFsN/KMMlbuGsmQzt/4f
THKEmHN+XEetBkJzdNNGGjgHvQqK37wgU75gQCHzTxQcFWd+RD23rWyyJwClL9x9vIqUpeq1OlFB
hxwY4SkqLOzKTqZMY8cWXECOvNOh2bcyhcSrhFdWQWn6VTMenpL0t4edumJBI5hvS6Zksp8U5Gnp
tkciJTEDKVEqrvRUX7n9BY6H+3zDW3zua3bVuc1ThcwSU6KcX4YTwE1dwPioHCXKnh+9jzzZ6/gz
IfuuQXWEYJwKGbW/tMJQmiiHCumtuP+HG7wxU89+aSYCkIJFFHRmQ80VrSinsa0B1xc9+/RxnnXw
PqaYby/dmt6LDkAP4+E7wdeWqJD2NkJA/PZRhnkQ/d5D+rRM+O1NWZmv0k4xYXcdTuQOgHhxlRIx
1yrgcFHC7QlVFZoxsXkOPPQxpro4tO6Seh14MwTko4CyQ+h0JkCNy4zPRP6TF2yPHDjnWBxW53xA
lFGQlUlRY8fOtsKe6KosFjJf+2W84uJ1CRyMexmp9MgRNK7cZd+MDyqkeZxxo007DePKu6VORHFL
RxENsAlHxBmwYLeNlBdwxhrKIwLvZywldYqUoRX06WQH00Cw93gWnnqvbxg0Qr/YL2f6pHQaIuj7
6EHi+7o7JdVWrS0RDnNbnPJig+hYInXFFyR+Az2SZy1okeY1SX85GPydzgEkPyLXIyeGdpWMsWuz
8Djptg9JVtksFZgYF5HSXm8wPtRGOWx6TxpOew4ex+fhbYX1eVMm/+gBxjrE+f+3IFp2N1tiiCrR
hh+eoNnm39Lq4rzkfbXNzt8t0NwhmLENfgtaQpimQFdpZKP6ZWjyYPoLvXojTF07vdqYxJPFPRHY
ZWejTjKIuGf+RAEIf4Xa0P6jG+5R9SskvVEs8Ml88pjQAB0mdYbzfeEi1l8nRu/KWtqLmR82wBjX
K2hDBtUvsCfVZzqV8jjpnn9suN/onlUz9jz4WXEcu5xFUTc592eh85RgbJr9AUDKwZOKvdz5jynA
ZZxv7OeVl95CxptfwhMmTHCtFeRDa5bE6d8ddQMhFi0TbVb5Kg555SXcHTL7JioUiBGLFX9oYsgO
OfBF0n98qX0RIHFoRH/6dggGeHoD0ioeIPB1TZVEH+w/fHYSkJ1KUZpcX1v0BCIcax94zqekWEXr
f85yd+ttXbCysv3rUW629rAlxkYf0LIaRiBE/dvEDLi+d5+DKYqgbyItZQFTZeKhB6E+oyjnWzDJ
jKKAO5W3Cue0yTAfC1nGf5tKVb61c72PGkN9W5hrX3eWMFGSCTEKSHeSuzze/ZTc72UNGPrzNQ5N
/zbRnHMR9eimK3irJ+yDPnmpdzOmCZPb1v9dDU5awD5WHxfket7sUZei+kjru0w3p1kxXQkd5jNc
dU5OH3KulpMjwf2W3bHYTQFjsaP73hzM7+W/ivfVUWmA5ojfNKJ9iBhTQbZhN2sAUt6SD8F0jLJY
iVAP0ndmWnY4kpCRuVb/aCwhw/e9nlb+HuuH2fpvdi7cANQSe53Rd9lmS/x4nEdGet6r6Ahw4rWC
nmORl6lPVwomcezv/J6TKbBXj4HdVBORPmrX2Oa5d3FzIDn65P6JAT/lNvCbsaog0/XFZJIwc6KC
eNummyako3qS8xTpP/RLHptDzdH6Zso0o2CTEOicgwuIpSvTuyQWZu48gtmEAJHc4lL0jg5r1NVq
SZGaAv9r8RDMLLAPTLwcxsvx+uEQ85rcSoi0Dl7kC7f6DkCWs8Ra+cOoMU+vT6IpDYO6wKMob+bA
bEzxNaz0VHkOBisarqTFtQwP0BDZ412rBFYFnsD4HjyAJ+SUNKWOv2Rjur5btQmD9cVzPzMbUchn
dl/rgndF1gWGiYolQZH2KOwz7y+MIh8+D9qo1EkHwtiQ3KmjTUUngZ1mo5qnBjtAmQhgipjTHaas
UrJPne6AmhiOcM+99H3zbFPf4gouT3A3m7CaRXyVNJuHn51mKxovepn781hnTAJWFINPoGWx/1a0
gcfx9B1cMvxm4HA34Ja4OJk0PJ/a0pIkd2AuK1y4Xch5z8drwXL4fXkrmVWqZnSJ2ybe9mthCNn4
s1B0SSRtT3XoRRjMig3AzLMWs5hGMUJOyGSqGDZALuZBohB4x4GMHL/AUyp8AWvRyomhkYvkhIiz
HdLq9jQ3ENw8fvSBbWUMGLfXVMCgd/sHoGEuPceKMDLCJnfgW/UDXOapzWi+fEbLvI3gC2GX945N
UUAw7NCrCv3uZsiI3gqAl38w8QM35sSdxVxv20FvlZiDDNA+F5d3TesKgsgt2I8jwEvOIk2uyHl8
MsnEUbB/vZuF00Pazq//z+ah5SAT10TemRpje3dZ5kQbVNC0ys0TLCFJlYhaCMOrxSX5SMO+dm4t
DxXO7SQTe2Dn8i2YSss3qGhBt0jTK8ObprJs6DAZkRaeHU4LETT8D0gtdwUpucgBWHS0J8ncIH/9
fQChpphR9h6NC4/48S8ajE+KdEfthqbmhQm4P3JBybGublNIirWFpQ2TdboQ40LARJzdq9OCUbrL
y+SxXM/H3Sg32k7miLvJ4nrlcOcvQ6dw9siL8PyjLgytP2fiMxeRHaTBO5n12I3IgK/NfyUESwwM
yu4QedW9+TqvCJfMChzAmAJkawgsF3Abvh1VaDTUe1d+PzE8rUq7QiGlbHo42CPgjWI2BygyzsZ2
KrHsFxIiX5DaSaZz1isxNskWtRUpc+hhnECyW5rGQlf5f2J+5PGeYgR7qoSDcHQScRhKMMxCwCuy
3SERDHmjFuPM7ABMKcGW1msYs7vETYv9Bta4+YvZB+y/ugauE2msoy7fyigZ6qfby59GTNjsR9OY
M+HrJiTKbXMz0q4DuOmXGyU0Zl4pyxzwh9MB4dx0F8gk7PXbIInM7E7MznM5YAMTEWDZip3iO9L2
ulRSsfobVuS1rugvyHRRjdhLouJH9SwYdWsl09f9Wk5ODi9+dtJ+gZ/v9cD9EBMfB/yJMJ8/4kth
tyUii3t4dKL26gZUZTriPIQI6t7wJBekWQtd6THoWuSryj0C0YCR1leWKsxXo35n33o1FyYeVx5P
6QnSos57PoBkwlj9QS9oQ+ql3aQB+gyjdM1lK6rseJm2L/8PGwxVm/AkNzJHkWzWU4rYxYflhF1Y
nocmcuZd6wTMeSm/ce6g1DpCyfl2/4Li3AFgoJHaDe66yYnH/kY0HLHlA2hlopX5hTPH4N11N08I
rsSCkgnLi1AMl/cvl0YAsrWfp1kUbVT3F5Fba3J6u4FBguIDSIPBuHcg8hGqU+OCoBrLsW0iqwLG
pXQ4obMyYm4WpJ1xUcTnSb62MvFn4dSka3DMzegLX8YbFzfhYxXE9h/pneoGte5twG2p8xF4Fl9c
GoANa1oBuRXEEvfyVg19xgSpG95Z4d9oXYYXgb49wUtlNRKFbTRp0IiE0c1XgeYuGj0d6Ys8azH1
8z882PDmMbmt2FgJbPDIm1wfHLlFcVxFLdTxUAYClJzVohmnOvm+SBfFtMSmHWrDBQPILkQIXBMs
Q/FY5zCUcmOiSuV1FsNiL5z+3JI8Fy40Sj0NPhgw40GO/hcFVEuX/Otl1p9nLhBmDUPHYNfe/icu
l56/hHPV6Z9Auyxcc7L6uREwp2GpakFA7s/Ly04sFjn/hl0ZgWIx+VjY+VMzMnwhbmslVphezK7h
VspdfpwU2xJN5XLslo7F38XvOMPZ4F7S+gNre/5Qg7bHsmburxsiRBSqQExcZxdLg4fCyGa7Y3hK
xQPy6p2tZGgifFaTkkC9UgrhIc6ATefaJ4vNMc8wLYDIMxanJjedLi+DxOLg1EP7ElnH3FAJYwGs
kryBhzlJ/zsaxHPCWMY0WD8XV1Gv+toUMhqjbGy6c8fMfKCrCT3E/fVqLCyp3TV6tMkVdXxSe8UC
A7/5B6kPs9Oviq85NQI3/JTMkPIu6kL+4fihoKEoSQqYtarOwJ1/QcnlWHUfKmlQe5J84xuo9bW0
Q413eDotjtH16BKUzPEofCVwLp3+ZsRfXhgH3D1vge1yM6joqZY5lOvkFW/rRXKnAIvcaGwksyHs
CwT9KgTLJi4BALPi0EntrdIqz9pUBXbcUvxvjzFmyDi/jJNf4AEFcxTX/atw3bH5Fq0omD30J4Vn
oGTTNGUKD4l4SA4zYsMk3oYrIvKEDAKVQU+eljMQdxh8pwFJpai89Ik8BOl0PJZJTHPCa3z8q8E9
nMdilJgiivAHRFaAAzGouZn5TAeQ/MsrhRFuRdtRTEOGZyxnboAZ3d6OMqsbZW979cNYNUxvH4lR
j7R6LRarnfyLyQo+/f93KiFi8zmHfQqGMXWNezuUNu7CAsesxuZoOxT0VM97dn91iZ8vD8vR9hNa
k76LB2QPqEC3zo3N6A49Fc2y4WEwDf7TKA5rfQfF5r6xdwe4NZoEMjDvXoUgVHgFjCa0DP2UkVuk
fGAVQCRRZT5R1aeFZLl+Th4scGc5tdoO+WV5lm66zSOekERYy3cglq5lmM/Cji2PqWW3T+/tIh2h
ocIWm153bFFhzpAraPkmGFHDFRwxA3NYpRtZLzUmkHpiOjjkZ59A8PbkL/2uJLjCkJPkRvUrquKM
WqD4Vw0QnW8gC0B8tUdpVN+1x7Ujou+Ch7Kef4KKHXp3nnX1/w+g1RyEA2X3VwmSSVaX5dg7bEYr
fuUraLZ0eRqjjazeFkXAMV0vbBoO0pyf8ilqJJpcjekAFNS5aVSgO1xUQPcZmiPwv9XUR2tUyq9e
U3wXBtrpSys/uYsgQ7nGfP5/uBJNyVsy9hJ/FTzkQd+fEAJJDPUBxgOmZ3H9/pNndQdZXcG7owfJ
d8F22aJygCwkfNE7ZI+VR/HnhWfb/WMZU19WJXLZvlCaoThVbVh+SeDoMFWOzCifBoEYelYhAd6I
iTn2VM6fd4OuxXLIPngQHOM2oMQJ3CYfjJUCUfn2Zr67mioe0A314lPulBL3aM7lPvubQSUKY3Q2
06y3VJtLEBSQ3t7IZ4FvUKaDOYfKa1sNwq8oxyvZ538bxC2SnjgzcioUfz0M9ZacKYv+s1RDtcR6
/Yxbp9AI4BQXrzDtj4djwa2t1e4f5eW1aR+nvsNBqfeToQLNuCly0T/Psc4kUK39TzaCk6N+V4Hr
yLDdsJmO7nPtuStsv9sSwgS6z1MoVBAFov2ZQvg5CpFKwNEEf9V3abcRIOvwcqu2KijaQQYW08sC
3p/JSbAuCkVw1Z57lV7u2nWr7a4bLFixHb2ZWSPjKOKcncwhzEXEhsITX+m/8koPeARf/SC2D/Go
UGndmq8c/hTJWXDF5Q0861ioiLM/M2Fl4MLtHXuOSij/7avYM/HY0xOjmq8+UHzid+XNpiY1t6E0
dwq8k4ZqruwBeBXqs/4Llj3XJLWR6dYJiRuGKNgW4DchTPQRBTHTqBmaDwj5lGKdzKHpjTF+FrKO
RAJgKWUKuRQqk3a1/t+j6TxpGyW/2c9sxGD/mVA4N/gJlDB/vAR9I4O5kKvaYzwTkX++aK0M1eMB
7d00Km2DG5j01WFTXu6sslLWRwOmtizxcBC2bQJ/pKCXyVvzz0kWufColFdZ7rRF0ECmpYf6qUeA
bMI+TT42LHKTSaPo97di2/UnYnkwfIEjoaFuyEV3lq75hHWgi9w4swv59SJBXi5I9wR+oV0beFkJ
Va6wyTSlCgrWJCMVzpic4gSJdAVdZV/b2DWDySzm7ZR/U91d1IUxXoDGuy0/LPV0aM+gQQlDk//Z
GLs8WT5a0ckaB68c6KvnWask8FBrqpwNAP+rT8Vkc6EDmy5m75exu4589ID+zcWSUIDeNJgT/TER
0+xN3gIA8jHGk/nVJa/zDD6j9stt/YnoIjeTaPKLztWff/iAUfFpp7qxnpVH6hb0NDFe9ag+fGDU
IaktD1Xz0DDbB7UhCJUPcVBIafihC2kO7AaJN/oJRobKZg4L07FUQwoGNm4L0Y4uecYAy+ZExeGw
ZdF8PrOeg7qiKyMkqYFF+B6g8GgkCGJcdAZ4HHd84QxehJYRMbNtM9EQRdlHJDzsHfr7NPcCNUwf
hPAeHDOs/NyhsL/5cM76Toj/OHnnW5TcaQT40Lvv2DfdCfB4uj3MyuuGikzP8LPh6wg96y+8K6hf
JlCnRY4bo6bXU6jx9iCHaxsYiof8YX/NSx7JdOEaOke0CUqsiKrSrSeX4iwopmh7Gu+ukVtqbvny
LjGhT/OWRQ5sp6ZieWy9h6ARrfx1+z+2COhJ4D3TqFdlgdTgDY4ZftVsvv0na+Ns0p8PByvLfOvL
tObQX+LqXMJDOY8rswfyEPNThz7/I3TxdxKzaf1SFs7deVHtSOktlIYY8R4M1Ki2Fueb/G3xaLTz
YXPOQ3qqXJFmPFn9FjGIeYhtg+csoBT9npGkp8Lp5UauZnUUrjDSXUG+rckItgQehM4i32BmPR9v
/UST1n2iYuDVNi6wl9D4K9QxtXCgZR/6WNh6DGrS+VboGYT6MKyEQw3KnV7ZIhRKyE1Bvss6qN/4
SCeFXmafddslENbShW+za+YOEbxiqNswe0BnVFhAiqEXjyBe7hchSn/X5Jkf/zFGK0SMnBTpAJe/
xIMVIdz5+qsBXlpn27DPps2fAlp10F1qZcAWTEB5Lcuw6OTrl3YlJLBp+l3mRR/Q2bGoz/MVRwda
VaBLyUYv7pY2R2mi19VtGZZf5TRIsadYcmFNV9jtTeDmbWukoNEMQyQYayrhEHFN99qFqhWD4mBi
m3a2mipojJIzs5t85CCtGMrQC3HUaMbjHm88ITLSe31VkeFm13/siuEzrso/7eZkAtyNiyhyFpRZ
dlZLZrUU1E3IEb6uF6SnpTLGT88OsuXnJcav/3i9nKiU2+hQYEZ9/sG5ZUnkgyEPBTvvpCo2YvO6
HUr78AEFmeTt+vygMTqlrhB1cMW8yPA2BK0/q0jEEwD9eoo3jZx9dWd+3LX4PtYdM1V+1ZMBcxiV
znXoMYd9E/ysZ81NiWAMa9J9qfL+B1t4enLgrq3E0VmX8qP26TRs27E3zodKca9BvOwp98wHt2mH
V1+P9EpBf4l9uuOTw0cCq+aXQVLGWb3kCrCvXBK0usmaOOubAI3DQxYCbSxv8Fox5LElO+R6X63c
QzwKC7wy6Yqi9XosfQbYb7nUY21iR+p3G3UbB3W3ODLQF9LP0IIHwC59lol8O8vhjsNI5t4dY8LG
//AunGHHx1+ohjOPx98042LaUpH2BbuAzS5F6fIj8ybbehkKKxEhYOyuy55XYqlGylnO90PrlID/
A6YKg20aoDDYG7tg3pRB6coFPsAOhCFZug7UXCG8c1JTrkEduXl5CZTnqCmUlbNSc96845v31m94
oAatg11+7RoY+VZ8aXCwHNy4AzY9hqDw7SfQPZ10/tiyY0lNjwAu2TuTOZx8QcAEYLyLrVB7R4pi
f1/feJSayPZKXQ7xSjK6etuxeHkp1gQUzebDGjjpdqwDRweR9IkXBChrAuSBrsUjPV36QBlzHHWk
4/xXcRfj+560zyvIYrVPZgMKR+G+V5X2PddGvu2Ffuve0iZcS7a2rwvxDyX5+vUW9l4/v5iC0ZAH
NXTF0KDiRrG14TtdtpG6OB5Z+ao9dN/khJZc5aywG03xeIqC0pyu6efr3sl0XlmO3lDm3NGDtlwn
ycLiTZTCYQQ0UifRk/XUjT1LMdoyPaVrU6AEP29vdre0vsMqvoofkwtnJ6jPZRv3U2XGblMC8AD8
IDhYQhBUqZjx/ycr4ttn9S3vRF42cfqq1RklYeR2/A//0X6KH3TG8z1dvSKbi6PxPSbN+EHzwXYC
jtpBSaIprD62fy3XB4KoFQZ4bxvn1URD6CeLZHg9oYRQLFnq4WoGtkaN/ltEcYz8BobYY2f0zp6I
kBMGEOEPnHxcfWeh2pE6Vy7ufhLvu2SOLPzgnMEQQvAK9QXhBlsWo/Pxq3uny9cO0kDxUtMLJkQI
gi9Q8S2o2asjc+SoepbGgHjsYsds6EDT+FJ2SwJPAF1pF39Bg75VloPE2oy+fy4RXWyl4q/P68ZS
Z8CIfY4erONIbOERBbZDiUxYGuLiT9UpsRx4jhs328qF1poNBhmkgjyOJ9+c2oGGz4fGbS3WJ5Xh
pkEpo0qb9wKC+NoYOY6KGYiGPiSXcAE+QR1h8cAPqq2wl8PiUMg2ubMm5MUTFHtfC+Dgx6NZ4nPF
yxTMwHPiEybGgbY7B7Ycbm5hGrPN7saeuXbITEPh2h4qfSBtFZT6B4WgnNz1OCHQYwFbvi8gcGLF
HwjO8iMRlhWafyMetedCkJfs3SCp4I7MsOvogyoV60lV40Bfj5y0rjmhsBwMnaRMFRxdR8pjWdKG
OVOhq3upRfbMZhk2Pi/n/Eyrraco62D/eCWyGRQqGhNhOsvkseJv1z9X/obyx+v8OjEXSQ3CQnH3
7iqTBWv468WcQFVR1B0KcUUF0FhpP33OBaJbgDpxI2OqNsdVcyAb2bAh0WLtwCys02t9PQFB9Jej
fAq1w4ByvX8bKPRvDe8I69qdxLwF7Dnau3t4DpfWpBHjdgE3a/RJQSkfoOb9Vkx4bE1SP8Vg7bq6
s/U0Hut2IkaNfz+HwkM2R/p+ToOWdX8hgTI2PdFL4HwKRg0DC/VrBnnF0KmFOj+Pk6Td7RJrfeyF
MavvXL3wrhjApf/jgxX1abJYmkrUYLXyb3Qrk/5CL27MJslkzRxBle5zhTVXjtGTBBSLMRepySmV
CkQWdwNN7UTKX9cj+ALjpmV/lUVGzZfCX92lw9oV1GQMC9X0jRES7e05Job9Z6UCfBgUP0htbhhm
bjKV2Q62Dp6QdZG0CBqzUi6CMKQbvMQzkuQ+ULLDJdWFgm1C37sHSnt3BVAUvEmjSLM1Qb6eltnK
pIh2q47qe/2Px9//icZZ7A8M6g3+m/05u/IjscT4hQJnIHO5nO3GMQHWtbsQE4f5QgBZSIdacsnZ
RCzb77CHW7a9yYBv/DSiCDSMIsmbYezQTQUNkdgw2EVOZYkX1XHx9HH5Hy6G9qmxCP75Uf1YDMmy
95pcU4AQ2JYk4egPkd+IsSvUmMrl3NikYDnOyn0vAKvYyp36Zm5pIz5LwkFcKYKO1wZP1tsKa/wD
/S82ZnBdP/PeH9xPB+1hn2L+WuHEK6V+/FyCEADLWMW5hcGmJcgZjqoZvqA9KsM6aphPujrZlT9B
RvLQ1Z5WbwzIF8wH0owRyWHUcArH8pha/LW0TVd7ymZEzU2/cMLnWY8RpuLJn/MLvlLdvu3tJ77N
Vr3r1P8Bkf4oxfX1VN0VaxWLNeo6U0/jXKG6qJAunpnDj3vrIoClhbr/mNcd1EiErmv+NhO5SnvS
uENIBl272VhdZgZd92YM2rGlipDlOPWomDIjZ8nakdb+zgXqpmCuyqyNjVFizzbyaojcb1HcVcca
5A7EljEZLI6E9tLPkF+pcb5RBDaM/P7INGqp+xleQEmBb5/Rt313WlEVSV7dmX1mp0SSLkWLN8R+
l7kKJj5FhuS5FVJTZBrf//JCRNXVs36ZERUeKtDCdJlef787qgDqFIzJRFJmJ86lV+FCWUwg6K1t
RtlgLjumXypyPl7TYFgl3OX7DCEoe6sLiAb+fqEpidELumcXBoArm/NzaKePafVnrwTBmswBtEEW
mIBs/j6UgO6QOSX69ruPrb0h7Z6A5z6/frpQ/zaykUe+OlD5ukj8mNHKbGlGyBpUdlTGtCVTumLN
0BuNudE9QqEl9ng6M2ZW6oYYP8elcwrcH33t89eYUN74d/XmlNc1CgTSszOManAEY1cTWg/lqX+8
hjBhII5dwhNyLO91oeyghFuD5qyVNjHIihdpwAKw3IHTtDojzBnppSqTNVus+57OldRrCDVvcDRw
oMMJu+BJ7ZKHWVefNx0P7l6VKASbsgYB0tpMo14+dHrLM75SFTKSfaeMxOzs6PoSOpkE9YqJ4ZH5
gR0ky+z+WNfspmFc/D5Lt+V/BFf8ksd4fgRO6bRWa6z1AfawYO/hCQ07T2C9zxQGKTROYQvGa3wI
BPfe7N98H4ztXhPSmURxohLwuHaIZDOpYWHuhFvDWcQq4rcJc95NtJ6Gma1x5rCoe3i+LliussiB
Lzd8v6+qV7+AFmL4XX/LNKxCl96LfJCIQOr0PEvynnYxNiUOfXsTCY8zPyK5yOPkKCGQgOmqiBXq
fUOj4ibH4j58ercj16IiHhGPBIWTHsHeW6Ic4XerdqTkV3sVYENuJ5MdyE/CjB9mmvYTLGKqcRAt
y/MrRxAOJFSAjGRcbtpIE5wBM0bGbocNp4GqpjCBJIRZW1r+TkXCZ83vq6iNL374Tp0zKqToikLN
JXi778b8Ia7N8RP7FA2i2DyvIL/jKUjLNzJp0usQj3W5NFItkj09L6Swvrlw/Cyju/It5du9CNfP
MUeCcHKybjb1TmYm+CHvl6x2uazm7ZeeK4v8BLi/Vch89acvHHiE0XMv6mkWAyUBptheVp4jLw70
UYa3e/3X2d3scUPZe7Q4eBcEtMHcOJXElpymo6Hvnnb2RgTDxuqWbsGHiMsdPSismFeQqEIQZJ9T
WmTs6EQ6V7zkFIldnCDz5Q4nPW+aZjMB5FBxiUWqXszUMu5ewTXuMl1VL2aVUjEQkGNFTOXQPxBu
ojiN6m5xKBqqkohKZW4HabDj6RfjR+/oZT8sMgLgdTsOH+6Z/iZbyca3FZh663c8FDSOYK5ExJJ7
wTo2O4gaqN5kdOncFfDljdB9EiihIa13+85dCUa19nvsXwxUN4nmCNn7ETV9Qxa1gCLjDfp1Jlbg
Qz1HcBYeOY3a6oqfvO6tt2ofkgBOn63X24a80Vezaw45YhTpke8coaKsfJ0tuMcdMWN+BNuh3vTm
AczmKwN+1rYxQL7Tn1XFqnKWxxLELxOpKGrLGGMlwki8rSJ7SycDbzMte4rgAFypEA1hD+IZ45+V
XLGBdiCZjlIHG5I6tdabivK0dhn1uYBZIytEKmG1Olos3Xa0sdKCGA4h7indE83o/Erj6iQYtEJA
Q3dcTXD3H+Eg/9IqRAqzChCHQ1n44FRc0E8mPC19F6CXmKEDyDsV1BvUD5tJhRW21djXQvbnf17P
qT1ohUngHOTW3oSpS/IsarCG+2EWttOdpf0Doq0gambcnEkJUY8XEXsVTI1Hiwn4Cxx899gbVyCo
HY4mGftcnIdCEA879ReFQmiOJbgD2HAETf7tE2gzN489X9XgiFLuZAkTu9NXmiwd6W255UWDHXys
AmwJviiaAqQ5DmV5O/wtilQd4q9TDsMiW5IFTdCTDy5TxoPW53GEfLqDHZSRpdrlcN6iegabW3y2
/FhzAykSpiZUNMNZVOdG1ELwOMsq8TAwe3W/QzpuIcp30lUzVlLrkJee0axAt6deER8cY//mKhqx
Mpm6k+XbsJO6Ri8unklyFAajJKP7LbW+UMYTXpkotC8XgKIS92tqDKmumBQFxB9e6d/Auz4Eox6Z
HhpnFCe61wCIY/Q7wkNoURcBbwvlfanIilEMvKxC19ZoswBbuZA9Y/mdpeQFn4hF+Z/2tdoG14dT
OYz9VeqDDiAnL68Z2jQrh+T6VQvg5JoxVR8eg1fe3okfpgOLXYCaOmi4RJkrAetmwGny6TFdE3Hz
J1N9TdJQiiu7exuCNtsCa+vBlXMsD1sMHxbg0s6sEdeREMmMO5XqTzaN2+lxAMMgHG0N8gVrUSSC
ZqhBcjj8wKfvHj2oO4ZruNcEmglCiswZU9jU5ls4ab6iz8nqNTkwDFSv00S7Rx2peS57xjihzTB2
BEFZywqTR5SnHzC7RD/86/P7U05iKkbNbV24FpAykoA1lTaOvH1rDJvnI2Uvm6HnPz9NSCFpuNwn
MJhHz/VItsy0Ex9IF0LFJTpr3RHH+zZyJSMBw/wHsAc4vozuzezaOoQEN0Z0dwOM9Ief8DzAM94q
yxGY4DKcyldQN24ujBo8UhcQk4fePQrLayUJ50mwrnRrD1rk8vH/ZNUWSt/dYZ67cMZiritessHS
Oj/nRp2F38IrrfJM9bEuvxEWRBOdxnVnRol2zQLFA6AmrDdnKC844++I3nG/zvDNrrpvyOVNrsaf
3ggatff3rBcpMFQqOVDtMRj2FhF/mF2oM4gAT3gI54bev1RlswHaFQAo0EkXwH6zl3wOt2DC6V9i
agt1T9U1k5un6pOt2Boy3pk18rT8KCfrqQV/uwbV9VcSE5FinRWwT6KjPr126gmj7Z+lqPGvk7B3
6yURoiQvyzBWxQhL6ewAYIQLuFMfRb7Llnco5LIfX3rZvJPVwmDU7fZDkNaIwLgtPRm+xY3c+82Y
wokogxi4jhWb7YmS/ev9xfuEOWp+FJh8iycFpTS1uNVFxdUTZW3vwi4nhMa4YdlYQQW4/R07bL5m
qy2ueOBylm+tnfF5UR5ODRftTl4cEZxHA2Eab0l8496Oj6w7pt4PjNa5lP9hsQ3ykEfUAXx2XTmh
HPpoxJ2NIyghIGQhPGTBc1YCud1HfC7jxDoPz6bcbTw78SpwLWPu1x+Moj8g6vgJwQXnuyMQfMvj
Zun6ng9nj3PhWM0uvlPJ+DBWwrbz9RGMc+Yc0eEzGGnpkjPgg8RC27CSYY45cBGa+bp2eBr+f8vy
ueUMw0w5B0GDb4zKHfbdSvrsp94CkIQZmSCDrFCyOej/KrZl6bYswKLvm2CYaoN0O44R2qN4hcOM
B+/z9ujhsMF7oo7Fkd7GSQ6YmxnTrorDbXwt47q3GNPa1tDod3UvA2ld6VaUPB6nfJ71Snpeziku
VzlrGxu77kczFUm3PSV+haOaWSBBkjt0Xqi8QpghXc3dW3ymqN5W6I4tBLWbOPCrJX5JdOJzXngt
6Q2ROqzHf8wpAik1QwJDiI9wfsXGV2229FImxhODZDB7xlPV4ocb+ea2kfTgOy5evzM7NXSdW9Wy
+M6bxbx0WdF1FsCvQc6GUBZyLuRRq34QGoRyq615sIn5VRReZYH1ptBihOSg14bLFedqU9lWYbKx
UYn2AKPQRJ9+jXG4vW8m1atO2VtAeuVd/KIFHqmBeQVyrsIyXQzSNNL58lh7furHMFfEubL3Krvy
i3Q1Ox4bUPOVhqmyUEtqjGRz8MvCFo3jL5hUx6zodDvqVPa1QuKV5Ph2eZOvYlLVZ4z5gQStkrlq
rDTiG7rID1tsCI375UPIu9fCmpS8pq2ECU0NTB8pcKClZanJr7K6urHGXyXqSx9BekS0eVz0RHDL
z1G+l72EjEBynTET22PeDF24JDLYvkjRzpGy52ZDOH9sgFxaUY/frPxYQ0YQcjd0IMS8TCl1DhRf
/GXSa6jkwS/E8IGTuj5vdD/jQ0wWyL7e/QNurjLrWfp8ZwkegVi4R4IChBGZj/tPfmZZgHf3phWE
SAQx9H0EQ2mLnEWGJh7yBW+N4rbzrgDgr3AiKHyyZMyp8WVrdUM62AcE4wPyqF3dC4bGnrKDhmvd
yK1spx2KVS/GZJ/CljCys+/sIZ9A9DBv4LUsvuTfP0N1AS47dgUEOg5A7ZyjE5+O5ciD0j3UmCob
XA1zW8SCRkGHYe+sMLaUTUSizqoCk7WnGUadSR4h2f5lVa1BUZTv1IuJAxpmgkUmV66GFdCPO9Ze
Xp+hqFWHt6ERBbUFzTHDaM5I8W1ih0SrLjZpB+C9IqpXwDErjtpfNPIEtKB/lIkHr5qm6s7Ddv4B
SVabpUFZuMWda+9hqqKQQ0nhp7sXVstm0QzBmF+DRtTRbWbzO/jTq5Xv098xqxdod4ViBggmvQvS
EsNEfHcQBouMCJmOXByubOn5G12FRHw7zD61ZcgMOV02XtsynQLUwe92MiH+Ts67oz4wHA3ox9ja
Yj9QgChjC0PN7JBk+SaCO2yIiyYf9qlu3AMw5Z2aKH0oP5F8LVd0MIDA9X6hQKXaSOITuwrqG6n3
AGMc7K6TlTCUAW0V89/USiYDLac8eQCEvl/i1xHC+IpT06f4yvaIis/P0omSgRcPYKIBQxmYB8Fh
FkX0lSigT0HgsBIKBci10EoSPv/5aTlpcnzQqDL6S59ZZ377/3tOOA3ELw1sE5N+Z09AAG3zQwm1
oSpHbyzFUKnHWncyj+UafPJY97oMyl+GkPlIW/pxqvJuB0EG5irNiIgUOYmoF3eSvQ2wW7FvPMmo
Lv/facsH+yrjUlvm70y3DxAiwAI0v9j7jak/8OBpQre9eXWqVBSy+i+khdwjuZNYpWGrqO1j+1o3
CqAR5Dl4NqIKfuiWDThPcCBHvcpWBi0W6bcxZRC7S9Bptq4sF4LRYZcAAtidAdBmELgkJtxwGjp8
iSX+WMt8JpXs531GizMSKEyjkgf6M5dWZAfcJtt07rNoblJp45HVSSpfY9k8KQ5RXbqgOUbyrv+p
++qp+YQRcSka9bN5/u3/xEIMLeuJRfKw/TpodkVvMvgATnsx0PJUjxMMwmT9F8jbCKFccCvLq3K9
Q5s6AAKCegCEQVcZKPCS7uOsPV4d+/0dQa5UB1nZi/GzqaxpudgI1AerlBZmlxbD1EjUu/WXBX48
q6VokiNkfjuPpzpqTqe/SdNZA5vwRQHjhpTfBMaOrKqyyP1i57hzWlayBxb7gDXJe3JnQjv0mvXy
gpEi7rmwO8WV6rbSy9opcXg8UbflO1T9j36Xr4VXh0MN5F0KAh+41kPE/Fw41RxdD39BjhHbu1Cd
XqHEEDUUktDgVLrHRP7lbPicERD3AqiMeUZabp1pTj5mJBgwNtXwm0Re1GraCqOLHgexczqgYqtF
4GW3vW6Dg8hnU5/UO2ADyWfrU5yGGdNVy2gAfz9IAop/pJ+Z3kgUg0+h6Nk9Q1PCSMhgnYI8Sl9Z
T7xD+k5eBl5slMEYkLtbk2yT9mBaIX82itt8ZkQr4aiPFzikamCO6FmK1EDrD7zpgY6ZJdgontHE
fA322Is+sGxbQx2upaStwXkkKu2z4zsQIhJWKpA3ewayswyQozg6W1rP4dJRCIbMQQOzXvhI9l1a
w3o3Lle5GPivJG6ymlvHUZjsOgL345wRi718XXRDkCM0qXlvGN2Hecpa73O3/DxH294MZ4gcMiaT
FUopb6FK49yNBiZMOXH7EFAfprJBYu6T5MIzxlHLq0SlFJRzMn4JZhUNxIBI/HwwyB2Tikl8nwGP
IdnsQQNQtLeASpgiMLgfZ386z0I51lvSzNAy/s7dgtMOFDVV+ro9I8bhJZTZqrZOo9R10NafNzXH
41b/NGIR5R/UX/khPh4hWocxe5g2GAw9DwTUjg+oc6pDKh8o7ukQ3WKxV+JUZ9WtC7v9vsbGZNzt
NZeRBqJYyQSUMvfIc1pKpZTHSUxNZnbyqInVXl9WfPxkxDaCPMshRsYDM30aLox0NLny9oAmDMSy
/863mY9ajhKKCURzkbOeSvKAsj5+QH84949cjfXJ+t/zxqeZ+armKfKvbeFQtbz0wPWU3sGKu3FL
qoGHAttwFLGbahBbChhLbRHkdAhPyYOf3nFr5rLMMKQq3oi5ocwvXnf5DAYOmwzgL8uHAUqMsi46
AFsLZ08Jx1I3jfgTwfUF66D8z1Nrti8lCX87W7i1IjSt6u6FLw0aAJNoNOUrX5PMKbgG8UaOfE4d
2wywHv7qmNIPsjlpNjjNVUNrSBrc5Cv7Of14Or1BC3DtfzmaP/uP9Hi7DEDdgF3rB+R1DBQR9pGA
VuJuNv0jaDtNboWAKA2+heJabi+FJxAahBv4ftZeGtNXanlZFTiaV/+F/QT8PSA21g0m7vdKGaMk
uomnI8OjNIQ94M2Owo6/TH4Iw37/NEfWeH7tNg1OebzARwQhByIcDMneVxgZaU8dvnQSC6OxdmlQ
aEzRjYokTCsClY4DwH2+Shyciddc28PsobrA0AM5oAIYKrGcCy1Ma1d97K8Ekj5dC6sdQI+LSsyg
1C0GFYkKcDcsznTg1BzNtKFGaJMdWZSVezXxWdSbBksP8on6+xjtnYusx09y1Wwi9hGnRaKgBT2x
XwRfO103GU2GLKOGbw69TBVtb/X+KxKHiN3gwDxSUZuu3qJyvne0QiIevC3jLi8in8n8i1F5ptvR
wNH3hQS7IFShXubJ94/3g9IXMPbUUJTjtUOOwAu7t+Q6jjCK70G0q56o3z0eDviDmchIClCb5IJX
dekbiXLkZQ7gOwflpgzqtwn9saJmHD77ZHvJzJfxbtI1FKlGw2X7vOD/jUdbDgcaBQXqVrOET0oF
Uuv6bwlhY5OpqeJJb7hJBxuL/StEQRc+4SM20iuc1YlIdDfp91h9x1dPMr7fisHeaqBoxYx7z+NG
3xe9EaWkWa1ZSrpmRzvqA7eN+HKQlv36HMKTG+OMIGF0t2MM9IBlj+NmmtjXsp/aIRsxhHvbEUXD
pqM7GA21PMgm228JLTFyadkRdOfOTw3+x/NnkDNRoRQWgqF2FO4/4ZBM9SK6bk/9Xep5oGH8l/VR
ULMOJOs75TSW2x89n+rvLWMMDL/WJzPLMs07kEdslOJWWT0ccYcUVIu7dsMCa19ZsQKnM+7B+PTV
e4Z3Wb5s9YmeuVkB5l4/DBGJVSq5Yx/W6v8k/+QG6jwFi1gdkx5BSsnlVLSdRi9HYSDlrx4J2KMk
PXYlbC8VxpIz2kqhak2rItxSMFbSrDQX2164yFz0PSvc7Qt3e2YmWWbepewfn6xS+0BNPl6+r3zU
2zTf6qAlQQOUJ0AE9NAMJhX8y1BMesiUZ1tV+/PmgK8EOgKtpoTw3R6aHa45D5N0RrlT1fk0Blol
rYMIvz80zpMYCZEHQBnF6m2wvWLVCs+Im9O1BfKcYyzcDDyApktHTJD0Gsi3OhzB14F5kP7f72Kk
5t9uHMEmTXTQYqcxjmzhrOMRrlrHnseIpgR2XqcZ8yxTnHQUsWI6vh9Li1zYCHHF7n8YcPtjzWmS
+tb1mAqfvS5jCqZJvVAQrTVRqCTendRXjHDfJystQtI3uYKurrAMZhnwH5OCZh04ekVTDyfkoyQ5
ko5IvhINzXObivuk8+sidhTNHx4SXqPw1CUeCSD+6UZKDYG0Y6l238x8oyKnAsGCdY8sOxDA9/OY
++DVMlpsslYEArhbBRAIqurKzB6e8rZZsGNjkHrLQ7Z5AgmOyd7dkKB5Wh/eR4PbT/kHZELv3A40
uYuXddyVNIOWyJDL1LW1kEQYD71lokwGYSv5+EZzdSDG6nFt3VajuStcBZUywJ5PoAmtfOfq+sxU
s6ccxl3Zxl2ELLIlWlZLAp6R3fe9RgdSogAy9Y1OIYmq63XghzbANxGjn8sfK0bPqvQHtTWPqrfN
QQY9EGuVYC7SbYt97cYzCzPmqkh67BrQ7NfqA5C3GiuEUEbUhQJtjlGpFePKSqa2aMxFWYQl5o3F
l+I6X52F3Qj90/SPoqPbXg/o+q/M1sQ/RgRtyFDMUasJowa4vRE8R2REAZxLu6PM/dRIH0Vfywmy
BlFFxAVcFqh+HVmVLkzLTMBMtS/duJs9nyPTXzWCssSqjB1lEd1abNkG304LT3Bz5ZOa2u182QNF
tpzop5AcDgatNoxoxa8NkPKJNyqsqrtFhLfSWmpHKUO8n4fX92H7Z6ueC96OxgY+23O1bj/9jGkH
FtrLSEqZBmzZlwT3wG4//dhg9LYPGqlXq9CHp/P6rde/u8fzxmjSu6RTmqerZ+QhjPDO/RZiMIUD
bWfbeWMwgbd5AKoVflRCgQdHE3q6QDaS+1HiGBXDIBGdjy8UPNADNByGVlpmyux1cHVqCT0LG4TO
whFoD+dP+zPIqaKTdiqEAvUMsbEoS+NZqRT3eQc05ivj0F78AyjbOWwgKqegvSkx1JuTE+ivhbuv
Fc1/w2VwtQ/Q9Cb1+kJda3dm3fVzBip9SHnDn9xmV+waydqILPUEDxz/B2AxLgjyMGZ+BF+jufA0
6QO8Ogn3mOTLWpc/2WpBq9l34kCKuBf61a7T0WDA6sPR8ATU+3nW1/lJpsOXhF5kwsmcwQJ6LkCl
V5Mpr97F0hyv0x2Vq0b3XZEHUFfv0Xuo9y5lRJfsIUvm8GxJ8kzRCXxttF7tZhA/R/p+vxQF9zqv
nS+0QKnxl6BdO01X2yLq5gTCdMmp9qVe4EDJsQT54NNwfnjzMpF+EbdEVsWOzr3a1CpqCy5Ccv+8
JyF9DDCloP6HD1c7JcbTcZV9r2GWqL/ypI+WZes88i9DFlHO5K8AIZgw70BOyk2nAOuQ99xrauoy
+7Dc57wIcjrSSyKM5QQAR77KiZDq+JwnVL42GcIsW+9/pJgNNoMOMkPfP42RSXWIAUAFO2Zg3MaA
Dzwji9c44QcL+B6ce3vOwB3KAyTqd4+VWDDZrSDauJGpOFHzUpIi+4Dt908Vt5H4pAiDEWg0aj+Q
PIDOFQWHSmUDMhwcrkM9HX9XdIXz7JFYl1HcEP4AkIiGcIPbksWohUrS8lJ0PE10uMAuXmu5+g9K
4v8Hqhei75NBgSy3EgKyklU0vcMaPMViYzpdASa9bsnPSrhBLaD5blVI2UTn14XIpEI/UTHff0iX
a9HqfdcCitozVQYsuvhSlidv3V62w6wvtkmfM0snurV7bdceV7IRT20q45hnxGGVi1SACiHXHyWS
79AxBoBjbDVPGNyHCRTTSCt3iGcEDEXBq4WcaNvFePpTkqETo2bkS/kGeI2rRRih3Gzt7MWLYNU+
M8WDKuqwBpYKLfuvi6G37bkHxga80dBWcqj11crGq7i0CjyeH0HsnOG7rs0/jpczS6c8BNUkWB9f
RRDEmUBKeCmfzfXxzqzbULRdRg3m3QLhwRBAQXPpN3fhlWELiRyVnvOAr1Y4LwX9JlOdTSPt9D1U
567QLi3J9sexDpBa+WLpMmnm7B7s//4sQMDXM44D5RBDqYeIXMiDsjoVZvhnKyNNZfSXyw6kwbhJ
6Zz5Yo/wrj8/Q+fEr3wPFoyVT8FvWReVziaFdx2tPNpRj7t/0ZNylkMd1r+t5VaPIlfkjLNwmMZ9
ugxMuRjtJ3qu1vq+cC7fvgpSQUkxW3vDht5LDcPhkvwIrGj7qD246eqW3s/WHliBFLlN8Tx/tw1e
G1S+OM4xZtK4qDz+TZMMWqQUDlhVlItW7zB0KT+TqZKd8ntiF9ovQWF4AzlAeRE5/EXH/2ruZObh
dzCx4KfmihvjM5txT9wfsnwhn/eRMCCGIMQrTpTF8LPn/PAnGMU9BTQ6fggHctl/0hteke6Xngt2
z4JdKnldHCeV/LXxHLRASKqemkbaNrvF7hsVdTNXE+kxjqu037kC9mOBCXrJMdKohcSvYvdeZt+6
uPmDBVzXogE/+PnzyEE7vvq5HJIbp9uPtMbphLNLJkQ6Pgm5g74RlH4vOzpp2dGaSs/KgGU/Gy1F
vBaszgeo3w17+OorLTgd0KQ+ktxLFcwul2wcp6nhMpICwGXsm3dM3TFQQg7T6tGfXZqOUUtAxwHe
zydkN1SBi1h1na6Xe9l5Ry0R8qXxM8P6M4K2crqnvClF6SyDIyrS+83vVMTbFjovFhbMDmZqx5q+
GFa3ZbNy/VbNRcTXDqRA5H3/WsXYlvRp/mcGObg9yYEWD36y0ql9VSZsuAluHux8kvBHCiLk7IMs
laq40wa5GwSlEyIJJzeeaMeeO/2h/vGQZDtBVeScKXdhqeUaTXy4sVjwxKkYIhMTKfWgMuKbdws0
u01dTMs/stOrqEIJY878P3P6k5j7ntlzAvvQmLXQNigQALdBJw4uNjmZsgrzY1tpqWQX0HLjo6Em
Yy3XRom0OcdTP+quz3ZfRdViWcp7yEdx4Q4PR1tlBB2ZG+CYcHOeudTHOSSOx1jXshHVKJdmn1AJ
eSNgjCwfVe4t7ZLKeoFwbReM/tR8y29cEExYBtGyjOHIPHc5Rs/WdMLIkdbPbEWWZXNBS/tTR5LA
VmlOyClZoQ6fMt40qt+QTA30Uo7/RmNtW30YE0xQojX5nwN0r5SoevR7kMLc3y+0DccEWE/mzGhf
PYj+ju1fozbrBqry5elE4ahezCBvOgQyeBsGBMR3oiLNUco44Ad1qt7SgMLUra2RyXhPcXcsE4t5
K4xOt7aJf3mbBp0CvswKLM05LqUL+WCCv3J3fVofeyndQZDAnLh4/yqbnJSzybUvxmZuzJBGUoqO
qupTyaqkYX1pgBqtqWpARiMiXwkehfODpzWSjh4/U86CYoRjoIhMEYvCb6WkoA1lb9gl1T56DndZ
8eVFbXQaPtSLFy16lq00HWFI9jbH50GGCGQaB3OeqasVdyPsdF0VLq98N6pyRsc6ELOeWvTqri2Q
nxPkZmBkkhQYIh44ssjqqIKZGpAiAMxgINKHQ7Ek4/EwVE0jGBo/WQZUZ+uOcwg6GzaSL7XQHYHo
9Hs9Cskg5dTm0BWOF/rOcR39gyZ8jYIkLNwBEsN6j8Wz49clakgQnIOyFxz83ieCJQdMqr9qjVcz
WirM1stFJMJmZUXxPPGSNVQfkTAk1bpFRkT/J/pjNCifqlcP1FefJwPxFeev0/2FBYxRMwf1nY1h
bdvVYk1ID43ODtyHGNgc6u8Py4MzSqk3tj/Z5x60KMtUVCYJn+dRWoTP4expS4YKRO+SRaTlpAgm
wJGTPFL8LS7sbPnX+pclZqFNC5n3LNT9IMg3l9w0o4KtuBucFc/6ldTlrYVsk8ci5kYJ1hat0Sqw
dt9D5dSBgcAQ9zMtAlhLCG9pz6dHeb6AEgwiAOEdh+h3bRmRUmBfrVA1eA1Tg8e5uVTrmNIiHaBo
YdzL3JaBxt23ei3kA/hKsiONVK6nnEFvxNiG2H9R1txqbUsOJpGyJB4/MrOrVrZQbCK/+bReFPK/
TX/2j494AH4iNaJi3/fGZuMrgVxJopH/wL1ljxA1VWhIDCJl2qb8tiueD5EumjyXA82jo+iCDdNL
Jtfi+q1ThHsFjSQO2XJymiepvAEJsRnmKDQA6V/gEvoTa0OexHNZbfi3TQrCyG9QCDuWcwUTueNF
TYVAPhhamW2fPuh2WN99Ze7w2GOGJ84QIs9EXPOk1xx3P6G/QJMXKgzYUuDRfgDcxk+sTj+LJHKB
l5lFjI6jxnhlYRbhbWU6Xo5U0HEXqwTp7g7DBkkLytLGJu8tjtLWOzQNClr8RLLe6mkSHHa6OTfl
bxAzomZgw+uqlmGJa7E8UVQpqdCMuQL08XXe7tH0tVZ9cV3/2mTHsScJAywMO6WoqgEgfuoeEA5N
oU2bz4KN1q/NyKaH7wCbmNJwrzzbGfJLKBdtJ+nfHM5FKWZn+TYrt1IYW+5vax23zBfxZOguSVhZ
cu6GBjXV0Yf6pvBhBng8kfMxuNeK5L1kwbqBZ0Iz5DREaNjQS709Gnqs67vI9nH0zHHMwg8hvlKt
OaFtd7D8tV/eb8jQ5AWYh7sDqI7gjtbw+3zwx44Xxjy9GOcZueuwbPRJ2h17swXXohNt6Y2nQf48
KJ3JR+ACShGiFio2hDDsEiEj10abxcXbmI5snQiRnTtWmXI2+3BzzNkE8oZAMvy/XBvTe4cPol5U
nwbGjD2YawMw2jvjjBrjHA5BZppZE74VVkDUeUy0soXVd2lDfnLJ8BcImE0TXwVBdUF4GM5ctjzg
4wLOgOL51urmA4TeRRAKKP5uylftXNWHAlwSHDtt/dPfxRAD/VptI0MlnwP0Xc3BWjfDtfpNXBnZ
FO20o66QVAYs73Q1sbF8SAxO0riDmAN7S1yD6QZoM8auP1e5tWBcs0zgBYR65EMACIlAWri3GqrX
OE+X4HvsvtXcl6OtUtmdIIubeF2MGhF+3E2nam9gsrF/r70tKI7wOaNI7subGzdBOKI6Z6Y/scd+
zkwqPg7vue2HJXLkI7grzBTkVYIny3yIUPR3w+id7ixu6X5t10Ty6XJar2y8QLFq3ccQDHt/oOXD
8ATbAP+sfINerhPquF8FVan66rFyky/QAT3v3Yg5kSGudXZYwlEmZ/ZM/yRV8hk3VuJEsitYL/Ly
5rpHrW+GRWktuGF5GF+HMGanwi1hDDrwlHYZhlkPPajzXh8kYuwnuKj+5ATrnY17alyTppEdb2jv
e0LBqiF1STh+OjexMDwg0o3qUENMQPXZRY0EaOdZ6kHJ/sxktXlN6mG5xvuPvfUbGgAWaGWprv4m
HXIgMOlAYnIaUv/yEVOfepxvh14I4mCppN01MwXcgMQ/S9KHqGnh5SQXs5W7jcOINJ/R1jubLKwn
ISs4LeJTAJRVA7PLOZsxZxMZnVZmYJmRyAT838755S51my4bvHWJCQm4V3fZ0u0ou6Gq90SlmX+b
zmZ6nyH+A0nluhc1R2nV21DWoUSJeix2+5McrB+40/oeFtIglr/gImpwbDb97NwCS12vo06txceJ
dltog3ywcE3RxqpggkmO3GCTY8IE/QEoXZ1mt8cchHl3x1yvYyO8/jwmbWssvnnUr9vg0M/J1/Oz
swUJwbNbQLVrmpP8NmObTTQgPzozK60uzmeanOBwq0bNXN8L7S+MQvSFH6XVa4fTgT4DpiUyltNe
D0pjzp+8xICGMB8q/J+rutDYpJNj8+Lg+pRENZz7Xx37Ppaf7foZ7vdK5A0z1Cakotui++esu35H
1qV1UJ0ga4hIpECFIUOqZJn/8r8LTPesV7/78sge/WALtc4T6pd1KXDcdDUVPSfiBvbSZ4+Hku2F
RhUfB+4qgzrSbpTVyA/bqB1z8PNGThRJAKjVkJNWQmLx50FWxxMMConuOWuG82YVx+nrQOgZeUtW
F63vV8WF7+LslTavje9WhRFqW94M6c2vXQnRiHNBK+iX1kRLPm/m37AeayCSLnxrpCMvK/0O4CoT
LKH/WfK1A92lETbL6llQE6Ejdxo/kqbB0r54exBZYZI8wHZJYTyw9jVfHbf8Xzl/I0ltOv+HazbC
eU0w4yH4WezZ2LDKf1BXR8w12WYDL2SkA10KGPw3ndZq6MICPpfEJueXvng/8NXoUVEav3FEdGcb
c/Z6vhMoDFVeo+1t5vuOcOmb41fHaOMZGaT0md6GLPHvGq850A3hVS+khK8quFFVw4TypG5JJgqb
DB+enGXq

`protect end_protected

