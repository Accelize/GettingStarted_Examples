------------------------------------------------------------------------
----
---- This file has been generated the 2020/07/30 - 12:16:26.
---- This file can be used with xilinx_sim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 4.2.1.0.
---- DRM VERSION 4.2.1.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinx_2016_05", key_method="rsa"
`protect key_block
u5LHwThgeDtC9gQKSBEO/0khBk1cdt9vNzjTjh+cLJYDr6F8TvfTkc/WiRI4yR6uV7xZe0aFJLQ3
VpqkRq1VxQ5M3EQcYtY9EOtKrtT4JiOZjD9hpIlwLczo6sQH8UWHMFuFhIE+39jET2fgU50Hh3YN
/CuZrKJY7TtVsLaHhQrSePlj7NsWa19dlGB7ZhWSbRy0EIHKc/QdyY5zBgK31wUWg4GsH8UHSU2F
j4MCDUOKGAbXm/5iBcTR54H25qieiApfqTkK1IOfhV8ZMGs+BB27GqYkpPtbRADPaGNOQIbitMK9
US6zbdhjUCwFCBp54nINR1/pmbqhGaMNUzwMvA==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
cHY6YvIgM2Zd1Q8J+jB5Ei7x+1QcKPapvlOsPFz8D7CVuEa2m8F1BSGezLHUn6ftf3QQeHgpseZt
X04q3AaWQBUOp05zl0Gy5dy0B6JgNwr4CuQxg/S2Hp4gA9KR5bePAmlKAA17kQCY1oiYxQi41aQO
v4NI9yOHxnp6+eYINlDEsqAkiA8v3x3wFqKOfcoE1xR7jsQsmEYTQ+EuQ88eX6pjCgefbIK8OI7V
OhwcZtokOQyySFz5w/vAwuMhgP1mld6lDpyU7PltZsVlsuJ5qg1wJnaruf1rERjXQoIHlCvoLh9R
Be0KNEMUAEnZsspL4vaJxmJX21P4s7UImrNsLw==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
U6R1VTUJnSY3ZD470ShBSyBGub9u3cJympj1OwD3hy9vgzDulS2U4fiVa6CscjS4Y8TX+q5//AAB
6asixdvnyZiS9kBZmDXwi3XbDM7GFZTHqgqWTJihrTRT/EyM8tu+txGuca7mRxiyEHt1EouywHbE
JQLcZbpNOg2nAXWdvrzx0ejzq4shFT4SVeEH+2OwNmOxfS2AqKefDm4mVdq4tnw+li/0uisWpu7l
/xmQ8PioS1nsbNBd1ACxfBbbiTpTJ7BwayWd1RPq9tzbQLAdDWxhPf8PG1flbmRUP9ZLn5Y/2le5
rlUOy1yrxX921j8f6TZTBu9lblgO10luOJZLlQ==

`protect encoding=(enctype="base64", line_length=76, bytes=869344)
`protect data_method="aes128-cbc"
`protect data_block
JaFQtFBhtFJVTxfQI8henex7afO3gi6M+VgjEl3sZ7r7fTSh9kZvZzgBqO7pmYt3HkhlX4OOIg2z
FDsSHVMh5XFECTsodFsW7omoYMiyAABd6nRp0AxkNBMa72uolch3uSJbk5VWcB6URnC4DL4wqn/P
N1sv+DnnuKXlyBudznTg03DCC6Z84NSvfSLb7s7gVVt6MWmpciJYtgP8OEFrP7Z+y2wgdLJTgIbe
KR0/ajO1iG5EDLTQ4J4yiJBJ2HJOsO+Vd2uE6+ofmhuld5/60Gcu0SQncBPkqUOHOQ1Ft8xxdLdl
6fbVEQXrMxThoVvgpI2MGWT68HqpF8WMnjbnCTmGItZnNUkdeck7AWiBbzvNSyYzM9NvRdw0Jg0o
KC2uf+Z9J3KnqKloegZm6a8tU8QyVEaJrf46bA2+5rzMstpvzaft0/1+6k5+SjxUPBAE8ui92VOe
x94AylLxj3eEBlBE/Z3e4wffZty84GJ/dBSy4ogrS57iOb6V94n7rfD5S3cDDD1MxQO6WiKARbNP
2t/sz8ZCfEeGz0PHeYp0qhz20UKU7JSRy5tCUNRm7U727m132Z4V1/kyK8PFOOvRn4Dhy+YqKRSQ
ZctZYk9yOl4MEOGi5Kyer65o9epoeXPJNpIREQOO5/+tCDN56i5wWeOATQ+q5YrsYqkXk3G3EkM+
4u7fdSwXG5gvvCBTJ1yLbKNItiMh7CVM87QWZUbafRlKBGcgFFuOpLDvAop/RHvcyVW2jaL8aBAd
NED7si4HwAA4CgZF8fxeB1F3xeBSnEiiBD/IuyX6ED9RRcKINJqZD8C9lBJ9vCNyC6KUwZTiTU1l
JpkMeexlyYLMxNGBUJfy33vAII5XnjSX/75esRzEVtcADBqShV9mq4vPF2lkWZzXqHL0fv4JM9g0
DcuelEqvRFhSxbNx5Knk0T4sWRyM/ZELVvbJN9sKMy20CeKI3AoG+L/6ksxjwvefPlaeXdARC2vs
VY8o8A9y86tl/O6T+UqjCx3j7708Oi9VubMpU10uoTAvjJBMFR9vHyuWg4+Rb4BMVEc8vKvhJIhv
E7ICma+D87xWKV21RFnH/E0Tglk8wfN5p04gmfrjGhiUUGfxD/zA2whhEXjgN4Bop/QEs3juF4dt
LJuTbPJojHLW7hBkY2LbH3o1Rp1R4N2m7wZwObngi/DFPBfWgpRymkYs9iRfwZ/jq1EE2wKiMUlx
6rHWnAUwXpk0iAfdd/dN675EcBxoH2K0dDW+EluBeV69nKkTNX7Ou+TSGT94TcnqslOE3ZW6m8c2
VcVj3Iu7qg78/PQKt8IRe5ENl54d3vNxzgGyuV6asi77U3nNYOtiQxP19L8PNw0xSIabdvIy3JIN
Mr2Wlwk3ctZn1A/PUXcKr5buP9FFhQm1HfMR+QFBKRlkuDqUopw2aICps67sgRAsxztxJbJt06Iy
m8+a9SCdTLIEFBand6SVxajBNsGiri4v8xe8nbHoVx2yWw5VjqhEMm1TQUscuHgJB8YWAdCzp+hf
kT3U9y9wP8MwuPKYvELxpR9PJ6/XmU6BRyOzfBPTyTIU6zzSlcBboMJTioOqN9bX/wfrbTiRM+qS
q09+GGFmcUkNXyALOfmjyC+Lk+YcJxB7MqgMgNVcCf2Pj6Isj3LDn43h49I4TYOZnfHdUiXSFELX
+CK6QtyUWAQBrC5BrUYnnMd99fPYW+ysEt17B/r4eDJ81Ca7QW85IV76v9xlSy2EFM/2OW618bJA
oCHr+ZW7OwxVCv7vHiTuNT53cBb4CFpfCvYMU3lPaTZr4GdF2WXaR8zYe8xABqU4ZpBKj8rRmB3R
AF5ZIm/1tdGifuONfmHu4sXOdGr0ZPsQgFUoIipn7oxPgWJUA/Vhs4WEvJTKuw2a4QW6YlTAWSXT
7wrlXn3yUVek2Smlfqq0j64B7XzFjeraVVdjkU+R2cjS4QN9zQXuuUgOLDr7WHAVTVkR3/FcV4GM
6JC286XbvIPh91LK+vx6HSa/gDGvV29rDHrGNU58a8NjP0mow9v6PAnFVTcOglETMhDhYBZsoBrk
IONLHELhb7JMCkZZHxbSUKe3LjShRw2v9gi5CgSLGMWzLmmiksnO8KVaXj7jceK9OP2gQKIgeWAM
j/GF+MSHJOozAKBodbWJsg5w1OF5PpYtffAUGH7GFVVET8yHWiZmGgaeI2NMFt6VO5LLrfKsuGVv
HGcL8BJWC/k6eWsN9ht5neP8scpQiKL6r3UrDivP2DvOBHF3nqG4vX8M40ETUxl8kTna8XrvzZSb
M1cqHLL8qoNqtBEfCBR50iSB6G3xd7X40RV3enBRUIEMH0cmluUg6BhJITJOo9XjWegaDv5ZZ8Kq
7bnS2yyOj+XxisN9F3Fqp/pKovNG5D6IqhxDaoJrRTtMsRZj9Le89Q0VZK7x93Ml6qIH6acLxGvy
izBtGzoXQHhwY6Y+GGfGF7o1nEvD4aZnedfiY4aXnTN29GZ4Q2dCr412HjRzl7YQffmjfs+weI55
a+GzTgUw9d9/elhWsMlpMVr5Jof3FthNKXtLnVS8a5L1b67EJkZr28CKQ9Hlz0cLvnjkP30TOzmE
La1XU786pGs2rKNH+wX4jJ94dt36OAhXwCpe7XRp/emq2v7l8SaBAL4yXBME20yFb3a5j23cvLZk
26qoSizDlqTvy41RbtXBHynXoMclre23Bm8eLl8JdnhUbgk6adIuTQRqO0zqfg2pBOjlbPnoDJdM
iLCa6oxwlyDcnRk2O9jAVS3d+XKqiXF1imcnhgfpc8Gl7QT4aZEQmMt1sPbf2C/vTshqTANgQNiX
YdVgAVfHG2AC6IKxickEXZlkDLTYy8WfF3vKJg1YiLjuCP9Z9qpRDhEAQBC6zGzv0ijmWXPL8mJu
/weA38UpjBfWaL1VtylIdSsKwZzQ1QgvbT7OMf+xwKf0aMHnAIVR0Hnouu+ZqWJK+4iJcgQzntWx
uRKdWLcWqWkrnqMNquFRZJ3upV5CpYp9bBo8AhXZ6OGqGB+Q2m9Obt2GpK1XmL6zQnrN4HghrCW2
1s7edV/Qh0vuAMlzvtAsPzb/ULAXKhnto56kgZXtChpf053xkAmNRCTDr3gPjyjf6OvrDsvlLKvh
HCChnNdzlDVlvQW6qrgrUFtyHkA5J5GkndUdqVw6gT1hj9sLMJ7jZYnQuAqNy/07rm/ODzusjdM6
cWvp65ySlzxtTojv8Hw6jgvID+rhuWSs7Y04QYLf5JPPU8mHA/KcHxTSJzQGiZViiHAOoLdB3odG
YW1+ujIhUZnJbdzmN24gGWlUEmPQetHnjmwn0J+efRewwPuUvPmALpC9oFMNtBUssms5rECFKf3C
NBXWKyk5RFRp3DlzMcnEhbdamo1UBBUzZ1D5cS4Fw//fA8Q/AcmbYDyp5umR2BpwnYRj3tADJnQm
pHzgOadwIcwp6F4BPTvoNKBum2c6v8Te8oo51E1+vHim+xQAivZEBf97BMYlPOUWHAzs0ZNjRg3C
nIqnHKf2rhm4ukOkVG+gfwkh6ve47ObrjijTj7i54/ket0nnOjTDOh/Uym408w7RjxuBnUD391UU
rTin7EFXxPCae2XBObHZSBKHNhRAzdxkwm+hhS5a8NQuyQj8k6siKWb1/pDYDSXvxrUmi1TGTaDr
d69papRTMBX+IsgtXRcCWrCRgb4kwilxe1YcOKyNaQul+BXAZiRwKmF0LHuVXgIacpHxF8tPM6uQ
pmkfaL2KhRsdj2u59iu+vXqYiILqS2bOhCNCts2DbktoQqXZaog9Ehl/+GzboNwleBwO/y+pSPq/
FrYcGtqPo9SIv63Hlo35tgrjIU/vwkjwSRowe0AQZCvySPoK+rhoq6uZIkiONaRzMuDyG5vhp/DE
xTyvRdHp+9Dio3f1tknHLAMvt53bbdb8lLz88Ernw6qxAj0pptom74bk8P8IWGvHth6VeEI73Tmd
27ZyxwLiFDV1IGVpGnp80BV8y51t81iSE/vvix84d+3o4GpilKWvTsaVx8IlnNGedWorcCNY1cKV
WDsXbQ/0Wh+rDkE6JAbtHYzYbJ3eJpiu/121c7r/504yA08zq+f+CbgCqAxhe2Rxy2iIOvQcYgnz
EZ7WodGgZ4IO8mqjsr0RkRajAJGYl4Wuk+z4XczhQ2jkBuL0prCwlgwpt8RuJU8mdFITC6v/31is
srlPXleEBTVXWMf5bBrLBx5VsBLuGE4RiVou5Ohq4u3DDrUJdBkv+ba1xuRFiswriY3Ovo+V0VqR
8+FPFyj/iikVS4WNWQ/m+qhSN0Wp2SbZ1tkiRvHdHc2FDlTsim9mXxkce3azcls0v4m2etnJko3J
20aftfE+cyQ458u5fu7wnCmsRDYJP9naLAp+PxR3S3SZl5/qWM+IwbCFOiZYdbEctFoZTS0Q6XEF
kc/Mo6KgakX03c97V7lkIFCTxVG4CRArCdCD9seskA+Dl6dpcybu5ByNhFUE/rakGZc8ArUXGUcJ
rZ0DD6Mv9Sr6UCjzH7LOx9i3tmvA0d8S+5tnwji81QGoR0O1Q38ezUIWem3Sc4A74L1cSXekbDlh
5yuRWJ51YmynUqAyV6aT3oOgyQi18LbYsFGFn62e/ePvqjKA3SGTu8S/RCwuPFY4rJjJOXwo0t3F
hPCB6RIhwq+aZVi0qfg1m9YX7P8ZW5+XWpsVv77eMxBlMnKNDDbTvsHMR2G8Spae/88ZudQvIEkt
GIOnEhfxX8yIwhxUh/g8zfFR2ifxCAMQ+TCxxnQq/ZxHg3d54ybh9fK8Kdx7eYBikkOz0WCeySq7
RFOeIDQTiHIUYHfj1/XrQLlXo7TZy1tTXr12kTXzP4AOCHjzXnXvj79VEIQbHBQVerGM8XLjr1DU
uYVqvkb5hLNcE5bswa0cYlxB1d+y+eSGdwYX+F/6zq7DF+5JHcZnb9AvklOA1lgtxmaBHEZH195Q
1vRdlSZrk/3Hcr+9UGmRGTwJpgtxxA+hN53OAHhzaWWbhXdfuMmTp2deT6yYGgz9fNxtLxgo3HhY
taWkKIIXm8rFlgMMtXT8IHsLvjJBeOJGeAZq0fGTefB+sCnRSpdUi3j3GPs7lOhh28OuekAYjeAr
P02WuULofPoiWgky6umZq4tBrTYqNRNa6RBLTUBI9xiB+EgA2607Q7qFG9hTtcv1/KGYDobV1d5e
V32bmu8fwJtjTwwJolJVEIGbhnsPI/SWsd/eZUlv/iVu23Fjuh6QW/dwqsDgkfP8BtpQZOwD67dv
LleSO6O1dzj+bu77BdyswMCNJAQcDvnxeQWN0hbhLICdRycaT5Jc6uIeQoKyQraZrszJ8b5tin78
MlD24VY3fesUtlcD+ipTh+rgEjNiHt07LWx5GnTFADTxXNjys5kdL2IAxYoIGj1sAM/vwOpUIerd
tycqFDL7EvNaY0+vRHQNejDTcdpxhoZIoS1Dto/vZz3R2XrdWTkdF0SWcC1F03ehHd6EXheWTsg9
YNkYcpKgtgWqEDWSiI3EhdRzWC3VxeBE/Jo046MtyBU7EqQlT1yYpnjULlg2mNyhjnJRautTgFBI
PsregcBWU5V6qxKsk4HTLGB/i2FhQ8qDN10GKtEtyfBARNt08oSYc/XDHCoQM/el2g1K/VMwC5DT
5aKL+hhEbO3tqrFUBqq0W0ibBOVogMNF9SYL8KzZ+5J7mYI0StKXabYLy6VWUaC6klytzvrG1lIg
X8UO/hwUqLJnowNj9bX+YP98aajL0+ZDcpvmEVQYRisPUo1OXIDPt98IocObOKpM4ZVFTjsvNyyb
zQcxYes9vrhIiMr7tsOAw5Q5I6EHbQE9BazfDN/Umc0I33rwO65fHlZKXZXUql7o0RZbvlpK8Uu/
O/adBPpOlTUIEX2Sf+uN7fN3KXyW7ZZPe9GYeM5fU0E6nt/1hqpX5AksH203/ho4DeAMAFubI7n2
VkGl7pwCtS2zO+O2G6FsRnjbv2jLjv4yLAXjIfUbNWCJNgH1rzxIcGMMcA2nGz6pbYBX+YEIujVV
zHS+XUK6oGLcH40lI0LRXltzo1FaKRlqfO8VDxjIr8oUVdnnvpFhB8SpfH+rf33tKMZY5dgweTLr
0kv84hRMUG1O9lsHV9XIaHqg8BFjvfJFxuQX2ycu6yQug9NU5qIEmMkCj5jmq+6P8G+tLXbHEk0x
9crBzjj4dfXDmvuhr3niQnkI9o6NKW4TLpt0Mk54XRXYrt/I6eZL2nTBqLk82MeVs9SUr3wII/V+
ZXL33M2DRpr9h+ojhWrp5O5xHf6KDRsmAHUMqRgzx/L8wCgrbhknl4Wt4ODcOGoMfhjXDIKgC+N8
98bLWpZ5L9YaSmStOrihS0OmKeQmOSEaMtxujWPuY8rwHbCi8KTPJICA/AJRvhb9PwVZ4Ml0vI0a
HadvjU3qfVBYwljA8F2gTIFaRIl+FESjvd536veF/cDHa/2Nf5KYTjVx8p2BzI6CKyRfnhtDxul3
0GOcoSqkfwB6N4O/dNpeFMO/hud/NUDNP73fWxz+WMCtBb7MpY3yGl1XzNUBWLqLzki6rZAqMne+
Zt3ihV2fhYhYf8TvUqNK1DDntUiu6c2ne2M9wj/IYMI3J5eZn5+PWFYWOXppEVeamH+5BT30mLxv
a6ylr6LpP70zBhkG9HYYvgE3mhn4jWFDJ4YV9tNGYKz1Md9jsFPlG0hXN6kfcRB6YJ1WioV4x/u7
SgngKK4F4fST+KL421kqidIAJaOJDNwVbayEj85E2n+ALIZD4BpuYujZxfoGYgSaH6xTUqyUKkok
ARBxZT+LsExlZ2OTr8nygboHIo8BFfMzIvO/9zw8LmLNqXhBvU59FofUkC/NKDCOKtX0gkDUB5tA
RWNO36emWIDbTOF4ofkl2x5y0+y2tsbSENAg+044i8eWnZrwfGOWTQuWhWnQJAjUhCtPjMBL5lSb
ijxeHs55x9PPN+Z9YkcsuAQbDojSKsHorpaafru3YXtbKCrp/wtIisW6yi2wrCZeTCvxL8UyiYTG
/PgMiFcVg8c5Z/WDdEJS90vaJAu9YgWVUvqaXfLjR9o5mGNZnZeUYPuVeJZ0iguPpxQbooMkPut5
3DCigssbxnRnS3x9FyH9ykUPvzD5f44YXrWQIugQ5X3cjSI8AjVPbD9IKtLXLqu+QhtMt3X4fpOf
IHLzzWzPWA4yvVFyAzLs/++TyUif3sJrHHII8PC9lz/5boyWBlAsrgsiiJYJ3xUu+HHH0D+8OKJF
aifGBqxj8Xwajt+r8gisP7d77yquU7JzDdQGmA07qJYKmtCjU5t7sv5e25ZqRdtGe07KZEZTexbc
g1ixGGlfbrRL8d633tdbaVZJabFTY5GOFnGI/Ry6KETF9JYMY750QVQjRnyTPZdaATz80aKDl+Zy
jh+EMmlQFLSyRBitW0GwVFKi0Mezs5kh9LwNg2+yLBcrILDrTsNMJJKkPg97LclnQ50viAzhdlHr
eVPl0hcZynk8Wwk6NREs2O/PWMrrDBYnHQH+rmEJ4lyIR7C58oVTgUesZ1p6YDJ1fuQMPii3a+dE
ud4JkfesmPSMXwxq2G0wW9eOZ0LRO9iM2VGRB0806a0q2s9VsvwuPvoUoGU78Devlo8AgKPHbt1U
7IR0VFuBuvsWFysCIPJgSVGS1RPnbL5eAl6fpTnCV7jBbGx2cGANVY3Jf2vlO0bBTimcf/O1JhX4
htgGRBC4p9FaUB7ho06SBzmCgNgqYjl4ZZ0Tj01asiqhKvSsE0gGvy6Y9K+zDDBzlHB3SaSx/VfP
Zqu5yURAdx3Yxx/PeSfpIctGJ/3/g7nh8YbiuLO6U4Q4opsal+fnsRKn5NnvdBORZ61LWFF1EN75
dl1qNdvVdN4KTQT3II1iYzekG+yxu9JNwNaJnYxUSYgI5kOgp54e/P44U+aTBg/WJFx2IPfaMGfE
3jc3BZzV6dWesFnI1mrNT5bxOLRj+uLUAAFJpIrJQSWr6ArtRlkW90hszzzy9+aHqYRxtbNqhxID
w+ZbJcwlU07nJVv5Gv6LCCEroAS4+wG1MTe0Qm/GgFSa+MSq/+SwEvu2W5mw9Ext+oQepLbNiVXc
AuXtbr5IfyRE/OI7CuciT7CcQkgaDJvZsNX2kFU2dTYwajgg2Rk3M7U5vXlcq5SB7FScN+3H3N+J
HEBt+JJ3Tbe++htC68lyC7XsSo1YXmP2o7EHZMDZXOXq4vus+1LXz539ylQa4OtBy4RmDapUnI7o
PhlQSPPZKo5OZWMkNOUCqLpHA2B1e4rqxC8YvW3i601I2IF2uvwqc2mLHkFNH3PnY4Q0U+BzWfJ7
z58eB2mfk7JuuAJUVK5cRqxwBaNSG9piudbH27ZXtrROz8uQijpcsaAWf/15yostY7JHYvTpM5UM
5pBhOorxLCeR+98xpTkF+1j25skrZQtJvnWROvcBZdUFQQAqaJprKGbdpEV0Kf78SQwzLKgxszwh
cQ13YCePU03D3pgXGuKnZ8/NpHRcvhn/et4wATS6YaPhsvT48HJbE+8146gMtBDmQEOTnfqg6s7D
draBMjrU8JdgLfxQyPQqBFiKTmvu+6VBYf0TT0KnCzL6TrWwldPHQ7ZJSn/5dAoc8qgzXiQBlTHK
k5ueTpAkWDYsQPlI2mAT8aBPzpADmPjJABI6+ONZun93I0miOJL9cz0Re1a9s+u/KP36n7AQ8XDW
sP6AS/FbEgsGGNqMMhJRnyJjPbdk1Y5FmW9eYfOCIfhpbC6e4A8KdUZbBgEnqaOEp3/hMlQcnWVi
8KvPaCi/qQuCiqv3A2f90DkWw/3pOLUcWu0/9UtROrbei2NYybZS24FVssXS02H18U+0SPzAY4KA
u2k1mGBfFo/F3EBE8CKCj8ogObYLtGF72+HM+LLMOEb3mtD/mzt62f/W/qyWuI6msVwvfua0Y3rV
sAjCvXAoIyaP23qGPEbahF1FBnNouRUrJLcRBDOy+TMOdHCsLnQNik7MY4DF3oVcQvbBj7DeOkzm
3fb+//RicDkmPEJTCnZm5UKM75cy3BLDrd89J/rIHmjHc6TCjVVCspHRONlFcUm6YPo+OXSY2smZ
2eygXD7f7EKVcnfGvlHGV2vzhRyt24YyK2/OxDWlPybDoORLRTHi5jT1jzPgATRBdtFM0dOoJPSJ
Ao1+30agH18gxJmY/7AX9YKofNdonmiDLWtj9adC6z/ePootSFDsooOgf2cs1uCt8IbVL7A7VvyI
n2No7t99zsvf0QLvLpIKQzQnakvjpB9zUtzUctNoK0iyJRBnOgKNaDWm7D3e+rHYwF6rblD2CJqT
0+JQffMYpWPbJy+mVc7nVQIGKgiwjSpp+WPwLniMeTrNLNuyYJMz6HjDVMUAF2B9DZWTh46xIxGY
SoxM10th4bu8/MdHuOWVwxRhCKKud9icnVoa/veb7pz/y3T1Jwo4O89yv24LZMjUxDyVVU5nzGVa
GznG7u/Yj5MgTSgBEfLaI8YIdURjC/Deat32XOUFDLuc9w0Rk4Djr90g5S/k0I6/8RaOX/43LRhR
8rJzYNuV90prSXVRnNhyVRQYLbfzKQhCqTpaEt3hQ8HQdbXk9V0QxEET8Iyb8DCjDNjyvg8FhfrW
hse7jDWObRj67VQEypf7B11wCmfbbePN0x8ePjpczTaEtydnTtDt//U7h6UFD3f/ofhUz5x3Hf6k
WkymdpJ7K4ajoDXxEHR+OzG+axdEXuPb6PXTEn7Fov4BAEFXgNUva5iCUkF0mO3S0MPpWbDXIG/V
jevPepPCt5V+RKJo9MsWT5jfV0mlsQ5hFS7G/KH/Jlpp/VmlMByYdcfK9Sja7beKInATlHOqHoGs
PGTsaFOztY2DkRB2sjqfwh2Q2iPgQS6Pkqh6vagJpRCl70n7eqztzk95tbwedkopEpE43nDN4AKk
xg98V+w85w41I+Q2aBpM9/69xZpIR1RXPa3HuXmgO/Ar9ZYGoLD46gqIYi8+Z3u984v019yhcMTj
HFxZzfeunbxAep1NbcM2ZRYv13S8Lu39fUYO31ikDoCs4el1SZjuSLUJPMqYyEXha9ccQDkHI2of
eX3AA4SXC66oSdaD+pl2+yeqFHwIhbseHd9stSg8AvwZYlODT7eHYOX6AOihFdPi6jciHBlL1HLQ
6zUfdxi1mCPHqublYppb33919bAtJLKwnCbz1d4tJu6TZCNXZ2+LrO1IFjKEzMSVLcDAHgHlg7Iy
WI4AqcxRodz4o1UP261kQrRtpAZKbLKdDhB6crB9xdmyyZ6MSe45xxvPFW9WrcsqrFXrUmjK4afQ
JSjPgnxgjZoixrWsLJ3GMc8MyIq/UXVoDEQcK1qUnESQGypotqupFPNc4IuofJod1hoM69+tenDW
1b22LOtQbPQNQQ9CitgnGmDJllHeGvLIfhGb5FhJcjnuOVeYdh0ZKKKy8/Bgeraq/uavvyWDa0R4
dZCMyjMMTLVt+o7lGYy18MbJnftMjXIhE6bPFaXSlbXaFwASRo/9UWNitLt/F09TcEk6FUD2EKdq
Q/+0DbV0NhEblI0OzweqYgj1HebFS1X2rggiQ3tJEFCLSaoK721aZQtBKXHFbhiaMBLTaMX6Dukz
toN3Cn53lFeACm2pipRItMTNeR52wjiPttM0ixUdbkK6tpYmAnrYEd87UeV50Srog+Z68O/oGt8X
9UlIIBzPoPQkizr5JfGeMYKfUAE/iRAjym5g/Qu+h/xnHDs1cumM9M3ndMznpeiQU2rxzLdeV9HO
t7riP3/bN4vlWFLlZxUZns/FADDndbSaocZ0H+z3ow5h9JP//PTlByXLEfrjKL3Sn6l1gF+7u/XM
MB3NZUmxujm+d17KvpVYvuukgcOnAL/H5xTkQe9kbYcoUkkzXxxnwnRJN5b5v7ye9jD+9eVf8jfk
mZ5OGUyEabZ8+nyC8e7DqV9X+lGAUyaqJPrBVh2Ox5Q7utID9wKiv+GhGwMHXn2LVuW8CF9c/Ovu
1XPeOPZDb5Jh/Le4fygg0nqWeGSpxUHDWoWV10n/UdR563yP02jWun4nNz0sMT6ir0SMN8PYa0va
Orh2zzgV4nE5O3s2z6SSHNj5P6ndtThTTIgcq4srd7Mtx0Wk3qD25SgXLaePHul3cKYSNO04qGQx
5veDzSJ43OD51Gzw25T744s99IIfaxB+LPZ4XmgchLx9TRdi0IJ0cVteXytfCdkFIyLnbYuMYwWU
NLasUdYUZkJOj+jLdrEREpoSHU6fRFFxdsxkj1bOjt0+ADxVmMhtpo/YD4osZpORcpceiAvJMDw6
H5K+L6vkMHQrmlBIowD+s7Ql2hQ/bR/ZJoggfbrIzaZ36LV+a5H9Q1IzNM2fRSYhCoGx93tdd0tF
xvo4MmUcqYx4WtMvJ1QEl1ZmqF985b7Ql4lYRRMXOJmZi+toOkgB0j9k1sCS45msak7GRPqpskFc
SXEiKP29CWvKKbeQAipQTTH2QkKHZKgRHeGAizMH6JGVpVfjmiH+kmAvLYH2+hGf0ajSxKTxrC89
mrrnARiJ5YYOkY8D8IRIdN5qaURWXmTkCjvb0TkWBjkJRSxl8zgFHF7kWZ47LgtkwiK3b+t0YVYL
1TwJ4T85NxBMD4YPT0yb+Xbr95BoaK1SZQ8k5+SEtbh5SWtpv85Tro48Ym+YgFchpBGd99Rf0p68
oriXjSGQos7Q9+Yulbi5+zGRgCE1qKXuuczZXrEmxyiSCkBKQsHRnPUxh6pF7T8vlRKQ1V6QV8RB
KMBVJoTRNEc+qZn03QPWPHH6DMf+qVW73AxZbSsDm0O41mP9z+6J0TuihHt8EFaXyew8ss6tfDnp
Sq/A++LscamKcxpcIByjIgS/1ZSt5J6WvVHVzY+DynbexiB9xunDc9m0qMvhlkvueMPAJc9+tASS
CMukjbGHdFe8DZu7NJKdCke3wrHRgis/L0Knt3HDxb0Pq/xAFDvg/uRlL2sZVdcSf7rm/5bYfCa2
hZjMVOTCGJQS5xJwA38BmodbduBRLkSFiw9MPIHiZFgmaWZQVXvE+4RVowwihN/ebzhsaYA//BKV
RXTMwAaZPgNgLSEwjYlSbSz8vOkzuuMJBEUgX5oCKiXeHgPXU69pAMtUVdoLmaXyl2awCb8WM3fq
p02bMdxiKDGVO7dLujFhzSi8BYFOTS3CFnkKwmRv+CNO8e6UlHukYPnRZn/3xQNjTNTIqh0io5nY
pGigUUAFRIHADpxV6ckJf8//Kdzjjc+Pg8w+6S6WKgXAun0iqSipwltcUHjZYqm6fTXnVF9M4rdS
XyTnieOFYb99oXpFYqeGZhsKO9VZ8beEXB5NiXAzcwC0YLrVuZe81fJBsw9b7Rvbo/XKzb+uhC0g
PmS8mr5R8HHF48Lwc0GMnPfxK0gAPGEit3c0k35/idlpnsRYajXuRwyLqVLweuAGrTaLEIC7iF0J
znoDpX1+upGg1AJCOuvLjg0m6u5FsFwh6MpEH8QBMkUCgYjh9lP3ZH/ff2DcDRO1XCL+ou/eFsPU
clVGRiOQUAG1Nusu13ZXBqKCesi3NHCKdT0zYx0iWzgh9RiZS2SgnZzpc9pyo5vVt112vvIxy01f
qf9x82u4aZnxxN2MTNN0cnIZ2bofVTuaQ5ZFeymfAVXLQpzG0t4DCfgGTgnoCojlcqcpgt45BS5s
qVC1jSQV6Zttcebj70bd0xHUXtfFbqpgQmevB/AJATeyuLZ5YInwN017uLzIUe9qFeQXOSp1QrsB
zC00q+oyd2yOisozbo+huOIakKiMjdhojlTRWsEw4rFhVF4zdQ0giTIWxYrlYXk3aWtuGvgQOEqq
IAMAQXk2D87MoMNawEvYF6peiDVoqW5FB5KPUwDbMea2hXRWMuvL62sQpXuOByJ5/tugqwnPFwiF
bv7igVHY6wPffkvIReTLKvxdlcPoQsMN9ljklRf+crLE6Kwrk8bGYoE/0wT1n+rW2IfoeMzWKJNz
HrxhvYM0HAO9hnePmUqea+UW83MGQi+J4Uzfo5o7weYoxaSwjl1J71+wrxs5LURexxpM+nj42lyH
qSXD3fJ+pY2TDubvYXuXI/cS/YrQQSbpB2LfP8g/wKHaQGofZ2btsZRulmdDs2ar/MHpoQf4kpW9
1ipLrZJ1onV1m4r3uwPPHUqu4J+SFOxr8Zk9PbBT9DttK6EecEQdurNuLeDT4uhJzncV7ktgy8Xk
W2VYEpuqW1+ZAvE367v6MIZuNsA1jclIXHTTYekWqBD5motf4XmQBfIOEBG7RwyOQAgu+jO7lVzZ
wYMYjTBnqyz5CUwXYm9ELi84X85dDkB8m3QyaU4pODsAsW6x0+EB1oIgk9H739QvR7YRbE6ibwLQ
6/UyjE4MMXpccFm3mGBnNi61hmSdfbW7lXL2RDeZ5LQYcCKCBRjgZXvzOnlrNylbx4tVuBMRPsZh
+MRbxwnCht1FFKY2zHzAaKyBkhX5+F9dz0y1qQmmwkQG2+c/FnHBwNQiLb3RXhzEKx2NF71MqzkX
PkT9zwikBzuelikO5lXVgs+pNwvLQb0Hf0m/7wpWYEROcrRpjwBaX0phy5Bs8/UBTmWTE5lRNP5j
z1gLrXKQyG48/AqWvqhmMxf8dPi/CDA7WxoNvewtQIxYpF+GDDAm+Jy5xYWDcKR/yvio5s68YneB
r4UjeomCC4VkPJ9XFYpXZ/ileAJd48IfhdtrDM32l5CpbfUoBU+ODYo0vAWePrXAq2wNnqyLz2BW
MqHcdzO7P7CbZeLxZvofQjhfKwd/cqWv2zE3cBsyJ62tJAtLbuW7ebLIf5PneZh2AgqnvwOrlZN0
8vb2QNJtHlnO2bsPEIEFmzZ08uRD6gMFQJT6P/kwYooVv4OsvMYXno+79fi2LH4id+McCpUrjP/B
7HzlFCbJNxy+AksVOkcRcv465JbDjkmGWkPiMX+MfVj1U1u/8j/zmJRfjkd5sQ+UlZmLUCEGh3TL
uE27Lwx8urp5X4ak0RKRvV/wa7smVGvzr4Hv4ZMdhIIWx8rz6TphswiVyq+pwXh40b/aaa+RrrEQ
IQrFjOtYB5B+A3OWe3h5w/Xd0MbEQ5nyFlAy8vH5nRJiZQpvyGTf6T+HMgiFH2+23MWn4NaPrCe1
dFb0mT4G08ZHppcBHWN6OjBhzRu6DMXpBtW8Z88lL4/ONLOBAWxnPT01TvSJQZ6S1S6wKX46YLck
dMwKrQBzjiXneVOAL/AAMz8A2EfiNDoanWasxBEH1uyMsNRAj5PM5+P5dp9YyzvKyEDJrMOAhcie
A8ssRj238ctVLP75cVHTATy5wL9g1m7ED71HiRK4lL1tQfPpxjEd8c135tr81382WDaU6yP6c5G1
uRzGnva4NNG+sOQkzWYWmPUB0/0SlpvOrfT7+aqwqTbaEsE/HpkYS5ynrBHdHoe2cKBdcU5LmeYS
IS0WAdowYjjj7KUgKceYHL5IVZK020+fCnS/0aTB5MVJA8mKsnRCrl+/qP6qVDSr6gCqhp+kOtA2
kAdeySR3cjWkOCQE3WMNfw5WntnSiRkb692jXo/tBOtUIMnSlv1H9DOVSmk41FFMWdZ//J7kBkC/
16U19l0U+utO2oEHqkQVlLvgluKyh/ghxiJ5+gvLJVc+qTaAD7UdC2cuZRHhJIbeuw1mesJDR7dD
W+8x/6qBrtWDqnV8AKaLgqeeCWRO4HlfwkHE2mzdjW+texQ6XEsO55o3BSq7YA9EcYoRhkFXwgjj
BvrLvpsPAWK5WxURclhdTsAA1khwK4Dw4nhIzraVuUEL4n8MOEQBp5xFNSHeNJAzsfWCXb8iex2D
3u1EGPz/4CJOidCgDKVzFMeMkE4jE3qH0bHJyWjZMF9w8IhYOEkGuaYaePffQMOdURtC4b5U+Q61
BQsZhhVg6rO+6SCI3NUv9rzDtu4E09owhQINVNwC3h/FghV2i8LyKTyQrHxiuA32Fa371vbM9IZk
vkY4Ii6v/vr9mvqtkCkpTSKqz5q0Dz+2hS87BR0bzX70115DnXBrRbISZDbU3b9rdYksZW77Wwyg
rHFaVJmRQz1OyqCV+w2no9b6fAesrQc2QQaij/hZLF7bqgdsay0zoV5+sjSBeWSl7dnAy482ELaX
Mhy7Xa9v5I4pKqGquGqxwcjCaHQI9/XKJhhKxPENPKxyjt6qDyr3NqmfDqbnO1YTi7JyzVtrfurQ
gVx/CVG9JDNiJbYNbSCWHDatajlRyRn98zdWzwo0sMkMP2++iGRrMrW5IzFjBG/UxVdQ2nb2ALyT
am07SMif1XFy3afacvuiRwrcoa/yQyi5A2VhARIHgR3QWWZVQVn4miVFVtxq5piw8YIY24fsawlO
unOkPiZqM9DLqK8ZF8RAJwl9sn32Sxl/v+AJ85aUEb5Xh3k7uHFbffQWbsRcEgLr3WxPMgnd2hTs
BNAW2+4l1R/WjYprD6ERZltPsRGzdMDM+t9dCJN5y+/mVyZOR3EL79Z3s5pNm0p4yMbo8epLxeur
NC4X4I+lBKzhQw8qtUn/o9kyZNmqKYPuOvccohfWu0qmd4C/jpjm7LMp5LCD+RZxl9yuVPQq1f8I
YpMXanuDZXa0U1nwBJrrsURRP8UcpwD5Cqo23bNpvCn5Er0rMkj31M5Wd4QUxIlL7rL3CKrpjeP/
1WiW4j37tYFOwLL/o5FQdcXypGYfx/j5O+5FtClHOytCMzztMMkjl2I2duQvXkJlzAFo8ItReDga
n1uEypHVoAZGk6Q16ycZCcRmPeJqK+SFPZbtbAP3YdiMcTZVVL6/lBhC/rDdq50R4kPsIxQT6g90
o7gfAOkAExYWjCMr9qcd8qXI7+Kdg1w9qGcTcn3Q/AZI+DUrEm+HwkP3MCu2U5jW/riK72g6UzrC
oeBeenYVbQ9oK8ewajYV6V708ZwoLRw5K/xTI8MDT0WnE71rDG0JfUQ498p8pkxt5lguM87z1dOa
Nwocm69cSL29JqQARUCHZIQvpgWlLm1+/JUlnRfBuMIZ42jwaNmt7TdUqnR7TEmIHsMf8bnapUZi
Y2Ka7sSXq4SJhJhcSRzl1S5njfTfsyKtS6169ZOxyHhcP7ojMmkhTrbeNc/Fkuwe1Gv+EPt3Abot
U5BhTZzasAHqJgmJ4+FdvKTTVCeD89agx8fZB3K4iT6Gry/OuQdAZepkV98Gaq7MFSCndI4jQ7M4
gLhXWE3l+x8Kt/Pj/hODTJsE60gBhOiiVJAq1wq4hDg4sGH9RNKYyN5V45KsdIFj/UTmAv0ZtIl2
S0IokJnGeK8TSQ6Cm1N0OCiIOW4G5aOijXLY1pIf9A/j+QYRDW2N8ejpfrt9ixx7Rym3Gx7+E6Ru
TG+SyoYM9c3OWkIBuPDZur7gLRtoJVVRSQev2WE6OtSr7h1H9u8CZARuGUdIAH9AwY9Tz/e5FYM7
of/zTWFhLZjbeUtZCzDZGpZqF1KVR2PIVWimyI7+wtF0ZtBXJMKS9z+L1Qcgi3b5l18YyRxN1u6y
5TX/vjThxPWi/551313AVn/YYooqkMiZ9QXywUJYHXi14/YrI305TUaZD5asuFWna0aoPLVoG0Y5
qNKHiu7qpxBrDlX7rWLv0ekz3y2ttALiVEV1M9LH2xsw0x/Zw4APjSge55hJVp3F5eB3QHW9CrVV
CO6FD9UmuypvGQ9I4mUcYmgXcIC7vJoALeU0QC7eo83dJrRuPPTtsTCNTddx8DqPT2BwAz9WSkRn
4LRSHXRJYicsqSDLzxSy3f8F7MH3waaKFHfqRJFy+P3vcVImZVRzoDnqBUn3y1AfFPydsdTH9aHi
BHQA/xaO8PdgkBhAtXDCgKY4XGPaT5J4K70Tie9Z6BErbz72qnW2baceAw2r2t/woe8XjCpH5fzX
1E5T4odh2ZhpEm29DYK6bok/Phs2LuOa85lUsPLSb+39tJ8jQAyADhv2FSWntGHZAlFy/h4Tzdp6
YqhINZgVadrIe7nY/v3ReF8Uoe1PvZezNCekjZGDaLDvUct4mLnO/Wye5vpwvD584dXFVYsAbzRS
r8sBbT1uqiDJg4QD/qjqOlqoPcwXAzQlgzxTQISC2L+5r+70ELVfXogj1rqCw2izpCM5vCkRvTFn
ANpg+aPuUrKrOPDHN0VqORQUmCdKOU+EjkioE/APPle4SRl5/NE25dtiX9WQC5eZ0vX6SofGNspj
A01Al0tquHw6riteQBVRDAK/fLuTfENVkkkpqV/+Q9Stnb0zathrwEan3Ho+tzSwikmq3Zt3UCFQ
fptnqsINy3a9rZ6WCAMnlVMbZzzWm/G32aR3vwUwHMhj/hDba/1kU4DCPH7lbtS8XlcInSGP7WHu
8VldXOqRUg5wnTkJbg/s833ZQayZaw4ZHyB5xXtSeuOmVeCLE4pSucgTHsVvziLy/uh2jSUFyrBB
epWOwtYGWb+d46uqg+U6zfhWdzvXd4eY9WIyJxvECumgMQC5iFHj33cZ7YmG/32hu3F7fIIu+mFA
FddhouknagZz1vmqQivmKlqt8mgx3W/2KeJWoDGOJnSCedDl1npJaw1S4ylfkPisVMF9oE3c4Uf6
JmQsGKxThLrqZwhADgKm6L/cohyEHj+r6WxBoDrhNcfaq5Xvv7n0yyy4Iy1c0eo5ryp6n/vWcRhU
fze/jPUECXtgpJoxdtXfrH2TJE1xfvtC3zCIsD74LsGCY5K8wnlFGfgTkLabUu9C7kiz+x5hakKp
7oVVJMxyABlnA+H5GhdTbUyimtnyl/sDe7NhRrGnsrTss0a0KTH85jGtxtWG5cQ2Pm4nTh3eaiUn
QBptdwExP39g43tS4Yt9+ns/02/AWRp04SBt6uzg91CLV5X8Cj7B/ESiq4RkubnWdGfUMgrXH+/0
bIAPdmW3eXfgJSpTjbMTaoonXWSLW/1uFqTAJEcR19i7XPGWKN3Ka3uP6ZMNgMVKD5pEbsr7rohU
w51iJTE6xAeO6xwSfgJ06guc0/KS5yptCA9URnf3WVPBWNvAQlbMdUE/mhSBpcU0Z4HDRc2y7TMZ
bM0FUBqLp41oBzTnfISjlTEPePhzI0ajaln3cirg5gWaoHwz1ztyZwLABjxdAvyktq80XdXweI5J
KU5w4ZXAlz+zafZmE/vKwubqJjoD8SAXkqJ9ZSM7GP0hVEB5LMx1aBcx4SGj8DjXoGlFYSIdVqP+
hE5YW51A8QdLkLbmAcO3+hlb4kODVuRmxK++V5hTGYIM1fVSznFGHG8NptDBufgqahYbE9G9nxqb
15M6/fMA6rQCnfTG1boTobGkzWqKi6e4DbjwehuM2byKTYXWlckkwK1IcvCpypKgE9y0hCr/mQh5
fMz/m1DoFWY9F/RarHHBsBMQI1My5tnSdwXNAtgfprKZ0535ecYorMKyy7Zc3xQqQ19uTUTGJynr
alPl/yJPpwQo6OlfjK6b30VOb3LffYQjWHrQ7Q5Z+x5s03iD/HGEJfk+Z3+WYNqHkhoghoqSkKoc
Qn6jGDjGaW74OfAQxnlYNmE7SXw3j2MdPlW7bc5GIEq2FfAToXgUH+azVkhdefYv+lHrEMHESpAC
7xEWam0wFzWd+8lpKKvDeM9muEN1JjZb0m8DFKNG0dfG/rZBPWI6ocALIfOVHEuD462o3No6hsVZ
sDnIdOM7fXrr5Zi01DNnCLE2Gqzsjm5zSwcWFztz5xIc1KFNvnSjjWWCgSdZApSyvrGLHDRvo+rJ
0Is7MwY2zW4HcvToIwKcffxA97jqe8mogiqbgwGf0gCI4pBAoUzV0JTuVZ0jhGYYxCa60Cmu6SmC
Cl+BvEfOxhXEjiA9gnYV2R+qVup5sMhe4gT3C7B659x9I8lKzZX+uTeaG6MRM5QS51+0eN2VepH/
8CIuTqbpEKm0PpcSjxFJA4YfkZpOS7HkcJ8uMvVxMyFSdnxfwknfCHzv6WnQaOU3kZaQFtoZok+A
jNlYM5GfamKo2yaScmTg5oZYJ46UV/O9BvD5RIDuwisw1YMOaW46Wu1Csuwu6SyYEGUM4cs7vXBh
clZ2rqLv1fMUhZeLc1dyTvc6V8zoGeJo1KOCzdh9hkMgbO3XnM8FppvREWPjh65Q6Ncx12Il21tM
ZDkZJ8pcVq1B/7URJg6alT5GnStxNgNL5GwfMG5LOH2AF99GNMB+ydK8uh0S2KPQy+MsqttGhZ9T
O4vSdW8KaED4jDCCyXG8l8VQWGV0bS2FlrtN9OO36ZI7eGYQKvzTn1iuZ2X7sLYOGLIdgp5GLmW5
P3lECVYR3Hormyyioig8XAKelO31dRuyWL6/JVIjgBVV/tqbF1jrcdxUydbfW2cFaiC8dURZEBJZ
iWspxmZ6MH9xesMUsW3uwwfDdHilr7OdP8DNonLkUILzAGydLo/h7IGPXrsNk8HvuWAYFLtqml9q
tYltJ20kbjeJvsT+AM926fWRmgNbyoTtMRuxifZ9jzvorhVyuByFMfcN6ZXx/yYb0fzqO9fMKZE1
iljqV/YqBtooHkSDUdlkLJHSh4JHMN+E23vniXNNqFXbpOhcbsppldIfvUegrbfNGwpkKrJ5aJ/g
lKXmtNyNezY6VDxsBqiWgR/izXtyJruZjfgdmqwN+oCktIyMQFoOXNxnChwKzAWcpgN4LlLFIsUe
fF7oTwWLlcPCKhJ6Ize1BMyaN8FtZyqMudHTFtFHa1HrC0P7Dk9clcT2zz8jhuhARp/BRplIQ3Km
DIDbXB8qnvTs+8Lq8jnlBYLgVd2fCAP5to7PaC0ftbG19qtCOnkHgWajOaNeUpKasK7edUKU5l9T
zMhXyhVG8AIR8zR66ElFgNQBz6ZoGBxDsr+RI89NIWeE7OK8uo4B1+RA0iH1IZmzZFcA05ysqeG7
aG24jRwXlXNABxeDR9YLBAVeT7dtNl+by/sa1BD4etFwS8yK9qpR44fQeqpXinnA4TVLCLLd+IVS
UM9bgBMwsVCIDkYHlDafx+3zZIUA6R1k6BoZSFuajzXeCMvtaECnUn4n3AyRElLzIYVFgmzD/Tw3
qpoVfyHXVlxUIB9OnTQUQ1ts3Y6R00CK1OE+Pxl4MBuo1vNf+BAe53BVYyQCSDBbMfdCaltx9inc
865j+WwFUFanKxCmDroiZJ4KZNcUfDKhdFwaWoX9faP+AMZ4qNKTjwOBpFALPrvA3co9BNn7C7m2
CF/iCIT5/od85uzeLOKDIb+LIx5xaKEzilujuefmETkuzN03q9E2kZSkjsCuvn2pwhhUWSNAJjw+
fPIKa3E8gnxfPY99K5taerxpwothznoTPs9ToNkWY372riC6/XN+kD5GzH1v5qXopvDKIwNMH0vR
tfl3RzLlNNe+b9zK0Ry9JPT8QmWm2iXnDHuTxqqM3WpQxF1BCOhu7VYr4M0FefTDWoCq8grnVMk2
rjuX7kL/YIV7Iw0UjuhW0NI0PrN2lDgXqFiQUbK2E6uhtw4Zg20EqnRtZjcP6pgw4xs4utEAh8ya
yvpmzHvN7244zGDymOymQFP64Oi+BFNDtMwh3Bc6WmtpSosi38w+1isc8pz8yyqGaIarLvtYGjZZ
OpESJjwm5i4ycD5SZCIftMW+zZDQpVin8G579ckHZ9y4978nK+DRKXlQbPwattL5g9CkUm60S1kB
F5emSRWmwHDa/lnK3k/satL1gJKroKRsPXyc6j6+VKItQBX/6crJWyKxQU/J3uGJIdALt8C56k1/
voQ59an8FcRxbO/hzE4PqoDLp+W5IgxXh/fnYRFeQTdKxsw4cZexeaKBDlS4+NUz55IbFB/EN26N
25nHSkp1/VKbyldpBxjWdQKeTM05oiwQw+c1G41w64y9LPUorTvLfHg9j+kwOfxIHnQ6oQj7t0w/
v6xTkNofT4PYHCpOAViPcdEMVt4bUTBLNevyuOQZePXcAX+kiAWz5jK6No/tovf0wAiOEHcae3k3
nMRprFwWm6t5U0r8Z8eCR0griFMq/r8ps42/w1aYWd61gqkWPfbRfSYdctZ82x5s5IqQkhmWc9tK
o67ffg0meG4gOJHEW0nOHO/Fu6K8PLVFXbo1Z/3kE+CEAwtJukzDlMIaZ/KYOgZidpzBGkJqQVab
vQf/vvLOAV9CzlRR5fiPnXQ30xzNxx8rlPS5iS4Q9ZHnrHggo+piDza4UevSrycpSRrLc8ASTanS
GoLmisvOyEGdBReekAyd7v8kvipChMlUuJr78DezvKjKDyTBp0dyyQimCc2Hewc3bBOPZR/OzlPf
Ixxujsopcmaxxoh3z+dvEFQ45B8jjCNEhy3CllkU+s31/9WxdxehRt25iNj/JN0+Dxra8fCDd+aS
usx37OFQqq+ZcPokxaheRNaFc3+kLo06c5QOghm7vggC9ntWzhcYLTkw1nn/HRAWtRWv3DFEeHGC
85Q9TWWiESVQeC/qGmQrLbPbeTvnjBMs/suPOXXrxxPz54K3QILpMyNC6B/VXp5iToUwIcDxOFDY
6AJYpgrBd5waKe3KlghWXj31TA86z3+MNPcJjfqh/up/5zWYaxSGv6v1KLC0+3Mkep86qWrjWOsi
bna+fiwvPEd+NGsTP1E1zgdI5c8PCFQB9JTwU81A6VlAmkSZl1QeRNSm6GC83JCLzRFRoBmNovuC
/mxYyYH20Dp0uwHwHmXdR0UUW6LbVlwMOdiUZ36XB6Kvk5il61jNjXmkbJsqrZlEmgcPRAofK4f9
egFYsAQK/17TYnDj7cZpavA4oS4FlrIRgn7oO+YiePSjFP17qXeudbxrYD8hLn+NM4TXkRGyZSPY
2OselqtoJO+hK5EyB5CheI3+LzqggeKXr9gWpgydNcrY+RiZCV3NDZCrbtOp1YNJN3qaoFfUXFy6
PYQAyV2EEVwf18oo2WapxuRuyBV8zy2Xyp6DjA+9gJ+e5x5zOeNru05IC0bamxM5UachEPurQiEF
N3XzgbhnyyO1gjF+w+lrxNoeHztGLzzUU8zHroDbK5Emat1W3aj1WHsDuyDoFDW/UhOFKSeTjipD
Bs2xccQdm83OnKZ/T1KWg5dJNRjCdwwZjv9bx0HtuhaecVWS5/fN1jzySq8HpQibIty+T+yGsYyB
RpwCl26mLSf/EuKExqV2lq+SqabXqBNPdO/dUGIQt142CxD2+cknYWcuqoNjr0kw7/vwaiDHHeN8
1onNEqpJlLM00Ru/yPUxQLPYAKV3RfC+fDnmfWB2ls7QpI6Wa+aldClzE1VSG+5uRTG7bl69b+mN
pr9T4nvYpvjpn/x+c3Tko3h128H+HPXNFxQMjZvSIissMaZRnJfeJYEhcGeZ4TavWhoHmUCz6aLi
ZecqiYJrtr5oD8tWkZXrkaTnlSogqrABF8hJUGGVViNkEeYmKSPCR/W6y0X3eMMVK4aFd0JZ8B0J
5DBio6c60GAgYSWK5AiyFQt5tSxc7FNWihQZHaj29cUvrkq5b2+QTNE+WVWcGJrEqUtR522NW/Pb
BVJjCXlWZ35vOeM6V/T2BxEAXrs24oimtBoSR9aBqrpREETNbOv2o95q64z7nycseKzuFP7nnKLY
aFARcnsasLEMu+mt6uMEt3JN7CdvbrY1RjZSqh9MDi2wHG2l2+8Jh9uHXvBMcN3SaW6ctjB26lSC
nuoxIVnSDpTtLsror5l171LsSPYPH9So9dA9S9aY1Y83L57ony9g0c5cPXYyNTpPBcJYb6ljPvmr
66OkQ9oa/zk7H2xvsOoab73tJTcytOHNXXU73OV6XKrS+z1Rg2xtEPdGhgpyMnQWcqC2/EOxBz7b
p1NjNv+dbbowWMx2lLXrM6KVrqI5lAQ5jlntI0uWP1L+PhC7gm+8VrKFH2LfBu3otZkPIRmW5VFH
DbAhJVsBL3W/aHeBBsIyQt0VveNZMjKxs4FxaX1rYJiJKUe/tlQ+61g1BI796qOfrP2YYbyiMeFI
shqytQwSizSmGKTc+j5tVUutOj+1ZVTGzmmiQDqJ0xvqmm+HbK9SPIh/m38ffQDN3PWxunEnoAO7
f2rOBLejsxFL11pQKxLsSGUOC1ievmZf0y3z65Km4fVDlxTB+PSy79JhJ0oKWnoWTP3PyrzfxKZS
sffjPtCKYGS3WVzbhcKLgw7NgG674p2oG1EO/NBFtAfyf16PMTJ21ljvx/mOsZ2SGwIOTc5qV3Md
WzVb5mgogdRGMlnvobZsea33BSy+ybuuyp8nffH2CeoQ3GbNPsFKjiAaqkXmLmiLiCUw2GaeNz9z
Rjb8/TSL/IQLlHhHbvI+LYN3ggVG2KE4tocqi/eitNrW6QDKGlx5QpXCDNyeIjOw2J5yRAMh3DmD
2QeQd3Ki0ElVtpagVWq/cI2EI0e3Bd6aYt93KNc/L4/etDcM/JvJyXSLGo6XX1/7sNXcQRJ52Xav
nmLCGELKTznOg8ul/RdVxetOw6n/an7lYwLZaX79fmCXni9+JEEqICNvF2clirFpDkXPQaJPxdXc
/+bmjGCsvv1wUrjgzg6g3JHAutbZ5eeKFrAReAwE7yocyOPjM5XQzNffpujQh2bCnrpNYKqoaip/
FWbZbOLcE8b5g2ybZenVfOKtSZzvSGFRduESKtopErk/Ll3rjkWzzLey6dkPeUmK83YGOpz7qbla
GNbRzWnEvrQ+Z7a/d1QxNzqkqoLJRbQVfIk7S+peXdnKYvxax3afs6WE7/FucbKHShYNC4DHDb9D
uCQl/VKn/ZuQyA2BYxLFeqQLWECqqicEa/IKBJfb/FAs3YDojFYDaroFrSLvCdc7Av7Dhg3tjiX7
z9F9faUuN8EkMs20nnEfS4jEQbB+pZqFJy8ouOBOFHPhySr1PkVfkomR4jzPLRiQsn4Fwq0CTvOH
c3jxufjxn1BrE+7qMZdKt4ISIRkLUdzwVzZGpPl8Tj/g98pMHeHY8dGMrokkJEmF7qyUfwik/ZRA
M+FAD5eiAjR4fTrONH7M7G+c+Qyzryez+xc/Ry+ux8QVC3sc4GiMWjvfCHE3MZr6vmekE02nf05n
vlua821UtRk/Ms4Pch6oYSDjVZ58GE8R9/ilc71B0NtZQeCViPD+VLDpmEc1nO6rq8Wc/9jqxNnL
aG+wocLDXhAkSvNeHgsFt2XPxApticsi0A4WbadNmmgw0YsYmri9pz23G/K4obnL9fKQefFVpGwF
nmYw31lbRx+G4GUO7In7uVvzYGxDOn63jmGADOCitQu7i2+G8lQsinydqVaaGn5U3K7GmJyDoo3e
mTF7LNo1+GOwJ2izUQTfSTZgRE8XRj1BxRwsUrVPG80rW7TNCSPqqksQDK4MT2HF63Rq18ZC9Ue/
6kLTffwignhZ5wOPKxHaM59bY3aB65sZJRhEa1c/zod4huhwa8yqDXY8hFhI5W8hYCxpg24UY1FH
JzGrhyImZQNK+0M5CQadOxvcZ3FFyq2jw1pEVx6BDe9d24GlLcrFQXQe92+s/Y1lGkREWOp9K8WY
hzmPK6qH7DQU5bZhxGSpzTvZSuLSdFyRUdFpT7upUsW1EOYdAkV9BD7SI+MvsaurdCKVwk/PLNcS
LJPquu2wCEigMG0xcp7uCw62UByLlmbrixnOI9Sk7/zVU0KxEWT970ig+1NypUX7+jh0lHR+K4EJ
ec0y04RL/pBMwubnzZqS2OjUQO2V+J9gk5pfk6FfxTbrEQO/wBewuoXJeFc1N5OJZ5eoxNWgYDDZ
NlzP0WG1Lp6jnLDchiIZbBI/hjvYMJvD9ZWBM9/Kgup2uEbaQdjW7KD0F4gX3yFVSoIWx2BGIm/j
P09W3lfhDS6og92FPKvRzzmhh2xAvqHHLn2abwavu+DjGfQ0gYP+AzyezOzbPbe5s1k3z9HZkHkZ
MYXt9o3ZXEdPXJS9Iakm23Hwxd1P2rVRszIFr7mGx9gxVVqMHeNG+u51w3+BYVufq35023Pg+yTe
thxXkAt+q902vkHf6ir6RQhODuIAAlEEyyKsKu5QVFXX+mF5l8R+lcuS4kw1YkhbG8lBHDZIf2W8
tfPhdc98aVf8w5NcJEYJ4U1lg0kgM8ksnCvJi5ljHCewgyHlRsQDddU8j85Zzq2j7i0w7mxr44jJ
ELb5Xjhd+E2lsJE9ZNLfJpD5AkycO3IeJDRWx/N9qvz9kG5PIUJ1JpDDNmIJW3B3RMtNOQSv7NfB
JcZghnjDYMaNqvaxz71N5LjQJk2ojpveuM2tpO/jFcYCrFnP88JJIL6e7/Pkdb/tzQ5F6NA6x3qt
LUTtCfWnrvDbyRnU2w8025HARlqqFs1nzihnMhOWFA9XbK1VpoACFYJ6HxxbQA37vivmRjzuXS+W
6HxI4N5uNrRVUon2V6chh/KLD9F5+ltvEeuPbuy9QucoX3HVtmvxi2tztHF1/8iRcXV3ZWQP1hXY
aAiU6Jie8E85TmE2NjMD1RTIn7FqSMD73eNYgByG0V4RURX10XsA7CjTlMwLhvMSBkY1tnXm2tJO
iteDbtq1Vj3I+TGXkF6PV/1Q+xL5qYCCDqOp247mRylR+shNQlnhajtBwVXsoSZuie/uq0fW2SBe
BVkjzyhTsAXW6JdSwRSYFYZzdToAhsI1Nt/LFQ/81yYLvx3AIP1jH7eFk1N1H2lJmryarhhSSxrY
ar6tY2bRUW2S8ZhxqDuzU7Ob3AWsw9WMrI1gaL5QiG9aoAZ6y1f0zeZp0bwJq2YVwDeqacmO7xfo
bMvUMb2NYfJRgCf99KtKeSJRZFnBTQgZa9ZGstyd5iZtU5Q8zj1u/0zzNW9bn76LEztGr4/pIvZN
/OxENP4/VBTN3cvh32LT2nlFnXMe0HFBihCowe5vW6CivUdiZs2RATIZoMIiMxe47MaH07GcFj6K
GfFVMkDiIhnzl0v0KcM/WuPmRyCLe2usBVti4yFTfOocqgRhUFm1ObRXucEGab7OmpVn5Bmi41Qz
AAQC7WhrYSonfq/GoIM9x1a0KxolnW8Itrvfxx6djWrWpzWMN06vEJ7PCnwBTvwy/ubd8lzk5w6+
EtQMzDNbwBH45A/i20ZGNm46R5O/qjmpmY493No5hPOK4ZFChugmdzRhfc18oi+mjQGgRrRPrqeO
PNhRGmbubfO8CRhPjW7dVoa+120WoOaRDG7n6uSVVwdJSjgtsOaTo3MS+de/hCkG15GwUBKH9GH7
VlYoDQS1y8oNJp0kxBD3OvX5VVcPGuiGZWniDXq9inEUtmyb9StWmIVko2VzMbN8MBRHt6yQv/2j
TeAmTJ0pc4KtcsgZcLn/UTRlc6ch/d0X5NQIcgqbCuG1zxLQaqoD8lkLUJYQBKXQpRzhG/ArBfky
TtiPOzgTS0Zyc2+iRwsXNB8N+HTVSPRd0SRm8bQlxwMgkGS3mxDSFfHZFEEE9zl4WJR5eKhqiE80
ahCcNzkyYrz2QK4TVsH6d2rUqPENrKZqh3XXoDTephQEe4fdFhIrNs1dCfMm6BoY5hpRwgrusWw5
MOJWGpi4g2aorgm2Ni0LxspH7ENI8f1LjOI2GnpTL+N3dMAgX115ROifi2myWef+cDy+4PZfyVXA
AYsXZJWw02SzlfTgYLa4agg+nUMqssoLmCTsc0vdYDJqPejoE0QO0NKg9zXXY0l2vr3r8kflIRi9
Q4c0d55cgTg4FfjTZ/dQht9xJP5zVg3nvRmuNop76fPbRTsr8sXU0h8FagajQ/wZa+1L33cnpxRI
ywuJtlhQUd1j7MDt4ODai2uajzRfo44CHYue5oCI624ZLGkOgutAUJvPwYgNZ3nJGOyrZ+Cu9su2
BH53SKBogtb3zXgj1/yTrHH7uvH2mgVYLjZwLKCHMWQk94MgWbzb/qbrKlZHa++Fqwcj1X2u/02a
B3/UmYkwzVL+gjucv6HUj+bF9qyRVg19ZWoDEeEIbpeylelNiUykNBNKyfCKh6A8AqijqPoLykQZ
x5fsyTiq2S+cDqJKkRPjeujH/LNsJJz8ABjM2JQpqMYKIcFsNy2MOEi1qcP/+0DzgcquOEiHzehz
UrcbcleTIARiLd05y71Y5ipOA9BMaZv9BPL7cSo3ifr4w12LxHaJRUdlgpDGt7KqVMDyvg8legDj
bFlKlIx/rp9YDjovtqAEIUG+NED1N1JW/3mxhw+PmEbyeLaDXp7gUz1iE0N0+51y5GY2hacIWoWh
Wv/Yk7cyAJc5vlbk6ESSTl04EyY5oQEvjtMDm4J7LgHRz5339GrjxoME6COmYkmiawZ9LF28SZ4S
PIl4DGi7cuGQ+UCp6eqmsnudMiJHzUoGU79GObwxDVXUMl1R+QO8O4DGPtexEVgPURZJjtAnpns3
JnimUal7m6vD4+LC7CPYUZrkfqXgQZdfIYJqyB1ZY4TlSCtycxkgUgV+PljSzKiiT6AFlD46fsR9
UyaMf1r+Kxup3Kea4Jhd1FvaLoD/lqm/ks1iHSCJ1EOweQEPW1VM9LiftV4QaEOFmy1as26psWwD
8w2sGSN0PGfY/w2jT9gLZ0GIdwkVFlRZcKrQc9lzf6XrT34i7kd75/EFSwVXYvkdOEsf6Uzsy1Mh
kAHQqqDuS97/NfWraefde48T3DVBSFYB16BlcBohpyxuPsA4qJcBgifhAMlaIvM8PwzAu4y/v+WT
Snq794GlSO7xuWRpquKiQVMkLxnIx0957inkl9sa8vWOcXPyuP0lW2giVAKN2IHrC6/8pCSVauk5
+T5SKaofiuxTTXO9a72n9F/HhcNKRSrgwVCCDPX9r6t2QFVoDq4mm3nycIaayy+LD7xVpvauYtKm
RA2kYr0hDF6naUq7Qucq7GaHLsK0kz9riIgJ3Hkgx+SwS7ElNfDl4vnpgb7fiBqq4Icx+wee7/M8
3/82bZlFthpZr/mSmAEk5NH1RhvWAmBJPFG4FxM8OgJn9BCdtkkkIQ7nXCB3wN5RIdX3tvNuQx2i
BXUyvVfQNE4LHj2hSn3PuJDa9/Dwvl7aoLna+llhLgbSkqkCG6AWXWiO7sqz4oNvqRNVxM9I5R/w
QVEskhkLBrtpLWXVCdJnoqNN+tf19V7R0hGsSPy/4ALz7qmyo75oQXEdKziL6GA6XCFGthTGC9Ac
751NxtKc7Vk59zTUzWtLwwdRAtQR8O2auSOSq+FseNVXaGUKRBkW2d54ObGpQaGlwiraUcrbgbuz
9dP7mJY2rgcHDCbmxxVNtfMioJrBBb+wE8SsB3fIApldR6xg61ZSwMjB+p/OjdtAsIGLBLUNl1WC
r0G4CMXfEfb2SUkKlF6hxCpHLgWQ8fzHD/hTgAjuqUmC1y5K3xyHSvZ0ObDRwYIkbXQ2IqSVN4+r
hUr2UjyTn+76mjUcycs6j6nGukIBAetRImqcnhbCumWTA8uNj/w6ruN9KNqFKSa98S7R8m4wSLuH
qX442+3d7PZUrX3ov9+W6/o8amSlwH3hdVQ7ndwxlRwz3PmWMNHkNqxfwPhodt7d5H9NzX3Znf1r
1GhiQRzMf8w9PCKPMdDsAEWvYi0W6SuxgZlf2ujjrvH+QF3FMNn0Lf6i6hCiIuLCyhwbi16/jDyS
CTF6gCnuVR6xNS1Uttms4HSFhuVtYUij3hMLHDML/giMj1qVUIdAh4ZX5ygrJbCuSPF3DozoZkRo
y/ltlrORDQoS1Lv4ZpCsJLkj4wWqsY1Gc6rPnS/0skj/K29W6vLZuyNgby+LHn2H1pRa7gNS+bWA
iAHgaN4JIpRz2PqDDuG0anIy1IXNn8J5Sy7NbJuevgivxn7LgGlDtT5J5UQ6Po0HNGUZFKig0Lzc
6V25XLY61J1KtjKqmkZNTBI8Td7fAjwXJJFZAZosRXYeEIZnzA3hREdxErW8LLrP0M8EHtoBzgz8
bnp+e/VNUYhx25ENkMeEdEoPbh6oedvDVU+mhXSI9/76drazuGPjeEhu9/UM2IlYEfox2JCVZk9Y
EXzeLoyOcDBVKwbn3HdwNFQgLxu+LXNq1W3E645qmH06m1N584b7+Tbe3Gfk2d4ZFG5WkBThiNg1
HpmNEIKS70EH1BrxhSMCUmWTigRzR3DGFLP0USmfbDPVgapjUk1tbtpAni7+KSuECvY3O0HNxb+u
PvWGgExEz/KkPFNnVbqlAil0q9rLONpmoAKHhdkoMrK1MJ+kc5Qp/QUMqVxDBBUMEx0kfIQahuyM
ZE5MY6SOrdclnXcIN6klNwCsGuk+okXctL+qrIdDashFYGXOjCl6nDZigAxSv/sgkSJJ7XWWEDpe
gIeEX0nezQ5fiU7xKvflmwXs4pp/CZWUNoiKjzmGvOlThUqLvN2qo3t95zw8efEhY2zLiXYt0F7V
HpkfR+X9TFowMz33MyuW4Qqfk1Zcdru0HS9ccFpYxpw8P46DrWWR0Gn8pyAmRyoKkwvwGgfQHlmf
NmLAchBGNjD1/nCbN7rw4a5RXjYSvoTgtvof/+BSGvCiUTi4NjzNyk3gOSs6H04H/1mj3PShy85J
YrXeAN5YE6hlUAOS9K1hBvfYEGXcAHLzIc+dBLlgRfeuw2dzQZ/vv2gI2jUeLwgkqtiq+VtO0P2h
YJIaJE5WedjLQV4LYbhUi3HiUrlTM7+GEwv6uFoMR4I25hf+OvXV06kbHpZbT8QR0jvvcRy0GHj2
vA43mnYA+/HiNpifJQniBzngpXdCmzxC+tQ/8JKgPZSjriYPCGSauKtEUPCVh51zUfiBiW9d7CeN
YZtOAVQoktwYfX4qy3flSKCPs4JyoqPU4FaDjOE+WC6t12ggrJl8EuEGKNX2fJuqcRDLzEXjQDST
m+U01xLZPTovXyo7gG3cPHfdEVEcv7d5qQ3OAULozwodSfw2OfsOioa0vNT9hMZb4RCIpfIDk+0B
4LL++9OGM7iTJI6b9w466+wXCO8LN6w8Wz6PxXb4nxycbu8XeOcPzewOGatlH06YpEqei1d7+fug
gwCznm1wH8kjZYMIHabuLNooaQiZHfcyDzJQD0Dp1i0e4DZRoBcH3hk21t2XRtqjW5qQ05Vr5rue
cMLGkv26wAXs3TSwphsMNyBIc4ejpJnfRxnQQphDDrl9E8qcc548kzt1yLMa+fIcJcbgySHI6b/e
kVJ8O3iH1tSR2YSMbN6dAikKwLqRMB9ItkowB7xNCF7UPLWYFpcWdzBpNYHCp58nVa8C1zZX023c
52IPrScswdKLlK2+sAN2avlhu31v5QyJmB7+zG30Rz57Yu4m0VuhMFtnq+aWEefWJ0EdxbjJ1Jqc
nFYnTEc07XspT9vjiijHK9DzolP0hSZOyjgiYtTH8o+BA/Afsvso3dAQGkCZRjqZGYJGsehTN/Wp
WcaeOTB1YJHPmP4oVl+hgQnruSWzhK1slM9E+v5bKvyb5zBg9m8U75LmH2J6BjX7hP/iv8nTN2km
j8yvbvFbHUkPAh0+3wFpTdRuueS56cZ7VYaz8JArlxwJ6dPTh0O5HQGKSua3CKanahOX7snaKNQe
yzVx0uizcdQP7MKNciPcgse7WYvuZL0MPqlsoSDNbwQaLkvW4Y/+ZVm/IYPizRoycHkicKICACcE
Lz9ZldbI4DwnEMBh0AomTvDKW4/8IItfddPA/4T5KC+QM8ZOTyYjmKuL0UHdwnN1PCVNZDzUbnsm
S7AJ+XpUaEjt4zm7QNCE2vke2QyJDEtKaYdtYDPt+eDxqz2sXDyWmCBIyUPG9VTEY31+oW/07iM9
fW+dwtwUFYkxQaImF5XZWDqLiCk4CpjMreyEB/zgOrGN1fCMKxoxb/HjpYkigcWGlaWfGmesPcq+
Vh5cl0aKIoSkQndLX187zBYgZNVu66c1p8+GP5tjxy7EnuPDvaSa25yBJfygF5BxU1Dzmxo2ndrK
CUqjGLt/tKjcbD4SrHqP3jWEh5rRHeas3Ru4iXfd/hu1e56oNt6ypzKRnuRYbfQuhlKxLwbS4ct2
SA74xkoaZxwh2kcALH+PCbEVUfRLTsduIymbhYNfciOELrxG7n9L6Ye5xAdFMKLr20pFlTBudTeB
XkwM4Z0qHrh2w4YcpMGBHzmI7Z8SqRhtDtqpBcvxrjmE+HWpVsNPY4Yx5nQv7Oi5Dic64ZwQ7IN2
+pIUik5q6y9j/g9s/5h4fb5pOmlPpH/X8bi4E3DicEiIau0nLOfHt14t7CfczNcZnG5jym16qCYd
dS6sm/KkPSHAKfSMybTrFOZM35ZLLlkAFmrA4iDPr1Oa0l6PS+SWToCUvMOALjCAt3yt2XlZeMng
75aO36S7Zc+HBpJrfj2xYPIuhTZYo1IAdnHrwFLYbBGdBdDZHdY0laDN9GJnSb/jSOYVmgk7LMf+
3muKZOxbj+F+dmsTsA6eqkhLPrizGT0/gWD+/gkCo4VEFiTQ2l5q7V55Bb6qZweeFLtBO08/m6Bg
hD5izIyf79MEJLRd/wnkzp0yk+j53mZDimY2VWTty9Z2JB1+YyuQhHsjximYwQSXUE10nIxXSfiQ
pb6mk5q2+P0r1Ts5emFWyywkcsPkgezwuCo9HrhX2Oq63ZsbYB7Sulz8rLd+M2V94dEAf9d9Sy6y
YfWgnKWXiC5CgQD/m68wgfsftpd6B9klBNg4ITCsWT/vYhmogGjPi74A9h6D5kMu0RLb2Xoxm61j
dK4hNW7TP/Bwa8KLHlpTg6gzO4kbldjn4Fj9AEHaRzfD0n7lgl+Qyki9y9xHBxZS5rJrlsmePznK
EpohkVk02OVqIrmPlBaiOyODOzZZ1szqbqgBDStWF+zWmrPn34BjKXabyexq41rlUfaqKDap5Tls
BMw9PmJYz+DuikFoss9sE+84FVumY9BsKGwFU926MIhk27qTeb8Z97V+WUAKHGiu94sfsLtYYXbi
FYoVe9Ja2vhGHaaFZBVYATtdXe7p5OpR188EDspX6ZZAGiRTKVyFhlqOKIlh1V8kX1xbZZTGqqY0
tYSHMrLZMeCG1UAmMK0olSBajF5p+7j6RAH+aJIMIZefbqjqNO3Zb4PkPwkdUC6g8uAQ3gko6Y0u
zLeVN19hj+ObKuqz0/5gk3JU82Fl70rsA71XgN5plI/QrwfmuKGCxETd0OEcfo9egbE+qJFWkPxN
5YrHwQ8fjl90d7EM+5acxzxUSrWKLyVIsLv80HkyJjdm/5kZvywHl8XwYuyiefFkupzRc2TH4OAO
xkazKJF2zf6ghXTTeisfzTyiVfi1LatQMURTJ4lWMiAxE7tGi04sbR1a+VUWYFu8WD1o/4GEpx1N
k6zBYZdnb4x+cUzAqmjUpUFGtJ1xEgZymaf+5Qg8L9BrkoNk6xqrXCVzHMNqPkH0sAgl/dZz+w3e
9RPGt+P9W3Shbe421e9HFGwtyHHr69cwhsGzocpwWLvFS/4LzLUwmTvwunVnsWldarEvajwffvc8
M9ixhT/Hv9SRPVmDMVd0Lv21lh++LATWh89cCMr9rgdeyFiYOfSBPKT0gmq1hJL6vpCHKpRoCqu6
NEkb96Uyf+iZBGthmbwbau7XESU0kvX7J7C9P5YN5XOKYXq1+2MHIRA2mEVHbA/EtHMER9Qzmvcm
YYyiW1QBOLPbTSvFCb5Zdu/3/jrmLOahnRhf64fo1Bab6gAtbLFDIZygvliqdSU7EypZ7XKJbleY
3ZKLB1QZaJg6zs3Mayuw3zq0XCT6nWo7gHINTRvb5d/XP872p1o1Sgb9FfBxkn8NowOk/XXDevf6
beth4D1DlAr3v5pC696XtpEzNuxDPYWhpHnOpYgp/OUjezXqRB3cVRCAlhPSRoKcmU9tgvK7eT5M
x4yG+5BQfDEyyL4I38Fq5t/Eq0hceUONX0NZgtDZhPR9uoMRMkMl7r1SdBn9WlUKcAm+zTyWS+A3
WWulyglTYQ8LAWLjXLSfs83YNaFCzrAQ98B2/dl0lm+4J2YR8EayiExzhOMmAVhGLFpOQBgVBLox
w6C3qd6epcHAEsJq4heSxuO+vNyEfNDgfTWZcEpMo98usvuFzqTOS9JSyk0pvQ6FdAJMzkes8gu9
3biSiZpmebdP4ZE70a8PqoiLgm91x7dltG7GiuTAC29Odo2dAs9vvnTsbKS0p3TuN4m5QTtpGCbG
+VixvdfbxyeePakN/IJkkpfQvtaVpWh/RvjvQECGZPotHjvLoAar8qLipGnUcwgpbWF4oR6+oOcu
xhUq23Gl+gmKLLID6XXU2ImNfReuYtG/PklEqWrHkuMmE+mbhIAEfOZahPtCSs6PsZn5D8vQFJmw
+X6TWM8RKvh25s+8rcRnqhyRB9FhW6s6GzTOuc9jwDW3b3ZV8J9JWmcZazg5i8B2cIvYzv2admcF
bBogsEYzWrlGruiAADh68U9UxVQlbatrGd7Ra0mCACugyqdQXB3dWlnCsb43OB/e+e9sTwgEVHlq
kuVmHgFl9htpBo+msYTEc51iZ2wzm7WDt7JsW8w4C/8wQbGykVX462VqDgZ3TSYO9JQy/5vf9c5g
dO8GCYhrkBEHwjDL7Z12piLooQp0Yf490uPe3f5Sma5je43xRcbvphal7l5bIxRCzgbvUQ8rKO/v
jbECEZPbcQ3H6KlCXwkPYc7EMoT+MipooLrLFfzG41Sve8NRLpGygqfSFIAsm5oKSGGOdUoGTOuJ
hrrP1AhIiX3bN88VM/aerTYSs1oR0lt08ZsfnBFUqf/Ns9MCb3lWga8NGLyOrqPpByyh+ZuBMX2F
2ZdkS4MvAGRyvyBymT6B4LNkeX4/8iAUbvZcIu7/cpKWmpRDIWmFQYVkO1+g35CK1OJbeF/Q2JUV
w4PSD6o/LxfRp8gj3Iv+RIqsMmG+TdD0vjsErwZsUukGTWz4fzVcOroK5/1lVaCa+9WkPwI9bLx+
gUnr8JJiXYsvPrJip7XHj9+5EmBCkrwuXqeywBsIJrp9OchV8pr+0Zvh1a5IP+8jx7slkcvo3NuL
0Cs8YjhSUax10pYpcBbmYH9+MBsHtxF+TFKiZS9wodjJpKQml+BWXVNdJvI4MhU5IKtkhMV9uCYs
4glHa2rj1M9Y0GQYzl8CBJC1ps/ZNUpCs9fgdJIqyjjeyQ9yOlTxu5aeshetegpqO38/2Vns+Os9
ZJTyJ3bnMqjh3bEp1yOL0pgY6NhvSGLKthkr6WWZ/2b4hhuDKSTfTdDPA2MkqQkvPHTYaEsNnj7U
b353Z9dI0VIcBs28SPIEQKGnvw3psHRmKRNaKMFkmi8v/eNrNYl+KTj2wkRSSXUNLZykvDJRXvqD
4S8Mx5DFQ4lOVZf8mcgcSYgO1NWMKRHkVpkVx7ckDbXVVFfL+rloODbZfW0SLgvtFCh2GBlBIgw1
dISLXipcMEainIbFr0raI18posCAho1KWcmnmAquJTh/7iekU7zDUFbdT/Gt8JfC2aKEDX61JvyV
ECng0U+Dy6+Zj6TYLSQNW97xADSj8TGh/TzeIez5Qx+3O1QAwTUEcksZpz8JTv3OZ+jv8SlncEJE
D1QOfcWIjL6sTL8Y2wjayb+9tHYnwLdWoy+HIdRkNmPm4CFAF5nN11J3Q9WdM3YZIT0wYDmUIVSD
GBMjJFyGHdGbzhXx37vfNhSWSep0hU4LOtwejNyEGZHOHVrIQX60UYi5S+6ERwOPlb47KhtANn2r
cCOVwZq8WNg5rNzkN7vv2OwJX3BWnbWsvmJySk0ZdHxvs2GsHtBl3WGK02ZBJqb50GqHfVomsxKe
Mee/7cYP095Dc9rQmM3XEKBuGNTTZ6cOiSABnOBxXNSBSkAIl6UnjSFY+SxAwNLo5vsTVb3NuibW
r7Fhp4n0AcEh+yWGr11r6TGpWXoMwj7tOxsj7+Gq0by+ovM5oF/G/K+sZVgl+a1kknFKEV4Un08A
778PXVG2HTDROGaHEA1cZDlhp2gTUTBIZkPTh8e+TT/6H4lnfU9Pv713HOg/t888SVyYWI1Ux2lc
51huqXZJOuLQtUHTlotaomIgaXFpQKSQiiU4a5lBhmhZELiDLZszd6xr29oByzln3dW3rwMgpdW1
aREjzCDMq1Fsz3sQUgzLxK+4xhnwW3xq4t+ho5DLV6lDKU5okxSG9qCv8xV1t2AqM4vwPbMA1Ac2
T0JogLxnQCj9jpO3u88CcOahAUok2NEgybZlA/DyUw+eKbQMIq7g95Um0BkUHT0Kt/ZAOmQm1+jW
Nq/gYO81sWsM0V7+79T8n0LBXniXru4MROK2NLf9xBZdGlQSBEnpghARDdetx8kiyQAUfOv9sp7m
ZBuXrSynq+6Bbg0G0vFhT/JtUmFsbj0panxRMQemZZqeL2D/PEBii9miaOKykxTZoo23xpR9R7xN
EGrr1oc6QhXmVoQD/0wZCCJBpfuyEdD3wRWdSsG5CYLIN0CsW5/QZn19qo2lPKRW5WFjSBlutNLz
xrRJGSiyqe33VRALDG+Jl4Aqp3Xrme+LJo69mn39aDvmEM1YmT6OXqbIe5YFjvYLxnuIRrQAsPt3
4eZUEMUmb4TF11N2Y5/N/HnwACU5vsgFCAXM7wFfP0TQwxNMaP16+YsonkKJyuxruGUtbEgUwtMu
7spgCIjQIwgyDpcT4SxmVo68KVMz1y6q11Li5U9IWXcRLLe6GpRwFRTqcCj/rOiS9v250+PlJ03N
1wCA69xwAb5x3AY2M0xdPY6cZz4XOayju27Gg4FeflAKXWtTKh3s+1ycRXHMF5Ipi5GHUmtFiSag
zDkZqMz1zq+Xk8QAWFmEEEdiSrMVBDETeedQi0LTniVPw/r6Xinljsfd8gNyrMIgKKSPRwabW+XJ
UW9xwKdKAYaTbBmw59UUyobQ0VdPUGKCN4iUHl9MWwaNu5DGMct2MDSt0jAqj7poYO6LTTC0haV0
nEiCvxr0zmj+D02Iu5XIG/oCgdM3mUIgbwLGKKHFOM4Ce7nUrDNN6kRzci/vnM17YcBwXyfKfei1
AW2pXt78i7xqHCqLU6HdxrMk3m5z2bt67VBP20IUa1TWuXE9OL9uvg7IQC5DjiXw0KsHaGzoE034
R+yJAVWeSmT7TctL2PKxQL5f8ozl60tPFYpFx0UFHK2M+iqRU9aa50O+kwOkLv81ZD5RdU9wdN1W
Ifhbr8xLkLmhcKfkCAILEKeRIzrPylzkdIZNciTx1x0PJgqPFUK9SKU8h6SJSP++sMDS/6UCuLkO
uwZztcY/LZJGIij4EU0MxvhLUuSyoVRiDzxS7KH+L0nWc8UJWZfJznEO9jPCeVs+iEBRIERar/6/
d9yqkDTqMGKQ8nEDg3vxdJ705bWEoiRUbG3q/21e/W8dXLnRUFfG3ZD1eq3prHRaFS9crh+HyGjY
zlMJQ2fgjzl87yRUj5tzRu1QCH9stSnq6rKlS96dfPsLH0Vb3yj6Y+I/wPRK2sXxFW+rw5Ev+2Bv
3iB0xSQ2Bb6r2UcuusmWoSfcknTi7cYAMz4+DiV1xXksJZAHvHh+XlZfRRzjLXS1OVM9BamruXHR
QnccQa3n1SWpb7bc7hdh94HPoAXt1RU7INy8JCrGOxnKJco3L1/jMTUtlFWVmM5rsN5tqSCnbGYt
U93ACkzxw30S6tdocrqDEqygpaCgiZRZBcOZWja08trzdGZB0jqDhlxK/bxQmAPWyQsmUoUKb8d9
BWRpVdkisiUtDJIXQqUNKV3l23/+3FWirPUmWBX6MCxygGCkiSXgKqSwmnC6HcMqN7wvgkTQo0r8
o04dDaBAf3NqtJN1Y4BhA21065CduEGoyD3ceCs11++sVKVlNhDIHRAn0ePFg5TTJALeJ+XIlpYQ
oWWJG62UIZzR6QtK30wqC56VKoihlIYlbWPRwJb4L5q1ujX/c7bbg+BwB38UcEqUxotUi80HNOlc
aoP55BDxkEUBZDswjwW5Bqtg2j8waBMSyWHxrqR2XuWwxVfGJYFxaCvqFboK+53qVHE22+6dcsBu
LPdigWkL0ig1mpMbULNY/qKkY18Kbtmo3mjFOxPyCSySOVDtFZWPnisBEYHRsjd/831Jwl3rJA5n
2I057KIDDMwPJBII6hgAwhqCZ1r0cPp4NQgAPcKa5pVo7YG13UCSQi0XRck4W1BpsjPR5O8dS9df
FlhBXFFIrNYLOemY3wyi+xUfFRMyHCRI+U1RmXMYQIIPCp/AY4cmUi69Pa/3qnX/jU3u5wU0vrfB
66KP+nIPn9mxPPWK8jwK326DAdc9k+2nYkawCHou0dWCn1dlCgt+zZnBAME8wYTa2OhTeaHtzpQ9
mBO1NZ7VI8vrVDw1fIkY1x1rwzoHL/KBVeAJJL0kgzqjWzEVyt3r0e+gXScK8gqyoSxrJ+yqwZmU
morBnelb3eVrBph25AVY4/sebI8GQqdigqQqOcSBNGPyVtXV2lCJDLP4eQ3oJ5EQohW+Gj6IbcfK
tCWBnj9jGJ/5FlUlf+r5QeikhLjIGHv9fUUX1J1xhwiJc/2+IHGtr5dZf5ZlsO+7rTTT5sCaVl09
rLIVThxmN7cKN+gyAnOMdYIojGsrjcjST1y6GJqrRDCxCJjaxB+upkFS1ZL3x3WNcHHBiLdd+Qfq
9O7DuR1CByTf+tqILSZjJvmpOo8rSXZxbkslVuUedOE/SQEPaliQEYc6OawrItC8P2BGgM6nmPk/
TyRFSEtfB1nQOXICbgohohmtrsWhDLZ7Ijr8SPfgcp9nyrwrRluCThYVJKCwFjp4qqFL1OXGfd85
+vDZj17yE4GULJQ4g/bVXoXg+oRvcUWbN+u4NWHxFG9EeaNjWLiJqCZGjBcVRcvGF4+dY61gSd/s
fzqnP+gjnEC9u9FQpOV79wVyZ4xjp1ugH8KIw095X56ko9AVva33j9DgtuGCAOk9KlFFKmOX00Nq
8GdOFHyF2Z6SfZ2JTgUeN8RUZa33iwMNjAcvSZHMqtd+nCb6/T/+28KcgN9FCi9Jt0+lgdXNQTgy
SJv89lJw4xUALGQZ8XM3PP3dKRnodfTE3Uy1c+Rvnnckhf1KTOWkDikslGto4K+Qhrd2s3GY5Lk4
xCmKeB+0wlj4Dm0Q2HTHnrj7PCFlWbRilQJOzydqCb6bfxxYXj9uu64mKj6m5gEUE65odbG8RwfP
vMjnbHoodAC6q/OI0+ZBkCVkm1uB/evglAn6XNpfQAb0664mVMUXmUYE25149C6j6484VT12X+Bo
/+Ya0L+6AbQw9rSJwj0lsup436kd8OyN0XJXu5GWkN0aRi+t9BJZenfy91zmW+OKYPsM/OsORqbg
dAiK/0qGiokm7o/178zjZngwMqUcT3SqqaRRa86qdDAs60l1cGp7yatxiO6v0KHekzNg8F+sP6TC
HUVZJt3A+vyj6AJMeYqiPjbe5Dc1tHd3Czb6jXfbBGWaaMFWRTDG9sg4tvHFoCztmNpVPU9TSrHJ
uRgSOe22pBZk8O5WcQfAw0v343uKj+K5+wHZIxTHGQOynC/Mj0z9dXs2zwJdtfEjAdx5ZPPKGLNh
Iv1XKFqA97FZOlrbk1fRm0IKpS4g9sK2i7cx7szqTxg1jFzg3M+YLLvy1DwpApKjqB44hc15g25s
7P7TN4mht8iS9oh1ypaaaLKfdkQiMFAGrz6hyxiRMexwvyiG+rX1axycyKYx5GFdQWXOmepL1qR3
C+sDFn+4l0b8w89HXTxW3iXx6MNTN06lvTkePTfoilZvOdUhn7D3NxSFips7QHYCr72acarfFOgb
dIcTiuzMiQIZH23oyonZrL7yQur9UIKCc6lskIi35VR/E2VrxxZL5DFQAFH9tNwGt8bFWYl+W3c0
l6Inrj6ciGOxWFk80vf3h9p2ZnBC9gnOU2CxD0GK84LLd856537Zx1D59+MlJH1v47sdLPPsJdrh
HeO9DlcNsk/ePxqOo65ft1IEsodfVnfeAAG2y2ApoB2+r7V6XBRWfTnilMHZ5t1LBbMHgfxL8HQw
sSMd/3N0l2iX0jr5WXRB9mWh5aYUufJQKocEQVJHh0JNLdXXeiv9RLkhx1sq231oUGN78Bl8m/bA
MTyYv62B4lIRTUbZiprbJD5dT/9MpF+yJ7W384cWc+V8/GLnKeOIkP1uPkzvKexBFkEyBJPib4Xw
N0KJLp/3UFqSRh1UE8euQ5t/0pDeR8v71VGNW1QH1RiKJ/mcrSmQawvo9b99vu2zjxJsp5DCQmL0
k5AbEFEacxKyMOXYAEZyr1YHk/2GfjWCimR6y+cpu+cPpv3cj/Rm+TZAZoL9A/VvZQs+20IuYHdG
K/F5Qain4YtXa1amsNWkv28Y8yh8WHgrVieKpKmTylC93m+DryIkzlDPSs/p4J+Ym1vyyOH/kzz7
pHa0A7oqz9WV3J03+WZ5IV2y9WNgN0LgGOQkCxdlNrZ0+IKd5hrkoLj0myZzE8HfHrjCnuVtvoj5
ACoKgRGwReL8+w96FPq2AHzR/nGfq7/1ADvW1EqGMv3A3NPQkMjkUUDcsPu3iwV82w/glXwiPXXr
mY6MJ7MN6cHtEBVz8VD7QGQzHo+LkB11luKPG6/T850a88GC/+RIpzUCkHvbNcQkMJoIZ3Qr5IbL
ObXolgTpF9pJDofc9QPWFT5zOfZsEvXEeL9Z6nUk2VYRQO0T9nJpZ0j0PwKl3k2+eufm/PXO5Tc+
gE3b3fzqyRoMIZi33WI+F69xiu8/U+jhYDvw70hEIQ0uYviDNA0gv/9cItfnNvDS6d1Sr8sDv8sO
RBlNvpoAbSVqKbBUtTI45ahG+PRQKmbBnax/mkbEOjAsOK903d3x7QXqVU0jo/jqJvOc6Ki+2f3g
RFceOr6+8pelKvPTjpblokkkiG4yXuQbcx3q1eO7ls2Y2v+r0dtwB/NjLjjJJfB9FUFDLQs1BqH6
17ozxKmjl3lfs2pCAqCpmi6faV2UsMr0btCNA349sxgtse/S0PhSuWEy+EUSdNwfHMjTAixmov0f
E37N7OlMvAi1LXKDb33BXglUIbRHR11oOGsWpIeQiP4M0Pifz3jJTLynAnPsC/ok2LtGbAP+dtjI
cDdpNzLAIah/dPJydMcURN7ehwGyn/vVy7z1XjOn1nDxK+J3mNk7NAdiAvXWKJym79kW3z2DCtpl
yQT2cwDAqXSfscUhSA7kBWrUBtNSxfaO8WsszhJHBDkHussQumuAJ+nkVQGFEkMcqEPVOuix3JzI
iGo9NYpnA3xJGePXKcLwKQCT5G7x9LcCn06O9V7lTjeGNvHpWH2KWpehiiu7EFyfZOFw0gmQnYFh
PwDXNtZjl7tSPOwdJlE2Sa4sz3M+EwIVms0NDwH49soSxdjyWxJf27FAcrZDSUKy6Ef1BqH75t1p
I8cwQ7qqGLzA4MwD+PxZa4bLZAEhIxVM1lcbYKox5iMPrpMrK0UYr7ZZUDP1LQ5Sfmj8WxKJ28th
smKJYZ25rzUNB3+TWsCUUK6OafXKy282HO5tBobi6re6L0ptDggZe8ppnfQI6E8sQjr1K0SoGgqc
vEf02X++uYjkymrJWDk5Btl3pgw7wG6gZgUjqrk6oaHldQ/ymdlsxp3wDdSsCWkMLRHX2yE2v1lw
fbda2nt9oGEAxgtCyGx1UX4N9ecyVopsZZsNps2v0xsUvEb9dKqRM+L6zg7u9a3bwZxdkHN17WeA
IUfIP/WA2BWgExMePBKt6j8nrfMXzh0cQ6Yq8W9maCCxI6dpzgdu+jUe57j+yIpSMb080GrZpNDT
2rc4VVzsJQvuXNlc01IweLOIrX9zcIE9l4x4Htq85ujuCWDogt3MvymjfkL939HYeMCkmEvQFNmc
3fjxQZm8eGqnjAYCQXhkg+Gj+GYQcvxtGhcCaWU0sBs/XcN9WhltL72pu+eOcmvEdiC5pTnFR7rt
onLOUOpu+K87byLGQZfCuK8mczf3dcE6bs/duPOVhBKBMbjNh1kazbF68j/uGfgdIDyHqwoXnoM0
iZSF5+7OsTp9jwsV3DlJ8y+BAqo28C4Wtq6aoGmBIktdyUsnvu/1Nc4g+oqeYQZ+aBHw5C6tLTpH
vPnHbMbIqAkIJG8kZ3vX1pyT+snh4BQcyQ/HeLYrjvqUCV4x3NwhS/CmIRMkIm6TkAC+FX8tC2o/
1xwVLFvATc/zvmx9miZU9ObVCA95NyZu/bqoDRvlQHnpnnKOKqUMyD+mqhhZPSrlwQs62ThUEpa3
U2AzAENURNgAor/di90yNOmNvXbu+R+TdPNGBCMtJnEBNylGE1BVb07jPgGT9fyyJf/r6ggw8W+9
OHcEJng/qOwi6mAgr4h6NAhwup0Fj67U+9+hSTaC8/MAwVtsQMq3Nar0uuze1w07jrV1iCPPWDah
l6AgRhMS5mPAh4PDup+p1OYtL2zw9XdCB29V/WQ9b72xl/rvHZ/57dILez829I7imKgStsIcEFcC
KJghbgE/1/fBt8yEI9tJle3eoxcFRLKI4HCHQw1GEv+AHnvMQaKL7gEjE/hBcjzV9fPHE4sSrKUQ
c+cBAXXEdgR7NKDHy0OWMkYrQufs8xig2otdmhghQASRaMwsP68rl1URv2SK+50E72Ao6fcVW6Lf
2NSEyl0ui/R56CQJ3uJDaW2fXu6Qkyr6Mv5og6x+8qORDb2F0HQcenhuYq9/AAomaArFNK0z/nlx
WMWCZ7yCstchyeIaaf7NCe04Ycu3Nf708Uhgeco1f7DywmHZ8+gKSB6xxCcR95sty56vT2t+gpKZ
RbGYA7rSpeg+hHIvUT9/m1Xwz1KVHrIRWGTmuvpclFlW/ns6aEJaNPyV5ZD1qANGIOxTIGzzvqKd
SLerRCvRugM/0JVdAIOX4cr35kH2RhutU95j2GInsE3b2n6TeeFdTDba2OaeiXyb0sdXSNwOu9T9
hfAGCq94CAWYnWbuoAcpuyNKB9sjusa/q0m3RELxY/X5w2Jl1mtt3roDHkSTRtOBR6dsyhnnxaEX
uRRwnZJ4ray/Jcwgpm4aR3Z2z/B6bF4ItZvz34MNvNjkUpCOYGh0mV/vYkhI9St7LrTHNQ3kAfpR
kO6U5B54oLkVSNGL7tIXpcOmvcO2lhwNCybcd1AZnZZy1xf06t/gyc9HfOE+6gnSMuVGTBHrsNBN
auptk/N4a/vKGHx/FxH8sRFmnhpeP6mmKBJt23eTB1YyRDtnCGH0cFpEt/WiQNnt2iaZhBS8zhXT
JhDESkQB2sj9KFf6iUWHtGnctAq2BnJhMBQ7kGVv4W6eTp3ZiEZIDTM3DieFj2X0EiiPxwgzua/M
LM09eow1tndpF8sR1nUoCmHINN+bAndaJPr7eV/07Z/6kf91cuiTxd3wlT1mT3fT0H6edsQtW4lM
Mgfqab7PVrKQfh6t3SS5A2Ber1/u2zkDHBwGilu1VZoZDmgJVCKSTQ0dngH+BqH5WLA5faYX0AiC
T7jyWjMoAXjjNRXQHjOChZdDIONj7wzBd0AcfaNzmS+omQRmd/ycwQyUZ0ccKvV1OJ46IxY2Pxpk
IPV3U88EKkp9i3y7VuW6cDSLX3YAsxyq+Ne9IWo9Y1YnCEUpoAbTjBjoyg6aQ2nTnahQeNaPm53o
V5ONyLLlMchOpvqpaBGLfM3m1JS7o1jN6Ikyl1w+XvF+9XZXU9rd/qHR7/sDj/g8hGu74zRq8VYR
ZkkTsyU/wa+uxug9wtDD3dX4VaRGxClsMIeHtqXoAXCOQogOxobfYLMTQUdtTME70LsAVHfL+mpw
aGsni09ecpFcaPQDd0XuV8yTnVIy19P0NF27rLNTDEOt8WqMzlUb0T11DJh10OsSzgOQtgGo5+Og
FrIknmz55a4yANcAKX1IbwMRJlDBm7ed1/EUzcDhQVavNK7RN7MwoqXgbxW1iaER734oW7/xwRCE
HZLl6OWoZYPWvGzmF5QS1Qw9IoZBqoDtJJ94GKmNBAYP1AZPwX46O6KO2SWjm6Mh+5Viu9yO7V+O
c7Hw9Uf8kYg7V8db8UFxexzyeSoAH+KpRkqliSDvHvfomrCElbYZd4X5l9/Y8T5VjcJ7YkccgrKe
828gjnUeNdcULKRJb3BkRKpHKD+dEM0I3oxOdmVh/DIfYYL2MRR9qrFQXzym7xMPveYXlg2Qdcwf
4beAzwD7wls5pe7XGT/Hxw+7mmUu40AEgguV2IvBCDkmgAoYy2co0t0LeJ04OCOTnpoTjMepAEHK
AK/pnxlfmL6t/1ucoU17gYJuecB5YEqhYVGyTGDqCevoF5J8rSDSV7f4VuF3c6A2JowTiXTSLnmS
8uPahRApOUT0Cuf1kVdciQ7NjSwCMgknR/ws9ntYmz6FrMANPzUq2cQZY2+Fs7Z/6J9C06nfvNWS
Wxd2uCiLWiQmTM2ydtwQDLD4HKA3H8CyHoqS4O5beE8tW3wPY0nlVYcfgj7BRc23/LkntnL3yKhw
0svekFsmisecvxLLR2Zj2X61Uw9EAdSh6WEYUDGG5hoC9Y9Q687im0zAqMHhUhPy188O5ICLEL/q
5xihC688tfDyMhELEEKv4Etq04Fax1nfkjE3obrRRJSxWuzVLNUSiwu7bxgsVxKxQu1D66QYgO+4
y5sAiUXRXmSWjpyVvABLmQcm4Hayo+dQkk+xL3TpoplJ95js1PmJfP+PPWpy8P6z7Ey39zDT3UD7
x9ww3oRiwgsevWH+C+KtasQjiwl8M6rv+BUY9C5KSKfgG4w8YQe+5zaENZ0DGz3r4weIN15cbfCo
w/efXltpFNitZG45f4e70tkYJXe+sl2FBlLRvVMn+E+og6ZedJY9mMxn2R/ZcX2L+/jfp0kvGyUn
gDHgd0dY2oykPzXEu6dgUkfuzruljL02B0O7niW77U8/fLNRcAfEX7jYt99FxXMMsxGppv3SGVnd
mYYGn1IgvALgdn38gw9oYwAtAa4tyBroCNct2slS2Hjfa87RZNS5FSJ+S0dka2oBP7t8itlGZwXf
nEWvxKMqBjEmDxUxAKxNVkVdEMX7+UgtOBBA4NE1cuGQGFr/WO68gsHsskVk8rIyBhPVSrjoyVYz
+WK+kHO3qQUUKotO1gcs6uQkYcgJctZqlJxeXrYTpMoS1eljDgbcYfKyFsEZ/l6hdbj+f0dJV4AE
YMExx2d75GRZCK16LnUyPTDJyl1bV3oEeH7zY4I559mAamKUDheHwfmKvtMRMA3lR1I00akWkILN
CXUSx1fY+seVB4toR0lyxidJ8kss7viV3q2jiuj2zeQhMWr1UOBSZU5wy/9ky1dFzOsMgT+GSkba
2sT4gT7vtqEWy4RgpoVapRLl1CqF++uHoB7XogzSTiD9BULc3f5oQFbdBou/Rx+jQmDNOTK2ipoj
5ceqts566KV3veeH5X9CepcnxHgGqEH0wsuZiOD5AtTJfnWdjQMusjOuicdWs8DJIXmVLiKog/au
vmEmSGIQ/WnYpFsugN5bKHLGg1RL7FYeXY/b0FLcA5hQY4HW/4RNJpbKwCkNWPGcBAD5532SEVkc
fpTsCVdOfIeOEi9yZURNkk9MzXC3dPppTTjgw9zdfKPKtJp0qyhlCF8FFa2j2T8kKCxXpXhya3r7
HfG8KyLO2vq8w9ijNqcSI55+NY387tPjz5F8va35IznTrwTvMbQUMfwMp3f/OXIOYUXSMZZzfSad
70Rzjn7YWj42b5N5kYgTlWEX2NXz3Q9NJIXbQspJTvDEqEj6jwHXVZeRFVc4lwder5wHx2s8Wa0F
M+yV2Bdg1CGAe7MGl4gQvt7aySyaVH4/1e2viVa5opE6rcxLxOxPPvjclVIu8T0+QIkxMjS9uxmQ
Eeth0NQ72L5c78wNCTeM2qgH+1uA0r2NtlnA+EdhyrBrDAAqaCcpqxMp7FoX6X9MqIKPI1pt4Kka
6nr/UmzNBMFZJ0JthyppAKzSVW7ePrsyA7ABbcl2JJBo0haSYFTvrDUEj1x1RGfyiQgiyX9Lmhyk
alPrz/p6wHAgJoaYCj7tdAGKzdEWKSHyaTi3AbOCejFkXmIoKXrCX4vJ6QahCLIjl0/4Kop640Nd
sXFSH/vRLyRf8fGmlvfPgoYm9QhNsuUXaDjuhKbaAsPbRjT70BWxrt4h7uH78RUzSe+aNdu2Q3OU
znMWplfcd1M6eqki01IKGGIWB61D9WnhupHviUjuw/mTSfZEG2R/LkWIJTslkiPUvF36G7yoiVg+
FGTVXrCntexN7I+JhcTl3gJZKsp/2h8aJckc5mq5N8Jip429PfzFoxlGmISi7kRwSNDa8rmk30AE
76OH3rQmHOp+IdpSvelX0qRdk17v8Ot39mM3cfCkUuG21n5c1NoKoQDXi+xmqRJKi0/Y4y8nF4Zj
Hj6Gss/WwBqfBgPUEipJyoqhUz/VW8RkzlP4MIlLH6YgsVgxn2zTYMVNPfr377GQdmffDLeCsyqD
HwdRB2fnRYxy/DJMcthZqcZRqCvP5B2eAUtW/Z4ykeuH/P31kWGQZVHRNdbxfoTkfxzgjr9TAKpn
DtJ/jzIMUoBxrwG4eKXn25AIcIRQOtM9l6kkscPuQS0XmsB4p8TPM7Lsw/quc1yJe17h5QrIEFrC
g/MW/I8dI81vvc3QksHTnZgLhcVLj2X0TRSpB1KLp5pMB1XhynmkvJ+rMHS/+RFFx7BuRmpzYl4Y
rUuho+EdJAd8eauO4GaFTyCNnd+/yFr5U7Ggs3/gieE2ZSA7CG/Ifp7PkYykr+9I3QJWWrz+wRcD
D4RRv+nQY/ITH2JhXOvta79FiosIaRQoqE7BvCynsotiGMfiiOqntu8vjrOPZbw4/0UsY0qgBFVY
ZqRZaVqNPnfDAK0VDv5nHQx+xNUplqInIYmDw806/BtpyqeTwZ8AJSU3M3fupgycZ1CRXki6THU3
eu+Q+FVJu5T/IQIFEZedCUkwvvl5bfp1CxzT4rTzgTSePJV4B/P+WKiw7LMg6Q7eOsT2IO/Mrj6e
d+cBHyqMYExJF5hAWj8xxMoDQYxEKI0EDSjBGWVNp/AaDBmZGPs5PdCi+DCqJVL4BqZbRD6dnbOf
DYcgvvAQ4aQHUDtVdKsfbjOML1XqzZET+zFbY+n3vzPIOJSv2V6nF/U6YEXhL7h/VlvKpI7eKs/Y
B6ssUJ3fL6A80mWzgadIOyPIU9vKRuM2xTIKJKfcDM6Ivri4b8wSPApjnvCubSowps2nNaqrMnZi
CpUyQ6fvNdaNDsQcE5PeX/llzIfJ+WjuP0RW+uESdj+r5DWJxYCiNB+npx5D3IjR8MeWCk2xvxUG
U5Br3dLQ7Ur0nKp/Ah9auMcvPW8czVHf2JB58NUxfJSKr9xgZFk2lQcRYdtxbN+wgrceBDrE1sOM
bfyKcEXekH9pGpIdeVZKoGsG2QFntu28hzERR4roiWJzeY9B+ZhJIAYg/XgOFmtQ8OtZIRzjrz9e
7VDCiqOryUMJP1DICS/33sbbzLgcj0+5vjyOxgFxLhqYKkl0UW5llkeFCdUTjHiKIr73jIYgtlmW
io6nj8mKzOw9hNIAlVepHMjcfpFqX+RbABOP6+mF+ywHZKl7YlHFFSZkrUmDCCGPYYojGdVkqfJl
ZmiuKaNk+emEq3LaPM3gryi7qX1lUXK8axG1/495CuSiqsryEcECPQs2I6xS16XhSpgVCgWJehJc
Rna8k+ZrOkdTR0VdZseGYN+GTwsmPseodxZlg7IBH/r8Lhg0O007GzKSWMhCZDEBqc+DtQYqtxMa
JfjzsaaQ1eY1lmfMiBPzyyy1+WFd2ENvK2MRryV9nZE08Nb6PRby5JK7GbRSeKlloEXTAjiNV8zk
HGxOScTc9sD1BhMNez1DuFkH8BA0JgmZ5GXk3gNoQVKklb8eTqvSxwmNXWATsNCBUHvgYD8MftNi
KtDSTeyUwNS/2cdupEJv96vFMfhUDo0CVaJVEVgCmYMkWvU32gJARVj/SWh1qu43EDioawoKEemo
Yjfvi9h0/fU0NQrbbXDeEAMP3MJtlnxnjvrqTOxYCb191alv+MT5LZzWPUBZtyv0HGINzseyi1Bx
lTFrRHgVJsDnERlYwm1gmugIF2YOQ5GC3m43zPrxReD8nP4rGUS+xnKiHGoxrMp/eSkfZVusTI3H
otMoSIR+L6a0eyPscU9Cnzfilgzm5eebIbJ/4h84Q2rMj0nhvMv9pYBT4hk0dR5ICCIsO59nfwhX
lXdvC1janojvhXcq7Crr8sBG6Voz9sERPR5lLxdUjNRPmedIByYAlc2H56LCou64owufuCtKCBFL
dlCZ6eiDbNsK4RxJravTsvWdgas4H/Toeu5OdznWbfIi3OxPqOvYv18hQ6p3BMiNdEMe8mAlrOE2
gezXKY8onLZY8oUb6BSAlXS+sYPqpiaUwa+1uxbGXco2EuKVsPsdUct2G0FG/xUwlDK+rxY3edK8
CIT/vSKfVWL9kT27NBHqjIbTjg8UQ5qEya1Tmt5KQTOqK0Bm+es/wGFUAnLXsKhZ0FfgUrA9h3bx
ZeMuO9NbI7FUrMKcJK5qJ/Ee7oMcQGg5svS+uKJ9m/3Z1YjfJ9pocVa2U/JczvRBTkvl4xzcA56v
DNxyWKR/p9BlCg5geuElcOZWnO9qe+a+Nvt7qtFmJ4kWDr4S7K+DYoSurzocKk4qkOws7oAeEvtR
fA10mR6AP4LW9ppjVcCglO7dAsHhToikidsmgLQ5ndICh3f+H/B6j3cZvGCYbVpsCA62dPh1NtGa
L8ZotAQEVQN1mb49kqmNQAwp6G662pZlkN/3xUSPn2N687bkruM8Qpstq9leh0IzMEB5G4ZCTDJM
0pCRrsAfcVt54mFNTvQwj5JYA3qAibfqqfRXiQiHjD05yxEdY4NuyncdUo70r3A3saitoNRImI/n
59tyvl1MH7f+MsfgFaAHzHJKeBHl3GLjmuHEONuj4fqjhfQ9lrAcM0YIWmIrAAVrTnrNW1S9rNe7
/JhNStqT9NRk46evoBtuCRdMhGhjyYc4AwhYLOLtLYQ/wirR3Oa5iMgZZTXESMpL6uyf3E4UXl2b
HYp2Q3EIkEjfzao7B82T36Go752jfQ76lS/wp+EmjJ15XAI8tB7rOqLPWSs4TtjmKDmGLfOll9hX
CPTJx7p/43Lid4pKInBjlNjE6TdpYjiuuFiRe1yFo/j0BHTaCRusnXNyM5NgOO/lZLatr8PCqYnx
L3z+gRzaO2tc98Q6CcnGDJtUgDrVfytU//yW15Rp/hIo35uUOQrc2tTzZ2NeT9QX03GSMqZB+f4+
XsNmMNNatzn+5T0W8vfzHjbGRGlMzXybVBUT7K061+K1fPegrjXU0IrLgo//Js59LiyQSZwAsUwG
wp0MMT3P0kxbFetVAdUBpYfF5B2bcnBTfzA90DEuLMFSOkqY4V66E2UERN9CNaXdtPxd76HKXW0q
JeO5jL8PNsm3IJA2zQjErMaVDngr5AjZ0tdw2Pbx3E6kEQ1/jC6CcFy4/f2Yjc3pPbUl9AYlnR7g
NNriVB3GHpgdbTQfaiv7Ug2c/N+qm+Qx2i2KH8vMCnq30GuCjTfBDF5z4Cpt9mWkKd6XhCri8YFS
DLBiR9Z5J0N8sYSGHeK2tZV0LeGCRjFmckNU2HJIsqUppyQkmRlR0/uT1rvJ/nrxbyNcZiAlix6j
vFr73F7HxJPk/iPfrE5/uy2QjwsfD5jGT26sH5u1hNkSVWZ3M+Cznm221YWc5Ko9doFTHqXjM9MK
E1FbddQQ6U8Mcz8hAd5pWo2ZgSuj0CsYvXFl4XfB2af/uEgCqomtusREutDiwQfhaZk2ShEHbo+i
lZSBpr4Lva78k+aiBcYz+5+Mi4tFjPWaurVRZGF6ZTPZ2QtCJ1VMuwJcZEj6wdK+4BbeLoc8edwD
kxc92ZlwUZb8Kue8AomhdAtPaqdNTBcupaLIxQR7PkOjZn3GCq3ZbuV3PXRC6kdszAKYwtRJc1hH
YRHHkpGWLM1DYu+0DNSvxsQGcPL0rNvBKkRME/NISXgqdtjcvAQtJULnZXsJeSAy+siOSOUxjkAz
l30sJZTkaa9qYGRFpePIXIohI3gYf7uzD6K4vbopXDQupBVWLdyEO6oDL2iB6idQPNeu0vH7m3Bs
F3HDGSAK+RjnkcorXep69ZmXVXZYqgEf20nkAAtEeuiKL+ExLwgJdXjaGUSzLl2ycKdqxr4XlKVt
lO9mD6Je48gY9W6EM/pRTAGXJSv1dfKiq+RUgjdwtgWfFxIOwJsPqsiK5Xdem2LjksrQ9+bDOw7G
DVWSJRVkeRTIwwZl9c5ZQ7KhkAzPEm2sMaZYkAB4vDZ5CvWkKo+UXGl6zeRN2VS9eXRwaXjqr60E
QliGGBmSJlhcGcBcGEFHuXhhRnhMiV5SjrKcdqzCtuhKte+nuWul9TN7Amf1Vh0YBMQOuDcdNYRH
OqfgwJs/FQdH2s5XSKk4v/zNBRVlgp8tvws5SX6Nx6YJjzfjUiSftj80FUU7phdKcT/CNiEPERvy
LMk1a3g904X//RgSN7Nn7jpUC6GLj7NBv3BhqP2YA7lTKxoINUbh6NMLJoPgXhzngcnF+j7mpfIj
wo8VK7+tMwrjZcefdwkGaefEmViLCQ+o2gMOqEPq979umS6jQeHcfyN611/RVjGq0XIUhCjitEDY
1S70Lp0PZnPfmLN0AtGeJa37La837cFUZPk0NDOOrX5mhGEUOYfIsim7/EIOX+eAPG6t/6ecDqOK
cJlxbBN0ajLwBaYBOWbIL5aqu4igfsosS3zQ+kIAX54uu9cNBa7aCCxDbC4ebqFi8NGuI7bIt9vE
yhDg4HMFPbEE/eUu8pnpahscZAx5Y1LZDqKfMK+aVHo2uuEiWgSrlnsligYV+DOI5Uq0z4fK12yA
6L18fX1xSp7dN/WLmo9mdWsQViFVNOTBD+TtZ95litePq7MvcoCq+gUaYLLTXP0DtksI01cgrgss
WNrk7n5lQzc++WXMT5WlCN5BkWJrvlt2nEgrZcYN9EGqQqZvrbgK8g3aWyUwKbnLMVDkuAoUmPwW
KKbyft//765+vFhQto+U0/vnMGeLmz3GO4oQNax5n4CyG+tMS9nhrV4LA3XGLQjVyEDj5VYeeOAW
TMZ/CuEJnhfPiQzBeAnA5D3BcFCbtnbQtd6Oqb3wyxV3iV5H34AzDthygFrSqCh8t1hUqwabFGcG
0kbQ3j9uAvhQLSFvKv9Ja2MSNTSm57gwZG86ky0A2hM26jcBVdnk5aKiMTy4cFPs0n5LTd515Nya
ujff5UW595xJno52NzkSy/W5QuUjf9Yib4hdIGp9WAHnDHkeO2Zks5Rf4A527+9LZkL/srhzJlaZ
LVSHbN9sim8WeSJIkdojUjT9sonVA/W8JyoqecKCy32x8VLuaSwE05WRV3ktrTAAwKRyUQKzjxSG
fPmaj8ku98oihJ4ty/d7sHRDm+w3ji1gNUwKNMW9BBDGKXxHZp/wsqaa49uIiytzit7jrIPS4CDP
Zi1r2edvL+ePsXoc7YutOiPljqgeTENrb+Z1nRx9R9j/TWkcXufSNVIqNLSsKUsQHF0ioyDR/2ty
qQnkV/H3p/noM0LbGKJWVQQErodYNqeC1VTUmmvyF/YjyawNxMqm/Iw8kIy3/QvmPkfCqmQ6Jg9O
HRJR7v0GZWXNtncA90AYMEyqrI7FQqwJ1N8BZE+tNS2w8YqdmrX2qCDu6l2mjp6pNrCTSDTpcnKu
6HKksOF1wUPy2kvdtOQ8snqUtOK33I36VYNHToS8IpsYGDIbjGO+1tJod5vlcJi7lKBD3xZdQoct
iJxlewtLXFfkT6CVFpql4OYfG6PljdVimAUKCR0vXKWw/nCq1oJXd9BkuFdB2Ifl7Rxb+hYTrgsl
uvZor1Ry7t20EuE80Ew9dHuNIaVOPeENBy8D2MvO0MZSl/KK6pVAkkNAPdiwf0aIaz5ecJocBsEL
PE9yRfHIW+KPZJpVl/gn2ygnKBzqkEMj2ASzM13RNWUi5B585DkmhXkJ293AJvqkAkowAPaW/rLT
IKw3U3OTVYTgTNBNUnSWknP84gGLVXHDLPLUt5pL08rLJSY2CEbcy3v6LWsGCkaOMIsbhHWzvgZc
keFVich+eH9k4Hyb8sp3qZBKHA9oZ1wAYSrF3QNjLcFb8wJqi3SiE0zxHLOkqMeUNiUoHqcCPaXt
XbbXxzaFwvrLqnK9to54HlKdFN1my3+THsJzpRtIMFAyaNpS4P1F8I0GZ9dcl4+XODHn8ZuX2vZy
7MC9UJBSdPpsBGXI3fN6luqxL6wilS0zeMrTXYIAkOzNlvIG5v7tJr5I82IPSVa3jK6pIwc5CBFh
8mAyA0UEsfbIWM+8OF0Aza3eU/U8E8RuZy6wJbxtRQdTwuokyFcoZ1ZPWr58dvvvwsuLcGhrILam
QnuGKHeyApqwBsNEmw3PuOJQUifG2UCeMS8aeNCe+ZVWhub1jJp5l6L/redMpbXjrp5PiOMAaFfc
xDUCQFPqCL5/uciMimJMXvlcbhxnulgPisTPJrBlcqFLShfEpTG3blJP1zFNZxIrGuCwtoD2GlZA
J0qRjKPgEEO+pEiCPjipKIHVMk757Di+N1vvZdW9jrSUvVmkupr26vgka44PCUVXVLHKTeBdBJV2
ip6fLkcjE/v0hGm9ykgWPGe/Z5ZplrH/oRgs11o/lcovzrj/e7GrWl0od/pv6bNfHI8ObROgtHZY
45il1YSZA4r5fX48kFi7+ZtvY4ASYpK1T6DrCEdB5VnQ/t6cP83UToXBCtJ6c9tQ9S9NirEk2dqk
KyVafngc2YiLLHiroeWPwpQLH39Gq6F4B8evCDfsGNFynB1hQUAS/7oXBzUNTgFUtP2nC+N6H3sV
Ncfm7T2w9SBL/nuUZJY+GfSDI3kE97ZllIQUXOtODMtwo1Bm3v3ld3iSOCDCP+LA96rb3XgDFaWJ
dmEUPOuNKTWe+7wv1whE0Wo9ellum55xV8h9He/38O2tHTTmAhl+PxTukxRlOnUgqs6QMJCQLkot
sisYCVcbDrpSW7bVT/UZWHw77yqdzQ/aT33IShA8YmWxAGB3iR58OlGmB0O+/NybC5lQpqSRn11M
JR7NtWK8Cmko1ij3xT7uuaTtXSAA77o+H4ARev4bdpAmgYsG/c8f9kIeY8B3xflgf8jxF5mPWff0
oR3JMm5zvFuUqCzyJbPZ/5+B+7RHJ1SouhjRX1QCzy9DsyiyNp/eOVPCYvmfkqdXyyoIGdXONZhZ
BbdHc9qMva8R+Rc+RPdVAzw8lVfeKcK5ZNjHfU8aoP1IGKH2Yc+8eZt6T8Db1aU0XLOtukNXbDI4
JRI/OxrKk1bZJ04RyCchUxXxhJE7eFS1AgJj5UVwcfHjVzJ4vY9Qc38yaTWid6efp3BQVbPagNb7
HxSYBDTvEsYE70f9dgPaH9opE4nzQqgH4LWrtr/r9KZSAk3j8Fxkt8VyqdAp+Sc4ZSrXA+oVF8d0
zY91l5cVuD+vXhXCX+5rUB1ktgnt2k1Wb60Q+7/Y184jp6BtL/+cCHcci4SLQPHRcgWXw+dwImG6
0YqVPYy6u+XHcF1F/yxa/MkkIFgLaZ+Wd2DRTYDqFwjt4rKaQbz3QOM064HSsGSOskXzutDovq10
5pf0ixgSMavx+w1s4N3W4eaqqNinD3d1iQQl6i5sMn0nnBiIrkp8U6IV4NSnM49PDjWLNyUVdMh0
0s9MFN4cd61UcwUgt5lFDBYePPGBuhrH8EVIFfwC/k0BHi+v78QwoBhFdQAsypCiQ3I5WVoGqnqr
D6YvlZrTPMpGMw8rVBFD5XzihYbfue1pkmwqxUFrduwuM7Fh5UwKYFNAd7jnMgEhATTlIpodpykA
0rIi4ik2kqrCdQWVKgG+IrAaV7Ap419576hf8/inoLIkkJ/XpCk24/4UnSeUgVwFqdkHD5XsY/AR
hY1wxj7m/kAeJr9G3mna1edt5d/cZvKLH18hTwWoV1VtB/s/ZI6uvVrP8KIeiU7gjay1Ooeg8Qi4
Daf9MhJnDgDKm8NJTJZECm0VH/mbtE5ZIJSa4t2KKrDwmPWRiIQEvLDFSpgVAZoRQVmc+a5+RdXE
AJ0QDUBh7n43eAOTU44rTXgjyM/lTjvaIIgeaVxbEHSZI93BCNQrbSSljoSrThyDv62zOKVhSpZW
XaohhpTu3oCjGZEMRhjyeDTYGGck9neJnLqKvl530D52QDsmRwz0bKTixFe3tcPL/Ze5qZUPVw2E
6y0Oie7e1EfZ4ioi5TuKLTdnRTK/F+EEQ2OmSJM3Hk14jWgXei4FB42biiI+KlYrhquOe0sYsjQC
o28evgCvjZw47y9S1eF6e3m0z64wt6AmrWt/2QA1wUfH6rZCNQu62dinW2NdSJSpuIo1uppl3Oi/
P6u8nBo4i6m/vmr1ke0ccxKlYl3CfKqjhYmI7NiqkauL08fCbjFFersNNbxtvuoJcDrmQGy1jzub
SS92m/x5w0Mr1eRG/IOzNZfWYhWxdQLChyWELzQHPe5m5VPfoG2Zapcr8ESya1BRD+u/JhajI+Ha
ibU2aR40h1ikULsfOv8Fp5GR98tBQUt3jbcuIJR8QZq8H1ZYmF7SMcyfHoanud9vzRTC/sPm7G70
ilMrci171npKHHn8vdhTmX1Nl21CAIMNqkLlWTK70POnoEAb8BGePtQscUs+UdXtcK1DEYvuWhPl
do/mhhiZToJHJFYP6raspv657+4DHhXrP0s9eS+FGAvBQrEQA2U4Q2dvrgLiAYaQOir77eIJAXbx
J0w3wCAwU1Svxx/bJJTFdsQ3ylwkNJKBCLF6DWklUoJRYarazQjWh4w94CKJGHvWL/myi5nod8qu
BxkYLH08t/tSVin6/EXOAADGzT55lnIPgNWpnaValdrVECJdZ4oaM8VRSW1j0XhVvbYc2Zl0K0Mq
y06UvpLJzWniNLc/jVWcJwSqiP5FVVbQkRe3teEZNJoBI+1VXTkg9qf9tMQI4YAHqvZeGp0/WaMu
4xH3Xy5lC4Vw5N4AaS7sQU11J6kHySCOEegZ36k1aVFK1Qz7mfteHXZGzdZA7AV0gtw3cS8fG0YU
7dDvK6onhiGBqbVi0CJhBQq8y5dFWi2FSWxKjMQCkhphrYRZFkX45+L+kKqdK3NYv099wCSeibFO
1kvORvzDR+dy5LIxRNq8JNUBCTwoeku1J3qQguMqYfBMz/W/hBmfq3+CT8InO1t9CckICeLWeN95
rB52PK8Dgm3XN/mYjuHMKpBq/8CRxamGvVJIXj1VXYq0S0kIwglQETtzuZ9gDTXsZD8X9rwdgtdQ
at7UvwllGusNFga0qdRl7sGAUveB3pX2a7jo+rW0XIOag0nSG8XJZ8z4mx7TZMXohroOT6gwJrd+
gAUCTEa1/h7ElPAKTLPSENhXwnkd3tyjUSscOf1PnzbbDo6r8GxjeUB1yqEvhE2g/BEU9wwuY71F
H57gQnrLYtUz535dIb4qMDlvnk2cCq8092RR3SmSqsZSt8FbnYa0HvtAjqZ6qBblhgszx7kzJACD
Dtl5CXcrYALB1P1pOt29hQhNbsqZSkg/IYOyo56NYyEVhg6jrpAtsVGK9MsVxOer1TL6udK19xiK
LLYyhCPAHUiUBgpBSz45+sZFY8ciJ/WIzqgc6EOSPSOB7KhcOOJciRLAdmK4WvXIz9DAPRPpTFP/
cDO8e7ad4CfN1ag6KF/ZZ21H7atopT+TD1gzUMCAmVw7JHy6QGFtV/siyateAL57SV7rO9+hUGn9
eTPLFYatC734ARAI0pXMfDERp+7yY93vCIvwMdhSNhXT/gRp/q0bDkp1gpF7+MsTOo1fL9dF9FMV
U1Cp0EhJAHreK0CiqE/Dx+x+SrlGgo2maWOxN38Lh6Mx2+ZxFV9nTHOAhP+zBn3PIg9sHp8rKj9h
zDdyCfBitQL5zD/fbvgGcAH8XbtrtmYjvZNaTCynVX+j+cG2+5cZ8quOEVt9kO5f6r6UUGLTo2gb
hdZ7bXibsZo3B77l+MgxcB2VjCzqOLnjpfyhyzQI0VRTR5uwGV9n95XMaKlkbSn3Pp4r0TIm07Hy
fhVpKe3H1Oj6c780BLUkvsdtMcwW+itFZrWpFzN6dLlpQJh2BZZ/DStst5Pjsyo6e3GFVFIkV8Cp
VOYdkTBwDRPUdlq/ESYqx+O7t7m8iUlFe5rDuJkTcvTj5fXVwKMJ4gz4oIa3dCna0O3KQU8ATunR
9zrwhTXGzEAIpG3caytFmP2gPK+h5yR/dVKDOqr+0LqDdtfNn6kMkCngKgiex7xUHDCMqkFhkzM6
sui+RBEPesLn+Eai16TJsA4M8V0QdjJLkczmD3FYHAtOK7dL9CowQU4I65q887Ejl6P+0Sqxbirr
v5nCuhs8cXtnomuLev6+1SxPJAvjZDn03Y1yCeCZ0O/M6o0/8d1JGoN/LqcfZ997NyDloof8TBXS
vTkmbuth8g2cM7m5x6nO+2cSGamREov1GNfAcnViuqz2b0xClY/GQHW9PMzEwAQdxvRdVeBrDog0
8L0TevtKewlClLsQv1BgUpG4+5VsSDgKXnssMh4UI1yl3FYcRxj0zmHQXIq0qStrwHq3o5OYDG9b
UnpoeYj8IprNzAJg11F/0lHpr0k/jczWhmf34/1XrppgQgJ+HDEFkdBhoH430sMUNKELQhwyjA8W
B5dCimoH/fcgb558UevD30P30TqRJqCTuKccWxB0TNrs/KO+8qCrwOq57jJ7S2srwG+FI7F00VAP
AQAGfKA6ywP/x22XUPJwfGwBZwWElx+JANKYMs/RoL4FmthTmLGa1Kv3k5aQUcxf8Q3FqWEPGKkP
eckJzkBZGr6KN0Jvlw2oGFg0xG1z9bPQv70KpIO+qy6Lmb2cz7BBnqK1UMdrzgk91feGyQHc4mBt
/7Dp1w0yPx1ArcPNRw4r9GVTB1yH6jEN8sBo0SuydZAkeQrLwq94GPKppHSIjwH0REElZehy09LD
/ZbZCcMZNd9UjxnHI145j3p7teEJrxq6Vqp7RpvGyW4B8OdKxTRSzvXQS87omCHI3inWI69GzcGp
7LWMwc/Bh2mcqfOGwvevbOg0qcjJdzurNdPQt08J2PpGxGKLqsIf3o7r39G7Pna6CsCAn6/44uAN
CDTiJ9yHw25q8Ig7G24zAxmtwoje2Mb+ddk1nnOcg6En8HD1jmumpuSgknx6iDevvX54jT7K0+wS
3GQLHtCxvFhxORDiHk4CyOGWQhYpr3EaXNFik9lPB2JnywJcVxmrjRVUVkMH6Tzz3C1kkrXpfhOD
iIB2jC+55aQAQO/1WR5kUTXIl/RzW120o7PRffP3eObnBGmGpftjY86WiBz18jwGnVRi3qmdsg+9
LdGW0P/bRQ4uiIoAdMtGR7HD3Weh5uV8OKTREncjeZ4m5fMrh9KPL56NLGfUSAT3I5C5bFbQ9FoU
MLI7lzQdYd1VXulsP77kD7j1O5yE1566iIlCK0X/jTFGoTArDfc7E3y48r7PRqcdtvzT1REGB65r
eEu/Xt+Uu/RcKLIu8W6zo6gHHS3i44JFHUEJWKNA7nTJP0iLFce7pr/VHEAHoeNg8tymkwh+nQj0
1qwzFzcMgw/udviJ/dcWzwsLz2jAGME1QhbyTq/BZb+xW9F/uE8D9juenn6UwQ9Ucw6g3VyvlK7t
95P9XsWJqi7mTDAwvrxNOIOrwAronauIvIYdMvcKfoQ3bgI4uerPXz/CPln+mgkPa479Kv0AFcIt
h4TRU6dM8MA9yDUzWvZy0dAWQaAjNHiuGETUEL7P82E3ButHDCkciexHR6XmJen3CxO5/l0UO+b6
gxt87rwluVNImcn1noDmTgPwaNPqZWWhzbVDJCICHDMl0sCpqza2+A1wuXVQz3N09hx2loVUOPJg
ZTPB492jGrs9jJmHWnYSIh6FcxaIVMSZy8Mt/saN/4cQ/LWQhdSieItDYBC47y2xa1jHT7HU+NEN
ZllMunHLTP5Zz8aPmw9oUH3q1htuzxKbWysIuBS0uEPMTdQ+GQDHVvPJN8i+I03JP8Q/EZs3muRe
OTIMzpOCERIncAY6fRgiAmu/5QqbbEMZLNlfOTESzqyB9qbEZrBAxm0lv6g+EZa9z+gPth+X427e
RoFRO98d7fk7Fpo1c0PK348PhffLKLu55rD51yLqRmY47B4KKligUBjMz/bc7lVxhZ8emAbHiaqw
/H05VERdnCjcayNplBmDYb6qfXEX6xWBYdsBZfmYSDV2gia3Anqa/pq9ayoX0YP5pxeSx9gakrOv
6oa0GnK/uJGIomTLPPaCGhd0Qn9WyNbahXFrOLULkJ6lUBGOcvjfKcuQomBrJb/wajl4Ah7iWeOG
d4nEYbfPmA3gGHCGA2tGBUJ67WDhZ1cvw4iYqN3HIybIm/hcIvDhnliZF8ZQcp/SwDGTxODIohBy
xIv0SLB+iiKWrxAieQVJKoExoyAzlDoxsIqud9OcvXsjivhGsblASpr7SgBWPA+rD0BJjhEWSl6K
oxaz2wOlIhhzFQHRIG9Oqm+GlbouffDJq+YI9Icnf11CszpmfrfDsUNeBX3zuHhSRfGdu6/jNsuM
oJ7uEZWlNNCJBxZbvpTlEYCxBhCeet3vQRtQVbll1FjnfRM1GvIlCtTxOuwbaRVSTi96mErmpebu
PxXZGRPqQZ7RTWtZBF1CZI02CW85soJwL3lPjr0+KOeFw9CjYiW1nf9E+x37E566kjoAm+LETn69
DkkWhOI+RtYqOMeFIIftMVz0WpGy3uHvj5cwBE/copf2MbW8pnsPrR/jtQ7xyjAxE3UPEDx8mGFk
RNoswl9X3qfxyrzUDOzOdCO0Asur+tbekyK852a/T0EEzDoeWw9M0VTzzySfppL2FrLt0d5cfTox
7Ar8Nnd/eZlYvNkafX41OGP6Z7NGf1nUEZ3QdSM5g6bJcaOW9wlXow4piUrFuPTkmY1w11SbIwG8
19+t2Dh33a9ixpspbuSP5ey03nhqAgRjPmHr9UV8T7AcXa4a8ngOaYvv8aS6tuKWIHxhgPKaIpsM
LB/54N7MLaKjVBjoiHl8JzDPr4Jzamv8JcTPelGu3FrdIX3NfM+IaGd1Q15goo618bz/UKPHgGxQ
cweU8lIxzJEb3kQZNWbjPTBMBD95ul8ArHHT0v85RMtk3g2ShwUp85ylI5sPhPYx5j9Ssw6HwYn6
kxXzTPsuaaGyaV1uph7A0e1gJviKzIHwYor8ZJq72QnY3CHK/1llPtA0v/nlhAQMQSjosqtA+6bp
y0cUdLmQXeXn5L/n9N1imKNQ0Q+9/OB4DAlD44mM7OH3fEGyat3wu9XtKAJFXYihV+7Ri5fLwFD9
JAk/F8sabqZEa6BFjnrLBqtkrveCO8y1hn14wT0Gd452J+d3TmWmGqgW2rIu8h+GhFWjqJnb/Dp1
c9VYnV2eo4jFCaEeOl3xaqp3E2Neu3NCMysYCskf8FFp8Xlk/BWcwAxTGOOVRxVKcoubP4KOx/TM
VMZbCod891v4MlsuIZYtPNqdjyvhgUVaWSkW2jJo9M5JqofxYKIieDE0QDpOx2w/UoeMyWN3k+3o
gCHJ9AW1/Eo8tCUh35MZ63OQpK3L6yFm1jlfuzPidlaZyZZ1y1yuj7ZUImQZ3lCo+0Tlcg19Ftpu
X7nFRbzVvcsFkDJ/LynVzt8FQBZLnutC7zLKhtDM57ubwYwYVASGH95fijrU7E4fjp1nxZUhXAVR
gZ/445gPv3+OJ6h+gH3QhUaX6BMJFVGymZcBzxsRXMrhpFwzttmgSxNyvjvu3tHwWQ7n0Jsgn59j
hAWW8lTbQVHnRkiA3zDbZCOD55l6N1s80KxNlVRlMmqGObWgGkm8vG7wVQ5pJAuGWSnfT5Kd7IcV
ScR1OvQ4prxi3TcTHa9f3EoO4bAIYSLKoFhZ71ET/Ja5NxOXDw2OzHEye3HspkZQ9T93JvKiQkk1
AVmX5Pgu6sT+KgTK9+bAHGeSa/H33xZLYpJVj2WyhgHy02jsNJddcs+n1U8EwxEB5J8QipzGHUs2
SXBFY33zysnEkdVkLiqc6oh20CmBLxA0sNdvwyG93kb8kouU/DDGqfZKZ8PB3pmEfdk0AIHNqHKl
WlsSsLNFmTFcdbAgAQQuInQEhDyd5V4ugxlq6QQeHirzRc5mFNUnwaYnQ8Rdh77Vl5g6ogSBgkPO
kpRux7m8ofGrDGlUIglamdpIsL/fuZbl2g52NywJHK/d3O8YTXcwoHvXodmf2l7B/UhA3T0/R5cP
PhOK/ik4FDlkmFVr2hT/VhxGlzMLvJ0phPFgOvWdkk2I4O3OVecqWEda03xL6Z2z9k5TGNqTmmys
P9sw7i87YAIk/6xDfc0utXLDJJcm/KDVNm3qROfUuC6S3DmM0PZ+JXB/FsujFK71dNsfZEU0r9oL
7Lhz8E+JWlJNuW0aqyetztp7SSVBfw3pOWE42d1Zf/iFuMFY+r3zZJPwJKY5v53lYhXYxMQqnUW0
MxuC0TmCv9mRUf71Og1ssWCVNFnF8b4j5UoCoUDJ6LwqLF7hKDqtOQeMhUlAXOxMZgOTHoD5fAMy
DnUenwZ1hj0dnm0a0jnK4I0PaZJp/ZBvZ/0NKcjDzfZ12CDB5G2haKLr4UyUvzaDzSEU/rTBTQQ+
oAQhZQhB8W9FMI0BW5Bf3pQEFhk0HANMTHphCXF6/LbAumZJGDM0cD5mc/TwQZzvXjCdKQn1AG7s
LazTCM83XiZ1KnAznvOj2KlcJQ9ZwaKJqoDdwQxsqBqVcn4X/r9KrOPTr9ahZi8golo6dG8K+RMf
y8NCUS/rqOpUcZZFQHwPGoM5EU3LU8YtXvhQCTFzVqyl06okp1KF6fG6p4F7v35pBfRalYCXFjuw
rGAf2lFKBzHuIvos9Jl6BulVG7Dfam89eDI8oXtG0oOtvwrb7GIQjrKQNPv8CxY+MKXP6l/BphV7
12z8/Csaj5pC1AAIgePKZ0FLi8Id/lg5SW1wMpC2SFMAnHMg84Ei+rldRGqMXl12VqyUv0lDunWh
JBSPR3/72MONBXUYYbgtZSFUIvhWvDnRv5OrHTHDmRkqBXQizqKOPX2Hv79yzuuXvCpRTn2N0oP5
Iey+FG+03e/0p8Wu7fkSGYIwYmdDbHCsMlPiDqKoqk8AiqsEYl1a9oszavA4uU+9khEkxchhIvJs
q5bplMTE8XH7EhoeaOdvIwdxHb+7FCzcD42hvyojlc7PkHGwaPhh14gWAgS93hq5CJQi/Tb8w9De
Ml80WsIvx5usRP+V2GLl3+STcnSBHQEiDVgGtjCwVPE7lcJ2yS9QfxQUKwe3riMqB7WkUkPQ2Dnp
vttmAtB6Pl5xmK+FXubBDVMLLQimCfWIu3sAcXrUCgk7ie2Fy6yN5LAHYpG2IcVzCt366gEcSG+7
9tLvid17DE4/kImWhO4h+nSBDaSe8eJ06vnQmzQOxtLbbXZO6uX8+ppfvFdNp5YUgt70EXDbv0Ug
dXxV0jjTQV6/DhtnNt0tS9l1EES3sgR3pSaMF1s9EDgolER5oY5Admn4cFf8YF8fAKq37Xx322e3
yGxlUmn6kYgaNFnmT5OGfipgrSeLTQEU42dGwrqXazGIMbMe6EyYviUsEAwz8xmRwJ7kfBq0c2xR
OfXaRzaU0oMQuQKQNijsD2xbgh49MgQiyryVh77R6jbHZK/uI68awSF3WDaQgwU7J6aADaPiJc1Z
ZOHq0n0Ecf+NEMwWZ7iawklxnRTnaQRiTAN+IZtSXV0pGOOL1ebPfLXom7X523oFzWlQBLvgr309
2+55ZfwsMqMTZ85P0YlxD6m/HGOq7T9gTBVgb++In6GhXlBfwvIvIKEmr2zcjemzx+nMsdOfB2lV
EHnP+KrltiBpUHXfPLumHZfF+E4CIzV5CHnZiQL9vg/eVILgKOYaQFf3mV8RNX0PF9q70GPeKye2
Z6wEN+BG/5oQgDNy7W3Ztd8S3Y35R1gOF8sP1+ydarhm1RkFBPJHw5UjgyI1+wzY8dZfCPQ3Tx+F
XJXGIYT1WQeyC4NxhhzansISCjmdAKtz9W8ghF3RzYNPV8sI4ydcKRk1pacbJrCXa2DoZvhq9dRd
APeOLYtnED32y7+AOShxksuHVcSZ1K9Qsg1L6th7bG177xQBJedr3y/TFLD63WoGH6gMHVhmHYqY
vCxdh1U1LhlGlA7pJXrTFoXufASgA8gsyED0HpSIzImVjFLgdfq9tU3Lc3jyvjXj3x/wofGGT7eX
SnYnFwaTCRDPhw0go0W38tbXZA8eqmBV7lnbZAW038c8glFO0YXY+78E6Woi3VfKz0CrNnl+u1bM
9Vw5oLVkoiVKURJwLrJELHROi5i1ADsTFk1xO0Uv/qMSOOv5u8ir8tyAfQPwaIQgZbvfUIqk6EeL
JMkwT1RQ7JsOoG3SxlqWEjJHcm+ovjehY2+ICYFU/U2L2kv1aRtd7J/8bTMDjJO27L8rA9GxVNNG
Esea4ijH/t1DS4Y/jZAICczryAdgAFQpgDOUkuHRE1cznnY3rrRmMTBc5KewoxXGlfgsZQB5zZND
bhGy06cEJY6Aws83BYozyc23xdyx4BrXjwbv0ZIRiqzdC/uRvGezqLzHEBruDmRDOh3P0qPZabYc
9AMmFmNqqHMrT0JqxqGjXUsk/Xhv92dQSdr4Vs5v6zTFi4tei8CQIryGkQASDqg6F+MJggcbV8gB
If1iL8y4MAf1egIY4wu80XPwaQ/IDFYRpPIBRfuNHqNgtQWwqCOyckaZ+nsD6ShprUxofGLhJ/r6
GdrViezk5CWt+8vMWQjrOOoZijCme0M1DS3cGJ0ylMRycgh5WWP61rthSLBt2JLswLp+sOH57XRl
dSAUx6BhVjxCNLR0K95FFMj/u6CsP1i6iAG/hsw7yiTSfyz14mzg/gfTa7RylS/bG1RHOSjNoV54
/sB8iRAUZNGEKP0d8T/TG8yxZaAeBuX6fog2JbAJR1EBN5NksWmCKL8PVVmTSwn5MpNrmuaruk+W
NT2Ch/5qcc9Y88NjPQnS7symfwsn5kN5lcoHsBuftetFYYC99gFdZiagOfWRqo+XIWiVzxccfTKM
xJlF5b5ORLEsYdVJe/uhZGn/JHgoCMhvny7yP6qADU3YAI9dHIvPJMRqEn4bgrSj/ZtMHjyGPnjQ
b03wMwHaXjRKK415y3FPKYrwjYjdniV2zW+xddzU806HhFebhl2bUhljAaS/PMm1crp9eJuWYULm
JIpazbVVEyTpzuO7vq04Sm8cDiEcbC230WS42QYbjN7GB0lmLTz1M0hZ9Ekh7SD/TgUTF/YsRACC
+3tl8PJbItO/yfhgUNouMH+heAMY2pX6vCY1CjDViirHtwSAXUdDUCBxkmqNiSHj2yQDDvM/Tzc8
nHN1EUBX3yBPMKfuLBep7kPOwBxHnCgJRcdCyStYhh/4fCnHD0hy0hy6GKFFsZYeQ3VozwFNa04D
s4Ww+o6kSzRt2UdysAeQDy5rTfK25+GVyMGOVrmUhDHmPbOGo/4nQ6/CA8sFPbkwezCGr1y5KMOm
kSAeE46FvpJiioXPrZlmifdJi6QrHI5llxhmDy6HKol2alIHBusjYINyVZSoVpz8e/4jpsJv+auh
ujNBfH40GCY4MXy8OM3qp+drbK31+MCw6oEQph879dqK/CHVVYpNeBOx2SI+U8XkNOYAbIfdkiPD
ECinF2G8ALFszAYruGHLTLU1aE6CBgbN42nAYyLyFjKVzlYg0dDu/n0FatjV4m8oskzCw5/PPjtS
RjSad9CFs8D0IwxpJXwUMz9VtYBXMKbi4JZFlHV0hNo/c3ZAQtMtz1onZExqU42TH6WYsRS01yX2
pPqjvpg6oVIEfpFSWICucFyf2REpwgKORs2KXOkqKYKBQ1kxibrUc1AHvxe35Vr3J6qZ9szbP3V9
cNN9O27N5ddezwtvB9Mq+ay9E0gkzVZBCyS/9+6ZzT0V1ZI3MgxqVay2WjwVtDG0bBUON4v5K4vs
P7n7m3HrU9WgPfMoIPhg7cp8NXOb++GJuVP5tGS/OYfF5uSoK/vYO8s2VJQ7GYMdHQmsDfJhiebo
VhyZikbv6adK02HbnsqULZM+5TlfKKaoBq+4OdUoHMnDF2iD3eNqxYpD5Cmcu5ReWgzGknU+q7fu
cgyYRr3YOfRJZPAGJv6gY1Gfz2qD82DPyh7/15xusL2JYTZi+0Bnj5ve2cvIna6yNjzOJmmo8JVb
xs8DdpugsGXi0yM68GM2+aO3AsL2Cdt40CvxviR1CZc8o8Nqj5oVtvu4ULzk2voVFRtcInI+giD5
elgYVFlPlJaRj9XsdZFM70fOVoISBSdRX9SDJYlzbMtbTykiAbq/vZZ+gxRT2QvuLhTt4qOE8i8t
vNAT+4XM5Rr08K7brsEjqeiD3peaiz2rRGRdArhDgiOV06W+HRbbLNoAf6CFE2DVeMSPygYl1O/F
NsfqYNHLD31+7gDnlyOUqDk51/hhgQf+p/oxUvWVM21U484uNSR+wHL4/D2GQJbX5hhdShibS62r
d0oosLLiYY8TA856tvAauHCeWN1ifP3tVjR0K3tqV1Ltgr0hGFQ9j/Di4TlJIS5vkdCVcghxWAdg
yDhmzWlBE4LNlB/bENzsGBhRkRKXqTZaZ3XYHV/EIHI6EM3wXTWws43WRk6gCzIIvrl2xlBUpffo
S0EyPj4Zu23zgVhySHTxc63yeZDs9k3718S8W7lvp7c0v1g2fLZXGEaKv87On2WgPTuV49x0rvJ8
Q3WZVqsS0suSA7Ipss6XGonbAI+4bUkM8dqcm7e9inLZbBqbtu+ZLr8bemfpk75JeqflcC0GqKZc
QdEYV6g3wI2acowBWtTrz7BrOXxshcesvL9mSxsLkIoeFBVPcauu+ufC+5x7FRk+pRHOAqczDbB/
1zwGTRUbzmyi+0Cbk9/YzdZ0rcwpIWVFjaoikiSUDU2mF4FhndPxzltv0H9/KPqKJ41OsdvFtaxQ
zcgpTsehfQIISwN43W+jaxYzHN/6lyRob0ZtF8jkVlK8xciUDm+CzwUvEwp3Au7sjHC1Ji9JI1Co
WtY8qB1rtF+IwxkngiaMZ/9Tw3y9wC4etf+lkcR3enJKHqA2V90Q5F6rgMadzKiK9kzILhbWOyrG
/0ucGyntpncLxfqkq8lmtzRHzsQeOIQ0zioRv3nKforVgiAY6NjCiXxESRGoNvKBhqpq+AYczNIt
RJNDKztds77gjNNFGBd5ZpYYxGCJ4RFrMr6PZqFsgKmJX5FeHVBaZyje0G/q3pIaN+tXE8t03BcV
CqStj/zWRMD6jTxJvngKYMVLE3RZw0aYQ9jpg8XCjMykS35MaLnuIrH7cSMiLNHVMayHj0hmPF41
Wv0ZqW+tLy4hLwlCRKtQks8cKydkiMwkbXd7lW9wOY/XNRePiJsdYPCL5jgp11A0xXQvXalaS8KD
N2Tvp+KOvQHLTMSLoQgD6/N7iP21Qg30EGOnihbxFk6xMt4AjOsF53WUl/amzuRvgGpGlHKsqvO0
3ByOogpeMg3+9m+1SwRQObkNjky3BhC1WKPa+odl9rK7wwxJkdejQszy366eZrdjw1tolotvH5rW
Dxqo1JjGPaeDducGafS49NBHqDvSsmpnAiDI555GyTkZKp2eJJD6kfV2GnnTqNMtzNxGcKT9TS4P
/eTZiCFizLFcUedY5JKzcyuc5WG4kK0a20OeItIL9Q3Es1HN06TG6PI4vJ7Zs0f3LyqSLbLO+bRp
KGxSUKLJ6AlADpLhH7uuSRadfRrX6/uZ8pE68kHnyyLkleHSHjzz+Y2grh+dBYUJ6tAHTIPBHsC6
uwFsYfBTBywIwvL0en7QtNj9MSIgIioQl6N2BBTZAZNaxjl1IkXTtcbjg16CuhNxh8yfE1qMMaD0
gGpZckA7vB2vtiIiSFXgFucDSCMcLpkcvIJCrvBg3/r2PQqIMCklnvglhhevlr4gSMevgKZIal80
q9ff+gSy7VfswZuvPdTHuMBOhCzaa/MXgHLfZcG/4X0cqT6PchPjiVnUas06RXpV1Cg0wwuyYBM7
NpvVa4hI7gtz94JRcjOzzu14dfnrOnoJuRuqS4ZlhkIa7SVfl9m+3yqdZqdyw1L5AB4lZgyFO6Nv
6Zh73grPFebS6Edx4HB47qzbcMgFmL0AnpCZgbaiA4eEEiubKGVtfrIRaZ6L/RGdE+EEFWRmke2U
5HFBpK8GEVtdALiYSjVr+bLGtwPgREj+BtSEtQktdizmkj7QDZWl1ynRH0MlCnt/GR1jWTOxBhCl
9p2Ai8MchlIAVXL0gUuSxc86cqwadtqru5Urs+9bMgxRBxLbqnmYHYES2xMifV/23vqbLO/mZ43Q
Wl79zio45qZxrbOCWmWO7rfzrxq23D05fP/RZhpNg0lstDvaQ5G7EaqMqBX4InbtN/d7IT0g/akk
CEsv2TyzUszXPyUlryZtqedBm/IcPZkv39hXQGVYe60wHNe3iLFxBiATdXbnYAtOPwZdsqiSvL0U
sXw/m3YtFcrG8CUWwO6NP+4+WuLDjg7t/gfhTewFc41N6Auo84StMhoAixszB3V5rcLAzzzKF9Ir
xPZ/NHT0myVGBJ+wWZQwUpGgu4yGeyPbNdgTzIoPiyQ5idU5X94AGoD+Wzu1RKRIYb4FJHQ0rF00
YGBCRQIZ7bctF+EqeP4AlrUYSwhFAlhrmJlJR3UsUYpNZVoFqHm3lneq5t2e1Bk0gcuGLtMM+/Lt
Xyh8gX3HgFgAzY7qD53Y7ftBDvPByWhsgLyzG5kbfO05SHQfaN3t+rBGuDh2QZdf8CAPPhmyCbi4
UQPg6pU0wkiamcCMoyFW70sMtgqy86OqureZ/pGZMU5jbrsfuwhYb/tx+Qc9GiuXMRNHt+BjkaeM
oETYUcPH7BhPDO13HUL26kbvIRi58Ig8ychCBnMvC/t3f8OLlwBHKVRgmFwYWKxMCPNUiS7dloHW
EmHpE6KJqUI3AXNIkaFfyvLg8kdOst7GDLoRYBn/fqmqNWPkquHkeIgKvTK9XZYif/dfzuTvkPes
dAjLZtnR/popJ3+3IrPs2VP+ilJBJFzBOJCNdpx15qPwTiAreEriL+KJO1KbM4sjEaIjg0wyaGOv
pB0UMqf7LuAF35PNMa/H+uZ5rEB/l0cMK02+XRTVBmIFyio1DxB5t7rXpgKFQ77trn67J7fWlgeH
iZlbGKzhoyI6kAdpljv0qpeK1G9Z2+4C8+asmNuBe60pCviQKtzYyAmnZSnnbbBHDbFqgVLqfBT9
VHOsJJGFK5G2eie3+29Oi9Z00KkbzPwJAANLg9CWOtuXG1eGaSKusMiPHWipJXDZKxCeGItDHk5d
8Z0pvXiKIPKDI9zvoAzPv/30okDgAW9m4QW2GzWLSakw0EkPvVkIw0aqBkLaWnyRyRkoBbcdvDhO
AQ0kXqh7f4vxTfFmD1iBIFuNrWeT5UrlwYp+o6D6laTR2JkBxL7wKcXImpazaMgcvYpx7ziV6cGd
YbbyLK+DLPbRVFNWdmVE6cZY0F0jogywkLwiM5B/I/hTYAfXrJjX1aOl6XCWtheIbkVsTVaqwiG7
3bSuk0G0WcdfPC/tACZVHoQhEACimyaJGmZ7ruN4vmfXklDiIOgUpmlxnihffaC0QKzjqATBq8Uz
elLIYuB1KQEqpz3gSD6Jhah2loK64QhaaUyYKvj28LpUKnTrowZC6IM1UpYMqLRK8Qq7jLLs9oZL
5gI4zXoXEfDYuIsq9UAqQgOqWi2TWJ6Z8QNVh4Dx4e0v791Hul/Hb8PkdP2aEG5uyKw1UlWSS2nH
5cxVWobUgi4b1RdxUqfDrCL3eYyTBOybRI85RJdhTOPeMcfRz0Cx+32sbiEhcVPFnY7op6lAX+GV
uGiw4FeI+3rnbRs5omxKvDdNTi6aFnW2tlIB6SdMRYuJbm1az3FVfVRNfB8NSKFbfyzOjr04xT0r
ed5SuKFURJ6oWOR2MAYFbndlru8jyYIXA4bD1tJaT1o5F59+b7S4UYgZG5XhXEaRIxy+sSsJ4qtG
fyUSfYR2RCVbvGavqwJ/Yo25cV5vmDAYdwd7qnFpg3vr0qAl7pVphygH2tIiu16TBpKyUKhxeUCC
cVW3B8yHMVWuBgE+gVv5RuhDZZW0BeqSyaRWJLW3mqzo2Hk9Ycti74gTMnb1aWCaFZqk4og0iOCS
46Hy2j/8/bp6VQ1RiSXppgfNrpcle6tb4l4lPSPw/9sk6HN749xOLmLctVUYgJG3/+vzQL6I0aGa
HBHm2aBvzckul6vUC7sUtmp5zG0CU/wOXW5g6KA2Vb16MIlyiZhMre+nlKRSac4Q8iP8Dhpa+B3V
lSzMnsou40MbqjWMoj1ShWkgQAOB37U99ps9Fi/fyEAVYwApM8n99852/KA4WR+BNbwMAWBAS4Jt
f6s9UMbrhNS5tlchkEkbW2lr8YuXBvDG12jEqfA4YJHFvxyt4wm4V5vfiSoS8eHsAcqjtJaBBSor
0HtV9u/7kZcxu46rHVVVivU+CwI/RFDuF4UsPuCzJWa8iNPIycXT700QRfRnAcVonNgjGDc6f0Ph
mC95WK6vJpxVYP4H68DSeOioIFIEIK4R8ddtTsnKIEc2D0gkkguihJbYKzxVhoU1k0JtM78D2bOM
itFsTJ9V4czsfrAbCMBdEqXVLK/lE+HPBY6VWq1oYE+Sp2F3rmhJYDmiC3Y23zGgVU2yOaXkoAkE
R2jwmhTc39tdWkzqg3xxX0Q9ZfnPJ/cutAKLnt6zVbxp2CcCzEcGl1kcu/0CKYeyFj92eX9tMRGm
mgZVcU1xLrWDSqb80+HTFdjm9yHx0nigGUAFlrx80OJ4RFoR+vsTdf3FuTSZb3z7Hrn8rb0cIe9d
KCla9mnSbmIYl8ZTZjF7ijL+2JzB2+PZ5iDv9Ryo1SfkS8+rR5D3sKD9KVMSJveFQt1b00ClYlks
O8iiVl3HyLQWl/RdlT/ohahLDkyGT7mPV1fwwg/WcaaLbRERrIe5woRfZikwyDjIDj9TCUf1VFeF
+I20BPilJ5/KjKPIWel+BdpVuYRH0m3hh3+JRwF9WTo3N2oTlxpzBlRNAfnZ1uE0ZvxzmNfjqhFC
9BkoEiymmSvsUHiQSfrXvNGVsgahE+//VOY2GOMOUNBrDPJg3QUs+Xb/1O45D1Jb5s8IoPJZlpQM
NrNNzt0wdxMIkZ74TlMDb9drkLtMk/8jJIs1dKhdwzn8pqeUuuiWHt6sM/nWWzzlwY/xoP1E/qZk
V+gOgHAGuze2F+i3a+UV/CKRGfxhOMlx9UI6JUeVF35895u+ipVX0w1UP9KCKc+NmUimwv0NNBZu
xkh9nVjfG7iyF6H/z1MFJUDi/7JCr0U12sjw6VtvjXIfqZV54RYXojA2cjhIjYSpD8PK5aw2aK3l
5nbidfMbsZOluQi1eUNdaoko7Zml1BcnU9ElW+qQfBKHrvHV8Zg825sOQ5Aamy7Yz4iZnKbHa98p
a6kYfvU6Z83fFFiOzI3RxsiZMEWQmcD6g2H6iuAK9HiwssVxcx9n9l62ul8V5q9qtYSdrUT2UF6p
2RCOLFOcQkfmRvwJ0fcl8XNz5raO9ZQV6JK1Kp53IzL6N7BwaV+SvWAlwAFYdkFE9MKRGE/29+Tj
hJfsJCHqTsZgPBok7llHl7f9lpSdVVKym5l+K2Ul3o9Ofpo0MbnhMxNjGPx5O9jeU4ChDRQ+VWCA
TgJp1lpkPfIr3iejZekGrKUM0CpC2xJu+6cSXEbqS3jaaW0WmIWLqE5hZpN3WB/t2jmkWuEPAiQ8
8wXl0yldEoQkOYKuf+kS9JJVR2tOfEYnPQp6X5to5M6zrlfN5mGGlSr4k5WqfSAaY19CLVbABGMc
ICvagw4VidGZyLzfi9dTCLu02azKxGOCS30Jjdl/C3wk+uLlZTkAFQMFfLt6UarHK/Xqkk6On++r
i/BSn8kPeAQTuCETgBcy7Pa/Z4T1BfIMV+090xelXrUNKotpTvQchxJAiVcIgW0RcBWm00alR5St
vPcA74CmxRNkdAcu+VVVlK3dk8pvljVm7MkJ5ldk5OYLAYRzF3g/Mc9YzcqeraCeKDpMltB4oWhB
PIY/5Ri9AHPx6bwXLqd+W8U14BB4X+rCm0oaq27gbo0EL3Isad8M+cyWhu2RycRxrPNIn45P/leu
BD5jcnz9RWKXcwKFHtE2pmioqsswHFq+Xom0ru2CjNMLKYmBdkbOSEm4ssrwtJWVkLR07u4ZNKIS
mmmlJJ0TOVLjAjD02VH4OqaOAwhPiwZMs4KFyINki4KL748keBpnF5tsTe8MMP2rj8aeM96Jn6ik
P7j/5htgcCej9lls8D6oqCl675MrEQL+THpyVhY2EBUIyYoroph8km+wT1KMa/Y4/rOHaulfSgSa
YiqZgoNvlWGWNAvMksN2KaIJcEiXwhSutA8xZ84abTxbskAOEjscobFo7+9C8f4dgrdswzsyt0PZ
6I8NYdSFB6HvOhZhtPVhjGLWpDcxe4gOh8PxnJiUmtg/ULnIZ7obO+EMAX3YIhm2BOFsvYf3FNm1
UYw+NgYpNha33GOXBpD7ZHTGscvqv5AA9v9lE8LpvVV6x/s6s5n3Sbl17bLbG5NI0dYD/HZEbEG1
Umwlg9X4gGEXb0tbgHuECWAzA3RqNCQnXzwaX6xJ/tqjNVhtCOkO7Sox+dRWNrwl3h8L9fyRa8au
wUUecF/3RrZtr5PIYvWQjJ27GiyIK/qbD5fT7V6vgvLYFjXYq3KGJWwNXUiRXC3wrtSe/JiBJ6i/
LnMQhkwOMz74kEhaEux5uiQFz9j1d4FiZ4/BzINRLAYwgqsjKTo8W7nJxzsmkRBV+4lSip+96b8h
AcDaWlPaHM6xnvdDkFAjxhHNQq5zqjK368f0ZomTjD5FMbzhuDk8U8rZ3hY8sdVVuJbV+WvJA+VW
lgAWEpCp/1Do18KrXYnS32i3ZjhnrPBs/3uKZhNMGaZko9vFJDVHM75MDxx1AuhUt5xPQc98zIIr
uytlU9LVI4wyZ6I44BH2I9qyq289mrvP3W0J+FOHhBaY9LAoGbVFy6yqdmW2BLpIqrFot7x0SP0t
vE+pyts67PufJBarZViVtu44wR8AZu9FxvSQCX/Ilyj/tjsoWs8THIwDGndJ/Cv8HvHJjt4bxIjE
pQEG8u5nsehJMPaEwei8XAjnNu9skI4bRknnpnlq3H7x+Dl0VS6hwDkssAlztlNQn76k2GptYpNc
7hVBMjB/V4IoXbN0NYpiysGL7BZm4smfQkY4cr3uN4pSSafj9yUzJITCbg+ETz48w75GrTk5YvCg
2z/6mW8AdpRZLM+8wBn4LiC1fYZnuC7POhFOAfjzVkj1bTt2vGyPpDdAULvHnNnjsh4zEP2/GLTH
kmIpXtcRQzROXpnk6grRqKMcx9M0yhMLb6RPKpgSlbE+5x9Ak/207FYUrLsoNqiK1JVpyzaLWAbY
auSYDFyho1kfZ8RHkGnI9CLd2gWpJrmlmvVZ0Ih79dtgC1x8x2VVAYHPjIB7OkWl/YlObK9CY9Jn
nrAE+ZlbaDG4VH/ggVLvVQEm6QounqsuNhpSfSNGXCcdugOoEtPnxUWRynRGVI8I3pnn3jYmFwWO
a4SS66mIi38ava/KHT+9CZ8wjOgE5SqCoBIGHALPZQJVhqDgEuNhMPlh59E5oKcubVicAu28wmpx
cfV4HeacHJXn3mLXBfqXVAcuCmG4Xg/ghIItUuhqNBH9OaDVcF29E9H7QwKvEtkU4i2iBhJh5lH3
wuUbP5BHvxGODlasobWr56ZSvIEasP8I7/6VnR90nVo30AkD6zLBtBN1Cf4lfMlPhMhSvNJbMsHs
42OcdRSsQqhZZQ/7vEeml8Rw0JQ/52lv0/s3RCKrNkms2RHl9NlIa27ziQdDGJbMc3Orf42Dq9j+
eHhIgdRLJG0/V43NvQLI2AnCfQ0+TLudl3CaPqDaF3IBgRsPOkn2V5Ceei4kJA7HNj1plNe0wkoi
KOm001K4cPznXDRheHoJIMrsCrFkjXCs4iYehm/vs7WPPzpWn3h0UAayMR5paJ7JSJrqUj5CzvKz
nDUUGCH1+sQsNliD1nlGtVUvbLxqBUn5CK0zTBlqyqVr697yruKieBu75vi7Rle+rRjRQEFhL/XY
TRf3NXR8z0Hixo4KhNMubaqvHu7cZ+RXamsXfMUexq4roBx4VKWeFt+Lgb6PksrL8As1NM6fxihW
kjH8On6MUoBZIvt9Noni34i06XlkRE8Eo/g//y6RYVq3Al1S9+Xru3Th5B04CdV+4G/DhAemK8LK
QdYrGwXkiB8lYpXKA11AeudVKTHxBfQn6B+q31As3+A3aVWBuwM1KzSPcbAhLSET2yoIWntKhQSP
cJoZmCHpBs4b91WeOWveMzvpTRbeeaTQJ7e83BmZNUAJXQyabDCMP+NC0vzWhUAt2T7YaHYrxzvp
dmzuzRdYHBTMR7+W7ApWxYefqfLNNEJCwzP99u4AO7gyryeTTtXnHoyxScHQ1kyw2THlKICY3352
kQLEVlZ00ApSl9ZE2Hb+3fDU18XoyBSoWtnqFTTGWpJj1W7HfE9BY6XMgN5k4Ig94Bq/m/cdn28p
bcaB28RIXKPbps0ByI7Sx1eJAZWGzLNOBq5z+5vHnBbNSJeWyu0dziqGP41yWOtA8lkve61XFajT
3ghZ0tVllxZQyiyt298k39Gs84Vj1A3flDuQjNyVm1fqK/6is22kLB7BbyP/IxmgGObsTDceuxM4
nqAUNm7ubH8QGNFSQAvZittVk7dRm8j7eLynsqLHNUNuX++4QANdC4b5Wnog/ERxSOJbK+y5ru8Z
w0gAvIHZ8T+8HdCIRl3pNlsHV5gTJfVhR2kyIb9T2Y5imq7kl9/j8fj4rcxwRpz9G8lmYoHf887h
MWBPb0OCVUI9ODVVlpYNGS1fCw24JCh2oDVRBxCKcbg1hJqPxwz6EjFU03iC4q5pwOc4U3JhXO5W
s0KrO1hp9m/sb+vlZVloXvRfsORV7PtrWN6HcCzIQYeIC/p1Gc6s17hWbyzlLj5jTP5HRMjDGn9w
ZiOt0soCX2EHwiqutDuDE3sCdVfLhfK/zPSlVK8VWqBAF9GsTsMAxKibDn3tt1f3D9tIknj2uBkK
RifRsRabQEAyeDFhEvXEfI3iubuDpgcNwFj3eYj3DIYurrIM7q3eLb4QOxbI5Rzd3jiXQpNh9PXB
Wo1YqdNVhZrlEXlz0V9xcl27ej9RxYmyE6zOD7FmGFtYrgyi7laPocG/cDW/Zv0AP2/VYxzJHHHw
QCzcEHNM+Wg5WdBFfS7VlbRn/wvAoWe74wiho6KfVOpmJ/CWp5pbWJ9TH0a8wNG1YDu7N7xDOQNT
stKQpz/075MXEiFg5mIihwCxmK6CarZdUIMaDcyOF0SFfQLFb0y/tRs+nUWp4v+LZKoV+uys+1ml
JBk9j5d5t665Z5rGgN6IBegUNsKFEhE5t42jWl10UrHxc+BF/0TC1Uxis5VYKbBQn6aDdvc9HPqV
5HqStmu6KRE+D7iJIaQdlaf6+Bc0p3ArufpfZZHB6NnvR2G4GTcqkwfBDURTH9QQReAY0a8gwBh5
Z1Mon1UHFS8JpWyzJ0AGWKw1A1InP3uwxVifar+seCGoud8KPYxL/Y/E0nifhXRXIeuGyYP7IPx3
YayvyDVZY03x15elQ+mrKhkLUCQ8nPc8lBFn5od3NRlPATnV1p43gfgC6qr95Py+pg+tovBhAmsR
uUbW2Lqv5JaeLW239mzaU6PCslJxOanXSff0SrYXF/kgJLVHkX2KFLJ8Yi3Z4FOnw7Qlns2n9JXd
lBhD9W8jZjz6IfoFRfH77ar9T+5mtmuH2LeR0H5g7gHCGR3F1CADFXFI5RBwKXvCH3O+05+rioyH
5pG0muIMk848MROQgRkgL3In1txLP7tRpizCJ66dWv17FQz4/pUXR8RHTgCly2QvLcD+ebiTQyjw
DgfislFJCXbmcuac8uesDSdKL9ZEKqZKr/ThI4z1wvSDflwB2YKzTdWx5DW2gbtIe/lHMOk04IQm
N5bSIDtf+hQskDUMPNClwNEeWMHsM60I0uv7Gubvk1/E/wcpz0wJ55QgN60/KKiTfv7yfcYuqbuN
Z2KKrO6KA6CkmLRBjmse53cd1yjhvohXoURt0pRMvXufBXg12CYJGBPl1/AyIVPRQ6IXb5IZKk9j
Cb8J5M8aNDuNrAj3ZPq8XLHFficoU0Or0wAPbYflk2Pu5BxII+HKZc/zoYiuLSMeMwhRw601+Ri/
ieS83DtfWioTD39mV8FhtXcHegj/ob8d5WEgFd7YxJCuTZipTUb2OHZc07XZDUojaTya7ySZFAJK
7AGFBszK8y3fB9PAfspEB2pdoLfwNUXYERUIM8LUqth29nicNz5PhgmTPLPA5gDE5kkdkQsNTM2Z
f9yxFcs/Td73fph4X81P6kJtlbCa7nlcOaL0O0LLx5Dy9/V7Pa17gVD8Fqb7qI80Znvz6KwLASgs
frWI5fSEKo9b3TAPWJm1pRaawWkzkIlfRsU79FPnGkBcfkCVzPNqXQYo/5znihLNZq67W/6rIYZj
QB+HeyBKB1qCZD0MjxEZ6duycWMk3SQrYHNZl2ZirHomSfbZpGqv3iabDw47UxpEaQKtf0BDmXcQ
CPbha/GxDGZBVfaKYtVwxFs9h2BOQA0QF2Hd8oDvN6cBlfQwkqP9o/BJqnoINCJ33KpoPSkSc+WZ
ec2iU8TZYk6wdH0bqpxpSrU5tbXTxeWa/St4SILT6U2D+OQoRXqsknYszKzkVRNfPTiAUwN7zX1J
ffqbKtLRwHVt5UQMyujFI+pP5JLaEwpRoNcIkqTDFw1LPQEUrqlV+VJjo/FmoKJ181uetOsCQ7Lm
gsTVp1Fi7O1WEacrBZlcKpYGlR19RL1v+YDGLGqmRmJ681sqB6znRTyzPGsjQJbq6T3DPDs8EQmO
d81dl2uWx7wxpqChCiM6+JXloIJB+lj+BuuM7dNK70nQSCuZhdeF/Q0nbA7xS7hLHtTTn4/VZrsV
3QL1JbE3NICbCvBeYFMFTBB7UIvZxr1jgpYXT2SkSv9/OWbCSfizJtEdmUh5guJvrf0E3S/jRZ3n
KS/F3SJ92thBGsTF8grA9sceh2I0frqIi2pmOFeauvt9zoOsrZKyb6vyHVkwP3WbDwmdTSBsTFQQ
RwOXz0O62Z1I1Nnm4gezm6kgxkEXIck3YdBpJBmoxsCMplOWnAZhkfQQWeqIvsaVFlucM55JtdoY
b52/k29pyhFVPYlGm+SmqtBTBHWr3ZBtAJNw0gAg6OUFcarKyX8jiTL2WfGdqnb+wVWNl5W5NBhB
kV4+dTfe3MiwkA7/ZaejQLgZ//cWR95CwJI8JrRZ44zxeYDXlArD4mwh9NF2Jxcumv/gNVokK2fH
hPsqHGEoReVSSK9YJVlfQiK1NV1s2v9GZa3oNn7/a0e2ABbR0p0MDlyRjs2jG+E836mtbif0FebL
x5ApyKFaXT+y6cPhQH79zW4/Q1J+bQAjlNViOkpaGVVBbwVFFJSGNn+V3IK3H/azW8h8167Wf2S7
XYscUJhpyfcCT8KYagZk2E2Lwmo6OIQTMUj7kC4WyLfED1YCPfB8rOpey4RqRUcjiT2xqiKzq76E
8xSdb59cejydjgWXPaKEdPeJd/E5mqbDGuDlXAO0xASqiWW7gb1i5ERyrwhsBI9G1tCLCYqcAsc3
ytDCQfrj6FIyJcGaCTKs2eYf4J0hi6lSzZ6cJwcIEZyt681lg4V5t/y5teQ+SflzZb+AI1KwWfXC
63auAcIQ394gWWUFDXEgG70kSo5Q12etT3BsgW+WuTppqngIA0l0uuILIdpqEinEQpUfUW6olmcJ
hvniPqnmv6cU75AXAe9Lx9qOPAk74ajbZDAH68scQunutDm8a9Ooq6sV/6eGjTDvFSXgA6c7ivHW
JxgvM2wtI2CYvQFRWg9fTO3o58q1tgX+6xVfycSHGu23oPtHDb2JOsJ7j9xJEXI2bWHyu4BJsQRb
68MdMFxLSFJmbMfRVNy9NwTY599w+7TtR10iIWNQcy7bWAKNrgVWHXhBNa/QsGJLaxRjUKQe3vB/
s5SK57BKupkeGQTTLeaQoCKJj25ge1CM125Vc0OK+xU+vTWFEZF8LVtE5bII9BmOM7LbvKSOuz/C
vkI1ua+Mmjrj2ywtPcH1Ts0nKA4Rt5UATYDXe3PCnWaSRrXamPMgdzVrsEU5cKe2dSPq90iEltpY
/IRDnn9at4jN4yZn2Rgp20KI2beW5285fiwVogNP9FfksiBoOiGR4ayufz4DHfwtWiYDz4+JfmIF
+r5rcyhgJg9r/fliVUq2F6C6JZQiZtAFRhIB0Q+0aoHY1bgN/f5hrCs4rxI8EBzo15Xe5UP2MpCI
Xg4dSKDNlLNF/6FeJljzKjjRfQ1MbXkCPK73eISeikb6nybfnGV5ZtfglVWB57c9CrewpP4GhqJ1
P0RqzuKCK7ENT17/w+a4GWEgWxVd3ejwQsXFFujcDV3Z05iieRKXogVvAus37PT88cZAvoqDmQOp
OVnXRrMXNH1NCDAb/YtnF55Fm/Z9HnyF8U87uztmzVUxI00GlPtxGnv4WhK6plCAZW/IU3d3/wmN
kmYQYXgIp7fkYj/J0xWk2EiAcz83Vizfezja261e4qwB2tdynH4omyzPpgs2ZcA9e480ZBdDpk0q
UQpGAPFsoS2tRmlrceUo/Of8MgP87raIZB1sVZQ44j2upcENWgzx2x0k4shcaoXSt2vdePgHcfHZ
GL4rRg6UfyWLThWQo42RMAvHQ7cKQjbJQR9dbVwSjQETJ3pii0yNkBdgDsStAdQ8CFcwttWsNbq/
KxUKBjBbDpUtH7++Zi/9hbHUoI7VAd79+PT/c+Cji/x5ADE3Offy299nXZGEFQo4B517gBIIMTDg
/TsqcNXrTiWySnuM6lKzW0gbDPQLAUuzPu2sMPGDrM4fg/bsiIruCXOEEqMZPS1aSKlrEiD+9mfN
852kZC1Uyn4tvP4Zl+EcAARfKb0rkUM/W1hFVJ9nOJb9M97lcOBz2uFGiJLoODqWbJfwxC4xdmbK
LWzSgreryHq3F4nA+JQpgi8f7eiQp+fKiM3LlRS7o7fNL9gb/PwsG5wLrLajjRZZ80duIzKqp584
nnM2VWEDSRlmqSm9CB34LXQTz7o6oae/nhY8/grGkb4rYol4T8oh1CnP/T6cHCFrtH61ME61CZ5D
oHzEIh1SKRImbW/tA9xJiymYeCmCGbGjL+k0vgw7TGKeDOPxJDE0gMxkLgRmvXBcVjNXbfHycECl
pzT/GVQI6Nw5pm1KqvMudObJDXeOaZyyLjtWCiy7FeLapRrwdfsXEQUKQevUdEAk3dpnL2YNuyOd
rkmxtCLhXGNg9peZA8Ll9K6Dz+taW8SlThFRL2zJmVPkaklTLrGTgvbOaTJ32p1CY6viCSyqzCLh
5rQkGq4GLFRchx1380RZaL7nXm87IwRTaKxLSmEvFU2TBQudFS65xVpK6bO9vpQClgosrgfaHFgl
+1XIXJzTtMV+YZJzODERcO+AMPvsP3nBJtsrYU4OKN5x1Si/OcBEvPXdIwHaeSdiTyTE26lui3Ug
2W8wM2YtOXdL1i30HUGDnQ5zW6t5ljZ3lQYe6W5TRZ5L64VlIdrxvhkjmTnHLGMA9Qk0SFFcoxbN
ozc7BP24oNW+BZbEwz8KeMOW7TxX4nslOPW5ixup7EG7a3UI9ppiEb4SkCgqolLC6I4vlM6uJHLK
zZq6DhGriyqBQjUyr9pSOip1G85PgO8JaBq/Y8jOVOgEdYNMT/QO4YBIS09RDGs3lwtuStWIZ27l
3QpjrX9TljQedy/94zduqaLEU+Z/HZqpFom7AVSPZ6sHHwiFLwaNWbQ74/JjRbdmZeeA2xz/U88z
BqXCTngxVqUVXMTOR7UaELjHGM9KaBUBgZUDNbwbWXIr7UZD2bJqIpWK4vji+bxmNPBTLaXUOdm5
h12S0415V3lRwkHJY9ri7LMkdbcU2FNMbpf7MeRsthHZ1sCrtCVrwtNvJuT9Zz0SEOzANhjvhM0n
7yLn1bahtp++TgZUKS+IP7lGoF4X7STxXCEUzsng9LP38YSyhP3OFwE+gDXpqoEHxgyy1xbJoHDI
+8+P0w4SkZjpYglic0mQeapU4v1hgZWWfUT4qSYKUJuOixr6rsSsHrUuDAisV+WdV7qjMRbvxzyw
aWI+iNb0YNSbGg4WIP+LvFMEhFX1f3RKSLgUMVxjBmHzI87ilJkp+fQUtLz1sB0YyX5F7LvlcErE
mANS85bMEPPGgXSDs1BWQ3kejvQ0OPcTfIETL0Kk9OtZ6YdhsY9JEvR9bra7En44piTG157I3HEZ
D/PzpYDMqmqx/QcD0vbAemRbiWzWubvMzlAhcZe46C4qR7GPwU+YnWYF+lWY3JOXf5BxX0WaiqvL
QhsxbnsN+ALIreKpquVnLiMZvQZyW77f95oJwFbBreo0XBlkostxTzuOCGClB6Vpxh0KaOgQoiel
OqmJaty1iveYb9hmlkvUXCuqAvq/AfVjbLIiheDDoeO4wT2aqrUJiIei/IpPvLGZxn9EWK3LDej9
RBxJt3tOjIDFEL2N28erd8rqzqJIihjiiKkt9JaC73kKM59XOfzd6/J0MtFFzdIdHh8+n4D8VDl6
8JK70oSdBdroZb+Bhf/4iLpbhv2qedTyiw9JUkukUpFHJGu73cv/fVh+nJrwJeswC8A5z2VeM+Z6
JnwWn7ASbqx2AQT2gZ4RA9YVicdgdeKYr69c0XcnBgW5CTG0CBVg3Rp2JaV+P3QMIM46E8vKid10
yP7jiYMx2QDlFNnZ8SEMVJE0MqGar+JeWWhLmx0IXYPFUhBlwMoudDo+WktXA76BKikyilZ3EDkT
x6dPhzhT5xe5pfd8/iLBLIUn7zBIn/KoTay1wkO2chjm4PHC8HepaWqsT0yBgg84UT7VBMC3A+ji
X3xqz48zAaelscTVCiPsYob3+Un4UxFaCjpCH5pwWfvPnoSVucSQmWqG1M0xpx/u8nZqnh9yruCt
G9H1iixuOOmj+Gufk5rYVzOQ+G0i6c+ZgXtkXUx5GBJsNRBahrov5o5mm5CDPbh4OjN0VBmqZouv
pUrD9FYTInecTccAQUPrh6ErOuLpYsWm0FZj67g9FmjQeiyzZ227Si/Ks+vJDFwbHP+feOQUbOGO
jvHGYNfPjDSJs3jVqBzUgLY748ee7N0WdUETFG9OTVezpfcsX/2zBIW2sLIqu7zoCXk0hfelcAcz
xNeIiZH6KbSEM1M1wiLV8hwnPsuUVVWeDJFbycMzzYZBfoptVHYTX0MT0GBeic5SLybjYxLtf3/i
KrtZnak/9j1stpn8nOQZIPV/YMJLbqBjZKJ3nmPy+qCQ5eZK4OzUB04Y8oC6q4n7SMiZyWKu9o0t
v3r3dxaYoKH7T1W8fp+yORKBG9nh/BX7+kyw4YbxMQkUyNS0/CgeQHpH0y1GCoyZldpJiWS3Mc11
+muuyJGBs3Up79qa6l2QtBlgKcXb+mT8QBQRb50uXMLy7jOmwE4UWEfgjABW/zmxzHuXewYYhEIh
K2HYghEaiX/Ppv5UHeaRQoaGqPzVjawt7YjD+fs423u2de/XKeF8SemDDIWpAe5Z22M/A85PlIMI
bPPbJxUkKdaKmKA9HiNfwnriT1U13wfmr7Sh21LBFVWrmEaXkGZLNFEZqwDeCDz8N3CA1fyVtKqi
GRpJJgP4OINFNl+gVsE+lCQj/Nzn/tTcK7AAQT8yuSXi6prPJP/VzgggmkxZh7HEPwAB9fBulbDM
n0Wrsr6jYvCby3yEgx84RwRt0uryNv6oGBsslTNKm1lkDdTABOUE6QeconOy1wUjPS/26Fj97nmU
D/kZF5k1S39Kt8dWN2K0WEj7r/7zUZmgF00ys4hGomhiDWc9zqI6ECnrEuJZggDpQ7MZG2SnTcpf
uaXZW1xKvIPz77lrG0/5Ofayni9jt0t8gYoQE2CRbMH3k+15DMHj9ZkisypNLl/p0GvFH8yXG60L
jwzdVYN7IhFpHg5YwkdoFB6+nTdNYBzcC9G9fEmT8NxjNaFXgObwSMcyPo68vTUc+kv8+ElRNAZy
n30DZNhPBssrCA2n9Z+ytyVNMcCq0nZo94e2jN3rwb/eL20ZpkKivA3iPf1dxaWgo8XFyzFtPVfG
5m6N7ZTNGC+Dn0AQ+iWexiCmkaT4vYwy10PGfQSi0Tok5P7jX17ncFn5VkcYc9LyvGMXjcRFLBlz
WFBZm7m8gTDC3wuWcKsPtMb58k19DJJnXh8ZUZoNwPoFvghL4HmJcQyA2aZmX3ruCPpVVV1Ssb4l
qwlL/DgOM4JWK9ikmxW5H5UwZR5XPgxUbWMWfHyAYl2vvtOm7cC2nwDaAFJxc3zgZ/HTx+QiAnLs
IfxKdmqb/6ukOQwuHKzQDXRzORCSLoHmzRcUf06qzqOjce8hU9TaBnObx41EsKCt0uerLlbQPdrj
lGPns2HntM3MDjZqmcypJi4kYJflcq7z2dYGTec3hi5DnGxEGHIK7L9NkbNmYinU58K9min522hI
Y+D8GPY1YkvMuSO8YZFvrOl7dLbaHrxdKhEDCO8KRWMjrewzgCZR9fJHitd5Ln8+RRA5XFFSk0PC
353xsGWXxLWsx+iYzjBxDAefyfW0S4PZrti5qO2Kzph1/45edflF9oWRKVzcy1rxSPqI66ZXHR/A
0yu0YfG5gZPuhS5vxufDhMc7vMWevuRakAMY6hvTJSoeC/r5vOX+48apAgNBBc+8EQKjkc+gePEL
KtqtpFlPudQEy64Lf1bxdK1tp7DV4sna6ebHpfDRP9EkufS4zC3IcF87RqQWSTm5hf5GZz/oecqA
X8/n6h+UvUCfeEIIYDh/bfOX7tjcBX01GRh1JzEJoflckpM4nxxPNUJKCkE9G+l7z8FAdNUCD8Hr
I4jnXzOjGL+tLqjRDjhaFaMwo3cAWaDRhcloBC4UjPwDElRYZCY3Bio6iv3ONwJn8V3SM9pP8ZYw
Pa4Vv7FemFf06ys37YgnXbxDqRahPGb7SXg5K+aM7BnRgob2SzoG/14/CBtqGShWJmrlNxHW4QvD
SYlkJRsXM3Ua1AJhUAwhAdUK4vjHsZv6maJd5jPzMpjRwGVshn40Mc+BA20YOty+pMqYBdzTMmVq
O30Brb7j7jryABHgNH+A+jvgXdVAWguLI0Ri0C3Ab+i3nEz6o4MQhZfgxLy82OKhxQj+T6YJuujF
wuuLenUZlQP7do7Ybyo2iIOSTVc8SlTSW8coKXvR/m+iZe4thwktTvPEA5kvbkX+Ai40G2BOuAjF
ix2efrY/hsGU08B0jiS0jltphhnzz/a4QAncOXjCfsy61b/UD/jDxKj+/AOgumwOpnd7XfoMDz2x
ve7lqKqanljyPUpQ45i4Y3RWpUg+AAJ6WQGGvfQrKURYQfrNr4d9t7vbAbgsQr1gmjdlcwCe55IE
0H/b0guwQ04mvcSeWNOoIIY7n7eHMqZmbfPR8q9HOOcJLNYpkzl01+Bc+aHZ8ktnXZ15ZRRpESQ9
4MFSFc8CKAuqqi7xYlx6jfaGs6pzcCQSsGkDizlagUDw8zMvIOs5hPxOkSBb7lU+aMPlxeHGwN72
Bxbk9XzWZBFL/hu89r4X1/L/k9xndmfsU6i4EbsqUbzo2AHF3DZTuB2dJmW8gHEgcTZPL5TbvXW6
8a9suEKwBZrFEeAXoPckN6zB/cei3Cc2XiQikQZ5eEnMmxbGEhL0G6JKv94p+QCjo7gm8/N6pFmp
j+iHdxChiPoh+HPFrerVm2pYNKP+lgAfuf/3ErX5sUI+U8Q+bJPm1LsMdxsDfXFBL0an19VGpcYg
UjCBZz0FwdUzj7QRgmie4CIlIAu4k+nOcN8zVEIif6fbWEzp3GATXLgc47jXyR7KILqw2vVf/3dW
a03Fe33922mabbXYYHM+3BGLFlqXXqVzXsrGZdXbg6PiL7Y2MpACmXJYNuSSZIMw35CU1AwtKlRS
CpDOMy/FNGUd/D9Wm/cfCcJuS8HuaYUQ5xkIxw+b9zd3VPAJQQmqeB3yrIpvPDqKjxgTbb4wYoAv
qHpvmh79oNOTXlB/NTZuFHyen9ztvo/R2PT658/jY+99kAzz/hVNk2bvA3c3kiIRYjWZ/DLLBaZL
OK2T+IpTJcFPe+3SYR80a5z/hi2wTxdh9o4fFM4Tzmxhs/jWJDvO0gdcMBcoCqoU2H8GmmFK9H7r
6KyS+xUAUga0AMZEqWubfG/iT8Ti4oEhWL4GIdPGfbMzbmVaMsWL0x4QeaMXdyqXUMgT4qoklYWZ
8AWC6zPowbIGCjFrOhOMdHz0HV4mqWWuLAcROzuwCa0HimfREZVyU3FtgYodw8JYWMM8anW/Spok
ROvM5J0SKlqXL1DoEX50EDXIBm0iU0LSSM+ew95Z5eC6gDokVX3y2YFQHCBLyr5Aizkxs0N14Ts1
5K3eKfN9HW/9dAnlIHYQoswcu9DVz7RogX6FrHjR0g/1hL8q22E/ByP16BnzRVsGmj4oLnfYTGKt
5piEvJ9elPK3P5l+9TQBCY/IC+V6cIImRE1P/dRi+yJz+DEQO4ODg4gQDsfYIs3ZY7d074QQLBdn
GYQW8JHcJO75XR6f4C5pWRP/JCDXmlIdmB7ocgKjt85+k5pRDzImn7ukUASwpNL+PIBlTPC1bM4j
AJevVnpqlfepv7KD1Seyhg61MXn9d+hl4TGCxpA80XZtGxB+A97LhmrG+xFQkvS5rGSChh1oZeux
THiiiKgq39f0AfMEEfyWrlmsXl3a12msFoWzXdmrLlXtxILTOvqAjqPF9Y3MYbHhbMlZ9ZgyGvaX
Ecp3t04lIzXPmhli5HzBGn19pE0TSsCDnLfMFkHd7DyjKQc+nhtsDvGZ3LM9o7YQJ+ATawaIq+qP
+2zzBb2esxcsjBjlyHSBAsSoXnKXTlsR1SzsY67MPixYU/pdVWxUk7qiA8FqDMy7VJyFz0HQU99L
zm3zhZA8+VirS9X+wL4OvKZarADhEF2i9aIgvd0qgA5w4eaxhWBA66EO3twaj39c1GBTEd2Mq/ab
i5Sy66AAx5i/sSSQ658UW41hTNRy2Avvlwmx0Z1Q8gNfLhJYyVSYXqvBondYS85KB9lRpg69ZLDh
Hjo6b8rZP42Y/NwXXDjBjXJV2vaIlHCpNKhSWNAzCAF7knYvawBMpg5GWZprDNbNDfmgKnBNdVL/
qpNXZJcf0flqrrmHw1wXZ2nT8CvXSU8tOEUGi4BnrdmByyWHJX7Lst7weeoTZzMlQ8hoqJ9KYSMN
ZBDroOSxn0ZMtfdTAsX6DecLCRDVBFO0ZxYyE7cD4kIzyjv2sjBo+evsaQhuNp2pcCMRU+19WkNZ
XW9tUgR0okEjYYCX9+5ArEr5pnEKOlwP5dDyRV6gIb03l9SUeY7t3qWZpDHPWgSxoHoUBN1vRnRo
C3gOouaygZhtu9ACxGhtCsy/KA/hsal9kGj6eSHbj/QMLQQm153TdDQegnpYXsJPh6svx/Q3xQ71
CVzY+Agu1jbpy6kqxp0iwVbPwJycpTn9q63aQY5GuUpgUCU9E4267frzEmab/2/+U67q+VCzYXRh
t9SYAcQ1NQJi2rPGuVxVT9gseZ/rrv0CVtj4Tsxsmup7Rn7hX//EotRci6znF7sccHPGWhod9gFu
U3N1a+eFaJ7JfD75MRDgxvH/dtikr0fIYL8upNnvURptMuYZv9ElwHaDDLZoR4TCb4OYu/IzLiX4
eX1EXvit57ela1OX1V0cLiaskPuBaiH4RhNVmrDTi0czLPLOHV8bdGZWc8Fp0zUorC08Ybn8z2NS
+Wu9RogSZpCp1E6MOBG92yRgWUhdtoQ/DTS/+BC4xHrviZfJViIFmzr5sqSgOLiYA3Cj3DjRLsxT
63qt3K82X5M/K2n9HKxTmgKQF9G85dXIDW5hfFPR+Xv+JossEXaFNHpxeqQ6YCVNuVDtAX4BBfD8
n/qCa64CVWdc7wqPi9pph0yDxcSb4n2OolV2ofpveocYpNJ5m7FJV4o302YlHcdnRjdDXIsTl345
V7pIlNSAxejnUYTCbS+kH4zjyp/05rCo+v7EcoAg21Hv9XBwlVtF7LwUAt/WDx0oUF79uqACJgxz
U6vrDe+//2O2hayd/t5XreeUtTlSs6xzWmPpxvswPAUQFoGRhZc7Pjvy5j2J2QvCGFp72HpqeNaO
53Zname0YSSoEAW4lv4qh1hNRR+RhUgL70FOCV0cT4w2zlRJyTAsjEWGwLMXNaQY7mHrU4HxAWDY
52pEZlCXhmO/9uBu1zK6Zxiu6zTAF+Ge6lsamjLwEZOnKZU59rd1TDI5wSTmH+8PDBU1wslBwAda
oYhPwo319mMfc3nMa6gv8+O4QNtrCMToVvQ2fiXBYBtWt8EPNmHXvb4X0Ar5lHflhKS6DqYqk5eW
rBKGESDQ28H4xY6Gju9GwB7AWQrDwCpArHOpB/NfBRWOybYUkDyR1tfSSIramMb7pgZK/kDlNwks
a7eCHdVwgEtivNQjS5MdnA4peIRlcX4GByca7oVi5wcA0aa+/jBImojRclR2ZHz5m5neliYfNv7p
fp1rAjV2qmfzD+bEAgwyLiu+ewyngSVHOn5g5VioJtbZlflwgEsZKryOCX8aI0PboX8kcRCMFdDX
CzBJ2dF3kJZ/wtATKMLO/ue/8/x5xIE7vrOdrUOp5XqeAAmWX5EzuJ0kmowm+VvLMraL1INrMlJ2
Ub8kWTKC0ComSsZNkDcEvaNhWvYXH6DucQGMjC3heMB4cnzJyN+VyiMq9WEseHKmoVY75qgI4grm
xoPehGDOPgHVompug4P95+9u8xCxw5CQ/CYF/M/3PwSQ/QWYVc2KeSXbOGY5IV7jj0WNFTUdrHnq
8ETLWJ+mbESnwyenCDl5+KenZHYkofM14o0PnXK4F9VQNd5KiMXFOfvuRFX6kfVKSMbg7bhGajZt
TAdQxnfw1YxafVmREA4RadotX+k9lSrbhQfj4dpG9fsEYM5egrGPWeAB932ooo1IU4jsTaqBD8mh
Up07NYLvuD9DMujpFHTDQI/yly+N/xIVr+qicNBckMgIWH9Z+gVp3Gh4o8yvMakBS+6QWj2jLvZX
uus0kxscgnzMsZlvIdZe3htiNAC4bNoZRSn3f6dzlmvyj3XgTxMsNQvMflyd1F77M0wsxAYUnAAR
PA9ye75F1im4DqFOMEGegxZ9x4bd5iLWYvG8dDspHVl0R/+DZu5E5CGfIHVEyzvrUfO6Ww9tge9/
EcS9XCGHgIxj78X0O01ZBNTzzXjaB9Rr7FmlpQGLFdTeonqTR+zXczSy9nTg81m1nm9C7XVCpZC8
m/a19yMVUCiXjeSfJ32xbUPTHRrpUG2j6nVCnjZBGRbImFWDizr8TPagddoXSGpZPWO0Si0Wj6Pk
xa27pzQs6ECqep0ZucVVkfm7nT32zBJPWRSNlos+lPUHnwSCSO5IuSG09ZyWGMACdA66Dwq3vHbW
AQypz9ZMALU0VGu2QZQwletULZ1ErXW2Z78VrdvA1TcxOWGclnZYGtidi1B6fQz4OH3PxNaZVn60
I65mJB1HM10fnjSFqerrYRABfgnqHal4bEeHEL5PYDHGIXMPBWX0qghHPujro4kzy8oaVqD0UOJh
oyPpK53ATQF0XQARrbC1J3rPOLIiOgL+i3c0rkuQXyCsq6OpGfGnXxrgpkqP9KTCeaKElJRe2+DX
twkmdo7y/hT3eA5YtB65ryuP5j/OVv0YDqRuegBmjs+TjsXoo/2VEBz1r4Pc+fE+Qz7OfPNdqnAB
XanDx5gJz/Km0nAKsLu3byfHqrSWj9k0jnMk6ShG8yCLmY8bSlKCNTIZ1rkQDxG5p+pLH63pHwN/
ZmI8hwIYSigIHTayKXm4HLH5gYYOVN2iTe5XCeAb+A2Gwc3E6XXfKiaLtJe7kmcwHso3s9gXLNIv
jOtAajT9e5D+38p4RC+xI6u4m84uM+Iib2bwRQTOuQuNgB0+iEdlEUibXl4OyKChZZaylFPsm1JP
tDyr5kxQvE4Zze424sUk3bJzWdEpPHp2AEJLJUWVnByzeWkqGBh6zuU0esgEgO0pk4CxhXRP3FRC
9pJsb/9u3/9Mc3EW0hu2VYYR5fusyAWFgqtPZdALxeLRCOl3LgXQhg0yRaV5c5+Qt7py5CLCZfQi
BvdSQ6zG9ank0b3m5av9+s70VKlxpaSno2zwKdc8AgQ6MuJbQc/LVS9n6QQWamv298RiCzQ2V/o9
uxSzpGgTRT0MqnEVv//gXnw2XtY8exKbu+pL62WUk7GZZzoPmJOPSLBDDBizAIxZIJm8V7fA1rhn
Ejs1tkqreLQPiKXXFd4VutpYZasJjtCT4QgU9s9cvT2SEslG82sqtwglqd56ynIVkJcz6Vk9w9AV
mZkyG8V6L6C3GOlplc2IiUJcJhvXJduT3DuTJ26UGRJTzEXUBIL2H1ckC7GXGmwcQoGXi0pXhv9W
UxNzSbJHeudywpxMeAO4i1YxrDNdiH1H4EZkU2Q07BGzIDOP1xKQCiWDcpTCcP/57NqZE8KPNy1J
MZjODGCa8PmLQXtrIWFfXO6fJ43qs9d1lYLumpwY1tkesrTd0Eh3agFIm75hPL3H0z8RW/F5VNmS
Jj0Er9TAKI3A7DbZB6P0Ab/whcywCaq2zSByu3Z9wnt235aun1+Su7nmFsnbNltbyxsiN7fdrlj0
ODiIcfjhMsmMlcyUWHyfiFMvmaWR+JCk57E7/FG4mUJaredd82/EfgoItzsYzF2FtoL8mYRJA3MW
yJqe3/UH/FXHdzrLkRR9+wp7vLh4M61Z5TDTQ5anX+Knn5h2gemeLVXLeR2Tkgbpjh4NgiRYxMeX
dG4yXi5paehkxOLokpvzT5+sRHvRMUBqvuPXfTdLXSNaYh1+IWfs/MKAtT19wXkjSMxUL6PJM+an
1useadEWhlRz6DzwBf19FVNnS5Lg/heTR1ardx+ej364bKvRzGJFX7zalnsYVQQA9WphkcpvXKZe
t9ULFcufUdCBYX5h54ekL83QsnB9RgPDkWDDWBJu5jkYb/HfSbY8l24pCAI23rfnMIOK57NfQglN
kdY3x4umpMsM8fwhshBJs1wu4DJt9RQ5Ezq+E9x5tceprWacy0RDFxC3FU/9Y9jEEK6UAg/GtX7e
cbNTBg3DaDW7Svs9o+EfWB8QmNEbEIqUVqbQA9FIYAI+PLJLXxhdMr9MKTVxhCNo20ylbLG6g9CD
6FcULDeGHM/+pEKmxAgqPuuKIDCea1W3HSK9DXZgAWMpc3QZAfgB6RJ3O31biUNsYnG1KZzTdZvH
UODxLR5eUPhPvNDXuWw1Te1tGT7zirdvmNh7rEMh/WqpCml2syvxhajS92eHxyICrT4Oru2iXivh
I7v3RaubbVAa5SWidoWm9k9yVeM0vK+BPzF82rY+9z0++8dcpeJyFLOgqKVeFNfn4ighvW9OAxee
kKaq4/x2K+I10AopFnkUL+roaes2dHZe0WSmj59bUQOh14UwyGUGucI9dHHWeK1VOE7iJSlaT8zf
Bb1dBrk+JhQg9bMXFea97ZUGrXZwC0fCUrVD/6yGDKdqu9du+0E1SDhhVyXcZu/edp7TAxH/G0Rn
LN8Geq+DWC+A8uvHdZG+p9foAAUa/v+EXv/NaHpV5pgTlbpU9V6DHSfzmXrR/m/lYDqK51HDmCMy
yiHb20yju5uUY8ZMXq31aW/k9DFtJ75N0+/hKs29By766R8J5bwUok4PjCn91wXtyR/S4BO1XdtH
E2iAF5pK7UX4FeTjTiv7+NSe7oMztEyz9vWG8C8axreDGgi6Xz7jMbqZ/qSYqN6648MPcx0Frfjm
PfQSIuudXwZLwTbveYLdyPniHrh0aDJ7VNrdKBsIHutbjANa0gQh2FHQEY8tUJDAiXK25dvLY83G
/c6N++GotjnqXUdEDXRQfHPsrAyrEjCJIyC4+FCdjjj/zd4wTD4/DIF1ZnKfDp7YFAk+I4l19AhR
0CfW9HiUkWTDfX7iWknjGv4RA9r31ZNblB0lWSh6WeYvmGmeY7CxprqqESpMFkz4Qm1f7ksmDgYJ
Hip0V6lonBISi32xYtpcxtnkcXJeOyFt4E45W50HRhEcnAPLCeyyP22U2x0FYuUz8HNn+y3PHh20
flwxt/w2n2uS1xw8rfOacfTFdicz4dfiS2vM+h+gTwjrkG3wpwVJw7vFn7hUWfRkVuidHB10WhRU
GBX2QKVtmfSFvYvAQehXkRh0+M83WRyYmHlEB3HDbSF3I8XwSt0wOUt5UtxjUtStC2Jnz3D72UvG
bq6olBVTWSMOcf7gbzcLP12ZLQUix973/jBV65VdR6Kj3uxKMH/KMKA8md9eSlyt617OqImabKV/
wl92dAFKZTpKB1ifP62ymKRsDJmVpT4p+TwxZFcMOnbU1fTorEUteL8OWsUS5kZvSrqiMZPyuuR9
KgUjkCPCPpc6f2jAmtytMOGS2uLLI9dPykpcBAipEymjFdsf4GlRu+URP8cVE9+ct16E8E4UOoaZ
VJVeZYtO+CcXYQfF0pC+ijVDX92Vpm0aFpxsdi7owHw22Pe9Jkf5a6G9v+Q7F+3rjE8bcJKj1a0g
YnJdFgbXavK9aQRK27iJYZUTHKzb4eDN3SthS1TLMXncq4k86rgxvRVGkk4BRfcIjiF3ptbbRIW9
CKQCsOghci7SrX6a++uKaCwj94JIfoOfKMatZfYSzWg1eyrAAmTV8RbEcE3p6WLqcKa2KyIqxn8k
B3Q03QpTBE+as5IBi/rkBYJ6xlpLqA5RUTy/3eM6OteuCWReCx8uRMZyMeahqN6tmCIb0RU2S9Oi
XnmKvImx9uldKXZlT4CqWxnx6kzUfBNBGPc8hzZ7W7ggW3PZkIyOAl9Q0k7aTvRRr/RF9a/HE+La
/7jSvOM8cM5uDXgo5wOCN+QL0isxamq7evtb66m8TX1vYCku6rShsTiTUF3JY6L3Pd5C9mKqY+/5
FNrK7nAt59cCV0Ru+ojaYm+EF9fAVrLdj0YTpjWoeVuav0bjD6mQYV4NCErR7CwkxFnRoqNMRM2v
3yyKEj/kJK6An2llCXEuK07IkrzNwnpP7GgZhmMg+QCeYOyhcNg51D+Sop/i0bLuo3QC8AzpOom5
w/44OGWSomfVEW4HJIDYO9hpvYFmbGvTjjujF/arleUW9m3zD7h2n9wls/5SXKVJ424tfSeeMn1L
/PXwjl9Hs191+Wwm3ewUsc6aTCc8j02uuGF1ZJ8sKxlJlaZz+a5EdlRCwdHRLk4+2G3srqmdmMyB
r7YEbQMSUiBk7KgD6nYN7RdvHxPJfXreGFZAsjz8/UrDKxhXFHtLP84rUgXNrTibQsGQlOt7hjjS
sbfb+NHSR1nYFETYh0+KTQLz6AEPY1DZnr8Ud/J1iQq1vXH6nsbxCDN3c2U6z7qKLTFxnxeBsirh
U4Qk3n2BXAh3uCxLkVkKJC9ml65qdzqFalpjpMS9JeM+1M3zM6QG2Lx6MeFFEmza9IYQRHtS/xoI
Zegr98rjQ2elqTdUeaSl0E7R4ir4Rp+Y1V3TfqL50fnXWjqWZ/vxoIMM0VCsKrPpxp5s4NB6Dmqw
Pw/3W4wRShvwSX1NDLfUBedhreHT8S2HgTdUpYeVlKabEnKmm+Ox65I3MR32QyZYUN2sRGOjstVL
yautJFmHCl+LixRUhdR1C2waYTq7Qwc0qp65Ux5ZrZJGq8c9Zc1yLXGybs/2eTGJBp1XvbcbOsT3
rG3awe6CiaKU0Ni95s+HLWuhH88hMVpPRI7G+57MuI3th/OdsU9rxGjM0RpJc6IhLSfFFUGpUmnN
XNcEICcUbIdQL7oOQGtYkdKONgS0kdOwxPiPCYrPYRFPc1UQw29OdDUeXZgKq+8xEbS8GoJj3UcK
IfxiY333RaaSVl/46UssC89BKLexFXo08dDt8qwb0Oj5L/iOZ0AEzAbRklqkBuYU5/Mdh6CULI5V
hkfyJwOSehmZifo6QiL/K87S70rVHvdWEY+n8qu4ZYzWWckMNK62Df5IA0c3RrqBp0yHrWHHhCbf
5dGIIZn30q89Cs9jWQOkLZe61dHXIA3iQEX/i6Ino1HLtW4NfGWsa4tpQJQvVM/RV2iERxQhqZa0
67y/pY8g+wrBc33+LgXqyEnpikqZa+LLjKTsThPgShum/IsmznKkpyN6XWLwtCluP9c41BN07ZIN
QHHy3nYAqSyPVTp42AxDvDJNw51wXrIHhYBJkNd6Wm2Xrxdr8ql0TjRqM2bwwfcw0X3tVL0tOm8C
okx5VCzQYcrUh2KpRp5JlsNi5plTSYOb2UnhNOve8Cg61P2BgwTrMtGjHBAHPMsW5Mer7z76Xou4
vibvg7iagQiiFEVoBFrjAseDd/OzicE5mq5cf7uMyXR3+Z38Lq6w2JRoIhiHGUqJuxKNmMiHKlby
y/6cBTlTN1c/JqLlNIrqOHGO38/d11n6pjYfRKAVHZthUNJDGrTFOiBScEqqOss0Nyfy7Q+tyPPQ
Xv/L+C+WMaS+4EGUnuajhMzMSXPGFhQPhPoeoWHA8oxlsXptrfXDWTGL2rFTCn//vS6IN5YTF1X/
6lvL3t5v4x6Dx6OcB83SHZi6bSFrrOj6gnsikTH3l4gA3sNGAdSI9qwFZm9ynQskC9fpmoxl07+O
Xf4UUq0uXpulIC4CdyqKMqGXHooOgAssxThHn6WR2RMGnVo1nYJcsMcRYPeYWDVSYbJLU/406wAB
3FCEm95QtLJe/Tk1sqWdQ53ekVDY7C4FFT7GUrgkbLPXoFoDPIVlGwl0T0v2kXlJlOq8L5glzBdL
cm3VeW8U/Uk8TQ8IeufhKAURf7xYtYWdDFJAWGx4B3ZRNXnHp4mzMh9cb75wvb11C89nHw7NKgPe
lFeVqUkOckIvV5Bsp0z7aXHh049jP8OhlEkidGVUopXAPBVd2N+p4mICHm4JhB7kO+9ZkagDatiz
wGqR5CIseZ1SspGSnxG2lX4ZdMUBuRTSgoMGFP/KmQuW4XaSD3S2RNuO8xtZ60dOOcTJTrf34IHh
4X/le5tPtINqwoT8woruLEBfSWPsJdyjB+GzQjx5orqOQS/b7CY7Zz4WprpL3mwuvkRJES7S1F2u
B0QDv4VUk3ypTs8+OohedyhqTcttOSVXMzl7cRbjLOJwd7ZuhpSrEt2QDNoi74kIldctG8W/xBk7
p/MKde1BoRE//PedoV4MeEN8faDoHPotgAs6hQxi2tUZYPfESikXtdGRgi1IejJrFflcHVKXrLVC
mC3ZTIuEZ7tTh6HLFTAz9chaXn9DXyDHlQEqoveY4YJd8o5XZuhPYKGQKL5Cxgg4NsrqJ6f6NNoe
IA1DQECVAaiqetjZVLUKWU2QJ+9VEuEsBDBU2RZERLxLlrHVK+HAoDojwOkbQ2Bf158k7aI3J2OW
OykIIMU3qKlG9wjDAbtSXCE4dokaAE2KbNJmKtV1YajUYw0zPXhkujr5sdeJjX+s5BzMEY9UWJJ8
nLd/0jOgIkYjGq5H58OFZ8TdQopm93gMBKjjOwaZZBN3d0OgBH0aLcAjx3kl5QhlHpXrsl5p70wW
nZHIYNarlKO30GimvQrSEFCifAgZqahR39z6IvQgm2nmeXWPkdhZONNHv1PdF4Lt5tRz5WZR2PCE
g5yQwLNWJFfJkhQYqA11CVUEp+AeBi8MJ39b2/3Xtl/BlPzfMrB49MyHhZTHEX8bZG0cbp8dfaa2
nHopEIMZFm89RsakLijkGXgWgNkfNiK71YnTPufF3MO6AcRQZa9dPCeL2vCajSe6aUek6wr/tGR4
kXRKN5GH9UyIELvPqBon+Jkf42EwdvRDe+5thlQ8TJE2VUosyohpQrvcvzNbmN9duG0YKiyp6gil
TYWxJHuwjxGnuCIUOoZ1EDRoEUokqZp80Dokc8GRPnguAK/kbEfshPG8Ss8b0w9GX5tvEk33jXh5
dDsc7oVXw//BTHSd/bfVgH56Jf69NGY0IcqrrLP2Bx1594Y04Eo7G5JZxDoZNUKswdrH6Gy6X6kW
pPoIhrSoiEY3sjufCFbOwjZV/1YTK0g4Nrr4vdNlWVpD5BiApJz2QMRhP/qrRGy5xc31Sfy/92Cu
8H7ljjBQ1aIDRvRL+fCvbCPFo+uz2P53n4xqhsy5y15BG2lFlYdIlrXADP68O425nIuDxHdTXE+8
1sCzco2FN4ZwHrElVQbnjGXU7fbfYrt2v+J4bD+0FORAiE+jYjiMsMaaqqQuD75nvdaA47VlsU8V
GFfGRC8/7EoHYJgfI7XltAsPEoR1e2MXuqMHz9+fOLVvhKW+XD+xTBZRF93u9jQZ6kYrnjWjkB3x
BXGLNtu1RTVA69oQKPdFFPItmNWcFqLqymE72SOh4SYJUeimd1FkqzvdZZw+XcB2pn/pVCZvn8i7
Y71Ks2jeuS0/0Tuyb/fBOoE56aU8Cz7gzlQfXvqKNTs5LKC/JigCc7VVn7FcF+zLY4s6QqUFmLgc
UQNESFipvkoJjyfZQd39kc2izoloHcnlW0USBse/3gqVlcHItqezVcoyJtTwFhKGk4hTYXK08DXs
ijnsPL9fr2VqUEFetZwo7iEtCdYd+hqvvLXgXb2VwdHSAukPTkU28TLb3jqdRw/paBN8t/FFZOKU
EXzxOhTHf3w/eG4awCCXMg/SgUX9rGow8nBwYqPjEjhQeK1uVqfPETm/hcNgRtXXUgqD5gznznWD
qPMz4K6fyV7OJWifMU+0AntjuodkwWb7ULpLehznLBOyVFVNydVUJoNglZ46jKNjqLuSNRQeSVxB
U8inKbO3ZouTMhXD+V8bwxsAf6DccZcO57wRB0gfnlDn+GcSkw171PQHC8bXtUyiIZr0WrC+9buw
UL9A+GhiuTEfw6q9kvjdEbt6dw1ZurT2EytFDsNK8HdXjyQOdJQJYihqxEuUGjDpifDY8DSP9+I8
Xs5Q1RI7pIASM+raQK2Ru0pXJTvdjtMN3dO0/m8/JaCQ4av+j51OdGF3VFIXUW2YeCS9tD43WqMG
/UKfbQQ8cGUwaGZs1vKrY0nKwCEIvKeOMgJkaNmeeCki62eMSUkMXGQ/Ue6jfxNeYHT+oeZAgZpM
jd25Uex3T0C+VGLNjRf3VieQVac88DM1wN6D/tpD8XV/9BkQMcALbForkJplxnoVMGkiEU9CJyqV
/Je9I4+490BcZOM6j/wAxSbj4PVhoRw2ybzSQeZDgZfJmxXKJWqbaLTmFAHOrx15YqmYg4V/uWLr
EbIT08HuLd0XOVtYZpZlTx2w7WNOou00BjwE4hF4VySh+b2cG8cyeN2h1ykQZik8LDouHabuU560
FOpG0V1i0P+NTKEJpnOgEf3UonAOihcwtmQ+kInnOzkeFDspUIkishuXzn6m+VUf8aJ+s465avoZ
dS4k6sHVdC85F8KoZJQYQv/hbM0TWKgwTTLy2QmNIpJ6OrIzp/Dpq2/iK6aroFWPTQR73a4I0Ych
OJt0niyOKdSFTqQuar2nFmmOSqN+HEIecs3bNm5+N5COlY8cG2sFIBdy/kOXouTayWtZkq+3zKmU
SIUEMfUgF+ziN7rURzAz/Rkqr5xfx7EtuFx5vNjR/OU1rrFwIYeIQkixsw8/CbsWwsfJvFQpn1b2
6a3hUbSEbWYWfd75gVQ6RMhWZUICcqeD6U1mU3hN5Ztoja0unpqKhjuT51NPeUtp8zR1IhYbZ0MS
U89geLimJC8mDa/nsKXRz/L97G8ujMVetjHEMnPb6gq7wL0g+cdKZ3SzF/3X89p1mMA4EDXze9LR
dH6DqjmspQChOjjQjIJd5GAVYf28sSB8O4ieh7d+0afzEysOQSZMjaLApKkhUW0x57VWknx14/Bn
TLzUX+/31wVZl37667Cvo3tDFwX9rxoTPCC3IkVCj99Fusqu6qMsorTDpEoRp7fRrCDYUtefKeAm
RhPqntMp16Ak5ZwJ/xgF6koEamW2N8yvAEEmFKsFcg4igVbkBewnMogNMsY8qx3hXDjUPUiB3tUK
oS3DOczw5n0bRbHISXIs/WV2wNW4vFaaPtPs2C3ZqpUsdzQiQmkR/yURNmJEhegh0YhZ+wSWCgJx
RmSwj7CEC9j4p+XxPbc0FY8sfRgXCsKI9CEjFynEcJYO2uIkqYg49plLdF36TwU7U53oFXaY6BNl
AMA1PGsUFZfMil60VigUeCP44CktVEG3QXoX3QpcfFQf6255fGa7c7D30NH7Q5MLJbz0B8GeDUVd
u1E1mBbn+INbZeZCErohTVvTluMSXotU6Q5s/qcP8cAsBgAtH868RbqzMo7K0XGIN77+fxUpmTrx
kV5/rQJdEBrTM73LYqlposbivn6dQBNpuDC4Zmgc/nFHzxRy5m3H1y3zgvI2nSopZpogo9ZhOLIM
gDM9gLfEJ4dObGJlcr9uDNT8uri1UUp1qwJdhiRPmcMPAj2oZqFTkmHY7ztmiuGbdTEqR0tiH9RH
Fy7Dz6utfMIzqPDLPU62GWvLEtpuFlt4qSGfJp9TpgNRCHZdLXNYJQXva5x/0qGbW6RfnLy1jXw9
UjnnFdCdLA3ITD2oy8lPOyBEMMJBodn5k1khaKPlPN7OKBaf+MQrXlM71p4aega3fS+8sjQCR5pZ
fdLdVF0XNnKv9HnIhYgKLSoFDpbsTpb3LRChjheCMvRPBcYjMK8ZZLIFCvy+mUgaFIUF48mqA8kk
sKs9wB4AyV06rvBTAf9lBaakwIJHoGXwcz9qMIciHKn9CTTMTPmTanh1s3YXMVYTsMgkoyrMy1Wz
AvGZ5LWExtKjFSeT2oCK9w95WJSdiYuoOb0nFgKqfa+4JCEOWM76y0OT3V/VABJbNQXCo+eQkFJW
gxC9myv+vdBIJ8KPt1eW6thKLucoXalqWi2igbRbvxIy/e9nFgXXvA1PkqfG2OpBsW19Gl+fpPlT
q4XI5SPcI7lfXNi69Xob4PT76HyBcNq9Bq0KpjDovxXHv4CFhF0bGPYYqiEbc1S+Ui/qPhs3a3mk
W9OKH8gayp5hXHTTBgmfUqV2FCnkp2JNAWsxl90QcvdPG8bm5P5+VQFSKvWpy1sOiCIirur3r7xM
ywC2sg+9TL20PN2pXSjxgmMh1QUCly60eFm7UzEqC5Ycuqt5c8+Zb7/nu5tQQs19NgOqEbXw/1eB
0MxVUahwzUsg89gqJ68P2F5E1d9MYZGmDxN2EFF/+Yr1Dr8OF0ZhVv4QiLNnPwZFSIBEtxs48f6V
opxZvhX8l7ra6eVs0kEOY09B/ssnKITIptZjNfyyQDWrypVEliIyPP7AdyPbwctaxvmLDdLok+/7
S0+rTWMTSQk+n9Aftr1iZI8EOTrPP5XI7wR4695dAvqf1GqWa4EEhpmKgb96+xkgqgsVXDNwbAwY
t3cG150oyxsaTiGwiDbAWByNqfcldVGezlOmXdeZKFuI0niDLroBQqsNB7sa3Af7ayIgpQB9cS3a
MJqBd6wUGl1waFftMJvUCDu5BFyqFKjrhZVVLPmpFrqeZ8Rolw26RyUyZ40MLIDepTDaTWj4e95N
ZIn0FMEMiMKsbAaK1RlLcmuo23FKg9rCQxlY+AuOrsbJ9msXxbL4eWQ5Y1NvHMA4KBzi6MGQFnsL
NsfWCBPHDFgqBaCuJkSQ+R40s2wlloPL3VFGUQI8ta9BuW67+DNl5A0hLghMgOiIiDmY736C6d/h
419I/v1b+83lE17VpttameXcPnIiY9AYubeTayy4H7Jv1umYRADjMAsEUkG83JU1RtuRIbZVuNa8
Zaa/WNVfkabPxj9t4bzBORpO0LA27f9XkYz/LBowSXMqGLn2vmE9OLtoGGqY5o28JJrC5j8gxpcT
CujZ3cvMWvxhDpCsamtAlvWUphapvbZ/GnWpsb/EnBGhhD8/GOjVxCa9WYLsqLr5MSJ3fO9w0+jF
Qlmjhjs83ugEr8buTBPWGLBcCA97c+pgOjBNZ75YjcxPjtL3oXVJq/juYyr+MncInFVVt7uMqN57
irVHEQmkZn4Yooya1k6A/yltIaysWLtu190L7+dDL/imsfuLoKNcsVKqNQPgV7mZW2YD9+3RrSTE
3oF2EnZ9ZVwExE/ExVcEtR5dOFZzHEfyjrz0deicQ3QvtdBulB4aTrdtl0k5BnlLDPFqundIpKEG
YMAMqPkDrQ0aA9DePdlWjdB8NdpM3BloNEccsDpjfiq4p0a05uRfrPOgEmqnbQSeMN9jkvW+WCgw
MhCinH/Pk9aI1NJncA4IvEnp34a2YffDYqjPkjzqBDRQM4YThdmPg0DWZjBWPB0Bwru08pnvntUT
40nMIiPXlJYBcOKs4l50MOFbi+3ZRlalPpDsFaR1pLOeVHDSFgFzMQF/+YOloDiORmm2oaijVXDc
BUD8v3EaOX6yBLnl0ylgIriUKw3N1d0Ae7OBCKbyA+svX4o4zD4zmiyizUAJrbGOto8riX2+kwOT
xYXsSRtEr89dbOnqs+grMKQOQN9gNf59hu+8/QGwddweE0CjB0s9Rv9ZRp20cpQ4ct94eBmzgPee
833Gy3uyTY42W7bnpOHaRqTZv8BqBO7MV0ZbcHMFeN4w5HH1HJccVlwXmD20EOoFRupeQ7pQ5Q0k
1e+Nv58DWCvl/kfsABsqI4EpOiudSBAyK+GxrA/pAyiyT4j1f/wbQOnjREj/cMcPuFgi1xHFrgzE
6yYjQXsGNTfIcLfor8U0CgBwicSf2XqjGr24w2s+oQKFcZ2DK7oojBcmEuesa+LILuAk46U89agy
Y40CzWJcX+X84EcN1dqu35oS/Lb9i9qPQqAvKB4cJBC0naFZB9soD95o2L7+3eOebt4hesl5fhTn
rOsJpO+wKL/l+v/sS0NKoLXMgNUwRK6rDznL1Cnu7j6gSOke18+GfSdPzyb8ueQI++BvBu+KUXKj
U/H/G9iZ6CpHyi1z+ZN8suRULOPxZK436aMwZK+OcZn7Vf5Trq1u4SPP+oAs/+gEuhG7f6wzdxzS
ShjkNgJf+CAkF9N+saZs4VpibRs1TWAA1Z3FJ5S3YcPPQdc9mZTeiy2OuKBpTDDHEyeDR4rr+BPD
GmB513dp2C2fzGeFzA6wk4XBTVp6gmSHG3FkRwAOzMnQTad5zNR7uHoRBSM7jx2mWG/6/22Oa8y0
3DicQ2VHCb3bY6Gnl4pdAPbd77hEGoMae4I/Dbjuq14zaNhs1RmIhRQg2+rVP4Lh79HpJQ26mPZx
XOpM4/k4t80ptZArCF+8IkTATn3BCNJynZo2KFmnZgIwvwXxrmjkkqt1JzSBn/PL7uEbdUfoxAkk
mvGLqlmqbQBVhDUqZSD8vlI0d3gsOyCGqv/UHdo8v0x9ROT/6BhXYFuQNTXGPu0kITnXhsr5UdPN
pE5V0oPpioPPiK5t3/bvU4yygp03c+6VQQBriHmm9y/ZrHBqgP0FXWSwnKxqu/EW8CoC3XCspRy4
uGgcuaunAZAJILc2aPSnWEWrcuDGrCIvSK6C0S8yobnsxbVNTP/AiGONW6svwDBo93GbZMXCBsWM
oiylrVWbBRy3o1zBPqM4dX70uQk8mBgIyYQ4nCiBz7PYtbNLLUnZVYJEQH/jJo5VpiewMCi0xaTI
dVQ082zODnDphiLoLbcD5ej43b2XiTjrxwLoPAs9h/OCMia2vRHIdIW87kUreJKKvxQLQoND1PTZ
mqvuXQ77rKTHf87LWNkjR9Ie5ANKxbnaLwjA4LrxnfkA7jWmSyBE8L3q96pKRPGAcWl6Sj3yzk1T
DiUEBvGQ6wDCZsNNnLa6MSg5BDZREBWqLF0dtrIcTTJCmdmuP+mqD8PDgU3s3MRXRuGKcmN6K2Ge
JDdL2yh5UwLmgKGaHECiwr5z7UIR/63vllHz/oBE3IWpubhcmcOOPIwcgysnMjVFvK4cL5m1B/Ag
KsAXxsww5WOfr1pzmssIGVQon18kAEn5M7bfEN5G79A49N8Euv0Qqh1gXYUVJUnXPmiLoDNd6v6V
DPpnFS5IEFuQ1Skf6ElpVtnWPDfi2gGl1EO3QzL+ydpLw7r5PWtOasZw8PyornVpV7RbKNU3HnDG
kadiwipE/pzmzm8u6KsfNTefHckUsV9rhhgoe+cZS5HVycwTh7V0zhfMdBqVV0rgsxil22x5SGQa
AyNRM+Tl95AF3D1kBsMwhBfbKQGr55tWssJqZYhDXodOMVH6gKCDZT8/dsglPjYcRYrebOUeCipi
m+baIbATlK0aJIIa0CdJDnGHvOzbFy7DTo5G7L7IjnMB8/FqkM2/8oVQw/SafAwDZOxQ6rl6VTbO
r1W+lVQCl9uQ5PArp/QZJVDQuFirjwmzFO13Iy6b5M6lIFh36P5jQBvCHAZeQ7tbXJED2MhTwF/y
hHFlMLqhU/2V5iOCcty9GO6eWYQDMYUQ+3gjyEpISnNYa/MSsYpWKLV+DjpmpF6F7+ZAngmvbMic
7jWln70MiN8J7a/FBj8aDXnV4Po4V0uHn1kKHhpTS3SLImSY9jIg+i0batHlASmSgWYjW20DAY4E
Lb2orjfR/8T0lFq2lvZdU2FyvM/GzIxX42A4yv/440xlQLLh/nPuDvRh3S7WCXTdcHH8jp1YWzEi
4AmbMLkbJM9GxzA64iYNaCVqBoJJLZtyW6ziGB4iERmzP7zhLCVpxKKVa6XlIOnxiIaS74Ii6Wuc
Iy7/GlD4TvOVou/ZliD8D/dQ7R7jXWWWfA4nIPiNpXMy2BIsPjKURrM/iy5GJD7+sQJnhO+Dq4oO
agotMQ5RSI3ZlIh68aXcjfFx+hFi74S4vm2BxZDq9kEKmPFsVIufdlRWTIdCnzj+5ifq85rV0VNf
xqYR+JqqOlKibRuaOzUJpWGBa5S3Ka3FwEoI88IuDHN3qfHN9h1pwCHW9Xqh24w3l3kRY8psIkDD
VhDoSvyN+EQZflx+xUSvQ3JaY+pWuabg9BdBHB//9Y7W8Y2fXVEGX+p1TUaMmhZqd0gYKgrmm2DN
SftKdgvT2YyKgFKUMfUn/xlaCbUdBB+6NmOlj1L1qQD6C3cyDFXmi6M+ScyvUl+gyiVt3lkLqOb6
O+lcrZJ3rI8SQRwpeVrFHjuJ/WKjqCbdjlUCJU7FpJKrNqcRoIDS/3RjqcLWUmWzPVdfjDBx943Z
rf+wFmemyPiJlOky1D75ugiBLiYaqwSi+ZjA6UuKfUSa9YyHzrCFGRyeCr1+EeJZkvGyOhV/S0GT
Gx+zgRiKXta4mhVqQC7jsu+mELV7iqJlfEJD9OLHVO62gOy4OsrUXmKl3cmabZYtSiLUrglHlmpa
pdXc27LlUr7hlREx9PEDKzJEJ4j/9etjl9f7vOv3b31p49NXUkIpUFPId4rolgkxBQH8YzuhusPt
qX4NGeOia9C4cvMOH/wpPZjrslbgaaL1dAAubqI8ry0hrAhhtdNGD2WURCq0CILrGw0we9KcogvF
+WyKZccFoxxOsAoRHXoSIVnzOasOdWiGkbn35rkyHDZqEaIOFcv3tEXBk38SoiWf5hkDwtK948ys
kGSVdtFUr5IqNJTCWMLnDI9quapQXq2dqIVM1JqvxExA2mIANVJSNyjwExMkcvaCy6v++t9elx7T
csCGkb3zNeoZ4IYnM58yhXiatETG292oMrFBgh6rJpgD723C22ef0hAu9X/Upp8hExjKLbbCrUkR
NBFqgbRzRXPa4c62vGkUAKOX0wwYic/kNseZH8CSgsQRqmLncQeDXtthStMUB5lWCukL8owhaAMT
bGFT6sOykcO4CjNC57zC3DOP8fnmWX2RkZ9tVNq7SsOlMWXbRYja3+XAd4gkE0iNSmFdzsY022Fe
umEVKMh1RESTBR8UPNglcnW+XryWtDN4EvFhDpcJGoquOvzhkE3bs/fLgVu8OIk1dtwH78A4yWGK
AjXc3Evhp1hvHAjFQbzK2Qxe0OJCRDiaOP+W6FahjEO8v+eaOkL4qE8O5I7xGZIUo3wxXGmerVFy
gLM4NSY2wXluxiimDNpCyanG9EWIxSt2lXoSpT7hyyYbnv8Bhz8m/u96hLdLbr5B35wOr3AVO3TE
ru+rqt14pGZJeyaXkAbPm1y3vzqRPM2OlxQP4PRmF3kzSMtIqdSfNKkmEKwDnVsSc723xodDnJNN
kGOwBy4RrlQkmYth6jcmhcNO23CbWpPIio+MgO+5Lt9cmFfcsU96kqmak02VQ7w71pPkV6mMpj2R
pBvm0Rvm1/+WftQwbejWjXwbO74PUdsRgsLoX5bjcAaSlUCuDE4VuAVprDOCAvnJz4JVjEWry2qG
wYY3nD6HiVwDLGp11UAfO7lSV6NdQq7ISfbhdRGGaRjM7yZQ1dp4p4OAim4mt2s9D9qL8Nku5oWI
+32tGNb1tOxwRCGkjI/ixcs6Af34epKQwylPaDOdOysfA8SJQ1k2fltkNDlqIGvRQpVRR+FWUrzK
G13KdMt7iKOfLFugD4USm+WZIlmYaN6YShY0jf6VLo+GVo53WpImEM1XHnxDZZ3VRdBnie6ZYkzy
zelY8TXolDvxf49iUasEbIxpq5ZhBAb3MhpkVeYcfK+FETvKhrRmBcAWFLIpucKIbwigCuS0coTk
upnVV5xKpmXE3VC4EaeJiJuTVBr4+9X/zqY2Wr4Gf1ERFjOBBq4MX/btIQAMr7f+Q4rJB7CP86V5
fPNpdveRvFoaQXrStCuWkyAQbHSobseewwTwj/cKqJacdv9S3YC8xJtK1wsKmGw+lCB8Jq+dLzqN
clvOQBlqiGonUeNntphVITuTdYgyST40xbJvwBDVlYqJH5+vlA4PJO4dxJs8qx/CwNeqgF5rCo7x
KaIOpW/pN4t6qvL8d2MNXJ+HJ10LAomqFZTPg2bDCnA5jkrFlk0EvHhjtpvwdiP5RObuJjwjtqMD
fFo9NHip/q+n+xLs4BnigSKBO6iLDQ0FH8lra8OyOEWl2l9/HGGtRHfCWtq3fo1GxOBwpaZ49OKt
pMtjTbj7OrmLj+nB02nNm+OfJpzBlMPuKhYUfJrbm5ktWWrGcqB3g8PTTsl024s4dBI8yTZ8qILo
X0cscPuZOfGnWfKm9Syir1iQNOMdk5QvLIH1LkBklb9sZnUtYlFvhFkLFrsu201w8KWm/VllYsos
zSedRefdEZ8hOq2zz97sSGqyGM0XVNVgRBaNyxdzzu/lWXaq0MDaNyZevyResoShCl18d4K+Lv3a
9x+Zz9Wf9VyOyq+w73HB0Z2FlIZj3VuJvhsMOX5z9DM6SYmzv0nHNWjqLkD6kXYRWpfLQB8rE/pa
L5Bb5xVsC3Nmx3jPrZ+Sd0B2qEXdw9kLUO5Yl6iqVBW0/uovmW+ae41YDQT6D1QAMWrhvseikpnd
OZcrSbcnqSrmwQ5Zb1Ud5pQsOlEQslg8kTMo5PE9+bPsY3YdKqshDB29NCjHHHA1nSXrKr18w8Dz
La6cVi/UXZoGnWZPkmoJBI8UTzDpqmbYm9czqb+HWn93BBIzqXjKcouvlBTXxiftCsYg4a66M5EM
c2gZ0M2oi9na+IpMr3XHU0AkO9ma4/dZdTZv1Bkrqyb42VNkMVQISP/1ujLbOX9F0Fe7i9/URdUZ
YF2OkBJVriNbQWPj5x9dxJ1X0KBwxWA79xrNjI4EnE/HD8JXwEpyHziULTugbnIUbl1LcTAYRwkh
PdS1gO6DwfB2QdUe3mX4cG5tcEAdfYP3rfrcEyLmgrDXHehLbz1RC2weLyxzf+z1/vVjbF/ucvBb
WOcniCYYudJO+rol//gtHrZR/WxqR2lJjWw+zvrghw6tL5yBovG1zfyXBugtMGvDzyM0M7apsKs3
AseMJUE2mFgXFJW4uOLe0vJ/CFrk6baFcS8i0HbDYQRRD++aDztsH7brfNbtgKv6ANaX6bzpe1qy
W/NxpgaPfcc5pNVS9w+fkRZ0CtujoG7hbTOOFypdQyOBaC/LbwnaIGPWmfAiIp/Mgrs1YpUOp+v3
r2CeSTUVj+g4dk5vyArkVqiGzP0ShV65aKw1ji+bP0Wg8daadCAO0vcigGLEJwe4UleESBnGdY9Y
bBIRyh1TyfZqTBhUlLnNLIH5mHxv0j5Ck54VE33pYPjD2DbUVbhBlRkn/AmX9raoYwylOWmm8LU+
aia+Pifzwb5m1usItdkW+qZZeVacL9V6JvmYoFChLJDBT3h1yicIL2nDJ6ndH6vnaN7fGRrdzAb1
7nFZnPecSprKxnY8cGSTJ542ONVUJDSYwMUnMcHMTv0Q8kAO0z+PFa4HAcQRWSmMBZxhiysXUUzD
XUcDoYFei+gmJZar72mXhNYUiYfY2N+XnEKqaE0XTo76hCiVEmCHT0dHY2KRn85Gr3sSXMTmB8Sb
ccjcoFN89ChHMlOkWiFzIjr82KEAgH6tyVM0bDyxafJXMu5oorlZ0rmbt9u1siVUhqVcTkGVu4zA
2fvLCgZRfRowDFC33rP9uo8H/iGzluhoDnECITNP86Cy23UNEvF8I4TSUPdyCb3uWvswZsJqoc2I
wPgUmr0vhvZ9RtTR2SlRgfU1OoabybFcPuxQTaBYfHljyLuO2Vwq+NUIIzAjG+UPpvshokmgQsZD
pV+gkLwLADFc7WOUV9ZXnoeWH2Xy3tIedw64Z/mRfiKKJ3TSrKxDo9opgE1T8z+B8o1WT+YuvJ+k
ETyVur7VEUFM+G1avZB1n48l9p+WaTKaNAECNzALwIA0+O3VmiNjmRM4EPkudsxYOqpGOsxDUj3t
izAVSo9oYjnl8CmnHzEeoCdN0AdfnyAfick6KpibV1s9W2R1scq6nTI7X1ZZ1Agr4BjoXN68sYNp
MimcgF7rFeu1tgnsl5IHTog4OBBpBR7wfJnM+R/ORSEwizirbX6CswgcqJE+0rnSnpy/DS4UTm2f
baKnIwN5QF7ApVzYmWjZaZTsMtDUs7rOhaIelz1KfUhprQ1TNTNiuH1lG9FNW1XBJVznBgeHpiyv
NxaCgvY3gnme6GDJ0NKPPf4h31CfmbAtC4ImnjEPR7gP62dUEoEF/TA9TDGzMlbS5F/BiXjiSsKm
qtEQ5ZCQhfGPoczNkvTTbuilnJDf4V7rgbIdRpKpoKezNZxxfSGpaT6dTsYQYIULnKNximYIiFAx
+BAgdxIcuooF2ftJJNWqwvfM5eJ78dGZ8x9vzQWIZvpqaoXn7wcSimKRu+qR/GmSpb98ZJB7VuKF
SEZv7KRmgT4q7pBCGzZmTdkcDCI0V05TyOVKHzB1Pdwg2lzcMaCedLmSCHuww0na//sqPxVZfb2k
Is0VQZ3lQWs87GWQn2UxFLkfDkO8lbPzbikNN1aODUioHgRDY0fVOlwuZ6lb4kVohypaCrwveD+S
YHIwfmVTw1yAW7TxlFk5F008iv6wJRHVo3ibZkpmARVYLAzON6aVyn7jV5SGyqJrgEQyBVQTu4hG
Kte7NQqHFvxOiLa0MBDTlfxCmon+nxVqe3iKQ2C7mAwakWkTIMJzKoxFxbPMIZ8MMXBcAM1pLGyQ
Dm1ec6BlIJVMlkIUYl3fB+Eb327wHB0TueVmVAi3Gyc0SKb76HoxRNtohjxFbI3hByu6KD6WkUx0
Zoko3EIFBU3nbVB1dnJwA5gt9hQgLMd3zh6EEywo6AjaopCwKeYCvxV18BkRAuTf6vaM0nneW969
QRlIi/G7WcK9cs6oefE4Yi873QFOL5RrZr/sKJvTQAyBFAlrh/b/EFDdScx33gUFIMW+bEddWKB0
RWZISgnRqd62GZGMJchVL8Q6JZEKcBylaCNDlH4MZLNkitUFhToWBaLBBfks4YU+jAK1qJpbc5Vs
Yl8dNLqbzE0E49TkCremao2jHxvVVknJiZFFT/j041IkzuXXGVDMUuFrqwbi8DjSLzYP8odHMTVq
q4ZaaomoY6svvthUrSbQTKsjRCbNW4XBPJqeCV2Pb5dZckeZdxu5YsdVmYZKKfmsE1Nj+MJ8TzGt
Rrov2qiTCtOA0r2MBhnVCbl6BSoIVKCPeCqQEvzUie73Qh0PVsdkw5bDpyxkye1CK1DttdZpv6H3
gxiiYa4rjV39GKSiE01qNhUQlaLeGfn6cqqJyzuWQGhC8aZlkSN9vKq5ftUe3kSCzEvKhESwXrKI
BbSufdVj1tg8XWHU3Hz2t72U1dc0Zhyn4V/UrNJYc+gej4b8U4h22gTacFZRciQnIeZ9OpngtfJw
8fdVlC6PPFEBKuCx2rNtgQs5EcT26tMH7+VBvzE2MtYiHB22XCJnOfk4rXdSXWNu0KBV1S39dJYu
yaMY28OxYylII73KH9knKJtU0I4MmUHhQu9vYvqLzJ4OZdLIEDgtnxklI8RI6c8QpawRYy6k+5or
+stPy7iBFPRxjGHX+bPEZTZuUjrxV2Snd7gBvMkC0EWQJPj6qQZH/XLzYveSbXFfHjUivoFwMmtT
GypgDCBTXDV8I89R+Gwa1odFiLHNWS2jXMo9EDqUfl1tBt9T202vhmU9JP5KxWtGbjR9Tzx41S5G
+ANrJBJulGQPJ6J4343DKkU7chANBKLmbgkcxfseNU4DoqllF9fGCXARANgxPGamAJBRzCEcdJNM
HurNODRB45aMshitXE1Y98DONrSoGLEvK7IX699143Pn7u7COjyyJy3Ow4abC0WdeF9Xx/gRWv0e
94otoclsdO1NK2MXGxwpY7W5fWMXfcDsyl2Gg47gcePwJBCDyM34hSa/lNlajZq1e+sIGeTtQugx
QkgFVsxZMu99QNwd2L8denSuISlun673MMrKHKEi5zZtO8QySIOL0AaGVkKlEoVCXAoN3+/UxZpy
tCjlikUn62AVhq0ZOLwqP0Le1EQBjEgb+y2x0ttKja3cwPrJ/nuER2lE0f5j7l605/Q/JKsMKs/y
XqyxaTGRavn843Z9na2jgFyAnjWioULtsQ+hzlfF/102USEYnvF2Ppw54j4gacz/ZpkzGqI5aODj
CRzprZ7E6P9z64vXDByeio3RxPfrFhfgCLGxHSTvfdJWraPBOSnwwmPOPsi+Gc0MepIyVwIRo8MS
rEvVNTzCUDDh5NF4T+oIO+Sliozp8Wrr+nAHbL93IdryDXjZa+912A0dtsK8q8fgtN3widvLwvij
TDfZ9HTWqVHwnqmw2/FpBLxxCa+sD/ESB1spBne0RcCLNWB6S+c7vF/09GUmQituOs7bw+EBLcS8
ZlUf5+9mw5DSew7iz2LCnwHPHraLb34W5Y5u5SvaD3eBMHAmsinrIMGugQaUNbTAvPkm+dO7f4zF
BFiwPo9P3rNpZYoC7FfGUQB3zAnJ7uc7VD7lAe+yXssQWRZM5sZ9gpM9WKUULv0CoVEcgEXks8oZ
PMIDajPbOJlo1Ap8AoPOlXjKKPXAtjSn2tjvhDV/jMI10U/G0vJU0qbAd7Fox3YPSVk1YU8aozwc
djcjN01kyWwawmG+HUNlkg01gXNqifsPJ3WEmpN77f0y0t9S8Mp6zrd8fbJVLmOUE48imP3MUACR
kFbJ4cK4RNdsaFYf1ensCBpG1TIIC/j4RfYaaFLiafzgloBrgBZebLDGi8CLHkw5JdX5fcFGrf/Z
E2g5ZzoXCjTVK8mslv+x5p532IaJgO2hSVE06ITH8+8F0Hkibi8kgBy/CxnpCVb2c2phtQagHE+N
CKwPn7i2m62SP285CcDS4u4lVD1cbPCBgdHl0WRbNA9az32SxVcOU+Q2NMWTu/VR9EQ71VqhuggK
Rb27nd6tnx+Zfdn4yaLMbL5L2ILyMD83XSdp4un3bdaq2TJrSG5kX2rnubYw8Vme6cp24k7LYj/t
+Ee2nAaLtwQxpO5NcTaQxpc7OxSWTNfnIwfw/yLkxQxefkjXqqKI4tmUsQJThnZvnYtzWwjLkbrK
aEs1qmMxg5hEUZAc60ZUKZaAh/1wNB2rFHJVKbdiWBynzA0Rnk4q5XqnvibIj6s4SjUYJ+ae9y1t
bgCK5Hl6pSsXsEUoRcY30H4HlNO0UF7xFU1cVjv4h015tlmwhzO+Od+j1PkrLH19/BEIBvcXzOF1
YsdaXG0jpFtQH6OpcgOfvZ3awJOIcKwGDVi7h7Zti5Dc4HAvKG2XsD8NFgeM1eCbC5TS2zp3tfsl
jDbPPGE1hbEhVe3eIdrMQQ3j0npFzhrSIh0vJA8L8fM6xU00Qs3C95k4tGJJUXqkdNi5QmCQWkIM
qaXfAKBH4kIgJoC8wDv5YVsq70RQVi8qwAtBvOFugncFZNQh1a1ieSlE5Ez587c5CLUKqoKI6FKL
M+wH9c6m7b7nJL0rmrdzSSFdr64IDv26lkQLB6V6YhCOtJnG8qjl9ylD+Sb0zXlN3hiH8veramPu
Wo14Rqtc5IH1SBfqEAcGWDgrk+jk/fQUZEfrRMBXoyGqgqpOCpFiaXBOA5t/sfHeRGVChBCqaxbh
8Nkc9kKt60MsIJXYIfH0zGZtByYjDgKL+jWFzItFqw5AwVngvgy2k0NL/hGgYiCzAN49XX5p0p0O
jU19NcFRFKDHUyQwuHNg3XOgpB5Nx/NY5FUXL7+/U4WF3WTzu458O28X35Z9hfLqFTYlqFG2iXJg
jwUxRzXKRxD7SmGkaGbG3xO0pfaBC7zH5zhELOZ31Dcq+FJ3MCzsbFKJXO+JGmYgRMU9X6fgrJ6s
WGKdPXyxPhojBgQAxRnW0B4dwxVog18ivhYNeLw3BXwGkUxIFz8x3VcG6hxSSBTTJnLc5bnBIkMk
HwShhnkk91OKersFqnJt5xEuPbh3MAhJLCQp2uO7Is9kDfY7H1Ec8HoxEhq+Sd15x7FZ5gd/RSAQ
kZrXE9rQHh/Vmuoh36oPWfKrRPcY4je18+sE49ELTTw1OaiVGNUYP/bAP/1sUGgJlWhdYu98nXvZ
OiHSl4V62S5BvhNAFODbGnYFsa8oORht8GpR33OiiveWoTPh8kDeP0YtsRQMwBXmIo0dj5T0UCBN
DdCQflDTeT5+era06FBGiPl1iWkMDoLQrYv5PqJuAKbJT+VKTs2OQrt2U3bNLKM7Sr9JPeEc8yTE
XI8WiHw3AbWtUEO7bYlRve5dgj7h9sVniF4XLDuZIGFPPoyvkpNJk6/MEx0C6oC9LNJiHz75OJH6
b8ZYKpYwYmGprmhrrDrMkt6PEa/HPOeUVmv+CU/TkgxRWnf1/+hrMdKFMndhP0+8gLIaRYzEOipN
R34LomDCFHOSfSW4YR+0J5AVbHP/j0PbwHB/eHSTxANSGoC/tHzAc87YEJ460LAGj6rVj8pBGgo2
HGu4hFtU/YhZV6fT0HZejzSFINEg30tBZ/RW0zBeus/HDMnca7K0tt2c/1MlJqly4ApVSwy7DdGb
hrV7863zSBWVoZTY1mZYvMpfGX6b0x0xWmu7RyIppOTcBK2Q3crmENBKXIgOcCh51IBbRFRH6sBp
B3UFzfGofEXmUg48l3YFs+P0AYaHeS4YW9SvtiNkvFxn9t1390hffybloeaNuo5PZ3MfQonacimU
sucyYJhdO4GQ0ONN8w6+sVD5UqaleRyuSwtVp7RjppXuwYIt1GonzUSnS+fHtzvkOwVFxNSdJ1Ur
vKeq/SZk+4HSRPg1wgs5I1dju5JH0XghSdsLXnvWDPBUIxfcX9DwH/4JATYKqu+BItb6A0kWRriD
tpnwjr7UGAM0VxddrW1nMLVN3nxhUU52F5X+BFGGm1VTZa2t0vb7RnTQpk5OCyG4gI0Ra006J/dO
vV5Ww2HdBtzbiGsSdqS0MQbzzBaU3mxzLQYyzRwkKe1gg6ZApf80sfaSXw8bfNb7gVWoJvmG35UD
cIiA9UEqz+tzHXxM3Fjs1qTlZuD8B3/YuhGf7kwRPjIc6krF23kv83hnnG8/VJMc0aT+oPyx4aWp
hWPc6J02GHaq6vQRjWjjxqm9OzRC2Jf96o7eGqSEmWjgvLs22k6BCxRxP0Fcos5NxemsD1vSpnhX
qI9HIaj9k/hX53nunecYcZ+hJZVqwFpDeNKdN0rj36jEmF//cD7hjdgnPvqO0cNfRBMTurbkD8UR
prQCcpHU39laKsj2ZXqQPP+q0abXWxjLHXZeD0M0yJN9brf5wOcaaDL2kiAca33T9VWvTvZ5Pbo9
u2hXII7vHkraxEPJx3mYKioaKt0b7LxxVgpQRNfyXcAfzqckXWAZJKE2HBM1LjnQIAbnr//S7HRa
SCQ+/zspGSnOVVr4fwk5ETnIH9yzcFgPxk6aTK9ZP3KD/B/ztHMw2762kXlgynKH0vy02D4uI9Dy
ouCYBtkaFbGXKTetGSr1XTzibdqNsgbgmMBkZBRo3xerwmZkfC48drJ4TtRTP4KvO8RWx1xNyCUe
P3ZcgzjgMDtSiIugnwlA359kYs4QA6nbMcNEfZCYlIcNQxIIzYSFVVmPNLTw3DWyY/d+4CXYa9AD
kAXTWdfnPQtWAEZ+hlX4pqCfbFthYaImvs/LM5RnwSDjWQ3eAX+1ITh8YyY9cafjXv7OqYQ/VMIh
s7spotfMEUPIZN1yMs1FzEldHDJAC8ntJFqq7aoiEyTWCuHtZg/7IEMxqtEUfXb99D52YCMXPmSn
HvZWtSs3KKTtVz83+CSpJJhOVdMy+pcLSfqMMNL61iY0ev3uwUxhsvcO03amKGCgMgcd0MMv3TzU
K/fSTncBYNLqHqD2FKQm+4yFtjOhr8IPARqqyonD9iofWUaUGtfbvoITYK3zuHaarr9ebadd6/9v
HU7WmyZhwQggUD5Il34bLbZmlTOyjWLVfAJgi6jJjEYz8XsvpNpbDd0GgmLf1HjDjpJhXRmSO8q0
jRU15Z4eCCFu6UfYoym0Q7WIIkrYxhe7QcqxBRkEfTEcYveZy0/x5Li2LsUcPYmF77l3yJY7Fhrz
Laj/gs56eYuokTZoou4D1KqKYFDWDCNqH4OUl9r4QhhCvOGdiPLogpRIqnVIe/EpNvNxgWmjrpTX
9QgoOVOcg7y4ErO6TM5Tl8u/dHY+8M/lPLdy0tE2ObTDIcaH9o+9p6Rw+y5AfPc8LGkc4jvummUS
Q3k2WIjeiavdwZAVVsUvCz7jmHTShhvD95UCJdNyzNGU8pgrXqIi17x4gHlI+TdxcUtm6uK/kG40
+b/xXSfed0Eh5yrdmey1iAZgbxU+536uX4/8OGfT/fZLgE+AQGyJjw02iBL5DD9zrNZGXlAdQE2m
2/zXxJRHsiQ9bgDtr4fw2fOWm7KJP/cgZ3Wi2lK2m1j389xPSu3VcGrhLavQALTh5i/k3LscUjHS
4qHTMChPs9031BRbD8CTEzOmwqtC5sgaTg1cQpXLGcxaph69VAUqYAWluVCc6tSEJNnulvnb+0At
L3cQsFmMQY1aczebvtkNH72nYISHRONJA0C3TOoaWZFduqx10uxfL1CJWV6Ujh67PS5k46fDrY+C
Ii5flwSP0AKQIq/auHM8VNCl1KD+fOdZmOnq4S1szSM9lN/CLv6a6fTRzyAteO8zlVrVKRdlihU5
Yfowzj8hLvYcGjfb6WWfWRnXo/0/2xL/pxrYs7Q+kH2owAV+hSUlNy5yA6kyNpJfehLTxJ3Z+kVd
FXxoyRHOhfJPZFvMtkdOefAQ6iZnItDQT3TSsRiEL5GzMZ6aScH/mfQwRjx5UvEOsjQM2Mwz60H2
EKIq1aChOxPNt0u7XNvDb5inhsIuNJegrJD7lrzRhTcIMrOV6Fyvf6WADnV06ERqNSkVmqcGL9oa
z34qkwHdJB05gyMI/vTFu4YsvBsg5gxKzE5ahk/FpPfKWhILM3OWOVkPZknYW5Ele4sriRB/+NIh
upCjeMxnJ4ltSgogECYMtchP6OlTNf0Dxg6TW5pHjSPELI/mGL6ZPk585Xb30Hebyn5kfZj/wSUY
RtR8xX9fh/llad3xbTuje1cnhC9+68KuLPivq4/SOxmmQ0KQRh+uWbcLafiAnfL+Nug6dPs5nkHB
E6bCnDN+TpoM4CT/1dNQDMSMDCwpZoUEPnWBSQLGCZGvdoGvsLSt04JDvXGbQCCIta+SyCHK7JQD
F3PnaIcpHw6K4daq9O9KG83TT9vDqp++SsPmn5pZu+YFbxDFUR8KsujihQqokqiiPk6ckL8EeqPF
kxhlG9M/fx1ui7UbsGpQuqq0/pWjvc//wtfEZ1xVvuPwLuuq/d9z1uTM3LqaJoAGrjapEHGDnQ3W
KsSdTCAHJoCg0UdIq4Q4l3pKFZ0Cmau+UkQKO+lOJZXOHmHmsonpOmWberbEoQ+iT5fHmigYnEWK
KIdgEUd5+xBr2uRfLCk4MRWbn3AUxtbr60Qd2otFc39QJOXvZAy0o6awdDmdJ3bVVX2QBJtj99L1
WtRMc5hFHmj1uCsartIR0oehImWncuUHLx2Wh03q6sSd0iJ+GSiqISbzqs/9xboHA4LtC4A/Fjet
QZB0M+5rehXmD/5cZ2pxJUAIDnXyV7fQa4FJnx0TJvpZr1tn6WcxLP1dg8xuntsT628QJ5UGzSnS
Hs/XUPgiA9s7Kc8w4SKHXXI0Fr8lO2tTdkEw5yNfYaL4kE/qyl0WkyaBQ574CwuD6Lp3CcpR3qCA
yhLIM4hHoWXuME9+b9AR99hMKdgFSdO924+AC4cBYUkkv+kXdS1hyPQoue4mC+SviAgPXJA7xO64
mOGxLefpqXnZ9UliwCqbtxJJLhnR6UXRBiD7sKjIc62x4Qfp6Ka9WzZdSaDCWXfQ3GxPHdGkvk1Z
eWFZ04YFC2fpVCupcGBzWG9JZiTevCXQ75aepHWqjhoqE2JoNB8ws+tNf+vsAgx8ukygW3TYl4oE
wlYQmGavPbiM/vQucaRWHB5WhMrO9T4BnEAVohv5MZshTpSjqNFon3DJ98kiHPk0xgw8ZfvRaELb
sh2A4ZEVUEJyCEfNFcaNvLm0O7fVaww5qovQvkmarjshUXD02HSw6HTkk1tsohTXJXXYx1scSb9R
fAhM/Laz/ZNylWk2XYxqSgmi6kUwffxEfDHjbbIgka5ZyskgK7SBdkxCEvr7W++Y5jRF1Bl/gl9Q
Wnyo96iHo10iejd/wTexRfjfTxdoKHjZxwCngWF2xxlpsenm42NR+FtkCoU0k8qaZKMoriYj7GNb
PlnlSf5WE1R9T2ie3TMk3mbtmTFTBQQl3RqM3yg6BrcdsivXiyL4/Xhfq72rb37h1CG1++0DkTVA
jedSupZlpELt6bux4Vky52noH1wrIkSkba0vmIM9Ho3fm6BopAYLu7oBBv4NtfRJAIGkeYNtU+fu
TSJ9+0EFEYmPybENdFIWSQ6w3EXx0wWKCloGxNxJaW6wgN5rlJaV3GL5HIIJIlWq4bF+ndoA7dC1
EN5Q+VKj7G838O+Pq3BFPv9I9bHQRCi+TSHpTPn3eGMcExDxhbcu2I5QbmVyZRRapFa3kZJyKi19
ebb2UuwdVLkrkLAcF808uf1y1v0z/N2cIY8JeZdb93r7TBKJOe0i74WSi/EuV2/vWydIJJX4QweY
UUIBeYd+aHVjDIyy9/KuyTFAMX+S9dhZjmiLGsuhYUI3bq237SxKF0eo0bw3QfMkMYf5rJoZOuTq
2JOxEEZLRDKMjDgWFrM7jrubdyoY/DPfpSRC+lcmIzmCtAA99MYr9g8Uy+RIZTEl0a/qbYxkQwYQ
enX4o+hdzVh5XJbYZY6tgvEkN+qFUMFLV9elv9EmrQYZDoaidQHyOt2WXxDkY7qXxNXZPqcrG8Ln
Pc5cG55z01WquM3FVZ/sQ5CMoiQBTZgjq+sBTSihamWELtPW1/MY8g+sDebU9c36aGbv/l5G9A5E
Jx4CiWywUUwotY0QYFZVDaLwO7NF52I8YkQT+2iBA86dtnILG8C+8CJfnGOqV06cIGiKn/4lgcPm
CGyIeSECNA+BKJ3Dq6wybmrsf0V4qvdX83nnTBVrcOInpbct5xHcxkfWLUR6yoS0xEffR8Ysj7c6
cDqLJCJ/fYqZE3YWVO0Ndn1Pasw4MLCIMQOf/KYiwu61cwPj2UgEQrE3sS/cT/0KH8aiKybV0xb6
haByJeL/jozn15sdZYznp2+03ZdxJTJeRw2BlPloCGBkc0QuwFVug/prGPzQOdMaKUTiRJ4hBK1y
JWm/WyxIRblp+W38aRFi7rZdyCn1s012BiUYe3KvtZX3yPeIi201M6M9i9Kg2fVqyELk/gCnXB1p
CJsjCP5npagOiHu/1miJHcmzH8VO4zWTknYs8d8wVyLYdTpDp9nEsJwolhjjObNytc1GzRhNLiJo
64C2HK4Xp5kjSm1fQER/zEMCWc3H/bJKEddrx2RnIs/M0AOwwPTbLbM7Y0LkDlZvCPAtBWs6zwtm
3e+O7/hwXl3Cp0FvCGgIrKKdG/96hwyWxkbooRHeZ7q6mwtAKQGNFNmce2YmugfoIu47Qa5Aw6iT
jnYGHXqTkYefHKxE0Stwqt35a2tOxhqb8aM/KpPvLCxHUB4ZBzTd6lmi0vYVkuSSqew1PC1ELMYL
wMH5YV7lO35Xy+Y06vWAgLstGiz4fTlEhtUUHWKmSlDJgFYJFl9I+JD9QNFH1bXVmfJMEoLl4DJg
EeZ0L6baZwOQwFAmFSwQrbMac6Ldz7qwMe+84SC5qpAKZzwvVBdaKJv80zkFUdMwteCvtcJY8Pqs
YnJHZFlHs9AypeEyMUzey3XqHfMcAcTMTnh4v9p2UmJdPQBUZN0D68W3H9Qd/F2CkAn9h9CZAfzX
6XPpDpM6PrNIWJahUYsHbYLfQ7UJiKOniSsWl/Yt06D0cD+U67KAzD78mZSpQOR3gb9VFvmOtGca
HiGRj2MQyni/1JHV6SHBcb9fNUuE+PaTAqic9zTg2evwxUskauBiDLiHkEq4uas4+LQRY104+nWk
J+llHd+vUHVlIeV8GHUBuf42nZgwCUuC/cGVez1z4Bl6hT1xTQ+AMvghao48UiNNsYTREHlYUCIs
CoA4oy+FVlDqD63WUdKtDWJUWsZv2MxS8Ka8geHqezaq3flibGVOzo3P5v3XXIDm1UNyk0nMH6cH
8V+N3umW+biqXdCVo/xpP9yVjUDBcBzL7WzUSC+zGO7Ocj3X/CrGYIqRzKcSBMcIRWPvzhTFzqsk
1wLekw5FnqBgtqYBibn2pJPD1Ux4lIpzeO+DeYMyl+/GperOO3pffDxP3WJoTsH5zfAHzCmPmSCL
RypHJMrJXAn/ufSdl/ephNMoEioHEP+miEK6invFvkK9+tKF8sVEy3Yg9A8MturEGPBb+danvEZR
gXSf0AM/8+9xKWe6DdyxWWy6nQRKfPIElks5/dE+Z/oMNn8Okru8KqRhH+81XNgZKMvhahj9RSTy
k3rsSlVRlDlIrOIGu1KQTi/GC8T4MM0zkRIJ6XyHRUs5i+Vl9AgR12a0Q5q0uqX1POkb4FlYnQ8C
wK5kPYFSbxDmFRcgjDjJJqEG+0BXCEgzJk0z6mBICmPZBxGp4RD472mcm4UICfxN1WDS9B7OGGG2
XCi54dMTc2XoOuVoa+aQjf9R4Wpvl4v7dL1age7ChiFYzzF4AGKB9KYsY6CKpG97blR7bYpoQRG4
qJ1ZeXDDdaJ8kl6txwPOQzNwXVEI4dd3Qh2ixZrpaHLkjEo/phKgA42UtbWzfTAjeygLikqC/Af6
JxaCIN9jlbRodXpqQBPOmy0WVuY7G1WXN0Jcw4am1yEFpDyHoyNY/7o5+ZfaA3Mm3U8mupz6659o
fKo/czzJoxJ5RVGe9Ig1fNHzCKkTsb0Gal+eHMXXvSD8NAfI84FFHCZaHp00q3gqmL1OJTE9W5dh
VLU7SCfMJTvvScc1TfDjGpZOIEw9k7mTdKuv7xKGrzafVjxV/tNQUOMTnvB/i48bhi3/uA8F12UF
Cl3En1c7rVb5IZnJJoE+dbVPMxBZJNGOJFCP96A3cDhvgcc+arCmVfxvztbmyBbqpkesVFSIHp0F
VPeK4PxbJL5Fj7Jb6ZDT6KFEU671/GNy4Nopja+ZOL3x8H0dRcQoriceIwtgbo5+NrgCM+mL/+0r
4Y8nDYu1xFusiHiqMKV8lBtvMOUK689aqbK90j4AzS6OJEjM9VNdPOOGBydVFgRVmVQX2AZB58XK
11XjgZXcPZRuxxJVGpBfFQm71vmf1EXjvVZO3tsmis64mVmYlY7sZvY/yU3BTW89oMV7EPk0DdkC
CzWl+y5NsEuay7gzP6ALJKK6q8R4FIS1F9UzSVZfxxUttcdIZ1ajR+jsq5+jemlaIYGIO74YlsTm
TwXO9BaXxK4QEAkBixKrZ7/enO9WyhYRbLX+3nh3fztMt2wabN9o2pogwDLIQ19nO02seWnCeTFo
KxB4+73sM60RNFp2cqrcGz9JB3GGj61/BpUAa2/bTFIKL89yAvdBs2XMqNlE8nYjpndS1Ee6in3X
XaefkevH33paagN4rpKAcXkdO/9x1FFwCYDaXjkVS7tN9a89btkYDVMDEsS8BGmVVH3kQoXjw/ta
h7LXuQsMhPqJtLk4jH/7Rn1uXDoFKOHNPFNeggCAxtcIghpaLaVBlkzFS5R207qWrO5UeaopxNxx
DvDS9DnMB3+d30uInNDbrI9C4f2ShmZ1/ZFMekZ2V9D9AlztRUDGuV5sga0SdrFtcwIyoqH72niW
c8ItsS3aD9DKHEFe3ioeEyRn27X4iaGC/ywj0jcsAhIndinNXEwMyAj+IRwKATULCmUXL25tk86i
RIHJcxQMFNWaTKOTmM+TPR8qrV98Sz/cE0CglZuWpHwmOXhChBbQKG/kXptnbqUVQnl1lXK50fEU
Zg2aos8HphpSAEehSGY6T4p+1MlT7owSPgWIa5DUG+5vTg62FKYZCQ9zXrwFthbGKEZxSRPIZQ+j
mlt7aoVUa88AZf1X9Nds2F9duJpQXSOuKPT7uSsvQJUOJUm4WeP45cHX6R8TWwprnKj9GveYRvoj
vmMG0fiH7RwKysuV7HERsHL7+u8LEeRAeuKxz1fr1Okyjupgo78Ei1ICuX2VTLx0WajARDQ1L0AX
F2DSYTFzj4Gij2gSNBr9rwPlBGx8l5d0lyU2Yg3VauYmuYmSvaKvpwlYHTo3V0LLQGLbsKkJ5eEo
pOPjotepcuzj1XWMbM8LAfbJa73fDvwMhlILQqPowy0UzOIuWY/mB64s1XmwTT/4K9IW2oVV1RDC
ShhdJO154n0q088zPbHQP8MKqp1Uo8EfezQH7/6njrrezc88YK+nRTY/lx2nf7kt4jejUit3qSUv
8QHr44KfT8iDzcLvmFzgzsYUQCHSDMqElEMk6rs4jt+lMx4F0xU3tG6ShcuzV0qSA+V7towzIxOH
srLIlmkREaykqVcnFtX/NrBMu0h0GEltoM5cVO9VvOnryLMoXd8fWWS6Yw2cKQkswEOMHbN08a0q
TWBvBq1OtNy8Uu3NSBdTvYNojyEEaCveq9Jc05LSEM4hIGGwgVgISFZV2LxgkBfoTWZMASpm8nmx
4/PylI9dJRMqsBNpX0pty5bht6lEUQr8rqC5GfNXXGe8YwFzKZVQtw7AXKabciwlpHKuauisGice
mytVXl1zkL365dVnrrtP4tFmNgkvQcv+4+ryWMoPJ/zHMy84GUofgTNo/AE1iXJRd9BuGiLboE/m
YmA38xv9nIPBz0yWbh4D/IGv/1A8DV9K7Uh2gXVM6uxLcayFmi8ljBT+xoUq4mhdtHre79OwlPuQ
zxJqOEAeLsMPgdZuvyaI8nW6qcI0pSM06QPn8YaLsdYtUFW4fE5OtPT/d6jLSw+ZkozZGBV982M+
J5bbJ2nghbi/VgH6SP1zSXC6b1D1z+D5zZNz8ugIqccC3tPrCx6158QlLKADaNRBYwdYSRlUW5NA
VThi8Jmg2wRv2gV37WGVtxAf9KBqObfBRGyO8Vi17TxLHZh+MB3um++TevxzddbtHAjpOqD/Q7gf
dvcSm1PPgpMRkOyalBAPQ73Qtwq/QCerVoJM4KfjINRZ9bh1R10lKHFzH+WeZrOwK2UBAz+i4+/a
edZnwdnrAyOoTmKKEwSaQrCY0PzQ2gRVJdfz9mHvDjWUMRLCGakZwUoWGMsji+rv2kgPGLOYY5vF
MNWlz5omq2y816mTz5hxCu5JVoUbILemeLy9XIKUX6+d+E9XX3G+bxvwirER1W7K6GW003W4nFVj
zcJSLB9WHEgpbwT8plvmlgShwezbiobYV7ma77azG4ottrOs8zGEKJAyfVvGhoLaNVfFd5N7vlJR
gWi2RCAf2H6s0WddUXqJUrwOFG6F7GKxvak1mz/gydQuGFmkUGlTj3wP9qRSKxuY2cLLJsMlC+7G
ZLiiP3hl+eyTdhZSlwmfrc0WkDrr79kHmcjyf17O7Yqt/yGtBJr2hFG2q0AWLFZce2lJw05oqJ8N
jmOOOFe0cZvxelrOvhanJZpKaV4aYh9ishnQGH1NAJMypQVODfM+o1Inkq0S+zsYZV9XZKtu4SUN
+Wog7oDs9KyGeLseHDIC3zbWJIWE9PBBFfd88L1qHJ4TNWEGPqi37cu4aSf9JsB6xPf4DyeqWhEh
cXgKiqpqfPkwB3CArhb7QGWOpCUipj354is0erme9973c+QXQHszbG7+H1S6Xu/7KvF01/HLriKA
GgEjxMAYvZCh4CK5bye8irmK4UXJCn+WegTP5UrCvybcysAj8QXEeZxsO4ZnG2rGYQWsAEmCPNv6
IrjMHlv5ETz7AURip/1u9YNaxrC8KAniiGWSiMOC5eRNJYOQFacASnVBgNvjikleZ9SKIQjtYs6/
obDg3LRXC2WKeT/ebRiNC9vukUEp3z7C2NBrKuTYzcZGzrdYeRZp+XL8mfAtOazVgDxl5OySdzzy
3GH2pFGC6Q3JXEe9WYay4F+408eYedE4+qsmHu3ejpBKBwjInCVbjXuRMOydIYiyEIXnvDwAW7/k
+S8TiiE6RuFCCpDB2eDA6DaUyJxk+s3a+JWbtn8O9O3zIKJuHdyxPtpGgD1Ln6DwZs0TMBXfLVtA
i326niNvh7pVXwQibEWXwNVsqSPy4BTYsga5yPWpccokVTyWAiiS8Gj36dVRGyxL2spUPdFHkIf3
7+UJxtKgLO6FQP7WUVckrrrLbmDheTcuvp51xs1Z8aeQKP2FTWRI088c3QPwyD5o3YhQ8T5pdJJ8
vIyQguKj/QCYULdo+JbKG6qHkMQAJsnRbo6V921NhvuDM1AZnF9CWFeSmB6E68zlL6iBrhfIyJ3F
ces/m2Jo+DyVBU+atGG8V2zlqF+VTar4qSvyL2kb7sV4mpItBcpUAkgX8BiQl8Yob5Ysi0JE+Q2a
RDll9u0pwOJzwTpMTR01GSu9eMleRZe2eFYFtLCA5L8D+IFwxev2tC1eOovAau9in62w0lzH0ERZ
Ydj7cN7nZnwyqQYTsDVYNhmmvu15KpAO9ZYXpdqcdfJ8GH21iafKNQfuAgh6mQmVBc0H+z2JSfXG
r3JyVFeQ9aY7Ha/pL/OO6jndTyNdy9TXQWoovzW15+xaWT5sB/9WOGRlkF6J4FF6dIDLu4kV0I1F
dwAQffIhD8R/IBrwjBB5UhW9d0F3UP6aYiU4kcfOR+I0iNgYqNdSFEUKkROgOYNIw72iJmfj5J1C
19OUiLgyfrp2iIyjYTIeO3dzZcdxk7TRIrDH7yQDKW1Lx/H18l5JIx2IYyTJnvQUJLun9ATWVL3m
hC5b/Ed/4DKCAnp0E9Fx7qxQZuvP9n/SSfrBHfdSaSY7ZpMQLrWPLKiBN/zwJSNSEHxZd3D6RtOf
XxFRlKFx/Y+WwvX7LIDxGjkVSnsbotiCG1CTR/1oqyYd0i5zkXUpNmFSQ/3q2+z4mJz+mirnODAQ
7Fx58bovUrZ/MHUalwG46pU7bGpouq7rbSxA3Q3qxWGi1PDWoNcJMhMviGaHO1EHvwFpP3JDjOCM
8QzfUPJV3us8uVxxtuid6XLlB4YTmO6RwPdDa8zqqj1IR8QOqyEHdNxfZY0+XuIHv/trgXKQOCp9
gQAXZz7BcvHqcLBuWRU8gmIb3GdrSJjGH4PxTEydUEUYuRqzyRjAbGvC6xif+/3dqKIQlTf11I2r
8m4uImEMaktzu5P/HsMmZBAF+MSuYN00kIhr1RE6sr78lr45Dn9AC640BIw9+JKRjjkNumipHzwS
Um0uaZd1VDH8cWuwhBrkaH3kx27EGXd2AZ0ir/w9PVHW/k2Jz3upi2BRcNyCO+M0X/lipJhwsyWz
d1k/VwInl1+UazKNikuQxBjovKwsR/BlMhXIDgdQKxyT8EZcHrbjOrOOHxZXNDzdHNsfGs8wdtLg
tmr0BtmYip9Tm0OOnTheJdsYpRcpuFs2CIcxiutbD7jKvlnQRG/tUGewHj6JT4xlE16/oFx1SPnv
DABSjPULfSVppu/9SYd5IqnD69P+8s363bGFR2gVQst0G/UUFLwuSqOYgom1fmilXR6FLKJuQvs2
qkTNZhlT+FcwRTgBsB7yTrV2URzoD9qid7wSpBArvN+4Q+RXZJj1cF1Ztb7wL6/mIdDuVKHtTaye
6mMN9ovlI1gAniMJ/kJRG3HV4FT+hLg9kpzdwYxqtKXmC2Hvo1JPrq8jteAxqM1+QCTZ6uydRleY
ZD8saCmD78kwkm4d3v+KHCWAZ8e8sRhrFO4UDjtC6TZOODOPvwZkk7iPomvhRdbrneLq2Cbxy1sZ
FP8xjAfDJJ6tzBALJ8Zi+/0N3aRIjf82b020vAMJLmKzcBThYprWttWwk/0NG/s7Pa35iG7yPT+R
/Rl3RUYS5xf6pJkHLgvZdiAvqaXTrZ+fvieQp4u3wLfvRCr97r1LsVfEZdo2IM5ak31cgNEI+v3Q
8hAQAn5/MmeSu52K3x8DVQdWJsl7OTDNwb2W+wAkuC656Mw3pJmMWvP+rbCHWCBSFTISde8wXxgP
/VZIxsfMZYalC940AQK+yj827yLx26GUAJSjpkjA5nPqFjqv1WRIaX8kVjcBtZqasA+V3ApXCu9U
WNcpt1xdg4lNBMm30Xru2gK2BZnA6RYpM12mB0ECl5It8F+HCsrUrJwdbH9eJMSTsSLYn2CWXf5m
0801FkdUUu5MATx+7SBSNBBTi4VCMTRBSYfs8ecpnWKK3z20m4Rw/XaP5/l19kax0g9Hg7GPbm/H
UVSKhN4ejOrSeurxXSQct7gWqCIgfTVb45aJYPtmXbv5+CB0ng0ezAKM9XX2P3M78Rh1/0tClw2j
F7LO6OisvreFWw81pa1sRzpqrETcrV9f/Xtn4LeLKO0DKJCmBaome47GhOj5irVvOpa2VBh47QV2
q5iXEccivo6kaUF27mjSpk+xv6Kqe8OwIrXm2V8hEoBxMnQYzYsSLhlI1zA9O7NiowNpfsljGjk6
u8P9X0KRe0AlGV1GDXWYdCdfNsB5kerz9eIzf1DkP5CUoNv9PXJ9CprVbxKadorhcxfrnXQwWVZg
vgkXg0DWGhvaoymDPUr7KEugc4OJLhzquXQkqlYaxLoN9ik7ddHHbd3XuzTghGFtAd3t6Ijn6MpL
6bu+JlA6BjPdN0zrH86Qw9R3bXPT2dftHkg4xiteyaNbKNyvxywxRfUDyirj25H21PxgZH4hfsOE
cjvedRpxtJDps4JzBU2IPHFRE1w0SILWM0dR7K59bEQrfaA/jlJu+gbuXhW9Hy2ATmT6yRRABXQ+
wpRdCWN8azh/BaffKfMp77hi+OOCux9ikUhriPgL3/MaxNRMSCl6KLy9INsQfKnTmITUHuQrXq5Q
s4ahRtQR2UV2l5+aTy/FyrWdZc7IMk+kLzyIt9DkkC926piyw1tvOgVToCfzwfF3LIlcleU3hP/H
CaaB6HR+rHgIULVyY9jYj9TLQklLkXsUn5uq0jzUQR7XVIKABQDcRfqeWuJ1Pc0Sg87abjhZo1ah
7HchuaXhX8521fynK9juNJQTkR/IeZbSXw5zrGfFV48cdqAKHAdYWSW1eCD9ot5jEoueg69fhhXc
zemHcNXAMNe9P5fkKMwxIue8sgglW5mO4G1g2CC04WqZHp6XQI8/XgISquEH36NRpumW1w0TZyF7
e7i/831F6J5G/Q3UFG8B1RQONbtB0r1N25NFKae/KH8rjx5ARCvMkRsGOldRClwN4pIoaMiaUx+X
cXGNP6bYqKHqC/Ad7HNX+86Xgbl54gGc2z2H6RXVnmv1UFiUnM7D9nUhMAuNQdkoZqcsxyxFVNFX
88ZdRuP6GQRMWQRR64pl0fcPAaCVD2EcLIB9kmEV+ipqE3bdZ/blPMZkjy+vesjl0rLncpi9imfX
/QQT8iNWiMELx0U7uuAGiRUCnVWGn6eFq1+6WOHrcTAA8yKaLKxEkEYw4TL++rIpRFFJT+MNap9K
qeqBQYqTyZkfvzeRmiC+dHaX2lUx4PcJdT/mybgY+R/aLP/+lshXJSOZthDzw7K8PsMV/syEsG7Y
sfkkFbIWBuUwh97I2GSp0tNAWt2HO/Nq6ArWU2ftq9zoZyQ8vVnw4ssbyK2t5vdGyN5W+m4ipzZ3
Hs8nLvbkLWOQSFvqR19McrsfDjHl1i77bb0XPklXpRyBCW1RuUTDakZynYT9iYHrDnHzdQ+wJTt2
QaioU8L4hE/9a+9qV91pAfQveHOmf06YA/dU2x93LGyyKc3Lpjw9S6e+oqpW9Bj0cqDmbyRBraEz
Zm7E4qbaal2S731LiD/slieGL0sxrLHFDH5qzHLQKBsZu52zHG4yt8OJ4U3HfSsKsaghBkpTXWIa
k6tqpyeK4A8AIv6KAXcVaSR74c7mySuRI0NuU+M62HEW6fhwuej8JGGy/HBWYFUV8/BGutIgSS8B
b8bxufWrTnYekhgtj51m2ghJNg3K56vtZ7K1uTHdc2zykorRnhQdYqL1pcV04ZAXiuukSDObsEVl
e/qdStXGKlW0norO5aohl40L+M70PgU+qKMahNweBiWNZQAuk0PUbHvUEeF8XUiPahz4DSPiAo3f
FowQdewRoTSAjYpFDBg7/TpW87Qh+yEy/47UDGs4Fcn+YWYZ6DQnFdl3tABmGykixFR2e3WYwdug
lnrxdmvGxGtiUNgYY6w8jmm+lrcx9MQP3+iLZs9jngHE+ipXpLwx5ON59lCM6W1DPHJXRmw+AXIn
gOhfDrsbjb4KdbtIMsrIgBCSk+EBDFD4u4BUMNiu2wiTC9YJpJcH8/jSfwcYsJa+cdZaAY5eqOg2
IqUYE2OX/V/FheZJPZ0amPecC9Axdv1VmhB0wO/pivXb9Bu0A0jHuVO3BEe5DvsXvUTCMpH95n/t
T8owKFr/zPTWRAVAT8kSgd8eCQutH8hUBqLv1HaWDQZD+47uNVI5d9wUgdh5D4RqLnc5dPMG5DPg
IhMK6B6nv32hnqidXD2PObppzHfDBxEhjCWx/qD3dhjO0ABdPyjOz72IbgStbf4AyRnU3hu5yq5G
T57gXLrSBL8FzWFQbuKodZn7yMwBKq+ptf+cenirBdG2hibQaVJ2ke1uVIrGpniiDXSSSnMznTno
sEA2i6Uwca1WXaJo3f8DkBkiHLvX0KqjA4eFc7TUKOGpjSLhGNWUhpg7B0Nw/yUJ8rSe7KJTQJoN
8WOmFAoHND72nxrIXmef6RlgGQFsyX2nTrBJRoJO6cV81NVDiXBwRDvAt5aoZLUw6PW8RBGOZwqC
V4j9TmQuybFYMdIjACQUSmiNsrbE2wI3tCjwaK3QixafJ37qAXISb1fBDyE+2r5Go3qNlcTA6fnB
cyBuMpZAlYkHmUQEZwRayjrCqaC4isxrY7XtOpHsEhs82HpL4w0noz2NsJYl6/B73pHUUTpVYlRJ
I5JZ/tntIHL4cvXwmatNsDssZps+Kkqe/XNf1SYD4v+mMW83Sraj+s1w6YDYuSEPwOMcQOnnVwGi
EyFamumhEkEZCZ3wP6r2eEJiJw9qJHuOpvw+QoliNunXfN8i4EwBfbMBVn5caV669gGQRci0jXJy
2PwYqNMUm/lSKBJxfc9qXUPPjhg37rrdEs96sTZvhdWXn1+GF50Rhki6mB8QbkjtPiXSyBMi7c7s
/k/1bOJeTA182E2FBkVIbvVu3z0m3u5oJ6ggrIrP5hbeiqPIJVVVK5cdfPMo+mgejEsrCKvT6h55
CF4ehamSFTQZha83B/5nQLfgc5IXRHV2HObYdMZQ5KLK7PMCdRpQf7jePmekGrtHG+0qwrO00MtF
GPIkJLOM3oB+tJFldC/atK6UE3JUCfkoGkPRjbrqiZeoAtWGA3goI6fdkfcrlhuJe4JJfx1Jn145
6cJD4o1wRxW0jpoVnjGQcyiBqaodHYkBWU1R/OcAYptlTnsED48GyBIlrFY+475f1d0uvId1DT39
sBtKur0U4g3VhFXPfN1Yg7DzyC4mQF9Mxy1I6dSfaPlA3/vhNVVXXDX4UeeFcyeVbkuubYCPNR4f
TDhfp4vpFuVW9ZP8fpW3JB+rulAaGzdYwnLqEmFIH35TsKUtEhZam1Jnr/agjNc3dXFsIEB2fxD7
h8O8SMNEGtC023erqzHnuFDdA38bmLZNJNKq0ojfx5LE6gnDXbc/xrv8N6yEnvPn+/9ZegAlz2nH
1CPxKHvT33ASY1Qx9PsFasVA2euVMoWzcEVuCYkVxxXY4nPMEkxzf/jtYbKcSIXKOE1PmC7pLgIx
c+Go5QpdHiRd+pFQ7suRPGoYVZ3lwYLVbnHPXstsPNhhx42SUCw9DykLPU2orz9cLGGNtsvOke4W
F1yEE6n4yWu1HWsuNMxXAkN3QcFEOuPP+Wa2cAvGSy5Ck+6LFnnZR5DRXzUNEsKgHwQVDXYu0ygc
t5PCLoKslDy/JfhT9gZ4bLXoKcwZumBU/rk3DuIuNGZIi8QjmgAqbeKewXgv34njP8cweLBw/ePG
2bk63r/I4xX+AneLP/TbLPX7QDy8/NnHoF1c5cuGJdA1esTvoQjzUpz5KcRBFpnzsawmQ+2ZJRrj
dEsqqY8I5bxUm5IpjL9e0oAUqiG6PMRBgVqoYzd6C2bcAyhZZmdDred4giCn+xwwSo5C0Wba387W
Eoe43XjtOwJAT0dR4KAniYc9Rdkca0u6rlK7wyfCNmlijxr8PuEeUvZv2MF5n/VayD89QB2NWZBl
JVbIZhQlwwEHX8+YTtSYKRFfU0bQsCcWqHbN1k3VeYS6wqZzqFiwiZ/FZdv+7Gv37HHRnMPspjWt
khZWGSnbfW1/NXOnOtcDuteAzb/wfisBY3qT1ICe2Og90HD5my13/Jkc7MtZH9lPZH6K3oYj9dL9
BSUXhCKOWvH67ox2CMKL1GHTunLQU0E/2nt9Ikzw1xnhKySXiVvXxxBZcKnAlMjiBjZqKEa9m1Ay
LrILHQmSCTwcJXvoWFYPkpAJmkhMMi2RYnymGEFW0pADGAg5EMqfsjg4vVgmnqFNPQ4EHS+8TsFY
esSWZ5APvO+/5+QvLtoI3tOCQS5fWV8PgyU1gV8QWA8iVuYhpsySSFqdDaDQonAi8zMzH6w8GdTA
rzRizlwLqKnu9sl4iKq+QU5cBQPEt5ufCb3+/vYShltrAq7h8Kcd8kmDanp9h6aoEZFlUaLBKM19
dKlz2IQiM6InyLeOPa+nQPcqQxMicyWICT97vFogciS9ntg3ZrRz3VVxSrur1XYXOq0yfeq2VW6F
iIzkPufGCyIacBNCMDMy3Kjtx0V9KBaDIipMFNJuitSog0i3LmERDYpFzXzCnhaCK3CnImlA4vQm
3Nbo5mSYULC4WJ5XnV7lSx0QDtBHt6+wFeLQ9kMdscFzFtpk4HR9XYz+W2sJ5M6Ix2CsPU8XX/tU
5OPDP0dAmMyAjZynwSTe4c6PSmPXAxR97dNLYMa8uc4RlBTu/dyW2c+VeS3oB0LLaTq9qabJoVlu
k4XunjcD4uHQSDiDxhhSa7Ptk1Ja8XungX7DMMWU4eUEI8AA0qhPsbtDOrXXxQe2FM+vWQNgwN1B
qCgDYgDkgc1XeG88NZaWLiMULZKB8fk0AZ52oSmS7rm5bn0y8s3rdqubc8etyOSc333jNLQFg7Sf
82UF5QfG3AWz18lZVpUQjDQfP8RK1G64NhnQXvpoQF0+YgbYqT5dSouD0shokpIUY9Duz36RJSzg
yjRmW4GEvGvM7Taj9POd9EMVXr5kF5n/JaK+poJhzBkuhYyEWcH083w57jLT5B4P62ea+3yXHEab
08ye/EMlTrC6+2ulSABb5v1/jGMcVMW3jIrrYYRsgIkRaEUIKuujEyB7rRgIUhNKBcALxSuw2+WH
2o2uQ2UBwV0zupgKwkCJT0QvrfPXO5EJqEmj1Z/XnW5ACWqUjEsdHl2CmSFjuzHgGwfMBJZlDSRL
NkRm5dLtb7YYJK2uJODJI+Nnug9jHJLet15EpLrUzheMyjjF2qxFMqWgsB/KkAI7neDsduOrtFIj
DRK3U0eQc54L+jBtyX3Jd78EwO0+HDUFKnLkhaGNWPzx8J9XNBLY5LlxxHZUhsFDYIWg5KmSSjKX
DXAr8I6HcSqtL047Y4VOM+wVW0fpEAfny+CxB//l2o7iaVbuG0psyqebr+595T/ApSjZ0K007Jme
YHdL3TtuwrZQJb5PBVV8WVeTc0DDLBPVPtVFNKsoOGWBx2chDbT9hOCZ6KXLJUi2FDunXmd2/chB
nYRAwxjjK4qkcBArcaYSWKRawCh2l3c+ZWCrtykje2xOL/jFWwn3iO5g0IqMVC5rKsQRNFZNtxuE
f4T87AT5MvQ8h/chBN99ra6t4RXfILZlvi9f3d8YhK3afa3RLoGUkh7QaA2v2KE9rsJ5R+5Kv2vi
Sy8xhQxC0Q3qiVD8XxzIYQ0KigrQETjGlUTR79fFr/Z2BwUERPOZJ6NiN6EUGk0UEskmjt8bFxvx
JiVSNL7x6S8tph11nQpxapS1H/p9yvdgeZDSxR3fceSUYfKDWDnRL0P8zaJlQi8suJhimXyuwGfs
zMVbtaUtgPl/7Ku/FieGHefKArxKuTzktkP/Ohr5dmOckBDO5DbyoCOIt+hjGY4Mj8Vd2V4izQCZ
6hNmUpsUKaTu1BI/5ZwSRnhalrY2SnRkGpQFaWx9SxjgkUS3XWf5GKLJTEMf32GJSfGP8ruy/7EE
kdJN8m8V8RUBI7tf2UKmb1LohCf0r9tArUPalBCQ6HH18MHgfUttwYhvv1pS9lIJKjMhpB/21H0k
t7z8Q1pdUM6N9l3oftjW3YG7fHFxppoXvfCYU0cVSd0nir/qeCu5HyK2REe/lWkT8kH1ZV9y/a8x
+s6im/cAamG30fHutpoxOGTM1GvyzBEwwSNRdwPNOkhRZopPymcU/qSlH1cOWW867Fu0bS5n47rW
Sx1xapt7UKB+d01OYJJEHuykJLNRP9OIn3TsgDQ2QFk5zo/nGFjAXrItAaVn1YeOZHFxPjknQeqW
0tqOrtsG0RDXuRnTbaBosGIMm6X/l8C+fkqCZGvTa8MFmwnyRC35+14fjYUfZ1/LIFscjnof3ymp
pYkC73aX67D2zWmQmK37xdYwUdc+mBFATy/vBYPT12nU2BSmgAf9QPGmy4ruEj2pmWYF81EBLmo8
kJlbw2PhiPHGRhS+KOtUk18j8cE+vOZl1K7Y6JQGZPy/HMNDOdscnTUHBvNG9jLKDLpxPEGUbt1W
MoGBTWbZU7Bgk/AHcUSILN6D1SrTFGSvQuLEHqwbHmr9y8KQAMgy7aT3CTbyOz623+kx+HhP95Ey
DnI5KRKZKDkMAoegNeF2rW9lO0kL0N6wGoDgHif4Oc61Y4VvWzExO+UdIWbDtOcOTjB/Aq9FGOgP
pAV2no+EBOg0kPMMUmVosW7bylTsIEaPjKiAVBX1DGlVHpn9EN/F2clcln0TsaWbejjRjv61lxt3
g1L4MQC4M+OXecY7eKc0UXMwICNAgti+hrsCxHaVg0R0N+G6bFKvrAi+6hkjQiOA7Wkbi3e0JkN6
StPntnGnU029SFUKH2oqBwwmK7gNICXNSGvWElx7prTlHDDoyh0qFGbiLk9jkzxWSPi04FlH76iE
9K+/9G/GUyrXkovxGz5PVFXRb1M3IkTrhBj0kSZNbxdNmaxcmSkLXEoaafdIABCOF1KMkXoV2Vk/
rprdmkIhLuOxtc4plIn9UWe2cI/NjRtEcwIJ03sE8QmDHvPAhQPS1KUI1siPCOlfFXmnMULG/Li2
JACAyrGjfolRkHN5hHd1FQHQvGuv67EIyEtG+Lg2a9Zracz/cY99c059xccAf49fsZ7mmiCK+dcy
nqc/pQs3ylllIN2d3eWa+UEbFEafZQvTOLv/LMsEV5B8VYKzX5icZ3ZfqLDSwx6R9o3YBhpfEAMT
jtJJgS59ApmXYPeYM3wJrWSOsNCxZBO4O0/ZDWs4KsMXan085sEn0I4nxHCYtTqqiJ5/dCcadUp1
cTyoLZg4ub5cGm/I3oYE2KDZ+6zZcArwu51kWjHkfzganDnMCCckfRHtS9Mo+nG+3aAJA54pAAcx
nyBNBC0qDLVD1h/7MsXoARn6kJLVTsCWsFwTF4+5sh74bc9vzZw3AbAYlIcpAxC5kVfsyBzU3Btg
c7nqpERmKh3mt4bM6uYHPLhiq28eZTqLlYYrYnBEyn3cdrrlgrmrDCUkZ6Kcxrwm/REqMgzZf74g
AHi0eqPPvnbPF5Sb/M+mSRnsBybWn512xakY5weC4DuOE154vjswkwpvhae3kq/qgAblZD0p5cGM
yFUoqssRvGSVqTV+FZz0jb0rKYbb/L5Zv/MKN08+ez/VyRHZ+86WVggH1Zd6tYR85+osh/hqlF51
ORJzGteN3KHJv0pjFHqa2etwO5192HvMgURrRh+u66xglJ/qFIBg8V9JDOaYuP/22zN1hRZzcDe7
93Tj0QpbjaXmR+XsQY+rWiv8AEmTUm3wKGoZK3BNroIG98hqdNAR9u6SFS4NY/lugaVcmyQ9cSJ7
ykiby3ijHCq+mOYEEFE6KSAwkFBRA+w58bfyVTX8mok4iu6/5c2cs7+lECesW2b2prYEiTIdWzze
Fjify4q+r8ffwABrhrEmBNyqa/tp071ZuOUdvfVygUNzi/vvk5YNoKFG2FI5R8Ad2Hw+Co3gEknx
8JY1Hp+R+S9865uvSyg5G8cpqxHzx4AXVXHAYA/k1cinjnKQRX548m9Dkc7wTsLcFEF2x507Smjd
L6IFSXf8MLIVfVu12k0EFbVhw4LDpdNXzvdA0CdbSQe2qeNyx5xYTRjRRhHO0XfLWCnN6nZRSDA5
F1wiLitFU5f3KXPeg1EfBpzAD2ZJ1RNmAZGTFxzgeGtF/BYdIdDZCNd/e10bevBWaLL91vj8JTf7
tQWCK4zRDQYnreVJ0rkYJgnXo5s3avMRbjvbrkNcfvkYSZX+ciFRDJkanViZTr96/QZ91z6o5Q/q
/SiNQCEUH8WAfYk3vqnGxYGJMb9P71id7Tm/qpHYr38V0dvsgwshYEzg4hY7btszPWU4S7ymYsVN
6alRnJTvQQ9iT/O7a8m6qIIQ0AqKGc8IN6nXvyTTxeOUXXg+D25D5ER1Qqi72RJC2l1VupVm8uZI
pLhJBlx5qWtqJ9EY9dWhwcl6ORr0zi8CkKJg7nFK2tOcT8cCpbHmmgLMyVoLw+onN+MlN6mNEU2p
gB50t04S4DcndCEAd66n1GWiT9jJdEvdDoKZUKgOZOdZoByjIRFA7R9AjGFYWGRhxtpZRrfUWiRr
kfw7MMLSVV6crakLqkCUVIPJPo32fXPM+2n5UxDbSZ3uRJnkPgRLqXF4hRlKtEaJUO/FO07snSHS
JeFUBB4tV3HurBgAK/X+7fO+V+VLyr21a7iB9Wn8+kSkccHS8gD7RR0KAQHNbT3x6PvyymgDjGv0
NaddnyRU6QzxMAbTImpPMgbNGSZcp3nWqInpl7iHbPKz9cMfp48WNjM4an7ZvP63XTNJyWMt+L9x
juHVnc5+cC416V2UnGZ+uHdJEfNvUzamsmB5aP+fL3epGweLwg+CsyML4r/dG0uXbEEG/m+XsfIO
2Puj4fZjAejhFOLdlbJQ705c7sHdqhpI2PnhJEPGmWqLK4JWiwGpsCJLPChcbindZy9/AT7J6cd+
l5jX6DTas2Pc6mUcAZ+oc4ttU2rDwdc2KDkW0kuau+T/6tzxkdoeHl4YZ3KCgAqR2PVbHjvtugqi
E0EtgobyJ2edXcJ4Wl2l1zb/ymxesb4jzxvebp3Nvj2pOvMnoh/4X7eI9XGyczCbDUgJzoMGRW+H
kvjG2oLxHyFnWRGZyD8VF7mkXq6Wn7yaAEF4qTJ5l3iQGc/tmTIHaSZ67YJThkb3JhpWo5nCtvmZ
3F6hyv2wiC7BJQJjFg9BsCI7GyrApDt2rrGzNDxSVMCqSRRkFeIwC8nCcwJiaWIm8jOBvdUg5DjT
6ruiIkzxCzsGvo72xJT9iJ4/3TgLyG9kqvXFhT1tHVeNBuy4vaT35TUrrJQHzy3gnwv1e4bXlbRe
5zbpF5kRj0jey7DK4jPFwcw0K4+HItVQ0gr+SKurf8Qq6hna1no5apFaxIS33eOhle0G1XMmfqAt
PQxmG6wbAsCa4uiRwIKMxF/cul1EcIRw8UaxVUke/bhgCEURIldp45CFpHg2J9t3OtElpxr6Ua3W
/7B1yZeVLutPFkBqwkduyY88Le7frGFBLTbjCRvllQ6FtOdEG0fFnnBjmpHZqD5giGBFinhSf8mU
WzwTPx+xn770qGiWXQ2NpZZwU9Xi0tuc5ghbXMxvfv5LhxZU3nlOY7U273EJ2JNhwECD9bDIsfCE
WHrc+rcrn9t8CqT/oKrkMqb+9fOZlWcENaRQ8Dlh9huAGQoXfNGa+gjVekux485Hs+/TGTe9DTUG
0ZMRZZJyXQn3/7GTSoDlciE9xNIO0Uz2E6m5uaxD4vUqo84M9U9wnkC6x01zM8XDZrLmtbWEpzRf
JRa/Q5CpDAYfrVFa0rOR5HyPkfShS/If1N2n73m22x3HawdSTy24/OGlUPlEQLC2tlhetfZZt9HL
kMUXLYtKwi6r1pRpYjj9A8iVsomALLYP88waJqZ93AKXc6WUWvgJ6tBivhMjs8aOHo7Lt+TIZp+F
Nq+ZKeACb163NBjzKKHG1Pfp78xsvvvmJWSro6N4ILemfKknmDc12Vwcd6PXsS6Ird3ykAuTWXR4
Vojbsq7VCo/qCEL5pmRYDgzKbWUJnOpCMES71N0Frj8VTyfwasN48xSjcRDdrq9zhGrf8Fwu7bHl
px1F+kEVDGpOpf1XcgIorbSmD0GAXliePjGahKnMPNZQC01McXEVfg1SGOPt+RHcO0Tnfhpd/BBp
kAze0lR77xj8qz2/a1sIWcUswkr8XrL098YKhTGmx9/QUsRtTc6Ab9fJk8akhb+C0cV1PlP4R6QC
z3qxcy6x70uaEIiRCOj15Bel5QQfKFbitsacbfKRqPoEeKMbBIDD/t+3YJZ8A9+2vs/MLrf3R8bd
HqO+T0oKQKpfEFke0mByMsjOCr1nLNex6s5WlV7Yk/8MoAifcXpyRNIKuQxHMlwvVR4pL8NeToL+
F2qCsURZH7oicj/puG0Q5w9eBTHce/NVNgEwjLMMvAVsmS9Ow+ABKiqhMdrIkdJR3f3hVoVpEmGa
qElqtSg+wEffV9PW3lzCrmMDfn9kWsOeXfKOPsAczS3Nfyngei82eTDeYA3MfZsnDNjNOBoHRY77
hHLkBbjCo5LblSh8iOfX14XXsFhqswcTnDtpm6TIg2dZOfwZhi+RGUboTvAeXq522N+TkwjF0o6G
O0BAu2vx7Ui1ECc6ZLFvhjya3l/047Yl96EKuHATRMCUqZnBbMtU7cm958a7FNqkJetWUGWrLF9l
FQL91ryu0osfOi10z1KhH2DXz4jhBKrG0ASvLbHIO3Wq1Myh35J/oKK4jvvBe7DWaxnUQq6zhv+R
uBRJR4btQEfwcKYJF+phsO1gE7XQ29eaI/B5HKX8kscVx3CEGxJVGB1BuzC7nmrj0yO00HMYxSq9
al7cqy3CE0werakFetrFk4XATCuGzLJ4bU6DoZvliqS5HtA1MCZdDVm0y4n96W+yKdi9iq2JIx5k
0GLA+f436objudxYXj67EkD6cczRlYxWGNCs5b0r70Rd6jRnw+h0/Ec374To7TMJzZ5Y+Zn/kYsg
Ah/rK0ec4h4nCL5Fh2q8b0QDE4EfSXco0AyZ5QKI9LbUQroCOSCpvIVVD5ox8TDh8rMwmJDaF9YK
vR14wMvJ9xmHSo/tto6A6gGSOnETgGsqDBzV3iQYvqflVbUF0JPFKBHKW9KBqbMkNmDxoaAG862H
ln5hICHfzNZERRJ5oMR/w0cs/U8SwzEoFgpEu/eJMo3tNQjOLZ8fK92dvsghxo7tczYwu3DUo69t
nJ59Pcyh9gHZstdRPxZdjOUryirIQgh1VA4yblfP1nOKLl0otvuY2CxqZ1w6CNxm72Ds9xh9l97/
xsUKbljVvyhX8q6MfEWOxBr0PzW+SE/DUnkpPoY1zclwQI6Mgp1tQKJwIQz+Pd8yXIZkKPQvEWHb
lQxrdH5G2NwL/CsYIlHeYwwdFYOiW/cfqs28i0VnPRNWC5E5ATd4vVBg4YXmXYVykJsBZvsiiwip
47L+GqxBtEc1sozw21wNFVj2EqXeYH5u2mVgmN2Xp/IW8V2cQSQYY1k6/tTBSG8wA32LG4aSUr//
06HPCHCpnA3xKHVF34OGJOs0cFGGMO46oTdDaoQ25qqgWDYUm4u4fQ0xJT+B94WoSJRUFQIRqEpW
S1hFLdCsOCEzf0QCG3mhMhRrTo45E/AJTEMGvLDcGYnT0OY2kluMIkcTehIKJxI8Jkvz1cH56E/x
jSamIuM2fVEpJSvCpU1B5Xc2UZVoa3naJCdqlXPxe+853nWe66MqCFWHRcqOl/MWx9pNCH+K/58D
hCGcPv0TgaswZWE+pYTfBsYMYhslZ5nn4H90/OHQbtLidbJrl1Ljd2zVZJiDdP+QQwf0uq+NkIpr
jMGPqlHyFBhcDjWpHj6xHeU+o7vYqtfpWKVM94vM7vdAXyvhN+PrH3pz668nTusn2lxfy4FcImuq
X+Yu9zPW+D8JCzCd1lp56UL8rH5uT++rYCj4nrXqmlc48nYFfgf8zgLMFe0qXWl3a0KVHpHOPXPn
05ou5gLb+iBmYZ2lPxmkwG4Ojs2JBt+JVlH+AM/OrSkevvJtAOXyC56rLoFtPg1gBLWS98Az2B3v
4xtOemXnnc+n1678kUcxRqvB45a3aXzqXpzub5BTXHxN6/gNZgGr4NVeNW7j50I2pYmEGcA+lKD9
wT3WOtdci1614tjmgqI7XTgmmRw+758SLbHU1sKwAx1lUQrPS2mKge9H7hNCMI0pXmWC9zy5CmWT
dDFDGe+n0zGRO2szy8aoNP1d8LjN6rJzF3zkbWbPNttsv7CVnIvzRHTLNRsBivMbl29VrkvrpDbt
9RPD9BWQ/cq6MppWs4qTuYUFI/H2C4DnTWi99gN+fi/xchgiKHgvVpZu0x+MvB7f2ix1PJ5dYsBh
mNuXyX4UlUJ4MtxwdabND7esZ27T0/jotqI4l6O0MpiamsB3zhgeMZKCl2fyKjXDSylzXvmHt8Ze
YJ2y7OaE5SrShVWw9H5pyZ7MiG7NoFlS/DWxqvT4eOc4h7STrNDf2zJ3jAkBfeB7o3m8XN5fEWuZ
J5gapHGzffgJHlqKw5sXKWsvyd5haOielpdR4lzwc+0IvD8UMVOOvSnrG2U5oOnyUb3h7ZF345FS
aY48xvntsD1Up11lYZww/tiHfS9dBUqkvYynr1xiOldwPx7jtyOi47bo3Swpcz2mZm00nyk0qIXv
TTQObaq41wUEim6xP94jGeLTm5Qc3M0lhJ2lj8WIkBDM33e6scIvosxqN10txQgnTHntoGuh7cJE
r7h9h+zwaTfV3TtKzVCA3IPLWFPIJVJ8CYNT2qJe/WUmDDWsQXoCXMvqZUlg2j2mO4Owp7VyoXA5
7OjR7hvH7TKHFAtrJaCB7ReYQKtIMM+CMnXAfgGq09CgdT1fQvWDEgO76Md9LeswjCJgUnurjhQ3
4wRX6YtuPBV5LsOkz49RoNCOc56vzBYaVK9eD3Y42kr2wYbq7VLplv9nNI9ZWWX1/7caTDvcRYfn
mxz/0OMwUKQ19QLZbfXzQ/imJuPIJ8UJpi5SFRORL/u1xyW1hQZ3G+EGUZcFFteDd4S4xqUkAkmY
0i+cYuxc/0JpQGssSwtw3iL6n3PsyEoW6pmENnW7z9sv/oq16IHSUXAXARZ7HCYAtyj1xjYsHkOj
/GTxrNc0k5ELvHKNp8CVj5946hS5skbbQIrpJo4NLga6SIqEk0SOy5THrYUaYd5HuqCTfo8Jt2Pb
N9zLjCTfd6AYUislcIenQ87W7sBubYpvB9qB8gH/IwpAbC+cguEej38pLhra01T59QVjWPMqGHVS
XoGWmzwtCfOPzmBbxmCfULFEpATjZxuqjRvlze7+DYJjVbvRbmj2h0PCe/5r86TyAeF8kCAcfH8o
vT0FKswCCcFTzS/8o59mgf5QmjGsvhGnWrneKg0hCHgTOB2nsOC1Vvd0qr9X37gO9/MX7vQGEEYa
GYvA+l5NF5ctghIdVOVYVLinmKGipTvD0d0OP5Guyvi3VQj/yQLbf/lQhI6tcRfBjAWUenOhfKl1
yhQO6mziNAo5k1K3M2OtLb4ZnNrAD8TWbiVrdAvKMfMMDBPCK2DT3CvQNHSe0XtCZSOgN9LBDc6E
t9iWZpoIds3bcWKpd6PdfXmL9eZFWiMAUc1y+sltK1RTD4PMPq+6XkJMnNA4r8vJf0kMvMlD87Rn
dM+qu7PGeUT5ofHmfPatQ065stlBMwy9ufudVRwFcaYhXA3hjdy0deqze8y/lZkg46oCURXFceQ9
qHrDwy9R/nWSTbsQ1XlCVKU5/3J1hKtfqp72KCRMBLEXAOGoeA8S/wYUaJjGMm3g+qhnwMBGmbt1
7Cu1GNj2+SDvGZGmWcSPLTW8bLJ4xCrls20BDDwhzar2yqlejZBRhu79NfJvMsLxp+5TVnuV0JKz
AtlO01c9UpTFthYYnd28cdlPvYqBt+QFlZTYgR0v6eU/5LW3qhqtJwbHcsxk9SNs2MyY9t5sjPi5
PzVAMJsZ/QDdgtpPdjDqqLQHHdxlFzsXt5iHTGaGPA7OtVKs9Ngp5Idq/GLWgvjepqY9oqCTvdGr
Kvp6j9kGAuPk5JofehO1U659GmzWshiERh8lyrYYysI0QjT1EQ3yDTPaN5qPUpOpwecNe1+M2L53
bOdPC9FrqyspljWpxjh7ikBNHBTreWm6rEgj3bm1+J44zTkejlRMtVvPs80basXGlB8J7byxDjkZ
LvpMNzsvO4xgqyvj+ATe37MlM6313MCFEmMjVESgobsYorhNnPHgE9yDjDfRAFDHypNNGPXs3WoS
1v0uzxaHpd34SC/LTkbvrmSbd+AIKWQuWvqokgTwfNIZ4WQ4NKeEPufr+jGLj3uIudQRKBRw0IrM
zHvDfkKy3YfKJ6s5rz0zYKO6eEmGc1/9AvpjgBGEknfctIq93GsFVm9ZyWS5g9wJX5zAUaALetlJ
LosW3pCFHCFRODZXsosWCDJRtvrLWQiROmIW1KAXeS5NQR7mYr6FSsCMmU9kzpuJC/u3E591LBSN
d+5aQ2lQkyZ/vSKh5BJJzRc8U3Pr+E6sTvkdlD7Y2ooq0L0q8pgGPm9n6hS0SEv3N4AGBcbPrh7Y
i633jg8L9UtAdy2Bk4sg75uuALwY4wbaokf8yFk6FpTHnCa1ewncW1MklYjIv00tBFruYxk9WVEP
WOKrlwe4tKkuMRA0KLGvosmq+S6R6ghJc/SiL6dVRHg0zNsCrRWHslj2mUg2WskS9x079FQn5mBj
BAZPaSKxvVliFpri8ZMf1GM/umqqaTT8cpCbtBOMPirwCl1UzM3ymRViZu9SokILmQCZKOWj0CrA
k3Vk3D/ypQrBBzvUyxqJ4eRzYs9z9PTOt97gy5vo0IE1jjO5jlqtCqYGrNLSRydtdhYsdWBmXh4G
2aZBsIO5UM3Dl2pWDbZm4rpNZQMFarwLnlX8FUe2rRjjMKIisWR4f3qiU3lQ8iaDhfUfJfNu4wyy
UnB4XSIJ07kGcOWyHNdxdZ97yOKqzAzblRpQ/1fA1V3wKYFYI9f+V8oSmssBa9wIEjbTdol3vnKm
cwqKvE4gUkf7i7iuNG4KM26RTIUekrbOfSlCgfkEbJJHN5FoA/Fymf0f4irhJw90b6VBJR+v9anz
JbqMV+37NCz+nNOGPR0fxIeIuTx0Fw+hLnhlWQxAWUypE1VIYJNl6cmPrCDJA1C/x4hBbVcl8pcq
gzNrZN3lQrr4qZdsQzqDVEncofDPw+Nvk+pUZ70UKt/eGnr4pJDvNYvL6mimUSiEb429Sufd6h2U
fLxYGYV9eP8Q5R1mrr9pxSy5olKGEQu07EnuPkYPo2gUtmwoHzDFzOqQy9Ik7vChVZt6Mnu4cyus
1je1XqQAVRF8Mmz/DRx0MWDhShTdKSWZN70dBUmKdrJY8n1IfPEqkR7Mn4pGOeoKbRfDWDoObXRE
Gc0j1pHl5G0NSn6h+zvCkxJaSd41J0KRSrun+MHHPmQpN6cnFy6efl8tQX+FOsNtXnj/jBHxQwnu
jucAWLhMk8Sske4Einz2w1T8mD0Ti/3HDZ8UQGisPfmLUz5bADkb6GU5wbpepjmhhjUlnmIU1UDp
h5yOiO3tNNhfAsay9RtwW0hugIxioFlkTBJfMwW7IlnBNI5A8KxHdZyaxfpIFQrA5W4XNApEL1WE
sdJcRe9UymWUqjZjiKz/82vU2LCKVKAp2SAhg2zCyJ8xUoObjA/wN3dvQpm29x1csyc3nBU8m2Ir
jDokhIGr9ZJZAb4gP4rKzWS7BmlHRjZ62TOKb5Wc4I/0dQXCbbI2iPid4QI3WyFpIy/BCusIbEjp
Ppad3TyOfqOOaLtJzy9Oy1p3Cz/drxXL6S9Nk07ngoxlnMp09WmLPBqFXevuBvEXmDFF1c6pBZVr
MzG0osvsS8oi1y9L6jlINXngStzvuFKgPlKEKN3+qu46xPNuORYTfHmo3Irgh3qco4CswbNaSHSL
z9+0cYwAJ6XW2ZI1YmOCr+BhhAWih+jR5LdW/Q6rT0c7FfMqLLDMCSmNoAGhUzB1Jz4J3j/eLA4F
pKyrrfgfPFZfooSf+wdm67uX9uOj6f3Nx9bMLEmFIyq29wyZiqCZVU+Oz+DuaVvSIUNF4sR7iioL
Eig6WoXjt4fnfuK5wME2AqA/seO3o4dcqA/A2ZTqV3vo4iXyHH+b16oXQQOm/xjI/Yy/X2m1fuWh
3mZKTxgwQyRT2R/pAVajUQKtGEZBrgJNFgA79cn+iX2mTJ+/4LHJv8Cde8/3bFk3fN1JUasNieyl
NrgmZebJXhpjxuArhDWpze9IeXJ2VmbzcIxm1B0VzzF72ZAfbnG2gyYIwEEf70LWdiepTn/4oPZA
0qw+ocIml6NAOSeAnzfi+HTABMP4MpQXbB6bd0SuElec9tb5Cw7ePASpttiFnqCACeTZqVs50uJD
60z23S0VcFgKfgk6YrO8s/8cRdGH2A7xHG8D6GAcMNjIUzzevMftXErxydJEzMnYMbrJnqB0/Bm6
2JAKYv7yODHsmfqIOHopWqOA4k79f+GFqd7grdzwBmqsVNrsltNNqFfX9XfHRvzlYx5bD9H2olGi
vus4JzmGrSvZXYWv80BuqAFtIUuDEV3E8JHA24tyHbiUaycOO1MM+QgVX4MlqXMUHE/uQU0PPiey
oO/AkT694zgBng2fbL9sy0fhWMdffOXTyjl0WICwa3OIwmWbNQVoMS9EGc4RjKDFh9IuJgnIrdub
lZVQc2FfcXBKYz9aq7szVJ8FUfcjwdnvd8+wqlIpOwpDgmlh5KT8yew+FLW2MbotCVaievAWU5HZ
mM+BK3/ba/erpC2V8alaNIwzHrhGix05nzSvV1acZgpK/WhqRp6fkUEWBpFGJ5VD5GGC6SkkQj01
VL7lrCTO/i/XFWWZi78rEPMAjnliVDsVGal381M1/YE9O4XRC/R+o3D1mcf1gelYnQhs/gd1G2Rl
Tuf2gJWaz1UwJaolYFHKIRpXP2XvhGrvCgmg9Le7qE/ulnm1gMGD2atIGrI+NkCIDsJq7k44utjX
W+RGl6LS20TtLyXNQE1lHYnvCYh9AyP5RKFZahrO+w7rbGA9DgsUYVGA1035yWpO1vwn7aw21w8J
uH54a3wi5htr2IxB5HqkPwU18uJ6876GOBV2dnEJ00FXoCiuoHz1GcWoC9ACl+n/mDRtP+xV6FQW
MECpKzD1wPKy+aOL2MBKf1hdj/VaQqmeR/m/6n8oSzXfTaAWJ+ZNEylQ4XEjlGNEa05fkXleH7Np
axnKNWBwDTGwV+70NoqiUY+z5YEKHCsNa+YqbQBITTCVZHN1YSTjjkBcfZFLirN8QSWyxZhayRIm
wY2oPb13SMMfnYVo31ytiIhSSBr3wFY1I+sPlSXQp2Go9x9CcApFKDvd854uIN7mQVVYFNJ5nNHp
5++D5U1dn+viBDGvu2V5RHuADhrlwsqW6JaDZg3/H42CpqcaCLtJ2ysSaza1JGVA/MGQe76Z0lop
QuOTr/AlVAVsQvfCBF4p0Wh4PRaDGH0qS7SML+28kTr0tf9rU+ABQHTkS1mHBoIeUnfcPZlEDYsJ
g6McsMwJeONUTDPuDkAmPzYr+rmj6h+BLSMxN701wQTeWmWf91PNghuV798mCm3Vmsqsn06Yc8ak
RVDsIHXDg4WAXBziB1raJcVP7/ZgQL7IsNP3gJgVtYNPtHj2VcOxvHgDbKuEKXZzVC+Z9NLhw+0A
71mD1eJO/nA1dR98y/qh+zB+MSbwig4NOSt4BD65dTyyFb3R2uRGe3GTadmi53nBfnTwLeIK+8pN
K167NVgfeoEdgPCvFAtOou/9CrqdqdZQrQi1GQe8jgm75fQB+nyT8AsJxy5NKfPvoRekxFjExRAs
TYm1KlzSNtnPhJK+r7slHxdx7wkKwU7zdshKHIQass+xGBKRop7efvADVAE+HfgeBx4CaYrKPu9k
FRIJk8EYonHeGMym+PgXUvymcbLg2O0LV/l2ZwQkybMcC/60B7MdvHL5A9fa+qo31CkkFtxdZQ6i
5Bm7UAQIaLQjZpFtryyPKZxbi9ZlLshLMAjD/5WOfLhzbLUwstAiGktVhBPaibd7jVoex44ejQso
FcBBHdDOO8flpAdrOJ4IwijBWSbKtF6CANAZw3G8v5BJEsnLvQTdwBvqVDeq90eof64ov4u4ngbD
IOsTew9Rv6VQZk3Dlbk11lKyuQrbyVrAd89U/yfwshGhzPGSQBhWG4HY6l25L665gLjBkyXmKcNx
9CemW0H8DEGCWN7P0jFwGx1rW4KHbR9RByp1PT5LyrCQqgvXuNLhGaq9VhDCEXJgRoOLVaI7dzaU
28PbPezFsGesK1QWqd2YsjXjVPgMPVGOrEoeQ1tlHhmoofa8e2SGAq2N2Ywyfoh4laOa6RJb7FYc
80SU+IkbksnL+m2Wwm0CwvvtH3QD5V55oM3mZ6O/Cyc2JuKKFdPUnRXoQsV8aGTAAeGkbvl9NyP6
p/kQYAFGvGa1kjLgk0dOoLRB9Xd7uTE8HCeSdyqp+DUGh261b/CDLQKaQ7FycN0UlnNeZMSojZk4
ezMf/SxVvlUJkBSPbDn+gw4PD6bLLUnPWaCRE8d4m4uVzPDBEloxIXmbbqORUkyWsHLYQ2CiRDKB
mY//UJTxSwzAuwe5suS5MwLRB0czq77+LpEfqBYvZtHSarMC9bIVx1rJ1Qj8lVWTk/oxlUt9urCq
ryM0kP26V5vNPDCKmDd40UOjae0+PV6CsEpbkV1kgtOy9hGUcV5DmcL6OJT0e/U0JlaWG6Rb0EX4
truRX0vFihaXR9fGRx1EZFG9SNhHYzxBhI5peQvMBhk93vnlVK9J/xsBBtlMcxdHMiKau4p3rOQS
j8gPAsn18t9BODQxDcTSrhmZtOtwdoy8yqinPfEIKcei0V1Eo7GONKvFlo3o2gPTIViNhoFYToCt
MS+QzVHyVrRiugwt/dLKqGsZ66crcB+nnTz8UbBnUI4lbmsh2DpaKYMijbehpiFTns9BzCH7kzRK
LasVR5l2tCObtijnnxYWnKtnBLDQK8Ypxcbe0M0E86eHSnO5rNysPhRZaPDGNsXTgN9ir3XQwuSU
0SYcAcdR4q1xnUxRwzptJ7M7+k9ZCJeFtkPDytMFW7pk3anOWpmHZyPwSI5IrhxspqnUr7x+uwQE
nxe85walC6vehhEwp3sE4dRarc8py3ZBdERir9l1U8hdfdxwHApkdVovj2FFriQzrtbE03zV1xxA
ijfcqfVGa0dBm4lDgVYRrDrKhXCennwVBuKkfvVj2BX1bYvFXk6Cm2NNdsIi0p62aw/tBiEtW+AU
ij7PMXBGuH/JXMehFpzzn/vvuoffkk9O/Vv40+7WvEywUXcITmJbRohOaWai9WMF+eHDBKNVxZbV
CpHBdAaUUqdkDt0Oqwm1I6k4LH9IaWFXte7qdx71504knSpKU3CYe+85Wcfg7nxRSR8Q97zWYemw
0AScuKU+goHYmo6IFZOkDSSHhY3/Bz6KGZE+g6qLBHnw35DLhzqeO2/ShQn+Vq518fIO6L7JDGEA
7HN5ANaPtkLzu2OeNJq8gp+PxzX79FSV1cW0PU682i/9F+aDwblMHiHBsOr5TniXlMqXEMH5cWXU
ADwT2XkJSSVFj2gLP9+8vS/w5P9Kd7Fu3n9fSmHJEs8eCBDOxj/cE+/3/SeTUBCArEGA7v1p9cdW
pKQT13gPTkSSKziZIdy7MGLsMWDXSvTjzC8IKAqD0YJOLVI5L1BP9muGzuRqjfVZTT7XukpLlHIa
xwAVye+kamOwgyxojXoIDb4XTl0KrwTiUngMd1HZLkqV/pFbYIhj+Bm1dklmIsv+V2Ap7u+hDWLu
zKcLHmLDn/ec0zHPz/7mcL9/xj036XNLYM/epI/3005Ye2277+ess40tBE9fVTXYSdvpjQ76gcZ1
90P7EqrgTlTyBdX78huM/HCWewFnsyJ5E+7KXCo8G04TorKwvexc9cWa3fzZ/yzF5zZFKxqyKke9
XDRwJYCYRlfJiNMSMRSMYWId9YczNGtoiesKSoDZJW/kEzA84D/dh/Ihwh1RMC2VHyFfGOTOjWU4
N64cqYKgGHlqRDXKZbVw9JR1QVXs5dI7IfY0K9I3ikSwYHSTlURqNHsHHAGBia2I1Y601trQiSTL
pA1B4/xNnz9wrO7SSCBhpRPY4WCKhdVRSCUzLTnPHEgEMoimzDyW5YzPoxc5gLy2OiE6TuUM4tPq
A7Sqt533t6jy7BsJzpAiqt2vb4BzG8UqurwPPCHyTJMhIF6/pgY5r/uE9CGFfbNY2bj1ammVVMnG
vc1mmxwIqgcQ9Di6A4H9eojx+h2C/a7DRngEIEeQ2tZGqQJzQ1eGW7S/1tKrNiG8Uf3TgE6GVH7L
3JVHNR/H5zpMMz78lA5LtqPJoAIVpCzHPHgPi9IuNBMvEgYW0Cmxt4ON6iq+xuog3bb24zArmUBp
dap3xj34qaZPvP4AcpX3+tMdXF7+NjTFYln+haHWrVQLEgTdpVkff7AF9JZ8CBVz/gzybtJ1Mp80
eufWvhnCJ4cmT9+RssNnxdMMUJsgiOyoqAnowAuPRoILzliwlqhC8RZm2lISUqXpJ1QRknavrafZ
DGqshuH1myUyDDXevRzaPpWUBUEziLRbOekv/rDLenWhOGGFasdcdlr36CGGVH7Fser2iCxyZiGi
RFwuIasj+o+Haww3Mr80PZsjyw5mfTotrmqcnBZVEi1JU6vcsp6VNfySwTFDb6ToTIGc7X8bLMLu
VfqaqVhv0gO4lnu9rk7ClnkrCoLUosfqz2l7v5S15AOxmCAetlbPldfJKn8Pp4/ykOIlbHCuXIXm
4yJWAWh3LP4QblUKWXdH2mrhm6uCzr1relI4gIS8NX01OrqkS+D6n0EPlr9tFSHxBlBzl55H4mjG
uFDA+K3LzAfi8BYk6xwym6QkpGysfyvQdRLV2gmyC3K+Q4KcNuDz9VPVMshooLDr/53IcVahln7C
sJbYbgRFJhO1jHhJ1Y2aFan2OY37LLgPKmQ3fhr1rgfgQ21yauzFi3uLgNOYmGrOxFkqF1RtAnCZ
rbsLJB0kArG7hqfRyylKfMj2WhMP0A60KgCPQ1rJsfKxtEhGO8KRJ/htFHPErx1C2rAvs191uFhI
58coi16cxwazhkdKbMr+4USVhF+K4UppmWGCHVg30Ng4UhPMzk95P9LRu84v7M7Pr1KzkaOJQ6l5
N2bnsdIFnJJMyM9QvYAHkZdEzySgYmRcm6pocXwATHndtHqk5r1B5TF4fea1XGKh/ax/HrbZPoMw
KhJOWa21ITx30wH0dTfSe4DrB/7RCD3Zpl31vQ7OYN0a23ct/pGqFwwQKVWlt9kKIf4RKGqE/WP5
MMwAAOeXN/xz8rVDH7QYhTEXYLPG7C5sNi93TCpBJHUIkbgwUYo+toe9GC2ObpoLld3dDZ+4eacW
oZnXiAeTW4gM26umQp+xJb5k/XWq2Ac7pwKDcr69D7DTTNmIcLrxf7DI+KDO1ah+qgAgWSKFrAGa
g8FxfrMd7UfNy4pCZVsA+3mr47Rwc2OwrvyJswtgkxcGPAyGkrD+Gv1e88+SeFBdHbCCCt/Y0gzg
bpj3wY32axQaYtRC3aEmkhJ6uLQJkzT2KTsDFuxq9bV0sB03dc0IT9YDCLh2Yfnu8/PEQO6bopnz
vLyh16kwlB17NDKqXEHzH4n5Evl1Y6foiP0bCzgsLmmUh2YkR4qolZwiCs484aD4VTlXcJTbK8e4
lR3VHnquDdjgCol5/38PPi2Q7ahnRlv8FPjBUbhtHIFdyYawsZu/+deWSAKO3lHhxzNPsL4o/rXS
zhXdKHSLJUq27WX4YJQixWqTcZry9xkSETidvzxgJMATDukUiPUuwEaFmfNFDWAxdCjDEvEEeuiq
NHpAgpFZ8cuqjlhiw9nmqPgbOO4X9UX2XU/AsLwcG80fUpq4GAR4885YQT/a2SZliuEyT1cVGu0Y
3LRSP05pRKIPQtY+c1H1iKK6s8YWqCYMAfCP9JTJHdZIQef8usNLEAyp8lJWE16/IGPhP3nsn8xk
VGHzpYhrzG2aPbTSjcJ8U4WAqhsEv7/lhDeR+TYaTxOUDtIKgspnX9h2nrANYzbYK2QwT2xrHCm2
fC++v8cTJEPpN+Rsf/sp2zshrNovCkXsO0vf26oDE8y+DzNGvg6av19AxustPgigwlKd4+WSu7lZ
FY8omzTAPNtVd4lQkOawFEiDm5dPdUTRZLQv6v+OWqAxYz7LuCAKgY6FKNG4FfbWNoG6/iJoo4FD
th3YAVa8jTYyZZJUOpnJFfp970ZBgPRd05yQFKJ54dZ9/9FtwJcgb+iP5IOs/4BRsyAMHYg0zit7
V3NdfBM5xLLJqmU7+VK4/u0RK95uZGcekhbeYAiHV6fYZ6UUjm1lQUQoQ4NLOsGozwb8zo7q/G/I
F9Bic/pHka7ZXHTu9RLEUvzVuXVYeR24/LjkzjYBv3Ll0rRQmfARPQJe92/0Ng5HG0MzgHvUxk+g
iVbh+JLHaWosaPp3vhjlMvHXkuooWyOBh2bBx/jJostdHYrjlocu1MsbAQLodgUjy1hwJfF1zsY/
5H353UD/OK++keFjl15O5j2LzEIRpjyN0sTa0C1lQGvMg+YPWXCcQBrRyKX7W6ykmWH/v14zYMtg
vnNys7BEKkmMF5D/p+s3Bexlv4ZFgV0tNPuXl8syBp4+jiPwKDCpobORVrnmcAk9XY9zap0mHinF
NZ/i0+GHmhMdbuKyr6Tc6I8lEGlORKQ5mhIitc6AnI8IL2tJL78agC8W2ROM+JMQs/w9XXt7biio
LftMs35t/oDocbzSdOYj4ZR7cxBoQvzgr3cf3ApQbAmLIIhDK+lRsJnWLHyTidf6nS7bvFAoZGYn
wTebwUYjKxicCMC5KznhjGdRC2IENe4UZJD7VO8Yctv8rscvw3jKBH5X5lb6t4ApS7vu35cjny37
6d0DB2LDy4T+5VG1Zs+nkZIFjVxcqKNQB1PAJXHd/K9uZ/rhRgmNKCtbw+JD5Hufzbt1ch22RLI+
Y56s8/+T99gPto+jO1Ms/a9jCNU0GkC4GYJBTrc0KfzOuUmbU1uXksDDG90OZZUK1TU0v9BE/Qlb
e5/B+SVdx8eNgFqjxzQ8hFW+AR/1xPqcy7r6is3bFoEiotZD4vpx4+J5c18NaN6LANKRxX0GkirV
f0aSUp5wudupmi1iDZ2/vjQlE1fM2zY/P2NOwu2fHMV1Hwyuz5KJP7jPjBkpluwpmLDTRoti69yO
S1wJz0Mp5deJWREFwNLx6+JbFyi2nrz2U7V445AGaED2coqsbiSS/tqpyd2uAXEsfLFICiu/8bWl
odTSWm5WSXlKEHfXDpKsaicWWGSSmzORYsAwpupWn8eyoNXd/Sa3GKiLlTXd+TnH1g13cT2SMotH
/SujJjl010rhpPkCA7os6heZUG+zObulChM+t84SnnSSH/TfWHBGGuhAmC7Ag/yyUF6oDe9Q+Z70
qPsP8uVEms0nHm+OuUlfqb7SfP6Yge5O+NE0qGgAxUUNa6iUNqtzXxhfUwMY6mwVyVeBHjgIXSCa
kO3DotdX9zXXkO1o/HmdK2llL6Gs8EzaL65eeNu7xe9tfwkRB+j9Xz+kjr4k3nSHO5nS3dzFanaA
bEJksJi79EaU3WAZUiu3lVv5hOUAJl4qgkF3a7enzbnXvtsxTYAsXnLhklmZhdrSirYZZqtgsds4
N09oNhgCBwJSSmiPiu9L0bZ7Imh0fljUhaYfD9TpT4esA95Ir+0ltjogFURRI57uqBeQ7H6IoYMi
dugs38wZ+m06q8o/GlNl9cGJxcAO0AF5jh/Key+UkPjLd+rHOoQNX6nnILliXcLt0v4P1gUKdKTy
fYLimrKgunOU/6g+eSNJxKNGvG8dfqqDA1tzDFs0eMT8n/tN9lkXZjuO2MrUc3PgdBXPrhavXHBX
h3p2s3S5vm0cMaRImGqVLhfSBXlo0r9/LobexVwE7jxcvLCX7iUKTqLaQhxkl76MytX2Q34r2IpY
1do+TpzprFiLmTpAR8BVYEU3AT0RdNnY3Kz0FSflhWIkGyomYFuKgrO7NU3VHbKPptW9CIHaIqFe
ZqBUFFAkxwqdsTpXTvdpI4c+WJHJOzFFuYTQzHWFrzoj0G6GES82bFtwX5Jr4/g36whky6j11Gpd
40S/lE5ConOSmYYTAPh1WUGJgCO3lsaA+Z/IDNF0/UTgstdD51j3iXiGJGM4+I65paqUeRGf8ju1
fKSunsOM2DsWuI3gjxvSJN5BIAHppvvKEPMUGAWEyF2mw4C4j6L8g8WXMinib3OvyMyUwZ8pHooI
GzoStP3UO8nt5nNxHMq6HBbgln4g81G/f8TxpMIKRdDSr4En2r0sqEHRjWEb3hZWmMqIrdkuIcV0
7mfkXzC2UoDGzoEMXiJo9as0v3z4OFc0dCO+axr4YOlVgtrJj+0nJzJ4zGdFDsUgIS+6vKM9lINJ
WK5lnavDe8FMbndyPe7py/tXDUn4+Sm3VYVV/SaNffKhkZ95HLASb/iRLLL49OBC3Ew9AD/94lf+
vkguWhlFiQi/8OyUks33Ishbnixjh5LRUdtgi+ik5+u2KI760EGgNF3Sbw7ZagFP7TwBtciOdvYf
p5HZSsBsp9/DD//vLIhYphrB50U234lz8v/FZxXjLbEq9KMdBkpawsDGrfNuE1t+HuhKSuGubNt6
AAocaxUIC3PFSrdy09disoOEQO7M7XaO4h9eDqgvFgoWI/rypxlSJOMOVlv6AYgZIdJ1KeFulT/a
aUy5l4N+tVMB/m4qgLX7C+q+jNHY/1tfxBWee/kyRK6xL5E2NhAhVHn35vZfOnd9TsDleNwOyaji
g7jq6oSuT+diJ/wEZDcPOWMH70Q5Z4oSJJeNTV9WV0m1RodX7MDLFeyz6/YWeXxZQk5R/An1hlKt
fNrNhbzNSwNA5YnNUCcI52XoKnukYxcPgw7QDDjsctrKitNOPWF6e5PqCSQhfPXcVOnTsOgVoWYe
ZMYx4i7PgClekGUu2m+rlQqSpymXBOo8oBQbl4xHdwQIL7L47b7fGCS3pPPBKrq8ZuyKxtJA2FXO
j1xw+2i4L2QAIIfIZsgPgCtYO00maG093SkXRjI5hmOGKsnTFhGJRyfJTBgqipUtCmIvz/sVJn1T
98DybXRunp3ssjWUJKFz0Px0Rjne/28uqitc/V84Rdaer3foLWrl54W1zoO4Wmt1zXHI6DJQ/nJO
+AefRBeAcV9VuWi3UbvXVYmcDYXFW8aEOjgKCvq95Av5nHfcgTNkFrKZ1igBZ8F8ri6//OUbBkSm
TfvjfsoNkPEwvNwGHSrFKtgKFIwtOxInXWqCtFERMfsT+qQ+9KcSkPov+QZzCIgST882mUhXpPgl
ti8QKUxOQ35whXA2TSoUhYmQ8rcmp+00ZlqaQDRCBZThc0dXVlQvkRn6sSDT6cy0etma35AVzD1C
6pPEey8jfDbuBOc7ZXf6WXRWEI8ZiZtct1OTFbPLLCbY91kTF4pl0IkIOtx6b6MQWRV1rte5vMzM
wGtZBMnbHi+ePywb85fqmhaSiiIEeufrwwjRW1/kX6PyuiPYMgEfKChfK21U1kNrJ8AcAKTMtWJ7
xfzoyZmCdWYbi2pmOueK1/+YaiK6xv2cfhvtmyiQr5UKcumV3rKopZ4RcY6mKcrjTizvZZhCPuiC
U9CcxmnAD4SeRQCFr113XUfYIr3xhNzBF2VzqD2orgodrfyoqGzOqcCVpA7yCylpejhqDsAFypR+
x+8P55tQcXMFQkHU7lDgRhf7NFtxYol5+Md998YiO2VnzWm1WRoGApCCBCc+T4bnSkGw0I44uQGq
xPXf5gp0nUxqvS6dzqMw2k6CZErXsel7bee4DPrmEUdhdA3B/10Yi5c3Y8pLTNl5p00SZfyspxR/
yhA79XErv9oOvBrPA7+hq48AuTs3/noluk8VbwJDNyM/5AtVREuQpUgn75z9DoBuBCUaaN1OBGYS
fqolqq/3zqZBJFPYeKW67GSSa/bSFJXBpI3d4OnCd58iwtraTMCnwb1/y6ioIyiddBK5spI2CNqw
jyVJaqQin/GBNaGWNe0CZYBtPG+lssvwMh74RJggCI10BLEO04ZxGhZw35dTeacQh03/oJqEZ0+Z
sD+YGHQyI3d9S0khQTnSaRqdDmYN+Umzu/U7Wti4yY87KJpKfKadMmBv4PQNmPQTg+Pi6XN372bL
l1KJlRYr+ckSv/if9auDwNPJeL7tpKxStjYgKmqTnq//lmv4OExry5DAp4nXBJbIEIcYQClLvmWg
efrH5WGJimFCN/iKSU6sHDekw+r1SL/jqRj0UOcLZEXgHrGYOGbAx8aRSsJeuNkOARqdXAeBEIX3
BLW3RjLBv6hxLKTUMwqOxkISITHy1nHRb44qwFY+fJOCJ19kpvjfAM35ylLWzUVRIHKj9UwGzTxm
d+qj3d6VZaWTB2qHQeP/25bCakaY+bbq4UOGrwsITu5ZohBx7kVammuhUc9wUwT1V1PlLW91lGEs
+0ePxMFaC/BvuqQzaM2rceleiw8qm7YRWggJd0t7Bwve0LLSVunF2gbYa2cMuatfDWQRw2mq73vN
OJKIyq7x6njLRcldpZ1NZKwLb0xybpepQVBbdewG3cT59XL7OgQHlFP7h2ApmUTq5KUccRRP/N51
+Bei4wRe/RfnvMokR5ETewqwnXJSgYXkXn2+PqqwGKj5qtRvQcbcFJvHjZqSz/7wFN1cGSMVymIK
6Re2eG9yPaww7JeY+JcjifncdOQJGd2hUlcYMuAM4fRGXpi8AoptU0n5iMRZ0ZN9qsEZTF/RVYc8
kIXgm5H+5JXYqFhbdS5ii42Ryn2dAosgJ57+hGGKTjTwiGppF0tF2Xei6jXtzO/mL4cw/nq1q0By
w+1GL8d0E+ut8OOK4iUpssiDp+sQjSVt6q55ynfMHrJWWFkCK2OeBNTGU+fxConTZBBW9PknEa9F
P2wOvbMueDk2MrG7qLozEyJt0XQnRhkClg4onI8h9M03Q+GzDk92B/9lajmcq0rcl5P6e2HVCdkS
sqKD9icpsOPEmHecJZReVnuUahM0XxYxAhrT5RTxXlgjMylbHJnacz8dyLVLdj4zDGtTPc2GLKTP
D8pUhD/UuTva2lYjy7rxYdH5OQqiNPHb23/NqEXxY7cDuJR4FrpXTKHvWSq1vqPrigTqlF4jh6XJ
8eIjC7YZZTB6gwNiSu6ep8pYRO+HtIAR/AHZjGgP+BeE4vxtBXhH2gtvxmd5xBuP4CPvl+q570Wi
OU0YWEOhIfui4D/RAbJjcu02sbpWPPEngozNV8KI199f0sK7SPUTMC8iGQSN72KqYSWIfLhU04U8
q7d+PLBikgqWUgeVLCrqHrUNuymkJh4kZH5x6P9N7UtO6TO/Cbe0l1OFMeX2KCVQxAJhw+qnGh8J
CF10u3mPydYYdjXR3l9BsB8xyYbdV/8ZqIkLws0NMIvoC9IScjuhY2YGuvVNci1YoBWst9XoCF6H
q747AX4VdincoFV997GYbUnEmsYn9GODRwjEbuoiopWGnPdMpZ0OQH8VdzfwD2jT0XCHjDqgFcd5
8+nI2xyUsYAQ9YzhtOTwUI2A0HhXpgBsO5loc7P1/Jqe0AJVMs813IbnhyV7Nwxr0emaQ5kwDApS
clxgJjbAzRE3vFdto+slJlQhHGjTFu/YzFQzykAGjddtRMI7fu+POKqIe2jQvTX6oFchGkbvSNVd
/SLv2OatdExbqjOR/pRrWfRsAgQF5W8R33woZn0AJMGSM6vTvlmQ3uNnajGelRk3sXlgBYG7P9WN
cJ1d4bnfjkqexFWd6DpEnTGK5TJ2UZUJe8iBlBiPVGQKO2yBzdrm0M1TihM8k53th+qT1Gfwhy29
yoI69htDllgAYF1NKkd3of1U03e45uWx6gUqmJUiW75p1yyuKW4mhcGmXtp+Ov148kRCGowNOwmW
+AvUoKWuZ5AqYwecjFpSRMn/oy+28dX4SArAwmK3i1I7RBUvhNp8G7joYdxHtfsHUhQWpfQivGCw
QJA2ZJntwaQKis6QadoYXD5kbWHDxOiXQHPJtVOV1HNVfOlZWFhcA7xR6ER1REfjPeBUDnnB13UE
kUoURXlSAbnB5lf5YbqaXSwU9oVWAm9IumhWIlqz6mjtKcuN8beujZaOtEIGuapCNZtPHMw0INhV
Jo5OK1gaMRsymKuHasDIqgZb3BPy9c4gXxjkUAxW6HHd6g1FKuNSpMBOE6X3obiX9vwpUHiINNG2
lIV+XjzShTxYXlFJZsETS2I9fS3mt4FBRwJbEt9CKi7gVOSsOhZhvj1vSmmAjuXyn5HeYzMsK5AS
Ae0hpXY8Hy1SkVVQHkKQYTog/wiIrMnHgJr/UGExpujZi2BNugz/iHr/mcp9G59TKlCEl/y2Zb8Y
M/oflqEh+DG086KFQ+9YeocvPdg3lTBudmxoD8U50tJrzXEyQCC8BGOa7CBhLSNA04jAGqgwixSq
avEEoxEK2wo/9vwVn75UWGwuk9vSQFZfSC5Gjf8pzfwhgKDvgVrrUe4I0+qz70kq4hRhBKEPnMTd
pwmqv+pEZUvJK0ogcrKMHUkxvZRZP/ZQF6rnZINew3HoXmpIjnPIDP1aQe0JkdqNALqX8rCE9/sc
bHCRMFz/SomJxqOr6Sy7zz6UHirsSesRh2c8WazFYl+HIeXU6SnUZ/33BlD/qA4qc0DYJPYYLVLp
gT56aYbdXu+dKiOgbYi1RVxap16AGzg/WLvlrVqn3UfnxWqYTmjM7/AMMsAlcidWS/i6y3JdZBsW
2mx5wglD+rC3xo1oozERY0AMvXbQzNWFnAqc51woRmj3f30aVdAozDGJe4OzTA8Sk1yt0MwJA2U9
cS9vvY5fS0pwja24dkqxs4s3ip1m59myJLeoY808jnnGeS7g9xmQQywwtI14B2AjHbb6VvbKQC31
AWZOl6O7nJ7S5O6E9OQEozQQfeceDE5BjIGci7q/ZXCsg9pOyTjErrOfkiCK4jxjqYRFp+V6Xfod
jc3sdQrCNOT3l89DH+YpcnBluFhwdvCvD/b3Ut2Z65oTvgL/F6Q/7JmybpbxUWzlcO0Wct3OIwnc
R/1g4vrxH52opSkZrLqF0J4IkK7iGUkA+r1EX+dEUMYy/bgmRKLRDN6hW63T29qjxqV1pT3sjcrA
+q7JfnnZIvsb/vIOLLb8jwKCjO1OYXwpED6MwcT+SGLnh401VEHysxu06bSeid8LNrJ6JmCX2KMa
6gy8zKL1CWxrZ1Pqt3QlIMojJdwkGryEYrOJ2ef/AvEhqG2BiYMdrIMkYgXVznsRHdetxqcl2Ywb
G8O1oaDMfzYI6M4MrsOqIi49KWkDcHfx9aCitH1j5pw6Zh6oJRlOFMAZAqM4Io/MGii7ta/2MdYV
YhpnEWpZ6a978St6gOnEifPr50AollZo1t62OuA8qdWA1BC0eMTz3NxofPCqcYsnu6Mjz1aduEhu
RrF7BEmX/PSBe5xsG/zE6Y5BYyCoc7lfFbqAKUiwmfja5h2uwv+qksgzK+FGpnjexI6I3Xd4vo9y
/iOCuqZAuKwDurAgE/vqvvVUJyk5ggcql70G4WNlddEhtsiVKlIZH2ac3ZlqT1NHNd5ZLjZcnDgH
CMZr36Y68NYnICgzlps9tt+c6qOZKI2hCCrtSbRI4O8dm2tQjE9u9MCspxxjo1QMTSHr19rKXEbp
UbCuNCUlEWNp5v4nh7XQycJMlv7PmHhhCNlTmD0lLZ2m05M3lBIC8br4HCMwhevsFEk5ZKON/3+d
JFKirAYRjOMiN6JZUX/lETU0uskqZkxWIGWYdqQqFn3iobnYil+/EIXuN0mAUmbaIFkaiJlY9b52
etoIAaCzCKnjNR3lbCl2wAXlEn5i75K1IPFLBxbfF5+Lwaq3+hiBWgjEAJJhi4n0DUeuroHK0WGi
G65PymWJF9zCVwkmFT63jHJX7pITXzbYvHPj6ApgVfLDOgzu+4NFpjXf0Ba5l7iRDk+Szrg+99P6
+CvBKAkFWHZk6ZQ4Vqv6+xgGheQfhp7AV66dmYjIUKpzJvuAwdKI9YQwHIVZTxLePuv0PZwCpJfK
bFxLstFj5wUOZ/Z6Kyre4QxRqNcg/zCz2ZutgtVcXXWrC2erQYCnVqtx8UNnu3Qx65q5bCU/ofkc
WzXy+MuCx5NfsdAf/Y0kblm8Tis7THs5NFgKu1cQMTj4K03tJC/m179AU75qmnkWYTkplGq3k+a2
wlS45kpn0RThKbjdXqaW0J5wAV8Jr817qSQmNgdJYMuE+kU4wPLHQXLpKvmXtK611QY/U04sFR7H
2ww8xBt4p6Lc2QYDiMpXzoQ37uDfh5TxpAK47Mjfw15rnD2TwsxxasEwyOpVFc9HMfd7IkgVQgr8
hn5hxAavH/bXNLywz73lG5Pxa56q9UYRuDaqC4H6S1ZWqdSnrdiZKeZ9BlKUYnPVJsiHd4EYHK0R
cRF10TklPdIkAZJvbnwoXDqyXe/fjay+O+YqHZvp0sDt8mseWaKGhs+JLxAv4pxNAI9NPwesFm9U
ptqvCLkNWvlSr28BaKT5cKmExJVQ+XL7cKdt0+jCZ9YOUI5MPb9SGfYCz36JhAH/7laCo1AH3iL4
E/LFSTyKMEAQZhcnq2wSINIJhvNnyKAF6iGK47JHMEnPh9CyrUq9jppvPYiE9HHJ0TkQoAb1ledV
Ak4RKtmtU85DEiJkY0IS/pOTwBctvx0GUmJowf6l5NdlQDoULUCofDKKcVQ+Zt5yxnfPKAkM8iS2
1EnEyNuC1rdhHk9/jXYTnRzIeAyYHci1JA8uX5gNCHa+vBhs/uX/SOHwVC5iFcfUe0qb0hhYP3oI
mNYNHiQC+PgoLNWIlK9FUlMDpTJ0s7dv3d3arflWpfw++/fwhVakN/so34DkbL9HuVbATaZdyTfE
Q2ViaUq/SfBsVMZkCfCdSJLu6NnyYG79+NHu4ma67c9Xxq1YnUKk536opEJn63VIPr8lDxW+52ZC
l3RX5WICkGFS1O1elB19xh4w4JnRGropdnMnSGMvetJ/sbUJHW6eaXtnF8Z5EU+PwTKxoUlQhof7
QjMsxA1trAdy0g2HovNiIfNOemWl54bkX0n+Ffq+G1LOJ2QNlo2E7NQ2Afgrkchjdq/Ylpn9c2Kj
5fY/+6YbR27RDd2Ddq9wLLc75iapit88JxPqLDE5mrq9VCIJayanU+If3Qt9CDZlu1tzpbgfwm9c
kqbwmxRizPZ8svK0ao2oFL37Xp/g12LmhWxyc0CieQYV3TQ4TXoisS3SABDZeC43QUuUG0Bq59x2
dtfZKCCReJRdf+YDr3G4PHWCTaYylpVsVTJtnkJF8cyv9uSfsTZgWpG4BBpu0amQho1PbDqbKkq4
xEeRiMtq/597Wo+4iwNstenS9utOxtZ1XQM/Qg+EYn2DoDFjHe3FKF+UkM8ITQZK1QWXSXLVxSse
ep1OXJmMys1r72SK8K+A5h2YL+TbnEUgUI4QxlU3+aPGOv4v8J/sKQSy9UwChseF7AZux5NVwBo6
ec1BXlyjfN+znhja/uCB7W5LsRhS3A6tSBthdHA9aCTKg0oVpBDosBfW6mw7ApLRMXKL7XRFwWK3
SIxgzE0LWyyVHZciALYnwtoYipAr7kRg79dTJC9PP2cS9Hbr+nhQxN58YJGqjrVx2jtEZGsMNnYh
vKnwKP80MNC6O15DoS6cuStHLMab9Zb8F9SWOmWnlAj7/YLOFfrp7V+YRY5xHDwKtHREQU0Yx5Qs
w3jKI2QEGc1AnZmjaccB+GVY+S3GhDxQyM9wVseghZFeA3S3YcB3g0pdQQtBVpTeiwUOg4Z4/kYz
L5oQW3NVrSjlxkGNuzNni/3VGGPHBEWJi2VHeioUaNfkfEX7NsOuwM85Z5mJNJvO0izYnGql5Z03
j4NsJmmCav7MxiOqzLNv273AG+IUGi08be0siW1r8cNvV5ZAWXypeH2Gy+6HnpOZN4RL/fqcZUdD
0WyJ3U3qgVvmMw5lWpNlCkqH7u8OgtmirZeWQJf5pIBUIHVfrUHfd0UcC63GFST99SukL5lQt/SW
+qEpmP397eEIGOwJVWS6rUufera0L/IxxnCMAZBFwIV16GkAP1A/nBPod46Oo0Jskzi45JZ9JZmO
yYuKfBO4CPrq1vJAQYyCffq/gT8rdZWXpmH/KqObwCuqkFGOO7rYCEcjeOlEeW0LQudZsMf2jOiM
XOUrs2RI0wxxubJ4zE6SeRb0KEvanRIQfCUgNJO09pCVyGApp7op5+0uBprc9Vd6JtNuqdqghtYy
W0e+jgQFOq0eLIguXtDl9R4de4bBqIuT9pk0hz5Z0r3mWZ83j+Tjh71NSPDo3xx+W95mE6LbJm3F
5+C6pazS1BAd53uRlYwWZkfbOVCZckTTd8FB/7shh/cxeCag+xFKAHH6swlUZ0kIniwjnU60JMWp
+Pjl3CeJGx5Kw9MgPEFzJLTE+lBV3RbUpu3kl4h0MZDGtJ+fWZva1NaWPrDLB/X8IPrZMMSjz7KT
vfARfBPvwlrSTsAs3QuJzptgUIP9LtJ0bifxl147A4YHYFZWfOIDGuTBFvrIXk3DOBDngAt1dZLe
N3Mwm6ZrikauR0SYf7g4aKkgHh3rrH2wq+11PYN9nl63h34e8tdZwvMtKm62MD1LU1PCu0ri/kCF
H5EszfJ+X1oTrqLLjjhbjdp+YItzmt2OkVSp+mTr29OHQumkQTgpTPnZeJ+dql/cpGsR3bfwN/t0
MHwFFrYpjyQyp8wNCfKl/DlPe+Q2OUbx0a7ExpOhtzQ40vLH8qfiLQYLtoH+xwz8SJd79b6OXQU0
xK+KbQCgb90jLPdglpeX2bhUJW6gJ2jfcQNyezay1YQ68+bW1OaMIirOwpS7pBL9zvsE1Mehc0vW
U8v2tSEgGVvuds8GDHip1bM0gicAjmeS/UnFl1T/AvOlEAS9Xomegw2n3WzxUh/v80j3h05t6NPt
EoTePmjeFd6y/MDI2lVTxK/yAfq0OpI5+lzl3IC47v+YDIOD7bkh+HyrK7h3MCvgU4iyeAVX8IvX
BgXc9m9mZB2oqcHfWVk4C3Olkc2LaD1KSiySKzcsBPtmFPGDY8QFE6vf9Bgop8JZpk487e9TpqTX
//39CwPt3eFqzKgk2q5CLoGgBrVhzJ5Fbe5iVIZkrLqbk4jShRPTHhQqJZM8t7pmshXmv6DgXK+c
V8x2Gwe9Fz1S5A4b/LZk+UMhf6RCcMkTRrJIWsscDo9885bjYGHXOzs48WyAccOqKvB+hAsEodlB
GhlpfZgDeHjXQac+cEbVx8/2ex8bI5fxRwtgJSH8tYWaZnmguKBmT3/wI+ZoCggJ152DW1+d6gMl
tP9gYu8WmUdXWHIcaCJ8Z2GJ+VEAYjcMkxN9h64G1OEoWeF9e3MvY5RPZeiUyIQzoP5euBSDVi3k
qObqOeHz2WtS4cqRxSrBasMHReK8vg3R9y0wz/ZcuP0Uy1qsRFtRgkpdPLsb0NB+sjcIL2wJdAhT
+V+s6ZC9HtcIgbTCA/5Y8qKEZtXg8yRr2d54wXFNd9SDLSyFMAlWSSOWfMMuF57Zci/ELZbVLP7V
u37tDtgk9Nm30mrs939/ZAQNDildlW9rNMlGwp+X5wTMcU4hLnLpay9hDSATxg3EdCBr0Y4raaTl
uagHhZSbJWaBPRrcHUh+bA4jX2aCTqdfXqeGEiUVhQrig9shfGI5+j2g3Vtzg5GeJrT5Tnuqc6+B
yGODq6SrBAay0nwilWLEPoiKcRAw7HqIHcZNzGsXj3quojPE9+786rbQ8pIZoP5Bw1sknGg9JW/W
Ji0UGltLCFkmOUbJvI1QOZloXGWN/IfLbMXSVABCYDJU0J81pFUJ3dEw470G97eXLaduT7+/4CXd
sZmSthczFgkoW2imj/IMBE7BcPzx5htS5aRDUV5gNlBQuVEzGOVnn6XIR+6QD9oGrAezuVZI6jMj
kKSP9xceqKvYCQBqDQMP+W34VVWDNHoYtJ9RAETHMmFJf7Jc3Z6wX/GpkvoWrXKty2/ksJmqBPvQ
nG/9MD93gmk019IRaUFddLDEC4fInpSd7vJfy/+ceiZ6Nf34knXSk603Pco07g3VMHCHVPFIW55s
BpE+6RQI9Lt5yNScNKoRKHZZFp2rvVyHoFNmJh/U9sKZzYIi+2AbmCq4xvFPow10T5UtVTw1b3fB
057TfFHpKklzO3MPosGNISxNti8diJkmZeYeOefc7lg5W3H0LVLWUbZeiSmtbrYwWWTsWGYyAH3P
pK5c+LIw1t7VUM26709PGtpY/IaOv9ktbgokdgFfPdZvOonmFytC9tykoNM2C9Bo+IwuqumiUl8s
WLQcCwH+Pi0AW/TTjPzu1+NhXsTl30KcGYh1L8iwbF9W7uGzN+gwrSz4YJlcnF08Zssr0nva6w/3
T7wjm4KX2eG1HwhF+KVG8sj7J/Y8GHsp2XJPWrY6Y93i0NwpN/4BmltFIGXRJE3Q2B4D8rkfPYf5
uAI7SH1UrJgiRG8iiMPh+Hyc4OJFNYRNGoIRRKp0Jty9vkIuh3lCYv0ZqxwtmpOOx+XyFh7RfPEh
8VjGG+g8ZoVRgvcGdsN+v1v6fg6TEupAv5JG+ZsBSqpSZwMYXWCdvuiaEoKX00lvTNsInN4XeoMI
+8czB3a5Uy6EJxBJvw88eXsQ+IyO0U950nUO0p3cZW+ofsftFW0jYfyTBkqvOIdmr+iKPtd4snCS
ycoi8ttPNz6zufUgxFaWiYZpBLICdLShLpNk6AHckELSy/PpyXZe+RnCUcndIWk+u3aB7Hm9Esjo
i/O2Ff3pl9QitR/gewYhmQ/a5jqzqoKd+x05OGEYrc+H8/w6U/+rlh3wevkkg/Wn6/f3Exk67foe
fnqVAPc+yW6C6N9qpLsc+J+JfPkNzD6688x94GTZghQ2F+/DzRCF2WeBTvmNGE/QNG1p4T0L6l/y
0Jc3vagkx5dI0dWtLy+BnhQzuS6TysdBPFruyp4uVQeYwiwevzgOFdfRWTn/Y0zNtO1u+lQa+b5+
cQWdxgLjMhlf5+R7myEABvv/U8VfuRhRchQQRzQtdjxfpeaxbgzeWJ3rFcwPs/L83EIaBk+vlFau
QqBOiifVkjXrcjHukUQMnUj+Tj92vDIZDy71EF49RLigcO6HUF5tIwdIjQqSibl/I4fFVRljg/R4
GO1KbDfl1rvEyXIgUyQXIHgoP2tuTS8uUZzTVjHNnYFOQAuTBsdp6LCMLhJAIyQrDsn9pVlRXCtr
bYvIBYSPJDhDTKXt3/3nlZMNTizdGTNceTPsMXv7E88sAx8qoK6vnLN+r8ThK+OY241NiM1tiWcw
wZUdha2So+4um2PYJMme8ED6+qVaB7WfiEynkU+FNPdHb8zyT7wAPcn83hwM7EMIra+CcgPkhUSI
pkk09eWVeDfkYj5NsUQLQYyWooHOS31U7h0fIkrHtXRWZcaMV+Qx8vgYjQELQVbZTWAvgEDyHauf
FCtSGn+PztNMUslG0qDo7wuVjD1cUHhRCLEAi9otl0S4btlAifMi7H4SKkfXLJiBC6tzVkVYTqZa
IwU/Dd4SXrt1gGLBVNZwUdYz3jngerHg/pH7lORQDhAguAPctwAf4CSCRooYKEVSLFcAmFyhjjrX
SRcCaGIUKAwrtnp0EtTT1+MEfRMMkZCnYAcQdm6TPc6BU6gjrPty4FPsbI2ypWv5Y/QtVvSvEMYX
jDZU1ulXl2oShm6zJVrOw0wQXRLF0YPJi5w1yKplm058xV/F51BbsElIj9BMDo9G1VTWO5Z1QKjR
9+gmlthX7kMU7Ge34+A2ntRr32WMFzv0BvXXAmCRXEG6wTb5yUB8cCX8buxtdwxfMIZbfHuus2dY
GyGbp4rilbzuF9ud0QmsYbS2tjBBlhoYFioAiU+bidIss2ZM/sUmPBeiKlR+/WUU7Yw7I+lAjOQz
CYrdNUJfpbQxRkC2RRSSssbIC1hruheBWF6Lor45DfELA+NGAVDh/eFsTHyVBsOZ4r4zcUM31YYz
7k5Xmuw0GC7Ux3ERJ/dgby4PF+rs9OfSmB8oc/F1mPgskPJ4ASusIWLksILgynhl5ZEGGpUxfTg1
q/CvZlK0wiJGlACMYvLhkCJC7ioH2lHonPKmRJPMA2Noy3ILD/DsAK17KwlaEhK3RhX3QRNAnUQI
sWH3N8rW7+CTzL5Ipewp1gTZObcvG5jhlsTbNhQWou+0xbLLyT1NJR8+9fyq9Ob1mxA1x2E9TuD7
FnSf/dGDW+4gEgI3bfCclzoEiyHtKw6szzciVnDBXKxdqRqAvyI4IpWpiTqddvPEWjHb6yn290/k
7yEkWWDIffuzXrFs39dU1V3zdAjDxTAc3IXyuWnHJO+XpStwKIMj36IGjmaNW0EmcSY/dpe1hE0J
j/odtgok9vwH1+FKVJmV7bohzcuNZGq2Cfz8BS28vSJs7AWxU+zAUJ9cEXRU4R1a7COeec/TVpT3
G8n7iJYobViALDv6/BBdB8Pydxhab6h5Xlnwp+D2JegL4MCuhWgTbytdmyN4vTBqAjamu8p47sP4
9+Qt+4ADxnc4ELWaX5edL8vJhXYZaLG9bQHGH2l1TU0ZU7hPp998WBgspR4msp8XsYGjv4d6Twkp
8rAXwZcMNYscA/guNqvjAzRSyMCHI+OiCDjJdKqrCt5IbkT0Tt5gdpKZcIPOGTD/GmxnVeA9Ko8E
7F3u+1oFgz9apDAzEmgYAkVEsP+kVSJqoVdk2shPstxWPvuiCZiedniv4ijhGXr50+7pUEbDPI9w
NgptV1EfWOC2KLfr8JUE/OzSCQTKmSPeB7ankpcDJMEPlPBHwf98xoAq/O2pfOsQ3WFxKjQ6fql2
Qhcl3HEMk/pxZHHtLYDsgL8B5QtCSPXZA2FKCSzQdyzhaZ69mVxcZeZ7JzQgJmcM/weh/Yo//9TH
iKPGpBwL9zPaweuqfz/bttdkQBu7ykp8jtFS1Q5WM8lSpYI4aEl07CQFopCXBySNNP3JjTI/ohv8
ndPaRXglP0LqigIsnGY5CH3cygboVCWc99gWC36SWPuAZnx8MbfonTbFNomGzoSdSQqfgsbLNA/U
9EUptxteUkpczqQnLtnwYjtPjxxUsU9knraV9/sTOykGezzqZL5INmf47EG5QyMjh1/gfj+tW04s
NBYpLuM4E5KrnT1kUOT5IOh8N+TdS2+N4Q41XkExRWzkfcjzHAbx1ueOj3w0Ch8ogwBd50kcSyhp
XlYgQr2Jaqy19N+uQ2fGdU/h9t5wA4ZUExb/eeytm72FOPhet1PvWv+abY2haFRm46SfIZX++Vxf
z9NIsvmGqtBpodQZKr+bt7wGCVT2Af/k43j7M8cRdMzlzrUMKU6XSNmuptfrTjHhHs4hRIoB8mex
B+hcUWGT+gxBiiZVR88/ngTZYViIOVxdBNshDTpIlTAX/4ZG+HncdK7gmJ02UT+HMws/PTFNpF1S
N+fcnCx+XfWt4H0CmNsa0ocYUGUywzjJvuPFcAJjeNkdEXPsLmy1Gs60M02tqiNdvL6EIb9vmdCe
AWJns5M4S5xSCkWTa118qfSG/NjYxtrasTqEA11CGEpWsFBr7Uy7YtOCfXZJby4i/sXfD3C6jyYY
wOqtQgVD4e2NXhinRnejWhmcekEnl5XemqP8hukC0ZbLD2JDF8jgJ94xShoj00OSzuD0fKHW2U7u
IzJLbnMTbkPkpumUliQad6CaqIx7VrZc8zSYZ/c7kHv0TXhEUICrog/GduxjFaY8/U3OfcrpsU8b
k/SgtTKYCJ+2uIRK+OS3/VvZgXdBrrgFHWcwbNxCtctuNHGRKg5cwtADjg5bK+GMBJRujwRMdxSj
adROtLebsb9UA0THMEeIi/ZKF2xXXQ7MOFAX3aMHmarR+8kbqT5RHbNRZ5qT7Y76JRF0FB4AyGHq
Mv2DeQoUwrjTLbmUdFZwelASpXucZOZjcra8fVkiapsAetCP69rdte2zkUm44+HSWC/BkAVJfKkj
1miQPeyD0KSxtx4iecBJIx+QUo3B39UIwb036vTm0xpleB+mDsyXOaVN2f7yGpwwUFoIlTyo4a3X
9Ftz9hPbViFqmAclOaacYR2nx/OuhfxSDp69sBh6fA+w1+c5up/fcPltlneA6X9mQn64KaugIqxG
lquMC3dzOdoy02Jj0zcB2Q9RaQT4HkhTq/5rYWt4SpqqBNZxuuGLM1KaHkiRAG83saV48WjqHiD4
lruMRYKNEOqL3JRo5F2XbbxU4R6aAvAzvMXx1R9C/g67f9yd1JomlVTFdESxLGLLYkSO+QDJ7ltE
FesEhGQ8edQWGGlb8T1S9WQu/zuEynB3tH0ZWz4Nki7Cw7XoBRhxwLc+mbNz+2C1T9qlcizGDr39
EcmRKiTdwblsJ+9ITwHAuFL6Yse4+45ywmWjHWZyad2erDRukB0OW1DSDY7CXSZa6BwNMWlCZWV3
wMXgvcPRrTFr67aR8xcyflQgI/zk0dptzj5Xm3asxP7yicEFhF0TlIGKcIV82kXcYLw4CrPz0qUw
mRpNjsJJWTpx6VPAM3LnW1bzWBv+hn0vBEu8E6gaFd0r6fvFI1irE5AqH0SkC6rjo2rWNDaBty6p
Tfc4e0y5Su6Bcts+Ok1G1omDNAj15BDBDwxe82W7vG2l7u8ZSxw8Fb8vtgPsnnbAGu9xjARjLSi7
AItuXhptPEYmCPjU+rQnwGsqRVIvxXfNf5wxaADqDCQWlpZ8Dbed2OsM2GIi62BKIPD29ISEl82q
xlhalNaJCGhF45A9o4tau1Uc+Pz0XwWxD87clQeJRhp/vMXDX9Gw5UoAo7G5OpV0OQ5Dw7ibi0+/
Jy2wSjeQ3l16HG4AadhKqPVO5FVENKm2yCTPwvN4SlXr3sxTcgfOIRcwMxJhZKIIgUCstOgQ/QO0
ORlhNruNU3CGGuZVyWLKpEiWwDLSU0v1yLwvePyGnnVMQ75JtiHNayiwnKoFLqgVDJKMVzCMcxuz
t6dUu1iTHd85lLGx5G5Br1n5EImRvEd3FsqUwWKVOtxsm9r+p9usK6x/m5ZcSqRpnL8MjCu9/h4Z
NXVMEcrspVntHsIJB9pakN5cmr8XQ6HNACW2s0+veesrud22H7RgPAYWJtroD/X5xjWeSXaGA6fR
waLSzBoIRPdx7IQpMDpDcNK49hLcNS8YUczuJgqby097Jn9PaK8zMzKuXkoL6vA1TNOGF2rP14qk
a3NThzCWr6xMCsXVOLr8OaudAC2pt09hg5SK3NVSBMXLqWfBq7ENRn5LYDN4/t8RgZT9LIYe3JVg
zo3UybTxdvytkV88tCzM5fqwxq0k7nyv37ya7qUaOzl9h61htCYJ1HV6uRkD5vSUNs0jwpbaFSbw
TvsOaPRbD2DMZEcDWbk58JNvUKijcvyTh/i+aFZ4THi/0iyffPLj9/CSlLtsq986zzhzK0iWhmwU
hKXabCl+raSUDrYvZoIgtjQXhA0beYobE8YTz0FaOG5u7lu99l6O6ghtqCk4cwQX9esKG+d/rES0
wpkuSasTYBD5yZex0ju2VWZ/vnhDluCsc6/uYD/5z7FrZIMwbUXEqrrhInm4+Q+aGmlRLq0ZXjet
Stznkk467Dcrs1JkFczM0LKLeHLcnU4WhbUJx/QhKC3odytCgUDRXBsA6F7jXrip2aQLuisljKAs
la7FIAIW+xBqQqCrqWRRNgWE9YSsMreLxCb9gAaDt+/O8EXQkkL/oYAfSoOGaQcqFTKJXN55WqRT
ghYZNDkon7qbFwKNrhJijS6yRpu6zkAIcdQafzc1QgkrXL65pQNZgr11UhIRxnNYytBvmqy4iqn7
PwSSdQsE6QNW/jhV4TH3Qq3SVoanMrjAvDFyRkH0QgcUFQWReP3+zq0wA94cHn9zSpvO90qyeLvt
JXhQqU2mS4+4JK16Y5A13HbZZYve+6hZMkLtJy81+FlcG0twjD39BJOT2sDz94PhCAMyQvSIfXjW
KQD/L3ZXfV27Vq+OFzmeIVz5kfnG82Yuwd2R9PZSI/+z3FF3PfLq4Zd4O7pYoLtpXMj10FNepLSp
NLh1WuzyfHTy/ebB4WaS+yoF0c/bJ1e6aZx7io5ZqcxLtn2MojoyJcLMyVgmJm4PipW+GOAXAmub
P+FbuTbVv7g5q7/mKlJF4nxICoaOSocUbyYt1kt0vHsbhgiN2GI2Bwr7SeFA3V/aD4Bo6p9Q4oyJ
2hb8D0yzYBlU0Zdu5jUvzzfexPIkx2hdndmMNuzk78pGkAwEPXdVizuM24t9QjxSHNaSukDOtpzw
nwrQDjnEB63SAgFEuP2ftHTuMVYrlM7FwbIlel84ioOgwdaPONOIrBuqZGyLs2cn7br/YOQkj63W
Fofl7e3AF+xLSIjk9vCoPDM4eWxI0y1TjqjltJLGooXwIOTFyj5F6a0UqJOOwiBJ7zu0g8/LjiYx
fwQ6pZMso+Vn1Lt3t9C/uSJ9xuEPyGEDmOgpIZVb3VR63hXOc+nMVkbjeqbbWrmQdDf7ABLQ5RW+
iPl7gyKWDVLmM8be5XT+zfyuuOkm/GcvDmXgIGrAWUTLL95ZO3GsUj2uRaehcqzpfjWbvwY8xmK1
jdVFT5xH9MMYNStqMPx5jJ3TR5gPSXGlovZbVgwIaWz+piBOY9DsaWqAJ7jGOeZ453XCb2DYJJnB
BIqXVxoeSF0q+4KgfnuKhnXo2rebeqXRFyYHVQHQp2fsHjXlBUoHmg30b81VIG9H2JHQkQeYz9d0
ZTKE2leiwR5EFKIQa3AyP8vPmwLm7eBM/sGsE9JZvHnRc0ihUGHZRisUpQYJN74IVFs2ZatIYtn7
yBGnEW1WpfNjG62PW6KmnQ21n8jP8KYNN5jRcqLs5Yy3KRg0cG2PGa6zxqoomWtRzbmfKyVWUHbX
Dc0UIrr4oaCweDKsv8K5+geMiSk2YyjerY7YSSFp43ms0uD6RP4gRFpm+iUQtjNRUI4fwBaLie1n
XZJEmu9PRNuQLE5G0r2Zk3zfLyvTrUyg/WZ2I5l+1YiNe0DcTCmmr9DegytoUEX1BVCFfrTdhwga
Qq498PjKLKQxU7eTGSHlTbO1xXhWJrPjdSFeZ1V4oBF/kfH+QgQzKz+rK2Cki1iLQuSPpukmthj8
fmevrh8DKy8HxSzX+1+5oM/4M1pndwV51S2RoGDvQ0g/hcQhbNR9CHE7jV7vk/osZ+yU+c3TASzy
merWUHdmGSx065alLUiLslkattwutwB//ee6Tk7gootguF+zTv8oFfzOgL/nuhwVKkGNgjCfuPOS
zVUMbzP1dHXl0dZ27HdERhTWH4ExE0WbE6w+cw5JJcN+kpjYQUxeRdbdT6lGBD4W6gJetmxcbtny
/swVb03eTBkL8wpe7N7B/tzvNj07t5INTKnG+JT7tB47B+pQzyvozZOlXlJy0BHhjKwJTpaHdS8R
ITfmt/1Z4zsisvdgmwqbIYq1qpXM4qcBWfdYukpWgbRk5gB27T+8pfVaygWUJUXH2TmP2nkiHWe9
DCPYTCVmkqKDPvKszCFdeX6ysGxn8lhLTdnRgekK/R+pk7WsRetMRvaOIKrk6B7sTsCZZtj5rGP6
FbNQm196dajzmUeNsjV3GOT2re5HFDbTI/MPLxNcS845FCHze1Ku5Lu5LdIxp5nNtng1NKRxTXQy
n5CSsTTWs8A4t1ma+n8kReXlNm8axtLwloUSUiKiMs078EUviZ7Y4MAiCQrjsxrFAyI+tt1oNkoQ
LDHYgoIRw4iHPSyJBdwROkJ1otn0Q7EkOcZ60FriFZC5fkBU6KukJ1fcbjoh5eOgOt76Hn6wQmVb
wYBxAugXVUyR+rbawAtdFagqLy/uEhEGS4IJZgE0HEOtjweCjaOQruy99rNt0w/idOTGNckmTYwv
GtsrN6ntRh6I+KRS6+TW/rVhTzYNuFd0yRekOtJJHlkLTRBzW8yhXKd3cxjVYjjT+DQ6HynYDJyZ
t3bIrOcdf7B8dN1UFEBdjgfBQFVUTtIlXsIscAJ//h7N2vqx5KglaaI0M1GMos12AYosJmNvq/pE
K4//W7RJK4X5AtTMkLltIke+et3U6Ad5/sJzHgFgj2NWD5X/M8KrjoYTBpYmWbwKmsY899jHJssP
wRqoh9blXwX1FHaFIfxjJ7Upjbmi9cTDeTNBY79RWmX3HqmVNtRD9Pz5vXcXx5ny9xwFM5CXkBpC
JdIKrb8sHYdjlHRGhf8QU9uWGJaJiAWTqUdmd+6n2/idFIEUtzvTAD8N2+eEv8DGIgyGhy1gnLIU
+h938ReKRQxkSiuDED5LZoWwXYc2S+oDVX9jls+QmVs9V63dyqZ/z0nZSgcernD95K+22bYt5pxp
BGIzZGgquITwYOZywVAiMwhjc7BzzK7EmyWfnhFH8cDW9Otg/j1gpS4D0WgJjBI6y++B4E090e9L
O2xfqKXVH2JhQwftFNobfbYUzww37pTkLNQPtBebe0x9kBo6+9vupWHbPATecdKcxPN8TVeHDpdK
UWa9pKbQOi7VBLBoaTxZplcGHcTMQutP3Mt3WkKOvSkT1UHFy8nyHyTSiOgrHEFaGEo/dFourftT
TAIW96qdeIPL1qZuRhUDXIyHxIB6UBR7Tzzw3iWGgIwZLaCBH5dMK6rgGfyE4l9fW2gUpXyNLmP4
YJrhRT9aFqfwIPDvNbebwnmGW2CA7xxtd9togG0Z7UzEcoUsj0Rl+88ee5x4G/krhN29P5v2xdcP
ARsDzFZ4shbuNKqOfeQ5B73ZQqym47Ch3l5jx64yuMMNhOoJcILS+vxPzLUT/xATTxgqm2S8WpE2
dRlNQK0Z34GPmsehBBfPNJC3QvZaVfJMWFo4a4W8XbyWoe+aiKhSywl1sBpq+01OrYxGtF8Sv0S9
ZQZgj2uuFAL78eZ4XsGfQ3WN73ntmSJd4bOka1MHis/9SM+W93ZxvC6gExBxJ0Ff07HOmZNAuNzg
OFCxptlbd3krFdjrWFf5ajkGkv+KZicjJKQeU7IGazLrk6ESl5aa7tCVMTAzoU2r5xlYZA+Bqbaz
GTcOx5YcSg/M1kefHyCPpZCZOPxHJiiceZFqYS6uhHcZPjmkFJMR6ofbGP9/ILhivHQ2ums62eQo
5eIlWxgrZDSpkMqyx4TfdT1ajHHj6JwVyGgC2tlDJJ9HQEqfnlM7qslPMA522+22BIaL/Ru/64og
zJgmvz3Xm0Ejw9yF7d2Mg9pJ4TWNqQiym1bXR88/nbzuNMTJ3lRoJGtYChb/qXSylEJWMy30id3+
oHP87JHx4PKmbxO2q9TxoQHe6ElCnnznCdHJHCPk5+0dc98tYFaL56m6roAGqR8j0dWyUEIbibGO
tuQTEmerbfSzpTMhUgNSKPkBt1/mYtTZosYWKbr0riIBn91hqVUjIA8tkawGrndI/0oa1ivSAkuc
JWZ3TOEFjm72+Hnz58sjbi/Kqh54iPbKDmH0YYGSj2sf/2VeYL/ackI2phEroX9jNJU5u/i9ooPa
81lBH19Ux/vlpJ5PK1bC2zplWVF38Gupy1k915Z0AoE5eTu/BB2fEisNGK/523D9dl0S2ytz1fA+
A09a4JfDfKXxuZbOkPRRJLe5E7wnlo1A01gHgVx9v4i9DP0MX5nJ93mFTBJxCjd4QXcD2k4U/jC7
HGQYWP+pwVsSrpT6O9t3fPmYjJFPc/nqPi6zvYgRC+GUxMmBAgI/J4YG7sjEoUjzE+wH47K+ShP2
MruJLfwv3wTAD/foggRsF7TXdFVFVbV1eauHDOrROhStYvICXujDwWxhIGk0Zjjbfq99bMfp2lWM
q7TN+L1MIWcoCp0HJ5vqroCmJcWiwS/UigZB8FEX2gtTKJwtKNQH++T+boxEl+FfrqWMztKxygVo
BKY0PHVkxMbu1lrUtcputY7FJerki1h1Miv7Pg2mXdyEYtkD66/gJ+r1NzQFyMP1nLwcB0ISUGTe
wTRNMHAwVth3GUVX/zupJdDczHbVdNBD2O1oEQPIt+cf1Utx58va9hfGVFN7RHQyUxgS6swKDb65
SbAU5Rt5/5MD23OyrGcrQOwVceD5JHd8y968uOgXzI6yfiCW6ljR50jZiEZ1/iiFXBW16Dn4chFW
Bywy9WJnK4pOjV1sxNJYFRb8PZAHN/Xl32fQLPk/qGXeY4E8QptDyVxAyKnBaGT51EDQviq0cOUw
zwWgiPOHQp6Mov6SnStljU0S4VBayRe9L1KakGnMBQkM4Ln7RHCYrsYR7Rx5MFXfF0s5q9NuzW/7
uJ20k9ueeyY0LmsVIvkDaJsWJY5R2VzosjDlHjQ3dq/6QZRVUFZEbvLSsnSAy0UOPV8fuCiO9Y4/
6y8x3RFHTuD/Pl88iXw+um4jfXe+hDWi64Rid976COkTF2NpX7uxIVCrdL6YFIAZmrjGVP+Pjhy4
nvt/SkB4cc4DheeyxP3gK6HIY4kVQuhxD5sVJ+VpjbVl3cDzCNEhvrC+Swi6S+mnOduViq9Q2TWg
ou2ADtRCeQGoHprzm2UrnYfdFjG7IM5pmykMhZpj01Alun7aXzZK6lQqTkAFyG5eRfMJZJwNamVm
bLPNse/DJQefx4oxwnlG8wY90cpXQyFpM6NpiViphTd2PTyzOJ8+6JK34BVOKuCK2ocp4X/l2AY3
1EVL1PCd2oDARHUZz/6i7QZKfQi+edyL4Z1eYsb2YD25sDwgTe7vI1HchlDYxZEJCcaHbNEEuwaP
QJF13Dguo0jzmh6QUtnDRzqjH1MvaU6nwx47NqO9LNG/P7w41f/XwsWvvC9ZIrkZlhME8vKG1QjP
og5NPxt9c0nVQGiIMFLpPDYMcTRILncyPPhw7xvP2hDBQDEbH692nvcaNAxomlq4+ZqfR0dxckas
AqoXfiBqMCvHNcFIzhCjh78vIMSaE2TS4sijEh3xsQ5gaxSN6T3FaegbVyZZuxunEDuvGDe0bf5w
qgHsv84a72pLY1HS12zMLtpK7ADy4K1uAd12DUpfJ13czchir+gfhy42AD9jRyGxxH8stslGkM6z
fhU7dFNhXoljKfps6z5bv9Yn+KBIOomX2bFXgH7w38NOApT0SnzmZnprWdGbYLnKx730MaSFdWGb
bfZFXLc8emvY8LWw0sKQI960SmZWKQ6z1uOS8yLo3fE99XmblNcO9BmoC5pzmvoLSUsVRCIcOtqU
HoxhMzIWJigZgpUNsf7QYXybQJc5atiTes4NflBrnS1WYkdRGdgqjTM5B/lVGyl6ZtPIeuibbasE
6FEUDA5rniVrbBqFhl2+LWIWPkjdC29duFpI8nAfjVW9IaIQw65CB/Dp8wfEKmutD2ywMvUZ0YIs
oF2tA/iA1NXDczlMJ8WlYxaLX6XpPuu/3JffKguoZBZzhvkEoYvjB+QdKZD6AWpKi9Jh8p2cshao
tL9/zm6vny6MDctDezfmGiVfLl1Ax+59wTYBfqECQny7vdpF9j5ckqlog3niORc6ml38yW0DxIz/
aoQpchwNk7PcCd4piMamyH6IxlQMfq0zFZGjKx9muWFqdJPT24DfTuHdUrXL/f+NXJKWurJxXH4m
O0Frrgwo5UAbj7BuymPix1v3pLsdaSV7wVjFM1KeyrEEHo5Kf3XrXQZN9sd7V6PvUAxZviiuDAMm
WnYblrcb6SAxvKxLIL9SCpOZvWmMZu+C9GhEoMl5njpYRTV+ScDXRdkkV9C7p2+pThJvdQnaRzZo
DKAYFPOzv3mH7wQDHskmicSpkvpSZ2BgXUb2ViHedg1zUeVFaOs4iPYodbqB4IAJ2n0sSNNHknBt
nr4EBRmjkc4QLe3DepiNIBmehuMO9i8J2EHFf8lfbDc1ahV58BnAx7zLQEeSOBxwX6APC6mdVTs1
nqqxKeVctiBXm+oTIestQT5zGyEBpk3c14KxzgMDodcqqGYh+PTGTp9/bDa5n8EkYM59iftPaBXb
ycThOd8/qvqq9XwVgW1sS+zrx5L4haRyGMxcbgAEYNkM01Spg/iGUHEWcCSDUJixLRzDuqY5pgRX
CY430FY4rNXLM3Ujjt4JhTgXGj/XWK7q7KwlD7Q0j5YA17nzW1I3QbE41b/ehw+Sk0mjtQtopGWJ
8hkuARICvEv2tJSJi8H7lQXaI1xsS1c2ri33xNInACdkUKSWsbGdLb2+U4TnQMWJqUrZHg4eBc7m
bfgmsqgI2EvAFvRm5zbMC/DqymR+jwDJQ9DXXFDbTWpHV+/rrHlU9w41EpRomXGGk0vgQaEMw/gN
3ezPYjth96SctLC4ddXCpiUJPaZtb6yczyI12WiV7wbkW1t7FvpjK9IJmr7AaDVbcD+nXvzGXYSd
BDDTIGqSBk5UHiDLKYKs9ckGD9kimy6vVmlTHqfjtjCqGrpM+tY5lA9jNzNn7ohLNafxlOraOepT
9Tj2HbUSlzlEwbNbMUoNvdTUEQZGqWoTk22U6TDwAOi/O55oB1QLqDfcVpF34m+FNawJFeiu8YxK
OFvCUYErxuQzE0zCKpt6gqQ/AtToC9LQ/kd8EDZVXd4YsgDa0F3WZF2saQMKhTdLdO4g5akgS8pq
5XiEL0d8ZhC211XI07NlwUWEx48XLY+cEq9olyDYyG/BM1XcKF0hN6rJAcpxUYkaFo1dO+B7pzNW
n0iOx6+HTr/t9PMEZviRHxO/4BYRw4t841lHjKYOXbD+obAPCuBIvWFMBsBtcBb69Rd+MSBI2oWe
oDqToZBDcLtvi0O8qb0plugvgfm0ds15Izx81rQKUy7TtZI5yT6ZQ3SrECG9W9u73509E5VyCGOi
8nu0ZW5f8v2/hGeObhtaITNeUheaGEwh43JvegvRoWegKZcPX8tkETeW7mvsc4u1vHwZndqB7Jn0
bIiSXZUV/CkfRPn+VUh8ofbqOzJTHg/rTFKvU4hoYDkBBA0th2IR1hXYzyl4d1LmaOcxnh+U8IeO
PLutU+nhesFG3HS2d9UgJFoZ28trRTNFjXMfgz1pkUi3z6ND60SXjOcsTgdn4bDwTeTh/CczqMcP
OLYjJvEeTkPwUEMz5wzg6Xk/O6ENN3/1LtXvfo/Q3tkDNQBeuCrnlE01ifDpTFuWuHaOhmnexahE
yIMTGieyzbH6lPkyTQKFQtaIoAJ9Jvk4lgJpFnC9afkKL5/Shk0DwAKEjLf9dt6DD9uoLUAM+cnh
8vArd4p+4BtQEYDOoqzqnuGfgYIBvhg3s3aKFN7njh6HbmmvhgY+LNowoiIe7+Ylu9KFKwryGU36
QG6TgNZoAa0zD9J6JfviDCFyCubQC4ErEe06kc9At6tYt8NZaFiENESx2bAVQLiNheVu2q2mTgWK
bmesnpjmxa//JXf2TZzCbJhioK+WmH+tcTZ1Td7ELXidgI+GyuMm5qxljLjcHg2XgLbhgq8tSulu
UY7N4VFNQeMeOGMAmhGvORuzELyEt0Iaa4td0aYGB5k+soFyblr8pOqG/SLaYzhI8ltHI+ujm2La
NcpBct4OOdKEy/mSG/rELlYeWSGn94fQHrjWaIl0h4etOad99/F75rCIpxrtsI98q/iLxfyZN+B0
uuADb3aeWGarmbw4JPRyanCWoiEjcQKGAl7pSIhJr9e0cs6kqSgC8oNYoBOWrfzx4DkQ0IqsUDny
sdjgm4p9w4lPrY4tsRO/Zwg72CNxI4JsC2MybZTiZjXKGngGNY3I2DrXBZH+b33cZthNSZkh0OZ+
XYBMRZJoPas7KK21cyg3/KtGFvU66Oai2mPizcHvRkzvpvuw5WMlPqGsnMZCAjuULliCRYqUXIjw
5d9IybJ2JAx8r+MF8KtBeVxcyZmdg7AkzTe72BeqbwFaVgZ78FRE3t0hgE0sS/dykemmwUTgJM3t
vxtYiu5nlzca/yUm+v4eQ0Vzc0jbGfUnyHHyIEYflysQzIi1gaIJym1I0jKpkSscWCQaqTWkMOGl
r8yYPuYsJlPvVpgvxDptXRIQts3opY11hsPp4o2ina2cgdjxhdfLoecxlxoDT2Rfw/CgfmqtN0F+
JIJmgVRAzwwOCeVrG4pNGKIFZ5KaNqGBqQeGY1wIMiGkoIiTtnln+YT0KKUk9UJgo3edX8TJ88cx
mPOAiJtSxBU3FUiZ0TuZ7Fm+vhLujptiqknjYCHAIan7XhCbvLo8qFcZCb4v1nkogTkq1TAZV5HL
+Dp5wR1lwMrW3x6nbPw/qvV4HON/SssmfqNtrR+uPvGBD8IJsDE+EerlmmX3kRWDRmzJzwScxkKO
0MRw0a8opH3cVvUkTl+Mzh3J0tr4BQg85fsaWJojg5Ga4zFbbjOfAEe5zN+Bub92sr65Zi2VK93r
dh4WBxp2KPHss0S9L2zfbKr/EnuJHYFkmVc6lTmMl3pdfoZbc4WKxs8+cjTmFVIQruGYrUtiyWjf
kbXqkHXPWiKw5KeQGRhKTMBIHTaleTxRCTiFkPLJ1QBiyZ3jRMEFyC0C4HLIeaatGr1gMF/u8zyX
ryEimmNdAl+x7drDA8PVzRQFTOatvfZq6m/lG1qmvvsDgzxAPlfVww2nlSug+aO3oHDNBLcBi6KD
HzviIgCjQttGxMNeL6Tl47vxV2Y7kPFFt4BUhzdPqPXgHsvbVC3vyvEQkh/+TGVvA5Bkr3POu5on
CxDHHBowYEbuRx5Y6VC6CkDAR8a+05JYwiOt6gh/VdCTRzXdBdEtSNsTaleo6ar6ZXut5ekxXJ0L
mUNshpVW9iLYn3kTe51Yp18F1fOYMrdUUy0h1ae6XO54sFJOjw7XDDSjENyKUFSG3K/HPC64UbJz
SX4gX0vt1qdBZ1l5XjizD3Vbg3P5oD0yifcqVhH2E2+mkzqlLruiljVllNQaIVf7+QdxTzzPthpW
c8PE+EpjOyI6b5UHXGahskfxNOiQYF91wV4zljLFLgXCl2GSIh62dpoUIq22TIAhP9mbj84UKbvS
815FFvD7VUHLT4f9C8Ms/wNHg23GIjk68qQo693L9osyf+KDAn7V8fRh7WgOX/Jjgmqv1QQx7h6q
h0nCDOcGbuMoTqSei20FzJ4tlbFzEZ9GPbqbsQkGDPkiTXikIT6wT9+qFMgMIjf4g2fecinfKIk/
j/63y2Tcz4u8ptpol3OT96aj5fuk72ZgDhlcg/6obbqUuik1oEZKP+dFvFc+t3eWjkIgD3bxyzU3
WSyt6mcf5mhlaC4VBp0hPjk92EAkU34FOy0UnvWtxeQ/AVyksTzWXP/YCn6lQxZ7QTPluG5zNIQ3
7HlFNIx7rqmkN+zGEnMoAztMvr569PdkkN0VHOXQtIVlzAMgpw7Sn+zJs4SejUPq5B20DLRU2/Cv
PzlOkrXU9Rqsy3gac2jUGOB3f8ki9GWBmPUCP5wplaAjHTNOayl3tHPZCK2YvHqKFbrZOr4fab9L
uvLS5eIYfVBhtKSsrO9HD4jTdHvO5CK4lIxbjUb0HGcZcj0ivR7ZTk495UatnPcio9a6Wk3XJomd
Ph9o52X2h6V7eiMt+A6MgvK1X1Aw5rCDNuqiNjv7rlpWOQzRzMT1LjuZGJavKgmMCXoG/4j06CXV
G9+xpHYUVumbiBqJveLq0qTGTtRgF/YHoglvLx+wssSLJqdHGvSwYwROgVfV3AZzCEAC9s1vrN7u
zI20FTS+CTVMerbDjmZDl9VX9C03LwllzTufG/S7NcFrhrLXKOSTpDo/6HpMrMWtg6Ii7rUDW+x2
YW9VTAJMIPAi3EIlS5l5sgvPaU4oDBJ4ZBmLvyEIFHbvEmBGHbDUOklD7nZwAO6aNl40CgEtHGMZ
FccNlTtNqCchFhsHn1ajVx9MaX8RexdZydlrlpSm3S9+Zk6dtcxzLDmRyCoJH4BcXDA9x17NMuBD
P7jkZg2UWwAMJC7rNDBBvIZ7yAc0vccZjLWdJW9qcjgyxUPuDcAih9LZAaoN4jURiI1Aoz12nQ/I
lp7NsA/qxLE7E9MjKIJXvrQjvE+le/BpyYgdAzo1o7XyTDcuVU66CYUXNTawcYQQrn+4x7mv0Xim
Kxl/0VlX3G7ZdRcCt/HL0V1UypGv37s/R1eQJNB/I2NuRtqTirK4j5sraV7cPO5Ksq3e40PTnp5A
1UHOoU2dvuAYLnXFG5ghUDG9G+dwMAE3c5UWz+Nj3IgyJye1HtT4iPpjJI35Ab2epgBEtauBCJov
6N8gapaH9mHeCoPHNYXPDOCJlKi7Bb88r4HKsgeFVrLP37qmJLIcq8thykZDw7eHgSsmnmpA3FEZ
qv68lzJnD1WOVcQzepaY0VFGoANw3klPnmxBDlBLbCkJMTSEiyXCK00NSQEL7hNgbINpxZQRgFdH
Z/tmoLoYkUegpySoB7C9xGXV3ml/z6Sep5ljmsZQR5HV26RGIL3P8svHBj3AjlPqCeaMjtippxLi
iZtW2OBGPDnZkJpbs0d22smoRtspkrbi21nSzT/if2IEX5CtNxb2wcXh8Bi4uggfEAcEXJGffek2
nvezD8EU3d6Mh3lnBPP/OFDg9qGyk4v43QpSdglYD33GTS45kf7LXs3aBH47QRrkptSGCvAL4upU
hd6vo5U8EZaK6FE7AoTxbqUtkSQEp+djXnKlG9Ugz/dFcjtXxcZp5R3S8PTGEJHEPNoRTBrKCQ0t
0Gq3iNZ/fBatQ3rDNTWst6XUZTGIB94BvHY7mSlAyKbPNr8muToWVOX/uE+eRIz/uWHes0Fyrsdq
3OoQ1JnZ/ZRN0XcEvJ1mMhKOsQ+DhJOHKuy8PCE1SE0AHxREq9wr12V41wPgByQ1RQS0p1KfdHwA
lP3f7/ATpmIgvVhGZAm7hcDvlv4oHhmGC6/m91Q++NSOZpr0nKQLOIxs77oo4hGfjDEbT7WCQQrQ
17XFEbxwKCckofe2fyh3RbarD1gcDel6I3Mv44J4B8RE1lgA8e3PIaKgFHp53WPgHj/r+IFH0Egm
YolsRmfdYPGXJNfGwEyY9wmpL5vpQC49ckB7OXm0qsIqjuS9szBSv1np0FiJ0cFbHnNRALIcMMBh
SgK5ee9HOairOQZ8M3LF+KbpU8B2qD4ozR2fEvvJIO0wA2JEkefReXVG+5YigRsmwIZqznjZN8Q/
vlx5ndivE1SVCfQZouNp1jlmTNPvqL3WrmYBkRBe1oyGojDSO6N+jgjQwnSshnVsXmgowEUI1WZ6
PRSexVW9u9xue3Ank8sM8N+RgX2LRsStIDfB0TVdcbVDKVVNjidVq92PMvYYifFsq7jqhNBCeBOo
oVMFrronW7s7i4+t13PWNW48VkCksZOKaII7XJLbVkfubzpPYgq1TO/hYzE4gdm6kFvZzY9vge4B
M7tq6x1u5MA9wmOL6OK0mcs/FpKlUjToMa6XOkqaYYac7MV+FdSMt/8kjUdCK38wxqsJX7zjf5lD
jW6boO4wr4oR80ukPHURxyK86CeMQemr825BgUmN9WoHyxXA+8UqzfWmkSj8wo0+5w2doxW3bfo8
CP33ata6iHIwGC7juzag308MTM3bGO0lI8HVAst/+/OGthLMowLvrNjUo5A+KejI43Uxngwlv9DY
fLYkvYMEbroCiQmhEJQzWcW317UuS34BCEBHs4SOWo49Ch3mVeKe9vfpcEDWh6hGpmqrKpAp8uhg
INswzmp+j/fUDLkZ927Tmxt9Cfsb6BuJFOwzJKZV7PAJHyKPmVbLskjPOn8caRc6QZyiYmaRKL2T
+4Kl3nYyGClyZ0eFj6PRahnneyW1iybUVjibNVRza2lpTFr3HzEN7ZADFSSCqHJCg4OKL8+L1biu
ggl8xuLhjnxd5R59oJ8SE9/iDzA658jWgEGMqtvlO559Mb3D44NSoEr57uYhJv2ls6Iho+J26hz1
pNp+BmI48Di3ZSyszmGXQFIzsrN84FYERnf8MbY7mPNG/u7CH2ps63bDKX0rExx9KFY6Ru3D5+Zo
ZnyOdtMbO2/SM6iw9iQjixzhZkV08Rxnpn3Vpy8kSzFSc3ai4kEyufVzLdHPLSEb1ZdpdFu6c8AZ
Rzt+wY4pfpZaC7pgGulNHM0gmpPzzF5zWuR4TnyFRNyN5MGW8CVjqEqdzdLQmUOTBIil0QVfOcGn
/T6TM8uHZrFVEazE11FPFweQCZJ5dfGAnr9SJzZHUXvRA/2ETdvEaH/Ec1wI+bKiw5LQ9LLAkpVu
gffyvOYMFhgUxvVuTUkFiUKH3GOO9rjztQFSxg0sv8wS3hQK1oyqngT7r0hxX2zq19NpFsw/TOJa
x7Z5C8ViidIOqZMkj/iB0GAS7PZFR4WkccjD+qDJ7M9w4cCpvNc8aifiTZHDascckrDv0XFgUCKY
jf24+KJaWbkjSFy/6uYDJwAjWfmbcUy7sieFz/mr7tsTf3RMfyGVC0MZFtHtus0rYeVF3IIqp8Gt
wKBh4/2TZfuH+bPJtQyuWVTAaGtTR+sT3EdgF38DmnpDnwlbQHHoHrdVpyJlxPN4SVS+OuDHAjLt
n4Sk5klu9AOOdkGknBwRx4IePoo5zbVCr1B+zA0PL1fqCNGkaYxW98yIFjmn4k8yoWeurpVlSmFP
lJZ/Z3YYXzNYcsBWu4RpCZKsFJaA+WUSMEeZYeNdzmIdtIpHGRDXVp2shZNAo+PzjJF2SMH/vvv3
3NLqJHgLnHe2FoSJgSQHFTmR6SiG7J6D6nCCY5NiGkhjUiaSuOpbDl6Xt1PC2+mm6CNXShz2bQIp
sivsyqXC4fdIKxjGnwNXYKmVAZIXXQavl3UsqkNEMj1zJ/flxcY5tkbSIR///SglRijY3KO2Hyq/
QmIPq+duSNml6u1VxGXDw8md7w2/T+ntXSpqsj6v9By7DM+EnNddSwGAE5uRlhB1K28wXWrHssLU
KeNEy1EI21lXZE6gO6f6EhFtXxqSdLQjrsqg1VLrzGl/OxC+9ELhuOb49Ak0+sbYyMHhzPQdUM8W
2nh0Q42o64VN5vntPVIy081WwPuz6/tS2zXQWHUGDbxQ2mlLJw+x4/6nT2V3WwjNxo6EPN4e4G7c
aJyo5kFkDfmiCj673d1RoDbTevHEvhe1rwWvxnYSvYJpqg7EB9BPnDFIvVtqlLMdZxCu0bo2KI51
PfmnMyKgIqq63H/H1XefCrhw6FEWkAzz1TKJ1sj92ZkN2FmoySJDzbuac63wBSTFniXNgpUw+aHe
RxqgKsrVhkWByzQdFJHSpeshtt3WfVTs/xgwBg1zLo7x7LxMneQFQuXeHCojYHoH4JSpoW/ygffx
Khx5TgMdLanInQBxZT2ZBYw3yO03NQ5vS7kj9aoF7wtEofSveSTEVeok/eqhpAbbPwIG9U8l3SJr
Mj7EowzFgDQSF1n+7G9OKBF5dd2SR+j1DDJ/nacQ7jQceuLtlypcO6S0IrB41N54SlbB1n/L348L
KZa3fekYYXO+sLrcpmSh3vpD2yYgo3XsxOVCC45kiu11Q/9BrLFDEGOMnu7bQQIfJxfol3n6dyMY
5CcqS2Tc2K6kzQs4558r0c/AJP99BK0qfwilby+cjLB4Yx/fi4L9JGtbeXATZ0l3xGN60cxeWTuZ
qAZ1lCRQoWBv4ulhHrwkW7uQ8ZC+yDk6BuYKaahkFoAacYqdqTva7jeWaAp6goIqEIogpIkvsCqK
CUWZ/aUhyE8RD7lrCyEs0Wkg6W4Ttrs+Y7St6Qc7oxNs8Hiom6ni9ggJIhAVw+Q1IG17Uo0J0rYx
DDC9/NT+dakIyzThrqJBpKb9//SKOT0aV6Jt3sMwtf/+sFnJXUOdPQYUHc+fFWgmhZuf+xQfhMcY
qJHDRSrE7BW55ikGpv2K2/W9a1bv13zZ5yccYNWZyebAykBxuV2928ecp1Sq/ngyWenPG4pLriDE
8e+0tT1sySw5voQkHixsOL+F+LfK0XZ8hQ7+hiI4NYMtOf46Vz8rRWSzfF+gzfrPNo6hLcObQ06w
G28FB5JEoXGIa2HTxqQC2+pNVIHRiiSqK6SAKOex59iMckjz5zd/i+9urUYRPtSZ0uDoEW1JH8qf
Rco3/Yz67w1dXuaa5OY0iriYfjj2SrAP0n+e7QhPlyymgsWF/XyyMz2H2HK5K89orDXYH+HSrLJ9
y/YKi+Gz45YjhRLAL9m39WM10o+7hMGoCj87QkpnfeSPQoMUrwNs4An+jCx0344rZgOxbR2LFQMW
UklilFHRWrl9PJGOqmzfGNu0XyQxiRvMO6SOeGmTzrgXTot8Jg4PEgRbGysuO84E/1eMVpmx0SYd
OTr098Koxc7twV9igdYNOJnBljMHPWa4/lfVaUxZLnPwMzKLmsYTJ+1EQ1p8h/P6OL20SaGmjH27
g/1QqQhzjePkGFFDTgT/Zd83otYVZMCUM6RxcDdWAFOFHyE7bw0WIdCSHYPmPiXihMnsQL1GK+/5
iKJuW8AAxplwnyfIVd/l3v65B8Yjm+jV4ey6s/o9VsZEiyW2eQ0mpCXhZcRnkjxpMMB701CnAkZD
IQ2EKwWl8p8WYFw3+DQ2B4vWkkNKXdqNj+dxI/LzeRSwCHJCJ+g+JKtJuto7fAgde7+TN11Saqmm
hnX9UlCTxoYGNzTwfoAtZ9Y5q7hASNQK5c0x0RWkYR9YNLTEBoHiEK8p/XX0zQPAY2e0AVdao0RT
FUaBvwJYxe77fklecX4xZGvP/jWaS10oozOdNJWsty/P7B5sailEss+2Yzr7iRgJ6mu1htdJTsAI
RQ/Kh0JG89LpiQJu+GOI3nnxHpDoQ9mMEXrU9aGHD5l8vbegUIsZdEPsd4yt2owFvC/ommVbs35w
fVFdLAcrbuBZ9BJcu0DJ9rd55xNkozWlHw/hoWh1gWUgdk8F366isxbwsBSVe9VlRi8pF53hdzSw
5zyZTclifsfW8I4X8QpxK3PXUmRNW3erxXe6WkELQ1pvdAYiH7wQfRgRgmWTPvvvWsGGEsgNQpiL
WtivI8UM+LX4KxoXuW1HzJJ8RtDmkX/cJTzH/SK/6qDDyYm5lb/rEuhJajXcPZydWrXAO6yfZQFL
iOiaGy6Bp7RsXY6f54zfcRo6gn+B5mguBPwI2EfV8bKEcrFfaBsjqGz8jVHpLfkRgjX/2Ofjlwwg
2NCO5Vflk64JbDJYTQILmPHoMJBQBtZs8JvIkfPhyCnkMbPV8xT9trn7WjWO8op/6LJx7+Q9zobV
r3OZNjIPN9QehNbT9ClTEH+80izilFEZtDcvXhvJ8/ppFL2EQ8GLS4NP2i2oMXaVTVRg+I+9Dau+
rZQdkA3jjs9sknWJEtV73EawY4/+BGfUuigk2j+GmOX1P+4wgfLKuck5S+QVLRSMJH5lviPtWHDo
LKAUIQTth/kfIxnSwq/aIb+T+FEQ4rhNIzZLfWC5aT91a9vjNaFsab8fEOONM399M8J5V6PZyHZT
sbNFGgKbJ8enZLD0tZoPcu0PU0JXKx6z3v0TNsCvBzyf7hYqx5gENFe752IuuW+/by2wNmqEN4wg
19QEjuB3l83l9rT7TMF/KDefsCoPLm+YOuk5I2ReeuXICmJFATSoWCZf+YAUF2Owq75xhMLVAxjQ
QyDU/Sk8D79g6mEZkCKd5owSewJaM6I3NHy9Rj4tLMAaNk32oyCzIM6rxcRRQc/mCXEq4y2hQ9GE
1Q7247pwVlHAvKeOLix+csW/olJZ8znRjRshUmPggqXnFf/Qr2BrXlL9F0XPO0oo06e63bph06BU
w95zSC28ltwMnS5fgYBDnfHftzp+wzCB3nhF1ZqWxRePOXQFehe32l/4DlrFxCdJVEJdGgoS3TK1
BLccIuivZpAhKq+l7kBpAqk/sgw2JhxfI1tvsJ4yYUNtiP0x0zONWcsWY1ce+hCLKeLiGWaNRhgy
9pyL6w7pykMMzwhXeNfhrIvM1e1t3X58VB1Y8WYrNc5CAPCbUKWlalb47fnGMHeSSXNJ5XCON+th
YGIibM7IsVoVsvI+I5ZFyLdVQ0sb5y/HkUXrmG/I8+zqabPWncJ6YUezSI+TwizBxGqB2noOoy2s
EFqFFdJM0hirjVraOQn5QRZYtlkQAYDwUJVLzES+FY04+10jLR5nUUHPVZ4fO2jcw5UdFRDye058
yOg+H4n3pwCZS9cxTM6w7t8W0cSiVAbWqVoCkJxvLnQ+zjalXPf4026igifR7spBLC9dhRzWcOg7
z+pGv8XjKTbfn6dsa+ByoXj569erKPxIkUtxA9SFxKbQqMRFQhxKe0lIId5Ex4HnA+00XcnXy4L7
sT70C+sd7OlJp+n0lFcBYq1Kv68Qdn8xtwhCTOmL3I0B2ZurHQWGn+1lnANj7fO5zFuQDngqqj3z
URLnbT3LYRPL15LNTNkp+xFnF1ZVNSXIfkRpENbmi/6UEgTGX7oRVB6eYkMULkJYV5451Pnd0D46
ji9NcslLhVSLfvoj9M+o3a/KCXhLjzY4wN7nJlFW7lUI94jz9cKyCdGjGbcf0yhD8CDkULtJvsFG
JwxBM4em/lncQ+dQsdmsum3p8fN6FMgAJBfMlS+ZQ/JB2KEMrxMQ2q8OehRISVCbc552QgzRLMRQ
F1QEmqLr8Hwehp3ksWPQv3K0WoWxFYQ94kUActDx2uDFU4kEC/YKf18dDZOyAiGGdIm76vblpfPz
rpQF/QxyfDVjUyzMP6HQzPFit8OVfcFgdUN7cigZWpd+us8b/A6JUjeFcTXlH9eTeuCEwlrsewF2
5jcCZxGiK6z9tfOborNVPbNKEQ4vyN92WkwDGIgVBzd6+/x+yNJoMsxXc2BPS4za1k2sI18pjkzw
SvrTeNYNN8Ky2jUjgIu1ZAHZbGNOCevlwPK6mpESLiYa67xrXiF1lZ10yhc4zv4KRkYKqGaLNa9P
3lB/6g+xCVNvHYUfrzjCK/zWowbxWuzGOftVaQC+KCnRL+DzqGpWxIywAfQol6ZqIRt+gnQ9fw6T
VwLq4jwll+oAtpiHol//udcMEvjtIMI/Hy8oag2iM2cLjgu+fOHNzqocR/3yBMsLXpTwYzZusAIp
zFhrqSW4FZ4vhjMWLA63+zpYCwvPNnxpkrFjL1Tmq4BQQyCCk5gzgcpnoaH2C2ddYH/gp6vUB97R
zZxBpZzw5CEjyep68vHJ+XxDDSxydw+ugHUNk8NeKqLvVSvLaQVJozGdgCWBWA11+ijYldRYUC3k
xuPWkQe3nt89wEKql0/rJZHf5Ey2xXG/lhXQSV0+aVRNC/JcHxBnGf4X3aEd/DtUNoNeqkrAFWLt
oTwBHcq/wqduI5Pzap//ld87Co+oQV7TE/BMODGmxeC7DtWDG2AKN9Z5PNURQUzeogVqCLPIdFBo
H8d6BaGpRd06tGfHec+aVXe9/SPGyW93uY5KsPoW+5HwftgPOv04e9ptXeYiECbC0QRHL1z8T9tE
WlBuFHGD6YUZr1x99p8Qybm0/sRQl9vJkRkzI7f2Nvg6JaUL3TSEfEX76ij1UD+/rJ1xwCXG+vNa
LDMXQ4LtX3qgNlctZAYMQqBlmuFQrWX3jYfgCm0YsuOzekOLMydLQ8h81ZtelgxGehn1nIgXYJmg
coKXloOHw5nbIxmX7r4uMFLpQLiHcHyIXqkzX+u20E4+z/noHkGN2OzDQVw6Bp24Mw9XlzggEygr
T0ed7hJvXsNIEITed8to0aA3lZ10scA6mjInfm2ElRGB6186ZeTTnAm//FN1E3BeVpe+cIdKbsWC
hoG9iPNWD7+ydjSPOV6NvuJV6aBN1/Rhv3RHFCtaYUYPSGcDkMD8WL4bUlgw1iQOojw7cIS53V7x
F49CeqJvCTLE8PFbXMai54HuJjqO3hbQz9URyDVS+3zAmbKjVs1E8s2HrMnxZSmm2RpAqlFhDpxx
DDLSJM0eL6hCbqDqL9pyneYNztau1DJ3khvlguFj5ofX+0gewC5WQ1tZiAa0YzmJcZ+nr9P54tex
KhSkHEAPHT37RwzkCDsBeSLy6pRNww8xZlN/LRcRCTBNneCXXQftfX/nRZW8hSmCmOH9u/Al8745
ziDxuDBkTvpYXA5yx5LqA5LrFA11GbORARd/ZnESsr7cvk00HnUku4oHeYvagf8pKoktruop4fVx
aHOOvuePvrfCEjV+zmjFDgHMR8FpftiSzRBxxwdwdhxJZyJueLOyRvZZwOSdO0EfrQugRCv4LNR0
dV2+G3Cwx49Vtb5DFyo/a/LuXz4JB6ixpsuk2D4x9vg6C+Lade+jAxdsAPCW+4Hx74YLs7d0BLCv
ABIxjrsOiiVPtQgT/aLJbcqCuMMF/Z3i32DDNSfbvTG60VR8nt3RGzUQ3cvSk2v+Qk7K2iZyj20l
HgL7qDGcqvJw+MViauLvU96PoIlrwn9Q5b9+AyKPUiexN4czS4EE0IkhdNJUYOJKoM9coLoWfCtD
IO8jzz8s6MHKnYJcx9BGaGR70Mw0AKG2XJqqU3ioH3DVVWFXTJ+S066EbWXKl82BoTvcamDmW0Kg
UNvagVruZxfAHGRR84kXnKzDOxWWV6BQV1eDWn8P0st7zdKTtToizXo/ayYgiDTc414FfZfB9Wlw
zAo8s1kmWQlBeaRRy1gMfoQ12MHru46d0jIbicdhLDvSmZybEj+SeN4W+qU8myZR9QFKID+0TNv5
88DAZ9J7uM1ehspC/GvzdAmd6+3hf1QwXLe+PH0L/JyA31UJtEKdLRajwz+E9ZqxkxhWFZHJ0MFP
ffF5CBu79olyMILidZ3/FJ05+HipX8Z7OiuOEmpJE/xBphYjjoXoARigkzEMpPtsPHiDD/dKYTnF
rR/bw2JmYfi/TUwNXr1Ox391kicp9d76O62LnOi8u57a02qwAFdP6uFeK3KaCwg8CHWxJwNkMKY3
z7nW/qBgch5iHmX3jCGcBVCQKYBiYY77VjB36Jf1mU4hpNEpn0FbNGXL6cy2qEOyxKyzhy6ursZS
xRLMcEseUBOj5lGDr/kwET6fN8oYc0TT9ctPlCFwfh8gr20md2+i23uLZTeL4qOWYb52hC6tLrUu
PDi+nvtj9q+nWVkpRkCuzFTu+bl2yCoIdsi0HtwfiFxRZJ+TJNVAMvhI61BG5XY/sB2pgHu3+RMN
KG1F2T/tPjeYm3LFDF3/mPsXxJiP7ThahDR8+Dj53n8X7jkHpo0HITwn8j9s4oTtfnQB8kX4V2M9
m4LC4pUWgJSV9D2Tq/7TmzO8uiTzfyJeCavjXvlyVBPkt5t+3AVzVWa2XJXCXMJZZCliOmppspJD
b+nrqe2XinbsNT1p8Dxye9n8LBJGMNbMxROGSaYxkuwnNRfy8grGhsxCtF09C80/fbaGBkGLLl8l
cZefCd2m3CSLvIW3U4Twi+BDKgIJIv3pTCVWKediUo1bjD+k1tMqfNHw038j1s9tzNqn2Lk3klZJ
grJtiGgDDEkCLC1F52rgZ4nW9qB1IHDlYRP645xqLKhaTx72XZdR0UnWucvsS7X/rbtlVmtQdLID
l/lkZBb2aU8iUCl3pBlzo8KghYVFFDWLrC1Qy+4H/YG7KF9jDj1H+hqgqQ+v+ehlCrSNx4gs9SSa
FdU9+TY//CLnzSlwr0u05vqXMwYmyCkzWMHRuXgkBPj6TtTp85QGnGa2KoSHNzMT/bfPyxY5Eabz
XH0tZajbVfKyfxh4w2V3M42xvWSsgPVoDM2p9tTUXocJ0XkHhur2uNefWiKY0wL2JdFSVWEkErPH
Ju5nBEHz8b/I9Su7r0vNqinmuqXaaYCML1Qa1+L0R6jolG5FNDskaxop9vQwVDa3P3mztZ6de1bH
lWRnBGIbByquSDTqa+EHCdh1SL4PZ0Y/pAWJTkRg1KoK+HyHwYDoZsxzewAYmtCz3qciqVxE4fAB
PmZlC7NUVRNVEQysUTOHMWZ72olmr5/cwL6HAkmxAilbN+wmERyl61fe26oRt3ZPbyqQwFADRaev
Udt9WGaxjjIdeNlvtFE/Vy+T63wxN+fgx69EpHQh+uT38mUS3oCGEkKWcGlKeoerXnha59+rsbjt
XMcVqtLBrbdffXpTAhUZdeVfhr5sksz7mRIna7HVCDdqgQHzmP3VEXSoG9D8laxER+J8ZBaPue3O
sL84GqdGSIfF19XY6u0j3HJ106MCHPumleKBnbItcYf9UjZmtQaVSC7YJEFKjIIl8YaMfH+MzVA3
KleXHPqkcGxt1iAUwT+Pte/oQl5LTPTvfMIH5scTqbGy9Tf4vUelc7LVDsTIPk2ba4nGrggYJagm
JlHhXavX/Djc14CD0AxPaCRwFB1b8DjAJJhoeyerYMTAE9VecfaWNupLF7e6ROUT4RYg9Z6uwA3V
c7gwbGbnlGcXESpEE4UjxLiojDJ3Vo1RrzVJMFvBFkIcskm5OE5N9AtqwRxQaIyOcdYH6zaifggZ
1GC7ojq/zjibZGjZ+/PvQH5Bw6SGE2rWglag63/suMLHW2HEAusCLuOaU/IWggRd8SGrnI4P5AhA
YfoDJND/uF2pJLsXBuUR1Oxn3C8TXQG6R63XKJObbffW5N2MfW18NQdDjALPFSWiWHowlsVilWwl
ut6gnawMv+isDgzuzPWS+TeRXPa/g6eGMaHlWM+YQbBgW4m2uTjnMwvSLmQ/WDdLGEy7U3NNfPP+
/+6MPG2P5GucxsbC64UfKwaAsTJGm/udpp262ZCoZMY+eRlKBictPzDNED+1F3O8rZaf9urhrg//
FcVQGd2PsxJ/xfW+HZC9s8RF45ftHAK13WslqK/dG2uSHCIT01Ju4hbMRGUB9Rsdg58Wn5Bv19l/
+IDfg8BArF++bjpYoo5XO68n0JcAf8+QRaDEdvgdtSFvqC91QMgaoz8pPZjDVHnEqVxAIJ+A0zjj
pXVX9iyIM/oOmAxUiCutRPu9OFuevjm2mCl6p5h/yhl5GV9j4eLumay4aD9UPwRJwfp1DkSwJ+Df
2SkyX/LGDCKq3kikZg+BYqvY9CG22xe26AkxfqrNW+utLXdZdKA+kewvNJuqU5wW5YYvSxSCyAkA
IgtyrMk7Tr9dL92uev/O4lbLB7mSMbokojCRkOpMi2ZFZxCq7Uus1Psu9ROrk1HwNcp3LL0/IEwV
zicyhqZRK0EDeqWZcaAL6E4IC821DhhPxHSE0AfXq/l9bdSizMxgdqxIzBrmtkrDxhPGkHxl2cUT
oeXcV8gbRC2mIVyNW5vduFCtKOoB7NLlqwmOQVwUHsvvpSulxi6azY8iuhSyUmVlVQdemU3/4LUC
yBNTszE0MvlMorTnD+3h/r1Qo9sjED2jGtaolvV+crIGBB6uKJ8rr4ToNSGWr+NNlEQjqSZmjrsy
EopIg9gTqoCmSDbOwZfwFFiRszcxtWKdQdofJiTqgKp3mjpLmxnVw1IwpSpHjsa8ebigeVaLXA9D
p1moPtN8posEqOtJEDdY55PBIHo5ccuPHo3r8tQ9pDDJBNpXWHvpnmpposUGd2y8/LZIQsc2h8sw
psJD6yzGj7Mf0KazCH7u+cCrCAmfrAADdnRnl2O1z50itXFY9bOSZrzJh75YWTnv5AP6scJZmB6S
1dcl17JEZDgIRFw4oM2a3dimPZsOfcqVD15DVQWYCxrNyT9cB30WqCU4qqf1pOcLHfI5kHUhdSlJ
4p8B2vYUKBL4b+PXcCBYriX7G71j1w3EvdBWgDe6aoKjo7zAJ1S4Ow0gGpWbTU4K7BOZMLj5qgAL
8hTmR4LbGv8sk7QdQ5EYM+FHHwth/hp/KJCJ63fQv7/2jtQb8c0GsudEFc/IexU6fjWluGpCDxUc
rQe5BXJK2U23bxC5vdcC9P7PG4axd6YsLyGTUT5Dss+qaVhqgTKmTGE0HJ+NmEb+ZwLzdr6qv01D
/9RY+Ue9oGllocG1IyffdthnoSvN2aE4Y6Hy+Gk5j++6xRMTs/SUK3BkIXwqibI39gjuJBqfvYft
VTDMqPGJvi1h3rBfxf9wOfQ8JZfTQp6b2ZyxbfCmzVzOfDdrLUIK4lrquScn/DWIgQG1NPnzSoCr
Up3KCSuqRPZTR5ydFWPxqxza2/kgnt05tw9DHR4ehDwOU5wUf3YYU5xXtSPAKfNhvXEFXb1IXT5r
sYgEyh/7k3F38pJ2aKlDQaZCqGF8GJQjVjcC5BYLrty0VSaxDU5eCFRj6Sy5HJIMMFczKqGEQxYf
dkB30Ed3w62TGoxH2VWuz33g+bnD9FFaLwno84pxq/v/zAberfeW5iCGoyKTzOqsyX42AkigAor/
MnDkeUoykrgo1n31+qgrM5+oIqqq1FqZCZyQ/zqwx5qF9xWU881i0iaAsD6lCWF3tic1PBZn34MS
L+8/zmcl10sJO5VR2KK0zYniJnPVONDip5dC8C4QclrAOrjvZNy+GU4rIKCQngHkJVRancoodhqn
FNeNZyOUnUub03QklY20/gLY5rV9pT1vbCCG0E3ZRENcb6qrgcSz5sb5WPo6rIlzyWlEoxw+aec5
JOzyk8bahJKo1ubc8I/WFzRAilmS2vxMiw/VwXpX1CVYrWPMBbVS/jyL4YceBnEqOHuaLn/M6Hrv
KDfkm6ZIHEu8ULFUQc01vuNVPCRrGZ5c9vGsk5A5AcjIKLOV+djQYMKpM94/nX0S4oxbB5J83WMO
sN9+lyb+eVE6tfn77w0rsiHZCz6EQu4kqD5nAnyfrWeMoekYKAx5CXwgQaiznKO3gvkH/+J+VVS5
hHz/A3O8WrduzBmaawU6SCBGxDmNfkVkhDviXJzgWI46cJ15Dya50BCgQs8a66GaY1IJwcLUoT3c
gGefd1NInuyHjkjhaEDwYdzSjd9ugZrlyOTbxro5x2IhHK1Ew5NySx8AAvuK4t/NF0AmzJZeEV7y
2EJeIdTjIlXd8XRVRfgoXgBpuHq03IBn4PTdnCpUZXejunruP2sE1ozf7fBsBZOjI5cH+FZMaxsK
KjMYiqWuVwb2UFRPn+ubAojjl4Im0vQw8RTaGhShhjY2HxikJoqD+CtI8rJA3QjarwS8iO+k7jJV
9KVD+Qayo4rqIgkoACY1LsPuKF2FX8qIB3FOVdG3dChRoT/IqKBLKtGUqTu0tCf91M4fN0sDlKP/
Mz1LUvDKnnqgm+4McNj2Inco2HJ2qEyqovqdeNzbVM8b+0BEnL/elsfUVtbucpieyZ7AWLcYpGGf
Rc8TZ4vTqwgnLR8P3VbbQQPpqVZwl/ul6lrAVwX8+ud31hDYYLJs7mYWIHEt1xYL4j+3EBPTc9tx
sQMu336oBqH7Z0ZfbeZK6Pmlnvw945jX8iYsucZzifwJnOnLyh2o1YOG2eg+HS70dcXNXT90I5iE
+3IN7ewYwcphyxkYx5obGwPb5AS33DIJ17hq+jEi7lLPHuEMmM7ed/5krWDF2dWewWvBGR/5MG0M
b+vg+sPHKdGsoi4YqBQyysNIzdqBmFyAyn5uWyWgGSK3aScyqu8pklTg1RlFIy1eb82cGAgtXMFm
x+AvRZ9PI0b2E5beRw3XnVZ4gk/RFVXOTkseZSQQLBZUMZ2Hd4rqu7pt2Mi7Dpe7yEx25AZdzAdc
TYyyQqPRb41066eQ7nUHMeBxsLDpy9/04Qgb5BXoSODLf4ejKJoU6fGiwWQT3yTwV7i9Qb/Fq/dS
9zoWQDzRZWESK4wL70a90SJZ+8UJsOarg8ewkle9rsw7Gj9Ie/S1tuaus1qinq1SHWwfRb1h7l2T
mWoxCKB3zr53km61QNa96IjMu8tCoD4qwdeLWk0W11CTN011Dtwyh+tnydS0HhXOtNAHeYtkjR81
tBkJ1GOYr6xqYeW3mqcy7p009czkChPwsAyhIy4lOntQXEJKWd+RJvc7ikPeD0Xntj3UHYYKnD6w
mUqkcMbq7BjJENu+J4Xf1NvQuX2YTzxlfey1yLBw8U6IBYOeg9r3EhRUT+SkpXOlWFLrsg5I+5Zx
aV7nRnsQqLcDz23Vx/h8ijA1o6eH0zX6IYDGmYjbI4kuN3OCpjDd6+642o+pKP13L43ongAS74lQ
EBeivkcQwSG3vaKiyfKOKpvaOrXM7cr532EZGiaO7qh1aAQGYcV529ul48xuQE//ewkbcQufSCr4
VWeqVFWtpjlW61nsUlnz/XtMcPJMEy+RuM4njwRlS/VpgXGr5mC+gytb3zWYWxU5MX/COzeG7bvt
C9hsnhJEIpSEEXmm/Kb2AriQ0AQRS9+b+9zEChUyG4JDthdL+rUc+FMO/TIHNufKUZHQge71owB/
pnv3Id3QgTUoKTB8tGcQlsgb2d4QZqKSVmu8zrYwwiftIqq0eo7uEujPoqL4CEk3gMY10rwKdWqx
Ix/oiQf9QGMRlkJRGFgBPtm9GrtcC4L/821Bs5+GAgK3yr4TJ8TKXYL8R9wOydJ6RVd88z8o4v0e
6+W4uj4gfkeUnOr5TYHy8fGzK7zJbzOt3HOiToEARhND5a8EWT/j/OTAowoawLRbpEkUvvZ8+Ofi
EaJcJ7paazyyHNsPG1jL0yQz1P/agOMG6TMHqNepu+bCIcC3TWYFY6zp/eR7ngcbXkWB9slIcS0b
74e0EY9RhYYsNo75C1mokougxZ5SVXTAbqvfG7tvUrRbTQhNsEk3oP4q/EIr5X9s+hBd4jKPHlAh
Q+Vcc5MFSGmbs4j6KjcicGSNRbyvBmdrgM8uii2hYrj9BFb6+eygP2JMPxF+INdXtUvFJWkm+g3D
GPPq+fj7KPNISstONwFrswSve6QNJ8EOdqPJBbtcK9zwqDZXNl8Erg5SiKwl90XtzUytv4VOrOl9
xytX4ZvhVQXhzcuvnw0xXMtSebZT8qRMzpWuTyc4XDi3ApGTB79XWZ66yCD9ScmTYoZxqLyenLE+
6z/T7UydNPAt4YkLBLeNsZzWrbV4I/BjSOM1WObteIEHk/+anH0agOZg16UF7W4+8GsFNTD8l7CZ
daB57w+cTChzcO3ZlQT9P2wPcEpaE7GP9hbvh4PsDWhu8Bjtvgri3TI8yE5Nn/ZVMaIi5Q/mFVsl
YvoAecbHLMe9xw+9rOF74+rTQD82IWtPv19ffEOuqPcvwhT0aqNidLe/xZZnum5DQqlTU6E3uQrT
yJSik2vOZvCYbC16D4KIc5jPWnqjGNeazLeVd3/pcS/ejiZ+a6OUPrGDo0dQvMz2h8WYOcaYQrEK
Ge3Wdl1feQKvpFWxayZyK/pmSlwNpjozqraam/AXZUjb3gIkOm5Kxh/TItWXiudO3yZ1CoJtBX/z
kISCxDPC/5nmKJvi0JysB/fGyu8rL37ruaP5OKePqcI93VY1H482IsTuZrQs3EJXJUcyTuTwd/2c
bDBmsNE1fO+GSwWw4zbIpZzgUrH/EQa2iTlVaw9XmoseX7ixV3VDSqOWkLHAMIHHTWBw7F+M838s
bQXdw3O9r8ekPkIZqQ80HHifb8ufQLezLaaKxXKFmUMQG7+qgYgVTk5jL4cRt/QdJWpWUIVEEkR7
E+eBtha6LCxIZr74h7fBwN+N+4toQMHmm3XWa+/3hdEUblfY7k5K988Y6Mm8YFJHQ287Sj0eiHJo
Jw2OMzTAWOM04UGreZ/kWvuEkCLNhC5mtUBkuQciBhQ4Dsk/bQxHVdKnKP92jrd8mqsMO1kH1oKd
n02XdSXIRK+KxdNurgUdcWAk9DGyfxmlrve1E1hAdiFneo2svgJZ3uIwI2xufiNz5RcKbCeLqc1c
xQnlYBzrZ4p0D6/EG9uyuJm1fGXI/wD99G4F4DcWxF8nwSyC+Xydw/tq3mbFp5/CFDONO9CRF9L0
kP3G7W6XCZRF53exU4GgeLzCFLLUYOAhRQuxmyuUdKV3iptYDfMpoQ1MFa5iZG487PgwCGsYjW6Q
AHlq9p3lqrbHvPurodj+cSaji8MZWkkoeqXBKH0qgrxuGA9ddqkyt1Qf3joAZZblfkvNnpnDnzZ3
q/4OreoGUOCFGnliuqFcG+GqRMMYgnnMOCx5lGo0YTFbVBhel+L37nbltngB2Q7CeULNfqrjhyfc
D1aEhO/2hC5Xgw0MBGcX3e/vs6ji+TKUzMNkXcKaYpXK6EmrsUUqA8YbgA0Pn1du8ZCXs3N7up46
yL63onxUqlY4kJEapRbQ6KNJ11/GmoLopP/LzO7B6+kuBIjSDDbqp6kIxzIyYv9KYDbNm2J7m9Ev
/hBGhZ38ITNpM2whC7+pEWABAcP+vABXLf7Zf7asATtzDvihjZ2P8IDpAsKl/yMCJrvdu14ZjcEj
zA+Ay2DKfVZ6pO5HFl4f2o5BJObIDhd7+fIovajES1fbYqAVhU0T2W/SinecQsxZBQbnW/KoOmg+
Vi1eMCwH1ONKLWQKRIabSeZYJFchGMQkSiOSyxP2p845jWEptIVf/m7m9tDbOVmklAad4mamEUZt
MIDmYz53QI+id8FsyvC5RCTwCdNs0w2ylmimH2MdE9IZK55BtRMs1KZz6nuAZjwec2ily41qGEDw
/4Sd+5Fn82aPnYbWXj65rX+AXOYEDaAR/M7M996V1AGbJnsyepDnYeak+ls4HbOiD+PSlgtLqwZm
3TKgn1VDywoFBUtYxPLlxYZado/pVwuQ/8RHN4RvIhFAKO+9ooQxxCwMFioaHSvOqoweS5LU3t5R
AlrNOmPmlNcMx4jkOnGxNwmZOH4ujZcjzHAGOOtTx+JHgwfPJvl3LMAqq6TUTW77bIqYHgkO3E6X
kx9QH4chu3ebEkrTlu/SXO8U43rRWer6HkiR1744VRaJm1nLSs5E7XRLvMd3P6XBOMmXcHz4Gpnf
OmTtBjwegCN8KmFxs5QYR2/l8yP4enayWX153YWLuy06JE3+6lE8qBz/dXrbfKLndS3Z3PDHLi1a
n43lV+IvTxji0dg311MQa8+385Bo1dMdIHHxzv/xAVQ5gGNYCcwGEYLlo6sQ7YpYhoo8tVDNXkNc
xo0h/LhK5PNfUDLRDBzrCnSpuRZb8aMomgPztwB9AtD3CLMXbJVBP2GKx+ZJVODZmKFRnPE3GhGD
tAylzhx5McRORyUvNdSg/LepcqT6q1zhzdKPRyDzQQs61ufZcBxNP5lNvuyeeVlQ6JsX8sHmZbxh
HvAXzz9ePM86G4CCvKVo/sKNBVSKltakyKeEBltS6T149KXKfWLuv2DOphyU4NL8BBi/L1Y2AU54
aQWnFWkkYw749snTOzKuOt46offU18if6oQlOyWdPg/ehskp+Qose54Pedl/gzKI2v/bAil9rUbX
e96QjtgCwJCZyU98zKuthB/Bczs26REXUswPFM0QyFVTSsJheVbNLaXTT4hR3KLH+rcgTiZ49bVh
vH3XqbO9k/QX4S9u5QLWExI4TNq7dtMNCQvoH3idLinQJa+JmKtH6Eahqnq2awyYRt5dG3JHhIuU
tHV+ns0IORwzBKl1hctoVl3RiHfGkEB9l/Lmeyw8+iCAomAdKzBG7MjZTFAq9uo4vC4m1Lw0TSEh
OzeQ+iu+N4GtR06mYiYDo7Lz+hNq4vvEVZfsCtLMpzJzyeO34clfYpy6rMPr4n2a/AY+R13S+tn1
91O3/PCH8UIOlbAltQKGcC4U0ImFmQ/pHK0CM7bMKxXkCNltYEgaOLq1sLudGJwAOLXsyic3Jjkk
PahvxbYDcXb0ao8aYDO7ajghnSj826pi/pP2Uo3rvvlZtdwvoxNKMZoPkfihtOwoBngagAjyeIFm
3qiEn99bn9+XVp1ze4wIFms8yLJAPDpcGQHsV5a7MWwjg54gkDRILxB5cnWLbs8RB7JN3fTzdgcM
jS5YbQ/e7DV3V7BAqpa9ZcAMLYzNSFlDUk3p4n0Tq5yzoIwJC7COY/gVUQmZ+X8xQEhXP79MyP6p
scRuUc4V5nXnF6XrVkMIzkxvD8PCoKfi+cUMvnIRH8nWNnx9He1FQxtTUxPCN6h/TPDfwDVjCKaN
+Z77rlQHqGKF83QYtL5YpXszMDmKESqLoSlkst9r7HtuyhvUVnpOaFqxOhkvzxM5IpmWUYxtDTXD
Yqf+oqiD2dn3AybqVn2KtPTqNC8B+hrrDLkRm12EDZliT6Z8CVu/NhGGrq0ll+kedLCT6QtfTg22
UTQvAr5+CQDK2mJJGGhc0PWVyeVJL65XCDhYOg7hJqFoxFhEXh8oyMSFHSgTz9o8aWNTSouzHKJZ
Vv17DqWvDbIrTuRmrx3EIM/Zwv9F7O0gwMI4iEX/2AoVRLcX2/zgJwkOtpZF+9AUqlqhsV5HvS5Z
DUcDi1TvF2lMpTkfMJZEZmiqM4hv75+o/xCOUACVFGkyoIF3dZ0pRTI0JCi7aOVH4g3a/l2GXIVL
AXY7PRhdJrauQ2azCSFNNNUZJWuKxyeMiGNGQxevgaJNWyVNB0oD0Cbe9s5YgEB179+VdxfyY0uP
Xo7QVVVY6J9v1N6LgtXFwY3G82r/BcoQAAtCU3tSSnpr8Pi2WHumrkZQ2q0uoXLSrj+IGZPUS5yq
jQDnmvKMoDsprvMhPsru0plYNHBhQtG9VtMeGBO9LU2JFxYug0SxJ8vCx/LnwxLofKXnKAOot/tC
8ZY/VQCLfImMa7GT8B/WPZA7+N95D3TlIuSE1T7YvMEv4Xwk9Y81joYjZrieDul09Ha/dzm3s9ZS
kIkukCs24Bjax+TMYGqX0pI2y8ozPD7H+5/02dKYdb6ja92hjOUYIMb555UeZyPbIFZSWs0dj7ou
Es0rr+jVLIb5EwcQmpu1hbut7tmMNeZaSE50zgi6j9+AVsdJpy1SLryjrLXyz3Ayp99acx1R6WFb
v0P61qYEdZKISp3ecsGJzecxkWdbpn2pmqvTvX0zVH37x0Bo41oCm4sz/8zQ0CmicQ8zEnoaq2rG
vBwR+dh1NWPf8O364CrvnUstvDDL+UWe0OLjEhN46+ZT2CB3JUJ4lng4pgdp5V5zijxL+E747Bd5
ih3xUlHAgSNQA5UopaxWL6Lxr7EWak6MfuRg4oiufxzrQzwjnXzVypabVw7CdiH3PSpiCs36FUAz
SdmGcaMkX3TcboZh1u4uRHoRZIYe38O+eedVteVjaZZhoxqtIVm7eVA3M4LqWLRvAl0UYYidtJPg
GbEIuJbXzn/FKhBn2Ka3h/2Lgy7RTZghEyryleMXAVDddVvxl7PkdUM+wkhIICV6nfoChLKnSDhw
1HODK1w+10cPCCplT/9b38+Sk0CT/aA8n3+Q3PvEn0+niYCB4nOtbZUdxJtTRiJ9KGLfwNtTZmab
SAF8oj40MpvXJHgl7V0VvrjpcL/OQhbThsEPdRFr9Edjjn7PCLJKE3q2lba1HglfAzliBD2TIDgW
w/mnP31PTNEerPWOE0/jne9aUohXO1CSaTMJR9h/Hry1BXVYp86YNG/774Vo+8tMkla8sH+/Dyuk
EU1JTp+NqrzBKylt6X2C8WjeeF4qgjQDroa0RbOjv3qCejOcqcPk/QYfiVRdZMvRIc+VJUMzv+zE
mdG7hVJvEfwGVRf0BHzpH18v45AUY9KyYPdGRq0geehbszoDtYvFqXvXXeenGkh5E8LHV3KgmAzq
IZz/x+MfrSAHvQtX8aKEceuwSr2OZdVs3/1o0OxKHZ+P1MwCr5r+omQ8jVP0HVS8mZn4okL1nC3B
3UkXCxwqgj6PwR9q72l03+FhmbRmZdkTWXaxn9yZf+QluScxyQR147vjJjVWLbeEY7zWeR+HiAlt
7roDti5PB+FilvoMM6g2STLHvhdLriLLAPyA70wvv/gWstKEJa3NOQpgWaFqQvo+JXhW+4ZniS+4
Z3kyezABn/xW3YxfrG4K5EuZ3QCZsAqf0+5a6IZgiOAYtBJv9L/lE8Rq4T9ljIJT/jgpGugQxMOo
VJw251yeKFmmOJH0CK3+M4Sy7JhrhIMeeDMVgym+xH0qhbkq/dfY1MlUnjRnLIhmzuN04a/TGI+Z
2KxWTFkOU9Hu8OTP96pogpehNSVm/ywgdg0AA7M1BKOzggnnVG9q0U0wp+fSfC/jpqS7+iogo0Z6
HU0rBbpcq4ucXSyD1hP1M5j3C3QrvqWPs4n3dbCLJugq0TKjzOaymagWSW9siMJhJvSmF3JRN2LN
TMI7/yutHastWhCVzNeof9KDq4tudRs2HQpaUFIDqSs3GaqWzgrIdj29O6TDvkHWjZ+/CSrP8CgC
fpIlo7tYZB9figLiU7TabEQnWYgrLjk/JFZM5IH/TYT9le3rqMVirXa2uKggsxsrwIt7CYDJvIVA
i/T5m/SDD15v+5rVw3mdp6UsU3fMUTXdLdWpkMyWLdToZC56l72HheLY+NNjUqqmy6z9Y8Nsf5Cv
F25OMAqGQ3sfB01f/vmVdPsGiv95IcaesAI2lo53ATwdQR00YsJXqZ6G8K0GVL3Ymd6KaN69Bpou
XPm/vUwSmNoEY4Pi1JwrwgmF0Vj9sr8UPmh8lfmKAjJwj5CRs4YJiUcmpIkoYTxvC4HGTCzfdAmn
2PbRt8pmVzLsUe+AtKlOMG6l3A18F/UCGsiCqwRpi5C7mr8H8jzQwB6jd8CNbnMnesGLjLFqlUXh
GnbPmbmaNaR7YX7xtUhfJQJrq5fkQ5R7aMM5atPNLrXFFrQSCLaYEoIK0sWS11oaDkWmxNgEM+NQ
QxKXDQIqVcB/O3wpZVDv5E0zd2vxVf9jgEPf9t2M6dDtYzkh2TWury7RjaBaW4yJxLSaYc2epzqA
AND++Uztu7hISS5dj12YCiQZ2AR49isHGmg5ZJzOj8OT7iIEaNBKHOaOOArDTMUTvz2T4PN5hIo5
VNpPM+0E0bnMtQIvap05qFS6L4wQbmBjjvIRv6Uk7CP0HPLlFcFUUJVNOOBA7pRNqQWH5WyNWJ7D
z+co0sJrziV7Sey082hPKB9qH7WjnuFY+8oe+wzvvO6A3QvmaMZPP0+HFCx0chYLju6fHdH4eYzv
8vnCvqRfXKmW/tRvZWPtfdG/v9fTGT9MRGV5ZK22Tk8j+lxmV2ptDABEpJB/5Glngm0me6ISCvhi
46PX19YxcbIZGXC/LU/Ytqpxh2pK9bW4WCVxH4VNIxng0DJ8C3aSsmtrJ+oTtyUfV0xySGVipoGU
JSdlwcrS3fE+yt/+ahpC2iACN3a/4balRMszMkQbM2DU7ycW4DzbddFQ860ebIueONE8bCmV0XqB
dV4L4wRDebw4YN/jYG8HcE3FgMrM4JieQkzb5rYx7pj3Tj2sBI1bZs/kVyH7pX2sQZehQAzLUvLU
aXZWegs/haqNiDmntSWY2dSy88+HHknAmmjLp9xS6dwz63EGkzJuJaprA4GtfFeYUufUipiXbG3G
OFUAeMUsV8kt3wQ5JzdvQ3GEnO7SMpyDTvEdIlZIc6sEfwNKiWqKSYv+050JdIPnpFwbM4g7C//2
R3/CvGNlElxsGct4DMF1DQyWTOn0uDwS+aagVST/nSmFAkIGp9lOFwjz8QBAX0XrOqiWIwePI+qJ
oHwFFSLIn/muw21wF+8Z2z12gLg3Bi3DvSlaTR5lzW98ic1gkQAqD16mUrnG3djjHRyk5b3zdquL
qwUoCsmjoE7BDE1uciP4+/Psq8EOk8R3HA57467PyORRKDsANAUfNV3phv1/FPlbmoTlx39WJ4jT
s9r1U4qtJL8EJUdKLV9gxpaLNI9tF6Vy6tXWXLzDY5gGcQyriMUNZwkUqkcVA/pkglMrKYhKeOul
9WoDHweQZW41bxlh+POWP+1nKOCR7fzQ7+xxByhQRtNIGuNMEhSGt819abWhkCgj9bnTAME8uzzv
48ANxQl3n45hxt46Pm2OF3MpUOUQ2PXG9mdmmNdvo6xAA253JTp7lkBknmMfI8JfYSFeKMQf0LO9
1vHwhU7tF/CoUrKyIJMuf61ak13huIfC3E/J/FPcrq4DT3VxCLlqA+k2PRkWhz/qQG/ylG2P7F6Z
CJNojyGZxWahK9yRvVkuee0CCXpAkzoiOVfzUg4fvfDTRgTJ+c0NYyg5F70JAZtal3D3MJJmTnEl
yG8hGJJt/KJqZyP9p0ipXjpDGTQkhpwpo4axdRVIoBPpWC7nxRqgx4YhDoD1oR1lyEHmPSqa6pjT
MQyGCOD1UDCKNsYR8r9LSPa56EsLNobHxaJEUhloYJkNf7oYXgZMCp/GRPdGHbYHIiKtIQ72XEkD
ujPatzTJi2+uUQgmBPO4rQVNr2qiQgI2WZYtSmCu4MgNRwx/8f/KAbX/hY6A11LlFS2p6hXDW40V
go/ALuAjk7NAghbp1bxkwkaLHshBWqpeinrSr6owj5y0EJvVvUiwdunX7vGNYaxrYGzkJSl9nE34
W6Cbwjk3MQibuDzssq/4J4m0DLU8lFminJDaKI4RFkDWsyqKj+bpZq7bXxXeFRa8aFdCnZR9u66M
JvQYqNuJQ9pFEQGCxtsFaDM0+qI7twX197gdpJ93T4e3RSw5RdA2XHXez4rg3eJI0OVAt/Sy/FL4
TYJaKMz6ZhDCgTp8Up5LUnPiBczt54h8d7k2EaAtp4zSDNsr9nV/OMPYIiZO92bVRROUGJQg9tUH
68YdM3n6vMemL5+2KM3vpVlhwzH1O/ul9wg+glcXN4yUKpdfHpx4h624ZfMzdoXtCbmsLHce+q8G
dNhtq0OD7dvOfcaj4teV+fFIxE5Z1NklwzDHNy4gkh0QbqNNcfIAt8Ug9emYyUXoryjXLwXVRMe/
F8LpNAEFQD7SWykKqgtoHvW8ZCsSSi2rBgoUZE4feN3sysYoZaOq+SVNIODNrhqyXD/zq6eVmPKh
95+ytHpgiEpbUr71L/lj/5qVDc1OLLsrulx7e9h6QZ6Vc9eFWDGtlfV3UZ3quUA4cVsSGiUOeZqX
FOCQGvos2AteOQoCAf/748NqDzcsuhHpX542yM6q2TTDye0f9CwpZ96JCzJZBjr0L7iv/yGkh+gv
t6KGkKmH1Bliziz9xZ6uAITwRV5hsZIMv0OE43N+vp0zharPFE5Vl4e2bFUuZViPT7JvDLudm7QO
/xTbqbC/HAwLQPS/dbeNzO6SDJbE+ooL/G00XbRnbJ+qGSsLInEbDXdf2jZncpJkMUNfsFn0S0Ng
8UfwoqNj8ma9NMUfgJRRvR0F4Op1oyZIvH7tVkonygGKxO7OgeIid7bXMmz+1O9qgALGRnYbXPkj
zMsHg6dLc8qlMmbybjZ5RmS6LxTpSrTp25w8E4fTnc6EYGDhx0fKJq2MwujY5YnX51OBWdpKqpmU
2KSBv5fpPFRAFnupVqA4OLIgQg5uvZ6nn3g+PoVLCUMTWynaaPGNCTf0zQGc0bzUsOQ+smwiWSej
DA0G7zlrpjMlN+l0yz/QNiFuknmTnYKmaDzq0paQvrwszIJBufLGZuu5Dwz3KeY84c2f6j4ozrUg
/ZcJX+qTdiekI2OZ65OKx8utc5VydIg1aBvI/mLFjOxRFz5tHJ320Drv+UModEJ9AzdXyTcD1qVB
5HENZr66kC2dDBZq0S/USws5ywomkagz9nPKMr1ekv9hXigH/ZPgB7DUNDzXDQ+i4zBiAdYAO0A5
DEGA4qJVWT2PRcfj4s97Z1+fi+catzCcMsgi6A247s+K8CO3/+3yYGqqcpdqixxUB8WvWkRwjYaI
OJ0ADMqhUfzlWcgaimlP8aZqJGGLX+sp8pgQL5huxfCQ0cPa7E7yWNzjXKr2/4Cp62v66S3sVXcm
6x8TTHXrdFBACz1lFxR287bNh2io7epA19OkK5QmZUZs2wpk1uU82hgD//g+3uwcORi0Ewpm6903
opl99ouCvgGi6mqwIsMD8aTHyX1WQW3sbw5JQwL5xji1N7tdZVidZnzP5YG6oQWgOREFn3IwlWAs
WXrEH+JOnE9AAgpTLEaUSYBGtBFEh8jP1YRHgJ5W5z15QLEbAUol7wnmANXv0AiT+ygrzGD4kvtV
UgFo/QLqZhT5tX18034s2ZFxY5t+eR9ZBVKduhKsuJuifrX+YU3VsgOTepyiMSpABhjKvcheKPGv
rk5KZ/bpufzUhcwymvIL4jiR+LLrKKMQtuFWYvtO1axEP0mDHrKzkjTvQhcAbxDz01bT0hGVC/SR
Cm/pPbyhCcfCQmRyNG+ziUMwIaqAHNNzPNcLn070BScPLNxV0XwRvjj+AqpkRqMetmN1d/jG6/6/
iFUNlziazDskya2dsDm7LrVvxWxn15xIGPSdo1BsFBhjHr2AcmEDqxQ5AJmkEW6etnQ3EfahYzy0
GRhvp78j+iWAWTcAU2I09QUWmpDFLhIBLjHXgliQSgVogOC0FC4kqaBmIuRpGahnOJGFfCcVQY1M
5KSDu2EpsD76UT4AuigKbC12pb4oJYcS1SsEjeOnK2HFU2yj/MqPdYmzfpFEkDWy3bsMgmxN/PI5
1Ff+4RBKrA8RiYNgifCyn6elU7VAbksHY6NeB0C+QV88SlTkN5m9xsTi8qcO3NQzrz7t7m/68PdR
5deMw12dsqPE9DrxPn0+X22zxd9C+f/MvdrtROo+RrSPv1xtdDtzoTqnEGSnugHAPmUQd+Du8dqH
1j3CFHGOz94XBj5Jq1u7j1JJwjFHfq7STJLWipaP2pVDyWaMmE0+SglfEbFIPJJ5uOeoypfbhECO
VVPjvM7eiEbjYCkoJVKE3ZfBIUjsb9YroRX/h/unnq9XXtUQosFttAv2CYassYqurucjcVEqN5eM
DmMv/dDLVbu2yV8iwxtihS5mDevUc7AwU0u/ATszoZg1Y2caccmE4nriO6DYoWjycM9LomqyCjFJ
FBtkUtAAvaThkhAT9Xy1fR8Yz4sRJZQAw4JpxUvlQA5yQF1kpHHQjSzaP7U2i8dkgFuxg2Zy+D9K
YCS1v8MDWW3ng6vpW2lW5Mk5jVGH/ETA9DkoF1ufYMTBCwpjhNGGrn61sZ90BWsnNGYsLXTSPNjH
EjmZIJ5iFiGrA2DpdHq7+CuTgPmRy99pExS8YoWL9TkA31bBgKGYzmt9nnKsNmVOAbPedQOeqhxL
3s0tXd3MNwZ5mtzGUZG+pIdUYZsK9mQr2AjNSb9yUSEyczxmrxnpg5Nbvvf7p9nHdeDgKGlhZ0WR
mckl1y4dkXKVIh0CAof2vf9KvaGYIJ3VcLJyWgMc73U85vSgLeJSY14/cW8StGEIp1JauGSj9WWk
bF5DGkrEDyw1byyGtTdlxU3fv6ZDuPHAarTRIgt+obHYyLsX7w98lk1qVSygxafqBEagM6H1Tq9b
wMHZce9NrSgcLhizOq0pKs+0K90lvbidigMexvlrGplCSRUJG+m4mXcQGbPFCbnaTZbpMEPtLPg2
3XS3FUN7v4lFppGR+fjZBSG2SjczkPLxmtCPPjj4NXaVo/QaSSwrlGAk8lDEfhQwzxhzrkG3s40p
XSmDMJi07UUa3QM+VHSniqQii+z9MUfhmAzAdqK0v6NpYI02yLB/nhggoTdDamuf8pLspFMVgnP7
O+2ujwMIQgFA5tLfb8xlp+CddhtVA3Wv+eIF81EC1LHazf4HG/vU9lR/CISndfuyQ+jeYoMqncvP
z/jgab0egCiH6ksg+d95hQbjl4IFiuZ5p/+7Q3RB+scJt0bobWAQ5KUqGdVetwO4I9pOSBtiritT
vvGWcpn2kWyB0iVXx7pa1sLQntOy7OWhQDG7pXi1y0ZPwa2utJHe7+Gy7o/Z5Ou5BjonKptOU/3m
TxjGp0Cegm+kLwoQbsdkEMn/anpH3zL4jvqYbuWAsDvTUXz+hVJTxHIiJ5d0b7oJwirgvicYhez9
AsqnOyIgMHpJYZwZ7zD69Hpkg5mp8jTNOYEGCEIiXXVLhYwlpESz/Vp7oZa9PywA3mKqV7ejimU4
DfJF9183bY2HV54vsdPtbLY2dlSdDVQ5s3mboL9XE7+Pyhu/8X/m67gZk11wxMsly6QZiKTemIpZ
VzynfxExS6MA9YOYdaTKSE5aVY3Vc83sl0EKf8OTrUydrKCOjUNKKV/j+ZnsTwvz75G2aNfS8ML8
xghLeUHqKrLmh4b9S0/V8089JfCRbIlJbCRN857ZQXRCp8JGDshQfLYr9efXPx/27h0Q4VE/owH5
iRqqAQbUawoIj+sRuikWG3uR9B9qRhlesVcPC4Z/t4cX82fRbr65HSiKHicsfxZ6R8mGfF4DsrM0
lj3k7Tk2c+a/qDKK5224ItoB6QdioTQRy2XlYDOm0hW4opcugXthCiRCtPlNnx94jQDb+j0fSB8M
Kc5dclGoR3XCoMD8We/m6Q90VGbH85FGWhIdinuxdIjWsxicpbvMnp6QT/pcLK5izUvEUY2XWPCE
L3FXaZY5hm5T0Y26OmhL8gaSlKir7Se8XJLDSAt2LGGD3QfZSFXki6XnV2vpc4nyGoEaCX3c6ytU
PHnuA+NGkrdeyPmDs8YezdfsNtnwj55KmJZiET7mtF+sTiQzIvadWiDLCAnyfR17XJsGMFUolAsU
cK8DjtYReDLuNXYwYoBLESWBWGyQFitosBMUJOhsx6lfcQ4CPeBLtwkhZ2GqDdNI3QqA4P3c4XtD
jZtFcRfybWdI0IaW8BFjo0ujR9eD9vEINWg9f4KmTR3NYANbxTsUtr2YL768aaLqmQvPO858hrkt
tpew9Z84sjpv43t2s38k8HemSsXJTks+WRpZM4cVnYfbMb0rVaDK6nuVeITntFpj79pX9E709B0r
NMsfNNHpV3jykUC6YFqp936NVGtpi8p/4iC9V2d0FhSoWhKdmv8I+CwH8I/P0lfPISv60ESbV4DC
6tgo5LgVGOJ45EFzq18IxTsnb44MF32OmuwNujpu2LbbHnY1NVlZzLOPM0koA4IFhvM2V7iRygJE
he3gYOaE3R7Awdf2TzDKhkzbqlSEmTz+WSzsTEP60MM5hsY2kBjD7EJNpq5i8TRtmEWn3H898wyH
mzCZNAJLwqOWIXHh/81DGGIlxJEW+qgJ8oIL14PK0IT1jFU51wmoMzhkkWyn5o9YB5wgI/VMEpir
kvdYMmmXe/jYcApd1nIV3EzOAdKDi+Pe9rm9bSvQzFFEZRIK8YpWQeiNpeI3iEzjR5H4l4yrEbtL
/rX/xlp1HZxcdbDJ9tdwRCNl7yxhx+/j0WHmw30HUcs68ADqt0DpN55heUpJ4PilI5864k3793Qe
em97TUBSi02y81Ply4aGHL5btEJRhq/jxRI2RQYT64hnQ3UAQBK8U08yOtJeci4Zy/ljKkV89z8Q
VeRS7Bgt9ZEa9zCWkMYQVuIhATCXKCdR4SwlOnAa3WRFTAn1b9GxKZfp9ATazAskAvNPNIqJ8gX4
F0U4lGNw30DFMJnoUyog0qKYe8055970j4+QMMrQ7R2yPSpp8Ewfk27dxOnXWNEKmcD0GD0A8+3L
l8hhO/ATquMcLZKpDe+D3ATHxw5n0tgruReo3I8c1Vvdfqafmv/X1Z8bJQhfgRKGFc7m6+EGE88d
bS4JcWxrOib/I8QkZ3mbwIBZ+Lqfk9lylMeabvrtX0WCw79qXm6KjX8mnlp3y5JV5PG+6bwNrD1+
thnYEHoQMwRv8DO2o5rjGfS/2GMi1yyPXKkgF3TZC+a75Of/qUuV07lOlmSElUByP55vbhFWsdDE
TqmoswUrxkkB5ruNtXlHAv63mFV9l0s3X/tT2WJT4t4xTQ4sodOTY+IYoVlfd7q+2OWZAmtxM2ux
EK9BJxZttwn/9GJ+dWccaMorbYE1Z9THJ/Q+mAE5RAVbb6drfTGO/DQJYW38xkcwLbV7/dEl8fR3
+qryLwxQOXdZPBji9muu1p7FLkr/GCr2vRTjLG+Cqb+Mj/k+jcZEP81DwbodAF5yN25jeY32zLxm
GsF0jfUBaWtA5MjDklgIhvT4Bbx4BOxS7ZM/+Hx8bJRf+PKCvGm1sx0fI45ISUeVxQqeUmbf/oNf
EzGUKb1vXvgs8MgtwqbOgiVmK+vnDoQxJAIoGI7XuK1xn91ZkXwXBsFu0MQx3K6+hxolMH6KBcoR
ZNZaVR9bYxqPpUGxes0cqtvcwbYxh36TntAN97mTdf49Q56VAL3QUxUqFedeYL8S2oLyDygShEGW
j5fylfQT2dYtQ+3MGJsD0pF4jzsgvAE/pL+kQmoZBlYwEgfYoASz/zo9UsU8/rEylPahiHmx6j8H
BCLg8hPOF7s2VjdBGCa1gOFw5ZQ3mB5Q1tpFMDyfJjihtdThujKqKiZd5lH2/x8Zse5BiaQGujaK
LSPJbIyTTwO1A5mreWO4wHfuXLUaLQu5HX26w/Q0bHnuNMWznLE7QZTfSjI1OuCR9HebEzin61rK
m35daRlaNVO8ClRHkCd1Y4qbJl8ZhEDuMn4UUzT98YI0SXS63O4qgyOkmadZc4nGnYElCfnQ3W2U
DUpjZ1yxoSNoaPhOgAmA+NPpvaBYO5kD/nKobm9IZWDgcTqaSH3aVtzYXCW6DF7hX9IGPCeKSJED
fCA9FD2/7K9ESaN5YMAe87EFmrclepaB5LrZEyABWlUZoz8JrjeFV0djeX+Ggq+ImQ+/uC94aHyl
GEWGVwqJddoNJP+tcDzjmljDkwrFDq6NFTah+SMvUh78YsgXEH3fCTljbxkpFCEy9zEgUepukLTR
E2lbYBcJNrZB6xcms+F5BOG0WUr7qYepfBoQoDP2uTa045iQ+fe/yg5Rb2kOgr5yaLtSOoxFCSHi
Fvbo/VSkT1OgkF9TPaC65qVihkxlvGRnv1hbxBwKD5ks/U14dK9KMZuRPiwIoDLdgYoYcpI4TfHF
NoH5Nf+wKR9sVwKJ2gETYGFRfvIk53nxNUtqqVK1FExV+cVo5aXPE1/4frA83mROLLI4Z/OgrZgq
KVTWA3k/bakCK1+EuWnkYKmmRiYqfYIb2RBgPLOPdBK/7DwcEjvdqPsPX5s2a4o8F5cxjvTRQ381
TFexUzuqmuPRGx8pgxxne//rnGfah0OtfVMpUZl2xmmWjHpZsM4sTNfk4vB+M1U6t+3BmdVGFmeM
Z6F6jSr1Ck3LpU4ncZQZZrixtfHSKuTA2RrOv9/t+gSOFLYH3bM8BZ8vIvOjlLCcEHHk+NBKnS2M
z5PF4uBOuWwDN7KGoB6FM9jItRZ4hhbBjFJOe9La0viq3fsiywYAvm3skJl0q1mYruL0qXQWLEEd
uoiZ7QWA9a1hrhjEaYCv7jh8molwqf+uAxBUP/vI1P2WeUkGprifbISp3HQHhIZE2SY/TkbsV2OI
A9ynwlApq7+vh5hgk0UjVXoG9NlkSWC7G5exW68IyqqjKCRgtkUYu2PM3bRG6LzQvNMz/5e26bRP
wBazmtx3P56RW2t8ToTuSmp8ZpmSdKwHy1biY4DQcmjdo+TpuIb4otv8EUzc/H58AH8zQAW1+OJC
xWgAb+oOEcMYFfIdln/ULDOV1lXEvEb1in02KUYy6Rj2Gkoklc7L0Koa64LFKMgdVeVJGsmYpFHm
DMq8Jqj2eI6oJjgWOdRzOofyrg4uXu94EWmCmVWk3Nn3KQPxETyKPqMjpa2WelCSQ4ODvCSFogBL
gSLOEcz2xbuBWmf6KsomurTuOsZhGW/MLYD4TXVdKv2kCqbThqSdQ4nCV4Vmmt/lYR6tU1gb8Fqg
fmNnBp1xQQhtdFde29rLQso+X+EYb6LGLf29JkxK4h4qi3NiP5xmuNp+mrpjOiHpQ+uOgyafuCtG
djXhCmNK1sijyMs8TePU1z9nqLuK8XxEhaeLayQrHpuNAb+CsZp8IZz3awEnSaKC6wPVeCN2O0EJ
RFOqdaQonIY5UCxJpElDCbZA+2bgYP7YBTH430cVINhtVeTVjYlt9DPntMYXXrdqahzKq1bVQYJg
xgwFkxi92oCXZFvFlHKDYQz+ba2Tih5d1BX8k0+kuiG+1vuSw7Ssd4Xhi2+aIMGsqwPYkLvHO3hX
vwWWIh7upjFyLmFqTDUEK58ys4UdR4LfZZmpeKaZfy46n/aaFt779cX3CPgV/PRvIUtG1U/xsJQ+
toJDNQjo3/FusE3xgaku+PFVgCyxbsIGhmzKWgTMwUidJYGZoJgwrT3ZgZP7eg2Tvvt1nQUnHUwZ
8nbPbgNuGt/3+CjFqm43t6jFmXBJkW5+WcmCLSGt+1heetCq6+owB+IoFezugDz4R/OskND77J0g
DcZIEzT+1q0oTQWHaxYj44qj/7qCjAsZOgHa/iTEfl8+XwdztKEnpruh8uFfeseb2AVWf2hp9/jF
1EgON37XZpbW9F/n1WyZglJZj34/+5Nz0Nq90qYBUpqdzC8hrJ3X8iiEMbmxB4VdPB2I0AVrNaNQ
cujzJoQ0ALTMH1P4VHaxAjuh/2+/dBqzgLJK/sOgHXS6IIKknWMhXdc15erfn9OWkCFQ3NFVoEwe
ACQGAN3YKJqjX5PsaD//CWPkfi8usKimJXj+srJ8Aeo6hnHT3mcesSA2nxFVIcdkrSTsA2iExssk
E6HMZ+ZduL1wzFbf1tHJ0yd9hEXUl9KcTCB0b5kvJ6BSOWw/nfaecnJ9XT6ffLVLWTSuHmlyz8iB
8djPq/15lapag/7ylQvehcEiZ8CMj6Pj6dV9k7f2+lnsuIxPvL/ah1kiOzcerElPKbxEy23KlOrP
T0YFc/0uPfV4ZqVOJJuPZb/vCLmvLons0fSEursWyopdBcUWfgMkpOrr7W03NVqU4VJitBFPZUwm
ybQuWMp1p1uKBAaVCGk4uRqEbsuJocar7sR99TM/65WOg19Oohdgb+FQqqXHRqSwOgnlFgO+Nrnv
eGIC/2TQ3yocvVH8nKKmZ1dr5ZfCG/Lg53v+PPEVt+c5WmPhE+mEzwXrZ3dMzcOefh5MxCoWKlD3
GIaYg7TEpmRYLSMsUYcl6ShvF8hnJmb8Fdbm9OeTrE3gKMsPyuTmESYHxDeiPu06iDlCu2Y2L3bv
yzwYW85ejpaibyiyXYvbZwfYLdB2Z+ELBmnAEhrNPjTOOi8BhWWg6k9LMnZD2uuRw+t/ySAPAwLt
F9d46lX3BbG20gEcGkBz707TFHUv+LfAY+rOQ8MVwcX8xrGeplsWDu8CwEL1RCz1O+n4eROhVe99
UVrP0U/k66oV24fIdhoXLQi1nnhbbsuNdndm/a5zeeYmMbCBord0zlnNTXj+F5IsunI8aYepeeU6
mGz9gEQaWbcxUJnC1rZCSeplFnxqxlhMvmZCkoLwB0MSmMwPzqgZG08JJZT+xpj+WxpYRDf7eb76
mw9wy+ORsAEh644r3AfhNYS6G9alm1452bh1zkYM0tj6tdIJDgtlxiGehoVLwFSGgjGXESxkbGGJ
7eg1PpLTd+OQoqdQooe3p4n4ObFz9YNfhJH8KGrDVMGv0nU49jfSUl3JWniBbX0iRPgv/8yxCB+Q
hxMXN8tAJbE3xC6EOpTuPIxtDzDEnIGUCdqObkI+VF1fjw4nYLUbJ+/IdGZSWc75Kf+YYQB9EfEa
+RVRbKWXvAPbDDLhviw9gkBJSUtSzNvzEX+tbUaZKCg/sEcm19LridJJ72gvEghM+EuIflp0Z9jf
ewJbXZIE8sj17CBgE/TE0JvOUwzJ0xIm6bvB+4lzKYpAILmY1Ftgfz+KG6X4Q9n3hlGsp/yNlbmp
RDccUCQw50OUwklH0qwFdTBRuHOmCy02NUJ13908wNTO0/fcZaXEmeSIXtg5tbOmSiqH/3VXo/ft
vNdVWnuSTkM6JtJ0Jr8aLhfK9/Sdz68MBypXaD8O1Bv4tzHVm2+/Up9klVvuLq3o12CeV1itwHed
d/EBcxkJ0KXbWddLXpvdc4KMhZf99UUvVchZvGWy/+9CHvU9qF5veexwOjQHItfcw4A9ZLskNWL3
eCPc0L+aoEnryuRd/+PMo3JJAZ3L68yLXkd0HnS4z+fjYQZwZ9SIrMEL13zVyDY584111JW2InhM
99MnODSOKR1/VAz3I39yx9KQUtWi8Y4tKCzO6pjPNzywPGKC03ix4owfAEKF+M32ZFgBytu35WY9
MVXUV9tdefw83l2DhnSDfdRhqtICPm+u9iaQ5ZK+wku2pQ7pAAmeHIzwsz/3iZP9gFTtCqKEjbFo
4PIkFawS+exO7A8O4WnCFFh0Z+0GdGX+M7KO3jBSygjgMtf4LyG9zKhK7lyQ5/9K/77uSez8YXs8
zEDxKaCdhcH2ZyD6JuXIRtp0qSXpcgKynzK4QtXnbhHdkbj72fRZzd0qZa//M0CBQjURz1fnG+bs
IH5hK8rxEEiBWfbJKU7/BKl2b1kSaMjkq6n03ZXf6zK65XXD/BjjJx4XFnmV9j5lQ7wDGxGT1W8v
u7GJw9K6rmHsdYGmE+E/FJRiJ2XJROZwrTn6iKza4vxL/0xgoT9iKKxWxiOygoy+FNoJ3icdWBte
RznG8FNRs85A1AeOzvkKHJJvgSGSZZoAnM3nZrE28POHT63yGVydFkef1EHHdebu4NO8yVuGKzPZ
eqMjEMA5MM17P/CyJTCVnSVVrYZ/+NEcHZ491Pp/s0hOHRMpCIHoZhlS5Bpg/S05PXse3dmw/cu/
0uDgIEO+0d592g4cv0lBgHISUK1bk/BToUfmZg3n/mHzTLdMpj/6yp4rVfkUxJbT62E1qFTUNawI
WqNWVvm/nZox8LCVaYnBIFYvA9XHULxzonVlfM0HKKnbBv6i62t6rtqT+HZJxH/UWiyrubNaKspw
NvCXn+/uA8WoAyfRN1RcRuYgd+kEhj/ZdmforRRbgg5l5qVAw/pBvlfSuQkeoZQT4FLn3QQ7QeEf
dG8Ov21z+sNpOADPsmCKOUzo+aXQTLy2e7op4zubjUgN/KyE+RDBdcft4kBVSucUy6rYzqb9B+UG
/QIiwpNNHprDzBHg5DY3uCnoKBohoCL5tE8TjvGYQUGahzdy6wnUQiuKRs9qtESZVmol5i+AFtvv
BF6eYD9O1liwAAXjMc7Ojn4NsHGoZFrT92oE17NNmSdR6kmFKgbIhrN8Z4WnImJsvoNUccDcOMut
/htt9bGnIMZ7IRG8zsZkvHABZN5w1smjf+/AEPn4Fo+VWNsgw83e4uTYk1xLhRc6VTW3HGPaw8ie
nXp7weXqRXkxE6soQGTt4Dh/CkMlFPHSW9H3MPMehAc8llf7sBnO2KIRIJi41nSrKAQG+2QlfWZE
Jg+viMPVJVOyKg1JrOOpeq3SbXUt4g+AOGJFao+ZiApUZUiOw24u4BCNbUFTCmm5U9ROIpLQn0An
NJ9hPeKbgA2aBz0m9yi2yuifNfKH02BeDamxFJiiKkNvncE4m4/0v5i02DCtimHvQ/g/Nbf/GhyO
cbpmJ4Yha5yaN+OnHqwL42RWYb/zsb278PJhavFQVqE7Rz2HdICmmAdhcOuJp1pjyMkU3/vZUPIH
KAg8fB3EeSVSMRNGIUeLHc+dz3hB0JOs+JyLnnvKHpFp09zdhsbzZSjNh8NPgubxpA/gpSidcXk3
X8WhZYjKYYz7runZrHGxwp3wKo9pAwUKxDws6w6/NVfcesO1WYfZT3xRB8eLXx83fLWAtSj+QCbh
K1yEYQtVhRIYcI4Ps6zErbER4BhXiFhc73I7ykCuiw5ec3jHjUkZLkEjbqIvwdBGIK+RItugjwSS
ABIdltQUEspX0rBIdjWVg6NiQK5t7/iydifmhDvEf/fUyhqT/bCo6g79jkQVfaas1Jhm+5S47c1i
c2zMDmXgt9VWnaSnGTrXShncFBRcojufwn8jlXP0bVeAstuCjazPUcwWB2u+4+0C4gM5fuqtIsab
WtGFu1QTAmtfhOauVS51cGwrqDFn1zDF1i0Wc4g/tgEgHYuUwbOVSP9+kVz344waVHuEG2VNgx+t
AAGATC8PM4UXnbUdhH1eomVLoyi15OLJQX0e5u7UT4d/ggJcUoNx5LtGSEGUYommRmyah6zZ+11M
Lva823gZv2x8q9ZLYjZkMhhpdgno6YEW27/YSvPjYT976tuJwf7LW3pzkS2WgxPA2YXN5IseWmyb
IIeH9bsAnnF348lOAWo63EdIMEioJQlyFkMsvaVrTi2P85o/fiSkUiZHF1aJ2Md8fL0/XMAn7rUv
bm8UKvMhEUutQh2sgPB60w1uIj4yhiMi/J0k6pCHNy3FF0opwgmtv/4mB4lT6tSR88WbA8S+g3J4
O7tjBZ4vqN5bJ8LOG1vSADdN5W3p1Ng2LAvtuokfvxHORu18IsONNcDDWMVx5hl5s5SVrDs/rSZM
LKw+wEgJPYHOLgozOw390a31WW4tv8lvTd5YHWtO9liZAWjSC/WlKwpRyHJL557bvMevYZqG/Df7
2pAMkvNHXTqskXzNekSobsFlqJcJi3qe8Xd3QNhHohnG0JdgNaH4SubOwjWCXEVwR0VMPTGuSiXo
ERxC+60dVY9PLdYzEUc3M0Lt8CpNCUEyO7f2gjxGZXdaHTFCPi0Nmg8FHZILwoSvp1NpkZ4y2uSt
IkRGsrkNB/Pa3leuP/nGKIGCu+cDX6brn27tqf5Si8kx+1VtMLj4nL3HKd5ebqwO1J2g8r4hwcUG
cVRJKUeD1mqmrtAOa5buERKpc82P82WeuS6a8wrdpgw5v0PBRo6KpHiehpbTKsNexaZaNEvFI6wa
mQ/YRbgzI9sEWvCnoa6OvC/4yJARvvmBJTFRZORTnoOPRuyz1Bq6Zr9anV0nvMgJj8RZ5Iwb9zkn
IMyoBTROK2KLaXmQodRyiFt8KBIdOYqWHaDEuZso0dVv6vKfuh3GlkZoOUZ+nzAezEZZAKaxIDUz
cs+kd4s/H9tmyx+1sbpHAZQROj9ZF+0tyU+siCjdGk5umEuH90NR77Qhab6rJjx1ID05JrxGek+n
aQXzMn0TvPZN0bhPJGpUJdzUVMAF11HT3YN9vAWvn/s5Zr6VOlfHWpkck/i26iImq6Vht1UMbEDl
nKSEdWw8uYwHwo01t6jBWLukoufvvdB3pqh2JSeMugqAm9u31TYlpEaBA/06gy+ceyZzGjzSROZy
tGimlEvjkp9+kbfv3MAWnhIMoxxLWqq+xp3vT59tJdykPzHt9nXVEJjWFYShwom4UNEgiBTCPl0R
1w1u4x9uKuHunNaTOyOnx27lq2YjIA1CpQw6YMsoMFXIi+VrhOlLnIxuljfBA0qS41+RyMpYUfh4
EzTV3CZo2dtJ57n9nH5vYft6qiUmEXdip9wmeJK+nLS0zSvSEKdJnCcy2+QOFyYKyG5okO8QAjAE
LvZ5q9qSRfB2Vx3fbzgN4riANk8E4vPh8oAcDsenNbwyxxPwmkhxwt7RG0wI9S11kyGkVN1YC7YO
BhcrDYxTuSmcgmh5wEU3vxny7vZq75YS7+A7sqCTB67bb6wBJlMgbRrR7S+MxiSs3y2UwVlt0cxL
yXhbsJ3o2gMz+8e3QSfOBADzDHHTdc+wr96yGHZXXWLCEkyDuo6CEbt985yu6vyPZ5WZUVyQUKBq
guAI1HQf4QImtxZAruc/MMEQZRNdGNilCFx97gb9BOhmZnVMhMSP363nwzXeNyjP0wiZ6KAGQg+/
Inx7It6gjpsUhEnQWxiDmLfjrrLBAsdzIDaqQdCd/WoZ61IjMC0KmefA46Dpd/QYW72gP0as/Pz1
43+ZeL7z3o6ITJdOJ83+7bVN1gahiTbKRE1KiPjMuZakbgUkC9RufDK9DjFkflcma0FQr5iwbY31
dvUxrPexN4Xb6ZtgZjLwtSjylbs5bNAHwhTRdFwnzU0qRrYXTZoY0y+ASvoXDWDYn7lT9i4TixR+
FVnINOkv9ixGbivIF0BdaH0cgj3fB4uP9L3Kf65FrHj71Xe7P7aMcMtEzpjxBpE+rTNrCdmt+0MS
NiNtclZqNkgSOrrSiocSg+trNhWM2mw7Zzb//VhWYP3T/f/BTO29ZJfXs4sSzKvqSlMF54ErBVIg
QTi3gxPvy6zLnsZGhu8A5RnWRq6zf6NmPpPMN8ov94IVCHzYynWxj7TSGWMOYOL5OV3BvQl8OK74
nKH/dp6wCqSarF+Co/bfzAM1gVaz9zQqxWqj4orrtj+fBWinGvVn+OS2GQlFAnBrf/qUb2af8Oq+
MvEmFoRHNM9dv9OKJCQ5Egl9WA8lkmFxSga3Gb21XE+2wTgaw6EJK9apmAOH2JgSOte0Qrl1gpcO
xAexbU+neKYHtsSGqK28hwJeNViF4awGlfPbJE1enkvQPUI7ELsyU+oLF0dwjHOjFGtCNuJ0UOlJ
ko8H8JKFVGUX1DN8ub9tMHLlrjzND/BQS8JPxU7oC4L/Xqtfq46avV1AYffyGE9B3s1MrPz42mNN
xKuhCimRjpYZsWcGR1ShDncZpOhF9unTZq4aAm8mvlwcVzBRHC0a9gebwgjON5wX9TxkOhwgB5pK
IPzTaJday6ODErgDOW2sCWsfpZhVhshX93wvPLMdw8GRGXESdr6kBLkAixBCqi6WsItgIak8+DvX
HI4EoQiZtGSfXOJqMb4VHECz98/k1xjeVG1LF1kofThbNO+Kxk86m/umnM5pg33sjlcxjnWaKWbv
vGBPla3L9sKWwDmKywXci+e42RNtEo5fdEHItLRDgcjCcNtOwdMha++IKd+HD/mCNhEcm7T+5DV7
Bw6tIwXDm2ZuYmlavN5fOh/to1rXn78XYhGjmU8p1TOheyJeau4me9RgTDCGQVzqonAouQW8Wp3n
lt2upk4crvZwtgnmwiKDqpHss9/TdTnaJ8d10lDpH5o34uthuv3A62+8b3YHp7CmzH0BtTsXEDUO
oko95xpuHUa0MRpFhWoG9gjXee0lWpiteq97b0H2MPmUoSF0JURDLoqAdLT4bQMyBKlYpvPB9XYG
Iz+mozjTFpM6Hp8Na6JfKJH8AF0L/alszCIZyTmq0b43+XBEjKsvJOuOVBXWbhv8g0ktc8/XwdeC
1DFEuWqKwGIZDR7c9wGlLhtZ4MF7u4tjP+WFYMF86XJgqLMGiuy3NYVeBYLPCyJX5eIuPEEHmWDx
NQPLOwQU7HlUrOxNj1x5bKxDsS1nbKYchXir9zlK3msNmq21SuZQ7E3epSHB0bDFzNmBvQr4h2Ab
BYpN6dPqlhqwV5uNhU04BuUy7+PgBPuhXuCYFuQgIR1IDyG/tqsZG0ezY5qsMAew+8B9Z/3djTa/
b1B590DeUX2bEsyW5T7r5GMSD2BplcCUjjh0CrZsZfYBzumUyOA4gp4vLqeehCBFyHMeWNAcDgXO
E5GaC3VeC/R8i/+q0maTh1p/KainTAX7j393d6/XYPlQTmO/csXxJ8WlYvSb2sezvt0Sxp+S8Xd2
b3n7RktDWNKPZ6WCUof0SQfqV258QuRZKXBtinaIVrc351M/IQHsb+qUxe3v7qAYnA4w08br/lvG
XedosrOyU89/yfT3ACs1e7kUTBh/2JiyurJbr9CBGwQ9J6QJnY2SKhSX+Dl4DzB/TW4bOu1Omb4y
3PMjLGYPCqOmXmWNe2qKSQpumyMplI0qdCjs9oKfLrThzYW5qLmITAve5VSwAE9vxvymkHY6fAKW
VdqoEsoX/iJIzaEvzTI7Ih2ZawzPtuwh7qvdrckzWSuu0ZYWLRR1Pr0xEGl7InBNkBQmKH6E9JG7
kQEfMoaghqKjZNmUHXZMiyV4PDRj80OJTI/i4X0IN9iO86/+N85TyM6ZmxdIJHwMo1P5wVYfjhxl
diCiWiwoRrAdTvxNQdvzWjTUkVOmldm6HDuQhUkudt66Sl7H7GKVppw+42olRtt4qabchytRGNe0
/t4z+WfXkyAgD7712qKqMeVDjZL0OqVnCX1xnp8PhYrCAHSbRoWf48u/u27U4+GNm3UaYxPrRrAv
ip4PD/RQbD1xfBe7XAAyl1ygodAjv9AKXYwPlD719Hgp7uaXFelI6NU98b65zjICSYedUxZ7D6um
qSxjil11dOetZZmgs+FDvXRiHkUX9Q1/bij3ysp9m/68+oUntOH4hjYiNYnk/cR+cpAY2frJelJx
L7oCyNpatLVdseeuhy4Gfm8q1f2sHGeN55ZTUZrazBFL8aXjXBwMBncpnlZ9d4mfvhOIFXBrFFBe
8lehS+K6AWLdt1h+VJkABg6mzjTDu60hVWlKL7F7nKtG3Ph7J9Z/bMPn573a9C6erCWtiBsm7m4L
4Hyrg29ESNl6MV8gvC6P8Xq4dJoUYs3oqO6g8eceYOANdu/WySaSaZe0o62ZHmB6BxvsMDZvpXg/
2q5vMdWKedCRTlcLwV9gbLSVe6c7pLBKGRWFfFmEKGe9Iy11WdexLKpmARhnLBXx12x2THR/mLVc
QNXvh4KyRZh9HrzzRHosdRe91g4rOUwIRjjMcHX4K9laChXIVjxXUR8tWy2GB2OLeqVH952YflOA
oWTbYu/CdPqZttY+oRFmk53LZHpmJEGmcPXp7k4h6udZNCAs7sOWD9z78O8swZOpG/Ay5w88/EJ5
+OykN/iCE9l69F1WkhNPfQi6u0gmMfpKheomjK9G6WnCssGkoosgTZZPGhzMyxcn3QPhDQKa9Nz6
g5vV2NLrcsqyVbbRWs9vjH2eCCbLJI7m71rdkUqD+3ANcW+YfcuAfcSd9w1f7Ju1W0oLUrxd1q4x
myVkEoQBWIJ/riIYLAxBdJk/VJO/YjKMAyVXn+IBxtF2eI27mfF5sUUE5BEQ4BjGV1Lx/O2kQm/f
eFDvjvJNH4cCvl+ATNa8hKb54I0b0z8Tu2QL0yWo5cwQ5zchYhUVviiFER515RI8yse+Rx4Stsdp
mCo9wrLXVDhVbTLd3TVmjY/zS1MfkFf8J6SrjrXjVrbvM5PvMdMkJVzMYjgUPs0VgofqdVmuOclg
Y+6l6sQUqZ+U0M91fIjFo2WWg+XczNy+LK7jRcdk4TesWgmF6v5tNFKwvolX3VRXhe0YrzfSmqTX
078P5zzam8dhnn5diV0C3OPtHhMVAungKX6YklgjfdWqhMk/gB5x7RJ/CC6f6nwWn/0aenJwqJMq
G+Z6H37XZz9IJeckIKc0GFByE25yhBVmkDxR7oO8fgnqhOlwb3QstFdI3yopSMvBvpvfzNGcNhjL
haBGBU0OYNUEkoLcDDuFzUnkIfGb44N6u3jRY/5jb9L1qkMAl15catnJDhafJ+OI9/7iIfqJO5jd
ScIz/lmlUpfRRvYvG8oAOSLCsFQ0RsIVkxIA+NaA57BzHtei5i0JVTGkbqSt9h7PgYUNstlJ1Uu0
hNUwTDH+p3MdB0Qvz2KqqwO0YJRlTCFFjxxxGVBmowdiPaLuItrjTIT8gBTmiXf1dpVv0P9lbQvz
MTmhfeuqPtA8zT2XakfC1/3hvl32hYU1xdS6jF3zwofEyVCiR/MV2kUve+8fR2/EQha9uZUVbNV4
hh0DPYq50siY6xRoF3xC8Yd2xzFs3KYyHgs4m0E6oPOfVxpBu6NLBDPl80hogZBedsufyok0mYei
ZaPv2sDGD3ZblT5Ca7fQGo0VY7hdkmurBXa2Lgodqwv9oZ6QsHBD7pzOhMNBpRT8awL4a7uqlxUo
4gARe4jjkAeJpxuxJKag2iUDQKjHqr8PV+ZhaiNuzGMU44RP9Eyzm53TJsHmPvtjhpShBLvXEpMr
KpP8PBpVOLnHrV0bATgMCwNCZrYhcM2tHBw7wMZmzufj6jGx2RfL8uygkh4p44ZT1iWw9PaL1vSW
Fojhv67XV9Zw7Fx4D1h2653UobgHQYdR1Lnq8/D0y6F2iL4w3PywIdMlynKtzQ3gMQU06Od0vo7y
JMx3nSx+NaZ+0FPFQwBFjJkxVKPMY6lEdPRHMz4aWAUanh5zcbH7XEiVFEWqjslZSCD7FmNoGxY2
m+H2U5p9QF0fyTZHeJCTqbwuhJLOsXS2I0PA5l2LUD6S3/3j3aiZs334zEX3D7AoMNEewCKPwz+/
fjztduyWNlfru9FjkpINSzAQzxvhyrdf8R/mxzjZ4/Ki29MippITpFeQjqDrzrZwV3BjrcpQ1DvE
A+Ry+HvQbw3KS1/A9agYZ3Oh+GZ193USkWcDA9F1kI24bSLKnAHjmnw5814TZLg5ZEfP2FdSHoqc
dwvpXXBk94qT4RPlHdxCA/th/vcWXW9P8HB6Y3uBveKPIbC0m9sBvyz/GPzuh65wmydS7aNY6E8r
ceWjE/UOErABcaiH0DtNst/BgxJRkvbt8uQc/Z3PzMZl9jwWEmR8LNgxtn3bsnDhTVymp6ULr9IE
+eYry2ZwsocWmKLFR3VvYmaIy9VH6DxszypoUUsJeiPS20xvVqfGglmpI3BTaTOb7M76rmNsMIBE
BUerZicQZNTSluo4BKUH77qYjR7nj+R6qvC/3Js+xndHyKTmCtQ59B9fO2URXIwsJiwgWPYlZvSd
tciy1uuejDSnC6cZz0rx9tnPCXzcrLCLQ1Rc8syurxeixtd0zTlmDF5h1V4b0HX6w6bgZEpVS6of
ztZ8p4AXchkKXfm59fCf/4sQNGdtD9Wpnks+e/yHdNkMkSK0ajPOIKYOK6DwaCO6OYh7HfRtsgUG
L3VcYFhmFfGSyMHZZI775mYnmENxZodVd42keUNhcZRtyWtsZj+yaJBmbA+THWZyjUb3E7zCEqRg
2RqpV01dMldtrVbHuDC/UPQlaVDC3QuWN8koNh42IP3AiPLa/DZJgIg7NCQ0ghl80Tk9/2qgYU9i
5KceKLGp3G3L+tuvU5ZjVOjG8lRyabFHOcthmpEDFqIMi+YmZt+YbzmaX5FbntJ6IyliVgXJMWUo
KuRywwZ0nzVnqknci+JWyrZxVN0nn7K0kisCwM9MLv1007rupsdVuuCaqHnFDtUGcNF8HZ6p1OVa
dq6JG5so5IcpExLRLChxSYmGIZM2PwcqpqlJ3UMwSMDxWk5Wfe0XC2iBs9suPMin0L/5iVG+0Jea
toxlJPgBYK4WBFP25zro8zVeSW7XreXximrgM3ZTmuHamacA4Y0i5mBYWCmUpn2v5BIpEd8ajTC7
VfVj2Zccm8LxCIpmvXD4Dr1RzHGgqoO20NCRfVvVh0Qjr8NnyPCN5277jEIYJ6iTyZRb+1r8hPY8
pybsFqJ6DegY0WM7fRBelnaQL3QMYLRZOzCK1Bio9OnMsxVF1fsHNepmVnrqrACH+H33DhEdq9RS
rhwJoUPJtCIx8W1PtLoB377nAp35cVY33HHQfVfM/ccvnFO3raA9vpZeymznrjN5l78a4IZWaOXz
lEaIzzi3ZGwntp8P4TdUO2cO7U+kZvPpy0AY5cddbgmJgaiOPVf9vIwaIKrYufC9oFpI+xM8L3VN
wTDtzNrUxFLrpLz5eqDpc8vLl2RoC3FuBtvA2DOuMWDUvvU7ZxfppiaajEcJLDabS4cxzXScggRj
FiNwPLMBJipxNv9e1K2L80Y+pBdSMCweq1R009v9zR6djY3VIMmZm1b9UVXFAcUWtK9rzhrV1rb3
aPDMV8sWQRVrvW+N1R2FeD5b4IBBRza9sSBieesNnpBoAheJqEFCDY4MlWlKRvpkK/JVqRqV6Tpv
teKW3q+Tj98Ra+JGBc4jfIbtd9b2KnFsRmr/T+9KB5pAdAdxEQEUQQp+dTlkdDUYGvunD/hVcmjQ
1NbJ2DWsgKzWarxqAoxOE0QbcbFu8k0GldExUkPNFCoIC8q4YGJzhcxpC28GO84pkT6EG467Jq32
PCdrDidc/TUMNeWKmE5qS8i7UxSyXvcEPJORYOefpMqzPb6ndAkpWdRXWjvwlR0yRRuWUV+tqQ5G
4D/bMSuA043//3a/Q5MkESO2JBkPwtlqqaeHWTnWhE5yIUwgmFbwMSDAxvaim5fGiK9H9HqjBrWv
Tt9bKt96MydBHF5MWiYAEIC/LPGarpRtTgrujnrSazUkwoSmiSKf6nxc/ae3ON4ODON2MROy8E8k
cEQMACG4lhJHXKDa1MgspEnpUtXo9UNYd6CZ/2uuWChwMJjT7UTlM/82IySl1b+s6aRLDYZCUEAW
x2OlYb8XkDO+kDJEbEfjLKLo+SsvSmfzX+Kp4cRBFmxatLJwCBeqC3+D4t0I+oWTmKflgPGMu9BN
95eEuZ2K3gp7zG6fDjm9n9hwUmenY3C2J/uEudicNv7oRSVqBT2KeDabOiFdc6WPYBipsppxi6W1
xIvvjOfGRAg9wuWu3u0kJ8+FFRYwRfQfRksGrfs7+wPjU6KvMLSeCKfwF6+/YNv9OPrh5rIACdNZ
RHaKlwCpCSBtGZ06Xwt/d/hD20Jxc7dqQkN0LIxqaauXfVPPJ347ct9LT5KyY7MN16yRk6qjcm42
z0BarrGtSoVnw4lW8X6Uak2+yCGrNaoJX38wS4Nf4CASs4/ZywxuvzBSbA0cFGmFGWTIQkP75ENr
Tsut3RTo8a0pfj9E03+XGRhkvy4sjBjCcPbwD63cFyrOP8I7rT3SWhmDtn5xi2vO/fBh+naqIwPb
E9ALavtyvJPrlTg1WOwtIX8OrLwiQLGlj5yWZ4MXNT6jPGhb6I27WSiVPLl6SpXzFCPQiUgcnuQT
8j+54y0o+qLAr3nMgKQf/F7YED1biXEezkolSxOhqh1di6+0d+pkLb4yb35nfTQs/Wzh/EE41F59
65X3Q6oqg2iHImVELBpKPLDfTBGWlNtlGiQblO0s3uKM2Ht6Y1XSnS7A4sHu8xDxIRytdtHeYXto
kjmggSEvCPrDO+lWarIpGaJFDNCHLWRdbxmoxla7j0kUOoMMbFo8vgby1A0D7tAlZhqGFmXpQXH5
S2fjRcE35Lfd20rhCf+KAk49Tcvdi841P/DRa+HjzY/MZLpX68u4Srz6d5Wnp+ykkXb8lWN1i6ir
Atj4b0rynUV7+XlRyAe8aDY8uGSZLAe/D9aoU9Fk3vLv2jtMZ1TzbmLCWloubpNkulBz5vppQRWe
fpp1Qr0wfxKQPgnnmoyyTieJJ0C/Iam3qEwZ3b913fb0zfytL9DBZwtaNOj1upq02AZJnvjq+Tpx
CGRq2rsL0FkeHuqqP3Mntht/B8CmTZwWZqJkrOy8NNCDHxA3Od4onQj3aQMDXVcO+u4xtqIJwsfI
PZnZ88MBArjHt+VZAjw+XjIVa1nCzuhzEizIPbRffQ1CAmuun+bUJI7QWwZ4e0bCLXseKVi0aFtR
wj7JcoTfXJ5HKVngqbO/c1FCaqLEGmM/U02QIeynM/t4goqwHj9TE7NheGQNeKSmLoLdWjyHg7A3
cigLLGdb52u5Q5VCv4qffDPnrUZaDpKNVc0JPQFAxELnd7we8udwSC561BGc1z3c7vfCmOyqXsIN
C+9Ajj0apxcX6eHfUDSHSFDqNihwqAIoKLfM0x5iIycp4Ol5X00jEHmhYuNBWVghrdiQGaVAtcG+
faKuRBEIDV+OJllNpAcxZJvKp1l+EJtnZ+mLByRVPTgYFS7KT243eslRcGEVipo/GrOsQcOUAobF
/2BWDSZHkIpbpxcGmbpTJvB8MtzgHKPYbZjUil20CtDpcf1LXE99VODG0jZE6lpIshu6CErwhA0M
UidoQSBY9iV2Y2eniTvhVxoa1IFiGS/wBtYX8JvKgoS7xZ2fXyIpveIEjmh6x+kGX4EhviCfuQa0
5huzLLYxa25HUukS4uzrFnle6yMsydCeOCdQDtpidX1rmD1B+smknBMVYcGT0kMQqQXg4dWpgMNj
tvtGuS4kR7q0rOJH3NFyWprd4/jrVlwex7ZNHGSAQYVhVHu9mvqBm+QGB3/wXsfEA3AVCroK+IAX
eTLHDbiOxbjGyRykijzrUyFNUWnJtfjfAz4OtF274e0DOy78VgiXEYrvqW3rKa74WS7+h/2ZM42p
siil/NFJoaBnr08PLiLroe+ygNfT2OLL6N7vfyQRhjdtK2Xo3sR8safUzVAzZZh722UTacWOIqyd
sK+Mvug5CRLy81bc5ZoMpSnt483h06tpIazqYNNYxU6D4a8Y5+uZZXLz0AbleA0+5ccPagtQcUU+
vM+umfNRdaYBaLuiZlU8DObAEghBdyNcBD2r3BNcP0YG3jD96ovceGYgwqsZeN7cG5DW/TbLLoWa
r01roLRxYe1EwN4ZZwHZnP/eV6GUEGW0vFPX8lMPO6G+jr/KCDxV0m1GC1vGs5PmNBnhHz6edogV
K9pXZyd8ThdfdC9zSue9eTZ+Hp0W9lfKX8X3KPP1UE9LFPpsvyz1tXo5jFBPTcvHtgxFOimbP1MY
yq0SGjDH0swet+JhFnt5M9paEtsqqoWaCjhzIshn/C82sPWWKyUWHyyIao3iYhtM9rPPjN7IQIpc
BCPy0MbosUFUHrB9SussFCPIPAVK+GlUbjN5FjFRwazuW/af2dmzyxGV1edlisk6t4r8bigxUL/R
Ce8v0BmKHrb11Gudu843DoNCty7wX9e3epstO15Yd2eu+dOhhzjsz6MHQswXfgN1jMX2aG7zcr5F
2AQZFnTnTM61kZTOysoyNBC2POA3U2PMKElJ7xP7UXNQaAIK88SDuQ6FWom4ufq/ELN1N7aBBpFe
UG6fQujsrAxOnvqq7aHPRem4aJ+oCr/NbusKwfhP6Jr5AW1CemuEyGO6s39jRNwat7qg8QO4L9VP
kxuhl99NVO+6nm4x+hFNR+aHXAD+rkUjXBj+VHIlDVjNxFMzjtceVWpV83vLxv/xe35cPlsb8tES
035Yg2KgRoy50A1vsPlv6Cn6L3JE9NT8Sb1K29UcU2gM+d8luE8PfM9cFIQFzzqi+sjpRl3TvrCF
nc08nDZarwwlFG3aTjifw3SRY7DhvG5AXzkL5AJPI5ym6KetlgvXrAjY53UP+ZODlbZoRPeqHnhs
KTqNZ7ZLFD2ePGNztvNWUJ73r32BfMMLd0fdIZsWfgwpagGfOCJiUPBNUwB+ks/1Qm7uoOWm3Qnw
JT1xgTEkERA2kpCTCvJDnRe6GyL+37JZNrxpl/AFrjrG2sJIf5Zpjsx4QCxRwFPcEn8fc/72PG3E
/KLVZvHO6nh2t8oC8knOcvChNvYasZH0sPH1BV0mdwrJ+EVnFYHa9MEBp7bA7b+R7O2YIsoHH60b
SgyZgJJdt7hgzB1mc3blWxRCQNoP8bJPVbkeZmLSO67f5/1dHL4w2/7usnAf8tPiHKOAMOcm9eTU
8tufmH8yzWBkah+n8cJLpF1J8QttMiRvc5wBmJ1taBDbGVcCIlfl2YtgG4qnX1g04xx3e/T1IAVc
54Fq2vsBgPKySe2brjJvKjp7rIxMTj+aTOQNNiHKtJ3oqmhx16y0G/hTVGQx4hy4C9Ie/TJyLtgJ
D6+1LXdJLlFV8ITC/GXTtRf4TFh1aRhIHPEbeJovgo8v3D/xtuy1AvAYuRRLdIsaBXTW8hmXdpl8
JAKq8d1+faABj7LEYr20VQVdSw+04P2PS4Zu9sosR1xE+Ck9V0l9LxeNt4p9HSu4sXFzTQuUU3NR
f0R6aboUqjKMZzzBl3vF+kvzRZ/p5tILJLguB+KVrL0+yBwS1f91I4S8XYwxzJG7e8kL0TIrY4iZ
my7lYrVq/tM+ikcZ4888N0p1hKGZnsYMfHEXuFse7iIexNCxODhglZGy0zjgdyF4k+1Eo36ugcfE
HYuUryHNu0PRKfz74wNAAis3mLCvY9Iq9wBDjNn9Ht3WNMQTHHpJ9TGcqVvFD8dHfV6q7AzMc2R2
r07kSM+PFAzDR5reQX9OECeCaz9f0rUrbpsJOVoXooTPPLG5CNQcEYMsOV0P+xYkeZuvUoX7Yuhv
8Dp5Zk4sXo1Mstgv6x0O97l2MS25JXCdx3AM3JzRyd26wKLG6pmpATKGw7+6BD0wehZuPdBdDRLJ
+h0H8amq8kNDGhuzh0sByk71bx++W51Q8gcnk9JmLArFoutit2ULICHiy9PaTe/LmREN78NZT9mM
RfHsNhzhD6LVJEdnOCJdktKMSAD9y2MfVEoHBcX7j+khwLOjlOc5ukHx1yCczb8YzzovFWe2/ZjV
dPMr9SLCxZ+8UyAhfxF5v8tidYVIPGXbBq6UEtMFKnnAM6nU9I12AjB/AQpLnDOB7au4aZCdGjkv
JG5tszCtY8hDUJ6dpRpZAepVeBtmQyHasqXOY0ojBl/fMdkxO2OnAT/tr3DsBwkcDyhxSmZ6irrZ
dckLo5eELmxb8xvXyWuH2+0U0VVQ1rPODqUPiy3TpG5BfYDxiu8q49lVmnGwzQ864FrQNRCknNZL
N5QXh49LlqIttuixUEJSQCSrgQ8P3mvsHB2eMmPZip/6XurKrs3pDN1+84Umk3GCFAydUzJ1u1vA
0L6478HXWLviYu7WvuMsbKEOghlPguow428bVpNHIYXCCY81z9U+F9W9fpjvHdW6ItU5Cig67Csm
GPJs4im3TDlhdGDmBGXzsh7ooT8Ec5f61O7f0kIF55aPoBbmk+90akgWmLr+Y1QoLQHMvaNlQZm9
hpu1ewyKdsiWzNjudd4bD/sV1eA/05YjJi5bO5xiMeEIuKjKXe+DT2zyaGKFaU3m8Yy9uXgBsspj
+T4QK44uQ2ETHfCwHOW1MXT3E3BjqW9zDgEzUFL0NJcHjKaRnXh32mbK5pAE1KR4M3PUuEFbJyA3
bKSZOE90LT53izGeR6wAdNFeUFXUN3IGLDzPCIS93uANjDQaHjAJHO6lfdCbqn42RkBvng+xW0JG
l+h+R+YzdRoeS5OtIv/Xoh126FUQK6ZhNczw7EWIsaLYAJC5jOLkPnyEkRmpophAyRCqRxraEpoe
hc//PajAmNYfX4Aod8Vox25QfbhzT4aKypHmgXkoTYkFMIHnLhR/GjZQiWjO9eNTXpUXmeVC/Dor
ls4e3giVgZCrNggNqhQK/b3VDahqUb5nEkRym2YkwM8CkTP2WS9/kpoce3RhNOoDVqvmfCZFQCbN
2buVR54YRCXqlWj5RCBmnt8RCUpj8GCbusdYjl9mx7rw/5Vnb3nXobSymLnywyyA3Qf5oKrWLKi1
LEsDO+o+xCQOGOwRnVw8n3yD+mydd0q3pdqPLVGtAJCUj2/S/QZVqjMyaex1G3mI6Hyh4Xmv33kv
9DkT3vhhAkqcstGh1BglhU/MbfSFbEtUb/L8tuNPq9ZkBiWiqSbWQQLR61E5nIAjeINpSVBP4Xre
vCs4PPDh56aNMWtjGIfkpW/OWnMC8kEA+IxRf/tE4fZIjdFqkay92LkmXrp5B10rHBkVVz1UdSKU
Zy7k1CvlJQYA59MZaMhp6/5K8BzEzYCAmQLNaqVuVvJv0utpzJfI9ogJAKHSFPGeYRK4ao1gu2Xo
7ZQnJNC1wrkoL7hvIuJsCnFFnFt7/ig1IhjWsNpwXIx1LfAMGIuQ1EnzwPtZAM0eII7NP/4PkSRH
0Rs/TlM5reLAsClJe6sCSvQA3qz3uW+DIMnZI4l4mxzIgCYJOyx7E5r1ot/OTH2NtjoVEUs7Q/8m
wJxUTIUenobRxZFWk7t2+3S7wOj+C/dQ+s3D2t7R9luIiI1snj9dqIb4AwWLYOhCWsh/mKcCHp89
hYQyahsJSG1WMGN8QYAKY3YNSudtE46+2MvZPR+ybVhoSv1iKf92JzCC0jgIrO5CHnHEoHFJhCRM
APMiTGFdAg0elMTP6nCROPHDQkGq198vJzHTfpeMG1s3TJqRUOOuCFqW24Gjd2r+nmIdOJbjmrAo
Rkg9y1ggwZjONlRhXcsaTpmFuS9rg+YFeZ5QNzuNEhY7faARRe5K4K2ajK0j8Bq6Zvhu7GojzmZK
ddpP5qkYqg0p10muGXRTxOM0Yb8TWWdMBFrbU9j/s8Q98doy1YylQZsLJdzIcwlGWOqNLb2FRJaw
VYMKZmmWvrNbx9JNcLYJZD0/BBe7io+p0lD/OWk6DAJuu1/BywtIAWBQ8K8RJunqJlNqIGZ/siZH
VAJa46EQZ4LOvBXOVR1JcTX+Y5IS2nJ0Qk1TklN0AOPh2BUchHANry0YipJY07dzbd183dKzq3Dy
3TQA1fd1VFb7DWJVB1ZMMOb7usuwYCph2+Eu9ZIox/PTRtfuaCvLIYpkyyPRNLnO1DijfB08nUJt
d76VkW7I+W8vC01lm90sLe1QB8wd/8SMpaomvS+aI7155+ypvhCihpZgR8wIBrHyl+alqaab3VRa
ei3dGJhPou/zNivxlJ/oO+hPfh7sBr3AAjpILc9vFEoozc1bbrmD2yqVbWgN8mLXiE5jl/QqPb4O
vNBwXqKQaCzDew6QhLov4N/nlbluD8U7mHNPil0HtM0RmaDIlttZPkOYceYObJfpVRwcL3YnXTsC
QxTOwnmNKUakhWVxvTjMZCLOPx5my7lY5tNikBemnjX9IjKV87Q8TDRqpJsaLKxneep4ohI/tvtD
YabN9mW6gmZ8e+mrXIy5zogzYu+y8m/4mgcpLspN2wpsmI5d6RFGDims25ahPsTw0tPGvvamY+93
8ywYeWKVnFFeWhjyyMv2eTZ+czY7B1MUQ9JfYeFFC2Mvulgbjyz2aIZUvg0D7oPpIa0aO1uHYJ75
wFufE1zPgPHC2/fZWcsb2vUTUOsz7vj4k0hC9VPAhvh6MsNz3mkzgToariss+VkQZ9w+90C3Ao36
uFWPFEp4qqZUW7VD4ZwubKB4uV5rm2AAWaeI27kpQTCcmP20wnHSGpC3XzhWW5P7/dVBEeZUojen
ncTexfYeCn9aYflGUhZcbp4JE/F2ojEq29wGHsKVEwrLk4QYOalZr/4IJhclz3imlaiHT3ScNAnx
nQjM20zMupSO93cB2w0Wb6by3x8109+tqjAUGNDFpnhxKuV1CCpPmukBosbMWgvErwf2Al24kb+E
1ljMtQWCjV1JSyFk+CVUglkbegsrhsGPJbDEx3/CzOeHAqrjKobTnw/kJog455FwFSrft40d1lew
P8rsh2TyGoKs8Q+1yys2OJq26DQmQw0GSseeAuHIqtWmGT4gjGd/1jHYt8EKN9DTQCfJNvg/dLpu
NWZ8r1nO50OGJxtVeFURqVPesSsDo+Uz1kcA/fKI4OglSrxkoyiaHF6lMar7qXW4zWQzfUnnQlh6
BPwkFD3XAJ4SF+OjQHuSx/cE/9VvZ/hPS/ZUFXtqmwl365V4vmFmyD+21ulEh513xSbf86C7kcIP
VrxaVi/sXy166lLh0D5I73i+acbK88MKBOcXwDVYpOBSBwJ3xrSNr1WhLmIyfag7SmmBwbSwc4P0
mn0P+EZhOioCvi/Xp5/hSqzkhhKXRrp5ffwaUl1M2xxdr3WkTPAvzKFWg3sC1DFNSudWnm4iylyn
DN0V8X+inbBZFtsI72Tq1Mf2MKLfd3fj4UcZ3fo4dvu/1FrLenhganrcNR/DMEnJUimninoG4L//
6d8gnkwv+PjQ+DghXB7cCAnFSqCmotmlYmMslu4AQY85FuZgLCU1jh/UuSrlVScSuYbEnaBAHXol
S9fiRZr4Wl1A0+LG8O5JRDvjORkJmj23qaLbbTAKGItbfk1Ok+lrK61TKZBDD5668BoKOghySIsj
uJuFcVWTgTlfLGgvR6evhf82a3xGAClQzSgS8kHDbFizmUaNmMf7Eh3USQfa6A7qbA79GG8nMNmv
baE9tOGwff4c0bS3Qq4SRw5BgM6wiqdH/ST8WuqmF0fzzRN3ewuufOGsdS8L9H7kqT8A4sSbBthm
Q64NQXwIRboUEtKijz/GjcNtnJOXKvftYefZnzeu3W9sPVNKaRYByhO7aZIIqLxEc9Jf0dsCswRd
7N4jooFwsRP9Bv2CRqXrp0QI869gkcg2AUsYugU7P0fGU4cusE8Brdd1HSiy+0/eJe+hBDMs1Y10
bPZKLIHb+VJ99f0T0L9JIYC+57mJBvISavwKPNKkN0/qZNIAgy+XKABvWyX3N4TLTCjlJP64MPIS
Ob2ECVHuA8IDvp40Z7bOywRrj24bS9KNxX+WjUId1J4DTP7CPQctKy8yshpq3D/g1dftFKKAQNvD
yxm4LSxTyYnUeYDme/n61TwF9GKOMB+svjBjEaBkFdXguTBAW64fz0OGUR0TYfgoVS/vqXOL1N3l
sQnTiz5bfBPHv9mxqfW6C34tW6aAZNFSpBo2pr212DXEzWT0zpY5bsKT3Fz93t1gvOezW6xAlDi6
khT0twWBaHrscPrZOAlM7pLmvymoQW+grjX9a3ZS+2fdIhL7Ukey2U1bo6bcGGBbp8i2wXKPhvOk
y7ozc1h0qyp7+gaiqCXTUtcPK+t8O7hp6wBN836osXOp9iHH5bKEs4LLx3JaZMXm6pRuyONecj8d
nj+eHtuv8N3/cAthVk9jQ6D0u/G27BhGWXXgsesGYSjs6M5J+QJr94epfs5477yeKTwtTWlAzAHT
NVS13aDzpiTQZF3kU3/8fzhe2H6N1m/fmOyXutUJDAZAiB2QC5owSEUdK0BBaX3Wm0tya3PO0RhH
u7GpDQtovXuOGKMueMjTd7vSacCN9Q6yr3eMAWOFjdOrRupepn/5uUp18ZY0npkcRHQxquBnfdJd
FE1NH6FpwpAw4+DrnrpFpR2LSbHumAw69KAkhjBwPIgNF0+ZQ40gD8xDsOtSLCzpWH3t6fjc4ftM
meyUpTdQDJswWzpFWJe4AMK+CvyFm3P5pxk7aieNmURYsL9BRbytZ5AeVMh9pgUAdart4kvDWLq2
XZd+woXITV7eqDXtb2fUjAUmCR8dB4HuRrrskdLFg+8oH1I/mwPgu6ndiaNkt7C9KAUrE8YNIByZ
g7dc5L0N146ZrQWTinUiIrn9fksuuNJLdSRIZv6cEZMAkdxgcKKnDdGrpwuB/bizeqmuJki48mPx
D4iStxDnuvsjsJ62DxkkoXjDFBp+ZbjLuiPWsHDZrQdXmJGYIJx6+LjSX/hNIgD+U+TaFnZpV1uP
BxKGd+jhas+boJxAj5ATT7Y4QVeuk/o/chGnXCNGnnCT0sfjNSITjmwhXcWQsaCFqD7kabCtqkUy
gAN45iIAmql1twnj0x3QLktQVnNdg4vdWtWUGLe/8FAYaSXCET2ldMTBTP8pdDY+uMJXxx1YRngn
IxoYmNOf91tfcJnBMrTkakYeqmqZGXkymLQ71BWY2HVGfQAxGXpYL0x9AmP7sO4c/AvZkWxWZKG7
3dxULt9hieokZhPg2IXun1NHbz9eMKGA0vHcRaqU4wk9rk7Mi2e3ClBRz31zl2O6MllzpXCEBfkg
0sWFkGcLKfg3UaAXzYY73xu+l/kSlL5DCvnv+H8PZYxdDPNVONhdF0NYlwI3ne1lVP87TUGRX7SI
RfvBAeq1HPQDrgq4FBHLlk5GgX2j0I/T2zQejuKcT8kIeY/TlVUqA+u45/LKmO9KFdyENMKv6qdw
54W7JnQozaSUd58/Kn8QiNAtPj75cE7R/FQqV1F/Oqd5xilUsW9Za6zymJkJ3/htWxOc/+5XjgXi
wRJwSyYgBsBsjUWm3t5i2E+EsK4LNPGy0AhEiXnC25m//LoN51UJ4f6J7Bexc/s6Jyl6xzmRbH1J
CYpPy4R4Ig0VhP33uiajApVtpd7tYGFLCchdslIQJQCTkH4Mn097rZfzw5i/DMPiRopEqBah6Wpy
kaYrXxKTTii5MDz1+TnWGvDwNhSrMMONjvnKJkVKb7EprnUwCtLa3dcumEjLvdR5AdNMtiVw+xHz
RSRudf4mRivApw/x5iQ5NtR8cW3OrvuGCe4sYqEPm7UESGC4iTyHCDcYXMI5zsgsY4cq9R76o/SO
YnutKryLmzRTw2S8vktAfN5/EqUsciVvGigFxJ7ltYOHImsFRwd8sTKYuznJfj4xSBpNTnjV3BGq
gD8jpI4vUkizX8De4WMEKhN+AH4sH5f14km27qoRE14H22NCeAR0eyZ4do9QtFvLkeGyHYhMnr20
TDbYHfBBkKfyw8bjaruNSOuIbNW1KycDDlWaT7KkXZzvv989IQBUWjVQKWwwTeb9jmRsaP2zlLqp
emIFKm+Y2pIhu+3l2igDKaEui7Nk6MWqh5C+1/5dCSu+e5d5DfFcttSxx4NngBppSNoUSrJVC7Ga
DCR2M2XT2MtjF16RJ21njDrl53qHb/0JjT7aQUpSrO6QikOKeIno7DZECcTQE6Xwbo7WX1qZe1If
KuZdDdMIb+HaE7eKe+rBi9CbnfiHw428Xl37WqDqYVTI3TPBgBiCGl69izj8mZJRyezTfdRdoUjP
SEt+VGsJnhk/LbJASvgomsMHISiVzV4GOxxQAiu9b68StBVYLErUv/0alSXc0YiS4apx0/8RPGHp
yd+DR+byjrZqI5xyWjMVCXj6HDHaCw7/C1gUxJtDhDfY5fFpC1VTblrwS8Dz0rqb2+5U4kr2/ewM
A+BfUt6Yu+e5ugmfvEr5MFeAHH7QaLIc3KP09QAzwe5j60i7fG+LJwMcZWPDO+7I8W630fvtjJTE
CH0CNy2eKWcnDZ6jI+vNlChtnOc9HyZTzqTWEcPCT0f+N5uK0OAmp2X4oI2iJ5V7lGgu875uS/lm
LwSCALnkZBy26BTeqZ7beSwPEz3p5+JM22GIZL2R57NNSCO8KZ1ap3lblbz6Rrkmt/8zb+BpnKNa
9jax5eoEvNQE4V01qmWKlMGbth0sqKYPeJHlPpVQoFVyowFGVEqhVKdcUL8ehawkDPSqH9uWuwPA
Xf/fWy4fbGGXFujxUCUVq7WWG7lV0ba5MJJ7t9doqetz7tqA1FGOqVoKGE+Hjuv8Auyx9qhRYd4a
VNQQIdgnT7oi4HqystXTpBXqSAFK9FqOEWcane2+1rRfTP7Kq//B5l1Hce6a/bZBrZ3tEcpyQ4MU
x199QUfwp7qU6Q22SSr8NDzUhVfClkv3+/98scR4lIoJuRAx3xQMDJutazd/VUARszOh9CedeJSf
dsduckPoBVle4XZwkO2Gr9UK1I9GjFl/NOm5aywH+eiesFs6yTD5ZtO9Vu60nzem/d36C9hIHQUG
XEjvisaKN2S0OxEhXxdMVr5mCSeJHbcxx0TMB0pQ2LZw6MSmROJW6F6q5NAEgQDp4VZ0UffICzqi
PUkUq6L5JQ8kJb2f/Y40IIOF0lcMNqaIMQWoPYFer12/Fny8ruxhMVZBZN3d4xzpAe0voRrqaqBn
oku8DDChmUehqbn66ZhkKvWq6VxMXmMPvcL99NGs60lnLwl+1zAqCM8m5i0cEsKWmJL/BuLW6ZyR
guuf/F51CwVOEgthsNjla/6wUGvO5rDifRvSyxSmWO0CTYRIKtB/cOWBdR6m9PvajleMnJGsVtiv
+NTIq4V33FrJ6OcJhlPOuq4yml/dKvPalMaV2ApXdsnO9jVKNxNepCumVurhnV+scGdD5YI9esTG
A9KJkLu+am2N3lo9kUWutAdYadxjBRgKzAWHUGoTqhGeOTXmJPhFjh36irpw38UfI3XkdD1pbGdx
VIkH5zWnu21a61KbODBilvH7qTEDYsgptPVC9Ver57Y4JNqlZ7vEwWPhJga09oBDSlL8FfCU2n8D
KEPOo/GNpwvjviWURi2Tn4YVuyaV5yZUqdMQk9DYZBxFObuBULJm15B0n7MDBtlBM4XENdoi4Y0/
dU4fSe+wlC+QJUXoxTfkASm3t3muiVL5vYr0a4oHT9Ej0Vy5v9aR46n9ajfNi1UeLL+CRY7Cci3p
bZs5pAdrKIVb+LjJDri1z0sHU8tRBc8N3Dmo96nGRsOSoDESpGd0XNugYaqF78lfHq30xIG1ONhO
/woEIScQY4SHJEPNHrS0ok9rQDfQZevQMMj7RhSEn5hgLBjNshPV3vfBe/plJQYdFaiGfu8lSSUq
FveH3MHtqbMzW6jsmwif6BH0eMZwrwZs5jw9Xa11OGjdSPedOW1k/7s0fFuID0pl1Go57nYRagRt
BtNwqxdkdw/ROA1VWJ3kHj6eKEtaICDXDIs3kGqfwmW87B1hp5knjJV7R3X/2+Mfow9hl3/+YjUh
qoEARby78QFjcfXonc1jKXWcrUQvVpZtwXMfdGKAgWfR52TZKtFvUdONA6ooxxzz2ZBkrVM6wcOj
YCbHPX/HYhErmcEMK9jw3O1cX7UVD63yyrt0vxCvMkbN54mww0+WBk0EjpF/NOT3tgWkeKVM+TVx
iOc3ijtnQj9mLukH5BSiDW6bcz40rlJq/2K0rJ1+iog9XIMRml7JY9jBiOmna7pH14sqaZF5q6oM
oz8eu8sVdZZTyEqXy1BUJVpyzWC64HwGHJJpmi3cl8fzPZNhm4QtfiEjKOBhAWjqSLeKg9Im6DVj
Jv9nAUm2eE2NpzabKZZ23Mh5gUR7wmbC8B0rBwDXW6h/HP458lTHhC7PUFHI/UZniuW2+sAoTqoS
V9tnk00jZ8LoowhMAGTo2Qg28CO/N00RtN2gyJK7yYOnUxkOVDSbuL6IPcx8B9EICvUnpQb4pcq4
anFznzkTCaERPyvQbxyjcATGticULrLWCzbPtQSQzC+aJ064+da9xK+1AMzpIcLxHvIsq/JV6Z6+
FnIfBqtKBLdgC1aS2+IHShQoEepE92o/VWjfeKrfTRsdTDe3uFv/8DVD5bIwqZcjwtace1De6rXN
COUqYSnU1okTy5YQrOzyXEeCa68X5Er55kWwMGZfoeTrbBxPlA5lZH+Y/9mVV6d4hhelhL3YTans
+eJqwbMlx/ioFJ8HVMSy0lusiOmHMK5s62vbxPMvsC4WcfI7zRVjbjlDqMsZXENo6Iw7yE7GAjVy
PvD8m3zJdFw6STmWzMz8SY548JB1LSp5T3yfeIV4EsXZb66mZut/J9pYRJl1Q3hIUnxAM8FjtAQa
AzBz6Q/SLGrjO3PVVPd3IKB+0eaOLmwr2bVfJ21JJBMf3xQAVZUK/Nr+/dHZvi3jX3qFAq6cq9ZL
NFw4/yn7V9LJZ0U3ATyOdnY9tOxs3m7/WSxVaM3cipi4dg7a4zSDx1+CqPmsZuGYDrqALxTsFihc
y/eAomSfcIEquER5YwA0rF1fTxp+nb3YbgsQEcAmYHb4cIzE3QDAmj8o5GJA/T9WOPg4tpcITAbe
9R/2l8DAC6T7jS1nRki342rPJkrTca6+43jtOq9f0qscudo19HSWXc/8tTRVe2UBQNa365haJbXd
vPD1G12ERjEgr5ugQxkSiVw9cgGBQJUils5ZNpBY47zF9+dqM48qp7aMVmjNd91LLBJmZD0ZyvJb
HVKLcvqe5wGvPkxi9YlFb5epi3IVBhA94Lwalupr1aegbScsPMpUPJ9Xqr+49gxtpgOYc6VPXA6t
LY485fPWmY/pCFpfqSKKsDURMkfKo237T04bFyYHdZ+RDUdMBigwnACjrtWog2/Zm8fDd7+Wbnqd
eR0LqSUKzqzf6eMDtlVyNL0cRmLoTC3XaBfiqduoSGtOk6yJrhwv7uhd3rNulU0Ved0o3DWkYcKr
F6ENAwDKBlh7Cf3Gshnqb+4FUazRsXDWCBTKSDwhpeKLJY9t4WxyKqLSNykuQjvg9HJ87mTR9TqE
9M7r9PCpnPchd1SLGzKJcHl470v/goGCwG+cP839xP/m62WshbdxiJxs3tTb4erlYmqm7XzcE4Bb
SqjRXWEhvu+j62vSGvlHVlhpFWQu+gK7+9wPR3CXw49cUVNeJ+3yFbD4NJf1DHu/JcB781G4XJsc
NUQQhX3UkgSRQA/Z/qPK2GqWBhpEcELv0Ewtc36VUAt9DxeAO8S+6xjGcjhGoQ0PFxIWLzolJM4/
6E0Av6f7OQJgpXmzgNEdx0O7Jjlpn5LLk825dvvK5YKhmZns1ztfYBRiW936wn+octzDA44oW4yf
fV9d6xXy6yKRuPE1YKrw7m8VqvccxE6y6/tEUS2mLiagGHaTftrhy2neluwUpINF4w0d/vuCwPg+
zHgABunQiGIiq7QQaNOGHblttxXnxI2Nk+l268/snNkK/VVobrwDqfVnow4AdYyWBSVpfm3hIjAF
AZM17ZDoZGhPLYFSSfHEA+FD4kxjHa+sDoxaMFvgMh7aRDZVEwWFnXKb9x0KW3rx+oZq0YZU682F
8C64d9/ba0WJf/tpOsHt77pBiyOMQLjt4khYIWJyxK/0mktZ32/WHAdtuG/I0i5qilhS2F1horFZ
CBl/GkDX4xtdExOfW73tbMiKhwOcebHqy0L24fENgn6J2/gzKH+1/EZuXoe8KdipKVcnOwx8fhg6
/PLWJEcblU6qTr4MHQ7OlhrxefL13KtS0OWI578lbwmGqsameCQdckPVYiPQ5BBgJapiPPVr5eOP
8oJ+kebz3YiZBckVBXUADLyWyQoK//zZ7mjijUror7hrfZErnmJP/0xLzE/6benrWoNJEz92I7v6
JyvovgFYbrc1Z0eDen7lj0SyZ3tNlA80D7mLRyY6sZYHzien/vrI0B3PRt5vNysUVyDq+HzXy8xs
tBEIcVNJ1O2rP51x5DDmrdwHCsiEp41y5AM/zVIAVQ8cMrWZ2MBxtx+BlhAPR+yYcdDkkuRenTRX
33klsrpB79vUMBI+OiRXXNVyvMbjQq04qio8JxeTXos3rx7dkbvcjBToP+9wX/il6DV2TDHJSOje
9zhbOjeZdrqmtRXjmH6bR/PLvqcmWMv7YyAV0BrozHWmM+1rzAxCG59uEf+5G3yrRiH1MTy4GYDG
jaqjl68Q2JKwtZ3DaYGO1oET60PDxykVBWzcYLHqRx7SyhQU4zvM7eTOhQuqwpyzRhaqBHnsrY18
uw0vpz1CqoSF7rVOgRhJRVNkEPijKnNGUezSvC40zh3b7ZDa/ExPxedgBxdBe2VpPsYL6rQa6N9l
kZLIC72V7HF+zrfxnW+sG78EBTYhsessE5dBWxZ+fhEgGJlNg13IoUFKa0r/s4BkH1gOPzsiIYTR
hrqgOyh7WsEpeoMYNa3k5alZcXpV/Zf//mXs5ZNOo/O74cQGvAtasYu8lm055+svKaWVDMba8bcb
q58WSW4N8HdLKXIHppc8om+/9MsXXeICRRWMgHUU0ZqyPj34eKMWmsvDQq6her7hNivkUGVfDMqg
mcJjLmq8/WZJtlZp5ykIzuU9aUOhCs2BbtYsIhxc+VzCsb4RIbtU0Ch4wFv9KocB8+iuOdLhe7i+
PHYxDy29ep9WA7042oZavO5qB8K64ojVZe9lmyLj0Tqe6quC6KVC6uNrharlmW5D25qbmnr1CjWI
BsoDzLjTgMfVi+GiAqC2TWFvKwXQg3dEZWwuEbBHDB6Fus4uzXCmGX6YTFlvhzCdiEEgS1f6fAmj
F5CCtTKlWeHpLoTpewIUoJtZq37QQ9VnWcJ0BtuLzK967h4L19aCUz98FwdhVvIcD9Cao3c6kuZv
rHPjo3jTtwSyXnRyzlKc8Lwk+2XWvtsY0CCOP2gpJBzHNTXOfwlWnUAeQT/6mrHTJlpDws7qBEuU
BdHYMvCpUbgNoGLAcOhWxWxDBnOGhAkwOyVqAB/Fbo2SUSFg/AQ4VtsQhCcupk1iGusVpTSiOQ94
YHeP1heN4to0t0oJIOUsmPosdlV4UP5DodovGUJzu3OsWJwLQhRpWUZJUT5kHNfxy6XfiDGVEY0c
TdQo1fD+FAfGbGQw8yHDnmBg48sUrdeRH7NoPOhvcU6PZVoGfWYfcdFZmYAelTQ5+XV6EiDTqIbE
ubXNvuVO9f11I9+U+mevj3kCrgmGdetEodVYjLvrLTv6XhdJgAviMQYgURTnDaYzrpq1PvePbBB7
gsMt5xUd62F96IhHI1Ya0QijvbDrdptgGX+0iwMkvjD6qMYKgAoYRaEHblq0jb98gJIFfr0cH8Q9
/tKbS/4SiBEYjS9HiG/Rx0EcZzYFeENDR2JQlRLIbA1ne+z8kfbuvgg28cGCSPgv2phwtzellht6
UiFaJ1mQS29hSZrrxcptyhwoULCL7pR1sJbQ4WpIlPn7efgjKMDO6fnsjxve6bZHrpHmiIdAA+Wy
XSSTZ+Hu2wCyBZzAlNe+/0gko1XnOp/y3ZoYHtnQH+tHZ8KrOo5J//9hbBh7CuVadLC622l/0MPL
oIKPrVFQ/OIKQoYLOhtNAO3r/H6ztY54GODUOdAQ6ryX6CClMtXkvfML/eiTCDZK+TKiUyRVF2Ft
+DSo6YxbzKJJVE7QB+2cNaaHhXsiEqGy4L9IgB2YZ5xUq7nF+jXwo82y74Rj3ddNCg7vDkZgw0xo
L+IDNDZF+Rvdxe9q5YpSgwbq7Ny/2/T4+dlTe+N6kZLil8Tv3AOUPW7RHVrj/Hv/4zW8gWgeOpgC
+sYGDJcll7OpWiI6wt0KZWjGWNYelmqSj5+QkTEuIuNizxts5tsFvkk+cHpNb+FhrZW5I7gasVuB
XRphK7lP8YQzeT6hmmzEvJZhm8wnk1vCjqitkV8DlYD5ug5PChjuAaW40/ByJ2xdU6MmlYDvbZ1s
tRAzny0Wkck1G/Oc5ZArMD8jrIdmjC+RC6kk2JOPNGI5BoUpDXdz3902KTMyYxeLIs6p/DJ2cipp
RbGl6mOReKA/EixjQMZb6q2kREv8PV2K8pJB8/x0EMoH+TIJJXs5siSGPUe/LWJDZE2j6gjYUQR+
v3EY9fG8WL3gRBj35RmBfJA3KAJEE1a9ou2jr+Z0BCoTbgVMl0lkR3YULZqrA0mBNTJl1mLo/rZk
Ee+4yCdrOi5kbEdaf/ZWXQjEVuWfjFLL4e5Mknk4xZIBVsHuzmEGcjmXxmO4NO4gQAvSXSMr7zPb
eAFYxabV4jvPPw1eqDY9Nc8rpU6UxbyIcsboPL/Q/zQsrk5gYNJqpMstxG5V6CYYTI7A1JokOjLp
kmwaIa6drUTevUtP5UQYnYVToc2E+c7wgOy5lbZ4qYKT9e7ltuBsh4Oo2bCQ9SIYRQVSDOmbU3H1
B+20OEb+2A84EPrlhkpmr1ll8VanJ6k6cT2DSkZVeVUSKtmw1otfj7pdUY0nqmN1Y79XJ9uiQmKd
JnURvVwOxwpzddH4PlRXbj2RakxhuMYfdJsCzWnSJ4mPJWucot35cnLfI4aaIa1ceojzGDPCuCRi
NWP52bxCJn+Dx8ZT/UzvEByqw6gVDwxQP7XnbpW4HIwyW2LetQWiw7DtBbmp34QaVsxZY061Xa4F
AF0g6Ay/SbdZKjri1tTd6cSYObayaN8kOOBESf8wvWFgXfvchJpUEFDIpUwqjK9mtntrqbhnUR0G
HLlxEoTtg7a9j8GqbZc85KLJ1tZwbUJXIlDZE7lM7sO1j/LHbC1wkLy5LK2Qs12q+R1K7Bga4Acp
upjXPAsxP/fGfIKPNFr+HECc+qOwb+weGNd4M3u8xUPSqIKJU7ofXhAA9gj7/Tg0w0HzIOeiGlEk
+Y38/0ZJpxjT3b6BUsL0/FjS8OwhpTVhWO+Qa5NWzJ6VxeksbWOu4OL+oBexLOQzfrszmOGxV/zj
GScrLcDYksauVa3NN3z7fzL2IzzBWTn4vE+9vLxuQys6pZDItRzhHCzkHg4jfvlPnGrr0R7JBcLZ
Nunr/oypUW6ON95mSrNK5xX2BpAEcMQFTPW28d94uoCUn5qjWAPOTZQUyKke7c8bJmV1IektBeno
CtQCg/9qm3ffUnHrKQzMNtcfnV7a747p3k/PwNVIyU0WHges4qC8GSuyr7yGq2rL+9muqigtdlo2
mT/w8K6OgDiVF7eU2Cz8jA9TgMWnZQWHx4eUW15GRztu2jv7MRLzs+Fp/vWGRxN2JdEH3ePwwI3v
84WOp1zOt8I4ThitAQ1TKLnrMRm560YvFQ4tDkQWRRei36tUJJVFIw/J7oh3M283V6qMCCBj/A1S
2ma1HeL3tFMvGbgfo2X0ITV6Wwgp6yph1bY69vfAIlAs5uSSn3X+1XUxJ8rNkeMiGYR4alcgykDB
kG1pFLPA6jtrYm2QHPTTH69Z+Cf1Q6MwGTitBOQsuBiWlVI/bFPryffX+jurSgYY+MBGaySspMXn
yBtXOs32XnVbVRu3ia0jCXmhmJuUbmqzAIHMS1luWQ8Uu2Jm7xpPH6KrAO2m1owXh1TOxfvT611m
ATrl20NtB5DgYTr6SfLH9zszZAVhsmzOeuvJCsl8/sN9MFx7xEky05Y0iPTALxwsvRt30nL0z1G+
71xIVRgWpJy94GDU2XVh+1bpNAZYaxgrBLXOGWw9VCd4vfAGmXhI203kTvgJDn1L2shjQsR9Uo2R
dfX0xo/yfYWyL3PvCOOmsDZnBhXY4N+ShLvrOJ1R4udwoL2btiX1NMPImwNDHqz0P+3OdBYmM6PL
sFm9qhBfKFgCWH+xfrvB4sCTWb42YYCVZD6dixJx8eOIlWJU2nwtDLIJ1tIpEls0NP/nNAO2/FI4
zHt9ecJbeSaQIzN8iCC0u5VqfEzGCHO3MftUMnXPwzGWnR4CbNz6sWITEzKWRy1rCgVwdfCZOMsS
uj+ZVR47A9Ne0WevY73vmvPMHItLRnwBqPJa31V2M3L/wBhu2Ql0iGNZ0gztVuELYjBZtKFvePqQ
DV/dTSosbhKvpT6PEsJ62dVa1KPIjnmLPzqqYmdons78xJkp8quUBRQi2DA6ZtLK/ZomT9yKef6K
NxH2/IBjIJsU8w/W/snLDu/Sn4PiA5u9FF2aNAjYkPso/ar41infM9fqRVE6LnIycF7/dWJBPpVH
68z2t9rqVI4qxOzhg6G/yUlSQnXSV0/pDfsNGRECbpvFYZjDacmfR3hPJlU8ncTV06tElMhVQppc
2cemVbzGgwfk/CSvUiKQrMvuasoTNtSeqkIAT/JfyvRaG7er/qoq+ENPNTshTnRrzIjghofU6QIJ
sgFzzJpwh7ygQKyZ3ChzRPFC82xM9ciFzGPDu5i1uFAcrwAW7U6SBY4DFIXv5xaH+YiraLRgnOY1
Q88lhWlLQy33fjuwch2ILaSYLWxebbxUy1FDO9Gka04udahZyP3Mo+1DZqMrCfj+tIjZtIpojdI2
wdPn1hFlwe6VmIrFApdfxds4RbmNQDFju1zaQ4t2M1fcTLoNjfBzSHUx3401NCrGm74CjMCKDy3c
cpWllxiHL3uBf1b3oyChloJZjvdpKetpQts3Ln5kUTWaid9gBWTsbkv2HUwR0tKWf7bFXftO3QpV
71Q2gR9mDUN9DmSRWvT5HPPPZlfYP6cM9TB291p0fsr/Y2jvGnG2QCqzKP3QmSxXQLTzoEbpyK1O
aNW/EL3zMBGypSiv5ofkzJBzzmZ4YxqF3/SsWaO3f8BThwhFNR2TS+rvsLI5bg/Bs0AlZHITJLMh
pVwg0HJbF3YtIfuHA88nxOvCdNb6+TgIz6YbB2uGkScSGaCKBtHcp9zR1AJpjPALwRocu4LBpexM
6kVllnxFxc7HoydDCMXEPWoAZldShwU5rLvJN7IQ5/3W2nB/Ymv7DHmP0vNXSSdrH0HRuAEDL5qo
oSZZDgQRUBcyYDr22nmQ8GfBq6gttS87YN4ZSG2ZyeFXclnzqbh4MdU3u8ehL5cn6irRueQMLP3j
Y+d0WL3ZmE+pvaNBDo9zVIDiNhJNchFHNRcxdi4vV9kAfdNVzE+hNW7g88swiKNBKqtC/9wKWOFD
N1CIspjMEt5SFLjdjlT8xQ5HPH0mYlvpbvSuFPAm+Vz1c1OoflO9+bZIq3OC8MuKC/phYq1itR7n
aAp38/v7cjPLma1fBB1Yh07hlknsPzw+OUMGLCtlSxK2aC4bLVYXl5fI39phlGvBLd+cu3yx+iTR
0Vtr6YlDzvmBcZmN+iNXN3Iu027bDNSeNFwQoUo9tyGF3yjCQXdsbDtgPW16Paf+rQNeTr1//dHG
iDUeOKUtSJ4grFdBTLA0tQ/Fl6C9Wl4l1Oir+qaV1++YSswHoKBwkkdWGXcTX+r3DAvQ/BMH5KJe
U/Da7AtqRTV6YBAZsDopumTzneR3R5dFaWFoBMbJwOxKLlGk2zazV3DUKa9ozSH4A58fRWNrCoRU
9IBIC1bd/rKdlzPp7DHZfq0YfCjfV+PW1Wv/P7LBqhKBHu58vc2lwRTVXBFISHAjSokjOGyP3GbL
EcwSiFElgN9Dib2WlpE43PPNae+b+IrRusSTfGEg5jUgzBOah63T0T9kVW7W0YykxM784j5FURW+
DssVYcaCprzuOjQH/+pXYZOnSACMnC0MzRzaAW0aCmFxvrDHV7O2/rmBhMZQWVVJYyVRxFykJdWt
NXg8UgeM8cZjb4fJzQmfb5CXfghOD3F+QZ+oETQusJA9Sifklz1SWZqY87kEcq1QaL7Ne74UIHtO
FbDGskuvALjvbOcp2ek1b0lQ7pfsMxj+LSCl/Ox52EnGywB+ZbqV5tLwGcD875HTJ8ADi6Rt2q+s
QmRQTCW9ikVUEurxLt/opYzwiIA4yi5BxL0zq11fXAEm9dne9OxtqNYk6h2WeLsiThyOjWk1M4Sa
aF8vHy8zfd3UdKUZfb/qMswM7fyeBJ9HAO3BGu3gh8vbNGaiY320Qi/A5RwvlXqkY9wU6wOQDWKe
FeOVzRqNuLII+O5w/9xKPd1OBy2BOZAVfLeVbGQ38JxQEgOzxI7CxozUZvm4itETDA+32a3/LA1F
hpWyu8E9AjZbrNeszEfMa6/Q+y1XreI7CwMkBz7sVZX5noE6cWqLe8Q+dVjwlIUIzRkwCNL/mP0J
iKs0C6mBp1ju2xpK0QoentrdkD38LHQ/HhyrESBL3jVcgd2Zr2mQdK4K/qlCf40JDWnwvadWoSUT
MjGJjwYeoYKx33JxrqePkW/9wFCKbsFDgr9JGehImSP1YYzu4KxhWUSbYZmv0J5H0xJgJmMsufuO
lEpdXSc0CY6kUwMySdWmNNzBSDadfykDl+ffIIuc3B2awPq++Qpkc0P9I4/e0HkXN3oy2DSRan8r
NiRFWWpACCmnVtbySFxfgyOeEZdKoFTq6xPxW4V8XCpvA3cDqg55weIrSrCUuZFQ/KlWAL9gjg5z
ubh+H+leXiWeTTdXpAvsjS5Jk+/+xAfqpKRCCSjc5MUg9YacpYTGmSOKg2G/p6HcRm4Yi7kqBEvU
JMFyKsOITrZQD2dulYf3j/+W4r3iLDNgwk81ylTaHSQCw3zsbUkS5R7dekkRgqrVikSQsOkyrx3d
Ku4fVXdFhR36ihJsvvctQc0tknpwhk+bImCe+S3h0CTTCX1nFF9lOAuzPdlgstH3HszXjNu6a6CM
1Z4jE0wDuXymM70dmZh9ZO5D9fdZ7orodxhv0vBfD/yLmA2yjFwTnSSN1uO3Y3q73zPS/KryWqYD
bwDQvqTtco7N714tDA9s0474pxXQL/rVU55cK9/euD59LActQ+XRiaaLLY1IVVEUqH6T/IZUf+nE
skUl4i71u0a4jQYPAq3ntlaGNYGJptGewn38X+AjY6KhAXBnR7uOBoxlAGgRI3UVoh/CeWk6UvZP
GYRp3qUiRNcXFk8YDj/XiiRirviD5lGTcND/Vp4iJNkrKniEf+nc7yNViVxq1KjY/8jPTGH7K4iZ
t2qWYEmsEg+TUW8SOpM7wdC69yZpDrLAvQrN+VxGgyQ50qrK4DLqX0u6IgNGmsCX365KuJTYr+92
tMtRVRxruIbqX2AlKj+txsitEOZrgorMyUY9c9vMPXw3FLO2HIaveKsw6CfM6HkA9zfaqjebDiQm
vWBVdLCY8geTQxPS1LwRwykrdz/fMRBJcsmFuN/RjaJQmcTaQwMmqtX4+uSAMoLjGiKGlXcUjXLE
Q63gAhl9CZJjVUY3Ybi816Rt1zHh4pselbY+xTVVVVJqJJaCSmGq8mRhmJ8MdlOntMI0URxAk/4W
OaY+99FgBNa7PF6sINmQW6PNddz9VcwZlm9gUUbcsL2KBc8gG42PvI7cEUPOjEyUbKkrUfjDH42v
Jo5wpRN2tyfuHCvBiqMGRjwVLOLczK8tuhLKEGppjgyqOUMnL8o7okAXKgPp2B+ccpj7sP0xB7lP
PHVTXDHFpUCTMkSZuVrBxnxTYwRnJ8DBbZucx+kEaldjEG4l8TIoVckk+X3sJhaOOce7ho+xdGqb
gT9MyhOCVYyyCMh10I3p6Tj3dWiWcO4LCmFznhrhgL69xNU5CcVmoBVipiIPTHnT5yagGjvbnTJj
RWSDJyPV6F1hIFqjUutIqBz9YhXEe4bkKiLyPGhi3W+1KVaQA9UQBffoqqJiBu7AYGocTT2lNMIS
6e9zgtdFCSApj/F2+oy1C0x9nxOEvZv5Wj8fUSb0iSLVz+/4W6BsRavpxJR1R9Gb5F4yii9ma6hx
ycBDnGtNyCDtZTTyD2T/7vnJo7T/PZcirPMjDcXycx+IcS1+CwF0xDrH1olzJrT5yDhSBYaFetkn
xLlQPq2Rpm6UA/UKwFbNPJi1+Kr//cLdKVbUjv9ofReey8tOKMVvOCkl8VXQLKXs1cZOqhwIyjtq
3e/Toagqj8aEMmLX2WAZvHP2755kiENsf/nMEZ92rIjZfFSnKgmwdDWSFt7B8D27mnBqt/FoUgYO
n1Xruic015DShg55x1i3/fZOPxd4503PFGBHNs3VDMN9nUH3QX3LKpCQlPDr3mq/K95+ztNDd1G7
ix596WS2GGCY7kfkAPE8+XdFkYZ3WzVLIYHVXcfLAIkF0KNNBSNy9AX583CXyoCKoK7DMCFPVKOD
RGcO3cwaDwilKvvUc+hwQaXXdL5zoKGR767cYjno0Y5ME2K4BBxx7AAAup3MKWNPX1tzvrvwn6Kq
mAJ/IFT5/5/dBDEi6VVhDl6OTXhXKj/V0c9F97qvRbiWjCzSEofvycJV+lDwKNvZxbfgvkEJT6vz
F1UvTHY2f//vjUR5fNIdqf7OMk4xFMqcS8rsZtUsK6uGwxf17GX+ai7EP95Ux2WygsbCZkFw7pMk
ncii0nbgxoP6yoZImSmrIAAVLEBiGW15Q6+HLRwnsLrfj0vcEBAcSQKrIfOYlV2LhPq8DAYtbvB2
JwWc2QLmLhUiMpBBVGJq24FMR/tX73HDFnqMzJ1ApvzpTXXZcVMS9jtTcslTiaC28TVvZdQpdF7S
P7fbDub94ugIFQcpSLQP66oQxn3IuK6avFUvLKjrOLXCt8+SnIPniYlVY5SBhOEIxdEjr28lkItY
tASV1uGZH6O2dJOv2dxbeh2Uocq2CDjeYQls00vMDpHmiOjplnKmAQb1vMog5YvbFKuqJJpKfQOY
MoZ9XuMCl1sQRP2NQcKKP0GRLI9t/LAKCUPzrpaZRq1Eyx+x+SyeUX5JVfnzfru+/wpUlg+L0r+R
3OVelSQ0C2mBZN0C7gSK7evwfDEkBqpMfFLRrwRmPEqUkq/kLfQ75loR+eAC2WTOjhg61Hyr14P5
UfQNtpMmR0D6CElU9vnon/N8iGcyWMBBam+6upni2Qejbcn5yButOTgFNPZUS4xVNl++rfbcpFhJ
AP2rW8L519R97iz1FAm4d0Mb9vqtMZv/KYHdPzFelNODvfd8SwHNTK5yxZxybg2pLmhYVBqroZtU
+Av+ifeg0VToVwmRjaiYmQhIBaN9kXc4MkL8aeBXf29SziPNF3XGHcTtsDeeEJTTcKffZQAzzFWk
Yz++Uipo0rrsNz432da2wygJsHrOhxKQ/cCQlaYZyyLvIz39dCRYWZ47htK8TRxiPqwBOy5SSLii
SnnBV/UoD702nWEdJVgDHOaAyfKmbES/qsBhqEzduW/KKhRjb2v5ht+eqSxNQuK7pVVoZbBfCcIs
CAP4U9FDQ/uPIgW4Prk0ap14oH2g1Fnxk7D+N1iLfywnzCOA/1Ql7e8FcW/xLmi0mM+0R7eEFzBD
AM4j8jGCGFigHqshdUTv1o2pwbf3RehLIJ+HbPGgq5XHWEYy4Ps4PZXCh60xUQcTLg/6gOvDNBL3
Nejhb5nk+xxuUmnuyfHOgFE+Ram+RkLJXQ7U5/cLnUv8ldnEUEJT0CBZkthNuU4mXtGUNAfH1fET
EPChTVi/lCDJ7tQIg4lyPV6gxMxzfdfrQ/cx4LJ8VMacjZF3cnZAX/fkAfI1aYBNz96zLF8+CtvA
ngdeRUJegIZUy76u3J5WUVW6i2boxutB5Msq/VUasbNb5suq0kNWz5WNoFJ4UF/yQolQv/k9O5o6
MqxYOcbpXL/5fHAyaSaGJsKOtbHRDg5ty902h2hMhbUpV5RGsJTUEDHYYxYfbgiegdgifWXujMLV
1VITw+Zdypi9AA9Hd/WvKJxq8nFVrPPCn2/3X7OxtcMTpP4E4V3nfzhZwxY6YTIw6HRWqw4uYDyz
Zdt8aER3rbuIEIFXUBmK9KSEhYMsV053bYdWbdAfYTYktCU1vdM0rUFXMXrvxSDKZ+ByTcjiY0Oi
+8q4FP+/Ov8gsk3mp/cWqnGPVNIcIh0fGkRTrmlol3BRDSajiBTsai1Vikj79mfebv0WbaHm+0aB
jfKEqTEW4mS50DLWshozxRGwTzs/7WKPhMVCylG/ilu+VCK90v3uQtpEv7d+W0Hn0KJXsj0Kw2LJ
WyWmVubScQl5WzLemiKAKvg8WYAex7TpJODqGTJKQCtbK4vyvQEwPqwvN9t6klW2Cglg6zDndqG0
ruDz/gQNJUH3315WHtwQSN7RHqEmo1WsLOAYYq/vncNTAXo3lfszaddWR3lFT8/y0PtnfY1ISyle
WyE306R0Q9blctIsmK/KLI3kyRKZOFgmG94gU5ltbmijqsJdipUxDHvssUee1jtzpCqnz7T48DJ3
vE89ViJECwf1i2m0M3GjJEWQO7Rk5KU/7HPS4cPpwUoZ2SEpehfV1D3qxjtCgPdiRlZ6QnPgBr3E
jQWKR0CyX5RMHb8PJXWvktZ43+gCmPVt+6/NQpPvfvCp/WUjaS2P3XEnTYeNsxtBDACDZ2euSXdO
RgQKzApk78qBxHN2KCa3/ECyN43B7brpMReTuYzsGhw4q1kO9VXIKTxz9ypZVodgAfmY1hGYOtVb
jkqcN6qe/7CgURcsHezbEuAEDoldJn7KUUsm7sJ6KQo45CV59fsnZ9jz0apwsqhK8G6J+Lyq5pH8
A2QDYt/UHNc0JY6DRmJ1655VJBVYA9obBWqvrWhz7eyl8sslqutDcTySz9GmA29yXTb7tpJKk1vA
ko41TkMqrE0BjHmNpff0ysNxuzsFtIRT5R7apsGDVqTm10PVJz7fCKiJ8DR9+xgejSwuq1ChSMLc
Cz9+wnhS3h9ov+L4g3AzT1ONHTppMmCYzP7uVaZ0BZrLm4QjOoqVZZgDVKP9wnJLnF4XmPXsi917
Qy6n+b/Y+ja3m3b57pKs/6cq72OEFHZYUV9I6b0MuA+JY9ccr7UQ5fWwV5npuCIeLUT+D3GygpDx
fagLRzfoQJd2DKjljPfsP2atcoK1czSczEF7DnNXrYoKjGKkmvlyIZ4WMi4O5urhS/2/353W/kVD
Fu4z+QYNxlHiWoylRJbfhCr02EnS5zg8yhYgABHXMHtb9E7BKLT0ttrZYUMHm/WLZvFb0Beg3koB
uIKvWYC9KCI8Gjihw3YpFM52oGbjx1P1x3OODSs0jZ3bKl23PYstRndTHMZYxEEcT1V5YsGMZH1e
UvyvZcRMlg/ps6Y1pV4C2gfPvD1CB78cyEnDnOlu44Gxm1Q/d06bimPE+APWm9qDYI8gCrsiK54n
4UngWSANuyMvHFHD5G+zWPEHMlhahnrY1xOGryRc6hc6DUXZzczo2pcP6SpKEk4134FZI1+Sw1SY
4NLgt1dOUJG8cF+usQZuXrslTk9MR3dC3VMXjhjtU4Rh6NdoAiNDmJ5sqHcGVsyADk3ip1Oyg4C/
f//xlMV7WwtO61C3voBUSsUlFx7bjUIU2HgZJfotrbfrQZJtlUHpy6/eYW5SJ2zgLntsEAK1KngD
VosCYNi30kFWn8h7pO2cGH1mN16NdHSaLHEilUHrQJGyp0KEGhFFlcTKWmCRPSJGy1GdFgn2Cdj/
DIBzis4W/pNvi/9cXXKcoNjiA2AV51xWEUpYxH+T7j8TEmpsvMVzJfdVVA7TcM1NA491IeWYWH/l
+mAKcLZDNW9Ihti2mBR7YlR0hNtnU6S0vtNPf7WCIqBXYjxKrjn1u+lNTP6tSZMD43N27Wxr9eAk
8armgsl/SDRqO7OgyfHLGbGsSRBVcNoBdH8DXjUnKOMM7vF8nQoucOsfbKdKIAwihZcT1rNPxzii
E5OtP/0YiQhZ5Z6lVbgkE7uCL7Ce1vhR/4ZvT2E4Oq8W8LkUGrUyJE2e0PV/yQ+ri897YJ8ikIlz
+GgWCU0xOd0ZjSJ14nCswwgCLxoWS/8+Xvapqt6RCo6Fpf0UOlVDnjht5pd4z7DrXly11n5/tgp/
2loZUyhMO3EQgCwNohEEda7Yb0Dbw1BJoGHCH/NwIlhhgM6Ayeok65EQ2RgIVPxbm4O40OcRO5YT
bDXkyGUBMzWY8YftUsSyHVf9XBbMaRXie5gdtto8pxp1KaxWEMCXjcXZ+PKcT24TynIIfzlE8iQ2
BbWM+jxSu8jv+0JxUp5lJ3PRrr4y+pGZmUvUq8zkPxIeDHUAcc8KUDyJ2FMmpP1H+rpllfhT+1yE
itsnZzj2OVkMOn3PACedbDP1ONQktbIXUgMLHUNOuhP9eeQnR7W1/C3LQgzkAQvGoHYVY1Oi6ucA
ar8tP/fkA4+6sv9AjUo7/OWgX//8PaWaYCVh8QB7W0zHsbtG+jWJsS7IfE41mXKlCw0W1q9rm9Hy
SePIjU1dASrSRCzw0IDdN4YRdHsVIctOHGIclZA0mHTctD48InM6BieUJzsZa2yXJFIq+7UfE0LE
F/ykErDnfy33TNNnFUymDhPqPULm6jMIlVG1KHogMlxddUJMfK6+cp82NLZrvawAcbGMc5fW6B5V
BmNbnwZRvJxxcH8EsCIYo4bmzuY2Fkm04nLcPxvPZNb62r7tJUs1EjyelHqjnSTmH6fByG7diO0R
86PdqL+CqhGTiJEjIRSFfVtDG/yecQzUQ2IaekPjRcE9cDAeo7DQWKkOhhgob3pi49cYSP9erce1
WEdMeNgcyRcO5aSwbGEVkXc3RFL57p+0jFjIm3S7PSpfQ5b9mELCOZ6x2KOhpkGD/8Z3Gz92PJYw
putmvsz2YqDQ6VgeitoEz7muZtdUtYzn3GKHw5SUYq5cg10X/H0ZsZ4yEjwCgBPt28aDja1GnqL+
RxaLNFtjsIKEy/4EGz/B/jHcABfYBWOdKt3Iv4rN9La/Fz7Zq3rEc4pvqfFeC2sRd13o6dFX0HsG
lCln56uh+xuDvh/HDCJ+dx0Xm5Xzc4Y48cDil/P75icfPMROfwAPUQU6YAMjvNFsPIZ8bLIOlbEj
xlT6TWT3kujC/vhMVS7LR0fdElYjsZNR7QsTEyV8znaXyerzEujP1pBPnLCwODFE0DHiIj8mFCKS
pamB6RhFdUk5zR7LiFiYlg2djqez+krDPH2z4v4lDlJKQ3F8dfFbqih0Op4RX8S6SqCaSzG/NCHj
nj+hnwTVoMW2fiDe421PMPj5GJ/wT8GNtKVhQ/xhV3smL0OXGlL9I1nUlU+zZSJillIsK4imerFh
sAHLxP7oqkfbAtUUpD/b0R2wANS4heuLj9UPK6Muc9tqrlL6vKSMO2pP41PB4IOte9vpQY6gsyG8
GN2Xvmw+MlUeeV3kUv4HjOLNskAth+aF+8oJ2vFlBAvZbMgaNd41YsWiaFOIDeObv57a929GZeeQ
+TtgFMNRLarvlGpYqEQdfBEA6qOpcUVnlkIBBnbSIm/2lAeH7+rsXg3sPK2/2XoYK/6pCwRdLGhN
U1wfZsZxX648q5kkpepPL+7nlDZR2F+9wa8kdFQtQcYbl1OPmL/Sfj8N8irX3Hdz6tXI46tpSNrQ
c/vE3nlnlhJRnZthHNbvZ3dopu3xmKusStbAEGmLBUUWRuVPsHplD09iqTq67dEqNtt37VKTsWn1
5Ii163wdYkMqG2Cs7zNcYbnvwDnIiobYTNyvAN8KD936IaTqLY3S+sT1Xi4ydwyV72CTT2eUzVgL
Kwk/bKdwDWbgc7Xrhv2bcLQy0vtrj/rHlkuSPoMaMuAelrEaVoHESxM9Rf8qZyG/2J/uJFpH5Fjv
QH8RLosCI1yydwTyamIWeRHB+bcANP/7Pckor+wRXHhKgvm3suK7ecRHIBomyNwFA3FRVyaoZJ0i
0D5QkNHfbQsJ9OqVuntOtEiiz0R+ZYGajB1lkw0YFLlpvUJ8QQHG6/RHMuZ4klINkzMQVf4uAHTP
2UWcs8nsPjL46+ujuwdtbCOlKHxz5EpeZgQdb4AIRii9NwwAUKQSYOJae6jNQnlIsU6Jn0aQ8eWD
Xenoe6Wj+2DePbVDaT1yco/fDIyYMk6R+HVq4uZlPQlMq4kimPC4OKLg9LELMRzLPxhriD+FNW6m
dTgacRQqc5X6k5XDEbJ3fPFbsVhXKYDm0iomoLsIUyL97amEgPLvPSvkooJ/s3608dCxnQkk/4y6
U0oTJoQh/2MLVmzcAiy6cwZP2rVAMJf1aRPc1ZvdDjbeJfgm3nXpRzj/gDBY5aMIS5ActmG8HZKo
JTgtYL3XfZ3VHHSRQ4eO0Hw5eBIRpGTQaMy/No2VrV2Gh1WZVoSk7Qq233sRRGkytmq+1v4/9xMT
SNKS59JJkbHeahf2oT/ObCaBjYmYQYzUTHVCzHV3ASd36ug0TRVXixihY73hgO/Y7NSNddfUEPob
f5dn42BHAQKoyK5gRHpsZl8TS60YewRbvcJP+VafF91v9lcuGDzEpGuLTXiLAPCxCxXN0oGSpnT4
KXuf5vHCp6qIHwbvndXsWkHlcjnp9Uw9i62Lc0uVFUrD7BTFJgKDhjVWVJErJox/heUZH3safEEW
D0WKR8fHf5SBisZKMS+TpFH6KSHJ9TR0EsJVkyrfI/HQTSq1mBaHm5qMKzhNq9CQvBBNjaH8xqwQ
aebxeCg+USj+X4Kvh98r5lcLpq7Q1JrGvjY2AfDfCrB61Q+rITNL+1frBBCYWQVz6db8NxnOVHlC
cVNpUMhqzMI/cJRFRDt+mvhqzpqqEba4dNXpghVXuUemVHLOG2v97g11fwdVZYA8aKDIb0wgzSCZ
DMjZ85l3b6ci8fWvi5kuCoWoU571m/WHgWCDVxVdKUOOFaA9r8DmkUgO21d6DIYCAnqDINLRs0Ws
1uv+7TfOI4OC3f5NsQVdP1UhdRk1KhvceY8P+2UJJuo24IqJi1jqhUwLoXz6ylGIqHBWzQPXWMXl
7kSMn+aQuD1X85h8aJ6Ai1IZ+04RraBxbE97Db8JIKCPPWY4BZlRjMBbpSUlTVgrcoA7ekb92AsY
+G/G4QaoSeFYsNSVXQB56o2CSM0X5cR4GScM59mAtsjaiKupSQ5MgEatVRpVAXfkBxtMJyAoXNQw
NkLOGKcns5OOu/HDO7jxftpPVAV0oH49WLrfNtS+EnB0aKvkwxkhtKbgHXvTKxVFYn9kbIzOwAKq
hpo/H0xNeUTsmHEYdBwsFvFy4gV284sQ1gN7UW10Lv8pUJ1VGex07CxARHTYX12Q+x/tZkRM173q
fU4OGq1OiSDV/jK/h9DYyxu3mFhfEgjHMZ5ZD/K78eudbIn+0QW3g1wLV1Dokv4nfnQZcToQKDe3
PF2Z9OtCqpKo+tPICtf9Org8J3AeEG9Uzq9Hx58NQvMp5+2ag8+8TcK7pABXHtNjiyLRlEgnXtdK
wV00Jm8nkOMxQedjzA37hqPp8dR+seK6wAO4ojCKNRi8Olidp5KbfTsoU52+38NlNSiUiWMyT1+7
z7hiHPbuJoRmbO2ZP5qN8WfAddCNUWt0CWm7E2JMWnTwzEMI3GIqLYg1/sjZeVWYysSrz5vFriQm
+S48n//elgLlWmNV5liVWa6TygAE14/5QxtFtlrIjkK+QPy7/1xOWiAIYMZWczklmDM7wW2/O7bg
H2oDIExk2Iv/vNM2EpHoD7/QiS4Mo51lifrs0JNE74wzQqKRleYBF4LfMn4eIa3h9WvzC3rNXu1o
hecj65ycQ9qe6trCNn2buHmbRjnQm9SYnouT2Iy0Ycic/pyrMEde9BUYBKfw/nInX3PyClEOZHZo
yFX72FpG8XFsr2dbpItz+Qaus2NZ257COYwRrV3907vf45QB1A2ayDWlyffPnelt5KNSD/9JxcBN
3+enncUmVzCl9i8xqx2Oao/s6P7LAx5+pzBmM1Hn+u/5afAFA0kyVX7HPqlUXJapGMzMKJa3jO5x
pw9DC4OoIwcv60g2Pv5Gjw4aUPGAPESpZs2pdzkl8X11GC7Vo3QkE5DnDjiMFr04TKgmFnFIZwYn
HkYBqfaHE3TgdQ0ADgGnKfJBHVL2/Ow8xrefKyNk2o6PDHlGLjVo65mgdeFFl4sQm/x7julwLIlA
G8sy+WB/bxkck86VmLHnYHsCMu3Rycbvot6qpTkjy1T5C2vfPCWDtH93q+EdmwLnrz5xb/pdqs5g
WIok6Dz5CeS1yEpBG/sG9JYgDb2EmmBXT28KAIUuW+BJzUd4H63xebP8ceBm1Tnz3ZZ6jXmrXG3i
r/1LBESeGb4qUCMKV72Qm4VsBnpoS5Cva/LGz+WzOVKUwiAd+oF3PkPeqWSz3//Oay9b16Rw8RUV
RbZRp62cIVzUGGzo+HaDn60yivMYosZupupfySZj1fqivzvrbbeLgRrIpW5cGdkVZxPm6FwXhsCi
A9C7InTJJ/CslBeMEFN6HPs/ktuAeU7XzLBi19j9iwUBUtTLuty7j3Lo7r48IPHJ9ZV53lVEXSe2
lGk9dQq85X1VkUFNdO15T0/HqxhrNnCYm/7qAEw4aei/TL3Mwpzk4d3Ak+289mkAxB+3rQauY5/H
QkMRdbzq4gepqjE2HOXYY5MsJ9vOEUh9mrBjnmqfhbk8jAhNhIUWK4ObmP3MXeRVumEsK9kUtYUC
wYOo5NJN3fbXnRx0+4uCyzvcZTHSiC4Dd6kAzPl6otM0Vzk+sfl/pOv/gT46nr9WIaLX7HsgsXWB
lpX0KfCGUanSwe9kiLOtlvlu4DFBkASD9Xr7bcXG5MXg3Orm+10Za/HAlL4HZZvOAq0+0nZmq4xl
KHq/Fb0PUWClxTjLS0pJCOVKUYoTBdP3BW9cPZ4Kk98Ggm85g3Xettr5dBLAlk8TPoOECl9UOMZd
ZGbnkZbm/xBaY1gHJHMWlkLi7hww6Ei8S0U6ueZOw0HYO+tIwxqYiDo8LAX/+a9YPIQQ2OrHeBmF
90DZIEKf0TWNw/2SBUuun0EBsoPpNIPE56ZCEKh+YL5jm7lRTMrU16upw6MKWBOgMOn8AlvRb0if
VOZUXn5DYuf8c0x2u4DA2kPuEJxx3QhhO9ggeRUBpf2j+37/dvcfqEIdLM+XxGI/cZE2nRxrqPhr
Y/7xBfOVeD158bXwfhCfa3/pXjw/BYNm1Ni0nLYZhK0OJWINlzvz1B1m+4iovcbNpxdar/uHfR3K
bhPAtCVtSauAi/L6Zw7W2rC1po5U/H/B01Vuz72bog/2RYRyeTr1GunlBYd9AebjpN44vimeoI2r
aWWeiDVff/nH5HKhSc9r935Z/+KzIghl9Tp9it8ghG3hiXMHOVjp1xf+447jclbrZjUInT66Xpv0
2R4KRjWt+yo6E/hlwF7oyxRTayhg/qVZPzB1Q+WgrU0LZ+U4efpZ8uDfv1Z6ZbXUMb8sOZl2nrH8
8JzLbFZaxP50Sp/qGsh7noyjpbQCgPh2FemJt9ueSiyLwheI8bywncpHOV4Lt2aprNtZ+a8RVeFr
5+JUIGfKKjjkvxiQHKHLD+3H2iRGiD6v0n5tfUOmlUZL0TSPFewyeX6MlGRENBOjvVkT8iXvJbBR
BMqptkHXeEBGsTjTFWyNXfT1xYt3xCovAyxJoa0Mda41gep29CbpCWla8Nmve1EVG6ZHZtu1k38x
icNBIa9fM+WiOoiAnq59MCEdMpb5ChvazhwwA1SBXybkbxe6G2pYlIY9WhfHuusDaFuKCZ1ZB7hU
KgqYO/H6929y4PKSR6rA68oK7G59uYLnOfLwPZZt52X0BubzIwbqRr0eixa5sbX7bTrofzkmTleh
83C33DQcCPrx7uSdrQLZEeg8lpB23xgw2F0GYNYy+8WBJOHhFKUe1Jt6nX89LhP5E1T5kARh8Rer
CDfa5c4HQnmoUoqt2RyDLCIiRlfDsXAiOeNJCzGzU55N+nQKGoZ0Fh9j2TXtkrIUIUi819Z8aCrU
ctQulqQPg3uMYqR4Wy+XxIXgRDeOiuYS6Jzis55/gmSNvgoJesozX86Bn3dFedwGOF1jbf8TF/qH
VYSuenrgR45ghFKBbNrLydO3l/u/JtCJ2Gea06Y6b2UIOWg+KsQDd37DNxWeFz2a92c5XD2leeR3
5aGwYkHeSeM1Yw/w81OYKkMrP4//XBdi5QmmqPnfdij2/+p9EmnoF2LBvZqo4LdbOAE8DLJkrkt6
7Fj4P9iuqdZ4KH6Mkge4f0tN9vtpbfEFHCz8llnBYAk0rVRgd0FcYSp6ElMuAXyBt6mIWBrcB4ff
2KjZnlfDJEVdgJy15gbn03o6oA38XIZkGt+2jMBLTrNdYzdpWiZWlphs1NL2y7HD7Ro75iS+qFjG
wbsIzvGRgCbNHcW9u9tnqjVeEvOoh0JF50Vf27pAHW3rIgdCowdylfccrQMttVedy53f6iGgDxoe
Od9oIdH3g9t8pvxa0C3a7uV7ruBn0EXg64r73JraRghIL0wv9IT/CRZ1QehP1Rf68ZKGgsrf533p
RZDP0LCI0az3e/vfKmwuDSIHKfgj6xV9dk2TaUTMeSqr5C9OwQQdtmE4X++4vf2Epyut+/ssIScq
9ezoVLZO2gq21cXleU4V4I+7SMYkk01J5ejzzKLFPIU8l859dL4FIpf/+z4XubGPHmE2dxN/grGk
vVmMHl7DgaoFdb7zJUsOHXvnvqzD4jIUuU3hUU6/A4YAWVxXyB87V2QogYdWhcGwXDzwdqxgKtmI
Mt844SAIAfdKKx2oifA7PosEFRPBdu6mU3eP3JkG7yKeNqJ3YF3dZXp2l1rMczxuiT+Ln+42dJ9+
/95ybotJGHl9lkpuQ6VA4Xc9tHhRxwr4FxZu0Rx8bzOn4DHOuurzZ3CWm/goCqTZuHKYdgXluGbV
WRQKMU8H8H+HQPAHW8dRv0whdZ5PSsUZp7LsEmGJgNNbpRhk1xD8rpyS4asJlmhy0A6h5bRVsES5
Hrgibn3B2CoAsIlyp8H9Te4xRYW5JvfGg+9bnknFTnWe2lJ5sATUosPmo5oYcKyf4NMOq4l12a7D
QezMrRWJDdvmQfWGuMGF4QVF2fR3hwpJrb2J6TPF7Mr/TTx8k4bzVwn9QHzdK13f96V06sv+kXGq
GtoiRb3UQy4ym+HKjefqPR3Pg+dLFzJDNI7PPZI5GrVfZOk1pyg5sBr2ucBecmUqZ1xavMApJC3D
S5fXaVvqoKQQLXIKcISbogaRZaaD5gwNV2GIiT32LkDYDs9vCu/h2vs1iHEx6g66PNS3S4OGdQFT
CtnB1Sl9pkH6qBSaC/EmrJqhJ5bTptRjVgemiINXbfMZfMQS3Fftin75lEp496aaIIbcpr52WifO
ToHaRTHJbf8yRgTtios2pF6NxuTiiQEm6YXMwD7kvLjZOh3iD1KQY7C5PrSPvM9u/qq2qdARLheH
ifu1Zrsx2UiFmWORvLyhTEveKL1wKRu1ieQc4k1ItEVE3gGNlSr5SqSI7FXJC669XtB0BXaYs/kC
DCQLOxBVWlZEVrOcj2M0tE6aiub+xai0giJxiCzqKDc7r7G1fYv1/VxSUyNjTsPuQBDsI0Q3lRpS
k4DU2l2ra/DTkAK9CXAkoL6qT7fbrbe/b8MwNqO7/vUCCejZfhK18/n2OVHDAUILerLFs7qcm/ym
teoXQl3Nl2ZjPyAlwSqVvOoJxyxd0P+34gt7kOfPR2u5ojumdj3/qoT1BaceaaZ70M76DLxpx/tC
li6FMWUNWY3QNvvzRT+IabDlYrtqupNYVznBn3Gf8tW5EstY21jbu3AMNcHMs7+JqNOHbqQutYJv
jEu0Y2a3On8EQUhQZdB4b6TiQKnA6m2V7+yuqjiW7tHonBKaf29IYLd1tOusqBSsthZvI/5mdy5b
/vxdI6btC6j0c2K7SBVU723pKB7zgA3rKSMVAeF5kHk9HABvfCTbDj1xj6W6xX3X91Bso4UYyVOw
cKTmm35lQub/b88+DeUXHuj3oHr8nhw3jQo/aIfL86QzZGdJZBFMn7ZEQbMGftEJUEEz22uXLWXT
ukWMlPP7NUr+XLBgobr+75ARNJMYBWg+UwerKwWw43fvh0bXKQZE2s2ZVGvgKS2Habl8Nea91Boz
kuuoCpwDk3iHvtG/kHKTuPLcAYXVL+RZGz29VyMLy9cHpDYy0st+82U+JDgXkDRJmyxFpTi/dI5l
Y0Vo2g5B6SSmx/OE1tKUvGKHz2pJbt1bmBSFUzKt3yToHW0/nMWiqoMmL2HN7KQLfRHBx/QvykfE
mxTpvQEo0cRF9/ybIpyQOt8KUReAx+uZxANk2af5ZhVnjCqRx0oluJ/4s1REC59JHCh+4qlGmXFm
QcapXXZW0d1aMs2IsA2zzJVCnv9W35wFYNLryAyTi5scNsTlobiKaUqhIts3hvvAGiEpTPCnzgWN
LmhXFGgFUdX3xcPFAK2PtYvq/0IIpnH1JeSq4VeSitfrPxFpI4/eF5Jzgcl6fM9+lOlEYH29CAfc
F8wglUXQp5dgBfici453Unf3AydcKPYtZkjaSh+uQ6vf5DoQAS/FBKEnvzJCxmiMAvFICzOcfubA
AdmtKNks+5wefl+HxPIOyVURK70ZnDzmxPJ0926yysr6XzWnl37TWS71A0+I1byNv86ULj+ECPW+
cDnr8qaGBRuxSucV7mnakpazQ07IYO3ECH5mbdZlXu+tst+xjeiOc//Rd4gwp0xHYLln101w64xR
Z0GjjBw66XXhqaYuQlPM5Q4nNQ7RhQBbqGo7oUauAFnRKvTrlTZGY5ziZU31YoLz3y7IBYgv5dkS
eomgX1xw+OHiREKSjP9US/f0//wYNguHI+yNhgV+/MLIzFb1Uye6Wpiz7vWZoXZP7FbnLvARwHMq
hFngLvPJM+Wp+G8iMiIu6gzHuBvRfCftxR0fqBnzVif7dOeReoxS8lfpl+sHetG3PzygrMvMjdGf
EDrNqTg4NWaNeLFC0MSAHkC/dcQFGuv4Dc0Z0jpeXTa4HDzPdNOJYY1MfG8je88hOssqrQ0rmElV
iVS2AzeRtBBmCg2F3yURHmXyESwyK6KXBQje5ldDPK1xvPi6AVfPskqZFg9NHRte0nkihIW3fR54
3lqGBI7LbaS/EYiUgvWgjAcip8oU3+b/4HMjsd/z7jVB6cO/8ctvW24SSgzwd9tAz94qQayV5Z5l
mjSwZ204g56JixZdfkneDJWYKhbetUSCJnSdEnBSiYp1fYoWegZR84qpiwTo49iwIg6imRQ8bQjO
l8ed4dTmit81pfzVRKyFLvQ0Ct7EDmMxGW7ky+sMZdk8OgRRlYd+h4eJGXmgfpLfubz/SRFTTPeL
O+cRoHdnvC4VFZvI2tQA5kHsVdwHZI3cgfqrB4u7hxigwYLx7jwsw43Mi+NTVGE6hmmEvqc5GtaR
y/CaSv+dVPZCNGeqNmZdXRCn6dUYYqQ+QuqcD/Hp9/KJxKjHWdvM/zv0pbWIQaDGYEBQBtPyPszP
BgQST6wJNTpdDaYJ4Hak1ImeL5+99vGHhiA+j2L0t1fVJjHZHSbaiPZsOA/NeIYr6bllp9zCNo9H
gX7fYGjr1HKhK3PxMn4GYr+6CmbyT+FPGLi3HLJWkoXBoDzNBBkKBvVQCt8AwQXEN5fZWhY9WKsp
g6KNoWcKffbJF3V2lFp7dl9d8O/Rb+BavxE3YAKELFIV3PhYhgoAfYbCsbqXQH7uEALwFNr9solF
HidjAOPcC64r4hffmQX6uKNXDLgJFvHtzUUS6ESLgYnAMjpsw4wWVRYouHD6ob4IuM/C/hs1RmrU
UvrOUJZS/p3gO0TVjsw/bdy6X9FXaz0IWsrPpy48xfmE06a6nSxSzXaMkZPtIzcUi3bxtAedCdYs
/YkIPAFS2M0a+4KMrY6A38hdlgFiEN3WLPOBiQLOJxJ/iOhvUMpKFpkn12HccFMk8iYta1QU+EJa
lrOYG3cOGWRb63HXxrWIIJStBZKk3zGUlv5WvTs/MHK2hYfuhRmGIrMrBdnQzdGPoHVBvv69BDjK
aj7wPr1sQuax5wUUXUMYgmHxKrwAYuUObwEPhviErlHnWPDI20FapvItP6oaKBLhVW1evlY5c5Um
9zs3y+caxh7/X8C8PSlOuHL5XHe7rIUqfmFNV9ch9MWJVsXJXo03cmt2D9qd9fEQGJL1kwX8jnAe
UDSugKuAp9sYL1JRV9omNs59OJbuxeeBZzVjMkkQSgzov0oYHnwYGhZp5aETXdJ0BKaMNlISPgKa
K+z71nb3jkGP4o78qcuxM1Bj93Ai5GxHRsnj+6BdV8T2AcUzHoWtvAQtgCyvUuT2Ao7CstAklkPq
En8POTuADregqAMLFBKIyXpVaUZRucgXeX96ZRP6Af052r/G4zcDKOuNWmBmmr12/XcEuYYx3Dg5
F+CEXhh3pQjY8YxtJYxw+LkpOX0BJqT3urpKPpjKx1Fm1MXw8jbPxtULbPWjQVCCagC8hjSFgn7d
SSDxqHFnsl8MnE9VBNciJzq5/6ZFH/Ehqf9FmXgsEV3kNR3Qt5GWCpohkDxdM+jx8SGQhJNK8t6x
PhJOcETLaV7kMGGOAQzMEaIRTZO8UbNgbm8iRdqiepZtQzP+sF5GUgFBWHtRGW8Wvoiq5BwRhvzd
k0AowCjeYYmm0KgZn2i51L7hCx7htwfMNTBnsnpul9lGBNP0MtoCESgymWz5alvTRth7us2l1+sd
IhgDE6pEOeIEqe1xV5IdHCdMuwBfBKr2lK9XanDsmEwdalj+GHsfZqM7WhWvudbJBuAMKod6EXsz
cudQe74ThThxBDKep9y+mxS2UUUxiWrTq2+uqrduPzcdTti0b/WHeNy5YAnpx387cHvpkrRVFWOb
lbpxOoSzZJewthfwL9HRgl7jpdLGyUwqs375LA/GcP1x+BSizY5uKGVJslPHxau1r6WqfZI5TtKh
CzyOKJSZ/iqdsXUnXlypmfLYAchKlze9bkgdh6+ZZa4FctgGEh7kNbS0+Bn5W7z67AQOX8ZydwaR
Gdg2PpbMwIMMxJSJmJODT35m3jPye+2w9ekNXD0Xqdi3Dg48YgQ1FKz2Cbedw5AkI53EvoTPmoo9
J7YmIIpIAGqyPxcHIzbKhe43KQfAhWd8ePVDsBUOT0i/4GkBDtU+xG/2upAbcNLojOYwwNiHqJ2j
921FxSC91nr88okvj4Su4foWBqaxaPxFn1rizeim3dpkiV+81Q/GbmIUsVoN0LZgPBrRpF2lDTJ0
IJcGoDxIlmnPhUIzcZ/hXJ+yu+4OkuP3pePJfGCPLE0yP9seE5Lfeqmwy6RuozkYgau7tHaN7E37
tbza2kxBh8rzpIgoJQHBieKa+/aKICbkb//AXQNplNnjLi/HgBRltTEZWyurLnBzyjGVSsr8srf7
5+lWr25fKRTYDeg395ih75XPIHVnsIbuMbjswnMFvGnNDzavsSZt2HJCacKgLUCF89kt2BzpvBi2
XK2wWuRqmDQoVrpstc86gdBfpLcmCttx1AmRgE3ORlIYzyV/wOvTFgcECUFGXS62roMyxv+wGtSb
r72f0x1Yw7PKaF2vtJVg+/8xon8eDgDCuqsJ6yJI8qFimH1u0dseaaAKZ2lw3cRaeSlPKnSWoWst
qDFeqOTQDJF6auiAEWPf0VhFAoAYWT7Cr0vo7qJoS++c31yUo2bj7rGuSaG2GyQMIzsG7dka+Rej
4tIl3zG8pOtFoHpU8riSNNvs0WAgn7z1yoVuLsus3fQOVddyVVhJ4VbZ2yCn7NYQ7TguaC/h2uVg
Ze9qvJ/uOSJG91c5VN1S8Q5KVt+IuTqcxeRguY5mm3q5WYSwqXuWl7gMUDnhMWL95VyPhrgWOpzw
wjHvkdsCv6oPvSzeYvdy44v72BUHZDDsAUNjKwxPDW1mKUh94wmigvxQDL0pmX8HZjV0GEmFetts
2cLEWsl7XnDnaeVvStQ093azAUcKScgbic2PrtTHynGPTlfij2E/KWesZa2Toz0HaiDu0htEkwQf
PJGKqFBS25ybhfwvw/3kXG3jgqqq1gDO4HJ0WHhqVK5eT0GfaQxW0cubDoeKJ/CBZJuBlBRV2FrS
JY0mPu2E13wApUgP8nmQaydCaNjAeBsjFW2+BVm5OrNKYqBQ1p7EnE94hv8LtE2s1J/qClWtiMFG
GSg/bhAzrGaOq87QsDbsSBK996dV6qAAwxcYcf+WOteoeOA7JYavynomlyP+Tq+pACnDxKlm9pBz
mYTQJCTnjomisHODetR4+QsdnTd9eCSaOCUbfZLrXm/IxuE5WQOnGcA2PgpFWZauVFo9vJOJNnqq
B7v5c/QinJEk41xwin94/mSgKWSxQSPERs4nZCW12qIEWenRD3Ccs6gV9Kt2DDTl/+7bs2+DZYKT
zBALH2Y5DbBf1SogFE55QxA26CIZzUcI+zJp0Cy8mcTmBuhmuES/ceNdxnZzTiii7PUUQRJmFMQG
AM57fWdW0HAZPkinZ3/tP6f8NL0DVy8TzUFR/fR4i3odMXmw8yTtldcX1/BIA6WM234aDbIhhPGL
6Tc6AQcyu5TXSCTm7qdFeZT1znfNGCo/J4G4CCDHpKsOCk8uqtIj4sIsOhVq3nUmuF23op5aLE5N
7u/oFEXcuoVOMnUr7rWPlXZaaFEduYlTVDFI2T5Vk5uF9qy4WvWjGpWvikwSDRSzFaHdcvH9Ex4+
euixDEbPPpe7z4bNNG7IfvdjvscGWRdMjDpq8BiLhzKVhUBG6QXz1Nu2WoQK2qz4HNZj4/SCs4vF
kqMwlU5qowKlpiA/xeNLUzMDXOPvB3ivF07B3hBtxEwJ6sWbKEEW1muB4iTnNRlHGGzod2x1wXCM
UnlZfYgqq7Mk9PYx+aFIyb+UOCQWcmmFqp1J12uOYNwW1fOnXaRh2eNs2GSjaf526WrXibj8TuyQ
qzk8V1EAOj2Lm81iuDzCoA1e111aBI+cYcjdjX00N533OyhadTnJdPTIQD8+QKIkf6X/9FYk3Kp4
54KZ3eXC90tNNJjkql3Ye1fshD65ffs7Kd9xHye5NZGyEG8Ej1v/GqJYHdsZqIxCpD/7QpUdvVuu
/Nhi1BNza4E2Dd/uybw+EtoEChFPugdhG0P9tjnG/6xCpWa5GE0HFjrnzs8lhBM6jJxM9wEmN/s1
RDx0o4HvVv0/K3TgX1DQLKWIpyxpp+/BwbbSeF0AjwrG40ruvrisSyTUSHSb3Y/0pW2v7V0GZ6uY
AEWPaOftXLqtTJEjakAYxrXjkswiSDhw17l9cpQRtBmvjNQ+ct7KQmXUm9YWkWVIV5ZsDrYhs/q3
uBhp5YciW5xnu5U1TufRjRIs9ZSdmGprn1/6VrZPEQMxN8fNhjavjYg/O/CelodtxyqsPW5Wj6AQ
mubS0Jiuoq11IeEs1zIPoJRldVGVDmkO17iTekd5wNIHmXpkk/p4TRv96MtsehJseAxK3hq0y8iX
oUUp76jx+fpUJ41SyCTkViBbnhe3SuclM5DfXFbl+evaxSE+ZiyO9qf9bBy9g2u2fUnjYvjPaYlu
n/9aHtH8wYODVyLJrcBDmRfxtgZKqjaFcuPiQnfRPzyiMHBet2auJ9KBo7f5cwRyY/7D2n5rC+cU
f5UXapU1yw9HVXtJnScPujFhkjFFxx2snnj1ZPJ6nx6X05SDe9D9tbpgNICn+UqgIl7Rx1OJ7MKO
z/1h4JBC0SpueAR1qpbm7X5Dgudao7NTYeLuA5xgm7PlU5ZocKkU3FGgP6LYBig91PgMk9z01xJK
qaKREXymVNx1Tq6jKgpjHONmLb8GzdQsm6VJZjDH6u/nIgRen94ecy30ayl7SFnFSQGNhkOg88We
ifN4+J/kw6NNkQKU+sa9EFlUt2KWC6EvsYm7XbQkiVWOdVIKXwmXIIktagwsKY9JQmXiXR+8ywvx
tpfM1Qb+N0VKUleQDiAM9S/yZPvJlHw4U5DS7AJfGj2BkwBgMzsPcyDsL48iMEuEKHuJs/2YvVDx
QvW+DgBDtnifOos2l9rxDOYByXG/FtksX9Pcu86lhy5ENBaUBpAQTGQTKUFzU/T+llPRc2XMqoSM
RjXPbIbzbUPtTLT9FGfKTeHDuepU7V6V3aKAFjQ5wkfF4UicHDgwjpQSUSS7nvp7eeMs2mh/VQM9
HBYNy1RZbO+tTAvw+Y2HSVcRlEKoWN8sWfPRhKbQYQlQM7SHHRYBbsJQSLg9azogSB40cwJK7u4v
fVKmS880jeGF4XDZm/C4cJ2Y2IAmtSB4UjR7jYID+cq4E8eoN/H3GVaZoTvej13e3KreTcTvRVcF
keL69nrCZaIvZMbjKAjwn/MT6zcp8RoemZ/1uxGM0Db7Ku/AbTv90T3BFXTgWgnBBUXVrO+/DsBA
og/eTr4GfhStZY8ndtPmYTq4SnqwHGntr1m6V3I8njCAq0IQvzEjP/mxquQv4yK6xJPiHWojCrkD
oTspcQaVapYNXM7Q+YLB53wUVEOjMYptdGhutT8qWJIPwSe5pLGEVceix9QNcs+vFp+Qg+bBFJgT
i9PoLZ3jRMOSq3lQ6EXqVSY1nvKQ1LoQ40R8QJR7qE0odHiYraypjXAs1AQUG/PorwMmzU5HfnRM
3ptA9cn0MwPjBEEJF8d4KuudYSHp54qYep4Pi3vSw0Tg1bXa9psoajccRwGbrCVlFq9sGpI6BrQ1
tZ4oQ+4IvEbMUkpLa8d8RtueN5rwwjqzvxwd6O7l11BOnrVVYSA/ssIUm8hP5MqU0sHmOjrVn3Zb
ZZj3X4sm3/EfNw4aFxfmZDZHAit3c7Sofd41hbf/P7jNwt4Do7QaH8oDg4rxBjhpKufuwV0y9c4R
Qhl7wZQR0a38qdNX8FfkEMUidcEA9VUfCvg5MSjVx+ZQrsNwwenfP4A9nvMbbHCEBkp8R4UZ5ZUc
E3zCU3RmHCAOczxnpZkSrZwEV6JuPc6Caju827OSNUEj96wQ6/7GUtR5h1lHc30B2FGauBlur1q6
xS/naNbFQ0PeGXMp4MiP4v6Fu941kDpbnt7WDKGGl/Ml/ApAfCxR8FdGNnHxjnCo9kQazxtvlXxC
BdUWQ7I/65q3gn4hFTtkcVQUtcS9SBGDI3zdJr/P2Ea+ZLYs1gPBqntvmoTyPvTGvmxj5GBJQpyo
tDOOHdu0eyNtjZ2C9aydTJy4gplqDj5KkzC03JvrMqGrbtR//CQj5FeIzxM2G6wJ+1+xbHuuh23I
zImfjpBXm6532OlJI6AdHID1LQH8IfbuONgzr1MAHpRLFbQoWUlS5EfyPPYaylRfanq2zSYQDL7K
/J2PSChmObu4f9y1wLvTzZ1miqFGCARtpccf2QUr8sbc8KcvxRTxFF0WMTLHw2zI3VrFa87XFogR
Q+AIDYr2nrI3edRYeZ6Ewoicjxyrwwdydjj9Ik7jPwSapZxwoJnJFGmQ3wC75hYx0ubNcROJuXgz
idNMDixXqY8sXeYfRFtC/9o0Pnl8Xludcbz/5tbqE96+LbaB6zpGJBs1JWyKT75Z1DLuwajVePBM
PsmuXefSRYKixwtiIzOmYMPJSosqeVQRlWvnD/Ib8WPS92fg2N7WoevDppBy6hix8CljlRgW2X5P
+ytfVe8MhEkVTOCgWlGRfJeag84k5/cVMrimHD7+JUpH65nYjXKNUOIVocXYT+sVFnQT55de2w37
3Yu8pYRpJvatZdvksd/QU117aHTk3livX8k5Nuxc0KGYwL8S8qF2p7jWMtLGIpE9FXb5iO/JGCTY
MarzigE90m2zCiMx62d48CoQRvEHVdjjTWgesRiTIvtmG8AGqWzmrMLDxTzSEMZGE8EW2FmU5QUP
8NzqFjyVicSvBig6Tss7QyjncsXrRMnz1bT82RibJJKUC3Q+E4KbXcRYLv7tbk/LfEDx5JCroPOs
6bCtt88kIOSW5p67WGQJqqT645J6QoptVCucWTnPaWl462vWXPeRgXHWirOONVbRB5bT4SfkxLL+
UaPlYKbMwEkrxwtu8NsAxMNxmFuS0SX12NKUE289hmwPENRez+dCvn8FRE0czV2gzqiVI0QARdTs
ZyJm5zdOHOKbvbtbtOBCPOl8NXbIckJkP9PMgne+yMpr9HkFDdsqIsXuAg1zbEpyBUjvOSdZTIh3
28TC01zlHb51eL3nUitLh5UDZ91z91tAwc1S0EOQCgh2ElfOei5nS4Hh29SDTCtDEIhKdbKtaHr+
ux/HTLT4OBbf7Vg543FFJXIFRh+GS8aqMZGHElmcLCvcwLP9q02m6vrvWR0pqi78MpnBpDlGNqdy
NbQFl9pFzjU5wVvsPWS/aJHXEjIzwY26OopvSXzN92Zjjqu+ABhmPPYRAnidBhgav4h1HMBcDuPH
Ihnx8AkIQxdtGIb5TyW8C2SeGL18eQ/PwizBfxAoQ5N0rXKsEruoeVmNbbdmMra7CsfFtZ+pjx4c
9qgktvtWEjzgM2GUJyCVx6he97q5GoTb9f7FS1yXcss7aJ0AaLyCOGBQAYgK+SfuMdeNytgMKK+D
gauBQWqBexJJNuFuW2cpzD/Q+UG1XzOMQuc5higceETg4rmlV/OXSFBWev7LbXmwpmRgPkG50VQS
q36t/eXNL25I+sS9nOYlczekHLqgVcrnPIWkdBw/4IOebCdAnrPs0AS0xesYT60zznWUNmEu4/yF
ftj5kFvk8UsDo5nEf0X+1sSdE96BqyqVPWmfzdoMby9SKpvBYwUW1FQg/fno5jSoCNgN65SRFASr
OXsgVIbcU95UBL+aXmZgLWLxrHDGOgMXsznVwtPL0RTPhQP4u9loxFzNj6Owkry1X/AWcs7wWGAa
DNRK3HWnVvIfX9kdxJtIK3YnHpDiIFnr57Y4U3PRMr/KTFL6ENaF+0cZVjBzsFTSP/vemdOFixgM
7zZAtKeEdGOav+FsrZbHTOle2uaj1zLNfV2MGHoJqh/j3GqWx3NIlPhpqgUIIQbkOS4hy7oLxQeM
fuWmcwgOESazGVyEDm7y0O+T3SYg8Pl4el2/OwhVvBF9wBSgS3MiZggA51kUKwWF/C1c1A5wRNPn
slMjwqZxfYZiKrqXc+E8E9MgMJbiFnyGq6A5iAsjdqvuRStbkMDVtM8VYofs1yH1AgG3Us4MJ60Z
RGkO77PH3YD+D1/brQxF/iQSs32Diac+I267tslOtRDxkTQRC41Oln3qtYlowlZQTrz+11lHg8qn
zoJu9xKpcAcpN7BBsf8RWzxPHOg2fCEY+4f3Nj62dmdSZM01YsnroeXK1XhXhzz2eOZI2Y04A9Qk
lfMW81zbZ5LclUWwXOrxlenxC7L451g7Bz3K4JrbGWamYNdYx4DZzfmIeK/sb0Z1q+sDZAqqcb5l
JBy3B87CL5YhqtHYGEI1brT+7eLG3T4NpHRwW3RM3Bp5ubQIIoGBQAX53E1TFIAQV93QPjYxue0t
DNLH7M2h5DSFQPUogOJyKGznugterBSyx0TtDefHhoZwCcgNzuuUV/2e/zWcKJjcQaflpjqMf4gp
dVN8fhJNzPYOt3tzqi0C/5DlctN+kR4h3S7n5x6gBstDiu7PL7jE7oEN/T9LIPA4lIGM6uGNQgZf
NHaH0d/bnnftbAnRSX29nUkClkh3Kcpm8gI/z9ztwryF1W8DoU4WQztHWIIcLLmpbB3yi3qX9GBk
j8HuKoV69MAA+vCbK8EYqx9mhU2DJNuKhOObOgzG7+uiJZ5BoIMvhLjgfYCsu+29LT3pW1X+P6tm
a+23ErPCFrMhIdpssw7wj68lw0mt/AGXNUfoQlbFx7NBQAqKZE7nkljblhT2AeJEW7boS2FYtdLT
dCzk9TBauhlMTLjYyDa9ZYLZcIfQxEZHgyirWDUu/AydvI9ncP9rNN9CWlmulwm6IJTyLqQuVjNy
wX9x9Izd+R4oJ2pM72hP68Abiht4yQU8ufBUwv/tc+tu/kOyyeooNbnIRCBeLmztf0zlW8UF60Mc
QSKKlTFFJag6Vro/ADjvCGwkMAZMH5xBk4bJb+OnfUCQcAHuhKhr0hypJb9PuriYankQcjUEzV3G
zmhdEMO4Rbws7AgQzM6rzv2bmpwovjZFi2g7kaV21Q/CodJdBLHtVQ6xX+qbioWNtDCZu+D8n37p
4zEfS9yvqFgYfXXz5Fmrr2XaS45V+0IOnapLzME3uCGOBPEG6FJwtlcZO5uj+7JIak52L+qr4XJq
nI3zVv4eTuh0D3xJtCob+6Fb2CdLyaEy84i7ai1464C0wZdvqRH6HQml8FUyXE/6yvu/5i+wiqSQ
uBqjEdUEbTIvWOwv05+dUi1DACYC8hUgOHFgfl3kqxZf34902pLFkW0CNJTz/F5hQ9UNosd3Apcs
1rkS8yD6HOdvJThha3bDE2QwfgRIGTI2dLMI9p7cije0L4mAwl/2jvAA/r3hsoYt5ZGGEAKgWmdb
qU0ZiE68MEhRvgYA2P9P/pINuGeADkKcyCAF701Mw/lp7BSjONaiibbBOvJ2XvI3KH8EyBeTv2A8
dTAWUlnl/owviGXNkCNUFZ62AtCS7Rv9CrSkdl17Kvkc+Fskxheo7X6G8EFU/6s676fx3gB99RYS
VOYL2aeDRNaCmf95NNiNIbT2//lzjoN6wRijxHl0s18+92t/ZSCt6Yhyms8DHLtzMLcHM0YmK36P
5E4elhi7yJJe6eXz9X9PyEtsxpeZAVFzIrHd2JINEUbTHSwAPJCtZogAXanUUyfqDSVHIVSn0tUu
bPh492Dbun/hDYHvxTkQAldziVY1HPWBnO87OfeuUZIs/jbJkLJg+JxMkwG1pSH34DW7DeR6/c1o
MqEG1DGf573TC4LWcui5jG2VFwxWXpgWJk1qd4BRUNDMxTECoSf7FW/cr88BvUaV9IKvtl4VZaQO
LZc0pjAGuLBsTYojCGFdponkHlKJGoOkj36DePrLg6RJxKdorNtlgBzBPTS9sgsq+6R4eGECBFey
gVfkkT6UJvLJCn4TZFAZ5ZXAWRcZdDFMgCHFfn5FfU4rZ3DoXSDplkNhtANDZv27Dcy6kIGi+feL
0p5jexnuDDarU+iqw0vVYPSAlW5Fy+t/RJQW0gpvbM8g3nKqHLq7boZRcghhXVp6mCqvjgLIZXFR
e0kxlt5h85dtoqSWw4o56YJ3m14wZnJXDi2qwbUNxzgD56ov9jWcx8e3ygTJJ+/uXWlwLbxHH0JL
VZUtCXPKV0eLZUAfotlChNF3V2FhAhmLI2RqwtQb+La2J0JIH/OtyUdCWu17ePuMF2uX/oz6RBhB
TIThOWSu6MYL5X7IMD/XYc7FebQPsGTbqOBUtlmPDYr95oQX4B/4ccvvkHHuJbzW+BrayWvASbke
0K5Ml/EkYY6slvFiEbA79wFv3Wg3kRN3/g+RMg0pV9mEqeQ4YcEQ4ZCilfnoRkvUzHzNugctOpM7
ZhQMIjmSP8pDBtzTL7ZhJlTIzixTHYKkJt3oWUoWQyhQ43tXQqmQR2TCW1HOV6bzI0iiV9VD1DJz
8Rl1DN9w6Miff9l7pkJ0Xh7ueSDOsc/Q1UumdZIGZIN9pcfUI1ZEVQEJA7ORbSICmuyHFpybCU6k
gFnEFfmB+UKGN/Nh9ZLH8mPaiJcLxOPTFrSigQMoiDakp3BgCDLrHX5AXY8ThnoUxqFj3c0O+Clp
tNMsVuyfohhVxq/ZTwESlJKsnFKX7Ti528QAb1CNcaCqwJSAYlcPBbbh6EfhN7G0gXAYaiQ03eV+
Zy51/+gGk86a8y8qEFJ8EU3kM5a6/jB4Oh/L3ND6HEbDPKNOjbkbKXUL+/XCTvOCzf10hINpSSYE
IQJMN2D7waplYv22EDrsHx9tUmiVCjO3/D4QBBH0x9YHjsu0GUADxzYNewh83QfamNmoNywblhjA
9Zm7t5ZG8vZOXFi/hRQQ2eEIKx0jGGXTPlfFEKIoGtAiY+x5aPUB3nT4yiSmvsKOLigUpZkflvfB
IWa4I5fzos7OWNPGsUNDz7aQ8ukvnsdiF3xF0K1VTPNk4/+mZXPJ4W01VER9l7QKCxJpFXpyZf5X
K5RYYa2uq3pA/bw1YBm7b5E92ZbdHtlt4PXubRGBqsMxTJuhuHIvFOWq9rYTzRPyks+mnE4bZbot
hWXDO76l7Xf9V7eTYt2x3sYM8NeoPxzHnFIisI3vD3hsPf0rcuv25rlJZ2hP1aEwXxofLJNKQZAQ
Yhg8Bao6jF0SB33bFnX5FJ/xJ0Sm6onAeS+XRy3nr2IgHQ7eCerPjo3CjSoY/MnOlm9W02rpP0ZZ
FUUmq1bzR6/yFO/0VETyc7OVGvEVmiSsuOCvzP75ZBN7vbONs8bwpHIZx5tPcV0qfyR9uvQzdoLB
BZczNXG2n4lssb2EJi3ySRJ9twKmsDZLGnFj4XKL6ACmAmdYvi8Fz3iNRgV762w1vOasSzVLiMHR
4MA99k2PfdZBcnvkvQVnrE88fnBvGHibrR/52tmI4BIqQeHR0pDESFrDNS+OO8zm+mEHRKqxgC09
XG1h9HROnP+Szi4ZVijUQRdrfSx7pzWpicueg4kRQ6RIPF2pIAm7adA+ZB8FxNYmRbzjHLrV+5kq
kD35Y72+xCQbwQwMW6Si/c+Xbrstb/74XtC4znGcJcFUDboiCRUmOTCT1WB1d4ECfKy3OUA6dwg0
QxUA9prYIU699X0wSWaI5+NImRtlc70TjLZGikw5x3iw6RTYZsfXGiXPxcVlL34MlU3U3D9wjsrp
rQv6Zv4s855wqKCcfHOYS/lQwsQb9p+erx3WoUfZ6klTOrZ3bNSJwAAQSeb1uh3fP2xbMYuxA5xi
QfbwahFLye7v6in4E6abTWB4KigunTN2MK+BQnUJQC2SzY+P7i2r8+yMjEQkX/+PWHkVCck3NjUV
kCsuAUoPYZNlryhYO0noElkuD8aa2AE9uPsNFz4D0MvXnwwI11+N0UWbpdIacUWTWRXMhvWwv4ZF
EzgAfd181vT+wlFO3NEpUTBuDLatjjFBh0Oa+dFmAEUFEQNLTklUNg1tPSwUemvQSlq39gt1siIH
HmoyvCi7OIrM2KAFgk2xVDq8iA6MuDuJUFvCIpmk9IeCCEraiJQr0HWTWCZREzsbMwK87JZMCpjg
gcJPmiztJBpBIKfS81cF8uG8pOP+Ce15BXB4ooDh/KijSAE1Z/qrY6zQzZjwCeAPSU2F/Dbu4v5f
gz2nfyKiT64QLX3btRvPZJnC4ZsJbhvSaV5pFSEj7kSBVaJ+Lhbchs6L79F+80umBI2RuyDhxyEg
KqOwEwnTqsCcSxGiXYUox0hhDK4UXRDYjgYLS3D9wOWs/yeXSMcd3nqffCB3QSeVJVOLkQ9oYioN
pkh9Ccgy7nrDZKmaKRUBnNTojpS1A7uEaujK1z/gd0pNa2ZX8Sn9BVbaSn0Z3SkADiUjaElgHCQs
ufUP5DRMeg5+u/MJdc1XGaI802UylgMXL/Vi/WVWfon+/v1c6+mroJ/NHOQoLju3Il4nTqsNWJ0z
3aMfWtmGHADxhuNwEsVpt/3CZ8rmZKN1lC3UBeZVzNQfozwPz4ZESL4HYADjBvnlw0wep9QGmG/H
KaLFhd9UWmDZbsgysgnuA3a6k5L5vFfwZqc431exobf3flWKZxBN9A9ch4cjAHoJhfpSwFYXWSR+
Kq1EGi2RcTBbOgUNHUCJsnFdtnZNYb5OqaJ1cLYX0Q3QJndo18ImxidR4El87cIV9KR3X03y2AE4
2YzbLnBNhWDLTwNJaf3rVXJE2mku8T4zE2wj5B/PnZ5rrZEDdQPy/AX8BYGCQ81OW52xHayX7ORN
qnHJN2QIjWyM2eks8VJ19jYBwEzUENnk5VC/+SLC2wZYyKYGVwB+7WbTO1z/H33pqxzmvh39gt8K
xwo6r1CB0ZPr6S7Puw52t3ZQfhe9B8x1feGFVCqQVf+7lYc7ePansZnh8kbtuVW0qL89ObzCFwIx
ZsLb9ePzfjRJZKvSno02v9rGwnYEqVpc98G8vwuAJclz7BJO9uBqt1/1I24OPNyak/qxgfqJeS0n
uI0k6gqCX+PrZwBA5BJsX9PklON9eopeR69XsrwU9Itb14ZZC7vL0jDZoFd4r8dApMLcTV+4p80b
qHRdnNNohzip7db7DEMKBqUqmVNEzCW3fObzcYQDLozNNiAohJtMiGDhJV8E98u2jaaycsjBXeE7
loswGBPXsQk8owqohKcTM9Uv3QTWvLbE9vRVYcPB/NFupDBguA8M1pYL+JXRppPa2MHwXZIQX5FS
dTrmHshrLUI+958jgqfyHmw1d1rfxPbUpzOeuhr2mrRTCJ0meWImEdMvjCJZh4zzR7WaMz17CU1e
nNvBNMzt/3znc8Rf7o0d0uRyM1L1Vzq9KwoN3XaKAaOcOzdIiMPbDtR/TarWsEQBPCdyJOtwCb73
knsVNI5Dw33PA6U28fi7UB2T2ZlBPaC50Cbg1TxnuZ+3e8IcUlX3DnaT09CACdhSCIEEM4qS5md+
nH1O1zXJ022mA8RjI/sXjp3Tghcpir2B4GBnNNAHS7GlsATsT9K73VwVJ1w+e/XFL/gQbRzPorkq
IBEV5dpDEBCJGSdpw/oXldN+DmN++TMTPA/TohlBgi+tBPJP5GzRG+FVsXyZ6iXNBcM0o59ENq+G
S+/oFhjjqLaIjrxHF1qWxBIlXEwTP1KxCnBfzjtmyYwg79IPUL9Q9fT0Gu4J+znlanoS5gvCYhnB
6B2l5W3GRgze2j7gjX0vU7flhfmgvacOUb1X1nLYGgE2nfycL3EDr2wWbygBM/VKLQHVbuIrEKZm
cFJdHhtnYYFPXES/e88REANXSLlJjRs0OGcV7KqA3bXae/xtS0znQRWFBi+oVcfwpqoIkX7ou4o1
gMGQjnVCVMgke38rKkU17AlshnkwB6ZYzNgXvNqRUzrSzK+6jB4Mvnv5D04mG9XntGckJVDxtAK5
hOcvnQlf9Bp6ZnhrK7nr/T3keQotYmtuufhXmo/U2h+AYqstyc8uEXGRutgIEVKSl+adpqYegL4i
KO3LCKz1qjIXeZwmHRwStPo5CMF8VDbjgrczdb7O/Aodqh92vg7LqjH7b4UJbA1Ln0Db9TXpNx0z
Hr6kHRFPkTHBSrE9hlHP7s9EiK9L2eNbXpGeJF0tAqEB+82R0OqAVLGo6/k8Mvm74rnDEoHomLE9
MtJyXatA1DdTApoLY8AgOjo8+Fc5WJ6MJRYMWAa8yQ3CuRLzqXTPHgN8QL0hVMxuY9DEy+58U76E
3HIhduu5FQ5sbFyYcf7eHRidkSjxrW4bpgsywwUAgZZvX8YR44aY+iMkpFKHDRZ3GfIgebyL3w7N
ik/mwPgnLqMGA7oSyU0ZWzi7UXvp65koYp3Oo38zGtf1ZPzEUb6+lR0THD1UwayL9v39lmNTvIf1
D72dTQVFx96cy5dJZxnzo7gdN0fA031lIzEi3PhXz/pAmwrwVTVw4mnazT++vFoCxpBR9tHcB73a
CxEa+Z7bi6Tr3uwciXNmwuNPjI1nDnjoCeF0D895UUtGxa0/Ve+CJTMzoi0gtgtp5QxWRsvParU9
rpgWXFnvJ+EFBaiY4EYFvJVcIrVx+ISnFwmIPabtqQ+xjtk5sxuQjPHsrkx2JEMTvZ3vd+S8kf5t
qv5sNTFRSw72/zHhYJZn0bnEs4RcPobETEKQefk952QIEbWu3kQERGEudeQq8PAGinULUNE4c5Nb
0tYBXk/GgbIfyLEDQsmXvIkEoWRi0NChIL6HxFfaxaaNmZ0oIRqY8iwnmn6jPak1/PrYu4IOALPG
keYRZSpob/2j1D7bS6H8U63vEM30cTMhvi9HjQKo67EpmDAva3Gh3mWjfKfYAi8jQ7CSI9iKRcMY
JUheX3cKNiYjlBIJcLXkYxNY/VhC0gHC2SPmWA1ohO7LFJ0vdOSeEubCwYwZG7FmlMcOL1V95g/p
BCzeYKqySFmSCa187iwHLL9D6j4wtbcBj+NJhgHOZkqKAGb4s7MMdO+Va04NJydJhsJ2xgZiwi7/
UuujHtbYlb9G5FxqahXt6IBsPIGTk424ffSfveVUtKSwNHdTV7UQP3H0F9ss7wxjFQ05FNfPwNtS
1idhboXIal9feoAqsqxv6eIIUeTJLPyodg0QGFObUpD8A2TiLWIyoidDUIYVbwIM1y4Y4cYgkP+j
uwitkYdkQudi/iEaubBgrpVeg5nXd1nCf48X9AGdjrS6zXzow/+k+7a19gN7AsyrpOiPH1SSXeio
LtyqyvOsN9PpLC39dEbJUaQcmb43Shk8XmPKz++LsVxcPNydHPvFpL9c5aGDMDjRfvakqWB6/fUz
FKFE4HxMg7+kJQ7GBgND9yoLHjyMIbn7NQYu0aaen8WKQL2V5fiNHxMix+sGp64pc+UBzuTLbbxo
6Cbbs/AysS9KajUiRqSEishbszXmgi+ZkosDXx5BWgvSSnTIIhmRFdKirVG53jcdjYYrEVwXHAVM
0HHIRl4xdq4eB3xWOq6rUhiWj8pgLZJrZGglDdA/90fsx+E+q735MsM+1J15kdmUkFbkpMmCsL5O
/OBpMczeViDEIlImpodegGJ74mdc7ncUXGiaE78z/dQdWgHsIKuYIubQL16qDp8WC2w0wbEagDQw
7hGSeq6GDC1uLT6KoNxONzjz2jb36Lth/pZ380ZWqz8a5IIFbZkxlDmax4HPHRFbBUxdVlnWqVqo
h/3qxNyHlB4yiRQJFMI/zFgNMgZc3FpfMl/5oScy1iJy+w0eqjHJyYEIvPqpenHjvZ85bLMSC4Mo
eY22/wKe53GWsecBpXMRhj0gfyj5sRR2C/YAZ+VrERG6Nhm2lrCbJXp2v6yVIXjv0N0eetCuFK8l
SEPWqiHLbFHnG68h4lq/arvCGk9DwsjHQg6jvHumcaU6Q1beADVBYHTmBx5m0Z097H6O27TA8+C9
yDtubG/AlFWHxx6P8xh3Vi779G+u2zalqF4mxAv+3dZZeC4RD2aPeFIfqlibDJIKNIcvka9gVryb
lkpHlpTJ2+m/lnjvCtmTw/uqo1VF0IV3qe8eB6Eh3MlfQZ8WAqbXLbrB7THaRKaHOKiSfKkAX2Si
5KfHDzud6ppoQNfb7IrEAurIZw5m8McSiiypAX5MpbabPfiY6wSZTA2L4j9IicvPTGeSoPTIQ1Mh
JCj7Hj82ryyOBYEAxJH4YqpOr5Jyge5mHYJkTBbHtm6zVJJL6iReqxoWtMtU9FrJKjOBVNr+2J9F
9sG+RFjzXQeRyR4A7j+oJyP2H6KbCx2GGwMFv0BASYJI0TQeZw2jzP1s+7OH4nJyTXcITH2l0f0J
kMAH9LDdel4IQn7eBbLXKVQmSuSgt1WKEJCQyM9LDg7yOR7RJaBAA/mahENbnaw5lsH1pMgITksX
CyxlU0GoaVU4qB+f+V32qoMKy5U1zFz4ljP3vZQNs4tZkoGVdSSzzk2TUzL/QfLpR7wEgVzUuVR5
5DB33S/aalVO+ZxTVJ47443k02tNZ6DGchG3tECS4LQYYG0/Z3GwxWOJ4uVwAvwm3UWePowyhLbR
rfuCE0AtIlbKdJndtE8fj9euNGAxR8vz0g8stV5AVN3Q07BFRMXa9FCt/aLAsDYuAE3CUCM9FwLc
twXVI17HJB9qS8WMWRXHzHeMpRMHz1m/pIafJSCCnyI36rSJvo1iCeE0mWyI5OvR5+JSVKBsyU/I
/tQadR710V14pOyeHEsPbjyA4w33uvnkwFAC2fGoeX4zSdS+matzuoEjHXHG6Dq6e2h7yp7JChg4
UBHY1nRQTtndXTKPHLTqPLaK6ojHqrLZp6O8JkOa6qzO6dRvgQWrkXV9KUrtGa8qfFUuHqCbcYZB
3r+79Y5iaBUDqt6rJHij+2RlqUCkl3w12G9HhsZb3eluTQ3i+mQne644SMhATGD0pZTPh+Wf9GQp
Ei6heOKder1nyWcvi7biUK5n5PYhhUqOugaG11twr7AtUYTMvv3xalhgmhZfrRdUaKOn48ziKOjz
zzFQzblmIHdyRJm3V6L9mHvsYK6NzlNQ/jIEdnzqsgm5WWV5TK4alrxXd6T3ghFInLmHRMQi8T7i
GBcT7ZBZx5l7ZFDV/Cjd79ir4H5MM21kSGF2e0aUfdMS+Uj2T6V6botDMMIOwv0QROjLOb8AKwZT
hDVfbU6KLtBPBjE0mJjp4JTPK+vBTce7K4Jz2H8HkDidWZqlo348dSaKJwpkm1v58iQiUfbm6VLm
9p//tE1eCJUxW0EiX+aa/lmqvZrIMtI38tz5LuXVw8hMjKauVH8N+m7K1GD8mPerNXKhH2SbLq4H
7/TBBJmOyWmuYYWZOoeXFg+NGoRTI3oB5Fbn22ok/IRv8bgo+9I7enyB3UrMSkHJLTPpLoFhzCwI
P5BpL8YvNsZO/3tWqGz6uN7hGErAynVQsGVDL7tXPP0omB8qsfLgyJNuipggy4y+1MiKod2Ppzds
JFtKLFyJzkX3t1XDd5H7CrNCtngmAaFqXztruemkAFgVtkCulMg1OUtDKK35+lNgmD3sZ4edP5GL
OzWrrTX2brLIAM3ObYLEGEDtNAYuVmagBvOYmVMNOTxzO40B03DklCB73TTEmvgHp779HdoR1XJG
rFry6jxOEgE/A7q5S4Wx2sR95eOMEw8/jFPN89Uo9D6WGvTWSRrsiPlQeT5/gWCP2GV3S5E39Mju
qh7rl/+GzLE6AxZH4zs/M7rjNgDrxSTEr75Ef0JVqeGTxqayfdqkVyPfci/fsxq5RC8bzgZX+/pa
0m/C9t271HO5zRpW3XakLr+OOLSarburI3l8t0E8q0ZIJMBeKgqWeXrSiESgjr5qb6bAmnOqM56+
bjK9XFVjYU0jDkkhBT+DY52GF7jugxaEWokwJe8nL9nSaXN7YHNXAzUtb9v+LqzpaqdUrLTfeZjH
2MrF5kpSziRxbnIkFWZQC3ZJb6y/Ep8frpRdnCyKYVwoqA3Pivwb24h42bv0WujbVTOmsD2Od1dx
SwDFfFcpEFGBEmvQyjEjEJFe1IF/tjQsAsK9lDUO7WfhARizY7BdUCRh3QrT/I6+Kopg64wB7V9P
GnruxEUQWBwBDFFuztsCNb1dbbuuiBfp2svY8Ka6wMR7KuuAX1TACiclEt1P+yDdSD/fiGTLqXMb
ePatwOut834vzrmAWRFOiGyQ2DlCa1/L2X5sWN8E+F2rgsabDmyX8yN8W75LJC4GkS0SGSY38yZn
6Sc8/BX3dVyrbNiHKwRSpxurl5GkcXNAT/u7Xs9kAbg4nV37ESC4UiGNbqcMacezw8jwX69uPDiB
OYkVQJMi+YjyPdY8y3blZhp3VZZzWipGKLBTALGUsnXnp6MDjBJOQYfMAdSEjhk4fNKGFtJlH5cj
qZzdm0Nsw/LfJQUTwUqtP4VrL3vUgavNyLXeYX+LSPgcsN4BxUl0HSMMaH9Ht+p7GpT5/qvs6r86
D3F0DY4OXLkIdlgBoBdxsKdXODr9XPwf1akjh48WJg4pqxitkW/wLNb1tnr2vXxRYgqYUv1nwkLC
1rlPp2Ihf89qxVsalOb8W5CY7wt7ADAo9QvIHp3zSlj66QcCMYROjNSincFcqy3JNOHENBjYguYh
mJXi8DCIMXKyN92lzn0OR4rcCdOgkuQJzmxAzwfVOwPjBpVheZxnontfJsPCIihhyPdo/gleyq5e
0aHFSZPLkyQjxpsNACBcbK2vdBdwNcN2K8F1IECf8EhZYgFkxQsvQtdnqdLBKvKgi1N6XZjGMrhz
fNpT3Pag1EFqQGSUdiTt08HMd6jHRdTSTiADiO44cU1c3tVvRyuErXLZBcJTvO9cqu1zEypjQNGP
gDtV3xaj+CagRhvHta0qYTMUDONuzoM4SFhNNnG5OfVJfeCiJ6iUb/VtI9DqCi8JfRKu9oijrgUx
g/Nk5yVHh458FRRpkscaFHpuycVB6cxZAPGF8nTUf+nKW7rjOww/8ezXqQ8eO55O2pqcKyw8oILa
JD7AAeLPtt4Mfg8Cts2ksdUxHqI0Bq7dwu0FobjMN6Ue4gBXP4X8yGt5Ae7qopVq6sLxVbsoCpLc
1h/ggxiwwMweq7foaYaC22VcYsHHGj4RaNOTm3KyVp22u7t2RWTlWbIAIcWfr7QDB8bx5Cn6fkY8
7AuV38WJc6YBTCM/WzF0l+MkNMljcP4HZfUHoN2NP2RzQZkPAnhw4EkXUD/Y+6upyXO1EZovDzIO
+0BHNIZevUHrTC/ZvWK3kyxfGfQTnhN48LCHY4O+lje5FBOy9c0FHV5Hd0TH6q8NS3XuFED4FUSj
3KVjXblwmX8xpW9dHj7jVVnIS5OckS087NF3nSKZTVxjAOFnk+eRWy7b9UCVRcUKj1fiYOn7lRhh
2nGpTPKGKQ+ygcvsyUNonD+B8CSQ73vIfoWxRziLRRL0pHnSoGhnWomjyXWX2VAg7I7zOgjzhDSB
NMk78sRTkIaQgqQas67wHhc7mrBlziG0O987inNM++MFudW7KBHgg1/H3ANyoi/If7CaBkB4Y/lX
xcd4BCDIvap2c0I6Q07WY0T75E+apCl65qpCszO5PL0gOs5xSd1/u8oVhQKAgWUBaQtAPRdEF+FB
mIfZUi3nXGo4KPCvw5ZvBcK+QiFj4pbHVG/WpnPNX9/davsRMuUm6332sCf7dg0dwyaxmpx2KgoZ
uhn+TPfobPrYzasAxW1yt1TquNrseDYjLKxkVIeHsW6ntiy3J3cNm71SgbtjjP9mykrDGHKA4P1C
QOu5uAyhv1sTE0G1zS7e4e4OupfYJh1OxT9PbXKosojfuWfHk2ks9bJPMaLCBF7NBAjUEFAm5UCB
Xxclw0kF9UhG2OATkrAnYGwi/9FxcIQWPFIp1PYm+OOfd3i6zU66A4h6FRCOBtHCPXAQpurwmZJJ
izVjKncdPlIV3V9zFm5mTqR3cSz7HAIdLN7w/5q1RE9Kd1G7NanKiLfugHbuID02rdQRT/BoBZw+
Ghn7bKIjTKQ+DS0ztnSTBnqkpvKSfDE7+/68H9jUqFrBW0Iw8sQ0pukptdgFr37KdY47Fbk9FkTJ
llksP21bVwHYgAFkB9q5ACv4/7LKj1mgec4Ts7vfWFbyE6YUuchFeIvTp8LA/cb10UNw3dE/ZvRn
D0KVl4NUaTbwGdbUbujGT2lhvQ44pe84qDz2ZvCYRPeKClrfCanG8iyO6ZQU1H3oj4I78VAZpPh0
uLe/wegwMulxyNODJo48VdcojcIJHrMWz08Qo+Akj8ZC8a56tSkUufsf8C2estdhIEu+SEZLatbK
O5vE9UuO+exL6r3gWAI9EWZUzTVQSLUmYqbZbvVEWwGsfO7CPmTV6SfEZzzQEmgQUbrkBMbo8LlF
yYNV2exlgqX+xXAjQw/zIddBcOGI2iaLZy3hc/WxsAjHwTNRY3PxbUqF9SmYLWxKCt86wyBpDJAr
C5BXie7TTethV3H58jeZOqcuQAOR5nggBWnsjWV7cL/xzS3Bsa1UIbWv7V/zI+2XxrVv04Zzk49v
8ypbHyxoLKsUdRtiiShL6YuHQkqoV+BxvrdtOtA9YJRlbMfHJ4bEYc08GesLr2A5p1rbJOtBATZ2
ZRV9yF9B5YyIOVZmJfKr1Nh2xbbdWVuifDTMZcOpzSTQ6AFevb+bnSIU30dIsKzbsOG6rDwISBpK
Y93yJ+GFE070pnF/+wZd3wZmcKFftZiALdmfuGpZRjqrKgXxIiOF7UZWnm/iGsOrazjV4AHPsYFe
NzozI84MrC3dwfBRA16m1BoMXxmAdUuhdHALprAHEuFVEoMLe0j0YGHB71knRWYwh8UEx0ytIkm2
dd91R6OiC4twPUoXiagzBvn4ybrKBx9wYybZMYNvkCpilbL7HPLmkxL+97T/vb+/4fsEVzJeLkL6
LZFJXStAXNxhZgG3JCbcMEjN9u8Vu8Wht0wVCmQUzbyVNYl6Lo+7EYiodRhXGH5dKqX+LLqdfRl6
3FIAvgylBowAWSZfh7T2GbmptUNqLGJ4+FGBYtYoHx1HHWKjbyZmYrDKas4shriz7SoOmQ6ks7Zw
U53ZrHisJwYJcvK5kiW4aMMsUqZ+YSldVyZTVXDNZ7BJ26ymFT1LuI27BEkJe03neRLip8OdQjwQ
tuVTh+6HVuOdcAbDmSUubtR8C3rpyt/yzzYsjcP7tDOvOGaiSLX8bv973J1oMQVCgxzKvfdCusYt
Rxl8wGD0mD10YfdpUaa9Z4yBR0XFAS34kVyoCoZcdMwRtaYFgnZyjzmHNOJjzbrXCnhvGa7F09kQ
oZVYAaxaumfPKfLR+Lb38Q4kZ8ZCb05ORMcZP75OJKksonz8YL8l/nOaWmD0QnrdB3r9ac6lXd5q
eCqc+ilunnmMy7cm8kpRYGlzz6VV5eeoMG1hsU8sCpNf2rBL5BvuNDt8HZigS4wAVI87nr1CmllS
5kUQNeV8v3WkIEYBia9RyF5ucZtqou9dkjSF+f7+b4g53n3eV4vvw9uF2XFQ1xpvjlykRdK7xJ4R
x6XbdRSPKxQCoNPX8qyE79juAUKsA4+qiLj8PzXSHiPfVEM+ajebYZg5bTDZPozdT0+iq3d/WUJr
5t0vG0ttjzdHDegayS5YlYqHOemtRCRnJon7/IOTXpxeCVw2mjaJaTsuI//NDhU1OyyYWGXwSgvW
6XbquTq0kZQBzHqWI9h+c3vsQOVrQKhmcYZq7zBAZ8vSw0S8paeHIYEzok1NW3FoDXtz4nqowxbq
keGDQsSMt7hEjRRUq/rCYMWkyJI3hQUBgB31NWWOD+eyM/YFgmafH9fMTzhsOUTEViiVPjqTRibm
qMyJIgOpxV3T8iuzQnkSRLqq1OCGIUxpDENq/UMpYjb3VlihuuIkh7iUZGk6yj749fBRD1lyYWPD
wwCqk71UHH4NJJbtSHvS4gDJE4MiV0N/wIJU4wyonoIusay5KB2Sj2y4P6X4+bSb9j3rsEDc1wkG
P4rSfy3mE/3mhxZoy9Wy+j9cUJkI+1G9mHwM3DxcOQzJRS4UYE0TS9S0vaEbMRHXw+1+b3t0j2Q8
Mv2vzsjE8Rhtd9U7yWbprUy1cnp22nEsq7BMbjpDztr22OC6QvFRoNAKnkE4JalLrj6yBWZGCq04
dACFprDirgUViVbXHC0AYySnNNKLJEIS3SzIcFLqIyE8/OtfDc0xa/CXvgCMowv8TMqjKvfSLko5
W2VWk0WW034QMZBaRhQ+2QnIc120PT52XRlRgqipJFx7NkIoLgb/9KqKRIw3CB5+EPD5EXn1Ws+W
xQK+lTQUTYZwA4gdvxEX5zXFtPNOA+V/b0qdg4+PLYpuZYWhigrKunKtPcANV4i7Uc3KzQB/1mRu
PzmVQdnU96pNrqBJLN9n7ccKNCI6C5LFY9WQjyNxqT3ioAHnkJrZ1J18GJBairUT8luCDzMTPnt7
f6MqsVMvRBfrfTaY2weJErzvYUcIxU9t2BciQGdogSuYe5Wm83YAv4tg0xEscdldLgwNsQfD/MCP
ZPR/KkY8iRdsd2HW2OY/Kyh2AACb+2HBneUFlgZolPnblIchDRGsT48dUsPq9VyPf6Lv3AbHthfB
CY4mcK4OAp2RJs/5rIXMvP2PrZ2I9hxnxkEStp5vT04lFMqrzTqehiTEnS7Popcch143RKJgL15M
TixmXVpH8Y4VkmcLcFBm4dMK9+FUIf46096ncKb4PC8zjYWQUdZ12Ta11ckOdhmVVi8we2ACWKrl
cHlYZLPMk4NP7tnPUhp+hfp0AsXKQqHvp0UcntooeU7aGoDgOSPteyyxewI4nWJkY/UM/ktzB01G
azPheC/ud+ms6hXYHLH/YyxoxgpoH8DaMpyEh+/iiaykDh9rJNU5b6mftVcN0QOXpyfjbm6mWm0Z
VD3t91AZTrNAZBsx6FJVkbHm2y/x7EvoKzJVUxExsSBBF1z7PJYM/6e87oV+7kciSRSB4CsVwOpj
g9j/j6nSpuHykNVC2XYHCQteNv9cBaItbq/inE1H6Cfmfa5AcsKEBgMHmNDLv4v56VcqgzSdhrnm
JOr5x0mUFU+X+0sMRgD48O0prUlAKwMDSFKCWNeUHa8H0+WaWwgBOgdFHONsGuz64VWMFiEYv1HL
hx+ZDokNehBL92pphmwyVWiUel+mr88xgT2pMO1pBPc2AqyTiG3vq/pnFzCoe5tjlSiUNAt5bs9m
CJmkEV9Bj8b7i8J1O21IMhasKVbdGInbaEVnccpo4jikVAgpgKKSEZ8zLmx+TV32ne0DBLXHkofV
bbkf4kToWJg66hIezSlwNzt0PaDKoNsSIIB63SuvbSZleYzZ4A8p615NylJEGPFpkWWM31lsdiMz
Mr8l47vPfdxAtHeYUKaq+z/SN6m20yWmF6CnXtGc/nBnyUTbFU/B9SniTwtIJwVgt0Yw6cHwcnwV
xNKSyDSDpe2Nrr3fiLvAvlfWEgCQYmur15rtvafM5v2Nqfe0dGdt4Ho3edQndGdH25SbGljKyFYZ
tZbV7+xAMTzRGsWHuUGU4rpGx7OU1lY3EtO+e+b9Q3DmE7U2hfZrMtNZTPQJBlWzwpgyc4l4/+jF
NaF0FZHIX0qDPGT5LUAIW6AevZxQ01b6AUROeS9LAsuzpKJ1epVmGObH++qjgMZeQenv8od3z4SZ
WaYCqyX2+ao8WdVO7ktYvAjbfLM8a15c7o0vKQ+Jr9/xwypFBFeEnq6pufEYNK552Z3k9eAw6t4P
MS44X2a90qu8YgaENYDUUI0/LAaW86D3mLtSV8WGMcy/R3gfStLsmyAJBTeNmY7aamA90g4aRUGS
+TQCfq/WfDEql6cuVuwJztSaurMoBUPeWmuWtlNS+Ko2tzbDlTbJbzM39EA9o+BV58pR0RbCu35f
mLRlkM1FovAnvDXVtep872gqNo6YYoQjBab+5q9DKuAiHLWR3mrSvK+JkImoeG1q+X1WMc8qNPmN
P2YIQSNLpOIrlexybWMM8M1tRkP+U4npGkP800K4MqN11JkMZSfsEUliIrfU+PAFBtAMCWb+mmVP
3qM5A4xvnFyxHCDI0jozm3eeQWF4HIcBzcjAqxiUFwGdTSI1hVhrifqrNaqYNNMNxHQfvDvvUYwF
VOYHEzeeVCpHKvLPVrYjRlw8rdDegKgcOoyWHMoq42z7ekPkgyfLklRDlvYmE3ceSXnHRSxrt9v2
SeFZH0jA42u+UDk4qptapNBa6d9LbZsP/ouGWH6PG4Bzhz/cpn4vudiE/OjxKwaacZqniWgv//y0
Ee5GCnkvpKCYc8wFgtRnBhqQhb8I8EJl1kbJhYp/xdG819suISuGZtXta7PuTDjiELtE7dUQWsLa
pOQpQu80I2jOJNQ6pex+ZtVuKCbQle2qifTScmDu8g1RUBkzg45nRula5vruy4wHdgNf3Mmwfwc3
aSQ+10Kia/MCw055orlnL4tuhtwmARQi+zf/4rHl++ykWpRurAmzYABPSYt+a1HuUP8qc4g6i3or
uYHQ74uGC/kNpukNnVJjFOuSJXzBGWGL5lFAhoyWBeqmkKW0q8/PjYZHYMcbWKv2JNiWTHAiSw8k
70JgKC+65M9K+XTgEsYGa9fTqQvJlBzVCEP7UFNt6R29eUX4IXLH4F7viaj1NN1a3dDGWMG5m1up
smWYI3HbWdL9O5LCuydwMp1GuBq5/oQNXg+dTB+pp5eKS6duE3IqLyDO8Med48zMLwlF7ZNAZ8pC
gvsdQli4v7IdEpolmhjpxReCnxmNfuCdRrIKeoe5Ay3wyZjMq0etMn+bTuXkdPjLaxoeUAiLonQH
MdseifdRQcGPoUD97tX9P9v90xatjfoa8XfPLsox+YzPehWMt62zsT3arX6+RiPiEwg+UNy8iYKk
Uoa1g76CpI1OywkOXyJWq5mWO5TSVc/H8VGjdLLeKvxxa2Wj30/njwMItdWSL0v9WEyWTv4Opl+z
u1Cj1VB/EfLAN2abhl6EoxptQnal3EtSxLbOzyDmYq9FLDiOJViswQMbz0rITMgoWO1Hbsv9J1sa
cixnFBkTSWke1/V7I9+EOYZBhn+RP0oyFJ9RHhvS0nBKukZZAioatfQX6X1/h7nXY4nTJoVVtkTG
eeNVqoy4q42yAmwHBYYfARzUrOpFzv68dExGsaEWPfRzusXsLU9iFX32WYLr+ZbNJAFSLsJwYbc3
GVHOMk9mlu9Cw8PLDM//t8ypJ9BNvlgXWU8cnR9F7/EeW/rBCg7JDIyPyImISsZaKXCIwVuOAH57
kHtJLfFGCg5366ziKEWhe/vZxPjH4JDZ+to7lN8dBMujMiC8czXwu/3buPe/wPIrZ+SkgVz+AEea
PaTrajjPhKdUXq5jh4Xc4V6C0bV71dvAFtJd8tcfhbiuyepZ4sfsefR5CPH9dfAcxFaO3jP5xVLZ
0IXEDgmflsi6sdCoueoouRqYS4LcCX3muXdcz1RC7rxw0ohnA+AnefTdjtJdK0y5MLfaiETpcjor
n9CvWS4D7k9XTUL4craDnP738yTPnYCDhKjBy0lvGql6AeCHDueos7qtwVqHOoRiqm6tgoe5i5Aj
93/6Alh3rAFwTN3nAEVVcjETxCAU6oqgPMFQC1E2JTxmKQPAkLHKnVd4oQZOGv2jqvgic5vLaJIk
vHXuPelmg6dmPbznEagRNhabMxP3/gFyQrzxrPE43OQ1t7449acEjHU4Vt3zk+CL7eD0Fej1tMCo
Y2l6GkC1Qua0Q3KcdXA42z1+fAQg7RK7mzlLfW3wH5hxN7OuFH28I9PY0grBoX9+em2Dtn1JBGib
7q94p2x+p4AC9ZtdCTzHa4EEyVTpsjcfVpTAWoTD2aoCAc+o8RVPCNotb36NuQJMk09LiVlVe5G1
35MugESAV4/lc5SDQHH5B9yKM9qKllc3Q5PSc2D0zR2md9E3zp91V4ZaGw4F3zUtIMh9ZQ5ah0MA
XOjhhMobJuigiAUOMwHG0V/Fh4/2Wgd3qX7vBlKKpsaWF7tfSJDUWSUl2UICC1r1R+9IGpOCnNQL
KCXyaVPkpBuVW69bsw4o7NtEcVveC2PPQHhW7EseuU33w2tc5pmrlULfDnSHCRrgsrZrLQfeaSn7
WDS5OnH4Yfiw5PJ2w+CCbVkegaFSwSxaJcaP6m8xoxQVrHW89JWRCnXsgDqPdDcyeyoXLrPMo+sO
ZiP58UdhjxPSBUPYMVt8qh81uCRaLY11fwjntgplcAfhYOBuGQm76hdsmQ0eJJKzLWtHaGEOpsVh
jk4ltciZzPQbJbMDYVec1gFkrzWcrsWjvvcUHUvJlkpSSDfkLi/dI7OT2AkmUQG804vWLbh8mJy1
iFfiaR1qHgbAlU3E+rePLAdD0IiV9Ha/9ahtqWgU4oaQnXv/esAAvGyudtSG2M5qdd+tFY7oG09W
9BjUSjFnv0mH24UZ/w0kYQixc54FEOOrNDIxThl4LACSRNJixSRORzBVaVkKYc+NfRcWYDY32zOB
58XtrbyKoa+pYtd8moegWr9Snw7eHo2cQaxb6DAZ7+Zo4XqDlYpo9uH7EcLfDBHUgqGpudITehCD
R5cRoCUKhYFr7shlYbzsR9Fpy0YxYsYtzv34+hskuOaGHLZrotTnWm2vQd+5yWjncJP/NezHV5xw
rhkzvIEboMWce1JSsi5VLJZv9xAvCaOBHX8gNRGnxzGfpUY38zGBJ1KmrqQ1x6bt09b69dTKdjEM
vbjMLbiobQAsi66+RX3UuVaelEafLLr5+B4sIoMCkYBVfdn5ZymSq4rDLKj7BFtcKFFqtEo37qg5
dhY1s2rkLQrJqK4luCmgksWfPLgWsLDYUuUgqsJm7i04pJ7+p+ZdDAlrdbsmAnvvZ9hZ3yVhPpLD
a3fvRUR7LFzqardwmifY7QHQWJIJ3Bef+0G6v7xxK0+BWfxVm1F+oQtuDPdanUMJyIHgKu2IVMtY
cCQZoAP513gITPOhsD/z10mMWRk2N8V1MG6QIIKmsVhSWZEYDh9oGlPVEgpX8Met3ZbKNtUEJDr5
LXkw7Naq/zvCcvHAa0KfVj7AwEawSJ9p06tt2TUZ8IrBDGa1OKylvcIWnKOxJR/y67tX3M10yYrq
uLYaRNc16JgRKBV7suGM1wTU8ujgeQo2VKz22rcTpEHvLu0WJIVIFfOgSRi2lxy03PWSYpDRp+/S
5BGsapLnPWVfDHNM5Ll6qPYAr0l5uVGonsLRTLFd3OliUXqAOLvb+0F9h5GF011GGqTQDATMLak7
ZCvqzQq8XzL7/stNFZgtLPSYmLjxAxhCKF4toviKWwn2OcKm/dNG1cCbisfJkqpTyqzSO4w5ipD2
w/NM0Atkg/2Dqw7M5uEIsyq0Zb6tmmVcp2oah1IyW5WGe4eJ0/lZ9hOLegjFvhivweWDdge760HR
rpvrs5QxwYwzQztbFn8G0eaalN1Zhf/8HQOQ9oKXXjBOMKYhBZ+1pLzjrtrm2t4sYFUdliHjf4cb
vD4b+1ycnAo/gGYC5lX6Qn49cpOPZW8U2l4Ury4HtMRPoXm9ZK0HX4gczuIqYFeF72BLTV+fUOaV
r01F5lLA9GUImlrZazSa1TnsOHE3Ue6iHLC6NfY7ywIvtgFkCKuSvNuWrkpNHpSkprEvTy6wI11X
3YNp1BKHjXaIRkVXSnYwPNS1nrkdIZUa3/LvXGQ/3LcucKGGL2yp47QAKRNcfTQU0mkyklealmJB
TYzTyyfng62n7TJTlRBLNcp8boIJmIFgmrV2gCSxKa7oO+ffCFeVE4bD11J7kJiuWvZnAJeY1TO8
fmYIhKmGVjwUxnHOUkvqC0qF40w6xy+g+tDS8/8l5HrfQol6lCrgAFyXxONpTDlHUcUSINPgOaf+
6BT5HScsPN/Ka50uF+BNqY5wI19ggbtwJz7eSrCye9csqQejBnTWR5YmF6mu7aDyTGXS04X8xSwF
gC6lJcbFjkBKN0wmTaFOSiyyGrbbMpjUENqU2C+qnA7gQe23fNi0fHBG9SSABjULb/KOh4luzp4V
czpKaIfrbPFEgLmtzxYGDcJMAf771VrQ2dRSqPfZ2VRHJonEdNk0t3w1s/qvYAOC+WQ+Ip7S+KJ1
6HEWW7wJtgMJ9lqvyULUGjjcIrd2cO+xGgUOu5PiPcnk4RnKW2GF1EiPaldlX3vqMZRNxBpOfuWy
R3yg1i2EN2HNEC0ZGvUTO5fJPEIO8KQvKna+WKGBGn62HpUG4aLtWnBEhfoZPlyKEHyiO28T7AHz
amghdkIrkazIj6mlrqMW7PTM1ZS6piB22WM7kbFVAbDgJkqZ92KQtS637T/J8axPk/VheMmdWDsC
MkHHhUpMaTBrE7vsuwDx8/s+9xW0VA+DBL9UdbEC14Aezj3WoOTCxRjnZiTMBMNd29Tah2Qb5rLa
0qU9o9lbKtoMh8skNT5GHhKI1ts9GpgZ9ek/4Y561Z2kcAfk46VdMFaiM0kivH0v4kUUUDyfH9dw
iKqZSAwYHRAwk76f2QzeSyEtgqBL0n2l79o+XB31yI8WnD8bCdrO/GCXVNfY74Jp5QF/SqATXxrL
3qLvDm7kkKgsl4KOMN2icesoY2vyY/LHj8b3pxJhHTbRhMzhgBryMo7Ft0cesHUeS1JmdtCLQpg5
TlbqUojP3StFBk2KiZKyWR0a52oWqZKaVOff6BfGUzFCZl+9nIKLC1PvYbnfc7ZQk+Wof/HFpl9Z
dcES5GOJr7J371BPTpYEvaUkafypuBJvSHy8EFpS8zUzosIuSLxRdoLA3NHkbG8/Us00VpiI9FJ7
NVwSs22GS2Bej/g94UiAFdHqxeQIjfrXOVPOLg+hTpzV5ogcU25Ke2Yae1lxQsyeiS8MKKT//1vX
69x4LFLpmuRbx7vlTdPIvAvxlG5wIgQ4S77DhkjlZVwzFSq8Gb21Hmd3BAweA3KNSf9cGWkFDgHL
UrDFxrxgTAUu7OZinupV41h9mckdSNZT7k6dikEnbLbggcRoLap/Vx4vFJaL9LmjAp1a//Tev0BQ
HVGmn/5lUNog1HZOjwD+9v7e6NPJbVJ9yjoOjqyTWJJQoWfycjqlcRMAbtFJX/kUDBFURrPylHDf
kEMMgq4Y9DHNMUSiEGPcC7gUi7dh2BaRgIRjaHV5gWXEkdjofkMr554iluaSpj+e3N3tm4hMJuAb
3sywEueI+Ie5HSg/d+kQEM0qtufW1yOKKuvt9SvOmtCpDzo1xCcToxOSs31pbzmiuW+qfTeitPmr
vn5DXtch03tNCi91O15BjI2MHfM8GwOlcxUDS3Z7ogIp+SJsyWB5rBDmWlCHDjNP3seA1SH29mlk
7SZbEsqlhyykVNfQ5ozw8wFNkoBmTOVvAZmdwNNVKtQyS5PMi1vSsOsS8labLTKdmZbT7ghPGqMx
rfCAIPfnKPD8vkaoN5R+sS+cVMvyC710GvFvhHyF7hLI7zPqYwZdD35+QmOJGsK/aL+H+8WcUlFp
5IaNTd/WEudKVKVoxW+EBwGHb/jTRAWMC3fJ2q37vlDxP5H5r4E5PTuTJhpOY9diJv/DMTQIlmoH
9mdJrCUAzx9cR25M9FfX4EASlcRS/1Dr58W0jI21mlilHSJM+SdbazKYwJwMIPUxk61QfuwSYBfM
VcKzPOx5Zzs/mk7kfYlOjRpUi+V2AscK9pjETdNdIHho1OPa9UfG4RY85p1cSSJXBc6EIY/nNXlN
iG6rrcfBj9E7q98rnsH8Y9w+LxP8FOKQeYHyoOfVAgOOHJAA4tU8TlQoddud5a3WGAV0iNfMav79
kHMv4Gf6k6GmVFP/a/NS19BndFv1PXvSfIKutBFmMQ085htJTOCxOTem55rCnrkUcxKTjz3uEqHs
3WKqK6RbnYhWTTRPc+bjAGSutUIiToxtDlhWLRl0PlKdteLk0fR3wFb2ewlSALAweBi/a2y+Y4P7
Wl3TaXN/70wY/fnc/fnfFB+9k+yGAxYSf/1NlxeU2sPvxt8S9zW0SLy1kv1z39KNP0+rK/DH3mO+
7YMhbqdoUqu6fWjh0xkg3heOyMcJonSvjs/L89PVEBgKHT9N4pEC07YajhGy2lf/BfEVwPsmm/Xy
OtU9+9+3ghf0bYbr/EEPK4Uq+ZlEPcpgOkBWEeptGfvc8ElDYjAKX4gbDYeon0p99k2iCxBWBn7I
gQwOuozLK+aGo3Z9BWvbPdfkSkw8Za/WgZ4ojeO7htpaS+FTp5sbcyTQaGLMWzgA1EJjT6kiTowB
J713Lf4SgeEj4EXzWTlyWL+kB9t/ACk0nLWTB/3LoEH/WWwH8Sv2X+V699XedaFK1naMd77X8Mwt
r1uvTVXZwD0v2fnv0+vtLXt6prnW/m2RM6kRkDi3pj+rWjCXS+G/aJ7GBX0rgvXn89W2cifHUbo5
52mvwVc3rINfT93pWk3uSXO4W7fGrpeknNlU97lQ38yCM+XNVbftNF3AEvihUmgdrIeCxwB5Oks6
oEaDWW/Zo+WqYTXl3RTCZB/sW6WYCeSsgcklBNdZqP+Idbto/6Wey0DITzDOt7AdfZBfPZpino6v
SnVcyA1IJM90qR+vvXiKd/pDBg0uIJ97I5dUdXxdOJWJRwjX7rk+4RNvA83HW+hT3vmONwWzTv0A
Vyr4X2qc/ZZFmpgswYEOQjKSoBUK8219Y0AfKBatUygW6RHoiwK2SQyB5OXufXQKSPuqj7+k68zO
Rfs2hJMzHlmaCG66MkhFH57g0I+jErVqJoDCmyM/a1mnbpCpaKhwCQKArz3ZIm9RlXrJ7eFaJSif
gMHe5r7/oNKVzJizuP2+m6deMfGkizAdq7Z8FkvJJpsBT0XLv5boMGezjOqVKgfLNhpfQSFp6CZe
88jpbjiup8Pt3XrinBELuh/9fZ6bTfHEuDmdiMzmr1TZpaV3iKCVWkgMXWJM9tHU1r18nDQzoXB4
W00M3Mq0vSGt6lkBQG1WfAS75mFNcs9GkzyxCCjeDt4ZthYfnxDqwz1sd/7B88aCSifrgvYAdd7I
C1l3f20soc7X1kgleP3YjrihtM2XAw4dfwcNPgpobIRsoi3K5ki4MDFhQcoChSrqZv4ca154bSDt
8uTRuq4/NI3tX4lTBymzf9lrSlowLVZDj3YhLg9ei7cpxccmlhXbAeF6SdlGKLEGV4xlgl20uSd9
QQpLptrlh1ATZ49zOcmh5RMH8uHuFU/JICk7T1P3foZlsHf8xb4hAQUsC38l1/9/el3sBGvmpkFb
5o/GB6s1IMyZ3GtqY4xol4GyU9mlaju2hUVSv5jri8euemwaVNT+55gDptEXNGROEKgSYNYCsL0U
nBPG11dWNnBu9FRb0FkklZneianMGpmudr1GvfsjMjuA9U13VlTTdGLjuMMZOcXEbPHrHYG8oXS7
pntpUFBJPbwCvFKh50VeqVa2zMh0Q6LtJ7eKAKIm2QtUSYkm9t8zyGNE8hYVW2xqSzZxRvtr6C07
Q6bYRlcW1QpQrXnziDRyMA2bUlz7TB15SH+cF7NzAyhgWo6T3qnSH7U8aalqcSrY6aHHiIN8qOo8
1Y6wpkRE0HWuLYMulmqk/B6hF4vdG1nnHUFtz4f4hoYHJbOHflwjnDwNrfsDyLTo2LRZ+WNOVIP3
NLzEMxWKwMIXvciJRPb5m1TImPIHRnY2uOj7mMzVdwZ6eh7jPDyIk7nEuTXr/OtjwNOGyuIHAf+6
wDYm9Ma/2knmfcGlamITc5V2OZKmeyQtVaLbWzG4H+uklNS0CQEC2L3Rot82PHXrYC95V/ogR8QF
QQKIZQkT6sGGGkRxQHYadMuujTVh4U+G+CVeFTztRxVn0Nh/mIYr4GC95PP12rHG+sFD9Xl5mJtp
kQ+yo4cWYO6ONTXbm5pSutJzxTzl9B5TGVhRcckMM4vri3JWPcLjWfCWOWg35Zn3QlLXGgOaV98B
0dBxKqNjmd06wjL0peiNE8kEV6IkR8Ztc9fQv2vccpZTUlmMiWfIhHblTh+n7Xs3yuVRVglsfVpg
RYgs+CXmOt9BcAMc6JDLJ9LvRBaIzs0FiXgx/s67LSdTfq1EDkxnTDlMNSG3avS148rbeApXi6BW
0HHso/PFWVizfEqlN3r25T/0RhE2k7OKRcAxPbDhrc+WdTQQ0GnA6BD56lsHV+YsLWWLVUP2FYf9
/v6jauFYftxhrXLTOCFEesIn7EBjxK766O6zwtkdg9dqQlWeEh88uYqcAVx+6Jnn+IR14t4FM8pL
1spICCvWbSpfJVea32bMsPzaGPF98LaL+f2tDsFXXuz2ny7nxDSxTcOsreSRYxef9tGOO8XcoVfM
n9h542DAGK0yV6MYRGWLpKfkw2wsR3q1yRWZqfsEqTyxsCAgq6MVGhKviCElYr6J5qsKprknmvn3
8I1AX+WPsHkAQYB9pP5tZyxrFfZdvtbhTza6R3zBYxvpDdbIHJBBlcCw9vKfQDyTFgSs26e7plNZ
GcR9qDwrOXB3oa/vRJAkoPsKtzLE2rXnR5/9RQ7Ei/PcBoIcf1lZ96f1vGp1+dEKtxNPOdKILgRJ
xwEI9cxnCsZvtgUw1ADlcR+FzqSU12eg+dYOea2pSsQ0nggB6bNNR8zA4bFhYPN5JUV4rCDnxfXD
ohdeVdxvet74heUeK6p4B1BQAxR3+RJNuxExq2tPk55+I+zIOHqeFb1BJutQ3xNHlL9HzHIgUyOV
BehIMB1Xf5lsH8+EMekOVu/BwQmcfrmAqRugdVUSyLDmLwrPpIYwq8YlRox1N6mAewELT0Fu+xUT
tloSK1jgU63oeJcqEwiK2TAlRanYJhBweIVYHMlWJcZuC6ztQ/6LisSYF2juhVuoWecG2HGvDVP9
zuQQzSa5qh418HK1I8q2kcWPeIG/3al8dHjltg8qJs1/Bm+C8/+t++so9lJ7aKNVzPlcDCNeuRkm
HXG/wlJVMM7UMtl66VmZnLG9JyvpKHQLXOX8MoBiWCC3nHb3iT7hTvyucVsUePsWjodq83uEXCJ5
qF6MeYeOqLyflO+JN0HhAhCNY/0ybJyVk1TWb8jq3U6m6A6NRZNSnzcG+hG21Uz+nFUA6ook2O5k
UUYk1rRP+BrR7L0AR4RKT9PDLs56U/qB8ZuzG5awQIZv9iJVy6b3H5OMMHRdzPxlTIAS8dPHTK5S
z+hcfDasKsyPEP9h4++6JcOYJFk8nxpACMUoGGkDTU4Ta47Njt48FA7qraNEf+wZFREU7yZzGUIg
qCBNxrvbagZL5NDNvMftzrAkm9zOCmBrf0ONwNr0nsKP+JDT4mmwgBtkuNm0GwtYbmq+4zln04i8
XmvpqZTj96bo1+qOdZOM0An3ZF1ah5IvkMErW1Py3IawWtPFf2ryBGDRpOxUhTt+tBO7p5f9nhtf
46rSDw81MOhg4AiIWfPJ88wTsg8/rG2JA9qqMsfuKuURmHIT5M3IBWgCxzM64XTl8pLHPGOhvqzm
OCENEHNGgAE5RGlD+QgAdSszfH4ItpQVeuS0+cWZn6gMzI8gG072PjX9Du1L+syKWTina/zJJiKY
M3dZaNtT05rXjdQRwQpxBbjtdEY8qabIej2X06HrXMEb71qyzWS8UgLkiFODyYZm2+UcN5VqgrmY
lfuVg/KLnsSxYYUaI9TSB4IIghN0kQz5TziNC6srDF9pTo/zHvE/78T9Jk4C0u9OCeBdWtz/ZaOA
14QYcosGqqcUdbJx37bG48k2i56JtV7H48v8fNKDe23SitFOgSHG8T28DX8bG41qRJ5b8nKS49ec
C+NiHsbfe+dm/0Xsn2PTrqmJf/UEBJdYHjf8iYL/SxSbQKs3CDsGK9lXWTvMmp8bXHvqEZfmtyCg
HKANwd5AE5C7qtVa8X9KFaBDM+Zm7kBm0BzF7d2SmSPnHhgzvCpRHRjoAwIonFj5digQLOTI4dsH
0Ir4gSMy/sG+sny1d+vE+ZAcf5x7w1t76HhlenMX5HuSj6OA9ByXagQDwD2bAZGI728YReNsewZ0
nCxyPBAT4Q0N5Nt0+15wTt2QfXA2GOrPMjuqQ8AZnjaEPqq7BOfv1V4ByTc+UUICD3nDXNtGoxOm
54Z501wRA1lpxuEUZam6F7qdn61/j9I/5SPcdNA1L4JKeRwEssHmVbZHuCycicNO6UGBp5ybCOSH
gG0S4fRcS2eKcej9OmCpqSUCY8TSMQD7fOHLirsUmKru4YJhDvlW6CYbiuotdYc9Upi5HaFhA/7b
uFzcsuXYc0rh1G6lPLE5PP4f6x1Gy8xrSWpTZ9T9weQxgm9ijqbgjBvQX+GNUDJ2nLLpOlVvbWtJ
PQPxL4t0V/lMvCDFeqZD/WWMGZxJ5AVJpCIKfN/ijOIu5tY+6Mj8I8WHbdUe4ESqYphnfI8ibbVR
vEkyKSmsetM+9vihDZA57SVs+vacfZ4xLvNseber4kNuANaahtdTOC11s8JlTSdMV3DMUhhSfDad
5jAt2R3mxh39W+/FfE+hIuJyvVxMSwyQxcors6SehBKpZuJ+24OmB0LtM0PD2cbSKbX45ZAUAQJT
Bp2gqbJB4So2tt5or9idLj2+uTCOu06vjOxqFPW1Ezgq8Q+cPsYpbNg5MdJm/CcF7PM07sCeKQxm
LAWvyDR4GoUF8NJ2iPTVuqIrURdpZp6KdgRu8UeyirY6HCnKfIf6nt6qpRfOtCS30HNgTUHS5wFA
7v3hqPVXmRp2xFv3jj5+FiCzkYFALPByZ3no4t7S69Il8S1uJSL73qd8G3HK+0RZSRxiAM/pLRlH
uSdwOjwWJ+702dm0qbcUeMkY2CmfAeTyrlKQ6Htw5342YaQKFYRuRF1hsI76Kh3z2R8v0Q3dhod0
88kyOs0mv+jSq2IGc2GgD6kLSdFyTttP8qF4m2mYj8hhCmBITs9/YQN/kiO7qZ0jCrSaCsrZmIM6
1c3jCUVZBm+5Iprn7uUI5/2EDqcFxEhC8fdV0KEaYbl7/BE8+ySZG3kYizNkKLWnejXqe4qRbqQj
8RLe0qxs5RJ6gszdWqL2WS6KUupwo2nTzVRE2+7hhqrUfPjPmuTNsQ/1VEfO/9pnX8inhmW84R+D
jHqj3FNbYO0+yYqfQyCdrOM39aieL3Wn35+S7asDOigKQiG/2lUHe8PqD/5OWpQ47A2HO20UaR3J
UnuDpqiP4KG6lYh30oO63jAHzRSYrYFQQ6lnQnY2y2dX/cLpvSmXVpsBiaWVB73l6UwW/NBV1IHC
GdHNJvDyGmuYRttPOsVNv3JHdiASIY2kbme7G85sRuyT/fARRESRrezpNXn+CYkoE5poZ/YtWgOF
uxBFqfAwIZn0ss9h5aVtF/Vg1sL1YnUSp9A4BZfcYgyT9Xx4WoImEGGfu6KsUE4FIjyn1qn6SOkW
0ZZwpHCA02qwOw3HjlDipxESYqiOVUbn3dfJJurmCCK41lCacwhs/QjjQB8iOxs9E/IRI6Cc7kxL
r+D249wB5JOGRiZ9s0Yin5vXkWAIeKN520K348ahiCYkcWCizv5ZLxrYobMPLlrPx1iK2bjfObE9
adeIUUSCn1x5dbkrjoxO6IRLoXjts37JcseSMEggR+z+5p6bj6dM2WeS50MZZ+MQhvlGfGImgqV1
nCk/4ZfILRfbGUzmuXJaL8OJ7sjQtV7pctpmLFGEVm6UN1i6d5zefPkQLTO4+ph/05Y3B+wsinS5
QCHOejNm7iKEPQ+0iqBdAK23HTloytPVlDkbcMEQYRBqq8GL9voxunge/uG/y0VBR3uivM1WIBm0
Bk/dbjF9DjFi+C54Sth+WSs2Uj/ooWdpGWh0ASxo/5yI5E8NZs01Ie5nQNDQLberQE2oboa8+9YZ
NOcyLRdUtJotXk4GIkewqit2f/uKCVXaGp5Yh4aLZF/tTnh0fz+jsO9Pr/RCefyD2Q8g1MEi2pMk
30zZShTZdjW/ptcf+08/niEmgbBcY9c/1bkRTJCyH3WAWBYVcXYsD78fQuZ7dt2oriLOh13cJHQB
PyH9SLu+uwvXaXc26m2I88BBHwASzxtWKwXT11hcE8e4yv/fh51tCu4j4V3hzFH4hY3DH38HWnoB
8Ag3KbSqSe9SJbvIr3fcp/ijDH70la0QsfX4SM5hTq/oJyLBRh13MUF716mV9DgFQrnpX39zhIm3
2hT0xlPW+ndVvNpb0l77qxN6Qv5RdfHiTrZJMPGWJeJ9jZWtEoPpGykzp6r4o+yYNo8v9/qvboVf
DZRW85mToYTmToiB0eNRdtdglrRW/2r579TKB/LIaQ6lXSDCaqgZybCNCuYoRzs6adJXbHmf+Aqc
EWMmRjKL/Tdqistl1+A/a62UJ+IEz9w1O7UucrR9l5dSW18SQg9I4A7saajSLEaY4X78hylsKrBH
FNDOpB5H046d9JYyId8xybHKt0OrxZmbdTjeDhxzPN+5c/as1ZPcOj5DrLgrHVl2p3tOMGp+iAvj
vqtQKwBE1tOLVAm9Mk59TL54woh907xo6Fe6TVN/etQ57ecSg6V7KQAUZeU2a5ad+x/l4bPizDio
mfZEeq/DSs98CFPUr1Qf2KLc8EQmJBb+8GYKu/Hg5c3You9B1iehFgj8kjes7ZQGw3NNYSUnOLqN
4FdT+CKIGdRr0BzD3DEjVcbs817p6cDH8XddRTtUTsQScVB7HkElK1wAEqRCqXGiK8ery0Z+djxL
yz6UvXLcc/wAtTLAS0CQoQNiFQNaHZTCmK6UwHESquR7V5lXo53BBmAkIx3fEED9FsL+cwUn97Mq
Jgx9bpE2PMFnJWi1GKRNyd579/981sO/d07xi8xCITPOJ3LxWQTPhw4LO8vIFUKUipsZhkq+4LuP
hJtBvgJRkUovEunPH83TpM4+eJoMVDNR2E2AHaOMZgvvHXLjgoRn8KEEEqTEMLGtuo9nL4dojdIw
OnIG5mvsOf2/ENDWxUdFUUkvwdqcVbhVmL37CIV0tGWYRok6Vg5xUxSt1MvUGWKYq/xOI2RH017l
/xAo2yJ5lEATFI/aJuRlFNCUs/YXtmZUD4RRbzd3l1+xExeBZHaV7ivVktC2EX8+ps5rG9tkrrNV
PbZqP89NwRihX6JAMQ9hyvm6l5QGDCCtuc70wsI735MJnJJzIXJGKDCyEtnUjuMZG9ux+1nfPgdE
CIrTxS889IO00SAyQnwn4UOdx3aj4xY3BrBqWjnhVzrfLcFwhhDigiD3rfVRRLyElOJAW3bYOL/A
rsSAWhgdgIX9zwBCjyb2xpqyYloWfPgxJioclUWIPWK9uF2QZZY32iC61ejou+urnHCAq+/mhRPT
XS6DtHaDfTF6u4JDWJ9QAawXV2ufYZRzdVBUHIQt3/ulQb2NE6ulrMk3YqbKVhr4qnNqdhDjD8HD
SGa57flSkpt4fiUewLzxAZrYujYZh6jOLIiDP201Md0ECtVc8W9GfcTcjrVVlj1ExispzVQ3IbcJ
sCJ09RVUtED1+7vUE282Fa8ioUYMG71ZuyJlkCpShtGsJrQMg2GicjrtqbDk+sZrojKkWd7Lrgki
OKeyatClYLqzXTpZhNmUPJe5flh/kpGw/tHtvC/BG6WHeozRw8olmKHqw9/7sJdnE6rpV2WOPM9m
sRT3wvLe5y0Of4Jxj3h+7IASZkhkqgsbkzzjmemfmAwVNLCRsBiXEz/MpGKylajhD6Ovb4hOhxe7
1hnd6u+GjrV9jMF/C+YJit2aLiRwzWKECQ5XI4CmipnLCp4V3CeYIqzR/wZi73ruZg8GP6lVI69E
s4vxj88RhEgw+clzryxS1mQofH/ll8+IKfAr4CLF7Xfp28+sku/R4pygUC47egzJtkItspCqF9mr
FqjsfQZ7idvKnHK8GwC8uU24RkzjTdkrgZ+IJJdqfP2Mbzjp8jbZMmz30/LYRPYgrIZo8sXYKBkG
0JJ3rgkulxwrxYdihMebGH9W+1nwpg6chBp0z9ibBF20LkkOVZnigunr93aFPIZSji+3AVChU4kW
rpihJblsomaU2zFif5xU414sRMloqSArmqssB1V5kDKvzSkCStuC3gH+oRq/KCqUdBSw4jkjtqKw
yxstdpKhV7rx4jfNQb+Xl4RBnpYgF0g1iR7z0V77d7avPDFXUT/090/zzlCcR7nyHdVD8bF3xMcl
HxaVskWMcEgPKqmVaaKO2pwadNhnzVBi+ZG88OwcLj20BIPKeTrrAQ9L8s1bKoIJuR1Rki5opZO7
kaPtNFTRjMpNjNDJP4cT/3yr9EtKbHMOs3lojFcKfDyy1FwF/K9dP1eXEvvTR8ERSU2Xxo3PkWDz
rED6lNaDljvl/64IhwnW0+0x/tQ8c9CmEivzZwx8gTicsSM5M/5kfZ2bjSfTfk94YzudzsdE/1vS
dTB845FU9+4EiEWLDbocrFImBscFlnkJQmQ6NkWiO+CcTcsng4za1K5wUmepHbXnw6HYfdIH4h1E
IXXpR4+lo6mg7HkeodWp14Cdmni7Ibq7a1AjeVG5wn0HnCIu004yp3gz1Ttr7MJQHaiQyzbKnLpR
uK2e4WkTFp3nBa0Ml4ePdaPKlpUkiDrRBu9EU1MNSarHm50nR2IHrzZMSu28bZlFqBbIZGnnnLoQ
NBcinw1QmOJ8BHdXG5i/CU48WdMiiZi22cMykvBIDFvzMs74KVfbeTw9hbAdJmJ6rHOZ7r/9V0MO
rSlf+i4sszsbcsMPJ5trIHr/oThWz2KnUZ0p7pSdOaZFRJSw8WAuNZA4GxlGsEGvUgR8qAhmHH8h
1eW6y0xnn+pjl84LC2+FLJkHg0mmQEMM/m4aO/7I1nl734gK5JkDYZyjD5Q9K4QHh9MFq7pbDtHI
mU5rTLwEpb8qLJDQBNbmZB2vZ+ay0Ti1QTu93Mhvms+Ri2Mwuy0bmZvAYwvnwLWOOW6fmUqSuOVH
nTTlaovTaumRLzrkNP4z1ifw15fwqKSwlwiTSkOviI+T0k8tGF8jufmQM3621tYGinFKmm7+9hwl
nPbf62jPmuMEF6ep927jZx3kRaGLcu6DC8IfbXF7zlst+P6CDn0NxjrWr8NdQRt/1BvJ8Xty8uT9
UilwRyYhQKIQLlGWe7JKRJ0OLkBf2+stGvVv9lvyG1LL/CKc7eNvE9aLIQh/JwgX/G31qoqztA2p
V7tCo7XctbURouLb0qJcgwt1OFXY9h6T3Up1S7ligCEzTzBy7syH5gAGZg1zLgGS3wsBFsCOyDPB
ttGx41c6/3UC/MD7qCz6y85OY1Ap1ZFlEgWFGR3Nw7oRzfX/UapRS0Sb0k6Y9LvNaKd9+Yjx2Pdf
CFYVIXvtTsmUKdjFjWrcyi0X9wNGCeEHt6LyCK+2LNBVkaj1bxWu+T8iGF83vCI8kWiZ+u51Enxq
TKS8fpT+iuINTYsxmW5SfLZcH9TmjAuxmVQ5Qf6/2McQcH/Fh0vrRUlPWc/D5UKqrG3G3TfHvJ3g
vMVQIsms077clTXDgxVSdSSbl/aCt/FHqWfnDat5m/rvgsRq+gbQxUt+zMrAHensGusKZ1kjXM51
cJPUfzvuU4of+Qh9Y3yB+3dTDk4LnLTToBH/PoeEdjrIoSlYvfUupaEUS5pTGnm4UfOYIBCVwdYf
AxtKOf/NuVNuFZP7q7VT2qXVYVJRdY9N/4EUEMVdGTwIvVHrD+m+F2wG66MSXa1c7KsKN0dV3TdZ
NwqOx36ZrCrciFTjD4jYtcb107nKRnD2IKQUxt4ZU+uu2c+O4DgQAw0DgOGcT1p0bJeorKUFXgxK
sBhigftZVv1hoIz7CuzHWHL7REiZmfi1QJuKQ6W9pElxeiT3sDKEH0H2ztnBr42W1IfbStnNb7az
eK+XpWJ5Fqs0WwX/wuVtq1Qo8aJarsvkHrsc2udznD7OvGl5vC7akkKE0Su8tDR8dai7wUmSRHtd
Ewm8bPPGv8GPxNGFtQct3XpIZQ4SRCzvnBxY+p0lsi0qS2lEOowHjQ6RXUvg+esDIEIANAHeIjB7
eGPpoQnttcQvC31r7vLkAT9L/e8luhEixitK279sVygCVxKPxGYaMK3xdZM9hUD4vIxhRBjDaNFq
jm31Edxzd99NXwOkSSpAdQpfwQdLSmWzKQZ0ctdf4y3SZcGgGVg3O14dngDornHCdPADCd7LyQ6A
ARlvCTqt2dp/WbFrm3fGeYiQjOa5TU5ZUVqxJvNVVms5YDRdQwEy1WEERsYc2JhvxIcuZ3tlccZN
TgNGcbS16rns2142dI+C2k4ffojPoJP0OvRy9swyKKZOmwPyvdNiyKkmrzZ1JoVIpb2t26DUK+XW
2k/AOuz7K0+8CADwkk6C76e1vjjMyya+DVfQxfrFQ0zWb5LxsIHBo9kXKpuODfFk6sraHffXRliQ
XtSAU0ajjKg9T4tPTMmaOyjhXvc7NZzuAdPji6aXNbWlRUD84FmNswp5Z2Gvy+egB7PlAXqKNg11
3iscbslbKemAatmJrvOiU0A+7bTUu9AOy1u9OSCU6qqOjASMT8W/ogPcOhn+0Riou0VQknVonkuk
qi+Pr2S6kIvvs+KoS4Dn+50sDDknwsdERLEURQOWHYpkrb7TaJxcWgx2ExS9PtwDqTKnNNIiFu1y
pVtJUhOukbT8mnD3td/B61C1BkfqmtRzGps/i0/6HcHPx9WSkT/PvbbY3001bga+RYkzQP7JZn7H
JKqcf+fZTnk8cw+XinhkGUpItwF4NsqJGuKLGaQFiJ5jM7Y+PNNBPKszW7h5IRdAVbvbMA5FQ7zu
iO6upL7GXFd1m878y4Dzaxdpx8/WLUw2KKDR3lg7Xuu3MAG0k5dmDmy7OY0ese/jBOh6X35NASTa
KxiA08brSqIdVKmUDqWUdjRIpsgvllAOIAx9WgMa5kHYb47QtHlAkMX3DlHOKUHBti15F58mVUwa
vVOhqTSxus3a4XWy4GZLhWCnjT3r8LoENJElc/kMY4CvSgOw6tEyIilWhAXcrLcwYfEKpe6QWBqG
6MjRa/L7kCBiCri3v8MNFKl8UEIVmgMLpWIWfPGa3OB91DS8ma3/+DKTTWWgXOzD4kVU+A8l5o9s
h3sjzSRGR6sBSXRXbDDeNnDl2OoRk9by8MqWQncfWxWhWNn3IWf+9cUZssSqfzcyxn0yGpPWiTzW
8QB3xoXfunmIMfsXnl1XZQsYbyRH6lrllQBzb3bXGt2X/hYjmk29QGSoLDNYOSOyhyMIqRk9mgMG
Gb0r2MTkPGOb527+URW6b3mXjtEoEZDfPOcdMTCY5bMwXApHtT/9Jm7031wydliqPXQORp2ROM0q
rwrNf6SkYxJ7nGnEoFxzhzQWJ304/OPVWLwqcnr8DXhuV3MRzyJPsX5wyL9ktU/4MCLEBDyvfoWh
7NXKKxImQ20EofOVy7pqYHa4MzAbcx1RqkTlOqscBPUyzWdU/5qR9RrCig5mxg3P5S3CTatUsdHd
/123Mwl8KUL9544fHeook9RMCzdLxo1ulB7sXv7ayhsxFKu2xKtZuI8ODwuoNbvvXyLzkPFrngrf
uVgAmrbJxJz6ugmh5HM8GStFzVwrfrclpIQEwgx5V456JmzcRHUfNysGesAVGcKwpbBZfT0+sUKq
KmsqNEM0NhGzxGnV333I0sxfKcajgAAPg6dwfyJd6FebSLEPm7pLFeloYqZsePvo7F+jMHYG2+kG
wAbpzSTyiumKYLZV4LWIvscg7WchCHglPcW2h+I4uL/bhHWV83GRDidc+TB8Eu3Vj0pHN7ksblTz
lRrho9RsqDxvuEttrpgUw/mnKKFAEn7FY9UPe7LiAVuWbCCV0WZlL3ZFKImbQuGraBMVYW/KWL5S
c41djA4Y3gZltF/w+nFVKf8EEwX/ZBhnZwslDDigyonFH9/F9RiWXi0NVXhemrLmoldOaF9y3I3N
YmVAU2EdAMw0Liu4Wvtrth4Ci3Ecp3HskvvaG5zgOZcubVK8rkktqfwxVnYPAWodTVAxaLtaypUx
XdX5k5slnFTVNXEwe7K1UMB8bv9MCiIjJrFnR5jws3Lvz9gxnOAvi/gqi+leQmdwOlarrAPUrO65
+NSaiV02gEmBgZT6NG5GPSYZuCSab2UvqVv+n+AXB29pEbZBP0vkM2cc+z4p+9iwqv5K4l6ocXTj
8argcdYYx+9b1Wp3/D4eNdYZv9m8xQk/AFgF7molDOEU9hoq/I+GmlrwOIzLaMjMu/6Zte9qBAlT
DcKk+VSkvBUx+bEodXU0FvNg7ddI6T/3YUh2FcVwPJQyWUCYxPYa6P3OJpMMVdJnU7zk86nLbRxs
9XNDZlILDkm6JuTWrSQqGKvP6K4qxxhl8AbqWGQ8BEd2WjyI9tsR1C5ZdF6pP8fvyQbeQgG3XgWQ
VJuxH2K9cUAapyh3maZXYTQisWgOIlAjBHDQVqUjNarES6ZU6FCcwS4sbXrpJ6DNH+OSPpcCu443
RXZ8dVIJbq8whryAC2qaK0H8uTClRqqsFPh2eYwIrVdmBsnHn20TnI2gBAMv3eMuX25x5OAZ22rI
+s+A5qp+qamhqVmFISkToApPbJdiQxW5xMimymz0MfFjbvveukUYFKxjO+SH8MNswBSEaH2sBQZX
FnbZ8yb46jDI9xhebm6Wgs2YE2H2sbhx1YshMDzqyF8sSuRovKOpFdwMxlc4VYG3C9pXs0Hf+A2A
jb9oKOaVl3WWm79+QGQNSDruDmCdCIoBZJqoT5GYrvBh8RMR0IwK/6I6vji61cqVmEBo24GWjEFS
G0UxKS7cWQhkE3Y2f+XmRp7ng6/UTnr80wuWY//a/V/N4bLrVxRdDfolP9Udd/6wXHlYr/wIRsJA
JU58c+aIKuniJnQPwS/Z5qJHx3KIAmd0uacYuqfS6db9xvB/Sv3vxN881D8b5I4KWLIQ5gHujbmU
t8vP/9iAdygjLlkJtnA7wjYCtPlsQCxhGVeK95Y6CvEL/Uicm0/hsHJEIt0v83cOSj1rTtLZ1Fnp
kAaRQMR2+MhMtZUzL9+nfqWKaCwmqLt1NKPoJ97fNUAIuQ2KbUWrfTsl5r7DN8ETVO0qqT6snCHl
cUTQNePGKeXccUwzFZcStd7CIT4zzUDHYWpVCY/mP4NhVQ+rZ8n0lOD5CgA98XjvM/va3em3573f
KroYwCkkyK/3IKyxvglZkz6NhlpS2LqxOtfF0dg7uugMT5ELPGpKXQ/q5dz4NgQERrMeQ5lngbyN
oOLZXo4mCgjjCD3onkw6Ow1BVKY7OB/JywL9SS4Uwm2UKdruJv5s+q7lKivut/CXAfIm5nKmSW3u
ZCiDfc/2VM1ueNJjOq+I90jsnDLIjufk2ia2+UU7DVtXqanCt9OtTE6IMuMo8/OmNrQ7IRaIkUyh
/kUHm+eOzIeUVhOQk+8km8EM9M2aEUox2ydRHHufTbugRA1I9nHh4TohuuNAs3JDKHT/IWi0wmE9
6ZuH1N1jGmwaYDSk8jq0mi2Ttn5shCS18jQj3z64pNtCLCmclVUnWduBWNuATra9O30VC8fwo6S1
Xbd7miDmH5d0Y7r1xy0QrNxxovw876FFd6JBsBGqAEl9a5dqkHjgdLOcrGFTrFo0uDsgY2xMmP/T
uWiRwB9Zf18yGp26GNkQ7EixKcmRC0r13aKkUlUKDnJvIuhV4PBeNOB2OHSZd8BKz2gkI3YYGjtm
QrT5ucsXxqMS2LaPRPYExwA5wkG1O8NaOf4t8SCwWXshINsjgsIp7yi8ZhupNLU9ZEWRR7TH/so2
ioXSCHGCorqviQvJ+y9uHCwoJBQH5ttsFlFA/CCc/dJe+hYwGrNkH+CB5/aXamU0ULTjH3ldJTC3
TduTW+vLj4wncw5gNbtUsDFUVbunQPYsjo0arl+oDu7Gswgm3nE6Tjyqmb8GFt5YDze133+H7fef
9AjurVFqKltnGMBDLQhGzUwLm4Q8vXfj3Q3Jr0lzvp6UDDMSF2cbkgxwHmQVpRbWIrkicTUzgCEs
hEANpHY9Fk5C4fCGuc/aing0C3p6Udtn/0QQKTJ8S4uRKrpaC59NZU+iw0bOtEK/NDCGPfB4Ly8x
M/EJpdsT+IuF96dbe99vrzrnpxpsxFls5ZdG4C3imTsVoAPRCXFiMqRCADPxBdHM5E27zrofQqeo
CddG+Fya3goZ8SsK4ufWE3zjBbvrxp/Uby6bQRBg/EAu72b2p7kYiLogX4J70unAOfGYu/mbudOS
rCfDc5KJZ2ko1ezYKFIc13UA0W/kvkwDpBWq4+3JAw5tMFIhyyM2ToCovGZHHAhnZ5MEM3G3USgK
5z+0hicpEsJ/TyGybbvENwSog8OHB+vtlzDIW/xP3/efpGQYkE7hwnaFaAqln79EkY9fn95UKQ9t
F7YdAhYrk+HFp8m0TpaYa0NqfXv/EcZTDrRuCt1j25I4Vs3DCWru2Xvcwtp+jnCBx/gEfgU+Gtev
tLeLgzoPYlNCW92w5X84fO/x/R11OVQbUjHY47ITZi468MiW22GqoCjiQ6gnQhL2Av+lHaM10+vg
XBYVsTHKx6eGzytnfSWEzjFLW6UcsfU4qx6+cT61pp8OGB7xOtCVxaOMsz/vI4PAgEu+SgYvFank
asUhk+k2ztTFJoSOOwenERxDvvKEHMJXW3l/sewhQOZjxwkJJhZH84oDnp4k2DzPJazTobTa/6CW
Me5b6sBaGxQiqB6ijTyGBuTrVRsRQ995p454cbNiCFd6e1b8DHPA9hmCE0RrqccKdgSB1pg1G4iF
Am0VVTkkTS7MmY28TFSSoS3GxifLJ1t8jmKhtcpD4+3ZADIilcU0jlOUk+aGlU114/dONjAA0IPe
LFpNMbMrAIyojiO2Pq41to1LgsJoHPdk+zSUwRtK8Oi/Lq2BzIsdsXluYNW01IVq1kZAxM5eTKs7
LCfBwmTCuENDnSvXAZVgIY9Z/AXUapI8A5gIDPqWQaRifuQYhlB3vp1U+mpRS+YLFf/OhzLOrQLJ
ajhBq80N8+eZo4LT1xYduaEPEP4r71ic0yHfalIMdd2cAw1m336Hg75uEKDJMM73phRxOa3IhAVU
yR6iVogm95N6Aq65OYX36xAfRcrUnBN5c3kiYzGAvBLhki/DzqWRlysKdgFaPVrdVJflr3m9XpQp
ZGHwnVN8woyfsohlq9gxPqedg6S7UqtMGNzM3A0itn2LV0PRBtVIhPenwiQjwnE1qavoI5TOQrB7
txyz7XmPY6fwasnbr8JDrreiBO7i6S7IF1y/6E0XDxYzXXsS8ya37u3d8o+2fmIcaIN1OUoIioFo
ZucmBxZxNH48G+VFg4D0zNOa0+bidMjzWX/tZ7SzFOUj4JyFaZVVmn5BFZ6JzVAnULLTAkmWafNP
+zuQF1lYhxewMDdqWJLj/d3dkif+GGRkwPgVZ5b3RGTdBXWApHwYk7GnWFKAttrrGtEDOqSRoQ5/
6/IElIIYa+oUnZfLz1wkCFYiVg7QmLyXea5CMcaI/un+4d3hndOPiesGqcyR7j5AIKYW0IIJtk50
h1HcwGP+dW7D8aERtegEv9wcaLftu2PP7izt4K+VtVk/648KSsbqDjQlIkZJ/FXiWxS7Fsmx9uTX
uXb+0+KquQKwu9iWa4mCBVNKDJFqdYu6pHj0BIoWVm6KtRxK9Ck6ugPnzJmO7TkqI2BeTPCvJY2Z
8Fsosr2F3OWZ1l8b4/7JUJn1l9BmZ+PIQVQzB2hLMTE3tw4U8ax3z4UC1+CRtlB7vUrzt1GsTPtb
j53t35h2YQg9NEbjS46e+uhi3l6PxZgo7bBf5CGUMMKZh4CnEHBGPmmUE0YshtPFKNPzsNv3vRIu
MKXFK++dWxcEIMpfW+9650I/WOUM+otlCGFcyfZPHjS7g73707lxuYWbwFzDQFodRsrPBo30celP
OCFN94BfRvIglR3C7YWsJdayxDVrPihAxNkxMQ/6JgFS7f6zgf9W5TLYR93WQ2bFUIDHPr1141wQ
rW1jyXF2MtZjfEClQau5eUGy/kKKw75rCyckmHbsWalavTQ1t3cML7WvMDxTHuS6I0RCT0nBNSl8
3He40LfxyIfp6M/qr0HpMt180NCx1MfrS5zQQNQFkxRiIfMTdKDT67fr3fkkFVI6kJ1exo51k2oE
BH4lxcqwiICVZ+TvgWaZClkAUExa7alMsNicMH9lIrzUcW0JY5dgIZ9gGaad+o3EXZHs/pta4Syh
zOsYA4oKjQ9jmN1m3dmCUeC/0a3glo0bd3l/bGY+cSVPY+IW6W8YcXNznvLPucEByX5VSrcf7OKE
kpLDylwEO9FD0XnLP1OJf/9j08qylfU7WJG4JxDO8COzpCgkzJLcNfnsxEYdBwdzPMCrhwCw6tPP
OkNJaSw3npZp166mCQoiZ4rBFO9G9/CMziwn2+6FZfQYLpugoitACXKOkfb8B9bqyR1MIfjoWSPp
UQRDIXIl5IRb/tDalhUvHBbvujz0u8Yc13Xr1HnZxBPg1Bqxmu292v641T9jqQrWgl7ns3cJRyuD
WB+fz6bNp8tj+QNOnTiSrP/k0gzpyznyxvyRmSqq3bqtHTmj/DW0aqFbaNp8SnQqmbN/gQTWpKcG
TPmzfDJW1ifXAljtqfoMnZ2RcptdlH09hg0159VnOmQpGIrG14hDwkcQHude/riq+kORJRZ2vpZA
ZA0azhHm7F2Yomg9p+ALl0fBMO79CO1zEtN19EdauyML5pjgIGJ3wDNTJaaochmWhXQUKWZhO1uM
gO/8HsUtZoKNWgv0ezmFDHLOy/q20tBxx5IO1aSPG1kWGmqrV5ncLTPRL/Vjn9OfuQ6gq4t0CQxq
wW+fl7Lzevc/a9l6aj7c9XA5bT9pK1hHf4MRW4eheiO7uOwEo2NwGOPAlmSW+NTLLmLxplgUEXUw
O3zkJt7/VsiOjXDg2Ou44xA5t3i3wJyk9u7O9xa4z1RzPQuQHsz8HgsT7ZS+57ttlV0a9xUM8/Di
HYo6Kh+i1mJxp2Rb1oMZaXp/btqInt8b2G94FtgOTK7vr54jswMVf12SOdvHeWpdQ8T+/3MVkfSg
iZmklx1hNTmLdXKTY7qsfYm4QqfydOb8ky3ok+vQhtIty0VSycEzCxC1nyawA0DmJ+tp3pUR85ia
ErqI3FarCnM1FRXf0Ats1uBYXp1Jam53I34g8wWdK/Rl3Wj/wJ2qPecQFtRZwBPRZR/7tOLNVZqk
IB+Zx0Vzm5OYLED4Jte9WFelext1BLcFVMvw/Yv56bQFP3a8EJKFpwlKTcQWk+vbgjYa248u4Afv
KPTEqOjeB1AjxGwONe1MrakFjUuBpWGMxFfMKcKrz7E0S2/1vFXvwse3p+ZrcIax4ln1V5GA1idV
h07fxgzZSK6keykaEfHz1d0uoWuJ7PoL5BDGE9oZteg3FQzN/WcKQ9bcTwhEdW3xen3eSk/gZXk/
VCYtkYcEXkM1t3R93dzhzQkll8i9c4r64rE7ywk6O7YtrRfD5AfudYY06mdOcbOO3lhn4ivGhMUE
AzyQwp4ERi1hWaZXhWiPY153GbBj+U4fZi8w/eGRDNH2OjjG56MPO+Fh59GIWYyhvu+f/HG87KAX
jq9Ug9/a9wqrkkIejIDi2RxybGLiVAkMaNc7UAV1t3Gi9a3gAzyzFrgE1yFj3tn3EpgoKodALf++
gdYq5W4WveO7JvFn9388Ap2sIoXuqVegYbTnxvhqGkOCbyc4k1KwY0E3sODOYKlebKxztmeD+iHy
R/zSFly/jdEYKCR8uGf/7bDX/QFFA4ikd3Urhny1kxkhbmuD/6oe7gjkK4wyu/6DO2HaVq46plWZ
uTB54w+w1A79/KYcGuokydcg/qI2gofOK2ShcyOUE+belGy/wAfcS6tH9DPuM/9SE1sqgyFMs0Po
0voxZRUnwg84ByVoOuQLEC4ex/eA2NsSJYQ2yqIphvb2q1Pf59057WZ5E02cWR3yJ4SfGbi8uOpz
xt4m3egY2F6tyeHzRe9981IzUT2mnacGx6pxlvkH+j4MCn5A491R/BmmJxVbAxu9Q1W4fICk4HzB
Rkv4Ub3hfW7EOX1bt1sm/z980BGagacVWNmlMQN3AODNj+GHVt83NNthi6mnXN61Vx+kjxdFEq6C
MFMGJQdv6WXh5C/NCLMDyDj8SQRJM3oiBBk9RjAUqNZkGdMqQKXp+jl0HuUN50XtM6Pp0xb9iDKn
c9AeDoRjZjS2rnX9eUYj+octDt4lSeDdBQ/PP3a7H/pJIMIT941T9HI0ey2ZWR708Aj4dc9ax6mt
loNKHdUXFJRtvi8WxnsuMPBt0nN2IBnn5G8hq6KK8U41EhT2IEMrQIC/5NY4DRAUu8Eg4Qxu7iwI
XtkTxHpHqD8Lz8/klks8whPSYfQ+exIzM3gi66ZBFwu1rP0NKFJCLqxmwd0Q4IyY9YfrsNxndlpL
6i2rOZQmfB+dcHcM3EYpgYC5FDB0JyxpAdeoQ9UzVIKBodE7veyEgsL7b1cOn8poJdNEhQOlR0kh
3nNklpIxpr2HXzExLkOcSxduFhOK+Fy1tZMfsjQDt7pYMufPw50Tz1JDKl0aJhE5owcdgZnygnTr
YmW/zF9cjM4RybzmGgxk1/Z6t519rUa3nqoetV6+t6+mphzK3U+zppTo8ZPD04p5ojgPmDPdfnCe
nS+0ARw+CyNVLq7L8VIS2ghvRBGuD0sgm322b1NtiS5E7o1ciYECJoBoizFYZl+5j5MrE0l9wlOL
79IFr9nBCA6nS2PFsSHmHZddhJj2yVxXFsiJvY7lujFZEElgFaJsDMpJ6qwS/0T9se8bdrhcwt5d
fUOIbMHCLHTlUOZAxZbGbVtmfUWdazlY4DnQUVyBWVlnO3Gfx2jtjZOXzefiGhbe7sVQWuoOf2gz
Uu8VH3lL5SjLQFYxECoP67tP7rNWYX8D0OknYonUk9HvHeld1dAln48JVka1gO33dbo6iRQE+FjZ
3Tu6VSygywnm3zvNrhbXOZ7dOTTCjTp50F1G+h1MhnjtGa0fF8zyqFvePO9m3yLnRPPZu2lto0gP
NV/pRDyWSNCMJMe7UrPOR+IYPkNmo54CYtmBxRXROwpHkNPI6BDovxjpDcPL+nyLny9+dYK/J+vz
G5o7gc50f9+Fn5kl1HkNyZ6/U/LB/AxW5nQBAaLZU2eoahuhbmC5hoqLljZGaHHWGCaJ5Y1eyETP
2F2aK1sQQywTbdz3ett0DA8HMay8P1OCxNQus6UB8FKJAbFyTafpZwTNizp5kNIOaUCKG10LRdm4
ftQloh1U4i1lJFmeSf6yIkSRKJtoL0BWhSUG6HD/5bOVggXVmEhR5aCT1EhUQRVYNYawEUjOYQBb
z8UFw/mWqOUIoFKCNuzv6KuuGVDupnZqvxqh/cjxPdL82aMkEuEqgd24/3BnN0dMGVjLioSD1PWn
sFR6uVmESboqkljskP0sHsvCr8u3EAqm+5tIkCU/TMvas26KMaJ+QuB2wu721zHYQN4ZK3HDUJ4B
za/A1YLjZ1xRl44lnsI+QkZvgkLjA61S2myeaEyhCxDXzAhZCMujlRkytJeqFbltADG9OxhHgMAu
dhqu4JBpXrworTrmhhhWhMqp5y7PbC/kotPIPYfvafL5sbjNfBSK5MHGcVl2UZNDiqnsH7FtAffh
kkitTVgqaqF33UpfS/9cjVPa4ykq9ij5Kzfi/1SXnGHdL3AIXW5iY1bWrKsVy1wtdhyPjb5slxMS
Kvvm640jJ4ilHZqa/dDHPW9BkHXNnMb09FMPuMqsj+/tTs/ODTqcKDCdRupOshldFpWtJVMUtcHI
AvRw7Hqu/a63Zs14psEjBFqfHHU3m9DhLAw/56tMLELbVRkUzbIDslsXFKJLq89R3fKlMRj7sRwP
SXKySVf2KYpsaoO6HdwViAjOVg9P3mavzyEPOjpUumvzT8EgPy4gOeiDenRqJVjYS5UxKBUlURrd
MM4XEkWXMfLihDLk8FCvhJYbD2B00xzGSEiZADm16USKjTHQ0OCFSWSO88pkTPuWWXIKznyqT/QT
8HxwFx9tHCD3ovMSX+drdFzmZD91TfnzzsOBkCf3ND+gkOmZO7eekuRB2szFl5N+lPknyfagdfh3
6YcLsYOeJxf9LS00iVIoxoDHLY0LPIz92ZX/phuRh+sM7StEAdZOQOtFaHyls5rkyf8bVuFoOBD0
5+6/5drLotv6ZsPEW51PpRw0ObbcSoFs/RPyiy5b7PsAYgzfm2gesW64VwW9y2/N/0x/4P+j7CND
C04wu4J+5eJ3GUdvqFqWXnyyhrmdLZHxhdaI9AlprarrHtJknm2Tzofvj1qK2695F69UZt175zDs
9tJXqmQwFkjee6tJYnmtSs+hk5XnfmIulsDQiMoI5CZqU2zU8C8F8Xm/pchBjq+ZCi/ZyczSgaq0
/R+4M+wtOl5RoajeCYn7FH91XmtpoMSn9+QqaZe6ZBAL2c61X3p4/LcyblvKOU215f9rEXSIsc+U
fdjCSGEyJ0EcgRgVPYaiqHRBxnntOEvAWTPU9h2N2deI/Svyu8hZG/FP9uqZpaE6qCpObLARg9dO
ae7MeOYbjsAfFzXvlfpByzvu9Z4SU6lB5MUfGX7LU1g1YVwn37UI+/T1Ul2jLMhVV2NMCFPlI7Ae
v7hN5NBuTEcCwHXxF76p9fnOtIW1zNEqFf6Iq7LB/fcj594HSmgC34SY4YAk8MH2rqlS33yn4de7
7SH42OG0nFXscV7VO9zrf396hY0nGhbCgglyXjZS2/8gl0Y7r4gnDsa6V8TNkmfyKKhJqBdZg37u
J7O9uJogfAFOUEXq85w8bsUZqHEKQ7bX2hyko8rf/4ZNdL+S4R+b/Cv4oVCV/38W43FmDt8gfR8K
uzPJkOX7ZZp/qIQ2Xg80OWVLQe3IzLh/r3r9XPy+umSK1psM6JAPrsjp58wt1IQWMPYHj4XZbMMT
tjNiGX1HbqM9MYEOC9v5M8Tf21u2fkX8DY5Y233vbxRjtXHc8qaIjw6XoFaaCehtR0htCWgF8vAK
JL15/G1AVs0Anoh/DmxKYheIGmXecAX53McaXZg4P9se7dvpsiJjGPpgn006sarxN05/f4LE524d
bYAG2AiJlOeUZdJ/r4MGSoGDWEVrEA3j4eW9S1ZrLsE+YiXYo36FsK9BhQ2Lw5ORDSS2uWCY4+za
eD4+YjKMAgrwvUDBBBXob1Mee+/VA7O7GIR+uOjKQ2i0EWKLPhlZCemKZ4kIyn9TpsnL9c2/X71Z
KduMspQzkoCRUpTYipe8H22qjgcvjBeuOIILFeYrfgZ3aGCwp18NIoyl7/qKYock0QRMnfNJ5Mta
0YVtlPhqDknIMy5PzdmKWhqz9BBalI1wsd0K47ODz6EfX6Ja2iaoPlsxdApe1EQU6ZWWOSmWuFCB
W9t0R6TTiWSN+w02M/vdFtUEgCA3uJpz+NzFWzhqy4XfIvmsEb6vqyV7fseTFfk+p6twraQ8iLO0
tUU32/pVm/PJ/Op2lacAjnwHFVhBdC2yvX/ZxjqlEhmkRSYlbmkxO6LXdJRIuG9rejZX9upbKwWn
Uv/xLzOB+YpX3nCljUs4iP5rByWFI/PzivtlZmf9+j0irZQJCf1Sj5tN6vGLbbGdtag0neq4NAGN
Z7mpcirSlimqp5hy6V0jj2V9q3YiMFk2HkDSdaUwccp88/X/7rZNHyR7WDBnWDE4B4zkiqDdYVkF
FcLVXiwKbu6g+w5wHbdlDjkjzy9hysWjXdyh1FFSr01WcDYN7U7TDFr1LWCBapjluYnjBP9tcbRI
eo/WC5hm+whmomxP8hLG/0MkyPhz0YvUMJ+Z0dOGOxb/8BJqBp+CX1nLppL3Xezl2fOi62kt86sB
oBvmtMqy4jfBRl30oMJ7uwmcTOdFJNo4mLWpNk78VCf2p2/BrwrcUbvNP7wL15vPBL8e0zr9r4MH
xOSB67RIQqK9gjnYMIo+xDIB5pX7zCy9qCkodh7TIuZe3e769BLPrhKkiCSYwBpCzV3PgaA2WKqs
f3GZbIyqfZwHR0d12mwFFViOlqzFNvCjC2cEG1UORsTRoKFauU7aUdtsgwGZrvH5lGWAr9x4/CeW
pGfvlvecEyuFgYuxX78ZJfTzoSs570dNlF0LYKaFTBuZpPRLz+w6/kqqiKriu210XRDwrKhtVcNI
uML9imhMBha6dCJikSBM2mWHm4L/IYmbshb2pOM1JsLt9XEXlr1D5HpXlcM/pF5ADHRyPU2/5gfd
oMFBdz1R+AE4tgnJ+XU/Ni2W2T7tMnqK87SOOIvK7xu4Od4oGK0DA4EWqezajliuy0sdmS6er5jt
I61I8w3FRnajyXf/elDVGZd8lNVkzX8SpGyhlSOaRU3qL3NEATTt7uKZA5dgJPvTFfEKrfRvatgk
SAYWiY1bs04Y/pdcroRV9qoytwOD43wZLT3wAJA3rXCn4ru9VDbucQpHWby/ioOLT682NEiihYzs
s3Ag8jiLGBqIwildX8XJ+Bb6Z2lPqwRgsyuplYXsagr/1/bGncFcfZEHnSFkNgjZdIVwsz+CYi/r
1lGsbdnjYZ7Yjn4RXNjRXT2oydzcyKjzOK05VZ/xXIc2e6OxYUDcJI/I36rimtW+fKLwBSQNP3yz
7b5ItF0vCTa6+gJ7oIiAdsI6B9W+hBSHvLcB+4OafTFVDoySqf+297uQK8bcelSrkwtlPvfeSyCV
eP2duquocqUFBil1tMzzK1mvVy6m4PmdnWXOtsrRlSQHor91hnnhKqMZQeYyla8pG1jBeQYykMkz
OsoKZDFmNomXMrm4j8E8vyxInupev/PfZaianBBytG0WHWfU1QRo6RkGB6DjYC23+0ZFK+Pu9pUO
9Ucb52z6RrLGXJ93XRJLkM5Z004Jl6iTLIpJZO/bsOvHuzvZ9fArZNXk1DwtGhv2BT1ckEIqhQUk
Z+MDI4ITjvzvar6O1EjEsV/SMfT5DhHmMhK7kV+0QFTY5e/32Xs3qMiaEuA2WfKJSyI4KDbUDsju
5TPE2UtLhoONXbxFWpaQXjpShE+jCxZ+jFG+sh3pScBgLTM9ypqTAvGIUnM0/g6CbigFV9gMqJc2
1HwtSnO+w6mOsnL9upT7Ms0oxnGX5egjq34M+6OKiAn9RjOb1GjyAzsdNcT9oTXBm8/gGgufCft+
cc60aMQngSSmMjPcSbHsUt/GqpgXInEgPP5BVOCIHAXls6pnwBpK5cOdkdVudKcpEXcFjQKSSVeI
yDyTu2nHnUpAGLM02HAWHrR9tTZeyzaKqxu+IoEpZ4HJM3CXSccwBeDie1PHLR0DZYMFSjXNKLjH
TIb/moNYlHtVtaaxoSbjqcumOX5OFP74MTaOpzNOjddT0ov6O7SfzEzSV6xheHncwVQyA+UQ1Ksa
tQK0B2NgBBC01kIAFSmAQFu2tKL9411de4I2nR3IkP/Lb037S/zta56dHcghq/axrQ8+mR73hgSH
lVwv7WJrVtBbaJTBBwYmwo4RLKHe5uao/7h5wga8zWHZdXeZ37Ls/0gufAqBEtvSHf5HS2Mc35Ki
XyX2w39WHvSxLYOrdrRFR9t/JbSt7nCiPFBCd3xEv/Z//GP7SBpCD1AG6pggeOhsU54hmG7LPuDq
z61qnzhh5DNOcjL8TmpGaNrPqcSEyohirK90mKiBqnLVqNoz/j3EHzu1VpSymMoFpZSB8/tIrC/0
zHfLv4Gmk8BuPwJ3ABNBcEFqVvZ9gVMEhAUGTbFDWWtk+NvGbZwSGT2QP4fMjaz3kV6o3L8DCzrZ
Sw2MAWHnZ7ernHMedkS8k3dsjhjHc4tornJzsgPk6F3aHTiNXtrCZFV938bHa/85eGKuFYAvTgNv
f3acDKVaVpbQiQrmyWIIWpme+hhaZCfQ12gsf5nQWzhn/9KCbfDdx8ZFh4F/MW23x9mL3c50AxFC
hblNFcB5twzZ9uHE6NuwkEW2eeBOoPXjb2oeNvVvrd/2M1Dv3ITJC9d5jKON85IFru/o7s2b+Hi7
ESM57mKWESPVfehV9x1hUSAI5HkYqAcJhAfyYPRPvc1wbIvi/9AeIPbyLNcu+c/RGvAUgaC2ksqT
JsR7zUxQ/Rx2X4PNTzGMfDu2nz6x8VM19lfku+oeTwsiNCIxtUAqSWGQoZXOd+VZqH+07C/bqbnQ
zNzLW3LEaPe63B6wwTiEOpfxPw80kTtU2HswIjL5W+qURYKnFQT16pKW1jEP+r7RLLURdOuXuE0Y
T7pC9REr951IXhwwho+ySDdl4rbHHYHG9byQKPSWlzPoUr7EUQJdxOeFbbNmwJvLdP8j96tOjTlu
qdXGQo0+oFPTQiofrJVT3jMUZ7mgElzsxsN7qrWIakmmBdPBQymX2awwSKz/snlBI1Q1cC0AyZ2Z
UUQwb6Wxr9foElFEOf3/4Yl32qICxLBLUjk0yExMbnmfchhBguqySM6TAN3IjD1MAuvXYW8nOZ0Q
T8BGi/F+I6LlFiKOkojfrC1Vl5HGkv2uhBypL9qWrnb+uNum5ujaOzRdEk3F+qpKUl4YYAPI46Wa
z/m1B8yfQEi9JFBe00MTOAjfFJERO76Z+2brnPcic1MukXYLIUn1pT67p7sANwsAsSyTE8AlHVu3
RWOi/1DG85qXT6U3LS+qiaGsZDzRDR2FE+9UquwUsJZZOTFCQ801VjEIpIWhaFZ6CJ2s2bz5u1fs
+dxYxb7iyaG2uAj0I1HdUrf97kLT9P+jXE3rXh7p7I+jHjzGj/jE2IyiU1JeFpRGEGTNWxkCZKX7
rt3A8dGrLppCGU8uKKFoWqsTIFd1ANgfHYjwVUujir6L8e6wimgsdce3gpspHdu0N02uI3fHpaTp
sH9Ef74wWapOjPr3Pq4BM/MqQKHcTFYZlZ1/W1czS6bJnJPWe2Lmvm9n6cjdewIXb4TvUgig5w1/
PAIOG0ik3VaiTtRfWHssYPW6l1jqr0nUj9ggZsaQmGRyDAZl/ZrXJAqhdPPLW1N6ZzcGsOiKoUIC
1ObS0+cmPrNumRtK+tTduMPx6hkTz5vLoEoQWFS69h0dqYta+c7HjvVylDwP4MrZIhJcY+PyGkop
2AWyKohIeNq/b9wZcc7iusp78wOFTt2IYakwo6cidUuFVInNuBUWSX8tUr0I2A2lQ3Q0odFw8ObY
Ipp1lYY0KolgZX3DmJco4ktvqZwI/xmgjBarioEgvJuVuXqEkcqrJlhnQRZVS7wU5f8Udd4lxaif
JcmmKEyfkahskWePnwjH9QcXqog4Ar/4A1EjYEhpWZQDWjrrvY/X/A6pHuk5sLDFpczfJQTPGXVu
QaM2iKMogqlKxwF8c40JRA59Qhy5qnTpgLujobx/dKOxPKCZng5MGq+R92J+yjPlw2v8XpSvSKt5
mMK0+GfzgxaRRARvLRaGaSnM9YXIgupBh+S2xpE3jADSefCUySQgbmk2qax2MblpA1sZO91+NP/+
oVfp7zOHm+OcLEzO3W6/7z3xn54Vd8tQRbWOsPfhTMauHogp69Z53VDCQhNx6DaNS/HcEBfNqvy0
HTY/tQfJ1FRugw5knsR8i1Ob/mI0HBm809w/3QfbRQjTAU2wfQAa2Hi8MCDIFpzn43G7DGPvT9cz
mX0hSOVq6HzEEPLX0zOqwpIdhj0ps2nAEkHN1SrdPFt6zNL64tNuuulPg3ajdXVaLsm4fzDbfkO9
YKqqZCMJgZqDuJ5ioseUJH3mSAEfhSFU4bdNPxof9Y/b8nsO4W5PVn60dkK7hdUtfdeN4W66ZJb+
uxtOOADi1q2LooXPI1zn/w+L71nkAxUEZuzK43L8+gFhgnPGgDaIH0YV1kuTeXfZSvyfdU03RQyM
Rdst3tC9n4q1nuukreCfQYIP6jwS6soSUE8YP+Ookd8RiA1wgr5dqOfAM1HzrMO0+0Y8J66N6VTd
QU/mfVkQUadltvGMhx5iGk3VdmcN5+D385/KTBf12W0ZUM8WcBp1mjZJy3s/IxbD2rXeEg3YgfiY
TGFOl1tParXQMXc441VdsaZPxMR0LrScYJ+mfJ6EJ91sLOhc7aSH/XTSwP9c0z04w5NAJO0R1Laq
5aQstLNmZyRuhl8mgS+wpnrGZBS69JTRStUrvwRCrsa2TBd5F0vtVKz6Bmxj4FdEij9nG04fFEiZ
t37nwTB03OxQKDhQxuOZkUqlbPE5pE8/MWHCVxu0eiI5FPeKx8yxg2bYim0mRnkNPEaZMFYyuIwN
yUtFf2vm5AimR133NdehAHFzgZsKblzPnVHmLye9St5qB1mOHBsB/i0quhauj4S0umJB9zmP6l7O
7NlQnljZwcOnDwSxQ/U9s3Zil0WffFMn5OXYjsQi+hkLgnrFkiEjPd8njopZvsMzoEs+iOoyaYbq
5PWYvXZNp4xDhQKnZGdrx4YVWuqagQyWVJLvQ1A2ylQ3gN4YCD9V6sFp8Rdnfs0CLfuBC2JEj3hI
Fj/5TvEwJoMRiaC1sXZJcTj04l6ccZby9+MdGYBP/sy8dfPfMlGMUiLNzALO6PmK4yySuD0nIPpx
wHL8RkzkG4cirpPSsMnZzLnZUrsiaVkzF3hnh4p6ftAHYfQEFs+JqAMCqKRERokAYGWmMcG2u3WH
DJBEWNHZQP0mIcjIgbZis3PWARCdojH7uoZHWkuu9qpTdQGzOLbTJLcYRacD03PnCE3uqemCaou3
frHgY4m4Utt/35tTTNyWe/nNckjxwrIPF10Lvs6g9yzCmD0xbbWKHZaXji8od98fSUExv/gec7W5
t3IhvyHeESm9inCiX9nuuD5xt5aKkasgCcydDXEYDtOrHDoyGtzIJsCJi/7NOlKyCxgT1ogdv/Xv
5dAVESyh/2fBpUYLZX7OO2vDImOPaqk4KsSjaNCObD3kgAwO+2SsvMjoh8kqqT5pIpOEE7rsgFg2
umHx30vgYSxah5Bi7H1j734JiWLtK7UlrSxA5Y3ai/LQI4zTqx/vHoNPaCw+/I++TpsGz3kTWjHY
AoaNNwQN8IDHkMZSZT6a/y8WzyUDBI7PbDYhKedWyPDRmb5XI0uaiTkvYhdJxYKJ3pMUc9VJw5M6
jIBUT5cTqUme6RepcLPAzU05Xt913fyQ5/G8JjkKMS80ph7de8vCIjSr/bdltL5TOVVawGRrrPq9
/nGhFtKQwzpzXuN4veOKVBHp9BuFQ+PHlGh3yLIUgU3mpWgmc+0Ligg4vzX0Kmx7QY2iaglx3x25
S3XR3mjSx2ZSWgQZkwmdTfhys+YAkfxHa/ekPB1mBZGE+BPoYQ7X5Ku2Tgo2XB1iBI49F3g9482S
+BR8bBVeH3smNFDDoFFLNRBsQN9GsFEYYV7DBM0PruELuC8fo/j6wCz06nZqTbcW8MAIcGGrjYay
q2tpUzcU1z3QNKatmtek6zFQfDib1Lllb5UiJfb5lSOnuYU8kFncII3awKRk5ROKA2LOQEpCvOK4
VGu5swnHUx6IaBsHHC7e6y9uLkwZLhtLP7xuuTRVBSHeLGA9RXmyv03+JvkjvA8FpubaL3UjoU94
YnuHOqKZEGzo3Q85QdJp/ivdx5NDZG0Lth0StxZhXnLvd7ImvwDsRjcW/0w/uo98myTvufd4QQh+
+B3ifQLhWQ+IQmEafcya8cSjfyASH5P1Dwy0rn8CDb3ImBht1UFzBEKEAH25PBZEUpLrB3Z2H81A
blHjShk/mu0nnkuawkiYpt6aPN35U2jdzmBtun8Rd2cCSW9HKVEbhMLT/5POQICZ4lTVhpU7yLYI
4IldlxDsipo/Jk3BljVkRWhFE6pD1Lgx78giS9clSZk9cHAEJr5wILMdoS/LNha1wavZrDpSqRoH
vMEZLdFJtSxD1tA0Fz0602zDEQuLEXyZ3tJGGXZfM7ptzlXVEB5z62d5vSe2s6YBftyhgf6TPdIV
4P7FD31Pm+uwvCJAQPW2u1epTsIKuDhJ7lw4RUTuo9tg284zENTNL1J/fJIplz9FiDBE49qnwsog
rlTcqDgTQHrRF5wK1LqK6gf4oQRtAaqVGkfqDmAVqdX5esSSt/BKvXK2Eo5lr84m2mDbwxGR4xZG
eGCAGaVwE/ng6elKm9L5WXzpemrw9cJcssh53vMfFClLFA0NUvpUNT3m1kuM2Jh6xkZvi4r6/2pO
ZqgjCRfcCamZMQmItYoOsb0mUMb7mKmndpGsFw1O9/QTJmxYXztRQKGZzHn0gKPmLLuyWDKtecbb
aaaQyb8Z+WxHFsU6ToXrb9byW+VHH9gGixfVoeeQV6JhXpPtEsS7/C+0fqMsru7xUNUTGWkNkv5p
JVgPNyhoT81qtqDuppuJI4tsQAfod7wHDf0u8oXJaBUz2FOLOfUKzDKOMatBMhTObvDik42SOmTF
HTDnBOMM64eRb8oNWPS06mMYwSl14jFjA32hYZxOisWCj+CcJwmJKJni51w3IbGqbipPDe8Xl2Ew
GP/lxCdGhUl/JUArpGh0V2hJX44C2hS+hVH1KgW7cBf/f6PfzSSrShA8g8TGhMk09wbgzwo8uMr6
f+ZQ94K02o+RcFBxEI8H2ldKW63N2OgjHCaMXJh3ftKqq9pdAQmIsdZSqsUuqvTECe+/Ytad7DCP
sf4aDH50Z8mS6clvrTraqovBnWcWDDbS52WME/5qv5M94UPia41fVlMgddUz8wpvcUA+wVoZmOdB
oto0Y+WJBhTpfd7WWNhTwqS3zOTL9xVzRv7sUYRGmGNJ6FAZXV3FqT6ys53eJ4un7tWVBAsQdWPX
ndoy12RRE+jgQgJReINxQg9SNluo8Dk9gp650U1T/+Xd0c2IsimnBqxKBVSFosFGLR1xd3/fT6Wv
7i8a3QTats7lz5WeKPcq0ImAlraHL9YyvLQLAGSJXF8B7hCH2eXls+wxBnyNFARRjATqfPUYIuGx
c6yRyhlXpMkx1JOnDZZDfcNcl3I3ukg7Zt+4PLVI5UpcaUPB0ZKIBfjBq4X5u7YbSzyuewnHYdum
9vJKoqJZBoHoHcAa31KImjgFYeRMjCCczPxQAd54FpfhgyOCUPHG5uLd8neS0cNTlOZxYzjH4z+A
Y6RLWNoXD3N7RC2xqUPl89An953+puSGY1fgedyYLwhCG4uE2DIF63H8GiboDnaGOltp38fI7jNI
CVke59mdPsqIbTVABGvUqyfJfoykaHBLuGtr4mmSHz7JHn3jHg/8a2uB5nwS0bmwqDehrSlwdEXp
SPMwLoI90wy5W2hLVCbEuNU58xk1WqqhhFlsR+n6oUw/0sIDHslrMFI6JSJxVpTkiacVdnOJc9zq
1zbpYOGqRd5tVo57pwJzvngw6Id3HFaxDvPKJCfs+c5uezU+ExAqpkwpMvHDidgYK2FVyoX8/N0H
+q4Oen5ppgX+4Svi61GsfXqB+45U0FPE0vnamw6Oforn30upLrJFr4JKGme1nLiWEypa5JlhETER
FO3QmA5iLADqsfRwz27vUpwiMtoqhzo5W24cg/fSwjExMru4CeYek3Q/F2R47crd4/TYQQkqmU3v
AXY/HrWblC9uX8QhTvwwn4xZW63nBshmZky1qVotEE/YB8BdSxh+gzBsKoxdT2nzcJ2qvEv1yP9Y
1lGT0erLYdfUHdAmAwD27+jHjcFo47NP5oRMys/gkBQSk9uG+wY5Aeql1/dIGa8e8jMMRkurA2A5
cqLMqzJFkJgpKYq2hdG8RNUlkE5eO8shvfcbW7DSEJSbVe6UxoaT2/o7QABTjcQxncAOmPsgQxZs
5XQDE5XHbaFOX1XdUOaE3g18WXfdq8H/K9MXouGm6fKeKzRTQKkHpQrXlijTJUA+pHvL/oYYMKD8
eBt6lOakNJRSv/TiACEIE4Jisf3ygxsQQ4ALK59A9+xGTnhYbq/jZWwYLeyWQYTjFraJmCQxDtqK
NMDai8Hksgia9CTKjIvPGR4ne+CUuQk/qVx5YPXX5rY7KuStQDGqiPH9Ue7FVJAMq10/HB3dhPak
G/KSDpX1PEQLyZk7k2j/QEx9sjuFP0mNBXQtNtovrMtQZUfVYN8bK7+SryUhS5lUJa7U3UfLw2pN
dvwaOmg74QaZdB2UXB2vOPVC+EyerQvuosTcYRVzCIKalBolFfj3JWnJ96s89mEdbpwgJW1yFWhA
u7XFoUNs993SHNb7mOdX5RikmLWNsevSCrKehG/kkhYibLBQs49H8WbBpmM2mMfh8/fwjuYpsbpH
ATsg7TJLHmq1CXs7MAuxosUlmqRkgzWCtDxCT3FUbTb9W/v0zKIsgVAA3tlskf3NGVvNht1ydE1E
5SCHI3O8LSyOuY/jGfE6CzHxymlqSrnUWVjZeEdkYvQLx4sHQQu/SU1lsn5YqyHTuDQAh0gax3Zj
2QTcvh6Oyj3PV2AO3X89xu6MHkXeWMd/whTP5mqvrtnfc5yQs52eiPupy/1qiCUsBGOSXmKBdLzq
Z5gIkeFUpfBEK19eI1+Tq8yPnclWYJKPsuihfppxl+DtuPqKTunmc+WZRYE3hRJtjJhz87NE5EqC
+3sUXk0pKDgG6J1AQxEJjX5BKhxmmdTk6yZSkz/G9REUAo2qFHyaRhU1XAvrrfZC5Iy61pE2Xvna
RG4SW1ksTCMNAWG605ostV4kg9MzkEY2R+g5AUwvvIDps1yAAKFdXCoAK4/ar/A45FqkUA4bhZ18
rx9xV0vDu2w+6yORsE8rJ4npQLmr+FijP6SV/uMoOeK0hTjdcbPD81Uv2LjDNPhfgs1DTmIjlPMt
o8PR5RmthVtYG7RGK6d6cv0N3nyJ02yhZZ8nl3FadsYKrWAJ/m/WkR8gfk2S5M0gfsbJruTW5FQY
GOTkqO4iZoxtn3EG4rEALTWA7IJ3yGsYZZ+U+/a6zp+/0tnSW/cdVMT8BHOJ60hZ20MNBzd0u+MJ
lPFqrx0XFI9dhfQYut5vyVNua07pqCKpTOirkNyCXGjAK/bcq1Ke6omynZXx6aiy909oLJ0FmjqE
4GPEhpWt0icsL8Uq4Vujv4dxFfgccdjbwCX5cMr0IU12d/NGSiEkhbcWETITa5XkQftNBceMNVgY
v/hN6YUQoJW7Pdu/qz+hAn/j8bLt+wR8NXi51+Fk6he3jipHbRqB0lOqu578U93QPKDFO3AbYvx6
8xtPGsXGK2DcYb4+VBdfmpDI5hDLF5Y5DZgGTeONWpk0zH/JvokxukfK00ErHqfD793klmwiyGq3
o6rZ7k5iAZwP+WDuOWLWythpsJ3SjZO5PxEv6ju6tW/8/0XHAPZAnXnoqse8fKiL5Jg1r0ZF+iM9
6fcU8wO+PgGvaq1+k9hSNc7admKDGjWUwbpg2W1LeamBNwPexUxPPnSfFubyI7wIGPIvF6iWy+H2
KKXarfDk5/WlRHXiV1QToM4+qhQEWuxJxjh0fe/CgKapbnV67Z+YroIeBuiIxqP1O8EdRUiOc3R6
hzeTh8H10CZLf0QZB00jRFCYc9E9qHUQg9wzKKZvkNO5q7FPvOXviGoZfrkxPwBXQ90RuDDJ5NGN
e02VNTIfF5wkZxRhwyn8MJgP+lQA4PubfX+VBB39WZkbgV25c/QfVtt7z9hY4Ahimfcs5bCpl0nb
dc/xJfQPogOMDKP7mxLpw+CrmOJ5Poef2w8eEk38/oudMbeWqxVE/q4CJggMPmBwZpvfN9R8ALh3
ubtZ+e5qcs4bRoISqyCXsQQ/jfcT2L6QUOn8nic98sbilC7nma0CiwlessmwWTp0rMsZ+sZmNtgp
GNozC5cuEpGIEoK+qv2BDU22RP9PFyiOb+3l5SCus4VZb6QhSTn8fjDfNEcjesBhWsK7ejM1ezFe
IwnGIKAVVJ4ECrNhXDdu/f6UzacI12+2dDJA2xyz6Eup2yxNsYuzTZLJ9h63Dt0vXmEzaYDhj0lF
sS0OIVCRK68yKGvEBB2awXmXUECVip6W2NADaTGubI7u65V0/Z3HYihxtfuVVxscUnsdMtyRkT4U
kpyKESNmTe93g4L0edELF5kQIRxUY5UM6KEic/womufII2mQXrayI3apthxT1oUwGfRk3U9FjmoA
LcQsRLZbtiHeX8NGZJAerkzGBO6eD7mJc3g2svcAwqcYmoWmThufhw7eVxel1SrgiouqVyVBUreD
6bstgugOKeW57ljg3a3sQ3LxSzYqvnPI+D6eD3lZlf3m9xqVkQlFgsOUCxiPp56knv1rctcpYLCf
xh/ishCgDpbSZRyv8qCHjzVHuYoSjOj+yuOZlboGo7L1G49POEQC3ELboX30ljCHS1tRJ7gdQ4TN
Wv1YdaeNSPVbTap4Bsfeqi2c/PLjnFym6sr5+dsoZ5yKxMGx+i7bt7ZfNJGwz5o50rbBwVYVQGoW
+XH/MFV9iSKl4vWQ1K4F2O5/hQC1jYiEK1P/MdSpuoIcQuq5Lv1UFgvXkdAvzM9U3nQ30gsSQ3yH
kAebzb5X9bt5K9CeXEYUFAqSe7MblAyRmbPq0pmZnDUust8hMYfxtkXix1KQYCgYGlkXECbFu04c
SXcHVNjCZWUY9gkeob9lQQJx51vE+T5bxRkuNywBz/xl8HUKH0IPb9fpfDSxWz2ecJSq8WNQRnNN
AD8unygUdwutXMvlaCjB82RU8Du4bkhZ+2U6le7Sgp1Wr3q1F8SdS2hUSbcE/w+3te6JwZtd4O78
hnOhY3lwfMbfPikQB8VYAnGZ8dbem0wJ3y8Asxdw1Jf8TrqXmr6Y5l17p34VtjWn68IKPXhGoRvP
NojS6IHSpylQSHh+5hKW8JfGLJq7C3Wpf/CUOn2044SZ3NcBRk0D2HO4AH/pVaSzTlVzZcRiWYm0
k8mxpYQKeb25uNqCtXngj3M5iQ8hv7k5akdA2aKT4GzzzAxEn8U6wL+Rm4pMhmsQpZOGD1tFY2ph
tk0oz3CN+L660+pkWblLaIhY8mB6Xy/rKAYPw/2CcEExY8ZxtRbXaC3yqU65MdWSpLSCJIjSGMQZ
bNuF3ob2IC/BYSVKXuH8jp+867veIy3PLD6LQww/3iU7QIX1otT3/jsq57lUeAXOKJI/CgpZ3hry
Na3apqgjF3cUx39WfQuJcwqxCk88eLuF/oiyNZG7/XD5FkVPMh5r4ka9r5XUSgBum4TK4pIGG5J4
161rv5acdPhFrZv6wnVy8YBfRJNx0L0NmK4lGp1BJfSvC+0pFXXS7wkqZvcIJwp+TXL/qzSUzX0F
zi4y8o3jo3YxoqWQHbb5o2q19ZuufjXcU7hIpiCUL8SKTAlaQmMi7UvO0EQ/dBlq239u7qDDFt0F
zALpr0Q5Ay4/+/VwShgCdBK3tIseEsjkm7yq4y+VlGgBvmgLMctwUP7jFrGA/+3nWSj86Zufjgv/
VxNSuRbua9X45RV+GegOvsGr4v7lk4rEeUrks2xxqNYDMlVNH/n2eLl2lpywinsEaqtmF8+t3E8y
b4pXfteX/KeFeE666OWVca2UwA3KBhMQdbztItB+z35GhRw8sedgXJ3GSdk09vzsSKpg2to9EbMB
xNuKde1JcGINv81l7NGvvsx0Ot4do8hhKwUebLqXmctjUSh7v4DGqySNlFLu0DZYJrLEwKjQ9gCF
iFnZQJtbGvxDLAuySuP+UlUFd4QNACJDORyN38/2vhqtxfeeK975vj/AqF8HfqgJrvW73pAP99cE
5Iyf7mpx3I3u5bgnDfoQ5gpLW0WyL5+OHKWwPiDJLQ602feZsZLOwE6cGLfU4wxPeTKHmkr8S2BK
Ty/C61iTz/MFcOGcTzAaqimNXtrJmKAKzXMFIzNO9C55ooTCwSNq2th5JnHhMSvi4ZUG6be77p6a
QOEfSdjYFEQeA8spiCeMfwtQgZ1aZ8GoIahW61VFhxx2EE6/lb2GneU4+ohStr0XRO4NRqRzVSxr
jzkGZhblVtXnoKBoXeK76uRDwJz+C53KXMKD8ZV9vxzwOklZLNnXLrVSDkdBALBJnfqP99damGNj
64dnwJ+bCV71MfoOsNIk7QkMEK80M8mAw/ruEro9PgrKaif06TI3Pls/UWpj1OdEHIaIpiiLNC7t
ZvbkQ2A9CEIDD32Dv5/7axNsKkFyWcUNq0fMwvgQrocqt1Rpl4r8WL//O2k/ILlDsJOaAPUUmYWN
5ZrjCmYlljNzLkgPLCpvO9J72PR2W21xPa8qCcJCk/tkUheyjO5mv+1iC64MnqTsFMOKH5FPYlPy
Ga193DDbZhdEAusWzYUZQlQyz5YmpY0F5bfJuShz8bG/10YFS05cQsAvw111h8xXWUyPvXgD1C9w
+92BweywnGp1SqrKElTZsK6RoFeSBMVQiwrnCYIf0AILk0eHeCLAEQNR6/aXvznTklAcBU0pQghl
0U14M28H55XML+ijzyFuwTK2pLUJQPofBvfKK3vw1Yr/2UziE+bRimw6vEjDTM0ZjUWM7PnZmwlt
RD4d8S6W1Dba6TwLQORm86tycjo0zRR9+HHvJBg2P1Sd6zX4WhJYe0nwS/pLiKla8RKG/Medp+G0
+g0IfMjZq+DFjGn2VDnQliLXIrGueNhV7xcyAqboU7WctX6GEl4iGNkgXewSiD9TJNnOmJ0paDbD
rU5D1QY26rvAki5vAhs7F3el0FxwJaMFgSqWSDKDItJg0jFxfkUVobzVjcd8Tm5QzpBwoHhCW6EA
7tJu9RxFu0qahjs0kKrhlmjCelKFBIkirpJ6LA9JBBFjh1Haco1hZtw7p07o2kksvH4TpIQ5XMEO
t6+4xs0mxOuSEajwGv9o4aRVyA2Ky0Bq6NcPNrwkNQNhq1awukdsVNCUoUUnZ/ovxcLqqoXsjbZz
6NGTzzbwKTLbaRFdVSZDTIycqtMCQ1XwIIAedrLj5E+68RJl17qYWg1hgTousRkm/Gx3ZW/uOKDc
VR2v+DAk9Tjt2tqYJj7JNdmlFzGt1G0GJG3He6nbLS94Ji4TIMk+94LGN7KRu6qbKpsfjv6tuiTJ
OlaSpI+1Di99Zs3KnT5MiAafhFgdJ79/hg0YfEod3OnJpY2OHj9O8kov7YLNvGGHZFzC9UiZ5T5V
HJsghn6RgeczjnM2gilk/qBGgHciJ43CG0m6AjeBsQG90/SgDkeVt1PFczfviiqMbeCdeSq9cGzt
OBr7/majNG0X9Ino/2MmJo/6LLZcCPSqAu5sOSRjb4khjv42r69xwfEV3T7ZtKtz+O68y7oL6nWP
/7vJexoXVdoE8htuzlfL/XDVAFNnmpPYhkRDEPLxV9Z5OIm6Eb8EMYQzF0plqLI/9qcghvUL+Ee/
hwJF2odKFazn9ZB8lIqURmyzWrqkzt/2k19e/KSOyvz6JEngsm9TOTfAPhhOSzJTBwCG79nJxbj0
ge2h6Db0hWpFPyRn9hDtoDGzCvdeFR0bfpG195JdKH0na/ryeP8jOkft9lNGNBOpEXfTHdbIUd7o
4M4cqB6+HFe+FGrT3LiyAuNUTuBpoMssXTcXdAnkukSrIk2hhWFuz9cw0y1oJT1h4al4NOP6r1ga
dbcgU5A6U+8+5JEPQxc1CW0lDhoWe8a6SfCAmHfLXt7OPW9QMN0l28F/Y0K5oHWG1sVNFOYgElSL
l6yA7n5K8DOViD6kIkQ/tDKRL4DFfTqPU0ZyUa9Xkb/y9D5FaM5P9sEXD/JsqBxZaLw9iN4O6Fw1
dkUp6ux9015HvZT4/j1pU0FJofBxF0ba+gtnvWxH5pZz3ayZwLOW1qg8ve8DJMCvZlxrg7f+Qlel
lXC5YYrmNFi1sPa7bpbpGOrdxUNlQa9/VafGcgVm8OCwqhh3LEyvcyiiJ+l+KOUvU1TgtA6gyssb
X5ub+JfSvLd8Wq/j8Fn8ct56MP03o14MrW0VfeUQUArgeE5BdNh9nvK2McCqL3TdcEOW8clRGgbu
NF7Vi1XIInEqJWdYrTD1lc7xWsdLhY0d84iVJM+x1RjC7d+y10uax5r3CLOebnoXF6rL/JxnbDX7
JTAV9JWxj+syH2AWUoyG3yyXjwp6di4a3S4oBQssX9zLV42vhi9HYRj7H5IzY5+u+Uw13xorRRuX
aEWKqMU3nx3IdjQXfFfgVVCBwPxa/M+P3d5fX3HBamDCI8ZE/DgSycRxlTIxWN0pdLZL0VcCLEay
fkxX/SO6F5RpwJamgmL5SCs28IXglFo7FeB4bM/GckeDKVLrY1fZg0f5XRwkcbp4gDqb8uPNQSkA
PWrX/+tY/c3nfVe67iRm+rPGf6ynRf576DUnNYQtgKFWqIellOgYFowRTIZJnDC79N5YGdeXg3Tn
y6UpgtQ7VnHQo83HB4MMz+ir5awME0Dgf9eynglpTurSlD8GPu1bttBMWOIQtLV8l1eYKBGsEevr
YTRSgqYPnUS4Len1Tf83/u48AGaCjmQDBWDCtp5YIQDXkFvPbkkyEnxvTUPgJPkNyeYjU6T10Okq
5N5BmD16nXyLb1u92ThQX51pzBPZLrTO43mMQTlcJuGk42Xdpl2q8b5SK/FyxzMytjSG6cCWcG2U
+AWizm8jO1gh29n/j2W+wJp0oxTMkQ22N7qWyzxYDoz9a2XxTBYGOjT5KTm8zHuw7+yrnJwZdGjf
fp1w+zrrAH1ZY0s8XrUT6vz5R0Iog7VyqXrxWzdT6XnNlIIPUIO5vDcA7kTtUba8oTHgCouDarF6
onlkEnfe4n7yHtf+ng7ZPsfLoP9GT0EtlB+unAwcOKwZPloFeA/uHn7OuoMN+pSgZeO4alCQnlae
mLBc0ill098QA5ot23GFPSTGIa+rn/3QjYrH9y0TNdtzK4MW02+X/Ly58bsM7rZ6LGDIEMQzVr/r
uNxwgtJdekSMYsKA1wbRBqNIhq108FcTFqiQ68CxFQfRv1EwaSryF1hlGAbQIZyHxNgb6ky3dXet
Bjt4CPOSimnQP4cNE5M4x6+7NE/IE2+N1cNYh5JPITbEPQm51zDX7+f732GexnKKZ55o/k3uYTuc
0K9BFnXepOKWuAJT7AqCxkWsdtV1tfXT7V4Zo1oHq0x5RJevvPb5Bx/RmdFJIwwwOLgIy5kXPNwh
Oa8zzYg7FnF3GiQJZQLpHmbvKrTMY2Sm1//w4wStofe+tnej9lA5RfuxlG0DhYUhVLzoVZdkvxSE
jXeDPLMqDiCzJXnA2LIgjzmBx2adiPYkLKWIXfdKqd9pBX9FqaUfOUKXqM3v+fW6EFkoQhmNAbCK
ltt5UU0Z73XN1DNgWMa/TMAoO9lYwrbIbWLZ47XVxcK+W+e5YiZrr++fZ2nb3HSi29emwLoArM4o
HmzL+uFTdpI5Kf+uZ1EtSVpCDO6oPdHTZtU2ZgpmgO+AQxpkZZaY7fbi1FgCoEhMPAFqnVrPvQG4
r8x1n+zq6WcHfkFEtivkAhpxv7mY20JW81ylTZgwPj0HXOCbwUd6UlJLG9RhsVlljRczBrfxHDdO
prKPjSnG7NfAlMz2R2d1zRi1O71HLm/SjEsTaq6o1/VbOylhhLSBFyuj1b5J6RvrK/tqmoTynTJu
gn9LTxgVYyjAXcTtL0G/pvDnaogaBOcRZ98K+H8ovJxX1CCCXDN2I+Kng3GEouCGYPaLBXaFjahR
d8Dnt31KOygEbaJ9T8t9MLAIV7V7hi20C8Hi1vyH0rlKhezyIDVIa9t4j4LTVikayQwMf2Ri7CI2
c1NcL75fSkpfbYMZpy0bOKHBdwdW1Y7cTYb16dRm80AAyRtUomTOMMPoDULn9P6knJIwlpuqENyA
N9LFxYGnlsdPtoMai+WgOZquPjE8x+yX9ZDgNe8fhT86gg4WZGnWA7lPKz8y5fiJ65AGTJUKfec/
WQ3gZmLTwhThgO6mnq4wD0oVA+1SoRt9j+94+gyiW77uZ65HYsz9TwU0EvwU2cAyljxIGh8hL+po
lO41ccGHVfD/xpU732eG803YldUhG4s1QyBhIZIRUIkgbyTyMPw4QKcFZvoMuylbSH8s8+WScnAR
64alNhUzM5/35z2ku8AZVhoQRHezNZJz8TURonsQjVMX+VqC25Qye0lDtWZzHQer4uwmG/kGc59N
5cwzhLCqdET+RkN2gcbbZYTwQMCl0Uem9BffL/bLPqZQlcKIim09Khfcb2ohZNklaCJYHNckzA7j
yG9WoUJlnSv0vGRDtr8isLPJBtPhjMRZDHbP3y6s95cLu2e/X/Jk1rOznNdzW8jhm1TDiDEJDN6J
iM9NQOntqiZ9QNwgQxLSRHPezZ1TApzIa0aBra0M69D/+GZjMOCpo6VEa46fb3gTOBw96iYL4ad7
it1zpob2CJcXU8qs2h/Eefy9qOQF9vyXmIxypr3lbF0eoXdUhExHLSeFw7/WtZmFSsCDQSmCEYjC
hWNwyEJtqL8tis50tGyjoLnsdeiHVFmWsC1NX+7YbSlHG5//JEhsD7m4VL9n9bTG0CYlNrZuPvq3
7PS5OeZwlWX1Nk6OS1lIJRryc2qzK2BIqsgPYDdlDzstbGwOJ1V93d/3IasNlRGSFyqOQaVbzKag
T4+XL6+Wm8iFvuJxO8CoPUEWNHulNB0APcrmmVgYxusDrffPMqCZKoEUNW637IBforWAPJKikoTG
yMwJA9RjopXce9/MxvsRpv9EmUESpN2aSzIHrWKBwmSfucMbPQV6Qpuu6sFGuajacluXI5K7vanf
GhTbB5ccatUgtYVZViVE9yfreNVQH9WI5xCi7uUk8EiN/j+sPF8yN90cc/wWoDcfU5xKl3nK9oTJ
l/c2/eM51PcmoPyoxba7lLi1sWI9mmnYQYPw4wa4ZOi9HDq/iGQAFMg9M9PjJKdx0t5aUOxugvF6
mu26paKaRXwJkvPmNFucm5jiS6GrPj1SUX+GK5eLTONmeq6Y8aEyWH/YZDMEHbRG3F/WpXTaNbW8
Qx9QBwjUxgl4VjFWC4NJlV5GhjBgDi+r4QQRyOdt//ZsLY81x8HudzWkfQCvuY/WXAC0dja3QSH5
6Qs+cOjOTWi05mpAGZouMfSZRCy1Tg13/sJMrrOt4U5w6CbPHsRVvIyWMxyLYjy+TJxEm8Cdf3aB
6fXQKN+dwm7Mba9cDCpiSIHYkW1UJ24LbKT+INsgVXHyL9zIcjgsQBKsYw2SXNjrLCfFcPse0LTn
UkzL4vyJnFA4822T6qcJ7GLyCj+2TC9elntJhFPOl00AFU5MlryPNbVeaOfG13AUxMgPbcdwWDdE
vc91db6imHGUXPo7ePSt1uXEn2G+pNuqnbym4CdEjO67POkayd/CzbRJ1CoDzY0wztIbwVH7XXzK
J5ICHM+dMudtY+qCCkP4kFcDgZa1j/aOp3VPvIX3XtjP2XsHgWQOsbu3zXPDJGnRWV4EyPOkhf8f
mwm7VvYZjoIp4BBBbgYOYxqo2fgAjzgAY1ibNoKNuVKsvcgKlmRt7bR31+I84KBK5zmmatHdokQn
NjR5wDi/hcLJDBhM8ObGxhke90mQkASsEVQxeZ/tvcvTJNxguT7hMhuE0NT4MAa7lGDpBuHIR9ip
1aY8v1p5hbAyB8jhPL9zj4AN4haeUYsMZ3QUtDurw8dKrnNt8dwtnj2Vo2o3+vQQYfROBVvFDlMU
d5CKRyuO+TJ94KHFZjD9i8kaWqBeEdtWc9mfnvTKLrfbveDu3Cw8pyo6eUymZo7Ql5oaMxMIbVeY
TzOaQ39vS95Cm+Z10NhF4FkMcLp9ak5fgSVqGjgQ8ASkBMljd/KUnpGirKY0xwvlcDfDCpc4FQrT
dkaDCS6ts1vuV3dOScMhqTS/wgZyxeSxTcWoXHBnUUtybKVcjYdTqp0D3YoCyfP64mD8j0Lu5FwV
DfRaB1piEBJN8vM07VPYfW192cBzynw50uuwKty3oIdLl5MGHKQqbaJyXsyUQbZ6yDjeOb5TenNA
lRkuGLuv3wP1NneQ9l6JEkmBkZGi8bbyHDtKmDTiNZ2sREIdtXIjXStWQzRCf0eaRJxL7M1Qzp5c
plGJf2fmG1dvMYxy40dB2ZSbZKeVaAXMLTYq68lunHAT/KLUw5VZi7geC/SrTdXXrLRs2cEMHqi/
ViO+wtUpf+L6sb3i8yOqkjscynMB2MRb34KrlH+fXR23ie7Xy7f3MDPD85GKJgvJFfkNcn5vAvU8
tPoX57WgKRh/arEBjDksvWhv2Dtc7gEiDA8QT7bDrKJljy/ODQt4DmuhE5WUzoCiv1A1YUzX6T1g
UwxM71WMHapp63FxUQaAy5Jm1v88rXklz0aCNDH+iwh/bOvJlhlAckLdA493niI2yNl1mTA+qWa/
jarcG6TL3GXKkgAr5K2OBq5tRtWVRw3ppk+VqYDwhjHOvGMLtlKJ2jkE8ZOQx40QF6eMQXcPM1es
wNG+8RltGaWJwhwMWle3SNguiDe4KaME/qJ0NOfOH/IdT4DeePWPYibkxpjM4sTk0/RAIpQiEKYw
xHvBLG3gtiHz/lM730YbtvGkaeo6st4+wj703gHV3T/Bynv7ADPWsUUixff2a9wDb4VjAPq6sHif
Y6Kxw1cCxNAD6hVuys7JJV/nVvt93liVp7/+ENnuiC8/bay7CcSzAKVcRUPxWBd8jHw5lE0DL4z2
UJm6FhXGPDujjrqhYO6OHMlZGkugHSFp89Lk7Qx7PuSNrnl0LGkRYcMUk07X6HMmozrkxVxqg4r/
4VRvtuwYeFlYQok7p+Al0tpQEMXWcZiEwtASPWLCEf/IwyekJ8Hc6RmqL6OTGWJxABkV7r5vkEV1
ttUe0Y2KY9/xvAUhC4rCiOllzj6c8E5ew2nwDO7ITsQRVlxsCE1xrqi+ZTxlpz5cTqnVGIPoPTO+
8ConmRhPuC/f9FBcCPGScvhCmeLp4OR+Dwc3OLSLZ7eZ0fnzh/XDJAMr0XnsrF3ueE238wmEv/la
zc0ya6ilH5JgiunIA0ZhpniK6jIz9H0llptW//7/tC7vVnuKiDjzY7MKKWvVr5qNMtgyWcSyajoJ
/aVn0m4m6ZTsVMO0V26a1HNNLUZ/68XofkxYvfG9+iF35UJwB2D8hyEOenq1H+wm24o0GPyzSXWo
bA9zgngRd0jvg6D4ARuYho/P8CvqSf9b38l6oH+3xQsQ28GYQHywwI2vyYdhoC55ytxqfAqXdQPM
31gURuUbk/XtSqThv+CH7zHtMz6mD6zyhX1PeRNYl6IWmIjG/2zMLMJfS5i0Ek/hPphgN16RPut0
Gd1otDntZpy8bG8B8+glt4y3bAokubtDg6vYCbdcaKT1/Gd0imE58O5VWm9Y3UYwGtZ51Jy1laKq
esTvHZ87PV1131pOimBB3NVtGI8lwkVasnACrueVob+pgFXJJe5/r2M/Bz3h2wq2dydzwtOtqZ2C
othHL2/4huamS9k4+dTAE+m6yyWPCJMbtelBQPHTEPuBOdxEP59YGhCj5mNLAAKbsvKuAxlDKnkQ
92Eg54bJkzt4gyx0IHYrBuObpjVWEc/iSHSNuuuIsbgTb7FeN3Kot/XxgyZOPlqVEUQe2X2iJX0T
O50xE0rtZiRAWAIaKrdXW/kakA/w2JvpSjx8dL7mQCKutgUoFRX5ygqu9PhZE7b6V12Uz3uhZJVN
f/H4LTfBSEFTHz39PsPl7iUM8mLjZLZa30azDs9B4aM/XKfXSkrLk7nBADvTcdy0kKtyldimPveO
B7XEWL/K1znP7yetMZ8ihb6+Vk75wmuTl0mP7LXDk760PFzek4zCkB9BK+Aa4rO8mGqJj97TY041
2JGU1jI5Gk9NjaRvOzZoF5iBWa1XBOYR0FAsg5+h+KJfC+9Iq8xovn7/nz5FsHzQLZtSvW4wdeYD
kIuvXT0zHLiM9RwZVCmNqQwIs68ypT3BvOLXXCe8pftA/NUJ6BVAuJJ39yM3byvOS5new7LPp/fA
VUBC72jQROYvG+SUA29OcUX77LRlHzca/5aNkV1/hK4DmYKAUqFQJUYg8B0oTW6R9gBfFP0PLh3B
T0GQURQBpJ/B4PuZXW53X6iUF3r97flwHfCGrfYt43m9D2MPwgOngegiNOBzsrdWM5yyd6eyy0u+
t8MnOUNGBH2d2BYWthSIKPdGSQQbb87akDO0MBnEC2Xzw3aNB8zGCAn8EbAEFOWpFPlYhs7bL9o6
Jn4HuYl15xOzit93XD804mmrVTse+heMgpVleiEGtgO9avvIo1sXxApNQQw0sO7ZqkexnFCm31SR
UNzAAyF1yO76InDICSP0AQlvTTbu3BQwmb/0gZ/pGLHQsBRK/87fKxdoO3p79WVzIGj9sKM8E8Ar
JUL88nIZ5jeH1uK+t7J6NRSMEXOnXdcUH4r/lJfR0S4c9tyALq0ZsZWIV4Zrqupua/10LjI9mlXm
XbkCMOQACXBu1zTnmZUdXL4JsWkj4zhXCkWWF9Z5tV6lTIHWBDc1hsF4cnKMMQ7uiWQMA/uxn/5v
bDZc5iuDjmIjC9YimSSAu9URg98P/h084lvfRRhKUs9VNo1qm3L1K5hEQ171IV6IsFp95XG4CM95
llZ/0Tfb6u9Zg2oIUARWoLoxtDKxYEqFoTZUJH+n5PPr/bCrVl8ZIi7o3qXBxlMbVaR0GY6DrH8f
9s+4OuijvNqnaqyXdwVEdo9p0xdW4ZDjKZEojnD6Sxk1kH44sExIYwtoX65r0kosx+JMFXjzsHLo
pGeyPG1mwVlawEjposkJqs9xiHOUX2sIFfZvqM2++7B1T/kcnW+6MSZMg+F7+Ced7Gt7gj7UzYXw
YP51C8Qf6vhATBVglPahnVw2gkFCg9C4mhWuszaAnneEiqQIZMbzvnN1Iuqrz0TnZHZC3iycU93A
/S9frNKXSFL5J1uXeZ06NnUc9noNiEBSiVTdsN6HAn/fSF/rBlA4gAaO42QaFCpRfXHrTqxFLtCA
oAWxjZoYoIW3t8SZ4B2PamyyRzEMtDZbUOkmPnsota562qH5H6mDNKi0t0m+7B2JsLJLCh6tr0lK
bvf4LZnOEWmThC9Ru5qfZV5I4fpK5JNDdSMRGyAP+U6xNHCzfXw0bgnGsvtL8Ftn02DFKWxdyYoa
9QOnU45Z5QXMCpeIduthIlg1ZUg2kifBWGNlXPjiWVIUbTer/ZO/4qdRTjNJadOFGXTeg/AEQ7//
jwWxgFrRXElydtGHExU9xfzR/TQ3ApuY7UZgPqzEcjEUZixthMhg/XNW9r5ViheQjtFD+97A3M2M
b5S97ARxXYrXoEPWv8XbWFa3wrXa3dbRiDreYVBudjgdZrWlHDV16gudBLp3jSs+hcC3fovG4vRi
Czft8gEFslC/ZfI2uD5TF9bq8BhN3dCBLpCZpcjgPlsnkrJ6Kz6J80ytNFL9PC4e/F2d5i+hu7bC
Qdu2uLzOthReAyG7m3npEKh1z5N62I37frPi5SDqFpQwla94wxaHYhu/yYbnRa2FhormUdihVPYs
AAFwyYs7g2gz4imSKPme3yTatZeoKgyJcdB41SmyK090F9h2hI8VDotchLvIIh4xOoCnOcxr1xG0
lZBHfh6YAWWUi9pEV5WehQLGAzEdq+sEZbDu1M0PrUAE2RhCnXMgAoMSOFhghY1YDmz8gcwN/kf1
fXZE8Wrjzjg7jfxw+gcuLv3wGtPsSdn2f8KwnZK/KLxCmWTnHMS93GRqPE+OMbQ5UD9PvWMUQLIf
WhqeoFYhYhQLcWva5Bw7XT2evTSg1ndHByZjVQb0HTY4br1e2wUXFDiiNVEW+8bE6p7BVfkRMQzg
JxDKBMHXKusGfROnj1PdBcMcb010EvModD7uLrRsJqdGgKTgb8tHVjmDTuqVWE25YabItLXvCOYh
gplGqm0gGtz5zPY2KNbXbjDxhNaxD5JaWFe/lRtaI95efefcmTOMG1vay5iR6kcDSWSn4oxOdZBl
T+ebxibab7licfiXlHCZrAtUoU/VedZErgU5sooxNz/Ko5Qr74QSOyjTZDjELKwKh9zo8fcorB7J
b2X11zD051RzHgJfAZfVIItgWHzQuvPzaFJhpY2WCuSeZRaJQa8lfS6lsz6yZ8hz6fcm3CR+zZi6
IjdurzVerBh0B2QpY3yP2qp6Sf9KB9DhA/ynLZjVE4gpohbuiWc5tKWpENYajs6JYRs4rYIdBeWi
ThITgnyVvXzhQU3d7TCWbi1ltNrGaZkZ+3wsHdp3HkFes0jEqukaZKubCZNrA/zEajjpsbgM+zaZ
BKLRL2LYVbb6d3vzuL8xxxI0AKBd+1iUoUTn5UyYqR2CdSsot9eUwyHb8dBC3iCVR/sJV5AWsh0m
3QXHNJ9a5UUAAExk1soAJwDWAYunYRLjpA4TaMuqF4Muf5wxx14Rt1dUj8eVAiuI2f695YaNVp57
emL78BjpgOHKAc/EQX8TDuaDXLxfAfKlsgeY3OjJWYR4da6JTpQCxHFrXYlUCGwqU/zMkXOEDrde
Ps1lUE3WDOQzVJyJGFuBPZVYRd/caPMbeMWPjoAEyOV3Dezxil2kQcKMr4zSir5DxQFkEfJbmL3a
gGqNRElRdV62Rps3gNzAqcGbC8asy+iZVuZcN+lxhsMhefVvB5AXeEmEvupbDMoWzy3tZ2Y/PZdK
iIygx31cIByEJcKRQlx1oRuDLPwHmoAT1TsakQtYFV+yiNoliin5Ajy4mUOafmfjGmdDqXf9sMwo
hsu/95www77e8hZJRFX/6inIDAFvHfJTfTymUVWJXaB+zGfdw/Awho+Tq44snXJZE3o7MS1Pj9uV
jLWdniOLINcArmYpNUC303qIXqM6V4W77HJXawNaZlHWJPdc5WiYB6ZJDpGDazhOI5sbimmgaZdE
u/5aYOHf9k8URorxfJFEb56oMqP+TDwAIycWSKWHoASlglpbqsRuIpH0sX2RPwVoFxk5wvxT4LKW
YguZaaNqdLcnKvuSgMa9ax2ZAq5ewCJlSEIYjUdTo+cbSdh2kWXi6lIdbFeN84tsmSqddNLfVMXr
foz4BtZfQ2X0IJ2d8eeib2SN4hkdZv9RDy+g4fu3ldPIIaa5Qjtwg7XWzfH66A+dS4M3ZgOazhqA
TTfEAUIAurgi7gr6gYUWnQK50NxGEda8BbdjAFbZ6ZJ1J4X3f621SuIPrubkGeFI96QOI/3tyPx9
4U7dAqmA/jFUMXIW2vzDwXKnCdpiJkmblZiQ1V+9dAqKQIQQw0bbVn7bDbDlerfxxl/AO6tTXsSD
+9nW4DobLsksMMtnVSXpkuoCdtDIVjLe2anwi5y8sk3CaHyPDV4Lcz68/VLrtQUlDkc/2NoBh6r/
C54c1xFY8snIAvrCgT3gn+atYAVrpzC7ZyM/haxjr3+E6rcezxtYlNFt85KmGiFkOCtIM1b7nVHE
bNnKRtIZJm0EroKPELAeRWv6rHiqR3QB5D5hoEBbIjZnvPXugKknm3q4SZ+MEAT1x28bMxWvBvb6
mFNXF7HDPc7BrbpBvcSoLh+YpjuYkJS1b9S3zkcb/ZNM8J9qoBOvR3bZfuHuTEt91An/U9c2CVb2
7jiBhIL0La+6GBMyVxH/VQg7YnrBphRw56Oa/HlZ3B4g0zvrmBrqWDzrqqW/pSGzgRmcAIkDwCL3
Fp011Z6XNFlpwcRiiV8QjkQXXifFpoiaeUcx1kOT6ytOA5SQ8o2L0XaK8tl/NmifHMepjKZT4u/H
l+lxU/zVEyQJmWev4+hkn7EoKiRg42Nn2idzOWYtExQVv0IEIAoIWnnt+Bh50OvmBB/2ZX+YP1tB
28krUplohsjAYwEyO3/F39xfLCKWEuS8DzaQuOWCqXv8HqYSM5SIBDdfD0gMjorcroGaKqw41rnM
bTjPWAH/nwF7BNJdrfXDqf4paCZqcF2sP8dCLEUJ62s0Rq7ilMmUlIKTft42swl43lGhW5cgH3O3
x3BFTz6tMQf6FsiPOFlbSYyyRNu8CmuhnxFq7dHNiXkZEH7rzVBylNSOJJahf1lnHRaN6paPRMqR
MwzP3uDH6MExN1u9KyiQYS337Bl57Rs50bM8in/ktetWBvzyK01WCitQQuQMWy6Zusag8+yz/RLo
iqPuewF4C7CtIyL31GLIUS4MezQqziceV+FCY5/hweb7HMo2D5udeuyxdp9ZbR6cmYRSHW9zw02q
zWL1Zb4fhjC/4VwBMHDB6uREZwcbzrKb9QoXAfkCyuMFQqUESWhMiRzthJhdzPaPBhPGDkltmm46
sEscX3bTXHVo+6Y6CRz3ZBxsSHFMt/CKsw/mKa9w22n2dKh95BeHfHrz/UPqwJCLTJOJGFerRnNx
hB258bG6IZvi46RntA/4rw5/I9zWoa05JdAl8+f5I2vPWGBfjnW6X088JUNRRBHpUeB+OVWSGD3m
KpRa7d5XQDNcC/U1NafeB0NjY1jF+RPbedIkMdnE0CnJ2Ez5+k6VcV0X7mkbZY+5SvEPVjdj7XSD
T/TnKRE5q6uABhePJR+7+HMEx1xG6rLUP/41aDdLrMol3v9BvVfN7rUboZeHls5e+MwdQ2ejKQPW
LeQQ1gGWF8QpETml+Gj3uRJ+B67+1UcYHClHUJFkwIIe/eXw917gEaI20jNg359GEEHNERHONB2N
n3XubKN9icIS+7B0IadIAqxDZnfXhC46XJxndgq/TcPQvFxNWfzkRNHUxQ6QyizQ2PZMCymxqTcZ
ZsFGms20mdChkLGjvsKhkHGIYuik2jnsBNAWkWZnwbphk0q/NipYtTTro4CFlXPvbmBCACYqHqe3
0Jl85GvdSDaTFNGT8Cd/+JKW4SziMmxf1kLug7F2TWkYlsUGTpa00Fig9zCsUMFx5yvPNX3Vs9PZ
jOhybw/F1+753qXkrvQ7nHyAEkCADN5UUfD8RCQkjlrFx3KVEAzwfwdzk43ACIa50Ic1mJrIputq
pLmybu9Ky3kLoGDZ+B5yX3NM29kVZ/ZKffgqZFUC9GVdgo7NTinO4W1YgEB0Mj+towtQCDOYXT2R
b/0at3+chWGYHali1OZsyRl7EQWtyf64fDrYOar8hkHXJLcv5CI299LBbt4zlGu2xcLDVT8YxL8K
FmGq6jvJMVZCoP11Js/UE4FCuun7chHl6g3mE3FQ+8LfPVPTA3EKJ8CxDJv1m07yrvSud+w9LAAr
GJVUgtxBs+vn+ZPF7MBLMCGZDI7V1qkizIPTiMo9Cg8wZT/3z/I7O5rPQSIu+RyC66Wn4JTPFYY8
JqomxtVMY+4ytXQJqajSaF+6DKT5p8wf0EJjNh73vPHcbd3sbJac8TaY7SJQAzJvzFhCqj+gSdPt
fl4M4pQ6QIr7getjfgFUigWQDxzqy8oN45LuB0dvUIgBtKjWhNo/0THmzwGqxI3N+y58EWvOuR51
0SLqSaUlFck7Umfpq2Xi8K74AFdIz79KN15/Hg+3uuHfUM5iBJT7Fg/KYlR362qr8wNfrE6qKQDl
CYFz3O9yXqcB1frpLn2WfU4hhoRPH37D1sbyl2r2JLV/k1Zwya5Dkma/m0zesNrbfv6I8WtczfFQ
pNL7zmktAt31D8ED5XPMpdmOe8Sp5OX/91y26HptfJ0o5AZfpJHRqcgrP1qrRYNe2dRX1ot3mWHQ
8hmR4Umis7UMuEoLwTEbhpP35wtS8jwHZ+24F4c9gkvHKu5EWJYs1VZESDfEoG9VzXLtF2qwaAb2
iZXpWzaWkxpjWpZTZhq2xQc3RGb2XoUebqa2hbQopI1jVj2OVNt6iuYxJaLH3GD7meLokAuQEUau
MPQHhSuqhE5OCW5TVdm6u+vpH3agjRXqvVXPUu159Rv4dZ8DjZvkydDFVPuHX7AZFO2XyRN3i+QP
t78C183SULjoommtF09ul4QjT17/mashUXA/ZDaxj9uzNc3NAup0/z2p9hGg890IkEE4JIGQNb0n
1noxpgqxViAWcs+nRalTl5UU0O2Wz9OmFb18k7BcLLI9jzURWgh9PnUqcXSyH38eAo9DnnMWhb98
2oBOZK3O7DCrleyaseFZMxPDnrwhLTAlHk8hJQ/XLVfEE3Bh89Qn4VPzAL3DtnSpJjAjhi7xBYvZ
0aMVO5/tHIgvOS3ZH+0nx7TVA6QJiUzI7mSFAUPC2vdm3ITYNHIwbLrmV/xGAAV85Fpwn/aT6EL0
yT0sgzzPZqVe1R70BNzhu5X97duUiwAJcV05r0Xl8gCTSXjnOHoFMeo9oEgi9mdDkYaBLE0rIz22
FcuNyfV5aZJwvRC3H6VoqLMte60N9mF75m9xFpUkrFOGQyiBNJfuIlOxQQdT0MxL/eEHeMv7SPMM
gUG9MHKNwYtsqPk1EOvnUCPxpgRQam7JSQzqX6BEu4uzpV3hn6ZF/856mhCIsw38O+NZeEmWEtU1
CRK/gEqwQaqsyiqZfCIjzo+hKM2WLCmv4eaa8K9pSxCobzzrtdbyuAfQkngVElJIqRLdwj8zLLeY
GhpyYlkugzC5CztB1MpWMy/gBK24MaSJWSyEQL8+mVK+bkj2YTKS8ptnavksEIbOLhqcqK6RhLmS
4uzhTmx8jRKtYb8EeecisdSCTmW+YYD+x9XP52esKv+4/GPnGGT3rl26mA8KQ+0dbTsKWD6BiA3S
RSdaTPkcCwPy42oYvhECwcC/Nhq0phxgA692DGmG5ZK2FrOPHmiLC0kfxedSztNkSZgsSFxIcUw8
EMSWSkkMDPH99OMAHpl+AxQMkyLsA/Ltuu99NRWc/ItQZ9XJU9vvK2sw6Kfh7QHEB4MFlxv/yONL
qqwu9qKGTVg5hx8q9h5qWGLWC15jEPaVVXrRFMx6gych2cSHqc19GqbWcQalnEys5r/H9ezJ9Jcb
HfNvoOqvf44IcYRsyaP87aykHgF+vABR2aK9XyULLr7YXBKfqbgXO9eRIb90SL496byWvCu+HSxi
oxOVV7UQTrJILZIbXG3GtAa+1OAb8s0dRuGZ8jrRu9PZFpnn8SKQfIED95lE4d6/sQCMb26hwVsp
B2kXNMYUJmDVDkH6oVzLs8z3pAPBI0e9WFpkRHPtCyzebj3GWOyB/L93KzWqbpJaw3oN5rIDkLIN
+W9yuRMkUMPPoD/l0/6Lq3L/ZhVbjqAaDm7HeZsKQdtNeIp5tXJ69g274aI5zc/HjrgeoGAch/iY
xk0EQyZVwiWpWkB0kBzCGgHKsnjTdDXddNHMr4zE8GQ0RUhPRtyP6sxiaorPCxA4pIvnrxVOIetN
RFclLOxDOeRAtoY5n9eQFmt6WjlMfWMd69oD6mhqGcS8Bmbd6tLJ5Z0+MG1X9wbo/CjJL7CF/YaJ
n6jVuzoxanTiZi+zeLqHwhluEA1SbEYBduV+hL/ca6IaoJqzHbRDi9woowRbVBklUpCwB08F/E8A
dOq+RajOPTQey7ip9XMRQI8Mza8VPN+DAmNnKTEH8EXiwycdLEkD9ks61i4ISzlbl180kF+GX57/
vVolIXQDjszz/GG+n9UDHHtXkNuouL5dJnFnIQtQse8a3g4lRvFhTMBVrrYWRjLKS55q9qWKp8LH
3n6jxjtcbUGs+y1okoAaP7clIkmnMsFddAQk5pDyeWMKfrw5WbMvVjv1vSTty4MrgoAdP9KHIKn5
SaWl+g3A86hY/EaEyH1fp5HHsPonJ+wHq0bKZ0TTLFnrKSll+k5gWb579LYgn2Xz12vexS9STa8c
srqI07ybtR4pgpHWkQvOsnxiRc3ydiIOEyubqRg0EmLTpuhhVKc9bK8xsHVUQLb7TKBRKwsvSgA7
7HvPXYvaURivZKmcVfrcz5d9f/+5igc1ho3GRPrVMj7f6K6LtggsTcjWzsCZSHU1UTeTur9p6VuL
b45/nquZ9F6IiNPQT2iGJwdn1uWfTpvtF/at2VKREA5x708qd0/inAk410wym/NpW8jRZ9JlPQny
jT1cMiqSVduugRwHzzyzoVjI3Tg0GV2UHnJUKRDopx+GIL9lhCnJuNaSvR7dsxJwOJTZRHhNhxBq
yqSb3Vy0WDCiw0En0m6h99vTNDxsW5Ag/Xfy8rRB18fOP1dRMYNx1pjvtULkmLirL4qJ0Vm2KHlX
RHwSXU3dVhd/aqep58xUTZeXJlDD6PzjAzDZ675gMMRI9DQ4i4d/YxRQzFibQTEGOiBX5orMPJ6k
QWtvVGzRb5GPV+1S2ri62yPHE7dvu2TdzD6XCOFs0p08Dq2KdaVXlY16WIYbEs1AnzOqZO3A64g4
zF2H/sxoclgKZ3h+m+modN0ybOKE4qkXceu/++ELNOcZfC2Pxt7naQco3n9Y9iEGEl0QjPaoNdyw
cRQ/VStyCo/Myys7KuCnMM+3w3XHprt8SpmGJrc3b6v3qE/IFXRHrJgYlWzoVT+/8AMemzsOKSP+
6gbu1/ktsy81+Hv6D9/GQGhp4/e2z3Wnnrx7oDA3VqkZcXP49ab98CQzc5N0LItQSG0RpSU+NT+A
gPS6AnL+ANtmL9nWR5T9yFVuCTsE35qK+4zH3ub1GMEKA096MD8B3qVifJGgZJ3OySVPaiPHlTFe
M+NYbyb9DPd6Vv0PyZJs+czxm8azyHWCV0NHug7RU8D84ZIHg3u6WdcVIuFNXIc86WuTPGvVfgvf
RgCJw8zJOLgFPP4F01xq1W8kzs4J3xk2adNnIBzk1ZVMBjuGE7HvPlGlzgBbjbQZuBHCWkg0cx5M
T8uoVjC+khxTL8baryn8IcBR6/LHEhq9qWKH20AfG1dEW0WLcdzLhvDWDbpQVvZIffo0BxbRvy1d
tbR3SnDgW30nrJgp6r0Uw3BohmcAzKeeZoLiRtmNPtT4TpXdsHR5xaRAAKmCWX3ESIpXBrpQnMOw
ZP9Q4ffA/8rzhrpE4c2OF5XaUaWytu17JFCddoFwNRkYKVahalYMZuax6cPIbpuoL2679LD4V7TO
/u25dRstD4yyyWXMkaNLsJ/cfSR98W5s+ooSU6bgwCIlnCCZMpSkuARyE1r4+Lx9glSWHujPhv/r
/nnGYa7zbZXXMsEojE2rpDsqCXxr+BhaLzs1yVNo0aZuhLPDGaE4EIQiVWyA2G9F9hT3ySZ0TpTF
oHjbGOAyBYJofvf0d4Z988XhGGOgzpvvHL6iq5E2yG+BR9OekFbNFxVbydHVfGQCozpjY+QZUwxi
qFZN1K9o39GE5/Rd/wpJdcaNJEvaj2tSQlFUpPxrY0ORtwzGye70Tc1my4h9WKZpyc2jtV2OBLLD
mJBw2QnmusQ/jqDZqLnreDHwsd3adIcNoWw2wDwod7ZLFCJvqbXiPtmbn530mrw7zYE3RZjXucTj
m2bu62vh7SS+zTNVvkwY41Asx+fWmCEqrqYz/q48SO9/BO2EBSKEC//svdoMN6VKEmqp1q4VfV/8
oN+V1VDOjW4RljRwh5XQl1Ki9RzEBL0/LHQfmeF3UggXpw++kAkFJax/98KW+B0Mq/igD7Wn4WBU
qFu7G5vZ69FloqebHZ6toIW9dzJFa5xbwmGLJuE7MevcBvjYbJw0XhYXQPBpLjlBpSzPW8wS/Qsa
hvek1n0GhPKjQL2jHZyH63J2w++6vLcyeorPQcMr4nV6vhpClf4ugUTsj2YAZtk+PykSxE3c5/Zn
GXZh4p3qxcbuhBxJRnQPeNjFHs6IAeKmZiCuFIQu4cWhOWg9fwLYlFSPmuAkwMZabZo6DgkbDR+y
OyblMPr31Abt7AEMoU/M1q5LHnTmvoucV3U3Zo1TMVLsXO7YAub6yGdlbfV9BJeeSQm4oF5FFmAh
Qc14fmQHAhfXr/r8xL3QSCr9a1DhT5k4AuUQNUZogixzGcFDsJ80FNqEz/tOr3hBJRmvWw3mRySb
7quwcTDBdhVysHuF6LsrMFx4Sm3UwzEjnXw8jBRhPhMgZb1zbzTF3/NHR2QldwKu5vG3KE1OIsiz
IZ0anLjJ53D+YHd2dzXf74YrHTdNoCawIToPqv/4m1cqfw1LxJCDQLHsVNRUjh6zsDSC3CQgBupy
eVnsfb7TuxwlTqC3mLZeSHuYFqtQq4O7DZjk9NC7NN9FUvOprF/K0pAuv3PZ3o6MwGZz+Scy52sJ
lnPaAkVC+3cph0lq90+f7/yMEaaErxOoy13Atl/pObOS4yRq1p0HnVg7vSHmAICW8n2i6WI6t3VI
jQdvSTEVMxlzS+CUo+wUwe6o2A+KF2QOLR18EmrhDjXvE8ynh/MnzSbZdtqasVmMyq4PZ8112ob5
sO8flTvk66j4fNgjPnEKRGnW3+Y2/kbgAq5uk6XIYNt0YDwpBoLnF7hkwK3LHh/0dHhTsPP8Fkrt
GxioPzRGcWhrp+PlCwdnkl2rphRoUklLYi0JjOewNjw9yOaI7poFZqZPSD4lFa+EYLCz3AjOUJA5
x5yMIvreyfj6nbSJvrwjipuTe5ZPBxMQqafGiQDJvl26yzTgIN3iz0A/AlzJpszSV0ueLB7aHPZZ
s6BxgSiZyuGbe+rIdC2KP8WC3Q69mSQdiworbxtSlhHhiSB7OY0M1XrldQtULYwkr+OC75qAe2i9
TMyLSnglE9QHcgwsxmKa2j+AcwRAi0lk0wl/OWkPoCs2uTwOQa5RB3mtMMEXQgxg0QG1NvZtsGI7
eD1hgU0Nwf0Q6Vwe96i5KyIq/lVNw2rPfWt5zow2lPG3mpHYx70L+Wzx07DYXo0nk0eA5cYtkTZl
+bcP9XmMcImnjXouEbD/I1gH55gunp1xlLOLXx+fUldhbspCPyA6asa/5fn8XLLCJetb/cEY0oe/
PkgAVeVba1XHs6Pf02I2FG/ERWGmOnZ9BPeFmFPe1qGjSEujg7ukl5p3FyIPXGBkGWAQROVXCC6c
J0Qu6oWFnHVTxj/BedGuZ2yy1oWQRrYKOU+I/pefmgeDlLxbTmJ5Pz0tVvEfZdJKI3B0ZJIdreC/
pRPRxOkxrUVixHJZcojs0wNQIsHIv0Fazbie4kqVbuiYXQyIXQyT+EwIqtiuoFNd3TxqCzJDGqHy
0W0HVSjowU6XARvJQMzy1hXKQqQh6UjsV5emn1cvHs7KKFWDyhAXiyhyA5ykWrD2p3w7U7Hhg7cs
59y3Q5ZnagobgzZ18g2fixz0MKgjwN4vTi3D+/MqxBYWKgQ2VomOlKoQjQPSBrKpRSaH0opVsCmV
IndmHVENPlz2lqssCTfPNH1jtGrdCCGKXvsIOuzet4g8HeNhsBBXjTZV0m9k5mZKLKEmIK85EUUX
3Gl7KXa8/U51q81UrjC8MAJY7gQEZ2ymdUoz3ot1N2KCDd4dBuUO/5k1LRYeueUdEUoRnC3EAhpI
u6Gw7qntmmAZ20P8TIf/4EME6hHw/+tlDDFkbyqbBa7CTJ0WvlMR+xP7Dl2Nkeo8TIFPv5KM13uG
u8TcoJ9tF6sURUZYwKorjsrBKv/zWbObaDIZmIq6TSMtt0YzpO4kKwtmGXJeDASwfQtDKJNk55Du
B8VATopANOGT6MTtVThg9z4TvB7HQuoR6d3/S3JDrHhLKkVbI7vGDUyXzI6RDNaCYWV+9ZB9kFmY
5FyaXb6t/1S9VKNHpVY6sp5cMqq08cACMPd24TBUPvTJei9hc9pDA3eRyXa7jQcwDDjl4Gtg5cUF
tz/2oSGE/cx8p7WWDXM78pEAQnNdUmudBPXCw3eji73T18GKuYIoE7XPx4Qfjax29CTULP17VSTa
o70RtXUTzCaBzZ4Unp8wuzBVL0pvD7YWfSo8CesXwyMClziMN0el6EkI+tmbVZQ0qJcFu4NTi6mi
rYaIfOsrzsokY4rXOPceHButnvhg16zH+b+TCSuIJ6to3mA+ieamTFNC+y8bUJrnB4HSPqukVNAD
rA5sq3qcPQStH5m0B4gtuICZ91OcX+y2PGymvg45bdjzS+Fu2BMYje5JX8O1aA2HMr4q8cfGiRen
Yq5zPRgTXx6ej5XSMu5G3KC70/ZYgTGEeCodEL41EniKhvn6lbjjs7r64dFfk55f8sFCAw6RLzaR
tyoFGM3jyjCCEesXdGJKyp19It9jGnEjXXMKEDCVMQEoXKSIMrJqqP5uJsO7gjAfZ8RqQBqmG0uC
LZ58M5hGzGv6/4GFixVcImHHesedDuWLlN10ZU1x0L3dkOiAAN/2Qj2fEb1Tq88lRt5t6pVqbOIF
dWQCsMBbrtlkXX2r9b5yzhc26HKzit1/YqUI7ckySocUPSKrUeGM4rKlsxqvbNn143QiXwdH06sm
KeCqdusgQtSYitdRrpPY/qXUWEyEUxozp6dJmZlJBN5zlp2tKTg62N+7QM4oiK3MDDXqzh7ohVP9
wigRP4C9flJFJg6E1ZP4SXxZdYXDw9gb/frNAlvvCzE9CmMNHzPkKkMXoGG1uv6ZC3R+bB28oHUQ
Z1B/4GxopezFxkSjA1QqRNFhjGfEexXDda4fYKKKN+qYNEFvanBAPnS8z1O2lsnkQ1H4SeS9JDkq
LXwo0fJLIhXAgIPzfdFvRtERHX9DAkp1YnJjA+xqeCLlnhrM5H5M8tXMWlQiWnpXCaHK+RFnQU7L
9q6lPAm9+PcjfeCPvpCsjm4GfnHP7mh++AkI1r1ShWJO9svkFqsx5WKhRJhK7fk+HvesVlylCCDk
Qze18TT6g/uz1tfGOmbFtdr7P3iAscv6m5ieKFF+kvnjTcjGspvtJRHV5ZUj/HQsE2SKfFV5c2C/
C6WiqGcYLDh8vklIXRrcuwSxlOZo09Us2SrtdtUvwRRNLKYFIRO9KVtOSz5Q0xErTj+uPGS3Wn/Q
SCZIybU6sEKtZhNz0eTqWznVuragijCq11v9w9MECjVXBf1weKXhMeJqBnO1m1iTKxDAPEM5UJTe
4+fHa6Ukh2o2furobXK/lleTtq9ToTSJv5yu31/NQK2T2XulCC8wSgTgFrvcweTlIzruFfJnYjHU
LXoUTbr0J7g015Bp0K3N9uWYcue7vY0gd9oMNkDE26ZXa/XQuY7BK0SrbO2Kx3vSG48ZmJGfdYH1
fD5IQnEK9A1XY0E8PLyFF0wzpF9h1piE/nMLzcrNMIdbxr80YPJA7tJfSDJhin/MBghhmDrdX01d
sttGOathqYcIop4qE4B1Qpm+RFjGv4fhl9o/a+bSOHoUxjHnsix2QRW/HW3Nt4b6roVnzC6sjqbY
GteSAb9NVGAevjUu5lFbCrZtgrCd2zSLNf4PNGnSRo68IOa0a72ed3p+ZwaXdrhQO3fGvH3LjqDs
fFbf4lQuij8qZhtXNDWGauobKvkU8s5/ZfWhQOSvu7VWJvLHelcPALjmWi1UTXRtUe/LQNpbrfn8
r3omznBTjlHyrOijErBPFiNaxZvRRvF+14tjA2ZwqlID6l7q8sZ9CF3Er8zXw86sNCSQP38fiE/t
i/pUmDZmSeYWk2NFiRg7TOUw6JyV2SnBGGJWwOzEG3/Wn1P14lidnC2xLTDLBJkl2QcSAiUvBtSP
lwN6PybUCrzJiFzYT4LMl3ogvTCCmpzJcIgyx8yZr91nvSuYD4B010kOvxL3w/0o95M5GFQXLPfD
5mgCJPOkWQqLwurAOQ6AEfe36wSyhQo8Bwjp3LlFxK54T8JIe/plUDACOknQMHoEj2dgzRvELjWC
kYbSaU4UEW97QID+4xYb5etDcZkNVyUXUwiY6G+GBzKMCeKFalbM4MdOw2K8s6LEO+odfhYvuu8I
8K3EUpAqeoEfVs1xtumeeHIkBCKywce1OXfrwMwKqMUdHUbuGIz2NA+w2FzCsPJLpMiA0DBoYGJw
r5DH8f3YIlQte5tHDfxOcVvnda7Dq62D8Z3kBOo2flFn7zYfXuTGe0R+uOIQuugkMX3ekqsM7gAJ
ggA2YCqrJl58ly8ohV2xisXM7kHtspRoJkA++gv21M9zTViiMIq4CFVSCDqb0KJAF+0Mp7VwBOJH
c+eJ3dxQN/hjd6XKoquCaSgT9H5Ob79C4OyGhvtcy6Gkd6zsiHZLOHsJSiWed535J0/I/5id+YdJ
qGhm6EKEZc641qGYLkDZvy4DkW7tP9NwfBK+uB0xMjs2EUq21DNINYyGNUVtNqzTTLXs1mhkEON9
9IALznmO3q/0nF4HXy9LBQlPS05c4oTBAFxUZ/eadSfhkHBHAlXgcYSHIlWEkZFTvTpJja+pRGdv
yVYjZCM39XMWJ29IYfknNiyQ7wBm9vs1yhMXl9Z44HqbDt/lYdTZNzSXthLPk61/uGfiIh40XJpC
pFrlEoz1nre8OgxY3Awhkqn0ZdMPrY8VG+LXEWNxV0f1Ee/IjHuJpxel0OUnvfdOplLdUlmodc8d
GchiTI9Qrp4pxs7f+JpxEZQPRjDVT9WasilIEcdsh8MdCvS61trvPKUcdKI8/dGiCMzQ+HGDuWxu
aGfBfBPZJV+CjHtXtf6pkTuTWcndVHYqdmFBVw/rmMgZzGgi++oAI2bNidv/n4Rh7zPWaXwCosh0
Vthw8fvC9wqHwfOtVseO6D8y9Kdu1wTgZl7K7eVOFeOHIk4ba1yuIqoRYA1JDwViNvwCu2G/Asbo
HiwaxGHC/dgDf/grkF9rzt7zA9+RZATg2fAmqmkPz8qjrf3GTUgYoeJkVI24ZEza5L+7mgPzsRPH
Dm6OPTFRVBjRBZFOKa9z0Xdk2FmFsYidOWTYQ4uFOMXu0oFbLHleR4EYutodERAvOGOptpYj+SH0
vpQWUvvkVqTmDhmlUR0NIppD07XUlvRfhkseb3wEatHX1bGHahUxvrAUtR0BnrrR6dNEYJD98cUO
o6dPY8OD5ewV/XlfAOjqoicJp2bIJtTWkroC0k06zI7BVx25lbNLf02yhOP7ZHTdKJ8p3MrNkOxk
O8ysGQbRo0xmJ4hDiJ28CM2Etsints9hCOA1RBzdrBy7ItjRKCmGKoTfvo/1Zb+GG1XxRtNT1iOB
ICNL/qfLZ9uPRtj66OWfPx76pEQgdiAfFgwNKDpPK8V6t9pSvglVMpJDWSrOBOxa4wXDrcOkMXmB
5AK0t2ZqhxWt/fA/XgJJKgsiqMk6CFi+oEawlNKEnpDHq0gX+MltFC/zwTcHmiSa2wVww+V9Jw7V
i0CCny74Yu3cVyVLxeYy+W1Isy/xp0G2HwPE/gG+XJwKVV8u97LsDf+NKwpX1J92h3dGCEVLO/yf
KQ2v6zrAlYz4Sq+or2Sb/Ty3Xwey7E+86WOBdlE0slZv2DRFyYMn/R8OnrPEe665cq9HhMyD02gZ
Vg1hAaxcrkp9OiQtrBulCoJ+AGZ5fal3edQ45jnZJl6hjeEQf8Q/WvyHwjnsT9F8w65oCTvqzNJD
K5bZ5XPmGMrItxqzwnTdLK22sfwVnC6g3LhBbUkmZSAJvl4YXiwAP1GXeFZSQwaeyHvNNOziw/qM
j/jx7ANFE0vy1HwmucFA7bUnWCj8mlgvPIjq7/jng3AOT78diad0fZe9DQE9LMiYA4UX6/4nUgpX
bLjhSedD7VZEGrs2uzq8nUyWSL1tGhpivST3GyHfYN49LjikOAb/Ddhzw3/1W66lGduh7IAN/1qm
2jjw/1hoYxzL0AB/xYPqoiU7OgeVECGnUMLmGuz8qwFKKn/q+po0V8flDaZcA/l3jva833EjpBw/
GpMUh/T6loqWF9B0s3mjDmnPvf1j70Ss5vSN7xwRisDhaL5IELyu0lVfO8QAMlJ+nXsPotiBP3x4
YphPkaeD1oOowl1pLHQyWRd0tTtUPwpftcy0+INUYNsKdGfc41HAEYfRZ97TFa8ydeRcO2m3xHJf
viGUTIBsorHOKZCS2CUKWqFtALv1o/ourxHTnrxo704KAhuvv6jSX0edLbHy7O1/554ulbbnn2H9
aWTGMEffxcTsJVip0dH70OagtR0LAtYET8OW25pQ99x4+4GgpMWgihyAxaKQf7Ggu7JTBfRPxgqH
ZBNz0nnxAkIJlEvdyzFSNQEwhu19mszaX6RJ/W4tEJrTLfGcKztDQXd6jdA3w2bku5+4Fahe8uhd
17J5NP8NxeAMlWJ36NbFg0oqU2UjwzXitIUWAeHvS2c6Ga5dhPGHF/2OkEPIWDMu3/wqRgni256t
XrJTfob3VwBUsHJ8Civ9g2l7sC39JEcrV81LfsQWbYOtflQUMieQWLPEDa3pG09kjdUdC9o1+J3l
4CVi/44CPd15xAUcaxuHfcIjwM8lJk/0OFQ3dmZTMZKm7ezfBZTugGkxIhWPquhDq+sxo8fHla1s
S+WlbMvpYYwbUS/o2InAWVbs26GwVpdvQ6Q1kBVNzcJDVIwKZzfCHopMX8BzdVAA2uIOgfvYWCNj
Mqfn6j6AV01Yc5gOX0QlOCsxJfZG0KNqPoV3j30wWE0bf9/sg/uIQg112iAdpofp1+DKPekYEHCp
MjGhP4i81rlE6xtELtYTDnszqtUofP9zCRA7JRoZnUykWokmscC6jlqoXgdsZ9UCBa+J5MZlzxSB
XARjOWoEUDoN6oVcwSMrTHwP3doUB54rFcj0qKVDWDu/fmUCVjZhWz8S3bBKCEyfKLyfLs9kpGQ/
2m45ok7P9ndH/xu77CUiRzhk53+Zq2W7e+VB6Ecmw8H6N6IRLBXO9HNbwPBBvLl5Vbp0OgXokBiG
5Z7PuBjs+2b8E2kEfQ3XGtc+UbsBx003aXZYYDKpSHiAHGkFC8ZX2iK58W8IOAxjP/FoWq//VpRH
gcxbMOjPYhJC2BDHVS+fUpLfcTJ2JedN+b/n3vrALVEGxRPJi3x5+jqVfm7WydwmePJtLmHbTwzb
ZVUL9paoP+Q8qxozcax4ANwjy+Ybs8ij+M1XghOKQtjY+CstMAl/QsM3oluCFVc940bxYSd+nlmG
mE7cwn5o6lDaffcSitZud5D72CWp7l0Za2TkUyRZv+92D5NtXsfW/HANVcyEPAm6zWJiiXYcR6ln
Pygry553Ld8BT1kLNVTn6UfO2Sxh11qyF8pm8qitkdeqjyZJgF2JcwyopW6pnV+uj+y6cpePPTfR
3j25VB2fNSZkCtNEIVkZZ9pw+5IsgSua/Qxtlhy5ICBY6G4UjY7vj310canMpciwC0pj4U5LEl4X
6fyscsxIZXoAdmGVqkGGc4WOfRpDa2MIPvSunECPk6kDAp1tPi9L2CZYoNpBDhuJwyUnvBcHELzd
fqBGJmxA6Yvezh5j2roM4nIxbiitxmnJxaRxgutdy2srfx+0fqn0Ls+2MQtKH3rN+piATCOREg0Z
2ZwvhYhy9lC6MKKAfXjdoWcS8E+KBbb3Z39KBeenTqKiL1E6rryj60XsCNjT4iEX96D90yPiYvLG
y+v35WXNNMHr8Nth4N+3v8KpCWegivuYgwO68CjO4YBuDBXfprHQe7WmufITTkrgfbhVBUD1iipJ
wCbc48i6Mfo6PUPVI20Dn0HGqipHKfzH3htXryxgGW1m6GcOcEjhRjSZ2CPKfPJTE9FqqDfmvf91
OTI1msnnJAU4G5doGrVPz/8tbvRShxsbr/3TirrzzGklx4J82K8lvP7LgdPuSStujNjqRUl67qUP
ZC+A1mrZRKvFRy7b/Ce1ZPPvXCrA8+Jq6K3bV20SOe8eaMGQHHSYfda5b9TVTtIlqO0+z87oF+4G
Pe1BlOUgaRvsa/9sHuNRgvvjc4cNFnEyxEoyWkvkVigMeL8K0wwopX0QLOrrBFuCYbCcGJ4mECJv
1EX8Ea6h5KPgF4Qa2BAne5iDq9YjdGKMo7KfmXPlIP1y0daXq1PDh2JfMOWyYHZN+p6bLUcE5Yab
KTnmx6hSMbZ1aNrBhZzDYCtS5Sa5JN2Da02aQ6TwKAANrpvTLhEvtQceNEIHXygoHq5hd9aSbU5j
ZZwZi6BHBmUJ1ifoOjZXwtlY4UiP1x4pN6tdj941tDcqKoQMcXD64F5L4GgR1yezGDOfhdu/aWOy
6H0RFqibwonTFwLjaAKnjqhmSQ9bHMm0rLItmqZa4wFuXVCcZGBUf79caVoIKs1aNEy+SCYm82RF
XNPrk9rPaflJcfeb4VdjcRTxUe7v9MW3NhpIv557ZBj9rRWF5SLN16XFdlzR/79Bk7t2XFf9uvjo
E2IgIIw83zDVOOB8OHt4PJu3YRXfgCrXcwQwKxexkESWr1gWTjCz/mvpCdNY882CPG9Ji/J+ifor
cxDRue2lv9QvWf2EeTG+5D57llm1+Jvn7JvnuQko3Kk9s4fsUcnX/wMK5NxqdUPuoJC0YBOPXRUY
fherbNAVkfi8GeWzCElrw30F4M26b26qbm5orlrcpFNS4M1UC0JEviAAB/UDODrjFxS2s8+ft2/7
xN85LspY8NNAHllzjsVqXBLRBGECzNAwzK5xyxSp8269HOpEqoxVagdV0Xygogw4o805zM4VSpT8
q5skjKLwd/Nh4uPIk2W8cfg79PTa3zU46NOe6/k78pYfSgmAJXvuJidES7s9Ot9SZZAeHNku5Q6J
9HoT1BeXaRHe+Aiy+TQuNZkFM0RVpwalAZVJRIG1xRwHUwUKjzn3//Su4EfBwE0o05M0vIdhAHl3
k3QjiHMeCG/wN+cqTJBlGB9W63KPMOqBETc8AE9/sR8ZT225nwssjqQGDFr4Z1ULXlRLqDM3usOj
DWs0K7wIh0vR9YvSG88zL5GhI5GeaN9UKgbJCNQW62/3m0+96jcN2mYobOvWfnbQgggkuXM6RKyW
TIFlM34dW29UJlOfKkBuUvzWBGFBtoQBByowmB4S+vARPMje9Qj86nGaqGtk/ySrmEg+O2NmPW7q
9Eb1EixQzgEYXb/8q79/yyTGuHpLgcE8FFCzL0Q+H54jo9HI9lzaU5RTd53IHDZv+VseWRzBBh+v
h8xIlMBXgnT04hzov+c8ouxMC2AiyL0nXmzPot5AAeeuBZSVo0knSYhvmHU56POkSqxnmUmhlPd8
O0Ok8wmmX8lCoIFuhK41X2iFIX1FhST4k6tEXwMysEp1LH1WIPeh++CUyUGUKiRXMTlarh/Btkw8
4DzR/HZqi0+ttk95yOObjiYHckf1MWNcK3M8FbipAiuoBr5AGIn9d9XW2TYRq9U8gO9NtYf9CzM/
h6hq6qoQIisQ9ZbHpwgoI2l4c0TIpSM2dIhAOQil+ohXffreun4RIPfNzAMAYj23pzLAgHecfIAA
RIMOaXgE5/uorF6uSELyyLqjkAP72/BScPFwcl4+oOTWp0ADZeOWNO2aka/tlWJNFVQwb0YUhxR5
53LygqG3zaibiCaM3oRw3cpCPyooqLI+PfS9r1hVHqRYtwqPuesRcGUa7A6rxpWx8BmT04x6vs/c
dmngJiL3ReKGDb+PAjVCbKi/5J00GPRLzaE9vR1rd88/yEPyXBIXukrXd/AvR7QP9pgfKK2kG7Ok
UARi/p7CksP98qOR9mmQRByri+lnI5nPEzOnD6PpOqLShi/x8hr/mf3enZIzNsDQ7gu49hZ+unei
MfGS/eFdDeYHVzfwUv8wFL64VYddsBqy/NGmeiXw9aRq/ChMNWJlWebjUGIWizl17gQ1jWEc5+HU
BsmNsMYSuIe4cbuBDjkgOD0kFjVUwkbtIMSkK/7pCpP4qWJ5TxfsZi36AXs8178rexNkJIOHbfoQ
b5poWOXYxcB22ZT1PdTwIMfv6VJwLZz3J1PvwtEwvst5szedSxF757pVq94LYBBrcvA3fVABkAcS
yMTyLwYvMf9o1GMFxLPNioqjttO0JRABr8LnRzrvoxEbE3ZraZs3wm/hlJ0E4CrglVNiMIRSpxEM
B9XBGXxO2+6yHqzPMnoeudsvy7/FJyYNggfQlHjaGVcztIZynn69q1j/Cp7okJjQji+gnGu+eatv
zmp/kLJBo+aJAcEhvv+ImY6kU6EHdVZikDMalPmTHFEcqjfXWqHFIC9lp1jZ46Jg/RMZNkvLKnwH
qt+B4WqkxYx8faxJCqvLzMh2sMyU5zW4rYWw+KBJ1qnJM/uBW6Uk8Ilh+1PMa8dkDvnr7YXzHAh+
ydfAHCVvoDPbKLM94IIB6zdOFvyPg51jtW6gL7AL85MjHe6Mx2vN8TlqqSFNzOz/4ytzzKtshICg
feFalPB33hwUvE1iuF1VWFDwomwvDa4mc8OZ2lDYkF9cQgmgtL7BXQfmwOtCRI9CTqJNCXdfsPPp
Qn9gzk+QR3LFsEuiLno+gCb6aDfxIYcKsjycVm+8DZCo0n7WhtFdIMDb3ARZODmXGoJ9GmpakEM/
VXqKXx5q8hdLLvV127ErepGMR65Ltdqvoc2C6jCbWx9lJh/9za5duv7+rnaY6EPvtf3Zi8xTn7jc
389px8pbXyDWx/OICjeqL8TFRwsCeoreMvgm2M7tyacUu91YkAdJrn1CLIudKmuCQtNYEQyM0NMh
0Ui99RzISdDxAdPK46k/VtWVyqeaXO8z4c3wMHySAUc6Nluxi1/hS6L8p+74Bk7Mj3BRVkEQw3nQ
NTCW6HxJZoR4KdzPU+DNCc8mlPjEww4ZvVRTkQdIwfsPx6ZIrgjQl52hU050z4wSBv+pkYN86LDw
EoV1HHD0WggCaUZDMl0GNTuamCVaMyBUdBYOxX+FlEasOm+57E3HreWrOC5gPYo1aFKI2Qeu4QDP
NVNruuVpNhhGOD/D9ap9cXAQd6gENfv1nBJie0IICfV+6rdDTSK8XWjLnEsSSmG1rxGOsXBVMgVb
Ow5pqunwAH4Fzb6cyYMQVB4jThCuFsluEQZSnbIHGryae63qLsLJiu1WwWLnnW355PZp+aJ1Dfb+
JszqnsI+PmmyAabqCETMTodQFs73aBb0KQwBLTI5M7sbngAa+wtwSkey3rcmlzLoEWb0iiMYEHd/
KwBRD57H2sDE0m6IUxlSJAwwkVu/BIjUxVN4guUf7zJzkU2zoCWfRFPkPtz1OgKoW6PEMTWglukt
xMc3hraVE80reDCWDkiDrcaE6hlX5EPAX7jzZXUK75lq0wTPNsVAc6V6+n79Jgk6eAq8F7Zb74dZ
3Xgw8Fov9DxpaSOKdkO+fI2S3r8BUGnD4g8rvg2UyLIVna2QRx0zzoKa9xaRLtNdwnw5ObYlQNRj
I1oZz4bxnMq+4Y4VgWeNi04Gi9AIG2KQlmk16qmqywpMp4yT0k+9CaLBuMQYdkSJEhZs1mRJ/6B4
yMSVE+wqH5Pg1fCdOkB39xFflbiqF961EY3o0TYDjSLdkPPU5szAz5r0nuP84qtLpNzKzjzmnB2m
hX6afnuMcw5jHrzUK9la37AChdljlQcg+yOWSCK0RR4d4UJs0v0JwWSlBdd8A1YZxyFeJrmI+0Ex
7LfxIK2tpJ82w9L5cZFZ0KLOq/XKnEoR6SFF/tNBc2GtPSSG5cRNN6l5ALX+NeIFCzHwP6q8BFp1
kRUC3RKrLNszRzbLGXXDV+bgunMjJIKYkJ54UHMIUFiEdKxw9WWR8eeFgBLmOoiOI99wIba42TGa
BdFLs1iaHIOWUCH0q1c62/S0ER32zaJedEDlknc8hX7LOTdTQs+vCWzONEheD9p4jWhWkMaweZAW
Mb40ajtITZjtqkTiyJLK1hDIDdULVtRk/S70omfphRQHuMHMEl+GVYK0EClHkhKJgrb0wAMzlH5o
6358Ji+gCKHnwu2xjJ1qoQnw14eu2dahjxoMKBcPxkUqb6e6EHAtjJhJwnY2fQNzFIwDKdyYji1+
z3LxVI80MlYscTz1bLKn/sRYX2bHG23P+7skgp2ez5tSUWRTt3cPwWnvqYI6VNnxov+KVNr62Fc0
nmoT+S1HPBOIu1SLJiiS3FxZRJqRBNEN3sMkev3z5eX1M6cfTEdvSjZIXzvy+l6bYikSZ/TIhztM
EMnNDGGQppH12ZyjT8IdwKOnx3oQ0gQgLgO0jz7gXdSraZbT7y9pWME3bRK3NHXKsL7FZ2R0b+OE
ed8qPmZEqCM5+h1cHtwdU7AVkxutAEjl+gRmezZ1EI3L9CQzxppOphPMOIPvh7Pg2BW8lAqtL2vT
lvg7mj/SI0i+voxzGlKDiogpAqzrTmsW7vR1NarHWWkD+nYLhpT4tY+qoogLkLmw49FYfzycGNnG
XsjzES/7hT4zbmj1aGg2H4G2ZSaTXHz3Nozc0+qEZ9KDufWhg2Es40U0/AJFmHJEZYCCHuyqZUGA
309u62k5G/fRQv5DXNyx8db8YrsSpB6YfwLGMr//uymXgsNjHSpJ/CKNiMOwn4FFTOMwSGlXX9x9
QENgIwECwZYV+5IMMMXvkSlqk/W+SyapM1CfxSIQohXTuuNyjphOC+GJqX3jGyODXcLvBq/3zpBe
3d8RVnzIjioiynQzbF4P20MqV7rMEPfyEMPuDQae6hK81+Qf6aPz75jnU0hof8iHgPjz+9FjmUGI
ks6Xgabx+MS6MZuI0/5gkLHDU8pV5a3vzbk2nPyXHC2mV2PDbE6P7M1qk0kio+FYTOUaMufbTxxw
g0wV/r94kn+7cfH8pg3sGvY+ACUiyM+9SnaGnnsQONYWMdsR5vt2U7weaIffOO6hbZFNhJHyv8kM
jvBmw5kbZJ0R/hkBNhXIAPuvp0GmbXejlXBGZRS8BZOxXFjvjcKS/1Mf/LiXttTeIyjpMn1OYK8j
iwrIfpNAoOHmb0Z9JxaeXUZdehBRmu0rchhkVQlS8HwIqBe4TK9GrQwKVoe4I2AE3+kONPGJoZQG
bAa5VcmLHqHjYmxfAGSMWWMlBqKi0p6Lkyk4J656MHl7yiH/ga+RdJbUlYtvZ4hTo2GXvfxOou6E
HIrfv9CBOTXuKxe4diCXgmhrmhrgpT8dxM9RrDM5QVlLiW4dxxV2s4ZrGP27T9gjCWPWJvkTvYFm
VLsQm1I4O2OFIq0yXR5ZspypPic1VJZlfcR0YsWgqOrw7kXiO02AAsxofUEsvzGdqqXZm8Iglkz9
s7YwQfpO+cJKxqo4kd3BInxgi0G/QHRw6TIMJaVfw9IAGeNk2HnnlyhjK3PVANWYHqQa4R1eaxFE
hcu3EiiNOCsqXW/72m8WyTAUfuLIO4BHjA/OLcuyKQo0UKaul6WoJCjhVNp/Ga/2Q13JmyWcvGnA
+ycbBodp3HxV3OhV7A6ku4GoIsuGMe201XEywyBxPZRK6dWSsTz0l73gwnLa4dToHcZwuCzlmVTc
S7CKEOJtTZ/TTFIeeeuzoyMAHjPsSG0e6+eIl7yrBdebG5gsp+rKXF7a2f8MPmG0JaqyCZC28kt6
B+8+9MIQotbdnxhDHymY5DVSfBhfbiBNWJrsipJI8SD5jV0Qavd3nGkW7UiOxssB5suiiQ4fyR0e
I03vzLTBFeU3BqykFhFOf3HdBKBf2HYBwB+qQwI7VacI/v7srM2bxRx18gD2Z3Bjv9b/ilRUke2T
zOZAdFRPTa2NpuoShvP7rAdTw6EiHRDPqmRqB+TKOy6553C6fRNV/kPKEcNz6O/iTPAF6I6+KCHu
62CR/W96hpcW9Qb1dCKe/Tcrt8JyuQP097nX2OUzHVXhwwyi8suhR1DX4atPwDyGkZ5IydnFCkHX
NPPjb0rQVgGE6EIhZFlvoq8LC7z3BdAcHghOAuXlgKDg/eD/1DJl9BlSdiwni++gsQr3f9Jwxy3A
Xl6rCpcMSnDxhBBUONf1Iv5YSLpTaOjcb/mx4kfOKp4OK9Reps3DwcNELoQskZ8+N+ejE9PC8e6c
PIFH8gIM4PPPei9dz1nrt+obleyeRigFyIb8r/VOlppNSYMY9aUj2FEguMa2B27QGQxIoB9X19DA
3imqtUEZeJcEl52AhnLD3zv5S6ywDg+DyyWtjLZsAqitBMY2LR04tkpzKWYnHEJ6d+4FdslfV47e
fiOL9A7ij+82HpY+8Q3cY98Xt7ART0DdD8hzerHcWs+goPg8iR7uKhf2q1WSNmPdRNPHTeBRBjUu
sreEhKGs5qOVzUnisuQEFdRFPAh5AAK0zi2hnriWD8evqicU25o2eDOmZyW6TYoA9eoIp49uHSa7
zKxkAblfjxMDYzRAQIafi3C6OcL0nP07uQd6GYbwjZbzMuwRXNMb3D2K/eTQomBi6bcyGU2BTYOj
8iGDBv/bOO7atd1Q5lx4TdhYXtw6mQXtcQjgBcQtxjdySWqHHPKkX0bYuA1obaJCY/KrC6RPj3OL
IAQBS1HvBD9SmpKs6SSJOXkhklWY5JK+sLRk4qDDRiqpjNcY/g/OhS2us6na2COi8TdLxLZ9tziH
nUYrruSHo05wIIGAaeVJzPkrfoW3POla3nD+jtrPAkIQX36I5PNjn4LXmMRIs7DYgK5OPagIK8eN
UKltOnfnwm/Dk8GPDSlyYZMsSo/jLYWsCLFpLRfBGNxibHvBSPjOyTZGW8Yy6fHmncsAn316yyRb
Gf+17EzTBWGb1NG1ut/12ENCf4x+wPf1cUrQlpKIL2kWRM8kYDG+kpU6kAxROb1i8/rU/UFt6HeW
Sj1cQBUy4twRgXtNv1DlUcz6CldNHJpTifVWVJml1agNltNEDRnLYB4kK3MI+Meo27CcmnO9Z7xr
E1lPt+CJ1/QnHRrEz8xb7h5S1++UB6uMvBSlOxZ4pSwLf4UMdA/cg1AGJupn66+FuZnkwDZz8RyD
s6qoN5ZoitCyEjJ/Hxui4ukNqqiEZHkqgniIqm9wjZfkZbSx1OTakeACMZkuqJqWAQ4offfb2Ejt
ev7yih5yRpAes3FVNm49byKvTUe2qFT/T4qn656VH1Jm/pM+4nAB2H6uBVnPX+2mjh/PeMioGpkm
3ZAU/xRFxKGqllUVvV+bMvhsrOOZapS5iTv3s58VreQthKBmQW8An11wcz/OtaoJ/5iuDY9LTjdd
CSJG4dSUOZ2nEZGX5kFESzr8tHNOXkQPmqX5RnYSpaWbFL//eU+CKsL8xS3ZzYK3wfRPWK/iKaVb
c0tq4hGCXd8FVJyZDlIqjliw2ul6owaFPAfmm7vLU4HgqTY1I7LAlkWJ1ahzZnmXa6KqKVS4wbwt
E2J0MxgCBYEwMFncLL816zTmhGaOuiNSuA1FQIeSMvIvQR+SmIGOqk/HMIjK2cCCvbwgherg886t
V/fJbL6gpAVsJRftzW4VpTYQKdiaPudUq4iZRWeJRGCg8LTY9aL7pm8QKluQTfBINotMqqtkZDr6
INYFdMOo97xw2D4i6Ur6dMya53I9boAQgOBO1I6HeW7LENQloPerKJ5wvxZPNzMXO9tPmC5L1U+n
RS8vWRO7TYdi9HNF03+NTZWG1n4Y/whAroABTmLBBk6FwUHs2rXB4SRfWwvxPo9JBy98LjPGi9sz
ZxylNrWPPiuLJCMF2d0j2ZNh7S295+uXG+KFRaYJ3NT/HjZv4fbl3iYBEwzUGK1Vb9u3v5xwhPEY
l4+7PfkHupZTUBN1ecj2P2czI57C62N+OF2aPTDSP6FANhCuSnhecN+6zBJ7OF30bJSZE+w516yR
CBlm1M3d+rHplBRvkDIJgWdcuBqvsVTNrQhHi3t6zhXFZ9xoToumAqWK9WDFdRkgtUVlN3Q7hvhR
zxN3Hw69qjn3q0Y6Qa3SWI/yUal2JebdktJkh1kjSuXPMonvFHG69d6NaPic2DIAHd0FYQn/BfDT
Bs9UyA7YJjDlHrWuMdyeo+YgKdCq8Z/DRcltqg0q81+0NSNxxRPSdYsU9Wys2jD0wLoO/FAqaBcP
ZiYtDBGDHoMv4Rf4drS8U9dtqiDbGwOHKy4G4ecHEexJZ6rrN2/gZYhGwquGLhz+LYnPbWbjjEhc
jDqHxlmbp5Tp5Mn+2hbL7T9GkVPFscBKiSYhYKLeGugoglo3I5IkusesumiexL/z2JwOif4w/ri4
VpM3qBv3waYuU/WgtVdwMqNAwSUUlXroFyPP8CULsuPN3mx8XsLOcC3GlwPJ1JkzQN3c3l5aJA8I
fvfxmJ94uETfze6Hh6su41SQqMdwKqvB7HoSuMh6SVQlx1Eq+ga0Vir4AjMc2dh01WiLDASmI8hb
j7RnirDkYyLfc4HyXU7CaPUGJTLk48lIweY7/GWR45mQIPLgv8IddfqYULEZOzdMDTfM6wafE0RI
4OSYl/ncfPRlfde146pB/y81vmYUgGFHP44MtJOHox5hXgIK9rekuMZFeVW0w68tPGF4TzTRPb3Z
1mnXTWUz8ukSXJbS/YroDWByae4eNoFoqrJdJjJkhCRwokE7uCN6xMgj92vxvbobLZiHhImcDmYr
lvXYHVBLG1/adX1zM+E0hfULnI/WhBPUT228LvffbWG0rxFigbZMwPeP6SlQKNp4PXPz1y4mRv18
8PYBoUD3U9G1K+hX1YlcDH6payafaAxo7WZpWhNwmXDleCvD6Ip2TzH2zkz+xSMeHJfFTpcxMdPD
AnqzCbuqx58Cm2YUbLCTNa+kSIFjpOOSu6k7bQvjfOGlh/+dWqAwhnIRmNRISld1Po0EItP8ECk3
NBQ6W1J6UBaiIqCIrR8F0wAbsA1aYKaL50GTt2ejGu4WwkXgbS0eP0lgzJGTvUTtEmgdRFF+w+GH
kGx5EwvrjJstBMS2EktArj5PQotaVHH1KIi4kAHrQrs5u808prLXlQFQd0bvAdkLYJgh53QilPaM
Q9sQeFGpj6OKGsAN/JyXAsDB6IoXiPv5CiwT5yhlfhBMEmdpgpDvLcHcQYczSLNiTCXJCdFZEROC
8mMmPgWjBjp03XPQpkGhBElETwaa5AJd0ZRCj8a3JjWCY2WXo9uNo89qLpgiGLALL/x7HdFcm28h
npO2veRa8rQhaP9Qq85dxQyyHCRnWHGXKvIfm4C63usme8YhlXjuAd9gwprXSodVGDxa0zd9Uw3f
KhzhwpWszc6IfPFagsEpJlCoWJxanTSy+bKJmGYIIf8nMmaqoO4iYx4J+lLiWFL8AiNOYoDX45WW
4LKAjrYwgWF5XXkURDn9gMAzPpahtNPSCe9fLvbdagK8g9Xy7n/qgWyoi6hVPOqnfnlVFoehGAoO
Z5RYZA/cio/i6F3niaP/Ysc4GgMVXnK3fBacmJOvJxSZVoV4ASJtPL5m/foji5b3zxEGAVOJXTG6
pyt7zfK2JQ5fpOaridBi1PjjFFjKldckHkxcipBCKaNXmcH/KH6bsqTZEt06RFLKUzWihZpsXS9j
PvTajcuBEQUIx+XW1D729x8XhM4YEaLdu22ubHD3NUUyNLCLd7veD25PZGx7QdlGUkrazQdfXZ7J
+SZbHUmr5xgfzPNtntfmaQQzLMz5ElmP+znVK13/4KwCD04jnU6Edxfd8BGRcdJWDo2FXaUkUtfi
5IwH07EhM9WibVJ2zPALTV2lHx3Wmob9KhT9IACfxmF2x/sitB3dTu+tVVRRkf4aIf5SNiEQ+sIq
NxQCs0+0HO1/MOi9Onp2BG5ugEplSyDzIDtClhA8XHqp3QA4bT2lkj9SOMA6rI84J4Ehqwok28/C
FciHS9o6v+3ZKFz6RLKBy6gIBQu/SiojHGGmt3LTWt11Q44XxCJodLegsJX7FIC7vlet7FtoGXL8
gIopHhwazA5VQ7xESlIFaeNvUqNcXAaAxKbtdE5XwWYNkr/JC2Iz+7a69C76+75oleRYSvf2KZSp
eS/bNt+Gc9jmhUjO4vNabhWxHbF4k/q23YTAXIXV0Hj2tmGgXqdI1u11bIPZQl+YxmFRsrlvlNxm
LTOzyF4ad4cxbvmGa6sxP5B00EgUz7LQO4LJ15wSoGylYsQXcmGHyb1Y7VLnkGMd36fhzp6j4IR1
YtavAkcDLBAUyOVwMOmm1Nd897bwO2sJypfsmRlyIXgVYKrjC8AcBHzXqN5+rORQ3W+ScuyrQlRo
RJSgx93fzzkXxWQpiZRW/eBgeNJSYgyghBV5H0A+N05lNPhSg4AKZkPSDY3iSUnCmWKdITOIgnfU
O35O1WaqPDHHAIyO7FQG9MYUT90jBJ3TvO60ns7CrSMwLyco3Mpals4EK3UIaN+fLW4TwCtMgnZE
6c1a6bhYb+GcFGnKVm8tfqM3g9a9Qduc0JcsStzCQyRElXrpIYIMugFmNBJbG0TNLuhQD+aMRCV9
aDHwUFqFzB/fVlSfjZWe4b/zl1oBzC8QnV0UNC+ZXwb90+OB4WLhcR0KskL/Qmc8keKr0DVVsv5Y
HKGuZQ/6yarF6l2cOWdaBiiKWpArsD+iCcIakjCqjE72OxqYGvTl6+jAsNLZ616i0+ZOl/QrmALB
Pw8uRwxPUBL6FtdLYqKvPA7h3fT3TundaXpELnpWCK61K3snBzk9fRylSjaVaG7Pa2wW1pU0rJIF
GHWHdBTDBSaWT1RQIQ6kyK8TVppG/BYZoaiv7aORUTMpyja2OY2rmI4o/GN7b89sMUPYScnu3Kfo
JpiSTRRewn80275ljstXes49QyuDuC466Rpin+dWVEZfijO8ZJqTNUhn4brGoXb8CBfjrgKAk8eR
WsToDWM191Q235KHixnwN9zGOaLEZSo1NvOIjb9of/EqOuhYTPs2oUA48pW8mmWbAPnMTZDHcO3z
yeyrouWb2lQPcPKqv2gjUHlLW3g3sEfUFz4B+0k3JT+8NHdAOeVUf5vTcHc/dpKfp9JH12K4y43b
BSIPwbhmKEdU9xCa6E0e5V18NYjgCtfrq22krYeOZDxHz76MIrdIox2W/3gW/ntP/pmdeIowudR+
2DC8Pg5/6Aq1q2PGS5OY/tyOYvygW4vpNiAe3Jk/W9JhAY+VspLX4j5eA19L/X8lho8xUvktP8QH
GKq/iorCJyrexg3rXnDFIi75HAJTneqqpB36ZOmY8PlDF/3cuVFf2gLCo2oE3lyR9m9N4n5FFeYE
k89NJidg7jQ43ZwwScSeJ4uj+lMopGxj1vJYHp3yg2nuPCGT6HrK2KIVQfUWoJ3CAHPb6GTz94fO
3c6/tNQkihpgG2btsgDkTEgqkMGittdTvMZa4qhOtcDftvW0d7F/qoKx+3wCa+CH8nSS0iRq5PRD
9ZdHhN0AUsBxnwHweHaDqiIRL9OOZ6XFfl3CUbA07qTnVMt4ZaQlpsb9r0/lxEAGHWLmn++u+i9r
FMBKBoOmda3naBMJWqDd7NrJHHgFSKogpcS6rSJCSjwdkJ4jy/Zgm+AmQs3KcuDeoV0RB6pmEYfa
xkVSCUy0rAwld8KQx6hjqgwH0FZFJskXlMPlCRLMTlwLnRvxTS8yocPyZDXQuLyGOBGRSAoMfDLC
Z1w+llKo5ZIzaVW/XVmLqfp3bj+NdFIdf/tATn9A5UjROf7IHAACy5jKyYGaC2/6ZhQLq2dq82GA
APZGnnk7+6AKqZ7qJKOMboEphVa0UFZqMMaJ2hX59qb22Qg5nLgyX+iLpAJsIiWdWSgqJZV9BIr5
HqapfOIQdqfDmTLGDUyAoTu5D1/0w6v27IDihTmT7RGWSPEMdnQKmK9WcgqIlaax1JxxAjtnWuRJ
0mpaXjniXzJa81nQwY0WURbPVLrufztObzyKhr1yuAJe/RhmUQgWgr8WCnztLO2BPc0tnPs1o+b9
nIEyEwM1tT1n74foQcPEwfAvKUAaprm5bohwoNBP/mZb/kvZkNS0LaaUEsNsfIG7vM4O3ZkfgBXw
UKdc15fUEamaRDzIXTZzprPKXYEwBU9ZHLOgvGLGIhkGcNXrFA2OE5vs+UUCO3RepfKD3LTwm6W0
FAibMt0BeZENW5jfrNsGRT+N/7lujpF4whzM6nWm42nYgU49p23W+qVvpyBGvYvoJ2yregRpB088
Codl3e1qepPBl5L1jjkvNl1g4OKaSgKfUJ4nHZtxGGrNc5KCTSWKUyxs2msElyY0Yit3njuzX3nv
K3imvHNuT/wGNdZDBLdrWo1jOQbVir+TOJatrfs2767oLrcT3cPZjjq/6zl4PMJiNKcURDcRnTSX
6neB3A8EcAz99GVNixc09xaCK9UWOrbqEOwzzCJSx5rJSegtmRHxnM4OghmhN0BaTGiJ84oNrNXr
Vvj98HiknE7FzeiqU4tF5Gecnbh/jtuJtZzfN4Zg9pZPRPbIixawDseeznXb5g8fi+LcolXYKRR9
NSl/ozwQfxRgXXicLb/XJjHnbAXvoaNDGcQnLc5W+O3HlJy1LduQmP7tiAmlDlhuIFQWqlgK0YyU
/g9clo8ALGOkjaVJ4p0IDwdawylHgf8r3FgdiGj3G0K1xJhhJbETp0nO7wWTyiiHRZ/NFZ8P6w9i
A42HCvGNRd/KqShZPd5ktWSl1du9BhdBGDqeFOq609VtHQ33072UwSvas9Jdf62PpdBPeqwcxEiw
OtDFRZKHvOcqLUtW3ZCAPQI2Q3SfvHHaIyDs3zE+srr3yWbpRgbLHFv8KBpLJyM8hBv5OfgO0kUp
uDxa/TBXXxFd1DYv6cZfKSFtzYMTafxHCe/vzplQx/hKcmAosVZHbk+BJ7g50GjlUutcM6D8W10T
IhjXCgmNdbM2/Xt/I3CSifJgXeqw+T5bKHG9nOlq1ka2UsV25LG4IRX8DasL0mRBP4ihyePC9xXo
MebKo31c7i58QeRn5yPmeDLzec9z2bkUkfGWC/FvAdFDCo32pAZfRCuADU3vSi/FR68KuK1bQZ2M
7qT9iKvVI+K0NLPVPl1AiIzwWYfmiFIMtSDLpv5X74mytkpDGdRx7RKtzBesb2CULlCFArRGOGrt
OjEiYA9K78o61os4RmhbH+hQN241gjI0e9bLNEGoOtWAPoCeF6HbQfkaqfoLIoXpr7S517WpcHoB
5ZcJAu34woNwA57hKrwcxWPREgmEUEWrlnOYNhzKjC7oeYJDwu2oxxEuR7U+FbVghzyXLhRdqNQf
DWvomPla6rlU3b9++n3o90Vhj0ILCs+1TbYwf2RFdCeLDDbdaCiEKerXYTVkAZptkjJ4t1vDrYRq
fgNuIur3F6JahIXW5S71t96zB4eCbPWeI1yDGfmBuk1tVBIEDpG6MlL+ZfUBOPYbarHabta0265P
AkUnMmM8NFDkmZ/LJ54P9YWAWYwfsqVeRzGYsZbAKoU3OKQJw9vd58z6LXi3SxSPv25JxC1tMmY7
KqCwOgLBZJ+N8hle7KnAhlTfKIbaqs+yqrQkx+y85Qk5yYujzUH3+S19KuXARTto3NcsXqswezZK
FuUOm/ezdZ3baBLcwcc/8ekANihmHeAClqe4Bms7QxRswes6/iD6GNyG00A1kemqUfyVUGM/1fAR
4X/G06NbMjxREBBLIR9F9OwNIgzGsfYkrnTVmq2lNRJbumai5moU1U1al/LflfElmuduShltZ1Rt
+gOkO+Z2ptmorDnKSEZLoUdB1fwZsIWYFIipgHMrge6xfAx3QczWW8MxdqV9h3pJEJK4QbmInc6L
eNka3eD/UMdoPK7GM/iTZADVJ2uMXp2C+yH1V+a4nFvjlmCSLNrWsmexfEHTushkvSgXIQgT5KZM
aPEHtGNPb5/DYelUwNHBX1x3HfPGM/cAFHgH3cnGETRASDURlmN3MFFqT7E0E2iat0ZWPjnP+JyC
B6C3+RRu+dhzY9aC+M8YuzVGD8xC0ZVLyVyjsZ1DofeXbVrWzi7zWNnBnsYEcZh+W4QY7+F+slCC
1wfmcYhs7j2MG5Bw7kVVY3it8MKsdxfCinWp1xobcgjsBxvWS12Hi9PHSHTif8Rf+w/Fgio51hUh
/BkTKkvCr9J6QQwsctbzChDIjVUUJmR8c2fVtDHXb0k5OUPI8Mrc3NC1tpVgqsRwD7uIMzjbss1P
Qv/IMZKASOI4xeilxRb1M4OxXwICNnMmXL6kGzMEDdA3DFnJG4KERmR2YMQU9maxPw6SnJ/j5IeP
DmBaidgSh6WL70bkzpW8ogcom1a1zMIIu8JZDc+2lKgwTXDDZeSD9sjNse9SsNywwNk7iVn3bI9M
jIU1ALqrOzEbcGaHMiz1/Dst0kKrwhvkFnyKeIJG9gVbY7CS2IjeRgi+WE0S3+fVH7yVxSf7Nuwu
lwReq0gu8+veihqKwBISg/lDqEcuvtu+iZNZ2Yxd5TPe/L9+FZTgwwzj+GOtm54DpLsrecDn22ef
CHldOWh1C8x8KRSB020e3RNOvKiE+XjSyms4W4HlxVp4WEofHL3fOs/8ZxSXHzv+Svyz5LKUJ7uT
VQkFS2VhuR7TLT0dFe99iDNfDriRFngNkq+6JKFXXEtxsPr+JkVNuitvkCx2QzUMh5R/NfZ64fSQ
H8cIiCiQpau03IoQRhIeDh7N/iDD3fpYw4KCAlL5pXbfTxaZqGg3bXOY+wJWBk1ig+zew34jhpl7
KIKqnQK6OGASIdeKy0hXgAjmFVMzVrtp24hgcqRIxc+APtw1JLQRD/HzmxmGwkLxCGN6NkA4Zf2v
Q2lTG+iW1MgVJqpZJIwp9ltXpMBJs3KYEmoNuNTdByqTrdCX8wH7+hf9+zrFJd2DgRPbl/asFsUM
YZcfcG+ffB2+LP+vSTW+bi0Vjv8LcVUH7gcDmLfSbXnX+84p65f9eE/nWD8CrUsuvqn81lb9+45B
+ef7SKGfeZKNLEylkx/MUcztN6iNQ+dfaxBxcLqJbfY5l4nx2eWyfmeJ18txdYojKoKbA4uZpnJC
obATc2UkFqMS1bxJZ1Lg8gyvVl0hrMfgiSQvvwWCo1nqVlZkJdko21VnYRsHPOao2BdCwHbAgrWq
jt66oueIC2BKhAi5V/U8FIkfg9xe/48i6Dk9g+QYVKD7Qz2WX8PZtB70bG2KPX+Sg0OckKyUj+vg
fPwu2qBoN4V076LygyWsBYXXNQva09342Bc0S2uIXj+bkYJtUrOrQCc2EylbuDKBaidzhOyuzaTs
OLfIohwdHXYEOYhzFLe4Ma9hmunNmaovN8C1ew9P/eAJBstBjnrFqXvqbrYGc5lXndBGmRcWxfFK
yN/vpx+CIJ10ySI78kEZsxPwQyK4zE9hrJ9GxlJsteon7TLxTbrGEOCLBSuMsi0m/LsuCFwaLNqg
5LRNLcrnImyFgsvpGnKsS2599Kl3nEOlZBFIwna5lUgIz9jfkR3Gz6wywHRf1uinaRUdkt4ZEv8z
cHnd8rtTmcAx3LwzCv+GXGlu87YcjygMA7VivI5vwW07ed57qyVMwMjxNSDl+1t2MAsqgmcy/gOx
Jjf9IrYxMXQ1uw8YZAWqU8udDg0i4wyJIvr+0R6bod1vVNpnA8FYoPSATwqvu416Uf7JuZh89WGs
wnKCq5QN4AvjiJmDCI2dvcY9Ww1goAQatpTsAOo8Hb42VFQ/ZWtHE1uTbCXgQ6tp0Op+kx26+uJG
c2r3raQanRl0s5pJmaQwf4M6d3dY+sBzop6hO3pV+PM64I/42QZ7weSBvPrXbkw1LvCzScHp+rbP
CJ+b4C41a11pS87Fs//4huqetR/dXqTD32sOsGBgFKxwiQC8epxoAx4kWTRsBgv4NXveXRSwGvvs
isQQmQA/HlaG2RLS0jcEKSRe0uCHahJdY1D4u2UwIl6dhD+hWMzwlK6I+fhl3fCrUlFVuqIeCSG1
qB/Y3q4gS8l2J25+IvJsVr/guZx9tl4tWuDI1+EhpfeGyCkiael13oukipYIzwzbrCJCUA2yXQ4d
7wcEGX4gKSu6iybLJo0mg8taB/wsWZ9HNqjOFmud0SisS59SBx2bKGj6VliBQlAyHO6qHEFTNUBj
wIz4lauYnQQfWsyN51X5qQdkmcD9id2Mve/EsLxVtYJOwGxR6XjfgdB2q14pATJ6Tgfq0F6Yss39
qWC/Xv6DrL1jWj1y8Eq9ZMOPS6LV4RYlBe3yKRPNEc+n/7Vo519xaaJ7fWkMVFOgTXy18ntvaPPu
v6i8UE2fuCWa+wvk9IUAcS6q+MQP1XHkJGl0Qp7tuAQzkO3nZHc6xc9LE3Z5ekZzxX2JUzrxwFIk
l19ftATgTcUHBDV3gFlqsEH7iQgH5sXNT858ANzcYg+Y3wuhs+thwd2bZLjn0QVNdmxxyyFjs2X7
65thAVviyJknnAb4I0CYD0g0kjFRBWPm+LaBguCJqNxSENBuumV7j/a5xDanA1g0NOJdHbtdefdD
hneJkmVIiHE3bzpHxn5k8MuEERTA07y76veTTENVf53JP9uZaxx0b/PHVW2k2u50Rw7Bn3jSqi5P
KvJYK5t+zvkEkgq3/cilu6aVpUatL8tpukWB2v43NxVPm6v5JhuszzOAYyK49aLGb5u+uXB+wmNi
fabTsF1UqeXG/uO0FFva/cWrwSS/OL7jW7MlwrCssY+iELbmaGIOiq27sKXbyA4p0uFhWyJxD3r2
ktieC4Wos9omPsfW+N820Ggr2Li6hm4MaDu6DcpufGVRTZwhw5kHw9c505JjTzMoZmOO4P6wR4j4
PawguycXFLKUlhhU+FbDHaxUkZ8x+u/qklbN2oEIS4DYbVWGeifTIkkJDBWW7kdHHOg7GmXRJW9/
jEnG8hMpitg+VoFqNZkYAn47O7CDNow8wq3xt/3w6kjBGAAqKeL93TTkKFgvz9i14BXxzbJBj6pC
8rt4e7xW13NvCzYTaHDSXdPqbmw67JhB0MY/5HSN4doQkF4JyEaOrd6KWWFOFimE9QyyLLQ1D0Yb
+vOpEVfy27SChPD8Sbt253DH9qclKT3VU9KKAfWXW2sk0BsJz0i3gyAg6ynSt2wvXcj/ZfPUdttP
lrS5jcsNd3M32EKrsc2k1ZMuwnp6ygq4gsrwJlVVdVA8U5MDvfPOmo54LB9AThhY7oXklFT6hmYr
a3KJ0TKjvgze9za9nUmtSolbxr5JiEW+cofB3Q7w8JjaTat64y5R06nhexfWGwhVpuGfngRAsrsf
XWIflDt4B1up0RVtiF21Os7gXH003K4KWa1UXfsyTmGEWc/84+VKEMy9ZN4UHL9NRAALHR4TZm0P
oby/kMYuDd3RGgtX/NLeqCoHjRO2TnPHf0yPARgmzc3NrJy9zjMkLdewzITvywP9eQS6zZlczy8T
oaphqXyLxiqDCyg/dB4H7VfvIPS6Nb5Xgsv6N1QbJJ8bDU5XUX1VgB12fcpYhV/d9SPuvuhkAEMQ
mbw2IpETzF4yIV0saYQmgTsPR29J8eZXuPSnhpZzXVsR6dt9tNqGeKfifdYxd7d0RLGVpBDvwNfg
Fda9hj9GdWVM0gmbdICbJdGieN4GruHPT/1JOrsQc/eUdjYlA9Swqg2CmAuTe84hpf6NqWJRHAC6
bAotsVsGzluYfTb7h7f6/JB5QVapRWE7tktYLcLDxbxRTDfTU91LOLSCoEuPF8WgNFnJzuhMeU18
7Qe0Az7UmhBn8oSeBIpPmWO1ELvyta1YB9kAPAmBBN6b9t74S0SlXwa0j2De/Qt3kpu4QQ/jOxi+
IkL29Wqmolg+Y1ZBm3VtMiTBKohMn8aZVZ6k6OH+5yVSHx0Onl7EOnkzmaVxwezEB6rUusTwtze8
DcS/OT77FyJNA6eELNIfbc0scsUwSAPiH0xFHhlHu4wo7L3+ygimod2EnLjrsOTMYM+9j16ssW9Y
6Mhqu1pODW93w2958tEBt6EOYEE868+Fu2kU5QqbyDbdKig5tVFYJM9MTH/49sZ3XD8oxkuZdx/L
dU55/1hUzuw4ZaMzdatPRTkUiH+pdBWf1FXi41RSnhVUJs7J4grz3p+TqL9wvHHRc5eVzWXiznxr
O2fNpcumoXaGzAsQv8wUlJcx54v0m45a5fXqt7R7jBZNMF5ORXfZyvA+eIcYCLGNtCuiELxkEsqG
aSBWUIL6vhXFmw+RrBmOZIINkWQKddTl/6fP1Oat0VxzDTydUjB+otAhjxgVa9i93zjxaNJUNqfN
l8lca26kWsCKJQrFq5iNTfYiNM5+ZyS5VP86lq14wyeQFAAA+c8KeigxWvMOwHlFW982BAxaCVOV
7S9BQOQaTvzibvB7qUUjECL4pERlIJgK5ov6KxFou8QmGk6dVGrPOLlkmFj5fu6ui8PtqGqY+luR
7RBzlBidTi51GoZSmsdf7mbpnJ0Gye5NqCLSO3JYjz0ajsxOADN5jtXVxbTUxZJ5Kv36VRZZD6BW
UN+0JQ4ovH6iNgBheXXxek0w2NKAqC6aUHLrU37eM9W9DGM6rNr2wjUL3cyvVowT67CtPh+sSwDV
wm8btWmbUqGk8JPUDl4ozHHi64+E3wt+wylTUkVQZyDpRycrPCcfNl/MNR/JzgXEWq9HVwT5hy0o
thXXiKyFQENesvbPvt1KfbYhc1DYDx5BmX4w9a/0382/81Vzc3DkRutRaXFKYMQQtQqV/FxNB+s/
ux8QhEX1Dn3qJEXMNLoF2tt378hc75IVje4EMRr5/0vpar3M6cuJVw6CzAm3OW2UyB7hRQTM8Lya
BxqJW5iCm+13A1ZkyxYDr7bVLp7QcVv/0x+MOd4/EIN5FVTKjfSvWAC423ne5DZ0kFSlS5ydWCqd
39k5qx0xfg1z+yNYEoOFVXRp9dULKIirxRLt2JAGzkTcFis3R1cRs0vOcUUilNq6hG28BX0twY/a
paToS9s31xCDy1a4QIjEmvxz4u2UXivyn+Hy2459URlHZbM8L/IbTEpaCKosGIN2/NWvEZzNGBM4
gK6mea1/x3o+JVXhtx8CSsPZ4gxV2lMv+3lMV5i0yr0mDrxT6fXToIfbocNvCETrtDrXvWlmSqfr
ngtmswx7AfKLPPm7/WNHZA9keIv1MRI9gq0X22GJHODcsaV+wTF+uwumjfjyrkzcYCJR/0I8Gg4a
i6s/dswe3JyI7eCXSIb4gypsanjkfuN9udl6t/ukBCnLTXmHJiXEBM5v1RSq6QaPJnxvfnQXf+6+
UyMqx+LIsLmC6tVrF3teEcIllvebousbdc8XhrJsWbSW7eoMYPwnGaxcYsqDY9iL2osLc4nsZzDV
Ga9Duz67wnfTh2AnKr5OUfgl8un1hb/z1ijZihCqW3Dy5P+1ioxwPW9jcm65l/teeSn+KR4w20Ee
CyLHXYQMvBy4SWS/FmIvTJB229KAp9w2SPOUHPR393AM0fzTE0QrQNcZDGypNQhqKPJUIMeqwVzR
+djL4KmfdIj+zgbZKDkcyt394LSynRnZSDGdOkSx0dQ+QGrBTDVw9phCG4YUX8PgoCxu3gue7np2
yKW8HKz3al7uXmX2DNViWX9KQsNZ1YlelJMNR8KQbwyIx5cbB4lKTn3K2XpqJ+NG3ZOE717z+EHi
cTFscbXUOj+CavYcG9atZorJkX9TIW4A4POUXFWZOOOx+VstbNbNW92DkHn8wJeFORYgiQ0LV6+E
FXjer0edwxgO3IcfyeqkQcJangUr9jD+KycQg/f3DT4aRmTCrPdk/uVU9b8y+DeLDQMjEbh6nd3h
sTk7ptztgLUDxIA7J/JJ5D5xFUlkV38aq5xf9H5AGSjtQYxoesfkEd7S2NWm8kohk0TE5bVC9/ve
WiMBOBRzCohjYAGITX/23cyQqzOo0fwpoij17hqEXEdkvK8qYp5NzQ1t1ScnAypBepu3gn/fxZB/
iY0VRxkzCXJFgdtUF4K13E5SgUAzPpznX3w+Hcs0rqIjOHKm+fI/vHSo2dIr5v6Vx6iJTuaMTIFW
drS93sZuCjyNSt9MZFlIUVXT7BNNClz5PhrCBDbqS95qAIfGYeU79R7y7mixRnJFKueFPXIdI4GH
RRUHJMiIMg/5WCJ0MyIAdduqBpDH0DAcVz4kaiGg/cm3BJeEVHBzuz6Pk1HV1y/CpmeoHU02dI9n
+bnXYPYWVoaGkbh9884/44fZnYwUoJUi7U8LeOO+CfnovRY7iIVACOM7NAESyF1NjWXTe0GVPgpm
gf2JAGeXKpqoip6pH9O6uqntZIp+bErGYYP10I3XDcpG2LIFIXP65nguV1N/oUNvsZjjfQUBf+Z7
tIJxh2WbX/hcqeEMTICWiJSju+T0a4086ARA7LYZu719oKCnYiYr3efpQ7RXL5lHq/LLPO+aDvQ6
mFI06jnGhHF88Exxu5HVRtzXlSj68Tiuem87MI41yvlEHlGp8qJAaPMOZ5fuQBZeumSkz6pOyBEx
tmGu/RAHyZRWoIsWZilWDE4o5gYV2CqzLiPiLmsxEW/ApG+M7g6aSKIwZN6HdRr3p/sUYB9WNCay
5l++xbvCQ1a9QXCAS4ovuNASwKeqifjrVA9HlYJa3ysyIxNB8X5p1zUVRhHeZxO3uU6s5rRX+FuD
0n3Wphj+04SHcY1Iu599d7ta9j1Oi2NxWxBBOjZSUNqJORqPPVM8bgqJ+dsUXz/D+3NeuisZelVp
vWxJi4R+c8fe9shmYh6KUPeCv4E7EpbtIVKIgjfeSbyST2+j2KiyLMER3gjuhEMampLzm4vExGQr
jmn78NVn1w46M/OKVOahVZa78X16CxHBZQoUGl69gYtMqpIXTI8AJSqxTEdoH6uE+QruKSU+f291
phg258RzftrC9ysrsHOg++KN0GEqLmOzd+3Mky6du9ppJccpm1X34hwmIc8gIGQiLfIHeqmzga0i
kJRJj9xb+Fylcmgj6XjZVspotTKqzjgF7l5bDCFQh0g6OnkI736NuJBXRR5oDK98EB6v8B0+V3id
3EmE99vKZku9POvzpC9xvYrjgJ66LPEjQi80mD/LjcacpE3ZKP0Y2KfxKnNIY0tvOe82iiQJBo19
8lMR9h+saXVZKwmqNAQkk1JMI5cyAQQ8GQMu7bv43llUpYdQd8OEiX9Ys9FeYDqW9gar4LeytPk7
izTzu6ZgnlyGBj7MR2PPrShpw305gux6S24l9IP/TFpVPtE3IudGzh8noxIB1K7EhxUjmnPZXdHO
FaEQBCoTcd7a+xaPLrJXPDD4aLK4vfTT2vDWq7aYKXTGfjbJwJnt1z/1xAlDADtTfdq3ml60sI/c
5XTa8CnzqL9htX4EDqYZuWEsNocYjy0MbPd+eQylP0N2TzlAJeiU6wcvwgQ8xZnstNN0TwJ9+NGx
utmPIAb2xECA5x3nLz4la4LQOyZZ+d4Wd7+jdWJYYVRGj+C0tRStF1QTdJP2YSrUYmicjBDTzXgl
01o4kqwHvJT7Br685Ysty1veIby8e+YS+Pv4N8QiOolU+q8eFkSK1YAaKJzxDijHBsmKnd79n25X
eYT4/It+umXzGyyb9w+JomV+YIli6tr4Dy8z4IxLwwuasY/JsokDCyw6qjJDDKW3pSzODx466F2o
LspyxEj1eCKR8D0uZSIygAhfUUsaAJ80s/+7b9/72lMP5mnM0yvkAmZqmSdT9jMUSvePhBVzwdZR
Nxu9ytNT53ZqmncZpNaNHRFK4m7LTZmB4oX/oxq0hActfodn+KSoqDFbkGirYVAbnp+kCIuZFFcl
vAPE0jofJLfvxc/JrKKNRmYwNDu+FVRYaBLFw7DiqcERLwJPH9XxwZn9uB3C9+nR08onRq4uLFK0
WiSnEPMAGXJRxH5fzzXaBp3VztgJIvOnOz8hV44FL0t7MmrXSeK6NLFSIJ9RkAnXnBEhWFj704N1
zKhWyzQ2gHPiuEeyHlmaNg51KSuMwWIP023Y10hXVVdQa/ol7cb7z41ckugMlmfpQo/6ahMUYjmL
GfDnaKB9uMEzhZ1Lf2hLA3CGJiyvxaYVRJtJuTXUL478A/KXpGXaXGJJUTLfCt00afKyP6sDrz9s
2eQvA6WtihJ96LRDfF4Y4io2Y+D+4794n8d5tQqUeMeBqNPleFpIaEcMnXU6kN0SrmGIAK0HtNhz
a6atnR38rwoiAImlGWXY0oLRpZ3FAbdml3fNmApvRWIz2t9mNjxyGskWiea1eSlxUFYISut+DqI7
H5WvCvZSf+RCioZ3uvPipoa4ymvWJ/gwx2080uQVpB3x6oIRdzx6ooiTBp4I4ZFyKr1Hk5H1Mv+I
kb34zgrP9SYV+wFY3KzE9p/HeViYkpULI3OMajVhO9IBj9BQaXTnUcV0RSCG2VpgSvHo5gLKoERr
ouuntJdiyZ3UKHNrtfIEdA50JNEk5UYHiTQEInlCzsk9iOWGqwodeCqvpj7imteLuCawx4Mf6jI/
S/nSXZp/bl1RBB0wturKPT1YY7Yq8TIqwkSV8TX2vqz7ctLydsvWI/tc4ojs4QjD04CT7bUov5Z8
oGEckVqCojnbR6hvfrOiZO5pVxBZrooEsxRwJm1jhLpovE7GQhu0hLrjs6UhIxvASHPyslC/LF4z
MgDBmpOS9HUAlygzvPkb2wjQs1KdUouF+hILhS5FAHnk6WxSqwpNtRB4otI+0/oeCsYaRImZbOVe
PPdvI210nt+C6yokq2jdbls7sEAAr5iwIY/XCbTKmUM5Uv9ay4eXQHv3nU6XVaBt5Cvmr2g+aOY1
8VKq1rHgvFQYSIOaH27w4Vm5pl6gBfaG3ON6vPiRlmjxm7uUvg/uBZPn6wxvRMsDKZBALgmGGVsL
tC+JSsuUM7UZNiK+DidJ8kuEJCpyZKJgYG1YjiEKIjnZbqZxH9YJrd40ssiDrHB0y2harzMoN4gp
QhF46rlWWvpON1/q3365SwQLMqARDKGi4zoEOAhf99IqGQQlR+R5K8z6G/6Oo8P/kFBnS8s/8TDS
Uh4pESAptkHhw6PHqUS09QUjZ3m3nX+zc1bq4RI04pk/XJ9Wxlgwab+Uad/2NjrZ22DAnULBtoJU
w6/Jnqh2CUxrc7eNHT7JOAsvn6qlgN+ZkQfJXS2r2wOiZqB1y9ewsm7seL4tQl/M2G9wozu0i7HB
YLxO8bDjd2kLYkstUbQ4WFJcVS8VtXyKW6UiPfhAMmBaV88g5xqqrRzHF+RCo9AYQOZ6KkoTGHRo
mB4qpFPQ3ZhYXWmtT1JMRUQVh2qGjzNTyolDjL5zumIfShwh2CqzsHN3ddy00QbkFfy9PGq2vBzH
PgjsikLc14q3wJOcHnV1h8RrrXt9RsQGHtMkGwok+jGG/ISdxPteiOqvR8CiX1K6xy/Thd5/aTHt
5Fjzh59Jypz7kktL3tbD4zb69huMYyER3lIak9s8R8HBA5HZ8pKGiioIqZhTpB5ZbYuDpsSHO3oP
e6H1ecXHAw2zo4HKSxlm0KdfJbnuOlGFkZG3iL0sGlcF6rismY0KopF2Pkq7Nzr6V7rl9pgVLgs5
iInWfnRfpYIim8tW7l4PLff34PLnI7x9YkyJm79hxGXHLY93bqe5YY3k2roovu4YRRXmcpbcpmkE
FDNKQh3Q9SdRRtylNQDolTZy/sy8jsLDdVopQG2KPw9B0gYcPiRdhxqYO9NsXic+pP/TVDYhdQhA
bK/HTHW/GKGNKyWkZTnd9dgZGDu+gsz8coxZR0oTp0mYrNhnEpkXWV/e17/PAh0y6A2ZaDiRkQ6+
tB6q3hUTrTyz6PEws/XhXeDTBiY/2EAIz6n2C0tIB8pLCUQu3VEJ05OpQm0orN11xsHu8cO2WYFV
JSlaMFbdeX//ywjGqDEL4Y9DVJhgDSm1jdA4cdXA3M9NOjev333cCBLOZq0YlkJJO7+HF52IssQi
3SB4LUGkzkInCpMHjVwGX86bZuwwMlv95jIVb2SU98KmOZuF39me4pQ8n1OS1Ulg4O9nf6vONEA8
Uum+CfeK8sLnLzL9sc/Cxg3PZ/TkmafNH65hpnwMMq+8DVTID9d9B4LHhGl15lrv4Tgrrx9tnB9a
nhHz6RpsG2bcdoCleWM1zzUfn8L62m++shnmPBuEjxGHhRYvO1VrGwxBja1NqUYzBhBL991K1nWk
aXhWkJM4sI7iJir630qQqQr0+RXSSDB7nELeIw6YTuDjYh7lS96g4NoIP8eyYSHlV1CzKeBYqOuR
ArGvWV8vcxUqv51Rsr4KlYjUpJDKij/A6GwB/1ZOVSB5meIMcHDtaPOJ8l/nC28cisUpJiZBADhI
LJ2Q8Px16DML1MvHKY+jWc/E+7pc/g5WXLMMyYj6CxG0G6wPciagWtVGfNxc4vcc9iq5wnnoibMe
gdYHxuI9IVvaVuuWxUrVNfKZ9zUwg3dg6dJwdbVala/JogYPIxs4W8fmlJDzIzu50Yr75NgkDvBh
ZnEeaDD9Z4h3wXWbXPUK6W3XLKH8ZLoqy9x8dHvldFtuZUh7rvuMbqs0TfW1/jeentI1fc0RwB/p
3cEtn4c2eYNWp0YuRbWEqxaPQjnVLTRQIIT4h/jj+Ae+jPNe/kqtRSrVvDwzKtxN5fG8u7Y5x60h
IU+vuWFVXLYDHRqe6nrxlkNldH2l9x55PVTt0vxvijowwnOSs+zwrIypQzVhkvEXWFAqtRuvnkSd
a58u8fQIMVbe/FX7jvTNtZQEI/n+TGzf+sii0ywsdtm7k4wfGhVFKdwZ1UxOF8W7SALXfqKODUuN
LDg9qmCb/T4h+pVYs7CWG/Ep+Kd0Xe8DYbmjW1fSCAGB6MmGDYNlVkiNmDt6y90ELNCWLHGY5i1h
In0WtCguugmcYMnfqWeWHy1Jxgfeaj0yac1NHm0L0t93RymfdfRrS+0zWj1bWcDEtNBrArmdb8Rx
siX8UIzGsfpmPAa/AlTaB7vl6nLe1DjLeS2+Cy0adJn8Fo1b3cOarPwVTaxtUqUs9ZpskXURYYGv
JMUoxABK94YLAFbxQeD4NP1k12cNb4YiMUAPNaNABjymeov8eZZt6+w1tek3Sne6Q12n7EHFsTA/
FRGo6N1Bwp5Ykhwkasujew/fNoD9Z956ybyNwB9WaFdKkZI0RpAp8D6bYfA35O+7Bh3NLfmzdbqb
SeTIiIHiEgG6Q5WaWrJWgznwffTPzVMejsRYBl+ISyIPA28Y88eoMVFHNQJhQZZp+Ei+IGeC6uqw
axDpK0coAeqBpUP13PBVBhrcvtSt4rB+NAiGS6B71JXvKghJI3rtLS4AWN10DVsUPaVyMjuBF0zT
fHP1BmnSNF8OgKcBOOjqftew7U8CATdisKSpZBfJOt27Oh8lN8D5kRMQkgxiAty99UQUM8T1m0zx
kOT4+tkf7etgTXcsuoLqgFPTvmuGPF/WgZNbU+uBEZlmlkeEpqclUWZcHhixGEgp7uluWWbClkzk
+QC295ZxlPIhxUffsBVmTxGsv/0k19yijS16oB4HCM9BvejikfUN+b1S4ZKNhFT2/sYMgvi+/NQo
8lOXZRbjByLkblMB1eRV1UD5x/APeSGAnOmPNlRyVQLRShHJxIBCEjYpiI/cJJxLnYhxCthQwmgX
N3M4O0ZpJHgr87xrfTnKDgUkNGgR8K1NAidnm3AER46l2uQUuhZOVNjLXzcsYZ3wg/+TkgS5Nn0Q
D/0c1sqVP/JyOTCkgtO6c5Kim8YuVXo8VZPuPPWN8seGoVbu62VT/c8rib6VbPtgslXmHxP42PRt
lCONhpBjO4+o4O3ItdT0hwILYMm3mD81ksgme7bAy0PjUSRTAK4hg3gHAyBt8rwUuAOpuW6J/U4v
+18NXvYX9kxjPV3A4hO/1q19OIOQ+TVMVap7bcEl3o9iv1gfIvZiIgkmkrWE5yP1O4az1mJHkWP0
rADv2hL4g6vTj2oDXpNxWBYenxrrcMZkVlEXNO9EEcCxh51DKZ+x2gv9zBwtCc76QKf3Kd4StnHR
r3/xb1RBo5QUSvUcU767DTXKUxDmKN8pAFIR+9lNTnRZZcDNcd/J1CBHZwbuhnAun3GEHmpS3RPH
MumdzLkp4ZSy9nhASMIIrY6okLvYXYsSqn2LVlLxWcnmMripdR6RWcVQvUmcoNNgHd5EWeYqum2V
MOIH96eCxgxHktmZjxvHJIp2+RS5uLjWX6ofpqEhZ6PnGLxwJQSzZM+mtco2MJ+tAV7Rzy8de6OB
Ok2WnZxIaJFiNpRlXqmET1rkTwEmx+C6J4mpT2+CGlfce0sVwYuUyNV6tWrEgXI8SG9IzRZ9lb9P
1SsF2oH1RLCZqm5FsXrXl48yKvZrZmF+HFlX1IXgLxIA8Cl89isGMx5SZ5Ha3XJoatJhV4bXY70z
Wq6sL401/SazikC/mwW+QR1jLlRtrjXbTRylg+q4gJReqL9p0lGEtbZyM5x/QrMAZT/LzP9KVNEr
d5tiCTAKzH55W/w1mMskvSuUDhSzMIpnGsAFCHKT8wdRvdi2ULF9dBgEIDbLvgU1r1AbKRMf8aGP
oDvazYtSXSFKgZQo0Joxn4MwW3EMzasuYXERYBhte3d7N77zbhWJeIV8r/zU8MvQ1dX9kru0ERx6
6gqLgbe0i/H/r7MEgcIkhlKX13wKG/dicddOGQytDjpwB8lysi6UP+kEn/4V0oB1NES8PG8WOT+y
jwDrUcddAStDVFwhcjQM1z0TQ5VMamE2kJnZrPfK+jvfE7cggRezP/quygo+Cb6lDsgwyn0Qso8Y
NQC5q+gnWxeJVxmHDvu4fhvGo3jdijvxs2PpVSzpkG5MS8NPMrw5s5gBKpWoUpGNkEoytJxbWxJI
2u8bczSwxWgORBkh3khAK+YVqn3Fm/CGtt8xMfxvFj0yNb71JRBYAp577bUW6GHljaCrdUuyl4UE
K9Hgb4eZHRg7d2476xMT9nX0DEjEqxhrJxWTMVTokAN0MA7E4RF+cOn/s+ZBE/lZFUcI7aunBB7N
9piPa5AichbkzlJydHJ4pjf5kUxEkdxDS2m/d0irYqkGruv8xJ6uP+L4wwxjEh9Llj8G/rA7Rhab
iA4IOeRgCL9jJI37XuY5F+JtOx1EkZA0SHImGYMjzINkOpZESL/QSGM1xBXa6+yBv+6qPP1PyiCv
ZiT/7/hM4MMEd1pu11YgcfiqK8d8p6tli1Kh3QUMGLU7flHwDSSy09MzX0A/3y3bA3oMxTRW8x0f
1wElgL5iGi7v9yNZP8GGTS2+UuT/nbYaVai9swfMGlfY4xOar8eTHmTpE8WeLyZJg6/aHw1LAQO9
eV9npXmM3Fvr+Fba7VA/gcG+bWzD2lKSOv4Lqdnw80SpuIEfKSYmXmllO8nxrA45G/siq+daOvFT
zB8VgQX+U+CA5E5jc6WXp+0gSjWYhf2F5btCJjMnwr5Se5huu4+cwd5gIpMOfifAtQqawO8mIcAp
Y2N74XC+P0EcsYk1vlOW9DzxpoO3VkYSI/yank+0PMoWHr9wsYaGXsaKiM2t8ciIy9zZrNHVGs0w
OqADVJ/D04B+ZhPedJhf4zknRyYwPAAcTDtNaVrTUgG6zA4j0xiEIR2OZs1M7uhZduyMroLnp1pq
eI4/zhmsmx97XoiEeoAl2xT37EJeqzpdpmehbcCY/YA/En6/ZqDqGslqQoX36ssR1Tpt3uy5bUg6
HCidVuvpbikAUkv7sQOY4ARlngGJSiV31oVu8kbp9vIpRb1gjVL6HfsR54N+9ut9AAPERnNOdAQ+
Dks7RVkBupAOPp4qI2CD59HjunSP7wowEljM5zHFl0LpyFpzqlZjnlQ7BWR/UVJAzu94BoNuWdHC
iSBOIus/cp6HaDJXHQ/CUeqPtARrDdCU2g2kzbSHuHlzbK2TTp4Ceoa72m3276/+8l8si5rShbaB
OGDxMT1jEO0aJgaFnw87s1gTLooYEcOGblv+V2ZIO+urNCTNaTKsqNrOvKdfImEgId4Amj75N1HU
VFF8Cf9BOeeAG+hMXbzxHVcWu0FLcvW+YWG6sqj6EmC4rhfybQtL+/rqiP1rV8frJLprAxcyD8Rb
x0/0LrzHR2ci8cJNHD0lWkDA3OcNtYamzftNgE2dCES03ooLy9e5Q8lSYaYt/4cUQhm40fUx3lDC
dkQQuGY1fSUNSKL2v9ghi7yL3Wlm1ifbkBc9TIvtTNopYvCi0A96aEHZaVmBDszmK1nvGJuuSpFg
MCbN9PYyM4WmnI9g0AVRuxi9UT40MIP6g63mZgVaVqhbDM/m29ZFieVMpQ20BK12Ek2EtOvsuF7d
LrBalmTJQ4txP9rfS5aV3iDU1czEA1gtpk1P7GYycIXURKDAFMv8orKNDw2uOKhF0Cx0LRg1wTZF
MrPZufB6ZSAiSpn+6VuVtYJyEwKzEhA3Emv9skBW5KpZisCyigQ2T6AnAYB9tup/5vrpAA29gd4G
0/hxp3HDVS0Dy+AH5PRo2gNroh48yX7CZmkqPw59KUc2/D4vFHkbtXz3tszu5CBEz0leKqeofEek
arOq6f0qIByKB3DW2zQFfpQt6oHdYtoMrX2RXnP71d0py0g0nKLVSRTOmk1uF6xduespx4DNxd8i
+BG/AGlToSr/UkbzAI0c1PPXbBlk2rQsdBDQ2VvlD7N+03/15f68bZKh6v2z4oFmdaCcPH3HS7cR
v9nIEZpI7y6uAt/iHVet7AXbMJsOWYj2sRVd9yb19dfneq4zWXWyQcv+QeW/HR4CSBO487cPEn4I
TURvpWpb5sI3qNYiw1nvSafCB1tutm812oZHIxAQhPpbb3udAGVRro3dQ8EYEE9tTFim9J3WuJaX
aZiJUuVCVUNScdpm+19IGwgURASQa1fEC6zBRj+ncjV3YGdWf38jb/j6UAnaugag6ZUOwAPLLPn7
lPnL76QkMfu/KnfEgFk/CX36Nid1U5BnhnsG84jK4A96q8KR+i7xhD7uPAVcs6pFnoGbMxm31mER
/+JfaAmDSdlNJYPEvIY4V4rXJXjItnDyGNTnJseDbE+w/A6h7wznOHUar8/Ekgbxeb2sC57mXAdU
BMQghXxadHneKdJZbiWpZrBdZ0vCIMogOdmB/fiMbKo/IB86abBW+pKjpoUZDWiokSnJTkBGK1a5
StO2j468RestFxl+ySvYO4pxGa4wK5BZn7sxhrd7K6Hh8O6eVLTKVXkeZ8Xzp6o62yVMwQQya31d
y7LZWGvAezTckV4YSOMtp8k6g84MbmGuugPj1JdLqVX8RMqIWEXHZKx5FoJTyJTCJkBdsp39slNI
Katm1TSJ4wEbglEf/55wxNBVUeeYy4DgXGWE9vPKWhVgkWNsaroG1D6mecQ3WqZuN4nuOLUI7EWM
bXAtuB1TlAmFz+QAmo9NU9gxgYDUc2D9pOrq+oeuX2tWwWqMJWTgbMe15945yPN9ihismQB9KMZd
gIy/vEqiQEG0WI2CyX4ANp1/U2nVSxmifsLjp9pV5bDR3fiwYC/bQChleteKU7W8I6GZp8leAAJ1
ViFQfHgaKMuglxfflrWOyKzcGVOeiMjAvRltuHKFqMlq2QfRrKQzhgzdz1dOmY74y8OL2MzUHlsZ
ZHY1SHvgimMfHDAgTv1CDCNc09zwlY7YIGH4YBKn4po+ID+PmeZNnlCis84QIe6+ZyJyxkRJ5Kdg
QAFVHIS0hrOP/Idfsr7qb6ybRUfCDENNTsjNPdGYqqs4NpipGsYgFdzW65kHNmyG6vox95OstBod
kE9XEj5BenhYANDsC9/uP9RRecVWxJZXyN/cqnqYr5MkGlTAxm1XEMtBKs8l1his0blxYqYr3hZa
ebdKFqZqQSqiCs3PPpE3UtQXssYPp8T+q77cHYxwkMhSuqL/r7kOOz8Cq8jbhCzlZRZasw3Hrb7G
WyxC+yIodiTjJtpsVUX0kAphdDyLHfiMYZv7YDRLlesM4dMmIplMXyQQr4+/TZFEppH3dGbfAQMv
FPfwekml+CCfBHDre+VqmRGs8gkIc8fCV5BBwihBYMFgevqe0qkeAONlr5swfQuy+7pHGOmDaiiE
LwzgXdf9tjaDKMYBg7leNhjdoo+Hqw5fdx3ytP1deoNWjcEo9Jb19WuVkQBo+axhqhDx5z/LC+pq
colwSRIXBvfD2z3t78uwJK062VrQmmsy0v/NjBSL7WRxbB/6L+Qa0mB4FzlXuVkplMglpa2tWCSL
GhyuAohVX3/P92Thlqb3Aok0xa/llPC7+f4zC0dnRZkojlDMzBDqdNLto6HZvzCvvYsXmloDd/N8
xKscgFaJDkHR6A98cPDjMZhVp99tVG5rPYVZTGEkSBi3j9zIKtx/u9Bb5bd0lF8Fust9A6RmVeAE
gFqsD48BxxtL/7oVqSit4wiyrhQvLvhJOAdafy8IJEczsIhF3ywe2EQubpkLEZYxqlwPiu25c4ry
kZ58stIfHJHcXNYfRFWOaw+gNo4KQ/eXMytKol8AnKPeFSJt6lUcq4Ys17+8CkI6Teb7IIIhOM8Y
XR7bXsnyWbejUCu8uMKen6jhY2iyz6l7K25f4IHVKmnH7jejyhSuWKI1xdZquQ6DmRFKrlDdseZy
5raAYskpo25jUqGnU+4dEKlJvt2S0fRpu+VkVkJH7+ZfoPFJKXGGiRHVJWE3kWgnAXbw0alXOR59
mt3JEr5kQ9zIp6M/jJRRd34lGGDOkmHT2dI+nVC6CHK9xhQ3YuL5I2p0wyWtB4V9YmDgS9v5/2ex
fcXHdcxKYCgR8kNLoiyq8ew12/v6rQ0agENIn9M7j/lj1+uHgwXLDg1EA7QQVcl+ngG1rG8NIrLx
ggY959nOmfgh3qZMowfki5A9sq91Z5dKWy6tJ5+Nm3xivbsWlOExfmTB3R2okVovv8337nIl7LHp
FBMQzqbdRe1cPrtsJO7yPxYnRq+TkoSqfk41QqmuZ/3aM86qRR4gQ9NzJk9XiIjrxsyfquZ23KF1
RpjEvUiIR4aBTTprGviN0UpQixJ2F154V6Rf7BGJl4dsLu5Becf+qUbl3QZQtneio/xyOZR43An8
z6jTn1rT7fkLhyj71MiUpccKpVLaasayQhLBkXc36ueQm4/jX8pFt0uaeLWLKeVKxGIOgF54OXSD
DbFZZ/NFfV8anv8szVcyrQ99Jj6QACVDD3n7d8aCvn99kWVQOf+HgcgzD8AjvDV+yoKKSQV3ud8x
n4CvyxTlNRg6E3PfwflksPIEzHzkHcWLTC8J0hXHr0KaLq8wyBO9RJ716dokkw4DiUO03qQD65LU
KtgvGbaeXhtrautC22cNVdjtrH4QUoD2lMwZIo20MqUqg0eUPMHM1OiXCnVj7UxF4hnHzLpSqTOt
ApiJm0fO2cRMf61s/pZ1KLYM1XZRiBn3TlMCcILx6u2r9NMFob1souLF3uKcUXwcDa/Tj4KifoES
Zfl8oyrbj+YvKpUHZKsW4DNhK2QfCWMipImHaAPEHtawkM3LnekIoLtWUdhmd753+ghfxBfzFTie
K2qssYJPyYM4M/Ens7iBNFA68ip7c8n2o78yzSRcbBj8gNz4xqoSjC3b5laUpwPIqWDc73HJau9y
24yoRezgUXBmDImQ17LVqH+QcrO2kjqSJsnzHyiP2D7neVH9Tu/Cz2N8KtrH1s/izTwNC+zmDg5p
U9QOBFoQDRpEMiZUpg/uFcr5y5+0Seh2oOHv5LgCGFWShqp9B70CGXO/NEJ8EvNHZDbGT+bH4bpk
/Q8sDXeWSYm2WC7EmVmJOjCUaeu3GY7P50Y/tSm8+SGIzKtoyeVJvBiUgX5OZmT9vNVxYAvP7TTe
ZZ0POHSVIHGkyTj+wpCugg+5S1GMkYRPThWoDpSa7iR/eRQsPnAoR9fEP1dnfTdx9z2XTTPvmbcJ
ZALyZEuf3X6bAFN0dJdUt1LMCiOInVD/PMxsURfHhSqGQbdxVBLii1xdYUFY3PThQw9K+JCzl8ZY
0dnxT6LrwefwXLZRgp0dnq5zBbF60OiQAyh/IFEgLIxtwcGE1KJRFHw8YnUTxnLERlr2TfkbCn4b
lbSwdspk7of5k1z7WF4hVoKSSsU914voqPVpu8Ievqe0K0vai7yehCn3iVRbuzOwiS0NaqnVXP+2
PCwKYsQvo581PGc2S6UFeBAFyb6Jwaqzp3r8R8bBh0pfwsdWPAae1M/8ijy3MY3K/gPqzgmhrz+2
hzst80u9NQI8dYox6JZUatdgBzwkww/NBnO2Li/SEKnWs6T/OX+au2hHcJSc1pJ2MbBnIBDKvIVL
HsAhCqh9tL0/U5HiLZBq7KTIYP8rvWYq6Jq2ccVQH221Ihp25h1JeUg8jipzbNwOeoWXWkVTb4Rz
b+IE8lK8z3uh6KYG7WKYDxkGcmaHgJeIvKGYpnS2dbccfF6I5CAWyH23XRqSLg8xehCwvM+tcEjl
vK3GmxB7EyLn633ELx04yas0r+Y8ReizyVPt0OqLEWJeOBpUdjwV99B8AgosRkxhboszuKs4rP+U
knCueYBW6o+mESr7SqrduJwh1GLE9b2+UI4Acfc9vgdcnYfHhAhDIYzhDzDLjVGdeMCmZGJr/Esj
WikxiJKUK9sOZUGGBiLg+H5bQH6URdm5ogEXtmWktfiCfGA7WLdOgEc/uiszK9RJtEk5tiFX8kd9
tG7nH2cS+q81XwoLu9QqHae+jGebNzmUcTHEADD1OhKLOPhpCcLHbbIyeb3IzU+TsDdMlY9qj/Of
a2vJknblgZhaVGowsORkJDwIYW1lpSOAED3FucUvPGJSd5wcZc7jd2Q90Mp6Lcvl67GubWbPkaaE
k2HnLpYA5yv3e+o504t506ECNUO252kT59mzLaSNhu6msUujLJkneLE/sEFT7tNxCBhNPlCMq/Q/
obxm2BpqAL31MDNtvXw4Ic5PaiLVl8f8MqTHHEIX1hiFlyepZY+eVbnvUOcL0UP7XBh0wbY4GZJ1
D79WkYAQqmEWidZvc9lwYr7k9ZYHks3aPap7dwy84i5sza78H6DKvmCoKxrtqEF1NS2HnCFQUHdh
atR+vh+4uUg2RlG7qW1MlydLl7s5IaPnRgwHs0esfHLYEkadw1YfxeZokx2Xq6ljPayCAk4dgSPu
Qnrbwkpdl/SbXzt4R5I6UGhWEATEm3IExTafaYNe7P1YiiIHjLpY6oNYf5fKuhugo0qNN2rntMmo
xUO/LhHIDmrC9ROU4wrRQbBvMq/3oZSPAEQG1KE/GRh+kHyrbihskuCX410N2UD798Ds+OynjTrM
HKF6IAqU6RjJMzYWpiB+tBjq7xuk35z2WMg70tiMAPfjMl7M+9bdW7zKHuQ9NYZwajjtl2RRS+3n
hBUy3e6NV99s1zLT1zV5vgypRq8tfza9YKw7TPD6NR9qk4Ml1xrzaEeY49pPNmYBAhwc4i0tR/BC
RkUJ4894vOgFhdmk5tZoms6wH3iyPdgHqI98jjAFIhGGUucTZxsruTnjqWk2pzGyMpLU3dv1WDZb
dYzBHs+9nkTK/1NfCQwWigy5r7uB3+96lggjbq/hcIB5d1hbYpTkuEKTWpg+8LfcMzbfsafbL7Nm
2n9KSgQHPSm1GupsDINdWXzofpBlRbNgo3zI9eYIR0GNdgPb6K0V3iPNujFwJX4Acv/YThJ5//A4
q/nitwDLBxgfBchNcRb+ka34OFThjecAr0u6QTAn632gRUlIq7wDX4wt080H70O4UgN2XcFA2J+T
bX61ySzFFFIFo7keBm50ftm7NL8pj20tcVhtwNXFwZRd0jECoVrqha9UyUYXQjwiyAhuwtzBR202
BY0HLj36DwZ6P1g6+WtQXnTw5TDwsubnmdgz9HuhcX3TnjWgE+efuBpXH9DS48Mugmt9+10kdTsQ
toO3tlHyDvJzCpDEsh+i0F6cv0QcNL98iGgvdv15Hi5E7nkQX/JGqq+xYKs2ZxYOrjnjjSujo4X5
WoxZeedE5ISIhZtSZJ0/CnpU6cvjiYcryRClpiU9/liENPX1Wh2XjIZf5evXMHPpmhIKj+yOaGp4
6ouwZbq0MVlSpJ9jUMq6W31YAONCalCYxB4wwnB9IuILUDQZUzjGNs6z4UemWOj9nagr5LIG19Al
/ZosWtVceHnSyTUIMYOBL/9MVfC6kJ1ldgXlo2W1E9HDi+tADICby7wuFHo4r6kWwuhNJcvvIY4M
y4qsfyo1TeEhET1QG5gHPfO3ZZRqLYcVWU2M+4VlyMbERtdLTHk+6UoOaVRHyOjgjjA0Vh1ZM7a9
5WHjpOsBPDSLhCGYXXSqT82oe/539dZpfeN81ERfAMx6LeOQdOqSrCGGDfg1XDQkia+/aWR3N8NF
y6KOD/flvDVDgHsKCKslbCbEEC0rdigC2yhg47S3ZmDlGyBJqLPzDG8gio8v6yyZs8DSfQ6Cqbch
NwjTxAXqvlf2GnDY3vSK71SMTKj3iK6J1x5mI7CwdubydRXVXAJKaEyOaJ238MxcVUXTrVAuwBrs
d8Az7gajnZQcGKzx5Z2aQZ5OpeXUpA/Vug+b9+QM4gvDL0dsGYU2kNT7qCqvkttktVnYl9jUWXRU
IrakZdmT2lFdDAQOUEBGqsbnipovmBFXbIeXPnicU0yngV/1dPdyGsBlg4k8eQZcT8mEHmNORKP2
e1a4yyxDVF5kIH2CTVMnksCf8ttL7TCNwl2G9TfhG/smuZ5IsN+iv/NaTuf/VPnfWYy7D+bmdzsL
7F33UqF7GxSAJqgrl4SfmwBAxxKIBKxmggZR5F+Ej9xa+d6VRai7zHSJVBZ5+K0U9y05jegoZ0df
lPxY4rq2gN1W1Pg9baa11I3mYQ4ahkGAeopgIwR6WmkqpDoulxD6VK3feGnbvyOG85Bw/hYHXYIh
hSypuEIfV5ToDGczmc3EhnZ2g9t922JXAuxbbEQDxDEvZZMNaO1/xp9oc4LzxvuJn/LOFOPq+f5A
EvjioPVDJCFITEVwy7OA1DV0ajow3WPlhxN3uCuOmWkb/cCSNhNUY4y+jLQ7uxTvol5FGphFf3y4
RlgO0BVFfAJd49cNvF262mhFFd4fNbQvqMZ5DageuW91MxwAaojVFTmlfAbvOCh34FLt845nILzI
tEE5qGH5mW6MOhM5Qd4Z/57TXFcGCkgXWzIE2+A++XKj2Izfl/QRDnwKHRcrg5h3EqLSr45YJGVE
kRQNAO8XyBdPygcNMhUF2bYtQHfC/Mk/lczaTTgcjtYSdN1ALuOfFGgHSbgOroBU8Rh5boHSVdkI
4jULBO91F40LGSbbapUy9SXCNN68e7glJIQUGvQ45/LERCZdmsRX7zKHGEGHmR0HI5rPS1VWW6/H
0eMgctN28UKobjckqR3vFWfip6G6sWuBywCGaqRsXoCk7j3WvhVJ3/ZdW16mCha6Ba1MC1iWO/PW
vpjH5dnVQxRbH2OKzpikmhcbA412/RyHwhISAbHkMXvMr/4MzKxElt2/JIYhcZlO4Tf00kwwwFG7
BlZxrl5yBWRReniWtsfmJq0R3MTh6H2AA6bif0fTIBnW22AaIGDTIQCdX79UlCO9S3UhbqtOnaqt
cmyHhoQweRnSPVms8YpEXjXnHssoQvGORK2VXWz6b0kyGrpUBBrvQ6YWNv4OQjAglhmaHU1mXwCW
diVhBu0TnZjJGCwx0aQdnxu1gHLkbm5N9wk/es1MgsDydRf5xcuzkCQfaRyzLG5m7ES24XPTA4XR
umln00+SZHFKfbGA6vhyoqza0YB9obcE7qoG3JqOec7HoMzPrU2TQZPsKV42ImX+e9PfTVTTWC23
5ZAKpeC9ndJ6xcj8Frjkhvgf8MuT3n6Vw1mDfaUY3dARjSLetdCMme5qxKY70segM7uvbnppYsWm
j9bZQ97J766mZduJYSdPhUPxRddLjtJa6QHqLWYtc00fbMny1rfFew5XfcRx0Y8bygKiJ5lTuoi9
A1bInUG9X/Voc1HwKS86AlE0bHmO2cl8pB0OiQzv0GbPiw0d0SoJHfp96Fx/BUTdibU3PS9vzLm0
WmZZZBmDFQMW47NpxiQjjj2U35Tv9tarrtj81XOdDWm5fGm3uxSDDfHn6d+k+5OcF99tfdo8UxiA
6szarxsbOnNRgF07CCx8SKIQRP4VZb0K9um5UYkykUQ43CGBbqGYpMHIwSX4H3QZm6ZZftSdzMsy
p/N5LpBiD+bplibZpRI4h6w8P41ueK4tX4Z2ARxy9iTSjStyW6Hkm0w0qP6MKz9BAJe7wcMiGUV9
TsWU0Zi2868FCOvmDxaJ80617ELOmqUhze8zCwXyIs0t+wHWtCD45c26pa9187kjPss1OrpqozFA
oRzjeXsioG85aftqxW3dkj7PTNBBO1dTZKgbJ2eehyfbY5CTr09DZ/TsbP5Ahn2CWtLA8ejWmTQd
c2hH/vdTwci1HOK0UNTKLb27/UHqRdEdmkIC9vJKCAe7LpUbOBDGwKz+kuIMuMq/9VPtbs8ygQ4k
BEgmHiv974SjNlgcw8kNJ8kEbJTnz5N01Y9oe7oO5Xsz/aSwzNJbAH0E5m3dz8z5gQqZSXi7KTAJ
Z7X0ZBPdXGM72M5XDOTijj9JG2eRZPcdXI601OJirhNvIi5lNLhogIZfmGnYxZwB7/SvJhJ6V7VA
E70khhZ46LGF4XQyBu8tytsmVk6Ygk90LAmM10lSlWPFTIfBUXY1Ifc7j+5nR/UmBV+jOrm1YGyi
3Wlr7fgFuQAYmGlMCQVnEfqb1ckb3uxqVSQ8nRTGo++ja5CQ0hxwlFewAzL9xWj1kLrvsbm01xPq
SC0Aqy1XEVk+26/r+qxoCgOMEw/yLxmqsrVD9TUv3gxszSjtekuueQXKHMXLhBRcCnC0LMWpiF+5
5FAAHeUVYJUbPMFrOWC0Jzc6Um6XGrt4fJeR8rAo9Y2qiRPEVgCZa9tCMikSWYLYudWW3pK1nEOo
zfS835r76wtKioLmIstZm1r5cfiUJAbNNgpAX+EOWlBW43SUpQx3CvQQTE7X9OQGSZlsG4zN052o
6hqcJHnci1FGgkSbgTfua8CoRDvFOqa5NAVgm2+ZOuhrFuyOtQTDy7lT45ErPNrneLsfhBdfDm4s
2b4SJTQ90YQB8IiQulrHOofGxzJavEdzg0TijzX4lxZA6I3MmffFuvQS39f063O4zglHMuDOt/l0
K2DH8AyRJHqtbEHvlivzI5X+DXkmSgu1+8f7XxNAU07qYP9DGicSOhl925GyWMXBrMdGAfoEJcXZ
EKo2RtUJ8+xZzdRGUtkQvDfCzwmkCf0N+kiLbxCj4RwXEfsY1MMGZokThWnYI9b/ZqO6c23QnRDN
2kSPKADr13gjCtJbRKxuD3elgAHCLZAQdLSRFgZnbL5JLRr/v5OFhl3KZYW9BCnNUTx/UUDJXNoR
SomU0F1VhrSufR71lzy9pJspHNuyFh6lTOKQaNuxoA/qgpV4wShrXW66F16eiiGFD0BS4enSWDS4
0Cz38zuz5tS58DJRsINV/g1Nq7MDdMy1eLeTA8hOV7xg5rQrm35RIB0vEFMVeMLqh6yURJ2MsBOw
hVPhtwSAR/k8lXHMaV1WUM8kcKEKONimhJ1uqcnBuBf5sdIvuvwd/j2ibGmkbbBKkCGAKaJDg1e3
6dbtjLgFaOM5jU5qaP271dJ3cFuLmfThOufDvL4yWaB2Ml8HmoXBklnrAHBXR9CIIoqyeFu/wA+f
mHFwuPesjojSJ0mxk5VHJSsm+DsM5y3lCgHnhG04Pr/g0eKw7/tXTIgqCkL0LTopRG4DrLadp08k
Equw8lcOQxezyG3TSV5h6T6QaR8TDkHXoNPZdnCPRn/O2YK7uT481gIeS3JT9FmUkAOJjrSVak2W
bQLtfM7issMprgZz1cMHo0Zm6tMSp5/NYg4RPUc2SEl/5mHyg+kAzNnvXtrX5P5uWSwceeUC9YjF
MPGPWXkF4DKqb00HPWOgTCQSa4wKRErBupEpnI+xsI8+fFhQkk3G+h+ijN7bGwHcL6eAkc63+Neh
H8tx3fv7fjDGZtI2UhaTwcET36sk8tMAmkprQTdBnrgGAkUBktbN8tRTVqwjiw9VWQ1dIxbZLTt2
Nb2z0jt+aj9AOJ1CC2x+oorkBjnR0N5PO/80GuoP54cnCbUxAaQBiZ+X69TQVrcTTr09O6VACvLI
W5UjHJanCD8i1HZxeH9LsJvElCL7jhekNQ0sUwLQhYpCDyVIypDYA+ILqsHXjLkFrKv458FNnKN9
DpB9/edLVvwwIAqaERhjH3wdvz3OS5e1h3txBUQz66PwKdtgwpXc2+o1nhUW6dmxSloFKYSDMVrQ
4gLaA0tYM25XVoSjV1q3J/zqYron4nPEu6LFmDvKmhnTMPlCNsfZm4MGD9fbC1hZZx67m1VVgmfh
jgqqMGBYA8NPJ58RfIGbFLNfukXdoH5h3Z9PktzZ7xBpHCzSSzLypEjO6EnGaWFgT66a1OAbp/mq
n9sEre41vF/aj2+c78rLzO8i0eOZQZ5y3D8sHYzMU6OFc1BwM3tSo1vOQGXu/gxJAIq0Elz8u3EF
at0I0Duf33Eoyk56bku74kza6vuRmQV8mwmhJ/taCZ05qr7IpIl9X+qN5YTCqID4q1hf6OiSoiXz
Vzlq1rxdKTASsfnyIY8Gu3pzJeC87YmTuU0ftptH4v6202uFTWwCu4WFKoTVfb+EGgORwW6oYl7Z
fG4fCmw4WW+jB5P7J0pyBBvU5+fqFW9LiwRd1PocVpLeqXiNlH5DJQKyOBRKsDAufEPOjH5DF5Fm
VjGotIGX0Dxbz5FGYkPC7cbkg2GPyn+uBZbJ5KmAvKlZlBOTA+MS+eEx+DNKsQBOZt+BtFyxI8qB
9RQTVIdeJV6oFyAVdenyK26WkauXNEGvKgaodGKkiJju785wZOPukXR8inDLU7Rro5sk0Sbg6w0v
XFzOtTT0rQBETeEy41AWb1ZCwXa/yamgO+oZogWthTYFpovC0q/SLz7nqBeHJYcs4HT02h07Ta3e
tQ6t+tB5YuGO+NMKbE2z4TtL2DUTasqYJw0dQStS/KFj/1dzM3NSQpW1dVUloR6XfM1D8ydiWzJs
D9hpd1jk3Gf+9xgilxPEl0mfb/0PH+UQcIgbbpj3bzfH8w00aTrG7tD447+tPRih4dHCHN61pU9g
yPK4Md+wD6nl+3DStM0A1CCgNxhkLY73BHLIjkDr95KF319CXbeFYP6Xh4MCEBSriFHe51oM8r21
7P+OeShhQXch+TU0oKrl2qiCVNxyFLcbaDzDv01QrwantLhlWgZ+u3PiZzBb0r3Hf8TnUYoH9OvE
/o9HmvXXIR/HFVjFb9KrNVOFraYKRSJGffAL7hTamzrPx8O8dFaHX++Kc0V/9sbUQ8ktbncOI+vO
kIwr2/3hpVdWB8VOqN+mtv6D7ePUgKDk1pdr00R0t/5AvTS7zgG01JS/VsRr/0FlwAmC5urpQfIu
D4KwKHC6NbyY6pQMJUIAl573Fdcyh5fpQGaLBBn5/OeXo2tZOD9KIOh9/gh1OKQDL6OEBTdF39gt
8QtFWNEzn5w8kljR+fS0he9HApyAdoY2xu9ds04xA3iXPQWL2KIXt4mhYuF7rJ06PX5OLrQeOeTv
ALAV1PRuwEB0XnBjwcbesGa/bbLbshxIi5FzXyMK2TTHOZYRXG3MJGt6pOBPQyb+NVs/oXYZoNLU
lJ29Gq+Wvf71KmMmpFnf+Kq1cMhtaqplzxqBRP0PfjCwMDCDlCApdF703sFJ0MJdpfV0n4x2HkVh
JbTMtmjU3jfU7mylFDhNc6YnP8XLO49edReGhIU4223yC0858w2U/5aWU0fG7EMSFSQJHO2IaDTO
nw4xawmBBnqKz+LVx5o6rzhp1PJK8XW6OVCkDkxJFZMVlkCtH3+BMp7Bc123KJqSpC1ua94+8jPW
Y4v7ynFCSiQ1JQv0NR2Y0leUjRVdY6GPh/NnEseJXOJTjcTEGAdQyPnuV/jG56MK9dT0WyNsQvwa
DyKj6U9ao1kj6LvYB95CeJC+WzHTIkhg2G0W5kKc305GLNwkWdDjG8eCeoO883aIHbTn183Pl8+c
IOyE0FDzRVNNpSIELgXo3ln1FI9F5x/WMw+GJP5z9BPD/SorRuyqtJiCQtNtDn9Z/hwKUqjXSK2n
ug3gfsz31fzYN/CU5J+8KqlKB/aiN93SLa8rkU4w81gSCcFi7EpLwX0AiuwgeejvdMu+g3ilugSn
Hd1ypu1rU+krb/te0+trgwKNpnzblIL4feemYgQ18SHvxodHhcJzDrGpY6ZIOvWHIQFj+2XPoa1S
+aSMwQbDHf0f7q0hmxVb+4q6tlcrr2Za0zVoM528kt5R7Rl2887WD/a5NwIs+ZYJlzJZZrh+ZUP+
3h8pMoTS8qZinr2xzhD2TFSz9WYBhpfj2URbUMYof84anrUTiHyM/gPUgaNuYQoLMpxvF8aqF+nv
7tYsaS0j3YqDpxWXv6J7xrfcjjTWdafGpzUiQbRbcrVg2/xnf6adQCN4dCQiwP+M5Je3t4McJNm6
k79hlyMufnfnkcvKjqmbFG7VtEOyDQ9YvAmO+c90pCgybDcPKsaFqVijpTXfCI5n0GPKxX2+10n5
RiVYD4R6+afveSTpPeZ2fFV+vwXMSjQdCSII+GmHE1PocDa3AqZE2x/wIEa/ugczUmbXOk0wA2d0
YQ06ojCSfwxMLT748aYw95fcVjJmQ1DW49G5gJdqKuiXVsuk81+mhi8WXpLtYX4ePiWzBsYH3TxR
N2eU1d/iQGkAAwZpYxRcsDF2wsdhlswpVyhN2eCJcP4yswhidVZaBo2vfWe1lRfHVZ83ExvfuJUx
MdZaSBHGz/X9Qq5WCwfPw/DNQD0UFh2MdOUjxdenGuIJH2oAP+63J9FgkgCC/HU8wUR6VZeyevP6
1wa/SXPmvDzArgBMfFVxSGdWj2aw9Gh1TdZ4Wji/pZz5Q/uSrPBN1n5aGm87in0t8Cmxj7yyH3uU
WK8FW5ofVEqL8YOExkLC9JWjhGAE1aO2KllXQ4SPx3RhN9eEc/4fKLtd2AVejTD6Z1J88IAbQJvC
cdJhmz3tq5GMvPtj/jeD7jyck4jefhCytWATKjuhM5FAPbLl93YHHxVnkf5ZnKNPR5dRHJsLwkQC
CTZfciHDCSce4QywbI12qEBoQaFDeJtpjJbUmEBpSdxgo3T1Y/w68N6E8p69v0Q3cQkKPl6dm/Qi
/zMTbn4RWgFqcTnkXmUwBoYlpL6AcCrTpiD5F40D2WKIHovraLeuVt3WuCnz3h1jHQ3Cfn4IAjeR
tq1/NWXuYeeWFZsWXEPJIGixeTymUz+/9s14yN/Lv00ryP440ZJy+HiwNj8C9UBo/d4C2yz5OMWa
lRZuUZeB1vct9cq3n6VDlsf+yYuinefGCS7MyGelItLlxweO3RHcErZ3RsidPXe3zHYShuxkwH1Z
wADdha9FUyauLafPW0ZGuBXsqbSVbVXwQTv7odrqOrbHXGIuSsMAGS3DjR7pjr0SFIQFAWm916wj
uKKCom0QA1OKu9SoQ3KmjP05CCbw4XpADsrk6E8FsKFV9NSvL2DB1eDs016k7CETIB3F8VQsjmH6
VDDz10chD77tERbC7AOd2Qz/hyRXt+phRudtqGzJsnwZJ3uhiDis7v432bXwPcJXQN2TzK2LPA1k
pPJtGva3anmty7E3PPcdwMyFF9U+qvU6x9jB81wB4CJKCq0lxPancFUT00S1MhPt7yoc3sscCAxZ
c61nNZXnj/xNL7H6FrxYNj6OmKrxJuF17FvIo57I7XXR0VLe9zG2041djZA8TnQLKSjBLvGqfHnR
8Rl8X8bOTtqsR3KAHh9+8nBV4wieEqle7nHaNvGK0xaJShsPmhd+9XLISibN9iPC4JHKKdnwc3tw
uNgzo2rhxV2le8PRPB/v/ZEScjoAmyby5dF+odLRkZ5XiFX0cMU6c/RI5JLv6k7Uhax25JAVXprw
XYs/Oj4CCM2QP7dX28GDS+izOnWTKdbuk5xRZAajQ9DtNdi3CWZYsu038HWNm5OT7hYQ3FBMfW7i
i9UjtyBfF2qjC/CsvVMXp7YH2efD1vf/ONDYbbJmO/x0W3x5olTl3ux+o32d/OHTc4pBmr4yB1Bk
OmqGvKnLUI3maiRD4q9oZ2Iv0lRlenxbeWomUvo2US0apXz4fVQx65yFrSaOauZ72JPj9Fa6Me3q
zDybaMdWaDH+DsAf9rGZVOUtEkkjXXXWgZw41iO2AJD078f6M/8jnfyUK9wKp35vt2xD6TI7CS3C
ZxB5dJD9v8Q8zV0Vk1ABz1QExb1pxqoj3VEgU5n/QWj0fiIJBF3bp1ie0VsBtzKH1JoZn7rRDkXi
u5H8YQTxK97qvGuxAhFZeO9TqDHaurBcaaRpom/Wbci9+ADr2AAzBQ88uYyZ27T4i1h4yQ7tsL9F
oTNuzHKgQcsiOO/sK7mGekQstPt6k+/sY90sPcDQ7PgsXqNu31uq9QDgxtuXTlzwseVUaQDic+S4
s64j/+GS4WnttTxTEudp2w2S/Ns0DtdipTw3liFpjDoxyv8E6giaX0W7mf7SQB39mycQ8rdonMpH
m/pSar7tZuL4Eq6he0otmrBARC3+MA2KvdJ8Cc5F+L+s7g3QAseld+O1IwJho0hZJiwNE1RHrvJ6
tvKPPCXiCqZfTWSF07u9j8NC29ni7IBVk2AeTmqUxGLDO3rAmArV33JDzY6rTwXSwenyGZjSZFQy
K9TxaXXHrNKC45vPA9URbic86mm3okGmh+1nqAsiYD7Z+C+5t+r99Dqy8FPHYs7VpOllkp1J27ud
eszpBFQ2jq7LD+0+YNDfYl//ouU6XsbWE91wj+7ZqgNEiXa/R7GS9CPT2sqdsPgAh3MtdeayJUZh
ZxeYTKa+NVIfgxirabJA5532u5lDw9n9ADTBH4DBxXY41eMNhFrowOEr4MHaQsqWyBe4beqKsb5K
W/ptIaF6CgKyT7f67rzb/WpNugDNtStds/guSoKlNsmUkuuEN8alprrYRJrTpOW6fgSdR1NNe61m
p2fyx6CZNboEKmA3K+8VbtvuRPWhibERZez6heWcZLRpSTDkPNx+2G5Of+q2giz9JHkYuVarzkmN
wfgOI2nvBjNMmV/m6nPGhNM3mWX5Yh9WWnTTCORaqoS6mV4fbwrVrbN2X7jZI1ld5B/F25sJiF5R
s7pCYdkpfo48u8U4xJ6ZRu6920rB9JLDS2SlqzOOOcssC02K45AxJfnP5Lzddk1mo3IEvasM+4V4
GtIHD17G1Jo3FtsgVMOavSEJxznHtQ86+cLXGSpj3HNGKrxQFpIW9xZFoCMj0xkAhZDciLZiUhW4
f4+Yr3cUzNy6pbqj0ZbZ9fowk2Gj7ycq8bxIzwfyylJ2WNdI2+rjfm53ppkPi9zkUqNk0X3XM9Xb
thGw/d3cuzn1rGTP2tBCe7gyUWmMynvmXJijhOff55BkKE5s/lmgqEpKG29rgyCo5OFKDmj5cKo4
i6PUUnGyk/fXHNMcjCW4gTk0yNQjR6XEapTSvVMttLwpM+ITXsows4NY2YkXAQpP9eeNeFPGbQAd
0/pCxgDNrMHjZrjQskNoayLc0K4Bj0Kq9SeUebfBRoKS5Jboa4BMi7/Faf/YSapFSGyQl5bAgNVU
ycr7e+V+osol/M2fOktPYbgkiQdfOG0GVWWTO+PnNKi236N4IEzmgrVhL4kY1EqQcVa1AVLhuMkw
O7Tsyd8dlC3ZVEuVEBQLLgsQTs88zzq6C8LjoNhomOO2Sb6I1RvayROnEDg2ZOzhzy9DZs9BRPYP
FPChBBtARJ9BS/MOrEPmnCGAOctytiZXkqB7UXQFjt0dr81QZQ2hJlBDpZRn0ojciRD1fFMsIizv
lT6JkS0Mt75itExt7/rmUH7GlKZXgJV+8rVH/zYJ1BojSkLC70pXxnDMMpvqCbISSF+s8RJ5lIpZ
Ut4CZYLcjGB8Y7nUCQo5FzhfWR/u+U6TQSQPrU/U+yfQbGEdJfgtgXnSdXn/sW94XXKiQ1OeFObE
tZR66XOeS0BgXQZ+gV0eU2wwe+1gRlseMZfsoWjryHu7UfdfENGAlBly1TXzE8GY86et9Xc3s3nQ
fqLkfCOZsnztkWeDbzLS2FEFLb4I0BPJIdvY6kPTllQ4o0TjceZHeJXIQed0KZmjMC9xEfyTsAk5
PFUlhu/LhOh8/NfFYKhlYVLseU3xwYCbOTxqBQICCXvRkTU8ksvA/qxAISdrGY6cVajnJW4jOdq8
XandjhsGXdB4x5531w8i59gz/H+CsRiT+Kx+sd4PNHSAC9abKaGcb093fBOv2qW73yYT3zpCdEQJ
oJdGZ2i/ueDYCKB+3nQXB1TiayTJt8Nbd5HKde67nv9Xdk/ifTa/SPvtG3lo+GKjZZriRhx2Mdqp
1uJ0RsRKETjgWczLj/gsfFUJT/g9vlEzVdS0PemVyKzULaoa9aKPgjDDqLqtt30OwnEgxlcnW4Ke
1V36Is6VrHG2dG5OzdkzmFWx1k39UTEC2plhmf/XjjLg3ATrkb1i3JxbEF5Ned9Ev9sOOiQatuKC
mNK/ug0WdcWJJxLwD6us04qASn9RShHpnuGwO1sWGFtkvDV9llrf9Lhi2W+g9Apmeac2LePGR9sT
n3qmjb/WHQKXJcZewSjkZYLLMUv10/ioDVz5Ku1FUYXOfgo7mDDYFdQ9ti2JZ8jaMuLhuSuwuVng
3Uz7VRuG6LOFJchiqvlf/1IQbNov/YprtZL2y2gfWQqxknB1zrCFR+UC9PfGllfyTsNuDpeT5grY
XHc459nqYV3YBiy1jlGu3LUzQPAW/N1Ivds/IujUQywZ14ceL5ztJt93OXTFtITXT2cCfe9VvRTK
InQM62cJ7wo4+bme1Hd9orza7UfZu+YcM6Ia1cT6eGcfqwUE8z+6JvNcjlAklG4DBdzNGoGy75Cw
OhGtksSSHDuHtXuOYd3XtgOwziE8KsdcTDodG9E5BeHBE3Xys+cul38i3Pytz2VscQ5A2qcR+4su
WIQ0T+IGZPGwkhhaly+lLwu0QSVxmGdPjB0l+2QqEicsV+89eQKLqF3J6jadMvXM9T4AXLPckor5
qAQOg5FKV5/bRBe93zR+dXQTmZ1uJiVRufU9HczR7XTT1ezzNKc+mfXb4DW325DPdDYJn84QG6/0
otsiZ/2+DsjR0KTxL+Xg055zAVHQmqGA4U1u6yKjvS8ItWS8MjqTWQPnyEORrR4PE+d4/VwxxMXW
A/b0hgSo9/qSRcMaiEfZK9a7eUvhfyGiF/BYJmptDuHeHGZH0mbraXJoQKynH5xbJTS026XDChFO
aoZXGlll0rhhnWOkZnBjaefZRM4QibaEMGSPWIoKqca/5bbJ+qjl++wDHjbAYoCjSi9+wg/U5bR3
HEIWEppTgA6vjMicdyI9Kc2niVjhU5M6ucxvtTf3rV/A1/kS51Z15a64uLgL+oei3jNCBI7P+s/s
8MJwWgYdR+FwB4YO69rtJcPViXfrOcz9jhmpb06fLNbxgnL/78PI3zjzXBTSx97fieQrzd1wpx6c
W55CacwPRvbPVMDG1rCIE8A02FRJEX2FsOH5iyag2pexjR1p8cqwC4JGoolWaQExQEDe3TYFQE8R
YDxECPC0vsa9e2Vo0DcZ8rF/BA5QCT/R0AbA8QmrQ7qilJGSvrFl/aYleWARZtjRJNuEitFiOzO7
bKKeJhPSkXtwnxsaNZ0GPRwwtyX58TA/l36lxWq8rbkuHzSDX+HLNgBQxYYt/oTja1ooqgEgs9T/
ocTLUVvkqoNHyvAfmRRZsppmdiAkQvhnWiU3zJPpEMKnkldsAAkvRDgeUaEIcPc0hO35rRyJYn1U
R343pZFXYCbXkZ3jKvzaS1P2nDlju22hgOGXWTILBTTHqzw1pgQ1MiTcXi/LSSLRTV/fodKaBflB
rZYSdvc8g6W3M5J9NCiozmBlhtXVc0D4u3zvQnDdqaFufvEeWLp/UcRTVROQM6tXjrbC9exBz+tN
C2sIcemVAqNSspmuJlLaGDY02XgN773kmT0CMR735Os6A259JVepuQgfDQUgpXQVuIWIIFNDMhkw
Csf2ZTzzeciIYQ0u9doLfn3pC0LbwKptKgX0laFVunIhQCys7k6eH6M8o8ZLnom7SCub+rpUJ6ql
1QzvK5WOk1UkThzuLi1A6adx+QcxE9rGAZzrPAMLXNw2LwEuYkoDlYsE0EuXRbWZh4vI6HkdNPYw
qWPkEBjCc6BnNdJ92qmHI/UVuw6phvijMvrCghLls72hWE+pnt3JvW0PfaCLo9p03MoudsE+SNJV
efqu5/OvIeOiXU+RSJrMdxTLJCUYAWdcyvRZx0Evu6ZEzr9+VlZr3gUDBHGh373uryC7fx0AnIJV
cRm95ETbGJ/9+9+xf5xKky0/eoVuymQDaKo2+LapUlPDROeLOGjFjVgEE94wCtAcxxsQ4XGEYrOw
4uWWH6XjfoFtNzKEnjvULoBZt0NiaRNmPGq4LRW5G9Li8pQjJ0mgwbdpQr0JRX799NfblK9Kb0OK
JeYFUBw0wpAssF4vZBENnndhksdTmSdccyPKHhE3rs65l59nutv2qFuftp675/O+b9b0zBc+/Uds
GnG3+Dy0zqyPZxQq+aQ4xJHvJha/dkbm5+IKb6Y676F0uHOAIwPhKvkewZozqy2C+HNypkSBHMsI
0yXG8zjNR2qn6S0ApNKTNu4KlIA6TFOMMl40ph6/2AXQ3az2etW2A/GpCqghSbhRvOHbaK0ce4yC
C2Eqa4TH4c+iUj8qPvty1rSATGWoPK56ugB5dxK2xNJ0rIFzJX6CxJYALcejHy9LE5QH0xJPXIy4
dSxgpdtZq3OBbB3Hun7QNsz2DkxqfQaVU04zbiUhMswkAUqCUCf9Lrpd2M0psZyEGdOZMdgBwZdI
381X4MWZCMb6LqfZhmRcqv40fzgW5+rQS8cFn9VA2rEkMxvouLsqKW6PNxxkgRnUOYnPRVxKpf3e
HEDjg62LoMWt0hdwcxL3dYRUVYVALuD9T/R2yRykJnvZWp9S/sxKOaUCU3mjsKj/SHe3oc07DzzQ
ZVwqBNmbcwtR3nOOwhyU27L0vl5XO+EwktJuQ0KC6ZXzF6HHiur4eMHEmfHcBcdLmoeYdw43XsGY
OnQ6NjEH3Sdukz+0maTg9bcx6uS4EEyHgw64jS0/zmCDwgVZt8mHEpYv7VAXeSsAWYbaC2z8XLtV
/TOYydALuhYElLTx69WCXFsLKY8KGlITt936kZ+V9DPJixPwJjD1aRY6rifvg+W1IAiO3gYsTp9I
py0EwY6BFfxE7Pb3MMBDVq2iEJEm2/dEwF478V4+fgB4Jx4iuldgN0Dn+WRVyMwRx752CCtYHdbG
rrxkYMy2F22r91fO9ZxvSWSIAJOy8r77lBaQx8T84GCgVtFyLCWZt2uJOxALRUOVTOz8VaGXSGNi
XuwzeAnVoq6ctFsaulHxc5VgOk72i4TVAsnaECwdhlrkIlyxi4fSjFMqxxMGW2hB57UFvFGvwnOe
Oz1yJD+V760KirgsWIMxFVeMevOT/IBZnZfBdc3FHoKDRxcK0/HGBgTTFH/GOPelkcAwvxLJ+fKS
6LLHiQW5ar2ShIm+fnzcEN1La5XlBsjMRGFxQ2qoRHqhQmu0rRCXTVZDaQrYMqCCZsVwIhLE9FrT
YPwxy3YGRU9Z4VZNBIZxzubyGcDIwsLyj61Qoyy95xyglrO9VB4BrEQ1AahO4tNVYop0MNhe+vgt
q85yRXud9DUCSKmLN4cmzqRZ6He+qE2k3g8ZJCv2NMT3cI0lV/VhmChHUd/bw6/A6SWfMqzxFWwk
4wwNpoZKk3ulZmRr76oc6fVPF+qf5fh85nePJy/lSRYgsKKPu3Utwa60jgKyFK7G5gWgK/6sX4mD
d8P+XQ21QW4hBlGx8uSNXAxpVKpCVA85jNbQQDz0qnXjG0jZElDWaRoViVh0PhCmulfrP2m9bPYK
rgxXp7GWf4c56sOEoBSTgqIRkv1dQctLieOnjonjAro5AJ+lu8DMK5ro5emPI6tkpaQJcR9gdEZw
e15+Nzmi3PIQM9Qicz9OgJNQ3P1R42VEjQW8j809DoBeqTGepbcFyi/W3YRxgiIFUvFdmn6wmET2
X78o/fTYRVirYTGmHvsY/iDZ4vAS6eXjsiDCDnDrEbGkMkAy8Mi43Y2cWJ1CGP4d4VHM8kJe/M46
NtLzcMlfgJUQIPVYv2njEKRSzfK/KHsR8NR/H6fSrUKF6n5P45wo0vyi+Z60r76SAWKeYy3FF32u
qBn06UF+4y2SAGWB6jqljUnqYkJgbuyudipoK5ftbpATLlA7gPRh69zUO49UFHCg/ByPQv7gHwSS
363CFRuoi04z153YpzTs8n7H3JMyac4fUIl+EFXTjFU+mW6wOwcCC8POrFiVcuNwdWNDSyzH9+pR
wqBKqmGV9LSk9Ag9XgOrXE+qhgZUUrQlPjZSZTdI5Dxti3q0d4G6qHSrFYklhzjCIYVU2eqmCp23
qEAHhdRO3DwWu9m+j2HfTb+jM/XpQFPlFdJL2sBIV+pL0pQ6T8ztkMfXOveiwsrDa7rRKgrGfNbn
628oXzp+12SuAxc/yMyyxvd+Wli4ieYgb7FY0kwyfdGXUicDuxevPo1nFiCA9I688zyHHm80gYmd
7HY/9O/vFgTlLfjMNTrozmsrCoWQFBP7+GyMxvCv0fMwn9pq/nSZACa4rZjcdnzBBdY43jxXtnZx
hujaZajj6XlTFOh5keor4tDNuJJu5leXXEyOmPyPgHOCdf8wn/6VuyOnSTxXSIBuJVCtl6a3ktRt
/gpIt9JJci2AAroULR8c7DRGakoyRVXL6RAwslQSIOJ0ENGN1BvD5gPN0ca8lNWOHY9BpPEdwP4W
VO6sEEXHdAtWJW2Ocg1eLZE011PkFZTspvFjau7wsWnaYabGy72M+lLynaJDwSBcbDakLG/bNL9d
/RrmQlv7OXQSIfkxA/kAc3EOHa45EbCzlndu39exi+m+Qf/vZQ6koEB2n1ZiTM+5P+KKOygM7qb/
J6qqEr5PAg0KXuo+cFHQTj8S+IY2ofGwHJHXClwmfIK8abRkmwnNGLlM1LaW3txz0QOEq2fn6+td
kT1BGUrfC3NUHnjIM931rcH/ezbb+n1DF7+KuP6BoFRGqEXTSFTN2F1XZXf+xxA3NN95QiIV6zz/
oyvRZeszC8jKRXtc2t3m5eym+D6oqnuaHCtFrkPVLQuK7PNo57D6FdSjK7fBIMSSMIfWAjPWOCQ/
4rHeVcRu8RF+dTgeiNBS2+fu3DZRQAXVXtRSjPpCSHhGG6/iwwmyzS2oCR1cC+npJIDhZjf74XHx
2OlTnswegM9aZ92MwWo5maJvV97RhELpjkpHbZCyr4oKKCsIuXHkBvwlltjmo2FDjEi1ophJti+L
rbcJOL3CjBvtG2JlAg+CZJELL2+3koWOLlyTVL6bk+7FqhWejY8JsdiH49viIoZXrCKiuvTgeD1u
jjyZq54DfSPM8NOc4AYyGDkKeG9vywTyru10DTPbesFCRZOZWmkF/tDGv3HTka4+VIQq4iIJakX4
856ntT3QKzTz0GlPu8lsRxx0ZVGIlqvqri5xpmY8CTS7qRZBJyFrm98022UbK0L0zjXxQJznqTG6
f8kL42DqlhI3tIdxFHjX7ddbGM0r9lHsAt6O5AS/DxZqu0y0nG03+G7pmjZgnfrFE+oD0QD/d4dk
43om6cn7Yh0hQXvkDM4L6mbIlzU6uwzD9MGP9ZretZU3odjBjVi31j/eN75Vu1wDwGndwwiB4pSN
cUA6s2Y+ujWmlLwmxZz2qVOamVkynGu0d0SlxxQy5b/EU44Qv8SiszMYcmuzLjBes9GUSbQNRkKp
YfCntTruSPgbGNEVooaPXtAnngeIwfO62y6DytdSLD4bBecaF19beQPPIdVjXi/yQMPDvG3iv6op
12i127iduHp26v4I+IRSUiPUOQccDDpzHCkF89BrEAMlFZELTBqvUUnOupeAZ9s99vg+bRU5v3eZ
r83YnXth+C0RaK0cgtGozJNX1CLGCxBJoXZ2uK5S+tWxE9sVb3u0NuHe+rgnkYouaqO6+yEg4911
spRcqbxsaPmxJ/Xzk/Mn7I+HX7jxdqlFq59zlIG0KoCIDpoJpjbZ5WQdb8kxPNY1abP9N7pDr07D
WkVTq/Rm+Ocl4t1ys8bEgaNXLJMm/nfazzOAQsxrD/NMYf6ZYz+02WYc0IKtfPauPWTUva0subll
7sCfiSWKSzAX/R4Ef7wEfXrZU0cNRV56ea0rsqiqeTsvcapOx/ickI/b2wOJoz1eNxUK7gnKTO3m
ncfRgoh2niHbh1QODjrwVtU7yf6XHzryh1RRudAHClOYNTBvKuzGnEzwLmhGK0C3BQIZShnTf4cl
LspzMlIBxLJekmPloxsOkVKXsMIgKhBolJ7J334Dq+con4IC0FsRRbWhi/c1nooB92cf6c4nWnwx
33P/Ta7mF3nslg1hd19wSWuJwzKygnK9O1ttGb0y7fvhPla74rITjVIKk5nnU74Fpe2/nnK1DMES
2jRd01i1q9i6eZr8YXDUu9MiMRqjfw1ACAdbgVz4Y0v7JGNl7iG33CaYi1OfLkJnyqraYNuXqrbY
hVgpn4GMHG5etfTRLp8Ne5osUFAiB5T6KgCOfu72t4DbIak05gOUd9bLSZEnMGoCycVJ/MnqPiaX
AHsVM/3/rWoOZRWq41Dc63PbcVzdZGNptpHK3aEVFDdtMnJieCffAGKU1MOye7NJunC0wSWl2Jp9
U9w5Mw0hlDoofJ8VoS/88gkhgudKch9Irpygp34tjNChIbMxYnhm4mss5gU+eVG7c+636WTjPvAH
UUlUS6aUWdY2sPXzcF6WC6mCbURB9UwYU1G9z1jw6fuUznKCvbfEUigMqCBAtETc3d2Hapgr9+/F
3oKJdER30/VLig+bRO9OljinF29j7rxcex1T0IgXTqafGFZSFKnBYM68gSb/FcULSAKBQiPIOvxf
jjPvCMPEHIMt/zd9Hw853MEsgnGMT3nS0cT+lkeBl8NHGPbMfZCY64nCYMFIkjPjaNdrrFzLA3HY
vOi8CaU4GYmqiAHXvkT7AJ0BQcSG01Xu9cbqAmp4oIkzVXpK+Mm0YRA4Ih0QDSaHMBZepARmGEwD
bb6xgaQsbyb390rY3jKKOHyX+hUFFAuuJRHAzLJeG4hBuI669vfNSKWyK1OuXoMBH+7pjsgZPwWS
+F1FD1y42AoFRusr+g/OM8ej7FqGgvn5+bPFTDPV0sPQreIXKI9DEi5oW4F19iTPFGQVvuGfipLw
JtpSlZO42SzZDIWMJtZs+1awOjTObU36Kxm9npqZgk0e6C4bQYErK+7mlOmtaa8WpqsgEGc3QvBf
lPSS3l5ALPbM3mtyj/C4UgJQOFCxRTv0Bv9/7lJLw0HYsHSJ0pvTN2UOHTi4mnQB//27B0NBh4X8
Kj3wOOszYVJ6k34CmlNmErZ8NcSGJb78Ev56Eobuk12CUpZdTVQ+Y+ijbowEmDP+fC8fwoN5OeIe
LXfryR2jQAyvJstoRt0TAa5GG9UXkVjWqoYZareMI98/7r8mFdqSt5NhR4oPTtGZpyHUk0RGEIW1
7jyOfIz1jOCX+TCkcmfuXOyvg/9kvLWGWj67/dpj+CzlWwZRWCOMwGibChXtFU9aotswlCT3Hyer
TsVZcwd/xc1kJdEv5fZxOFgXwRhYpngj329Z5HYZZToB6qEJh1VIO4KnqpcNyLFFzzKjvXY2y09K
flb9tkvyypEzBTHebRKO9PawD0ZOdR0JEepWZh+LW5Zj4TK2mKh+Ax4yQG7nVLMOKthhP1I1z3dA
Pk9svTGYZPvvDGogcfmtg3vpuo2uCdKlnpwf08boDiy0Cio+q3IGgb1gCfjGt8DTK4/d09GodrrW
emrSbnwTsGvYezq0HGiAPAMWhCEKfj+kagjuGwcpIpOMQ2B2YU7vegj5a+fybYWNuezv56pLFEAP
vRIwMk0mWHnWVLOsgox6JvW+2uehbQ2HyiJAEwBvNWRUp6Sc/kVuu6I+szADdjg/Mb6YhQVVWpQV
4BLv1IqKcRkFXJevdRh6897HVkF+pd6ejcCMvpJ/39Id+cfQBppuvQd9UORSlXkw9NOcRqlqMLdv
x1WGK6qKufarvQBDMN/yxasMiwoCdx7GWxxLuLXz0YOpe+zX1+vrp9yu8QW8qaALEGrnzxXvShO7
baVvw6yGj7kEpbVeKM4EwDGG+SaSyva+Pyz2JstKba/adq+X+639wA7oa/LzrNM1xjnBFsLgd56P
bkkCNjdlZA9F+QQVG5URRjH9GZT6gDUvovBnu9yDZmG2c+8UsRsGuATgbDw7/LdYUmE/9GBBwxzv
fSgaH/q85LX/iwIFdtmFg+q1+5TkkS/BoQa5ocLtsRZkuFjbAEpkD1e+hjeTJAtlCaOuBr0gVeBa
EBo85vl66qLoT5Dbq6pp89ABl7E0F/3KjuKhMB/ITOdfBoG3iAeFbJbKdxPofxicjoEHvcuHxLv7
FntPN57QB/ZJ+sPWCDNotBnxdKYYwSjrq1I/5iqfEToJa0LYx8EoXo9Du7W7lDX5CwvM1ER63Ddw
vsusrqT7ROJb2mN9KqriUCCMF6ga8E3FMz94cb89mftfKA2UtmZGbYqkiqbaeDrLz+CGw30lh1HJ
ynyeI7ZJrQP1sKF+OjQsGf9R8T0XnZcc47dnykcoNPrm+nNWIAwn1pmaXkL5h+DHogXZJ+fVId8P
OOLG8ThQw3THHYEvL+9C7sUtP9WivWoi0ViZ28ddJ6FokHQ5fTGOj1pC4LzIJXOla3Aitbr4umCu
nrtaGDUk6rY+35V91NVIqcULZhKS5wjkgHKt9VUnJeMCjhRzGFMWVcj0dZwa4nSAFsmhQ04SaXYJ
qTqAd1unzTwjHdxQrKEtA4fLPrG3hgRWVxQOsHrBIo6wCI8ZXdxzZ8AjD66geqnnhZy47CTsDtvU
+BfcSPwa/J7TaEjfeyLOyc41Yujo6L0Nm62grkNFOp4mfk7vpPyFg+ClOmd0GH0D9/+yGAmqIiGm
f04K7uTfJkQ4lNxQfBxSbz910mDIkNTYuiMr9HLkbjPMdZbnPYN0lYSlY9uwQdut/2kgSo1vD8uu
KM32oXNXh1tAppdc5LR/NedZIzlATPmXUtZKmQm9HwcohSRIUCyAdmOk9lyWa7vPuBaxG2gSbDbu
ht8eYtZ5M+T5QX12O5k/oukcQjSYis6PMtmEDdsEZagxL6/Veo2a6Wbiwc1sd2LZwidtS6J0eu/0
HCmklfj9uovz11k+p6xKsPiM+sSZi8CMtDKMGODc2EoCHZIBM5WESvHdxFdB7aJmuDjEKQHTVAyO
w5eZInZF2yUaMQKgFhBP+VaKalhx7CmSpSNSyy460qyHtTCuFfe1ei9LhENWfaBYSg54hMSPv202
5C8xLee03BmqmEXkmkXu2mv6xrPa5n+KM/k/mRyAu5pGRnO0+gnIjPFxPnnoT7s1jwWQf05hUst0
pL5NgBgJLXak0zQa/MnwLA9JPY0gHWOn0hF1PeY7r3eEICAWgGVue3T5DGJkbRnKvNfS0DDKNTk+
afNddO5B/gTdtP7Wdij1FkOYZnOBxPNSzRGZvt7wvhqGsOqzPGO6M0VVri5rDxckQLsqObFUXQQ/
CLaZmMBJunJYz8JwWBVDLlDTDILm5WnhXo6vUVXko66gmDWApUGnrNBNcqQzYYawg5tWmoxEGDFJ
JZidmbAatu8mOgHmSOOxbChXIpqjPdoHpGyDb4nEW3laVr5ytiOjAT7S7ieQu+WbQ+EQXO2j8XP9
rBI4rVEExmweiXGNQni71KECmRQTiwqjBJLexli/yu3VX3desRBaBEU4yqdo1RthamGiG2llWyUd
t1k0DJm6SJGUiPzngQDQZmKusvXbYrifroFfzayQJ7nL3s5e353NK5WAxEC/cWl53jOeC4A7LFAj
kJNstKQruwGlnbYPRNEYaVs2eKmJ8Eotw6RMzHH8QGcd1JeX2wlJWgeeB8nmqaJebhPc8Ji3fLkA
097zzwI6yipzjQ5HY3/lMRh2m+S1/NZsytIEmb0ksB8N2ojDLPxkoZ0Izsa4C8ATt2CJBq6bajrt
miBB1e39/B8WZDL+chiAefdyy9vpxBciwFqOACGjiG54WlCdjkUjDtzYNokqRaNSMhTIH6pNvR0d
OVyWSMpP0Aeww/PZXfbXxoXm8dXPexBXz2tZodu9KILDej0Gr16A++16FTgiBCgEB7mhSICRaK1F
Y+IyiOzn74HG9PoStjkE0dsSazPHz/rz/hS0TjWPa4YFTJ/1c3w846StG3lNByCGrXCshUDKK4uI
/hmBp5HYx2pZq1vzNDyMVayRs3JdZj10mQ7IwCgCdvGyF8yuhoVF5zdd5LBPuez3FNpvfNmu+nqC
2TMgkc+U2B2mteEA0m4hLnAYDO1anN00/Ak+VNT0XRfVQeXVWEPNXufGJfUQve0Ce84YGIKnq7XF
aHJZiQgXupVhfCo1TQ7PQS7SynXW4xvJXY5rZvIQ702MBHevJ+pZyhjGLBCTvWhOIhJmH3DtpuQM
z5zWkDmJe0jyRpj+Atj0O4JSyQgfX/QB4lb9+H6WmjSoKc2lo0Qtjmg7vRWHCE483MFGe5i0dg/h
ZhQdh8o0mpMCvakRHl33SeTOVS4br/w5DvTQM8I5TWu4Zw0GIbBVwU5UXW5eD+1ZlAe3t26qnwB6
jZMq2lRCAZcfgI+1s9x/pQt9AhcfMb3mZStO4+6u3/clqCBlWMCcOaaEZosieY7dMwTH9QUiZ6+K
7qE2wLfoVDQ6NXHzsLecQvdAKwZ8aIyNM5uFMJn6p+mbpVYrtF/UFPAspghsZodobgfDBLUr3SyP
eo90aqrUEXPqrAqqdJhB6xPynhDIYWXQjiXXJtN47RU/N7fcSwzObIMb7IZjwZW2YScZ/rjPBraM
VewPG+fS/xfYb3cWOrzB9gqBkTjYff32quw+UmP3qHZSb31CSPWZA9h6HDiBDUaH7etcLKugy7uw
zbOUiU3VGl6oeP6UMZ0S4p4iUYJbMtph8zA+VXrn0EIxYHAnY8tmXZNpeDwRvDIcAu7TQsb6sOXr
otTWnP5BJLjzr0P+wP7wSmTlOk6LsvaKWHL+8o7MJoFvNaCFMvMeok800D6GaNHmKuPdfQRHiDJe
4qdJlMK6oOAhGaJ0QQQv5Yi+EFpzfSrcfdLtl5wQ4xMS1EboV/geM2Q/Oe/mEXPGPZ3mFJD5G/mk
Nibuv3iXmsesrZuDHtS+VEE4ALcUQ0mBPR0mx22tYCJHLykmtvCMl57H1el1eCaR6unY8JU0qcO9
FU8r0pG+Bonfh23IshsXOsnVvgJT/Ir+pqCT6OegHY1O/KPbPZInCVVWIStdHxFR9WIuSb15Zn2v
GhRX42zs1SroaVaIzU3Xh4Ul9E/hRx0p8FcJU7rsnevReT5h/yfQ+vzsY+0Mve+MyBn9uCu2aFz/
1lGZvUOWcMIhnODNE0c5xia0QIRYW3G12xJ2V6inde08AfUaZHmAN4Ca/AklPHV4CpvF8ybTaUsq
dZqZ2xKAgcvq+Oe0HdXxF/OOosU+rlIoa0R/G4O2fv+Tx2z5YjL6OUFgLjHu/mt0usIFSRqGtycZ
rDmrNmZeKlb/CQZsm7JlEDRF5WMNp5zJNQBjWYlugRMVHMp3SOfNXtflhQwgFhGtWsMN4mOP+kiE
gIariCtzPU/YKh9ORBcbdJCOxgUkvPXJ+2LmAf8qt5LRXzqUmWWNyLupuq+w6RXirDxfxj1zZBfq
dnKdgLIPxMugcvH17+z3aUFcXf0RqPHCk7/gJgj/9RWIYgR79iZBT9LoxYMCKRjyTx7pR+D9UiW6
NzlCwYUcqhZYn4pAJiNI24KgRFAvBwyuCpaB/viDolKGy0VARZ2YrRyCIORRA0zi/Acykb9L0B18
6L0Y8nKJNrkWZnRO/3B7ZWX12saW2FW/sCrH0Td0HMoGtS/lluMvU+mtnJYtg62VAdj2T0lPDNV+
dLzCyRvoZXcfu3PeOjzIhKv8QwUYnwNl+iG+TS36R7Gw/1k3TOyrCLYicehVgO8j4y/Dv0Yjlxw8
I73krxzHQos+8iVWU/WbCN/tCjrZ9PiUg33mZT3takNcf3zNmW4edzrlf+0upfWIAcxKaJJvzKrF
Tuz+xX/06XHLrJ5ZvX9KjVG8jG7jVCDUZbvq9pAX/XOpQmTw3G84hsKq9KEmkv5L04A1P6oJ1FIM
aaRv4ArgmzlLX3E/A3nIyC3QrJrUlXLTqqE4QPfzrLohXPW4TwmrL9eWMVKRXugykLmJMBbWSaeW
QTTj8hR3k2vYw5Sh/8GTIJDXVCaNONlKLsuNt4zHuBw31gXP1pAE4vNJ4NvBx5aw4LikM9w7UiLi
UT57XGbKXI2063g+9WDROWKr9mM17w/3cWiPqf+rpBaZzLCyWtysN6lO5xpJitdBr/+3TQpvYXvJ
45ogM7OZ9Rl3n1sz//GnV2AVfCLb0OzZ6OFkVAoi5trZkkzlNkE8gHU+A2JGb7nAsuruWQKNeHLq
3Ye0qoU3X0fBmxdfX57MXF1EPCJwtDfQ+R0Fsb3j33Tqvh0bpKIk/kz7wjAGreAN7SFX3maYu3cn
v/JEpPntpOvFthmPCzEWAmcBhxN0Js2opQPvp0TPektmUifFb3qi2GRe323NLcHMa2VwEZsxgAp1
m6111v0B9WEAP/CKVsyLV11qUOTh3Fp72ctVhqaQB/Be5NG2rGeOgEaqWmaqiKGSbycxwBp6LrUh
SjZMJwaBN7Cuu/B7zXTmxC89E7iof4l7NwMMmYA0VHJm8/cBehYgK6+fIpnoX3+BOKcUZq1OLgrw
ejbxTUFeJa6USiBtpeIKaT+OcjdkFCzU7xKIxin7fRVXuivuxXTuYYri33B2JkKU6uo8B5eQbPRb
KnxWs0ahwfeIcOQrt1b3g+QfRnB08z95lcYT6mVBSoAIm8JYSXy/mXZyw9JahU5XKOQGIxxHODDP
0wEXLq2g/dbva8+rW1deCvUBt4mHcU0EJU8brpgV30GyMLr8OXtoohOc8kD2j94PyGa5LqgHHgxg
Vxb47REIEG37UQ+7bCUV2OnKWMAYKnRA5q9626vjSVJMrVPOM5ekiddFSgZfUspiG/tUQSnClFlx
hTD81dC+0sTRS4rx7FK9Z6NI/bceidHQx8gRPjqVhZsj3AHWlW3y17o7TqxRknuwk0zEta9z+c8f
O505faJleqGAC80cjAWN+BsQ/fS39QWae5W4n0hic7/G4XOgF6gXSsop/nKPNfBYt0lTgjCKyFAZ
qGxZK2DI61YNIpo3bdEtXbWTaj1QK1PvrRDggOXqk9+6zADl5hM+BO/VRsB7U2LoQxqWK5cZZAMA
PRzCUm8Js7NKbQ+3KftZoswBhlNaBjfK0lEJnmYvzzaGlwJNYTldI3ynwhv62a+/PbdQ4VP0pajG
0semazcTxP5tqvgwLTF07zLLJL6qYkVhl0yz8R5BZQCef3D2ImrbwuJ0o/CXgt6q5971kB9f4ytz
eB0asgDYKT39kJJ05jjULTb6DQ9Du6Xk19aznZWLyuhldpkDXvr27DSBRJdkkDm4JtAmvwaqIw6V
bVccmc/dXh2Ui2Dh18uuKF433ZP7TXrpj70YuCyrOpRkNOK+j9b2/lJja4y1/mtEpktXTtb4r/NM
n/fNoZQfQAj7Yo+xoNdW1xLRCIaY8BArfdJNQKstmjCAcTezFlfOFcqoIs6V2xU/m+3M5T+yIGRO
0mTbFQAt+M65F7JEmbZiMxR9P/O8gxEdYbUw0oEqnWLULf2XL6TYmNcAbZZMMErN4Ya82nH5Nuc8
sWuj+xnsjPNlQto7P1GzhT83FNwBTvaJGUIRUuedehx1h4W3LH/qKpR1Y20zmHtZnaw+XRIh+ic2
mmKNjxQ790xt4qeMDhKkZ0dJK+83mDnBMzWfg2aGZOAwqSlx72UJtBHtGNN9kAwa7Jlwccx01EiW
8xPuA1Yr4fyrv8PjV17xBQcJZjv0Rkhn5bm8n8R/i5poHk9sPQRIUZW4BzdluUNd9eHwTE5rd3cm
rYSOoMgGIrZArh3A+MV0S9gFe5QvY8SI4eNk3VYLkT7uMchXe5h7/sl+NOqE9GePoNiDc+v3fgqd
sEU730EMv2li1TfddFSd5zvlZoxjOKuAwsIlOXudMjYRPEywmlJkHfp3Js+pCAxERXfQcp033s6i
gDgjHWgViwdR8nZZsbdOmJkVBaz8jPiD1Fz/7mEkTot069tkaSRbphYCK0xDRP8uEL2Sv+MQ5i7L
chiFJa6YP22+kQboU4YWIBNcK8NszEo9wFOcJgYfwwX1jcC/T2dLje5QznQskaPtQJpdR9NOz6OJ
q2HExbLb/VNSTIuj6Qg0TzLmza4Mi0CxRbttpkYvseLS/xStvxZIKIYCsNuEeiL+Gt74RWfnWcob
JhY4o69jcLbEgR66ZrEkL0YoEyAMHaEvj4XTa0m5KHzvBzYQKSAhBpVAIl7SE8GPDRAbQl4HhEQO
QouhHgMvTWMdlqv1UoGPEsx9b/1GP5yDb/tMi8YatxwpPJB9Ogeh4y/KwOaC4ner+CyMgvH+dsRQ
Wh07aLv1TlUjwD4wFJQF8NHCyvUVDAUa/aJyBEZceZlqF0wdKcUSYpc23d69ZWXbrUT7yNXzq4eM
eMKSWv/1L5zNDV8D6Kmge+YRoOM6ZA90EHe/fGMb+aPs4BPjO0QOtpFg70dgYuowZD0OcHivMddM
WIpyMrDi5/Vr7NcxrhRX3c9GXiKVO9W2vHV3mbnN+7zQNuRPolbUYhycjIk4V/kD+bgX/YhDoL0X
EvLN7YvbmETcwS/ShOJL9yF6rlJOxN0fU1qyw9B2PMofn55p0msiyz1DBfR1CjHGAHGYzQW4FP0r
DXciQtNuzjQr5yKRHLmOjrf8dh1XDWH/iroRFVZLrWcYP5nXFwAcOiz/3VZGojKSU27/Q6nyKZDC
HnIJGhC5tfmETqeC7dvfzYDiFWOlWbgGP6irQt/j8mJTK+w0zCBM78e2F6/7G2aXNkbMDyjsYryn
fZGsI9sqghvAaQx708NeAgigNziR8HAisXaoq4lPQ6MhWN8nUzMXoaN8Irw3aA6LI7+Le4N2oo7/
JJUwKAPO57daLFy4RpklKwN2s0aF8AEkDUi5VuiW3QnUQIVcic2WNmFWfc2xPQWz4ej4DGZU/Tpc
33hvPabm8SZZeQWFi3I/PFfdx09iaovo6Cmx5R22ucnDgqc16SQhV8EM8CVQULG6nNmc9oVbkAj/
QN3bPhXifB6WLcUfjus14aecytTjowYGZk8K1m5cGOWPJnuOtLjtko5Xc4mJTqG5BmEde+KYWt58
hOfSOlqedRcmnJanra7GmcmTcvyBkCp0JssWbp/ytcu/ehU7YdI8N4x9xl3npJVgRHU4jtwVs+o0
AQEFrpwO3nYckm/uzIXRyyDV43IZ3xSQGcBotdp17VjmekIX9SkhMUH+BUj+IoYDyyTKPtdVZzUZ
eaf7Lq29wK+re4BstFSoure9rTwDahoyVfrqzSbJ/9oEUuaVXKO1nmoqwEz1678CWyhyWvDLBBCz
x3C0gzVSYdau2JGfrnje2UBv6mgUFYioi55AhQTyrbXc72SzU7pFdIN4ygxBFR+wBSothzBthz8c
+9qYGL9z/ezOlguN8dg8E2i6GWuRBDteqbu18CLRMjUk/B/8Wz7O/6GZT7/1bB0vI28EWPIUNyW1
e54Asp7TavqDQ7PKM/mY0s509rVgc/OpknRVdJjahEHPmrV3er/jnPrphU8d7R14kqV8c017WQdR
5vpq79gWsqiYSsiKyIpkr9py+koIcDkEIrcydbiALKAMt1KIBX94LPoez2r79ADrt+iFtVNX6Vy0
Kr2LAcBbzY6CC1k8KJWlLUTqfMnn+PtnzS8bD3NnLrA52w0Tqs9FAPLhGJY+rb1huhTQVDqRKCFd
+fuQnxn7hp5Xaw6Jwr9SaWzwGUDBtb4IWSOzvPhT6FO8RZzM/Cqv1VxTG67whGBCZ5QhwvLqkCdw
/7OPk+zucRSQVWByetKIY4rA1xzaXU01HaTCZc5FVHaPScA9KhFNYjM2bz09P/1uheoCn9SBmQUJ
ssM5mXdFVAUTH2GzYPBmwiedCFn9HAwQJ9PkZdXdZhC0DyfUcwE3sjld8yMqDEKgbrSJIXTtdDt3
NRYsd4YZ/MofaQGQF7+2F/NNXfTBiNFdBvVQMs8Kxl0M7HYSShFMNKRCaEAozfze/Hah7Lg++/8q
zHOq+rJJ8v1bpBB6QHXw/Hn1sZzWogkDD4buXy9lEKwiVEzJ/UDwpXpR3PniLtgL9BNz9yYHCS5G
M6nqqM31XS+7n6g7g0RyhN2QD4umI4gZVQhG8cASbXZfNKfNWU6rtNzbEwDf4nhC9VOzIh7jIZ3J
ZuIllLvFwoIcfziJMafYlPhwuzkYoDJ9LyALTe7uCJ7O5IkNM2Zp6fDweH1NczlBN0DBtr1tg4EM
9Gry9LzDE2QedATiQfTXX+jjHOqPgjApQcKcoTGVIXgqu8AcYKhnMW975MBYmZ+rMGL4HcCl3ZuX
M3KpRH+O7V0s4hTFX+QAjgpsaR5dqRqohdwIvVghB+7vgktrbH6N3IJ+wI+jinqotSQAexJoLuRe
DUDp3YkzkoNMJGh/+SxF2htO9l94wSXGuAlOlcvegtkw4IlBgYmP0YMkq3EQPjrUGAPBvzMs/kr9
sT/VSBVMctxcXLrzNoc7DPyxvORhtH621ymPOy6vcBeti9CTICS7Weg+5TEgZ7hgbOoCu2LK6hwY
AtXZhMwF1G7EYPkg3boyttQtBrnlg64f+sRDmyDRC5VRpfJipvc80FaYpflHUMrwYNHZriBY8ggm
NLdhUrgJoVQ5KQvAL/xRjvNdt+QBR4lIkiNlRdSEOMyV3X6xvW+RkVFDD8Z4eGuOEUnyNDb4uoff
yhKrSNtc4Gy68i9V3ik+AZiL3bvh3WscZRH2kuAonsIO63UKDcjl2fGJXiAqYAfV5InTjjBjuE/1
7pBldaXMM9uMa9eI/4zp2dgKfz5qu5ytu46M1YWtlt2/HB4bXsY4Zggu6Kspygunli/qxwGS007B
4ZVXgDfd9eQ6dC0y1608WjXKuHMJxeVwbGhSwdJfRYMV3/n1G3/4kKL4jmYtHUcYn9L5j8aFFDH0
2DKTOX5kNvr//VQHiVDiX2mQhx5vDR/cIITLiA9aVEqEqyCx4EfGBypNuDomLcUhvtPA0NP7Z1vs
AEBTp12huCOzJmdX8o2+Gwj3jVDDVb1B0ZQzDV51WLAA/MkpvAhOr2i04SRCGxQYrwJqE23tKS/2
5631hX7SvjGrNzDGoH3SOFmQxW5+bQRpKduZmcq5MI8XOIwFhm5m3nNOWf5mX5rTkC08YakdMQbr
f48vyPTxnWyOF+J2JqMb4aI72Fq6kjtUfmW331MMw+HE5rx6rTzJWtju7JlIZQTBsdm4VIWnwE9P
+AzzQqlzry6CeDFsxT9XPDva8rXRe4ykOg34/oZIativzR32oaBZsmJ7HCx4cYoNRmLeLAY2mGya
iPQKe16qxkKkYVERjhmCzVMtck2MijW7TU9ersRQ8cYU3Uw4tJCOKJLznGmCqxkxDxtqj0Z9UnEc
8Y0t1bZcLuWzdOTqcWU7i1fTPm5vGPvzur+LPSltDuC17gzgoJQWMbsp8EjuYaKdsHycAg12WVEY
irwCSR5GKCFe+1e0rDTbcZTfewOxIU+9f5ZLLWT8AilOvxxQ8FpjVofXZj8O0oTLMucvpVhsmzby
yeKFWdeHZnAfPKTOYedVuJPurfParXI2JDNj6pFsgQ5I40ocAgXBqQjArWJzwwUa0IgXPYgLrfsD
Np3K1iuDLRq2tDVl2GTw6kbYKvJbpo0y6pRhe6KPPBmOM3/+NrqTjGPa8CY1jaU4PH5T7T2FhRoi
2uUXdUT1rSBK5O67ewqSOmO7L3FEx5V3Hzo7BwGiqmNRgckBiVBdk7uAfRse9A2yGK5i0UbITGxl
tzUCwP9NV0zbbgJi3n/egNXNH03Eqjz1IMZ40AQE6kWEV1LUvQNnc3HfgwT/N4NPIZVf1N5S9ybN
iHrdjgHPJnX4NRgDmeWFBh7Sw2G2XDL2H83qWMxDU/fO7+hsQ+trH8l70NN+2bETixyH1attzQ35
4kS1dBSzrivMLPF9OHsPO/nE+7ZOiqgalIvveDn2s2YvhaF/pI/KYhtAHCWm0WqehGowkfK1ndlL
5TCzv1ZZNXI7fDfiQ3CnYRiWUJRGO7aS9SuJ5rtjDwkV2YWMDHIMit7qtrblqveo9V+za/0lp2jv
APVsAE5YCM2IERjBeANMqYs68EIQFEzygRnLeUnTcPEFkNGlIwEU2YFZYsE0Gb2y4qxy0TiKDFVK
DQM8mlr8gXonCbP5+n8mXivkC1FrDelM3GWwJOzH4CtqlwtmMC+6jDcb4sVZ73oBTQVVPrrMmqti
zmS0kgVuRk8l+tQUfsJ6eLKTJUkl9r3MkjOj4p7xc2qwukXC6RxhFM/Sq65yJzUTYMHB1jw+3Gj7
SrbNYn0FMwrbIa7I+2MgiAtb/0TeLVxAmavv1AIKTABuWaL1PsbM0zVSBBT8DVmdcowc4ozpqWum
krTbiyrAG0BqmZhj+WMO5iOSJYloF7WjrdlV7eQR/gOcsobIgci9QDyaSqLEkjuce/ShVH4vr4qU
bPV0fA4ikpz0ArVfsC78xBwvBEwfUvRbvuA0t6G/jcxte9GjVOE208HR1K1pBo89bB7XAl0XAb01
yV91vztNefY/Uhm4c8Q3iK2omX2118ZIA09Lcr9BZRpOiukTNL17ozFmPhtfXoTN3dTlkMhOqWfw
4UH9VInt+MYvr/8FRR/U3fr+uQomUrhFprRtKd1UT+NdtQZb86xratxs5YH0e1ut5HhErFKfkP2k
P99DjBz5FP7N4sgBiRA6U07zQI9CPD62zvAJ9x1ZzpKxGjXC2hN5iGZbPj5APziJuQxV4Vr90ZCM
K4yvGYfGFBQna3h0awS8MwFYZ/tdZeIfAdF2NX/WFiv1TFfeqC7P0tCMqwV7y7FN/7vd9YjCF5yT
ZCLKUv9O+qeynmF4Rh0Q4Jye8Oc+Hl/EkuBvKL6shcn+pMFKFm2pbf+ja5f2qLEREBpPXje/wjwi
ufgz7rG6vB5s0Luccm5n/r8QuRRGJ4E6CXcYJjeCb73FBIgbkn8yj0hbevZYBuY8bVQbQDxaAa0K
xoM7HPGYPWn18/d1oxUVC5vR6YbLLdi4U7tB6XbcBtFzc9rqLKlv42tlO4X1crZ83lCiFioQy/J+
sd3oPJUDql5GG8Vkw6qCyqicGZ1zZSn7Pj143x0etf6a52bDBbXJgue+P2Xea4a/7C84trjjaWDn
8mS55fqX4URLl2M6ooIXvClZpS6PU+BreL69llKix5LYymWD8GPyRDtZD6aP26DzNTs5N9YfajDp
9fCR0WDWJFPivF3MNGCJ7DyLFOhx4YOmJk+fgcU6E4PZPyFXxTbu5v+vKM4zzNPEWdPxuLzWj2Oo
EitrLc+FA784jtTAaFPIddPIlfwMpaWWm9hqrOZM8n9fdXCij/frhc0AjuM7ofJ7hSaFpb4qmrRK
yza00SYJ2LCRuqoI6Kvw932gJnXvUwIR9zGpV/oEXrcOWBBtMvc4DRehZkshDs1+fiCwzU4KDpmB
Tz155NsM89kBH+mqUfHN/eVeNpw1HOkMuMfPInI7qwWVoUdDVw9sS3BXKB3Y8P5eLUvHjjxwnpH8
gSxd7eDRTHuDOym45iKbqzYe8K03khZawePmjUKq35nI27Og6BHE4hE45rLSL3k+tjATf1xBZbDM
c1DicDX+j9vMcPz0MKQ2mFwqOJtkVUl0mYcz5Jm9kEaIVu0M9x6GtxF5B2KXYkUMp7VM7tc5VN7O
mafY2KqTLRzyYYgdT5zjzu+YsmiYvGNvaBcxks52LLCtJOW+G5c+7/o1p9TWbXr9P8ApLYG/dJP3
NA5vLa9XahKzXhftKNHn1wAmd/r3JZy4Uveacq2bj5L+duX4G8etrEAZGrZVHqYzd5FNFsbmXIgt
ElXYkGCSlyEEHkAKsIbjpWFIjHme6TyMIMyzPrYRHXp4O1zyADi5HerFlohWhIH8ydM17jDWSR+F
w3ts34C3j8j1NZj76+kI/O+Sa78QN2QiVm7qqJKrp0r2q11QB4apj7GrXhObjDF94isdEzKqVvqa
1tAAmdVWA23YjSRH2Xa1Ij8B6+sv9LNt7YupRvoBVqs722hqamEXZC4DzZGGh+igH4yd5Nu+5m4z
Cn72+6hTwIcR0lwyHNevSnFFgswnASnbUKVzNYpNlkoOyHOW+ddSh66IfBL7Ti6B9NoZ3vWQjwhd
BViUY+DWhyXFZtIz173xmiGL8juO+JrolL2DqTzToTlSsFHXZ+9bBQCt2CuVqdhT7+zi/+ahKI/R
n+kH+M5k9YOvmK25rmCtzruNUAeaOrFUlXLRwHr2A22ARHc5w7AO+9MPuSR8m2jo0QoFQmwymGnd
jk0X0LteA49/GmeKJf7RGWkIF7U2O1cDldfTUM5OAtf1rkWJtzpuP6Gl+Dl4w+wwxUD7TlGo8ZOx
5Rf5fQ4zFeJb5uwHmSg24vklRVZvOW5Rqg1CUkR4Eibu/jOvxudAZ6L9q2IKZWXt5BTv+hMk9utf
OWgqtHaJveH/sxBVm8TCNeKZUg22NuB/W5HIZbFBQR++R/FVfchEwjfat1gKjgbfvfp7bN3BqhtB
b2uUsTdgpcuuGj01CqxqnWFscYEBhpt8ReVTXp5g4Vcl6D/0ku+AkFWWzKDuS7rZM+h2XSnI+i6K
asAs7sRbqnamG1gicWev989clLCdehkEq2VM4Jsx+4OocqqmihoUzAkdSMflZY10/8NE7oCiIWqb
Gsh2HwRMcfpD2TRsieqGmeZFXDZddChvHae6150UD+ccNbjmTUo4YrjNvr5IhsBKAbkN5D3APxgC
znVcdxI9pLP8pRBPpR469d48kN0iiXD8/3+U+slzDdv5SqZyiSBq3bB667aEP9Z9kOqshdYPT4EF
S778I+EksVFxTnMALgiqL4rbL4PFw6HGwLiSyD0SyB5B66RFL4yEwoX+d1le/iMieaDfmrGB/Pbz
oCnNaMaYn1itQbE9FaIfZje5zGsaIIEraEQ0KJYFLJQs9ClF8dvKU27GVCVlmFwXJaomtfnkbIcE
S+cgLRKPcKirY6rFV8cAwqB8mQp5YFpUIs2FoiW+fGTQZGpf5VtpmehKRvas6JR+Co7fapXrBTEh
fHvpp0blOtTPRxhC+fLyF8sh1S22gcy20aNE5Nuot0nfgGOMpr9wdJfI2kKQatscGvc2F0uefnv+
R7hD7c3nGyALO7WyT9w11bK1HYVUl4jrUVH/W/V9MAPSaKXF3/Ggz9GNl40HhmaAEY6p1gsaeEY+
4slSuRK21Fw57r9sDFDf/OH6SU579Ziqos5HPM8oi6fkwlLbW5IIDBM7VKJPJj3DzRfjFwkF75PH
x2aODvZlP/YSAxzCu14dL/LIXr2eMT9pwVS+aMF/vlGQDbpKV1bldvnCUan+SAyOLPJigWVJRgw2
YwIpYMvIQnfEq+7QaBx8ArEWiMCYqMHY4HShK/UXbhTE8GfWSake1w/IwinpnCu/db1h4YamDSdn
or86FneMtaU6NJfdQ3UC7tWBRCPDnIfDgryMZk6FxM0e28/xbSKCeNVn7hROjXpmoBuHBPfUOVEH
dHJDd6363EWRUoF2Mf4nuXe7VNLmnoa+QBoxRO09w1+SeR9fbG0iLa4TOQkkbUnbhfUiIyQEyIZW
9GW9HBPS/PfqmD8abayz5ILCSyWS/vtrW0eHvSV6pJvOJkFBUcO1dDwsAvJTIhb6/hTQxW9bmZOL
BOYa0SRmT1O+wD3lq7Pxct5SefcngKjrvNx0mhV7vYSPWGaX71a7Q2lVthypvHr097zU2JaeJrRg
3HdyHx3MM9xkblzgZFevCb9WVNOki4ycywO+PV4S+IwmGmPorwEoAigEKjg7gW8XHkYgLJRQ88V5
YOaohN4ig1YOPymaOD71H3B8pJyCd0tXeYwDyyjs4K6/lOdNqZlOanbPiWqBQCT0PmueqRqKEB5/
CLRNV4oRtcRlkBwspZm1/cz+B+tUV4DbOb9Ym29/eLbhLSo4uSHkOMqHaeCWTcNVPvDj9Pgh1OVq
bp1LOWbIuACI/Rp5/W2eCh2fnZ2t5GrwMS2gGR1lpmXbfzoJ3RtsXNbzM0LhdBaXxf6nyzmkVcc0
XN8FNmI4scFRBnC5KrGmcY+N9pYh1mFU1z1nziCoG7CrKH/YugJgEvJZKePGvRhX26b/ceHzyygn
3LT4RVbwLxOiixn9/edZ+8VZxRsXIaRmGGklxPec9ttu9TqzhWhOq/b2pfnnxDNf0iCLHYbO6+Wb
PcyDkFKUIxn0MrRf4MPcLMDaXhWq39CgKzMLtbuh2lrLNPU0ieSnKmmLxqa/1Fy5v/1AMCs44yfH
1aIMY9FX401eZGsjEoLxXh422beTuEL+iM/z+HVNzhZkz5fJTOGcLsvpZqmkWItmwL/z9+xpWllo
KZe8dJtd2SHtcj9daJK1QZO8/fXEVWG7GdNeijJ/3v+pRmtdFF7zrK8z7fPluCbjbgTCmDjw3DjL
H2uVHXK/t+LbKh7hZgHxvinMXdzrAe56rkFDikBdRRBB4Pdt5XqyugwaS35yKDlUz63G7qS34Zds
SZqnWOfl1HTSRWoaRE4q/wh4/yrVSvt1AGqVW/qaxy37dcApAfkKOULsWnoDTP2ZlKBjJuktNX2J
XFINSQS3nHjX45VR8W3GOmH8fAwJ/Hg/M9CZhczXYZQTH4WULi3ubaZa/J4r+EM91R5OSdQ8V4+5
/kwVuSepkSh+rp11YH8/3uiybQUlyTFBy8ijCASAvxkcgy/8IP9a0LBzWqgp/LUEZ1xcDnoPp/p9
/2U5iIuGF2im+J5n+m2nUxTHLfc5Be685JXBthlCJP8p4Ff2i8s1i4QW/NUigAYn/xRb0K99Yo+f
W/luBzO2Tg45FBBaisS0jlh+Gvas5ruHqkHdWi+hmb3cySclOR0VFakHFrZehOlpriMPdUHq/v78
ahOvNt7/zRQHxEoz7HEoUd4eW4l2bpB87nSTEgzhJzivNoiOjqoC/WJZuNjIqi4ngzRAwH1L+JYS
CjS1JqlIO9CBX7ZReCZLFe3+MXvpXjLCCs+Gk+PPWFKnTEbVbbVjXJYPtNsIUdL0jr6HlL1lmbkj
AJOYI2MpGcT00SrfY2b7XRwmWOFkjIwKX6h/JiugufBQxq5ZRx61m7i2yLAhfwSYPhF2GICulotF
1ZzF/VhHzTVO9Po2Gy2ryCAWTofwfCiwJIXNtppCguRPTWtJ+fk505gMk+m2Lb9/KBjge9cM7N8z
RY1TtW9fW8gqeBMbTpH/wKYHns1iaNkTjFEPYwNxFIU8Wm0AOojjNic5dh9XznWLGHaAnboKjBz1
yl0Q8DbmnZu1EGsyQrkyhKwmhHZGVo/hT0OcZGXAmkon/Gtk4clGfVb1sdyAmvwNmrb4mH9bQRa/
55TzeYptR5j30327K68sqUr31k3i2M1ZV3EqGA4nzwXG7UFouov26TK5//2btvGg28+Z56jnGdLG
6lAggJ4LxDbOuxEIn9dzmxA0ICGAESzAYGg+/mXthHHAYCngfwIgDKv0RZ8AN6spE4pdWVws3hN6
kYlZksnJJhTH93SWoFxELh/Mrh/B6CVa+q+7CecjLMYrEmtwQg9aHGd8wn0X7A3/p1iCXlz+I3CH
+6YZCAogrf88mAlAo+gg0It2s23Q8BrJ5bpXDyaNatIXn7+3qekzbvYSFHGYIBbzNvBSvD4PSUV6
EO1bV0S9kamDKr9NbXh7SAkFhJ41HDd8/XjLXW+rDtMH9ONAuNarKmY4WsSJmOPcECz8qy6p5D0O
4s6V5WZ5RthAMmPl+yAV1QgWdYUSSfDoQ2hhJiOiAUOLtj98BklEzNGJD2zYilcgHxwXqjOTzKot
wsB70oM+Rw+y3CKp0b4JQV1WsGeNY82iExHFFoRoxO4vQjI1pyMOInmfvsJTIHje5zunoEfGWib9
SVl5sdLn3pfxS85TITDkSwtHvK4xogHGkjUJtcQMHjObotOxytF1UdkrUIDD7I5X9RGKzor3Kuq4
UVJONxjNrKhveLvXSYZdpbgzIGj1gCl4F5xVaV3Mjp4fgfmTaj9hE0IfMncHGawUpMtfTH3EYqlz
gWtfrKm8deNEPYKZvYhPm7wKFM8h2FETbWRlWAhQlUR7iDSFmYDabV7BjaeO2bSaCv2xaQe/ckej
QTy9riuxFwDjRDfqhTz0GGKMKVIdyBje9XIyzAYlztL5oplH7UFrCAd5SJnpjusWUzTASCS9QZtj
eALnSxeuPq7gwPN4h5Vkqh9id9Tt+jd98X19uJ2W2z62RxY5d+ms1y4Umu2MQU9ESOfQbfVAb76B
ASv+U6jaJ6z3Z8p7A+bFP4qnyRorTutLeiTLL7cyDaHSziZFDjCRWfyl2b7Bd07H4rLiPesnecjc
40fPwt7F3pj7pe/ahD+wHceBrUXtet+HpngikhRI7dxajc6C240cPMH1FuyTvtHP1hfuUD3d93iD
O4pW+fHvo5dgxtvysOXWIlzAuv6uAKDC8X2LGhvrmvCiBhegSBeutfL5/wms5pjqup0+XwbzECYV
ZrIyHZ2UssDNahnV9aslA9mZ+aMaDVAPiPKh1aTv09Ero3lvDd6HDCWJMKtQm7MSEv2vYHxoyb8A
sb0+U/zlQov++c36m1x2AeTRrx5xV+4gH95MQdVDMJiugX8d9cH9XJQRPZnBDHyNRnyTOHZSXflP
MFmwFZ9EV3sNqymQ8LCu78c2j6wIy1ij2iiGe0bogRKMu/iFSloS95qw/tIepCRBy7BwWtm9oL1P
50ZbCbU+G7yOp2KaeHazR+8xxFTvEBqpnKLETPcCj1y1Zbgz0XajijLD8Er7YKvvFb03aVVwxQM1
283hvfOw3+8w6Pe1IDoVc0W3Gs2KLGKsyiS0+XvKvhKDPf8t+I4R8Rlg+s/N1nE13lMQsZxnMljo
CzRG/1if8PmpiJO4K1S53EE7DEo0redbuLKiemSZvBEeRIyeDDJaSHsPK+TxJNnQQG3vfvvMafJR
+mTzvNMkNP1/Lybh9VbUkGuiNOfp92sMd3BIGSENvyXtHWyWTjoo5oBfm7HnmR4za8wv/kvcID8L
bLtIcengTXKT8XC9c8gp+jCUW6QhPi31p7+9fPDIODLovuVVsHb0RkDn1Z9IHwQ8isUBQFc9Z49v
zqMhKIhNJewRbQK26RkWQfQkxuVm2sBV8LaJqhR48Ulb/8oESgC73sqxqG/Rnjhar0xDjaync12j
UpxidymaGOib5ktOulRA7OMLOjyZarOP1tgtMaBf5FIIpv5aj6+zKxE4lrCWVjYZpcd9DYrj9FTg
p3t5Y9ENYQWowBCIlrAKO4L0jez4WkV90QFKVdbnffYbUTCRGC3n1YUeibUBvOm+FAwPLco3Zfjc
KI6qfseKwm+fAtGI6yGFRlL43xJtz5efp4kxGv1jMBOfUBHna7ekcNlPBvDjq6VbOB2lxcx8Bdpw
LWGmXEDQyKrIZhjQmjK6P3ABccC5cix47iyQXeYISd8avreuCG+W3e6/s3/E8wFQApEXNzRu8eqd
40PZXo0x9cSup1dn584cKNuONFs6XIYpM0ZHof25KJQxiYI2payvjjaMRODyST81gWgHGXt8WaDf
NX9rLqavYM9cGIDGheh0jk8opoS67bWGvDI9Db/BrCrfuyyQql4iI07zCOo+Bh15lnRvBEplimMX
tw9XYFsHb6EIMF9b8J9Nh3fJ/p1Fd6gd62WBbUw6zl+rGV5c76Zr0+ALa7RLcXK+XKrQf98DQsPQ
e8UZ2m5leuWX11iQRrNPotZMY/NrVj6fQqD8ccHZ5R5D9cF7GnyKjnmKBYh+/nXd9hn+XPPHe2AJ
PuI8PbojhB3krJCr30HgC+SEegg1mymV0VZMXC4KwHEmZAuthP+rJrCqTzlo9OqKUurV6kMeZ/kG
m3Xs2rbh+TdnMFoFHAuLYuwPiLLZ3Dn0EPbkOtd4qAsYL4bQ7IVcaBzebobjAnoP0PC6JN+gK4t7
9HDxcxRk8cL3YUs99xLn+Bya/j2O7AkkCwm/K15NP1OMU76hDZYq+8KpGu29K/PZR+JzlzqIZcpp
AXYsdxqDSz7vvuiliRbaB5nNOojUeg+P9x59wOjOtJzpNeHRlhYFrVZZExKJS7LZh6k8L9e8M0c8
t6D1CWt2i/KcoioCMOK/Kkb//+Y1j8kkNCzLGTME2H07k40I9WfGUa/H3PvByk/9uDJwsBOs9eox
zYRXS9gKp5gUlDBZX+iRfV3mtESPzKBzFBoqkFxyStDMpCORHVOjPLunp3SFILWdUTzNaEwo6k7s
kEAMl75yzKRFesY7e2qKItIXbNmkEGy8ANbKjs8eeMWbv1ryCj0XTncihlxntGyjsPIKTLktuC2R
7n3rMuRkki5UcGaJBFoBsmWowBrtqYs+nZYegUoeuk1UtVg+9Ar6JANlbSMDxdRMXy0WjXQCPheN
Q6tymI3oDuuZWAeuapMnAAEsbLxwGAoXzh4RQMZDqq1gpA9v8xTJMHgDGDBxn8mKcL+n9/lw2DQw
/G/V88r9ftlo6xXvLQW6KT3ju4KpQycX22y2cNlrPiicmNiQM5aMQUmuYNnVtCfcxo55dZLiWXbo
teQZrc9zxRNV8kfL2HYuU6Jo401dEdC+Q7BzaUohZ/Z8+3q0le8Jgt3C9ymV/3a3DG1FCqiIp/bq
8IygW+IiVWpxSDGC1p6Z3o739khaCO1kTAVL9LNvtnZS44lA2h9OlT3eX8TaPiH6L6klXutGoBDz
IFNlTloZ7S26c+mxFxCd8A9Xi7F997kXCRMazk4JBrMKL4sFnnF52PFDtCcQ0bSrLKvjAPbfZH1d
PxBXpvv1snMzL4ClRKYArOLvDm38MNbX8u6iPtPh8Um+K9QRs85nIuS41VS0os8kOPAMaqeg4/ho
UQ9K4bfG3+xAf+QZiy2SF2MipVGMWvOOluQkUBFUZHcd9+rFKn6Ph83LzvTh7PougKG5nfUL6XAp
vhngzr5rUpLLMqeWG7OH882yVT06/Qdj504xcD0InTVVJkdEySNGpu4t4wJxZrGAVh12MyXRXJ2N
F3YGc5Zn+yKmsDMvmI7k9nPlQgnrWAu6GhCwFM479Cr1a+LD4ZJZrtO0wxf5DC3ADUSCMvmQrMWM
KRLCc5pwImqlYsoW/9rR1InrV5Dx9FSMaHAoXiyUHjzVpwuIDhjziHMVdxRHuYaZLKe8jZLlaC4i
yVS1URRvds5hDxNE6RIXtJBcEQPR7qOe4GdZiBqVg9MfF4ruaOp7iF4EiohTEh9oUtSb3tZq10E/
Z3FmzGLYxKiaHemScgHeVlWeB771WuxaclYFWu33eGpdX2qpY5YRZOUjG4Ny0HoAj0iL36i4Rugm
+mSl9LQuxBdE6kFw8gC3nw2MdZvJEruC+R8uoJ+4LJm9qcCjCtMtaGJOLZw+ycQ15qTJyaa+17Tg
LNpLZYsnkLK8CNKYcw1DQtYTc+zpV7aaqI3FTDHGRP/DqqZIpeN/e4ZtXiWSfja2NWafHfOl9VLv
WEnMQTg2G9oS2aulfXZ7lA8x4miB/yiG9JvFdqQqoXP72oYXIFcQkpEINNkt88EJfO/N2TAcwXWw
WNon7rxMA/75c7AZ1ZOXFVLny327EtqDRsZEM1pktxHrPt7SU5OJFJJhXdsCDjZ+n8EKM736rAab
Nf2hPoU1z2e/bJEKeyilMN5JBhXckgHXNkdp/k3ZtUTkcXRe9rWjrTC9Nr9r9nE4rrRcx+HSwtCa
PuiHcSZdffTg50S/seQOM2KTQv6QOuJO4CtzPJewkZBFCvs0J2IyxcyXbb0M/ZHqh0/gKKJm4dHK
Olg1VOaQPzEzFxBxn3JI/CQyIKyuTy8NJKsQvQM6bY4HDYNnAE0Yo607W/RbxbSLE30OzKR+QiTD
QI+vBwfDOnvYw2+WhfMOhgZncgpMtWz3ZF9sWck/jNjOKnt4gJvrIy/LTFf90Hejg+lMhsaAyQp9
8sXQWsVrJud0Okp+LtuG3os/1tezTuF6Zdr2Zx5xnBnLcDkTEFwdDT/OynH/yALq6sUqQOkpMEV0
90KY6camiq5nSj3Ba9XXKsqVQhNdXs95UtSkpZ6cM4dvXNUi5Fna4J2Vc5OZ9aGyx9UBHXRovpoW
Kv9qtUpVRGQ0nBKmj12hmuYDhBrOXCIdSfs6pa77hstlr+kKE/R+wZP+7/X27wbxL44+jN8GWU+G
AwKnukmZTRCh9T0+3ZAmPz1uBxTvcb4o4tgHLgPC/4atuumF1c0Z7YZMU+sxf9jNBrLRXqsu8qN1
m9e1K1M8f7UwFJiBhfGnQ1TSyV4TM7JtvPD7U8kltANe8yoJ+XyKC/vutAS/LDzF7i/3YynwAjWZ
TPwvHOo4mo5QKjoDGa2IZo3Y9egjQk6dnxnANR/SOCxOc6nqTcSgAhHKeoXbWBNCRvsOnKrIWoHo
ntOelJpHIaSohB/3Id9CU6n2oxZSq6PQHoXbI3Tp+IGk3TEHVlVVZRzShX4kDuJ7uR0YoYS9fZOd
6U02NHkx2XQgyOvRqD4bdH1jCoT7WfeD3fa2sVzljvhjzvTEXy9nu77FnbQHHYuRYrpchZwAzKdt
jYhU0Wr86l1VXhjdV1jJYEg58lCgLIMBjaWGsUGc9k4w4tFmsoA/QeYW+KLUDOxFHtEXBIXTMiyW
WY96gRpgbEtLGd7HcxX37EHrWppcJ0kGYhjBOHE/7SkIRcwJOmOaBq8kitw9R2CvOrJsND9Mcl4E
A9AwY9xroO0Owl/ry0HiYjMdQDwG+ybh2NDsWB90Hd53vft0OF9OweJcPdQwyYY8sCwRaM/fpidJ
lumepyyiriHL+qBOzMZInQXXMN+vr5mdJy9cXAw+AdkBkuCwU8t2AUipBL9uWWhlZxui4UIQ/mNT
S2E8bfdXsP9+ZnTixYpEJMkrc2p6/EsFrnGUGbJ4mc8aNMP3AKZCRXX4NLMloWk7NFh915zkTeze
fL9v+dV27wPiPhEKRgZvhOzo7bB9KIBStiE7d8R9DRhlQeElfYFoBo5Upn9hxRU7nMck7r5iuncc
lR20piioz+U9Y4ctJOOlRSayoENjtnwUxU3wupkRvvnli0aLYWZl6tQgUUrn5vlL7b+DL7A0AqhD
BFByUdh/tKqVis4VwDobmLTEUcdYs2rpkKCaWXE19E++XBpw8H2N97731IR2+1fXN1c+4TdQB1NR
vsHvVyuAVnpNlfNWO4+r8zWm+OxMVtiOfBKAzeUuj7xy7LKAGDVrjjboMUac6cVHmsVzO6ZundPK
4ALR4xD7sWcWJzozIfjWLmTlUn5JF7TBs2sxs6bg1dljqn+ImOSiU5aij+6WUp89sCPRNWXFaqkd
c8kgTScPiS53oyHm6W85z5p4bDmvIfeHN8CBRa7U09NSqIKLjz8X8B8WwCmMy7O6+P7f24HWEbJO
8D7wr8ONdJqr0X30Md/hj6B6iX6ev/n+NprNiu4kQlVIghPSm31oXe45kKIVqjCLMa/IM4WaIgGn
bonN1MraGGEXMqGxN1wdz3/4SoQihWjh+iRsNhfp0LDkyHV2oHLQnsChnaVy8gZLbJiJ8NfgLDBc
g6K9J4NznrbSgCM2Y7tfDNghd9NbvzYAne3M+0VgKSJA+uE+D/wLy61bCDktjOYrv9IJeCGYsH7q
Upy8QveH12ho2Vz89ye2FkKXTopORSGMwMPAyCRRfcvmMO/hR6RfBIxWVKChEHCeXSzK/CkR1Ifz
Hl9T4NKE6ndTEWWvHIBsnNseihV9wlmh3molLg5v6/7HpWRUz2PztJGd6ug3ohMbdyNJd8OIVjQ1
TNx0u8Hq7Z2dMnNWPRctKcdQ0MERjNv6ebYOwDVry/egi3h0xaFxdDRw51I1a+3jeT/MO+K8XJRV
7AnddiQ+OVvi1H0uaH5bLkNVwdb8dUpTJvYbjslONPS3KRH0LGFZrMbndF321MJsIIqDCElGAvUG
N+HNaYBq8/coUcR5acKk5gKYb6T3mJd5tLSETRINI099uRekp0bkuliDxcBGfwwHq4PVb/uyu4bj
EPiqsoK6JB1o5ygDen34zZMhGHh4ZJs4KH7awUV7eHRQluMtKtdsFx8KBNW+uZooLKrbktVWbUF6
lMzMBMPpv6byZJD3rJS6cqwrewR3jDG4Bl4Oyr6F5xbywJZG/g51QCVdTQTbVyBBS4WuNmXBOuni
dKc8+gEQ7y3GLbaKub2FlE0pq3FmznrJhLRn+jdMeLR41tf7Yjo3sJqxGYFCOSZaTZEaefjhi0Xt
IiHbhst/XL16fyxo+fhBz7NjaIfi9aSpILTWpBTosz1qGOqljz6ju/OYggV0asz7QqEk79339XZx
j5VAr1n57ttvXj+PYCIfL4sdlU6NXCWO7Zk9dpGCzlLCaHQJVSziUCzznTzVz7KooNJyFT7TIJ+v
B7LjKuLpsWXQPD5LgjPdPr/tMJspzjEYpBuq8y2TsSdBpYXkyCQ9wEnBER5DSWgPe2sFqt5hcKkW
5ua7DHOuJxqvM+NU3Nz9LN5EHIXFHvXebt04eYvqylLW6tHe3Og0AG2nuEjAAEcQoDixJcYATt2a
7xj8KjXMayhfsitm5cQ6jOX3lv9laowG6mgOSVLTMjyxjaQ0Tw8qIIeCFibiFukU2QeTHJUScDU3
4r6Lt9foSUnmgc9AAO2FewLChRfyGsGmeQhwd2n+KWRF7zt7WYrBnSXH7417aVYgZvRSk88xG781
EL1rGx0RGyyKdSQnVKh/N5i8APmunuRtIhzV5G1nzuu6YbgvfQ7iBtrr0tpAuPU+mWNXEDtJ/iwi
P0NnNBSM6kMHs6Li4LwTO6134jKYH9V/vdN4VvyicpF4iS/PPr6q6vfkCkT8vy6YauocDmOj4eEC
1Q9hymJ3V/ubBMT6LfKJRlsXfsqLyjAH7IfMiVd+emTWHPoqmSB943R2bv2oyPaK3p13bJsK/ng7
orXFd3ETI2DQBpdDK+3U/p4i5l1Jfk2Aa02f7qE3TZrjasBCcYOECUpGMfdAsYgozAIiDddtDD1s
tnGxk6eyRYk/p28Ckf+pL9t6AAAIEPS5i1v9QhSp2CUObhFSchYtSAiF5uJsIeSuigLFW9D0N4hF
vCxGrBB5N09ihi7dybUc7sC0jzoD9/eWlXNVfW1cX1ayuOB3reiPAwGcwVCTxVQ6PDCuw1GZvsyi
7AUGQtQfiapZaOwq8B4etsWX/39h8/lxacsRoJzKxBD31kRgUSQfgcu5tezaE/WyvcuTuoRqbkdT
s1hVehsZSqWnszB0V6l9saBVwN01EZZugKYKspZDasIStNqRAZDDD1mklgDSOmPhYd7GfQrqgF19
vAYiPpQW7A2WfcqnLEN0wZEQV0GWI328ALghMjId0MeFEzvqax3KQIYG3891w/IoO17weTKE/C/U
bBWCytlE8OEf2axIle0atoPNRRgpq4vO3ILpFd0cydVlRWM1kJEogj6EvXTsx2vtPTneGjXykz+Z
tpfrtSfxrybMkvzNLl/K1WQMjX0hC4uH/1KETzAXhIA2rxQrqxLgx+tlYnIidSaEUMlLY8J+RMzs
FBNeuvBZ4Ytv73ZvE7MQZkB1UJJ4mCQzs3CyJfzrt/Tgl0Ps1QA087ZpuI1erhB7P7ZeHW+2la8X
5Z9MEivkeNSO/T5wK2xKotWhqknvBzZhPQPCIihHwzed6KDOqmXd/1WWCQs9dAKkQ5dhkNLHCn+L
npdMYSog8MjNcxLpCPho+RP8idXwz667GB3Y8iYcyNPP/aYWHy3Bx/NIupDOvth36FgdOes9kY4x
bptxR978Ouvcuy2QOj1ozQQW2VX6KDtxw3qM47gfQdaiaJAgpQz1ne/ZJ3Dx15j8ffyCHanzI9+n
EsSKuEanWVyaZG+M65fZAlup+43AIwxT5XKInQsJwOJ2Z4QQ+QnZ4pwNON+WfcPa8FEFd9kA1rnY
UnrRr3y/qE3dYAGkxJHh+QmsTuaoGIK1dLj42yFaQx+e5ZW273YtRKuePG7VSq12Qss/nPLBqKNN
w26KDODzzdlwa0o0eiItMWj7bMXJokm53NCqewxtito5zWf9+m/GcfUZUYIWhuxBXhGNwODbMTIJ
saH2iIG8d1apDoxv7258VfXfHwwE4rXBJt7CXEZHdcLLwBQ/puY4tw8p7KjWjfhOVzY17UvsuiSv
0v1OiKM8ze+W8OjPsWbGcAxXORC2Rv+EVd3H9kObANMJSwjXzW1YpWxxUbKsJD+rwBe0bUE94kdx
PkfOSlkI/N78y7vHacjR7YWSnf6HRuOKwSRZPvhD+YwN0X9+FkFPYb70GCn17ffN354dQ0+8T2jR
PE6UJhMsM9OEhkNtFQG0d/ZGnBet3Lm1dILcLKpftd7YVyVzJUtAmyBUOZvBwvGKnlzzCGbF8789
SaBugp8mCXodxcLsdlIb62EkWaMdLBLfG6QeSUieN4pGaS/thogE5vT9dAZckqVVdqGzwcLzX1/8
RdUONA3rRovHl8RRHWI7BFZo0tk855MMRNpmZoMs09RWr4GP1LAiwqivyTA/hhdjcE7MSRcedyYa
VC+F28s1xtetVozdQI8yIHGi51tBJ3EigztGRtQS2KmDDlc5y/XloN1r6xEk0xto93P8nZijGwDV
Q7UrjsEu73qUG9v/B1lBM2NvqKvMNn9BogstKMxDeEX25XWG52hbcqKNsvHDpPTFm7vhhcphOQNT
yRPcp856i52qsLI5B5UVth5O2oq4JIVv2EyIPsMDov6nN2uYcg9IcK9ar0n567syNxVNwo5Pq4HF
rYO7GBp9N0A1nIWPzhrFrJ0ZroXHIxJz1WaNWP7fTyumC4g+mjNW8ui8X7Dq5UW6A//LRSHSwI5T
WFgbh2bVWCUImkU+/uVS06UOwvT14b4xKRIb0GPjjgsk3ub1OLF3rQ5R1hsY+R/nBTkdW9ipyWbN
CBG3orrtyad/bZd5MK0ZbG8DW+F53z7fEykz2xh8N8W3H9FG4L8QgOkbncrLVYwkSh2Y0pmLYs7W
jz6z+BeE4HxnG9yMvtDLpoFJpwsIZym0emuEUL5qH9nqyuFRPZNw3CYUrXV09E4JclD4JmgCF+u9
3m9sBZhIOOqMoeIQn2A3owkKNEJLIKbfVlHqfhlbDKR8C5Bu49QLaHmfm7QwPfisakkOIlT4zUKg
bfIsLy8vGEPcej9Gly3QXmvUXarXGhMeqCOM7Fpe1TRy5rWy228nnkWkf7Rn8A9uhnIqGlQ7OtTV
XOSHfbT1M/YEySG4LVMbA10NZjS7xMT6LQk482X0vKfb1HQxtlMUJo1uvAVtD2LyqGTJQKRtgX4r
emxedP2QjA1LvDBSi2BAKesCsl0Ud/FiUVGoGLZTtcY+xqILm0EcD2cVna9PoVh7Z6vTYS6QNwVF
A9koGxehAgqLV4/9I9zugt3zTWBWoNVLwXB0FTy6Fwp0xuabPWvGkz8k4Lxi7nkkd/omUALnxuwf
26E3b7nmEVjTfiHqFDW9u5sCqpKKZS6YtrGZRqdDocuf5vvTWKWlMHCyCMhNoq5GxHzuIC8h0nA+
HnIxdQ/gtoXCuHPE9wwSt3GCADQPNzc6HxFx6MzsnLMWWPo09ZRHkiihuQPU1tmXn84lgnODWjqt
ptmeNje58u3hBFCryzSzGxBdaWEEdaF90diGlqwSB900nlMMjBzL7mFcLkpYvuQBhn4CmUxE8e3u
CL4LcOZoiFMA/mQYDGzdx8k/wotKGszxHf9ouKQIfWvGw2Yq2beQXYRzvq0CVtHqIu82N40K6OU5
fFs/0Qv+YFQkl41HjTLW/CCq5fzSieyS3aq0zE6L4D6QGIDp89W7XRhqwpFW3eSmkEUE86CpHMtU
VN4Qm4I/w9z6/y9FVO3yvzpgEUFEh3KU4Pkrb+X5BIaUq3J85sTUPgaJz5Qy8E5GUrsa1mBL8KXV
Z9KMYfy30o8Hr50KMJhP0FL5+o+WkPx4HP+LuM1/SpBzj3VlXHEk6N2Bm3S1byCCy7zuqjjNqm3i
dkPGEMzEe7aDz1gzOkS5clrB1C/w8zMvsllQFw/DStCITQyCIt5jlSUHvM7g8kjXJ121JagGn2R3
WZP740S0zdGWob+niJ/ML3Z9+kCHL506PJu7GPtiaSRY7MIGXfM7jS8DkcJIw2zpzUwTjYpqp+zi
J8omvXvO91IBd4IeVbIFGwJh+Xa6RagGQzddnR+jLIVYo6vGEyTW4fGrM8qxBHTFNAIKiRruTZG7
4kT719VEt1ZYqQ3MZceuA0uf+IXxAzMRiNgJ49WQjQb5wPVPIUe7tTtbaOrQBcrYl9ujOECDsO1H
Mvqn6LVMGeTGRjSA2JsV71skEEtfU8y5V8x96BZr8g4wJo7F3h9//zXC9ddCW5Lod6Qpqd18JkTF
dbNytrqOx6m4keSM2h+Tl3hPdjnXhR/aS1CT5OdqVHTOdvA0pZGdSaTdN1p5MnCtC7c/X5nT0O5x
X/zwHADvpM6SkekGhlOFjkulrJsHMQBuJ90Q224/ww9nycDGaNPO/vSs0OWsrGffGmm5qNvh2uaQ
AIIXqeSSnfG2WJtA32N8e1A0ItqXGwFYLw+hTLgY5FJYvO8LFOqChs5jmFKXXud7OtDlR+M+aS+I
i66BvgGZ9biM08H1W2lrJ37ETJIPrcChvPQFuLKfq+9nTCd7x7p1OZKhIWuhM+WZ0mRyw4Z32bAs
qDTdon0G82irSEzDg+w6jPI5gR/TjTc2eY3lhgF0ZrnOAn7nZagwkBrU3nNmwnvpeLEYivX2jQv9
PU3Nx0jUFwSPvdAiFBHYGBBna2LZZEiPLwUBZcaFHbXbpZQTEQY0s3ZxOBs708MGMCT+VV8Z5yDC
llD6GWuj6H+1lQmSl+2aE2HI3O/5EtlSGH946C1Oy4SVG/G3ZhbtkXAvlfoMxzoLK5BW91rqT55Y
A9gbKK5H0yKcPvlAHYybJCKqEYqyxvxs1OZtqLQ9sjPL78jmgZn+w1ax1IKJJagbPekuJJ5C3KsG
4/tcoIYuVqUmc/iTdzXw3j8NgpDooC9D3Bi51rHasLb/UvycmFe3Eif6R/0FSZIlipS0iS0h9xKw
KHmQQixR/7NtdEiYzh1j2Qmo63W8pEir2Dqz2cAfgBtYngevnBMZXuPp9yjiS1JqhPKMltMt7FFv
R8X8Ai4YT87TcNcR9tFpCw9oe9e8vb5WB76ns98PSFhWtl6BPh4FzadgogM5QCF9nkv8Fg5buG90
jLszCL0UXxt+qX3TgGYkE/cPnfSJVYgg9ha8NwhDQKRVzPkS7M0nC0sVrqFF5VE6mRt+8RUG2mk2
UNMLXRKH8r5KZJGM2qhvngcdxKD5OWCVw80LjCbge2r45n6Q5rOQ2fSlicMKLMc8dqTFxA3GG1Uh
PrGbl6/0tMI7SMyLU2rRtWfq+Ju7JgiQUA4Ot6Y/80zmwBroYnOYPIRoidhW2seR/4oh8kY840pz
9wRzd2/0gdBW2xOyoBO4DR4O5Rxr11oBuFtZvE+oOdTDkfH5NQuGQfWOTf3eVTM6s/zOZZ/COflu
Jxpfv7UrA4gVR7Mmaqz5d9AG8qidNoTV7wSUhd/5/jVMEiESTqMc7ZRl6n4F4B51paB2rf0GR/vH
t74I+4RpPXLjmarmhUEwWEZ/Q3lRcaHBTZ0NsmMakMu7suESmev7fgHvQlW8W+FaXXa4kX7IYiFc
rclvUFYd9N65NbiXxxpuEgNS9gL26cuk63Mq+PZKCv1G1gHd0kqMNQpcH9hNqQ8uUXI0CtyN9z0x
CvG+Mml16MMifGEA3iz7Bhxn9bPFAnREanq3dbDPbrTLMUlZDsQlN0jD86LuVpNTIjlWrxSXVfaT
JX8O4JO7Thk4DY/iwC2AGh+LAPT4EDqhuSzC0Acr69askvAG0jDooG0eL/0tzb0RaRNPq8q6q7T8
U3lMl+1IvcmZDrx+QEreBWaCuUAkaM5N1c75sFsXlqQsRCT+WpHEuV8cbNnYs0QhzHr1rZcrio0+
vAXK2nXAZL0suK95Qhm8VS2QL6C9Kaza/7EmCffXS0GLVeJDUZANvfuXy5cnr9k2lFvRNS/mDzkJ
wXcbzJs7eSiANOWWTesPhCoM83WJArV9St+anss0otgti95nDXsvlYGvKSnfM3PoaS2GH6RlW4pV
5wxrgVedgB373GsvcU5ubztpcX4M2y9J7EHRe4D9O44doVLbrx0EWM2ELtbbXaQkQKpQ5MRfptUz
WyYD4dOfZJixOLmNGw6kOAkCnp9jt2UbIjU0OZbhx4NCFvrHU7q1G3wOZF+uo6ljaJAPIyCYymCb
zFr3FlNHtP2SV6NFukO+ZWbsZzbLKZ6IZknfC8DWRESDjM5cQZzmgfO+1/Nn/JQ4PwY5y4LaBUBu
Qpa40livQbKGjIXXTdgzHajuXDogHsbd0CrO5IXjFK8bdl4EjoQOmZjwstjK/KqudRA4yYzi8u5C
M2Z4EhqE+s+gFjaeWaoRZZ/8g+LaIWuz7v6we5vj033h6xaC61FCY+BVjEYUzyNjn1hjaO5zWNbE
ikTj6xXjPwU1/C1ZZEeI6+8i5H7QzZDdoqc7WI4seXBl6XxI/0/adbYyHR5jIfKmlbJvbTxsgCAc
H6Wgdli+UggXdDRDEjrEU3g/brSmQL4UqbtuO6Qwzr3mSz4rERHe8vJWca+HFI3FV3y/uSAHdpgE
/E3HSyDW1IMBpdNG2T8cN8qRklum+358NWMtpih9rG0INLVuvGpRpRtpzcFaZOf5t22Idi6iu/oy
q6Zr/x6yuZMiFK9M6HtNBAVRlOMGLUxVT3lhKwddBCP23gijIx6l0agTFGqlACxiwgBpk3b77n36
h8kMqnZnuohkquMOqs0chyVlMbFYNJMXGKbr11922Pr5Kkdf/5u9F8m2EdiFXfIlEhVmAQt/df3U
BQJ2gOmEwXv8VCPm+h9LxzSGSFeXFsWYNnh0CCjgpRGKqoPq1vfqLDBXB4rPGt6YrDjIYvnCeYpm
nzocKaqp2mQxMK3mcWUcZq5zapCqY1utnmGXH6CQwy7ZG0rer0cQU/TW862V+3yaVERY125LVHbq
U010LUTz/ctbnaGpF+29xAPFzhpOxEPGyhtBRjQw6zzfof2bfMvSy9E6b2weWf+2qSvC9GaU3mD+
AvwArvzGOSX9sPMmrHKgSWauDC13tmHdCRv0hASrC2TDCRW+UntalUTGcEjxyb0+irdI86yCs7yO
KNfV4Webll9DxxTHK0VpX0DHegPAIUgzxBMv68oNMX/T/GTe8eRyMXY5BcCZOUGNmfL/WnIKC0Jf
c1z/CL6Og/Vk4NST0EZJ0Z+AIlDxpb+RpkITnbf5sCkHNS+blw5KeSddSaxdQxu+HspJYH9IVAI2
K7YQIvr+VF+OL909/6kcWeE/6amIi22Ce6zOvb03php8TPBxCrDZTBqmcitu5QSMB8q7D12CBFNQ
Em4ZiqweEKvPgo9yPZtNu/R1mIjdqmpGSLwq1Vm0fhbJJn4GhVyIyUSs7I36BXwDA8j8VvTFFwBY
yF9tY8A2fqAoh5cdvf/AtgMI5GFcmLfVPcHz1+CJ8uUNKIZnIr6V1q/XTVZ61zkR5bIeICLt+TbV
bp07Od43XzmeLVd/m1efy9CKGJaM5nJCOAS0L8bIYTz+0RCCHh9ACdttPWC5rRXUk2F3nI7XFUfr
sZmW56MuZbFhr+nm8JrXeF8pucrYyOe2H+IP6DOwgJf8f0FdaHpsoHccAUZWBpPlND4SQYar08cX
8dP/Tz0F/1gFrRATg5aXAomvJ2lpahdD71BVaEaSy+MVnX16/7YD1kkcBxdPMV1ges/I2hwQCipl
WK68kdGK9lTCtarCNVY5IOA6y0ceal9eCZzIrX+9JBB3wMJj8DfKYyqs6/a39v1dUIcChVrnPDLL
+5wSKClytaURab4T67JJMRxqtE2vw+/+nQBAm55USkLZ5P3J9zNN3ue+EsXis1/tRT6fnIIfOc1D
gULvYZ56O/8SB/kP8ed77TP9A9LW20FjZyruy8D8bREMQY+Ptl0GCL6hWId7TR6pjrPjbaEmCO/S
CHGGb/fVY02MLeGxJc/51t+nlxB5w2e/atn+rm7lASZT+LK51bE3GCHL4Vpj32iYu00LWKQlpbS+
2aSKgvIEpsahG6209RFZSM2bTlKVBRmsKWBF6YzWnxWMGoPG9n/lai0d3BY0QDB4ZDkc2n5kRBfC
p4Ng0oN6479os9rJmUihiMRbxJKvojt/jbwo38p8AOp1ZURALYtMk0hQtR6jKYol6q9Gm+K53ujc
f201mWiRl5hil6+Nw/i13uQVFGuM4+JWaFB/aiSWmgOKZz5qqUiZUsOPDY24+31s7eKQwNRN5TqU
LiPh89fQmD3nCqhNWHrufPxKItos7i1fjMf519sgiG6S4sgAtFW/OJFJESo5WeyUL+Nu7MtFITMb
eY+GrP7F7g+8PHx4U0qylIzmk+c+SK41nWlssbeDlY4jn4L668BjmnEbKsWGK84izQ3CFeubQm+o
Cy7YnfcixjmA8Y/SrhsK/V4/5lNosNHjSdwyvasygWbYnm1zFMP2hJ9sEZ+OMq6SyF2HqlerXUE1
eofYDRBvMqWIASf56KNKsF4k62ZGf+jgCcG8Zuo4ZYxH0a9AyhCg4p50DRRAka5fe14XZIpr96tE
BCX/4oggpEJ9XtxaErKKFcNJ7ZYB/GekAz2NLnncP2pZOf+5P3XJFkFCLzOedSzw3JscrMxYSqI2
s3+Fyg2pPVUqNIzSJf7Zck0stPK42rdNjVg2R8WtaizUq7NIrw5FCXgKgZJ0ny/HJVc5YZ9wjbR8
XXC3p8Oge9YjROS+78SclZXwdbL8HRjbtTrauR6pFr8/nOGWZJn4oauDCQSVDnCAaaxwztgMU4Mb
aaWVePB2KYsX7cbuv2/LpjIj03YSgSFhZeJo1S2rRsX7RGhlkJppqSrubq38/ebMNhxPXSc02QXw
b9VV9rpCEKEtE/28AJRwlJadN6rb1rLBsPnqALzVKjMVNtNRvF+4M6neSJn+vVwZFiEI4Y/cIv2A
5LStAy3ah4f6BBzoTo36EhgExknyykvsz33Weuk/adNY+99Uwm7qlBoaVBzpRtyDr7kqkg1mwZrc
LMgxx9IcZtNIbfWk1lRS5ylrsRuwGOkwqBZXjS58igYDHBF5ysb66HHSXXU3DZM/aqEb6IXRj07z
CdzsI7WhpebRzWRG6HlAR4AzIgvOsu/HEqZbqHAuh3L+Qwu6ZJr9HyID7zNZGigyaa0HIlnJmWkn
nOAHtXroCXRxmu4z0WoiIcQUqDq4HhtBY5NRQlOKV9UuPDLAsLY2WyAr1pPBGpIZb2twiP6I5XDl
f2TN/+R4xMi5rPd7cGxzcyQmm3itE1EO7mnkXO3EfO3fV6eO0ccjRGudQS3+c9+aTz5KhZOfxZn6
FQLyoxZ/eerAvi9TGkwsUp4c24nIaxlMa/BnfKC6Gwl9/yFB+Hv7TzZ1r24ME8kAlNPaBbvF5oca
rb6ZXiavb5Jk/DDsvWxy+F7PUHbb4RYNArkpPuZtZrgfnypdaXYYIu3KsJR9OMInL5tSpcd4XhhR
OgSkGOv+szCY5B7OEb4TbFrhR0Y46fItcmIvRvkPtRuBzz64a6KmH0Qs4mdyULefPuXkQgdUZ2yx
/nleGCmXyM/EbcMOf5ITPKfA8RE7eoa4iTlSpt0UeW6/gMgDSM+IWq7TNsWB2lH+9yy2tAYin79s
acsQeiNHIr4MYi1Z8+4Z86G2wB7mOLIINomULcV8PQ0PU0YsNLhuaPj6bKgvavls8maF7HBUjlRA
HQwfzE9gb68mIaVB69n2bwUR+hm5qtL0pB5+MZD1Y/juuTxgD1SFHlPZs9j5M7Kq6ezedzTBJxS5
/gpJ7e2+1jawTJ94WqD8hlAg5h3YW5CJN3y7rdH0Ow6luSfd7euaZgy+GWTzUWJBOxU+Rl7sU7D/
aTjU7s8NIQbiW+f3rVQTNZwe13Qiy6XUPazVk0N/EYkQOQi4/G8RBW7u1ADQIxfKEW7jAMWEIhJx
9y62pNvy7ZMt79pccFVQuDpsNR2VvNoASu2s+DY0Xumd3mDennGLkqOHdLtdsIm52FQlUm6vLoJJ
RQ3ULD+vridYydnSnuDbfvLMcd2jfVRsDP75AQG1SOtLJfm2qA8XyVb3KMTRoXf4Bi/94/BY4HoJ
9RpvAPaWkSmwG3Q3J9vR/1fvC1RY4uHVlHY1+lp843EG8stAe7E9mEpN2DXc6a7aS0YiMFtFdzfn
ghxJXbf7ShL8xwtDXoVwig4d4DyQxcWP5/mLOI4CLk1ZCTTd3P/K3tqiwSRtOpuzttaUu+iww4FT
56HLmk21mHWsCx1JiT3kZ45+yzdxnkFQl6IzAZIj7S2qy01M+X5T2UOc0+aeo2OGRCTB7XEglq9Z
dO3Q6Je1JWN2DknzPaSQps2GR3IuRBswwR04loIO9SOm8G7SrBQQ/JbDhCRJPMpzzGniH+dt1RHk
e5XFpv6omhXnAS2eRi1p84a1mBz3sEUpX3GmuKA/Oy7Xf5dCzyjQFCuUD7/L/mEjQO8F2Kl2l9d5
OGnHSMWqV7HwWqazlmmCJ7QD9h3+SglowDTaQkwRl9ecK9VH9arOUMnQOIemBKk5qDqeU1EMRYQ1
19Nze+SgEClCZUtNg9Ntru3c/dpFZeVg5L03G4ltQQ5SCZgAYp/9hUPIBsaR7zK+NRr9o2OpUxbx
TmaRtN2rLBdkJHArkJlVNq5l+ZhtWeqqZZQSOrMHEog2tD9g/VV3UwCX6bxQq3fJ8KuEZa44fNgU
xLidBvskqifLB1yhK+fznMRZP1V9mmRG8HoYOJXP2D21PiBDLilfRKxzEnYbJM5fMguLc427N6UG
kzX52j8et71AMzv2/Gu0sExA0CXLWQjXF9zfQres3l2q7jL0HzlyCcsNRxBEAMKXqavZpLQ+71BK
dnblzWOzczlooZ756a/dZR7dFczBb79T/1vtQ4C/A8fWg7cNUPRZppmvpUGgeLJNa0ekfrE+QUQ2
A0b5LHEvSPwnJ7IRVLxTAjQ7YjFnWpOnsFieq3LgHIu7Cg3Cs3uQLNLUxW5JutV7D6w/l+oCVjwW
ame/bCe/PejGLMONlBMGyUJYY8Bv1Ii2QgIlC1zSedEh9ylN23q5WpnhipcOBC2fg238fzJHh6fS
ssEKJo6D70Xw8+1Qa/QDxTAaLlzTr0G9zU1KvDvN6g8oIwTojF7Jmus1lkc1YSP4x7CX2cuplPAX
h2QEESX6IRRcEjeEvZ3ahiaPyG5I15Vr5MafAv6ZCEoOCUmMJrEx86FCdR7iweEe8C+F+hJTcUAX
/GQB6pm+r4m9gpM0Hp/ftTsqRA8l8mZzqeMgSjPOIzSdcAXWlrCz0/OAk/D52Au9itSAurgzgtIP
mSW0cTU6qDTnTAr2IZQxYj6Sf+GeIo6CFq4cwhfUMUkKZSNOf7k7KqqxDmuHAy13DWKOaoLyg+QE
PSejMNobSXhK9PWgdRSdFG2/uU8/+hzojcy230nLWlE8rdvaG7QFKJ3Oc/r+9MhzKuN01aa/T8al
GVE6vAmtjo95LNOOoRQiWExBXSf/rhtwRbJN5bIki9f6Sb/5c2KJ+Yqtki+y0ra+8jCRlvcOghNZ
HCktunHS86B2bwoNQfq5h7BInoJewOolWqsqLQlwwdj1sbjiP3p91Fei5wUXwtXnveE4FequBYgM
3dqQ9GUzoXFnO0DJALLGgITLoKSg7LGbPb98Ztkl1tanVvZumpugyNNiQ2SXpq73P4r6yRB3EZJa
dLnuitmOPHy8hV5CBKAKZnYmTLasQtJ70NvUFeEnXS4Eh42jLSTQigSzBBuGdGyfP1ujKlgj/KhV
Y+qnts4AowrVprm5JRVF08XGJe9tLuoAQ+CMFr0apHYKThej3oucp2W5P2wAuszBTSswul2IWCdG
Asr0oHSAh5HTgKie59XJW2b6YrhWZV3j2ImLYcFI8AjbD5MRy4fv0sZUEtEYAVwR3NFzb8zSAbpv
XJrVilMquE6x7qsC297qnPn3+q+tzlnbEU7FtauCkh8+PanAUCIUbzGiD5QsaQro0KCuvcOGY01D
axCskWOLVPJuTjeSXDrDE3EFSqSgy9OdFp6xq9SfPsvHtkuZvd/kbRsqfLwpKR7vh54AGETXhFtx
TucrrA/7DsRKovDo0thtpuVSzip56DJBnWzlUwRXx3C5b8V6Hl+h3Kh5BP4+dXA4OgBw/6x42pGb
eZzCIwlIRpZnOWCoJrAcNcD2UwJPrso1oam9753YvC7gz5niO+f9tJGXYCBygWgJdD51apG2bD2L
yQvsn0npph3JeX3X1COnNGCvD4qpfZdKw+qjFy7CV+ROfp8WMGvADDpZ3K7zgv1WPes0mf8c6dTa
W9rurlVEN8hJbrZb2arTcGogAOYFhzLPvumeF00RaSu3aic6K1Od3C0vJuE8huA6D9K9rCUrIHOE
TL4FQuKPtGAWM5HQwkXLhT1Yh9GVRnlSe2a3W1xDvz2r9l4TIfFgy7awKC7pttNS7I7DNewVZvtM
J1W0Yhn1haVITcxeuuXaMnVqFnzsoQI2XqriejLbz6sf35nyRKVTz0fT91pPEjR0vIXmB4rvT7yk
WVelxqUiEdr9OENsfBy+yHxFuVJP+1p2QDpS6D9NkeKhZqRJviW3vEF1kg8j6vEi8iM7ORIrvRGU
n9OfTgm2oThPAlT5u19l8+B+29rZcHD+Mp0wNpKSp6hyvWjj4WFIKAmoGHq+Fkvaz+jTOQegjkkb
r8AprgUGO7H7pcZgP8u4d2kSmcBYWxbI9fgcuSSWM9JgtIVM3oRW+X5k4g8ylhty4g+iIkB2LbCO
jBT1CyQA8IlSm3ZIw+coSi3TWk6grxZiObqw6ytNQ+KiqA3ChrCpsNcIrbHiN9lwuPJ8vRlc1BoT
IKJ6FsWl+zvJKkkJNJlqgwWLHnPlh7EDVIDp2mkk2OmXhDY3mpxSzrYdTzYaG7YDeXk38yynL9Bh
bFvs9kWMnGfuJPIN6NDqMkkJ+FMbXlEs8zj+Yu0sUbr+v1WjnwWVHOADVzvxgGyDldR//BEka2cG
GdnU6TmzIuwEyYQ5Nf8qlttUvkEw8lwyI5yFW0uqmLDzztKKLWDsPYjyUEoTteKAf1/ZooY8sFi2
MeRa6csHIppU52lq21JcreCQwQ69avIcLHcjkXotN8joRadYC68Ha1/tp9+KeGt7JMcitRekvM+1
LCLCJzohM3sgEOMWJ1QQ0NlcgQb4sYFDoKA8/9CGZIGsmp12mieZhmuG4NoqQoTmsZDCT1hrZ2MQ
uxED6lN1lEWn2RLF+lLjvIXksBXK2JUkv/Wu+PipKQjOH9E2v9VJ+G+XIJY7WBOt6TkDvzgPunGb
vG0NCm6Y9pq08s9TPdbcH2WcUzfz+sQyL5zZZdp1TiADU+MnMb6VsvJWrMJB7OMt//0u43sfagxG
dMHN7WmNxWvornjire4F25ADl/Eub9MdbG2LNrANTWJSkUQtxV1ygqFNA5CnmEn+60Dtxuq7Vq3O
dyhCgyu61pIL4cjaxgjLj4+1/u0JbS/qhDkGZ2/FLvIpOQcDqib4cFzAlC4nSoq8lRhmE2SaSLUz
nrWCvucwAV0ZTODIcR4gM5iQclqNMy93x90IV9RNwu8IODJccgyq9h1fvdArjj+pgU1wKqooVjJU
i4pq99BvD/oN797VFdOs/mcyMsBPUY4IFqIznX9as/D5O3DL5Clcs4L/bnmldBV9Eugw2AixJofh
QZIiscnvG5Pw+QU+QJuvDk9ijG9YB9mAcUjmWjYPdHy2Y4hxeelyr24pXK8Drqtblvn45fAVqdKj
SoU//3g4Vd4i8Ac5TI+5LGl3yPQ/qnvirtFDSQMcL8HZcz19RCjGM+KCnFXg+Q1Z2jteiD3Qtbzd
1vjWsi9j3TagqsoMS4qKCtAQFOa8eWJu1ZXCwNja/77x2XIyp5KqRb8cG4O/+h6R3rObr5+KnH0W
6sSYuIqupvBi+I2i2fHmo72SrQ62CIICDEV/Mf/LQkKDcjZFRdFnJjdHSdyqIswwft60QkBnjYoC
UHbgV4NIhw8ZWe2OlxnzyFXzCLrz2XPJ9RHjIbE9jQydIJzLutLq2ZHoxv3EU28GfWVFDVieVUqk
m6bmwRuNDwLeB51ngatDU/oRO9r+TKwy/mbO+czLiWMA+QmoOUQ9B5zYYgVHiwnzGvaK9DuPXUtl
TF7A3bjCmURCKjQcO82TVSKvEQu/sLV11GhY7JYrzFGpFujhmFR8delqJA9zydZJrChdKlIC/yHI
+IYGTqQrbGjE5d+qsBcp04E5LfGOON6dZwcVS1kFm3kkLF50DFM5a9JNa6Dzhk11V1iQ9toCRK6u
2QojdmHLQ3Y+hZMJGSBhoVye9gS6N6xIP0haf2G7UH4ZLTqFMaFmXWuQ+BijW+SC724naWiATw+b
8/AnRC9QAqjmzY2j6z8Pq1bPCxtBR/jFqtOOrqlVUimZ8q9h8jt/4qbNp9/Eg9QcXlv7nNFR209m
Cui+a0+w8ssiS3hfUTe8c9bows5YlZsW3Aeg0bgbJ6hYyKAg4caGPcl+V75+ueFvXNNf6seiMdut
B1FFYnNw0hG3VcqVkbhCq7UhkGX5mYY0dLvVi4zC1xj/uRotjhR5f5R4zAS2U6g/Ja2o/+vELFyY
cgPjpx65Z1jovcd+SOE1uW3WTDTo1A8RzvO5EaFqQEGkToGYQUrGcbXBP/sEENMQt0fD98eb3ERi
bHwDauC8jErCnTXSuWl2st8LFKcHpD16gKf3yRppOFWUSpx0roLvNP0Nr8SYYgpdL+GMc8NDAmJa
fTt/kcMFHB/20+9vQJELMKgs21xIllIvAv+lAOvahf1gaA7dIjjwCGx4XTCD3WHPbhNlWuYshJOb
VAjgK7kerMpYtvP8Xgj3zYu28o8YTx393XG3jwBu93/KW66i1ecQjVlNS0a5ILXbMis4GMBalfaS
cSY0QCckGDOTnZw6XBpRt+pXP/sn3soTrU1huwHkTcJFHkCo99NKuYi1nNz3pKuBHC1noC3zxap1
wVeQ/F9JgkEzAIWs6AoJ6APB+omBkAM79QK63eyq6wrrGyCtQr9xnRpIajBOKNhwAWGJFBjIenwH
9NZsIj/y5NiKmR6XomiURVOQJOTl+tnkmauGo9SdZMcKW8cTIZiRctdjI+eqU0anhSvWw41U8T0q
rCGprbqZoTJJsqA7ItueT+ckQVYt2Kb+DDrBIxNvOQNDBRvHGEK1p34kYFrm3hwaaLpELg7MrORA
qiSOeVw4JqWDfRQAQk0eAAVG52adypYi4qs7kkkECY2hsOdM4GtEQHhvbi0wnhNiFyTxXuyVIl9+
ADwBIHM7EHiRgndlZXi7JeFcTLydmFdorPIZcDcrZu4NzRU0VFCH5YGSuuJG36GTskHHgd/WHrB5
A+ALnc7lHKA2qPWl78Y2SxeuY4S6tUnr5SpgIVLEDBsm2/c4lRzqwfEBWUt617pe5H5fZyyPtPCs
6pI78wz/+fCQ/APkrz37tietvTNcuqc5ybEqjeeNBTCNlwQNVanDrxlauOlVBoTXn81MJ9j2ys7q
hkIM189vMoeNCyuMzkubh/ZNozBYvfAlLdZFZw6MZ1dNMmsm7EWjvjNZqLoD0Ki8Xv6a0yAInUUo
8uQG+hIO2+nCO1kBKE5g6GyBCKUAB3NMffuNaV74ONRjw47PjCl/hscWQaZr2c+gHu36BLUykJGR
OKeekaWShpDVD1/272xbcYcyXH5zWd1zQI80Wysl9MF64bgP6GURq/wDqMuIgB3X8KNTEn/jK0RR
y42TJksr9kpPnclqD9/fB/5lawRzoiZK4xbN3+jOFGSYwECKLbCGFT2HSSz7AskaHU9m1Km78hfq
slhaFK7U9jQY3irw7UHoS2YUrv+BpanxGGHi2BiTnXFIradR2neS3NjKDBwlDfk8EsMTcylUA02/
uVOj3l/ywZjE/J5brbnehDSKHsUkK0LNpZBny6RUlf6RxD+k4tILc8UfhtDfu7vHCDzJu8VyG5Sk
088Q3nT+YWT3yz/CuPlEFhg9ut/20jENNfxep1e0lvXk9Qg6Qhnkm0lgakDVUzG1Qu4bVuC5vSu2
HYXIy2rlB3b1mGI1sJEh8axOjvVzWyiQxZNcsmeAGKjLazdjTbIFXzVUJ6Emqqt09MEJ+XrT9G87
dCrG/ITgmxO1hi4umGOD1TzsA7CynWvNB8ZFm5ICm5wXHV6nCseOMH3P0d+PBkeJ5Ah7JfavXUYW
+F3EQbjpVeOkDMnHIz6EIxqJ+lcXKVHNeZSytx4f+YmSFQ6IrKhEoBYkBOghz60aQkKQe4GEFpJp
A4Ki/LlpmhkKeTtgRJH28iIaRaC6Yxuo9jjri8mHpfVXPvZPemJyp0WroLUw0PqyuURpCFr8pNIj
h8PgMf5AYvAjDuH00srz65HhD+uw5zrMe6eURpnfq8KpDPVn8RDhiAnZ13tdX1qHwPiIpA58mZ/u
4Jg9ERoQcNJh4UP468KuJGvToOmQXdkGnuJOr9z2r64H1VOIr16UBnGItSsmDuR+KsjmYZTu0kbo
jrOMPsPZgvjvgyRdHfR78hXbW7vT+eJL+0wZKQ+zc0nXl+FnAV0tnwDK3bn9am4HvAC3QfHImv2X
6crwvCTgqIWJCfp2HwVvWtnjcL9pdSCmIj21eUnjGj3zqlfEWNL++OleemY3eCGSopwrPYhwze3P
m79k/zYJ4Z0z3Pjs6El80/Rmn3LGEcWhzde1htmr21yhHIikBnJPR0HpBCIUZl+VXG6iVblYhwMJ
2E52rJ+m30BpVUFtnINkn5xz9ys2M7aGvVDKGHdcq8U0ZyVH2tSZYjjMiucaYvKcjDRrrX4rArCg
Lk40KqwFngqdZvavLQsW6PNOorjvsfcxZyF95RC6Eg3BQoSXYXsy5w4cOVr01ZakmQ/nESd0EhJK
zH6YeGsqYe5DGN+1dJExxLb0GH2+C2NNqlT4TvnxeIti7GrNt4E9j340hlOwxjRkAY9LcTJQGOHQ
I6ND3zpWT9/P3qDMkTTu1DDLkrBKT1XVM/ONqnAUd8s584ude2M5hKkQRGShzpXfBWJEVi2bXoLx
wpftB0uzbkQbyoiu7RdZCdwY5Sdnxbn7F++5uTcejh3MQNMKbxmlMqOQlIBG15Qhw5KSnd03mLEu
fJximCroNjNyfVdk4VeRSTQy04vgbJrO4c5J+MrF8VqzckSkLK+eYVwJjUvNvcyXjSSS1jflOmdn
b5H+yuG9ZwYog8ipI4vtFnxsmk2hqsTjG/Bpj0RfxWg7bv3AE6dld7FkgL8osGQpKl767FaLLASL
yEbDZnMTwRxB7OylzIsZmY9o2pgs2nZ4ntvZN3B/q0+PtuCVWjZR0D7zMKFnQjEhDYQXeQCqzomT
09Dlne7V2XQ+IPVgePYoxc3kKMJSMaL3JXIMXztFJDvF0iEmA4B3uto4HWV7YBMYEXVxFvbUJNPc
GEqCShykWIHaCBEQ3nTlK1f2Scdl4to3SMKMr2uai7+Bv7zx8sI4RkRPoYcPdizqw7cvxLIhn7Il
tRt/xNjI+QqtNECqVK3K1B/l8kIAv0PP8BsvBbwm7DbJyAfg2TvOZDCh4MkyB4/W+Brwjj5KdzZM
+42zoYciMT5sWCwhTplbH1L0HlARF0kHhxA5FIvj1LLs5pJA72A7Bh8Rvsu7T55/ZkoHlwIQbeXD
LuwRf1zOIYOGaVwcwIjod0smtX52tzdoQIYgZjFOFft8FFbVgj+m9lJlIouQAXVp+cijH6q751Xm
tVNs+if9i6Xnj6N1uxx6BHFcOLpYRFWGOuDa9ZUw+TA+FtZmXzndxKFpOqNJnFAC7U89TJXQhFif
M4zGh+bFgRrxIZscrE/qGsw81M4RitVomsLMKRVZJ0zGB26E/Cilf5cIMvAvPkvlyshCtb/+sJAX
e4aOWghbdx9JG19kH6M9X3LveOmav657OKkKtiSgQLSm6cbY+hjOnSORmc1Tt0bBI0z22t+vXZsf
30aDEqjgjZ7NNIQ3cSp2chBp/hACWgyYow3TYA8WGwZ9l5dH8LjUaJNLZzIfq0RczMl6aVuLTY2H
CDdFyYOPDz228ndDJYthv4R4YDkV4RI/TXw5ixYdt7KuoKix81Pue4+vSWJNI79nXtupbZk27Ncx
G++a3GEBGYKCKhdPy6w0Th3ELli8npzH1usIo5k7o0ICpCWdqcLCShtr+CpBdRMNiVgvJjHihZj3
q364E4k8q7qXxC5Hfu4l6wPrSIa4PLxn2AU/jQjcNcXguVqsydFQx142jDJoJm3yOiUI4rMPN1SM
x0sOSA9JMsytOA6s1vWmzeJLsSRAZ0LTqUKfxA/QE4sNgkgfwOVMd9UfJrOboTVjMdtGKsFtXAkf
3+U0PZ6C/CwRKk6LxQne5HTWam1DYgvIoYuRnuT07jj07p9VPfGRhDl91ka3Llw4yFbK++EzPL0U
GUFnCOdv8BxeQ2GbkDc+v/H2X8cjb0mH5H//j/gOSbd6JDbEPb7uT5Nd6gIQ8hQF1RsW8VF3B6Bj
ixYBBbFkMt4M/fwTMQ3TPEE6tonrqEuxxSW8HQrSbVZQ/vDH7hpEI3+5WbGjzdO8+ljzMftOrGEl
+0hAHdUrrKGTkt235XS/LtUFLPIMSHegHQJhZIt1pSFxqT/1D3KsyI/vBUqyOpIceNuPiTZDJsgg
UCyxrYVRE9X2NPlxBV2eRJpVMLMqDGyaKJQtWtc2ioGds5KOjOW7IXKon+A+rw+3a6JGa9giK7CA
BsKP7462vD9gPOP3MkMgjC5NigZ/r61MrKvkUTlyHwXQEWLlWaDB0JuPyl48FW3m5KEXftDJ44XV
y8BrBd3y58z/va+D9WZFLUf+HR24YSPs/qfX2nLakVlIZ4jsFHrXi0w829D1vfNnDwdmyTEbO1KZ
myTeEWDrkq+1TzK/yOUis2zhlALumwXK2WCmxleVLkALwmZG5gIoha1WbvWC+7SpRbyzoRTLwoCj
gaPS8vlPshWfKMB8T2vZtG4e/hMOimBgThm+Nj93o4W5ZDznjb/mPWYkc5vCl58swYZ7BZc7Doc+
86Nc3XG03k+ymFAwAp8iiZlDoT44rApbKqEIgbYbZCbi3oePSnHDxu3XnT9+dcvIj7V28iZjXSgs
fg3e0fHq7RyVJjgsjUEyU/PINI33kun9uVswOJs7Mhc62GvmIyuI49qzn4N/dtoh8ZPJRWeEm2aQ
Vs0tDgoWwEryxjbSinzTlXXmbdr7xxgdta6ZVGXHqVuWLktpdQRTrwi+4JkHM4vHYQoGFjOnNCfO
F7XH5mzlpioFjYnIqtx+hiAYArEKwtbd9noOlfxDpFNfASwb4k6zeyOWYdUG/CHTRk6fmtzSmjcO
0aNlo2R/MmqNYI9m8cS9veHWqkmWTepavoVjwuKL9Dw/B0MhLVuM8vVOwGZ5FeV6AotxTFUweJlA
+uClsPk9N8mzxNxLEOomf+LgqYHcHlTysPtCUsmKI4ztHzr1GanZc5kGXibRgCNXpVx8g0QKOFlf
42bdwVs9tJrOT5bK/4/6ynQfJlGEVeV67pevXa2C9H4rwGwZf2KflNPDqyOPCtkyzlN8bKps9tCm
mTwGZpDS8nev3llvkI6rZYJrebYEHQVz7krx65eEpBCu0hfMa9pTRbF3Odr0RMXTn8NlaKa3Qfk9
ULisHxOLF3UOOD+Inb70ZQKdHQRiE/Nvolwo5Xq8G7IbVyMwsrgfQwst8E36Kjr+kocEbFLrESv4
aNnL5yyV73lYm3/lFGBuUh4RktUxwTQOXJjh26Z+qywrCZiqx1jGJM/qY7e9SMy9/ecj9rME5SNd
B/3f5NDqTWp6duJ9zlNyCqMcUvKB4Np44a4cQlAm1OnIEqJFvcOE1B9bf61Y7M2jYuntmBya8dFj
t4A/cl4Q8UIasWf8zzN8HDw1EKWXEzti/ckE2wW9KzRNw/qnuCWXBIJiJzVj6OkN02/k35L0JL6a
0/jGXySMowXjAGr4kej3qY0pQwFrZa/JX7q8AQOXQsQxbqF5ioFNciYhbi8L1aH+RraxClVDtOGY
iTAvl+phBf7n/67kY4rl+sECrjRXDqlYTKCQewSQRsex6u1WCBH6t/A1kxcBa5V6IvLXJFAivcC1
GqfCl6U+FZ8j7ZdOtZ6NEL54/SjaaFtbqYd25QOd287Z8CNW1kJs/bQjMi4sdlzVv1iIBOYoPtdB
3X9xfavkLsQr+tsLoOwnJiUkf/Fsnceo1zZMdkh8NtyyXe99I5j4/+Nh/FDAHhMlVzTXi+iXgpGZ
efcdJsR2GNAXEJ0pm2Um6WLmz8xIZ08Fdrh2p4Uo8WA2JnbFQd7W+AOA36yUgHzAjDLfUTYvmzdc
9n+X51fZ3xVQ7W+rlYOLMYhAQuf4qeJf+W+nhOUK3gojssh1DgEWbm97i3FSQGKqitCyxOHUnMHe
Tr33br9AQ3no0knhAEYRQaeWraM9ySybA+kzsUcK/gqSetuhCt4q8Ch0iGWYOfeqHFc1UP4tRNRy
qqNPJcdESnJs4LMVE2vwN/3HDmR1o9eAieHUJl/sZglYyaR80kXSLr6/wl7gB/8xTLCG4+S3db12
pzKnPAy2JYqb0qjfUPRZ8sH+6ESa1mdZErGEN35hicQCNxYHfDKV5ZKigp8RaddKeXje4Ge/hLcc
2HvwTYrzL3ACoOv9F1+fGq+u2+cMHlOz8Xw1UcPZXlmUoRh6tcM/9t4Q2kppVJA+KaxHhRvIYg2z
aR5GuZAjUqmWNe0Lr72RLbdny5WWHAXQXAsZ9StbujCkhbN7mBJ34WIQkDrOLfOeIcdoae6Ezyga
KkUEkGedH92I2xgGrwm3qEDMhUYZMMskbv7UrOCVmuG/hp540iNGXCdPrUtbXb+KtYanscPmAad+
EryaSzy7VWE+m6d9eT6cpCveCYsU7aGjR9Fb/aMZpOi7sSea978+1mkTmFVfCdXmBLUXXsw24jzZ
SRWcA2pG17zkYD7/Lv/WWkeZvz3HJvTsFclbBbB1lgYJ0c77WQCsFpEyHMOyOePwq5w6H/ZhHSxB
w1zzKawp2+j33CraFgrrREEKNJBIwxXZzsTcq+yioms5Ph2KWgrqpYeTNXCYT7xrSbH6hrnjqAvp
42WlQ9KJzl34zjBu4KMYk7rIg/Kxz6VA09J1xfeKFMbuljYZbwd7nWs/ektk16A7UwfouFnNHmz7
dh+tQaKfF1MwJr4wG9vgn06xWOCjwlNykw2vWQS+iMXKL8q04pTX3BNvGAT/yD+uFGArGW9svooy
uvgie9zwQ4KtfBNEtuM44Sc36c0ABY62TIVJ3EdNKYdGTTyoffdL+odgKBnNVbj1oN/B+c90Q+pR
lG1vIjBuOS8jYZ9TzlM9b6ZP32C1r75BDhg42Q3Ii9gfLC9wnr9qpoeyGtQx8hh/8XatGF5molJA
NJKL7AzYzRk8vQcT9XRoZic0JROdq58FYEaFmdUfqSX08hfxIhVXaQ5xSC8XIiT6/wYlh6iQTbIY
uLH+/P0gunNlQViIPnn9Hfz0PF4nt3K0IPbHLlN08grqiDZDpgbC/KjKKVgR35Q6If3L6BQuf1QU
Sxl8dqDZCl6iL1K7wcOtmOJg2Ake5HCchsdvEhlrqCUkRe033zAeDjBO3pI8bsxwEP7UQQRzz33h
Z06mm6fnf/7W9A32YIiZ0IaKvjGDiuT9S1NKSRD4CZo+C4AJG24a0cCYVzFwr32JGgGIpEZ9TrPj
gblNB5dP34yFvlnCbsNcw19S607/ivt2Y5M3CgzpWOFrrO7PYvRZob1ymbPZ3CGdIqXVxhnwm4Pz
qBTKaEbgUj4xw5IdPJARR6zXgknrvGufiaByKvgw1mfDmhzA1TbcEJJl5ceenvYLwmw/8NkF7e11
tZDDrcVQdpBLh0umtiiaw3mncwtXplydkbc6xpoB17ulcQzgvcRfpLCYkMVLk/CgNGr95MJh5O2y
AtUjAY2oGY2tui9WnRkiVE3AmNfTMKjXHVXmZBRcOIX9HxWgIXUU8uDO0F08p6AQy3jJJsxAghv1
uHSEIYS70mOfJrwbBgOE+px4riUcw+5FTB14KomQY+osXnCzOtjbk3mJLtqLPb9eOWU2IgIRgoaX
aznCZSVG7orEB6aF9fczFLlkxx4xcDdxOVl8ZUj7tM8xZfSbilU4/SZN1wC6MFBDsMkYNPhrq0US
ZCGQnRIvKhVUHonVXIEQvUmZ4lBWLe6iVKnS1pT/Re5NU5DINFmu/4vOvvLPz4XNfmtDNXzTXoc+
212VO16mYNt0KQsVyBRlnGoT3Mup6FQejIDkQ/fgwqSs7f3B/lmBvYinw2CiiiKRuAwxi2kXX712
RHuzsCvQA6KREM6m2K6xyNrJGqNt7WrxrcYR+bP8H2iSsf/4XqW0+HmwsDURYsUOu4K5PEDuuWsT
Cz/5W0KunYMpIaiAqZM9w8v8F8jsqGd3Su9Ddy5gzie/aNCMkSrXJGT2iNsm89PFjtVGGjci++wi
kcU/y8moPpGdXAAtr0ibwC89/YnmUXWBuKVVXcPEUmgkii1CU5Nu7bv7Zn0QDGxuZ5nwhWckpJqs
ia1ClFUSEnZwnrPXqHT5W+FhLUDn4mFaCp0KzZ/4pxiN0K3k234/GJQOCpXjo/1pQGNGBvi1yPWR
HcRGEw0RrVDXtbaBBwxfR0LrMcYDMpNRl9nN5Wq7RY8VJx2WEhvTM52qrXk/d0jY9lMVilZHErdr
z4vTuYQDUs9AlDlHsZiiqQ1tkYdf9QUG3f8Jrd+75GClA9JjxDpA33hfEwCJnMKUA1YuLwHdqN4o
XaQ1MI1CEdLz2JY9x7FsnyO8jzug6zMX6pVasv743vk6mVBjub6vFHy5S4BcuA5SEcsRR5+OldHT
QWgBdYW0y+njVz1RVicdQIRanMagtipANM7uHVLo4+OfV0aw5geTjFqT1Zm5nU+mc6rV6vHYY3SD
7rJoun5yvCAJMCSt56im/WmUYPHChzGIw8rZJzhaVYTXK9w9Zt/s0xBUZ4yMigymXgs1CJxIkQVO
9KSe3c6BsUO7/6RH1X/TDxpjoUeOPGNBj4Ed9fuAgyb7hgUMgbzYze5sj3QUTg5ZZQ+JqBAH1c3X
yog2YOeQ4rLwlftoLgwJErYAgDMaFuDjUvgZLSG2yxPkjJKpqIDQkdmZ2e0GEFahxtONQmh+BzsS
u4ClqmqeJnJ3sCY/N+6IBDXN0fuUQ/qCmSRZhokng6YwqqWib08/VGu13U0jli23H44qR0ifq531
baRp1DvBYhUGoRrhu6Pll/5K/e2LE9PXWEFZ0BIgBlJlEyOrfTL83b7kSZcIDXP0vYpRiRhwUYft
+CeHgXuBYdhroxPH4IVCUiB5/iGVP3ideIDis1azW6i6nhHC6j9IjYlqi6fof0Yae1Ria0AyY2hC
dG0JTRie4LGaVsZgZS/6TtFpMkRklxT7H1jdRZ57zizxO2gRz0hQaoa3xEdUPA1S9+qJIW+Dre4s
il45HB4AlYigSrzsBUgb3wZ0pWL7qf2ZwIvNsIXFeq4YUufotM9frkN5bMjztrOBLO26PKv8ET1Q
/STR2hygm/Uy4oa6XfugAb9eHmw2Jqkdu1BHhyJeaou/Cp7h2sbkO0+gQuB8UFT3MP5J2MoxRyQK
dI0J5AXHAmQc1MKoYruB/GNIbrMAh9AdVvBoFcHu2TeaVzyCZn95sxp2wGXup+xAwcGkVmFWoj/5
JpVy3heFu+qrF5TO4ar6sFVUaYoQhj3DdzEUzgpz9ARkkf6MxBYNmNoQ242x5KEmqs6zH3Pb8YpJ
d4AjGjqRmEwM+8gnkO7zhpv/mO8ExOYHxuYwXYM2+8zNcXwSw42uZsAlLAAEb4WMpz1fGXFg9Fye
GMzYv+tRkC+sbBFxbJ2l6KZ2+4H0Y78UrDB7a7zb6NqBT9smCsV1tq6+xQBVhZbkc4bJUgHAPX0r
CQlRu14/6Gxh0cUBCI/3ytbAKUleZEUT2CHYJXXxEMM1ivrFf/5oSlJDaTbjZ6bvCw+BEijuOSFs
rI2NpU/c/DRf5iKoM+IADx2Z6E2jBN04rffSUAUd+FjkzvKdcpLxnOTMuOPNyHtFT93KGdorhu1I
6oKGOXDXt3DxREXQ9XAacfVdaFkMWolRcTogwM7YWq9tlXoeDky8/25nery+o8/3sR1kWSztRIdC
2xxPUNgL2XX7LDB+CiWisw/yVKAq1EI8uS7XE7BfFbOVBxLwFybOhJuA+s/CrBaXC5qh0Q7+JJ8R
PzzXO1vi+PDQDTUDg7wYJ/ji7MXcMF8UhA5oulj1sy6v0lG35JgzNEZ8QBA8FBrr93g/74LYQjUj
g+QiiDzvkAzDEYgYiQ9C7uh42abrhrh03LBw4gZocyTqyi1Ej/ZkWrP21p42qzwnsc7Zx4XfF0hF
87lLj5DE2//qhQxSATynBQrPoxhXwSVsc6EESx4NbISZ0soydZOlCaundpOckZZMEShaYQijMw7Z
p7iS2maiiCkX27X+CIs9nQ2iu0M5eRCwG1c/P3he/RCB/GCDo/z/2Eof5WnyZ4Bzq64lJwNLjpOw
OHHqgsLFSEMN9C9Y6CxZ42lLSR/rVrBanC/PG5960Svq57ROacBRQfge7VH4FD88Cq2jOthHtk2K
m6ztacP0Zp0f4QeG4ewE7yD+7S0iSGZuI8FptxcUiDKJHHvjbHhWcm7v6qS/2SZD9mUrwvYkl5/i
h0xa9gLJ5J7nqllt020P7r0rCdkrAbIan1tHClg5HZXOka0Y2v0SIG889MUYrdWde45k1Eam2A3U
oyumzv8dsNSiSolYwS6ouC7TQQEB99MY/9TrDw6e1d8f52hR769bT/KKqDuFV6LH3TmDTAQkOKRH
FuIasNhKd5D+qeSNXcNvT5CfW/q0rJVwXhI9YZgk7TXkpSPGwPwY0W9KY5DfFPr4kCq0em3EqXak
OrZmOMX/s0C0VwJVEbKucxHmS1bJNQNcuxEAOXDZDrKuTCLmMOI68kjsYmjwMBX/QFSbp6hQr8mD
c+A24ZjM6gGzyBafKaZcyEjQbtBr71Y1r7quTxyRbL3Lt7Pi+PdKFjj97UUyx0QPMTr3rH52ugNP
neUiQXmiyMGbbI94BQRQnAXVoyvMG+vq4ECFikP8ramAZvAEGNA0hgJwy6zvPI42AQ/wfgT9+xZ6
odMcFMe5xYeA6g+z2aJmUkwSUsiGGxvodVsfyBfqtHSkzDbNxWJ/xxzWXAeQMI6S49Px4FfHywKM
kXHgE+Q9lEw9MDhLnI8Ad4b0qipGJ4jyLIpcUEyhBbVUW33y+v+xgshgxmbzdhUvxgwzr2GPFBK7
lQcSM2jw4oeMb9nlHGO1AT2Ipmd0GbOVCGBd/dbsDGZZGcO1DYV76uQA5SSsq5jR+hnvOEKYdEsB
KIXabusoDRn/kfoDOX8evjRaFqgVNoBF2C8iTsoSW09ERs561ZL9O0Z4vPFBlFRPoTPKyixXTTJi
b/l8OJ2NiWn7LeYh6yEd5ihweCDlTSLaeiGKjsoMPqYhtaZUiElgV9g9ZvC9Mv+1WFCPT2RnCynK
Mvk/vISOiF3JpuvlPQkWM58g9e20MqCJzBMA5Iqe+M4kcDbEQhRONLBucZbrLN5VAoYM4r6FKp1Q
UwNxu3DM7vhIXA34BMcP6FH1GqKxZjn874I1AIKCM1TijszrNxrw8VULf/oj8lnwgenpfcuszRo5
F9GOW78/+AhNFP3tnieRF9K+j9rVdBOJiKFgcKS8dLFRm4ZYgts0UYfudvzXGUAtqJQvxI6zGMCJ
TKGZEMW0UbiFdsmok7iATjA0C6Zfmnphy280RieJz/8+sUf+n36xeNHB1IDS/G4AUZ+sSfplVExV
5eRIotyACi4RGOd+UdRfBen+iBZm1uxlf9L2Dc2Bm+Hylj+gkxrwHdp5Zz/4sh5dfHbJHAmRMgXw
98sbuGsZLzHVHjSt24OSTtvzCvLwEEoTMsHWIK/jWNDAIo74UECo6DZsgxv7mrh2254sR3J7gzA0
tIFz29W0k5TWi4bpQh+Yki4YJKZv97YiWqyyvpKSHdrTM35a86zFl2fpep9bv5ywfWbQ/q/VqgzZ
n3arGEhuQpPHOS1EyiiYM268mjlj8u8n5miBYUa5sMLoTGZy4PrddhPHzCJy5ITinpYIrrDOodny
rYzvAce6T9ZHLw/4BbrxQWYR3dIlenE0SQ3G/uqUaCCN2FH2bdTd4dQhia8Ui429PUHaSFD5KmrN
NjUCaS2O9KyPXzgKjLxyO62fN4NGoUnTJ2fCWdx3I46YB5ZId2hK+zEcSK2LLk7zZH+WYT7MK+Lu
JkxOjhPJ2a9kO3HY8+SYMBHHz3WH9/BrbSqFZeYZSGz1GjZE4TGSgn2JUZFo2wCvbru75eDJ7ZEl
yFsvEcKiB7HsgDBttThyQD/EWyYQbaIMc2LaDVA48qnUjJ8B/hOezuL/xg+wcNaYzlQiV7p4plnC
AdUVR9Bh/7H7xYUrgAfLPE6lli3kd/6SOFV5oj3O8aHkGYwCWqmzGYF/fDrBOFO4YVFSfh6TpT4L
ZiGXIyxrDVa0kuHQolbjCTynk0K03akaxy07JQVljRsAGAhHS21vP05oCatDtRjaOVp7a9QrjTG5
QIiS4iZMWRr8bvEsTZHLMMldbgg2t/7L0wY2aaYmUraDGdKGTCy89V9CNnzDRg+rVAUMa+jWY+A0
6+vU3vwdVLaZd0hlMu7/rJAW3jf8X3/ynV3Nwf9A2r6FhbRFCwd3F7/20N+QFaqLObFUalvW8fbb
S/zjHvzvLF+UgczE5Gg32rgVT+Eap/rRRof/CyWWGLaK7MG6RDyUZJl7J/+wudafGtQzFSixJhwt
0nhjy9thjec3PmGUXwZTwMTHCgN4KcIk5TtcqeTckbo+C2NAsyqStqs17zTq8qjD6muDjn6hus0R
CdVQmjvw0zmyIYJcy3s2G50YurIqXLyErb7+6nlXmcw+9mNinABBCGbcN1njSKFeZzGnr96NjL+M
Ccm3uhE+ADIPP5Cgso6pKXUCE4mcWvBiTM8m5z8LdMFeMLoH+D+59FtuRxDvTS+1Ed6znPrVEswD
O6BcqGnqpTaTYizF8U1KkLah4O+xUXx/TVyp6GhIjb9p0I/opbycA8yG0jk+PHsDN9R0Drulb+Uk
4Dr9THjEC+xYA2Aa4ZLR84GQrcb+91mmLo9cGBaHBktOWWBfIlyLDUswn4+xDqAYKbF3otw/SfQc
DsvokABDIKgoygGDGG7CU+cGA6KSWlOwc/ZaFmu5cu7BKXRYrh/NDP8FLQiG/Iu4Ol1u6rUBrkAt
QAXFn9f5cl+5BQjZJSP26rjUruTrP2g/x0zKnnYpIK0S3tWDB6d5q7PCVMlHa2Nrdqyf5BRWEUkt
1pshIgCTIYAl1E7qV5LAlUktKMGiDt3h6WLDqBgsAWM3X5kiKya0XGQLHlDRdOtTrQbnGBhB8JWF
Iap86rlHYsNKXgL7xqHjcc1NqXVbfYyFPFxF9Mpy1e3kpku/7WyAFmkL+vf6B5G7Ad1Dr4b87GFY
VI32/58qrv2PhIKQVR1xUpV4//3pWIjs0JT2TErVahvosdxOQYqmmMFNokYCcjbrM97JsnGaSloK
FoYR3tPn0o0FKIcwYg/Y7Rf5aeOz7Kc+HfRcvY7mwf8NfZFVmvDmonPoy7tv/Zfrrxm1BDxUZU6X
rWPjEr+ICfUBMuaAE6HQ8Bt+wHwO8L4szIy7xIt5SbbOG5sy5DrEJoK4XaPHpJUGHqCTve+gzHz9
S9Nh2sLW9ULzHOQUeE98nuoO1G5166cNb56YHb+A/zteVBipuOCZp+zlxeUtOsJp5ZGbbkuBEM6X
SfmwRmyrh6/X/XN2T+2LpROrtYJf5JZFefpkekMBFmDN5iIaMeOiCkV0h2T9J1AYGpl1zzQaPzKt
rCm51BqIdd/HR85QWb2+UGrxP+8EW4r7vrnElrf1wc8I8+jdm6VDEsXEIv7E6daQ9kTVH6eMDoFK
j9DbCEwdnkkOihogSyuK8Pg4i3FN1xBQDRJRaptriEAx7hRlrHuakESN7nnK4dexNzEwIH/M88xe
IqWsSDiOK9y/tMJ5eA+9l8vCfES8gc7nRBnvsSdUEdzg72IOlt16S5gToL1pCswOnEkfGAQhRQ7n
skQFcsJ4KqwdclSGKyeWOUhZS+IYmy1H8GPnL046sXcjSgan5c4R8oggT2ZtkWcQOHmeL1H/tfSP
xm+LYbtj3XkQUMRZL87Ap0c4QxeIczSnOiv+6h7Iz3mJ2yrjBZ/o5oReM5FKws4IsxvJAgA98Q6R
L/h8vJ/6T74LR4FuVnlHj3jzjVY2cWsc/NpN17Ki+2wIHvgHgTDh0eypxywSdILQwxvCMwqg+BdO
cw+lejNeJ8YxH621nRJ4fgdDN0w8HzcwqGlSHOsRStU2MtkdWI99mWW34J9TZ3Pm/l9crPusUDao
s/HP2td12Ki45LvVKQe4BVQI80L1qzQNRPQ8NyhVSDA6z5bGXEQM4XA6F3GXViQiFspiyJEmMYLS
FDSsrxrVzN+63sc1EWPB0IQA3AGr/c+giB+0p7iGW3puBDbYRpM4INghzSxT4N/Puo6K15buy6Gu
0tFVoKIbx3ivVXUh8pLvdc6aaaq+f11ccjttKhw99N/3saZz2LIGt6w8IJKrQuLMiH9iSaCL0ERa
baoKNwRpYvCreyFYLwSAHw2cPPW16FUN+wt055krDfGiY/cMewX6RdYyjovI54/i5Us9XDvyBAbr
WOVxs7FRrn+pD+AqF4ThetuD6TTKY8BOnyjN4CsMHrzKB3jbD5S+Hm6AtlfzkGvqmXTRhdZbeMRU
ytfBURVVCW5R/ZihDKRmcw6ihadGF7krUuWfrHI7KZvX0NjsFs5TFW3d236poj+NrXHpou25Eqbz
RqnISXw5L8+ZwmDId/cULaC9JZ4ZpKxncV7Jj/pmvso+TTfBzGZMkZWcAw74KcEM5M9p/2L5V9PF
kK9iH4B4hDYLWysPEnSM52laC6dqXVFANXkRRDEwr4F+MbucM920m/im/QoImmRgp9ILfNMpl+kh
mxZOXPiw4cO2U1VdJRK4TkOXxeZX2eDdxFfTVaPtJrp6GfS/TFRdnagGo4YR9ZfMMrjNSIuPxRY+
HyHAsoaTFBHRgzHFyozkh70xZ1v8JjuCSIYXpLj354uUEjyUKy+LDdT4Jev7qSJtMcQlkoQud/5a
OQ9t5jE1ly40mLVG01P/0ylP+4OlWftnobAm3R/jDJh2G58/sZnHropSRB+jBZvOphV2urXn+5TX
jPs52XS8+H4fIlLv9b8VeqdOhpkkY9OMm/48SwFxF0Z3iZlfCKUND8cipIG6dG/MTPaCMFwAMF3v
xS5GhpIdy9aJm7WfMozMULeqTxZKjbdObcv2aUbc4gI+TeAOLCe5ylokp2BumLJemrfW0jg72WKg
DAeWJFBk9DJO0PNS446zzm/D3gfypCOTm+3+a6BAKkOsk2aHmysusp2sUODuF+jYf5XXeq5N0WZQ
BjWZGMsn8dlUntntI7catt9GXl6fCjc4oKxsb6IOrCIJKvtI5xpUFObjQXcv7D039kd53NlfM+XB
NYME7jx4v8mW8oEtpZAmikU4gwZFo/i5XIdZEvGrlOQSWD6mDAwV59FQqvF+/0qFk1yIDD/niqWJ
5Jw/JfzEdVr+JTB2rgvdjKZ9R253LEpL5VLiPrd23EjrcoThtSRH0a66lL+bDXfVDhaLj+t8TP7h
NxjQnGJN9hysLwEIbDhRIPLH46OHr6wfPeSqJZ31t4L7jp6dldOtjXfVrjz/bm5w76zK3j2pk8rL
Hqn7UeM7h9YHO7B376os53sCBd1zmmqnDVUsFxRWjJ4QxMpNo2s07LwHKwRZ8nFqofegA53StF7D
M/eRFTKs6iU3rkd1JTrLidi92fFXpv6KGXo4UIL1u7R/ty5GR7TWcpFaO/u+K/9HqVjJPSd4J+No
Lnz39psXmpEjnQUG0urE5YovSWy1Dctoz+0t2kSpNavx5i5Paz0VDMro7y/zjw5xk4yYpItYsvea
l6p89UPmvqE4XXKAeCgbhCwgs6QJ7VBocMQiN0fWv2ZZuWMPmbJH3ZOJkYWEECMpMqCa7AeV5CdS
esrGtHJB3QatjGGDYg8VJzHG9CbPyiBDomwVQa1yH2p1VQC0PlNM2U5T5ByRYIlkX0BJCY8mV6VL
jUL9/xitRtBblkQr1Jon00eNku1XhEP1stPQ+WfBHsje2ANu8M+5QsMR6bZb/5P4h1Jh6PJ4efIX
25MS+hxGiSLiWAVxog1dH+/tg0u0ZjDoLrzjkE36dMFI/r7y+7NkicSZTZojYO+7dADXl34x8GOA
mvDkfZaV0hpZJwp8Rdh0wnoAhMmJ3V6ODRL+6q+3ihLjlfwYSBIUVX48soPCeDgBhxU/a6qSN298
17DP73f6dsgZdQ4nv/mVnuG6q0AJOXEfPnwnGtnVjKAfty6AuwrGiJsqjQCR3Q4opTHBKnjy4AB4
VRa9KSEiO4PQJH6xfSsrEqLsEe0bmwGG7i/JeOjPHn+wsGadeFN+IMEtJU32sl51sX+wdID1LqQd
xJT8HjNopRZDik+7fcAE1J6MG8T2nhlSNYd+9mymsqS0kiQrcwReEKx3hpeR9/bTNp6JALv8JMxE
xiSq5ZDNojMMkLSetvdqrihy43RMGfZynAE+NKXOzt4nQEISYjK3d4apAS4ltompEBqFt+agNqqP
vPak5UTcLrfYbczj/ZGL0KWbtRT6TU/ods1JsOMPhKM7Eyjbtfjm7OD7rPvAHy1c9BQaf4Db/Plr
Df0C+6Q5QKdo2Htfv5jX5x0qGDMsYbgdoC5WMqDgghuVVIcQoHA328rAfbKmMykY9pUVtlzU0wJ6
2I9Qqj9fr8d4O9TQoWXmUqORPbyLL8Dd1JVjh61MHaxJujrCzHl1KraynG2wxwmeyBjFl2uwmiTs
oUGtTk8WO+g92Ief5Kc6s4bQ4CJtGw6UGaABITGNeMhkRvIQ3Qflhy7IsooL6p8u7EL/7cU8g/FB
S3dRrRFUK6oDQ4Nli9t2V9F7L11AQNFGejPTdoiX1gLLFeV79YF2I8xtTj1BckwVz8cnO7Bkz5f1
roOEkju++fIwYFekUIfZaaRbniIVjxwgVZCjBfaSRu7mmvsaTATvpM3vr5hZrRbxOIRxLtRELMCZ
xwMUFXNqEUfD30aC0DdcPvEnmj1b4qM+wo+z9snvPVe0A69d+HlrqADdph5bYRQk8jv0cGP77RGp
IfVGiife3iV7dyMD6k7DI9eyy6RD/zNfSxJSv6CFmMWZx/BipfIyVSVl+GnOOYCkkkX1geZsrrGP
koib42VQVVpqXxA141dt3xQNnjqNtHnFovXRBWGdP0/Zum3XllQgZBVBfs1z4j+YS0XL+jAHiim7
ymCBXCcF04qbcAkN5H3slslgdNbTSTvkbUTc0HVp8OunAz4/CF1Gyvjkp2+/z3L0ZiD8z5uin7Cv
LijJWmioL900hnDxSrcu/b9cduHiLH+a0TLRDAN2HaJKg8BUbi0e93w3vSjueNmxgjfq+SbbxSyS
O1xGFjTlALADaa7RBAjEKC+2TWnryG/TOFIPJEb5nW/6BEa3dBDkigM13jDC7AIu9DmEqNa27Okv
i5vHeAQhJBVJvP8TfNtyLpyzr1jwcceIHqoH0qNkaC5rQg+5CQZL8QCSq9jnEkFbxwFmsr3doTJP
9vWj0O8/7sMkWNDYX3fJxXu1ZkEgb/PyCvYePVQSoiGjxHcJMIdvODG6GvRLLEOIjcsqegTv3KUT
3JUfvvr3SKTAThLyu4Ov4IHhXl0NRl2UTkf9FMJIJY3wmt5ky2LJkrlh33aSRSLO0ELikFTjj98n
6KYhebDwVhtO5VKUsNyaKV2ARaEHnBxmqd77j/4nsdtgZI7t3xenlBt2mZ38msFEt3ZPgUh0iNSK
EXbte/AlwMlDVOWYAFh4IR/s5yR+DVyBLWVprUi2KsvKMgyX6YsSxKvJyBYs7KXqmk90q04qsQpY
iMbRyo5FlLZNlNh4ad3E+yqQs/ijjGRwoZQiOG6WFBVGS7fZiztAQ8cm1eUI3C0HCSyNFJwnynAw
MWFZG9voOIVs6A5dipATuo76C7kPnUVMR+Wa9YHfNiN7USRq0pWOxytNFWxZQmqNalYAIBrwY+aD
QSlYR6q2QC3cGt6Gl9+nvtwiDaMYr/PkedqpuWKQFSonFlkJAdLlua8RqZYdo8NHS88YSpr0ovfO
8pOZpnvdqpvGqoA5ABsheQLJtLIayMYkdhTXSizZRM5hGg7/8jfjfXJzpsAwIl6WC8LmYFKFVBqn
E2FsQnY4iJGbZZSkuTK4OcSLAdi73z0C/B5SmMp8hU9Gk/Le7hYoGyrcO3vERW/xCs696NWfWtWR
w5i2hmcPGcvIpi3//cKjWWc8ugJyDqP4PKHKfcS1H7nYQzC9mXBb+L/I3fUB9NrgP85Ax+JL3PRq
1vEBbGztl/OkeJHOQiCgzM/Ir7Nr9k608cE8w0itL+QqoMA1VQja9tVJfuiLe38cCHxBdxxB+AHz
lSsZs4Sfgj/jwj4xyXagPFJ/rnlNPYnRxR3bUnrgwPO5NZ7I6mOU9rqyol1dkr3z6RPHsTNn0kUp
56VUpXqHAnMnwihUim4qVEwCUAGbpZMmoSj4ce3AmkTDv7dKvj+Q3oNozQxZMChA2ZOZQlPoSC+/
o/YFlSGeSu+YO27ti3/1vZNbLtOIOZsAaL3NeFYENY0UC4M8TnaFIoPXToZdV5fapMIXuNn/ndrk
2zAumvMVpETdoupEWVg6JJdszIQl48mGN/9M7PhVrONoTwlxL3yjCCWt6jHa0BQFXrTOO7LRNaxq
1/wOj5gs+j5dM0dG9Kt5QrTdnFFdu3Sk/3NP0kpSsxnKUEoyLiWLMq7iaQQn1pPJ6zdN8xLcIZF1
fTwedFJPgkqOoyRlZV2bWgu4BlvL1zVvEQBZLAngDxY66mAQWfsMzSBS/BGprKp09avzzT3yYP10
gG9tcF84CoY4WqjrT/D9Ph3NILXypKar8oD0g3PY7NPyOwacnojujK8mEHN3M/6UWYVILVJUJ6/A
BmSsmz7cOlPXAwjT3W+IG5SEetZuWoMyNU9aZPatqf3LnWpiNaEEHzGVpsIWpa1FYvTp8pJNqf8B
ujb2Jet6GvqqhRe6osVKmfP1IFZdezX1d1N93scnNjclZL/HrclrVvl9SDcIudmoBsjq+HudSYnG
/6QxTLwFBRfNNEhLsFRk4D+eb87M14e3nsAZuXC1rWGBs2moJaYF5hX0540XIBQyNCMU9sJ267Wl
2y+MMxBR3x0sT2FU6Sy6HOpcR4yvvMb9afZuHH4qGdFBXcpYrO+76wNd/ZEpzMBGgkJOOdMJtavL
8sZCvy4LSrCVfldTR8WXNE7VWfLBoPZPBXTrhdZbfiVtWwVZ/CpsuZONRlwEAjoLVFedF5b1Wo0L
g7ti4fdwB/sGeLK2sT3dKBXCGcWQUHGTjiojxvPAXTeolrytiU+RXywT/W4Pn/pUsMylnQIkzh/i
4TPVSP7YlwMovsXoplYpxb1+y1dIElmmPjg2kFd13yuCaZ2sxcGxCebnW+BctBKfeSHPxn4oqbys
NtoAnRKdQxI0RT27u5elpnSbcrMgLlM/q18YMATDVoRCHa+k/luj+WSx8qRR0JbHeHcLfNZO5NnJ
KJxuQbzJpJggkFpqwNXQ5BCGFXIwhX8tOkS8vXjaXji34hsTQxtdM6tm3/RmXIiZM+0pHcpUQ7VK
vnC1RTvSTY1qu3RwrfIDv5XVondz1KB3UIfHs4RORf+Vg79T0sqYUjUHgAvi/e1GLxtLJRkb1yPg
LkJ07lgGZwVHmUdfGCjQZW77J2mC9Ufzw5kfazleWmh1cS6Dcp7yj688tP3YW+34FHL4nwBeKjfU
CwRoRItpfYl78SCxvlgwmumXhpLKtn3BcdebBrgqqkPYfRz02eDj3zEOhn8sPq3akpJVcaykO+/i
hV8I3vk9IhSJ9TKpXmvnlfyFlGjkJhHUPxuj+8sQgyXHR3/skcr9zu8DCT2Hr3vy6lb6d7qf1pU5
fdfGarFB8ai4BCGHlDq5VoWyk1Z1+jPFk9qUAvcdpjV+hfSKst4CCE9M3HBOdLsDqEYFewtexRbF
5NPAM6Roi8dFG3BlksotT+JFZvSIu9JRb4+kOlGtC39mSBf2F35BIHCCKXXEWlBvCatvXyB+Hwjo
10q9BvKKXgdCs04AClPVBD5eDZbvKC2VB1v62ywYAsDtQPQ44tLXX8oGMDp2lYvop55vewT0Siyk
oU6/2/3fRMSfd5gQWKdggN5m0mslcfJvFIpxMrSKN4u3OxK0dRUoVDKQYIOnGc7Ekit1x49CXHit
6xoFColnid3R87tzJ5KjqZXWV6wr3VxGO0ycL30nXFn8Vm1APNv0XNJBuq/jAF3GmkP5wj59G+SK
FWHUI+zg3IJ1n1VG2CmYjcFVhufQP302et5xm9P9g0aZTNlay8vmKHIMCk4auUjT5jVVYomNCC2n
mhaysluMExL93zNh8cab9IFyrbAsd04OcvRybBBHfUlkSmeCTx50aD87pQlSCNBL2NyfWKUrf6G6
7oCsFdVrVfwiGs+kJ2k7+0OoS5K5KdXTr7QdM+1l/0ttK8J5Xvq8Ds8K37/2PPPwv5B/VSCRPJ10
vfaIWPARWnRfpTcPD6/jPoqDcW3cklOmQscDIIvSp2z2MLZ3iwKi4iVIQsU/MQCfSNG+5kKiPtew
izP2F3jXOS7ymmkSHcaMMGz8HzVbCd4GyMwCDzEFzeqygrikzruxW6sn7DSQn417N4+sWCxoIEeE
ScvKLcjTF65RxZwkbJf5TungGHLLCC+z4x/Q6D8KoH9vAGhx/Dj6QgWtBgQDdjkYaItVU76g9JaR
WPDqXhzbjcDhRIJ/oiUbY55ojQv4OSk4DZnvuvj3wXo8CJ0kUI7qa8NnIGBFp8BCrUvbbHLZRKLD
cjdHH+r6PMD+nIrZeRFe6yQ0VwjVP2CcskrW06RZylv0FWsVA/w/JywyOuj682bmw6uIWCFllxo7
3ZBZu+w8QrRtgkitysRt1LSx9bqfciYFjxkm+VDzjGXTwRMRlsyfJNUGa9rhwNsci4l12cD3ZezG
uEc7NcbqeWHjMZCJetcM3G8oh3NDeiYzHfRjGOFG+Oaazp1N6uNwVYaUHOQJ1iA7MEj4uVGo3KXt
A8HM+5N1uXLb2bWvTIQVy+j5Y4vp553WRms00zsgJsCcTIYlSCGR4kGvn1E3oByz7K/NpylAmlI+
C7e4r5+a/FQ4qG5V7uS7lrlrG7K/XBR9/PTxjvvK9antQUyf5VHOsGIUjaYxg0VoFFAuPcd4LBVP
4z4lQVSGKGJv3eFY0tTUyEeHXgABLhGHdlJuWFQipUe/MemD6eE6Z2cjvgbKzoIEomFbm9o1ONKk
/ZArqTOH0Q4RNZ3VQEaqM7NIzH/JP7e7boYhq/5+2+HqzDPU5Z1/okZW281Ylun4t9TrSkefRw2F
CgpIWe1XA5Y8L1RSVOeRGFEReZo/G9pmh8RC+oBy0HCYXQ9ewJ/YPr/DiOX5HW4FqdLCOeirZ293
GJyn6DVK8PrtVBb0UCBuC/CDQHm2HDoNTxM4RvhyLP9+5c64kHGUVNVp3J2bEyNBhaYdiCU5o3NB
lOQ7sjSkoUsShO4nWCiMaudNLO7g+tEimt8jpx/7sb63oAhhflf+GZAP4eKtz/n/NGA1qQZcXgOb
hpXEj9d4CPlueu+4EuKO5bX6wW3xIvdtRuM30VNNE55TfW+A9EzoMvEArCeLXZndHGmXk+Uh9Z15
T/KFXHPLxlLYNtLYsWXmeOQbTacDMTThLTr6KNrZHkhswqTLULGhoWGoGTbwxJ0yKNJYxfjl5+md
1sUJK32ULA9L2nMWK4HIHTSuPJ2cbSwyEflvO3tBV1IRBWgMq7REpN2SAOzFC6xPp11wD1EQzShJ
mcWsp7kKXtmHjYln48Jg/WQR7C7WBTZr/Z1e3ynJ46Qjtwr5pFfdZRafbyGWb8leitd0/patfNdv
uzhegiytVjW9Sc6L+WnTdVqKgBxgTYvEpgux98K10DWIP17ENy+NsFUUeZPK1gODhX6bEnas8bG9
muyIhrEA2eL1s545cFO27QwMCqlAxVB9kQThRoJlH+HB+5O3P/A18+56AhWPpJjWE2vZlIp5ge3P
BD0bcU65r1AidPs+xSrDcpcQuQmA7+acLXya5adzehsHqSLnc6O0vodJ/W/nRJ5aoM87YafNfigl
Jlz3AUctk3Xg5962Iw7lyVc2BAdV6wPAEy98zZE4Cpcgpu7j4LzGMlLZRfgg8HwlCEIjgfKi5zq3
u2foX+c/HeOP5LX1JaHydXjhoGlPGqub1/QkCeq611UURuiZDOiwjcobulQF5IgVxzkiVAgjq2z7
PONzcE3RXZCqJqFu4ly9Ron46H0rVEkkAuOyEDM6BAb1NIwMtw+HX5ONsquBrv77OaRyxm1dje/N
laN8n3V58QGLqWgCAbH6xrTXu2xYihS5GsQ6OybevSo4BLZw/ajObF7CXpqKS/w9ULfWtiaA7PeS
paQRXSuTQL37z7c1u8W4Scts1IOg4tULAqW4rovzOlw/tMlzgB1SzjSh8xgDbK+Olo9/aQFOuGaN
sYYggyxilUsARny+GNf4FSqleh+oiS6Rxr+2S4MiNmzh7+wYiY8ltaKLM2RtRRpNwQVwdRFahK44
RsG+ZN9lmm+Lf7D22DLtShf6+gcNjmmtmFeypNcG6POGSniP96WNwiUiEy0WlqTquGI9WSEKahEj
tt6HsTZE0qkZovLyB0VPngc3slKumRDXeCmTkOm+CjYVJ4C/zvk8FbJ+bsAlDE8Ga9FAS3bHLzuB
ZaJAkJ8MQE1+uTy+DhNxkCAsRwt1JdxIAGz7mrJUlFnObPUk8Rw3GugmRJrsU/iJpQ1+AOhbVZ1C
j5wYgvNPKHu+kMTV5gB/1lwIYH95qJyacNWKphFlhjyHTjGb5pACWc2O/IF5o2JooDogYnbe4HBr
lQZ4xwBPhfSpR2TeD7HOsgaG8EEMPHR8wu4vesvOcfOrp+rvGj3xKVvTZAgMZXBJB+mNY5xnVrXd
er+QM0LrAitQNnJjHzbU754d8NPHAui66qjCm7a42/HDxPKMdjEs0OvelEMY625gLrP/zu27arqD
JySLHBCngd6flKsRcSz/bcn+kNTK1j1yuW9mje+ZOodnhp2Yk2dqI7c3eM7uMljy+P2Mm9OMXHYd
W7I2B3CZ1RWjlSdfNjGaDVlBewYf8ojNHfORohey9xL9LF0zbmokRXxHVO6MK8+Ldfcy+btKcRvM
/K4mzCL7uYbfzQX50obEHh/vESnTkJj3fl4FRkr/5Q0uHadJ6ZKgQyP2GRqB28bo8gl3y4+M6GjG
JwqrdjrqmfiI08+u1ikY6u+hywcT6Cwy/yjBQHEUPIISwG5uCyVq4pdn4b4VG+w1XZWGv/Vpaze1
EgmsT2ARtOIiQJ9E1k3LdTRPCxO9Wk4UzaNEEXfizozADw4qRj2clD4WsAOeIf5jzdwcQWCu9xvT
kkoL3dZWEKL3l9IIzR9zQDtZeHiJawPG03ZswR39Gc48+bebprcqXdPMAtADiaCKYW9gt4pQKMZR
/ue6t7PH/Wkz97QEUnkhAh0j8TPshunkGbX59PBbzMcGbkbQeVlvsp+6Pu0OH8n90P9biiEaHclR
YF72I51HCqyIX3VIwNU0lEjF6/WEWildblfxrzaWMbPbROv7XaDGX07ufMoqrg7IIR5IvK0hb3lk
BioPC1BB0KFApPiTtWFhlSE6n9OSYDcDBxLurXsD2y/scoDob9ROktipGUH6PNUlXsxBzUHoUGRT
rGrQTmIXh71blf/ARy+uHPZ3FnntEhXUttRv8xLF0fJsb5Zghrqe5hAJ9IGGnIsLW6PIatUnBGjs
Cr5YQkOo+M5TMjVlNaK0OC1uzDicJVB63PSNGOsQxXG1q5jn58iBiDLFCsWgAz9HDI5hrKbZVy1q
GBpoNHHkD88X1vvEydQ7lP4L2O/knP6X4rUJi0C9aQm3YiD//LFqhetv9pfVWIrCmJgCyB+sAgK+
cvwiLh2x7TkD6XuDkbarymeTUy76PXYOJReGP3ZTeH+bjD2xl/hYWHoVvX1FafgOJJM20OxhLODB
IuuiCmwXh/iPr+DloXRr3mphxKQiBTf8/QjGiV/+L/fRDuy+WrGy/bbJ3h06uCO4V10OUnrDTTnu
hV8VVgoP8u8BD1Pd6cDV8lZ6rVakUBscPQLHLTKjRMHVHZKwLyEN2QkmYoW9jWDW5aKJ4MuzVY7W
uJZlggevhhU0dTTPNYyBdbKkGoubx8VL7Jh6KMOjNG06WJyeCgDwgqLrv3oGY3L/OcvVCCrTOnEu
KkR5/prHQyPoksIjpx3yH+iA8wTm091xF/mxnnUE/wkbOFU8DKhnzOqW2K0HlehUJCUo2GuYjRSJ
UbwZVdr/PCAPC5QdCmIqVGzTQpP9Yo5USWZzfQh+Nj6z5sEEx4IV6RtlDdt89k7X3dWCgPlp6l0V
CSPF9N39SDLSZ9kX6/zXmIvhNt4FpDaD8D7H2V2r2v1wWcoqQB/3bnyxhMCEuB0cPqDNTPSQayNE
heMBWcJgXg9xtGIzU1Qz9klwf3s1L9jC4vWgknuUmVvGFHnAnXwtnP5BW+tK+cf5RBKk2gBzExQ0
ObZdPBCzdmA7P87zWzazOoypVQps2dC176Tdl6LOYuTRedPDLtFEIPzzgGNQ7V1qsqTR0TnN7VCE
1O5AgyJMSGyOKYmMSiWeiTM+9hW0iU70T5S7URhd8jQQmqKsyDjS0TP1QB6ztTXScv4uIn4BQB4a
bOb+gT0byYEDxzX9rWJiq1U0GOnabixqGk/wp9HmmLewEoUCif4ulu/ME53BNq6BryVOkfTCslyx
Brv+G+AOwBDg97I0zPIqDFxs0MnT+T04IFv6fXwT2WFY1y23DdkU2xp2mV5JWVjKu8RVnSttd5Zm
ZLsUeWq/FWtds87QfBnC7LOwWvPFD1I3HyCz/d28MUPSEcQ8ep5ywc9DqhQa55xfhm/YDXzBF8WD
pK8+iRrfwMm/ZKs4b5Np3VFvhvWyfz2P+2X+pItUpJ2CPVZ8irj2U4cTNcJqmHF6tCtpFUDrKiiE
BXcC+uW07+WT2C2VvWBF1hN46Grj2BjmopD9hgafaNflcNdhDjuPMRAnhTMkJ1lwpf8y+7MEwrsx
Tj4nSNiIgAOZv/2urNEjIEE88FphZyngi/VSloTcf41cyoNddkvWihxM1I9FP65OW46ahDaGUJyq
l06z1Z5dSk5cXAvJmRTUdZWPfy66tmJZrnrHmQkwFc6FeXf1Aww6PqH4YZCIdUYk6Ib/oYqwyp0W
mKKlC71KYzZmcVDLpUgqAsmkVI08N3em+PeZ4AQ0r4olH4nb0De/FCK6XTe4KdHdneQW7OTtXS65
5TMmxnkhxma1qZNUizNA1j1SNiSChzXNkVb1Iaks4foUqpYRG7dfSPFwpM7Vl2wz5Ia1azam01i+
e/IhQ7M9rbM7Sivh+mrixUlFosB3Nwt4IJIRsXc2Rl6yDHT6/OXpB1xp5ZyIuAiqn5CLaQ6bhrUh
vJZmVdsdPwT8qKrASH3VLJ53fO2Jk8voNkb9mDh0XFTVv0qrAOYIC3+I/gH2Wqa1zulkJc+2WuEw
A3L6Xwf6CI2jMi6yzDgvP+Q+w4jPTWz5rIP0EQNd80gYYy02Kau1bDXZeCdH5ovdbju0M71NQ2YX
ktf5fL9VnCjqyjVravYbEkXRUtKWa1mpz2LPXMqNQv0G8hFoV5AT2V3wKMjFWXu2aMFUmHkK18pA
6aCBFcgQhm7W1F7i/FJyjjUlCQyYhBnnhAblf97qysyrrhnNq4KIhtYGNjaGFbIUn7rN0Mf0mutu
KO7McEicAmuB0zGZA4tAbM09TbXPCSK84MidbYnMdxvS/qezPDeQce5f8YCwrx7I5RHP3OO8J5PY
P26DObDJseZOuPItRVLLMeU0ksKivSKswznD6/NJMy3APSwuisErQ4aQ3KPuQcBO1xOwgX10x+1Q
1IB5W8qmJTCSUogr8ITrkxomdbvUoNHIeX+ZfahEdpOKNptzRPwi9oxERmqLHbDaMZ1xJA1G4kU8
pLZCUsYgL56JsBIj8/d54usTpBjfQ6QJZP/AKtdGKlkf3NJm3iKuAET1SuruuFI0CvsfgTY2OfDm
g7N+UFrvhSBqvpIiDnlkw1AppwpFvmJM8ctNKdcnKI2RhEV7Q6D81AuSIBtdErfg9YW47X3w65QB
7Dvqpijlr22ocFOvM39zD9QpN/Xz0jQKuQwUHvhP0HqKcyfhqZ81HDWm8X0tb5RFmDSxDELdZogr
61u49i1av2S5Em4NaSbNytmD9E+u212qFiDPDYt2Lh8OMVpoPayDvPzzM3yWul504qp+ODAzPHCD
OxyM/TsjV2bOKHw9G8TFT5McZjQkv8tlKB/TQWTt+5WIwf7NAG5FXR5XnnEhe+Vm1Flpn8S1mTUJ
CcMUOWnuxb/niQ3B7Hs8fWhcFx69YG5BJZx39Qm64k7Skar35838HNrLLWM/XoPNpsnMiQPXZEn2
yKWtfv7aNi2Orj6Xw2aResE8TbudNY64DqNWaEjLRdMlcQmWcp+DGiRB5TYErgirlcTEz5CJ7Tet
snxdkxq/fy7L6xzzFxAQE172aKIoizsEKGu2EOjM5UTwEU9Nqs9CbqAGRAyLICpakQg6waKf8BgF
6peTcs6KHOgnGAXhcfBtrk2HLRQNFOPOe14w8+VB/CsLgZuqeB3pFpIkX24eq2WwSDU1uFblm4Hu
L/fDkEYAAHgrRYfeecyoi1cLNVb0fZaLcOthwr9cj+bhOGCxmeJpByQw9vJFVy06vR3OzhR6dCWp
p2mkSS/+5Q+4grkJnEyq91q+dIyS/0cVpixVF4KTvs6B0JCd1XmeqrkW7c6kiB3Q1RS7s6xp6i6S
9WsLkPygetOwqynQkHclxshYz2JgFy51YRNw44d1ul4mZYg/9JAdKLGZ7Su7AS9y+lAPmewPaz9l
vHt9Itz9Ll0kpkCcfw4vanJaCOzPAVlGNqcyL1Hcu18RPxfo9CX6Od+eAwqro6YC+Zr2m/gSlsTx
ZRtlEhWDdqv/ipwMT7oqV49RpWvFAVlaoA2kJnmxtoPWiDT31Q1BYtvWjAHKbEfuVeez5y0c/tzH
+DPFvDsosiamIups4QnNvgcj9Ybzhcr7LT6UW0oNXWQA4un8vvTHrS5rNj5zHAU6Bcz7IefjH0ib
sGYwm2n8NF/Sedc8h/UInpS6yXsctOJOtfNQijrzBQS1UKHxPEOk75OzJy9UgdxdSV8AiXrQ0yQy
nLk7lcRNxKnc/VIAUmpfdDMBDtmjwmQQrFx2uy0ybzMGo3GeOVlNTmCXn2FkwQscaylEGJ6WnQUT
IcALI6xDM6g/Yz3c3WvxGucO1gg+t2n6arNhAP56LzsYu198cmY4UAuCe6VlKo4HG4Z1g2B2iXHE
Q0H3l0abrUSq4s8312a8gldkraPmnAwNPQgU6EsIFSSRqqZqOurncd4zxYVOsYZWrtkxTCruWWQI
R1iWweVH6ur36KULnhdMYhtws/RBnWkFT0w+pj7yaUQbcLnyOEu7GQfAtHpFVgY8jNwGdUbJ5IOR
BgMR2doVW8cn0a9u7L8tvD2lhpDtmip2PUDIlrfqSw8HiLZQrclxPCyanHsjVDQtju8/J4HWDP+A
PqsLMgGNWrf9JpDB2CM3HEamw4O5gQ7ff1MskhhKKFL++UO2iuX9TClu69MLmJ4WVPpZ10y8wndC
JcWnX1aPTSs7ny8j5s3pLzDHCpt5JnYfcgYcmFMkeHmB5N4CBVk0q7vIFxcM8GVBMdXqLxaoNLsp
ymC5rvM3zleiQIUAQDtfnuRUTNW5lVBpN3u56uLVX3ZBsz/49iaICAWF+jtQkJpF0T5+Hy+6uGqW
JewvrTLpnrHRAZkB9tJ01gGbAERktUaEB8AodC9IuIikOKZHcLw+3Cw09V/D6sswJapNW3Qlyci1
nnomUlCuJPdWMOJC+ScK02oWlDHiahyq1lozJUVOtFH8gGxe09Du3pz6q99mUvD6s/1Q1nypSQ9s
byyCO8MS8FTBqSddOO628HIXfJapHuJgVcUxBu3phmxzOdWg+jBTXWouyK6KXLo1NaCa27SMP3sy
BwUHYdtCkm4LF5l+r5G5ukvmRiAc9IL9MpoMalE8Mx2SVOydB6Jz5g+z2tc+KZQMXU+T/kYMIFPV
0t7nrBw8n+PXNLn2Wk8GUKkvELMNO0ipe9H4iZjFKjOFtSFk1SYXKOm9fBg/Id9nnLjOqTnu8XWT
j3rplDpIkzxhrfWcKUQwpgqvcSu9e8JPVRXBWvAtu2lqTJ54XORt2nthOlFOv7xnOWL3ZnkYL4rg
mT57KF2hwyLjf6Hmn5g2oF3JAgAZ/eOO+lYSmURv3Ka99VcMUaPPXsAJpm2m8ycFhlJJacKYj8ce
MjzSeGmFeEb+A4u5WzsAIze9ESLIUCnxWdsVGCJpuDAW519NzWZIjTTeKRG1g/AwoWDzvyXMnOGp
MjqUvMdrOELdjCtYJCjVOneQBk/+DT3d+33wkKJAERzOeGy3wMyeSI9lHg/OD//oLolWP1Dja86c
BN2EXlu9O1BFCpUUeI7hXx2vMzoac9HL36KViCuqEJI/ie76Np+uVomWuasY8TPCHlmNfqV3O2Fi
Xm8vPnOfZ1woEwf9B1Q5T9u91FhHdnmr/rDlRTvJLK9cd5vla1WeOtNkiZFK1NzE8YAoa1Vpf5Ya
R6xnPsxbYTHkqDHJ2aLkj+mqn1Ml5GCIr9DW69Fl8K49gZgITP3020+PsTyBn3mgD1dqUozlC0nM
XC0pVabnMsdvrGoKHchq7E7AwVjvMx0Ic/OXCBn+8is38ZAtDt6U7IBJO88PUfzQdFrVH0PuVpUO
kyqRlCQUUI0s6f9L7JNotVcESjJoIq57svIdiMmYb6I6gq4SdZfsdEe1VreEYlWGREG1o6E+/FIh
VK1yCWRL4BJXC72yswkt/F14x+BTUQnaa9K+q6mr/UiMQdwryVcmBkMol+HxR7TVTwOUmOPCsgXP
/mdVZ7AWsLbSusIalNbVwA3sk4YnGZ9fvlxp4KHuBqXofYlbA80r+gEWMZJEMh2JuMa/qOvWNo3D
4Sp/Pnsa432o6Tpn476f/Njh3T7lsZCd1dG5Yp4GGhb+a4u9kzDW1nzO5hiMPy6sBEf5Y8+RnCd2
X604XejOIRNCkuV3JrfZpEX2lefq2TQwStfWl8oIzgETyqsmcPqVe3N3QLuwqOe+pQFCgjIAvRZM
+DW1DLPN27C2UJvasONAc2I6d/hVy4IrZKqoqsNCL5YznWiDdSR8mZhJoN5LhR1INRgoRnK7ExEp
vr4WvDwgDwMOaGTC5oVWMgLt9cidOBMT/3Cr2ieso1lVVq7e/jUeJiLSGwqcwKxi+F1gR/xHU/V9
CQ8eGZhCrUykQ33FzFRnmL4TICoWE1k2VshritBOAmewg4l31mo/sGbxQcPmYduLJ6MXXVfNTKO4
zquVFps5dNX4J9aqS+g2wFEK+fjJ4j6A6a+dEsOtY3VMkqWXAYCl5cybFnoEBPP4Hibb4/BUc7G7
02au8R5sEWuu7RA19yJ+EOTRCuqxomT5ijFthlOFvRse2iwCj4AX15xZFlu472OYlmVUiLDf0RiD
aoTb6NO1RKM+6IcOX7opli9ypJdlWxCJbSTL6inLaJ/zQ5/7weP3y60aE0ki5pmhmfi34+PqWOVB
khjS7d/j0IrzdlcH1CMYcWhKzoU3ijc9UaP0irEZcWUO9yYPPCDg5zsWtP7cdHaaCKvgW/y/Zy56
5YwzPNpzZNiH0xwM0gN+Sq+U6Ho5AZeezKqSYcImFIwZfJ5NQQ9pwTeh8xjhlynowj/WOyvSzbeU
GjvqFPAyAv8Bb6fGhEjcRSiwCF0NtAIqXt1ZXnJJ08MCzqjgcfLDiBXUTpgTWbAHLQMVBJJ/vfCJ
Znh1tRB8kjI+VA92Uy3zbHppJ04pqwreRoMVwOtBmjGEiZBjvyKL6OYDnNiEi8XHFkMvsgyl9Il9
DXCAhcjQrn/9ZpbGMj92wqYn5t82/WQ2NdG4E/sjBJOCLnCdTJL3XEu10QksBT3iTwF5hddWp71i
aVaLuOoXbajvVpY1/OUcEHendK6QD7ngknuGO1R84GUjRajEOQcErGkCxJVlWss4KNtSYj5xrErY
AwXOtk4Sb7vjePxZ8A/RVQMBuvcWrrLU/WWhJD12S8XDdx+rbJwLWUB98ZSrBTo4ybJAdfN5f+QY
ToBQR1BYAmd8n3GxT0yYiKDNd8GiKK6kwCYkCkPHVbS9BWpcxyjgYEMuO2oumz+ZimR6uI6Bl0jP
6jeE+Y/Enr6ZKfp7pLgX64r24Fje3DcnCkU877t37hKDgnAkS/1eN2YR2QbbOl59jzsM0LuzCgc8
k+tRLclFacik6Gx40mkYtzB7+Gh41+4ReCR3EBWXG0xwaw1SmbFvJvXoWAP4uSHY6qf9gtEFFpWE
gXwjYo2zOK5X2im1exeUQ0ouZnDYsWjR8zJZvqBz3OWIQy+yQ2PlgYRL7meelI1GPwKwW1uwgpqb
hy3bD4BIaSwa7oc5s0duKNlfjdjTKkFh0Ye0wuKlEV5PkbVvYc6GDZw5UzSIMV+wuDjjhrpXyQyN
hUOKphxAkMi5ZWdJHia7bo40wZjCFoOP+X7LLlTNq/ylwA3KDrKXE2QjD+JRFbqgu5NIKHRl6hj5
4ZrkO9a36QXCP6E8fXuj1ThY9Ax3PmE9b1aov/q5vyIOmcL2DPfAWM29zcKcbcqqvyVkRG7fB6/b
qilq7x0ZWqnYZQsr5i40l3eeLU2l6xw2HXbVv/Oxbf3fEoR0Rho5vlkuVxCEP0bBsM9pbfpv+g54
aglp9QH/vTkItlHTuwHfXFDR9DGWFlFJerXduy4bbBd9+HwgRtj2q9kbA9IwPqHGLBkmKiORdWgu
s5oITUq3JpyI6SRH/5/f/mS8DKS+6xxii87NaTJ2xS1SwcEwLZGBzvXE5Z3LYcYZ7rxE8qiY8nDg
3sPC61SsLbYi3TqebESYeLXoOAiJBWi0m6KlBVyVVktqcjSCPNU/nRAI0KAk0McYd57pztlI1J9K
g0to8bG4MUXwUScb5kPzl3WnqB/yWgO5xS7XhI6Mxy4AzlN3y5FtXNayyD/ENlJdGGSPsCyTfONa
HCqBJSO4cZmutUM+g1xfVHukls7On3ZPflgz2/Fnqq8PWH9PGxfAOiOE8g/hJgOn9YgNw+7teGwD
zRd3zXUZi0TuSSDRYIajDajAqTs7uGAD7fuXnz4EShh6ugEgA6Fg0+lqgHQFJzAh3cvLlN+dwcLh
bzCz01fcIZj065w1MJLPkUJ9l2nircoH2jhFe1tJLrvzSuus3LLlYG2LoF2rlurHZU9ukymmqKBg
0aZdyam1UX5GHmD5T3aFzL4kAKt0/hIaGk1mxVbuEv9+3TyFSPdlcwTd4nNF2VmyI7Lj1D0AeDsO
gRgWg6VkDKNSX7XHSSUDUCCGuMFXb2nI7WcaK3XaqqUJ0xX7foS5T73BU10X/ZHXtwcq6UEmQCKp
SkcSVbDfoo9yLvxjV96FVejAE0Y/4Zeouqc//5dCVUQIplOhTOMvm+Rveexaea1rDBEcX5kaTMFy
VKrWqcLonuuWSySMHwAOm+rECPpbLXdp3BsQP36hIllg5f3jF1f5ulePAap8/Ir8lHlW9ZlB56hH
Dw/l3TDAhlYQ/c+NpOEjj6uB8sEbLD4uziIhUqVwPQEJtXZAXiUzGFAnjVjvIG80f+69699mxHY/
5WSLQ64JhXiSnQrjZxoglIDzBmgHVr8o67Dl8Xx4fhPUrrCodl7NnKDP/BAnxWgSHwI2CwMeRHDV
wiaovD+N5+adbjKw7SWKeGhdYaH6+xWwAjbGYg6eRweHidfXgdVsN60khqzuHIZVmrQf4xQE3SgK
IJJwYDGmdlvG1hC8GzXzRx+PB6UlKknqDuqbCjq9Rij/OtdM/0YsfvncGTSf35RM5yZ/VqepH5tI
9QWWPnIAFUtxyAZWl6ohChQLt0XIMe3F3JCrIf2YAc19NEGk6yGI3Ie4+r/w/kuQUcrRglFdMj4u
mkI5G9dteYUdufF4Wj0LCejlNL/XdVcYTROBYENqN/YF6DUfkx6K3HekkHX0qEDhDS3kK3S2+UFs
mS1A1rIi3kvNXj2c40GMciy4t/mNINSbRs21BCXF6xPkkNC4wsNzTbMYfAzmd0nRvqKt3y8cD1U3
Gi0dguz1l0LSloLE8AgNodFWrC8F72IbMyZvms6PKr88VDzB8ua7Ur6lZ0icYRa3I7xvPCoUYLC7
+n/V9hXHBY3KR1iKloKapTIhEWLVJ+jZnmanvULCl0IgE+47Gg9FJkJB8J52wwciPeFYiCmxBXIf
hCW5+V3pFdLfzy9zioGnwYUElvnS3XWC00UDdnuuzGmiPnr2vTK1fsQRt4JyGIF5tBKam6ftiWXm
tcx1IqSMXNbCErsrdoeSqkzv/Ubx6xbvm0aqvOnL9ZUxhf7hPEnHpTFrTBYZTC/Wpbl2t5HkBAp0
ks1z2qZwc3eOJOzSrO4zDU9tMDYk+13/nH7mhfqgBnxbx1R84Khn1QdUXT81DZRjIl/I2JP0wi/D
JnF+lBRVo98SEdGXgbIBSIvm9IEeGzM+fTE1G5VaH2TzJvg7buW8rOdzYQO+VFrNgY2wqbCaYcBJ
ptUhr5mawhzDhucbsYz5hdI3TY14vmQsG/bgoEL18EIhHgCX3jw5UIMsvuzsQ1rBZ1L0NQMyJtt6
E26gpIwkWHLKLmn5oop+nDSK/gitGaKIpbv+/kczXXo5fI6Z8VEccb4LOm769cwxHvfnGYV8n/Vd
FB9tsGfBWVZbSlGlNhFQJcEp+FQvLT9EjtHlc4lys2RdwFBuFPKR8kELcIvCYecvELg5CvE1MKsi
qaytbfRc/ndKR/M0/DQReLDIyRQpHNKgN1bCqnI/mVnPSVIUMUgLKnfbyBWo7nR43O4ncPQdqEDF
0Wq0s3iz09dCBPiDDf7MXF8qJFxST9RQRJP2crhK5tPO/EaESFzYNOBAExblS+vJLrzZTsLBBL+H
kXpoda3ejcEyD96l7vWQquCjY4I9A8gq7goXGr34JVz/mIIprG109wtwoUWpvBm1TLIXkp7lJUJD
GIdjyeIWucOmhJdwXo9oxXxGOzi1IV+0JF3wpo8VKKwlXnoLcaR7AEV9gmz+h2bI/RlCn3/pmx3u
uAF5dScCKYdIYK+6IZA5vpOiqDh0Tw/vvZVmSFWa/6YcFKpGapy60hDIb3SwYs9SCnp25cmIy18T
fGmQzs8az19AvMqJ/o8wGjiN0sjHDRucLxQgdfffwXBU4GkIyaR22BcK4TF7ENBKQacN3OXxKtxc
c3+Dlm3/5GnndmwGzYSf4Qcj7nz2xGcy57a/05RsMy5eoljAIuofr7pbPAt1lj+1e+GRyaeHNykB
kfrpO1LGY0RrA6uluYbOrrWQE/cR6NnnVV4W+T90FUnKGauw8nk9jBGSpwoaicvEb8YlQEYmSSkq
awNp5nXdpssqyWQbC7t6v0LJPCzzI7jC6o35WWbRk7t9LtPDRPCdeYduiO5uxOaO38SWjtE9nzdp
HYrcfT8wxR99wy+gUf60+wPjdUeX4jNE8OM81Xht3G+QgeIvMuRFYIJXxWxf7LxSbgSo+Zs0F2h7
DeamDsxDE5t6/H8eLYgVfEbe+n2EA1DpeDa6Ww1+mNni1uzV+e3a124eQ5FAdTUR9piMQ4WllIx5
zXu6orsD+fGt9O/+Nvw5rLoClEjYbhPmwOOw3oTlHY9tNZyCv8J9K58kzKlhUbAeohw+rff74PGa
DLDeuGhngh26epKLFhzgr2ALQGwIuL0E4OL3Su53Cs1aAHToEllx8JMCwdeHtgIJq1hJNi6eA9ou
ipV/doslPXhl51Yju8eX0HK75kSiWYX/KNfRZeRYSUP3jJVLbLX0YHQDTQU+2Z3/ZxlEp9BzivDu
82Pko+g7XY05PxKUrKzzkNFivwkSWRvsNbqPNEoxO6HEwG0TbI2yPXJm8GB9WMH5V9dIunYwJYCp
ey3MQFfrmDg+jeT6WrQ8G+oqFpNCWqCNIG3N/AZgR//HmMNn9chKw9K/OWhQf2FDN/jTXBbERAdM
Kd6SHzYXRuPi1VlnU7KSSgAIxPCGtwLgLeLBp4zQEgbzlfvNLOat5eeO1WNqTuIUB3BlKROd0mhV
4AGz4RsxDK1kHEgc489UydZ35d2qFPj8dCuyrdS3dR0ThMoNgqVJDkQfY1pU38TkNzNfwLetziNo
fWAwqHDizI1pyaHo0Pg8X56fNPZuGzcwgO8a2dvltt5qI1C5EhWBZJZGdERs9jw+7MxY1rAlrRSE
WBkWcFPrNzxGew4uEoWiyr3Eg9BursGNVHJfQLNZm8uZUKv+ppmof1BrdV7boYfWXHwkw0wKc6bR
MFo1xuG9B2LYgpHOjmSsmFUSo1L67ERTAFjy5wX5YMmVym62BYcsRWuF8k/2sHHRs/hXyo6hqQ/h
VQ6YznH/JzQc+uzB1rkfim1F/bOO5El0iPG5J9RYAdvaJAqACMuGAAgrfdOtf3TsebtkjHRo12H8
HMBs4AvCe80Rw5A9npTe/VUtZnV4oEFLGUKkBtoLtmaTqGHUe4wYEePcVFtajkodADS8rrdlss1r
nPg/vAsK3ArIaiwh++fbTZJtVi3DXY2X05fkW3Vpyk5KVGbyjJBPkWICyHnMVIy0BSSDUIODy3Tz
tHZb1xB9D1/EPIQBfCKATVIYWYxq09zauCorDQqsLf3hJjhgUsDz2VstuRJHmg5titzhcOdw9KPn
pGaF7gl3TNkpiaZI28Q+qboR2WqncKBBwSSM7/JfpjBaztEV7W2gvULVunO3pWo5D+epD+Jyrypk
dScwyUdeKNDRv1HpRdAimCZKsLWJ449Qy2rFSSUd2urxvDGTjuqE4AlLx6BDqKtnkqvArBZaNhxK
wM0tDy7AOBIZ5oOWIj3D8SUjAj5jgZSH2dHrXcwUAMOOji+aUoGv/bbHcDvP5ofdSrZpFF8qxn8X
pac74SEKEepy7r85yB59dDfGgOsYkNqsRihhQQEToCjIlT4ibN5chGfqnrgDcsg3t4ujiKi+cMj4
67ttR2J3Z9f/6SIYhLl7sOdID7ARPqwgKXOOUGqq6tSQ75f9WoxTgyn4yRH4rf4vdrvbiHA1F7Y+
OUCWSLPcIfPuUSlqlwm/0O881LFlxwF/gxhb7pT2qo2gO3EYA9nhzIqMPv9UeqJLx3taQS5Pr80z
B5KqH2YldF8PRWTo9tMdbaSq++VHNiPM+H84T2GgfiQQKDnWU8k/Bn6caMmc17JC2vS2qfWoZQfr
KeIUCkxGrRyxKG11O3OdhLjNqYqwS1EqJYKCN++hW0bXdzO+LwoEcRRID5TtpTk8Aoh84epQgRJQ
eafxTUoayYtKItP4HbsTkIodG3CUt7jlwPLHwgHW9nssiC/0SQc5ZF8HAy4bt54F2GJrrMM8QoIo
StvrdNTV52LaSFfArPuB91zOSH/qmSej4WCmOgG/+Py3XtJSXvxQY6pcp+RkneK4DQdK3n+eNnNz
oxCdDFQ8mfSgLJybJlBGZsusqeSY8AAlpVcF0wCTXtnkRh6yNUExWAabXLK7FSAcbLLshEDrQz99
Hah6wbjwQTJ6frvUt/12zL7+JvzavuyX+hbGJbOCQR305EKk3qH2ZOmRxV1NPEvOBf3S5vKPRMSd
wxGgMaKf2EcgMj3O2O9zbW3jxKLi67G97PDmS6G5EvNE1qDnbR4klWLgggoqZNWlpJP0cxcMpGsS
FoiK/gX174gnMmQamWCdSjve7n1lu4Ca5WomRk485WmgOBhD7emt17TChGyTAYqjsDM0+LuHfXK7
auu408mvJudysHkMP9XBMtsJEyccBksPl49wBYCDsKGIZKxLSIYEH1b9nz/rDt7nOPwarYA/wtxi
3GpHE6VgTAOFLyq25M4+sqldb/Rtm9Ulp4/64oTrvyLp458j3u5ZMigPSN/WSzEPSpwEItFYkY5C
mlbUdW6vqmyU8bUDP6nPlR4Jy8TJToNuMmSVx8yUYYsE01QhVTbLNJ5oGH3rOLjHdF9UfK1fy9Dn
xNnfYFqP8yGybISodgFUIvRvD/XKTKd7yq8u7/B97PwxZectMGxwOne01fuwl/ZeTI/ijaAs5MRT
6O/tSdqo0zPD0KwgtOuBWdN4z+ZHjAYiJmnV8o/ehqy/3nW/GKBuZgVs/SPvflsV8m5XUq/vLVcV
cjtz7gVJZHYZwmPibnxF7QgD8Z5sYlrNrkkLFymY/KSpJ5nvOT/351qb5V1wMJgZa3uqQcTmXu7g
LbxqkD0GuU/WsI5aslddycNL6j8sEHGEusNGscy61YxGqRUODSvnoPNFeunxE3w5QeM/cUPD20m2
jii00aCZvRIggSg9kG9YBVRMEtb00iQ2rxMZa7zVOemMSAayQoF3yjgtHf/3Njh3UWeKn/aI+dDA
+LeB15tuTWh//+iBCDtA1QwFyHbIlKts5E1XJxkNhTChvxMOFRKhXJWd2sPRJz9bEZb2T9t/VQo8
kUVGKgNJDoTUznpr4FCIbtf+Dzn+1IBFFY4gzmmjosb0t907TNrvXLjZ+L3pqrvgrlEjLl56s2Fr
cQr7uQ4dezmR1383HesBujvZfbIGNn25tjbpy7C0njmTwnolm7vl95qWaj1dyCLk3TA25JrMMg3w
lOUF7rrHHZpfJWAhJX/94zrmKGxYN/IJwODQSAuuuhpDijGWvV7l08TjtqBKL0/0xmqjs+rCgVgR
FSj3kme5vTgjuEhi1/vmEw7TptZ5fULEEru8hgNqJY6Kj5ntfE1/15pDnC9FEpZ2BmZ+2qj/H2a3
tarvOOJFrsD9fePAFpIU+aYOuEj3lBJHso73liR3ur0Isw9rp++4aurboX8KIdOr79Rnleeu9g+L
fqpYQxN3q7ftfEm4ZXl+SMb9fsvr5ABfEI9lFRdnnbWMFl8bKGbfPXR1C7kiomxsZjdmGzpheOPL
w+4czd3vcRwtAGECjAFDzngH0cnjRFB48AOLbuNVltSgNWyJbSScpk2Up77mp+z9gjK4qwcnZVjH
8wvteQ9iObI3K1YGFLJ9buevOxD7zqYxQZguwUGMgxzvzVlQeChCjJZxIj9YuVQgxYZYBWiefCOz
5FPZS0UId/2bT0YJA6RWSQtmVwiOvRDlyBHX693Qy5aL9pxKWj/9x5su1xpNGOcUIuU5XJVa+WSs
ox4oLT5nac4Bv7mZ12aH7R0yk3AdXmmox/uj2dDKCvHckzYdsvqKnSwtQ16DK0KxAMfVq5TZIs1T
81PC5Ex1y1svzbFrlvh2fjA83fhLfiAjroWMh4p8gnXffR1AAdkYjWGv0lFUnEh1bym2kEL4/Cf2
g+JrTu1OXsoGzPuSG2SbWg2nhO91x4wMlP0V9IkxinLhD/LmHvPlSZYuO7dvNVF4XqYdoFlJcRoo
JXswrreqXCqrRR6iQe36dE/oBME/l6iC0CCpD+9ZNBnggYQguZB4JgGf3oz9zC/L1WUd7SX6QKut
fRD9I+KeUKjapp6ssbHSbNx8jGoEVbNag9/71UJT/H2ullY03tKeLLjIOyZaUmvnH4jBH692wzoT
u1bO3qXW9zISUVBPoWdyEayYLxOznEn7f0w9IL5FK+c5HEmVRx1+DR/WTOpn86S9biZHfXD9vFlX
Hzuef7b9yw9WzJvCKt68TK/L4yIpHu8alFC5svIO0HYtwvKCZVQYeRNJkrQLJoAOyDIVLOb5m4D4
KkKYd7x83EsBGLvsy/PPkpICKIgqA75c/0c/Z3BLNS/5pMHHmyrtqkFl0jK7CXPtE07AfqYIkoAx
6Ndu8PII0ryI05b4U6eTOxXQAZML59ZMFMZmGi+eLqHzaLpGoApkrKW+O9O3jJte3Hn8CHmNVUxY
OsBJ5QPSt2urAGFlMjiD3/akasM2zTa06wS2L1Um56iBriCwVUZSDA5hs7wWurHAoZUT5JGq06GI
9dMShmyA+amGmgfcCFEwmcPbd5v+QQ2e376hAyMvsUlKEVDmZUZdl2Cxqx2n2GDjsZKUrEUY2UNR
OzZ3YCjBUfvb/22GTHNS30ifm0EY3d5dVVynkSQ43Q+ncZZLgrZq7KrBhg+wdLlJnPJSdIxWEGcO
zZKw0FqqqN+sAiF0uv7YsFP5JzQvyCfBXpdJkpl8PuFHkZP1OP9xHroQrB2eqlPezqOMktS9ZYOW
EkVL33wGqiMwZqLs7x3+z816PMgoYq+nQ7cF2HRAkats3pHUpCyaa2bDV6RDTm6Jj3Lic98eNLXM
9RRL62yuKjESACdZdt2oJsJZqoOBklhuuPhrrTDCWlFsPCgreQ3/0sC+9V1UU6FaBnYkMihWhTRI
olSVyL2P12JMiE+aEB5wgZybLK+iGI5a9HRFMRsTI7Yv+7XQ0X2NFa2+SqBgDqPcnU/1IRwIJQaZ
p3KnfhUkw0FvWZSBRAX1t8f91njLxnwE1LbZR7tQMnrgu0IUn6Kzt4lXzIvuHU6m5ospQNcU+jxp
XmRmlM6XDUCaEM+xCygouQqt6gwn7I20LOMRu0UWQnwshrA+CF7KxG41b5FlbMuxy9mJdG8BmR+l
NXWjgsE8PvyY3u9nLi82G3WrdTCMNnNACHIstt/qyKwgb2C0c74u7uCWjXPWn9LpC9ypXz2zHAWZ
Gff2mhuTA2Si1pV/+q5peQ9NiRJqd+Frvkk7Lqvk8ky+w3aY+MdZxxMklAjmp/gGmuVauY7y9too
3gTpvR97JEmXGORXxNTgnyyH1cxECpbai6k5GiglQLQI8BxbyocD1ODIyldx2BZKtyX9x2SZXjrl
kgo3nFpKCQqJ8aNFp1L49lvV2/yOnS7Z6t0abgsF0uU/nbLE6WS2gWXzPPzBiSzLxaDDTnwGd0JP
aBCqzz9vQ546kTQoamwuYkMbrOjlVNVQaYEeoTSgUKqS1/BQ8MzdP6fBFzHTlb9yn4u62Kw17rj+
tKxkUBymIdb4P1fMhZBFjB9cB3PuV/jvjjTaYAzogbESCGaLrh/nfG/TSM0TrjWQ6ZAqMjPXMz5A
kssfybHGb6rv2F62vJaGJqFOf+IRYe2Kxp+ZKvXOrozrRAzVmrDNrJTBd6MD5ua00T7RsCKFWkJT
Ap19fKI6AcoUbqPiRViKJCnrrxzqx/xpWA/WLiXFfEdRGPreNTas4UY2aYPIbSSgxm4QGY3gfVJf
0RY+ItGL8ZWaZflN8YCpg/4lT23Fs9jRQGjLooZ0/VyrgaBBAKd+eyGcjWlV5cjewKy3gaWz/c8p
F5eroqTqTuwU5S/H7imdGCxpCVjwSoXUUW+vRz6ApsaS/DXu5jOG/Z0Skdh/+vxD7NrUkq44RSm7
fn+x1pu8EoQOSc8Pt+asJ2Uj23KH/qK7wwN3zKv5Wkjyfdk6aYqwPQnmEmkbLpBZB9DKUJWxH1OT
dXrI1RIrd3+XHAJgGLbJt3LeDT7KLmQARE+HzRhkdK03TwQbKVURvUKlykSkIbZjOeEBgOCCofjs
7elg7k7VeDe1j9PNsA1qgrmnSudB3ICosgMQVMkBJna9k6lNOvQi9bbRylbrMIseE8o0Z1HvEZu6
4iJ2gt9rRtwqpqxoc6eCS4sh0cHhJOHv+lfPVSjbE/p6bVrsF/4cbvIOCr9kuOuHc209RAwD4BKB
Scwy4qqBaB9FsqJj+A6uy/dZcT6vHoEcWpDrJKE0a5fTee0XQ9VynRn/ZQzD/dOwblfH+VHItSHC
y755qZQMTcQmR+/yGzO985o7K+B5ansJgWMbMBYx0h7GDML1j+cs471aoPUWNp5rG9UHTaaQ3j3p
84iyFr93y52FhWiANhzDPVFmEQvptcohtCZ+exW3FNvLm6MYx9adITSMkx/bw9bOk8wIFLkMsxRp
B7xjyDze6l/fkXcD+Ui+13eR0M6MA37E1K29iIRX7lHHwyOeZiLuYULYXrVJRyKXSkYe6oH1VsXw
TBYg9aMEnVFItSBV7ME2h6HxEJiNNt6s19htszH/VaQOPZyJJnWmfHGjngI0SKM8wxSl3nvO0mBI
OtRMiZ/K48dh8zu4ovylCls7TRhjEsZfD5piG7PmTPxboeU0+xuQNEFIiXwMdgSKEWJK0pCP7MBI
SIdn9ko2U4lR/1cAOTqnjRVl8Z8J8uq8D/OGqwouJFmH0hnI27DGerucx1flhsdbRjwASB+VOU7E
SrjDy0N9P26+FEHE5/BKBdrFfZhrPlMYeUZRxcy1BBkPquS4WtGhl4wKApIhkFUT7TgdhR8HT+xM
GbNvaePQosX0LcwdPoYl3Kz8s/vLZz6/ZYFjmpQ/hwuARB3DKH6zhkh1ATLKQXZhP+wo0i6sAgq9
dBuw9LkqqrHMN21cTqUW/ZN0Jnt6I/MLaFwhdWxsQ/qtQUJcPyXkexNnm2rsDzX3cEByrbYsgQwU
wFFzmkp2a2TuSkZ1a/U8r06Anz4HMH9v+ERqb1uwDOaryzM3/IOi+hMN3DLBiJLtPz3RFPi6GyQY
kW9IDDoApv6Ofk5tS4JQ9mGhxyf7vo5v50UbEDfZm1xnZqNzDjY8ga4NKn1VBCUV0gg57HMN2fzz
bMUFxQaicfwn90Jdbd9FFBAGOQlGKBGxeiHtkKtQFFDNva+ENOc9jS0JWKs3onTWuVq+Ti7HH2sE
jofryafmazv5WHpF2gAfdFQo9zJnU/qV/1mKXAh/C0MnAHcCLiMOSVG19vpS9rEA/y6uxBhGP3Mi
XXsmCr7HXwT0Vq2XvwexmnXdAmLuSbADJTtnBLZkzxTp9YHbbQBtc+OPjzvhB8IXfUaqpS7mFWhH
RuoIv3LzZjn9L9A9jcDqQCyLOoUF/6/4dzzopIBItFRc22QYjjYECY/FFi5qeipgdelB6BG+3S+9
k+32oglmFZ0g9YKaqxU2EWNHMsfIATD035bLDN6cAHTY11kScYse7hC9JOAe43Dew/VMfGLI3JMv
ZnNvPiHLlQLh1zgQfO53Z9r4UQXMBxugy2hsbR+n9gotQxRll+GyUthIRMnNXIHPUpOetXoBrLwP
If8UUabA6xYJhEV1xzIKVSuV1rYQ8b31J8wP+aBrArsm4k+Tpu7lbUfzP1nh1l/E8GcZd+afw7gz
dS0gCLX8JRJ8b72oY6xHLMJc/30mH3yiYdUaDYNRpFA5ZyWcZYAjPsDPxkKHkzi5ruFwm87YC6D3
buRhkrEoeJZkEWHk1Ly5eL3nZmNlPY+m3n3U2uncymNf3wugrLnYNufzF7NcS76ydBdyMa74WhGH
Ynl6EKqOT6iHBioO3ERWGiBg5PAz5asm+krux6+ZDJ6uS5cSSMeqDQYQHAtDtiVXwVDOAmRxf/9f
vntPny4p95kEOxTYVhiPGguhVsktFdYyV5JVkj1ETpMC6rDMC39SW4C35KW50lKRdUWlB4fe+VXX
XrSOtAGK14kuLpEQx82RD1N/vSIaCCEcRxYyndw6kxSsq2ihLugKgxsw/ZWNCRMg4I1EIOxsEBBX
RapCRX8tOne8Z0nnywq6FFGBsv0GwYO/Axvhe5B9jeZf0UjkzrqAUlWUhusONmFPdbuh+bYtRyDq
kGGgdlW4Yqqtox5qjl6sSo71HpOzqBv6lHCbDDrR3oIYmzkeF6w+0UQUNqxvMz8Bpw/992DPpNmX
laZGAjBClRwcrUuOuIUH+CDEm8NOqDoJWPCwvphG5CAFuGZ8DmqpmOOSri/L70IWRu3Tnl+1JfTG
i3i6cRWCxJBCLMDZ9ywS5bvU6Kr7nqtSxV3w7uReOnpgSlKITaNQNrCv0FpG+nh/LqqWmPCpiU21
hLvUJZXYGQdBZeoE4Se11SVD1a6AEzSWLBthtMOxpsPQEcm8L9JPdOwB+hslv5hHj//UoKPs9xg6
DY3xzUDrgJxQp8OCGKteOutAoMsqKEn/0ZVdzyo5Tzg4k2Nvo6KLUXZROR2Z7W3aJZy6h+WB+ms3
bU97ytKx6GTMMdIqJm7kw7JRhoFLvv75d3ErV+vxaLUpIH4bwhajGy3AZKdBjX/EQJzs61Q0q49D
Fwga+/yfOmViVp+DIJwy5H2ZW0UPbd67w/s2gQrMMCFeZjI9kdO9F3PvMq7GP9JihVLU/WMm0IpR
A0otJCHJmcY9j91OrxuZ86Za/hTTjHYm9l7DDWc/ydEHcVt9Xucky+GEg0Ms6JEJrBWxkRNQiyoc
zsdVcFHUWgx2B4zBJ7JBvHExB5eroSPn6FLC4cUkkPTTZv5KBY1F3wOxt+4gK+o+q+Lo0reyxBIf
b0h5qc4zot5KJNzZkZgawtutuN1WDQ9plDcRRuJ/6gLxwqdGrR+m96Cc/2YiQzoPrY/QcP7Bxmvd
ojBZhKdD5GvVVDqBaZMFIrqp9Vcn5z5siKUMbiKmyi8udKhngTKv6WuKmZP4HtyukQ86611rh7Xk
rQuTtB4oCbvjYprbsiCHgaEm5cHlRcZVH6LYaU3OnJQdCDiOwhcVWw8ODkV07PQy+WSQlLNeUYWa
UFcReuZ6HGt4NxO5uFsALv9Lx2/Z6HyV8Q1X6WgReJDZhvMQhH9iSyl8MKaZAhspySTa2y64QJkt
rR6HjvxgfOGVDtJyp72k7z4nuivVcdI/I2d6bkEAb79tn7rfkqSzG5zfA4KfaobVL2Y2Ss2oaUv5
oB99blKYZ+gkO6XLFvC4xsCtsr6FRRez8ewwROdMwux4Tc+Rdh9kK5KtAiA1uJj4eCiY5Mc+Cx3a
aQy1WmYjf4nbAggiv+49MePCYKpnCkKBqsH6U5edbAa2AwNHm2vRdKXbMjNEGKrJbTcTRK1reh3q
bxTlTKSoMas/iWRbNY4bY/Nmo6mMJVh2LnYs2hN3jIw7BXlmLq1LonhJG5h/00x3AjLkPJeB5fg2
oVyRYZqqA7nydFLQxT2XtDhf4jcSrCQhJwvZ8PbT0kLYcWUH6nUCud5vuR/4DHUSpZ4/QRSiVD7P
MLA0UHHizSglSQtGTjN5/X4fWCfIQZVvDWl1CJSarYOv9jU7O9kaGlyQs4lWlO3R5/f/DGUUKRmI
JLXigVaUnb/AUCTIAwVQQyIGUqrFaqO9Vn/WlziQC4PnpQXcNDoNF2xMkPoYdVe/xBbc91iin1OB
e8xewf5DwxhwtMbMe23X7FveFVa2sD92kUKZNUBqGlK+kkivEI11Y4I2EtCLlYItpaxH58YMISGe
knOM/RLnGp+mr5osFGXJ7dpWBe63JdbU0VV1gNwobFWtZXCHlkMJqY2f1+PY/gEpnvF+6Kqom0z+
SvqwMc/f+UaLMKCnL4FcFFb+GHeJGRByqU+I5kCioE8kY4Om/ilcYN9UhMI7FfpYFhPQf11UoT73
VWAMXhIpMDCXwizw6tK/ausm5TQE05RkPJI2TOcXzs4Vxlly+O21Sj/z2GJVWOcOl2Md9jV9B2Uc
QrWsXq+h9LNLaHNxWDxZueVzUIcA6p/e26hFhMW+UTBieUj3PNVjrUQKMTDEHLfdv6+ENR3ViPhQ
mA1/Wq/bn5iXDE3s5Xv5rOi8fgCj57pvr9DQjsGcaASrH1O1aDdOfzyxJW3a9Lij5wr9fi6eVaKR
HcERlJ4K7BhidGVkGh5TiOzyoud36z1YC0lPXZX5EGJ/2hs9tyzSuPK4+1qP2yEla8Ms94XIVj5/
OIKLaofPWJhneeCWSQSlCUWPJ0CPLaNomBWgMDKYEjF/ZdmC6XvpRENgOO3JA9XBoy1QG4NHj9g8
6plBRi1XsYiQmMmuqONXlrdlv0p05teP6F5K8y+Uos6qHPPpYPLc8spfTKKKMqOBsO/i/UbfX4KS
9teX59yjq1C8DZTB8JZNyBRtb9O9kIp3wmW6l52SsXwjY+9dYw1ZOqFKwteCyCpH4d/t+Mjn/TKA
lQduI864jxZBLSxqOUQka9QuZWn/RFnMTAWFzLwkPBo0b2eaVhGGAlvAMunm5B6me6pO0Izeephs
7ACluj8Rkpl3N6emxwDp6/h6+qEK1dfxxmuh/wbTltVbk0DgUTUJLq+GGyiIYuVW8ej2wGypufMA
ImRNRUXh3C19vR8rKQZq5l+oC6C5WV/JwcFR40IwF90Pp2eFcFLAv3nX2X2x2owg46H8yv+wXeFi
TBn8u8GW+wBpIkPHgM6P1RJiNzhYmHU5ZTq4UEKziybFY2KHfmg0efzoz1tWkMlSTt6l8B6nOfNf
qYsQRA6ymr5G8BJllemxj2IeH0wNh5tEkdK1DD7wrxYoJzfrCPECu9r7tuLMakPRz2XFKVLS8YVh
fHNDaUIvxTrvwdrpgRYgkp4E5s4/Bx6YOBoI/TyJqPTgJ0EglViJv8q1ivoM61KIe2AGk/yiR0xv
3S/ln2RX+Y+66JM1Zu+T/QF0dpa/OAB1Cna8D0rL//8U8QvLi6e5edWCir3nMFAHzeXbNV3sS65E
RjINxNSGaX5Kx4c8p2Zya5RMOgVLIthn1lAucsVGN1yucCW8L//EF9itFOuaC0bYpyCsrB634gpM
hJoydKnuu3zFAYX/wryeHLkJIXYpzN6+EulhEecE4zgHi4MrB8HFN4LZEUMfWTqZb5+imrOUAye1
ylYmtH+mY+KEgXEurm+f/dBTdoNnl0yxdX6kRLyt8V2syPXzi0oUmmwu9tsTqRNEAuQRWoEVm0xb
NABRkt9dcmRTbLUILGEjgF33PwqF4mJ88coRNfNvtbfK+/AEibTJnVuCOEpqJeF3pK6iNDM8B+O8
1CSI9vyhuwrR/MHY9EhpwMUC1BRoSPV9J6VeQPm+qcRh3W5o4e0nkt+j/u4maK4ZHjurJsu1P/VC
uTk6BpZdWgIoaSLk/rslMlDeZINmZI3amZ7DcH5B1GqkTDi37Dy9Vamyy4Gj2un+nab7sRKpBlB7
FQek7k9DXNq+aZSrN9dAkUh25pXBWmtx/WR9q0nFwOKl7dsCFspLVhU9HmvFEX316lb3R3PENN/P
FT3oiOOMhcr6AiW9caiKV8Hexss+xRuH8xihGhoVCTSJdEsIkiombRFJUihGFMmEi2f8AJKLeO5O
W+cQqU0cpHm8oIo35OM44Wn906pe4XU00W4xmWYyd1KOk8Em7z4d5yw7IGUvIzwwBcc7RVmHzMpd
spfpK+MvEFgm8yXrT4P4CdKPS3CrR4mbSkG/R80n8yTCpTbjXrLHuKPTqBM6vEsaxSKAlM+TBtR8
h/LowOv90lTT+q/tPvvolTmEgKXc3OpdpIo+XHWWbIETag4P8I+TezKD7CYHUyOtjJkHpAC6qVvl
Im3gGUP28omE6PAzwNsMlXAK51Bs6wzGz9ngUc5/Bm2J+gGWXzsqxSHQ6NkIvqnLafv+EDEdfBgS
ToW+sfUsre5ULbQKs1FnWH3spe1+qnyaiC/n8GOfPrlFP+ZxwGl/VcVcJ62lCa3/jhJ41XBOBshq
GAxxs8TYmUPEfGiLHHx3W8VXGGdIOjk9Zx7C5SS0mqw50Wlhkxc47oEeUe3k/k9/6kWI4I7zW+iA
GLcqQw21gbfvfgRa1PYWFpLZyUCU1hsulkVmXijlxQUQc/GaXXqIvaYiu5IlCsDkUJx6WrmVpeiu
xGGQ3QgbMCj0UPuBhwV/+cetUwFypitlRPTq/06BIM+Nyn6VrkvWKU6ekK1IRz5kW9cgKCDb/luW
AQCF2EfCOoYW6m9sUcs5yCJ7HpOiEPLn620OQ0rWiTGvZHiR15F7SjkINsoVsd0z+mrpctyJC5dQ
wVMbpigZ/XvmxckcMwRF5uAqgDZgQqH0B+3/FvkCPlA6vouBNlkB0mkAzUVNUkmuj6B85gVKxRnR
4OCZeOWvjbhSQ1h2Y2vMIL/s/W9MAXaob0JJ5WPQlWKdJ5vB3MCmBN/siuLFi3RD11PAiQG53pCF
XlkF1NkIQiV7D4wBKDOqcDWIVvDjJwSwjxeadkToI7nxNY2n/1AzKOaQcgDt4QM2aBA60beLA0d+
nsWJmjdmlpgYJa8jRFMQYeD10oolStLGE0BcU46mcumGgBzoGDxRTJ/o79fszTe7xlI/roN6BJVT
cUzjeQw3e+aoh9vSsmafHhbJ30MStLydZnmw00daKzvVyAFYGs+7Q4v+foiwfY7GX/5XE3NiFHaj
sc+E64p49+hk3dPRPaQAKF9FaY+x782mrUV7PTo26fbJTui9JACd4sWCqndZshily0aJHBguZ23P
WIUSHawJr4ZhcXXT8Hc4Sa2ywXgkK8A9nu3UJ2bdc3+o1bVZx0gla0PHB77BJWavRKpP1k23FMR8
/XFJfJOVr0aEkcQDBxBwbcvgy7ed3mECVGIoIzc8gQAK14cJsyr7LHoM9XT2uUrDpU8jw8VbKBJ3
r01lD5zX1G7WbvXp/3iHzsPlsG/jySu+7tykyGcLyF8h+4ZXC0WFCQ2iF/oJlQF6eFb7iunwqTpX
cke1VB9s82gAG/+O0M/au7f0Kwoqg6SW1o748N78T/AUl+Dp+ZhuT3nnsXsOjuy/7nRUMIxqE4YJ
fu12SCQGEdKf9n0qXvZEMcoKrGy6fF+Kf/XhjI40et+VDt9evFnyMY3zgUEIfZaMozMFRrUx0oM8
9skDCsnHkteVAVYOXgE828QxbW2+ayR3rWgavaBgbTXvdJDYbL0/6pQpN2meA1vR3A4K6lnnX5Ae
MILIyXQ8aQwkAagMyAYF4vrPgh2qwDYSqiMErGw8F7V0VltcxILcd9RAxzhmUO5CXi6pJdpQQYPq
sxLNs3S5+leTzEihb1vI+Fa2L4BwMYhjYhMUmDOgcw/h7loyapvrDr8z7arStc/Rldb2m/vz4WJc
Wo2/pAJOMoDK+9Whs3MiEzQ9jg5aThe/o/eySlNksddFEikWct9HuOO63XLezO3/onwk4YU/2hIK
PEvSdkiedX0FaXAZBYNtaNz8lU3YoE7MJj8EkMQIvn57BG0qfBKz4hGMnmOKZyGH7rh9uYFPo3+A
1NpiOeKU0OV6nYcK77x0aIsAN0f8ebe+vWuzLsv6ChKKtTuHM1Cb1sw9JdTQtR5gTjV3/lOPeS/w
u2C+SDJIoHzV2MJVI0NMRPCqtAYwB2JNGgRY371O9d4+M6DzxBJpcuamsKMIW9xvaTN65fINTHKw
xaL8xVe9QXpFmpHDtItjdvjfuvl2izWR1ZyNuTRLG+xhJOAKRfER8wXAPLJ0alqK+vF9buBBwylO
KZbcmRTRlEv9oo0hLorHYPLcPm1nevvUTVkAda+ViWOxKBVqpUINzq1Yxn6/VHaHL6IgL3DXxZws
d3UisqDE3gqdnDTBYpfedvg/xY73AccgrKc0bVh4TS7vyH5wRqbYZfCMEBB9Yne8qs9oOkNWCPwG
6QI++s8Bm6NErTtcz+JZVtptMrr4j4rUSH9wp6UKQZ7uSKnv/6bE/EtGLrYclLE46rdScpRbi138
CIcEyki9FsvKwAxrBT6ucjghuTTAZSLq8gyDqiOdYxF4QPZ5JfWdGl6FY12n0IeWi6Cy5ngukZrB
lxggSBbTqA5ickHVrDWvHUJBJ88o/VOqA0RTfn/47Wf4A7m6W73xeODRtAWQtEl/Qfo+qr3IjCkn
/dT1XsGUkpxolvC/jjDQbSACKSlEzzdAASe6TIgbDMRauz6TYTMCkZ51r0eUepslTSdnbgWhnJsj
qBb/vzoB73dt2N8pB0trFYWYxjznqIvzgu5tiahJlZ6zRqy4xryrUhbg4Y/IHjL8IG5DHumepC7p
VB/VD5UrRHc2RMm2+PP0aZwV9PoDY5y0XvzMmqK66bK3Fhvmqz735eqMed7Fmwaz04rlbUKO2Dbr
QzPvy3wea+ZYl+gLbAdHC3Y+O8UHSfvVV9mz+jjIco1spElGcvsLcYiAMkc0A8K/peaxyTRXiZRk
uhxspPA5RpTy22xo/XfsLOggUHFj4lVvLCJZI0tmSfDEZB/UhLHMASNLxMO0+Bgyn989W//Ime+R
wtbZFiuidc3UugdjgFBtFtBqxP3hSElNIfENAfNBLUSpeyDUROvZb0vAESgYHk7hrbvZZ/fW7D6F
dAWGR3J0nCJn5GB7c6c2AZaxF97oUmWhy/4g/sF8waTAFcEqIX7BHyAA8SBUYAEuV/Xxt2lgM6Om
VX/7ag4Dv47WQyexi+25qr9TX3iMJqBmjhK+2VjYGdoHHvL/Id0JSY/GFNIf54srt4KZFCDfpPoT
fVsfv9eFTPl6Vn0LdeGpneHQFsv/LE1XaAdknJpkBte83/mo0pvz40SVX3csBwb4BnQAJn3Ut/ts
mJOnwJ0964sZRs87tSFuP0f+/ycDM6faDh9GohB5xS4N4iMDI9I4gVVL4lvBNCCfh7GhiDgK21ZW
JMomsL0Qynr9u2MVuHsO3fAxdGxv7X8ax6GsJxMDcGeQnbUSLOcnqGanJXbq34Xp0WyKNvXOIs5M
SCIPS6u+qtKTmc7I51fMPvk76V8akfi0xU8RsapdnxzxvrVk4liyV3Lzo40fWVSDfPh/dbWSkZNF
y3VzfoiKq69d22v6h0tjitjN/63xIAfHcuhSwGNoPfQk9vZJzf/HJSfLE1maef5WTq6Iegwx6Umb
OaCLDGG8xhpdQlUPbEEM+dl2kdxmZD0UH/Lt3BwjsF95xc1ubwq/4/t7ciwXN5YVQ23ZWjZi58ko
uy+1q2Gql9XQ+5XGQ3gdPj8LJ2i1IpHrEvorEGKNU4u9bs9H/IVzrYMZcVmreA+DnkPk7T9D4qo3
Ga9EhQP/WOGht2oAC8Rx9L6jo3UwKlOayo1H5TF7V4IPU8tppfEVT5BGGb076go/tzRax9PZQsO3
8X7u4/bjrsLFlyyVRj5XkMl/1Yvb8PniKW94R72alP09XIwW9iXD8soLPwRwwUfcLMeHCRcWoIyi
OUH+pnn9a41/HfDFV9N1hi3eFG/IiLxMVESstKHvGjdqewT6ttEt7r02z9LwvG75chfgH+VEPLT4
n4MoAuULAMS/+IckLonBKNEsA6oTiF/JxhBPkemcelkqKpqT64CDnVIcctxzOzHK/JI/p14AwDzl
fsB6yFwEq/V3+YEZVxk2iPZsATLnpsGDlXUZoy9mhtZalVNuMzNBl0C5ZA+Zo2WdlqiDG9OKQumk
Hek85J1L56ZA6kaMik+eVTkVdzSTSQFsiJdQazUOYqHWPU8ju/mxykqnmLK1xzwmgWDi9DbSW9XI
jbRSKd9I7JVR1cl0fFtf/5GPT1Q92AU1uWU8R5YS9EVDj1LAd1W0F5E2oJdeYq8ankh/+zmkT9og
NoHfzl5Uqm9BM/JDzmp2UDTkXrBHCLWGFBuXXi+DAJ5kQyBRFG0kcm14JBWPDP7YuZctMw9Q+S17
1GuaTXyh1F1en4mxrpmnlfmLE8gQMaV9s3ZBQnzJN9TFq7Nsdnew+MZPhqU04tsEpyRKEsBYxxQP
NNtRHyoYVp778VMEv1uyohasg1UDGDmIFI2XUDX74rj5F5ZARe+NFJQZoKxD0qQirHS1+xu86Jbr
T3t/yAspjRJ5KD0f9cy3hXZ8C+jcV+zYZCrPWAopxwqQfMgTY7kdZL+SJfLvVD3Zz61HQl6IOiGU
ozb3Z8IwKbSVqb3Kl2DbZNy6feZQhxUcu2lz6aN0Ox53zslzsDMbTaK8El/TKhQhFVZ9BJalDUPu
jGJnRVO3egG304G2TbyprzzBNcksLa7y508z26pRn/I0rkOjPBDwKWWS1KescbaxKEpgq/jfsWlI
1QxZsk9P1VgbGJQSN4/bIwswZt1hqzY5M6Oqq7X2shi2SJnyUALGC9f58nMulizWVmjyRdaud5nx
lwt4ApUr89oCllru+5tyZGt8t6P76RC83x9Kj0iIM7CiWKIOXwpSU8u51Rr8aLBJ+sHF0bNo58Lo
RzRxR2LbK9jmZ/Lq7PIF08kLn7IYRBMIAeDT9AXNmTgmmy0xrUpuyxhVsIsA4BGJhhAv7Y+sqn0B
JLs0FQx9wKKIdEWJXPvnwYWyrJ2FhVIncRQf+Rcw1nredh3wxUBzQ14jh1yiHoSAAwmFZ10A/21b
6b6gTVMDqnOyD/Dv3kts961GcAyzaWsYhys5XaqWRgHq3tqzw1XdfpayyHYjngXihKqFNtg1CV2d
Ku/RFFAI/xxQSlKzJIC17Ipk6ga8W0CWYM6SObm+vYRiXcdW2VWUq61f1NtTWuZGkvU6VNNe2TrR
MqLZkzo+0GxSBUYfK56jKbY77r6kNfHutH385DZfZyUVF57RznXr0TSnpx31sDT/6MSvaAwr/OUr
c+Fqm8wn6CoqVj/jQXPtBwruBP9J1qV2n0u90zMFH7hVQLUukA5gSMozMgcnvfDy2BhQYldCsIor
4cWcrigpgoOfZfa/ms6F+F0S1u30Kr9TwUmiq8eoUHo5IpVjyQdH/4Dlw3UkAbs7R1Cof9FgXfsd
U4cZv34xV8C4fxLHgLerLxyoOUiq+aR6aiB3k8mqMvNXcPLoumU6MLUcOoZuf7kMuA80CdglaOF5
lvvrOoE1IcyAqAqnMGLRR556/SPjcvAPnRHBPRwb8bUqkUeSp1ZYPFnxYe/zAfeXN0pvsmO1OxsH
9U/NMrctBVA5u1zWx1i9APymSHo6nA8zlzpNids6uZr5q5jamRrYB1lIg5Z1YW2g/IzJ5xZRxwZM
iS9Dqp3JM6Q0MNTI2WKMSP6NPhl2933lrUQGVJ1VPrGKltZCVhvCSE59oWTSaQ3V82UzhKPTjSZr
d33gxaCU8YY9cBDXF2zVRjjkyJ8IbLHx2t0JhsN2c9xQug2lf6Os6Cq82rCmRHOzGU5jTCPX98jQ
ycmCS+YOYNGl1bqENq6YmpGRxluQA+bokbq0GuOsNq4Rgv+lDVbLGysnAi+3AG/qDsYU46M092NP
Y5w0o09CdIsMH8ppdV++jUcOjCr+aVPynUv0hfekYKY0ixj71laKcYd4jTh+hMaMadijd5iyvdR1
wIBW9mhnn+8lHkQjwFxzl9Gd997QBme8DGMXS/H+yvlHaN3bOWQuPaIyLg4PXAn5o7iNxUoUSslJ
a7go8dOsc0RoQewoeucIGrrB8z8VvPMLYFolqCSq2SU3A4eLLNByGASMNYT6/3yyizaTkUarImAv
4sO5cfdodZs/EpQcTm/LE5Qk5U7TkZj7KBoDxjvoK/ljSEe/ltDSRfYp9XVBoT1sT3eClRqin0RB
1AXCh0b2PMHY/2XeC5NAjAJxuXoF8Efzs7N4IxufvG2nvMSCEHpBYqpSn4fDDkoyhM6kaxvNQiA9
fzzT7+mIKEq5kgicm52pUtLtQW6sxF86MYd8AeJUGtaXgT7XX3x8VlbBw2ShIAo5tvXd8vnWMmKH
8yyGt1IkpW/NYK6QpKpAMqnWVAyMPIJoZwvArs/Hxz4SjqkUzTdwaK7S++ypZ7w0ZvZ//qbCh6N2
DVDLXuSd+7qi60mnUMgHdeOIU/tGw0Ah8lYpw03D/VIh4rt2ezrbr2lzVLU1tVxBISh441Y/3O8B
r+G/UFFcNCJBdOQqDJiFJ7nj8w0RDbVSFD2DH6hMnYgwi8yaYfhvULJqM98+b/j2y3pCJQYA1H3a
JgbCWGvrlCX4aaKlDrQeRaJxKban3xuZ4QyWWN1OxZv4xxuvdZ/62/9Th+awMwaXFR+egqWCSRXe
Vlt+OXC364C7UWKd0sh4MiYuTn27w36ZHK3ACrzbi7eLHl5LkDfpJWh52qfrCCvMQcScfeadKroA
jHhrKuq1IFe6Gbp2cjN+CbqjlfLm2A3OUu3Wr6mMDKos3aBqVVBTsxauBdyG83fCMP3fQFjBiH14
Xb9he7t0ojGpGWGPXQM4xjBrlIbU2inTm3h1xqveNeIZn69u1FH5LwYXct4piqs6ECmM2rOEhoL7
oGiWbYRnkpKqGXmrLnJFzEpAFOFsq/PK7zXDWAiXWAx5YJ6xQCpGIy69NC+LPfD/5bSenACHXLjJ
ftIsIUtSwf+aVq4gHguQ7araqvz/UhfUmcs9krvbfk1/awemoXkX3GUX02CtjhzGT7z6q2W3FA0x
oEf8uu62jn1k+TMVuE5UfSYJUgB2eFgHavS60Koe7Yc2MjA3PfT4GnJ/Hye4yFf5/ElHcGi6C2Nx
XfPEC9vlHiqaCqelHPsAkTRk9k61oMpLvCc0kxi7eN4PAjDR0/j9wJgJDSewIJDeahHWAiuKw8g6
6Bx6D47Abn3W5/zM7Uy1Wmh7aRl7SY39v93l8WFYmnVNg115pGubHOrgeQAg42nP/Zmcb15M4a9O
9ZBXUlHnZCGQX6J4PxkyRzJtNB34/O+3TRHx7gAgcGeSEzltwW8vm6pRCpNsdu9kjSfiHcbW9/Ls
WiHjrynqwPtUgqLvj1nTdZFd80aYbY8NtxKZ1UtBPtBP1y+7rReJbQC5WRi7EbPPr1X4o2n8gRoO
vsSIbWUXKML5XEPzWPCVHaqJDdtLrLE51HK7CEJNXWRNS4G00dFeLLJ3cr/zZSQh+sYItq5m1TkS
g3I0BX3HHnqF0FW49tdL/7LhbRPOEHGS36n5ve2wf1Z9sVBFdFNAbKXb7su0M5WZbSuTcJsv9Oq/
vFIVgrkUF9M3LJuy5dmu1fI3o3c5HJR0y6Od6SS8XE2eGKVSmEV8aN09HGWweN9j75+umrBdPWne
GjUxKZ2o5i3n2//OMeqzkV9tq04LPCUP7U+gnmLN3l1DFvOo8dtJxj2vVGpFKYBXN+HL/hh3V/i3
VS+LrjJVbwo9bOKbJZ3vME4YMXtiGgQmTZ7zT1q2nw9xoc48kvAvFRyhEHWHOmrD8T398mgoklPF
ZnB4f8GdjNXzRKPiuOoJwYWpsbwvZLsTBDij4A5hiaZz5WVpdpSdkB7dS4i+KQtD5uCC88p/pFke
gsFkLJvqElXumwYZ0KQZj/J+8ogbqvtkeg4vhRUY+FCmL+rfIsRjtCQrjqdnSFpTUwqfOQmXPkBr
gQm4TqOhrn+pRtl+PIcmkA2SchsuH1Spj8dq9QZaLx0dgKmrHyyEDW/+PVSEcxeif9x7+uh5unnK
BapaSsEKdAHqEBFHwn+whaH+/10gc/K8etV/+orx8sX3WETBSk9lDG3dLayxJ07OGRdkpk9mNhAW
d7SQz2BHH3br2q1bkuWprEnq8YkUwlkzOOoOG8b9neMwrwOVxaRDEskuEAZQ4ZBoj2VB2o3nMyzi
qsOo4GaibiBMzwlIYdEmYgMeEClJmEAl+y8O2o8UqZPCUtAiUf5ImB98khBnlfIGVl/D0LOU7JXI
AM+wEh63zUkvJYSztZisPvGgHWm1ikwM19Hxqno1KW/8OShPS/EZyKssEmx9pjubGHM9rbXTh6z4
JTgkIeluQcoG57BobUduVUmJFGRTy/KE9iVwq9DibfQcbpcswC1AsEym6j6Kx8yxnWjcz6U+sb92
shWkHRCxU8apjSpaNpa+KX63goEowW8xtVU8ii7CU4TA4kOhDfi+Ow7k+pkL2F266JN+m9/aBt2o
f0lFt91qWAXXD1aMGjcIXEv3hFbHGvuwnRFtBEI5xXM8QY/T2cDiCrVditq4gRutf6cLUnKjdz7n
x+0g+KvjJfMSLOI1wDPG+Tgi0YgmbdLaVQleOGb4BsnCwMtGu7b6SVJLg62N50//EG/jBrklgpr8
NNP096GVH1Xm+sOw0jnPKT4a8o4uCNiEeN4Nyabxqh/HofwIAdjqF/erd8af266AVcZzUKl6GUHR
strkZ07SOVzQVwOX9hehHmP3TEK16rBW17ay+IhZBTDZ+r1gMC09rJaRVeCA48w7Ul0zLDJgTiWV
R3MRoQcSRkxwmF2TSh30z2/5hp/VEZaTIzmcezj3By1iIbZzCEwjZB7D2UrVqayHBqQw0uPr3JmA
RUJa2SjuM2QkbowzCII0p9HQc6vSOsefpbUYiJKhP3xASofiY8diQVtU28oHBA8qz5EG8OruYE5d
jP4OAAWu43BPthbhBMg9h+eyWaD5M2ddVXSUhH3tmlS1sM7px4KoS+afHvAFA6D9Tj533BtOwLPX
cOPKqCSga3Pq2sVwELw7nFseJiOmZhMRTCaoxqM22ut03mDWH/UFF2lrVT7Wwzjd5Fr12JgFljdI
BjwNmOoWNWS/ZJ1VxJm9Eh3FloO6/W2Y5HIBfG/W1bmiluMhYoqwMjyYW5lqmCSxASngz9HWGH3v
Kh7ejBDLNUYB9QU4+HDWWVqbbdzWUF97G6Axyjn1P8vUhh9vQdNMYM7aMUoVB5BJyvM95PFFOHqU
4cmUQGhjJIDLTV9AXeAQccFjJE6FqjAo70hLCloN8mWvWvQTzNJaPV3WUERwWUzz6J7tDhCAfkix
Od0e6iMIpQOYIEwg/fLW8yG1M3kHnpFbCpcnqcpgM7UfcMFvkSqBWvqla0jIbv3sHuksZDj6eAai
dCPnlYS2rGP0eJciFRPJN0AxoHdgaTbAnDzr5EOvaDZO3E7rNL2X7/4DFNKb+olUPAx8FA6jsM5c
WxtkZ3lhFl/RNDWS0+7rndamfxAdYgYvPHR+CA+sFgnfrvNHNEW7jtvSEObppzQQLvrB5KkdPpv7
E7yh3Gli89Blu8LfvQjIMH+DK8UWC91j8oyIKmMfZVCJhrl1OwF9jcqMdhNNO5ysLKqfEBmpdEyT
8eF1tlNZ1v8W68oQU3gxT5X9+F8Ofjt4PeJPUkK2DKCpaS6pQlUwgeyz3XiPdiLy7JrD1iBjtwi4
IqQVoNftnxS0V2MxDxwCs4yXSxiZ8pF49+mwGkyfBzBjMUwEUZGIaiLl41cCf+YYeGIfUFYsNHaH
HQzaFHwT5b2/keerbsYJb2+HIBv8z7YpgKvTVr2ZMB1dBPKGG84uIwplADnLYYXtII9Rm/Pm6dOx
4Y+XMaZsDmNKmc0s1X4uTTkeGQ/B82kcjvbzFwdZy1eKJ4/3t9ybn9W5yuAqjdHwgGsuRXI4zmlY
5okyWcOucsAMGjWzlxjpIfxSeORiRYgzBXkb5epD7OHPHB+nMb9v5i4KfjcSSMSfm1XIBXhvj51f
lMlh73lIIOZDUUnEDNJvTior2+OOut5WQfP385OjVy57DXvmr48nNpqv6k09GuOqELqBoAEDAsSs
owS6GCy68el9tUpuigyGUP5doWh1fq0T6Z28lt6TFuq+IPMMxSMcCSRxqp9LzlcAhYhib6PHSm87
SvWgI0iq+/yB7QJ7rLA5hZ5CAMu4ne3zwmX9sPmGhpwhcCBl1/nnri5gAk5nf1aiG4oTjPhciSoJ
NghTQpNVpiy0VEz2gzxXX/5Ny2TypDzrBwo9si47ysWAqmhLXFtdvFjy3EulA5SbD3pPDsi4Kquf
p7yibW0egLcw6eCLM3tT2XT+519P5rmheCOYEno8Ce67N6dvTim0w1/qOLk8orQtVn2BtPmAM5Vg
lkKy40qgIlC0rqNtEvWZJptwBEw8HT6iF5PkvfG9OVQAHaFRSs3/AbHS2XX7Poj5xmSUlL7qe4ae
OnUFaMDY1VbBNDGataMYP9n7RaioSEMyL5Bcn1fBCsqN8xZtZGhHF+1d9djDs98KlnJAZqn6w4c4
QrdxwHFxqY3+Bkq+xR2osRILy3d7Bnxyr9D3rpMAJzICda2R9eH50T5/esLVnjHJXI7oeICscmrS
bWjnRTmaq0KbphJ9LRrliMsIiwk2sr0HTfLzMnr4WfBuW00Q/jajf/krLHUp8H9E2rvu/PVKsPk1
KlxTn3jjRm8pJoPqfZo0UM2+X1s7Iodim9GFjyeM5GtAmxkc7tImvs9Rn3jkjWbrCcYqI82GY86d
8XlqmSmFg5+zJJ28pyVa12Cwh0odHF8z0pa8lClJA953x3Y3F6wDlgoRGBRdT0io5OaGh9XXpojB
6zJyhBXGj81uNvAIn1h0pHkARk0NoMUA4cxm1/TfnoyvKU3rDgHKl5rjTf6ZPjlRBuFiXU9cwX4e
w2QAGksUJcgpXnjXW9hGrpU85sCr3yTVEKtEkMGmEkATsqtcA1tZQAF91fowaqNYh4hiTZRXJBhN
mh6oU4tSlC5aaVnJpv9WOALRU/ychwxraZY0ilvmKSwjdQ5upfCKngBOG+ncBypSHA8Yc3ImhO8V
mE3hFOvSOusKvG1lu+np1rsoUlJAeAsIJsJ9LNMIUmoSqEj7j/5nB6Tf+xPWxivuX+hKFmthZREZ
kwGGJQZwlPO5lSBtlNmhuCOlZJNuaEUABmXA04p+BTG7q9CblHZyZ6Ol/EyCAhsoz0AkvYjDkfNg
WIXWsoG+JXHRCnsT9pUnhs0FWCpb/TdzzTOEceFUQtowGc+VUHqBbBMEBnNJBS7q8Fz20Kp4722h
xCp9BU3RH6fO6eWPjjy5jwccJJz0lXV0WWEnRIR6Wo9Kit3V46kPoxSUxyyJZfiXpCPgIJP8/P9L
K1anoQDpqt7C76tLodGBsIBxdIHOt02wGhk0ynTZZCoYPVGrxr7RYwfJXrN8LL+B/28ME39aYhuV
nx6xlqoh5Oqwft9TXUnWG6pXMzQ96SIrTx3j6rmjsE+IjqpdFDRAEH4L/pXYnOegUNne70v9ZEvZ
eGRjdYgbPZU9EL55SUXXXEUZGXLcGII8rl2zylbeRadXrFZ5jhbHmmSx4K+AG0y3ZMw2ZCGQSJih
KsfLfIWT9GEHv2GvID2WbA2no+P/M6EaXNfCfpZEgXV4rkfymDnxy5kwY+TSSyA/KiFRXJMYMJV5
GF/efH1OiBPgsjQMvmD2rmVlgLj5Us3IVA5kCMRIqtJnq6TOwyBifgx2GubG6480CSC/PdKRZdwg
bTvntkEnbdTZWKWWc1pjlLof/ppiF0vH0yOYm0TsWyfNhBTY6Ef1M/r6D0UiZI4YQrOo0tXkue3a
YdBX4PDv1IuTI4CxIuzB4nL6t+xLvvdThts7vI/lJjpziIKcflNVeGylkx82Brm+NhugmSSIEXQY
xVjDqhzSFvYVEnxsJJ9lGzp2evvOjCu7GktI4E96tyGWAGpazfzY70GcY3qS7hOkXzQ3rAyGECIa
Y3om+ztnPOTHjeSg9cMsVbnt+8cQau2jDH9yPkZRl+HHkLrCLNGOGOSE49GmdhoYPastcSkY3CRK
rtXHGJDnrTCVgZfW+4STOPflZoFBLsQ/CEcg8GLuAdXfri4OYXcqpBpXYw3xfGYVVm8CX3LjAW3E
oU6hb7PUdaxg+5PIGxwxSCqV4vNfdVEgfhnd7aO79k11XYRnS/kHlea+TtJXVIyIl6HReQVck1I9
seg8B1ppVqT8TIdHE6OZgMqj3x1ESMwBYsGEjHFc+k1s8pNrrPdDh1atZuHbg3BqjasitrG634QF
zHKqMHHa178WJvdLVN1HWdMbwczq4wqUekteOUGL3UHbPOD/EDGcLsx+8IYdK4qhgr1lyDm/NKv6
l5U50xlYZd5QT3/GwFFTIFynSxl75hOI2qxqSL2C0DtvDqAJGX7YMCLr42JpXbYhQdc5anFx/yvF
YedSVz657PghkqAyTwYgJi1sJXvF2i13/7m6dHBcpMbubVxZQjB/OOXzEYkRpO51aZQ7F9g4PYkx
sQ/KFTux0WyF7pHWJjCNqmzrBAkZGBwP6wiU0UvnaVdega0GxZTF0dkyfGLrSSqsihS8+GOGorYz
bvnqI0KoyNYqtj8ZlAMV+D65wdMhdRIPVcJVMxRiJFcha44UGp85TeUpdkQHt7jc+SB9Q9iddRn0
kVB0pdf4Oicj2DWsqLv37+3m5LtriYljVRyXSWUeO1LTxMTRXlqhUtF5hD3lAOOfmj7Yf1E8YR9Z
tBE5lEvmWn6pS6vcxXoSSZN3yR5xSom52/HTV3xEB5xMWgjOoBe/5X+Elczf0TigaYFlIysz4uOF
ckyuIsH6Lc+3tArFgpG0L84qtULAZTn1O+jh9Y3qMhFbU4ylP9B9nySI3i9vAfc0p4CItBX21VcQ
EZqCUjvPEIM7gdaILFfmtbZOKu9U1gsZ+snt2Iv/VxJ2TtW7RbqV1gCzoKfzo2EVb626mJQWuZiC
kzjsjkNiytTdaLvTkTC5B6pKCQaJN09RdzWGFBxgcFevQNm5ermbGoOVcW42eDsuSerKn7VdCPKl
a7LHhU/GS3AWJ2x5NgfDSAuakT/d0HdIjd+nNwDpYJekC2rf6OQ3eqmMIhuoyFIf3JTo9ucBrKHg
fX2VQDWwjsg4YjJtTw497M5QsTzEU8aIFUWKzsqO1/2ChcDWZEf5LvA/fssNna6Xk0QWJKkTJ9cB
1BdGnCk7GIsKx8lujKTG/ysrduJ6TIzzll4Ioyvim+scjPy/8nvg8wASnTmwoW0tzdf5FNFTr4pi
RfAfL94fOXP31tuG4CDOn16cteMBIKtOESNRVudrG6f4KOrxZ8ms9fCQGrKNNhTuPMibQw6YtGVw
KbaBzPQSx1d2xltirQIKxFPXh9jZOtjAtzUGkvyDgKUunRdnV7WuLOwYEuAt3H7HXOorpx4drdtt
UyD44xgB3g4DlbaAQwfNnY3lGZF+79ewddL+aEFyrfFTw63+SRtdB7VV3/lumU5Ca7IpclhEk7g5
y/U2KM/Ov7QDzN9EhyBe7s/E7lnoBBfuI5F92a0poNl6vlMfZGac6gNIdt9MML0EuCe0OMNspS7Q
CWowlEPpcx49QrA/EIOEQUpQznrM2lPQRnAiPgjdpmxaVI6QScbCUFRPQZq/poydnIwn80J/dZlM
cuPtmJNZzOdzosRYtd3FUUGgBQK1XIg9prdt31poi+DiMqeC9pTwK0KYgmkMW662f5ypWClm8j9e
G0ZbdXeApOEdMqb/I+RPYmHSyzPyBJscPmFcCUX2p2PAT1pdjYZ2j905c9iITnUYnbc3xNORbrwM
fPXJtumWO+nSHRjWw/60R4DVIvi86DIbpOpPlQJFTijE8bofNesESriCAheeCGPXCW0d3RWL3vnf
K2MaB6NlUG5ciHiff4cmIfBjqWiNCt8ScGaJ1iaKkurz8qkuDljtzEqNrJe51qb1GJnZYYjyHlz/
mgnNXpQiUFqRKfsUvtQ2/QkO5uRT1pt8rTEsxGrcY/FC+InBWgU4JpUs9kb+8yo9Mv4y6L18eypd
PV/7yZttUobZL945hvAzlXLI57MO1rD1mgvdgBbXcUYu2A/RPCcJ4Crj3fTG9HqXh4I53yzWm6BJ
fgitkP+Q58pwhdAyTsOFmnC/D1U4yIBsojMmPcabHMQpM9ukYVbw98brP6VQpaqSTrWHf/Hf47fh
Dc5dhQAKX4cyLcG8Zvb1CBgdhD+cB+KcRxhOSxdu5cN9Qul+rBWCm5tuGo3M6CZFcWr22GhtmT9M
kKAc7ZHPyuPEaPSSONs8NbMQgmgBztI7/M07cG3w8MqmzL3SHIQK9zmP6VV5s+adB2MvpsWnZ5Iv
e/qiDjE+t4etkllv1Tc1zzfCbhAT6QdhpULxpoHBhpSMvnDyqRfON5Xs2QLpKxngAmeTmpH/TasN
zbRFRffIwrYpLyO9/ld2fALRQByQJMnBFF799Ux7vu3l5zm7r7OBCk0IMea7m5dtWmfpZkIJUmlI
wnJMfLJrNPPvVNyCo0WYw/YMjfl9/CUIEBCLG/x0CQFOpM3KkufhdvjLBrccRwNSpZHp9PFuA+dN
ZNZMKW/onPTvly0VSUpYwVeeBtlrdS5Bj2btJM1L8YcT5sQNL5rZ3Gljp/8L5k54kHZMrD7NbHYJ
kTzCq5tw4UMKPWM56bweyq9ObjDhqXeqiy6Vw/BAO7HvSa556zFqLWwDnJAmLvmlST/UFldmWAjc
h2lCWYdzllU/Lm/vYBieeq4FboWsm48GghM5gkN9Gw2GmhHFgrH0TcAD7E1t1pUa/d8KMqeBeYjU
DeZ4yNwF5j17/9gQdBXXg6ZWKZlBEieYIVp9tc6R9A8VhB9IxU3zgjx+4EDnzgIHeo6rxUEHrzZB
lsT7r4NcXoHQHrk7vLwQ7z+C33FJADioLe/odV+57PC1MR7jtzKmeyyWhvKRwPRt5M4vL3s5EGF/
aRXL7Jfi/NxX2/L14lL6wbOnxOGFRS8HTPy+5ka+51qkP9xjuWBBx01Uwwb86lAYIYZwF8K6oo93
1UXmbvxJLFH08aciTVpeuAl2P1/roMwVjB8/TD54+1dS3/VTktJB6ZqRMjKY3xFLe7s10WNKq9bF
+DrQF3EQgPECMM4wuLp1pnCGHOUT+sVv1WgDxdGFu7uCOdISdg1hB66fCWh4PaOpjbVOMsp7KpRO
VKgYWBa9iu0sXmiL4GOmTnzzMvdVto+A7/RGYGgAF0l3UEjR+PRvYfGURby55wgmqihH96x3weGr
f1H4HP4ZwwFUCPlnHQGldLOqnRqu7cxMr64JJDlA7sJPXENSWGjBWBMnA0A4ZyXQIp0SwDIdvClZ
EnLCp9Wp1Ahk9sXOi+/lExrfm13PmzZIq9HJDi8kWHTIllZ43VAykad8B8CXx4ekcgGBm0cCXc7k
MfNqWUrASFYnudbaDYC7KHI95CSqsrLbCxgIc8OD4Q89POdwxSeYwdktGwhNzh+qwOUTBvofv3sJ
o5OotTEK8y49np+mM77tvtuVA7fEjOTtPybSy/VdIYYmG5R4rUtghjhK/MdBUtKT5gdA9VOnC/zN
WhB0RSBIEbi6f0BQ+C6ZYaPIcMT5vy18PjWkyyMVxEjd5o6cS1gqgmgmC4QQbBVo2FeKaw324aDz
s2kMPQjXPebHCqwYGowMwxNcdp1FMsonxQxck2iCjhzRLZEO6a/4MSh5LRDb0PuaOtVoCxEAeq+4
lDe3M5AW+kTGRkicBr1FTxNhHVX8JTMYHfFQJWKulEg1C9W6N4y8GocL06cotl+yMGBQGp4xnvJs
YqtgWr72oNQybQBb4dRK7zdywFR+opnPFyqBRdYJKlUdhS+r0Fbwl8Bj+ezNZAMYyix1Inr2x7uH
yh5FNhurLwvfUlGPJ8wx5eHfZLs2DleSVLJs4n57gXLAk61dUwLOzRVOjBUM3nO/4un1kuI68B91
x2UmHk3AaNmD1i5WoTgz6j3po9RKQHmQQYRV5ZtWfINFbuC1eAjM4Ssz1T5Xc+XJwSs1EZPqlsBJ
HQBe6RBZTVlNdiEiRxyxswt144p8o4htQxRPfI56sH0FijBg46VZy4yqZ43nY7HpniYuBDVHX0Za
zZB9yh/+CXk9PhN6nnm8b1/uo1mcmfaYyyJ+QP50P0f7i36QaLRM0TBmP+EGFWzhXTu6dPZ/Jrjw
uFC9DQjmi18fhpTPmuhdvx9QvSv9eFQEMKZIuizMeaOnaXIA7ABmvN8Ntds5DGq+meXJVyBojZJx
Yu1RS0N883RNHTfHF6Y0U6a3YGN0hO8y1BsjX8skp5+BGSkSXoQYzoC/ddtgoXkubDol8UykE35F
CI6KTse1w395MG71/tLNDFW4jBz3idUSbCR6QG7qYmDGOZiSvyRptFyzw/xwOl3ELgvnzvj0lUJ3
Dsq0NAnl5qD1qcE5tefc/bnPyXEDSxmFepq5EurtL9BJ/stIrBffQ3FEF7zIRW+ZN4tyYYHyCkXN
SUTIn6+3Ksy+oJO3F1RK5dwgGPJPt7PZ/a9Ssdmits5AiLgtlRKW2jHTvbjgspZacItGJmto1fRE
7EiEaELa5FA3uNVKVUxUnRUdiMkNU2M725AaEUmnLVWXlNpms0Ya9KOA+/7+a6ZQ/KtIWbmK83Tp
UCC23+BmdEmmGoK6bUX0sJRcgztOjv2dGTqPyAezeC2mGnSkv3CKTDk89b5kfiY1cheXkflSOTFd
qT5cNgFVFJy5HT/sYQQMwNqq1R4Z8mHy+zCtUlc57UeVro4EigQgDRGwuHJFPtkzaqR66VMPAmaJ
JJ27B+sZy3zv5u/UiIkbeoud/PfbNo3znfNX8mNw2/g+q3GvGaythxXlgbZL5UxAGOOS8FHFNyrI
yy/4+CeEBtgpHdxF0CW4jGs9K9TyK8SteXz5ngqFM/Gs3vKKyj5M9CDplPf+mkS404+2j01ajCFp
YIojYpGzRKMg8smqjc3KPwrC2yE3xMmEkJL/t0Iqysxa8rFnyJitEsLkAXTbszOQGaW2s6c+hy65
Nr66+b82lASdNBlHJIg7VzedQMzorke8HOZw3n3qqRSJ9DixR0Zqx7iB5wMe6PgfqRM3mkHPhnUp
0JoURAeS3vHToFgRwSDtNtMMu2fRxddhcbrMmOCBBaghG1Dg48Aa4Ue4XKZrf9SPsQruL570tuFk
csEEAy1hZRj8GXEXl8cSC0RAw+lMr6AAcZFq2uLxxfsUXilhVVvdqIGSt8zWGr44S88gMPbekbA/
ljyVDxnZL/FkjcIrvexWjNDpzshonZfpM8QT/PN35fo9C4/3ujtLRbn1MJZLBfGOsEhuHWDtI0GR
AIZcegWabOlJTBGrP7OL5l4McvifbYgEfj3ZQ4uYshL6Mf3mbOb8X7l65IGe4ESR4c5DOZKybnw0
c/mii6/e/KG7PjXcaId3X31VvBgAeKqlUY6NPpi0f9BWg3DncExNjDHTWeTZTDGtP46ituFFaTnV
O27gxzMKHdyoT3IXZr/raBpf1ZhBTpHOqL90gr7oQ5yx8VwklRGfHEpMCQn+KNnRl5dykN2GmZmF
mm0HZdBLO/6Ilo6z1t/HgZn3P10/qbTXGIkMa8RnJIigi8T3iCPw55DuXvKEsOir/haUuR1FrgnK
NwAJ4AiPBHnSZh7vv8MOxommscKbJagOc+IiMSK8D3qQf9RghmDRJLrexoWy8MF1n/r4To6bJ8W+
z2ba0cNNmmp/GyVoJ27yVqYc3N98eBepLHCP8Kdud8bFbR7XQA5YT91KPeUjl92L/bR3C2zqtId5
asnpE/eZBM2KAJu3ybiFB6KdwVYJiQ9WuqQvEfDUInxPAy9AGrQYTm+qLgo/By26sOggJZMzm7Wd
+9dS08ntUknQ98YnmLFP3wa3REOY+48WIHi9GukK9UbuPy+TCeh4glPXJhtZHqd6ZvWz+pHDmoVZ
0kaq9fCWojSkcwr5WtVfWPk1NRBLsyi1rW17c6+0FCdwvKtitEqOyidm7T9YAo2aZsIMo//8uGO9
T+h7Ko2l/RevqkiJD7BvfpsN1kRuoJC6I+SIesLav59jAKF/ZCud5GNzDaYmK7qJxOosXRfG9N9W
baMpYhneZbQiXd632jIIkaOLr1QgmeoHYGMJ0f+EAPfKqKJ/SHXyhGdPOWIVewwT0S28whWyPWtB
ZAPYZQOM9V0Sdgv2P5pw2kk61Q9xZ8kWmuIpVQQaNWPO9qI4TtCWc+knOY8+nEl3OmCIVTgr8s9I
lp9yYiUydd1xBcEFl+6fWVV549O9iF1I7ApFL09v8oeYNlBgSB0+wxRIUFxC3LQhZa0C0dQpPdy4
I0KFTgAbBkhjAT8/0V3xjTNI+thlxuCVJXprTrUrOyv2x98682AIkQZigsDeT3EJyKtyJy7bIsNR
OqQifAXgEhniQlyqWWnk6/V+FGZGhuNKCdqlxtqwsJ83Rd2IVwMFqFJHGEQK/0EpLol/94qFMXU0
mBlhYonutP3Y+LVyArnfMyqhKzFsXm6DH/I10C/0Tjzy7jronZowrVUHtBz2XFIg4i4I7v/qTZO9
Rm/M1w5pC7DtVy9QBQFEcwFcqHFYoGmYLS1C0ZgjTxBl18VVW+uCbwkMk1y6eAo24eEtn4VQ8soR
dmGP4JB6boFNGUBe/5iz7E0qqy1rprB4F3Po/uCI1z8Sm3fNXEfCNCHodDfmNhdBqrsPJpscKZXu
2ttIqAT4ZCS84uV2ZeMv/gV6vn8vd7TN02PA3BxxS+KoLZr1OYW+lXOScNFTAQrMNDYsZSEezsyk
0o7ozxw+bIP2fyxsaeRjfOaJqElQKRLJcyR+0mvIg5+O/iTa79C8gCqLaCBOY/xXNeIgGOYZI0rD
SI1fYsGG0HgN/VsqleYHc0+fuhPGxb26LsDe+hmC75XHiTXuHHSCn1CLUHYaiv2ALxrRhmcnl9eI
nDMu74Bqrw5AUZdsjBAds/0gJltgZDpHjx6lveRse5aiZkEPJGSq82UrzlFdOnG/BtV8+tGnOXFM
1uVMrND1fAIdHuTJ26JrTbGm8EG8eQTtE19Y8k7Z3p4oOrAiPdo3ltsihOGeG86eE3u6ipsCQZ1v
864xUfK5cRpx31oUka2X+sQSOT9nKWYh9pCLvpxRyaS8ath6aR3BxK4KyYn6asFGUKoh+sI3Yk0u
iV2KpxLKWumP3T5GTlVcH5kuAQfxpE0kiQA8LVglz/dq8Pweyk16EqLTw+eDvqwQy5K1bRKvQxaL
S9gUbuSjMYDsSIrvocAjuwjqcAdyHyUIZz2ZKbx2u27dMbkHUud6HeZ00duySStI+4VIeuRkXvr1
etog1AaMmp2EbKOPKMDTSdZDD9k1oU8V7F33HQkg6UgCMkKxWeu+7CIOYIRvRtqpU+eIaCX48LC3
6XrMGSjWP4mJdVYHThQEqOgXwWFyqa7WWzXcpBWmwPIDjJI1IGkglTqK+VcAbgs8a6KZwAQO7tB4
COAKy32D8hcebI813dkylHJ2gjV/W0/LY86uf5LnYFnRl+Mh35qKRsQ8lx6mRxhnvD0c3WNWNlH8
86CZ8o4ougKMjU9TIsKbtMoZ9aVX0Vo/0MArc0VDxdNdEkBP4adbGHNW9RR+FkXE0hpxeCRhVr0u
GhKpJbDOY1KLFr6t4FO3NDcRtXh6QCakIXVqf04dGGg/m+cO4b9MdLj7UY5V5pvyaB1W90ZNqEsW
cxTBp1WdDuHhhAKMVmiCwd/pXBOK/98s4z72PPzd2eELxNL3GhrAfei6xKo8EKfAz3Z3ceSuJpBi
dKOmCsqkbhuCZ/nn+osdnZCT2O5ChR0wypbt2Twe7r9gnewtac3LFf0Q8TncTFxFGpLKmZw5ZN+z
j7adMoIl7FHr/km0CB8MEb8m5MywxAA35d1HAEUWmL0dhZm3gJb0Gv8yIjgrlz8YMSUmylIyrVgJ
29Yyr7uwBrZaIBkX7dNvUHWvWgi7Li2QXFj8jSW037sKKO2HY/6FsrhJ034f+gwFAlX2Wrf+l89K
AmA0GxGuov/vhE88Geh6k7R0yvlGtodeAAZXzQNDcePvdm4oshKH67roq6QE4hpe24PMLCD2lbh+
2WogsGiDqJrLiZJ1XOOmKp/q62Z8ftnWa9VewJNsx32VR/MKzWQ1aBvtneIWboEpaBm9jv5XJvpF
zezeh5xAP2VgSTdiupRMYYdEP44+iB8zlzKcMdQK1JgwGnxLn87tZLUpZbRE1qCP8HfngaoefB1d
vQPfZ6sHzKfGJZUm8xIm4bvqWH1i+NoxSOaJAHANEpydNdOxOCUqy6JeHn6szVIviBvuQ4B7IMqL
K4BTEPnIzrFAj6akJv4kzbMvAsegEtmaArYhQjg0QrFfX2rf0vlGhB4X50kZ+squIlsaOsByxTrl
aJOYvuM3/I1iLBDsDBJQJL+gtrvlOLpvGRtzmdZbIPfeFfflcP5s3RyeV0I82iW7d7zy9BDiOTdN
H+4lfF8/F8T67NajAUBySN5UHLOKjfV2aTuoo0N5fsAWwrXEqb2Tx6WAW99eorlRBNS9Ouza1/R5
Cn1ZRw7sW8SPYNatzxSLh7lzcflBFxn6UuVjBLOfIS8ZdyQYm8L+O7fFulbqVYYfoqjrKn70xGTx
BaQNsDO/6B695wJydktnFWWOp6Tb7t8eNvHggNJFmDZ0Uc3bd7q92BzsKmc4CY9nwU6J4PJjLmWA
04PhFGrjgc8JAaSTcso7q0Fl6eZ3DpDIhmsCc9vpqA7zSsIoHq7xdN45XN4FjKEozEglVz3pXzaA
dyjgacDY/7STeT2w8Be8UZcPIgPSPiZmcfkXQfz4Ku4ZZjz7G0Y35By1Nj93ytwQtov+GE+4dpes
lDp+a292XUKsyLIJ41tSB6g8IRYQQRyz4QMgw1kT0v8stmhAd+RtM4pVPvB9YW5y6xBVdDRCoKxF
fDSHIXs86em+QPvLb2TSJsLlfrte/LvZJNV6ERk7TkxCSbbTTSYkfQLbmw3I3/On9oPjN/IxynUC
7tY+8lJSgncsDeAH20tWydfzYM6DjRG5k8k4oaBNgsbI4FzbT19Loo58loTmLWM6f6TO1iuKXIn5
IsCFdBLiqcg06igIYwqI8P9QiHVpWYeuFXXWJ7Z2e56jykeKSK4H7L0+PPU/LWbWstKL5hlTmJoj
kI0Bs0vhxM1swiSqvNiXY/iSnP0WeLQ+nCrirwYVpvBB0N7aq/Q3RplJDCv1gNBpL6vcb9+B5x/U
o5qSOYSjJ8gRZEMEDwy8q1ySfYpjAPYzUCDiSLkh1yT9fcXCrG4KvRNKYd9mKG5SuhDC101eQjg5
dmpgA3AbNnt0vx54MG1NW2yKKe+Qn4fTko3A65codeQsBra9FVEqfIIAMaNljEVJ05+3uccUjIK5
K9nJDeFVsJbtTDl/w9xdXMXTBK/Bzoc4ZyI9AUENPBRUdFbAIvMSLvQKIBiC1hc8AYkZxLoIihEb
009opaOolK2eTym449f8Z8jwzmlZfNlUValFUWAhLwdPoU8vcTmdNkkrkJLfR98a0H6DGyiY3YUL
xfLvbs8Z1uSfbVfwJEkBC8ww4hXkAQcLPHAPhHIeR1t+6DPW5QS58Vid6/exi1TMM5+0evQl9/b8
bOR9P39t36A/XrV63vjOAbfwGYZx6ZP2H+EHEsgJrJfIN+0bROTMUnRyuOmLY0jd56rVRNWXruXv
6vR63eojvxXPPliyk/tZzH+xHEuAVUrNj19s5SCyNoxqO5/aoVtowP5GxF7pu+reP301JKVAJSsL
h3CrphlpLLKD1nVpw4L1fxEHmCtxYaL7iFmJ4+Dw4zAu8RX+j8WpIjZWQZpmXvCte15UzyDR38wt
hs7WBl3dUE3sySr59MWpLkQy9VnVk4aatu8Rq28gusWwCNjR5mTx7bC+C2ORgKFJMYY+YQLd2BOV
HkRycNuuQbgynn46+acQgS8cbjarV3gLrx9PDZa69zxTmU5wVNhS3czUJ/TZwMDZtkbobesVC8GS
cnfDEPUQzvmblWDa+0dRMTQOALYJCksrmMh0tsMjQVfyUsoSVk5eIGdvKvpBUgFpCYA+Avz2EvaQ
1wSOOTmGAckXz2ZKsf7ApfOyXaClSd2+0eEh7EvzajaYTP7FFe+d1HN4TLHktmZYITD/u/vHjzIh
+QMiXER0OhKWdvPzuq3Q3NZInUTYKAdEP+ygURbT8NNalmJAZAt12FcYWmMACZwhhLjgVBhIFSiI
wkt+I7MCin5tbKENVxWO9djhSVzlVGpHobzrZHX4ait4Lb79+yV0eNRauQUtaj//vfq4Pp12rTR/
5ErGNwoLQlqwiKgVoW1fxk54TxwrlxRsLY/dGDZF1X2gurR+LuwpxCcqQiqez01grB+aKLJbrlb7
wPwoZI6zbGrSqO1tGyViVN4L3+EdThEprOr6JMYg2X1UyMpObmVfziOC7Y9gkUunR1Ep0ULqnPrf
gllXLN3zYP1zkJpOguOMP0mdKLBqe9kG64L4uzZEDL4lt41L2q2BmwErG9mkG0Hl2LnjEtUVr7Jk
0q8a2JhRN9+99PKHhTVivAH4hVL9+qz4nDPNbeqxeLNkHKKFhfYA2+rdIPXmFvWvTypVp/5VTN+4
cDZSFsrVsEEE/We7JDcDqb4JPYM6BiXUhZxesRfA1G3g1i/ixjZYHduO6EVEQBgegQjVDdM0jsEr
ReXxyNpCmXg6cWtwzgnvqQsqiUHUXIDX/e3lTOXB8TOlmbiv9IK5XX7G6G5GVXfihNiUdQmuafgr
sT8vDKyXB/c8Jq19CObKCftdsX8i2fTX8tNshtf++uXyyyHEjTfLcGE5T19a+dMvh3YdtKosne1Q
+8/19BHUVl95GDXGkMASu/arkkcCiuxm7IU4ScPI+6Ynr9z787Xlt0Qf8lK57wlLwSJ/m0eEDUDM
n+rqic5yetw4Dqg2jVEsqPuDDJEZKal0Qt9akTgSaVUCNKBbnxSNHukZGsSWZD8/a1xHmSgi9JzM
CCdWTNBxRoyP/BDRsnQQpSErFeEQuUpz46VvFCUM7JoB23U9efWuGQJWrOIP5Lki2d59R7mWoUwo
bID9tcfHR6kEUIFzh5+bC0/8Qre32Jo0VFo5Nuq8pnv9/oG+q8+JM0PyENpJnK1gjrJiChrkrO6b
BYUx8mZ0Q+J6KkLKo0W6Wdg2jEyIQ0Rf25IG8vCFUknSIt0YFGxtkpzBHufk/w/jUuXjIyiF3tj1
SdAkPG7rUvRPWRHuezNJUQZ1GfzCjY2tM1ArMnG85AFKI7ni/yGi9nLQnDwliRlccL/1ItURM0IP
nPmGwoS9zRHnWa/TFpKehu3xvsVelQa/kPqboeR3J+2MeyDQnWulDg0BNBbEz/0h0Sfysnq1kiQm
4Tt8wANoxVTeNBY+9P8gwsDaRCgaK07ASiO0NCseGKe4Ol3MG6hbhtURfgifPRidxR0KIaU3lvhI
IAJTwhR4GuDLRTZHrmWtUH7rzGGU5C8TajrkMoVcrQ4A9bKl4NmypEmYiaEBtN3EYwjytIXnM1Lz
xt8QvI5v26hpXS8oMi0Dahns0wGtdfYelb7kUGOYtC3bm1Ohemlx+jxCryMzsnW3sKL1pTDQ51T7
e4yPMuj551PWawcfomEe0JycSRZ2v6qpafFRbLWpnNw0e52HKan9zJTz9/Ej9CsdfeZE8ppB6hQs
nVzwG2Mr5o4AT9Uu+3gPSFfp/63JdeviV9oKrJcv5nfVLrEpprPnAzBsHob8GSVGtYDjo+YFlRvb
mPwBSkcTn4MfKAsWUlJv/8tHiIiVDLbvXG98gSWme4ljrrL9JEj3hFOKjg6jWSKGXtB3Ux/d2UuM
coi/lZHj0DLMF7rflPZkM3AVtIdHhuDfHa5y0sLtFQr/GhSTR++Ak7rLgMy+8vMoQWGFiKuakosM
i8RxCSiNvjlNxhvdYwXnpyEf2KLXEi8MSv191qOXuUrHK1bQGtPePhh1U+lXMMxV5Bkxxssl20Cm
eJgAP+iCoiHKajzreJHQpRska53ZtB7HtrzkB7lJ3R0rozlJH0619tESl14kD+9Zeq8FrplgWN4R
W+DOh/2B//Kh9soIeABkRYgekrN4jK+FymAPpMsAbQj7J9jCMVkJEHjWG9X+oIRSEdL3/dOGKXz1
OZTUZlbjAVU7b0rQh6a2qdJWEbbrsLTjOxIu0QQ+osA2db70RT6dKtk0YuUSVYQ0K4iEF7mR9CkX
TzmD7Hd6CY/7Xv2MXcSkKmdayJLw0wTg0BJyTx0QGf4YRqoNp/cRszPkiazm6AgddVjeCy4gB4iK
6m60mtygmOwfO+1Y+nUpF5UNLpu1Ql8kY7G/gJ2SYm6LBKe78lQibLqDzE9wNrH4F2UvZnKS8NL3
sIe5Oq/26WDigzmalR/Io0u+gy/3eBX+sCo0zVLi54QI9FextfSpZFwHHK+0doYHrwzyrOToL8Fd
e29bPNnyisp45iUbGtnmpcjFNx2nrTp8ZwNtkgxCzHejNgm6p2yLRIhHudYdiT9+tb8FZ7gBV/G9
zfpKLVIXFyxQqNUe+14WYFktO5EFihD/Yq/rzcy/rkCumpVfqYBGYh3VQFYR7JnfxdWLkfAaSS2J
8GtI56LSaXilreM53IY7SqyJ62G02Qw1N16KDP71Mfgi7V6K1h4ootwXIKw3ZWDv6PpWFPzJDWEV
KQEHj07xHrW91udUlMxcw175SvDZJxq+WV/3nFYw8eVNtztHQOXkWgZwbf98HU/cLkVACwc5NbEe
EnC7iV1tWJRLo6AsH0ofUAtD7eE/gPEJMuJRqv4UyrPKVs6CgKkjigAYh5+97wJUY1xWnH/CjZNS
qHTLRdEq/8i3s6aT1rfspu7rOUSL2RKZGn9T3P/VC8vatBHWMsmvF9AXdrzCbglPok8mtTHrXnGj
8iN8SVpPaVNqmE0vCpl4vOmt4bpT8Xpq00nWFG6n9LJMW6C3AMKoALDGIOAo2DTFxakMJV2F6wZ4
to9REBCmTcflQu2gVKEyJCgTTGpM0JhR+X5LbavvTt6vCt5tpO7CWT8Uf2CZ3MqhaZ9JjhTqGiyZ
4WKrrPQ7KRZZq5hTEP2v5j6KXi0XsTEgoYBlMaQdT54p7olXKDMvMeSvGCAecU+8b8rMnNw8Neu0
ou3leFtDO5tbi5cJuoOAlTaB/uLffOMz0TYp5Z6Qwe2I/qN6qTr/L6KaLm4JG1rLqLt2cXH0J1Dg
jFeiWj1iRSe4Hg7Up7yKO3Ve5S+oTWJk9DnGIkmtFH/QT9zSYCSzpD3DdkXPaGL30CoShwO3fgC4
TMBJm2RYZf4t8rUu7gDyieuaUYdT/cIpOZynY9bMDreD+3GUROiBA+NbZhTbqeVOanwtp72tBnYq
g1D6SoBV1OxyOMrNByDV6eBUuNRSE3F3HeRuYDnKZKzvI68rT2U/rdkbcHzandjMMfQrE7bKJPiJ
zuB6S9i/HB+X17QymhbcuVVQP/gmcEu91mwTOcUmJcEwEKuVSNHRlHzv6LgJrTu3jhbsqt6fpAib
cXwi3y+A1caKUaWyJgO/EBPveUxk/LQr63GM6MxsslVJFbM98bX+MiRj49AubC4aVJt48lo+pj4s
VSBHaB0OaeSE35IdceNRrA2fJi/XPaEjrOaQjrzVEQQRCAWJbxiwrgomZRy9ZGse2hyage2t4Ymo
ECIeamtorcinH0vWmsCvQCeDevlNxs9tyyB+QLTqCF3FBOq10xg+aC9hOg/A52IbJsiSz+VaCxm4
ZXM2FGMi4W9wlsNgm5RTzZ6p93k7F0qy3n5fTInvEyOfNadVoegOaOZsUliwJghLYyTV/5Cb+8+U
M9tyOQyKXr420LiUEF89UTYnhhGk3TriFQ43FYiQBx7APFO+IG0RPnFnAMqjupmYYhP6tsjj02Xv
Eo9VvLbM7dd1rkEbWVe/gc+hmtqkzGHkEKxw+H0FW6eUUFmS4tYtjsKV3RIFzcu5TUeOsxpWnE/L
5reZ5w8G5E7wfdio5cTLwuiiZFyaOoXBywj7Kde5vPXCTv2/vn0YQLZOL8PHeoAT0MkAWrBG/rM9
VrQb70Vc5+t7awGToQ21LEsP6+NGTIoXRXakSMx+i4EnSRlHKvKLNO/geTTaGZe9pZiRr33AhRTT
Z3qbDY1us84330LkdHSIvR+EJ+/T+jimFeI6LnXbCnZzTtsZn4tndiuNYagBED6SmrQHeU4MSnOq
IZKUWO1qWEIdsQT30u9goj7SP7KovGDt10DoOBKRNCnsHa8gJvJy2gdkP/0npaUIKXaR86HuQrkC
UEizUxmhNnFUdg+opRZPWre51HL66FHmR+MacNaEHi+3wveFH9LzLqBQuCn9ppaHhPdHmlmk4g6D
EcrlriRVHzG67qlljT4vedzEadcf88njz+4QEymHWSaL2t4bslHHDTFVHs3ibxLcrDhRnEwBuCfs
8T6Pd78HiX2vHRmL+1esV4t6pl8hszeLFnW9lEoLYy98XMlDJhprpCYsQkgDUVITtwickOPczy7O
y+zNPPaeShN8xym+LlE1ZGqbh4/1khq0w5joSCTK6voDy6zj6jVWsr8emYsYKdlfFKtctgGivPjY
CJK2ECHxks/qIjTQKBf8MPq7/oCM5SBM9TatCWr0077VBYNklN90Au7J8/IMjhoUctvokg23s+bm
4B4v7dfNb0TS2akQulEWzt3NaR0/WnYFAJI13xBUO/4Q+RkevOKLQ+OhtX9hutKS3A2Cl31ZWAkU
+uEXtzbGaYkUYOyGRImhg53/3vlZ2xTjdUJayLbXSAa4XlHDzq+Z/MBR8km2wxqY9rSPFGIlOU/3
rrron1jC6TZ3ueb9T+IwJ17XMf2uaTInhwqnXUyda8M8MHQaHELgCI871SZB0fg0CIQXoxvFfoLu
OtN9dZaPqG0HeMuQskO9Apisjf9xh9nasoWxgac2Z9uucb/Dcz/X4LMXhncfTRfr4YobKREJ5Q9i
JtGiVGMwk0LdioWD1bDAOaqXtlOAHaxuS4Vd6yfSWCbOovC+dN42mGKycQDyexkz0PVq/pE5OV5e
uXCZW070uaZnJpew4n6Rreck/I/GDfhIIXpcfXQXEyNUpswhWQeh9rtaOjRP1RnbC1QjpPdtm3XA
8hJuW+Z5i6BfXSlXUrfHVwwwk1eRVowEZxb2hJ0BU5W4eoKN3borCGshsOKhT5vxpzfxpOM1zDym
NfZZ2q/MNkvYKD5D98Udvg1I8FSXEW2IZeYNpAW+Q3bj4wm2s7J+NczmHONgldoNknMED7IovVtB
Hk+OCc1mBW2uaG+hfQOROk8v0kgrrXQWy2/SM4643xYOZApuKbcGwVvuU5Z1AzpCbDllCG+a8lDP
3QTKzQ8m5ZSpceGUynbO2IKHo6g/plLRVAnD5OVN7Dx7o+DOlwPuabqMiTiobbF0GDreClg4bkav
jeZtnzoKUmItyP33dx/sMkP9u0AFHMLoJb4hxOAL6yk7YHW511wL/oGljxWkIGSiaLwWa7AsyPbQ
PjXZrpUqDmfeMZr2qnvrDq2KeRytMfb529N+Fho5kHaoAoULWIos1VBy9FS2ENA+3RiAgajYj2G0
Ahkf9ph/TP2oPgSxCyZwEcvn1OoYqRpB5JhwoPSuQSmI1b5EgaqL2QvmnkLT4lBiHgd8l1Q28hpT
v07evUqKcmlF3ujdnp0Sffh+ltQE9aWDbXL1gTPx7r9t2S/OmVYDGRX6nFIbjLK++zSGzVFMjdCM
fojAznXIjUxQYJWgcmJfK+JBxdSFrUHKZzZpM3+TKgErCJ6TO2w9fCMc8iI/AvQscHJkryudJ0jK
0GY/g88OhGqLitFygdTkKQ+/UhapQ4jfDyQyYinu0lrGoOMbI6LGFhebmYhG1OS6lkSpDuFwm/0O
ZJfcIf7rJn+/lBEdlBuBlQdFOfXs0iVGDxoObLg0A4rD0RzwJVJQ9Oibw2UywdbcLmlqTugWoKUJ
HPLxa7xRaKBrRIl9xS76eQipiS72KvERG5sEJFfQY/TvJh2QWOkkDBd4zITMxOT6m25+Fn3WIzH5
elRVWSFGkfmUjVuEhdaqfjy8hu/Vjb7+POiWXBMmAiYSJ6jzR8KNkahPXCmH7QixKB6LjJQfJn+U
PHENECcKA4POnTSa3hOvvFoPdvSKhaEWGQyRJ2sCUhKKjOMNyBmkDi+3EokCwMSGnS50oa5w1NUV
RjSicb6p+s7t4pN0/x0mpwkDeW9prRruxmYuBu6IrudLdZRETXkRyXepsDO7Ov4E2rw6A6Yf5uQB
s3o8CcCv1p4Ps6dT7yJZ/Oyo6rDK68CPVHbUMoHr3+fycftiPEKvvctBEpNpCllOdCzpfsVXZv6q
uFDMiwpUDj7LeQfRa8gAV0hpH19eLOPMfjbY9GIgUkOQoCRUDHMI0U7fWG2wnzQKIk7T0sUjUZW7
iSiIlOcRp9le4g44PwtW9WHJc7phRm8yuE/utQuGiFaICywZnczCspg72C/EV+NqGlU7mRJUV3TQ
xWBIu0ZmhcWdU+zZ5fdlOWDvyOWMi2EAJmgljO+BQhgJEkGw4UVCLmLzIpy7iMyiBxRM0BT7v3vM
BG9r6yoP8g4xtaFu0EuRUchyy98SRFuG6+FImndGWeKBP7oQwFnYFN84HAu7o0POjmFPrHxw2HHN
0cut9lNOZ0kkhlwVqFN6Bli/pC2LYGp5QPKX4RpVvHNXx5CG2JnnRkndwW+/Y3AxZeOQ5P1h/zUX
KwMm8TOO0OtsSDP8a3GjLjNGvAUdQWjcBp7vankNjp0flYhXr8Ac4G5IUlkL2ozKXoiCN+RFX+up
WQ4iqNMRBSvg7IBGSwbPR+UYvTc+t5i941vMJJSSerZE1GuZZS+0IX3zih62EVqOJtKU7fg1A4ia
RZjDY9jEe1dUz3KJTbabK6Yp6pMD3MAAjmrq0NS8IvnXKTE1WRmpb5lzlWsT3JEjefuz/7cy1pKM
FRScOXh3HF+w/Tox4SiH7gT6I42y3RxDBazLI5p2uR89353oQW2F4Rs7o9LWUrFRjMQKvDnNCe6N
nUiKVLIdJJmoHmOkXbeRiR54WrvAQDliTbDVKhXLqwjrbr25ki+EDBIPtKbuQ0u2QNEZHN5ht01Z
fUnRN8Oz4uH9ho+ATkszbIzG2yg21MsHsZjnYlN1FIHPQRsvJwVeB9Hlx8xaUuHAF3PkXtNxlXiG
W/e5Vertc/cw9tjAIRQUZaJwvFS85cRPqE09JTkz8zrXYUFFtGPAh/hoJQoUxEd0ro+j2rBnoMaa
gsdvkYYwqQ9vQQOVfBxac31uOdQGu52jEBRkyGN4NZV/bZhBofWjcPfrnEDVbVCwj3fQ+dwH/NEN
2En9te5grVFxI7rXw6kOswSuk5i8I95W8bNsszh1b78gz+Tlsr/CDbU2pH/ng9FAfReoWnR/W6Vd
KTC9mW3GAMeklKvA1+2ck/AeGv0J5UEFxiFTaI9tfxt9RQdtPPxDit5dd9nLWe/5ZoOk5cZjk7GU
KE04tnhL0F10EXB4afUD/L38fqn8tDcWEitzJkrVLdES4bW7oXTvczRdm7f26ipZgh16FgLVLOFz
C5A1CmAayUS9AZpqaFFAHST79zaRkmuqIkMBEPAUg4OGNtjC6ZXjurpeSgm+UiZgP4NM6P110GN9
mZlugBz9prvbbtXpPzDy4TAcjDbEm9+0cA90wf1El13cli6DsUTtkwnc3zSiGJzGgL8vlkPLpHuP
1mw2h7F22vw5Od858YZtcOzzOWDa2M3MPk3tSi7DmkEmqm1yT4kJhkMnPjkoTrT8QReOA5sijtwc
dTP/tGk7SocjZI6wpKTuBxJBOA+jrIkGuH7GB6LsyEfm5wM09CWq86nSrHwbolLfZ1d/um9r5XGO
TSexOAfQ0bYx+nj0z4EQkPWlCDy3GqnVfvKPWyhFkKK+B2l13FL/rT88dl15LmWr+pJWbojLclNG
1wVBFtNSPOZxAiJ7BnD3NH2FedElBydk/HhkXSOYTbFGB5O4rtNIpUKs8aWnqVE0BaIIPpOatLr0
tV5Gr93M8w99z96G1y5sBdD0Jz5LF1BWBrCYvsIC4hCXqOPbSC8BWczS1p5b4oJBLqt/cvz0baDT
sgq9yjOoVr+UdifhaRKNdIcr+nKrov2SrClfBCz25KwUtAPhDsqDOuVv8tDHh9r24wxHNo4C+6as
ryAPHtS0nv0k7Rt4Wk0SxPRRDMEcbFF5odnKLITHV++1/BtJTCZTlZRFFc5eCS6r1hTtTPFiHwDw
aHrez0sHgWYVEwzUlu9Rvh8POirnRa+kEm+r3HJbmhJmCQR64kSGWgwP+tVHe/JegyK4m9B+Tvno
rhSEbYFB8VbatO6MOftJK2c9w/G2zOYJyVap1yAh6quwI3IhCbfzvvPEE2BD4jrGAULq6ycDdgKB
Ck0KsQ1EcdfcOHvJNq9LmRhIz7ALf2CGV5Xfe0un9qWvwc1SpasdOuWzr/pt6WKM7umikEeL1EJ7
ALS74kxG9Te5RSY9Li0TzPo8uGAkOZraxwo3mvhmunMangT6QcQ9Z5N1AFHTxmu2cm4xAL43sMxO
ItAGi6q8KbxGHceDuJiY/KurPpZjLCcMr6uBLrtz8ds7LtxGa1uWkBuUP4KM4R9+ZQ4QEgDGDNfc
CFFPwj5PUk2/53AtAezHAoj64a7iQ9wfjyzz37lYpdEXfnRmz/Yp9aiBHllVaW6UiODQ68Ty2nSS
CYPjQzD6DRq9V3KaIreCsZkJ0mH/LNRluerb3uKW8K+eR+ms3+U3bOhhWvhjutnlpoSJKFVxe551
FQAc7X+6llSU65oWdVkDeoCHVwV4QF8x8jUCaUtWjY/hZeiBgTfecpyt4PsAPiZVuIWwLtCzUu0o
SmgI0mvOGHPki+Y2H/lGwXgK34ZKeIVEDuXfDM7zcbpg5L9y4qK9lQHWLakjuhcOsmfiFCCPy4xa
RG1wffRpbowYVTJZCmu8X90EjQFx4/c0wjYhqMEF/Lzqb7UBVAo6t5W54xzmM6n4B1FZcX161xZM
MWZlN9C8EZOIMbsR1e/eVIOwGxa+uwcOc87oPv839nN9RkYOiQu/4NMpFJuJJbiHvOlWlroKT1b2
0trFewtfFtLpIP7svLyt9K7KLr4JzJmrNWwg55Poqn/egLUW3+s/LjPrkJdVwLKcl26V9fnWufk9
KckTkEXkVVfvMAxKDjPRMMkZFHZBKnGlHn3wWMsI1InPjn3d25YpeLZvcZ2hdEY44gqPb6nkGYqJ
NzqzkCp1G6P82qb1MHC0nL1cmTWBVt26GXQ0Vpl0bK07E9ZqHBLuhJ/eP06hvMPEcaHGN53buLMT
tv/rXIrCb8teYhSR9GsIJokslm/yI9GZSSkt0P5gPIpD0GH+4waYjVt2V6YfMI9W5QT79En/vSBS
aJMdIfAVmJ+B57g3O2BNlzv3ThjBqjEwv3qH6xXJSsnYF42GzP9fVrSUf77KVzr+S8p8eQT1fSML
Rkzn51Pb+RhkFCjVgNh+o79HPbZxDd/F5Gi23PGqZN9QH7pgMSjaFfe8VSIfTp1t0WaK5uohH8fz
0xYpg0PseN0BkKIfSWDgcOxqynj7JVxBu1XiN3ZaJmBIRrpWna6xf+xWWNjRuJUTB9OzG9ksAYLB
QlhXhJmU8Ixpj7P/n3SkNDzfP3WGg0UEmK0/yeBMCkMc2fy3On0NeuA2lLfOb24uLAZR8MM9rAse
McLXcilcqCXePW/zTOYBVXSIXYPPGfJhfa5GqTQt2KJzeC/w6pAdQBgk7v+cWY2IgnrTdkbltbqp
qNqb8+QRTefUy9WBYuptF38RXvV3qv3IMyS0F8Nsj6cMoZZd4xLIRLvc5psdkOW5m76mj4eBbch8
svu33g/KDeR6Jp/pxsfmkIFIKCo5qub2/GX3G/XHmhtKot7HNIo8Jy8boA8V07Ik8ZhSCE1GDnhb
6zprE/DYSDyNV8xTGvzZSh1ZeYKArIZCKwMlPTAWlIFds5KKEbnc1ZWvlkw1iujRvadD5QKIPlTm
AufRqHuKUIBwXgpHOlP6Zs350xMyu8vm21qIhs0JU3s6UvcTrhObncuSkEtIicpMzy3uoxzqhhBB
fQ/IEK7QWgdoGq0najviBFmfWW6wM9EtkTLsXhZag0eZj7Xj5Zj9qSUBfkBmUt/O+rD/tbCIayg3
ydWJpEFaZuCKSM7kC1EYuXH3DaxuH3B6NTVMLLtQ7eBHFh6/9ghVcGOvBqS33vyJ7ckNbdBBTtw0
rnQ2z9JTcpQ2xRAtPqcL5rGcDkIXsBa0Hyz7njr+gDY0yMYhqwCTuTkDJqTFkaCvVQfT3eEfHKSt
STJEAvWpn79sZmOhjXwAyUzwyuYqNAcYBeXedQrz8A/z/hVdsDOKU90w/YTWgJTEMIJmpdymWjYA
rQpkHSMC7eD9/3VwEq/kggqWr3ZwJ/iZHckAZMqkUZ7+JdxCkYBcBBaO7hLNdV6jLSZk88qkmaSm
Rg96Bc5oYXreEifelNN+w9+VDRIRn8vWiFXbBqmvMS/+wABDQQBPWT7eCPA0Yqnb2zkNF5pYjkUT
QezRriZtXRvckm4r6Jqys1Wo7jI0tFOZl//ZL4iofLWaCq7OCkLqovst179mGvmXsWAYil9aVsiT
qMlZHRgYW499A+xOFIQZ4Yr4NVz+ggLFINMlkZ82U3T6fP4lqbdBJf00NbEvVp/4Cy0TeMdHuRaw
totfbAY8Q1x1xO2ikGiPmV5Pv1FCCVal1f7HEBxrONU0VkeDcg7D9XgIyQibFxni5WmA+3BCkDdS
8GUnMJtayDtEmz70ZFazhhdkzXQyTNc0fqNIscaRVVsrGiPPiBjVSH4F/k0vXnGafRsy1ZidwT7z
65VosdiQbA3cMGJCixZ6OyW1EdzBHS3i/fswsvr5YIjZu+TKxMFjl8k8XJyVb5FjbGBLQW+INb4r
Mb7adHqwrvcjaXXJK6Vzw/69WUtrkoFxUkI37Ly33p3out3/fvbIy0r+fcBHl0ikZRH4BBUhqsTj
r3f/608tEN1RS6RkQOov9k2WKC++jfKyN7GNrbnnd6gLUz5la/v/ze/4idGeQiF/QfbkSuz35kYH
1wEEqdloXmY5JVRsnmcI9cof/zQ1zxXx0gh99Wxn9U/DlgyEVyeGF5fm5zpRDT3MqbiJz1/kF0Us
1wWrN9t9pBQROOL8eHvGgnLg4BorIG7BLmIgY3zS2Ti3n7syrTo9EypuA4mBbbKZU2wQUDgOxomD
5Zf4WOeExHd/3hK1guCmUfuk3bKPatwkySl1DsdPXPVfnAGsV3nZNgAvfMD9gJpCAsrE79GFbWp/
EVlPj0dj3PxS/xcqCGuLnwlJkJbzBcKU5oOV6jw8ZeLZJy7gkLgmnj6yUJBIVsgzdwolU7Oxspch
N0uJXJ8AJj78Ph6RXSXSzGzMxq5UYEzEv3HWfdzoMJ+nq2gE3r/OixoPlQyY+kU8i7HAxAC9Yhj4
eIGpS8tPak90Y/VyzyHr0qXVXgYWRRUc2/l7wTSg4IH31cTDEqd2flnwyvBubqOluy/4HQjti07T
9QPBV9PPR9IjKtBrkkR672V8AJQEdcPidAgGUVJMlMrBYVhkWmoSo/cM/wG3Z12c/Cpvkq1Y8Nkv
siRUPDO0tP3MmB1UlmCqEFMHKqXrAXJDzux/aqs32aZUUVyyXROtsYnssY8Z8+I8fgs0zbif/f00
/bJOjjZDuqphtnIRBnWtfwciVVor/D5oz+mSyYbckEEjqECGz8Up+axzWF8qZE9+Yh53et92xHnz
Z+v4E+tul81rC0D5SJ7kW2WmS6VyPbZRzt13Dp0HOwDSSbuc9f88AdjvOdG7ydXc7cF290AOzybf
8DKrK3j2DH/WSlPaxnpuXFsKPngphRDfMR1ZmHKwLjQpINiQ+4k3bU4NF2EKvDVQ/NkOLhcMakD8
ulMJK+LMx9QEnNPfeNFxbRZhrF7ykAv3Uje/R4HOFpMJ8PJH2w+5RGOqFUWOCOVzVIUcO19xX4m5
b1lZwXVkHq/lUqIecYWfiNhkg3YJ6z8tjQlLne1E6SCWfSUrDFzELunkjTJwE8C5TQxRC4A1tYI5
TxwqHFjezawsbUWCSPtFVLzqQpQivsMwGB9Vyxxt7XAoW33jTx7rbgFnIrZSFCv1XCNNFPHLWtji
8U7qdL/iMGqtQ76aRzzMs8PYOC7rkqFf8mffhZ7CBSGHfJ/cY2B543E9iW4Jc/7lIa2AKL+YGhAO
PCg30v/JI24FaMxPEa8QzbWWayOO4UCwolGbrwNzKx9/lBf+30O3UhjtID5Ia23qxQOUhUMTfMdw
nFfOsrfc5hFw5eBoXEwiZEEW5j/2aHJl5NQwgrABfSEMBc7mLCvsLEbhEhmCpxdb/I8bsPObs4YA
WiyBxg6zcPN4q5gxHqbM6CaxIpOhYWpl03+C3TeWgBX7ng6u7JxXJP/tDpN8m5OyiZ1m68zSIkSM
3uf4lRuZA/0SojK1NiNpKy+PGmpSgqvMkJYYtiRjpM1XMcOxcA9WpmgAQiNi0O09MIacni5wF77L
fiMGQdAqT/popYmdxIUpF9Viu5q4ZLAadZMc0nBbec5UfwI1u6fN/GTFDlcaHVOHzkG2CF9YK6MB
ADCkgf0+5qAYAKMo48PL7j4IkgiUNQbMBX3RUt7347B1rJv8niiMP/apb3KCzwBRQPn7gSyBpxhU
AlUBoNyzlcKEAZz5cZ6iyySgrBBQWXdXWW1iKuI/wp1BubAg9GwPCPaAZllhYIdYh+MZNEeSxZu3
SY/DRS9BeLqBWhLrlx0Xv0rn0flsimepf5OsOpg3dxkau+pYx5oQ3HlrsgZar5mLRe4p3d88n4Z1
L9+siS0a7DJ0dJAyvldr4suQt7juBQWZ9RkwcwmNTBZV3xejPNiyjVnUPbQ+4sc2kw/KxlFHjkW6
iXxQrEQTuGc7soXuOdciILochedHCZ+lnUOPs+HQ/X+Kbemz5fqGLM2L7GWxpmLmemNct9Or2nA+
ZAc9vARqtYBMqI3bXmCYs7FTgeONbeZaf99gSRt3WWwERfoKFyZqwO+ou5kP6Aio/TyqghsojTu8
Y8EcMYWmEe6dUvEZcgjz5jVCyci7egzoLAPf3r0RYgWFxRHqEtjKVC4ZjJYWq+hrgPFf8lDe1Kzp
IFLfHMSPbkYOrjLKf2ytGUhdXResmMZR3QkB8a8J0tY/XPsbovq81+4+HNaEbD2046wLo3lDYa48
u/iOb3C0j9MlMtP8k7AEwgNbwxPTlt5pMgr7X3h+FzOjgi/LhKUslDz8D0lHHUZbsHDFDctszMc8
zItWLiSuRcADIFD186P5zy6CzAYjU0VF58nXBtD5HIWKsHPEKK/PHZ1dleyaftm6LzDaHWn6Rb9a
4UHS2pt8Dpd79XEVbb4z9aMb31ngC2J7tEL1PkEz1fNkZbavOgYrheQ10V/HXS+n9CsmT5BDXU+T
Hysq3GK2m0rsd63IFvp1zXBzJTeCgE3xvs5rPJgUrJfbBa2s9520Pz8Z+JEolGMdEyz9VrdONU9a
QhuYhYvn/8cuj6w+lnJpPyDBhqRmOPcDXuWVyqgzTMHnSqZ+a7WV/k3vqi6xBv83vqmk8HfPCbgU
8a1+Z0AU8lBy65hScBdHmLE19FcizNly3dLizWNcb69uqcH/3GggC0oLNnGr7kIaQYKAFFVBFeq9
yeknJroNl6I0cbb1D1yWTrCOm/bCY1bkKsohyc9dA4oz+V2aSjsO3d/wZO2syMTwOFS6/KDlcInq
KEPDHG9Fa810S45MSKt7iEmDM9gIIXnOa3+syWyImfDH/EEKeWNyBva2GNWeyNgAg4pP0Qgryok2
CJbuvxKhf0gXPnShL2NLw7qNHrddxtCUcpvo/nPQbXfCmS8B6ZMUpTlOr358DRv8W8bqH3BJd8Py
vgvsfyUsO5xiIKX5d6jh6tPSDz8F3ZmpTK7006Pirt2Cf75vq14nCOk7e1lpiUX8Smu3m6n8gFNK
Tf+5hN52YIfqfXcSoU3PxJ6IPx3Vcy+uNF2ot56f47/BFKaqdPTYWUuQIZKEuz01LAIlzmIUSEsI
yNKF0pBqY6le18Oecb66kMxcK3mNnm1IvaNXCynklIC+Dng3+aWn2khIfiZFPh0kGMDg2fhE5+s0
tt2XK0wcMEUVVcPKKkLTT5QBDN57evxUiuOXoUI/pK4gTICmgXriuwfHZ7XRe2WPXnX9oR3+5P28
mq56z/b1Pouo8O8y6BG/mmrhfFJlGTpl29nxbAaRjFDhHnrEFotMTsGbDdSeMLQWX+WO1/cLTPbJ
f8duc79y3sIznwYiVsjj1o34tJY0eRjkw7AEPW6cBmtI1/72ynQZPqiISypKdYj299wtRoc31nH9
11sJylGz1eaWSE4VpHaSgQ+IULvtxPaYlG4PcZsGVCB6dKLvvr8IyJmbEPG+OGmYcLQ0HUfWziAd
SFuAKJd77WSF+R8TZ8LcrM6ExAVYwA1Y4BElyOgB3boc6NF4ROwlTE8IVuyCzBLcRHTn2JV4vXLV
jW0+ZAaLslzM1ZsKO4DkrS0zT1v//VjM6EpnmA6CBZbFSotY2+XLBwwC6/ss9LQlDWW2cuSYtOMU
R6JHgwXK+ktTdQGpSDMKa2uI4cWZ4jaELIQQvcu4R2DEylzgbp/8M2Bl8zGPm7XuebVLok1rgYW0
q+KKCBRlKL6B8G2SPb/N2K7nP/dKoxfjTd7jLmZKM0wp7IT7OsY3ABDLiqTs8gA6DSnPQP+fIXRo
ors460ohtn80yep/+hZEz9BvTZzAkmQO2J0mlO293c6md2/b//iyHqIJGNvqnjOWqrpUJxlNfh0U
j7IqUgaZ1DwxANrSn1UGIcVb40xRdcHoGoh0WPmjCjXSgMVvwrqew81twCM6v8084k9HSTnvTPP3
UfFiEh8WZV5GdtxLAX388hLJURlmoAeKEZotoh4IN+R1fW+3WbKB9KEtVsXXu49UGMCq+sScQyeY
Dh5tXxZ8oTzkY8i6NTaVHRCzpKonmAgzv+SVZqtSQb6uORI59Tz64e+9iA1by4j5zqvVQPknmO72
+/HD+8EVw5azAYl9oEMj5LsphoKWp0+sQ4rH2JuwO/mP95kTPiWf1GXT1UptEmVa+tebVmZHh8+/
LCGbwQ+qZ3odYJUHrw1hY7bUd9VRjVVdtClZhY5/YeYnmvKyYNS+g6ml9lSdFL5zqcuJFboDg8Xn
iM+KVtyU3V81xftHC2CeUET/479u4aTMekSFrgX70yXz/6zNkblc70GXQMITMbeCbIQHQtrZPe9L
dMHXSTnBcwD9yEwnGHKmQhgQ3rB4sRb77ukPkuCLJbttVGpBZScE0CSZyoNHbxNwRYjjiPGT3UBH
CX1jg0FQWchZmqHMq57ACONlsttl3GI/J+RUlQuL9jYO+6jDjGe2bxPZB4L7FNypSp6otKj+Fg5Q
JRzyeu/MQz5tvCmi842YYytzk8yaQ80JxjCioJevQDOrPMBpcDiaZ4LxKuKJ3a9FmftN+FQ3wTkV
Y8omBNZCv73adWABpoxgLFlUYgxjlzlaxWugJkpYIZ7h1Wj4nufOeKQhYckhCIbwK+MD4f2aq0db
O7lRAtOIaCNQT8lCE2juQ8FHaE0VDQzWMvL1z9YnzMDC06wNqi+jd1l53ggWG1QYRaA5wMxA/lxT
AOUit+wF8FX5bKYMLawoJIbeIy8z3xU7bjztrnw77hQkqVr3VM+6/gQ33/8TopzMH5S2H/rWNvOT
ANOD7M01/FUAXT8k9zNi/DRZ5HkFOxvWMWibwAOMdcXPmyuMwQW4GTTy41QoCnsG0R342ZDfQhCI
epThlZ9AAmxiMfyHC2JQAvMrZGeDHJ307ffSBPQUF2pj+hF+U5d42YFglMUQCwi+slAH96RdEtZB
fVEBAHGNaWwFnSsKCRYY3+6NRpzrdt3MtNATxLSV9tBMjBHndQKRWKzwH5KBcjeyDtZjWcrb1bz2
378/7K/xvficmvBDu92CbP1OmW203m4c8BkYhL+lXx3LbzgUksckFJk1hJX5ClICGJUl1iT0x6VH
kmU/2PTZJ9FHi+BGhK+G2hxIdrlhgDw+yx9ynBped90MlQ22dmSlbpcHDxkB6Z7HKNYhzKQsxAvt
xjYaa/Mv/1kyRWXEs+F8uqmc9zpAFdvxsEnDCb5/qbCFl3iIzR2f6bGodEwOto6LFAfkevRc8vSd
sa66g1ru6I6XacMUAh+Imtl4YnGHL0yZH4X0O6qtuazHwZJS3VpdNh+ILWsQlvMViakcTf1k8/VL
4or8R9ypALcDCpT1jj5w1e68l7HefQ8jAmKJyMpZfq4Pb7Pw/1hLUenv0OM9SigGjUUWujJXtTQO
KwOBETLFbnzJXepnuybWYmfYL5XQ5nOJ/5gu7Q74bPduhBMZPjsEJHHfjQa99HIZFNT5GHhJyVEd
OFSmavhKiIbqUWwR3uJ1wr9SJMQ8Aut7V2E9xAkhbvxpzu1LExHVh/mOudwYrZ2L0c1vuNgEucRg
YkVb1NJtGzo1Ks8l3Hvsdzfg74Su7DlzBC06Y4EELOT9dJwsHGudXzQJRJAymu26UasQRMMG8t3a
KQHTgtVo5f7NPegYvYBDPMtvxBsyfBqCIM3S/8cUiiMoUzRMvHmBK1cTGV0tFARK+4TvgMKsAML0
caBHdDbsX8LIPbJ6+s/lxvAP/AvW8C/3R3j8QlSevg4blX7NjOzh1ATYmT6ptb6Nby3zMZtGbpS/
ZcI+NcVizKiZ6+rqnWue0N+p5sA7mqcAYC0N0pgjG/6fTOEuHmiINwF8x12Ltb3BDu3ozONGkPuV
oDzwxz9ewAj9SzLOxOpzPZAFWfKitf2J8+bsJQjdsKUBl6MjLrhhUhkHooM1BZ+XqWaFLT6KiM2A
El7cDcj2NHG3qRMUaPMCOS89PeMcNCR/BfBCCh4nFAyprTmC+9HDL9CbTU15/AocnK9ZEQazhEB6
ZrbK6JQWYMro96RhQyJ/kzka5JpoOfGSfxocSGLV8JWAKJ1pgeP8fSnak1uyUwcJoQ34hDmENjGc
cCA8ZZ9uqEzdc4QKg0jYcVOyKxRrwZetxiOR3MIR8IZBw8jeQtUajHleNMv45AcPmpUc2xSnDdUr
ddk+oep2AKL6Ii3Yf2bBKcoM7XgVB6uuypH95FTV+QeIB/iEhe6wDnHtm7IfSRPV1Qpa18foaQqR
aGDNIukQwEFyD3mzix6xj2rmvXKBUAvQJpdhPxxQ30gyvfjn8EkVOWjW+uZf5vKTHXjwXMMkqFZm
YjdEt6y9y/P9pwAdv5evNnuWfjJfUlxoIFC+qLE1evmwjxdSEgwMucK+ziOr4qtJeKJAC9WdB8ys
6dLMl0bHxcGT+hoiED2ZLdMiEslM04seOmzLbvyW0EMJlNPbg9RWJ0ZhxxuV34Kf5nKB6moR+sGu
utqqgBXwE868ue4yKabOuM40U4uZQArPSwunGWKlh6PfWhKhNCwW9HZXt4C/BjHUv0u+iWDZPYMs
eJp8Qgz5qG9Ysm5vcwWO4bpc3R/Gyadb+gIMmUIZCAt0GX/6x5E1ezf4O/lJYOzXXaEgw0cyBvpo
4AGgvxpictFdhYrkBpZmEQHCBoTrFTiU71FBIu5tfGUaZxPUkozmk4r5kVoSy+7GnRxXRF22xdsF
E4zqnHYRtqaOi/a2JX50nV+17PQEIF3yf9fdXW/Ogrzo2bLaMesIOCoN1MdxFtMo7n1TIdEE+si+
tgdDrKri1p4sQDeuZg4cZIO+JFugEo20Hqfmd0RJpJP8VeArEiBP6lgoq3ZfHuxP2zE1irkO0D+x
mMSmLWchLSgKxqrUDr+ooG9815sa5nK5cDAla49dVB7tmLShFP3/UBPxuOymMACRPdc28lUAFSaB
Q88xVQblW8xj978IYXv3T1QVad+DXhTKBgx5HRR+EX4ZRz5Nw3qYUYW6gBv4OYN3Nr5fh+7b6jFi
vB+82JsWX2A40ApYYTXidbNSdOXoJ1+bCxGOpCCFDoyIYIuyrEi2GuyrWpHJ501re9tpe1fLJmwL
6CIEi7VTL+Uytn0I1vJg9DmpoNo07nWoDnWfR29h4ZoETJJEFvlVfavzZWDb5noagEKjs1Ss9H8x
M7LjPbWeckij4SBNhv4cczIzdbIloa7bmJcTAxLN17EF6r9wQs6w2d/X6Vq43Mgth4SYvz11AnZn
GPXeAyjEuxIqGoMRMHi6dMUurK2JetRO07nhBJA7gSlXBnR39ceImPBFpWLtsuPd/daK5doEHt3U
hZi18116LYRPM7Sx+6ww0b6ROIy7pFi8kQFBCG5gPnBHJLKIPyodhU3uLOcHFVoFO2NlmWPKx6sn
tjQe7OzbuK+VufOOmOEQjcmjktxnsrzAm7gKNZBf18QedtX1QPC5Yly1ZFXO7wQpZiZ/CIec5T21
Q5IKHXORg+ROQtBMN44S/2p5cZ4ySODxDymZEcP0qJz+cpqeb+sfIzB3VAvC0eeoE6TA4REQsnEm
uXb7KvPBcXqlPDMkLirGgtYC0kdAAARJSCCmzKHqTtvLHTYetGO76SbGEhph5JIz3gK6d+v5Wjju
Jv7EgfTjMbWuJfPMAjFRmpsu5hem816J5YKQE/Hz9rbCgMK/kzSHrRaxyyRZqp+QqWzCp+2HfndB
9ill6AW8//mYyM46Cvgphtr9RrsXxKvjkAp2/ipttryyKfbzIknQ8RRP5OKf3d7MkWgCe2qiPRQ3
SrpfPZtdxcc9jHZBG3J4snnu0aSxJkYWarBeh19WRDNT7GgudOx3KdRObx5maXbbnNT+Lt6Y6uGp
TF9ctObrTyPXaBBZUerndL6Cx+t2uX1xDA3YKWcdl4ctTQh9P64X/zZiTrKudkOYz2XmJCoIW0v0
gfiC90bVmsBPkJ3LOPaGFyPvfC+l2zSpcGuQC1G3vqlQYZE0eL11urEPVBygEie371UPLUmYQaja
z9j+dywUGxCA0PGY5wnI5AXuon9yVX110UiiUZMua8hti8Cb95T2bbrkjyygt3MzIgaurgm0izRX
U2z32Vr82Jpi2OtLGZ/zWF87prE2yUZdf68dT274qCCOsYBB/0HVtX2lyro3NXoq4DRtmHPsLbTy
EyEKgjZq2Lkpxq62rwdXnqvYlDTH5AjezIoo0MFK0xyu5Xv7SYWXzWfKoX31/eXOmd+mnLjoL3YT
Kjaj4mnjlHIgA8JH82fhxswTYI108oOPaTTtJ7dtI2aoCKemYkvnykvwLL2/pg7+VS1B/ILOg4y3
MVbSngYZM25+EuZRC74Hj+9jpZDNkstpwdmHJKCXS28VznuXXQRanIhAFfnbN2USKJiQ6YuzvHwx
iPv7AzXjcakZkDqM10M16Uw4eS/CndzEF+8hBMDWeDT3msY+drEpOAxZVzTEx4vrwtN8NbDw+b36
+ZjG0Rg3kFollpuYzirzIyyzxS0mZODz24f9otjXOHkCcssLyZ2K8ru6ZGtejH90audIUWme0tUN
z65Kr78zPWION34Uf44mccixeZQEj6AenNlaV0NCOenNVguqxBg3Ttpv3AARP0a79eVzD8CLB5ID
vDKUfqW/4zALaHs3UpKCckcYBsCxFhZLYAeyPkF8frrddPbx0onPkjs1LNFsxbWVSER5oxbJVd1N
xSNT2jtvQQQA/zpQXEz7bIqY+AjRCxidY9f56Uei+8uzHGcaXkRxvLyvg7UDBbmBeu6plP+6AuDy
4QAkw8BbcKLVY2GaMqsvfbNMv0GE0cXM9sHFWubt54UXQK2Weshm0iu072cqWOQiETbpHq+ssmTX
YZaToiyCPOrIlqMQ5/9qKUu5a1isopcsydTUx3/PMwQb+1PM8UQ/F72y7bx8liaodd9UroKDWa+t
sp93JInS+p9xTuVcVaAg5YLyRCMnA0vrUpLMhgPHZiDziUER4xd40lY+F0VnFqNXp8QywOIAxlFe
fflju5lfzfwbj4ASFWloCyNN55jQUbhH8oE+dL0FKd+2D1dKLUnc0Z0DDsigMScGnfYeymC1ELQb
ZvKTJ+JWFdRpmfC8NvFxXDkB6LeP6K51jF8cxYMQLWyZhTUtutPvqQgki2lFYbZtt+woh/sEK5Fm
K2B4oZ/B5S7mu2EOJ/flrwTWybRq9vmaBiHA25YmSKsu88vpFWwiOnSWcpAY+kde1YulzOjcZkeU
6Ke8bjEHcypWzv1HNyutwDwxxjymSR/8ER3fYzVhHfwlqUX7hxOu0u1+dbUs2XtcoeWjF83wd3s0
1n3hGFLnu4fv6xqSvc52VyBBEQEokeAyW+Rk8GOL5oQoU9mrI/1uOjQOxo0cuOwTPpzU7KKVKnJY
gkkaDaNgPMip9GkibJ4nWSAF03mDGgiqp+bCFNu+hUT9QcJGhIxe1gqeAUcNvl8diXQ2lMH9vUwV
VrGkOzDDO9gXv30qUJgFGXTRIRDfgsBTVVNGA6/UUy8HLg6kBZnAPneOA3dzvJJ8SGKToF5swMXq
/SDWAdfJBHOAlqL9YyE/cAxesuYnO8rmB0St5yQg3PgyPlq849MYB55JPlAtpQ61/2jx4wsquffz
Dz/lIKI+MGK1GyNrV7YZ9x3RfeZnxZNMPV6pnNY2aX8N4xQ4EDhM6DeN7obkA+6DHkwHdwjO6KkG
pQda/O2Nlv78uEIOD+5s7gTVKqMjGNkZpxtAVdZ/OgkFXCPdo0/RDe0EOH6Sfqzyfh5mXGuvXqMq
HpRQOU7nzDTYpdynSKMOPMk7AHUEXgW58VrIu6QO2NdBttJSXEJbn4NUjxIl1Wmnhl+KIXZmwMjl
aoCCKAMODNDK17uoVjtb0dBoPHNj4DkE9EfjjKW0eT0nDkihbxwMgr3IndiaB/rS08QbWOA4L3ft
MQSgoEmHxat3VYjSK9U9xFboAW8r5FN9E6BMIn+4KqhI8ePPmAqTd0hUBRa2oycLLf1evDmhVT4D
rGoeGL1t/nL8Kne1zQXbJmU/iGt5lngZKBvGHotA4FM9kFqCtv8JiJFL6iqYArqmEHrQUDdMf/WK
CYVp31pbd4EirhYkFq5V/FJH15N4mPqKIx3Vv5ZwVZRZStQowvFfzGg2CMYPvUEOMotqXr/clay4
QQi6DcjZv4/A1wpzV0kivh7r+0ydf27D4DZ30hs5g3KaeOQs7nq9dZZba5ozjqno/JIrkK1G7CmI
1j91BKFbs8z8DSespzrXtYoJ0Az0Xs+eaP2SeedfAIUaPXEtZU8djeY3MmRp0Thk/5Ez0rRwUPAt
ZaylWo9TUgIPkHdYfgq34vwkW7zCWx/LBndpSd5p/AJ7tpvQn6wR7FztZf4IuK2Oz9L+jrTPtZwx
BAcX04evkbhuCyGCVtcXjsvfWRxcKL0LiPTkzXwfxEo3geEpXTwPhqNNNaqWF0i6UrhXV1fTAc0r
/ZopRlC+k3O1jwJtkK7IMytNEj+fYO1luxOX2w/tg3UaZLq1pySkdT96OS0GC+cTgvbllReJkDGD
N5IjI5CZtmx+J2BG5Kq4zllWPF622J+QiTCkkEEM2bNgvVvEWWMB1Jb0IlWrKDeYMMQCd+eQbMtC
yRXYsiItvlmvfT1GMr2Gyfkrsj07bvTUc/m2DRcKBcuJWWKOkv6IkAdSRz7CVhN4Jas4LhJs1gsJ
GfBXOH+oaJpSGXt8+lHWl7UyBskQIdYU5+NlPX2vLmxA5Fbh++XqHd+0FjY/uPhlg/+9EFlhCKl9
oigIe/wP3Dbx/cgv5gkBHls03rXzM+MmyfxkVzQ0SovC0fYBOYC1XdlcZHRHO0jk+TyEf0adFPki
f3MZq7jPKPFcCA3pzS4wHCN4Lg4p0fe+BC65uMtRnYdi8dt6VLAzMlWR4+iUnXABuR+umejcr201
louKiu2gMuGAvL1M80VW4jw3bOcqKgGCzs5czp+CIe/2h3LJ6uP0HOnBXrg07Pp7Ovu6h/ztUjFf
98dov47qJyHVKfkFdMtdhWrUeWAIilonriHW5x5I9Gj+PBP4adQGNV9z8lDNCy/W8NDFBUFwTmUI
/OcgTOjxhLS2gMNLUjyXEbS0qyaLERw1qxKMhOWg8+dN5hDYdMMtwFFvUSK8bISq37zYkZACO/hL
KlzXOPsjhAC1U2M17ByLbRc9GE/5vtqLjUjrc4NWnOWOoBrH+z6GTXxN/JIfmhHe4bM34ZRPUKaI
hBwEcpSNuYzmMOhKwaAJ1IaYLXHFhdxosvDsM0uWYwv7CI3ijt2j+IADQ4k2j0RCqTbBj13BIhDL
xIgZtvwy2mz2wfwjqWxYa86Io5V/2mHnTde9gmRbKxXdsp6xsAVJhauFajpSQARF/HU8o5IjlUyi
Fxpf091HazCoA2n5Gy8Ao6gdZW2KD7MywpdPSsG2YUQW2Xz/3wf3vj7Zzx/IsJ3jGZFqS6jqNYPQ
wZNDLpQzmjyW7cXkQHRlBzvrYVjyDoKZUGcRF7nAA3eLGaG5rBp0F/HwrQOJPxS0d6x8lrR1tv4M
mzy1ad2qBvzr0rolVvvFfovPIZQg/cOIziyPA6+YvK89hPti2aYKNwi7WfkdIRbALmDCvXgEhpHc
Lh5rX9OUcOLR4WgdYfS6bVS5XCsmIAqkb7LkD260AS9MFokjkbB5yonQSIfOi3oIfk49XFqC0drT
a/BDaGCbzVoLn27VRLSoMK3hfTSrQNyPz4YLJRPOIakVfucvmT9siLa6H8RusZ+y+bLIlFVPyAYn
i3vfB9p+Peltb+6GTUXy1jpHl/tzpFa8nRGZm04C3qBmOqv8JJQ2NXtIhnO44t61YbGY9eu6bVqc
CdbX290kcluS72ncY2M9lYUzhFSJ9cgkQZNywhOpThp5H9VR0BKweVTxvpP2fyPahL3YPrIOHUdd
qV+7AWHBAz38OS4bGMoCJ3MAYsHp4I+dYncBRFthgLzjXmvFvusht93PQT76kO0rqowiHR+rWuZF
SlBzOnd8KWHdzcf/ZdAsdYz5o5kSAOj9v0+B7eEn6TDLRd8AHIXwnXvqF8HkiauoKJCkRVNA9/9j
Kte0rvenyMFrKqlwDBG5RPGCus5+8XYdt1ciMdOROWHJuBqGDuPhZ5jM9K2lmPMhY4mUDRDxm/Q5
98BTDPQzLy+C3kzTpiAM94wK8/t0XQvmnJ5ewEC3ytpkf4vGYpKgaj5kg78/JBLSK/OB5lg0POSq
Pym//6Gvepv8zjnj8Bu7cBiMZmGn1EQhs35Xs0BmIQSVpVhLtsdXy2YFCUJepo/G+gOF1O44d7wq
P8PCjKlYEA3/HWram+qvSN5HK7bUh5seFxbj+o5ZzCgHb+AlZMZ7SlXER7NiBy3u8hAJVfIHAJ+5
Pz7eFJigF2m0USa/iEayyEDNr/R46S+GJLNYs5DJVyMhyilI/nfO03a9SVGjGjEW9HheRBfEP9YE
JYIgtsApxxWu8mU2xARiKmnL9HfhyUorMjlBZux5WTLEcmLJzpI5+al36po/auG0lqSan9kVmX4B
w0PShzDtr5aTluKVJnX0spVLs+xw58mc5DLsnwhCDmU3PjnesoeoLlWs3CYIbTn0s4d5wOTp9tao
ao5uiVKzc0W60ZZJh/d3lbd/z5KL7bJ9t6TLIpr4Eep178zD9ncf0tkMPMNswibSq5rENsP/uriv
OJfLCharOzPBTaskcSovY430+Di6xIsYr1FRY85qw6cg64m5GghmVl11CMPDLp+wYw3pN5EA4acd
OOBBy3E2e5BQkME+77uzkwBu4lKSLpfLvCP8qPwqPBct5d9lCu4wC7oqL2A7JqAMmAXtTh5hwDdO
ok1zwlXrlujjd4/MLUKvwO6RFYOi8NHaxJ5yzI10qchbXiiVQ9TgoQ6P5IfY864PHc6iFibTmocz
Kk3C1mhyFREq6f/e4/mkIjUFMuxKm2NYaulKZR441Tl/6qR4XNrDsoiL/BdF4mNeptur8rkqV62E
Dl+gE8NUCF0D8HecidWisjE9FYeERL2SqiLVouYjUQb5Va9xTolO11+ZZ/+0aeIHpCUQfOhmeMOY
dvCJFNoSTZ5hk3C9Qc0t8UQR9j9nhy0Hq3VMsSvLbsNsGofZgfTw4gqb31VgXvBoy/jka9/p5huZ
w8zIcmus8dTbLFWhXrhIrzkelen/Re4z1w1ZtpC5yPBgaY8PvIcEJ0Oxx9zphtReF20jHVFqb7y/
0dppKEF/QAK+wYGJ+df/FUjgn81wugSbJXAEo/RJnBN1jmr9rJ681N4/7RcxgF/WwX/A/k/3PdVT
lI35EPzwO0k6TKQ/G4usg14Gf0Ryy5XKf+RYAOngEN5ENRRVNXnxU0vL+4dnswZlMv7rQ9Nu7CjT
8o8MeAm5nUiBYmGKKfkqwkBNaZFccCwf2uErmPdGD7ywhz1NLinJh7633Jv9OKpR/zy3OGxGNQx+
XNsB+h4X2lDJxWXL522q0899Gr9CU6aAjGUdY5v5V52tTxQKWb1ksvIUWj9jMptCJ4XRshFN/IUN
ewoe5sWVYGP1GB7ceQP0MVOUyuY2VEc/ofzOY/y61eyeOOgAHQtlelcho1NdNBzPBjBX/bBZOljx
KQsjWPDXixOf6EXEE1GpR2woxfqcR386Y0H261x4sjC+z6AilD9FNV8NAvYu3u8ZjTjM9WjxtbvZ
mZZrL2MoBjwSnjsM5e8o5lV4Y3OW6dtQZufHSY9FTWwQKUmavcnC+JNbkd7off5vHfegIDrYILa0
a25aNUEYLtvJTXcqpnasowWYKFxfKJg5h347J55PHBQmZsf6rcW+JGD/tzvFpzqE8I8gFlOJGxSU
IRD2evc9wpfby9o9hXx94zaDDgKpDWJnbyvapAutYwp+Y2Ll/SnDa7WthG91Jo0VT/9NrlRPjdLY
263WfGgM4/b33l60kAQHFzEv+zk6dq//DzoKw9iIidgF1ijvjT8x0MzaaPkGoqnY1mMbj//N1Eo1
Zr2sPLW2hR25zULWE6n/48f5TXs0yMvikZi5H6uiybw1OC8mEowCDLQlzcUgU9a1J4/Y6MveHV3f
lkDVhbgSdBVQDCguEUEii4nExeTDTemzfxG8I/oePYuTdeFqwI8+YZa5V15RVJ8DI1UdIs0z7UQ9
bkvU12te63PN7lms9wXwb2HMlL1J9x4bjYLh66pXYM3+h/jIQWNkjfh/sRlDReDkoO5RYaUChsBz
rL0SPnPjn0+pYlQEacAMjRErdmH/S9rLQAtFwAbDyBDlZP63a9NYb+pW9QJ1ZtuDu1bwDEylMsrR
SWLt9ysNptTZvoEamDF7/lKcNZ/rqumpEJVgNLX/UVgkUwjNxbpkfr20f6jucmAem/vUPxi7Nkxc
PkLGpHaUZSH9Zfhp7helmQEMSZeVZPMuSQIxLkkHq66aRPQZi5GiKdDB1U2H5gs1qQ9TCdkEVtjy
L2XOXiUuWgijQGNYsfwPfsl3xQYoULMMIAhG/iOvd7zAPyLPAUZbsKWNmwrYjTa6abPWdwSQxzCy
5m9RMkLA2Oa1XElC5awWyz8UZDtSbpIu6L6fSDq0AR0eVQE2vT/ErsMtgNxntwYB9VD85GouMHPl
s88kz9GmyODfN5dcPNfXUiPfljhrQCkng1G1CerI+OCiQmmnvnpQ7VNtZeGUK6d52ZutAQecGk7n
OMS3uBsz1F61yYhGp73WqS8zv5Ok86Fb7JVUfPqTrNpenRyULuph+0fcDc1nZSKVqqK1ud+3cF64
ceNF5DJj5l1HCW7SjcwPSHN93Y4f7ScRnHwzZ5I6c7l3jX4WqzfovSpHTsPCRLmwBLoLbG9+khdn
O8kSI8DySps/vQrLht1SAmOxpryTXWtvg5f/+baluIlY8Ax39y/CJjkwmNkpidnxp778q9kkqAIR
B6X3iyXh3yad6eHuExEEFLmGegOY0N7BQNhZUVBkfrZGvRUL+63dqxpyIwNTegKeil5HYCL+Lp+c
QhZON6/ZrVRmSHnG/v2T0RWScXp0UAnBL/arOkYfQ8e/gpd+YOqgcCVXfIEsQTBYxqXtjSBOxxUH
wcKljWvPCu8neVevIOC//zVXRmTzs10ZL01scDVu74txEiDzIwIiwNcAdsVIQTVGWkWjKi2uweaE
Acm704VyrWbwP/8T4ILibPmCGSpzLwIPFsezToTPN7mC2X9ieJacKP7hcLs8uTEDW3/C4JEn5+nx
Bh6530xDDkzSCPz6gz1qVn1gw1YrTD1vq3FaHkgkW76eg0qy03LOAWUpEgR3bsHaPYzbzE8f6g+K
7r7G5FRaZqXceT2bhfIyg+kJ0OnUn0BqgDkE6hpDp9PTMWAFFasfjKiCU71siinzIHb/pQ63705c
7LtYRqHsgBbqD4qFb9X2DkUw0p2qzX0IJJB43g/cEGlcKx0qY0DwKFt3MD6PY3MJov5Z48h+sU4M
UdXV+pIVjralyDmCv2BIO5s8diXY+MGNqL0OOMtdLM8feN9QiiUQtJavBu8EP3+GrWyiKxLLR+NX
ikiC+HCeMDuU8Ht2sA54SrwU97Nn5qtNJOnM4C6tI8DFOnD4M8loT7XuVk24lNbEW29/ZKTsI2AL
4YcHMhlZMhVky1y3P3xA0nciiU+ZugA3XyuI+AeRilSce7+kebd2QdrN9KiCITwhqEZ6wWsNFzNe
+u29asGcslgu8x6zAETzVTP/Mb+QFTjtbKnQ9i9tCq9aEd15f/8833eyYTXI3Z6zyvz3HVb5sWhT
ZYSbLALSZReksedf5Fg8W9DI4g4nFO2t6XnjXH/Jgexg9up/lLsHswoMyEmSUgKQWtQhB+Nx7kF+
/cvJNvuhv4lWaXGWWqN5FEfSKrsCU9H7eSrBCWhq2WenYOCszAShtw9fVH0mFYKdQvPHphsxJHI7
8uiAwpQEmO2KGoa6uNjMDkFngU2RKkYhprspe9KgVTVaHwhTAGLt6Ot4Y93xYwttQ6EPgYlx6ULA
Ojkji8kCOiO5EjnbTWjSBiVwzwtOAOu117Y+c4L4fShu9r1hMz7BLccIHDCFnRAlNJmndGke/eyw
kbnPU58DtCQCr5Gml6RX5Vh/Oo1hRmwpLs/t5QGauBBZj5f6F4RisJ7Yf14uV5gZW/TfqOenA5hp
00Q38KqOHUQnYn+Q3uhqQxV+PXrJR06LWCxuYD+PF+KCKR+fSZyu1jbwDrA24K7i5ie5QlYMBCyO
AVgU50xuNS5+GPfAp0oz7YB98NR3OiWV+0gNRU+APlK77etL5c+PvAq7FLquEpggvkAhXtO+xgCN
WPed2L6REag+XUq5ds9h+hNuZ4AjXDfq5i+MBbGghtYUnGqdfflJVg12IgndOQ7fIkP0EmhPE9J1
ix3MQHbtDW6vRwIgzSns8Uys8cHP7P2fmHwOh8Xf9h9rDv+Gi/5FLsMupG/SWWR6CfaygbbEYq11
jd38w1DfxJlz8RRgqF3t6jD03CZ3vqygcFjX2nQtKwFtjgx18W1THs7618QDISNG0WUlEULbB29O
Y7HV0wBjFiRo3cgDW/Js8hRJyrJAEA+AuHGDf3Mdwfs8l8dW2mSJvuoGGdlZDF8IKRWRsHUI270p
p9OeRvkrDH9y+Xb3FI1f85NpTKNfkAqMR2SVaMlzkmOhXCHFQAB2pWy0k4tF760AWB3JzV0HJ04E
x0SZwm5MrV2UtgnIOjfw1bJA2BjUPY1G5IID1QxPyXCiD8DMyATae0xakNDLyt+WVhZaNt9J744a
yPKmkJ/7JDLVUc0gKPsf6A4iTEQr6EIOFb8wVC12ZaVi6VG5WdBCsiJuf2X//UwqyvOHnhOeGRE8
eA/BGsuG8lnUM/3XS41YRqo1QPtCQq5bxeq0pUE2JS8KD71FNWPzZKoo61fSKKd45/DGsGWSoWVs
l0oMmsmWOD5BoY1AI/t5ARlXEiMR4LBfShODTx27E7sL81wQEU7IM+6WL1eFoy/hP0YtFteGF2nZ
YaU4B9CbtL/hOtqe8mY1KZlvSft/w58Eh6K8TBxlcTS5IrWiunHFwyiHAh4noPJTEt0ilG2+dbqi
f7MvPfW1aV7/OvGlUN9C7VDYk86+UQO09Q1NFiYDtlgO5vbRuaYZmBelwwP7Uu0P0TYzigg+DtSq
eQrZr4RCJOKgH3YjHYU9cE3TU8RdE9vrh735EMdkJd0Bf9LxpT4f9GoDmTGD3j/wfuo+6apfB9UH
D26k9mHqoP9cguyJX52OH6wOLjBpbIEzQK+eRM+2tB9XHJ1h3rZOPAJlzrqYc1D2M1lOafnm79gM
lhplhAHNrdZRtBuFiBTCsSxUaFAsJIuw5YPD07ADH457huyN9H4klzVTNBiVSbXaXj1/va0vAJrM
k3dk1ps2xqc37ctjZZQTYgnUI7jcVEEoVjj6/ZwPkb3nJ7FTM2arlLVEqzFEckXZ88cpBUt6dlVp
oKLZMIf/QdyM8pKpYR9sokBO2TkiCxuGBSUo3RNMkDuPXBoDz5q6r6I0/kBr22bMbjprCuH0KmDX
2tAp/w/R+Tjwj+oZ4hK74aZEiBiJy1ZExW5DKiNnMSxGag+uL0HZOA61NAWsqAVDh/Csevxb/zCo
Ud5wze27QlgjWGZG430Ej+XldkYOAhU6NgVevpOR6SwOgHEeHPBu/sv9M+2X+FKBtJqA/70Z425V
gFWbkHaog9P24hGYKo6HX/EH/mQYL4xYloe5nphYWSaY1BEwkiDcUGAPLnzOUimjMaLCjMsJHHKa
U4ZDAdHMJU8vvIyBYBRxf99SuYTP3xK8aPNl0AE+1qkP/UaPSMo3dSdeg8IJ1y9QGwJOZ2dCgsHi
UOFOJuMNR51wJr4a77ONgwpFhBGfP61KwnRGp4o6aI9+Yqtxr4cNpsqWP4CslW6Bif1dnbX/ttfw
ewjcgPfZXm4sBMwcGCE5leBzFwJfnJW5h8J2raz8u50n67u7IZB0M3vXUOTxgPEUjanwje7lCRGs
0Ck70Usmh+clZQ4NgcYL31+qCqXu9o6zmvR5vwF4XD30ndXedKz2j/8QQk3rt1PhYnn8cEG7S9Td
sz83XHbpYH80wS7zcqImfl2AFsiZLoqbvEfI3snd4Dc4qgUK/OLl0wk97fI6JKyEyA8cEz6fnwof
FJ6CjsHytxx6h8EXAI1ezcYeN9qnXlcgeDbf/eTY3S1IsozHswJEkyeH4H0MacL9TXrBLdIl32h2
7i1pcSkwbrsaKASkXRZxF/tG9/Re/bsJCjKhPhvi8gZkCfDJuJWlo1RR2RGsD+qWEet1xfiN3I2U
K4jkQFKL3kbJDzVEi2rkB35t268CCaSoMNERyaFP6LKoI6WBsN/Hc/RhQY/MYIInsoU+KjDYVBYV
kuaAxxG/yaGo12SJz0QlfIx9y5QJPP8ThRyg3DVVZ/0jKTsmqWa07KMDEslC5G0ua+Q6XuO7G+7C
IMkU5Qz2kqDf8XedKfnJ6SP0MfH5J2Ny1ZprQh7MgSrXs0q8iBzoarOpXJmCjcTJNRoqxH0GLKGs
GDYM06CliUZkNtYYruARHSYs6sIkBdBTo9heTCPM6oFTYRyGTlyD+em7oi76sdZXTN5dBbMo5ngf
b6PvPvTZ/6lMnskLX57eUFBe5Wz33xbQf6E3eE2Lhyqn/H40YZrlvIRbK5DriZeFkSzbGodJhT8D
Lh55acxxhVePpvb71StCWCMJBk0QOFbi37JrkaxPZZbry4uwSbPSivB+AERDUmRJchJF8HD4j/Xb
KSDyjRyP18Dz1+ANnVwE80tMGyjzcoWuRU1GubU2TWPRnmsMGxPOYCiUHnh1+C0X3ONyw5YHpUqn
6LPrxdOpEP6eDe2kclDBwi1NhYUlxzoE0bSIKUk0/sH/2lzvhY9ujhs3hP/9JY5n85ffSvcEL6kF
NUuDwpK71KVzEiethBvfs3bK4bWpqli5ddOFlaHMQnM9IhTgpN/SB3Pi0K9IjEZa2rmf5MXmS3Kg
vJdbvCkTr2omSirsXMPaJUHv7DZP+SsMOfxaTkE742nkyocG8thPHv4DT7RQhMiPGD7mhB4mLISM
h2GMV+rm+aJdhjl2kjqnR4cZwvxRpd0O+obykfrmX5actrH46aKBqEUU7vId447aAHpY4AxGLQfc
3G/02OT4f0Kc2l2kyE1hBbghPSBrQH4Dg+ZcNd0EDe7orEwF/lqOAQ3Bv1FoV4KJKYI/a4tkkwPb
4sWmgoTYy1m95NTSAZpi8mUjWRkWgGzzZw+0a2G8yL3FFGbWzrBHNao+YN3/noTWS5KC6cMGjD0S
0rTMawrNyYlNvPvuUvhhUIla4E9qhwOJvfCQni8GSvBewNKgC/EwMnYEoZScki6nRmwGz7IrullI
IztEgJxTjt6tRdfHnAM5U39kZWqSnh6rdT/JZWcsotJdFhB4uLtrLN6V3UPTV+PWir1tKSTReGgo
aQEWhzkNz9K1tCwR8nL39pqjzGr+qqWnAMCZfGeD5SqWQH3EWhDb+MFOHQ5e0Pdg4GYTlW2+Lgmp
InZLfDadle1uMUhA+VKJ6SL+eXVNIm4kCKvcuU0jzy2wqEWvWBUG1O0dWZxojDciUQO9ERpmGov3
j7kz/KSY5YuuoZ34HbQ/YqVVxeXJcAXAlDk1WYwqUkicd5qePsKYjuYqkewHHHjIW4EUDeejzTYF
7i8lcaLKMr/QTGOefkw8x8GGoUzStwdRlA48GGFFuDYwatz0yZsh9ic6wRA567tt5vIgobvZ8Pax
XRJhdX6uk1aHwl5Ep5f0QPMIwAuj+PRmSewGKkAyB+PwCAsz/RsOR3aQ2OlGI3Ag2FxYwNJawM9x
+cbsBJvmBzOlwR1nQ5eCibiFBic0P8o7qPlms8JLr0wjYTrN66owzNr2FMkwsi6b27c7KnaLFpHx
l9q9/ZmxOzts1Yp6VJl5x3Qfrt5O95pN2giKuDuWQgDqAUhs2hDe/Qq/bSzWDNW72tp5/SMKZpTb
iRY1Nt6XH0IaFdMOpf+DW2y9c1MnS3fqhu4sqksbwPLqe2cybJJGyywlRW0fnVdHszaW9uL7X9pg
NNFRrdVOhjFAnOHzxduBpgMxYg3jiixanxHtD2rUcsjuxB4qDxGj8jDXkL3B/fW0c/jjoOxxeRGr
ShvK8s2xe623E5cyci+wGL7LsZIOWG73yC0YaHIY3zwdo8AcFucYvUB+sKepxrCPxuoFj8FmyK3q
tsWz/KY4qGyQguDRDPeaEXuZSS7EqcNj8ptrInr/a5bsQjWY04r8oAu7B6dtPx4PuzZLnrgz85zI
YV51n1Wb2zIdI3GqYtBx4iqBHjoiWTEyHiEoXRuoCNqblHvYdnWTYuuris8F0cOSVLHw30NDX8AG
Lr0x9PwPoqFMtKOLp6v6nZ2WiJLdX0i5sTQQzhGiNWoNmHRjPq+Wr/0XfCwSHhH0SppssZpB6SGU
6zUO5QtPNoMJWrrpMIZj6CZmVf0aHTHVvsyb0wprvUOx1YOYHJy4zOAH3ghvpmtfh3BHqKVdkvJh
JYsF7ray3L4WHhnnQWQ3PKelIOj5vgqXREHoRy+rEwt+3ikRb0124cMEZ93wREEUqu2ofgzdnLN2
RFnY8k7nDvNCANhcnj50GvOhT0La1c/iG7okxU3jxzt62kNKqOQ58zzyKx8XCi80J68tJULE5Y+A
7rW4CHNTYgxjIAqKsndiwfmMeVcKZofXOkRs8rXsaCa7fBJ0vNyd+BiGRMqveKgYnH/nv4DRqqDB
UEcGTh4UZiPJWKlhxj3msoXLk4h63MyPf0e9gzK0oKRHo1Xbx9jRTkF/17HXHYYQuvGwUCKY5Uho
JDwKzWEVfffetN3C8w0lAiEmeN/PKkUFvqbRQ5PB7Mfb2kfIjNuQ3fpnxbWkFmafDS8w2EjfMWov
7D2qZ96fnM8OCVJxdeVh1jHItP7eWXAfpT6B7rYK9HykaARTEq00BVQGMu6NgadAG5mzgUDTCl06
JMaIiN9Z4jx6k1Ag7Ebu2lXCvdPlko2ohZSdB7XLtCQ2Mn2Unz+rxy5HqO7JFpLYCzW4q8Bna9kN
RnguJjyZ5dvTrXVxBF9YnjZ0Dotc8s52khxxPAidXqvdHQwMtegGIN2w6uVsdVVXn10PuWjnjuH9
GzfcvAzjxp139bwH2Pxy+z2hDoPWXtZnhHR7e/GP1gVa3LSXE7X+51akXJjply1uGdNi+EKihGf8
wfjUZjX+L/w3xrWcmY97FJn4Mz2LXrIs1/kWJMVyZIjMV1XDWBtBmLAW9jtwdoeTw0g+nQwssOzb
ZtHkBvn4pK3ulc8GPC4T8WKh6zW56ECoFDsP/EoZtLZ1w4PHRCCY7jJMbU5craj7BAwq1IImYH8r
OLbgSD2xJHX33L9vNaRAvqkBG27Kw0+Q+GheqzjTPRuDXBNm9V4En1W6jcnG8LTbNQRK3O2ez6+l
0KmQR2ZhRyBJ+v87MtSdTN48sLR3Md+LrXWgiIeIUYFUyeHizBTI5hrNzj6j/EsFMKowDFX/pyJG
BtDcru6EMsPKQ9uSI/qeofLdKpSvaKc/Fld2ZbWwFv/oiFb7/1hSf0juOJn7wh+yBvCKs/JVHb2N
odmGGvRLvQ20qNXXJwnN8ks0BGVvuNsiWs2TdW/5o4CcCv9IAYWalrX1ueRHOCsQBXgW9So6VcZp
KQ+6h7PFFkeUpEhCWV/n0QLHwCv2XwP4hO91wvHbCcNEY9ka4Q0HknzPFSiOGe+74H7bP/qkxopc
50jyhq+4tbbcEMP/n13VizyeFnf2dqFZY3rBQOuk/Bm16mMRCeX+MoHeFT+AXY/bpn5kr8MBXA0j
bb3NqhqTfs9+FfU04GpDdxnHI57eDwYQVnhdn92zZrd96j0A6VUcEIV2NtkYvHc9PLhmD5aR167n
tcCxOgqzMtmVgu7+M37W0RXk6gpl15xRQuqvwmZ5uw/kkm5VW3rpYz4UHNWEYdG1/kz5qqKM2AAl
mglFH/jpSrlQbh5Ls46SfuaBuZa8SQNP+Ldk4XtSP3zDwD0QEI/yqAfohZh6dORWDc7L02SYDNa1
LiJl5rjDBpYMwnUuINhK1af/Kty2WdI4Er7iChK/tK/LGxTjA9daZpdX16IrX3Nx60ZMbvsem8PZ
ryoMJNky5+59UJU4zAZp8q/NHBp7lH3D/O+wTPGNc8rrFy/xfDlu+TGQk8adM4jj9JDPB/rrwWYi
Ja5eCYgnokoRHG85grfRFMiElT61is6S5nIAqAlSNRVqrY5+P/R2pePAkS60I0k0wkm8yba4KDSr
3ae+LwMLoHlUel5HRRgnNFFA6uEozH+WUe9jK3ri47j/mjFhxHkGk0wbv0lo1iV99b4UNWWCM6N4
aFTYe+6QQxUm8ygqBPi2OUWaldCiw71elVu7MINAJOBr9nfhfGE53JN8xRC1oGjW2CGeAg4Mekl8
fndjGdFNfKNxuZ5dN588XFvQ+PqoEptLaKci2T2blwEvRtl1Yn/6ur8LPl4S7uMSdgImBawVNtvn
OoJx41f2EDSVVp3daVdiertmgCYDndIsag18yQsf5sQua6rElCD0J8wwLDTk/6rEGsobLDwP27b7
AxsqyeNgv8il0JxA0hD/4n6Otm+C3kP5I/7fSRCCvUf8q2gJLZJVOw0FmM3RfZCCVGljaO/9cSAh
yQ6KQvkytoqHOQH+9HRn4XD/Yl7uubHDh9k1FKcm840LcMhsZ32bUL2s7Ey4rZpXT1ASGw2PYK05
TXEuslqEqATvSbNR4ElsPlCPI7ACM14MBhGYxOAECRveEJB67UOPgoU2udZNa0DzzhlUwyqEf1X+
MWU4Whf2dir8iYCWzC29gHRc7SARdID8FrJQW1dkMqeM4zbcx+xE52IOiU7AdpJFz7wukCfx+ZRY
XrjeL6x0fP8lHCSkNTFdxYTKHb3cZFUTH46dUxovq68EHoPk9B8f0kI6TAs5kHG9wxfFaVYd1qSG
TJT20s/GtARcPdsk/UV4dOk/KuJXmjcPwJnyDE6KcgVqFbcgVJmx7+kQnYMX/HC/EpKZzJ5d3wwE
DstVXks3DADH//WF2McUkSL/U3dOYc9lHVymzypGgwmLmo+Fym7Fe/j9wAKpAgzSCxlW6YV0qrhv
8s11Y9IDo///yevHLmQAuBW7+gcbbkyvFSiKgabLr6SBhbOFpOouaWhxBTMOY3BEeBPIk60XFoij
8vYSSm8zICAB+di0Us0oQGp5q36Yqe/0WxlxS09Qi1IsGwSBzMEYEG+gAQugFzsiTNQtuZYzALtd
SmdCwT3OAVCUjjmDeaIDdsu5sdw4AKW3B6Heo98C6ry6m8jXxL4IevlA5NdHuVNzNHurtMSQ373l
2OcsI37WBYUiGUrhBLJ32MwsGXUgLhAGNdlsbNepk6MoKlasdSwPpD9qkrqIg9PjdbZO/ZA6+sqq
ZPdJAlv0EqQVSL2Rj0O2B42TnSJEXtLT4pFwhK7dbwHNTmiHQpBpaUFot7Gt07eiEKxXZ532i6XX
zNULDJyXZZOT38Udbt3WoZLNn8z2MBmxi728ii2C/HPqIYfebrdUyFDqZ8QqPLF4EzTeQpBf2eKF
f/hx/iZsByHOMkjop6LdV2Zrj36nYibiwWMHFddtCWokGHJlkh+/Itu7cFSA8ElTjs4huEK4U7TL
MRYG+x03yrO70Cvj+CI/BjruB6gTCW+WK0Jh50+tAEgyc+dJ+ibb3hh7NGAtdHZVs36HEVrOZ9Gw
Geq9/0IY6EYmDjlMh/k8v97Kom4jwywVkOKXmmiLI3ZOjKVMND53xtbYsBgOmt7XGF9kPzTuMZeX
A1t7MTlj4QrPkVt/DZWI0ecdIhRvcorFzLLWxRL+8ouhJk5+VOvjghZ+Lqz++HEyypDSd0oV+O1P
BlsNZkXqlomNV9S+2KhbPubnH26sIfmrmCk8TLIqtLh0z2Yo6RaEnFV1iT+qZWtkTAlkYLvuW4S3
P3SVwL7GQBF50IUpUKX2DvgxJYFI8ZckdNIzhR/mbXpKXLDyJnkJfroJBp23RvJTs/XuwI/T6rXP
PHro61DcSNG01AFkJC0CYteKSgYTlDgWPo7Ujd+fKabpcOebrWX80+EFTl29VcIeRaZ0GFmjivb4
jJygIYfkp6AE3NgARqkeGVf5ZANzeGFkUvh7qHKh6oPB0EZuiORYEen92xzmDUZvOiirZ4X0SL9u
0MoDF0+nfJbLd9q+luNeC7qEJqfRWE66caosB6dlwML3zX2S0+Pq2suPmBHsa//qtsT3yo7e3ge3
mEGDh5xz5kDZo1PHjYkXftfKdNW/yNsJ9e/YzseKPAeJwJvHfeA80xHumJE/hFIT/fhkVN6fH5pL
xRuWdJgDjWZ54uWc0k99TGEzF7fBrCYNguu+mgfpO/Zl4luaiNhRCt1XIflMznpMX1WVMNFt7NaJ
1CNizj6x/rz3Ml1OLFIeHTDjvbtRw59nnChPtezUvi+pzcF3vGPOW8eGIWfrAa/+EwbQJp69BfdH
ZFf7mm7Pzfo2+/gxRQMT0ur0nhLSiw9kpA3vJYNvNfDR61bSpk8F5QmqINnBbrX6JFv3Z/ESoxPH
qRTFikMI62cOg2yh8VbWh6gSadyHdDlvgqACpH4CjAICsExGOfy5D19nkyBAtX6yisu5CeVCiqbi
RSZ2kYjWbCB3FmyKGaw1ffO7r+uXJ/A9K84LWmgQOwTkCETU4aTdEKDM+YyfY6Q0s6tsQ4+vAqOE
v3UkNLOBpsJ8VO6xJE+cTZEz4FKPRZ0W8nNUUgUDuTH0HPjRM06zwzPvMag6wqDbD4Kk2AIPN//f
A15FkBjssesxnaR4rrhYaq505M1scDUNEH+VT85MVIM5Fr2KeASz2KbGCCBUXn33PcGHZ+COxmRs
onTk9UVO1YBC1fBJAGDXOzq+FWlIuPYCPubo3rYFwRXDyeoBFKJQoKrxtL3IpR+8Ub9oHaWB8SRr
02QWRRilmTgstEvBXpSvg7QpsE+1kP3jKWJjhjAdKNV1XWju9tuclfBecX3VVLEvXDNf4PuZtTjR
Wt4m61RDJJukgtGYrvYDJXmPSV5WHC5bsyWoESVFwdhH3JnC9IiQtJ/gJQcT3gAxCM+Q3hs/RDLn
iCrHkgDNeFkGd4hRD4X2C0lZRsNfQdHG6yFxjmQIz/h/i7SRgv+f0f/mjH/wZd2Fqrw5C6ye+djv
sS+hCe1iIAYlo75Ps4FIbIDR/xV8TwJ+VlOoChEhICaZ0YN04BH0c2k96k1vDfAWg/rFgti9j1yv
YZWqx63iEe4mjBURb8sUlEAhu4j30BI8oGVqA6FAV2qxsaBRpbJ18ogki/v/B94ig67EfDvvXZZr
CtCMQvu+l1BMPJliFvh/yL6pOYAbiy3X8nQXFmG9bnpV38lgBv02Za9IXz1un71CHvFd/+We/VeU
GuJFhFRd/D4mdfeMMZDKOu1G/39MAPMT9ltd9R6ziwqO3xbgAYLRv2VWv9E6KI76iJpOJnfjaypt
9AT+Q46aYw4rhQQuKyLT4srxhWcdaFTKpD14qJqRPYBhFgqj/TSMe/5E2lcbaoFWnq17spdT2sC+
DK8As5hEx5W+VSN7ZaVfA51rmBCGrmZ9tVNJWu34EdVQzSu/WZMTFv9ShY8DbSJBHTbBzMLqjGGI
3kt9kVWYeP+2T6zewG0u4krXRJnEDtwvJglFmjae9/03tlWi18afwajwJdsq3eOgD4Xb1xQvQpvL
47oCpbu9xi6LQIQIk1Pr9fHzgDdUMiakw10EMA++DNfx/bDpOWJ/xy84uKBatYgRV2jnFWqeEeyc
iWb7rT30gx382AGKtvU5ZHcZujd32rJ5HJgc1kq/oZ7yFAlRr8J9Z3D3jHNWoR9SBBxLSQFwmFUC
l8V84bwkZNCpRSorp3MGtQiRlXY/becF+izi4iuxKCYDxU9XIMtqu23CGSwTD35Bxc47lnvOAKAS
bvMPCR5ofqW2MOR4YsqiIIGkgX2m+YOS2wtHBvyqHpElgVxTHH2RuNszCq3FyLZCMWZZDT+HrFGU
ebzq6ZpDzAPteJOKshIvXW6n3IqPScKNUOSUBE6kNwx+aqLFMD2alkHInAghry7PyfIBq36sbu3g
btz4VQYoBbs4PklnNEMDxKsdIybT8aYda2PZ+Ol9CGKcdl4AV23UEapfQ+i34Px5oFXSrVkNlYsD
dPYud2Zx72/+J3bkVqswRDK30IJKlvrcY8WD6Hk+++Ibc1PCKBeCjjQiRKRNb2WURrf7J4xhcPJQ
8lCj1Rxe+rQR1gbz1NX0FUvFlKSmWGBvRLjE2gY44DY4KNF2nyB+Ez9Gbr+eKMcQhj33neFC/JQ/
zAeirtNn7sBGtgI83igAG8o0akpwWdNU8/ZhPmF2U0ODOFbIYVf4+AIYRPdfau9H6KyybqP/O4RM
VtRA/nIUbO6wL6kHevgw0HeK+Nj4vcoawofoHTBIzB0jHPDQ5vuRCCmD7kgZNP50QfE2UqCwgctF
LpcOThi+fx/s11wLrpaAzxWxx64U7gSVjLypT6yhrB3jZliid37rKkFgMiq9KWUiTsb/XDOFtSTc
xE5WWHdt9vr1jl4DyR2quQWQ2/k5i7RbwEjfD1jzLSTb/YvcUKdKGZT2ZqGkQJg2lW5gOMbpmYgA
3s8J5Fm4bTU5Fy2kGXUmWFdqzkVXWx5bu+HTrOsgUiiSVw2HIbnjOCNXY+NfK3Txv6YUFu2f2D0q
mhYkoauD+gZgMDlpI03yl99sbkRXJRRp2uVyHGhkEosWPd4jVKjqV3zcvz/r4uft1P6MI7iVIJnP
7nb6NZLLquQHUmDBJC92+2fCvED3PiBbn2bjyloosba9aOQOAMtH2xdy1F2fvtpTjS5s2HzCRFQQ
bPYvbqKC2P1dvHd6jrT1Dhi7YEsfUVie1T62xjhkeeJnGCUiCObEqXVukAiG/IYzr/S8I56Op6Ad
K/RTWrMRL3dwEBr3UrpOzpH8pmW6Ps1t8Kb83l9li0U/PKIJoWFN60jt5CvamPioEPdevpMywelO
cn7oHv3VBTUt3yxjkCg1T/yFzMHucYgrNF6flwIHssqvOq1NFE515U003a2QsAR91qp+rgd32mZx
oheUCX5Ken8FChHgrECQorIiJX43wyk/WD2fiWIJSFHUYOLS+PER9O7s1yE/Mo9ibtbMg1FQwc2t
f6fUt3YT0eJC2dvR5U3ZY5su30Aaq2sMX1alX2/2OKldcycP80J6u6CRh46i2oyI+yIDtciszUFT
0WSYTDxu8DSwGHvxr1ZZGiKXqGNJcjbn/rCOqWoBmNKhTK4c2cM8KwrNd898o4qcOSb+svwVKtqw
b3HhplMJ+NBPlT/Nv9UNQBbCiolx39p8bHq5zZ4tZg/JXtg5MGZf3mointXqN/5ZWOJwxiBNnUtC
V6P+zgR5oQBnN2JkwsvrBC1KrxTSewGjPmoWgDhQ2YMPDmQtgndlLL2jeIKNRx2nYdbQNVXXY9sw
sL8cS2v+G0UncWEcSLfoIPLdb1oFAvhyWUyB3vFitnN4b1y7iKtMUly+ba4mrVbjMu/8ovOpiD0s
hJnz60huXUBqa9jaWgrKSQtmxbDUoLvftSGWcfDwD+m3xKBX7sRV7FkHCqknpmISj0cCff+UZ9BN
qB1V22Jtu55GnBh7v6umq6+HQsKtPlm3FLhMxR2GsNEgeSqfx8VsSO9ugn9/dTgP/UxlMrdj0qwZ
6Rowl8h6fTR/PTabjPdnqB+vTNtvJ9rJJWAyJ91qiA/ZfgrSC6thE3FPsh2zWwMuNGMdLWuqGIN6
Ho27YOWT/Am637tgUdmMx6WL4tFQ9lWy4BQCTfZFrHS2PpE7Z3UOra3eQGVW2YqCnhOQrtdvH7c5
LVa3kjgLtoQuHUuSbqq/PcJa/alA6iXZnO6YhmBboOhmBDqc1srBmAs3nbEg+0H/jn92qMDwVgW/
WdhBySKxBYOu07kW8sC4RAPTEClSCx7oWFv6zY+DdNROluxgH8OkG8Opic9psd484ZERKkLeGorb
sIa+4RiRZNEBcFsT2aYbOIcjS186iLQbpzj/9GOWCqnmlXaECIupTw1o+PKznO+3H+dMVzOeIc+/
pH/P5jt2Lx5GSJtLcTbpK68p0G2ITyNmVhI8e9yScb6PMWTGN0MIK/B7rI3ljiMu7wNRTRXs+1xd
F7SqOFO81MOVgueuqlQEaFmlyc9FRq+lxIyk3d6iS79JpeM6VJYAgse8Nt85RCVfmYuKHetCWEfL
fnyuSZx5m3ZvIykFI/JhYGlrVolc7lUjeB4Wje5acf9ahV77L5Demq7iIWkX4C6C93IxwFprQerj
0Dt6+FvuUetM965IIx+Ml4mLNzQy1aM+nRiE9tcByO8snesQrqADuN/mxa4DVWtrgLlR2H6HhblU
X+LZ0VENjBQ+HMS6UURo+S4VYMu5kuqAsnmFhjYzFheAPC13g7beEICTZnukCvRRMOAVyojlWtvm
rafafxiyUrPIOx829UXNcEh7I/kCQgaTd8305SjLuik8rjcz3GSNbjQonx8H1ssEaAarSZa2wWM0
gl2l4tVuoDL5aRfeOnenTtzYvluOo7x37eiXpzOsP69oZYe2haAtTAyCfg2yyWIaQXVgz87dXjRf
RT9sWZuU5N8jI5ygWRBqxIe6vUQMc6YVciOWTVo9wB57feUJaqHmunmPSetnHdvQ8MpWLr9oQ2BW
amrqZciUkS1rNMSXc+2LHhj+LeA3cfmvtP78AaBK8fJ6cMItrQeHg9g5IG9cEuP5wWqkaFWhJXCl
e1yseSwFe0LY6pGwW2YXVG/35rpdUfCMYYz0SijpXwfZkTDtrOQcuxFlLo1uTyrNp7yRV4HsWL1G
n/R2BIJRFjE+fS/imDnsEhol1lagFIiaN+jCvbNuC/oj9P4+CXxaHnUTI0tyuCRn/6G5nLJVtSHR
9I0luPdBZou7minKaeeSOoUTLwGyolhWpSiMSXxLMPoS5gu0knNDcm2eXcQtn/bOJLeCe57pt5hh
C/tzagqwWjIgMbqrBJsUjY43ZVztYas33T2vcoeakrJ26pLxEwKFzSIKX6LrpFpl2TSrtKIrJaMV
Hxzdw62szPobXBOJWQHK+QSP2q0fTX3i6JZuS3l2bORERvi0m0/CzLTHJkyzjHxeTU4L4zZsR0vr
QEoTOPZ/WSvmJC4LWmJY6ZVuPL+Qy2lxzvFfvIIKLZlzal7blLKAQES0yGH/1sASI1/NoVdqrhgd
ZFZdIdqv6gnvOqsZuP/01L3nyXWnc4iRT789UA7qd9qw70FzjspvXGJK77SNG3NouHLc9Y7Z14S1
JWs0u4r97VG8RF5aT80VpIIv4S6+/xt+gyyjStVFuQrnEBGcbDbaE5ubEkyS1xw+u5Y05oMkFP1P
gAzJJCnGb366AKz1wv5mFQjGLin1PoJpZi/qEB+W0ETOtgwroVlOGgNcOjWtgPeS6SD48L/iKlVZ
YPQFLvL3Fma5AQ/MWpwFG3hQFJ8yWZDwi+qr/RGDJx7zS34zfbgVGFgOG2P87X8JxQV4rxb5970z
c+0Od1/s5dETm4/ZXF2x9nCtNdL33TFk04tD2Qmx2uZPKaEMIS6m8L+3nNS0g64G0d4f73hBIe26
Ke6myU5wX4A42VVLG3ywPsYuRpGLErxUP73JHIXqKeMpeR8NMUZW5c1XX/P1NwQejjxgQHlJIRo3
3wPaxyLwHIR2GZvFvqiDeha9iR+8zTMm7mFKj7/VKkYzZmUUJN6x3OaKbfS6woVF9rEfUhvU3LlI
zVWMKGfTIgPhqUZ8aNCPlGCW8gWnKRwFteBakL7fz7qNxyuNBXg8gan77USgvjcElne7rbsspmDl
aeDQ9F1N6dd2i6RTVx0GoJTmoegeCvncCTA4wckkDioy2kp6o+w9BFFpIESl/Ri18kWFrpmKpds5
xUn6ITROBOUqNWw+xXBoLM7qN2VIEv4iaRhraYlR+pcs91lMFGr1svx810jGfmw13W80nGT3i/ac
RobWFOMVk/O8oa8H4AoKvVJAtLa5wSFt8wO6Qfq7JdXZ8HCiS5FETs5Sck2g9kpJoU8TqBCZJHFS
Lu6iN2GvpxtDBSSYl9O6h2hZtTPx5AENnt5jovQEpy4FOXdflBCc8BHimVUd/4keqdOvjLvcFIrc
I1GBkt8Lwht1zV3hEP5Q8m+qi89hKM1mTGMVW4WcBJYA/1eeovnnZbkEKjq6xfr9cuRF9e481gWE
FK/n+5AoB8cd7hSQHUOKSm2DVT7/mfksPhl+RgqaMpK0AADiSNoXB/XHmoqU+E16wZjTTcNdSn0b
zaljUV9/jaxUkfDlUNHh2k6DV6TyAymt2nPkocyMvbSip32Eizh6suwsEAcBIrYFQDjD6NDsh54B
SKrYhjNOJlThEsdHQJvtulVxXAhNT825O/TbJu/f+1tobPfuwauMMQyD9lbup7Gezes57FMmrSd+
aqvW/ylnNYw2yYy4+Ol2NZ4TCIRnwqX/NmIfOWBGgvgEeT43S4OwCbK9zpIZc//Jvg8feuPMTCNB
AJiRF3LysiKy+SHjYkW5lt7GfAfRnKdQqAkkyXDIID1GdGSAHqe54Y2ZeXe41UKXwcdKoc4O80iv
JwyOAl5MnrkJTrdMJqqLPaK4+vo1Fgx+gZImByQq1/dw0gPltD+m4Sd3SB80iYs5G/ScfoM7p4As
mg2wYted1Y00/dpOiAhVZGeqynRe7njH4zDV8jL6hz344uHI1cvvoXMW3ZJQVGLKf1XYvBtQaQ6h
i3aZF/IkFzz9NGkIEMvYnmGPZrHIo8DZf+qN9Or3Gv8GFYVANLPDFSGLEeOOMyLd84gChQ24h4Em
OPmagjNVY9gjNamPq+E29ZhUnuZZ9IG7eSAKuQ6m8/Ij1xIf0KJdRujLmjsVXlwlqmaNK2IrAUdq
v4xGzPLu4byceQIocb3V4t0v3Ip/Y/q15DWkMYunDHUQnVXAl/mwkpTgJyGVuD4E4TbGZ9SJHWBJ
jC3EZNIsy5XbYhp9m52onJ866qWD/EjI9QqWnmt8meUwaDWOTHizR7yHI+kV82crI6nl5p6wI17F
SGHVYb/12RwH5JX3IRXDmjCSDmspZZ/VjldAkz1HZ7NnkkVBEF0rU+UaNCJCRhzA8ZxncRvC1owy
Y4D+fFoTz434pnmHmp3FmTt2T4RTUI43ocDz5s3P/4/n/JA+eC0sDgu3S0VCUbu9XmiyC1L6eVwh
kAz37aL+utI0IL6NgBvszz/18Zpi8dwRsBxUY5XDqVF2gUW5Y+eg+b6KZKLug4yuMXopB83FEYu0
qrS4OljsD/aUCov0SBoYbEXvE3zwEA+V+cyx5gHfTzwTc9ak3N31PExDC7+bFm3D2+QzzS1ZJ5at
cpUiaPCmqOsbHkGv9F0EfEy19XYUNvSxSKnrCJHrgtTQ0KQ5UaFLWYwuXoiOr4FXqcLtbZMPc6Je
0OkJW08hxSfWHZ1hLmAnJdKSr/OcS/n1rsaTnhsmo2H3J3c3SYQST5x0tMwRp7xEvB24PI5kvE/A
q3f299CMt6LSEorMhKmD3uvsXYhZVQ6gtRKnPpRp8ZHnCn14o+67JaV4SwePVhgTmLt/Ri6Fr54y
I5P4tAGcpVeMm7qTIwjmFUtZ3+j9e2025pWzgdaYvwE0MyV3PxY1Mx1kTz2BdnmMn5N9T0uMNLmy
69fjdjrbl6SQfWg5WIZS8GdKNj6RJJ+Y42Ewe/szIRutaguZAvlGjLXF645pBAdnlORlq0QQjenX
D/eU75BO6ZtgSglZ6WGFr7Cqnv7MrZWcHumvXhyEkVi2Ii1664HltRPjdXG7iKTFS+7mfbRjzyJX
07ibUPIPsAmZfrtxVer29BIXEuDjzjjRbX5zkd537nB3fusqtldps0DZdOBPPP7RqdppiWGbo2h1
n9PUa3MBfq7lvlLwxds3m7JqglyfymO7C2gJdqOsJE8yLpwIF5fxveW88HY9xGASMiFxkAkI+3cU
6nDFcQoo9GSRhrseVLqciBExizd6WaALBO0caiW9k24ieaKczOTjyeY8rzswjKL+l3uI9amA9yqj
YGCFEdMBcjn6NCcBi1mndJFnOjjjoICYnRq+oiUAF1dHzRK1FS+ikJp5YUy0/4EBIiY6lCc8pKLP
owxl9mmwZ/zPzedj0/AqHgd1G2CP0NN6XsVafpua/Tg6b/1kZe83LToB04y/3ponWjIfRrnQqFTC
gKn0nB6SK8KotdF1oNpUx2Cpkq6FcG+Q7C+hjdhzgj5+rUEU1SMPe40yBzLSFvmqqyHcNz1xcnjI
xjCi2ZdTYvXYkRICzG4N6iSoy08E/uaChDKxaZUCpaa3F8gYR9fyXxqoBNP98X7CuzmhaxSy/t2X
oYKSe/N7esoeZfBnD+DH6CNc9057/iB0bqPa3upU0zdkcBnuU/w2o8HwBu6fQN6n5Tg+Hw26sXDI
jDZukHhI2ftRVoUcYD9G3o6R/6aDoRBpRmrRFqq131e5Bj95uutVLtcV9PA0QBNLR8lYo5thqZNf
jBX+ByJzU+dPaXvBrWD8If3YkcEHojEoqL7hhAdlxtOQ80u7PJ72mJ9+UyeN3NPTeUzUvuFBd1Rf
hX5CYhD3uJWjmtsS8QGhS3aQtm8JpAi5uC8/948SLnhbDBoXf3HD2jE1AMV57XDfNozH74ciU2QZ
xMs8Vv7dPvvYPQGGiD0d984JILfu4xsf6Vp06XHElM2RkvgHsLP8us4nPo2i9/9IhCq6n3QKPzam
nQ09l4HNmS2jnb59ujFqRQkCDd0MIz1AzG86j4D0OJELLGXd68gEatQAMv/f/SEzsE66qLvkxnBy
98kFmxN/PYQlHKazxS9dQRgmNyI21H2rVVjIW60GhGIR9yK/yA7iIlh3Zbby/G/k4gykv89RG/iB
O5n9NaI0vvSOlwGpbIT16rn0UhPhL9SEunG2IYSr9RvLb8jYzWkxFZRA/9Lk0pC8ons1r6/p/KZw
jX47M7codRCgEiVesOvflihpRXBKIpu8apgxNB15XuxQKCxQvXXPW/ob1Xgh8rBBtbBs8RuvQmYG
siePanqFbMXkaKYUClhflobMk6XZ1yR8Ze3+gkMQhPQsfkXIMRLiXdFTDQAuXPXWNdvUv8j/0nqP
6xB+hh8L1dnROT8V22W02VFy7D6fVZgbuNlhnkazmM3I4KBoDPLnC8lLy8e0otM43jHc/JA+3iQg
doFPQuKaCN3NJslfCpPa52qs1N9YvSdlNbY/wbylfS9brWuLuqPHkTuJoN0XcUiXQzfk033gaUz4
ZHzdfhn/eV5mwndrc16StHUW7SBn1a4oHJoGx2e4KiKrmQisFlOFw1nJw6IDPqsH+HAQIdY+MCWF
38x6aytcZNMeAoPLEccukivKWRfbDlzC1WmZRwx62lTJETVD+dk4BEKAyvzsmosywGUnSh0tp+2k
9rTS86pv0d3vrgB7U/kiqZYDjYOrqjvsJfPiElZDbJpQMTVD0NF9EtI5Cjg7v2Rgv4xECn5LZBHt
7gfF3hk6yIWUizRv3zotPmjq1ugfNA+HGMzCe3WGN43j9rLNfgtKn0VuLo7eTF31w+COtTBxl76z
me2CHbKSn+I7lr1Hdm4bB1blbfIPBKle4jAdbDkl7Soxd8lyyP3YHxERxw/QuKkV5DC22zM6uJeM
jiQ/OsEHZHjajXUghaPbvpFlSHOOotYGkHJ6sVV5mh4XLJWET1ldQFpE+Ss+MDAI0gx9TDaujjlc
WHWLk0eOv0TtgiDO94fbn7NpadsgXY+fb0oh0z4+CoBWaU9IHiSh5TomsesssqqDXMjXiZ5haSfw
u+Usg+etF+h6Ofj1qSGgWCRBo2YL3sHfBuxn4sVygqwJwyGLYjXDL3qXedW+5zNTPs2R47gG3RAa
xdzV850RCMv+k3KiHf0Sw/ZeiGJpRE5+hTGdayUXY+Vdi4WgFsc7ScN4pGGZE4ZZ+dhwy/fcv6jl
+UcaH7y8p7RyA8NnIX01ZeBsLNlAvCnRUO+kPBBVuT9i8uGbGN21ZNmDWb/5lFxiAhYHwKhNwt1M
/X5ZMK7aozP9NHMAUrxf8xx83CSIkPP2CPvnk+LU+Ix3vp9x2dp2OHPf8lq/YnXLnNsCf5bKyHGx
SVcaTYWj+bNBxDs7mYi25b3zNUvz6yRaZ8F890p1Jwlw6kwXsYlY5haQJSf8Y6X+sgxWi8KwEZlZ
3l2D0+GS+sOweLVgltr6LqGCy+mqNXQkm0EB1iPUHrQt0/1SDoGJvAai6vEMNkoPiEMYDeDhPcLW
RigiZXCgvEZDURemld1CO18GBwO8ocSeQ2dxoz007ly5ZkcMe1qLq1M3TmVUvMZNpdedgLncmSJW
7pVZ8s1RXWHiZ/oDp1WiUJJL4PL67GWfuTdzgSY3Dl2DmOT8wVaesMvQHAMEJxeDmHJZs5MtJhzG
G+4tRHMYJ0t2C5L80a1xyef0Rm2sSbZs0AEp8AYtr4o954uX6jvAB5G27hqjgo7GxSiIPN5A53W8
H9SSlHzxJzz55MOWzNcAOr6FdOAbWOni9T1xfaL7dS24MtEPN/CyLx6UGTUZPohpf8/R90kpO57H
QRp1tcK5rMG7xZ5xqANWhoyASXBOZ3y36jpalFzyzL2P0EBhqeCtdCrwyDJW9lJRj7KXtAP1Zx23
seoLjTVZBL760/XrnEP9ANmT9YHvfvs39T5H6a5SQG+9q4OuFMUYIm8lxsZx22X2H0qeeKVoJ838
o2WpNw4m3oIbMQjfY7TtYafD0HFRJcgrwBFHecX3TUlXiXPphsunAta/ELJGPvDVJCRCT8Oq/u3x
WtOM9PyeVf3ZABkC/E/n5cjZD0Kk2LPKQ6se7s0XNAH4nL6tMpdME4uTSV49lVcE077evLLPRTFW
sR/zfBb/I1fAvT64VEO8sE8OXhWTfBVIr1nJPQNzaFOamhLXmMVUTeuvb1gHYCbGRv2pR1fcPD6y
RrL5e4t67zaR7tyVjCLJYNhUt83BKTp0FGX/+dLXM09RcnTLMn/na3pcqdWlhzS+DcCqD+eqEhwW
F6KxxJ33+ZadaYcteHeKsERsg99kg2IlcU6ql+waJdQw4mNo62uvMfMMtu2ZBBZP6VPf41tlafB0
27F/imdNN3Bgl3tt3kG5DqL1vMt9t0qzuai7PZaVz2cikhVCwTJzlLnUGVIFaSZmbOQfwbx49EA5
a5FspoCjoTKrOra/QZSsOeFCriO5KW3Ed1bLO3FWMzzGW5XR1sxuT4fUwg8f8DmKmj3bCeN6cmFS
5hcXjYyBhSozF+RpaIFPPbUB7gvGUtQr8tN5sTWaKsiN1Gd7UrTs0X18QHeME0/rkDYTIAe26IKI
0SRpTYt/8LJf765RLkpDecJA1TK7bhWcDatN6VjcypvHnkT60qccb0a78mAQLr7KI5amRg0bFzX8
ua8zsAWAJzoYiMdVUloGvxktj7zflvXvg3rXds+Iye6+Wr62B90kEbhNHMuYoc8e2QIF0TJ8R7n5
BnDaxsG+86LnPCA7RgWtMPsjvI8mMGQVEfGZH/XKguWKvbvqosJH6ENAS/CNxWVBfYtsblIjLOCd
VJiB9VuadrNrB/ZR5Lf9UUlf3XAYczIQhnWMOLpt5S+7ex1LH7AHGuYVyJdk3lN/GL5/sAvS0nxT
f50QgGSEONGOT0S8w7cL24arg+fTDDZDadnzuvJJCsfOuurp9zUfcvAqiJ3VsRTIfhmd7QJHgRm3
j6hpPiO0R3mcm5fMZOMfRwDfHjT8No5souvlj5z7FMkxj6TU+2GRHY6iOkVPu6gkavzuBiiKi3Ly
USD1Y4vLTOc7kbbqNwe0XPlTWg2EKvDKNA7lNQtlKe7yaQt39eoaEIGW99OocQVVQBNm9EBNZpd2
salEvdSCH45xUlG6OHcTl7OFJJ7ZJsmreEFSNFZ5H89qeUmOd4VaKOb3bWRs5jABBcSJh/2z3dXC
TXM57HtUGw9VPjWHTFXB+ToR/vFZKYNPBgGfmOuiv1utxe/xDbPbSBma3zssFLOhU5ExxRWvhjEI
O8HnEvo5UQlLFft1YYSwDblmodluPAJ4y6ojoqDzna3V7779McJWNpfqUJsmoRVJz10fbb23+CGq
fyIs6wEnKaCmullRk0guogYbw1bjy+GePjxy6I4SXUxpkK1xqPxi4fo1MMnSzK3wFVdUkVGo3KGe
d2JZ1pIsUsv9PEfPu0dV01t3PdpLvTW3pWoO+w+DzGusCMbaGC7N1B07YZLbGNv6Dt08aExV85Hu
8tafdd+rBZ67XtNWbHoyhGoxPGLOm42ae3GyFilFcSaSOHWKPRN3zQT8n/wfC5usBHbnYJ+2gNF1
+f95Ay+kFQJrdPLekkwEoCHQ0/2irTYlyh/Ezlf0NYX1kJNHP0PZNGtJYiJXA6hNrx53EACSyAmq
3qDhFYAEwr47bzElyEIahn7J63uwfJjvPtjHk5dtY2nI6DSt1/Lz4OHXodCOHytS7Qb76WeeEnN7
BysAo4vRb/AroM68g4+VOxDwn3SYQdw55Q6L4xUrnB9uUg+x5rNIpoCoZ/bZxw8jrp+/BjHt5ea/
s90Z2z9atSiNX7OhpyjTisjmlJf3XK36jeSgXjoBQNq/sXHIZ+xPVeKbQRyZnzxWpgXqSB9W0LyK
pHZSZ35jeWB85WEW00LwaLtWsVi79hENI7L5WK1po/H9126B/CXbGseLq2vrinLPt9EvNtLTekV9
JGH3KdT7TZN/DF3Ib3VVt4enf30vMT9qNkQl06PjIGLbytp6aoz0kaVIe+cHTzT438SEbcDPQTEY
QCNJ+qlHayj88W3VGVvt8gKVEl/aL91eHBedtEHVy4BbiGYlzCOj0SORgeS/dt/rdL3nfJVy1kPE
fu8vwSkkS79vmKEslC7CNXU9MGZ82gyGdDeOU7teNffMDTsPWejaK/Skxps62U/A1eOSGVfuEmI/
MpdyVySImbKWsvzOYSXCK3jia7cIMTe4QYKw8cVn4+eqic7/YoffIAG8b6lkgWG8MJAmg461oZ+A
Dr0/sHgyXCrpqbW9kEqlPg+LMzgAuuX4vwAZQdI24axGdeVo0qnpXleUAImmSENaxP4nsP+fGdUo
Dcsh6dFOqT2Szfnsbgfxslelc3dSKFhejOprr5uuIPHezpbBlWMaD8gvRFEuEJSb0IBJSSQtGPSy
YJ5G0nhis2Oq2KpfTBsV2Iq6A/41AfvbHGVjNOUZ2yY8Ya1am1pqr6RaaOWw352qrs9fy6yIJF/w
x/ReD7Ii/bj5wUhyYaH246OrMT2mwN6oaGFb0SDC6aI6V2vzWjt7friSscAVviIwNIGhIdG1q9wZ
vt1gHaCA20aB8krOsdpco8MlpUTlH5ShfdrADz73lNUMWFwbVSU9YUoX1o1yr8gqVUnV6q91hrby
WPFfbdEh9CDktsGLVnCtqvOSU2iAFE05IGxI+AjneoxME0N5/37Dsf+he1XMxxUve1i6Q/LNOHW0
1s+xb5/G9q0YardcFkIW5XymX8ihH1fMrIRkdaiU7HauObIBNfBFchXIrS7khbOPPYQoclmg06h2
7pxG/Md+/+7J0paQX0M0RyRXZdEY3eHTDRP/+XEAYC7WsNT3dEnq7afwZNN6djAUSoFzRqFJ78Yl
norJcDuS3TS1MYxSxS9FecRLshvd9sQisSb9oeRxLh3w75kJ9xfeCfmFZC9vpLfa8B1aPLQMaA8g
94NzAz4tKfgLTP+bAA+2rGOU2zDmqMQ2eYv3ZFeDozg0QM8Z2HntuD5s2mH+eyDucLCsOyYA/kop
2/wfxNgB5iv1V0g7ON/z06tncq+hxJOVTDPnzFa3Vajb4r26su2mYGWzCZcfrDKGqZtNpgSvVcfb
KxJYQS79nMOM3m4FB6B9SyXxS9j+o06WeJ2CzsiY8FuUodhTTZXH5FwbG5BJQG67oPdXCya3TAoJ
MOC8PvdA3L7eM+FktQgDcD1A8lZ+ivDdNyfT8jd04TDDNjzhWczqbx71ZVaJ0AJmy904VNmMoos8
kSdgg991Z7Ze09v4YWwtH09b90dq78aQLXuF8PTXY0xQFaJpz+f7EwjU1OhaNnEkXIoJX8bzXVcd
n9Yf+hecxpIQZHWItli4rMInShVY+P7AmV/Jhf2H8PVuyqagHgUJFqRha/MwKx6M7/TiLcUBs9hW
9FoaIJ5PGC8GeWr8MArqvgOhAXelmQDuHK+IqtJUbBG/8VFyPDWSunjXNwFoJPoNWgYxCJhA/v3i
rjQp7eAEGzt+Z/Lmyj+CuDLCzQp+wrcW6YFiljDV3uWGQKeMjsy4fpFoO0iCNa8Fla+k9T4nxSIN
Uf+1paxCFq5ezZoNMINSKLHkdauW9jclZb3js6T0bfMyb6fEkFjh32th1t7UD/+Tm3cMBqDpy8+7
gGoC/yiV/6UR/58by/PInOrkLDRfPJQodZybZUaa/DW4XVmfO5VapNc49lcZsZwMEi5VWa/YOBim
j6QB8d/pHB0FrINEx2nDObjIE4POBxDm6BtF+en9FXTBYulRVHja8Q077SNUZBvNoWSnsx9lsxGm
cgs0cnTLzImWdlfmLyUszsuMAS8wcm715rssYL94xCXdClWg23awaBcdlQAQ0M55Oag5yCuPHy0V
ioplMs5yamugyUTvb/DjS/DcDPT+/cdD9P793IxLXmTaeFQdOfFspACwl78BpOaNbccLh5U6FupE
hvRgg+IL2crQimbOGRBuTAKLBDDKPA9rKAkFK7ZVs+2wP9RVHY8SZxvn+M/BoEQ3F9Rp7koGJSvi
yz9vzieJCFye9MFakP6yqpmJprdm7wj/jgXVYeDoanKkNpCK/QQYE3NsyFFSC/A9XkeWI2Lo+rkT
QlAVikiPXDQyHH79Sa9p2FneCfOEyUast0zhM5gFLe8A1wIvT+jKMA9hltsl6f/0KtJbcf6Q2MNf
a6iGzq34FoUblcfCbMYUaMMnxaT5E50X8hlysKeok7T1ysLBA/L4A55NuN9UOHHj9Fu3v8Ylt2AU
hhp16n32PhgJAPrErB9PLH6GJazcvrmqRLw6e91ti1l/24xdazxwrcFP+4/+cl/FAWaNv8cDSLcK
gbZLOENoNo2xNhTrN4fH20k+n17yFPFEpTMKRi9vXxTyFQtQ1E93+TllVzxFaKfc17L/fuo6oUVJ
Oq/uddK9mz8PrQVPAD4Z5DAXJIOEu7oiNI2weS+zQXHkIXYa6QeKR31QjHEcEQl/nrQNi4+eBjyi
X3qKFZ9ybzMkEU/LlCfCT19YERVacknMNPgwZyBpSDvxMQlRyBKII1IVVXBlq415WNydOXMMI3Er
IVx83eoSvRCx4b//b2I4cuhXr/VczSclrPN3uTuNWLwkFT3DJbyUnVc+XS+z5M7eglnHfgDVrIC6
K/QYefnxwJXca+xbmFVQEnlVaF6b2vMXpm/5vsMxjEmLqQsnGbhnRxtxg4N1KP4EODteVZHiMAfW
KVFnuOA4bwzD2j90gyR4MjEtqGPIwSjs8eD9OJ/1NNUayVSE/6kBX4cGQvBLuPFlFCFHWKiT1SMX
H+1IK0ixyRYp9cD3kALbZ+UQeZn8D/2YZAAicxH9/4AP94Wp9a48TXH566Jx0HaCMatWwjfj/cXr
r3uRo6DBjBMV8+ms1gE7jvZo08UeAKZEaEV/faZ6t/Vzw+rSpNxkS1JEAAqwXzKabRcLp6r9GQI6
cLB5S9bFZncVRuXE14rhBxGOqP8xdQX2yopMS7Usay3HkOy10mYjoCJahWOGtxBWEfOtbjirFxml
5PAT5fbHfX2YqumudB8gzC3sGg3F0tPktIVrYds+Pvc6tvprkbWdvxmjvs6F+mhRqDUHh8d6ZvMy
v6N1CqGceWZY13+t9gMdILF9OySxYd05MXlgqIsuv/cJGugl2VmMImFZydVg3SpOwAFes9Yqrt/b
XU8hj4lwqhn4SDwuIPJAFFUlP4yVxNILAEhlpx9uExnOyqrSrdg9n04qIA2VSxXt5OBtD9a+lIWi
R2GRvG/p7u1VQd6peAlq3x+4Y53Xrsfga1FTc1tXNJEgqhmMWXz+kA0vD0XgEjqiwfRXE7zOYNHK
CPy1IVHAJDlZfF6Ff7yAJ7NBfAPLWIk1BAYC+yn0QUXfRBlNa8w/SwXr+iJ+uRZKQJ+qFn9Rt+oD
wjBrCUJHCzp0H+CebYeLhL7p/h2Gt6qjN6RS/wRC1tLolNYw9zVbrAvk7WMJJA0G72ZEeCD0qfOc
Pz0aLXUsfSz0pFW9VQF+/TO+ZuVWfXlg+RL4bJrdPh2Nw+Mcpl6mmUSNl9k+BGbJAAbhcKW106/q
MwJhL8gpEGDsn81OaE3J27KP5nYNrwlbcy6x7TcDjZ6QJX4/H1f4vdzW7U0M152LQxM9gUPMq3De
lmPgEIBXekgiqpArbu/fhYejr6yGJH/Kc7MxgSyz/JBStz7hBnDBPCIOo/CPHUewQKrJatXTJMW6
HZ21JJocGvc1JMi9NfIaDAOHaXx/zj/2q8Qhj3RxuhC6eLKWqJArlfx+O7MoT8OpXVb0YjQHazUP
bWjGSkDT2yEjXj0aZAd/UXBLHM4hoYW4Gs+GN5AmaJgGXOdf+m1Fxr70wlT4s04xaZibBm19SoJS
49elBuWcPNOuG9Y90obHLeVIsVme1+jNs7P1lLNjBFJusPKWof95Zm8oFkUolaJtdxQqWg6qNR7M
nZWf8Do9hHxbOFWS7NtzlvAcvoMXFsn3pQb1HBNJuy3KcAhmsNXP/ubqzFLuvJkGo8Es35Mr1RhH
geCEkh4DbIzfHa13ZluHX7UGQwxNbq4VJbk9bT4WyIFaICECAno1Ly1mmjhOvxSLIrLTZYVhwkno
CYTFZixDNy1iJRza2ZoOStsapS/LrqvzdtNjNgG8maqhD6OhueN4/Y8QAfnEwj9lbsSsUN8bUXPX
pjpsMIvGdQ7X6AUoRYirsulceTGHBanCgwj9LTTl/+MP+78uJ42t2tm9CdXVakv3Djxkibf5pj0D
EytJrB0Z61oPQYA1z6COtIy6kMFkuchAyKbixU7VgEaEI/JcLrBJIoHqCWIC8VIqSNnxaJxR/Lyj
QRQ7X6dF+WSJ/8zEk519IlHwVhBLFCIZ61nDWAlgoK3Yan/sNpbXyeVnPfP+TzxGnRGhiElvlJjI
1OyQQdinWXgqkPGCUAFJO7K5IrWRFRgz+f3qzhu1D6i/lz/iFfwcy3tnUP1VNAdNdFi7sFMIG+na
VQOPLO/GvyhxXWONT461JuvmUq+O5y2va1y50+fDVTsoWDhPGeP195yKqtgqCGz/Ch59BcEraHwj
VKBdTRl9lnaVRRRWkNmzWm93Ut8w8iyaMoR7sWQX5TbEnGHzzLgapO3cIy3x3cFgHE26ulUwielJ
cMbYMxv2Kr3vOq3OmvxjDpHLz7KCv9K569CZ7BySD1VIZMgkeYwYlIfRJvR0Cqi0bDSIH8jL8gBz
7pXmS+pjVuf3LyCyk7F4vXq2jsphjI7ZYQf/u+F1e51CDGOuSXBt+MNJU8RTxw/Ao7twP9KkK3+B
EbRX+R3nRvR5545mFat/7SVNJ7t+wZlMUjpJXdHNA2RfBaUmDrR767amEE8CH/ngZ9aitvIoOC98
PAXbBGUapeK77J+6I4ED9sa156eiFVd2Ebv+/CRJ4MgLrq4+mMBLn+/YCqnqoFsKGr6QWqCdhVfx
U3ZPTtUkC1cG392YEQpBKtKL3lXiL8KDPdJbRnYVInqOr0SJDwNVLkawt13GMGrjwGDTfuwg8Qh8
E3vbwujo6eXUFSJnHkE3Gxo9cwEpEvaq3upH+UOnSO/jOzKuGoRrQtd7GcSkMwGgpaByRUKDeHBI
ofKLpmH1G98VCpEb/QRdc1UwKRc57SKSdfo2FalHYNQWTu/zZ35fWZQ3OIL0upleeiCOfXVlvMqf
W4HaeMlCc6Ps9nZlVEtmCZwV/pGJfcWa8Un/WzSZtnjBeWfcl1b/86R5JAmSZ4o8ia72Y/zRj4ux
yufqOrRQDiifKna1rERGir0UqZAj30RzDltDgX1y4ibgxSBYm+pjjobGEubMJSs4UT4nMdYMWMq/
gGMepMtSHw2c8MbZBcvdq1D9y27yJR6VSxzOCWV+b0QleK9TXRdEA4oVdpwsQNhOPKpneFSYt+L6
XbM8TuIeWUhfhZqykZD5Epbu4NoZG9toq8Oomud3/zFmcziBeujvjQ9LkP/dN1qtPpn6Ys4RJzEO
yZVJuBJPmu3YpIm5uYUZPBA8dHKalmvdmOk8i/OlroJS22xNY9IYgKmEBXKMtyZ3n0sSFsrJkHyS
NcJNoOP9HWiE3WkQJe+2Nu9RWPc67VmPrp3bP7gRxpDC/DiwAFtmtd5b3C5qY7oX8DdNsR+wfSzc
Sc7oFJLzkLbr9S5QFEmQ8G/qvxWXXQaXI7ttgePgl03dsnisx4U4xkQ8rAzryHEvuRFPD/hapLAm
g4W7qb7p8Ji6bI6Os3dAHFeBFoKwnuDzuQrccBsdQv1f8R3P5+rCMKhGBFWAbdm66DDaKuKiRxwh
ZowgEErJzwzs/OO+rMkHNjPSctgcjpZ57J3/+yjV1BBdKtxBfeklNS3wSsmkP4SI6EAuOADw14xs
tQG69aib14ZHwKHnYVLUZE0HLsc1kv0HNykDEkAV+rdcsfSNXyBcSHh7gnSiYTUSK3Mh9cfCratv
BxiDxWPaKZDP2ZA82+OtXqp3vBz7yjM8DLDxt5L899NIqoY+ZBsDF1BjXHi3y5g55tiKqSuE9/gL
JIRoDzwo+p7Sqvz9E+RZIOCK0NLLlOQrbIz9ZbGn/3+ZKtl5ApDxIUHeBjvDPxEJulJcxN2mpXMq
8xwmehWephSu8yJbwNFXkbhTppiCjuYmDuY2t/E+c2PQGtOgDGTFaBD4cG6oAen4POWoQMkwSp6p
/lGukMzYH4zGhKHXb5iEHcX30ko0dZ1P6pFfwPA/z5qliG3R/T5jMxfI4oQaKOWK68bhv1Ijamat
pceXVNwMOCDhqjXZ6qmUAbktV3Z5tylI+s6ccubaPxFAhkMhJrY+t1PBigBrcwMOWq38DqThzvEG
uj1NApn8LmLLw5D2yMcgK40yu13F58TRr9rFDfypQp79jwFgZ4/tvnTcfaPxSHFv4XzOmsgkt9rA
wV9hn0EkndDUqCirrUAwKItOYOTu4aE0aGSpLMJQxGuGG+0tmkXzuw1EqqxyTwXidgQzJK5jHcAu
OatpDfpK8qNY21SOUfNKBdUH0CRz5yniNQpMAhGlDN3w8zuzBmmOm+dF6IVhIN4jM58pADu4nt27
vB/8RyFViDLoYV7eoWFRBg98IrHADUceVBk62moXI1KnjGxkanphjshNFiNK6zzDTAScIcuR8Uam
au7JxYojtGFDJgZFdEJu+CVPZQceSXLR8uptIT4e4OmPolFcQLPanQkKRUWOxp4RzmiBbKNFcZcG
TbkhJlh2hCHnEb1meZnKrvXWPjQtDi9lYAjn5HlgccjlPGvjV73yvANrSq0k7eytveYtGCkaTU//
gOK8kmu5MYYy6/KpJmtdxgX0y5Naa2vIJC7/lWFOe1mgfPlU/KlapsoM3VB28CbWS4Lm7TXMBYcz
/W/zmQ/kDg2SZum4OhWd7u82fNiIlbtqG8DpW9HhvR7sTltUQlm25y6k1YPJjPZAiL2oprYLZG8x
dBB0bW7kkwS3rnQCd6w6VT42tzDK6oGmOsjt+at8oZ4qHFdWpWUoiGAbqadOJR1NpbmTJN/m+FgV
bFQvnuIOWlpn7GVXMIWXxhzSTcPq+4JrateiiUoCawdLFiLVsymGbOpoNEykEZgOrAknYTiIELvO
AD7xgGkmANbFigBdAgK81ptGlYwz25tSN3QNKwyD4bE9gQYlmvaR6rKVKaFLsv551Ltk2kasCM+K
WH9yvbS03u4nDkw+PsvhZzhsrl9zV2r43MQR17+a1J2Zhp/DJb5Gz1G0VL1QzTO95S7g3Vjk78Q4
T/yiYCDigRge+7xA3rF4d2OxN621ofZHD8iD6lN+/KSVLz3lmnE7EprF8cpGwxI91k3m3p/nawq2
60ZrFoHGIUBVWn2coR8DDIUFNIS4IQvLHmMP923pAAnM8912L+FXSpP3p4CHQNBn2ihcYKNYafef
rr06hkjvEP0WxK+96wKpHRPS4FME2SHBDkHxuIbNd/rNIuR95HWu9gnO2+2hxGnBuRbESx7KQ5nu
dh8MPCUH79vNyAgRIOIrP1jFRB78VTK8HlJalmg+PaZm2B+3JS9/vPS2XUtAKk8Vw1t+ehG7ZP5x
Hw1zysbiwbeoEPjRZlP5NGvy3hTq1WXZk2eAf0hotD/bBIJcgIMCdDqRl4PNmPcKOixU0bQf2Ade
uLc3K9fES+mVpckCZrpgbwcKMuxO4USrmOqSQzttvthbS6RdUFjzgfC/kTGR6u60qaSiiGPsUUXy
mZbKHv027FLqP90UfzMS+PDDjOzHGNkEe958MK83b3FxqKegIG6pTpPycpU0EIdvGuhIOO+b+Pw4
XskPq7MfHi8TwEY5hB/x2nSm+N3s9aOQ3/DtoMtZV+aId4I6Qy98yWZgrZ/S9GTeOMpT2hTLYR+R
FBAzFYxe0gkIHGvEwxpP+Bz8B7IwzFQnnp0K2yAr+bJCzNoPP9q7oue5K86OTqjCei26/GxasyNd
QF/IcphL/QiWQwuV/6KU82ebKtJdZJ9ILr5UKFBE2CPZE/XGcBJJJ3Z+EKVWpdJllk0+2B/yKR/F
4PdRjROi4nPKqsQ5Ry6uva0+MX5LRYsi7GXYnShKgpTKOskxfLMRAPpvfD9YQIBq1veloOhclev8
GyG2zeDobRG8uoOpiFZeUfz0EKqFEfWxMpYALUl6VSLD1pWkWzWdtMemoPwdIkBOVzrGoQclEum7
B5qhk7+h8BtqRkPfLYSBMd+BKCtJDpOpEOB5qCR9yg2/S28ts8lRgbMLKcGD9FejY9int/gBmbo7
0MO2IHLmVLg207KhQnS9NMIAu74QHcoKEfqtVhUB782yZnRryLTaY5j2j+IWsWlFXlAb9Sk2S33W
a6bf03aAHvhoGG93LJCNpNNEaYBMRuCDfhNAeP0G8MzV5Q0BWE0hFj3iGfet6DZfctee8XHYlXRU
sTbw+T3QER1arOF4ePnQb6m1l5usb38RK6XvWbhBCxQiYFElx7q5OEUyncb/wWaG2e3nj1q+IxE/
8hpUOVoPvgm2cYvW5Lrm4G8XTr5mfsXyQUP0BUQYyKAINzwZrhAj8L9JmMLhJSE7YOpeQ+lqXJgf
Y1kvpgfKwHmagcmZDkzZF8VciPw7KyRiJ9V9BSguL6Kjf+JveGA35GsOgOcccTqqqp2wRro+UMvm
/C9n+udN6p6YzRlEVCiw7IBr/LMtwPUjerTmxN7eB8Nuyug457KxHFN5s6JOV5fgnBG/4BTucJDm
0FwdMONIh6o+hbMod5eWdZzq0RQzYholgpP8avEc2aE7ynuHJHGrTlCwZkx+uxMtyD/0OCuUjzUQ
3yY8x//6UUmeMEjjK8BSkcGx2nOKqUWaGgMEOkQlrjSVJdGQJ+lG9k1kq2jluBdGDxMuF1Zy1FSU
aOHwwNCIywUM7FkK8ZoppTARPd5xnYPyWK2wrHGTOG/I7MMJ3/+L4IrA7Q6n6lLpPdZJqbYLT41z
Va9rI47SEWsDqtr+8aq40PhWWl5qzWgjl7IkWvoe+Um9hFONJjBfQyXLSV4zV9pyfJlvf9f9OW7X
G9sj3z8xjBoCA6kER1fGxugGu/h8hfwnPDMc2srLXKE0J00UdFCm6SK4WayjoE5H5HmSA7n4jxSE
r9ViXSGxjxUE4PIakgiiuZdMv1kV9eIWIsgqamufpF0RRSY2UrG4HRHBBkF+HUaLtBy34yieO7aD
XkM/ud12GRKH1SAHsXvinFbaYdYm8mc0KOi+kFK1csliS6ESXYWTxMPwG8aRtIMmt0oi8TjYsdck
+7piyu8PHlVPw8fNSsSag8OMZMzGQBvQSC08AKVXTufMD+Pwazj8aVvWn218lqYZEXd93T5CVhZD
akHLfU8al5z2biVaU7ZMNdI9U0y3emj+NSAwO/HOq1qTQQhsaC6s9cnuvPtGlxlALgoKUdNysojJ
LqMsXJFbrxYHvAxmH8tIc6WjyMXBjiiHaEUuPbMQngFlXb3tvbvLaHrx/71D1Ad/OaFT0mZkHljw
PN2bd1tQiyHTxtgmHk6gDXLCYgoDHTT29rv3OyJYGNsSMuWmYQyxgWmotQaGV++sOm3tEE0h3F1R
tmOVvaSGNUhFve9+TcGJhk0yQWOnBoI2m+PeIgyNhR9LXkNwiEYhvhmFqEe+Lj6E8p8HM+LIQ8b2
pS4lcASvjKGiqzMTNihcO5CpxenyT14NY393EgeZimvOXoyucLWGtL5UbaOySPFS0jFnnFwyUGIa
QW4vCsm4e10J0pndZdnCaT6u7IMKhVATp4OlOyLt3UiQD+pRREEnUmubqPjF/Bny3rcvPP9y1XmD
+o9zSF2GEfRZdHwhLcns6MqdYroxWsDkeBhn4D+ipSxdsFpLkZLoyiifTDi4RRWvFCHt4qncB0OV
cJ7ZwpwyOq3VVJltq6O1Hz9DIq/4yERg+vhvCf60pcOJDpamedN9yYddnibdHAe7soJnfk1HFh2Q
agjAmV6FmB9cKBpV2NwzpfkQOTvmt3kNpek5LDYFhyK764zSLfsbnazSxoQ2fjDIFa0rw2L6p14h
gBPU6xqjimiESo1EGMpNSfeE8iAIywFW58PXnzsjkxRsODT0lPybCKXsqOJSlNj8UQTq4uHOqjOi
EyOXRLUPc2Mzki1tCPLN5N+nuqLVErHGBay5I0Un1QQDVRQd6vtOzhAF7xXSXa+Ofn+55TMxsWlV
Wy9zPXUP0VLgYooJTX4gPe9AWmtpfDoAoT1In2U9jE/iGkGvQ3CdLa5wjj/u2N+duT2qKB0OHTIA
Dk/lfzKbG3+5I15pu86yZ31v+tlu4OyWqAa2T57TZTrdpaJ3o6ubVN7MWi1usNgaWk3zfJqUGCkB
9GrNnII1ceC1wScCru7Bqssoo998D6QRKUV6ifn5Jj3HZFf6ACFhytM9B7Z+0d2AY9SUS+DbO+Wy
oyPsTpJblUBW+7LwTSPPfCgg3Y13uFalzXJPoOyz4s4jKitRdrqxZJsWLFikKG/fT7+xQgTNl9y9
cOpDpQhNeh3igib3KzPEfqyi4SRjX2Jn3vmSJAtF747F726RSREyf/0oy2ba4bLq7dumKqW+ubt3
q2HKJn0VzOAbbhimyW/f7JTKXN7tdcZjCgNWHWNLGAAeo3ycRnYoPMB0rXHIUhv36jNnvYLspm2s
HhTYP0txjvJjX7Lz05rB+rdib6hRKaG6o2Av1wly961a8jAM2a1VLKTn44gKy0tvBGhvdZE5yFaN
QGaiMjo1yiHxGBp7i1rflm+HrJnqzXN/J24OogSy4dhluMVHAD7o4fttWIbSuSXR1HYD2LSgKnmd
JN8YZ8Y4hYo5l3LVLTbfSgkVK+YbraIp7tbGo9wCvams+LL4qt6V+f2HqHTfW7yFBrWMAHgr91pH
pHGhffqc5qbHf1tbIu6mmT2PrvuzP88qwmCvu7+5uYqkrqace/slBzPEVy/MB9QE9yeCn66zOf9n
qhF0d4oKivmvQVb1TaYnLCpyWubIsNqc4P76rGCvawTdTm2L04zxIxDRf9AjvDvoYkQ4oeIuyTs2
4R/gro85yLYPBVQcPRm/ggBRjQW/Xduq3MMJiqUOqvS8NLuDF07z9tJDP3adzpX4fBUBY0IAiXqM
Lj033WEs3PlzRr6Rll7rRIllAmVtV+kOi9ijfzsNHYKx16vqsWIYdCsU0RM1zOLpzFJxYnMTPJ9V
UsG2rit1eHXw5MCz1x4TGiy/UKcOSJZT3T0SkH93G+ccOstI1cIyHABreOYL8JTFQlz4ZdH39fJU
sgfdADV9JXz+hXQiVblQAzSXf2uJxtalX9eVroMQ7V2aK3GoQGSRIg7H+GkYT7PukbX2U7mJNwYe
q7qv7oAd5ATdW5DvGn2BwpNXlH4/NQp00wE8PdkjtcLFBJnVmGZaccxpNBsykhicbVfd86Zi7bSn
A9tZb1KW4cWOfw4BwVTzvHx6YWekT2KV3XOjEO/XkETz6Gm9t5iuEdNBBBZKYh4YnmihaB3ROKCc
FzFvUG/sFm3OPTC2LS+Uht1mbD55Jhet2Aov1GiDiyMikb+0Oq5PfDtvQpxIk1Feou4BeoP4YO+6
McdiqQ6heNfY93MoIUsrvyCDbExU7ZT7LKTOnytbsw+BHyuivEzzXN0QzGsaO1wwPxhDmQ8RzqkO
Oo2lwYCbhC3a/QxtYCafAm6LHVu/vQNu8k+UM5PmHpxaELVuDDFUmKnTxRhk0tdB5EUmCHX9+1cY
VAJxwlpe+tRwv8t40rKJIQxheCJsNZPoenBZFZI66MSm2OvwaN7VD6i2vEH3LRmtWDgPxP8VDVSO
qmZWma0wBR1vPUDEVNRGIsoKqBEuLhtzFiMFJ4IZr6TIZHkiJFwq+NMWNUvHlaBRpTmOzwhk0KgT
D/GCn98weERa1Ns3vfbuOWpNd90BLBdlNnZEMpX+7xWFv6cSYEpz5hqvqs64qtFOubL9+NXuvsK7
qPeCneDNM7HDOxrdoLw7J+/WF3h+eGCey3ltvKwj+o8F1VaV008fa9+3H900kbrwN2FTB2fKnXlO
LLPHDgsPX915YVq0tvA2mLrr72Zm6Lcl1mYNUHu8HDPtmd9lMkpBQCsijQgk/d0rnMNotLmftbL7
Hy+LDEUBEoCqkN0zQ2FJVaggmFJNMuCtS0/3ujY+3bP24Jn+Ndymw1Pa7h6fO5qvMevm+DZm/0Jc
vLA9UIm32TsiK7lJvf+ev8PADUALTZc94wc3dq3X//0yrVHY8NWuVOiW5qp+r0gZndjGvJ9K5Yee
vDss002o1IbTjUhdGkH9Yh0gwpj1m4kw6Bdj3dL9IadK6x6Z3eAg/JnuC+Bw7MS6FFwCmBnuwuGJ
BThA1IuRA6qmcCoxfJgLlOtwmkPzzJdev5CvQwy2C5PBmeGPY4PMrTDfHw7E1S9gc6wpxFslOkUo
TqBMoZZlHa57wN27gaNu2jsWAXaAqXcNZSaeSKmOlrsZ+xs8WOrbtLzk5Qt224Mty59ZUosuZKJg
jY7B/YjLCVwZScmmZU9SW+ftxYr737FrSSeeYWK+3YqlN1k7BpfXqTx8FGDNE3j8IAl2Oodu1BoQ
prDf0CUpUvYBVDvufenn73TMYcF1FKQ2xubH0E37rENA7rOMVfbLGjbBTYnDoYhtyBx44UfvM/wA
NL60iLGi+hFovauV/uP3t6MZnFVVkJzjGKrDaD4GjEIQslHIVk31h+0yzAJFays/dBvgW/mVcnCP
srPz/r0qjo9V599v8mRY0AIYI3r8kNoXXQPVZzom77BKbYTLvk7Pw3HSG95Ekh2GyLqBmj+xo6CJ
u55LuHdGC0OiwcGnkDvQBeboy55yBqKEAsRX2PS9KzbqaWnmMEduPRcyPJcVZrqGPqukqyVZLoCy
UxsVFVVDfz31rjiCREfN7rgYlvHuf6MQ1c02QfupSoXnwB22p6/K9BQy7dOiCyECsujU9xnfO8jm
F0ci88UhNrvOTQ5+W7fZHNacoqk4EsEgRkJrXlysYfHE61/oiWx9XMFMfpusPs3d27hn1+xNDcKe
C8OHZMVN2hMuL2i3W0gxoqvK8FAQetutgh0toyENwYcVbiYlkh1vuoDDngVbaZD8CxeHv1o5CeB+
dGtUNkbZJ8BhBh2yEPsjtY2BjhK3Y2Brwe6QvPgV/yn+qteIqoOS8Tjd596HuYBOirXVZ4xfcy75
ZfemwHjviDcrWshj5RxKre7uyMOoWv8BSCjzg0DUzGsgGIDv5QOCMhfWHVSU0znXx6hiyxZFncvY
YZMOSGpQCkEiuoFZAvV7nDcISWkUWNUvIZFrLX2uQcJphYulIAh66ZBhNYM9MuCrGScubdm65X0p
3g8k59NwrK8S8vCEPFywqjKzY/nDeMX1bfl1fRBHdIg+83f/BvPQpq3p0fA2cBG0QTHolgdBRGOb
ibTb+We/UBEwsoFmi2Gj1BHdrr3CU5zOpriOuhGPQ0Es+JSIoiyYVypQtisOSLm3ywkgiVm4VJvr
rRBcne1JXND/1LFJZQVXlGE4aQzMcgcChzelVu8TfolWQgqiza6r8OKqkXb8y6KSYG293FnNrAB6
RFYaUI/wc+aLraCWgtdYAZUGZilczxFrMQaD0PiiWQqqWodQKJo08Rqru/aruZyoNh/7MEz3nQoz
DNKF09seB2jYfFR7iq5i3Vsqst1QcIRbnPLTLYaKJg9eoyLnEu4TdbXSDXKyq4neAu1rzzZg8rQJ
wH0CY7gLCbbPrUmIU2G/GQsl9OT8K5Is8WJkE2T4e0r4RZ6dWhoDMQlv8ZikbF1ka+Hq8CQX3HWe
TFcal+mlA2+mxUEK2DYX8ufglgZhXAL9l+re0LBvMxwL/9r+mTeeZkB2NUe0x7rZhm4h106E5hiu
kMFemhwpLDRk4Dpi7w6aVl2mBqEZgUKKqCNf04+9HeFVsPKRL1uKLd7dzHcXwrwB2Vvv37qca4aw
JUcm2p7SeLUiGP/1IlugHF71l6AB1/mufrR92+zcWXYs8rnKt+0X9ah3xJV+P95vn+IHZ7MhZF3/
0g04Rse9AgP8zpD8GWiEkYq0inamVBulhqQnuz7nTjS+CO3XGOWQ1dBK79SyCuYoMZbTFdQURGpO
byyc6Eb9sB9yTVZqULU5mkj/yHlpvt9Ad+gDlxu8716zW3iTFcWiG9COxDIYpuQJk2XJm4ZKOQpv
0ak1K76bv76oHp6KB21giSQDdSBtdRnzzY1xp+tz4tdQOH2zXBOGShe9HXzKHS1Rk07jWJXAw7hL
pMXfPABTDEITuv0mfM8Pndq3B5NyLhj68RRrcv9Bc2KXO8yqGmyURg0gQLF1ndH0e1WAf9io3Bv6
YS/ZnNNM2k2m0IZSQDwLCLM1I/ZNZ9o5UN8SZA8UH/rf2VKZlP9cQ5Oxvo6NCTIH7YJ9FXH2MAcX
9JBc9e6muQMo38K3zAHnZ5RQJSRKYoJHlBkKBO5ObX2CvF0A4PBozM8HVx2Pvyysz58/lTW9wApk
f1C9NBtaatODSJAopxs0ZhoflWfl8R5Jv8CydCKiYVWklEmlmWwH3M3Yg2CLvvMP+xVXHjBohIyU
2g5xnMl2qozZrficicQGP50Aj8+sTA1JCd9BEL8SVFDABS84l27B823IDnh5iW8772oENnTDBKQ7
pudiNuMHN5mMpv5vptGs4xzxjULzyVzxkuHN0JjWONNK1J4T2aWBkC6MLvAbzuJFCT8PimmSnA4i
K8oh/3SGOJQWr0EFogCKnkBsQiWDq6YI5V3PxZY8cpaFUVHg1+5XAEcLbbQa75Smpeenb26mDbgW
Fryn50I5GIegqjGhdlp2O22xvdYmW+7+Oc1cw2dRP6XCvq6b/Pwe7dq5FcMvejk7ZlxPZCqBnspP
asOJRtKqw3DMRdujJ3iSsZ0GBNDzzDoZ0fnKvHM6U/uhCbRHRpSzkgM524jH3Oa9nGP5cDsMGy49
yNGuogLSI1/kJKOE96hVhpE3/zefUcA2r/KKKogxibMOGILPp/RFKn8k2D5vDzsvLlW4g+VITway
j04HqYp8yHR7go5GD3EzcqetEeWmmS3IcSXKc8OseFYMfgB38DjwW5ND5gTswDXn5y40BKSt5LxY
vAHY6BqKWC7ZzzGVKPfgr1wLZp3qQhAzG5AUyvQb/XXIVQB11ypa6tOvW9VqXMhgnVipN/mjoMHm
X0voXLqmEUa6Mh3lNmUS4wgtWxZc3P5ROD0Xa/pFT4TW0L3eE61J7AeXL6B3bGuH7TKJm7tNyQrV
MyHGyKh+ISBBz+b35nab4wFp8yO9+KXU7aovgVORZw90VLZEVr1Pz8KbvRyAbyKm2hRBFbU8Wc+s
bjg2irqJhwHquv+PbV3KegtmxD94oGG2l4jQGCyZcxkr97zKT/HlMXzjS3vRb3R6ZFcq7sXjlLd5
63XtxUddRsEq18VKssUJq/GZiSVnK4yygLrlM6s5DSSEqbG5tocMHknKSpztmz6acevpySoHYjzH
S1SKCON8ZLtxyhtiLLXI6CByfmfZPPkCPjgfaQff6fugS26brUEf43CCVk5ZMULMFLXYIHClkHR7
8k8jw+TNv2Fy9byCrQPqIThc4yuReIBFz3pE57h0AgmL8JaAwsJ0sOlDA73HfaUQ+EFKE6xsvGxT
Mzng97D3XyuW3xH9y8mOxxLOvsgNVpOw+WGiSB5SsTW1+yrveCmkwsJvfxpOGALoUUENY7tVJyT4
n1JMezgYvxCgRCeen9JBsGAMSrM6/LO/ud73bYKASHWcZYnHbUXr1WtCEfqcpjQDk/yJw73aZ/56
lqlKJCk7+X9ugtMYyqvWqIrhZ1avbE2pmIjDPPr//exB5Yj0691+MgzOC/a3dgU5Eq/wrBfHwmgY
OqgvAQv3fmreMFGCzjZRuLn2WwJ4ehX5ahQ7iZtq+GBOq0j4hFA0iD8PnkSHHPMxCeyH4WXYgVvA
62mP3qrd3Yy+4UsnYisiLt6UhRerJsDAmAR4MuhV1sefRPVbbcim5mr7kUGC78a8WihjHRO9b5y/
F/zjYxURuvNmNlNVreBssEP51ynHtM7xtnNf8FKz6Xp9h+0PWeQYkixjtz07zV2yEozoKSer6HJR
FnomyixsqoCsJ34+NBYiXjm3AxhWswjxbgVdYjQXerOmYVqKT0gDJIgITOXiBBD+CV1d6ci0vlyi
iWE6Uw2/+p2/IXqoaoRjLt0YxbSSAogRqtr7bx/yiXiiTOsk7XehnlGlP9oiLfKpAtIMsBu/X/2G
D/t07TxH97TIlYzFAptpVCT7yxnNjVJSRlEJX2aHOIB7YF97EIjnHWzlmxgh8e9C4S3QP2CkXjBy
svfj4mVbBNo9elTR9TanS1deHIgEjIBlmjypXw6FcAfnQCFMoVckgcMG9HYATX6SYJbOdDYm8icP
3FbkXcpsoJ+I7WXQ5LdP14wubQc0BZXRGFfX2uhGhQ9337sKRWC7WmHJk4nHRkvwhycn5MyeQSU4
jihrKWfFIKLboC3UzAgkN+HtR9O7TmWZOfH868LbgwaM3Q7vEzVELk4XnYr+9s6KB5RZK29cb48U
vOODeY21+J36I7GMQ8pf4RK9mGo3bJ9DtJIGouVd5pRWIeYVdTCZoFA3FzJmtDo9o/yUrlRpq+SS
+6miQ8vOw6j3ukO+L5ZqouMUvBjsl+r2ltA4fGiAZcoMWUr1NAmgLYeUEJdxrxInzeHC+oXNeljh
zZDXUT0VjLLz9nc/0haPop7DQ2HxVtWxsMVMA60AxbbiOQCO1SumpfKD2zEY/B03oRjEISlOV2bP
YXROUw5b1HvgkpIJNYXVlA00upOMk4Zepnt9Ayyc1E7wfcDh9KKQo1HOdnnGPA8zh0d77HwtGnWf
RpH0JoEqawSfA5WagWvAHHfcjFkMXVIzzwj5+kgYu0kFDTppZ1UUhXet2ogdGLADXTlt3+RVaoKo
hViUI/HXaQPSqk4+OgRXvjyN81VLt9mLMqDV3kmuevg7k0jS0NG0zrqe64kgmQXMJ0FQrQ+CHIVL
8VBB8eJe4GshTYT3p5Zni9rLV7RFBRy6FSeZKIMx9qML/mbAYTuOC3ncQfqIHc8cOMthPicQABKQ
LUqMAxA7jgpZJ9UFNaX1IbpFEJ4Op4DptV75LaUAkf3LuVXi1Fnf7/I7xBE+Y+6EetmMJq587zcD
Ym2EAePStWpVVPpfwY9yqnw/j0HMG8Nh402EK/bdBTEhTdGNTOvI37yuI2EfJcjTMsnhe7tfBOlI
mQtcFzl5vn7eBjWVJzNNPEQCW21DEGKjNlyD/ErZ0cwEyAFaYFXR7aVwUL7oHAdIwyLrEtJYr085
qts4L+U07gcrRu3JgLkjR/nvCHXFuv30WOfh9LHie9I2wg3xN1WbsTvAKhdHzmBrrJdeaCE+Rhq3
K75CYLXPHQoMje24hemdecQJSKJDLn/5gknyw9WyHV3erxPzNwSsN/hramkJOE6CFsYvGA3Pt6mR
Qr6S08PJLPonW2cJIL0EE/vw7/hwtXfcuC/RowcHXQEygLjagFUvJNRGKvVwoZpGN4A2ZeBUOZt7
1CG0GeacQVfrZniN6HtqpjIZsLEOV4a3e+uyZvdCYmZzRAJAKwUk1/65j6IgUKZ4RF+ZuYiYM5gW
eI1UgWHB+oHAA3KsY+2FjoBjpgiUsApzk77L2oDRygRwNofgp6riSBxBdeSvdqaZdJTcqZGi4P/H
WNX80McgJculLVHRijuX2OED89707uIqUFySu5hafnfSffN3EEidhrfFxmfeUODAV8Wie6NINYrD
O6CbK5BtdqDETsbKlocVqV0HYehLg9sLkinrTosNLW7bBXPSoK3yv9SboENSykCg42b3bFCdRiqM
jM+RWrP5OYZitO6ZqlTP3IK3F174FFW1VPv2PA7hRcYfQ9D2p30HpweY2Ry49FtCEZN6a6UbB60z
1N4mYD3O7f/LRh+nvPg84II+Zlu9pyKJJg9yZTp/3TvbNQNx6Ik9eKfEsRa1tmgK+Nspk6Tn560f
vP9E2dd9N3KabFFt+DOCAKL28USduHWajqTNUrlgOLJGPfBqrn9rwkDdrSLLtASrRqfdgQdbd2Ql
BecKEW+t8l91ftbOFGOdSuQ7O5ldp7YS8jyD6QY2P3t2tePPwkEfeVJeeG4KO7EbXqphAzpBKYTg
mZPoFWayifgi9YJ+mjmuOgqC0mphzG9lDJ5sJeoy44EM1pBMIv0TWesNtlNY1vduqUqLbMvhoIDN
NJG8GBXjS1v9UUjtpvdswf6zbIy466n3OV1AgQt1iaSgMVFqcpo7LKr6kwNxzP3RCJJ3rjVCkz1R
7x3O+Yi1pkoxNWFRKNJF2nvDh2LxSSa50MBlPHk4Xk/Mi3EPTQcWSufn4OOS/JOz5/bIJ9tfVRUN
R/doWEM10yvO7w/cLrC/fSq1suc40mvBJqEtF80GIHUXArII9DEHBCqDiNUMUzpGBN+gZ/eI2TIM
NM6q6jcV7SBeo2SpNgyRXYKJcqrJQlgeL+2uNytpie6u1mAyoZqroE3IC/LXAaqJCjLV1AxyT2KV
cxh6ojQEKjYXQ+7FybevhBcFdlbrAp51Irb0LVI7X7lg54uRp4huqym8XXVwE7n3CI5ay2KQ79G3
AjBoM56jue62I4P+sWGbzhgWcvkC8Q6T1JAy0ihOWslj075hy0kqUFzSfxEtj4e0sbh0oWYO2OZP
ZdG+LCDsYUC8N3E+JtS/kbfFF+9EfWybxoM6I4fjldLsoBxyGl+WMhze/qOKboMK1lKuMZU3FdeM
RUG6VUkBy/TGZGo+8XFeyHJOBQqt6WUdkA/I9RGM0XobbI+j7XfBYp0J5tmm+EpPLAjBV2pyJPiy
M420M0x2pdRG6mvx6a+46Qz6C9grlt8XNfbYwpvjVcSkuLR9ODVo1BSuYdf3SvbSvP6SssGfAFFC
Bin4kWcKSlY0Wv9JZJ9VgPYi+fnaMfL1misBzE3R9tTZbgnSK8hC75EnSaJBloJpk3ibU/9u0DT9
mBwdBHwMk38TkKFqGDmtAmnBhEHQ2WxIkKEFBC0rYS8FANHuXia5q4IsqV6Z9ycEJ7MmoYR1nHnm
AWL+Y7kWSFK+VWpaNh1nb7Org3rFnUgDS8w8GCbxIU/hgHsrSCRt3mIHv1r6zalXAUzMsUumRL3A
YncN7NXqskQBfrqXL1JwsaITzmz4MPel9PGiO9dVvgWcIw98aQxDJQOGYamnL+IcaB14pUdRP61o
zQkrs8PeWWBb3MSKqVcO5pKA8i65vjHY0W4+QNOZM1i/hmbI0xxetaBkOLiWyVUyg48s7euFJCSl
vSVtEhKx+5c7kDsgmjpPraA+a35kdDjXyKJVUOm3xDGFyb2zLqFb02eL7IpInGoUenjRpntbY6qd
sCyyZBdoQo7pAy1kb8x9I7woJ+wRP3doeiBVBzzWRqM/6DCnwKfSff9UL98Ex+rsQZJ4v5B+kyIn
roEgSmN68F2Nx9uUmetsdcn+RAnfOAcbbKhpoNbihCO5WEA8S0ssz1B253Ld9LFuPdDuEb2zmgls
Cbwsf67TROVK8uDKekNauK3KuSO8zXzB0D8dZpOFzPaastsrZ6OpW7Oe0a4oYji8ffci7dtp5rfS
QmqXakbHCdK4gFBrkoydkt1zZyD+mMj2hdC9Ay61oUBtsgE01BUSPq23Boc4JhFnFC30oCOtgjD5
wkEOHMYacJB6nihBYMP60RtaWQkBhtsbKnIyCJkdvOG6605CtL1zyeUvn4WuyDq+XUYlMEI/P/DV
Z8M/CQh4df5SqXsjx3hiCA3VLx8Ss7GXSlbYCQTvfajDzH5IRlHsqP+fgOSa4MwSJIn0Uk9sngTN
tMJVmpPN6TyQmF7hP7B51ycw0nydBcupqhsIhoiqDMJMXkJ1fX1OJZl3s21xHYmfSZJF6jzcHDdw
K0uUpSo2o48b1su4aK3VrMn/rC0UromKpy3faJZFtqvcKdW10m2+qCSMzQheYAVahUjfWvV8krvI
O0KA5fCvz+SA8sE6N9axr4y53esq59WUK+HpqxJ8MKeDOUpQX58jjMdRfeHrOw76bg39ECfL/jya
IPkdktM3HmTAbJbr7AMmaex9rc8DbHQ37wxtp2szfHYeopjCdjm2IpcgHsMSI2sSUrssKkxYm4TP
0R1qHcReKg8yyfyrQ+4axFz+sD++wwXKe5kOqh9M52kaGs9A7v1NSZvJ2wdcCvmMBgy1gxL7/+Q+
TCr+PFvjcngLFOTvb4IfPKOwbVqAWKWclx8BESHvGrEmomc+SYtsxw65CBesgzUn30rMpoQ6mSxt
S5Lm+5n/dhGUw8Hjm+24EN2LIoHkN6LfagDHWgTq7XMMpcDVE/5ngI3sLUqqcgWKwmqULr0Lfm7g
yux+ckeiADBaE+QTdRmMoTlPrWoOBei/64nOhF7Zm+Ks4upLyjQ4/Na2Rwg6jSqsNLA9rmgcIw31
lwsxiZoOZuUBIf4N2Lkfmz6DPs0WA+3zD6aAk98R4tocvos4ISWN78gO+Jdm8nivodsqkb1Nmplj
wDOjkB4tzhYQ3rBa9hHiCwm8GY50gEpo+8n912xVc7rWEHKBWLBFhItuOh62CxaBMEhbcAXcMNgz
ow+buL1nQWb9sFGm6LOUKLJvxOh7hcskb+/V3WNU5vXtLhDlZd+lFhXOYZSwjilojPeCI07xXdjm
hP+U5qsEcRjrwQLIipkBZIqlAZgtqST8hdkD9KsMPS9JKESQhpc0npTcEcwXLaupFn+hpyNOZrga
Be+nCAAaC3mDucSDAYuX4WLW6+i0F9YY+crW3p7UM0eQsgwBf+q6AhU44I2H/uvcSGK6EYHn19qI
AHVNixfJMJXfDDsSJDZ+0+W6z0Xl0FDe2QQD1yeSmlfGt7iClrvlgJVbigcbSBe5uvSid8c5q/5j
v5IhR4OzsvWyuzoW5cv93EppCcX68Gt1zzXOUHM5f+G+x7oMcoTgDv4PKfORuhbrkkVV5SNdAEuf
W2JcPF4XbIH4AmebINtozUe1bJIYdD4Ph/O0bknPW4WK/YhO782ESinXvPsX6dOpr4qRqBiV3pPI
rOMWAIwijXqtC4UJJA5VErvFWmwnib3o4/V3NTO+Emv6Zx1M7i5rSBPm3bt9N7xl7ozgbeZPdeDc
jTj43ngH51CavT7g+FctgO11aHI0EEooUyPrwmfzYkbuJWwNlCxITro1X6B0Yml+D4IAoyMSjzdb
2g42pNALBBOmGs+CbUhq58fv8BBK/WGv3jRt8nGDOO8vG74bl5V5pzRkDrzb8PzFopcEFlu1VTAK
oBoUrsj6UtQ9wylsaBzlNnXVD4i5dmmhuYDVH5tU8DUvMHZwsVQxNu6JL2s002G6degXa5SHHc0f
R7zRNO44ExgjORyGCKPp481yP5aRep+WPXV6Nrpd0VRjE/PXPUozXVFgAauKQ83lV+Sc9PluKlIj
edUqtY0fyRUgKFzgAtRmFadAhh/lITzu8a564nPpX23LWSOKluZ4dMVNyEJTreIAf/J0svg4yR2L
KUWaB2X5nmNiuAW+sPUQHdRE9R5OL82e9u8XXDuhfCx3r6lzE+A1M+aVxpeNPfGG67PiiJzODIQs
AiB6UddG/jkhAXO9lE6KBF8VEmXrgHsM1bFSMEFtp7VtI2tI9eyM5Od/AQnwGVTY0ZigaHImb11F
A2CowYqFty8aMq6c7GBh5N3lBwZwUMDIbLtwHRAbu6A/74YIYZ8wouv9GtWfGIwyawmgTsId3f/j
eb45HNTq6xlWsDP48mNzQmy7Ll4J0z68o7ZZvrESB7Hy9XPLOAdK6q2kOhW3+8b2pp6eiiuezmMd
ykNX4XRB6lYLufqnc8cf3n+VV5SJGjVTDLhyC4+eI7x0Sgnbc+7ANZDIdpTsky9xoUQw8JfAQEbn
QKJk35vui1W7UkvtOlCefbS8OH53tGdSyLsjEL79LzQeXbQQmq5YjqNsA3Rc41EZAzkeObhVRZMN
JWrrVO26KSOv47NTthJXNDPo4GEAEAMlnZ8Qd9Voshj3CIlGGRIIQkQ2U6q3UQ/LiSWshJfMy89C
w4s8itHGt8j/0VVxGm3mx3eZRWBfAZZuKpkDET2ImIdB1VGTdRMPJH3gCA5Wb/1R/QXmQYTf/Z+7
Igj3S32LLemCehQxrHM2zNlQE0aW2QKVi6TajQ848ONQqkr5nOuvSIJtGnspsUakVJLKf/Eh/++R
z/70f/tjaOnqLYv9AN18ZT1DANX5pN0cn8dyMSIgObBqUZcRGk/X/0Uq2S0bKfWcVcdWQhP8uYVW
6goUDJIcx5VolwfDa65FjFX9E9xJLSxpqLjp3c7MxlFgLKkODec7kg/GuZKkEhPh3HyvVdIwi+2U
8AMLpytMnEZyU57DyAYts8j1J0ZY13kTJFUwvqY2qupZVoBZedxj++ZkCOt4aHxbE0z36ELK3son
HQDu9B0OisQz7bdOKatan96d2ANOsXqCjQFpwGia7SdqoVRoFY4M877R0KUTvqbkmv5VhpodB9cy
u2Rj95DIOiVzvS4wT+tcAdqPkeyN/Phehq4MGEol+9bAmLyNeKBZf8+whpnL+tNofCCtfdCBUtGf
IhnVW8rV9QFga8/2gFBozR4E/PIb/e8w22JC4VgpvoQ2pKYtoTzxjEdnk0vcVPbRPrT1fXOAHaTD
kK3dDM0O4TtQwXtz6Kvw8N4oYIuMoCbbt7yeTN+WTOkJa1FGek/DB4rrWyuXeOvbEUgnuycnH6+5
5fFPnxHfhuJ/ewNGserDVBwQwDz+e9R0XaBYGZR2Te+mWHzucXY3zknMuWipXwrTgMani+ECYJ2A
mZBnSlSyanFq1NC7Z6ILXky2U0sXaZ2dqMA5B/c0VEGiZm9/1kbTM9NwoOIzdRfW4jf4Gm4RxqAW
vnODq6z+t5cS5mgZ4n7n+9EtWRfNofv5VHzQtsJ+3b6EHKMW6tPY2xfdghIaxpsdMmgUhHzLpvc7
RPnd1nSgqMBbJ3enWhk5+52nlv2/Jnl7Cd6jx7QJNjKn2izkaHOTqXAX3ky/fWFWax0p/5POO/PX
yoHfkOEI7zv2LWLl2kGM31B5+PsPMrO3WeuXJzcpzS68T80i4JAQ8Err7EdiRqYmE+fUhrb2B1/L
sWufebckZcg3Y811yK6C4BeiLVJ/8hpMN8pPhmI6B1QI6x+SGSWC4dufgq2UsMT//cdiE/z49tfx
/SIhTuumMiu7o2/TGrMdo+Fu0bagUqGBvifLB2rfFFUbaokoB+fxQXZdp0OMCi3fedpEJ7W82DC5
jgu1bLXzeGAQ0ol/GAgAcmb+JbuNh1jOey82BHiu4mQS5PNXqJAEsQCJPDxL7AEXtloO6sh0/ARG
HBppXmp38mlFAP3xEMuhb74S6QPCdo34JZmmq4ZcCCwPidBrHpIa8rY12kjNuiLEtNJqxwd6a9wM
34IKFqN5FryStqNrUQzNje7fTv6VvOWd33Qy5eyoVQKHyLD9VRBcYHafVKpQ1gGcuJbyMSGihE2B
E1B6ueoJMX1MK1KjNTzg8N9vOewNJKJKrzyi4N0AhjQN2Fd/C99uCxcp685Ie9spUwA+lvKoeayB
H3p8XMrWBVQbEja9R0zprIq8BJxGNE87gz7pYkOVr3/xh2hqIn9AooZoz3HkmAW5jdHAgLcx9E5+
glldm9h27UxUmMzCkHX9Ay+7gcMpAhvyftReWTcVZUXKyl2eOKYSRNtiK3GfutkAgQNkHejOmm6/
Eo8q02PuZMexOxVrVUGqLpe4C1Saabn9n3s73CEbPvKAZaBcsNW4IW7RKxNl8rLnrFO2/VH0hwhM
G2DYQbhNhegW//NifBxBUeXaZ8XNnY3qV0GPF/b6m0Ljgh0JE+OEIBsz2MVu5LfXjPJdpsYEE+PT
GVEh+mWS/fT7qlEx0388CajemRf6hciiVIRWWoj+62SAUMDbv6vhVIQcTOXkaiJK618ygZ5BLkNJ
GFkjW8X7UHzCtWVB2Ss+umvGwZ7SMFXbUCq9Gph965GWQF8DzOR+1eR9HpfFTKCZrsWr4h/6baRI
+DE6jwA1QY1gh5fiJ5K+TlKHDFs5nN3QUhlCBoXiHGIqP1pYwlsLE3kxWmNqWLHvxzYQRQVtMmI7
k4gI7zDsnUF2bFF21T688Aup9ROjBllDKKhxssePzq45wDrEFi1ROHgXIPPjZQi7CN/iFjkIMamO
U7kXdaAZtNe506ogze2VvX7AP3+oMu1QE4vK++JtR7jOoNnFuNH1YeU8xeat26OfUm/ZvwzIwy82
Z6CM/9/NLHaJBh8W/LuBi05utoI5mUeZ+xmjs7AETv0AEZIAOn+XifugSd9xa+ppDp6MGUfJsFRK
kqI50bk3gI6glObKW4IM5X7iReSA7rHlaxOvLb5NT5dxB73yfYuQTMsT0LvYgCkUcqRAGw6WBUPu
pwy7vfe1yKYh4fCyWJuCFsGzNruyVC4guzz57qDgnBt8KT2oDj1F6XxrzvJHZYaViBuen4KAnBwQ
r9orAUnSPbkVUGROzuJm3H+Ha7S31Av/T5ZC1TbcTXfgIbJAp8KOM1Z8r1lGt7o3JQ9QhmKT1gdS
eNrnrNQqnyX2rZ4nstx4EEPWsnzOekIAMK/XY9tD6CprZqZdzzYmEClCSxxqTZlBH8h2A4I+Ft01
dr3Dt/WIQ/aH85uoyf9bklXtRK8N7iSoZVCnxZcpSJAE/rv8tT6YoMz+bcr6laHJ2hfR5cUtSrIv
GeDbTNBt0GnABcoZhNHRlD7QkcQEvxLT5E6FYWCzQnvZ+9xoj8UHE8fJ1xUK7G/c7aiDyg21C0Wx
cq4BDiRAR4A+ny/8ak/MJiRJLGz9KY1V0bWp9iQ3F+9/nwaTQIkXCN5gkK5LXO8uUoH557ekACmo
jeRTUkz9g0hrUGGX7k7KHmOtb0bgYUkyxLB4VTTxI7ll3Pj518c8/4PvAzv8xhZ84ATLoWM2Vt/Q
A4/7L7pAINK+tAZ6gadBPJyJZRNZEdQ9K1Sl5ZKfZHxn5rTBzUaj7T9UP+FYmq6e3G+eDNqeoL/f
XqwLKfiu9eo9s/QPfIP4juvgc1HxroMkv4ix/7HL9yhEHTkvChMkjlsUL6v5TuwKor8wglT4eifC
CLXfV30uMq1O7kLc6WOY+5a8Lz/jSDWjKJ3nXe9+TJ7f9HH4VXpdxiQyy/ji+IIWrCKSs/rRCNm6
9gFz72g1+dWk1W1iaNOBmi9Wi66UYNLbMTc7CBh5ALlToaWk6HpajJRHPiYJ1nv+nAAQf/Bnu4fX
Nmm4zPz1EWa4FvPanpj5bkArnCNoC+q59ygVXquNvlPbh50aqD3uwVGQcY06zaT4VKtxg0JG5p3v
ozY6/BA5KA7/rXyc4QV27mBG9kECFtC8Xb7USlR0EFq9pvS2nLuHTc7EPc2+M6tRg8E/+IfJV9ix
Pa0ezUbZU8vQTdB2p8bOErWnF9LGZCRE45zTgfMOuMbo91eMpZUjfktb0eT/RuYe+F8nM3UNKxdc
WSXW5RsGZ/hjARFfKl/hO2xnsRsr2tZMAQtM/Zq5z8mVtp40rdT9hhVzZEEASfm6rr10EVbH8LzO
Vnrl+xGFLMGwlpKwGOILbINKkoxmzGbWeTJUAVo7ZSRC2yLQXrlz+cYpfP4Ny77MCnZfvZq+o5f/
K0TO8dI4y0vqr3ACf5VDmoTF24eLgNwi5xq+C5Xh9CzV5Y3Q82yhFA8wzjHcqEo0/qPCRkyAB0/e
two9YZMqYlStoRXsqUcF3cX0dTtZXti2ScWXhJCjOHOnK2eCwPF6/Sk+ZZJeYEJnzB7BQ8xtzBTO
adIHOuyZtSnSZSmfWPVFIfHUAoD6BVnLGmXvM1vYznokl7ciX/3LogczKRjDCjD9DPiZU5u1rcpf
/85NiY5bisEri+MI65//T9GD5Zhb5OH1DE94ODBHf5CFvHIWBUcHOjPGUXhqDfcPPvZQtQ4VqyMp
Q3umbEhlKJYyHd3sWF9QKV9H5a0V0U974nsJs5hcpe1DxrJmjpGL9TFUqqw4LVuH2tq/EH4FMZKG
06pSh2fqpbvhGPesPNAByDo1zgvF4rvXpxc4KHCwnRo6/j34zbdsCl6Mnuo7tlJfVoy9hvLeXsBe
VAy3xdUcRYZf17fn5esMP26f48G2jt4om5xiqkM0EAfIEgfVXTYdzJ2m6qDBhgEuaDo3Js7/RbA6
LwNJUwRFOcuAb75vcGs1QxRFI8N+3wAf+qgosQ1sVB6F3Cl73tiCEQ0DtPgqLqGTHkhsyrrEx5FX
syCi0C7RMPo+U7+Mg0lF3AEgcEYR+XmhOTuE/t0LoyrNPJkux+T1KneGQPMqsNbarJt3ujlRP/u7
KRm89FakmufuoiINEjxRCVw30HnL4oNnN79rrkBu5x2UTcNS4sYB4cXsYkZIGId6DN42RVsHhwjl
/HSMcSbTJWTdzP8rPeZXQItdtVbA0lD9dBhtX9dhY9Z+2rck+Zrjh9unOm16w17V/VYgoTG5yNRj
hG8+4+XAzi7MAIVgngiSvBLY1R2Rc4b0k0sCpnGpdeKew5sXz5/mFsDDiq1Jv2tJQVTqI0336x2G
QB/gS2etNQiAIQaKX7tUCRveKcb7f/jQamRlar/kU7r5UGeaqhvF6nRXWV3abST0arxS7v7su2qF
YtY/ESWAJ0hdnch65aGRkXlkJ+9JkrbYjuf1xRlSAJJT/Nd1lKRZNGj+bhRFT2/lf64CiYz/5uYS
DJD2gAcXtgAIysctaWRY9ewOILvyvq4HnFYUIiRozMDlnIYufdEOnf8/O++Qf9wbtfA4hjIcffJm
jsot8KA1yoGR5KSLwOWbDufTXgTHW1Oi0IMiK8Ln+SeoFtDVZyAhCrISZKAIxi1XA1hSWBXGuMMQ
W4Lbe2LXx9vdWkarIgfw6923GjQ3/LSWM5oD83C6XSsz6hpuQWQ9uuypt+U93PXewdLp+rnNnchw
Q4OCTshgGNoVmdqUIXM6XLu9NsF+VempGo9QooxcLTthGIb1stcau6sBwaH/a8UBcDx6AQbLV4z9
qy+0JNfRmojaiUZny6Snt6fxuz3RCC3G8qCabUxNoXPFezlCo6kfW6Hhzv0IsDvUweZ2srWg2vZP
hn58bnDvP+sRF+Ff7d05phv0F0UqdTV1PjBDJ4EnPl7yuakIr5un5IuAT/WT+AMSDvrxzKihnVxd
NAN6x9HpXMg4z3zmM3fSF1Q9Puzb4vWQKUctUtQ3buTScbup9LwDV3UgrX+3FUeREXrWjlvDOzT4
VCxFRArU9QGCPOf05/tNwCnqw7IagdCGSRbwy5tZhwU07AK8Y7i9xVWdis0zm4LpFqCPCExtoeNe
jHI6d8DCx2VFpAfz9KPXPDd0cPgrqlgPcPV9SY1eWwQZ3DxR1TylobFeGcdZIgorTKidpypKWi8a
rKuSFEkzmqZwinhClxskAk6M/JjYYyO95IAiDp5TwLpcGOTkIXrkDW1I15XnJWI9nEMxTdejprPG
i42Ek5kyVqlvDXSw2capC2nshgWGTPbL4k16ISIcTwzjl7GHorePIwQ9tlxcteTJPOXWR7OGVbkw
Kz8Pq6UecKGUPEXuGRYXdBfRk5WxXU/9oQfU+iQAl4tgrxYtCYGw++Ile/qGrATIzaNKqle2mahi
xl+vxWXKijMWtJiQd4yaAfm+M9jVIffyz1pPkNcm7ZYyHy7XOLyfwKQUykVwNJ6WBYCE7wC3u3su
frEkPwWlQ52baRCXiSOkslsVBCV9Ly+Hr2nndkbOifJfnVfwcS0OFpa636f1qJU5r4zyg1QSl6Ca
2dA0gHB2gkQZ8x1HfImSPGBqlCpz+cUbQf4qnEy5Mna1aeKKHpxPl0gAew0X7+OhqAbK3vLLN3hm
1IfNpp6fVFXWCueSGd4SyltS1wfA41hH2qf5UAI2AsvLPlEDXTiDUyxY6h8XF1LiSsZ7jE6TTpWc
9BsL9aaVMyKohexYWukpQfJFLo4A1gGTw4F7kAtNQnI6AwSTQuaupy+dGEdshdlDAQRy//oXZB1X
aABk0nrgx1KY0qSXw3r9N/DdTRr0xZDoGdCq6widsqANimvF8GUm7bk+X6gUFexwMBFfUb3S5/zN
q97Tw+YOtno8oYaCg8ZMJXhuZps07dpvgn8Dn9eQrKjiUeXnIHd5+GdWgJyNdpzpdVo7+jQbMzM2
VMSatD33+UmYGccbksqAGxo9kwFl3KcpeJ5Vo/gKGrYUchuADyCkAv70NZe58qjY0RQIEAs99D5q
/rYdYZM2wWvE9Z/79O4lHxjGpz4VuVp46Ufl9hUrHvx4Yiy7X79UfqSsrZvNaFTRbFdKZdfPYbgS
DWr5YdyI+cq4A/gNsV4Tx7ldjmG6Wu1tG9Rm0rA6asonpAnQSPrVdkOsgiSs8IKcbmFwHxvhqgGr
FR36FPQP5p/VI+nqL4XYX55Cpv1fPsmszG8/aqJ5Zoe8ohrlTxrxhOoC0Dbj8I1Rd4RjIXXH6ncv
LPvIP//C+fxaF620opkjgjwzYp+S5luZVRhMhGrrl1dO6jsFuHDPGmKcMHZ+y7AW8VQck7h+0JHX
Zr3/C16cXrYVLOIRZa7KXbR9hUFaVAuhzkbHKIDauJlX8aPVVyvBpEmXu2C2DmlEEjGTDN9PhMYd
qcPEna2yad1GkDplLb8C2+b/DtZG2aJ17806A2Y/f1v0ESzM+8yUy6IBeBhUOn5lxdqaJhYvZq+3
USt/gxx7W0R7gPyxukOzc4kkCqzrZTV24bH7lpEesFHC6MMm5xItGCiRmV2WY82alGSIuwiTRTkj
VSFi2xZNVdmhAf+2ehJc85qAwCifzT1Su1398brCN36Ov9U7tPmMenIXXW7ujwxcQeROgO9WlX8S
4N6bWQLwyf7Mp46R+62lgehEXAwEuHvBlU0gWmLP7f5pMounSZk81btqY5vS8GmiombuK2ftrKQz
mQ6I55wj3TNT8B8IActCBUZpAJD51rzrSpMAyqngc9N3CE8DafHxCOi9xQtWUUX/pYedsY7I+V43
hvCiOTayBpB/leTq/vUHM3ruk+TrOosQ/KjWSB1XkLMUL/6X7FOcYks06UYAcFwICmUYS95O1F9b
5NfNsP9CmTUmCMWoVVuhl7vF5XrxV9hxlNve+9vGaidSKWVcr5OnEOZNVUvOL3lVhHcxSQiSKjXP
J6dkLLTW2E6ACicolr1Z9o0S4SjUZ8yzGBA2RSmSIl0b5CKXLz2Aaw4h/7TKfmOjv/GJCzlATCmD
Cn2Y3HxYJG+2VOvPAgfX9fkNzUbvzqtB2Lcu7EsFe3UrA3ZTSANOqd6RVdTX/YExt1TvuOlPwMcF
L3dAh56IV2kEamf8AUsm6nKA5/Ev54adUChwIodbme2i9FuHbk97rM2AxtKihFTHtZmUrf7tj/pF
I8jJa0C+5uiIzDn42pCEuS3tLg1yHJaSRQeNWC051+xmkyNf6G9LsRGWQWWphyg1MTEyns2mUYlN
9+WQ8yrGjaTBH1H0uJ+I/M5DVWdvkeewSrXYM3Yf03SzqKl85JlMjUeBuJ8Rl97fcPJsZFOUUHKp
UzmC3Izp5pzn9WvUNADzHpN4BkjFERr/iz0GAZnSLXx1js6VSjMc1xMQEjbqg5zOmCNXPMYfAX27
6QCNeVKJQndZjg0Hp10rnNpF/FyfkUpDwMNVwqCYMmBpcFbsMn46JXEKuXTxNNJGtEXSPp1dWRir
7PO4oDxUlHWiFFGVZDodP12cTk9UlRCi+GnqMyKvTJfD4wvKP/27qPTy01HjTCVWM/iT1WWbX6RS
UPGEpiHTnLCKs1i2rcL6ZLUQOSr55A9lFr0ksVC7JU+1LpeoW1E1BWZw3ukPeEWZLzgwVi2ir852
sAotB7NN0es9zejdG5QQaDxdTP2T2O9mxIZl4Ql0gAdIteb6tz1+FUeCr4PsgBQqkUQkdgWF9EFW
yPmihk2qmQozowFabsOIM6AnSZkYATpYw8YE7dPH1TH9QJUUGEb9fkS7bWHeZOwbrV0fPWMdelEj
WZ/hCFIi3oDRLJA8knGf+zi+ufqGzme9UPwOgtdxrVDLAelk9p0FqZ+qzCjs6Ci4ayZU1+/vrO//
jB6KWFFKRUbp+sYdloNOslpr2IqEjZNyH+qd29U3TpW8BbWhNbn6cc7BRWbVH3SFfNVnLxwAlXV4
mzf+5bCy4/5h4FKHWkWenqxJ89M7DFhax+Mt8MX6uqFDflFVtTpbqmZnyMA3waxAKq0SDfKftizj
UhZIpiHC4vlLb/MArZuTZYK6t9lQEqP7a2xjyQTbWSAmxbPT1Z6o3CNeiA53DmOBg/jMu52+UUY5
hMc7BRxSx2A/RmGBKGhPlXY1WdqhLpnuRlRg8qKAwqBc9+4a023Ex/56lxb7z5BPIEOJvdy5/hUv
dMeLCiLAec7dK5Ujcvm0mDVd3GoBPKo7HHxaM7VEM+KGsf3SUT60oY0YZoCsgEhuQ7vmyWesm2yk
MVv9UjBoFbybXpGB7yaCTEQQglujYLn/YzkW5gcjsDiv3m5A/KLvQp/qUDSbyqXTD5/lK9/DfNkN
PoETO+vNzZR0wjM2tTRcT/KHYFNhCUu8OgsuReiBekAAA229xQtZvG7+Ovt0Vq1HkdK+F0h3O9E0
ekLp/byfHd+upjq639Kkyiz3AsHwd4hGFrDqEwOeBwfiOiLw7wOx2liEsPLngYMOmSA+/BBzOYkj
Ga1i9yz7LJJRCyBmMPvCI4QI5Bq/wUHgCUmeAEsKTwC4+x6y8Kr/Xg14rjBVW2MWf5imStsjJ0UG
GnvoaLCFicn61HW67wAZqlgs77vig5/SMsqWOKRjA+VnXZ46dLbzPi+o8nQX6BuHI59ZLPOrUROj
eJf7B5vxA8Zr8fIGJuqLMuPxvAmNCIExfwnecB4l0g3vcuV8Hs1pUxOFjgT7ISGBtnticj4+vEAO
GDVkoj2dtRsAhKhEqwAEQqfjstgs/gDgIYgarQhGMteAjOZdKfK8ZRUhMT6ADo7fr0G2QJMLhNFq
O0bkIE0xYODBtIPyNAeqiQBmIZbO63/w6e2Aa2+PkUMfYM9/PM4xBxr6NQ5Tfbm37iKbbqkI2/il
WxjALM5xI65n1JKmLJx9CruUJzFdPTQrxzMSEDH03sj5GvNxS6a92i3chA0I+7yPxVcCej4ppwDt
SQIqxWE/Lqo67fnpfOt6OYUVKRJrANwauKbm0v20Y1UwdoeeK1oEPpGnH4mxPf1wG9EkFh4NHOCH
t5GaJwIOioA/vFmZFAjfcWMPvxf/Czqr3lT8bXV6QP1LwlHRFV/bZts6JdCQeUUejMEwJrSDZnp0
F4scqctKg9/BCndrkoGbm7xMGbHh5hVMmjCZLF9DvAXlbGp3RBBSJnOHlnACwjW/SavU7G+ol7Tc
K/l79EeVQTnglgdI1kE6lB0nxHghlmtJHdk1zA7Etl/ZbuPge8J7EuWBygqLmzGdDlzbJHS7WKBx
/kMNPdhX/FipDUeDeTQliONRXtOSL8xs+S8TZUM2fIFmcVKM6IumM43zRNpS9Z0CMt8L1S6CKyw0
be4OD9/Y5HccsoiLqRym/PhPEwUyuv9t/QrtSTqjvLHT21eComoMSq+Df4HihuIOHGYGhH/45ta/
IDnLnsAEpWO2iLkYrkbs+AsUdkKHcEvSSwiCeyffMleopg6uCfaci4ji5GoWq4X/1irepJRmzVVD
w+dBOdfTsvW/vsS6hjpZo7SgjkOXtZgvC0ItV0fESK+xPEMQzZDgcEnkJHQMgdogn/3ou/vNwMrV
BeHyxEZiPXWmkFdeJLypNB6ULwQ7ILqeynNd75K8jiZ6RbVurjO8hrRciN2jdBLZrxs47D7V5bkf
pv71CmFXXnQLpElOfbC6M90d6D5eyYgCQ5ZIMjYH9hvOFxTEMGVe+2Us3DBwntfHld62wsDALhXK
Bo8aq074rBdtX86jcEfPlG/ba0ZU84ErTJds5kMF8Nc0jdpHSv7eeFgrDgK7MIS3XAZxzdOwRDKU
rNjL7ezY2uNlYk4byco/D2aXjYME/8AlYHjAHcX/c0ketwrMvmumPjU7lm//vU6oHIu6Ua5f02zm
LBqhogvAM6r4x5SeXlPOJLVDnKgXnaxeMADnVN/GjKDa1JnDnmD93rD8//MDYAMQM2LPhq4iepo6
ReEcbPi8rokIUfZrVwUNZohhlWR9u84gul7JZOnZ7DGd83V8nAdE6Lb1x/hoaJEr5bbMcHJ9uulO
reV5nyjEQkv5JmyH8+weFKmqRTCeQKVqCXRTc4+FltsWiUxdbR3FeTXzT/6fIWl5G1NvxeyNAZ06
xHj7/Nxsv+RFRFhXE8eq9fZ3iLH0RHhlUqWZDt1zIQVUa8Mt0ZmuF29Gb9qZyCbtAHH2WIiI/P8k
1qZ24kaUGSNe6UNzXl2sdmYqEo3YQHMURqoBry+S3WAis2ScWP2ImPrHOmGoYi0AgFRY7dBW/bFa
GlaVgPdEAnF/RPEJzZfP9hBm9Ycmba1a8eNKnn3uK6iJZgA+Sz7kKgi6urmBvBISv3KkrKuZZS9N
mOwDC2h9QpvZzpgGCr361BHYQ9RPkkj6EQlI4FWGQrJma+BC/74f1ChZRdmUnJkoSnjorzePBZ5D
SnZ1i0sVwez4JSzvGsvZoMLsEukiJeWtPmnz5CGHyEQiwetzF6y0ZBo4cHwWRhgwhtgiSxF0Cdyx
qJOjzl3TNupVvgEinAbQn44Y4U0qUXe2NFgmhlBpfz9r6QboIVqtv+0PCMDLCZht6ksrBHzLqkYi
Jd+gZrnvYAgI4bzdWyANxRSpH2j23eABRUZNP46pVHI+O72GaVlec9+r4e3USXUhXfp1St/UllNs
bh4ASz5DptGLC49DJiZeE0TbXk/bewZsRFGY+arUUuFqhxvoBWvDhQ6vsGyRxC0AbTjmokXEOLid
LXTxuNyvXNAMCGpEoMa+Ykdh3o1uHu+gnLvHFXwdD7jf3aKLR9F7lpckRuof1mK91ssIjHZoJNkb
eteLBu3PObjwaXfnG6TUmNFeoJwNQnfCHq59XPhOzOjFsVmU/0PJ5P77XIDNtpguE7MMIl1ywZjI
gkPWXyY9eV1V9pnnTI5TWldJ9bFj9V/NgOglz3P343sSjFJMdrGCA5YhaWzJEPgko6/0hvXO4zIG
IFWqP9Q9OIXYrcWRbeRsk+zlRzILeACiw8yGpVskzsjFyWBCqrwXit0OxEH6lF4epWkFxCugFojE
IcG5eWUJDXjiLYo9PzUjATf91GaPQaGohdRjOZefyqZEwXjVrVbvdLCiFBEbWx8lMxW3B/HSO4ir
qTuq9y48A7OcklAJNZ8xE0sZi5gQ+vWcbp1gyHTjZLX/qDz3US5L+rET+XosXmuesfHuAkZpqnrc
iUN1tasjnYOsCSfG5UnQ8JaPAJLcnPNbAkVpqGlmcAvRFb/CA5uTlCRbhV8UiVDMnrpVlHkvlPoe
U4L9/LY5KYUO3P9dYHCNbdrkodFbAAhIBQqO5EynPwQKuyD351VRmE7m2Sqd++Eb7P1lscP6yBag
HqSqLHwDPSuyl/IGPDs5LaD/lqCnYIGIdpm6D1CtpQAzebVQCfy9L3qFpAboiJ+a2+RCthV2toAJ
WWUNGY6buOKrbA/Le2RvibRqwpbRyv1FUx89V6TGB6yRUDhqLEtwTP4/M/KfbhhTM7y2FAg9Kxin
yrsKU25ckJBUCCuiAgJlM+cx6DoOzbZlG1ddwVNIRc1ffrdG5rexES4oCMeOWf/m53VhAYi4gAXx
7x4Op/NM/JsLInFHrMUMHfDl6Hzm1mTnSSuOQV+f9SKj+nuKog+G0Y3AN9gyW918LDM0EIpck/r2
eZEvU3zH0B2EsOGlKCLUpaXG1jyhEiKBJr9x7uuT9m1YrbZeL5dSeyQ5mVtchARnCp2yM8S83Cd/
/flTieySBwHRat4dIPccEsAGLKQqjFXaKRHM3QjazPWABs81/+lEEnwIJbJGqampqzBlz1JV+Po2
evkdGRSk425t9BKonCKbLWdZMevenQzG+DMLp6JsaEmqdNWovN+Iqjpt61bdlB6UV3E0OIWfa13s
kk9iaqNys3Q0H58kGGe9C0zO4/mSnsRf2+ps1tBRa0v3LO237TDWa0N8qQjAqMCbNPaE5EML9ZAm
gM2JyDG+xMSTEm2NnkFQcICeNTtnkCtBVYS3R/8YJIZEwn7PxOHdbepB/16JGOJh+Cd3f+//cSIe
SVjyIcng0ejUQmrnHGz0twIu6Z8doqkuBtdlWECX9UV3W8923gGvVy5J17yGX9Bq/ldQWuIvQjdA
CXAPnqULh9qOw3/86J03THXpfiyvl3l/tzD7E/ldt9R5iYh/ib2bLkl4ux/c516aS5F6h5Osv9fd
rvsfkHqSOvX+rw7tKfmf0WNFCD8e/G9hISZ0saHoGRK3L+qSgKS8hpOhyQFM9GRhAobVqlL6p5VV
SOlwzA7aisk4bGYyOyvty2l27P24zySDz1LjEi3J3T+wTMO3HT5Qb5YqOEbG0qwezBME62Msb+Sc
hUs1oFGAX893e9/SjKxF6nuCNbsFNJKRkcZDoFTao/MQeIAPH6IQ+uT6Or+0jkqWMMUSTbzMcaiv
mr83SnxsvmMqk8ABcPlG8QTXGYD9dBJ91tXx5mY9R0XV0vcvgyI+W+33Xi/bw8LJXX1yR6XgAcbs
AicEw2faH/0tf7ZN+SD2ZUeoqdNnN/V52Gx7xiSt4GOlxn/TBAyMv9+YbYAGNSu8icaBhXNNK0+C
nYvxJO0fuxIpyXei+W42UXtu9knLWUn6fKQ9o0XnsZsdMUe3aX2f+Ctr22O64fkT1NNyiSv7q4u0
y+SIuS5IeVOPd7R6k+wYTp27PaWDIJ6JcR8a2QbTd+tV4rF2uqr+RE+Cd3Zn52HyLuKS7iv3FEeQ
ClBUO3zY+MQ4SpkfePFWSTSTS1ikwbfKpqeohL0Yv4/Ef1oWSVDWyEX0KGtzgceqD0ecqADUxi6c
8fNNEbw1U7vZCiws7jlKO4Sryvr/KPN4o1VSopdknGLmNc1lWyr7EYjT4YN/m4kQ/Wkx8/LBj7H1
jOeGRrDDPRUSkZaloSk8vMU+Re7DjZT/gyl5I14290MVjBFng5r9cz+bqe6T3vIZHOonfNyByUJg
k2bONg+WsmU1UdIy+i4oRQLHR7GYqcgViu6cmo3O8v5/TfS1z+/m7KAbI7hXmIKdUfEH+s3QKuBo
VOT3ySXG/5GpHVAI2+fGgluksl38SO0ZUbhtBgqq5dU14cFNHuC4lR2v3YSfhhjk+vfbGszQ0lta
12u0WoRLO3mpIhnhj6tIooAcpLfQq7Xynrsfr5hThAE27qO0bJ7pHAtrVokiZEreuipMPu26w5Lu
5B0NwyB4kQiiMe9fwsaqqyMl1+d6CJr/lPhGU4MdL8mL5m7khMI50gN15aK3yHJZqfxyT8CnJtFY
2f5oaDFfrQ1a+V10lVE6MZnizIoRlIWJpS/JGCFl9gvuFTL145CPqlGpEBz6kyVPGmb5Zh2IBfCS
UlvWfAQ8L7qvOp4uboHfgnL5bmmbuWOeWzwt1IfMlK4nwM5kysWz7ljiPRVY7IY4F/F6dNc7pRYq
HASaAk3fF/ykfBVXzH+mpgie9Vf27mM+ajDLu4XvdHv0lZuEVVzoY8CM1fcOGtLvrcJlqT1GtDfx
gFs4OLtb9N7meKo8E6BQqg1/rro3k2QJqvxdvUDy2McYJtLVd0DiRexyuudHDkW0QwHfxjA01gd9
FkzUuoNZreyqA+eRzk27ve0SifWt4pHs1vvvXHxvROGG6pR0xAYLjpq7Wat6VdGWX+TqazE0K94q
qLofrrz9NU9Yi3uX4fxJcniGs1/iNOG6hOcf+3DatchHTFAV0k0qFOw205e30mYLFQMpaX1c1gAv
WlBPzKL0n25WdBR7i9mVpsOs5pbh1FFMmHFD21qvPg2EOFYL5nugGw95VPnKGQTr9gqJM/56Lwmh
wB6eta5YuAwkAi6TmcIYwa7leeSDAgbbmerwP7SsxspiAR3WWUm+CuSiHb82aBXpjEegPsrG7E7V
qhDueS7zTDBRollvuwWRM5T9itmjpt86urwvIMPG37QTbk046Nwr0KPHDMtDU4KS9LxTL0NpwLJT
rdX+gWKxxJ6n/nma9V8Zf27/zG9UwLWOGgoi5tpi4I2QvB2zUp/hnGLGGkCT3J85KuVN/Wd30gGJ
obbF+KOPalxMYYZZDcdpJDvzeTAhTzu0U8S5ENcBAisvC5Jqjt3XKE7KKwK67kC3X49Vch49fQB/
dV/3ULUXfVgf7S/YqvbTGKoDkbprqJJNlDOtxi2BygPaBMHHzfOETRvBdHwI5mS5slTs4pz5UIeL
laqi34bvxILhZme24bBwXqULit87gJ7BySBvdKWydfqdUJjNgOiTnXleeqOLzjXJ2Sh/jlPfffmR
jxWczahyoKktNOT4h0ioJCrHHHJxJaFuFdPt4ejyXXRUpuaCCkjmlyUOt9aKYYoeJGYRhzKWd5TM
QcADBDw1cDUn8Y8/p/ebIIlc+fPr16m9RWwH5KzOMX9SjjRV277a9Wck5iyqgn2iZOmCQZAckwnz
A0d+4G2NvxgfWstuaju7AKWMn437fs0wCswbkkMbJQgdJC+tu9vA6sO6YqPaIhxS9zdJ/aVGpXC2
LLYrjO6vC1an0LAcTeZKCl21QXUpuJ0nxZpC5mzuBamulnAAvklHz20tfGeqnG/XgKJ6s/Zxy0+v
wiDTHpghMB2uOcnFDWO3e5Nw1CzJW6pvBpxEr8jlHdpdUTYUw+ZfmPSZSk71yJv+3QMi/U5eJa9n
J92hdiHHABlEtVn+VG/YkaLqzzaDO7DkDNaw1+xf6Fy6oj6BXUzAN1KhTOsa9ql2yKpeKtd3hsTi
IgTUB4TpGLqbJH/H32x9JaIwXvU5LJFEqaVljShsqvdd2r1aLuNyY7reD2hAdT/QvA1583G53GzM
DgQsWGCCOy8MYZT1A0mzvT1Lr6QrsFZOCpBwR+rZzipbMvGk7fmjsLkegiC5c62a01r6dmnMPOrI
po8OsReirpiQaKSyrupyY3jAK/QR+yw9rpC9LttaK5pH1bD5tDQ4WN7KXk38zMv6Nn3XliCNkQ5S
aOJS4fgzrRFY+25xO81aZrKm8gE33kOi2Q8q3UBxfI16DPyu3ZsHsAZ5ex/nyuWPs3sJxCFSJ7QK
mSGpErgJZV2Gx6B/BCrOi83Qd9puZyIh33JMDVCSIgW2PbwZp0HYS5Jqyd81o2P7Igh0ZEWLMy3/
1OXXZ5X8waRYOSpR+iRZfoM3ECgLiPZc7YH7E4hzWC+Cbk+6M/oSeptSuzhkK6KDwgG655M6pC26
XMll/fCK5hmLE2gErdem2gQeS4vA2coOsI/SRYuZ9ZK5HAp5c5eXtVwabOqsv0CJkxTdcdQELSJx
Y+CVOpnImDHI8NO0f3KaeDqnmgzbF5KClvWaPmmIls8cxTL+dHuBDY6PSRQdQlFOQeQTl/7tTRc2
XNZ4QT9wTvSaadtqmsBfIVQ3rOZRgvxIaLs67fuDY9RZFXjYrBX5xDFfhoXqViCWLQYwqT7buMkg
YHoEl3R2QZHa6rxGA+eW1vgZxSgThzHNYLrcpf87pFnIFl6EpmZYKXBNkAsp3wwyCuxQ1OnDdlR5
R4Syf/DjyC4aTln3FyZxfLBLCvXEd/Q4GUaZtfl4kYQUXNHlk25EfPfwCKMEWcQD85DMkRC0P9gq
dJxCW+J027Z2/tIgdPfJJaUSeyaQN2gn3yilqLA+2nW8jrZ+QyrGVtFVPFWcb6QVjzeyKNRMx3QZ
+oy5uKWjunbf6FJxgkZeigx9BuuBczImr9ZvMRUgGJV2N7yM68hbu5vhzEpDTzSBWS+aFGstHlBp
nb/fzMFd1OjGMlbImQ5Oo/Xp2VfdHsYFW1g7S6VPuENX5Fc3FSFK6j5Dg+oKP+kj0zeqneBel50P
qn28jJEeA8+EjN8KzbaAB2YpUdM4E1zvTVBM2ot7032dsPemuc1QdMnAYRbsGqHozobkPuepMV92
t1x53JPnH6b/L7mIeKFyZHpNIVvCTbG0TmLn1q9U2kDm44MLot5fwwvMJ+V94MrhgtVApHyNifuq
q4+PqXCP8dsx2eL6RvpRFpBZ+8/O9eS/PZLAVEijR4UxpEnJ2w6dQtoIN97ulYc9XFarRUsujTsG
PSuMU1yCUM7944g3jLWbvzSzgXfykJASsCdCb7acvpWbwHendo53E0+tYnC56PJIh0ioloWIraV9
v6M5wC+M+00/RVxbVWZQtq8f5HGSYV2KZ11lVjKoO39J2IsLUVbN7+cmcjGGm57WGWf6hjh3wbjC
iT/+mnMj5QmhCGxeRNvCrpQGwVGWR8pD46ILsn1rOqeY3j0UhsZj7AF8Za7HfhysIu7ZL3Q4mETF
Z8vxwYf7aiTZBjg6rChOJxmEPqCGVJr6dH0J4U2NYVCYfNZed8+E/LVjB117c9LIEc+btI7IZOnG
qJJThWgYGoJJtOfv7+4j1pU5vkZlKSFro2on7NHpBIKcvN8EAkIUCe2Sp9eWUBx2DSCwHhxdcfWk
u6FU2Jh+p6HBRnSSoichDtzWisF2np/YrY+e7RzgyksWBOrcxG1ECue+5smbczk2fOWGkpa89rKR
I+amh9b5LSnr2dHBDFFBQHllkklOL73HeLUos6J6yeSLuPd20R/OCKYpEYZRZhfWd/9dFiAg09yu
p5ociwRppRswVzCYXiLg6mkCVfl0FkJOxMlX5C9pDk7d11F4ihoZtaWtsOazryC/5FuQQUv5lyv3
4YcUkUgae4bTNWA08Qv4GOam2cZ6CU2LztAn1E7HPrkWjgvrYv8/vBGvLjeCcZyK7pLIEVSK/Vw6
eLxf4I/bsMqQ1M/bzu4uQEt1dJaXgCSzSrAEntQNA3JA6Kc/RKOJewch6GhCuDd/xcQHdz02WhPR
06u9miSC+L3PJY2tGA0kb/AZG+j3YseBd6/Fr0tkJ8v/FmpvHzpJB3vZwXF69PVCQ3UjLHsac34z
bFMfflJT29WfdxISg7PUHvDR0ppvOybG7dV9PRtcS0DfgF5M8jC5UWumK/1fBwKd7bvWQXWFz89Y
u8lB7svs91LyA9t44daLPjxfwGSDFowMfkxmz0hvjmJN3d/XoxthEm66atl2vjeTItW2tvsgSRpx
rPknvQfbTGiViNkZfeC0x2MYFB5IXfQNJymvn9hvMZWJDqGd8tAkuzZp3sAdR52rqWE2HkshFmgl
eLsZxugiuU2O3vxTBHoQuv1oUyB25Uw/vwIMXHgTUFGdxpnAtkAjnSnqCAEFAOREjpbp8NL3A0zI
jqvAyCWSn/tM8oYzNDcAwGKqfzetc2DNSrYjVX3WyIpo0nf+E/9uRtohnpi+16GuZVJp0uvJu7gf
HBsdoUHLTxJKQnQwS2cv7M2AsyaCy4iYSTobaxLxEWr3ZW3ShrCXwZQXzCrdVvvL/IZZakAxO+Py
qN7VLej9yb78tEVKjAR0+0opNw0l6B0kmBzEV6BoWpx6dm8sNnBGn0da+FwIv8w7Tnnn1XZZSKeL
zboUIfS3N1UAM3g1wqV72lTedBgc8sZnLm3sJYY+2DNLUs4BOqNTTS0Wz8qtdPm6/gz+ruOFOoHM
0ULyFcwjs2m57jxolBm3ksA5VN9oYyeOWHBrdFQCry3BjCf6BZWEFA3voHWboqwLb0CQ8PZrHXAR
z1xS6Nkh9FX6ZEAYPK7ZND+IWbiI7irjBOdpSwrK6b6tc+fh5ZS0s+6vl8gh3RXkTxfRRLmIIOpU
OlSg7icBEPcMYBgdQJL/rtAqpmW7TBEOajN7UBbhbxJCozgG5X+IDj5Y9InTsG8XOFnZHHPVLoMx
WD3XiljjAqQ/pjB7qYQd+9cd2d+NXZocF7sss2tVYWRis+MkMOtisyCHj8bHh59jqREqEYLK6vJC
5e9EKOX8RMgGPAsRQV3d2Wlm0cWkbToZs91f1r0vVTcYn3u/9xKxz4C8sd8IziMtgoj55jb4YQjL
45Ky4mFUDxMHK9klduQzOMQINniuPybk2dpr/eewBJdXZWwP68VgekdoHfY1ECS8whs+FqeKaxqj
qIL2LGQmYMJGuza3nhcZ4bGF6UF5fH4nugvwPyUnND3ToYqub3pGw0YH36uTQOpXODU5C7spFl5J
qhBvW7G/H7PzqKCxpAFOb3WRqcT7q9CeGKRoX0AHmgRm5QfHa4lkncsJgQ5W+eRVZFSz8MRJCMpd
sQ3/NSiiDs6uRbcdjkyzgjqwNrv9k7k+JOSgM3qLaPef32csutS50w6ApMaUJeAmvu4ViKW4V3DN
GKhphTIL6N1bH+hFg1GtVM5KBxBrycbPv7JSBWWJdDmGkNfVQyufKmflX/ZH2Mo/nrok+PLkEkMi
zSLWlOYPC0O1XbpRVGCUAMkBceeHh1V9FhDYFVfzudFVSujFljdoAiDr3+OzURWfsxkbLOGuzc/e
BDmtoHuInZ4jSQVc1olCbFD9yLaR5ZZDTiPoiKbTz5XSENAHeFrlOUe9kWuOKHY/8ouy0Yzl8AiT
zMqKaMFC/niuo2PDkMEmknueCkTQPU6v3XCuhPDepuA95PjgKpvVXK10p+9W37Po2qXlR9WoN5m4
fEcPJXqpSF3WiHxMNo5wAymqk+dCGiPKTnwRUj5jiNm8Y9AM8f2xGe/sk6/+bciJbvJdDREyrpgG
V/8Ntu9e9PEld6pS0mhzTT8GlBPD4pLTxNm0DWv2RzvDrKZlbhTfvF+IhVnKOTzRbEsBUz5wS4OU
qaTFebF0G6PvfYqZeEGQPh9EJ83vZwW5gSQ1vE/ooAAS7gUoIJ1QeVfL9FhRbC+ovb48VNwqAgZA
R+ZKPEUmSAGrdmo3NtJi2NDo16HGgeYIJ3Tz7IxugrPsCVODjdmPRW3iQUpQWgTnbnaZgY8KkHMB
f2wuPqjCi1T2Zjw2uvqkG3cylIT5j9/Lo/DcOyaopl/rs6qJ7qMoJFmHZOFvD6cljyLrnJOtlh+8
SRCYeOiyQmRQMvS2/0duRmNK+fMZTE2eIOqIfzihA4aij1Be6FJpOJbYtBIcy/m+EIfVnr5q6feD
EPuu+03gIYFu+6zYsPGW7gIw0ibLy3qIgvEICcIy6BxEEnbfTaY7R8PKeCHKxAgYVEvuX5Q3h2u+
zuyq5h09116DvjvX+Ri/J6MgSKHWo1jn9iika8lnWmEhpdsvdS6u1vqFEI3isG04cBKOvEJKgDDj
T3oOfI8EF8VDu2AGPFblC6SM+a0agakjWgRrDTPwmBS8okBX1JQnv/d98rUMk6Md1nK5iEt6H5Ce
8yHhxsfCy9idXBFEIsvOC6jKzwCsV7qvCoJVa4j8hash1Kyufmtx7Jdu0LzHfQoBovlmaLjtn91i
Yanvzt1G2+/1k/ErFWDN2L6sFuCu4qLP7FTB6+2HykT+3dYLqjI3QwQEsZgofYUOyNfm6FCOZrMv
X6MsuA3GYFgxpZnZu6Jty5jyZVrH1gHjUAfuawiNJtSAII1ZxAwIUslI/uW/5bqRFo0Lp8RI/JbP
noOPqO/eNQeY6kjfK6ROKlPCJ48fl/t6NWrT6lS2Itvv4q0Y+NNSgPMAObty0Tg7P6en84XhMYWF
be0sx8tCPveoZNFnYgfeJN8vXNyucQWxeOebR8Wbr6AM8JFnN2Jc/EpXmnQUiRJ3N3VxmRUsCXtu
JJaD9gH8K0S2TxeMV7IEEIRNddEUNQpD399/sPl61v3lE0ghOXdM7yDe2v8/sZiMLhiKNzjeWKH8
SpBduLFARBNNeUS4SDFUTXwRc3CDtz6wW1OhcJQGygvhqevngWHd5F2hfviHif/TjV8Yit3DYdOD
pJQDghMgbr/Jc18EzRBnO84bzp+YY/UdcxpZWj0wDEykFh3XmJPSFWPHt6AlQKW8vkO/y+yKzty8
JYKY09Ru1qGz0N4t/SBA8cF+LtI0CCndvUVu/VhkVe8koxkKi2Q1HsMgrqWL3ynLEk2JSZxxOZkL
8yfBYwk1PpyfU7qqWkvGWklFfsvJmoYpn48VDtUD4Jp0you/D/tBdxAZHqVqOUT3DBc61brSWmCx
tSlBIQKpxSPrUmJW5zQlxvLiKdsSuJ+5rvlmNbr75uXzPquqHOqzAixtiRHD4ixkiJeO9xAziOJH
ImpJ+ulXiPR6kYJsUDMPi3ffkhRU64rA3xAtHN15EMxUeDdW7BsIhq4EKCOwzT1dMpBMdU1DhQL4
x+SXs3RZ50v0ZjEo8jCFNk6XSrBjz4xsyWuw5iH2xikcGNS1eft+MhlyyrDPdtszmDUK/UEgUdSD
jvWaCh8hmH5VPdjEDgIS7VC3D29nh6TbjRwHeSkMZRTSzFuI1h3Th68B9+QSGc2OxhPDuLAj0UYS
Th1qsvJPqSGtdpp+CxKHa10Zpwqujh+RkLRKF3qAS91l8i4kpA462aquU3CG5h+uTNIt1Qm86ULZ
3snXkV7bt64EaHRuGKLT4Tz/K3Ek0ngIqBE9MvsehVWLL51D1LdBLnXiLox6ziT9DQMF7AMVB/K+
uM3IYXUC6jIB2+z5c+JC9cQRtq1M8A4YS939QJSgTXzCKqBU13CRrhk9tDD2vwk/AxFtBqc+l9l5
jkjWh3a2O6LJLJEgpzY5EUWptOKhNl+zM7QCi9vINofzHs6WtjxxkqJ0hTqEmzZdp5RZu7rgPT0F
SCXJggUeitd+IjrtYDw5IbD8LMmYsGm4IwpXjcQ9zcxM9j7YTYryzg4bjs5DYxTSjHwdt9cacc9J
EUe+D1LqBfVfeYFNoItBylDxAoj7JEqHb5yG+IP0+JRznnlK/zEwXe/EtovCz2Evv7A/4VVqarQS
ASWP1ZrG2WtKbIQRF9SU63cpKGYxG4W9QSH5qRx2prusb/7nL8VGh95ou7KjdDsd4fkZWOV6OpO4
dJguvptRWn019bScWESRIsb42kCka/fYzkpEPq9am1OdCFALweZp0UYv64v8r/3s1eoLC6glJ214
tU3bTnn3H2DfkYlvUD4l10IkYoKHOaI0mwM/iyGLmULWGgv9iIlL5GQ9163Sz9Aw76mFq78Xx9bk
6Ed88a+QQrKJlk+PPeH30wnGGLzTrZZkED0X7pJBuQ9O0Amc5LwQ8tmKmkhLgnVYsuECzf7IR0Uw
WCF3OWeDLrXyLlHl+vrKw/3lJQN6RKGv7a2XVcO0Uf+F5JJeia9Bc5tWg5OdzKxlvRgBRGL1sL9q
gTdvhUiQVMUsUhBfOFUhwohYHhIouCO9CFxe0mrJl1PN93v+eQLD0eTbCyU40HOXNE6pHQlaokQ0
1WYUPSpslNTzMmFViTVIBAo46GB/KxYtuIxLzH1ZzSQt/wQgYGRGvGyWHLDaFtObq6W5sQ7c44ek
2FB+FPP+HgSfL5HXwRbu6p+8MEPyxO6q8sKrDUildsBNwOZ1UIlatrW4OqzA90VfbXjHAZiR6FYe
Fw9z4tezBMzqNn64TbRN9jRA7ZZ8D7KJI3JFpmeAs0cVEgf6gdOPtjJqdsFHnjT4J9HICBsldXh3
0fk4f+Ubbc3oI0L90fGjQDeVpQqLqBKu5J2spW3mz/vbBJQgxiwupur8E0zh4DCVPBPnXLEqHXNr
3TDK0dStJc1pevPe1w0tAIrsRyYD+xYTDdlpm+TRtnj46EjwHAt2eLYZmKvS8fysgkt50Zp20eyB
a3/3uVV3PJT/LbSWFUqg7q92A40DL2qeiFr0+DK9r41UJzEAugrHHaHnkDsO++AgHb9dHp7YulEp
EDaFRaUZ0exPqljUvx8Rly6I/0rJznoOAugmU/OxgaOp0Za+chSudqrZWnreXyuw6qgjGJwiDJzo
SHsjDkumCC6rBtV93PeMAsgqpXPJpiHFMeDCWX+lvTAHKGQeNluNBAUhAP7hVM9uIb6s9FADjPIO
Yg/IEVcYVdSYBb5ojL2XQwRqAbnDROFtll7EjJyJpeQqudWt7z7SK+1fmhd3wKcUmBXouACJlFaF
3IaB271tgTILmG4aw85LAAsyZm2qcg2NsUU14FddJWPvB5OPyR5a8AknOsPI/I5iv8Wbm5q8K1so
LBcpiOx5HuN11hZTIFkQrB0bmu8FJvfsbyNeKvUytiec8oun4pi48d9cKKr/7SuwJoMpjy6fc6tG
lpnHEoXwlY55/cAZSSYOpweXyQJRcbnnl6G4p5jgvcYAWqWXJzXn/9C4k1+9iUWVQCrHzxU/kTzz
v7HjrBatEyJMynBOkMAOj6CSM/3pvy//lud2fqwl9Ai24iYMRP+AVZv5gu3nyhLRu5dfFgZtlkxR
MlqojESxT1zFg+JZ58sVh46bEbWi0yyOWmDuN7o1cD8T08kbsJfqmrNx9nEXekyKHVaGW/mVnt5w
0CR2qeAm7Eq3d35RaN3aJQ4cZjuMZccSh91rRUWo89wrYWVsenaxhriiGfxmDZD3Jj71aiECuwQd
oGFqycyofTYpL8YRYU2lI+o9AHKhH2/l5lepnreHLP9WLGdUnMADMDhOf6akw7RDtqg9f6VMMsw4
tJ2xJ++gbv7nfupXJBmYxPcqo2ZUTXK4AodpYIKWPWGP6kJeH0QisXJOQKYLCFvTn6tACRs8IPJR
e+MgVdRCUu2td7ZLPXcIKK1sz4mEs3dZsE/Zka3oWCP0fNTCv/E6ss6qB7U1WKg4MxWudMF+keC2
v8HIdafE5mvKeGQHVbgQOPsKVD0qVOrHztICa5sxSIG+kCYaFtnARf2rexa6bdCCIAv/VEYetzpH
IpJYkcjSwElZzqx8txuQg/zd05xufZS7LNrGELZMsOXzo20VvoG8omkh5sQ0alqafaLKqo8YgIZ5
9JNaNKdHttJverXt/6Vx8EXMgqtyqCW4gmMtih44sBaqVJ9IodmBa2apwlCtrBhZ9804SyQlP5tc
+zyt1GOKrvvFiMG1f9FUlbAsr5HGLTpRPPo9pu4B1Wb+AGOtTVN8FlddljmlAR/f/1hg8XP4snaP
gDb09tfYuBSEpk0FCjfZE5IxoF8K8rrOFjLIaLms34eVrXT+TsXlccJfhccu+fSdQnq568J65IJy
SE6nj2APT9/lZ6r4VWFaUEtl+Mk+vPbgO3nZAIrTo53+7I8H+NhmnGFwf0KXMJNWvLJK3UcHl2ri
1gOc1Zz00/0fHJw0gh4eD+4HEqSOhJy1mf9BVhQiGEfP+Vn4h1Buf/lP49Vrw5ZI55fVP7z/PTdI
xEEWzIX8IBs3GcyIVyC/azNUnvsrhQ4mSiJ+cOK/OFL0aAgSQ+E4gqmyoEFl2sqyA+W/YSy4YBhI
73p6ntIsmJaMoY+5io7F4dkxPfK9nJcEZ5JlVwuK750Wk8CjaChzKgHAvilYQRR2SVlEANslAhzT
d1q8Iz1nhrwANkODIssoUQtPfm7pkKvuRSJp1+LMBKqQnKuQj1OiLr3KSAzDAbCrpY2GdCtXPbkV
D2SEjJxA8A4bpB/avQ2iZ9Oz0IcNAO5vvWZyzDaPFISxnAjoA/52dtcw1kxEAgdAbr4Nw8DWGuTK
cvKT7V20JgpOKZkLMPRrY45wMVxTDsi1MxV0EvctH7iAKEck80Y/0nALKVahqu2KVoNbzyKi9/7L
sEQveMkiwTjEM/d8BCet7COW+BFHTbT0dMV+m6qjoQe62UhbdiHLhqb0XoqfH9r+ij8wC1f5nJSP
9SuW450cD3UJTvsYzo9oiHS5h/O/sWhsMBrW77o6AxM6PVm6m9zxd9+cCLeDGOTFtKP2h90SAZNm
Cq1NPFhfFZWR2/0u2OjRg2tG9y7Ho9vxjRa3jdiDxOAGCL+VEgV7RR3QjJXFP5oMyLEcgfYqUks5
Ju9Sf8E1zbmQyhhjYuh4UdvXosjnBINWUQRG/FMw7muo5L2ALNBhC0ssKsPWRs/soTyTLYyp1pzM
a0pFuckadjmRrg4Ssvg6MgOFWSyMoTCGR9hQDokfnk6jqrA0RXpUirI5ejMgGOjjcYXWN9ayFrgo
86dAaAoZiin44MFMqz06UwFTyo6ZE1J/DEkRuu6ZZsPnQXjG7o9DL/1/hwMI4NNCx7T0uAwc3nSK
Ud+OkFQByfeJBQDA5KmiswXFLWoEUuOFuh/R7NAdvwIg78zfPwP2vmUM5Rkl9usHvFZB0rSIEC9f
/cjq+LvVig22sigmUu3tPB+r+URRl/m9QFipIaGwkAktEKNXyp99snlJ/B434HtrF26ueVr5/M49
Nu5pumhZIih92MMxCPfbjiyfr4+p+u4BxcY3vujxEaUJx7H8Q7t1OxMJpEouQ7T7UDzf3xFgSxKb
racVOCWsCdRq+BnNmZNjkLwEA3DOWo1A0eirYU1MckST74AypgR0LVNgQYjk2N95eKUQR0nFf2Ka
ZiPjcJ5dxeshv870UBo3bBQnlDJ/3EeRMD9ckjWeD0snacvXGmIjR9oWOaVUu4na3ycLf006aJ9K
5ASCsRAGgir0u+5zBVC/Y0K/Rtk39yHFaYiZ8CsAvsNcS+r1+m/zZ3ltlll40Ifki+Tt/YGfYDp3
vwophQCOQ/Yds/j/B2y4YOnjMJIJdGIL5rwdFRqvkEVYCrFuPbF90qHez6DAaxTHJthfgl8Q51eJ
aEotUTUUnA+Tjg5MiASK7W7Mc9xePGYWUkLtXk1y4p6nfOp1DeIocFLzphrmpplHG6Wbyu6n8SiW
IPFlSH2b1+ZGqQeitybpmADYlZeLtuimu4yBuWElXl1GGzS+pS1v74uIPeRlbvb4QcLPPxnDFs7S
55oqM7Jw/fmkhTE+R74vycO/affAM/wWpn72TQrBmpNxnFBPGpR/U+GEt6juhCFqzm0LoSiFSBr1
e+kbnnKYfeuWPCxPtCfdlIeS9gomq1bY6AfNWtJIgsmqeO5cvzHg1FFGYWHOzcl9fEuk2Iot6NnS
W2h6zRdzGSWLCPtExhI8IBGgo2vJISiGwrbeNUPIFmutLFxwezltR+pDMdtHrBALZW80uQekIVhb
cOccw9XkXQQeOTfQhhRkTg88JGBHhyI3VGKueOAODVl9/3UBodZEeWmrIDZQr078efkvWVMpt3o/
o9UGiDS6U3otYL8hgblDOThgPAXEGrF4ZXFWYFScy2TWe/l8fkkuPMgbNP+HxeONk/rnIwsNWGh/
VySx87PUuTPeB7AIWM10mbisewfA5hOm7MLIOsy+dCyUdiJGLE5qBodXhXCZhNKdofNPViYa02Cu
gZiR93IzVOrVartjt5ZtE0+vpc3+Tch+p32JZjMa5N91QoJQrJScFUkmqb/jbls2joQN80GTJoIm
TY6KBa/n3rrVX02MM4ck0kkEukC6LgJV4m9zclhpDtQAoQjx5vqljjdRFZDZ5j6gTRCIZ+FhHwki
zdgA2KFJbAnhWlrYVOqZ7ODuuqKBN/Ku1yIMCTnNLclixkw1+yg2h+vbyXe0c1wLx8NUafmTZ9ty
z9odw4BdQclQqAf5exwli2iSJ/0GzQLd2E8OVZnBgzwQDzNhMOqWnfOHWhUhNgUC6OMpkz8C3+dF
qZOXPZd06lC1NZucGZgAogXt53V+s7I5WlwemoCWtJ4eE/d+Auu9bInuleFdaMhiFcVG6+s3FzZx
6VV2PhjEQiGTbUrQCD1Htr+5jN65E+BaSClk3wIBaU0FsvpjZt05U90RSK82i5jmIP6PAPVX982+
DJYwSroStxP1fttsLDidIC4PAP0gl980Vj4cQqm2nqto5WjSY7DNCv4Xmf0k7BD44C8djwztpHnn
XLKMOVgs3J0fL6ROKixVzPcFPHVDkEJJepcmawLnw4QaAtVRHx6AtBxXo7TiV3SzcBOIAn99SwT/
05l390/uKQO5/tk4h5A6Blri3+zTNUoONJp8emE9vlfDrZ7skj02CkeqyhR5Tf54VSIsf9o/Ke7d
ZbF0Io9ky6M7ZyJvBeRvloRMAe96Q28s47apywFX8FqkcCjP6eVsUOkNTSLuGt1vI1JYFin1Gmad
jMxrkPrOnxcKH97zRNVyQhcvav/oIgqtgZhzYkvVPzfMbeByI7qhhWEFwTUMkbtHE531GLCrNLMU
Q7c04xZW/J2yfQgWpbrYCqbi/gynnM5mMb87AfDyPglgDQH0NMwoLuKCzcbigtxwmDxWqbzZSSb9
oD4VD/6iEPRJ/GvT4EwABF+HRmIQgA0NLH8e7bb8ahPVYK9M50pWESF4uqu9nUV4RHOg139gv3rr
9vdcB8NWGqvoSkoA/8EQGBVnh5eugoO4alig6/72RHX6hyEPEcRfKOUHaGm38OKVR/hjCQ2fiFSt
KKKaTIUw9sD7MJWvRlbFkNxW9Zr10hjK9k48WdUrORmkwBFyAr4QrDOl5v/McdgzTVJgvtxR2R2g
CZikz1OTYze7N2ulnCPWWvm78nfNZmVt0bf1+l8BvJp7kYrEwSXIicfGYbHbcpcJEeh5xJYJ4P3F
p/DW5yEYejpOFZqv7VpID+ktM7IdIjeCb5xg2xxOxlcCHpwXUfW92ytafBHUaQC225q4CQkzrbbM
7SQb1WHx19r517TBz80tnh3+0cHqyn/pppgWcWUqD3YXMaXX2n8BjYfOu5NFBGFrSMRBQnCSPUh3
a/qNkSxbFBitSRHwoVDenxCN6+HvxLkMCylkR5l8a2JmTjrE2XBeIDe69+0ONumEW+4beFXx0hsK
iAETfQT7zKDeyx8Vv97ZKo+BD8tjYjWaIX40KEniZYF0/eB8GI0HWhggD0AV/+wABsdlgaj6OgiN
ZVwICPsML/SFhun5YrWXBBKWFrL8h+EwQMJF0L7e3WFf+aHleqlvwoW93qG1Lv7gmYIVzRbb+tUK
maSeeqkaJDbr+Vjy2ZP0qVCFFycBoKfXLBiV4LQ7Lyl7RVrVFjdC/0j776tXUr1Zmwj4H7TmOa+Q
kBXV2HaBbQo4Vv0YGsoSdy/S4+PpiqBHLCODpWqEg88/MW/G+S3pFBcFAdYIbnVZqtG8BbOBmxda
CHQTNwRpNXCYlNvE8LNUcoOEyy7x083gKwdegkxIEI+7UMGRm/ojg4+ffZD9T3YXe8RCG/ZaiFez
GEJc4kiYEdby72gIAQsNrKGiSYRMteyTFwgVe8SVGYGpiHTPPnGQ4f2dncxLaXXOyjqsai5nKWit
w9ulZLShXvm19I5TjOCedQx9fDLOGUM0aUZzv4VY/tgcF6aLv9NJIqPHjoD5ubRcBWLt/cftUJhP
5YAvCJQ2vACOjQAWN4QhTkAX6ChVIB/voZHjQ+t4VMZxR7bZPZlJiZZJFt9KSYTyP811SaOO0Bn0
YVzuXxU22LJYVSNL8+ADDOebvYgrSOJGDO2vEV96Lez9MKI7t2x1pBqAC6gY8ntGcz/eUKYqYbiv
jy6+lho6h+dw/rTYXlbnZnJnHvfUlZFrqE7c20RLzbIzGsv7ECoSgGbXwrAQklFGOuObIBvABZNj
x3bXPZmnqIaRzBiRdpzZGUkNbgU+H8+XzC9SMThIWWvO70pZLO/JCGUwyyG6/Xb7W2Rh4261qkjl
gKeJOYpaIk1mTi9HHpeOwGfHepf6Xdm/Ey2wtBiQo2lya/8V1gRM52/43iwsyuzDWIUL/MkPwzQl
0R4bgjqySnXrAlmrGfe+jqnwJBgCdkIQS+i2gOwnhVr6uM750gPCl+p+Cq4UhqJatHsIrwrhjzdO
uUr2QiIesURqCp2st3Tg4ow/SUY85SAeGYHnJvgzs4uXsaj3zZ49ZGXTenoVJCYy/Z43BffK1bxj
AGKQwJZdImM3sby4Yh3EFiyIeji0hRFgBWYuBhqsYqWWNc8VYUlbWvFKL64k4BewQskYTtryX2mP
Pf14G6rFZATMv6XDmytVlV+IqJ9mabhFWnKP8xPgutvdEjsdRnZb+4Q7L7dQjvSfZC0P1q2ncvN+
r3UsLv6ewSB2HGKxFe/0qwPrwEnuqWVrqvLSaBySBx8SedIqHI/XJgsNn7FWQn527DTR34ZeoU4T
Jyf9dlUTnvbRKM6S/vGZb1Lgj7fkVkxBnGNjrvBCumlTwoVxdZ+FS94kYKU+XMDDIgmOeZAkg8Jd
6y3GM4jSQ0rq0SULZMRkWzb/AssUY2lqV1ZIwe5UssvVzRaxL++MnSdbfWwdqDti75iUXo3jh2OH
pcsyan4vkFrfAmOCGQsRFy7cJpnsITl3XX3bZk4abk4N8iBLvtBXdS6OIOhbMIoftbVSUucnMFh7
Ni3DSsZGYPVcG7lfLtG+sNLklVJZwWkohwMb2fL0+F1+4clkOSnxWvzG4xnMkZryMpjJ+3rgsjSr
aTjj/oX5puQi2ZtQneh89weXpg1az5xCbaR21OMPtqhsZLvWwNcxF1GorSBiZ7R3Jdr7xkr2q+UG
NX1FNbAx9ADMoyGZZMqsy3hDz7ye2ihvILw5AYKmtUm1gCY75QmwuVmAhnWNAiJX4Z4aqd7FO79o
P0xsHAGBPDeNIFnLA7bZH2WTJAOR9uYRDER3xuxknheeEukSB0TUHz9kClx5nIvSbLR0Ss+6XtS+
kLaehZRyeGkC6WJTvXfxrAjDpT796aSLIYtKIcp+XQsClrsAucpdli8aDETPZA9fS6WwqQbmDIP2
WR6dY3nU+bgpUdoYCyOGWJG1XM6w5cvKm2AJhqHa7CZfs1H+x4hZdaFkylo9N034WlJ9N+J43ZJD
WUS9xsfrUEYjEUD3F2oeQynNM0phzRaF3kz5EiCZ/RoA3q2o15cNtINzQRYMdxCssHVjvmZWQLJG
nt6L90a4FOYHxdTcFWW6UXpu5BkZlG8qhjt4zlmnvZH+TUDQD9uX/puBGT2TWbFOBlyMpWdfKBGQ
ew/dsN2+3KNt/6J5Fh+yahhOu/zx0T/iVct3ZMqwig1MLv/qOMuGKGz6mE9n+h7BAvJ0GUcrwc7q
hrKP9KbqaItjDuO6X1ilCvrKd1EFqbGYNPkYApIp92gPVBnDsTgopWu89LUD74gg3QY68Frs3pYa
w0Q7g9UQ/4uIqhweL3qkEZvqockyPkDe2hxkajCypBiNnQ247BRWmoXR5YsdJ0BNKxXZgNeXly7+
/QInEbcnfzQEoM6uBPR9RZcEGc6msAjuUyhm38bQvaa9aLE5QbbhrffgGwvbz4FJibHctgklO1cT
YkVMTDm+lqhyPOJpyWSophXAVXXckYn2GocyuW2P7ip3Kwl/0hDaDo0EOPP7qkqngYEehIo1OHxK
2GKdsQOmC+SSQqCG8FFqrwNLnrtxRPZ+3xg+KtxY5DSF0PfqXIqCk4ul1DwO1BAJ7nATDz3g27ZF
jow/ECyi03pc6ubWvq0XoeE60J++ELw1B4RKfYibJPV4vc6OPlymER6uORxG3ev5+9SCdqEkU2Jo
kWD0W4ZapyEJILsDoir9VkbnlLGNYtmdCKtObP1XQ7U4+45XctGZD5eCaiOv7zFPEUXO3E0lNf8s
3AIFBCruzSdviXYBWWHOKozlkYYNk6CEG2Mn985SIinHdgAFaJkrmwhB77huX74QTZ4oqXidm24m
rGcphEDXV5X0xOKmE8ZBsNJL6fj7EXpixwRSlrfKt7G0G87rUJrF0pehxzGXprTOv00AqJfcMP+W
2Dj7CelZzqzw5PysXnDdfC4a+lu+Vgp+umMevxYaAP7mm8yrXNK4EANl+k1jugveXZm/kdg7b+yv
Lu9eE7KoIVXlRBTqFHIv2K3eCXzIPSXbqTCTZ8Vv4yxHom7T3nsrvvFOOWdUT7iw37CVvul6RXR5
+iUNgbDuANvzEdbtY1txcuYX07zJYVHE4UX8vQ/bGgyk3rhqL+0Y/MglIgqpoAjvY/8+unggpny/
wjzGYnHF2TM/HFO/XA3LNZb4aUjq/fP1sUfonzIvSCMoQbZFkhp5PjE1+JB5cV79Z3ONDBLRfBal
98XsXf+arFkDruuXDkBxTDhV4HI9XBabE4MiB5EFDP9AHFxbhbdLCmjOKUIE3vJc1fmQpoBl5nva
QO7uENBYNiT2AC7adyxKoSHrIAzv6+7rW/4uiB+74N93YLeqnxG/oA53sE+lcTwadUmtShFQJ6WN
ovyAHfR/7PZBj1DQrHYulg1kuc3GIszDeP/eWTcbtSV1R/wX3L71bLxO1Cierj/p8FnnJrsG8LQK
BKPLlHMM5Oitcq48DqsuZetlCmrtJdF+/BNsoxJD9AU5ATk/5HWVOt5eitknIGsR1q66Lm1p0gqa
QOupduYo+KPhe3NMMlXi+iS4zpn1S+M7sNZ+Veg8m9E7VlyKjD+fYpxN8tqbzGDirTbu6ynKApDE
L+I8xkMCynxawW4XtV2TIkJsYgO6/eJNSvL7rqFNlVpeqy1CIICU/ZECV0KlpN8YiTavlzO6HHwo
ru4kUByhDLJRBENMD0wM6Vma25l7gh38ONQ2wjimMgSy4Di/yNu2KZsH7VcM7U9Twp//JU6zJ6mU
bNWoFFYYMe1rYvxMdDzu4mOADiYZw4rQMCB0ssf16N76w9mAfw3/398DMHkBVsYRB/qphMmFW6pm
AURccuCP3/QBIM5t9pKP69LUwjicZ5b2xXZVOoEjkU2QfXhuB02DMLoxAKUBlo/7FxF6jfXsaalj
HvIypz+WFEgj9Xyw6V+68sBhCrqrxeAzoORmbqqANAuvRU7fIb4JjGLaGQCl/Y2C3NChxh1V/DCm
+1fqZGp3IySyAEbzhSBkwN3T0DRXlN8bnt1jKLa861bGhI1Qgc8mNEpKBJNIq1z2bmVEO8YoFMh9
bIbFm4+yk7PPsgnvLo29TED2zMB5Pv8/OoPxMe94Ld4MfsVm4MygmKZwG+Cd3a+3zfoeg/0e9Drw
s37rFep3H0vDqDmppgFT8g6w56TvqoXOM6ekFhH6r24SwC5T/BJW9DNuROdAZeGt40v+hmDL+x7F
GmB5phQoz7JgrnZWl1ISu8V80zUYteu9CgWu8UVq/5cgBVlrhelPzu6pWl2VDX+t6BuF0P/H3Q4X
gUpE5Fe+SKYM4YHS0zveCxvrYc8tJ0zFknS4CRf9bE7KIGnH2kvpsk7aiX3GQ51Vps5scS8JbmUm
52dF0OS8hsJlZ6ayfhOhek2K7Xw52h8eFUGO6Ul/zLRoDNdTIzgtB7KIdlho0VZBSq3AJHGM5ERB
knNa5Ia1iu8XxHzrg0yl9dSf+whF9b201ck+jgd0PmQaeaUPUpBYaLBnTeAC2IYXhqWtL4Td1ID/
1CfQediVvTnH7eP6zNZLvyLAZP3jeldSqSzNPHNKZzxn1XeogviNdKb66IdQd/zZnWL0KQAceb8m
G+7iq3MiMroSJzyV/0oQK6xyjZJz6Ko5ZlDjEHN5aeM348TvJC17v7Szq7Cua+ByIpk7J9BBXnaN
BRz/Pa6zlbTWtDN5Rx8UsXsJQG7yjt4IJ/27DruRuRubm0LtL4vnEq5VsVWOLZivFLHdwyGN7uAZ
gDc8FyxUncD1BG3vr/2tAP2RipwPGZmzK5oC0cWsj9cuss5VcAGpndRiVqjRbqiO5f1DG96TSPKp
UrudnO0xeQ0r/v3YmdQNcdHhkx7g2xWX0a4bB3KJgh1ZNhiqYs2NsVj2/6kB8EOJgaQpGPYnKWgG
oGRV1wRSThoMqEyslVaIdRV1xNzLUppvlJ5zrhG513LNCff6wv0MSPd/P0qs2k5oYeacINlT3Nah
uXlopsJAy0erG7p7b2gDozX/ujDYowGCsPPKc2oA13FWZEDk5r7W1lZWxi+ET7Rl0MeKwjNwq+w5
RFvZPJj4vEY0eVRCCN2is8NtOICDqSK5qvPtnZSYuFq9gVDflqwyWQUp4hzRuzWSedq9A7osjYot
W1FlkxHnhOhzIofZO446kfhfpw4xepd9zUKbExJnp8mp3KpL3K3rLRk+kCgHvxk9l1QyXaBeZCsW
lZFfKCqGvM3oAXLhXSONSbAnWQelnuDTiUAST1mYCILtyn7moWF6MekO8KPN5N6EvWaQnG+ow0Tt
VvPz5hfuNl7y5B4ADWmPSZa+r0JT3jMHj/f5QZxTEeYyoJZZvS1elgqbyBL2qKmTdVa29DfV61sE
NOcSZsSGYmsAD7xMP6VXuQi3mszVtiVnIKakQ9mk05jgEzIxU1wWp6OcA6se24os35b46AzKq4oP
GGM/o2HfsKm1fNRaDaTDj15SeTbioscmmhSYx9IZ8XxZ5LZ9O6Yy26oHJubbGSvzhjPJqRaoqYzS
JfDtjvzvDL/03BkX8rlXRfQuQjhhuTev/mfZpEFliqyU1hMdEm2K5Oa4ISkrjrt33Xl5ETDQHb2m
VFb8XxsxfTzt04UIZEq46bnueN/xSvRNVP3EhieBoXBO5EPys1GX+oG9tJOYo+U/UAc+RGpBoE4W
ad12ydYMZhluTnvhM6EJgMzt53/+skA5lcS4v078MKwF+esm/xQDQXEySV5A9tiofOGFwljuMe9S
iKy1hQGXfhm/MoEI5Ur54WRanNjkwMxHE0BNexEb+CrSFW0InOBwz0Rcty8c5L/K66U3w+mXZCRb
YsYzug2KCVtPOzTFuZ2ejqh/Cx6ZrdU5n2CX10DvzmxrzDTl/Kh54XSyrytVwPYNSuAPP0IMy+P0
Tz4wx6qFWFcBbqNcZpB96kaidL75ek2FvpuW24SfTcU/CcgQNTlJjsyt9pLZ/t725wTz/Eo01E6w
1XBs1/KJ6/D0OahuwmdpzBrkRzw1KFmoX0i0TGG1Ox59qMxcSRzIu6e/Qu4gFo9VbSOdXdmSLiJL
wZY60mtxBr1ZmdgOW3u36NUO94zPgryk9ez42LOaKhCtphQDgm+ez/mgOrtZDh93DkChXMVNTKTR
3nsNFMKIcq8CkQAVzlGgjqCFdjiK5rpSDSmYBtGJPRZ3taJ5HkLB8l6r0xfcngTmMzSfeCkSTnQ9
RnCWBxgvCCSjo7a0JtGjOuVpPiG5L80X9Hr365LfAy81KGSg5dZkugP4xlY/KS5R7mPjI/tmvelo
OtFbxzQFrL4IrfzjfxZZuQ0Rq1Nw3R2OL6w4znEscZdCt+4ykx4Z5pS2C84+DEpXSqRbWZek2V5r
h7/aqfT0MErhSIQhRJmDdgeXoTbBmKppJ0B8u8AfVPuvbwJs/afPaOB9fhpJUC8LDXKfGxTWGic5
Bo77w/Z5Cbz25fI2xt7b1WaTYpkB26CPGSWAXKDP6irZPvPUUESpjoKWdp8FGiVAPdILhbeykHvC
0jIrPHKL8munXFa8B8yHUvnvYbbXfWVFH9GJqch/3DKgClL16HP7C98Jt0T3o/qNYMjl9AcOXtqo
w54iMTQ9bhVo/0DDjq+EVgk9NfUOflf18A4K5A9ln7JJu0M8uD3SCAB/1jGU3FZmkz5pWCG/+X+H
5+Z1e/HSZOaUCfMki7Oto8YlbOcmcxWhkgOIH9yDAo/IZ4bJSjwKXpFUJbK/alyrDQoNFrfG79vR
JJdHnvyTEbqPrnxdm5ZuF3WImgielVUqlkBf7P3EnIPeUKZ0Fi8GtB54IsxKoOKz7JU1bGa9vvrX
XuZSOCdeVmEmBF7+gVtcbfzNO4BDIPurZnNrNK7MMw724Cl/yuKgFMVZ7U7RUDcUS0MUnsqNcqkQ
wEjkACM13tRUmX06KNvrfANzVlrsm1rUDP2hvicStI+S5w2sej0vG1ssA+xpejPq/LmvnlWcvZE3
rF2nL5TLNM5RvS9zcnVcr9GSgmkR86y8dajmp1Hal3fK2cXsPOFD4dQukgaLFM/4lVzQuXQnaXjV
nKgcWMywRBlBI3iG9cuXI77tJMipsHzpjjr5QDdnRHIqxclStS7E177bPRujDIxlQM4FQyxQudww
7C11gFv6Fl0e5NFWrXc5HG3wiTgQfOJyyaGADSujqJarRc5kFLQL1zdl6uWYZAWAqdfgmAsuGvoO
fCEv44IOT6+EwcPZFkXwJboYvUCITMdNnFiz1As7GoM+6Bx9Y7SzcYvgkjTNGtoLH2KqfKhrXPVf
aavOVUrqEyf83zL+WLQFqOejyiVF2iMTkRP/q4ACbuEC/OvxqfWuZ5FGjskc0l7j8THWHt+aSRWa
18XzbFXaXRy8ejS99jLVNoCuL86ndLHM3rfGuzswzw86RgYaBK+0tKEdWpf/ufMGbQHfxolhSEg6
H4bJv0URVP6nt6JNE9mg5/cv9eG90PBrxuVqn2hkdj5i/4kAE4SwhMNL4yCWvaNJJBjCDdgpnzxd
1bLFb8jO/yRTlAdZeag96VQULPV3WF+B8CS3C52h/ttQ0i/PsuVL1GZsRcHRHfngaNW42xyP24GG
SH/2JikkU9/OwGy25OETIRNOKXTLnrYO/ca6Y8uFh8WQWTORpoZHH1f/o6vLH+ZRikT/SqxSDJJA
NoZ1p/Vumv+71u1iXNLk7v8iOslJh4I/pbV2BY/jpqmzSuZxeTcGZgeQgR7cfk0g4RvOID75yclG
NRryTIP+jeqXvN5f5khapN2rJuvE6IpXKxc88zyP7hVnnWhpXzoG6dIgEXrVZIJ6GwCdnTB4V3vc
D2URudhfbrmrj8gWy7r4ceKvuuMCq1Yk6gTTbinenYPqfltpRMxLVllYFbsWCOklf7QlDit5kYgg
BOU8sspuuMRZPQVGkIZi9N+jaNMkdOAkwxeJo2EC/UA/wswxpUCXGvQXAy+7ZaQ5vqPv93bntIB1
hAJydp9hm5xURfv/+UBQGs4chjAhU116QMkXYdlsDFEwP3NKky6rZAcLFSDWJaQ9f+Xmv/33RWM1
Z8ixhalXoVX4/aNxul7VfHbHuGx0F/5Xtm/AtmfqLOeHAlllXNmuiSsT0v/jzB3K52YepznppaWM
Ve+nX3AMWefnqLcbT6bGd/n7ipyBRSwb8ItloEPARhKnVH6e/1vvvfiv0uD9V+0n1B7ttkai3t0+
vOe7P08DQSdeUxLaTW9oaboNlljy6blbj9hWTATykM//sIby7fjSDjp+/Uud1HmNlPpV/EWXvtwj
JP0V2ra99MGFPbQRHaV+9aRpu0yeYWvZjxiiDC/N1Rs9K61pID26ccsUvd5hHoCh9QcAEc6hUHIv
qNzaj6lcqNBFaB36sNVVyeQ3WlNWRK6sbNMYtkFZVwCagzl16BKzXwJZfQAi77b1i9E6DpDGXTWl
AmRg7Mp0TjadQLYgxHvqfeffllpst/oZRsC1TbM0AqgRMw3fVUAnipgqcaRQyogcJ9wl4HHtKe8v
LeqVc1+LbJ+/kLOuqMh8gMg+xhdtDae3ojaIZNlmsqFQJ23ktvbaPWiF2eVAmzAHSlyx0Iuekq34
s+yY7XJTjbboH/KaN2U4wp93FgfDjVKDBT1PlAAEJUKyTWoAXsW5Ry1g4FZnfygLVg9cJXJW29T/
QVxB1r2e/34RcbTtrHzyWx6hk0f5s26tscHQQUZmeK1G5CYtVHlhJyKqOXkEi2pexOOVS+nA6/6w
+n4/JCMh8PZTxMtbNXs5b5oF0FwXS724T9WNQ0gcvzE1MJdgWuJVGlpfqIHi0wRoQLC+fK/9uxqu
8EWjI9f+a04yJ0lWxcSbB3sMAmUtecqaLnr+tTKtX+zwq6y3T/3riibfKkFzvq+zPan6ogJQkiTV
8w4DWD2U2ArrrY6E2Iuk4x5iHvpprY2Drf9ob9ie64H1p++8WTdyc2WVm5XPge7B62EG16O0vNMc
M3klj4cHcv2M4VRVKcjYgXT77mtgSD7rbNFqKMkJNEX6Awna0cUnGTS0CK3h21w2NE+EfIo9tLoV
xJL0fWor+OstJUSVNO/bmpHHC2/yeMFU85BuCjw/tSj33nnG2NIEPf3kNjhyvsdgzrAdNrNB5Fv2
fOAD6UqTyMXVuUcJ47biaL87LE+Z5Vp/MFYAre4BP8DqMEaIZedE6og2mejzrDDrTduWuArtQP4q
wiEdgPOIrGb5Rf4w+LNlAUb8iSdRP8bo3BwJuf69nJR7wKJqMCyJTv754y0JV8qZQmrZbHHwHHBS
3jCYX8GR9IVICu2oghZCYRn6DX8eLsOfs9GGzlytolu8VzbNqpPKiPmLDMshOEteVRm5k8xJitW+
0Fehob60vANZCeYlF8KsMkJOcDOjKxVvaKYdLVt3bAFoMNBfMyIDRsnDQR+vfoatkhH/mPaUJu62
Mfq/7UOB2YCignPlwj1N4ALq3KZACOlNr5POXm6bZB2cxQrrivLF4y5hx/DxwxEyaYf6kO4AdOCT
/UCoE4ySK1IW7zkf7LCqXkYIuIe717DlqvHqpt0+fK8qosK7EzEBQWj2Yw1NjST5iFXmBMM/uzpW
SN/Xif5AYIzgQs6y60V0wLFePgac0zNproJdEPgCIKgVBtgvSQRXfQHC8cmiKoUInEEvoH/SJKcu
EYVrd2yVsbqhp5SqvSQ1x/Kx0E5VmifbPa/iE00sKXdq2wVqTDpWizVIxxtn4EeQXdbUt2OK3biu
boGB+6MAfEdXe6DLSUh5NEeSsteFsxJnKLE49ZdybPpMozyDxu608CTF8lohE32cG5RVvfX3o6hw
Hrh1uADTUku/JvJFUhAPSltAlV1zw02eSMnJvuQMuuxqvfYNpg6IjF7DjmXEGI62Mdpggge1D85v
LhyUGBj/dHaP4WPPtAVsK0zrM+uKKdI9rVug57aJRxCUE8H2z4czBeVNxRtFudUIKl73DotiY9iU
23PFaceE3S5gctNCG1vigGsUQkc8xiq1YCQeAAVwiuEL/kdt5gPazghMUXusQKg9dq7PgVmFI+eZ
6UQ6uXdixmTbIYQ2F9/N/B2PtPbyp/5nJ039iQz3yViz4MqTYqU4uPT61nwPWhG2uNtT6X4Ha/jL
Gd7ffw/N6UxgUAFwAjJRcKhqKHpqzyWfB+FrerfgGbGbGr2DIIcYyc7G5XKV2LM0KRyWT8mUL08A
BGYAu9nm1d61YZC78/KxHDtpbvb0fybM6smVLLUdpW/+JQlU5NF+xoy8wih7zSInNwkkQFFl392z
V0I83JIkr37iU+ECGA8zkjO/aevdziyyRH+YkDX7tJAGZmGnj7dYtZUcj5Aqb2jAZjP+RErS4NOY
IMXvXewguLwj++afjPQsMIF20Ph4D+lA5n9gfq2dfcPCg+rt2ZPAz3tbvSShVvXzxZ3IiyhgE9x9
vn4q8qxkAYlNvdLxNM4e6qVR5HxmsZHFGGY9TrU0U6gFx7kR6lBDtrDCToJ4i08mXCQKYbH70iS5
n+EqrpbAs4BAlXUa0jaLruJd8q0HFGUisXusC9miD1hwhfHyb4mZ1OtBtOk3uhI5zOBfMGaZpybH
tuxt2z4jR9yWaPu6/Rqexc+8S03nzaTqAvIlv5SydR3xiaxE1gq16pf4iHjNc21EQdKnuasumMje
J8hSeDX7L15gt4iXWknfjKZ5rWvi4dazjdXk3mohfPrcs9sUFR8xEv0FAtG7D3m1MZZSb8iS3fsS
C3gnp53nwIMTUmJXsoomaHxt74cwzq68Puh3MNf8s34sCo9o5JxaODNSGLdyq+c0aQh9rw4rqiid
qGxZQAespCEghU6HinSl2a963OMDN/z/Qvphyfv7HGR7AXxL8Qlt1QeNhP0X2OK9Zx/pMOxMQGVQ
ZOksXlKW+77IqwtFIZnXYOfRRMPiW3b5c1Frxd9a0W50pgDAAKvQm320M5++mBYSJNSjhgrDTTnR
g2waG4vQU22gt5fBfHOISdzpL0P1MyrDd3umdGwo0nEkyfmqbGyU9I/4MpJpQSNYLHUp7ArBkzLW
mCYpdpbF12iwmNoeIs8xO/H8/lF0+u80Mhjb268pSllg0cFfjfUaoJhnteA2w1DDonie9keRPDHI
4pZbduUm2X7GfIJN/NJP7GWB7HaR37ZsqcD4mLI702K/yR9oGwiPW1KyV/fufvtn0KmC25cBtAhT
aWNIEqoKaNPPPWrUjxBzB1PU/g9F/8nQCD3VHFQKPPpMK6QD2DPmU3mpzrKPImCGc0bEIXc8jD4v
1uKq4ez9nlhTn25yYkMOU1KkUsuAiEPJMOgfyzRQvmfXCKHyH9bOxEPmGOa2fgH3osIta1nLeWMM
RpLA63DtXBYRXbEuZLYheEX/BYmIauzYYHQKKqzbkgGrCnvpn/vN3q6XcTqaQmH/0Yv74CKEA91J
X++jISkYBY5WJjJPX39ldafIEgYPifJ1QgynHLoigsPOZ35v/WqYBqM03P7Ye0xarFWsrRuMdYcY
/3r2ScmcoPUrf9PRCggIBTJuZDjh7oJhh56ZGL3ozHjFOySy32SGUXZx/uCzuiCOZEOF214j2e7i
jty7eS7BPAK7aMSWorOO18mO4+m1vVxPh7K4dbf1rXFRl5/E84Nffq7Ul9PSJpjoC13aVD+MFrib
nc13glz3JgFPvH1F/GUx4D2EOSvNMO16ws7Xx/Psl2WbL7V6oUkHWZozom79+CYQpfH1pHdZIM3N
nHHCLTs5M+ZiB/f2Pz9v7y+1ke8PF2zjd2v1FSgt0O0bJCt835xn5IT9YVzP1sLPMEbsjk4oNpXR
6RkvHKgpDc7wJTeZzOJFhsZA8QooG/o5QSHbgRLMV7bsyDatx/Vpwf/2HNS1D2hTj7j4SIK1VNJC
CvK4fp44G+WJyDrnzhMB2GE9rFX0jVt2jRvVHHzdotEtO/L4NW3wx57ulYsEwYQRHH/TMmsLyC+U
qNwR7PVacRR3yUhcl5j2+XqEyRdmMh0v12NRbBD6uudi/GRQK92V87wOPbhylba5WTSYR8A6jHry
vYkSCddWA0eyvI3UbYi1LpurcKUXPyg1+0pdeGOWkQl5KZX5mSX3NI+iVaoKSdCKaYPtDJtsuIX7
she0vYab614VWzCGLFm9LwzPOviGHUdjPhPqOFfEEZOS7b9hhH0U+aDqVX9tmRv0J5YFBffixItX
q1Uxp6bg9ZPVTlhLb0sU6l36Gx9QkOZu8Ts85YvnbJb6KXiANO+z18jdJfApaBjlsw33V0qFdojN
th3lIlcmDGchh8GcnvrNNgatfT6Sn+IBAFHBAq3daqaw2+NRgO9+MNwSgasvN1be3mBd0/RYhzet
nVaVgjw9Df3lYESbawBh9C/UjhLjz16VF5rFglVKteXTgwwcDKNRi03bx00LkyKLMxsJeL5u3U98
GJh2fmAuT2mTkkiGmTcf8gHg42ECQ/gJPGWaQNorjwQ8o1g+J/vZiDIYhmmc9KMwuzp5IEMOtImw
TROy6Lx7kRV+44KVzkDvJt9VrggmfMKtYrAQDFYij0p0AqPbKe22ePvLmnjn/aTvUNCNQKRVuvVt
/gTNXJQ6aXglr2RW8ENW6MWUEMFSTjOlx0ZDeoSieOpYFqSmbPq1Z395M8Kpk41BaiVPMpOjGwoY
gShIwukG1n658hJq3qOFUYNKDoPX6EgR1Wo5JWwODlieMRx56vntqTCg395nDJ4MTmIeNlJYoNtW
d6N1OPambJhhF6lrlHcadRDdH1Syqn1UT9itmmgCa6qqaA10HA+SsLLC/1lhmeiKTMNQvDNm4Hw4
gBMEf/3ZPff9KPplM/kX5a2IPYoQiqoQC31Ijncn8huf6wB1wvja0FYctu4snAvDNPKJeGseGNPQ
5/DMaFb6r3O7n4IeV1hhuqaivv1mIcjwGlUBZ2jpYOk8zfCkQJNCF9fLzsyUKcMNqcIzgwQaxg1N
YLRwlY9Xih/Qfz0Z7nVwHw4fNFHH5CekTUVhtC37t0BE+Cb6t4rh7RXyV1OT8fWs5huLYCOsNFUN
hlbKduIhn9VswWkGELtvrTEfNmNGeYYYAKau3Q4rfLQ4r5ztF3yR14a/CA68VTtEXSNzd11rFh1+
YOj2hQXNx7LveMUZVD3henXT22hhi7XAMHdYOv8j1uF+icdTKvIY/Ji2heq535v3RQpmSmRstEzL
UQcUukKqb3uYhfgN44af7928Cr2h4dXIHhY5yqrPCDT1zZNPGmHHHcqek+jpSf6/yY3vo7i+lui7
tKB8lP4E6ohFpYWpss3vF8JGDsDim+5R9YsOcptvBocuJO/5tZVZhVLAoRuqQCxfJF/hps+JoqIi
txPdleE4Ya4wYfnkB79g3mAK4TYgskifLPEa4nUdoQmsH3yiJooVUHjjQwSpEYiMGp+wV7fmApZg
fYksOecl37omLMD6BlNMGymxEXMPWNJBQK//kYsSO+chPI2Qkbleqhd/dWa9Nfnpt6iuy9Z8tE6C
JEHDqNI2B0IrUCRygNd8oRCZBfRXH5Dib3TBF53r4uaLjbRPHKEGK+kGG7YiaXBBwIpB6SEEElAO
lziRZhSjXiY9dVyOyIGdSVJ0/h19+ID5WCMnTTaqMtn7Ig8ep7r69l2uaNDZYPJT/qLljHh6Q+OG
+K9ieOEEYKiGcQpGE6l4xlW3+TcZ+S2V4B7zBeds4GxtqxUvXJjyB7DNLO4uPNpwlTuZCDHr+kAY
Wv3IW9ZQQgf8fqRQxUqoJ+QfC92/8xtmJY5CCSPDtzTW2MxWyvaQ5emH5bRdwS+gPA/oS6xddVzy
jn28/C2RTTHFJi9KGNNmD1DqSM/o8A87uUaAlFu0VkupOMwU0zo5aUx+cop9/5k2wf+DZkOEJISB
wKiGugGyAfsNAbMrsoZH1Qbg0Pu0XxxDI8GHG+bTpvx587lUhdJ4dykfYkA+yUNRrsjdAycEV53b
L1g6G6ElYGRBNq2m80A3JWg2HyIACZt6Ap5SVM8fRlIKjfOxW+ipjiEtCiST1ChndfxioJssA7RY
G1b485n6rsVcCU3Qffh9b2h2WdPOlQlfRFChuqfHZ6ChvWn1HGeiKKfCZWVOxuHSWJ7AWE4lMk4U
hrg/Q6XvzoOgxP7985UHgv9YaZ4HrOcnRH2n89i/pne3NzpAjLHl1KcEFb7JH9Og2TTWifQ+ijT4
mgm52R+ZpJfFcW4dv69S8ugOxoiTVa4IM4c8fLf5qlNpw/G4b4nLWDay3oCvqtXNdtd/NvKnoQQa
v00i2oHIzJzbi9T2Pk3g+t9ik2c/AeVRl7jgq00/eAsDLAknGHuH85DoY+5QxiNeIYHWkXu3jhkS
xIBNp5AHPKrG5iqLVDBTcFfOcFWW+EEhw+BCykh+3/nwjf9oHh/Ckgbizt0fPwSOWgu9GYrxiOAq
bOvyo4dmMvlWMh75NCwBjr9zorMFPcWLV6+GiW6co09vUPALojYMQMkAW6p7APsqcBIo/n2mI5rF
5HkR2mz7tryv6XblhqpPaJrnOO8c94hbVlhwUih4uZhEpLulq97+FuHOQCz2U79PiiHyo8jbjZ32
gDK6gfC9KBuCyoGB2xCWdjkPv/xaQiNM7yVuLsVFHf6CNeqnZ67X1kfc4qzROP4nq0w2I6HKXIhx
vdb+OjTQU6mW/Ip4oBNh+QbwVGsdtMi5a71VNsdEJldEazVOcxlFwjwbnXaVuQmRXVdz04cipXae
My+NqOuAZ2+N05tpQk2EPdPX/sfMvmKJ+3S2BNoRdp715flbsqHGIZ/D4M/X8oq8BDA2KQnLS/7q
j+/QL0AyfsCGNwKMdIH1aH8Id0GLu9PG+1fofsIyLWxES1698eoY2X/iPwR25JRCQuQ1+B4UfPq6
yQmtzCd4ygnPApD4AWJQSoWrX5ddPqsfFx4MmPqnpLJYb7F7aTK0aU2YQnS5RqmcAo7wP1q/1Yy8
K6e+/G7qOyGoUyaWPcmS24Y4fkVGoE8505ADaja/r+/O4xVKWa/JCHsr1ITkHmiEYgvCxkxczii9
buvrMetnaE9mjHPqEehb1wZbESBdDbezw6OmHpICSMcOgMJcCSlPa+gcPFdkdvzHMwPqoKEbAB2r
B5nFC4V0TE3qgBrGCxRjWFGGK942KFRBj9LYD78tl1dZc8C7YsQvgBBPicNX6IbEffdHIbz1CSWt
wygUlF6m3j1EXfzqkx+Jry3/EIZyjdHn3d2xmr/YMQ9VH6ZI146AybsnQ5iUc8f5K6VY5pcXYK4S
lLW/vkCHhiX/nl3Essgz2P9sz+X62j1erJhEehRHLHvIwir3EIpof4pkki1DfrEwSMwDB0ZTzx5F
vH48NSn13ceDarJPlVEaayZhoKaBbeP21Dt2dTxPli70Yt2a/tD1s3uaR0EONlEHKoWD7TwViZ6g
tUE2rzcCCFM9WfajgaXqqJ3YDbB5fh/6GSTEaaLJo7U8w3JdrHhFpmBAfZ+5QIjkSra30spLur3T
atsqgz6UgWK235CrzbdA3iBwJko0qwFke14V8kSZ8fQ0StLT3z3i76VdtC0Rd+3XHr6Gtl1VlOjL
n8+3pIZibssfCKlCz7hwrWXcQdqqqLe0NqTEsbit70Ag1BeEDtnhSVhPUos0KUjgBckSJIhjqibe
MxM80LZahHcZ5v2zEe0DeMgwg8wdT5lzLEKvH+MHRjmc/HxukBdHDq3sG6HXebMyweS/09AYYW1o
NMclbDztn5ePHEEGNCeMXCr27VekpcJ6bdUwPs6BNc9bTmXh51Om2h+OQXCEApzg6r6uYUOfILVe
TWpC+pr0BnQ9P/WAU27Duq4idAJ7tWmCPokBKzySK4U9A3Rx4luQklsmzqJhh9GGrrrN7dgQyTdo
ikVq4CY8NIuHMxJNcJD9cJ2FXukEQaWSa0sWwygtu1F+i2qcX6VMHnQlQh34NXVooyBIl/o2diG7
H5Y69b51g67UkThh37jI+/cIIR3ZEN5g+E3PEF3+f8SyJ2oMSXwSshhkfVy4YPl5wZ2MJ3qNH0z6
3D6kOTuF8CjpWJp15ZnZ2OvGKpdwsGEB2zgSN5yiKHDb5sbaVllPddZ7swS1Ai7WyXvxW/to7X0L
QWVPPchR24Ny3+l/kdmk7u/6rMhs0was/p1+LpnAkPUzMlYV6yYPFruIybs1fK/6h8LVltayaONL
+YRnxpudmcWLC9cCj/NogBTTyGVeby56GCHXOW84+tVpF+b9aK4Sb9aQtVGkgiOQHsPBVgjLpMZg
E3Sz0HUiX4cGeXqjbqe7FOmt9+gkM2paycov/koVQ0C4gnr+PSTZrqLCS0eDhKNNInTkByfNlLRj
Qf8l9BKMIeLMpMh22z30rQ7CXiXAjx3XhHw0hDGGl0/OtIJltGOMn7ho+R/trBMUgBq1MykvKQRH
rGZ+HNkdcjWe1tWTDtsFi2gorfvb7QnIdGWHn67UJF7BZazBVi7ooSB7HNgu2L9zvTJqwNJJhVfV
rmFl68GONPX2mqwlxN790ukX/8QhoMvBGnRYmO7MHI+2m0xcDLR2fwpAW2v+LrM4lcIBrJWHxMYS
3nDScK9jgQ3TX+VRNB18RxkNQMuWrnjUFOOKgHlg+ho1bwSarGp1o8dzxmTj0yHjyglW3vMa1/a3
jAL6r4dCkxQNpk3QF129869yc9jpDO+UaAaKlc/xxtHVJzPDdcY7umyRDxRqutvFYCQSV63ytAbm
dhuEoyWdPQfmt46HhJ3Q6lXJKWohPy+CAUEmk9MUC6jyqlhUuy83Ar+n3AQVsMNU8jq8CvXLhIiD
Chh+lRnvag0jUvl+cWskoOcXI0u1l02dAuNuYgmElaAYe6Wotg0rbAD3LWjVHa6tSDvFbjHx29I0
+DFxLbV+ee8KYfy2uCPZ30CIFGedWaQ+Ugf/XHZV7lhjloLTjO4kd/Bs1t+jOQWIDvcGB8AQ6Fu4
SrvnS0bIYs0882I43ah/5LMY0KEUUCWgKcdffZU09Pgygq00DrpM9HmG5N8cfYPIrZ7nIQc4rjyl
T2oDbZfqzXJeqC7j/90Yd4f5u9/VP1MmJ4STp3TpgEklg3YqGOO2Ym27Ca7/ena4jwWqC7qzhaN5
s+nYllosMqy7fR6ePCF5E7VA52xqHcGjShoGxHGqx6ck9B30eISK1QLZJz18adkE2L8ZJGq63QQ3
0w2Apl6zZkV/+OgQAx+pr4yAMa+xfq1o+c1n0j0ebOV3MfWYW2WYQx43Ae2hR7LpaPCEaJk5k+aj
DanwofEhmcG5tuOLpGp2OWjeN0CSvMDj/8eU/3qQM+08Y8GlQj8kA7fHzAWp7aLE0Fz/q9SNvfL5
d6q9jLkvGTs8mWrqT/hJ9Joh0geV0wskYNgPCJj4idPhNimdK9zqRXsfAQo1Eq+7qY1CUBaB47FB
3kYIsd/gqf1pyDgdOky6EjLUBoPUQB6nI7aAf4q4hhoi0+QzOnp5T6WNcYM5IJVt6cwqclooUqeB
CJpMN6JBXEkYbpt/ghQzXryokC0wuwoLtOJ2OJSampLPwmVARIAWLvpCqjAcxnG++omFdRpXiY9W
NDsXNyyewbcxAZTizcQz1BB44GGYw4tkNFGaLKIwJAZe1pUR9Z7CDOpdZdTEftMTbYZV+6FOL5m+
vQig6MItGSVbmACwBCfzVJ+3o1vDbNZ29WiV9dWdiwEPV2lc8VsIVPijTHq391EfPd+4ttcku+8e
+cM6OK0cZAYdcvqNBuEJzwPXZ/Sj4uVCbg7EjTS0h4hRtsWjutNs4iTMZVgPnkI3kPl6TA9T/nuT
LPZE6FeJCiremnMDwfDMeznNrh61cjQh6bjn4tF3yObgOtOE6AvPhor6cyWM6Ccqgd7a3/J+guJ3
ZYx4W3eTynDr/oRxPZuEbb43OL0RmJLTnbdm5p9smQGAcyjSXFbWZRSIiLT/cypnkGhvB9YYyrlI
5qW8+SliwONd0jVFpwG5Cm81aKqvLqqboVKiSjdqq6y5u3HgHL4saa2pxQwtNYd1jO8g39+e1JDk
tJ6awAcPbGVjGLKqCFnskoe4CCg+Yy35ID32QAvYqlFdDuZM21TkK10A4gPnvrSJBT47cVs1Itav
Wad3bWttUHvOJNUfzh4grHDtX3RyQ1hHCr3CBHyvfmYqSOq9kPIrWmrXOQdh4owj/P5FJj0kLXk9
AfAJqdIwwDu2NOCZa+Tsm/8Ay/H2wK1j+C3l6NhZzichf9QmiuisoxlFicCEBm1wXmu+qJmUl9f4
lrkpSm4b6XEjYxaRM7i/F16A4Y5ZjCy28+t1Cq9+P0Iyo+WYvxTuPZT3gF353Skj2JLhdPeuTsiG
IxIrEYJP9sNu7WuSYY2aFnSjQ76Uvx6j/O+Hjf55U8DHmn++2rjaD6pI1ia8/k9eP9SlL4tnsk5U
ZWa03al7hF+9xNcvuZXSebQWwmpUca9Oy7cu4kHTJVSxY/Y4GMTI/ayHpIy0e7u7ILv4kbbF+0cf
X9lt/yDBkOStIIdjtxJObhnNrh4wjFi92+C3/Ct8faRKZx5H0/C/TRZ39KXUtA4MhTO7XDS9aIpD
3GSP9UbPcz9qz2ei+8WVPJhJghGld3o4QfGNK/2+CmI2nmHDlUPnyacrIC0RoGAUZVVMbfz4vKMI
1Co/os2JA3Ae74UrpsizfmMZLWFDXqi6tKyWVLJi6RRTKahM54qZbRMzliqtJ5+tUtq2J81LlklM
31uMRv1ioQ3QOQK0qcTs/2nQKgBomh/lvCK5vnAkmRjvtcWm/57AdKov7eFo6gHMepsAVgoVpA7+
0oVXs5mRaWLBNqbrvHKWzllfHz4GTg3LTPeBXut5LmPp3JVZQXiimclGcJDsYTJjHvX0Zgz5eV7b
6u/OR8D+Q35JN0ZWARvj7+I+u85w0UPy5AMgUuvXiJFAZehPPGFfSyX/5IXSqhq6NdzTV6HMLESF
O/9v0/cAr93g+sizZSKYPRNDoWz23YZ5HSOzXQCpTcxzvhXOn9+o2Puwqk1V3U82Qsieac4BeRrq
2Ljdl/UrXcFY1Z2rgesgN4D7KdxBJhGXpdhX7ioWOU9ukJuSjzxFAHCp3cOfzW2uAS+o5SOKQNoP
PcMK6bneHIS/cq4xW8o8pha8+ls4TGcqLn6c30Eb1Pr1QGNc9759Zwyv4wcUf8Qlaovv4nM3C5V3
FSEeTas38EYvH+sVKQAq0HZikR56hAdJlKQJCqN2QCI4vUqGUK+XAyIgmG+cjfRJVUrsAsTd27mv
1Ebgeio44wBbP4h84eliP8wqBw5x+U/3vqnvJozwJ28Qz/rwIT4FHFtChzPsBCd+Z+huvB/QDmjT
GcOlGMgbX/AG+fEUBRQBib1uSrtcho0XfAw6+xZSpuE7STq1apgS360+KXkuj4apmXNzKsRfsa55
msq5c/yvaeRMw0pv6pkz9V9NvWFtYPj6nPkKRVoDIKTZhdcENDSl5WMad8J6esYtHN1RZTLA5Osg
hutRofu7M9Z6JYVDLsO2KnA8IWPARllHALCD++uHf9ZvdYGAU+kCuRr2QgzqWnnv7FYX1u66WUmD
DkOQAoK0Z3Wo8eDvG+qF6GQWHd9RAUQfkTXC3Ext7qve7hDWKviiL2Y88++blyZWPQRo48Hy5fBb
eeQMdFWnSBlukPIqHVVWxmeMczCK0r0NoY81PxeSwqNwJ8OvD84pgod7WdYDwJ8cxT55XWcEPVYc
Q26moozpzfUUrN2352j34zoOhs/ZgF3P1KFqGS0sF1GhjmukiAufoZDZncyASWcfg8twmnnORPPb
Whb9LzOHBWvm7qyF+puRuh0Bb1uaZ8TxaOHTFDn70DJL51/3qojVtDyaMKSKgHoBO6rA+FWWeIxA
pxSxv8pWDEoSA3Rpjk/LAY6Lx06eXiX4Hun/nNvs9d8Bq/AKfJ/DwyECPXOxabc6wjLakWZKq0zD
679Khfi2yGKNB+ukNgdFQkRvp5P95ZqhZCTBAE+HeaGcL9A1hw5dPx9MPayKyH7me6rvLnn4x7lV
rj3/g8QX+C2orHl+9JZsD3o60KTRcpxvLXSdmiBetAqzxBI2OIHNbonhIoJvqDM+QZfOt8i6Ugge
+DOneyblsTC5exoUSAY4I21IRuUELhAnyEUOXn0mziSm3Zw3V2hB7D3jm+P5OlcVugrHrHfykZ6D
jtoUgbhTR23mYbnSyMVqdhxhlWAZTj09ZRmdc94Phvk1XmowAeYS23FvhHhL7hugud/8+3PNxaFP
gC0tGN2Oyhmf2ewV9j1nNyQnRwMZJKEwSMt0P1PSmCSWrB+beIwiW2J0x0QxkQSj3RYh9jdn+nYO
5Pvr2YO/xs09cM8+8u6z4qsIq0Cp+gtwX4mt8cSDVLtvZcCmd+PVWtOUKPZvlzIzfNgeQ343cg9m
189t7shj24WNxZ5MUYdOhymtSLLsZ4oLjozHSci0hZOmobVL+BlaGHIpjJRVn8gHZPW1XVsiGXjU
fl2ILqx6GzejPa2AdcyX0BAQ0G0c5yRD1v9RllmF3nqQeKxC1UUrgpd13UM8WEBDSapATyiSVtqc
/B/pECS8yNhxMn+o36UbnhHJAmbdPTZw0OlN4NsMGpNwegxNllLxjSHdnzjZMAI8g2hS9WhlnOm4
baaiq/W5OpKRBB+3JAGoKz/3K98j4o9zsNqdldaD9Se2WFcWEMnXz6djoR2kIi2WhmdnRQcxzzYr
nm+uv5eXPbY1i/ini7o/dcfG63p4OSDfoqshX6903jQ70Om+kfzmfNpeWn8HMAaTmA8HnqyopoSP
7Swu/eDAG+zG5Qi5+hhYZLSc9Gxl5BR2RdjTVO6kUnmy4s1JHHY9YoMKI2sfOjEk5oOgWJh0so1l
tT4jWgRTTcnvA1BmbcMw/jPS2kyAOKMl0Jh+X0WJ19+8Uh1qTOdIfyMDGkq9lqqOuGuLEm1e4Qcg
hFdi7t1HOSXiYooPRam9SZBQ4nCfsFqVwiYSHZwJZbPFnl+sMHPl4hyJLONVA0CTgFlikqlRIo7x
hJtvLz532sqb4+nWHX9dVym3cxxtf+0f/EohvwWFlZfXuR2/GFjdfhiz8j+w2P33kcD6Lgx+9iZ2
fyPnIlZseP/7mrMnVnGQh+P+czfhqVpytSHkrOJOvVvhXZPIneqf3enAF1pu+tT/JnI8esnl8sya
5AdI1A9B34kWJEPg2idC9XQ5cLazobElulwIOypYZuSbyqkUIaDsEV34R6ytw+LOHP9IQlQbmQM7
1/6Pyltm17FAMtUuc/F6LRpF3T3D9uZZUZDL3EYpiOFA0GvUmwlWlcuyrAe+tk3QfsUH/zM3AtSz
T4V0k3yUcqXExwSyT7xdy3ZAmyEd5Ve6xifr7AF1+KuzXTrUcDbp4/Uxuj/F7U22CSSeHlDiucFW
pCbVoq5j79WUv3p7qhQlfT2+WJ9OY5rPMg2EySnp88VKtIu8nSgVjVmCLowaNDBNPXHswnAXF/Ga
5O3WQ+sddiVDW0pLo4D2Cc/OCkuCKpc4UCpyNX5u/YJrGJdduV3bSB/d++CCDhvBL9UeI96fgF8D
Cw/dOiUHJaF6NAUrRwuhUjKZFr30p0ym/sxJvfu+c3kNatCw8LVCsJ3fS8C+LqqPn/dqP9PtcgXR
poF3qqvdN9uXGsOwmX4pYsBzFbdCBdR3btwnfK8GH+SmJWSNoBogjCseczxI88k/wkt22MrrV6ah
N/WY8c/TmLSOdDOsniOmMDb+zrQL2f4LjSmeuakyli5xYrzWN1mywQi/pSJKoCM4HHZQkIdMLiMq
HlcEnP+nLX4J8i0UGqu4Uv3y3FrYGrKVb/3C5qspGsgkYra6P2GusauSXS6nuIVB5H1BdAT7x7oK
qvn85S6WaxeS4g6H5ZsCTzg7EyrYRRLWPD37xEXPsGHEPpp/ccknuQaZ7vuj4g7BuIOkONzSPFPw
cZG4Njkb5eSCSBPYkPy/3R41PIKJ6lcgG0Yb07jh7jPtPOdBMydrMdL22qezsuoWN08aw1bzFAzw
5314spoQtb9BUNG+d7iJdmoIED6mhkmMg7jqnIuLESmxAAxpcdcBG1No7INPsfuy4EwwKS1SJsDx
PTZDNbUIthsdbhDL47pfUW7VsRW2pIFyNlAvLLdHvTAizyVjkeK6B5iHxxIsIV+kw4n8wxmZzg9B
mrXPVDYLZ8414wc9BMvwRF0syskXDUNrALzlASFWmRNKAVuvLjEOxWaQl2hGej8GnlHBxX6f7Wzo
FSLRPxlz6+nz6ZIu2+XatASI4oTbMT0k4YpgaLg76fH/7Wh87dPeqbBCTINL5HUXCzROPdmP5gAH
EwvsA8Ncvgk9mns33XNfdKGqgOt7YM6bLleqmFFrrR6SslCoMdyzivacFDDJYl/VoAST0Il2kL2Q
DfxyEhuRC6bCeB+m0d5jkUYD+8IejTMm1DK0C+M4omkUIxecvwBnr5wSgTRSn6GWJypFYB75sDiL
iWogBL+9SEITFCMYD1Yyk5TPscZM6z+uLFwGC7AZ4JVsO4ZRw8o0GcdVDd/ZJnqBnx8wOyr/CYnD
usM5UCvEXJ9lNxWQxyKaz6ukSAnmcx2T2d1gKrmR5cD8zJRy4e3jmBpbFC4mkQ0DJEsVmgx0wurw
R6mZWl3aku+w10zqoFVbzxXtZeEN3Sxdsf++NG0yNiPhhc2pjbieUwHrBmM28K2LhmDpwdlBEPO9
uk7wY+ZnI+fWr1FpJsIlJp7f/kcJmWJLCgZJR0cAHlpS9C0YZwTjNTL9RNXdDZqxqdh+Ti2qX/95
a3uB3WHA1Nvbe12C0S2rN64F3N2UCi49l4nYsG42zyXf/Js5C9wfK38VSi6KEJ1HRKrLY/98eHGQ
gXCa/DxdCht16Yhx19YaawgrzNFWZ6cbt5rR7jaoXwyW5BJkRJXUI3QVl/2/+ogDjM/+KnVORy+v
516Nw3X10w0xRUVX37pcbX9cqJzTXAqAfC3/6b+o0OFlGXCfwAZBTIvCX6fiGd0wHtgFyflUMEon
p59eXZxvXZPaAshBH4oPD99RG9yMf5cxH64b5A5r++rXKUgBX8BvRnVajQJKdKbbcaoEq3oJ8XPK
Uzv1qldmZwILLW0yAtDjBMhjSk4Q847z/G/8fjC2+v6u1qD8n0uMcEdQNeYoGzzcp9dtyJyOhmm5
VT+rdTte3JnnlKSX6N7ChkYjWmHKiN85tQJUtmCGdmvrAf/q6Ias0eYWaYLhxTJBwK5yjYsyXM9M
ZQVXOXXnvyGbr70TH3VH2bs+e680omiJ/Y/gNzIMN2JpWe9SYgZTfkeCicOgVOfRQesZ4Xa6aXPx
UMEa8Q5/0xlLDXYXFO6EpbSQp0vg62vp1xqCnlkCLxIqSgBYJ5dChaHR1ujF/0Q4RrddfYNmpka4
tbmpZSWj7Xg27Wrk/+GuJnhkua7HrOXOAuNfXysB1OHaNzEfk8nkiez6M4usFBVOLnWgxUwerxaj
IUiDyYz3u2XV8OFeCqFakTXyR8G65cdMOR6JqHALyIh8HVaBrgJA4TZUJ5vohQh70SUC/0ISqjpY
0RW2A2PoH2D8609+UEv0xWaXXTb5T0sPT+7jHdv3/aXVMF4nIjuFoWXEoHwcBirSk3kG3SXVRRF/
jO+2y3jiEuZbsJelZMMhYWzMH0LZKGfgUW4T/IM9pcd3InUpq1eQe9EzsWdAn+Vz8Mymm3QhWSU7
8O4+pODOcb7D/Et2y5PdM12eVaabrTQskj2PuBnWNBO2oHsmEgWjDEbeXcFAKcWpBuc4KnJ26TB7
qJnnMjUP6J7OCt9wDd7XeutZu0wsvfEHyl667vLT84uWMD5GJEmfqykenV3iZ9PQ0g0z76FjQaDZ
ZtcsVmCu1SeLC+E6z5XzTfDnwJfaM9uqi0++g4/kIM0W+HjFa+pVmZUkSA/OViIOojkElu9gv9/K
qilMIQdCpfVf1jtJmlq+TveqBd/4wObKyKo8zILOMAgr7WqB2L/Sr6DlBhXhBQB1oY9E2NXx5uxq
Knhr4Vk5rX9ibe5bWRhcf0YQT4uW+5Gw9Sg4lUfizx22QyfeHg816+937HGDXGjGzLBmP6DvurVz
VGmqOcPPkL7L4gc8quNQGTZ0qvCeExSAoyNcNzxxGNYAz1PGJbz38mlOoYTgTYgTGoCrZYiR7gpT
8pI57K4/ISzi5vWpIvoC2rhfCdNSbr48oyd6IWxxDwEyYeEKRvzxU9yL0l+0I2iFSGxJRRgcHdcc
4EzOU1jFkFlHZkmzNP7VOn2y61/bO8PfOAS/ie9kNQQyJkwm88LqxIfndSvOotSK43PzRLG/i0ua
IO/6TJAVR2qhVkqJIxGtnITw1h5V0yP9o4YY6xE0wV1lgq07N5I5NK32ztgVResp/GMwCKsKTbx7
QjE8Wo841KAuNLgLtKAAm2gyW8eIqwGI56tMk0LbVW1LFt1ERtm1l8ap67e7CrgrHBxH0iqLU/9w
kqlTSFJBGgnHpNfqsWbuA1hgi1xKPWG1k7hHIOLfV1sms3YGD4XNoeqB0TQhd5LhPQS+DC27DDPs
woi2K7wjwKyd8be7fk/D774xvR/PIGNyzJmst+dwhBa6KnGLQNftFUj4tPRY0Jw2FuFLJ1SV8Bc4
iXGIAHPN/jJGlDWrPTey6D24NPGnvAUrsfARoeSIAdXeR4z/P9cEC3jyHlUwCLy0mMnSLSqDgz5V
ifPvj2yNuqOnYSRS7XQyIjVozTEa0MgpkqHabY9vQ1hM5GQ5uwUiXfcqHOYTrn0+brYMtaB/BBue
IxiSvxhrYZCE5BJFKasIrYogQK9D7vlAkJRgUKwwbIxaTE3PZ90d3QZc/SSdcQsEJ2F/rqoePvI8
WIk+Es+lgaDJd8mfwLuCtVBCp2/wDq+aDEJwndDIyblHF/Q11nAyVm/SW85qGMuKH2l1b37nbE1I
sfRm/de4KWuPFh1GDYtO8vLDRrSwLfAqSs937qo2JdLIfnz6lEQ+XhssthQsBEDVukAXlgxpCE7p
DajSZjGPHMqJbAAlcaLTaGt6tfL+24ukq7KN9mdGjQNviDmurVOuWC5NHYNpzrq/oK5PtkmAz1Qs
b0C+PUa+blmAjAufO1rKDdwBZ7dxUE10dFQMYGykvAJ4o+KmjB5MaowYAhUcMCUJGC82gcN1RFLK
JUV95UzKDLF/ohlnNieIlpGleN3kbSpshcXr06MItsFCpRMxiEcP88xOZm1dF/mxAH6v9InAKhme
LYFI5k8L6VNocHys9EN0PcTG7iLbDGzTD4ouDY8q98G7TlxSurRGQrKutGRAKbYj4DfPZhhwnpEk
yoTdlmPWIc1p1ieI9IrkFefMczr8z8ScPpuJ4DQRpwUIu93DvMVFvo+CqOy3gE7NurReEx3nKD3Z
tqfZGBoEl5fHjcmiIob9zv+ILG+YEkklP3fkg7Mo0tT8t/mFmN1V/mjNgy0o1NCGd6FZlLtGmuJF
ZXZPFsgIHmi+aJDjxISTM5lHx9CQvHxBAwm/x+i+Nj2EsuqarMTE6oFSPyoYpSKNSS/ikNsmFtOv
e2IewyjPIa/i8SPE+SHihftI/OCwgXB30EDsGh+efYbqxjlXcHet19U0YNGM8Wd7HGkCM0wjUxY0
VQMbZmDD2vrj/dzGN+O0mYY+cwLhOIxY0BzTbAwNfSXYiyNmTluwEOE/Kg6kyZsLIYwhZNPm3a9p
ZaPCrdQWkopnTQNCxjjhq6zZv/LralEOOTcntgi2tbUPoP4LSQe2PUbNjbhIy/vPhFIA+d/DVkOj
WvF9a9HCSDeX0UonTJ+8S68Zmg6VuO+10S8ACihCOzwvx51TEkuuSFEZM7Cs3MnEf5gUXQon6Yt6
OLVU50OT5f7GrjSs6+1pjWP3z3awryNSOt2vGwU/N9mU85U/xgp6vlfZ9TeZg5Mr/qVQtS9zufSr
Nu+uqzyAYP1hSl4VjSOX0OAoFoEelBx9curw0MSdv8/M4/vkQwwtbx4qa73K7rror+kTNluRBd4p
2AttoUbRAPyJDyIzg7AVt54kqbSUska0nLGpGbmroCx7tn7pg9Ueo4cwCc3NMuKuU0KH2qzDzkB/
9rmCjX4uf1WURFMw6+bNbBQyf9FU3pkDVdek3Fei9w6P+2LNPiWbJjQxBL5kqoIBba1xXdlMZQ9t
umMkV9lSATWz9JY+CD28zylV+UkFLYDV1VPUPv6IOQXT4pjeQRNnbG/wyVccEE2ckVnW2DB1h84V
BXZpCc8H0b/VBXX5YDfMAtwzLUWqMUIrYIuXmbZc/95+o/kN+Ot1dulBCiMQgECPlf9jzCTSksWE
3hBA15rSn5cnAMDUwrvwO34tKV53ZT0yCH5ufETae7YJ1gciIHOZkElCmb2NkX00ZKnb8NojIAcd
kxtjQRO0Fd1OP5GqRnpmiKt+6QELNzz+59HoI87ASzEb052XVTLYDg78Q+H7l3Tej96KyJMkIMT9
kSAk1apeyVb2EmUAj8FmX3HrMZWB+bDYg1kMQ6c4+rKwuy6SEq0dlbqU3om9q2S2+vFcvfh0FLTm
+ExTk2N4WMXadb7m7rjvzGJjDqNR0ewD9xhAsuFYZ/0u14LTh1ZYweJQm7rj17M1Vli1aysTmFgU
maY0zpPazV9QXbm8HPHhBbnKWCaLpWFlXh1w7OzizhUHnEpq/nPgMsV+uu5045MOSNqKkY2W5iQG
5Jdk17wd5w4wwFrlvYnTk7yg71Wv3etBM15K3ZPt43OoAWm8d+cWyMhDNZmYuTIsx4sXnOVxwnV2
B9yf2uTptei4RX4wU83CpVxt7vpDx8q6A5q290sGK852KixN5UOLNF1iUA5GFXWwuD5uYmhF4paf
BMb0cSJEZn+iC2CZy1X3mIZyEWJe5W0QJWjYco5n+bREcp1OmLFo2UbxG/KZ9WC/jGpiR/l2Qkm5
gC2ANDT9hdtUGwGveqEFWgnIsSUYbTp/1ru18RTJPbz7A6SaYGGrW5txNExuD7Cuy+zW9WTNOsit
KWbnCMP4bQJWftyPAyRUdZQWli+4oyTm3mHgxzOEQ1vW+r0kEZyBL0ggjBTRNpY+CX+5H4NkqKiS
/eJpAVguesPhxRwgBkfgQHQ17ZqCGzKvhE+Ty+0CaXAJbTs/rmfQzjP5bIYy0bWjHaURoc3UMRfy
KULp9R2TbJ9MX2CYIiKPyzXBapYqQU4WatV18WHyNjfJJkf4wdhDFmDxcSurWMt/BWfCmn6ltc/9
CBkZ24cznNOffBlZDf8eGAIl9yn0o4pDX13jprIK/nhdJqodRqDOqA9CJCYJaL1l4+jpLOG03+fE
UqdY+LroOujrQgU91/4INOy2Um3NDP5/mvjc1GYfw4isLaEaci/PxY+n8YIR24pnfVVXjUoFLty5
DmIiBkwDIuTUaT19JdUFPs5QDB75zpc4R2tLDMMBg3j9dfJBRrwoPnas6/anyyeNRCdcZEcAT6io
3lCL1rssZmizU5n9v0bNAPnQU1/MR0Gg7CPgHjepVoakby2sW0ZYr54yaaKpdOxYxt/YgQeeoXlA
zuO1pAyBks6DndTWREWWuDn45oOS71fluLeSxO4uBJXAzgzRN3gjnQclShoxGzix4QRsKfPZl0sA
ZXqhlUyvL6vSbdHa+L93FATxVxzDf4Z04XkKtuXeqUuT7hdbzMPffDtAh3H93U2/0vTIp3DO4W3X
+smDmxCX7YKvdbmQz1sdWA7bawiiOjJcaDEAOhi2BrCTqN7ArfpJNdXxInaeB/wIcj47gsBgM1Or
kMb25VGQsxMPeoruVDig4fBqCDE6OYil2FqeqPiC13w0IKm1vDLH0vVq8MvIOe2TckZessZjyqiW
77o9m2C6zx5wQ2n9S9xrnduCV45/XAgi5qHcnCeb993iUUPueteoEa3coQF/gZxwxOvvmIOllGvl
UU0IjwF9HH0XaGeraWjFop0XJoMuhY328PIS+vmANNKJz6Sm6gytkPDRfarsnDsEsPyvy/liQVyS
YT3YTrFhvnH/rIFBowZ8EvezyyuR9bepFm375QXbJbz5LoeVisWHjzZp4+juhp2H6zCYRElrwRAu
OKYRhmQnj8CAok+vsrSGK6Zh/uWm65agkfkfW7t2GUatXetsZSGMcDCFZvTEGdPO/Qy43c1lgf8j
ql1I4ljWTPoz35hKHV0Njd5ZlUz8KOb7SvA1cC5t04mtYyLDGrhcmX0j5n9QUdRLjEmlYDQ9R6aI
yBSCBElrOCuoIqulwJAuNSfrCGa2N5k4fffMeLbwjEIBwFKrLz1AsMxsDTghdN7E7c77c9tWkrvC
P0gRVNVMGP1d7Tcdxa5AThCP0MrCEKT3H16JIL3bjoVgCQmSPG8GUkP14zqAbqQiGSAc4XWjW99E
j6rWWpkhTY8aWt6n6fIgAYycxm7njnxjCow91lK9SHjCdxLR653gvgeilxISYMp85Gw10gb/7G/Q
KJhtO8Vr9O5ohancF3R0wxIVwUR4ZyJOYMCY5uCJ57BCqvR3nBDLfSSuzr+4kuPPJqkTnhz8BjaL
lqY9drpJjWDCOEjRzfEkCm535LgcURWJPUd4y7zG9lYWXPobpkPcFET/4F7pMmYx8EY0rzKvflOH
I80QuFokcNTs+CwlUwL11NdnMj2ejaddM3yHF0PEIFu9jspoNd7jQMU3rSCbjR1MGu9YHNH5vZrl
5cdWukLPckwo27CTdiA8dAUWvYpzybaCGMHmxjy7KHZiKDR5FOSI3TlWKjBBSgxn/YID/HFBDrJn
cG+UCK6N9A50GIwnqWfUgTqVG35hnsK7YqBLBArrJm+uvX0q7Ae/M8RNfEd6W6gIspM8/9FTHk85
NVce62bKms8S5xchIyhx+eGm4OpsZmmBJ95Gl+0Ss7M3wqJxAAnjo/zOuTr9IWl+a1mIpTcbUX16
UV0lG80ibwd2auProWuRxtnqmZOwHLNaIHnlneAfGs4060CKh+TSuuExAX9mUav/6IY2kAwOMssD
KvdgTBBOmsvlPFvw0choGLX0ElnOnm+jKqAiIRPwPiXWWJqqMnM5EKumJ0ASsHBRRK8LxQoVI2uV
3AAd3TVHYDeyxhmJXKeGUB342YzMtyVKMhT2pD+JsoV/J0SvW547eQKWw4tozceiKygoXeRRWVgh
EqLo0hiGQMaEgyGMaH2tqWjFANmmAMCgWXspjZJqBrWExqkky5LLhQsHE1qg/CcbljYjkPP64k0n
TKDiDJt2u1b5XgYRcQ1Sbcp2TkgDCf34rdDfRNcaHafcXwYjR9dedZyocKZ3kPqnpo8C27GTwdmf
bUgWQ7/XLQNO6jARVadZK9NhUgMJD3qfohUwTHcC+LGjJsd20YyhLhBhIDDpSnSEmqC/gNpnA7W+
kJL3ew34dKZ7wgnsuYDnjvNuKz0wkghl2GZIFwJm6HnIurG4uReIyVSiPCuBoFlpthIFFmCnS2Wz
EWbjLhWzTIGNFl1ArCIP2P4qYkPSVPF3lr1Q+nzHs45po8LnXc5mF+1sJoPs5b0E+0IAMyp96rvg
oeFqbm3hj658fbplVaTL5gvsSRgecmvvPVCL0MIaPP8mBiftd7+0AvqP6SOGpAgKzd0dpdKeV2kQ
tANl16151287QDmwyfC+4QTbAjW93V7WKJDoD8t6C13Kh37bU8jwBtIj94Msa1tlWrcRnAi5/cJZ
tr+BCbVtA4cT3hU2fLf9fJoaIWkQmLVZnrplhawzy3+tQBWFkqQS6x6Vwl3c1sRmem5y4iYGhDl0
wrOBDxNR/ONbu5SlRW353kSTCF77LxabSvARxHmjQsJ4admuvDGsYCs7sMKSusMrIGpZnumDvmtD
g9Jnzn5lMPkjTc528MN766emK/VA6nzagGlrVq6qgMADS+vhmMTblhbw8+EsNNOVQWrcZH+MjTWT
9ZNsNMnf/3JDTYJskQfrds2/FOA3cQayFktjHaX//HJt+SdTbDUTRIb5SAq1MtG9wFlzF28f0qJI
rHlumAkqnuz9xPArQaFl3Mttyj4kFH7/edu76L6Tb35NvwO6XfbU1OKpkp5Eu84LhvzEzk1ANf9c
98UyaZzlj8UbSGzx2zdW452TWDSjns//0+2cNUly/zisTXmcJmIZBULxb6iy7sZDWxazCQOwSMXq
N5lM5LajC96Z+4mygfx9Oaca3aAgE/q6a+p1j8ChhbKv+RGF/MT/dkIHcLIjG4Wion+kOXxVLlkA
L4zqQ+/25UOf7Ixy8GbZNXsPfSYiowLrkRPOe/mmaHo5dTsJm/K6QgUh3x89tY+POsVagQqebjk5
6LrJ6iTdwFCLtU1MyTLerR+vQ2tJyTaUpajEa02U7JGZTFmKllueyq3QurLnNSc18lL+0jlEA6PM
74ZWIEorH8YRNiuB8sU7U/Wcq2O2dGtZ4P57vAZA/95h7BcPLeBZ8ygUx+WqAg3YYrFKaKy22nv7
ULbZymNDaIMf5x5nvyW9hbngQ3fzTFAYePzRgi4NAHrz/0tNpSqH6WNU8sR30wgOzaJmNMYqY7ul
6jyR/0jhqt/32qqly0AtdUOPL0Ehp5KkLY8C8Uj81ubZ5/IE2XeVhYsXyQ0a/v9WeOoaziVSs2ER
f4LeUogQm3Icl3jBYjtdMaCL8G/Esk6pYXx+vFpPoIrhOwg1KLV0GUKdAxst3SYUEZKr3daSNJuJ
OWvU16kkoFy5sv9+bfJ4oP74L3Fl1exS3phABdlhG3YjMLzqaKDYgNaqOxWI/lTxL4+JFkf0DAq3
u7O+CB+tyg9vD4Zt4rqcJ/FiPforES8mp/m+5iJPdf4Lj/BVBdZhoGJcKK6zs3uq5tXeUzEkJ+Hu
lWSYNc9M97GnO7OXYRm7fyg+HbKUcL2JRKUHVk/Z7hNScUMraMYsueRodC9CRgCxnC3vnTy/smjG
D1ukOXDkSw0BS9P2Ynh/TeM5PlisZXpOMqX14Mk+fgltmjHBX+gx1MDlBw0lUPtvJ31YGwMs3gEq
y7YDOgQG+Q6PbbrYGlExcHlFdtKUKZ44SNLPOlj3/WUwv+MIeY9Wf+VoFgyQ6mwH0VOcu7ExftaM
kMK4lxwl+EC/6Dr0MNWwKiDie9qVypTymT+4+PcaZDdb6n0Nn/qi3/5SASWMX25J2luVli/h0b58
QOSAd4VorUm9OXX0jg1x3kfTSfY85vl8G4SsRtuoKZ8I23iIj9BRdjfP4nXOICvycjw0jGwIwE/w
LyygCH5vQnc8CM/uIZ99Fhjw2w/WSzTT2QjxNLbkdI//TOq0MGxfnBZc+YP0dO+Xf1evUyzwlgqD
pkruIMh/DbkctCjsKjXBIVQ1ztcq+vxSL06Dta9m4Y20FPWobxJLpkfAE1DR1ZNCZhda+nPaqQoq
9VwCHu1RLMqdtCNc0186PVoVZ7tyPz1Vq8bqYtzrzIFBeoDhTxVh2hVG8NlQUY4qKRGiiv+DmW8g
q6gscp3bzAyJuGi4qU1TrlVfcWOF/0BdRI519KtkJ3EBJUhunhR6iSzs2UlyTfuwWxH9LFXXgfZV
Ve9o8n3XNG3dd6ExglfzvXdRfhbq+kdagnm0Y7qcHakKetBr4dWVOA97sPuKERiphttOo8e5KTEE
cAn7dOtzaQKq+ifnWeUEb/++ljQtgCeFRvOOqXLqmKD2q9mpZ0UJ9mk3TThiyuf02sX0MF1oHtsc
G6JWracyRDZWfMufpELNlHvvJtzgxEzL0tUYwKE8S0/nH5ThWNjQ7v6aRjLOkl7RlI6/qjVEecIM
rs9f+a+4ezJFh3i+21m+GFHOYIfMteARyJSprAEvZ0fv5tQt1aSSQPKAbpcHurKuUM/pNiIXx/O6
JC1W/pm/3NL5C5i5NQJxnU/ZYYRLzMr+HpWJa2HdebwudaG/fZqqn2TPzH23av8GUXaT08b6H0Ge
bX6o1fzDs9IJTNDFiVLUlWnVzRDEQh3G56XAMWnMccvC3uNCtO0m/9fL4BeeaiDK+PsNYDvb0c6V
Wr9ptRaoN/DmabIR0ckEHlNMvnFQHY7Qgn+nj5Wb8jVv8vYsrdnRMXpQoajVmZVFs6PhTFkzVIaP
3zkmUarfqVkeztcZMnb44t+2hYzp5T3XHA+HuioMIKnokfVflxjltlbAsr7jxJLdLv2FpqiKqpDV
WVzf1VZ1v2CxGlRnIJ3GsiLJ/i/XDIsxO2jkrs+JEcsFqReQi4tMOwS/CaSpKybA2gCUqhg5nHdh
SxaBUvbXBCeDGWgD2nIf+uW9Dr/uyaWmSyn4p8XKHUD9x1CUtC4eLt01fY3/uZTq65EPYv/7/DW5
Q30+3ditMXbH8yW5c/AAcCopM5N0ghAvapibBGKtmtLun697ZZ5IVvveWfw8fAVL+EMDOWrKqo0+
lFhd3ss92e+EYboFI3hI+ktgoK7UORX/L5bNZfeKS6PtNRb4+uWmbnRgaPQ5Sakk/D4jUyUZ5KF3
PcpGeLwvkef1oxU/yZTXCAvCIgKWr02qlL4m5hNwNN2LXE716hKNmjX2aHGfZIArZZreWCIgXLE6
VTNZjmiC9nZig8Hkv1IGomj26U5sb0owhz33zVDrQ19AuzrEIrOnkbYaagWSvyAkJQYB1sKsMDkK
l7L1eAjf5zdky9YCCIazlbgcWP30m5cvWF9YiVYxiIAHqjNxiBPeZ9pdgz19huo5N4YEUqnIpkuA
poAQO3BiPbU9p39rbWLKuRD8EtHfDkFz41XtbHoRs/58KgSc9sWFenEc3W0CNgnQ+s3zjwW9ABVY
6j04WwRVGarHyzFUdv/Aj/CeS3rtd6e03rhtf2vVFV1LZcKGqJgC+L22p9cBxEs/ayI6B/Q3DfSf
OdrnoHCN5EANjGE9rgVoW2ETm6zroIxXPa05iF4HmS4uQBPx1Le4XdsWphoKcJMYoOmE0selcsTy
Xr3PkkJThzI/tqrLgTtFhome4ipQ72W9EYrW7CTfWVvV6Tc6j8iI4uz6EjsdEXyPjafe0BNJr+8R
SG6zGqXuYBACL0KMisKGQhyZRH5UgVyuHbY67rUVqBLXuCxpr3+Csi8NEycPETXJiac6I6QEcuT1
bo9h8BVwZ0odIaVdWfjrVGAWCiokGVTucIdnCyAazKNYjGMyATM8Bu+xqdJJUNWyRq00x+DZXaPo
QWUaQabLdx6X25bpNWy+rglshLRJJlCrd083fY5XW99dv5870MNikG37W+phDz0sIxRmyVF6Rmp7
/wcHETh4suDxYQW3Pm5RX6cyH/uspdxf7NU2NqZn0Ot7RiJvAAlzJWD5eyb3KTp0tzn+HfgLQsNK
WF6Nvj6eVqkVVNzei076uhzTm8+5livJUIXhB3Q+kjvROzZlX83UIc2L0B59s0s0edb9ocbGynpn
5LTmQcDiXxIYPMAdzpzA8e8GlAadf8lximJgED90jW+3x3lZJL64F5xFoOCpygpu85zaNz4K9ghI
CFg+IFUBG1FfF02VIRUXJxX4JTmjwT6NKIlMX1CBYB+dKDdPKanKkZzS1OuqSj4ZdQnIki/F7ZA3
gdQqhzSzRh1D3xE5F++kuXTPec8RyZkv9hEIGE8xg2luicLkUmGKJGC0okcDAbxrHupWmUabz4/z
dFS/sJiMdR+3sUEkAqoAGvQD12LMVylkEOs6cw2ynH4lzZqUpAbMIeL8wteJ5peOWj99rUGlIEHS
qV7qrW15wLNafZOlc/t0MFIdNmyf5blGYkjpgVYHV1ct/T+WzjQyRNGmbXjEr/LIPVEwHKvH7iiq
nqPoTAW9ZHxgXBRSqab1SLSNPc7Le/KbELuigJQY07L9bqE69q5EL2pTj2RtZB3ibxNG//lr83+U
0GYaMeiY2zr6j17FSv4NpCPBTbud2hJl247HbwJ4pfFV5zUqeUfL2SvbufxD9bRwLH1kqAM1v/1c
suJ08kQynq7lg9J0DhHuv3AdKgGaAukZYQgny/MFoA2+d3ZSnUznAwCZhpPCPh21BUEICtpxoQ7N
f+iGXUCCT6ifQ+78xkanL1Bdr/J5hL470Z1jqxyblZQh10952NhMoSAqz3QzCMiu9cKed85JZiya
qa+nY8vBuX6NP+PXI/3hJ/XZWt+qksCJAbQHR3hr/H7MeNuTSOn0Co2mfUxHVtXKcoNZpxjO7SUU
bee8aOo41iHacwjK19NQwHoIbUiFnt2B4igGPWt3DrM4btXkxV8SPihwXOp3g4qVwOF9mmrw0Jas
yqEUo5HL5fq+0xn4FoHGUEZ6P5nLtri6XlidWPtu0edp4mrLgobfSESF8LhmT/YzqYbDqzmUx1eZ
i6rQ+2BLsBg/gnHgFOzjRT+yuGEPll29yvZlQsmjiLuErtIOSYCAm2smk2UVvomXi25cou4j7szw
RNa5ThSMAsCfE3+NNSeU9XYip5UWNS/GL+LOmbLTY+x4VkUCsCIyLEKqyxNLj29xnulqDUo9vzrJ
SY9Vg4ANZOQvGb8ZTbbudDrKsmnnpd+G9Yh0U6wEnWdreW0ecvkm1OkAgVKVFLOg+LlAnQWdwRwZ
Pnh3qZUvkUVEICR0eID58IUJ3zY/ZUtwaol7oKV6ba35/d+qKqD81NwhjKjss00pfBaLdVhIU08D
G30/gAhoy6YCw9n/m6E+LeuFSuyEzKGnIvvbUeJvkqFtVUbJ+Cf1tHqF8j7Yj1VFBiyFWCFB9zyu
DMbFC2IQgoGg6zLnVEm45CdbEcqV0Y2jFv5rponlfFTdTmWJiDFOpSqwg32HdTYq2BT4R5acCEbA
Ir2K+4DvYd1yV8cGYsAdl+fW9z+sh+z0yztWzP8hYj2VeSJVIZD1JMMXYy8IEImD5upqrY2a3fre
Rqgn+XfxUGS22CWfohlqesPSI2j1P8erKMTBuQY4QakwsjQ7F/FrfSF1mSP3sHvnAYwrcyEVcE7S
EURIzhgnLGVBQTxzIiKPaLBB7hXjBHmx+oRJfWDujrIHJLKGuTiiiiqqnD5XiDzzoQD80OvxH+B4
sfjBQxsayPxEgCH9lhUdPjE6RKz2yh6dklKBZKio1qerB057B4yoB0MWkjK27kMiDkIL1mygSWRz
kmTO9JiZLDxCf2jgIv0NA6oht7opblfVLvNNuczj/nXGMQa6+YFtYoYb1x8RU/RscK7GyXd8dyAd
aSKIlR/oDm2FlecZ/7hUIAZnYQDHtGjbPTUkqv04dwyOMKP3lGLaaQ1Sa5yoVdSX0wL8AejGkdGO
J2iDEAEveuwetpT247+8oFsiFkwECZaju6A570p6MouHUTXrYWO2uITrBsJPNDzV94T4Z7vtuDya
ONQj5JIZnbyz7qdwPrnygk1laJc30xXlRZXAmVcMR9K2D3LDWJVSyGuxAliRqIHfPRVRxHDoHmOt
HUeqHe3Hj23GZ9yhUWxBB0xAlOGWHtfnbFPEtCvNt8a9BN4Z/2eFKNZV7Wq9hOJvGF4z/S3BR9CP
ak+JfinhJV5KvMh+/sU/bJ93j1z+UW4UEbbF7OmiGoj4MwL8S0QVRk6yRO89r2BS2I6AsbtHWz71
tgZ3yOl998rAL3gksJJC8MPNDPCXDXIwobAGOo40jHMpsc2HuO8q4jo1i3yLofO9M8vBHPuxhtqR
ATHQHu+JQrMCTcIlxQTRjG8u/PKGnOj+pBdPRKfVwT1rgN0AkIMIkIGjUIlQSBncFMlCOWlXzhhd
1pB88r8YowEL9nfWCViCxb6CZzizVwyRJIL73M/pq2B0MfzmAvaQ9DAhUgzETE20UCxlGWKnGg21
VctGdSh5DLEVI0AsFUIvI7tSv1CQ9Vg6PV/PipVJoR21X5LoE2O1QP/i5GpzSISnVLOBsn17rkEP
Vb59K4RtIT0zjoHXrAMcwDlUMwhpFZmxrwtf+XDU0L7p6Bf8WuY803s4SVIGVc5YCskpX89AmLM9
zdJB4KUkXGhgkxQ88S8YYD+URA4iYae303zOcDBVQTuoX2kLPNhbL+oEvm+ERK0MwCS2Oks+eoVH
M6eH3C4m0LazdxG6U8EU6EBlxvIJDE5WENopg4sDJgtoumA+vTm/Mqum6D4oXT1EaE/tIDuMi8/p
qVU49e+eUni7+4ovzRLNHcbCp32rVeoPOz8x9a0z2l/EWBdO6TJ6qPpgcllold8QrrLgA1piT/TK
MFrCHiRPIblu/yUR160iAbmLzzWbEJMahiq1KpUDOI4yhK6ocEoLZky1+Brpw8i18CKRtpCRgjoY
QUrhBvLfsthzlt/gImActaMwoovHMWW+HIlHBMFpDkF5KgbKoqps6JWS6LbFJoZmtzW8xyk8zZwA
5EfiumrmULZXC3ik7t0KZevrYvzeZ6nO3hSjKG0Znv/oSXc7njOx7eLpJI4PGmdKM68Hu5U23eY5
B6Hlv5JRSpKCq15tyobvn1WuIw+PAUb07f6p3Cvc86IHJR6d1IkjqxPetkfSS07sORNVLNKuIkLv
A8dQAIGym9uocAGZraMivY1VzvnSkb6jg/v7WhLeETB+3ZY4tj9wobvClWCqIcJ1hOnqwsPMt7NS
3hiBu388XTow5bXxYHQ9CTmGfQ06Wh6Z6UKqIyPvlLjgOGttjyUC+PF3myxxdHFRYRkqo2bMe6L7
n+A2gz8XuMbuEganJmvbWaLmJZNYkfRLQJ6KNuHaUWrkTdQ0L9SpDME9n3KZXyy2JuZpqZr7Uv5t
T+7oItHu819SlnRdh19ot+fxmWUHmplt4gS0bACnuWQ7zSB5U3/zpoGVVPCgpkYE8r18Ecb0J2YZ
nXXN2tJhJ0YdNLvRadKV/kR+x8jrJ8wwpCzziISUMIrfuKxdBTCwKBu57JgAxPrLceo10KvYsD9h
ZymjuSzgeuSMeTBvuoM5+HpS0Vmj8NuTIWrsbO8YQgOCmYW8ouQwrMTcLfp+BxOl/VVWP+CY6bEu
7VnLRWUEtggil848jyxGc43eoOKS1EXD8cbjJRAUFoOKIxxW94oq0AFD7dnuxZ8kGiwYkzWdSGf4
P4deedfXbIMn0I/0u9S0o9Qi01My/6apSGsFOWvagBCnDdvfjNSAVuNDCWquVwjpTaWHP0iOC/y+
5STU//VjzBVQg9dDCuWZxcYLOUbyrOZqKnPOf0X/43C9eFkb5vUd4U9e0FF45ykMPAHPS4VYKEyD
ZYJSbM4L5o/7DfzWhp14gXEEmy+oU9L8xrwJ6317ZQ72nx/bOJxiTNki4f2J0XYIAxoyQTdVamby
fDXIHUyQJ4SirxJJeXU2l90GCl45nCfJMhkPHdbdXMVbflHcZyBO1BBe9bkhhy9MAbxnIf5Vd4o1
Ck7yeyPGOj8l4dS9jmOwPNygWbRHHbJcYmpZPwmv/N1OKTSiO5g8UCasgdwHhlXXBdBELjN5Bpd1
Wt5jsFAcbRdUVwPmNO3bxUPJ2vXsH5x4olwx8OHqwt2rgsdz1vTamTF8CXqkf+IrO4XcgVGILaYj
qneN18pXoMJ4FmKqZoC7lhH8KJxt/8Q3yKW1n15F4vifYTSYVTpxg5XXDodBcjfR+N6grnQENL+8
DDpUcgToXrCB3J+pHTRXowTY3z+J+Q8sho4q8OqO9MgoA8ObGcoo5QHQc/3ZLfT8VdfN8AzrBIaA
3dxBo7WV9TAOY5BFek4xfoD882opTO1JY4hIB0PVpdXrHBhn1ZTl17nJMHwrVu+bko1MqpPmWUcJ
LKZ/5tYW2/zwDkQqhN+90N/i+Jo7rerjHaQ7W6iAtHxsnDy9drEBRjEdhYyZc9BMWzRdqb+2ys7Y
ZMqToHTo7hKY52FWFLpUz5Z0+KkiDeb9U9mrZDyDUBmj44xljzBYnGRrGylutkbwHIprDzkyTEoN
4/8JyzvLDa05ezF/XK+hsSHIDLhJoceYzjwgRMgGbQhAlMA5i03IS5jUDpBbfJzWS6U6o5tT7owA
Cc6Gy4ABj65KOoFMKCcTbMMOZoR5rVeUCricJ1adSmqEN8i/dkbXnZw/nGRyy8inE7tGLtCd34bI
Dv1D0S7SDSDCso+wPe+5MlRCSTyl5Uw4fDfQKEjWyYzteY+RJ19faOEuHtvHwp00hFBbLIky6Mbv
b1VwyfiXGhG/1ap0OYkBM525inUfZCSae12uGi/MPzSaSoE65SGDgiAJreW8LUWTsA6LZy5DI4RR
DN60oMK4zkPCIbDXSKh7yR4Nat7avDBQ9zK7fzwmfUbbn28Bq+JvyIK4wXmpr3vrOMBmsZc23XHs
dOQ2j3E+AcL5BEVpY++1ExOEGfZPiIa27YHj4zbzmIt7t0FiRhnHIjpwx42T/mqXJb/eNCzGo4zw
nIGcF8Y65RUMlFfgkkAA0NxznkB3ZiRHYRr5R8M2uHt+8g8xD6tP/edMJhjClYTWwew55PWlLCPY
RlhDnM5LmESD55XKeTUunMi2bHOLyGap5igkveLSUG9VeE/u8Z4dueSfnuQwjBKIJqxb0bEHVBFj
rX/1A6X2QehwAOWIQG68eYAScKzAb70K/N9fB9LNqXyPJdph958SmLW8644GnWAN0h6lmGbY2mq/
mq5BtuOuDRS/HRB8qScpkCcWVcJg2+wfU2XgVzZCIHzQnH7o7/BpJ8wmI+Owihda74h4XUvGZe+1
5Du+aOa3kIxBsRZqPiBRE37MOGvZl+WSoxZmqgQE+L6VZndKkt0LagIdicl5tL3yLuA3sBK6L5Ld
qu3M+7UYhQ8QnJiLodph5LHTwXjJVKtllxdgxMrzBZc3cUfsINlBsk0uFv7OVKzXVYusbZSnYdIg
nX0RQQDXJrlOov3m5cIq2BYHytBS0P0x0nmVf/E5v99pTIBLTn/EgArJM/LBhum8qZi9OLpOWP0g
TX4n6Z1rqwL7fRZHE0Z1zceA+2Jxmt5UunaF+vwQhd5/uzqnTvoGdGaxMdi7iEtBNybzJc2AmwHt
PqaixLDu4pJZoE90+SVt/tyWss7g1VNM8uFHZhAZgYrpXzz+EMig+tFwECm2SYCNACbMRFK+Rfif
deO03pWXZPCwGOzESiumNSqEe6Xsof4EyxjgtOPk2g3svFXnfqiOnh8YXiulwcdZegXYkC4etLcA
EXP80Ic42etHhHwAfsuuqx0Kpxwn/9CNFiJh59Wp3zxgJmb9NLXMpQ1eYa5gJCB31Oo8A4xbwGkh
polvfel3T64GoFozdw6EUSdZuUIDmXPECPijTRvPxzaifaL4gIM/PoTjSEl3gWtzNTsit6pchSqt
Q7NOHOaqgBQehbRe4jil6uFleY/C5inRoO1vnwZDw10SapVRN4d3VgDw1K/mI3FXczeuDLKmE4uo
oOK54s6c18l97rxb8ZFB0VNXt5pcihmqKk2UkUjg1GafiCrcK7DpzxmnRd/qpg4sDpVPMCOpRNVG
OrGTkvp5tjHDlhIYCN1R56NH7a+2IeeWySh16McAX/bk49CYg4ViKhHYDuR6zFkE4ZZxYdk5+MvJ
14iqqm4n4aNgQ0RPHmxKVvpJHGfvhjQ12k4OSjde8N3rjWdjhrT9bpiqFovF461hSpRU1FH83xHF
1at7gda/l3EiUJzjNJVsDyv5sL7PmLpESQKimf1sFOXtUWUYSy1w/0AqXGlYOPDHE1O8+FO9D0Cc
fvOzZZYisSmcV3xw3BuwKlX8x+aSd5SCtC13iKRXNMcnr78puTXTO96oCNWvIXGEXUsVPm6x0a/Q
VWTGEVEatpcKOCZkmuAQGycazqN3xezjvE8buBdHBZrRgGiBPecBocu2DngVeytLxzaT181tVz+y
S/af8Px7Yl9otaCov25Mn9VdM+5IN3kU/9KXpcLsOM6hQyxzea5jZxggfHcGV5jfTHuNmwzku14f
W0UNt3pmIb+j8zFMvNpRNjifPpkKapkMy7q7jRRLp0hIHzJj3OYV9qrLznhrcYpZpxMCvbs1LgaG
mkqROnnUAZp88aGcWRw4kxJFTkkvl9A64y+aXTPyUKroaDVFeEvagYtAksEV6Bn+IWQc025HkV3D
4Kwz/ZiMDcYzDrRE/mknTRVtcVtBioGyKl0U9H6Xlpwl8vocsHmA5DeYY3Gj23VAK2MAEZ2cz/nW
EZu/dMnX2yWmoNH343kaPBi77AioGG+jhMedvL/sXGCoBv481RG0EisFL/1CFPVogaeXEZiqhUCS
d7IqQnk/5tfxJmg+vpvuF7dwToN19x66TV8rwOTgCzXATb+xHfyYbnvKujwx8hnf6eXvMTvfynp+
8YEyuVaZRsdZV2l5pvgFxA1v58MMD0eVvDm0PsslrbQT9AYlAlLmFcV/OEPzAOeWZvk9pGxfkeYQ
+R1Bhfb907SQN8I+xHKrbewt/G41Sko5NaBssqZ1aQtXaRI1VBX+9ohewgcCnCv+BYAv0w6cVOEd
QSLLhRQL58ZB4KNj/8IUGQCMqW9Ju8/PTUvF3w+EiJFGmVET2Z41NPHLckQWRXMqXtc3PYjVuvhi
UHcX7ixWCyifandG5TfC+xsr0AUwFZx8YBFfS53rhPQfdrA6FTfcez5Sggy/wURx+aNjzNFTQB26
O1izmc1ZerDUTGEMg99Cnx9nktgEmfP4/fDdO3t9W0G5wsM56uFlot9MMEoJOCDIdZCO/UwSff5y
H7yCx0jMGtBxyYyPwQTSxHOGtTFMo54c/HNKoVqsn2ofjxznFuLJA+tS3HwRpNyXCyUBSeq+NvBq
np7L9dgHspSnE3g7a+hBxBt7RU0/gLn79LX4tf1KLUmNwI1PyQbL0mmoIygAOtLnELRUoklLn02T
Etmj94Qj9PFwyERxxOJNaGT2ehuRoxV6PIQWmQdoUCKvGAN65zYTuk4gMjW4goXRdN05qUeUllC5
kuvjMV/6cQ7s3yIELlsAjTPW595S1vs0rqTazIXz0zrl5JfeMMKj+dSb3cVyyEvlGzpuWtaNIb88
Ekss6Z5FNQdlpKuBvy1kPWxqt/DRxqxd6GQXcLj9UCojq66ccYcO7yMAVxPvl4i3JDj53p2RLY8/
dWEEIK2BTwUcVZzJlghEGorWlClqlqN6Q6w9dWFVv1CNPeTLZP34TBOoQvmsmj3DrF4oHKHcpBAV
hgD5LxeicUN/x1Zq3WdK3KHwVrcmCPGVvBCdx9U2CDZ8ChcbusA3AjWXvB5xW3Tx7PEZtUvIQzDH
0hG1I3tCWwt1AjSDMaocRsnTcO/euChBzj7WI9Vt18WIoKRjZ2JqGI5lGitk4ul+gDt/MspSn0zf
wsakHhlE6Hmt0ntq9aT9xNzmqtaKozpcMHpo8ZuJkQ6MjaOQVsOkBy4FZX1PFNbrSc6QXhZwgV9O
xV3F7khVJAIOrNJBWWj8r75CxLrnCb+sZSRQtFRbcKUa1cmRkLDNqjwBidRpIh0YdFekZpaNFvKl
tW6uctMjQFoYTn3xNqSkPKKNMT+nkshaFGw6xEIiOhzODT38ABa+HUx6JUL4bMQbdJ8RJD9MjS9w
a1xT8ZLRMXxI1XLvYAVREB+sKbkc16L0VdKROMkYYNFSVdaax2+eB+/v+0yUstprSavTraChwI+U
aw8X0gyQPBUG3Fyp3/iFlTrDHX061mUh0KED7Zo8qgZNEGNEz7YQPiXChuxJh1W71RM9ez7lS+dH
oZkLZ6KyyPxvjeBEVughFXX5LU/eDFfyIen8GbS8gN8010qssjZ1VpWc8dzZtX50AoX1/b/dWCI6
G1N7qXpMmuRMuKqdVrNz4iIsOq+WU7xbUxGoCro/bvWTm6TF/3brSr+ucCC8ydMG0ivsMnN3Eji1
qNVhYRmuqF1jZ1i+yJKSU8G0le5d5UxofHizHxY0cfn+Tn2ZgZP9PPHeBNGpRZrozKiIymhcC9FC
qdvtYarc2S0v5Xd7wGkkfcNpsctCO81zBYLRsGtwD1Vyu1R1qqLqDRZJp6eDwRvEtGeuIb+4wNpG
E10vvuB0OtIbm8pfDkIYd0QKjjkl7NNBZrXBPnYAhc0w3lYH5pWJ9gLF14henv2XnYad79xkPT8C
aS8JKauX2y+UwoolEsRBRNTXUx5EHjCI57emBi2EF4HmMXegYLMy7GDCdLHQ+rEGRyNHcftfCijr
hW84hztKuIqGZnIqd3ho+rrwBPJ6VrIOub4ebNECYNJLCmtQeFqrUkbh4nfZg+GTRr4MoUGPm5YX
si79fkN9GfkH+xg4mU+qYZchayQaXQEswXqemszvaY/eNxj7FUCnmCM/VSHr5kew4JJ+yntLtEGA
Fa/pQY6BHwvas4qL2OlrdBmAgdmiCiWMQU9Q7z2uz7leDWsU5aTMleBmVoecqKTeMjdAeE0Zf5Cl
Me0mvCCTg3OG7xiqAO5GVkSND8PfAdvq/1cPC6Pv1pVzmMwVy6OS7LLMNqC8MujD7LthILDZln5X
JzznWHTQT6Fmn1ePj/3dsRt0IyEsrOAY8av91mck89DARkE+4petXQpcWAxhYc/N0yXYypl5dHKL
9MS9vfBlqDuRoobIEz9gdumAIJpyHFHfr0bQlsBjKjLds6ZZ9V6RtVLnNAujPbQ0qzsUpOR3F9nk
MHPcrZaAULHOqXXXbFmyUAswkI664ZLe63eJdTZ1M2P+AwBUhagvfRz6W0SNsMq8NiCkTLDBiNaa
1vRu2iV4hO/hxdYGzmQGUsw68fVO4qaL0gVPIySVlnnDifKW+VWE64MIiMaTDcJvnMqUwfSk6eZg
ib4vDXbqaF2+rfglTnjshYFdndPQuJ5/E0f77keLd+MdEophFpoMvmamAQ9P8vUTSh5MzjTOEO9z
NELo/lqA298BfftwwQUv1tMsjr9LhhRXKjZpb0FIUNRhD5LZQcrRYjozuGA3LABgjau+0sFJ+EvS
FM3v5JpetzjTETx85NihvLTi2CtmIpJPqSG5ZenMXBnNvhB28A7iIy3vVvy633xRaVsM++gXwyNV
Mur/n9AIZWQSzrD2qbcB8T3s2FG9Ir//sXCVCu+HsQ2+/rUiBVD2yNITAPujkkh4kC29AlZwZ9oy
A9IrIKj7VXOxqOTDYVbGKWyefImsypxCVHDfwB56vL6eQwyH90WJkY+wCgVnVrHnI9QEkd7UkjIj
5cCLNGnvwTOZifDl71VYtpYeLiOA9Cy3GUfVFdgeMbUVHL8gcqChRpAqcH97Z6nYZjB/o5mkbl1E
zxNm1A48LRDncbIZQFGqhXHJ0pSY9pxC//q00nrTDNW0aCwky+9dgZWS+UD75cDefwYooLu5rtPt
qz7ZyNU9Q1UPvpEzSdNk7Ee+euIct1voGHsx8UVijFxvbpv/aLrcIwhT2E3qddFWwo89sIWW5JaT
UodHuoShBTAQ54x5ORQHasova0nnIs+xQc8Dl6qldAzsHf0aBX6/U3gvrtFmsnHqk3VdqqQdqhmh
foocUc5eXDcMzIuXpsXu8bsx5aKQRDLmG4AJyxeNvhdKHn9SO+6tEw9kIm0TBVPhZUE0HG2smTf2
iGrKiUBjjXuOCR48iKXmvDWTK4yISZBvovwH2CgpcWs10iXKUiePO4u1y88rEz3XUVg8Hv0+ONOJ
oVyc9Lew0wvGbfPI1DzbrfngmOb//oidmyU/2S+b95+/T2i6AI45lCLS4gV05XbRfK8xBFgFHBz3
uU92fMRr6KsAj+oJjRLzSIzYZe6uulk1IT+xF9f+ekx9SDUOF1BW2P7nl9VOxjpRt/lUPcsM7+By
haOatnT8WLgGHIPk/P5qHDGXTcLOdJrc44+SwzH0vzAeo8gxLrpInbmvHLINsBHYzdgxXsTj8h9O
FL1orpjrN7eYzGDUOvUcqEELDKOEGbTcTYJSx6oZ3SEfnWdKCO/tCieHMuh5srBvKS6kyRgVFOAI
sooEki0q05AGMl6T508KFJvvJCYvdtdAp3q4Sowbs847+ybqfWU/jAf+tfVIfXf5gPg/KXxjl8sO
S3wkv/EemNIVLQJ5Lu5H1v2t3eeMseLyku8O/rByJj/SgZ7QL/jt5lkpQiNOeb7Bh2leg5O8kCHr
p8pDz+VEY16C3pGEhSMTdMT0AgKp9GvKhZq2ckPzAJP5tGo7EsBjB7LHei2Qe1fBXYV5E7eFdeZc
zXouK6/RYkWzDfCR9a6Gb0pLTq2V/4yd67hZsxLy4rTxPjxmWR0SGTPcnOtrCfsrGmho+UnixbY4
iI3rWxoQsaDQU903efWeEpywOYHeOF3MKT8Ff9dTrw7+MJBUta+rZG0fz4QVEeCDrxui6c8dTGgq
KsP9NA61dDMNmYWkWY0N0fj89TNh8LCx9UFaJZetHYpRQ2yf7rRES0Y3XAh1v4mt7GL39uTx57T4
oHtD2jb/AUb4/BWrqYjvgE+f6RXql4eOqkeZcEtEFhgHCWtL0EVvhSQXkd0fEvgCWRw6Abg/B0nG
v9rPbWMBrJAc6YFmi9YGNPDYKmey5yq2AplHndUXpSyFNIQFTud5eX8E4dXWS8SbvvNhYL7IEJAI
77QI6K2C3AhHPUQrxckPveeTdCrjRNJo7Ryr3OdP9QjG0PJrtILFOKmQHPumRauCSB6inqd2q6hG
XDCCJcjqPZuuUo5Fux3V7EQbWOAOFp2KNfehr9UJfsiFAGbB8x17kTuB3RbWKeMbdOz7+oUBv1dC
tanqwEbXSELmy7+r1jcUO2srWyWKkPaI1c3tbRaAGKy9a4koa1QLCcXh0VRtn2dI/vu2/qBl/mxL
AiNK0FIMaNLcTVWxNS0e9DA/OkU33itvT5zpTiyGYbd4nFpw1haqX+jDioiYDFOlIthMJGHNzBXJ
xAk2kfrIic4CwE0I3a2oJiuMW6zY613adb4eHv+nSFNc0LsTH6IW3YPXe0N5cQUSi3H49EMek6w7
9DPUue/ZtPss/KsmwcW5Cm46MhZmR2aPw9KZKxtL8WZoWzYOdBOWFu1OF4Yh0o4Mo5CRMXb+TjXR
w5J1lvkipxHWObdKmlTwYDklaLQtV8rgRer09KgHKL0mZ58Gu7YJHb2MG+lWs9UJwMS/XF+QdqUN
Ws64fyGp0sCKtLsVMn8AATCRbxrTYSOxf0VAthsnQ2QVY/zWa5N4xX5q+ibASliTbegVXB3vDXCl
tLg/ihUS0CMsqs1dwYI8X5Izs40FlBe/SkDquswUkmZ2NCx85qkWfULjNASAsOSNN6OU5kBTrwU4
QNZdbag9QlD+qPbrN/XeYzqNoqMejw/KlceO3kCKOezC79KDuQRb+QVpET/dL62RWs6cMIOInfj1
X7u6iCdtX+MEhAqJ2Mm1iSKfoGy9RrhPHqCxmnWNnf7wjvxFaCghKKzJJZxaHHrOyIVPURfiOQ4I
0rqPaDaXrYs/JFG4Oqvv1a5LsR7fsMgfIW/PJRnDVEKZBmbv8VCZ68jaLz3nkCgxqp7MNGQHoaY3
JlMfGdNrwlY5I2T/dbkXWRAbZEc2Z2XnVLAXGGG6Tohv85t133Xa14dlRcjIQT1NA+5JRwT/Zwp+
J+QqiEh7WP8px5rGae5Z8oiKK5O2ttLrmWZIUanLLuIFb9oDdnGdcnarsUk2lIDH1UW5UK6dnqTc
hcYIzPDFKQOeaU5TP59qsmfLthj03NErtO069aWSSlmuwtNC2Rc/H72Xl85oy5DwsAzFs/ZNMjWx
wyyGbnpeS64dZUdAh4l8a9t7qjjlzRzUxQFbYn+dfuCxr2+I1CTS9FsHdxD950AF9S3f62iGpTRx
DRXDA/SpKQVyxV8aMkouILuHwt8Pqputpaz+1NxS/FzPwZ0KJ7qoEqf+/KNJN+oLG6Au5ORKeXcF
T5g8QjO3j1Tk0QqfJAfF5fg3zrTNJ6hzOsBBiVsvW9ZiPi9jLSY2fZHgSxJePnJ2gybtl6eV44F/
LhP7rufpEFARCJVib9dQutQegiUXwSwN7sAGliFaYVoD2n16QWhJKoY4RSOkTjp88y5Zq4iz3hog
Bq0SL2UfzMAy/jUHXAWBK3yJFolz/sQmKPmIw5ydL3ba9U8ZXo6nHKlcw2fxh3UNTXA4P8BJfUJO
yyd5Kal+1JeY81EuCpMwFYB05YvAvJDCSEPN/wY6SDqYXDmAmMfTogIF+PtW2ju3/HnWkDaW7dpK
R2uKCrhpUB22wUjlrMjxy2aU6Ryqg1ZekBEtyeqTK9IeKFnjur2+YXavAp7RkdwbeOoukY8heAHG
NsWBW6sgLbi+y1YNTW+ZOa8FgO75FTV1Ap+YPi871yh/KD/G0TCwD7d3QzCFAy+pQZHNS8gHApFF
NgsjI2HlUQ0WnuIXh+golaU7hCer/Vrq+VIn49uXf7h2PQwrf1unW+jVE36F26TSRJSZ0Gti0+CI
xH6vkebrHevlZlKWX5HccLq2Eq1Vsz9Z/UTsTSRItZjrENQ/kdPPbCTLmIQYruZRPJZZ2jLRSpXh
oPM4RHMRFDVIIgPv42KCuvRNQ0WWgcReHdEHILrgOOx2LsRi3QzZriBYRxQUU822N0WymwZ/LeNa
QOP5Nvsipj0OS74zmJ+rvCkHDBmu8+7HY2iXCaP12RthHGvKSVq8UvDyvLJ/dUnqnyxIlSnavDNn
J0+CaQQivVzl1DPzrR+fiAOLii/YbIbRivNXAodPi0BF58SJJYq1ygWMlI8hezcPnuIir8n+61nT
Nfk7pwTpR+QKAqCRF4tcy4SIxA9mIsDQXaiKEDnGqq1kkvopq4k11utyXM7ku0v4oYYIbFw7WlhA
8ZpjNcMAUTuCg/Kbjsd3h2fXq1lG2GrAeZ/NCczVUHX1OXs05GEqBHcBAw7vJnoAm0d0ZUr+LC9k
zbUilYXxqepnCCBqqDXMCGEz/dhqNO1pOfgziMaOGsXhAspFtp9n7Wv7mMX9qjWF6PLMWE/l0PP6
+trRqGcdu9D5RwoFSXuFazIdUL2UDKnhOoWa4MngxHtLxtg/NBH91PuLH2Cfdlyg4rEPjgrbHYTq
B9KgXTzF0kkQNRNG/d1W5ZH/9VLhp+h0vTI2q4IYz5uAxsyM3wbuaVSLH3sqjEFZ9yFr+9wLm2aJ
WDfTMe44LQncdIZfBDvv3Wo9Rsjx0t9uCjfacRjg39DLalG/cXRcmjGWJlUiO3BypO2NAjtO/ZEV
/+cFFubrKXWsx+0VMWo2UIjMmyS8g0KIcFUl74ulYcSQ98Z1lNOeZ05clhklKOFyKUM64Y3ux5QV
ccx2OSd7r2PSC6cmfgRakGNNjPTxinIB+kUqMrIcTawXjDnLOHLyE/MXe2RR3fWa9YOFIMKQZGDK
MCfhQzO2bKvKqlNaVSJRQY3XmN5mCQEovpgrOLDq3VRX7DDEmwUWL359ite8PVHfEgAMooYA05ot
Ea2EC6Or0I4SuCmda4/xEBwXBKSnja1Oomznr2Cek9jPeuaMWM7siw6LiiYAeK+6EiyJI6QkDA/i
ZbcMl2dqZz4jhjSO7K26feX4Y8m8jhUoSPSUUh+xYyIgPjnsgWM09t5EJyNXIlL+o+OIRwcuePW5
DelwgAN65yj+nhJ+8dxI/0/uDYtC16Un/f9INH8FtrKdkdsSEowF9o7TKet40ecLOwALxpjwN7gl
BB1vuzytlDGJZIUh2Jx89V2jbVmialYoOuQfBgGDA9uZfUav7ud0W0xZZ5rOhVSv2AUKVlCZdw39
qRrZ6tD+QvMOrPrgtqGmJZgOOXppFvt22vMtJhS9jWoJDRcRKPj/AQ8CuM9OfCsIa8oRTK5/M9sk
cdO7TN+S8JxkGXwoMB+9Va9n3pcSYdbM3nN6kAg4OOQTJgq+P8+X8TpL0HSeAfYSSFIYwcACV73b
2pP36xts08SRH+Rcly7kN/pH1LltQ+GUBQH2WXfPEeuOdFwmOypseYFyAFlp6vzLlxugoXsb0nQg
hleUmcf5imxhbIoCT7L4JbEq9BzI4g2JQIHYeaVv80XbeL4Ao29edyUw7mOq+rcZJ8LvDNB5/43C
mj/m6TjNM7/myz2h54G8sYnKaTjEWNoTsTAwAXMwZNk/x54NTfheV4ZmDsR0TG0CqoTg9JcPfmbE
WQhXdkyDUgEl15Tb02txVxScAQgp2WAXVxhecESgJ9awupSexuxaKoC8kMliPwFOvHIma32zprMv
gUy2MFIXaZFwVAAb00GIo83U9zxTF5RkZj+2t4Q/S/zTIRwuObdZGGk6Ie3l6CuDRNlrRzENL1My
EI/EuB2yu+Zav1epCVFS3vHCUNlkKDf0SdoWNU/9rwV+ZxQ+eYDEh6vl4czWw2w0eRgls7YgJFko
K1Mf7lVGzg76n5H2zNwLhtF14ksnKLYwen7gerhXYyA2GWvA2oSlsxY8TAxj69ve0tuwpcnXN8n9
eV2HK8eLl3PwlLaG9LwT3B5Gmrp36Scmb3Aa5xwuAxAeHCo/kRLCPoCsQ8iZ/gxVnhdQmAnluScM
e9YEqZ+FxPvHuUeHCwCfPneRA9wLNIrls+1JZXPMWx+FVCeuo1/eZccQt9m7k59FMEvQAAsIeJgT
WJL0HE2x5xitOqrgDokzEN57FfOL0pE8e6khtQt/lH/ajBYU8lxQyNEnb9EIkAbWxH1cLDR2NYUG
18b/hid40VybNh0x9JTr9gHzNUEFm5n5CHyTai87ebSQZ+StqtiFoYXUOyBh5Czew+1k+kKdBO5L
r4NsPjGcMBwPujYhM2ZkZ//9NX1KuqsoHJtLsgoJy0hr5SHKTrZja5t4n2ehWfK5KRAhj8m7ZF5q
+fXe1mzj73f0TYO8hVUm7XQ5Sje1ZQW7XqE1zQg0V6c6TxuZEOb8Qf6chK7ondYqZO0f8FbnPmHH
C1GhFCHbVLXsoG+thhdnW9HjDnjQAP9tDyU7oZkkjf/GVK+ThdL8fx8aBW9NACfDvFKMVdE+/0UH
ipQf0bDDJANtH+49uS88iiguzTHUm4WST4VoHEuCXx/cXx/vYx8duND7LdyKOx6SjxXUJnIp+19q
08ZN+CwtXt5y/yVqwL85FfOhH2dXLLoP4mQhsQk3Y3MtJyUek5Us3y9lb65ccpQSjY3k97EMJVwg
cmbDx9ro2ue8lOrSvnYznL990qLCKBzCuRS0tdNUqbIrbg9f0S1V6HGxMC5KNGztfcT/QMWaRHj6
FgPGfWHtGWA9U24mhg4NYTuqSQ8D38MMsQItlecPuBDUMVekBnCO+kuV8go9fNNLe6vgJ1BVb/Im
RoK8hN1ETdPpFabmpNqJJjdJbuFteFu/gCcNvuM4UDrJcPri4HClKWhwNA8EWBDHCw25HVh9mbU2
jfuvZnqO6G+RUodUMFXeiJn1gqug3ps7pt5xZYSQAuIqb4uYIjjCGpxy7k638DU+ws79o7VgoFDN
hG5jyQEsSWapK7Rg8Qju52niuMdZ8KLod8y10JCVC0dZTkq/xd2MihQJC+tJmzfwYzwkn2bGRa97
+yVxTVVJwkm878dcZNwQVKqJMqAc0VkJ3ZWr6F21cSL25VJrF+TmIBQBgwXmwsjW7EX+aHyHkomv
u9v2bPKU+OUMi/ozbZudOPptoGMGSvkhoXY4D18AiRoczo3IgnxOJ38iysAKHyBRWhyA8GHbcOXn
QxzkbZN0+a2Th+2MPV4eClPoG0W9fjpMe1+mSO4mmNKY1HqFGkfg3jjhtRDl+BCOBJvuyiNH/cfa
mOUMRL6I7AOiPHyxsu7Yz8tCfBcG791WHAcdofIb0iyJmiBs29lc342xW28aDcNllC5DMrsvOK+f
6NgrER0UJpk+Q/rgyTPjtPDQGIctK6glIjbK6SzPWZMnwfDmWBLp36YnUPcKUz+yhGPcu6nf9uEd
T03wkCgaL3YoxOTtOGdOiSsvT2UpI5tJbtInKFVxchdJTV0kgVRw8VLxwx/SnK8HV4vPPSDxSZd7
D2Cpi92tTqhCWiYh3GUZgNn9zPtk5p9jIA0ixqLWXvUHN8/kpchgDvteqacMSnBmUzTL1KJk3sKz
FUVP84DNpGqxoV+9MjEmxlbrXQ8P9sTeHulW8Aly1LmVVlcwjqatgjci8TA1kAVzT327gb7oMBNb
DdVAIiR+34Kv6kkcx+OmTO+bPVclshMu0m1QggpaKPsCYoyUmOba3FoLMdTfqDpM3MpRULvdPpVM
jFKG953CYlIVcPYDf1D6/SK+MRNaibL4xGwjoGWl8JGVT82N3kokdb9TsKhpVXCJbx8qksWQB5hl
D8XcVbpWDjlh+f1hC9S7CH/d7jBF5jXXc3zENfZ/774RvpepErv5q/qQ9bPYOZEYu8nD2kPeic2v
JGA2iKdLMjQ9KBZnFB5Obe9IKYkcTkC/VKI9xd3Z05l/72RfXGKPufvLu7kYoGZM7hCYyAZZzHxH
yArNe/BKatlrKv0g6DtGpT33BcRPvtCcrlXZpnWX+hOyyfSluGft0uF+m8Kl2WcTo0OLj4KSP7i9
w0xKP9lYs5r/AvmSlkANbtnvs1y2NjH5vTtHVBnIC+AbDhR+35WW5VMrxfCPZzNzdvstdRvCxzLR
UUl5evo33Vir/HWU1EPOdGVaWRHnudNlhNOSuApLDG/xnpSogzaT/5cClx766d/o0kp5foYLgUoH
FmKU8t70JTG031bH+hMdPFT3ies1rVdz66ofCm2dod/3JpbDorLXoi1c62PrkRX6kpBRComTOtwR
hr4baedvMEbtFsjGRfr/X+WReT3LVWXdYH3mZmgm+la7TLyVves+rupCVY9T/ExLaPp2R7wm2aT2
yO2f94gM9/Uei91aEgiBOJoEdbJnytsJ7XubZ1K1I5neOdUmP7FVgSA12cvNu+Dc9qkTpFzArlpX
z+X/WYX8H25LORHwveApvhasRPQWa1euxyB/FEhgZa/Qz5OoCpGBo+rhfFqrAdiOki3qIOHSOMek
Wt1Wd/4MvRY1WUMS0m1crPe/UalH1ncIUvkvR0Of3x4540P2mVxMvff4vu/BpyhOsYkeQ+UtQlSn
GP7c0AWyVFWsa5+lYEGcPRQIXl0EL+BSf6fHRpiMlsQv5eCq3WYcZga9Xv/k3ZbwbAiUON6vS4xZ
h6yGt6rCqarGz1+4Igw0ikbNmrnED4o4jtfsk63NrpezFkpR/zSBTJcdqoWW6famxfFx9BlPe10d
PGpnZU5N1RpAQ0we19379K34ogwAEaaqZZFRhjErThizjg99lFnz13yqIrOGgUArnkQocpqERVap
OYW3pEAGnB7x6xiMwxEMiFasvHE10TnETKarENwJGtFrR5Qdt3XRfLDWl6ISNzvo8z7EhMMi6t35
/HRM1mGmATmKxO8rKhqwzIfK2NIipwqFAnuv6RFq4+aG0HH5z1H803ldikUnNN4VRYVNn/wEuOHf
TTSbm66Tm9kH3mYObgeUoFiS0ksi9vrdder9f+HCxpga4Mg9Q44SsI9ndWsUGc6dCSF8JrgzNESi
2c99dd0ZgfjLuHiTQGir/W9C6sLH8eB7KmnFUKl9hRxbLOylmNHdkEddiT9VcYpqA23jLNUDd1iO
db3GErVLXINYc4jq+cqp3bH2i/XupZH1vFG7UWJijip3M5Ipw3nNrTMcnY8YOBY/tmjjo4QrCzwk
JrUUIhBaFNdKAgd3O0bve2PXu8HoI5IuD9mtfZTLKZO4mysGdoeqyjR2QJm2rpjgvYx6j1OeuGYE
5N9NyaJqfazW0p/iNO0TM7vVfEoGjNceCTBGmKGe4r+8lNNhfSsJrYAK92AIpvXKCh68TrpQMJuh
NZFap/34qukMqQ+2bk5jNRdGr0iIFL9s9ghq6zSqUVzlgru4dCkzC0ofcmj9hD9mpVa7B8usmQkM
ermfDJ91/ixPOe6kavI1Je0hOcbsqNUCjJ7uCh6NNBNlIxKOEokRykEkz/DDiBnMcGN9bgXffbA0
GE5MXPo1Q4HpESZ+ietLZIMlGiFnb/LkLrc1dT03xuuYBwW/1l8mPusASSNxuheIb6ctyfTSXMVF
h9lq3i9xZs4Yd0oL2H0glBZ+Nzb0lYLX0khtyO89MsD1XXImtSRxSpOG4c9NhOsw+Bjxr3Ra9fW3
HUK/8HbdhP1KJ7SYtllbIog2ZkZ3SmXHvICJn7DdSqnRn8EDQf2MFCbUHAoi/Mb9vL0Vxnz3Z83R
gMO0uyrS6CMJ0dvedNU8l74qKSMEAoNVo5+ZoGmp89B3rEvC2dY2RMaAZeI2ArHNnOZgmBZNOPXz
1wzOhRcCIDMvDTFp1Gj9XzmceLZJuYFOZyPWH/YTCOzbj9uEJIaMWX6ZLR2m5aDzGjcHI6peupPW
Sy+IFCHY1TAAC0AdgX4LymsRRiZmIeuiifDdc6E0D18pwKFhBfmelONzao3i4gZFFJ9R2WkBFhwv
MTMK9qcRVFAe8yusMLCG2c1iEZv3XqhDDk3qqunI+2BXpQW+l6tCRJdOqSBgb5sJrYhpJ2sEGrJe
Z/EZT8EggbcBUvCM5rA4SdY7oVD5sQSioFYN1lYV0SAK7YWKcRgbpg0DTtCqqw7KdBiSrDluBFyZ
LlR4AwYSoAWbAIN7FqF8srb6jnaurAl3KKkw5QN5nB4G6kOPwCgq2IyGnWkHI2R7zGZgDEYL2/TC
EEA5UZhYhl6aCY8Y8qZKl2J7HOrzqGTIzsq2bqyO7nvKFj0KFq6bExwcRVmbi4WvF6I3Y4SGBKT/
A9STiZQpBld99Y8jcz9D3w6BFhOHDuZX6sxqsNOQMmVkYx2RorgzBywUUyFU1HiOW1nO3e+OKWZy
HPZnZ/6sSBGBgIyAseSzMnYRkEkd547cGPyvXEd2EKk6/FOeg990HpHzPR10Dx02i2akTBdSK6A6
QmAHSu0o4ptljaP98oXaikwERyVl87xj8xCKgGEqHt5AfaG4xKv/XKE5iZ0lm7T8tyul2CxG6hZI
pBqwDEx8Bu7qepT0UmOGx7vQryYwdWKeWZ90vCe31lgNcrER17pAGCKaVU/NRZQP9l+6WmsnQ1JV
+iMAVEFwr8Ma4bYFrCCLi7IA5H8TkhuD9DsRyz44ZkEOI3z1H7hSJebuBUs25LAQOTIeF7PaWCk/
/Eb/WDFExtaY3B5rdGms5SyaRJAqTbMOF7XTqN2dXXYMzYmXoYrPwQCZVEo+THau+ekiuYiih75+
BcRmFtbzPhxkUa5MgXycguz/J97yj1GJI2qXOR1lU0I8XzhQV21dO1LCuZRW32WI75EeCfTjWZKi
ne0lUlYyEMtcYe4Hb9kk37RlTj1RNjHAJ+eHMY+DAIZfsQr6slLF+ols0VFkojUYp/Bl/BCbHUbB
FFXx/ocTAVIZnVaOTwaHTuGA8ZM/jNCwBlvrr9aW918F990Qn/pJpzRX8722B5ZSPVdgs8pOANfr
/k7Gu5DRLoR4Xa9Qry+ny66HLWkMy57BZj8PLnekYCtWVad0gJW4GrB/uq3YWI5bsYF1R2FUDc/x
KVtNhT5byzg1rC9Tqa2mk1p36cqdAojANgmvCfDBdyAmlJYgxoECti+1b14HDOhTt3X+izmufdfG
npikH0tcF/CjSXl3Ibs2cm3Z/4N4buBF1gM5+3QYMQtbNL2gJcjV4wGRaAbu3mqYou2xJaOnBHuc
l/BBFPXxbX590VB1jISXYLPuQ7yqe7Xq4YuHHKtl8/Z6QY4t1u0i7Dq4GSULpQm3G7VFik0VQK7H
Y2kDJnvaqWkKwJT0ca1sLV+ewSJvYx53DdFaqv7uMBJbY/2vXILMc78qI/znldBQUuQEb2nnf/K8
GdYGle68ATTCLKHICAIUfY4pPpChaT/h6bWUwYfKHdXFqQ7NqIE7Y7nOpQ1Q6dq0wi00rKUW+mZ+
7vG5pPrsqLipnU6LK9w5/LCR402ZoubinGUqXFlVUZvv+7ZYO5JEXBeDA3gbrrFfMiziuSklEIiO
XJqtov5hycfz4ZFyOiwCU2hGGgnSGT0e69QKWVChprq8smXdUXIlP0Z0+lk2Du9FhRI0JEmBeN/d
GDkSlCtWM22Jjor9EZ/0oDYSe4WK5MCTjDoaDKnxziBGjgBHcKmu4kLRXIK9b/z+eN/BLJDVUMVM
CzDgwx6r+kCJhB4SGZdjfgd4UTDvtrIhzwupw8ViITJofve7FWKTcAB0+x6Jv+7M5+AjN2bXdIQJ
C15+7yrNH3Esw1WXxYyufCC3NwZ+CFH2WK4EPEU/fjKG1KO8yZLSeYC8FdAI5+mb5zeuHS6RQtbD
OceiYcT6whBuFtqMScu8g3h6QjmB1xPK9+EISe9TGryOvVjorS4chZ8qWcKEV2Oyi9CBFRyD3nm8
v5JB0+LA6dZ1w0TqT0MjfAFATZH1yZmXVdtAp+BQ+fHazSyud72JZ7ALJnH3/1S5o3VpQwRVj3Vn
qv+FgJvEYpcNWEeiuIRgIGYl8um6yQNXEXhCwRGZpD4c0giYZ8zFsGad7r+5UJ+HiJ+PNz2xvYWO
ZgYrHuPGkpiQ3SFzEDSyDLsnJukzglgA+X0GP4hh0TFs1Q4VtF/YqcN00wpDirmGImNtFFtVHF0T
cJX6kJfn6ea+CBzg3v3Glka583Pz05mRdD12m8FN/iXrrLJ2jDvQKrEOCTsO3kYv9dokKA0STkkn
RKImFmORoqEIH1eA2Rwst6lI/xaOsP30nua3Pw0MSjxxVQJf8JWVfFXFe0XoKFC/ER7tWPkmVDpF
hAbyR1xyIMXQTrWe/8XBzwnXYd5ZYqFpkQWkZ2LHQlzWSnU7zisyvIUv8+Fp9KwgueXXLtGY7KXx
fWqhbgy4xGKm1Xi24nr8bBC7FCnxaXYkn9gjvIFmC8Jnbj5ZRahVRbX+M8Fzw+HOsB4lqtre0uYm
iVyyzRgyKBC7jtduz83+x2mcGh+CQ09/zjE9tZIjVl1oWTDwGMXqeUGETRUusjb6IO19cCJCjzDF
0oL46k6l57abnJCnJis46qZstcOFdqGN0iG+KDlRiZevDEg7XH6Gzx5kvHUZMnszEtoUAVK+E1lc
sQCeLXkWZ+UEvkC379u1v5rEwHNxAKp6EJnse4YubrRdDx/vXfh3Ysi0oGrz4hzhOQF0xWLfF6q+
3XE9DNdkCT/GS3EXZTj430XJ7YaaTwD/rvRAh8xfeqgMHc9N0sHZ3x7YEivSFdgWO8wjdQTdOmz1
LMWfoCLVtgh/J4DDVgCgKNwk+DURq0xFsljFwFSvzEU/yWVbMBfYOAyBD5DUyt2FKDcMweWVIlGy
9XvE9JNs4IBM6qgEQ0ITj5opygQuGhSqc+xI3/6aw9lT3Bmc1qMLQWTYq75SkvkmUwtU8z+xefEL
PvNo7Bi4kPryMmrRsdPavOZDYhbpjNnxWwLTgygGNY9b4LeflbPPzfANdr3kei3b7mOxykv9TNhN
BlOESVr59B9CuhO4ezi14DvrqNpZk9NqzPX6QbZRR6WX65zLgfvJ+Fq/GeLS1Kfkc4olGhZWDw43
Y0ugK7jC1iTxmzzSxs/biiH6Y13EWvlXTsgOEBMUp3NzAk4Ak6YjCUXT1+2Zuu5T1V38i+zYiSJf
sxwWwgMx3Yd8LgsaF+OOBZGnTNi/AjD6/ChWZXB1KEbGq3oj58AXmYWTI85utjMJ720pBY8n9YoY
hyg9u740buGj4N9Pt1TIez81bpxLCmNxrpTMy+/9BDDj0OMqidTHiGy79KBWXKIP5Wb0kTRgyUQd
toZzx03L6JmmW6RAG6guqIXCJY3GlhA4Kag8e2jOFtJ8r+aaJ/9bACinUvjC9BHZfFyyRyLhSbui
8T4glz4r70hOLMse9gkWHJogRtWNFxXm7C7F6636BdqFpfrlQBuv91wzAQYMXJUKpdnY3EBgwFaO
i61Yd5aA4RPAn+MX3S0RTBRxL4gozx8OLTheQocFpROxfilIYC84ul3aljYaeW9avkd5KVndlI4F
6Z6j7q+KmnnML/GlTdDAa/wJZdeX09lumIBbPoBGux1SuNC7uUwIIb9TXRDBvtiqfNgUlVqGp/sh
0KMH3o2M2IB1BrV4nb1VqI6ng++QqYb2nnGC7qbj5t8nO/lN6mI13HkOI351z25HMfOx6XtnAFt6
zRAd1vzFsdtPH+Fg8sgo77Ndf/4k7+zzp6D8vxmCODumKddZjEQGqb7lcdfiQDmZ3nGMoku6v+63
Y85WgEF40Qgt/WU42N/sKEFCigMOYY42UwONhHeoPZtBjGymmL6c4FnQ8MnNpuCOLNn5KM9YFnh8
5d5WqhcFiAY6nuN2mBebbcBPLJq/o07npDqU/iRWjRAM8XdCQp2T4PP/4d/5kmDc2RNOEbciMw5Q
zs43A2QIhwOOl+l8gxdksOKyvQt/eFpxzfmmGgyCT62VGBa8ZoMcZf7tL2NshFKdgqX3rHIdXbkr
9l5KVcPabi9dvUojMhSurkxa1Ld5UE0DL76ebKmJuYopBMd7s/fO056hxVUNT4kxN7sEdVHxoMWX
XOm3qqD0Htg9jUcMmlT2/7IYq+bbDhDAhQzOtbQVQgb35fKhEBA6QeyLmiwqjS+mU8/u0HqO2Gn5
t6w4ep6rj8sssxD4fWSSEH9u1wp3hhnLonPwnmRn6padhjR4QQwhj4isdjyy6vYbBPCh5VexINaq
EmiUGFs67XWq0appvTFLqapUixMbhxd0+N5LojB9etfra4O4Kf7PO7qaNvGu0edFrhCG1dCLguDn
263XcXEGw7EQzorbzhjBo8HC0Rvjk3EHdSCSsxNBP1+CcAjhTMXRFl1zEm5wrD9fD++r9oTp2TCX
wf2owSBwBier2OTjcanAegQ2TLR6xsgg4MiC402FR0ZfTd/4QecYpobbqpxiqt/4kV7Eskl/eEOZ
wKN87Wz5nVVG/uM/bX/Hl+TSBepOzd5jRlcwl0BA02cp1dERdC2ZREXzmPu9xxFms5rFVJwkIl+b
Y5NV4MujApEgBE/QpAJA8k0qhKhfPm7s71QZByyX8uZC7bD3vjg3J0TsrxrKojz56mTbAjDUEYYR
JO3iDlrLZJ7V5DYsj/EDvLy+jdAmEOeI5e09ozOITWlaiFbEcshg9Ess0AYVQkXV/DP8wdYkSC8U
aDOVg2FBR8x0PL97paVJ6bs4/WunmBFwWrWHAuQiRSNZaiZN6Oxs1WE+qNYzo9o0o/X0HeOuDxFg
d6WeUdGRtszDCW+1O1m1RZEbbu1gLP9ahViI5Sb3awsqSbQQ605ieAWUujjpR+9rgWB4QAXnAYSI
fm6g06oNWz1CAdRsSGtMTui2LHJVD6w8VbyQjYdTpVcmkRxtIPCEEpls+lLm2eVfgo8PIdwVHk7T
i34inN+1iH2pYDshfVugZSUfaLaE9jpQxC6na2zxkR6VYdWdHx6p/19ieuZoovll3DigFTjvHY8l
96Aj5uDg37PLEz7p0j3HC1a/s9NtSq8hvUku21IWrPy2TA8nAGwNjdf7O/ov9YhSUwVqxj184pUZ
yWznYj1lVf2ECTAvUn0nfxp1DDNiiJ0w4akvCIcHdmEjpie+iaagyI/vf/Vcdrtcr/T6tCicof3K
UvU3Lv1/OUsQrZz1GHhbzN8/miKPaX87MfTnEkUaCSM+/6URVJMqoZEZdmpq4tsxtWNBPwtVK79O
kciLPWdnQ2v84/HRFaCbp+qFlXoAOueFGWORyq0/bInqtlSJj8azfOQz30tcovRpRIJLWmRglJPu
XZEMIkpWbgRsoT6hKLZpo992kLJ/cjFC26NzerZ0SmFpblIw6saHvLr/1D2gGc0TqjqSlNrUwBvF
4S08YnHY+CPPdCycwbuZUvWvMi4EqJ1PKByvBQd1/iWD+PH04NGpHfXns///BZ9DAUi7gYdOeHXP
Rs99GGJ0+LOdnSU6tND1cpeXI0S78DxUPFj33Guuhxc3ArO4EMhizsr4Hq5iDe8+kDr+zedqT6xR
srx1l/a8NftaVmTcgAToi7VZaAh9mwKGkF1jsmvMzCbF8z5fxZ92oLvZCqmGhbQRjBHTmsMsxY7t
PGbIYbBoBaXz1J0r0R/D86Qo/SrSsg+VeCLTZHs7czaRSKvYCdwHhvWB31owa5yhaDOtK55dL3/G
ong2gw4nKwbaKtiwVWCRbbOMXn1o/CW0lfJM0UMpVh1C497IpSq0VlxQEZfUKRJo5rf5cboWD3ln
x5M/czwi61J8xVOcmwjn6WTsW7cI7T04ZafOcKYtohkBdeOe2CN5y5uWZdws6ww2Civr4XjzXdwC
8FI41QJI1zagFN5gEv1P9L9yCOzfAV0JzfmLosgtiNGIYZHvllrlErZqTNJDNx/Gg0crs1Z5epTy
BNOPepEdUSPPnOgME3Z6h0MaIfmngAjK64muSPtKXeJ2xM972czvaetC76C5YywTLYBZPHgTlA+j
HmTAimnlnJXMPR6bRk5g1z6BYNu7+TrYOYHCPpwSOXo8QXkP0Ybx0xgHDg9XYiLAF67LJ2ZYwfA9
NStbrUVQzpxcj5lHOahMblfK7orOBbcT0Zx8i5NeRCQonuY1wcAaWj1NNdkgjc/i5odAdbbP2BPS
sZei2oMiNW5uEABpITzWSDypNh2tqRc8Qt/johmVYUnhljkfX2H3s+SdSKC7cIEFQS5pIuJ04TDF
vgoCsvku/dCXJDdlQaLwpZzu2togIkYlyXf0IIsuhr5H85CmJNaAdp/BrbPrDTtIekRd5/J3MiED
HHNItBGNyKS9Jeub4NjeA8d/DdYn66Hrqiqkwb2CEK0nSeU4vrlnnMPgcqnsN3KLWvwxPtwh6zlO
atBKE2ZiV3AaRkUWGMIkieuDeeCfzd91R1Dla+HxPVGT3mdn/kIi0f4AOWIa4Mmkhn1vE0pUbI/T
79/K4iGapqmnaWHDu4BdQnPQJ5PB1ei5a6CigqhKY0M2eFfSYDK9UQrMOpFF0P3nMqewzi5p4WMK
Ne0Y7EqZxilQuEINNizTgvJzPL8GRk4B7nZvfmAaPNdcNNHcYLMdYx/8WCUMrkRorErrIE4g1ibY
43uWwjj4vycGWyMQULOTWvMkALTUF4abY8PMWyzESRFcfJpe3fxMXAmXI68bORgvwoimu6ZNiK6y
x4sojlW3fvLOkjLQk5JHfImKm53rC25IibK+Db/wqWKYfu5vIPHiDWTraC9P3a7+04Xoj91YGrBc
JJ/T9vTEGbcouHAvxdnFkRY5Q9WHRSZc7CrduLFIoQ7RhR71+kQ+O47/inmNPG8D5xwcwh3XMGHk
6N3I3EaTXgqvkW9/KfTUrf3xgYkdK8Kk3zHx4arGy44HiDQgAAE3G+nO1lmzLxbL1ePhLktK90fV
GKy4/gZehYnNciGyI4uL8fujoK7NIopwKiE1JngpEEV4wLA/OaRVG55am4+gr5tRZcExqFPE+9op
MpRhIe67dOpYRtwRpyjyYkPBIADI8/d6Ne3lAksqcnHmytWZG+Jf7n6A7770o8MZwLXwG+ZXK3qB
mNnP7l+m+uYIr40Taaw2txKQN9v2adefgQjsdbmHGi2J/v1+V8uZO4XPNDKyxX6sKri1qEBwz0ht
OCnPqQD7L5r7Qf1llgOGeQevVkjQOBHe1sBg8W898t2OG3aSlNGRe6c7CA2Qn4/cP4WWuhgMYGCi
XC//9fcp5aRgZyMK6QIRbrR7Mw1x+i0fMHswnRPXC1nKN+Ymf9t8xpiPetx/S5mbJ4/YE6IyJb5r
jpNVbDadWKS/7FkarbTV5GB+zyLm5poO0/YTn98nlSbmcdnPxSQf6cVYdLOLEbjmT+vrJ+kok0WY
fbYuLunPE7wRuy1Sf9llswMT+44HiNx6EWZhCxYVi+KubwbGFy6FBAxhm/Fu+1RsxEz7hycMJOD8
To3mhbe77RbZXpHNlwD7RQQRxFPTSh6fWF5t7lgnvXIyPAuhtI1e/bZ8XBiNcy2JLBdkXJKNX0G1
ksVAo2vt3WZkgprYVwsnbGNV2TlqldfuLXZ5f3NuBUhVwUjBHgv3bYN6r+B8AxnDNGfEx0L3Zez/
PtUEwkhr45OCoolWMWldGxM/UvgdhpJjpjHXwSVx3EKhIYsHD+7UJu0/E34u97v+V3+43yniBRLY
kiGBnZo6tdB93SvimUEpPO5bMO1Kujis3FoJiSHvWqhM+ZbnkhNBdgoZU0JrKfWYjFkax0/HugFm
B5otr81f4wNpwi/o3ZVX138VUsGarAPs/kZcx/eHuIL6MTppR/EXHxsMjL0xljtbsWEdj3Y7UW9A
cO303Zu2+Q71Enc6IoGWUEo6msJt6SZFeKFls2XQEdcVp+VHtPa7bi6IGLP4IMqeOJbGN5Jq40FF
FoPIUKtoDY8tsC5elNQUzVLx05NSBZIi/RcgZ3Wx+C0Q5ra8MistcrYVR6EEj7Vm+QPIXQDkI+KS
Dnm3symhTElcs+0YWDYYYT3RDLIdRWpZXso5Em51eyZAwKjoFwhFCwXV4/pSGnW026cusSIHs494
2SO6TNussS+E1DLXqkAVpD3uxgWBKRnQRWmXXCAA22oxq8L2JwF2y0MA4jsZ8tXdkIyNTXMJpLRZ
z5EIYhagAHZRrkTuDVAHm7vnWlzpECzKals/iAaSyQKDVJI/ji/OXmjw7kyo+CPsp+wjUaj82pgA
p+AVIhDWpZYUHLJRXd9vZMb4zwYtYe0+13e6PRqQMSjUSSiHU+CuQ0vt2PkZvTDGQz81ef5OmjK0
CprRM7jQHOJBoUn0P3lEtIFjYLEiAH1S55mo9INUF4+FaGwEt47seQuQvDxrIGHyeGCrTq7fJYHM
cObbgNNmA9rj0wI0PFOlwsFakjVsUf5MQQ59sSGy6IorYeL5eSxysuIvJH1BnyjfghMhIvbCGrXN
1CryXTFFY/+j0wNjNA8EsMy97TokZdJ73kekeWZTCt8PHDqtgJTmPJFgZZLq5IFczIGXEAKCoNOC
ZJcWeWBRkjErXHrvwem7gu/BuY3VgyJW/ErR7ENKNKPBsoZuIGm0EizCoKOxTibdDAJ2oty4lf8t
muARLiA4aLoYgMEZxAf7PzBbyUycAt9QDu4lAvXWinRh06M3ObZdLG3+SNzeV8S9mdAGOIHGOzzc
+dOH35husAG/PXM/Mukk/eQH3JUy/TNb/SV9aw3AUHfIdfBeSv+DvsOFbIGn6eXS/AA421gu1Fxn
hSH07xkYzWKzQdzvePKAXV4SORaS5p/1FMNtn/Bnc3tWYGxitdV6meNgYsEJujigHkbjHKswwjNP
42ByHowWY++g4ZeXOqRQOZPqJLRAJf1YKoDjA5BMbwlWQ6/Ja00eMP4H26PFSzW4UKZcsiZ5t0AI
N9pnB1C8y2xjZDNLjF8ICZGsAqtH/f2B01lMycGv5E+R9QqjsDOAfWdvBIM/ezsyrdrNuvK8PKWo
xnmLTSWVmi1W8glOGz54JsrAFQ5sjpdP0AxLkhg0q7m1lTFgFRwhObR8LuSzHMIUi+HLHOKVYw+e
6+RMhuXlxnm6AzlEph7XpmaxDYsS9CqyTXwohOPs4C/LclOdHn4fIOuTbRgYaoqxTakn/ic1DFbx
L6LR1ZOLrcT6/TbgVvZUX3aiJ6Tdl3GlBPSIpVbfht9kGj2RwVlT6dJP1Vm6crzTJSlcsF7+ktKJ
FUlQxYFRBbeHWhE1lKWVXbwY3vMDECBapdu4oRUnYyndqNdnxFCGuo401EHz+f46zMEdAvQrpVd1
spcE16cXcPp02TsxVvdlJ8azPko92FkFtF4ud8Xdofijl80IWTVvTzAHOCMQvY5yFZ+rZNtjX1AC
EHZQnv0KQV1eKnxcbCpXNWqQ4tAMgqt5SzV1SfSZJ/mndIb5H+Mr7CTiVwRX5EjajztF+GYqeJxD
mqaF5aJY6VA7ay8mDgmJPaxVAfNOku280L0gitDXRfuZZ8HglL0yBq/2NKz9MeRSVHnMA6i7aWSZ
3NNlTcZH6uQJLpDRgngwPVgj1dFcjDEpKzjpq879okHMTSyVVvX7gMbnfCtiCsyfzx9zE4oDPv6v
6h5O4Fs9kTfMb9Ruih94CqaQ9qbXGOHIcBQT3TwKDJKJNfyMX8F+YE1w5I2qT7CkLc9+ukCPnLq3
uX2cxBVe1wgg0eDo0AJN5mQG1Ahx7jAhuDkuQu2HwARN88GKqf5YrpK++kLBoaVu4ebkxrC7Cb/h
0Xcrf+MBULMXHl6hQiD0sfgNufE0d/SrvtaAx8ShcemNmAqdER0ZJkEjseooxwyNZ63UipM/vDMo
fFqTIn3mnF9eOPXTWv53Gu2F7QXdpbEFLT9YFR+qaU1csX1mAbWbK2A2d0VXLLiAh6ecoaPMviJe
TMe78xuDBUCWg2f3ezqjE/H2hhPKis+GUMEU8aSQM3L1PUEq9rQlCQXVOggx8MzVyml3ZUMsftol
xq3fA7ciDCRV9nKe8ijsUNSt6rqsb4yr+RgcYSads1T7COl4J1QbdNYxNAh5UdELv+IQmH/BHfdV
EocBm2CVXHniPPF2t92Bs3f1oRkLhi9h/EutPDZdU4ue+fdJeUle7FqtZMGdE1g1mDHajKIXgcnR
2p2sPPsXwrAbTupsHfkVTpxINSb+8N82KKysNxmXYHtd4hHx/hduuahXXY9YU0olS6QCNhsXOfOU
Nm8FaydCdI6knCtKZBmYvxpEfkaKU/e/+snfWctlu9LjWD/yPsIvhcZcqNeJ4nnbfj0Grfw6TSXQ
+ggqHWU78Wk+HsZYED15OCrX1Oa5XhbeYvAAFtrCXZD9a9JLqH7s3lvoGjz/FmbhEiPvfFTrmCqT
UmqvfYd7a9MTEcTmWQOhp17Bg6exMWAstSVMNTDArGPbT7aw+2Cq4IrxolgSSmO8OGULDCqtZPFU
7W8P8k3EJ1iMokIsuXGllR1n1zDa2grVd7USdapUixxon/2yrHHglIleW4fPd44XVoyyF5L1Uo4E
ViaebuqNzoWtGEZYBEUsrF4B6dcP5Dy7AAUApwvbtOIt1jJfSa2TvpjFuePraPeDQ4JYwJfGwRZ7
bolAPBW8POqj8Zoq2FurGsCpR0hcfYcskxO8VBY+iPwRJp/rwIX5RB2SFqlm0sOadqu96HXv443f
hnUajcFOM9b0oH6rhhc+JE32MX5tvuh0QuBNpxO8inXNlmZvnSp3FXxkEaebtTN4pFK+VwoyiAP1
3+xkxVb1IN5/h8ayzDwzwgsmnvRIx7a/x7uoAcQqn+BNliNZaBeXWCPmpJd0IgCWjv5zcJofXU2b
OKSecmd2dGDIkJZA0XVpqLJs2MjIHddsNAKr5rXOqVTOVCRO4Yp/ZxOOWINLS8GVnj+wDP4Zjg2q
PUMeRDDcHEMauvuonizx4zvDVUzZs6LXayOJ+7E4YyT79e6woKaAsZABOcl+XIpaKts0RXP+B25k
cO+V5BpUKt9xQyn8CXX4Jjf0+NJ8HO4CBsVXo3RbhEmRyPbKxPOxpaeH7a8CsecyHUygxHHvgWWy
y2NWMIRxeR2xCjf8NFDInOxpijq06G9SgaMRcLKMukacy1gcXKxNyB7Jx8Ml3WRKNukgACoQjvVk
frxvD3Ieyt0HxCTukxsRzOMu8KA+FR/qSv+gFtpNCLfif3TkDw8Xr54nxQteV1ERS6Bhj4KuCBFz
fNNepehs+wxkwthfrJIQgIy8iu2l5SFOz7DBvq9S7jZzLf5ISSz16VAI/MsAf5JQ52FW/sl4w8Mo
+Ec4KlL15bn6px/MT9vNwDgUR5aA4KlLIzx6xGr1Vfgpta9UgYqfsjiz5tnYKi2TE1zF9GX7L6XN
6OU9zrTQgzYHX2XhKDabqOU5T+QKdkFpVg29kDJYUEA7zXNwbPi7UnBcmMnjC644I7S8DiEal8HG
n/SzD9SeW4aAsissPEbHNLd8DbShEtStO/di3fVCz65t0yxWGnUM5s/wTmLdQevbWjJ85oogdAq3
WatGJoeCSdm/6L4YIu/u1wL8QAfJm2fESpbhP91ao3fDuvI2COsKLcErM8B7Wd1kF33zGib7TUIu
NaoR4ZgzECiB8uqLYhUWF1LHKJCarm0w8e4DKiGkaZAHCswUBs1NtIXsx7zy+rVhtfj26BUC1K6O
GL+KIF7ObtFsRNoGDzbtmASgHtrhh2DMr6VZrR92NziD/tii+hobq52tPvLlKQ+0//ImvtkkeuJN
kbQCqK+RkKSlEGacHlskNPO9GLIiKjTJaWiutoLj6QtSmaRx2jVTgRU4WMMsmnIagJ27ynSstlbj
Y4Hyg+SSlrq3f5loHYy4xcC55WAOeiQKEQ3uJyjFVYTHR1lMy9WJ/MDu9j1cBM0L4/OhFj6/+A7A
2nXBJsCWGOVQDm+0+C2XYD1qjHnLPjphnqQVTgH2z8Q5V64LZTM/HTejHJHvz8oAW3LO1LFvtccV
nkuNx4QHkWjlLf3BcTqW7i7SHzOsr1pwn8vnvgU4UckBlMopyE6+onhKLCtW4gGo7gU/PG1jfxsq
hsciNwAHtYpMJoc9K1MuQ3uibtfPY/7eNBqIMt8dRZH/Z3kgxfafDTCM+RL0OJFddzVLQW00LKyT
Ie7occPIx0XwA++4VbS0BOi8l8E2wdrsorMDC4xzGEbdJuju0tXP2vSOumCbDgclXkoKYQSAT53Z
KEXbKCa3rDpDAh12RI/YWsJo+85if8WIyDm+xhWmrisyILCo4jLHHkHJbM7YU5enaR78LZZujqHk
g//AQPJnwsFL5SB0Np/xXEVxLFQNIkclUMOUEbcGQSRD4aKG+Fc1ESAEFrnsPAaSTzk/FtKeSLMf
m6FyJKvC3lURHvBfI8gWDkIbxnaV2KUDjZbE2hP8CW3E8s37vcIufiNtdZzTMKpdmAQg54i+40Rz
oNrqTUCNJwkFXaMfp/MHGpaI03XCRSjkgC2rhTPFPjdF6Bad2L7IjTjxni+GB0Na/nqACe+ddFpR
5BfD5XGXNtf2q9ifK7k31uwkjCJsyYyECY1kpfybRHMP2gG8B7TjY/TtNegmmboRiGXstbm2fOz4
o0yjXU+dNjO1SGUbRYOpuhnYCIndhEiqWruB0SHp4Uq8cXoQYvOxriYM5MPf8eItkR5TdLGuc93D
khj/tKclvW58LNMKBa+ym4YH0IkIpvipMIW8KEbv+n+s/gF6mBXvUrklCXJIPo1d/8vSdw72wY6L
rWQuOTxCCUNOAV8jCRMISogqSHhF1PHLRDg9+/4XDTr1K3pDpHsv3Y0hX0/0OFNrWEsjygXN5xmc
ru5A3E7U+AIJdgru61MSk6aG5Jnv/R5UOtqzuTGC39Ao1A87AeZnUWNKPUxJvdP6WV5KcBvHTY/5
vC1/3bdlhfcglGKBN9dnx5QLMEXj+yBla129bihMT4/empUd9PfrZszpXrmBNefoKia2MgKuSce0
lhPkLX/6y2EGLFn7sjjTPsnShjKH+sLl7PAhXoLqzYvguyJdBctKUxPiy1a+OVCt2stZrw39s+TH
zWFDIcDCScKVDR7u6LbjJrTTS/OO9HL9b6QcfAxwzOvq0Y5RRD2aWA2R7zW/4YLlJLUkRi0BeK4w
e5kcIrmmQM/KjfUZHyJ8B1aNpZyjyXJv39zZ4IObQjuY3n0+5g/FM1W63KvTKDwKhu6LmiH2HqkQ
NA2UQMsngCFWmOnohukppbn3lMmniVWqVmZOYYUPI8WKc0rZk9gQiMi73t4iY4DMgyp33qYJMc6/
XtRZAa9lDyqheD9vhKLMjvnkZ9ZCcTdky7dceXa/z5Z+Ar8qYc1Mz1wIEmCd9sKJ/mbyFrBBKWcD
+NHpZzZmLqxQDShGOsFmdPZmNwZ71Sp11bDKNDJxPG/D7eupW8NiR9LnkZcPJDWptSIINFSehuwA
NKmp1gMH0SLCc9wssrSspWRHRgQzDRdwT6xqVtSF5sH/NtfcViqlhlJFundYvzuIfnnQZVWf1cN6
P5u8Z1idAzJyvwecUowyH0AB8WwrJgpTgNc+jHF0BVvd0nNupWWNGZt6slKjFXH4vSguJH3yC+md
6KensVb/LQpvlCuzFsG2lbzHU2T7Y+xO5acaeGm8Mr8XVoov2BeT3e6EJYrywxeKEgI+rZtVW9Nn
RUwtZ0lOBSxCz2fimf/5cRMjjOEcl0M16XgDV4jT6ptCleIpEvW3UbDXT8/KPqqNZmiDHQ7Q0B6f
XGpw3WYWgq3LWKzRiBaO++XWTGpD9yGQe9jczV5sBDyRQ6q6JO4OKHr37BEp4o/uImP3mitW4Clp
lwBrBBvsC/EjO5j+a1CPVMyyp1Tz/5bLUoPGXx+ZyqiY+tC4O68aa6kr56vKB8Wdob+7dsNAPF9f
RA56eYJ3+piumpKIyf67RWthM1K/kemeZxX10v4BwTt+b6fLhy+Uk49X511A4cG80Tauns9/xVfQ
cRACUhGRjgmyy0EbvfYwadF8JtgTleWut98SnujQ1wKqW8Jwk5RRQN09qlcviW3hV+lbOjQiU5iu
krzm+ZEKOgItx+4eqLETs9hlW3AgbX3OE7Pn12cvSbT7V218oAGXXShkp742emx2N6VLAlbQiZVX
DMHLEovUCRX5m9kgqcXPd4OtnkoyLZEh438k2uCyeKqGNsfgfGK54rJLW/5A92g1aKRZTydGY/10
Os7FsUs+1wJGOvS9Xj4nj72o4u0NSg7yAl9nHIKSk2k8E09fjKMOdalF0ifireoKmZrgOnEmVfQq
zQ2Gv4m1S9BeGpLLWqE3FLkfolohR83C12u+5QQdBI9hniGuqdAMudU1s6ZlMIbG5CXM1Xo2RC2R
71+8bUq0otI4SB/cLec+zgCryM/PAWi9Qo4xwvX7stY52gffJZp7QdoQQZqB19rmzsimiovCxjq6
k8TWhY08MdNTHVu2YbMVVBxZFrGxCsIFt3WiKlhB7jl1WI+GY42yJ2DLpnAFLSYrU/ADp/sfn/dO
Tl6cby3A+voB8VBjcyYMYl4RZ5ez28YGBbRSSXfALxhPSbNAXjqFJuLId5fc2abaUza16UzxMyu0
MK2Q1yublU1nvn1GGM3OtH+YaB7iFliyKoO5Zj/+xrBTO5UzMy5kDjLLCT6COuwKZWLO/aqwEfF6
9/TQN82LWLbJbKp0tmnJi6PrOkaFZz3J0AKWd2uffkmYChlxSun5C+wwHqolZ6R536WtXYLwcd2E
kyxM2XOIpiduDOraOhv7cLPT54ywGJnobEl1l/AffBIjnJjHKlSM5us8IiYnUxu/kZNddJXxwi36
7ZILgcj1xzY6aMy8rUC/nJ0Sv+jwv/A0qIQKuxN9NcfRHB9zlfrraPPMLOz7G6U+DdjFEucS6XKK
92RbVrv1QDWK+0j31WU0Ma0OijYAoapRH390gyBEdlZTDbnjMW3k16PiBbMw04JzgI8RcYOBc72r
c/iqsH3TrzSeyCvxlGBYmjhyHyX2wD7SuN1s6oaqWElIhe/tiuGKz0KDef9dzI9mARIjKi9oxi65
6AWFX69MRTufFx02uW8OwhUCjQTUSN8fMETkFJxmqC/+NTkdryQ9b/FpQ2nFycQkEmwVL4ZzomXB
RcaAkxm/jtnS/F/jGsWoVJ7mOHnVBvfRZgjINKx/imYszh0W4BlfIQ3IPqb/p2ovTb5wgnSHRzEz
40MRXknswdCsnAvJYaUE8tIhzeReH4X/WyqSAdwQ9FTqFH0CgAHazIGq/Y4nlREE1QGnmOOKc0Y0
RBR5ZO+DpK+pYy83QWEnyVPGuWYTyrICYPM2E0SBwquOYuUdBYrzBRYIlbBtn/kjJWH24Vcl5SS/
7fMc9O9K9edT+F7pufe7ddi/5GEXd1MqAQmEtMfJMN1GVNSMlB/7s0AsEkIOr3NupuELbltnFz0z
6PvQgKcv22lQ4w7FMUt8N5/TWKOv4xjqMzNvLpMUYFh+mRG9zWCTEvRMdnec53s78jqYwjN30uuT
qGGVzje/Gm2BXlKCG33lMP55YU9yB3exOrEYqjFiY0iV/7MqkCLZyNZJLIcuLfMfh/ht/WjMARNM
t/EJTFBDLcFWSwMuidQeidiZDO4oK8b12lhB2yNEuRQqItt3uaCI802b0n5i6W8/4LRjGjHMPsqY
TMmD1jT5dDuefwzvm3tw1Y9I/RfqBwrEZpDufmmTYl0P7DIRm6qn+mEeYcp13j1+oLgvErD7gj+p
SERFwyO4QTGj5iFo+lM9VHXiSaKiG1SEHGoyVxj8mRkJfDTaSocLkxg8Z2O2M/An8eLmEOUbfBUL
WXgZOjyOW8gX8nzCAJ65ppZTVswnga3L59e9Yf/L461/bIKLqyQtHpHblpIVUBHfh0GZt5g3DHVu
iF4qxyw7GWME09EjZMawRnXsTWrrVM6OXbZlm20jmQXE16OhS0/PYiGMBMt/dPQLztaSIgGfdRvx
isaSPlK4L+1FJaINtquDRlCA5wM84eIlQKNKxtmePQNcjV/cgOzMyte0v8GHFY/PelAZPmdZMMEH
FrT/hZNitJwKG2aBAsmump2MuhgHf1+joD095XdV3YB955KYTXxSoahbU6gIjtOwD4pnM49i21hK
BnVlZAei19LKmiYnICqYGjTsPuFtXaQOXGGSz7yH5jCtDb1eitvLC184L6TDPWgR6wFX8axBJkUP
K7br5nSiPaS+TwrnhHzvVP8ZAr5LLV1ehxfpVt1a/3N6urQCjiyczRlyUvxG/JmKoGrWf/3gRAYw
XP07OH9six+3OtlsqV/t6mDyhNV50OlpxhYlbtKdNKJs5iNzSxajjYotoyoOvBUVaRfBevPBz73E
bQm+DQvxGMCJ2RgUgjyBjB5VrBSikc/WbRkIQb1SbkzaYOsr5XIZQtwtOOO7bZ1cRxRNBYEcTyF/
rgnzL6/rKbTnaNkHvpmcL3hf2qB8B0aLWVfsLDYxvC+Le9PIeMUOJ0Hxb2pwFnp53zOsdlXpSLgt
NrV6MGO3R783Pq0Qy5W2kjwQJOf/LcHW7nbBZwo+neBmKlAMY27xHEuTYt7sJtz1PDFHE57h59k4
c0d7wXTPHMBS5u5+4OmzKXTh5BxHmrqeFOfPofMwpqJjZDkpmZVE0M8z/F1uplMqExkbbbv9drE0
WGEYLW1ewr0THPUaxUH3qdcH3imhOm3G+jdUwXP7naIi5fqv3H0FlJVnDFK1eu6sPaAxh/pPDhgj
3P+2W/PztCZs7Qr/v5bioQmdt1mE6iYx0kf5Wyls7ULFFa0PhaFRvZ0+nZTQFwfSZnq334iyaxzU
7M+RhNe1qlL7hUYnrmsC3PzfrEV6W91U1s/zH9IoBmOk0JkUvt5zmSpZdZz3+dnSyLfSmO5DPlUP
c5QVnykHr3pbm6RLOhqSrb1WW31KsgQfBIM6yyQIrdz4wn8Bqs+4mL/NMQxHYWqqTtlB/1v7/TmK
LpP4Cq23pf+rA8GEZ++yR4rHIeJ1hdoWo35q5UgKc8P38FlJQjfperj8YCz6SiJqGiQY/RZ181Vi
kWRVgdYBWzJnI9ZsOX6OzulfzhCihtXTIKAQf47CvQlpxvfu4zEQxM1M2X+biVq/d8Vmv/X7Y3K6
Rk4+sxrs/ryurUjG1TD6pD0yVXU4f+rz3A2BF3gTnkUIlfbm6/qtcVG481jwnCncaeF5OcZBbEj8
OXMCZeOSCM7hslkJPBLW98U6f2vmlfgz36WCJq28vymlQZW/2qcZkH0uQqY5k3T7MtG7At3XN7jd
CusIfijyxF/98j4MywjnaQAaZHJZTnw2HnNQc/crRK+SIUNYETBs2919Wz9uHH/XbdnR81rEUpNC
dMU7OaJZuRnb7sk/2+zyXrwv6pe9c00CyIGw35xoonBgUYZdfH/NJ8Kt+Y4BLwzadZolY3MUk0K/
wskutV9N+ZpSXAm1xmkgn4KmMH4esp8Rz20Z81EZv6yS48+zT0RhBRmu4LDc1tKh3HPeEWGQPduZ
eYpw2+3qleHs+87ZrOCfW06DWgHMzg0hEAegVzcPbr+rgJnRDtP/P/hZQjsyeDq53e7MGtwpmI9u
K//lYglMqe4AZieNO6/VEryJcDpAZQKC47FqzAwo+/GQgVe4uUZbkVvvlKkrpRrIJAyWn10Oo2xl
37ustmJ4tbIIJF8eFgxvPRWCb0pKk/fPYxoAKhGsKQyOuODH+TnBLwZzMacQtPRDsjX3KDytbTFt
0qdXGJAoLAqxO6R4UWV+mDjnwJGJsV7a2QpdHhwASrrQRACRCs0MQHA8hLRmCWzbfcYBxyhaRMk2
pfL66/WOL+YdaJeTgO+7mqbm6It/bSl1OkzO5G49QvX1Hel/J6cFanBFvvZq+1iYwY/rQf7U2KB0
HmrTNXOikhcZVEQ6qeMe0vN6HZe5W+rdaBnZR1BjELBFVV6QbJB2a/qw3/u9SyiHw3SXsW7joYnp
SkVzLd+Zm5qMSO5FGdgjNgLzJIoFhVxdFNMSroHMqpd3JB2sOXRj/AaIQdCj+Nk6jH0awEIdEyyT
AWwSBoD+tR5mWuTGoGdK2eS+KmAReJLgZxDyVZ00s1WEcYg4GR8XeMOi5JUlUExYUGl/ZcYZo1ix
7BvO9hrDk9JpQy+qoGXLY4Gkacj/1/bl0at4sjHGX4AfOGi6JJky1tmuQri5DHOAoR//xw7UBmhP
SNt/pOTdUsNs6db3z3Li3La5alnHw8vImdkeDAXtpOL0SkjGu6xW/I+LPmBntFgZ3k8oS1fFNBx9
nOkqwUSJ7IuBbBsqp+nhkb+JiRfpwi2PG9VEazGD2O5kvcHrnrpxhHK8PeIapdnvcGMS3VGgCLty
Pk5KF4/6/5GAzXv7WkdiUhUqz362OUFMY372ZoKBCHNEnlWyMMKhpU60dWUoQlOe7+LSH7MhCgjG
3UQpXF+WA+/9rrWlX9yB+h51vNWOcLsqplvtlcgywb8iJkV7uqpiFVedhtwN5rVvwdDYirhBuB/K
hZc6yO2aDLrNSo3wYYzQuW7RVZClq0WM9bvX/tRujjhaJZ2tAV87orkp4LVfgXLAgCyIYMS47uZz
AH+K4l/Q2Ud2ce6H0lqHRKMwO2Vf0r4guSwpALinnpNIebjUOSVTCAweSKpUSAkLvisY9xIGOLbo
QKtMVqeg+2HequMyhoFnHq7Yiqip+PyYRmVqbfjgfmXB/1fJq+pRJICYafyPD2f37tX9OGClWlvj
SRT+wgDl1os/vzsLUnIt1XRT9VAcWn8ZFSxMP/icynoamOwoTrQ8/eFfNvUTxUNaP5eYg22yM7SR
OBMAxFTMi/oBvFFC4NFXHlnmp1SVEpyoLwqdzBxZJJkrhfkaO51nI/Mer+v2bDW0WuElvf3k6VIY
FM6DCm4leeCxFyR7TEjh2qxOrvPk5t0EIAcsZ0z41WUIbMZQeyLrbY75dv8rwHPK+JvyIL+BL86w
dDc/dfMhBjy1jpE9/GZ+/ab+UYRmzcprxU60ZZI7RJzbx/NUZgj5VT6IsM483916es8iRA8WsCJc
QBogZujzsgb8jW2CnWaWjbewUcoMl71rSEUdd4wUCuwabykb+6LboaeRWjQtAHKq61hhKGyOLQ50
Zd78BEOtWFJu5y4H/gzF41pFBEyZntaTvoOkX8ExpQ0/JCWKFn05YtLBs3gAsivz9rptHvDXPdmj
T3Yt38zT6/4lkV7x1aBo+ysA3ScmVXi2Eg85cO92MHIJbcXXCIx8LCrddZP41QOnFlvylGccoE8I
hw7TiiJ8wPz2aTLIgz3ZoIqvTChB10AP6M43TnBMsD6r7dQqDec1z5hHW/R+BUupwNpCmIzzbgFR
z2wTndcpSU2hkkTzRXY6PgRtlmio4LzPrftfnql/gipOkRkoqntsljOXLhFo2xY03vrBdQSdJlI6
MSLEbRu/DOBrBMxcsQM5ejcylatFiOYIyeUqPHOSCf9+HlINFCdhxN8o1SxHmKeKP1QFS+C3Hqnu
dfVF7ORHELZ0Wto/dyOy5bIhTY/hyJJ6v/2nhTxvWxU8geGuhhKWL2WKceBUcpvudgopVZHp+2iN
7NR3sK9AsgsrrOzWA/MVSy9bXwDj43BCMCotJX35wD+S847C7WlgQm0/csDZxM01mpkjoVT3KxvB
no702RHvAhcWo0t+XCuQqnwm0pNtcYavCkCKPEhPwZPyNIQgS/c25UdEZit58Thl5bAgNRnqoTnT
EXVG/86GnCpD/BnwhOEyA36TJz7cYmnQxtVBplYVq9uOMSiCEPQdFYVeoNlfZjSY1aHhfWFO1htw
QjpXGxqPJ9Hauu3wUc2tLt0lVDREe1w1zsC93v2m2lIU8QacNdRTI+zZc1gb20gK7Lu8VcRbJeNY
bHQkcJ395Co9c/Sfpom6R1CUAGCPng7Z47DMwcN7qBzXXqY51BJOMxK2JpZ1SX/zmYkQoseX6Z7i
mOfpSbZNOs8UAwrZ19JNy6RJY79FrFXGOhU29DkEvORLfHoAMW8obNCPhqIpmFW3nczyfLls9Hv0
sOf6bquZm2Cboj+79Ew7seh28IK2S/+uyhEAG2b6xaikoF/Zc77ce+crKEa/Y4XedFiSpxVE40EB
XfARl5ml3KPwyRXU65/d3TMs3rA9mC9yHcXNhNSgDGSvjWAayLrVz9BdwRiXB7T3FuGMExuE6y3t
Z1RA0rC03UtGMkIxgoVxRr0Q/7uGDkB0MdEvtSLDfsbL4VU5VR5Gck8xId5KC0tq+Q1i38TIDb7a
/2Hufc4rc3JiMEAYcCfiXaTPgWGQn3UCMCOu7utfxreiIYLSBJBpdUk1e/gIgJFegF+hga3/PueW
lK7EVQ1qJfw04J+HOHNwQ7FaPhDRxdLJe4bbO6HvMtMIQNhdm41a6xosgo5iFjcwrQP8tH2i9MOa
ogS032Hk30sJ0Rk6ekzQhBsO3qULGTjJD+eeHhurzgGu4nEbPbXwYZE2K2gCaLmge9ozyu5XrUAN
lu7VqBllLA5Xx5C/8XdQtKfq/7RYIe6dWlEL2XNk1IKEJ6udradaNIhAasEDEJWZG2DFCr6LtTO6
IkymRQkCe8lTBMxoZ0I6AmA6As/mZd7Im1HCGDmIf1C1+c3phsNgHCPy7juvj/Dm00zd+Jh/DUP5
6DQE6JAMz5ADSJqLXEV6Avv0o7zG56T8SBbWxs2XTDwioHBN8S3236A7fo++C/wR8KR7sppi3rld
IIeZjWVfDceg5z/7gVshcrrpS+AtFXMycDJnto5A+Us6cghKY7j2U55jcHSJ69HQz6iC6AtYu0PO
Zp/EGwnNNSdP/Uii0T0ZgKlpA7pZ4g1EoLbdlJuecLOBzqsf4ZlCzujPnP6y2m/wBp9HdT/XCiQI
cocZ4TKo/yoRTxEBZUOdZiHo4dh4LaZcGYjMBQ6MSCTDV35Xl9HuSTFRB01sWQAvjJclAk6FX6ea
WpahrFRP09wfY4cKD0cfRSbXr55fzJubixgKyFWYdwNiumptx5x2UkXf3mHR8+3X7Nh/j8YY7+dm
Sz/sFsnZM0hW2V+0RJ8pJPjPCmmb5TAa5fbOr3gPQn8Qqx9xGiaWANL4jaCaTrltcxCrqiwcfd+k
fpHwAq5jfrcWlGqc2sycW/B8jZcT65vKKcX+QAvXJFU7KMsq1NUBJ1G+X08f2NpynOk6n/OFE7L+
Ofb1Z0lIFVsX9Q8V1vuCxcF/B92oA6H64UAFhrYMT+0grNlZnz5IiPbALHOs6Y7lW5KzGn6lhjcI
0Hl9akB5ogqahHNR6PCYRFDRJdAkqNUgJFVoi1ZFBIYg2DNLHExmJrK187A3TvN2qT399YgifXTu
DcQiRlfr/lg6a1uoVw2f9LCrCbhXjQuS9XbL1gBXOUdfYOf0ALmKwmqFaQ/eJMb5wHtawYSFjSA8
25o9Dh8VorKydnLmIxD+GncCTbOVmhfKDUh35bk+nTe8YIJ58bHknFS7C67boIhibgWQbA2B3TdJ
YoDa5DbH62ltKoIJ+qRFj5X2tTe8xlOKITYmQnGKGPZL7Uwr20ET8UdWV5qCLfQCTUQLND6jvn3t
C66aei8Po0ezNumI5KLbXKKUMDWnoBqe90VPcTHC/MqJ9YIT0sWSVD34e1yf31C7otnQB0gP4J4i
KClCcfeANgVfYDHRC3C07WFin6NiIcknoiNKKpcmu7so6Ys99IO0qJkMbbWqF7IaeyYbFTNVf3jR
FxfCs7dXMPvaTFj7gObe8XqdkIcFRoUCwRz5b2DnFwLZeJLZhQhTWB5HQGtsiwiX0jWvcf5G+xOF
qW5twMQSSFAYBHKCTytHpjSY+gm5hzIwwxMhGbaqTCKc8mJnY0nkY8t3WH/RjF9V/PHv8jnvQXgf
34t9e4G3lN75E42N5cMm5kSJLyjC/WGb5CLqdOTV7cxmw0BvqFoTMhxBPNU4myOU4I5icPb3d0D+
VvjoDXZstqKzihY3HcbnTKFQecn10Hm8CvrJ42TjR70oD0TMDbzjyIU6XAdMZBphlmxBEGrQrwR1
H4WyCm9rkdACNeHF1dVTURZBeX73UbBXTtzXcmEJmiXQnSaHGjF8Uoj7bohx/MZIT7VaUAtkeZfy
nNLGiz/REJXZ7+5dbN+Int2SVbBTGwzp1O2fEfKXTOo1aeeONDkgVT7II4ipYt+3x1N9jrXRWqsh
GEEC1i+sQ6Rsoi7S9hA277nUGRNN/SshO3bYDyqfZCLmnMyuDfxZcDhl5FYfGyeP1SEgfiixZP8T
fTJ+SamGDGBmDQ1jomlRAzJjEjeKHTX+ACRno/miHgl9WnIed1Qxew5+MmICHv0Mfzr3RrawnLk+
j6ucLuQDmPt+aIJ2JczVqyizplVtaF3dDpfj7UqkvGvpxd7XS/J1okA+EfY0rX3vpOZqu/U1j7NV
HNKxYFh2aFgH2ld2aFuJbQ6ZVnlQL7Sv5tFNVSteVtifdPyySgn3snilwEalCbdIsjtVtUbdo2aM
xRkMSa+4Ozjvd3+NdPAp/GLMYf+SRHyYnneOPBBbzLVY09F4c2/xbk+d+dHi6ulyAvzq4Sypz2Ip
0smCWr/wQP93XCNwgcg1KMRA8T0F2QbCnLo2AEyxZOAnfB6qxCrVaqhjS84Zrjw+dSnDfRg4G73I
nibJylJD9L+1RV1BX9VHklPn3Vrh0SJbObfdDqrXSPyYndLdyqP5UxpTl8EwruicCtg+hdhqufq9
l+1cBbJJ0LJ8oYkOq1CYsKVrI/NlCj5/i8+y+kp32tMCFLUkW1jrn99bv2/7raGZ2CuwG7HyTNrA
e6Q2YEayS5TkUfc9J0r015Yl5ztS7xzd6JBWXpNANIgy/zyOb1PsqSM4K/oKa4zo7fVdKhkApi/U
gg3/KIEeYCoJQL5rBoduOy/8dtvX7Gf9Z3XIZD1xMHHTqo1AwBUP9IvH8cryUy7pcVxTSjtASP61
mfpWHpGsoecRRIpLIT8uc0pruA2ZRlad9rrAU2Sk+oCQKBA09Rqc+zM1SRXNtxsOfSBzYERYLpH9
0Nqlg7HWEzMOaana8HeRW+180GjtA5Da9/zctiURYiOf1tLjAiqEjvu0RE/YfWMniPWyx5AcUhdE
yVcyzP7719VM/I7B6LGCMM5WbC45DjwokThqUlrivR06UoNtfU5wtYKquq3r2aTFC3N3okePqTFU
p7ocaUWxCq2dUCVW1mIwcHKAudd9VnAKYufwP7ddNS+CRfUqDwngwobEP4G0sAubUQwGvlkfHK3m
LzCtB/Zuqe9Fxq2u6pzkiwJCx8SOCx2r+KP1DSehTPIiDYkHmWb7SXxIcxry3vB35yjA9XGgJ+Xg
0i/Nkxv6bkoIR2+g7KEL2lfG1eFxqBNAL1MgnWbFeffdE+vp3Ks8+2Id02mIPln+oe7G+X1OzI1g
kCVJmvlEVJaYdMpUQQ3iTyYWGy0NPcf2reUoPyWYmM1D+HEgdGIEpEoLLwxthObbJfqsA4sC86SW
H81o6IXs+r9IUw7eZnIx38Ux6VmLPgUeJSU2jO7gLjFXmVi3jDcs8RdyoVg50/hiHfngS+DXZeEO
MsM108I0k28bkElGmqlZe6hXaRmg7i5KkvBaXSBghLXiIWf8ZhXcZIRe97Qprse7OJdJeElt2g7C
ivKnAO71Hede1GAJivmuRzIykQBIv8z8Rckat1fQWhlHroSRE56+0Llcs4HEFLCOueTyFraCfvWh
7fJcczzhjIH2tRFcIZ7CZOvBvjQB7YCgXGGboC3d82woy4xiiwmaTvnkjnq2OPXB+gFFmlIKSKaY
nOJduYgA2VSDd3kJBfHsbDb9r4vaLzPJrhBbXN9ptdhI7nHQ6iOCU5rZ597y38XCWO4mt1OlRq1B
m+OeCZXy4+VaHU/hvQFb+Zcq4FnZTlgv6cRNP7b+JGxGrwK9UMEG87jECnCsUH4qZMJZrLev+eib
1xjXqsFEwskpLYunssP7/wQk1UlQaqxP7SWZ/O/Y8VMeqi1VV0i/G6AR6ygdox27eTEN7iVQ9IZI
IJtQ0JGuyNrbKa49a7S9lkO86lUmBHbz+iTu+64bFJWsblbktitGXmJHnV+/1dpgVK0CPt4bhBkn
sCROXsLoco/MrX6KzLvteiDHcNN0oFj4rC/K6QPrn9BKCX7KNJyqZwsqLyefV0oaAWFryHMh9V03
DWvleOE3bNa5EUm+gsvUfvEvO4Sy1zHe6BOk7V3KBa1wMMgsBIU1uMNG8Gaox8+hHIgnHtDkurhX
zrCg4usKVRDu5UpchiZWuGedyk4SO7oB93Abjg+qhS9itDv4sdFouq4XHr41pZaX3hg9FyAtK+Uw
fLWEApweAjwZdGmnUrN/b+Qrj2lnsveuKilL+yjzhgcG/lmJ4J6rEkSCYAUrHpJS2XLyjIjJpk0I
soKn2O4jtJltFEcnkvy4LKYQhx1ho9gpKfDLETXS4Cjvl/pHbmNxnKPWk+nY20IBakkM0OXEw9Ls
+upplN8s+tv+BCRcIsBOnvUqrM+GX5/UCFTk03nsoP97D/zOV5TYtJl2/DqUgv0CBtiILhqlc/HU
EAw+cxLUNZY7pFgkofQxTID1mNviM0Qjl1u6sxtonJAIBWYoYpzIv7+T9KdUDXy8Hn7iOGMJLCe2
CbuqHhTwstE3O4dKruMqsPAygbuthzKip41KIw7iUgtHgn8IIVnyPqLopi6IZPLQn5k0IwhiaKoP
wdqANe9wWyuEWH3lmkw8CdTGCHLCqavGVKBf+htrMoDtHwUWs2eJMvUQT+HfBVKqXwJzIOGelBXU
Bg56qnqjeOnptza3XSViRcZGkSvLX2P8fE1xCwi+Lpn+9Hq6YhxrmDg2kWlDdqJdxz7kC6AbR2ei
RuA/QHVw2bigIZaYStklNmfXvPweN4NkrPevo4NUCDIyF5NnleNdK2f90KNPWTl33sDqqwSTHzmH
DuS1k9wrAqyIAZN7Lx2KOPrkgSgd77PD1v214G/WjS9CefI/MEkR4ZtU6a7WaFFai4vGKf2IZGXs
L91xYoIM8on07vhmofUytJXAGbC56RtTKqlYDZMc9CujUDAbTZb9YkXF9YVWrzOZJmPRWUWjwcKd
e6yRDDv/AeZ+wfzMkuLGW/nmVnQPtTV4JrCctDDvawva2GqjG/hzyHQfymuuBJNnrQA5WnAJeB1A
WM3f/Z/ocpnBwhrUDfTrFtHQ2tO0Sle3N6Gt8vdm8H1uCWUzxGVa7T528biOkte/5gvUGIAETrXR
O/H1DNtUAHEDPwk/LaATQIZDzx0zXyhXWgMKgdb9KoBhP9XkiwrFbTj6bR+Se9z23n1Bi9mEEKgZ
Cjt43x/3gmFHfdstr+ajMYyp96lXRUEQn+9aDUqc0z4HTtPyWllcIz24FPlqrRuCBOVZAWT2KSWh
s39C3pPwH2w5qyuyYi5CQP1vvUYSpmaaocagQ6dvByFI3PDYrYCmR8TBJ3PPSR0sgrvw81nsckPr
f0oRhf4ZhfbhxG3Idrmb/j7q9pvpyh5tfuGe5OK9MhCDzdjLWUxBoK3nR/6o4/46o2chEg4ywxM4
d/7h7ylZuKph/8tDEc5R1Hx1S3w8wnv7xhgzxaJPqTneEKAsLuSv2Ea18H6Vtv2LfZLQVHJ6EVDV
Wgy2BDQH1zzuZiFSXk7eqOihU3eqGV1YVbwCKBK6Ycg7pIa3U1/UHczgdZkxq/a8sakuxZBNvlTn
hsrXG/ZAf93KJECwKSVie7Zm8lWBN/WoqkdKZ8kXijXhRKvFxOKDuLJviUfr5m9In9b132zU4U4V
2RIUb+wvv1FKXkDYqL2kGHIRRxfgh6KSfLI67IZ6KF+ErLVD81ocLKLjUbVL0+KS1NFn1w5dY1HJ
JwZWNC6DHsda3RG3U57O3QZqX8nsj2dGyMGD/XZhpZcrvItawXxrayxbgnOeEHdKFx4Lz0YtlwhJ
U21cyuh6gjR3EVrP0CyvgPxHYxikQKqXd9u4cZv8ztJutOa8xiRgewKF5ihmkExy9RsL1FZncBnd
XxkbI9ZV+gD4TukMhbMROzlNMHTX1o7D+wR1UfkGR8Vmz4GUZd8KCuZ372MFlqIfaZA6qu65cjcr
CE5oIDiiNSpE/vc8T14wdnZyHqnUwg7INV54kzrKs3iFuTrUjUu5PrG+zuOORAebO591O0+E4VXl
3UAlHbbz4tBqPk8SwAI54ipIO5OteBlE1RlIYUsh/vOXzC5cjYQbvW2I4V2qyX1oJTztFTwydoXS
HaHIGQgLlb/k9bahrvWDlbKFqt5jU5bo+MF1H9USfmLMUAusOlmWf/gwq8SsIdRudltKkrMME+ie
683HmJECIXAf4qnKSufimVS5UlSf+u39pkh4N33epxl6o24YTpf0Q76KiCiqCgk4uDmQrB+Rva/N
zb51j35bcVbGPrnVM11v7Af4jaOroHofHom/0pocARtyS1vjIbwltDFgpv5POAeAezfd7G4WCkEP
1wQn2q0AdmA8YaDDtqOceVPme5yBh90zOM0er0OcOCcy9WL30gIvjYCJ1Ulfy9b6x8mkpJwHCWuP
jSGAkADtLz1KLKJX4a2nkKN4ZzQIev1cr+5pQcqcJiUIb26GrR3PJb0nPtBEdCVttmuFfJ6RD3Y7
Rwfh32RzJ0xmANszfapQmzvN+Sc12eON+UlRJQP5117CnJExv8zcY1YcxNyo/kTqGx96rPznP5/R
RH8hFPwcJr1UgKaSELtwPXVHB8iUi54JAWDJJaQj8ELhFQN3MkoHR7IKbCR6zpScFgZTU5/nIn5f
gBUXD34LCwx8NH64bOajxC2vhz/2hhgLjL8iS9gUATucsONbS0NH3PYZkjfjNgyPuZ14sjjEHzUa
S3o5g+SvaAslAdqZW4EKkqHJzMBgiqqYMgF88dxQftPOWmuNCZq9WCCner3lrHZdJmU5rNAzxrXY
J+QBAFsmZkMk69THJVE/RQ5/wwTYNLRSVZojUUwZO3Fvhe6sw/+deUEwYeqp96WL0f84Xk6P/bai
ZJzH0Cq9MhD9/ZsPT0U7kVPkc+229vYDgpVE91PzfUtoQ+uaS8fLImob6lRtv/En/IngLfQPezCU
VomlVBetEgVzsVPxpFDlVgV0976Ur18e/MuJSHopARxKAXMCsgug1E/jFOBV5CYQ7Dpi2/LRwRHe
7UTp6XUWVgqnf3Jnxh/6UcL0ZzCYNCkiLkCHibwDEG7hDcpv0l2fcbJAqEnpRgAuDtHT3x4vSZkO
AWpmiFSI+L/FzhlisYbauLL8p/bgL4oxMS05p6yCe75L2mQ1Nv2eIGrUq+6+ueGr37LUDDNHOWwx
CaIjlNYZaze4QKA4+/gXWLSjQ2+xXd8H4bUnnW0/XpQBnCWNN+/rqnKvMTWGTDx+FhOJVY6XxPEg
fzeQFGuJS3md7rrYkog7VFA0J/yTs5l1Bk1MrxeU02N2ahk3XKWpiCvWwUrjhEukGoyWLKvjWmay
4jbluXWi354epEjOHCgoTWl75fd2MDUEoapSBH/CJryl79gryhZm+JbuE0mkP1X6XAcBIQInhvl3
46p9yNDmHjOz1nRioWbT/lqQ4x7RIs6XZ2LOncYD0IiCrW8V1AGHuQFxU4LLMe4p1BWmFdDPQmqo
XTIV2i76icqHSWhcnyStdZQ1Khxms4nzWmnWLVXtOYHgAv8vejuqcPON3HLvDiII3Yvi9xxJqc8R
PlfANDzKFoBNJgSsJBszTwngDBgLvEKGAt9u5qsKE4r/QnOdZDPRkE+kdkf2qnoCfaSes8jhx9fx
MJ6Z3JpD+hicw62Q2+O5ybzXVMB+m/YM3fG6nhWqXZ0heL+qUQpYnxMovZVqzZ5Glah/K9m0BDvF
mL89cFuM6jnDseLgoDvVmAtHqyAx+iLjATapMKV9fnIGur0scsDxC3SoHHxsKiwrg2CKxv+SqOAa
PXFVYGMnNMf+2aynCDyS8jDb1YLtwYXJR7CRWksQdhsqNr8XUQMVxR5o8Vi6EUSWWlhIZxYu8R3K
pP7OEsGk1mY62O18t9Dky92oiQ/C8hmEgMySDVHK93sU1SQ+85QZneHB+GiNOe4pHbdCuQ4AGgJr
QJUkU1tfa3zH8MDdf7N0NsH1ohcgHDHEfUBKNZX7ZV++jK6kpSAjYlsgwB+xI9/4MwZlR6YIC92D
GcigPnfSXmnwpL8KOPgN1UmTNjqZsQeMEACcqrRSf56f2Ef40GLaL5tCnf0TSONxVMg7Pcr0ZcDC
JLG/X4rBhwxLYjDWw6JhCjYAl/znRU0CGljahjo7eO+uXpkT87eMwaWRz6igkE+zzeUF6N6NpTRF
yRLmPzvLp8jMI2LuNZh7pk91cmJR8we1YB/MrZMN8pc4OrQJQE9Eg5I5MnT39Mg9mT6m50rdv5J0
Hy++Hb+DWxC2Ylw9wuFij3if5xs8ZxxxVnUy7vizgfsuDYAXIsRqLh7Y49zKWg/bmJWy+xJhKNBs
OqVeIACf3bwwy+xKhufI5p6BU65fnziVqYZBQshd5a2JmS01p9IYHSDo6oLDcwSzl1nrYUWb3OUM
+MbmCxeUh6MyIighn0fezp63BOOUsUuRekYXmdfmcqIh4MHcAficLf6daxqQsXaw3yBGXdjihHb4
6beQu0QAPjmI4tTMyuC3Wghc0A4pufWnQ/FF8VxB3uH9GyuUyP5QJ7hSbIKMQOthMz0YKLb0w3vp
AAy7W3Gk82pj9VnT5ZX28zrb7+Ohb1Ce5k6WYZBpVcidr5qGH/BtczV7Qqloxf0EmTCE3kUkm9qQ
/vrgRzSeDksIIrUFvFat7h2W484BrI/DUYQM2eaWsy6gpIlwut2GtcmkvN0QLSeMglmJNuahPoNT
3Itjo7Sr3JifmI8yassQ+bAJBlRboGlVUz4zT9Yd+LrtdPAtWrMG4KtCiUjFe3vX64T4fruvaebA
Yvlv3sydTl35dvTUwyxLfnP+8wvxoB22gMt9/EoloaSW08H0/73ZunjTSg+2qWnAs4TRoOIzPl7F
dAqiGcIrm4WB1Cjp0DNAqmpEuqdGLm9Yd4qtdiXVw61PtJhQ5M/sqhqRF9vnwrE6/iUiXOvkFFJ2
vN0OkYAiAIdJvvnePzhIAcaGsadgnQMyVvuWURSSZFXEh+6xfK0Pa1GeI03546ZoSTslczMt2TYn
XUFe5S/2fQXymf1abjQ4M5yrniqo09gkW1NSeTpltzUP8S+mD1YXu68GaWya2c2KkCCOEV5eRnmb
16Auw/zk0EPukFHELcYg8O3KMUx3WYunw2v7+T6/dqGDXoAR/fkA1mw1qkudGv+1B8ddwXumraZT
CPi7VfdhcNG/CFc5m/EWgw4xS+Eq5J2HZJicjc7UKgWrwIxkw3zDTQI191cO6eCKWejxzV0fX+Ov
poLhuohgHMmcH17dOFqqonABNhli7A1wk0tY3VQQ9kT1b7A2lmsWxVgOexA9iy0kR/f46OT285Wu
kVuDkyuICphGrED8AusURQeqHxU6qHq1ednEsnxZFOGQRjJ+xY2Uipxr31nb4Uuk16Ul0H100O+i
/MzHZW4Pqg2S6nQOxBzOaSoY5QxPfojDg8XvOLMcDUBWS8aqlUBtfjBF44yaixFpvSvAUdXlzgS4
ecalKWj5lvgYASnszOBDZRDXEkqrkv34CEmRQ+U4AyB/5l6Rslr67sVYO11eyPDKOu7gJP5lEqZZ
Q5XvzFkm8RqItnq+XV6Cs+j1wxIiBKB4WCbIjgCwjUWeOeP1e+JH2m+mXMumxjqsjYLISu1YcsdD
aLN6l1roC4coc3R8M5++UhYBRU2M+p65kwkCaaoDQnWx9d51Z77l66wFXsgAloGjjkaWEY/iN4Xi
jr1nz4FE0MOeLIkHzd/wNFRxIOZzOITx98CWssR+CfuCdFC4uZTTipk87OGfywY4oo4/83FgYX6P
XIfUy6s/Vsm6JnrWwJoIslwniKvFGtqmaxXYdeO25jNTOYDMAI/MQYSYNB7qiPS0kCoRHjYfgqN9
UGyS0mV+7pDWN7uOP6hB+oGgKrt5DdnlBQVs5FCENTRmQMAQAHFNbknAhz6RefYF7wi3v0EGzzan
t4BBQogwanczvfot+nJyXLkFIkor3UZYIQuJYfB7pTfQRa7qjfPMg/repxiwCmw24Rl5kAH9LzOr
7PJySXTxvbF5oeE3U/gUe/ix1NWmRGlH1DLLCps67XVFXeH1LdbzMmmwZwweKIGQDM/eaTG+cO1R
czfBYjgch6z6J4VEXIj2ajm83TWtBZubXgqvRiGAPZB06hEDynMr2nAB83TGDuegtOSl9G3du2xu
E7TQQIB8/Dos1TZgwmi0yJJ5mpzNstO1f1YEofKKQ+pZIiDSzX0NLceEEtgJFaw+lnwh7EoXsNMc
XAxNNY7HTNgiVduPtaFYKpy05lorlEt5pF3PMfq4Qi5WQpQz68+BONlWrsYKGyYqXvcL5KxqVpb1
oT4sIkEiwH/h4lgAol47bYU+Kgc9dMnvyeiIYAPmbzaAcKXwJ7TvMNIPAmURgWvGjuc0wzsP4Fc3
x+GrU53m8PCrbVFz3w/4lfX7+4OXc3xdAThwpnDz2P0qh1yyYVrXERuJJSEBZGl/0RJoMJcZhlPm
SHUk+gQLFTytW42PBWl4zUNBDCFZS9u9MI2Wv7WbOvgyrJF1StSUy7QIxMawDuDx5f4ctjVvYyWw
UGCpUORsIepvB0PhgkWG0Apz2zwRJr/z4czd043JFc7ilPZ2nTDRGBEqbHC5OEqO+M/ZDj0/xV1f
hMwf3AyabR2w5X9lCalmlBfoSxHX9ZRvSc3miM4yd/9/SWWzmH8ZiYaMWpMRejcLGHOw7U5C8hK4
j5sVrjCAUGmp+qMA5NnPSfb3RNeZJZCZUSbkmLJp6UOWxOgvd6sSP5YTjRw5PFZ5oIaY+rBzJbXS
/P+PQy0n5iGN91Ukz4D7PZ0pn3xZsc7tNIKDDFRYt2l/NcG29C28Hk0vZ/kldIxMe2wv+2/e4L1P
TkSn+lW1u56XF9qJIuExPjxSNbOGO5DyFK9QQAODCRkdpWB+ZJ76Fc6mKsLPOgY5uCkPjM1Z7EFd
GIsWgcr0nK9jbO+IzJJUrW7SF+USuUSKyJGKPt4GLiWtJvFZW48f1NOspYqsEDSCteo6nUr6meJK
3tekZ6TZGADFVN+iA5EC4cdVRKolvh+pCE93GhIzMvm+2+HXDBzW4oL2HXy+WfiEn9PKMykdgp01
lMvEaa6WGILywYS1Oj7MmPv8RDtd9A23w3FERZ9I+7t632FBCBtLX/cZpegkyS2d/6iLfBOYFfbV
/JiEhaN1DoFhIqQt42Ug3HJw0h3bRTFSWMT1RsNuHh9SSmobI87Y5gN54jU/80MeIsEzzjufh3vW
/wX4VXHPJmoFKCroPmZc2CuGYhxAN8R1qDIbXp99Uw2usoottJa5xGrz+jr2UmTdFkiWthtzVLip
oruQrIRqJAJsq39aZXafGj4HRAer3mbKmCgpaPc+BgVh+Cco6oOOY4tIviUaDoWzLdoPZKZNTjhL
U8ilrgaOf+4igqSQSsFz7qkc8JskD/Q3UzyZTm0bgHPlBWZfRJFb6gv2Qq0YCc/ok9JY/s7d2vop
5NUQWLc/vP+XOqLtYHRYGaVn6LJfaYi189s7aPl9zMR2HykbUcZS6r931f1APn/ZbKB+j0BPv6Yv
8VsQmfIWSVRKTYL15yUnW7LFz6Dg7LokeT7HMhYK7xXk4wmxNVSa2BY91zh1PC8DP8lZOygqYw4O
yK/WdgEe0uzKNxAVScRoyh8d7uLphWEd1AP6a8JWSbVUZNzSZQ96xa2vXsPzpeehXKRi+U4uk4Eg
+Y9GYyXi8ucR8JvsZDU+doyEzRAPeOV2oJkFpZS6QVznHTfquduycxJsGwsCAvVLm85Z3lshQtqJ
3oadrS4Lp8N8U7DyTugN1fsTVRtOrFr1hwHKRpbyUp/16kxj14CySW1ptHvOQUxSRBqrKp2u8hwm
0VVdHt+xvyNb6yZJgByU/JtJd7RlquWUZBOpp12blNv1pLV1eHCxjh3FsdmfxU531oIEFibsvHPI
d0P6xQApM4XVJ+PD09wYxNg8u+nZZhAHJGIGRES772AOAhicx1teQW8y2RTawJCuS3Tx0IB+qOIU
L41WgKOFmgIdMmFgOMFOTieCN4c+1avbcZ2fOeWU10PwPx/5Nm3+26u2WH+N4I64Hf4fvB+CGsVB
LVxaSp1u8EZ9cX4eedbtMVL+VgI3KnTGQJQu6Lq1bnDn75dxpIMC3ZTvcfnmjtxPcX+ct36VNLHM
Pv7grQfB2WZE4d0pR+U5/AGSDT+PxQVaroedenOJR4nPBuIqWEVymHERc8fOmtEFMBI3DTJgTFu1
WjmenSaOSfEuRgUs9Jq+vxzo97Fgvt4uefHQRuMBzopn1cxMRPWvHEcol32ABGu6WP6fOBmoSqH4
62UPiF3xwRt05AH3lpUmKPqcU9R1ctOGW0b1eGG32XZAfJ3nm22g0PWGwYHapHObjjWSxL4CZjjP
RGDxTvZUUc37Szoby4xD9Ny4NV5+V/8xOhAUYm2BkiqXreAgKIgbu36GeN9NgPXU0RLmAVPVUiia
qvoelarKISSk2tg6kjUOC667Dx25BxJnxF8aR9kybzU74tba3eD2NIGYPvum5J2POaexX1B1JBQm
CPiB14+l+4LCdXwvRUL+vse2vPwp1C6C5SoqYfSLQCWItiE0ycjO7whDGc8hKvHYbID8bpUWgBhI
MnHylHSkCKgcJc13NrjnjC9T4PDvuMYn4FF+gmXugtAi6Mzt2KpR9TuWLzUv00O1byxmFUsjoHeh
vjGgt/pAWNIvAUbvMWEsA2MxhQWMxI4w4zUXCUq/fvUzkaAH3VIMxHjqbT1/DacAqCL86yK00aW1
qGpwapUXOf5RsWNNDR2SbFB6xfHxvXxMpQ1RcXgvqtdFyvFonloUb3aMCkj1U6O3MhvzTHU9D0+i
wA3qjWIjpE777AgvgznjuCeQWQtPXcMk7CVtin+GZ5t30VFOapANAmYMHzXxby/i9gX7POS8r9Sb
5GbKdYoF5e7u11JfnlbXyjRKLCeYKDtJFmIue0iLkGlJXfbIMKy0EL5smi/2tzRDSl5UYrnWWiG/
sMcrCtN4nA+D0CUJtp3/3uYY+n3kJkAzAAfsmldwOHd5QKCzZ/x/3te/WHMCFWdI1hRlWzBDLGoE
3+M+oUgYIJ+zxHpk8wvHME5QVIr1qDojbYdngsuWE9NJHHcmC+ClSckkau2YR1p5MBwkNs3UjLS/
tdv7vcDBHyXP++cU16pWVyIlPKw99msMbp8Tp9GOTg6RBnMFI5weW7IoLdxRevyukBie8Afuux4k
Z5fUZhw6h7JxY3EXmhq5EzjUZg8s7xoOvg0JxMKor5AG9qMfJ7tfER4pcykppxPvGnyfLQiiotDU
oEA6Xbc1TPV7SQsDtwXiP1nukZMHvURN0uAkHFT1qv65edP7S8eFX7CiiYfXWJt+r6wWJN+FUsTq
bGxQ3EUuDPf0IDF3P4HPotBhsuaP5p+nfqckFk/pYvpZEGoY0BflFuSksxx5bgbicUn3rq9ZCl3C
Y+8pBzzPXvbuEyELdev30HbsKR2QZzDg58DhpNlo18boXweR3y+w296EYFJzrajm7GVQK8qTv8am
enyUGu1pZNCSIHon3QeDsmTosAVwEO5ZjlCkUi34hRTbMW8IJX3m3HqcEhBwPImXPtbOr/0G+blB
yILNafa3mHnJ2N8su+dN6OsPHDka7lTSRh12P5FXyOtmT5RUaIXgEz0C68vvnMXKHN1pjYVFfKHf
LZ/T9qUbE+n32f59TSFeU90dI1QqFddNOphWhBp7nchkc9x/pgl3fJpmw+ka+39VSpcp3UgbcvYb
jXD0H+BKSSKG5uuXJSyMx7aQ0sP+4Ynmhr+/x+Z67QjiXK3ytksarx0tWwh1oJYP7rcCcd7OFBHt
HCTnM9u20kmr3HlhB5wbk6+xisveJBu3E1BIkhn/uyD7k4n/xib7XJFXmeFkZKI46byLmJ9Wn6IQ
aF92wbMVUpteBjNd30g2LnLhsxitGDaqLRLyatH/IoWQYqvxln2qS1fUL8Vx974XZRIIHVCJ3iot
3Ha6gElQerOEzGrJ/pxRn6amzmfAml6qdOrRTsHy8sq6GsXT0DcRLo+sO2WxEYBB1R+IZfUCoItb
QCQffHzn7EOIdWu4s8EZC3Na44CnDhMc/RTnSjW2TodaFHbZDUnKqLDkgvHYGa1By64/8AvEaUay
AiHd36tK6ll1kOKAeBDOtf4l0ut0tQ5eLSxgLDuA/YH5tMnQ8TaZt69NX+eHDwtM/ZjMNWpDlUWl
G7mCeuNKESlHdy1t29Rs84uLfD1g380YZU5AgL7S3Eiv0iAuojv4395IfTfeCSafGuJXz57iD0Oc
WSqTmegmsqqtsBpVa4whJycn0/YveIn9UuAH3/W+GK6J+/1DU4Q0B10avexVokh1jUetquHszKgO
JGmeV4Uo1DqOJh65tZlULmVKqer6Pr8qlu7BLJb3AdoJ8e4bgWEJGwErxkR1uHzJ1Pc88EcHMSAL
mjJe/5YAAqDGX5Hx2M0FHk+f4ASu3R10cuH+39f3UIbku0scJr/B7Lp1MxCHifVS8hzV8KySr4Jw
Gzrbb7MwzqrgCZIVrZE63udOazOfc0v3z/HgTP2XOdm8HS+2E5dkS4DIRGSmIsq7W7Ol5u3IkXP2
oqu8dCCjI9QjGlWGAv86sME+tCVPlq5iFQpaWjfAoIV7aCuvTgd+hYfaJAhe+mNXNbzQ+NWf2li/
z2l3jWUwoQDwO/kbDZ5dwdatdGG5IXTpLQ5ODwd9dEeuaO8/SdYkFJIVQhI8E80/G7IqT2qJiQv6
UAPllUCVYkhM08qOUD05tzzWpNIxcmwofM/9eIomr5mmpRCU2lGtadUhEFizFwcaNNrqObauW4Rk
pMeO+ZEZeh4gIVcqByZx177vYudB94qGHvrjesjwvHV41k/FM8SJx0vBgFXbB4CWFxicErCysBvT
e7CL+ViRdjJKzxv1G7CL+ZVLw7r5pBSspqnBE4Tf6vypLpXN2j+EBkpbfBRg0GsfQk24twVHALpU
/TXIwPzoNytFLKLhzHs2/gb+ZnZfUeNpddMUYACFaVf6D9LHeuBdLeHUCmNuQ5kHhFsUJk2a3FMQ
myD5lO6itN3dUP2EUmC8gRcjSYOQw17a5zL3UEjOMJYkuarhhL0aPiW8gWQNJHSA2xrLiMZQEZrM
+3k1kmcqnAsIC6lT8x4mknsjmO/2wNtNyavKHsm7frscwYMtWD01h7/fZ+GHdfWZp2GrbGTY33QF
s+C9NFi4ehPiM078+N8wzydM9eSavDVc0y4TZ5giwZ0B7n40oA+CgfM3q9/S16ghdUuWL6sGU1Xg
/I34qiMeF6QQYxIL9ICjG8oJWJ0CxF2DlkX90VzukKMRMzRdqP1J/v13NLotJUGTVrsZqpktCwNy
OP7LLNTJdsfI5WVPfiSj1uJHgJakOVF8KAIOg3lWedsVD0uw/X0WTW+c6JvfpOTLWDMhOKimKHM8
ycWnENR+ouz9HR6+IXBFleku5yr+h9050UexnT1PyXs+7SOcBuPyvfWtURBg0nyo6D+kB1ae3neH
HAnJRrUnZz9yi7PghBQz10D8HlxDXx3NkzK63ZsfiTl6AuCc+U4OZPvJq1VSpFd8Qc+M6dw+xe6D
riTmK7Tw4+xyARQJagiBL12gGYlJe4hyp5oPdwXd0rwFPtkcU9Hyu2nMkELVMKQEZrVk2iFuqy25
nUDzrSyYfuGl3HEdBYofpEdmwsqqWdi4ySXk7YUdnkfZ+T+qWufUe3irEpGupMTMMkAulJXPUgPh
BYISRok3KDOOBailu6WuMNtPTlNx1lnJdPJTD2t0U2ZLDEWHaOJ0jxumRt0K4Z74EhA1Uzt0hTVH
Gk6k2xrJjaRjMPBcbIZlIaTzUQw8rFR0NIv7b/bUaff29nSEpg8MSUChn7ZNqMlwdv8rRCwslMaX
KL85Y7vaIOyfqHl9fVOsYmx28AAmLl/eGyCc9gXSHEzP4LJMUMn54d5PtmddZx1A61qIW5h24xeg
w3Bt0iYQ+q+4SZF5Le4uzlDGVBu4tdlpGsYIIfRQB10tbfJ6TCLpAbZiTZnwU608UzVR4qdt9GW2
3advZbn06+4HZpq365Bd8zdIrvjHbpxi/zZEQ62+QUQY+t6aOOziIwc0mLLppmdCJtQ4Iwt5UHDX
vvcj5NoUuViaztUkPEJHFxEilBlMFqwf4qqZcGBWiBMBZAD/C5lbEk3MGBVvhjHxEqXV4hKXlvaZ
p+CMRCHsBu5OJI205d/Bf30z12MJbI4ezS5PTKtjiu0Hlt1hnVvh7xhho+ekmslIdReIBlUXFi/y
MVw7z14/RfgbHsHT64MZYa9pOEfw28tShfW4GM83G6Wu+VKwOi7bPZnsmOdBPzz9psp3Qob9iYdN
IrfAPzvy5gERLyPdgHQVVamgklaRTVb2FchXXKMHiYw2UFouvwCnoxqzrNCcnHu06OFSK0OZk6t2
riiEbjwf8gQnFEqv6l8uoQOvJaCooQOUWxIDNSum/C9pb0A0H3a+k0U/hiyKBeAVIcskGTRzqALc
mHFnlC4lAFGf2wb7BgvL1LGkMzotIc9Ww+f4c/uZVh6xJXSWgDkKdCl/CnPlvN39aEJliTnZbeff
wLD+1hq5iy6Z8nDrJ8qNXpP47iQ/l7RWm1lwmXAcoK5x69o+HdB0g97/+5SfVWA1HoTFuuxO6QZj
EkQiZej28KtDtdTUvGs8OCVH7MPM1YH8Wc7/tmjL9BfnvmkfBM6raaLNSnBA0Y0pZsrlIr0IV9e9
8KVsUBBKRsz6oFKH57K1/T9Sx37jn7FuXpDt7uGv/PdBwMYS+AuNsdQEOOVl4ZJPOIZ3j789Pe9G
NOlXNbCQgUpozAbZfl3u8YVnMeXIGKfiltg2s3ktFFeoOgaZLiZRJUlqpNiINvrcwKhYLYv8a31c
5CZPS02g71wzKLFaQnC8AUAJQXx+Bp+YkhCLozST+h8nnSUXoU8JiJiv1KYBKBdpih4p00q4fDR9
A8xS0f8htC7siUmG0rHaEt9FAQIPrPVdvNlNZkFFk/PY5fEWNa5EoIqq+F7ssuU44ZdnDFTt5HDL
9i7qVT1ypg/g5Met46pTyfWZSub0xDtbh/cKOaoJYzP4OT0S/aPrCYIWvDE0p49lwb2mWUWKlxB6
yCNEy7Tm22T9zJDLZmTcEG+M9rUizTeI7RsOfu0j0ftqJfsd7ls4hzQiunnfwcA3zjBZl1Eu/Bkj
Cli/8P6WlQgiOCu6yv2w3MP3HmA4HjZ/ij4SuQdCQTbwNQUkZ8QlwbVNBvnsSyaR5+mggM8C5sI1
ucb1Kh/aYd2LnH8lQ0Hg+GEgc9+yF8fmZUoP8gAnX7kHesAHcLy3HAJPgVytlvbHTRzIRGka4AzS
uXb9LqOSfkwxlWfLs2Pt6c2E0vMG9nO4RfC9hmpx+4e0y/rrykLBW+hT90TiAg9Uza64zgrLVseL
ZeAcDiwF9rn5vNYdkOIPibqepGt+St0g9PugktS9zwGiaskM6kuOLok7cd5MGTD8uolHsoF2dMpE
7zB0t0LjfKT9YmPi2Wl8jYAsZeYyZkoyvT+wh/F0uYO4hCYWrrU+grc/jxK0I1f/O5nI+iti/5AV
j5gp2sLAu0SggeY/xGAz2pCJjZV/XV6KVprpg+xco4Xt96Bd/GczGhtmqm8mZuejRJ8oOc+sqbta
WB7mV7YRIC0R1C1IFYROueSAHqEet7nxYsNhBTK/oGL22EkIIDqSnZzxWaA+YeDnIN6m5Mj8BYCg
0+z0MsN+D5+UBwthVF2fW+DXQws4lUegvWvoAqKIWQQvgvq7B2Yz7fIw7g+0JgmuiZsW6Ebe1k//
GCfW7ubdjCErMaMfg8HOg7ju6TRuw7ScgbB2bctv3wr+V28mVnwyoBddb+NwliVWhU/GFy1l/c2w
bIKskesetg8PhwRB7CUgEFi2WHPy6LfSSzRKm94KkalslpBc4SHlEP/oA2YPesVwGOATmYYf7hTh
k4akERMlEgQekhZnzTk2gepJRDcCbkphHISWsIJyBJBzKs6YN/p4l6Izr6rPf8uMrKnzTcfz6382
uLyGJbLFkFQUDmn11TG8SAQTlFNPBzrFCzU+uk9NRhK0z25aaZLtF+OXdguJ5C529Suqugm8jl8C
L+fPZ64pPSg3Viyu+o63VCrMwVjhsBrCuXzhdGUAADtw4YmvNDClj7d6swbSXI2dYlcMKEY9BbjA
40XdJ1aM6AElE3ElsjpkUm+nwVwzbKQqlOBwsbMDpuE35jHKTMQOm0tduARrvgsPtFoz6z+yXeF4
Ux1ohbReOeg6MAY92RlsIaLfHuzsSKvQajeXjB/HgO1uYjZ1jCxCgP4KYcq7MW7iKPiTRHSLJedD
fNhqAmTLvLr+bex2ughVxYS/TqsS5G620w3lSSU3IpdFioCbKZWvhwCIP0beig7GA7d7vw5txNWF
Cus6By9lbBzHOMerXcOIafjv/lS9NzldXOq1VjdGMGZL1p2KA9Nex1FoqnY5oWw9BrfkIBkwv3WO
DepBA9/IcxRBizdwdxP8aQVamAL2E/d2MToVnqioYzICCElQoseBsveEpnxWqZE/+aJr5sX6tA1U
5DhzWwraOnH7NT2tGB4hR0PiBVm2xclhKTMQ3i1dUfHQ63atoSw6dVN7K/tK5wsPzTsIUbvPhdLj
M/a/tnVbxUP9VHiHLXDwlXF69rgMuochj3UMNPFBOjmEqDj2Cvzc8lJ4vtMXWHb0HTxTHglL/5J7
hjmq7o3p8JromBvIF3Wvc5ndQyPG7HFohwbaKnJ1czL2M1+oY4BlWaZtdgAmD8ledXkI8iPyUBh3
s9w31KaZmo6zehHlVAi2CN+TxlydtKp/ivmJRHKcQNyaqSjWLzsmRFWfEd7YR5R6pC92WskIadhx
GxRUfPZfFJp6eVl+MXZXNAfZYg5ahSglQYKzodOgbJjDI6geh9SBo7kvx1z0s1CTo2w18pJ6rW9y
iJZQOSJVIP/t67PNfZWZt2WFBIsu6oXsr2IgGZzIPwFGiK8fx8SFQohrA9x5MbUkfDnstmM59TVu
SVt9FfxEsB4HRTmVP24Hv0ZGaKw/N96uN/3Uv0OPC63kp2bfCV3ChHW4DrBx+u77h6IW3OjExXmc
Aowp57y4x39j7b+PcAe9SFD5MABKEc79jpIv8NnGUZQL+FbvztDUmpF8undgrrmm0p/TqwhGfz1f
n5GAxsspPPZtcYNYZLTNmmpySKQCMJgPx5Wevt48RnZ5Z11lOA+98rnO8PK8bMqVmqvKe91VImD1
AAHefLlLmf/BkEHEiK0l5ebWq8LA0/uI4GkveRnvpYDbL5kV/7J+sGbL3ZGqDjm2BLy5166qFxH3
3xNcseqeH7q7LPyyJ1xalNtowWbVe3A3ibypVoFUFlr4yl3zepFz4C+92ut6CxQcp87cO8e8+OG4
iTMmRVGE3ozQwvpmIyaZcLI08cab9wseC/CTphtgA8EoYodx+k33x0BncHCLYZnjL9dmvfl4E5DZ
ltPlT9cpuTPDvgCTAN6Cf76EBiIGjGn4NtwbKk90Xblu8PylgQdJ/I1Ud+2lHAkizbpiWohut6FS
XEtA0n01LbwrOKUvnOjiacL2UF3KedhnDcBWRGRfsNdktrXp4j0tuUX7WmmboSPiJ7SP3V9ZRFpb
pyzJdMGpRWPYs/I93KcKWLiseUZBqBASFDf1HegqFWBiuHtsfN1o99OmEfuHY+sHYvUtGhusOvtj
NqHv8aKsb//ffgXRcHVHvAz5P3c1z+KqxTbx3ULqHKilyUeOInKRSZ/zB8UG0AsUdqTcwWkQ47e4
YDIfMrEnydQ6hR/tDFBXjKahwJkGRXfxfOH0Trt86UphCmJ9u6JkExKBX0YyCNR7C1crXp/F3usy
wZTcCsZvoq/EiFD+NDQrFIy0bCWUDrABuR+oArV5A4cm0luCcipP2ouTAe9t6lekoZehVJIqmX/X
dEdGCYeodgHH7MwwPQDAKC0qC53mobuSsfSjlW3pP2sPIKh1ydPMuR+4ySmadcZEuaEH3bo0cgR+
Kq41t+s6/YvIu62/b2RKfT0qMd7SrHMlfAUD2OXDiUAMX4UjFYoVsy7UzysOgbWXazzQeHbiUwEs
TMiPOuICUV89pprPwPm/is1ZzLIIQI1BuDrBqpcRexbJDKdRNNxCeWxPt5TUWDCb0oPP7gO3jHxx
E9EX8SA+DaetDWYUHXa3okDfuuMb8S9Ui2sh0/Ax+92fw9pKxwJvexoV36O+sRit1vC8ZFcWdpuz
8Xm/KU74B9YvQW8wMn+viaogeRD0cXWjBlIFt7bkP9BjzgXV1chUVAMWsv/IydOyR8lH2E3amteS
VgAMDLVDmyGWgZGAcG/is5zmFj7WPYjvocnyQSeHXDz7+3MwxoWfmDimgJ0l+y8Xse3L0HVW6RNm
xnuMu0V0sB/0sVNXkIPYvn10Grnrh8Ct1Tk65dsnN0GZe6zPwe9h4vkBM9ZX8ikJxnWyBAb2qD1r
U+Fh8qgLRe1qr9O+QJpHuS+n7EPHNybfhvd06TEAhP++OMPs/u6pqsVb+ooVK+/WdQb+9lECwLHR
7ipKnH+WXecQRBx5owk/b3olJ5o4OmPJPmyug0KPj7qIuJBYUOZGmD+PzR3tZPJ1DAhtVbfRO/Q8
F0ftj2GZnG6j8g2qxF23DLuU8W0yrLWSGjmU+wakeRrtTgpSZA6gD8X0HNycS9q6ollxC9OE7/1m
WEWvN+Zz8KyINP8NO6/1f2U/5zafN1H1yhtt31r1/swB2FNYtGLfeF1YIK60VjfLhqRWfCf2ETj7
MxZtREO0SIeUPrl7lPYT+himOxv2v8v85Og6FH7juhiCvGriBfl/isplPVOxoVOf4u3zymBlqSLE
OMqpTKGnkKak4z4iW4o0yq2qBOsszC942/riXxlo8brsnRxFBYtsS6q65vIziXtgncXJ7BPjv7TP
g/KfHmBiVj0KMafM6sR/N4U1O0NoZhFvFHI9A2N92EPpwgne3OUa1xL0JFrzzbbrpnodhtUc4Rq+
u6GRASKYecCZ+53V9vp+LBdzN+UncGF94CcegAagBIG1qstVOTb9gYVikaTppOXYYlSuYtT40bIb
nDZdMO6c9vTIsFW6nC5MelUg1GugLd6uiLWVl5FdQx8rHWSEbO5BIR30l8jBAV7fo1wgWbLNPMie
ZTTVbr64UoQO74Gua5+WnXujULLOIIKYAjngicCJgI6RBSZ4QUk58dIYz0ZJNNl7NWRAjIXG//ir
dz6BAQyPuOxkQwrH9jjFs0sJZ7bpbjpVANFpJCQC3ghl3PCvOJAjv2p61Tgg+rsD0EHEQM9dMy9D
z+AUNTIeH7Q8VzNtT7Z7sLFgq1GGAwz5SPFoExzwGfzR/HxeambF2m0QpIEoOc5UGxwFyjo3ZiKq
D6fHVAT0Iw1kzvoMJduzoUki5pFLEa4R0IAeNYxe2Uaj+4f+e8YGIKcXUHjVCf6anybzOvkztpzU
Ifx1FfEliKewPzim16HqoXjdYa3ybaU7UPZApmD+TYWQutKVEmx7OqanUGLJ2wjmbYq5msLxALX4
iBuH+h5YeARIF9sFa7Q0JaCwRPWx1U74SuYr6Fiddo/+qxGwx0RPKnc2vLnpN0jaTqDhW5e6RPGI
k36Bejj+h9U+MfJzhI1Qe/zscMOK+iVVtk4//ZY4ndbnVQlomHEjhfn+ANvoMluFfeEXH0BmivPI
2djaQRq7l2+adQNyciuASG+snGR5opnJKgaeNJ16+YluzH2DNwF1FgZlhaqfE7uFOS4amM5qIzXU
azIZl/Vl7xzqaSrqql5yRCem4peHKU+Ee8E1yShaFMiHHfSQUdUO8RO2FhcFUpVUuZeTSJOIgkCV
q2TRsAdNs0lhBB+6YMmepppSZ8FGpoXHQPsqm1FVO6g23ZAME8PvcbRgheZwDsFhHadoBGRVdYj6
okeFZPe/PhnkV8oICVz09md3XY00ms8f4dAqXxCI5oboNjrxoN17yW8Ykzb6sinOWy1TsSkwV6aL
O2Zr+4GEuLvupS5QMkcNBwpcxSMAuBV7/O+7qN1Apbbjj9PpAyMB3W5UpP8LED2EFCFS2Umt94ai
LuLnxaPozkoomVKgL9VniJzaRXlWJIz0oszvEDCaT1Nx7JWmrvSpKTGhnztxKjYTF/DxNnrxBCRl
vOKWzcT1qAKGVABIeZqCkHqsj0RmvRX4yEm9KJU/XxKsuhIOTspvDkbJTYpnOXhOFmI2tpAnyXqA
553uRjsciHEbK2ern3p1POr4EEuCapN2MagWBPQh3w6MyDxr+sQ8g5J3M0eEHn0r9Z0nvzEw2i6c
1LqEGjfiP7kvfllJuiYNxYvc1x232u9DRJu/OqYoJAgpBYfsh+fZR0CKutm+aRHnG3mXPeCdRiCr
0QMTulgaMtHF1MZ1cxkueYZZbcuQ3Ys7J17iCcptvrGG3dQrVMfBrfcHOVqEBHnzddboEU9mPQOR
0ZVwc+cpO1t4cstj+nsEiDe7xD63t9IjkT4NToUyYeSe8AeHmU7kQqG8WzIcb5AjTtfWB2Ymgdl6
hfs5D5ypP+x0UIx5G23AWI50YpR6i2TLCl1CCOO7BwjDNQ0w1G5bcJ7kE4kpotf4gvKxKdtZklHS
KzpA/PzWMYXgVdLIorHZT7PHnpB8xfPmudi/ZjZEvgbvhUAqSOPxyzyXazYl2UyUx76ViV9hYP18
Irma+nbQgVldaRUs0zJ+n1unATNBGsLJayjxzuyePU+1/rZ/Myybo2Qy84qwP8p23udTya+QhxQX
+bvwyirZm3/fbltGr9+C/2Q3WoE6BO6Zq1aOVM0vWu+LDMwp+6/7BBOCqxl460DxGU2KOb28ad7E
YEHyF7mDexnCarkE5afyqMFTWdcCtt9k3rzKijgPyXgetHwA6y2WorOBo0fGkhy3uf6G/xXA8fDI
chB0rNlI6oPnQHgiFAb0duHbi64DxlJH3RNMX29VpOqf9e4ASYQBUp8Bs7Q18UR+XVWJwSoedznk
rW4rcb/HR7/wPiFvm/yUlcnROmLRin5u0ZpMl8jBpo8yiD8bETe7HYxsygbkShd5Mu/XVFf7Ov3p
j36WzWGXePdtNoADUVQrj9D0w6BLO7gZ9jhu0ExdzOrFgyIOH2foy/wCB6pAU9+aZ/Tod3a2QVsx
weoI0NodzqcztdlmCwwTOEXu6OX1KFWwSHW658FDHOW5h8mx0HieJ9GXmaY8FxM0cQa9lxIQQLR5
YufGQe7Px++4K5jXUW3pHAFRJhfmoT02UJ5OxkHiojIbaworcQrncx5gW2YPN8Ao6VI7U1Zpx7bi
CvP2ikE0R6i2f93EHC0NQEL0Z4AYVI7viFC71eUXTKibhrOgHK6dGyLUEY2Gu4QLTdlb7y1cPqwZ
UMH3kPQP46bRFEtAB0b4+4HH5AUwD436VmNKLu8U1V1EU8/Y/tZQNDLEhnJGLREgvWfrRJsNL4n4
1thHm5CKtb7WPbEydTksSMkIFwGvl9HzRqdEXQ4Ixu8Ys+IM0qK0ST74AKRpHy4DBfPAth9KqgGv
S7XNFMAo4fqeqtvl3v6KU+aJcGrQb4ol5Wa/k2fH2Wsgl2UaGZBWsswoZnzF4F5wX7S0wfD9DtyH
Zs3xp/96Ng9qS5rx7Llep2v0jYfRpoB4MmMpE2jinkKiRt/gtkvvrW9Jz7N/AaTqntvWpLQ/WeUj
yJ+8zWXpp0b57tRoRv2zH/8AyX70pYKjJlFPMx0Sx76eyFCX7P7gAzzPGfdTWtr2Ntmx6LukXego
oQOAO/8JX51shDH7nwR2osp1KcFOcgr2aerQVunfa3lg6sCu1FP4KilG2TnVoKVfVwn2J2PTBQDk
Sz+Hm3NCZYycC6jodBY6wiv2hQ82TSOJsX49Igb9ePcvlRdphPkQC93quLoR1PUqtJaHxMjn7F18
UY8jNVkjEcSKN/1KBACq/0MpUUX+P1Q/2LVq/nBxtK9PXAP3kT5nGtQjN5RP6/1XdFBq3qwHEW+1
BQKZVXzcltnyd6UYb3q8TVz6uOx4/rUHB93sFWEUbxQRgywJeRsbUGzs2O9lmG2YaokY0u+haEV8
HEmFJlZuzlvktUQnLk+gRuvQR/ylJ5AYZyvk0XxRVLSkWgLhY2FmigaxBF2OH7hLCJPy9VcbPmqz
PttpZgplNzEItb/qK/acWDhbmbzoMxQtsUIS17PaEJLHMIk0PunanhjC6nvb9DMpenr98AeEfzZ3
SyAMC59eZD+PRFfB4PokhudOs5Utxqd17BdsaSsNYuZdlndQuntpGhoG8wWh4mcF7OmaJj+NigPn
6PZPMionMVQk8jINb5ZWrnsZHCSMF30pAzoq7gm30UXTwlvGGgGT0iiMAhJja/meRAFyXKT4RbEy
IAfda7C/EvPEySwUwgotjQJDW6i544z5zoSRNF9dS4i2WXGgrbHuEzuk0Yz/jLDqIVqBBcvcqWuw
qTsQXOc864mI4kkMX6F6D1NYnbF4O2POIxDs3XieQNo1yiieldgGKoEEiO+Q4Oq7+FhdAcXbAawu
UOmrT56KdiI0VSm5rzTULvcniGEzflnoPVxl/8rRR8rFwVQKQpmeCs89qV2P8EAPJ2/WnQRmgxik
ACVNeuaSyEA08HFAbOV2bAObe7EOZVz3xy34bHKBuWBSp10rmHs6laRVZhhMy8kTXjMjq/If/eqC
ztJgU4FFfT3d/YiFG6aSmsaBn9ypR5qLHTjaEADHaJWAfovi51uD07oAsaJsGzaGDU9fQWRFsHbE
cEueHVoLLehOrkmEeJ3zfUpEsApVCV4+MJfnFbuTP+ic6hAqSMg6YyIpdpGICE6tAF1IXqZApDFB
xC9nvi7BQjwM6/+jCsH+veHxa77qk/Ct4tD2AKo/mE/YDuW1wOpefU14LeIrNFRmdJ5DRKiMWSSu
XFnXD4KzWYmx7TsdhdLEp2bmvYEE3YJhekVBacHP70TukelFCUZRC+kmPaJ5wFO3qSi56MR7/1Ue
5X0juqrtTrAwSsUavBeNrtZGgb/zqElOf+2vfWwzVa2S8UyxlkI/3dhaCWxQg0ZSbZ4DWqB/VgWy
w+XtcReT7tN2eG4S+3Tum0azZx+miLRYldY1BkWP5s3vXLHpxksXu5CgKSXs8b1ec3Fdy8BJAfa/
6binFA+9Vk1UyrK9IdQT9JdG/b6hkRbQII7zoirg8XDoniD1HxiAD6Boyfz6R0otHrxUnUVQRY2W
iwZCJM2W6DNxGwdvcbZAW65UQ5xdl6UCRN+NcVe1CHa6PcsHLGB/0MSx9YZ/Tn+FFa1vjIxGj+NY
Qx6MAxBqRBvJcQtnlBulKAZyLDoMFYNVKPwMnhCTNSoGGhXRsyjpstxV360pquZyFnpf9cnTCfqL
HV2cXYN1N51DRri8CgwFnviIvwEdr4h8MyvNFwGngj/zbQ0fCNojcMbuxeqLLNydn+z0NxRfotD7
ehmB4KIx3SsGeovaGOSMYspjcGKuEbCXSiDRw6hfHxgdlDS4G69vK9BccuZZbCSzbbwYqIVa2YC/
nyu/4iNCBRCinHOJc/DjIkr/pnHWeJq31oVtSkLNeqc3zv344C7xmyqF6Fhg/esEdZE8Do6lVvFA
y4C05aLKP8/DUIhRd5/Tt8wk/ydFexDU5wz7g9enhbNZjLHCPV5q3mjfo0ApTcZO2Ce5bXn5CMF2
mK9xf0njtAzyI/IQT7u0IqXZZccSJpd3pQhmjEByDAiBxP+CHm6mCRn0w0Fctp4NQEI0l3emuCte
pHEzDyFm/MtdF63qybKzAUrNLKsfl3Qrk8SIErzvuG4U3xqcmZZSXqOrOsYXOcvujZFJAVkEfg7m
y6mQ6K2IZE+9KuRN6XMbwOjDa4NJXHLSnCGviZVDRqihqIMrAYrEo3gWqwJXety0YZqBIakRp2K7
UdTLwX89ldUQTgxR+a/0zyC7kDpwykw955hcWcEX9sgp1r9Zg3Ie6zCloENhj3mpLs4WSeYVd2Tx
qXwi0VHy/e2Az2dgcXnbZIR2V/bjYbWE/52anh8/4v0yMEvVsqdMp5oWWli9xth1QaD4tHsSz1Hq
3Em1dL5BqHyOBRG8NahUQpQ1l1X/MUVi+MA4lu2JC/hpJEeeWhLUfyLpCbONo+UtsBCtLYXVKZ9W
oqQZH5Xc4plY3DsNcCnsp9ME+H/+VvTIc/AG3Ijd7Ub8aKkTrK2r88f4YCTvdOE1IGDxzhlC//2i
zO4EehdI6P3aHOgaISQgBiEfHdZ2TpoL22n59TeFF4djVO9JJxl6B0FyjL1pI2eXNq8j2a0D/GFL
NEOHi/b7ocyXa53l5Hf6C0BIh61qxOM37JtK6Mhc4nAFNS3nzMVAv5wIU0ZvjZv2pRAazFqhS+Un
KP7uXrHBLtO4iccsBfhrrdDnjcMraudjRrLSu/t5mrhXd1dwTzcFgxwRqSjzQEQ/DoomRcybCTSM
b132ziYkm/60aCq5V3SgG7oda8TYInfVEsoRseyNuXZrdyFFpSafFShMD9MuZet40tcD/Uufyxoz
fwoxgmxgaIMyOe9qLNBQc/+sQZDA3FwxGHQQa1TISr0EDaDkaQbVv0idDT2+MlCTPzAG/hkV5bj2
PCwfN2VUeQUUlcWg4V1WTLEsqEWiJmY0OidQuF4slr0H38tZ/VPzExZ8u78v1oWp/7pEnWo44Q65
R7/W/8Nt2cC444ObnsaM9kNLQn98nDiHzEPGQeYW15Wpvbf8YuohXihvaS10s68IUyvDziTClpKd
vYdfaqM/vasConvA++k/YpnwxyQNEQ54dhwuBcLiPsee16P5DacpHc3ai8J+WnuTiWMFLqnBDijI
MRzHCaw5wTL8yu6nycboNgPuFNLWYlL9w6AVXbyv1Ae2JTgJHNs289Ta3ywCvISvCM9yJu1MYkEp
87by+8gsF+f1+DPenFNOv6aRgx6GZ4R5ackStqGbBxN+8wBBAT8xAwwaAIsMYdLwEIgG9ec/3+jK
/M923GVF6ALspImfLqqXrK7EqazGSOLMEzI+pKFQthbtFeybcLlOU/XnYlb6Uh5J+A3f2xuwWgah
KRuRX0UjWFJDl/fIVzlDv32A/1iFa6uZ03XtYsICaZ2WPc78tIZrWBA3BOOwTfv2QWSZlEu9nDle
Bd5RyCEl6F+g2PGJR3O0RK/CJcjHIq0HdqeKiibw5VdnX3kWAo/s88PPlfUmSZpDszuD5LlJoTvV
WsRt53OaAdtSG01Lyy7mmcoiLJ3AED/mKgDjGEjmT6HWInsSIULuqeCsjaGxr5PzcMh7VHB/bGs1
RvN29Ml1huZUW0YLcUYBpYoKNWj3GDUknZk72/AKjpfK+t4glNq3/CvzDx7u3Yr1Jlkcu0vWRmCm
xu8fhTk8n2YA1QnY9TCa62NBccoADu19qbEDDfHUm6pmXkV4vpVUjP51DuAI/KeHz85agLJewwwW
E1UJAAjxEgNIcrbMu8ZHUCZezNiwRipDy74gSgII52VSekI/SWuY94R+zoXnM65mcQ85EyvivVSP
TtnPfg9X6yfkyJbcBz+cYvu5DS5em6+pp81gmj73d/1IalneJnHfFncHJpkIQIlE2GkIAvqFdA0K
8To/DTxHX8hFVmJigBnbngupd3SmCtDAxPmQ4RNgd8V2pqsiA6UNe5C1vIhguV76MCjc09wPBOs0
HBK4qt5/OCisldlnkVNwBfxbX2lE+iuP+kRsKdOiAk8dnX0pxFJnC+jnJ6cT1C63MFghPsWf/R3l
xAmc2v/reGj0Q5in7m22cz0jUeMBasetuO6nrtj7mThTAqMQsNUmT42B+a1A/x1IeZqLLnQQfuls
qNyx48f+i/FGeQeVkeVitjoUyuiIfmbDEJQ9rYXW+ywQifeHDYzYwbblAyMArXsBECRqX2ilwqHF
1zCsT9iKo7kp+/cEiDPuCINxMZsCbwSCECv7vUwcVvczLqxL+twILlbTyF4BoUYYbxKOqNqWMtC8
zYjU1S/naMfi96TIJltn4ui42ECAbH6AZTDbYOAPjzpQqvBwrSyqYzmJQB0nntgVpCO7niSG3syy
SNucFgJVtg2XEZNrve7z1ptjhke++kCyx5RehKnTwyrMdAu3zBHF0/fWXJXXeAm6BW44S9id0/sP
Flz4BA5VCN3wALURr/Yoxlkmdr05iLMD63X2Bmyd7QwwBsU9zkMeg7QI3fltA4/lQbRcI2ENXYz6
+1WvyL5L3txJuiUUv2Exr5djSAqfvqmKjBX6PTRN4z+CAg9T/uqhUM5GT4YrqDK4xXh7tx6ZaUeV
fhlOclGbNcVsJYVegGcbjEG3IYioI3asK1FRqnZDJSqQoFZbZw1IoKcziz3O2E4Ry+v3hJA7zoJU
tgvInN8RpfAPqRyzDk73Jv7z6d2EhgDWc/fAap0i5jtTbIAXmmoVyO9kv4M8mGh2Jibtg6tx/taO
fCA23Lfv7BSEAm3JsTEokwba6caXYjLu+Q4iPSS/CwMQ6N+STS7sc7wCbLiS70SevGYhZamJ7ci8
n399x73qhL3HGUMaFjmRovo1GAKCkYEUKxhK4E/gXrOltY7Wdlp8QYNr2jl2i+7vI+EcH/rfnkMX
SdNFQSnJdTRm+JyDEUFj48XyAlIkv3GRoIMPdsp7KsoH/qpxp2Cuk1v0Wpo18DAg2KpNIXtrygVb
D3uQ0awmRRHRpf1gSArNGsLKFUbtPETJbLrEDUQ42mC4nz8s2kvG4jrIm0oQ1v86M5GE6/VvH2C+
u1t/Sf/rn5glaNTmJGnfwcxIhNcydpCjwcXsuh2FA2SXm31Jteai73F0Hdm09so/QUEFaMLsODsB
QlJUgWvzC1wBWt0h1p7ZGlljv6dhHnAgzhsbJ9r96A1ApyhW51mNSrL7rQE22qDqvrbOq5FKuYmE
aCxBZ2AoVFUVWCrhR/0QpVzHe9zEmKSED/1SbDjQHW2somgCmvq2Yjbxbl0vQRqtiy1hwkzIAIoQ
pUL1wP72FxbAAczdMYYcVW546TDSTmg18VdBUro3Yh8c3mgPZh7TX76ONsy4ZFXPLNm9MiEanKhA
uyxA/1EIlx1yhGCfAtVINiTaMVUp/UZFD4QbLvPaGndBDcdt6E7qYjyVdjbkMoThmUCr5iu927/y
OAr9PkidYApW8n7Ku83G2dLEaFtaJxhxx53KGSHSpTyLRX2lcIaETSPCaQx2MzYe2c1D5ZxbIS3G
FE+t+zo7y0KzYS9MECIL1N1D3jJMc69SR6yYZUN4EgKQbw+Xh1abUohQ8txrd0hAPUI3jsPhK+Kh
0A67Yz77qmbguHRtEUzg/aGDmQWof9NY3vTTxIQXfNi4zMxhnGkdtGsTU0fR5sKz2DMLeHFyHpeT
Fql6grKRX76HFoRVezXDqqWetT7z0KgumsWyPBFOxOpLKZWRgCJ+T2FpqtYkapa1sYqAuFr73iY+
4xuYwoZ6T1x06O8X4QDdPbe/GBFWBr7f05Ek1PeXzSQEBiZsDF2hVRpT/SAha0+3YNtMLF6YkAXk
OsfkYdJX0OaUrZx+Fz+KQ2h2vQpz9vCYrH5/+GM3pXhZydbLMomBVz5mssX6FAQixqupqhatClv8
O7L4kTn1HmudDkMpnvhvPCAzjSrDwvr8f3iTz3/8H3s1nvCGElsr+rX0eOrrylH74K17wMyWsTQU
mNNpiccQ0LuapApSwrzmv3bCmABJwxpcpJWEyYXrvLGWj13q+yBcidGvUw815exJ3X7oE+c9seND
2s06QN4RBnOGoshUnZcR9lmpPBLTkR3iJolMpp0bp4ILAkAIrvGauaH27HRszJ/piXMLngEq3u9H
KEWhKsQq02sAjA2V33cyGyw6hFc2CJPHdJ5W2Y5PQterM7i8rDtTQXBk/RpxTCDMFQwxuHCpFovB
k9tjC3ThF8H8liIclqi4MgYTlJmSVyQfoy+Te9Itor8ESzITtXOOsgDxhbKqPvqgWW7DzS+mGAHj
GLjsop5i+f7TxB9MT7skt9lGADq1juV3+l9u3QSsyGMA+9cXAfP0N/s16ZoPOL3E/n5K0CEMssA4
dNm+WGlzqjjMUlgnQN60DV4DzbtdVyVrORIkBkI2lqqL6Gh7ws02TiGktTdK53AO6QZmwGl4isp0
sbo8KV6UIUewuQJ4pC2p276i5b0B6o+AfeC4RlLb2bw3igQvpPsqKcRkGSMoDoBE78hLsUueMMTY
Mg0817wKWeLCdrvnD4zxhzScWJ+pgFdHh9Pz9XdC21eUccbycy9+EDBvnrax7QpucwsYm2Th8iAc
Ol3fAftY56dmSIapQtW5yQTzBoJiOck25+8bKC+gCFWv+j7U02Zv8a2aSV7x444K04O4+QNLsX4A
TlhuetnwqYulYyU2AUXVStl29ld34MnJzmuAolnyP0lSENNmuV2IC2TaSB7rKX4AGBVX4qwAGgbZ
D66aczIFo8r/ZV7846h//MNcy0n5VLL2IZhGba/UZgyoFhzBmERRRaLYkSFRakdX92dzQlno5/7f
kRsIL/l7UlV0VPf78SwwfH1xXjTifCO2ud3oLZ0wyExveWeK2oWv07kxCwI93pwBawbMkJCC5YXn
VYjmwsimixg0kI6zvqFx5g/Cpr3TbxZowOl+1Iu8KCMVYv+zqdE/sdXzPRJb352YyHUMQmnuP3rO
8berkcj7Me/u7pEgJJwZQENg5ZhCxo+wPMh/gYT3fMIeNSIgvytNlTlrE2ZnN7APSsCGLNcbkORo
LOgB+kA6P/cBMvSa67NOpBR8zVcI0I5PRmymfoFWAvLV9I+jpUs8V0a8s3sPIixh1wiDpuEkNUiJ
esuauexC+2FdAfGvg+OEKIBvd+Y8xAYVWeDrqH+N8941t38X9BkKTk1PdYtOxrW+9pYhHbny4rBk
7illFYgD85HCXUSU5g/UunSBKxqrBub5IHebAIk1ZQElKNj6bqbgAYRnCyAH47PzRApDjX7mD9FO
QM70yJmKBX8Je63hTQX7hLh2eZYSkMJAuNJ5pQXMmBVdlh6f1x3gaNB0QUG2otg7a0+RSlsNwZOB
MSwTSNWJ22yHBqcGDFqqTvKLtXbLYIEbTJhtbdiMQEG8zyZsD1Rli/P57G6Ip0OEcoEtxaYCz2JH
7PlHiORhnxRriq1CqRgi9h3mxWoa6EecvhmPmzMWJ08n8L5ZnjHB5eRzzHXjEE5FU8NsSE/awqvJ
oOYgJngBTyQ4VuHlFT5kuKROtYdJDDEFX5DOaBbVVWVizFoM6+VvYNyjjGksROa5mYfe3UJstugM
eAOkYclo/dLCcFajTiWBqs7yk6nHJmD6hl+LvInarcO0x5oiuWRZuwq9+ur8AITxWbiqWPojyov0
Bg0FC0b2eozITcFPjg3RQgiQkOpaaryUZbBm5jIZl29QoBfJJjDLVZn/84ZFjvyqb0HGxhE4HKUm
RoEbzXU34UASGRRzygJunXoGutz1E/2oA+9PxNYS6mzkNrEpUaXPX0aZd/Dqi8D8jSznZvYoVFop
3Sza9F9J2paxis/YGo/lyTy69tPo4Sd5dN+qGuI5wcPgwhNVfm9C564BQ4V+GVgG4uIyHe/Av5v0
gkk6bpLqG4ta/zzhU2gUkqnPPvH7NOyBU5oehhQxIdXiOYntIHtfaKpXnYSODZTaCu/CIspibdPR
eriWP689vWVZvDAsFG2W6IUJixWg9qpxHrQabfOnTL09cu+JdUxMaKwJhakiSE+r/EW8u4KocdmT
tWdmGOLPy8PkpZYoBXYrb/ncs2qJZLvMr2WihchsC6B8dmCSGLC5b7KuS9Oa2RPUW6eh8ef5Jamg
yRpWWuglFCjm89S0c4CZew1UqzQcEl/GvBv25uMJ/O1WjGzXu5+zSxTa3ktHBHODUuVwOHa5iSqZ
wpX2iMrAAdBZzb3Aih2BreDVoEsUh7qB+ynFKoiphJt048brjiYAN+aK/6I90yhS244QJIFM2KSv
/yHujnXNt02XanfA1wLfWyV4vUwuvpfyJQHJZylikvMsmMD74FQVToon0gxn1yKmbes0mFOkR9MR
NO3GNeMNf7n3/iM4ccFHTPxhG1h/zSHENo3h/b6RFPpp/Hns1hnyPCZUFr23Wfsy3NFY1J9Cauf6
cyu3mNYKNyHBpFd4Cy6tP8l9tss4bqFdNZYNJ3ltCIwb2o+FTKztakIQDCAfX+wAqNjZzEyZBChW
NaVZSl0Ah5YAXUz84kqxj/d2PF0676jO0vneVKEJx3xB4z9+z2es/rI1B+AyVSd8ZHzJmr51Fo8T
bLTgBNbXGZLu4DdmlwapSAFQXKwrhAlL2301H0Z1sZXIk/XVduvo8mUz3LaULvh0IcnCppEJSiQF
sTzA25R3I9zZupiol5G0ztJRderE2tcYchdMCujZsCkG2D2Y427RKbgG3ltxQBQ351OCMS/Ll2Y5
meOPN14ItVtx49nHth6SxMhsUwmZK/z9oA/+mZ4zJb8g8Ef6iAaE8w5ErFHk9qJzeBdgGkc/qKaI
R0I9oHtyO13QLG2a1tX6HpdLsBe0xFE2xrlDbjj9s0IVd9x8hkY09UTgNkhhGQOqQU1aNnfex6Wm
iq7G4uehgBE7L+4sPZJBvNoYz1kNa/6Jtv8Fl/H7empCeHJewofkqZK54JNg+ImRQprXqIuqcHQ6
dCTeg5C+4RjnRYn2knbz1gU6JBtYYm644N54ZYhre/Xz21p7JvbuXHINWqi95bUfFJo6fZxReu5G
0c24nlMqOdPY9oxPIz+xKA/PpLGbRLR7bT1csMjw0JDuy46xk4e1HNXZMaGGEbazlxRv+jSMNLGr
3weFgtHps5H2yUwcriHBVEEv0rspVMMuBiAJfZrodDSLS/HFmNoyTQVIxs0NYLmAYCMMk6DC0xoe
3MUEcgnaA6bqeqgLDYB4bWuxEpUMZGWz4VB1hffldbebY6mdcDaiDLQSrIi4V6nqDE9L+srPu796
vteZwg17FDOJa31SCywGK2TGIE32xOQbzEYL9I4ImV1oAxcpguDfuGszsfIOjEtUtkOcgEUFISeu
187dNigStKHnH6CO7r0iE7jsgf92mUUyG7B3ymNDF+mgN1bZH1yV9j5fi6+koxCCGU0Do6OiYkJC
Otv+ao67Ii5kLITqHmzupF7HVtk4vZIu0gyOz5zR4DI08J9Jpk8oD4FHSSxrV8lFqWFb9UquZgWK
AOiwVHw9CjvclX0oLU/iQ+AUE3s/eCMspQbJz5FS5Eko1hR71HqKMxyMhPEYdJ2TZoBNK7WJourI
9zIv4a82Of+EG0lFVkhsd9iGlFeT7e5loXAHxW2DYVwQF74V0XOYCuNzCScSOYe+dcAPWue95eCF
M1WYEgrNiz4x3Bpt51YlQOMZHJDtjBtzSju9J3iLtxn2ryUthYgM8jXzCYbzoHDyimeQZpiig6dv
9PRUKl6WV4JR7qpvytAfMQE7WRwIj80/ewc/aVInGRAqaeyIKKe4TXPMUjxHclu8HG7IGbdzoVuX
1N2Cv5Iuxq16tnxbo5ZzHPd/I8xxyYkgmgYu4nAo1i8ArjdZX4eolUTMuZ6InAbLVKqrfAdF6Moi
98tBMIH8dFyG4fXV7MFKVayxxvr79tM3Co4cvSDki05sKk9tTJqNhEIP0gRT0aqMGhTjdiTogWdb
py6GpzGlNFAlZvhuJ92bV/BBJO1T/lWj0bHSXFOcTiQO20owPKeCuRkqUMmhzY7Ya1Tq0QBpJZF1
Iz+Osaq5Vb9TrbgEtvLi5vlv+QMNyochXfWFlDYtDgYRzFY69rf3MF2nxmeauicE+3kYguDYFGbH
3MQQAimNs00RSF1Hy+CWFyi8LqyJJiBYv4/OqjpP9eLRNOB8H5PpcVYhwcURosHHxDBNzWho1Cp5
80I9bNE5QaRDRrWHXjO6OGeTeHcG+qCWu5LiIZMYWS6G/EX+d0QMQMo8IovWnv0PGP0laY3i893a
yxVa7z9vfGKblB5YHIhAqCqiN1GZhwV7PJE+9opJL/XZpVAjXV5DlroYSH3+ezHCFYtqlpjzlGAc
jrsVxu71ObFF3uzmrMxYtdGTPRzq0OAThcyjkZMevZgIy/fnrLLgUTYcJ92mvVDkoJFvhvGF5Iox
9fQvXHF+kfTDDnfAeBhB50YQyXPZndblwpRGSPOSKV1Pki10gFB3seaqGMQdL4NNPojCQ80Mn7dh
0eX+qEyIYmLUo09Qa2gF8S1Ad3rcFZEMkJbmnhubdsgCo7uHCyL0y3aAcRmx+qFbqNUEmthrwncZ
ATRrblObrxdbeHvpW31n2UwAlxNPszl64+C+RfMf8c3A8O9a9f+RyatoSpggGjUG5u/DgWsDxXIN
JfIWi3igA6DDkdTHSDAqCyTb04SpgLWdQVGp8tyQevzURIobroQc91zXK1SvSa4ievmwWok6TgzB
Iflwa1+01j6ffLLesQAbtZBvtHa6vLmyTH16o3wmlvhc0LhgDEoQOxuNE5jmLL93NJZVSRo0mSoY
wx7KxfFSMRjSGfcBE/YS8UnB250e2wgD3ggLj5HbThplz4b37Cb52Hsfv1QMN3LtQz9HvrIdBi3/
7mG/LaIaoKYQi8nJDrxVEokrFk+CH8t24ivd+J8dz0EFsU/bps4Rz2crGfg000RwWZTQl6TJA/Ts
B9DWjtGkq47Dre/1Oem4xFz6YZDe3RYbaK4lBuN+V0dbQouBClAZI71X1tWhO/zAAOzvVG8aJcXb
oc+rn7sFRZBOgon8JoFF8wpBWKUaOqPkfYK8/e2ITV89TeTGyIgfGuJxxzUDt5b/TW/SvAl3jR0q
WAigbX7LdlYmEVruG2jOIez9Cw5B0r2POp2l1IkD5ib1l1jXeO9CgNgolrejZELwS1tdwnB5VG8m
QrjabdTh5fBtgLRwFs/ug++w+qixUcCl84kbGghFpz3dXQpYzAUaFUuFYLYpK3YlE0EDFvl0H4V5
TGPSZ8wMfGKc36tbVie3+CeHP1LO63ppaftIIUI6EImecNgf0FGgjQ/hwooZDdKzKPds/XydeS5M
Xz695htJHr0J2MJCdMqeN8fUXc5AX3ADbUPjxJrUfVFsDYeNK5Aq58sspgq9S+hyZEOUCfABsqXE
N5jWQePMP/TyPhP1GaHtBPUEMKs41iOofjFX4rCfura5q71ybnvj234WtPuN/95clc5v2/Eh6Qyj
0Z25/19u0a+ihNgKkYm0RYoGuOlIJ1bg1IdqLa2xMf/yRl4lqKo+bmfztOMTkV9dSGLQWdWXvvCY
AY1ppeN4UJXXq46M+bpReasM3Zj9PVvQi1jp1L0crcAF929lIMQJPyFIND2j0fLvQC9znRaN3NRO
6T9xcKjGXgFR15fLVQdnliPOe/jHA+3I/hMvvt4m1Z1DIu4fWUJvBDXSF6VPZsL4bxFkz37VrruL
4WEpprgnxJWJFNBDI/ViHWnIt7JDfxRFevmlBiQVKJ7/38bHKKADLal1PYaHQjF0C+S7HzYvoU7L
ATg0Lj8jzoyoxVJg2+aH3VlHE/DpPUnIsidINCRrrILf2f8PBgr4cG+JdE74cUgA6Wf46ALoKuoh
QHzTUoq6DjpzT8h3IBBJkvt82z/jwqv+Yjfue2aGOSkCD/Gnqd6bEH7tHYuUmgSOqvr3ENI+teqK
FcKTpKsb61E/Yf5DPk5k4sSyXB9mjdBbJq3AiSK25Fb+k1Bl2rR4930OtwrpKu9UCYKXCUPsXLSf
Dd3hX/7jg58zXQAVe6OoZqt2xq2XR0wUuNgBOpHEcmP2tcA0heNVi1lmFt55qm9t2EeeaUm7r2UC
apIhWa/mxrKUj1gkysEw4c2g7FJhWBUHEgAEvSRqLUMYODYLU295vDQmHPJ9pAMNFVGn5qblEJsX
cXxjsTQ+WZbiqrR9fFPPkfui61ECkmZ3RKMq/G9HTAcvaGkB1qoPpVZILpq2JV2BMmepUze2r9v5
TrCm6bOcIp7ChmrJZdjq/2ej16NHKmQ7gqTcBJSQevLh0rnRjceK9YxlD4JSh6KWxA1heQwkGX3b
rP8SzOboU82PNeKzv3Wg8dtmJFAxglp1Mv7Vr7VqOkRtwXgw++pYS64+sxv6HqPkU5FPrakaB1oe
/PvUTLVjJ7Xw+H+/ceo4H/krnhdfdBJhjkxOVdtlaWu28U0k9d7Tcr0X63qCPkS69rix4OoY6eOA
gj1/6YiA8TYrqB2IUskYKPfjC7roLbpwFIz6Ll39mBwlUc0QBU+XgzZ/XxiGqhDMp+2xKHMyOFou
QdUz6bZSLdszGJZGP8Jsbr1bGb5ZPmgiFwbQem0zK286oqCcraAElN8M/sh5iZ/di5un46EqE0AP
IfB8MODZhQ2s9uhHvccYRFfr9GFmxECMPlWE1ALX+k+XzWfU0NyjddInBq7bX3rJjYjpieDEymbt
3P0yG4hSnl9HdHpBBASjqWLo0A/nwMRLkT9O5IAcxC4BtwSwuSv6UbEhUrdHj09nGXTjOUUVxqf7
lAnIBrhajRMbfWjonsNWZJGiJupqkd/eTeviwUf8LHuyzhsYUgS/8HmS3bE0YdEzgJm+hhvLuO4Q
okIxEVAw7DBh/CsInELuRUhRP8E5YsBNBNxKBIaknNrnEOszzrdgl84QIJMegSd9KViVeVsVsiJC
xF21k/oLN3QUKcw9B2qbCYmez2ZjLGWoVjr7EftBjN6GSs4bBwkuGE8mV1akjeNiRFWIuZiMjkTX
fALro9omNgWHL/ZA2/BLIwib3SvfUfdAu10Jslj0Mv9LcH4ntg7M9MeUUHDz9WngO1dHJovE7BQl
Kule7W51YFYDg9XH+1XMzTvf8N5B9mn6lynNA5+iZFyTV3WXmBjRHCAN/O2bSWgpS0pOZTLcJi5E
ZLS7ZVyov1QIuskNrnnQDpqhMBUT5Zq3LzbHRF+WCoBtSVWM7mV4dDy5Rd5U0QQI8vjbeNfTf3M9
tJUA/UmlhnhHhbH+OO9iVoLNqStzlxNIVDmSlPxRKDJmkIQKo2JjiYOYLTOytz+wj8yMDx7gtR63
ScXDZXoXzUK/K/wCgRIbMTFyW4vFbszS6Ez9vOwxEdukNLwoKMcK1ARjb/4GOG8K4QUIH+tYUYVs
YFkc5sXnLBuiYjNUwLGSE2slALKKMc34kyJlJZptMyFQiwgrPucT7uj1lkQsMuN1MvNhu9NTkPY7
DOKtp9c02dWuzKD7XKCeZ5DGu75F6nLYuYs01j0NeYwrnpHOYgh9dM1SaJVrBPqP0/2RdfBcEvSG
kkIwyXRM25NrQLlF61bAjqf6s8mSiQewLj5zhk/SLBcW1+9AtszBaEMPOPUishqlyyv4H+XVlcDS
jol6gGk+cB4bYKu0vDrEQc3ti6ga7YcQ1WMqqEgRcPFJgU6tR8pCyAxYizK35YVzxabMwlu6xSRS
xy4fmLCYidDsj8yHA733OSimDn4UAPlfZWawmL/BsK3gnQwAHEyiWHkVW4e4SWIc28xzNdQ6niJD
1nQFsFBmcyRTJkV1xplcAj14ABF20vzY3Djg/X5t3QRNu8PJpC6UsenS7Jp7auKa/TQcgoJ8Tazh
RUN1relKweDJfIlIcxw+jy4F64MuT7aBizZb7q8jS2ft212nGn+CnFyi6QoyvQtiC3qfpr2sy5Mu
W7TQy+3brjdJpHx7wASziy5UgN3/wkAN+nI7UfJTv2wU7HLR0wwD0B0jxoLmNP72NMTKMDPEsopC
jEFuQRUGeLOKy+R7jeM6YI7CJrYk3JFtoBAN3+0VeJOAUSwrnjM33AhbNlryg+24UFZ4DYG4E83l
oFTvw+Ir4XvN2SOSLYe4BESlwhUxYbRdJj/HLZXqeIDcyrGu6RcOeK9Ko5RNlU6zT+08vrAJJMVp
8cwsiHoMKY19DQhsKpdvsJ0k3xCssUYeS3oIqHPqhbf3LYuqE73ENVc673HF6JZTrvoplw3x2pSZ
IsRh1lx/4uoKrvOWYJRzIXH+ScVAiaqI+0CdZ7pNWK/o7v1FrswVRHU+kOxdYNGduNwHu82CaAP3
bsKhXCgxxa1Ad6gS9UCOrRybdsSIM2UWvhdvn5YS1C1FE3NVkeDxNyxWPhxhFE8qD1iPIRaiFUNs
hovy9hMFOplRLPzUZn794nIYYqkuBU4n9+zMWuytr1OoDK76bgNWHI87KyD1RCMRp/RPkBMunf0t
z1Cc1lm1wmqVt83HwB3fM9gHWmasx2niCWB7QWJsKoNi70MjSawdQYbrlxxCn/kKigDM7wQMMBkD
2ZMdooxpVLIc9sWvRGpIVAlENQRP6RWFxrx5lOiUUOgMoTC/R30UFc50bRKqav/uRSvOofTks6k0
SPBSB2UuoiRpTDpQpHGMHLpgm2G6qk+eGZ3cpBt4iHgOEUZ1EnB5elSKVzb6ILBaxHZfizjA41B3
lKLeoAdN44+tUXLkNPyZzlJtzT7pXryq72pghKYz2zM0Voub/OJ3FO7KXGQDgBClVjMZz8CQqJwL
c9BRhDeMRF+iu4HAHgDlv1h8TwvxBleRMj4KdLJ6th8ctyVG+Mx+g+kcVHSrDDnO8cAxCIHUVZiL
ps8fouKhct3pPaRZWayEmd9YZR1L/itg99ITm3cTLoUb+76byRER+I3bKhifp0ptarimbDI2ld4a
x5v/nLz2Le0Dfx2WFFm2uZ7Qjswwcf38BXLoU78Mj6vn0AtO0eGtgr0dWggF8ge3ffuK6nSZmRDe
copPHg9UMrhwHnvHh5jdNWRbSXuy95R1dRLHnNCWIyVjycht/URDMZ3ZXOWydkruHmS29xdqmsSJ
lAbTBOQxK5BKxnvnaGGChpYyM0rCb75d7ekwVRa9FHAjftU0lx6Tqm9Jy1Tw4FtJJ5FYmMu5MDjt
UmrtZ17bjl2uC4lqf/QPDxzFZzdQxnjpObR4TmY2P+JVzog01tIkEP95E7ezPnkIip0EJ5bj4Lh/
T/XNOYmpJm4X5lr/GHqWebqSFYkuwIJO6zttArqSH08oxC8VemejvlDDmlTn7c1hWfG3UUJHS199
A6kXtOWFedvKWvgjMPp4qLr29qUkxEgX7M7vfk5EsS0w+PwvSFoq+NX5lFoQPKfqg16AC/KfNfrg
W6OLjdIJ/AwhjmBFW7slBhbnUOE3OJaiOcW9e7hlwo3JrvwY9unJBAyHtoUbAF/3e7+46iH3RzI/
DhGjgWjGEurLEa95LfDuQWwj9V9s3vW/61B9Lh5XYcrfaCkZJ1SWBbP/KPL3m4Y19f+BFSL0Ut9G
G0iXmocFwWQLXrIotSx1OTIxcn8aDR906PBEneP6h1wv1pnLzuX2UW6dmNTaqzPWyq2p2DnRbwID
bz2V/AURxHSONKkDxk5rotcOeBEeK6oBGJCm9vjZNSHAh7b4bI8j9esGSebqZVctUou8bLfVoYnU
Le+Avq0XsdjHy/2DoUqxz9GamDmgCt/5Kcky0kktqYbizr6979Ul0iaRXxeVP7HmaXERW+79avsX
X701yhWv+AX2aJUvfdzG310x4Jj22lmUr76k69knUQ9QqKXT26Z0ebquGQdjxbuFD8NfSczpJqla
PQYMHeQFCP1v7MXZxqsy1g37Ln8bXZy7qK9yJAqxipFeO6WC8vjiombVVfaIaxN7yUcLUskJaVEH
lldO6U0i6WZcSIHFtsoqhsj7zAug0O6oVhO+4cEEeV6ppieaum5Bo45aS2uNKvn6ZXUpdZXnxrIg
egG19aQzd/fq/sup0h9AogisWgJkC3prK5TFk/KhzpYTwhM2gGDrSdQ72oKfA+idA9leU3dl8bCT
oY4IxD0gl2YVkrTYwXYVg5v4AOdcvyXoAMLbP7P+6bGYE4/pCboVKubhAE63Ff/XysXMkdieW5CC
VXcqZWFUHAZP9eEyMKEvXnw4s9WZ1lCKlad28IdqqSKs+3wMiPwahm134cTb7SOG6aHIPZb5vxjZ
Q4oLc+LdW/PG8JZ6sEc/NYdggMllqQPTpH2+CbarX/Krdzk84EMFFOq2RowwKoK4mZ6M0dKFdIi0
FAAfSTZD895uxcvHAIJ7h0qNSmBsnpbASsUQu47tm08Cff0qYb4hqZS0jkEyBTR/yYx+eK92ctTj
+UbcUvcyxmx39EGANv2KxxbUlsN2+t33CkCv3IRya08IEMCviiZQfHAgMpICD3Yz4FM4wnCnaztm
VcV0fYqTp354Cix8nY6apQdSSwina4fNPRkkj2u+jfIlKwYTskCQ/xY2ViF+MKXZdC1iFJFRx2g9
P8t5cRkbc3/NGKEvQgQvaTWAw6/M7JSbH0w9U6jcWUGTD5nlGnCRRb7MESY3v0EQFpOvcr3n91mp
Tsai2Cc2Co7Ky+WZXEMK9BcLCPYZgXgabk5w5eMIagzQqIY2rDrbf8pUjjWFcmqOYAxQxgpQhKDo
YjhMnFCqLY9a8i1P07t5LMFLHqS7QbydvsSfkALzX+9D7i28gMcnYfW096gadmiM764rn+94VG07
j0ibMUeRBHlExrscy2f6Pa/zqL+NHUv+A2UwZ0qjDxMSSCSw+i+qtKm1/sP07MafNM6iqyojqOcV
BmDf/wpBcWa0OgoJKNdDyzJ52tBfJ2YplCoNmLlwdYzV+dyhjPEO2Ohv26990iEfJUvuVtiBSC+8
ss5sOlDk29Ls7ggiMf9gCuetWMm/fsuvwgHew95aDoOFz1pApi8z+/rVqk0Sr7FYdiAyhDU1DyDq
nvennzdZqGcZ0TZBIt5+HzVOwMJsEwNEFlGUS9tOSIf4l8vxGCnZXn9fwXapjQtRkbv2CFCMkMbp
tz/EThiKKlH2O3bov8bhCH7ojWGNT81Eaipx/Q6H+pwACO8O308WH0AoXyyo7nwzDBMCrXKoDpcF
5k5bu+Knj9zhwPZngc7jAM7YNjFVtoNyxZcYN9HJeozFSzXfKVHC48BIR/u8KB280Gr9TQ6XkaVL
jG/Bp8dZOXD0yravQuLqrBHKeUPQO+RE4XKxGvMqzaLE8UcOktlc+8BtwIPJoPy8m/PGz5fQBHS0
rLsTLTBHTnvxKGlD9W21W8B/RvYSrUyctKMXgadAG4Gwe5rlP3ukxMRJWq1xqMrtGG0QiYpdn0iP
TW+TQM5zEzQorUcHru7kdgrl5vkMVsgmwaxD+thwY2Nau852LTDppMlKlnxoYuCG00H8Ex9Gf3s6
8bFvWv5iO57862HNEV4aThzUArZEsDXIQp30Yl5skkf3nBz+45PQz+ZRWszZHYcROt8vQeLrxz53
vSAMywJ9Xl/UiJVaZnVWqGemTJCZOxPhVMnB/SBS8VmweCKcCmiCeSGL/JYxNFR9UWcub64T1hL9
SpvPP/8+BCS3bFyqyr9CBwnXfxUw+ZxIQxjAJ6DIN7Sklona6qQrtqhzEQ0D5E/C07FjC8lOBxk6
sDqQafE2tXUWlO9DIGZUdoKl6A9SxreaR6sQm9n42Mw2lPxDsLvvUxU2ov8L3lGxzmhF5/WF49lq
a0+QtT+80TQJjXP6f0eyBIcQENV3e3PFjdjYAcRhK7GKy7sk7XrXu2VGuiwAIbY+XqSiHLC75vAu
51hvnbAtCLoQxXBlSAUxuOoQ/eqcISzU7SEUWEjpj6fDCw7V7FcqvecCiUPv/8YEzjhdh0dDyRHf
TLTsRkBQ1SOUevhldfXB4OCfb8TgHFsKLaKcrS4f9AViEUwBqxU3Z5neXXkURxSuQbdY8pBkA0Dg
ZMg2cs86QYSDnwvM84C95fPgz6DyDJ9xoY55zmU7n9I8tbCYTXA2pP4trBkvigpOJJZm0HqVwDb8
fXAjboVwjEN5n7l7v/X67EgbMRvcJxCiEc8/IhnKgumEzB9oUMIOinDHeqnYkw/G3X6BBOvfUPDN
DJ9HHpKIUguPqxg2Zj1ZHzHcpG5vO8JZtWoBS9GNcP3XEVxazMsL+G7+3Jw4kMPYj4NztmySZmyG
egZFbVB/ejeqEgaasguR1o5DKLkZ9Tw0+x4WvWGTTNupQPpa4zenXpQTddeWn+duqhBZl4jGt+Fp
tGDyYatvRdr285QAsBQ1MW0wdr2UYIJUarcLEGc4tSkNTo8IN764jNO7EAiYlOx3bFjcP5tIWKUr
kfjB06ldra9EDCOTxkg8akQoc5gF/2mdzz3kB48JrtKl/NE8eldC0eOlsD2zfnbbVQBwp7wt+2xC
l62aYJbIPZftXaBNF35bKji6ooiYvA26ucdbYBn8pusFvfmeLSc50HHXSjndaw6IA8xxMwhOuJzJ
rfraMWi4H5j/Ky05T00/Xvbyi473hL1FkGs3xjCTm5EDln96yEJTqF1LPkilD47eQ2yGEemdhnCx
Q7xiBlVfcyOndDIxwkLNivqNs9FB4bRj5629LEYRBbBhDqu14q2VgPHUXJiu+YhEITvIo9LN2xwo
pc3M57a+EtsCKNRGbQ8VQdtLOoTltTM0hxABgjjTaMGCehhc1gXptKDaDqJC9Sun4J/HxzPvXTtE
9lKpHx+JpL+vhWM+DXXOKIa0UF+AQs3GRnhhq5QmNfEB/E5uMLneWgOXAIV9Fkouj5n9E3cysWoV
xAuZuI62lffzkD27+5WZAgCpab3fqQzZIktFXY/uhxLSY+5Si+4S302XyjsA09a7nK+adOb4pRv8
QEj1BdFQ8HQRbFr8Sd0E/z+DjQ0HLr0FoiZOCch+/3k5hXI/wSfidwQY7y8GnSnuQnKJf95aX85v
FRmnt5C+9KC12YTj3qUCgsffElEYbNgsU9ZjuhuVd9BbjH3xD5sj3Hbe8JVRZE4yJWBZq+7aqg3c
vsJhOIy7FyAZFHpO1r+eFcapxUIOiOaT5TDMPIA4jVbo95S4RT0ZJjB9SGbM/w0axKkO8+3z4PTK
SZuPVn790eKwcAruI8n7oRxX2AuxSb227ee0/5KEruM6R/wyt/E4C4mhoJdCR50ZmR5y9kjZmLAk
5ibxEcvjXHO7tm2zqp7zYbuki743N5ReNdw4p5GCgLoTYCot/a4t6cxUz7IXcled3SQOoo1dHncz
jKhRmmRoxW6wph7/UvLBu5c+pRCGZvfMDxtLsSknXbn+LfzDyKY43w4wysGbMoZ6+noqGTwImKfn
7OLd2GD9o/Lym0mYTDxezsE0TI2Xkgt7OoMqtapXv6Vh1F7jCosXkEkFFEA1BvvWL8vRgquU0oOz
rPjNWZYB+FsB1fAr1V6dGedi3/zfLiBwtmDGY63vnRnCvjm77vQdKXd1690N6CP5uKL684zSZ6+J
wLjwE3QOIf7t7q5vgnPOYq5+lkiUbKgCQOhia52anInIs/U6MjCIiUPRWaomZgpUMxaNdAWT1B99
ECaH5s+pwgSIsLgD+yj/VnZOfoMJLSDqMDYJ9mbNYkFbzInOXW8vBEzqaqTO90kDB2gh+GlcIX1W
wmkCvJyb61ROLZImy8FsDRS1Lklq9dMt/RgcoT7pbFvuLT6VVqkGvdoiIM1TVyRYuSGWv6F4lkbR
1k8I1z/aHSDVidnlPrN7pm+y7/2biKz41zu7GoNSAPrdivw1uyjWZCHMuwN++iiydFcRJ3yKnnwR
/HLKzh8lRL5Zviu7QiKLe9U22zkGMGgJfBQvRvLE5hpgh4Zk9pq4nsWiOdEhk38/D6su8rYxj+6w
pOaxa9mrYSjGqZt3nFMSMrBfgoIHBvLYJ8heN+JEBp0GDt/qEM05tBRCYkgnKAyt60WWW91pA1tE
wBqGKVdU7d1ccdmJFngDpFS3xvN9T/VGG6C5+Vjgm68quqkzdrxoAYwz/qWIA6OX7LfJ0xJu6Qbn
WKoRXXb88x1w+sfbbH8FGzRtiK6aEqRKkFC7pVTIKo0ip4e0QbLVyQvZHs8+lj0qcniVory6oRGW
kwprP+Z8EXbfgar4AHilj2dzmoZBim39iMdl4zwmkinTmFF2Tg35stlkXmInZjlWoOvSe15txIDl
kki+ANGhf9Q4M0fc6K9/VBliNUpPxe9gJxVOcfDWaS/tdiRHyWlSPvA3pnTcswrRUFQbiN+2WN8A
REe+4kvWNxx4EnPbRwabJcg1t4i3UtLEUQWtSO09H1p2A3cxyHo4EIP8pByujQt+rm4i1lOmOP2f
EJtPHk16loXQEqQw7fq2uDlY7i2BtsxaqhoLtmBYby3GpzmFKRMbaeXxeFPKS5jtJxt7kFlZvr32
hkjhmdEiaof1ms4x5FrlwjfEJYO7jdV4kp/xAKTncYAdGi2AmbtETxw71nzYoUzTC6vNcDdF8EDQ
3AyVurdR/nHR6B6jsqf3rfgkGAtDvOwxyHs8yEcrm5HkMlCr/dqec0EAjl8NwDcKt06GrO9tuRLD
+aNvPrzem+w+JfJozTg5sH3e7te4F3LZlYs/r1LHmfA/2j4WXmvrdKwJycfLpSiLGLucEajaQOjg
Xz2Om+4K7lkhFrBzaWFQhwt8DKvGK9X/8P+ED6D8vLTB2QSmmRatp2m+X4CNOFTT0ARl/ZkrV+Cb
pAar105eEwSPfvtVkoxvthk/q2gTG/0QXyJHn6KaFaqI4zT3MaktzZ32PF4aE2/vwa4aClL61U7Q
glfO4WGBRjUU5JrR6WhRQZYzVmTb8cS7dRtPuk25wwVgiL6bhyNkFIdLoknbWqyRg114kES6JyJ3
8FtHdDKOcgZIQ3tsT3wecDHbfShJ5ryCZEfP/PUY1tsZHE0LMTtsetFSWf70j8iLrLp6uRmZVtD/
LUe2/2tq/lmBiZ45NH8U2slC62h5eoQcpNpLvuxvrjvcHjUg42Z/p74kinY2OM1LlJo7l/JPa1QJ
t9wgssYMPIpSPJf1A36qOVJucxxGn7XO/LZSKFtWPLQ2W+g0U6kv1eQnbG+t1XK9w2HAGRSFdk8d
cqvBikiVqZYaUxVxvBQhN31RtRnkas181vofk9XA8N2/V7JcFGqc/Gn1wajh8ykEpyA433BxUmN7
4tsCnHY3qQmNgyxGFe7oCdLPBsJvCvLM7vnxUV+AUtzRQD9teITi+hJK7BL3P059NuPEbaXqenD6
pS9obay8e9s2jSlGkf9hMOUSm0fKjy246zWKhpbWqd45oVoGWvWiKhcJ2TPx3r1oBJRSvg17hjp7
p6IiWLb2k/SEe5tIHbkGlX1xF/opDPn0WUXrROeHnPlG+U1INxscVw3slH3gT/+PeEfKGY6K1HAW
7XC+xFs9zVmtz5nLTRSjAPZnouoSmfWfHQEYbec0MTpeYakb9D7TaDUR8bjJG3qQz2cSzD1qLP6s
MBncPlF59+HJoNfwRaH9UfHRbcEtzjH4LcVAK4/fGUPaTQqolHdVsyyvXt2O8cNL7GO/AibWn9Q3
Jx3Mq9XmDCLKD0ntZCAmVyj3s1xZf+AqLMmrcRweRj16/UglGNn1quFMnz4wjHxCL2umpE/QdFeY
KLfUyZuV7ODegQqgPZak7jHvg3zbHHF617RbpJcJIqLITwm3io20+wZEjgzJ9WFBRJSBPIhKrrrv
M4992Z7/A5hvRV/fU951vkE3wZNeheL+eFul5GnAH1Ho6sEmsvc2JX5/w7C+Qzwb7ITAJzpBdF7F
IUQgOA3WYAzbijrUrUSg/vOQkHG2iVk54i5ORFAW/Z/pmDw/wmaQB7XCygUjcF7117krO9YSOhd4
V1/dA0HQAKFRHkM8BzCCBk2t5zUtWSAfbTmmbpOC7+uukbec4Fu8ekrkmTsdECxtDFfddnt6TqE2
4Oi3nRsDrze5GB8QYzcmg9OdpGhHuwmM/VyayeqKIwVRv7zXr+5tTWjQIoO+Gheyiw7mts8VGwLz
XZ2FMHVy0aA2g6Mvhu3p83Snlrj30C1Wq6PmLh5uPP1z7qczaQR6pUUyR2bNkLqcq6YLzqt7f0ao
VdJVVPCBMAzfQsPPre5ZovGBIMnjq+wogA565anoFQPlgHJjWtHFoa5M21yr/uv+Xc8zdD+9sSEJ
569bQg1Rcuew70oU9zy4OzZfCGIPfLL4Ecg9wUViOFAyuk/+7Tsz0/WZ8pre1BFD9GkSH1BayLXk
JemayppJ2yhOnqx4/VFPgXgCzNh0l/VUnm0NWqdAqiyh2p4MM6JF8SgVhh08Kx11jPvHaoomW4er
vd4qMi+/NPn1zS7g/IZAjY7OAx6focxXbYYolrYHcBdcx2r+oynkopBbvHfz9nOhFd2lpZCm78gk
sp7sa0pCS4seMZQv8u1Fk5x+xUS8MOO2EYdCBYEHCMNwHl2Gs3ZQMi5RA07vUdnnYeF2Lvf1Hyfv
7AGuF95r3Mgl20AJD/h2RixrQvhGeEaRpir1iRNHkTeT26oM38L/rRxd6mmdpgF81DQxn8oWeJ8w
egydjNn3mbYKlztZPdQK84GZ/Uw3NHK1qkLrrRUm5WxwWYwlYEXc/yMNs8OLulGgWx0N29YFN+qE
dON/VM/rUvz+3HXXN4pDFtjabNEG67b+ZOzvBDxxs0Pz0sBW1ClsY56x47xaJlJpT4qDN8wYtjSM
XrViwWA5bDkpJ+yyhksdSc57dZmvJIDFI3PH1b2BI2dSDqn96GQ+qpmfStFNP7IoAPsfTmZP4Ug1
QWKyMvVkAdb589BgOz6PgdZo1ESOT+3wOKzur08IPXTUGZmDcB4rIopwxwIGyNjecEpqIZf6SxiG
MrCzqlZ5DVApoZVVG5pg7hFjCbEe+F1ZIW7QmBnUdAu9BlXjR2aK5UJ1adPYU/ryM1du6IHJwQRW
VZ/yAjO3/Eiw2uyRkWMqgKkDjTq+xVYpNDJchQA35o7fpkHRQtYsidPOaSVXlRoBZS/6apkf2hcG
iWIoFn65c95x+0KXHuIuFcYnFzdVl30VNP1OGSHJFk9IztPl31AsXPF7NBk3AKmkQKrXluPOQ1Up
6eMdFp7QN2XjbcIed3hF9bNazFIrRmsP8BMv1zPahM15SOvjImjRjgK89WkT8jxAo0/ekG3ielpC
/5WDbAmcfcSMKLJ8qR1dc7kVe5R+Hm6HXaXeuI1BqEySagGR3IXt2DdK0P6nMZqXafuWaJIQyoQJ
7609unD8RYIsqqtzs6SysrLokRk5HlldetQcEQ1vK0NR9JGll94D1JM5MRZrZN6eg3H/ZPq2OBYd
VJuOxd6Urkd9hpUIPfaDhqb3TFJGrRTx1zlIAqTx8DFBSjRylZrvhiWoKp8Kwc4Tlv6HWX/YRSSp
PstcDrBZQc4PVHnbTsMrp9+DwwZOcQvR0aR+AYUidJTgbCqyIrRIcLxpM2cj4x85uBW/QnOpzPWe
pguhAygl0bGDhslvMfMCFQg7ZxEGWH1jl4mZm6jY5GT/pQi9BCMH7FK8A1OppBUqx1ptEDAR/kOH
av5abZmIgWFm1dXb27ZtF0KruhNkkWtwGknqqHQkCAsuIBbGYP8yQ2xFvFyKH2P3VvTfLxOWZmxF
6I1z8we+Qa6GHoIFytyAYbGd6jP59qyO5s2YeUrRXSRRGNinNXQP/wGcwmqSNdNXQOvYDOf6jqj/
Uqsjj+T+vCdyPhW7OlzMK0czQ6ERuCP6NaWBJvuTx535490GKoonuIHjUczKoWSt43B2mKAMzeM9
bTJSz4MWpiVKQBXlyCihFKlENLYkwYJkTGZDjyagMY2r3qysXKL6s/gZAanvxeXQXZ56YHNIV55h
IIotXUvOnN/JR5F8kAqUdPySIziL+2s0v9Mu9mEqQ0B/HrIGJ6bw5zBUDnVTShNJIjD4ok1DyXtD
RF/3j62Zv3DvrOd4boJuxg3X2gpMf/2uzRW2YMWLZM9Hju/ReqwejNMs1cnAKlfyNMsnAqtvtE0N
buDKs5VzrRhe1oTbHyG/EKxUroraMItdMKAiGaOwEyAt9r0xjUfbDQCGMu7I22phNf3sUMHi3Ir9
jTbX/z+d+cYgBjIW1H1BNal4Rjb6ZS3XDNs2LYdkJdk8dlLoCrXsdqwfeY7i4d5n+zg68eqH1Y/r
Ub9zTZoGCHiXO9FK4kcNzJ+B0uEstxOU5JzvCinEMGpj0vgv6ufpJ518zXVpF2zwvqYiotwvR8Mf
DyrxJqmX4dBqgpr+uXizGq/Fz69F7uKPqKvZS0INgCUtHPDqFej3VYMYC0N8KSpiTG/wnmVm7alq
cfEN7wqnenUzNyqe73Cu6p03WJZe8IkbPKBNOs34AH5iqsBOwtRjTpUV5glOPTLWwA3pf/99yYji
/2xKzd2PzRtVbj8jmNMKzzqkYmp+/Gp9KSQ4mQfqrjMhzmgGdWQhh32ixsEfujyXa88YHL6fAAko
IQuXBD2YxjRV2zaaGiRZ+Wj+5NI69Gt6aY3CTqlbED7gCmkzse0dB1MirG5FXS51i0N8+kCj+KzP
GPdMevilpGywFCalULJh8GpvifroQmg57cPYgSVki69IZ5R7qydMGwDXBeTLLy4yIERLQOWZkSq8
7MOBvCxtGghDtcHPwoHI2VRzWZydWEFZ3xUBem0BYc7p2spTb/+0a+NkAOTKULgcWxNligFBOp0D
pfmAj7KlfEIfEe59oeDbmJCSt2azaFZvBEszNxi6TJX7MvN7NBGGD6mxDW6EwJsRV4OUkbENXAog
Vwn3PjSaSCtgF6+VVzhfBLDNxz9V9ocUj2z7IXYzmmyGCSNx47QJY9sN/e7Mv0X5ravDrkkxZXWh
o39crWN4q5pMaMSOypeKYIlcicE+bnWuk7q3B6DlCU28+6w5PENJBDRW+cRywnbCuAImuXRmZ7WZ
f7M+9gT+5uHx1XrnDWTfzjzhaTLWaYHYwugyvRr36wev0TPsv80vul84nDnPmwoy0Tmoxo7Le3pp
Q1iqWfsdVpLuAXCMdaUwkYXNW4fctYnN4/iJugGtgjaWX3WWajWyOyJJAomHRh5PSysXaM59c89G
p9JvT0LFUeaXCameRBrt978emtd1reDbnIFijR2meH7dHqguwfwkKjfwSOwvzPay7ODtSLM6dRdw
jAx8tAoO/RQG6O3f8HXNg5rY5BCZ7Bhjh8vKDNb5gpZD3S/FtgaDZy8l7ayXcSFQZuojhytxnb+Y
3y3i5Bn1+qteCd5TwTGR3CtXYvkN/UwunPwut6kZgjZ+5mYqj5sZ10A9eoHzWXx4WWMKXnGoTvRe
hWP9qqyPA8H2flfHfdq7Q2sccI2U9IRYUqAC7VARzBYinnksuHdFCxOx9P7oB5+pvpuuJ57y4zpk
aurLAqid6VYO74TpyD5ZYUS8UmTkdktpxRRDwWC8yxHncpsv5OvoRZQOEiIVSnvpbzYwMXbhPB3p
OCtkMHlQfvk8LKl5+aJoNO8AcyfqucqCKMEv2IYCF9zN/Qe48TqidIIPC5JWXjXNyrIx+f3zg7bX
jWF7drGvSFnQpjxLuYPLlT23W1BpMBCYnmczDPOBCpV2l/Uwdr0Vyx+/Y/pjF0u5RuWFdEad079i
absUGMFws1ssvKh2BHYkGlKbo5cFI24by2B0RO+wrh2px1yy5ibk9KDYk18GmMwBvB0uRaFe47nm
KN5H3/bTiaEsVY1o9LMkKxwgcDAakPYvWZAmpJ7PJTRTtzrDPynmxczp6z4Un+m67qA9MShlQt1m
+wR7fLWxtQmd0g6B0VJKLSAdsBuzkZZywW6oC4RLCMbgVh7CCfY5ad0N3hscvJSfa+hX4aXTsSK9
4VFULJdGuK2ufOLSJjLvsQtMyeYj1FK0mjdtmg+v5LcVgKFYaO23D9oZNlFNbEE9XaYE5hhOzSeu
Md6f7gksm0/hqL01eqXiFloZDabllyQSmFLcsmCbqqw38gwrrSNWE99+UBhfGt35dbMKbScvOihJ
CC/pWpSkckwVQkhfm3LdWQNnxSLlrRjr8ClZa/AvBLhp8+DMIUXxKd1l9Am4Hnljkefl0S0xZXwl
oyt0cczF1fLE42oaFRw0kOMeOnvbxtiSgMgYqoJW614DdxtmKftFXcC7cbfZLAo0wr3wkMAPxCmn
srJR5KkgtdUx05swh1DZPT4q4t8KVytz8b4RNNV62FzFbtsYvpp7FP9ezueSgnUDODq42PZG7zYK
j1ixIdzEzNX+EWaq62cpd6yy+kGW2l+bUA9EwnFag3n2ciroRxekuwKM99B/uQXxXqmPOphaw6y8
pan7GTQVN8qDXvIRC2/oMvAruBlL6ervkGSn6+tr2swcTn+QPBkr5JupjjXldCNrGoz3Io5F4ek+
+pVcnaGrSOI0EAOBw8A9t9YYtLXibWvhbzWEhUgU1sX8/hRblKUHWEJ2pQtmWJfTjfh9Jk+bWjfZ
EMdLw9BsS4gtaIHvsAVNAbDpkHR7KEAzq9kpku7CwTwJOgPpCSnC8fbi626QTItR8gZCgy8xVXPu
QcQ0B6cKYj3DmyEDBTeVFI+lBLAciTNWBOAwcdIAuUxAlpzgqmzsKrlJyYRQq910Blls23jmTRh4
lbvcO1ZnfM/EoYAHhH6+TQSQJdYEAQhyfPGg8BarJTpghBVMdn3C+GM+a2nHqDPiXP/C07lWWGTi
WedLQocebzZJn0oW/6NH+AFBx4zVzXKx8bTeBbJJFD5TdPxinJiNuL6opV7Kdc9Ed5eJMesXjXvw
wOCuRjMk7n8JxxMhAzHisgH30FyaUtNyEoPRHTDjyHbUO88A1Alurs9sva64vmIO9mbD0y8bKzcc
OK1pQ6aRyhK+92wHN4Lxxy7S5UX4QOdj+QA2rsyIGnvuKtCbP1pDY7nIkybqQxdNw8cR+3WYtmFZ
tmXPo2MipG5hi7XffDaOWJbLiLP1KxQe+N0DmB+E31KQuHuq9UQ+VNO3949fmpcmyd4hW5twZrOc
pyyq+Vj2dNnrvqUhQh3MMRXUj5j447Nw2A6wojj+6pfq42h/W0liJA1ngPvBK83FRPOK6oAc7+sd
T8fdITrU5GpI4vxLQfhCP3ro1RrUGzoYPyxFsRqS4mLnjEg0FlzfEHIrBTERrsqn6NZwBszkoLy7
5S7s9vLvoLLs6aFv0wK8khJXO6MOMGfZYZOa9kM4+TFbe/HbWXKJ8Tk37QmwCE/PURpGYXb8MrnR
WU/J7+nYU8BOb/g1RJo2vFXcxLgXCGfrFBz2L/yYvewx0D/CGxAB9vyt49QUVneaHXHlnh0fhJxG
l/PdZhvqEnj9z5HAfLdrwfIOJLHVfOmOKnISZcWFXbs6O6Zbkjwa8uzRQQEGVWfCUnyBa8vf2TMu
OFCrwVYEwpw2Zpax3TnkI/bWT8Zj+FQ9LbyvrsNNvAKKETi4T9+H5HGfpv8zCmKjmxdf2eV9DrOD
X/v6F1AU4GtxhofQMntb3Nb2x0n9peKCpCjr39m/oQ69x+dhG+PNOojy703/9A3sl5dS7i/kshgK
qb8+9lTzf6Ja5FKYLLLT6jrgOxuX5z2plbatgwkbkegbjKtS2KdUgyEjJxxY1lR/7pKXch7XUZ68
NatMQWEIEU+8qZijsUy8SmSYe6u1fb02ZNEGbVjhHNVjkTU1NR4XX6tzjH/UaypJB7GBID84NKTN
l+qK9PCrcLW+3QdxgGB/p0wdu2jXllH91A6JodGkLhgNqMj8q59sJBzWeHiPppFBTYtRErmEePeP
y44Xn9mQeFCV2xDN+pUCWETPHmlJzhrIlyegEqcUId8BLswvd36oPXK2+Ve9El9/m8gEpsYObr/Z
ubB0BEiE+yNyWtsxsp++dgjr57j5ZUrfOkONuL21n7xpft4LOISB5t5iu4ErSb3l3qVHwHFBQw8g
Ol8XvvAkmNUHCvCpjCbCH8FVyTxmnswe4p+HIXLjQJJzB3UmPq3GxuO9dkcXxExkPrsqDE3SH9At
cWaguTAB7h60m9n9uP69RYXTZ1tzhqWzoqMEU7p45vPQ1v4QU6luPMV1ETp/+kEgMU9wEM/BXt7Z
BJRgXoL6ftmlwb7707NIDjmLtEwYri7Xa2adrKV1wUMzcF47+8TI+YDn6JPQaedhyGNg/C6JjFNH
XjAnRUiEMFTAaIoZmZntIt0JY/ob5VTRWcPHUPe7fF0+w0w4eZmRhjiThvDGMjFWJm4oltAw5cq2
OSmmRAENQr3+XZdbVOAAFLRPKSe2F8vaDsWhz2AXmqSY1jlzBJChFKxA+vOOaeZVv0lszHAVUIAg
AzvtIfM5lti+sWuzBer5RZjVsux5U5wJbG8OcrRCGcfItSiEQjBpTYppgc/yy8J5bqDKSTbjYZMp
7LUpOrQQn7Lzi49BEzsNdMUH5MezZC8YLxDlfUhwUS/IG+uQEinF7b8TFsMqtf1DLriNvlTQOAF3
2UTdWN81gVP3Qm4qxN47afKizvHrAkwxHX/EN7a/PgPgVzdnyuQG0NzGQerN+bAI41dKe18DEDi0
swvtBD+g4FojWmxsK2ajg7CoP8zA3cgWallLtk/aO/DAwp3FP6OK5y2pxSMADMm6GNGWeXg5OD4r
c97zMBlbU0kPBBDMLu75Vln4hSLMUinbOBT08iuy2FCanSax/Heou5gYocwBtC3dUEWWTInzHco+
Tj3EkGlE83HRwov5tzshZq2qQZL07SeqM4CPzMtXKFyELIUATu5K3Zha5RHgs9BFIL/Za3ubbiZq
yW28II7zySLbNIWXeAaheAv0Kx70/K71qiqirpgF1SKQem6uMFiIKyPROhtK+vZGN+ux3rUwSFJx
DOesCLXWu8FYdLLBYb5C9b0Nz3hhqQGDBs5qDGyp68w3aGrHAV1LGpxlE9Kzs9Rjsnyz07ZmRE+/
Nc1yYIZB08g6u7T2lcRyU3CzGSRe8LCZalCRS+y3kfXXN5n/zWEfDaLiGe5VSkTNtF1/zQpD4Z1Z
MKz00JGClGhpK1TyS1IhsPlCWG/T2pPcRY4Qev9/20LpmO+CMI/YNpqTzLD9ZlK5Yp+WyPe6pxIX
u6sRCiV9Uu5mWLYUefNoWAmpnLqeZgHKH+60HnBa+XEg8rViFWK2QXaI9F6lXl+w3tIrpLTnpBzg
uFDojO9l6KPIRYKE+9nMJJvmQVVQ4eoy55cUpeonySGeCuBaCrcwLf7HnstqYZRYITJSgcFczTx1
KwbP45ufaQS7m7ObPku2sZpAKPZsQDGQ8ooxNkviVb41eUAWaXh+SOKIE8u+hJ47oLkLReMktDI9
i20HGkb5eQ8BAuM2BxXzDiPgqUwcMZRCjqFunqRmVScLDRX5sAjyNPtNFu42eZJEtlwn4SFxKDpL
SB1bu/Zz+kttD60S9mDbtT3JZxEeGCAlMNbA71cmEy9A2IePo9nQLLfWeQQtXX/attMqsRlwAOul
4lxsTMxQA4EgFyDv6u1hk7Mlr21GWBZIqykY3PIyKOl0nh+ZddWsha5PTmU2BZ/g5C++QCuNxXRH
i4pXM/Mtsrd9RLrveKctLoxPaRM0HNU6wcqosad6IljrFupbeNTAJdfMa0PbBRA9QcFQHC4isxMz
lRNp1L/lRw9xWFjhB2qewsGR7PIjo9oayEdfe8Cu8xgH0LEzA8E8LkL5umcuw5uTru4Yc9OzU37B
4xjTrqiel+d6T+gig0bYnkC/31BbkLfO0QRGrBNNM4ISwOTzA6/swT8rzWXWgTYnOK1ugYyHzMJS
D0s2lalpjj48FiDyMqP0shk11sVh62szqZBP3PCPinlqM7ZgszBUXwvc8TpiLtnppjE4k3Km06hP
zXuRdbk1vU5VMQrGZlEk1Nwp0TUNXBsyvmTcphXx1VvGihKH/KplZXsYBIEEPDxBiuZ/zHHcw3EQ
Qb4iUM/0WkBT58mFuKlNf49EuQlhNXylsBaD3f0/G4FoAzp/bR6oSctKvT6KvK32DLJnl7ZfaeG6
vYxYay+qnMdX+MTySNyoXzC3i1v1IbxxZhRFAUBq3CEa+MTp7LF+a3D/MEXMy9pbI6ZIbqJBHmBz
uc8XEEipW9Wsd+pN/f660W/o+UOw1DVPL6eIexLYrJCxHLZTU6u6naNKJpaPgvX6DjwVH3WBN4pt
IQXtAgjiSeF6ulz+qculkqpv/e/x7Fa7kkQCpG0stBGsOd3yEVi8n57J4ZyGtKYUeH+FI6uEq/6v
uwKgJd9y+wygo9Iw0KeLZRe5tX5fQfWP6F8KMPv3qnGmOTUieKdy3aOtK9hThs+Ej0IU9Wn88pv1
LCfccYVMq3BqbkSKtTn+tOW52381BIIvgOR3rDIoBTNujtV1W/5qNpIwx+aqZwB6MDKBSsTJSA2w
bV39nyvRAT9HxIHGxE0l+YdO+ajsVrSy5uuiBKTyDPe5T//TirZ7nhfFsTlxjoFWiUzWlkbqdK+T
SfcVAeTGuEdZCuSRpHwytZ3BXmLzg23UFi4Db/5r5O9b8z66Ig14cDXsXNAbdDSbcA8u0O8Mcbjp
F3XvBkLvmF0rW7us03ICZJiIdzW2Mhm6IPxT8nRiqr748sf7MOw/32gzm6Eowc4YRR/TDBSX2lAg
KYLj9QncTQm0SJPnGTUgFdb88BzGvzkpM70B8ECDWldwPhLc1I/O3t8eio+PEg2Wi1is6MqGk7gN
o7wxNKqfh0YLA3nnF+u1FH5Umdi10pyKSDy8KUkKOXXhIc0V048D8DdMMAmDPkOXWjzWLf/ezmGu
e6d9snQ5inZOIv1BKrGB/lv7IRxBd2Epi/djYLIzQE9abdR8nAWKfnB6wD+nDWO4QUVaNISKTech
2sI2v1L/PWevHo3ZPtuCOWcgOFF5CiY2OzRIBpeEDw7lCM3MOcTLpGZXl4zkcsLLBgXlzpg9dsas
nWmU6zScleSymOa81M57dVivXZ4UwKxi8sxTndrdphROrEYMGZHeJpRGbZUsbUTofbz8ybO05Xh5
J/ZALCmWyOZ5fESYyw7k99OI/4Kc92FdIqUoDf0/SBnyfcXgLmeOxcZC8L3xaOkht1wB7EUxrcKR
ob3SErzGDvxUchNyn+523g5HcxtxZylCZYBrNm2JeRxSzO8Q9iAhHfPRaRp5SUFuyDz/U368pBxi
0Rf9rshX/UlJ3JfmX+AitEutZ8lhUl8wQM5kbEWxpOEy5QXnna3879GZlqZMslAX57MYlMjN6/D/
MKtau9dBD2rzfiyjhAN6NkACP/grYreuNRbJTwP83FBclnFKAwaLFkE6KdkoI8G+tcNHsTsxpiK0
5AxIaXlWnbFWVaZFrEzloHbdPPA2QQQvSydTFde2aq97CIDtmsI3i8PoM0RVSJoFdiHm6DIvZhbJ
qD0DYVqTdzQK5V3ptslls7iwZUb0jckBJL+P4M4WKWRh2k5Uh3E8/JYRGXkHrQCg1CIftKQJycbw
y/NY7bwRnzicFNsxUOLNSBSIStSPjgzZVeeOxAfQnlxy/Xu3hepGsKTrNZzYC9oxkwPz1/2rCOW3
jxTTMCjAxxvsp84a7mzs5f2RLDVUc04IZVfRXg1h1AR1pAzNSrDNR9bYb/FzpoRUSLUmYdb0DkB2
hkYTjwOtqVDfFgg9yJOquhrThL1d/z1qciyjKmm8EIvmC1AXreQFFrVwgilgoksNbRB2z6V8v30r
+RongsU8yYiYlrncGlB1hlmofbGXHtry2XU9wa7moWuyq9qEeIRjLk2JTTj0QZHmPUOtQbU0wn1K
2n0AGQQhI62mZoiCidlGPkX6EVIjbYHVkoNnWfe8ovj+fI7kFRZMWMoH/kv4piQCz387btKZjO1s
zuCNf8J51htEDoDnkU9fyqhlinoRGEXnErwCzSEi6iwdWtOBNvZb4E5+lx2u0U5EjN0w+bAQOLYV
DIS3oXPZ8/4FnwjICyteizzCo/0wwLfacKnduMO6cnDZRUgWmn0SuSNK52RXNsQOH1LkMxSMHsey
HEu5ehNVnNHVdzRMlEk5cA+Q7u+oDQj1wQde77+/+/5ugMmO8HnXI5efHJKZ+fUmuWwbn1v0Zb8i
8xey14yaeNVQ4wmCsEEs47VynKuMXeVONP7KJaTL8npx1Ts+YcBwaY6+gxKOFgdM1UBcA6Oi1kO5
GBCDDaM/g2z8rrw+7tK2IrH52S71cpa8Gu5/ysLsSPgF5P7WvDt0/V7CnrfI9KsA47wIxB6EFevA
Uoe0Fx/J3wfUEemPV2vB/4+5FUNfNHRFTdXEVipK5YUHbMhDIl7M+TEhBD7Kbx8dJrjNg0yKKxfj
8AtM6sa4qac4GKRsiIiG4q5NPgLBnsjOjsZ2Gm3iY7vAW5YOmxM5C5jr5Tl1LsXivLdgBcRsZ8Vd
kQwsXZqnN6zwHlN277zKB3nV0kANEwDElJUlntbOXrcvJxC5v0j3vsvUxdOxM36k/4a6Q8k395Zu
9501Pccy+bBfTMTByvuVqmxfHbuccZlHWfRzEVToF3Nw83uHNf6Nbxs28UbVd93cghcM9ZD/MBk5
BQQVI0hXXVA6f/wXwzk1BU6hY4K6EuGPeydrsctKVLGB79wBknHdmYdTRKVxIM6vI3PyTgzAo7Zq
lwMA7xuwYrd7/KI8+Hzn1lTlLT44KhGbaLLoYM5YrNLPrQDb2HXIfDOJSQkxNLTnS/9zqinHwbDw
Yg6j8Y7Tw/353pPzLZxVmkUcQFo3Xo0cYihMXOzA01AMhc+Qw7hH6rKBQ8AF00y59dV9zxTaBRF8
AkP1DqwwOmLTghFQw8DCKh8TvlWAe+oZ35VQ/tlCRtOM+G9d4QMP4VAIKCn5D/NbtP89e6z0IN+6
iofjk1NtyuHaLIIKv/BT4guaIbGPgDPDTDqU4BTj9n9yd98DEb2UKqXzWM9Is0ZUyoyOCHnEaU6V
Ss1a0zPgsmW0PqPgsQuCEsNWtHZ+Zkti/dxtBcCRTXPVTCXHXma0A6fHuUjq7JLL+AItEgpa/R92
RPtuFDglma/v2CHnYbbveAe47HG4DVpX8xHNCp53pNQjvh0THKcP+yM9siTS2JOfxpnIDizGI6Wr
5lnoKgaMyyCGLfhFQPyf+gJX/7cpV3+josrnDFKVr0Y5rGkgUy2uRweXU2/UdzZ2CPAJ12IbgEFo
yDAocIhxm4q8nBOc2boxAK7Y3aCfgPwGSJlvnQHN5VP6XTXvme1PtLNLcQH6OOVGWqfmwc+FbCRj
kvwg0upbTMVc87NzPpXbhOqThQBRJbv0g/TPwEw3wlXlIxq13aAwsuoTSdySZJ7xj4lVCcBlYAw6
+xAEme1Ye0kvqdkA5E2iO4GQOu3MG3xTlkoxA5F0kFu6bsqc98k8yLV5UZuxE8cFxvSUMr97aS//
VCgzAa7CAodiu1bYL1q4NLP+jGLrby5VAyff4AaDX3RuYzn+xC4VYxTJF78htxT3QxjZmuOZTWHH
VNd9hWhm5iOaTpcJGrnVGSmr/GRb+vobjHLUJEyIZmoY11O9ROiQbiePyAVaeZDMEmENZw3mp0Zh
pOKelcS2HfQq0LsZVuej6EFO+nH39ETIKR0z6fkVUmHLsYYe1saTLCMcEgojV7v9OxrKciCwCl9V
J6Tl8DywIAeS+0vqcvdQMqPheSgAGaGJR6rWQ2x6n7qjq4vcc2UCh2Jn2vqG3zMQEr4osXmfykBq
DodU3g7bOnSB8O70LFVjWAT2vvI3dJ2ONfQSdCAs+4h/e13ocYkqo7+qmxLaLpIOp4J2NmZxCfeW
le45EyIQ3sqVgMvF5alINqHy4x1EJMlqA482BwFuZ5oZqzjo49XcfDB1aHu7Nq71ktEZFXHgoWxf
5UXqasJND37BQNcxRKe65j5cJk1PpZWyEkKLSqNUzPxCIFDI7/gkuy1fxCT3xD0RubGrtVTsqoSQ
OJqpg+RGEX66XWV3F/F00pS2tY6Ab2VZKeBs87h3XFOc9H1lXU1fsOvnQlrrMyv6kHkvDAlv04Jz
fdvEqp48gpF+nPLtqEj57ea98BatOfhk2bL4+NBeNOYBEG8SBvteLva0J/cFncWYhZFy6Px11lzF
jWmFNyPfGNn6+CdFEpolpboNNgnjx4IbGg5PDdD0R3CH49JeMaY4xdHCFYPs93TLb6mS8DrpvK56
5crc1pQR6rTML681JH0gAZ+0ueRuURkPWPT9m4SnHrd4G+K27Vgiy1sN0HKheOG/XzkAC0jl/r+s
dbL/yAoja5E+H2lgIum7WA5DIkqMaZs/2h77S2teLkFstzgtgNugKNSAvY9GxLFiO5l4rCJyojkI
TulCT3dplDO317I3TTLENtwA2WdkR45VzuLtxw/MtSoFUcn4JawYwvqY6g0G4L7NV2sBxumkFqtK
SFd2N56RkHAUjtfLFMQrFRWUUz3f2g/+6N6SYZHDC7OFiIk3D7U7FCE2KVXqHr/0grr2nhB58hOm
xUC9lApIKT6CWMIrmrJvOYRIW3x1nsFEhHJP8OGfr0/X5CTLNLAlWaymcvhXwz/f2d8R9CnInfuB
aorVEsy76xGKTNNXGKZdUwyP06MymTB7SgF+6L5+OypCxreNxPAmxDNnG7T1wT6kS8GxGX4R1lkm
Yr97qZzJVkTPE6XAFUhueK/qnSqnG5PTOe5U1bU59UhYBjTWDgArE+R5G1iCj25OSt5rVPhfCGyd
WM/CFljSMmNlMSIN/40cBLimXCygITbUTNCnH9yR2M9zs3C5pZia5Jnb3sOhKStnfj2dsMM0yMJ/
CoMk5IngEv4Kd1tYIs91jHmWH7JKfb/F0NGD89FqFByXja6LyLnBuafTNbP0+wL1kYyejFx6UA8n
nEwWkg2RY2ZEQlqlF2XZS7/PXBjoQAztYtHtwg1bxq+pZbehSC3k6bOnp/3LykvtHqm4H28NV0hM
B1aiAwFB2hx8a7Hs3A9TSaLA9zJvm+9K0oW/0pXjjFMrj4GGSRE3auDzl5tWwhEAUU8yuBmHmhD6
1GTOtVQHoQctHn6Pgy7vmDBVboNLCwfLAjVe7mDB3h7ruU6tVfS2YjSXPOBSLs3Ndh6TtvKkEojD
tjoYd0OVocFps75QTNYtMB1i91hTPnvD98Z60Mc9UjZ3va9T2DoOXvb2ppMLcOwOC0KFmxLuNSnk
zFm/UrxLur/x5r9XMlf2/SXfXn4wpSpZVOvQUpd0EeheO0bBA7XqYMLN0TzPMFuldituA5+voqlm
iFHdCFUMXm9tVy0evYc0XELWxPikYHMLqcQV8Q4KhFOY0m3UA06jkEQaEZ+W9t7YHLP1FPxdezW+
ojsQtVw06MmrdYYMhHJJm5ud97Mu9qUHkUS+2CHnvEwjoj0jnacPiNEvgIw1i+FAJl7yIE7Z+KQ+
AjllHGnhoiquP/P8YdQjLHsl0ihlDJlSRcJ4+ji1YqEUA07cWLuTlOor8+MHB6ZKP/Ms4Y2Ke9Dh
BVPF1+s3WvOdwhWpH8DEZpXidg4+clPlD0uQguRcDqNwGK5MAqCVBYi4oZjsl5drGsMmU/fTw7yb
O8v0/ywM46fY/b77419wMrchKmRsF7MF8FB7eRnSG3hvp3wO/wL1s/4G6jVZikBBQmzI8mmiRyqi
NxtSmJI8mlUj42gofuhjYgDs9SvbapX56bCAAhmYbF2HwElj5EGg6jkJJfyfNpsvKH6n0vGXguQw
UDhrrjBwSiuhbvvOyFmRODFWQl6wAoOwicPaoVBY6ceRxBLz3BFal1T6srCgsNVQLnlv+MgI0BLR
xpQfZI6meJbVUBY+R2IqAum/OxnVnVPsJ/qv77ELc0D2cY8EEeJTy2jh+Z7cJ8+K3Z0WvF03l40v
VG6W6DUWPKI44jg+GBEsfg1ZVI9cdyCpw5d1vvJc2Xt2MLkIMgNMOqra0K0u959Har+M9AabXRh/
ZxIysSHDs4vvy+s/JhqRtrP3ZX7a6zLevQSQv627+resaOVNNAma8bkRfuR/zLqQosy44kwsSTlq
GVjKjy0aWmfqlxEwJMmyVYNBryS92u2KacWuv/H6lei3q0h2qg4zc+9zeU8zQCjEcr0uKh3ENxOI
KBPC61qj7Rzd0jWhqIKj25gEAEI0bNlOAdpOr5sChf5rEdeMbJxp93zvjqZ57dVuvI/YElEistNI
o8ZBSEv+D/AMt+IiwYW2ZA2lMM3fX8OdOOJsYjk880atnmWLQRR8XMarfqRoXHIWYe36yhaM3en6
PrvF8dkATyY8SVNpPiDDiuSuy90GhLxDlCPBeh3C7XamfELxegmYQju50PASA+yLiLUzMv82xD3s
BG4IlnkbpO28XjtSADTCsuOS0p62dMs6jxp66E/BBV1efYs5GQYdbkFAl8eSV20k3aluNb/hcbme
ZqB7NyVUCsUr0UzInlt43GbwIzwS40VWlYNU7MhOVYFsLRWW4RCk9appSjzPRyrLLLzew6BfIGPi
k29afgwn7Tfrqu3v9nWgMjitOn0M1moOHEGuTgT3toLMEy/XcJO6Nq4pE7J6qX7cswXp5ScybD3M
LsWO/A6EF/qaFzyU5vMasf3SN36X34DEb4HhtV/IzvWMI1mF9r+SSu0Dm3tREVQvFG4o3dtdKByI
8agULim2pXa6rmdUO6PTMkHvPmJDjJFJ0xRbf12vMxxm7NLBsEcnK/FKTnfYihJqOOpGkbe23Dnn
1nQlTeD/z5zFgW5bC357n3lJzxhfOeW0nfIVvlsSxFXEFdXURPzxg4XLjMKUzfhCXcjJfGJhfQW5
MpLLIXKq2Yqqgu9/19FgIDesK6CECzYoMu8dS2f6wQdiHkkKZ6XvLaFh7bKGLbrc7Y8w3xrLG58G
5F+/PmjqGFFQ3sQaSwf4ElV9a7jLKnavf3T/E9rk/K09idM4pk8PdTJqQpfYEF8jvqioCvJgSD1O
9CPo542TrS/hVub9WiEMu96LKYtad/sf4DlUqSVHMSsHbrfDKX13eMB6b3c8pvyuDN6x4aqsY9mW
QB+luQ8O5MUpQN4gOmTv5VGIwiob8vV0gf9DjMFGd+fCXZat/fncdBbEoTqZbm4s3UanfuAgKwLo
wzf4dOpnZaB3c0Vst7MjPVfIjKNoL8heoLvBg9qZB/UCLRD3K0UxAZS7162yNHljODAyKyJI7H0B
y+rEO4LPtLT3C4ziBLDuAEEXwI3xPvFG3S//oXvzgVaxSAIdjtSHWBMudCb6Xhp0qhrwYHXq36HG
ydrR82WVP7dGKB9T5OuqQGoyWfpGyD3eXd8p1pbSq2g805cwueyUd/VOYUP71l7XBwDYiqlcmXXw
3xbz7I+WVgUUEDiFSKnSJmC7ER12UbzLwfjezih8tCnGfufCFFMQqvf38Si1GmHMaRL8TwthfjSZ
k043eLFSkjIS6It600PhKl5GpIc0OqQhVkmjJWAdoVVRqxrn3PVwnNBm6v6JBIiOsPhJ1MA0iYpo
LuX/kZM6LyY4uO7+2km2GHZCpwTKcUsBg+KgFFpvBMBuFaugwn/tV+NkWcaY5CkC72JZmtHRSCiC
XK6G90vQdumX3aH4AtT/uPhpvhL75pKi+taWrV2GBrdKVby8IZoY6wsdD17rZDIsxNTQCaPVE1OF
DNhp+X/BlLI7+fZumn+yHjT6oOyLdCuhqF826FtZfbfB2OfusAztMj6GlkQaR4rhwkfGPG4fuB4V
uJITN0CIQRV52hI1VKXY84k1GxJ9xQGDWYLdJ22DLcAMABvgtb9J/53EjNHuVGjrc9lh71RRe60y
0smmcPHNcitGM3qQd+ElBif/2YFmvT87GukhHUVLGIAzEOiRO0CAm31/6mFj9F4ZrH+TXV4hTfOE
xxXdIdJfhGsA/K9PFZZlhbB/h0F9SicnUrhbKgIU94xCNeT4qZx2yvHE/naPOBTnmw3K96naFRtZ
CU0FFCwge5htTKeACuSdc096/6Uoxt//XbLL/azd0llzC4oMgYY+N+I4FEgooGrnofF0kbL9BRqI
fIIzd7EX39nqLF3FBKVM4W6eOIP+he+CfKYXXNL1bp48nFUQ7GrvzXtcJvdfZnAmi/jh7OJes+Rv
V8/L2BrPg8U5d7cm6fv4gouXJf1SjVD3abo4ADxzu8DQuv20+59jHzRy5GmhJIqLFvjRxKTSgS8C
qsELr4QEL9/eu6yf9LkiCWf1dozwlfkBKFHPmY1KuAypZtP9SetVyTwgCwREEhlGkQK53dgqLGkW
PkTETupqbRaBhcd3O0jAJLUk349Kh3RC0gLwe5Q146PAdAKbBLrWslhRnV+uT0VEKTeg6WeM20mP
NcVQWRoorfeCeQvf1TqriKcdUpYzISxk6K1vF5S8B8h2BcnRsHrIx5hyoOn6e7v4fALcrx+XLRWm
dqIQhwleY4cRvPXF4T3SJpDPod4wXO4lvVqlei2pUsY/aJz4qb37MO9SH45SShZmgkPcuelGrDK8
Z4weUQJGul05nIBPOzH4R2c6fwqBgheh/on1WjOcFEAD0+tWPX5MzlpRGsxZvpHBOuFId1L43wId
4q//stSqWqfmJLRfohTOU/8qx4QIQff2hHEFWc2CKTMj3CCagT0CFwAUBQ9sK9H/zwBwJGT8wD+D
oFZqplU3LAQ2i0oy2lmpFfHhz53wonxQlsnkQIid3sMLgiB0h+tg7dh/+oXhznpjZnjq1v94eysF
KWuZsSYdUjhtfvc0TGVw3plQnO4FHCiKFPG5msb3uncdNbe0dY9t0bnRBfnUpt/YgSpqNXR4q+UQ
BoqCFCyRK4eJSp8WowlKHEW8IYei6D/P695PxMCd5iNHdCLKB7rhJ2bw7YbtWHYeOFgwxb1k/HLC
3rL1CInvRbdBt87Gn25pIlQ27Q01o1lV1fFgSYchXRIoURGoKFFDCHAiEdrbSGd7gepZLYzWklye
CnpCL1IZ0aGPZ1ZRu1PdHhGVteCuckFHdPnRqdr6+U+Brj9GWE1TbtGHYkI5g1k9LTaiQ6G9/x5l
1Q0aNgZ3CiPrQBcRIm3RIEuroAydEgSDS+0Oib1HgBVnDwuXqHby6fgWuLxCaiaDb6d/ZcSCTde8
x5/kYItZSSQQrCAqixwY2UhvDkQPtSb0mSrdKgz5NQBU36jepnsmvsYO8KE98iDmTcao9g2tADrM
WDYpAekqI4JiCdp48uh1s8dGRvrV+tUS58ajeVqHJZwZIwWBjGACaaaT6PWFvVPCX1UEElhe0HYg
YIxGPbap3VSQHwKAZTR+JuX9KMWpA33yulT2C6T6AhE/jOVNptMlRuq4OwN47RfIVTe8e0mP6xsH
zbaZXy/RgWqTJaUh6hnXf9uevUl8mu53+j0ALCVEUdgxtRK+vPSPjAxlZp1iS0au+KNWDlksBMxr
wZW9eXYAr9v9De+UXlOm9XxzP5AEWVT5R8thB5Wps5TedDQxgCeq0spv+Zop83R/FGUkTX+4zWoQ
3a8+LMgw1FB3EnWpAxu0afe0OuPkOs1qjPPkBYqY0hPCndZkScQCpI2aKD8lwiKNgRozV2/3sKHL
b7xNonWf4irXcabW62+DfYkoLid7Llf2kiOT+OEHRNg8b77wkBLtrJBfC+o5Edpo1Z0AE9GT6Ke3
fiQ9cq4IBT+nhQoTU2oJTmagy6sk5utwgO6l8AibfGaqiRnnSEiwNHRPDqX12wWDsE3b2E50o1HL
aVtbkLrmsY9Xiz6CN6zT0LUN92WjXBrfz8fmnD/YRYFm4WOQL1ayfI3LEFvHQZkA/mrW1Lfjm8bK
HmxcinsoJ+sPXTAQ6uW4T8KX2dG4jcoOzidcRqp57C1mGUuXMHbbs7g73FRaYClrQ0N3u6tIxVZb
5gGcdhStyPylwyzZ3J9NjLaXvbaX5BcUh41x+e8W/TvrEoRU/WWHA53U4Yz1ZV5503vMH9yXYrFU
mMjisf6ThtCE5Ji4cwgR6YJMCNWQW5OWkSMEIlzDtbyy5ojJJxXbQ884FMtbaP9X5ibvLLwCLMVg
QU51nCY9YNLLZxX1P0fle0nfO+VsZwNdE10V85WUzpgPR2SI8zCDAUSjFaMTGcsIYvZxXXfV/3k0
3H+Jj+q9uugq9lMDnk6vWp1UZ2PIhAR8h3KCKoDJoyheKIaBx8ci3+YPW/fxUOBGWUA6FtzgHow1
y9QXZ4LFi83nktivTYLYwuStf0mb9YNxLX6AwqkTYhe4OexmWfkP1YghETdteVD+PnujSOVr+0BX
Z0MaUrjwYG6TpKq0bHX0m5owHRCyXd5KJ+RyHoFm1HxZQbuBzuv7IIE84JnyDg/ZpyjSn1qExTW2
RGeDrolu3NVSaJCI6loiDlsCHcQxF7rK+gKqbgmBTHDnc6sXeJ1AVnX50X2dGOP9zxHpPV17n/el
RDDD4YzQiGoJbdVzXBqUT0Y4cEUYiAXJN7RuXsZOKreK+eZsHbpNeILXqNWBeha89oMQjyIG6LNP
psGfZKPn8N1PvSRVrWYn0JWQAo5LBngEQlJuCUfotPIZQ7tB4iQf1+rkuT2irNLQAfwlc22BbdJC
8vc2QJbWlSq1wwpDhv6aux2eJu+ASOpsCQMFc50Oo9sI0iNW42Qq4Xx/2Xi+3vhqzakcWnkHZpkz
v4rimBUSz17nd+S0lgrj6joOdvZ+WUqTDmKNUxnY774kdYJfGg57FXAqna+nPLy3+KA8b9cBEW5o
zYMdPKDgxPg2P54bGRS2XplwbagHvKkH5tAecPPrAMC2Y0FuY894r+84fvOEqFcrbnmPzbt7ukVc
I6ip/aQwHUH+QCdStizq4zEjjMsTEQv2e3jD06iV3GD3fMUvdrSDa2BbcvJSOMb/np3J0+/TYnrZ
jb/YKWT3WptgfCPf9xEW/mTG/s/dev6o5RIjHGTvWnY5Yk1bxzQ0NdCnKUdNXXzGrX1RmwFgST+J
zg6O/SAexggk7yK51BZH/wkuwJh14EoKE9LuYnOHiYAMe3hZOv4JIbfJ+zICSfGOsvm+x+RTZ3UO
OI3w84DGGwYhkkTiK9aNeiUc8OU+t9jWTA/YPTVIoKvAzniZQtUE9SBfqRwglNERuxzIbKYP5c2g
H7VAkx8TKh0axVx89ZDacFj4GtZFks/c6LhDc4b2uFHqaTfCk8m+hxIKTm77FBTX7WAJ1AS9C8kr
LsIem02n1uEG3egZvtimJphtXCQss8H5PdmqgbZlhRmQ2KD2RRMUJNlYMIE6Ee7BuvODEgamjgNE
EKDzLnsQCHsUGN6sesPv9MD40CKHMCdiCyJEFl10RpKLXT2GNaJ3LVoqRlnRCB3cyFasqrsrD2c2
ZtmEPuFMT+f83F6cKDnjZ5O3pnXGNNCIKUEjwbMBXP5vPpZbNq8wqi3HFbBjOEP3MBV/Wwg4TaPt
qz083YoG8ju4d2/LCd4qy5iLgrrnOgce7rtfCsOpCBhe4zaqOIJ/wXmciTWB7PrOCByc9GIQnYSq
yM2SXfcSAbbkjXn6nDSJIyuQIes1TsiY1jOQ+rCYHtjonfAvEx47AO+MxL/tDbc346XjfnhVZFBn
dUXSqNRwFtOIr9wCEkafyyMqdDJ9jEd7UmjG1lr/IAsiitavgoR1RnLESiwVZslqCSfYbof9JIU5
65SQ4qXpkKxnZWG1pOljgVXl3ryA4L/O7NL1jL/yVYC3IB65t5Z+iQxv89NAJ1JeZTN46KNrhUk0
AidS8bbcw3JwYrRx4J5486HsJE2XATtpGW2dZqePRnYX3wTE8FMij2oa5wMag7MV3SoZhHy6A9GU
gMOc8ClzwItpveYdUJLK07ewcJVnm0oTb4SuuJiM2dafrSo4q0UCUJ/94hEkeRIA+huipXUhy9V8
6KcWzZKPRoZg9EqYXO0urlOdpNBPRSFcIeipnIZsMQ58BtaSVoCT041FDmJfBTV2bSMS3J4u9uTR
EEgl9IFftXUCF0NZGmXLfy2E9ItPX22G4h9Zy9m5gTuw43tvAKCVRdzQkqrTzyqDil4ZLrYoSxZf
622pNo1LeKpAnz46E4Tlq5RayibdwMNaRKEpjte8jQQx6K6WzYGxtioUfxU9mXiOlKCIJS2nlIUr
BFwfxotOcOOS0C+eYYlf0FkIzloUWJC8geudwI1/cfzM7jNhElS6+5C8bcJkKF6oVQJTdf8n7Tms
EHrgD7PeYDbBq7hzx1R1tPBeD9gsHdunZI3UBrayTrNTRX5zaHJa9U3XPKFOjErJWAbkYurcthyV
n7pcZWueENj5l86APJpmEhfhA5dYv///ucX1mkag2mBfxDGR8R24QUx3UbwRzR9KZHsxLo7hz7bx
8//a3zMFjeHhF/Fudrr9WO1i178DyMbg75xVnEdIiNB+HjTufraw139yshAALGlZB+7tUAQYoLKy
R7stxv2g4A5AiB4wPj4g6jJktVmbn6mn0ocU91VQE7Seb/fUqR+SCY1CufJ1Zq3atB0Ks99zV9Rb
TC74VUJ8j4aD4AIMBZegMvGRJK5ezeMuxK17759v5NAGy5r2jPrZRwkPSW7YE1ggtowxfVLEpYyW
HnMgsZOKzWV5fxW2QqjJbBGvN9s6VOixndcnEQtrqtSQEPKpSWPWE2tJI4xeN7rQ+Z0T7dCjV4+C
isZ0gCwYjFuNxlctu7v8bS5L+Z8jt8RTWJTamC9cVx4jU5427Sh2jUa79SxDd/VzZJ3rz4ND+vXM
l1nn7pjKbRPdONcxnxYyhuIOQDieraqFpCq5NRlG0MzCcQtdMWvVGrQSS83Iqzub4fJCffB50Nc2
st0ILkZActrBMvrPvcxzAjR71T7y8gfgHd3nUPrkWvJK4BZQCZXOLy4IEEagUKRkVvVWClgpU0hH
MgeZI6hQthHDsPkTDwYqK/Cmob9toWD0Kx5P02AwpynEWpaGJ96QUaY9DkBH31peI/39jtwZid2x
VmSlIidPgNNkKNaPLp6QGvp7mzY5mDrcc1PW519ljhGivKScTo1eJJS5GNJWavEvUSl5zRaREcDF
TAjcBoc39zeYuFL8X/Xm/V2LVFM+da7WsPBlB/rgvyerhbQKDDd/Zdcqm7K/7b+yS6ipe6VWQEFQ
33x+yqSNUdzKd7PNqm6b7wCf7DvUnkVykPOJuCzThqtCAssAlTCrT98O5gEnomNc6t0wrud83HGo
0Rb+y56lsmuQF+9CGcY6jkPAYouVysT6CC4zNY4KoMkbXWyerUVG3i8dEzvZNf57WNPfn/xVY8e1
QmnuYrWbNPnYKMeJWMkB2g4UZ5/+lUM/AjLbV1alB7C4rXqUXLMQoO4Llj39ojH0sNA923EBJBIw
44vZhEHsRCwdIoMA0glFuveWE/aNY68bqOVStazLaHWFoYZdbw6ZUaXQaneytsj9pwyeB6lN2wxK
XImL7zPnxthg8zgHLNh6wvUkAKbKQS8ELQ19+CgtFV1X14HAlcumy15lbs4WBJzqQAij5A/ZJHhw
23JOMtcBIIn8LZyRqjZXoMR/r/ZEi92t/SPinylDAHZzDAa9JTl/evHfaNFMFQ/FhBoMyY5DFLTX
45z2KromLRHZyKrhmDf7bUfJ/VQqLb1bkmYeUdgl3koS3YbnOfEvEZ6EmKDWq9tevMwhBbZ8BXW6
OXZRyOsIuf6fGlPvOz+73CkfByvEL5+XXEuyj9y/pqXwjerYoDhOTkBoiofbj8I3gzUBjlTetzxy
j55FPTHR0X/Qp0/svr6DHuAjN8JKOVOy9jAToXFjmVLHzK2KZn5y5aITmVUARFJZ/yOxs2g9Ad9q
dCp6bm+iztrERbDESb+STlz7lKOUv6WshEMSxlQQ263QzfYbwmrt0hU627B+BC+pdJN/9SpwFXKU
NAXgvduucbh1gkiTThuenecRizgT1mCmUMjmaqAong/qcbzeiLOecfAJuNGPddyA0oxLqEbSsRms
jo3Ds7JFPXRFpBZoV0tUeL0KgLNqgaRO6FMY4E7HlctTgj1hBS8E498+ar8qEXDnQ4hDLkwHEqQL
GC2x0k4vUkFksM/FGmPBlMoO82w0HeU01fXoB0zSuErIUyZd1yEZbv73ZuCFHsLw9xnECzTyZ0Zm
cnVo2m2Hq08GDC1ypsSbm4gaHyJZ1wd2UYsKEgnsORa/PRN5sxf3Uv+gyi46Ab0K59xVK/4S8MDy
Sc1PmZdWFfs42Qop5da2LNgpLJZqc7s7yH2mzBmmVzQ6rXq8H8LCnkRwdrTZPlKHdXPZ66LQj8aD
496Bj35xXXL8iVr34vmrehjvoVpGu97Ge8PAKIT+9OTpYJZ9PgHeZ3vmxJzbxSaslMw6HfS9sfE9
NICKbbBx/LkJ4VuCAiynZbd3FXqx2wXNDfUpB6yHAhIx0k1eoZQxaC1E6Yex4MBGNhQFHk0MaFkU
mSaJusx8mvICl9YUWLv80vXUlupt6JuBU4EQWAoYk9xbsRdd2PcgmEWhhmxBXULZk87fNyQUBNij
SWBJuPPSZm5kqW4wK1TN+oYMuD/i0zeyzFLnLGe2/ReY+ropwGavak97tg6Nw+UE1nok2nV0rDVt
CtwRNlml4vz2JPUJbmXvNMtZXZWyUX5YGTesmcqSgfsxJFCEqF/Wr8bBZ+5cRg1qh2ds9ScxWfI7
MM43Z05VSiH03IXgK00GJXf0WsAyzYAn/679BhNByW9wvp7Ep56DTYuya+vW0pnYzg803yMAvvaR
69vcjMAh0Li6jE/PHs3CWeOu4AiAiFsU+HEKabL/BWEL+FnQ6j8lvHeQtmlojY1BDi110j/ek1/0
z0JRFqNLA4aarg1YI9Hy2wjPvx1SCYdKC15gxWB7/jdK2DrE+vUL8gCoZDsfx/apVjMHFVlupofB
ifHMtgyyGGOL+xxjq5uwAFPk+HuO7XXYhKbQfIaaCzog6J4NoFX6tr1bcnMjNJzBpzw7WAPT1WO3
eubg05aQUIKONU2Q7fYB5VCQ+fAJX2V9InzSeAZGus90wtJ8Z2In4hlRSIzh3UjdERK1PIxMv4WD
4XnAccA5t936zvkNbf1Ei3v6O9zfHc+hWMbTTFZeS1ZkqAzYucAbO+NjK2DZslqrmyJBFpQTnrSD
OZwuGQyKO4/YbfrBb7aRrM3Jexr5Its2YG0XKB7YiqSs8KtoMSJrC9+BF2qNJc6wCSoZU9ezaYks
yG48hfW/lpRoDGbFtsr10t3aak5ys6o00bPBvsB6Txi5YAdrKzE2ILwMwRltsmJDAEQgYpp2z6qe
SSzh5271iQ+76TGWuULL1M1/ZFs7e/zeVGtYIdI7bympSkrzjE8SvaGYoUYpVZP8/50SmujOhYX+
FiRAyn1bx19eHASp3xExixED603OqcR1uvNdOWyGiknePfNgT6KnJGhhY75KZ8vFzAHWXeiEBRXN
8rZFsXje1b9M3zOvFU4Ojjfp7Km1PBBJFXYa86bd6tOy5qc9RrBlScJMf94yi8WnMh404H/6qkqS
R1C+HZaUQQg4vC7PGcvjZCqnrqkRha6ekBF/SAWCTgdOl0ma3e/IB/1i+KdmjJPO5P7ulGvEANqP
vE4SQJ9tlUesj8wd6ZdK35j5zkI+o8jus4/NqSqALY7avNnWvbAOgOMupWBCSxrQ8lQYcqt+jlze
CFLklZqFJwMeZR89yjx3YRxotb+Z6LRXjwVo1uC8bqDDfoB3UGwB1uMiQsifDjj/e4k2uuFb2l0Y
vCTMNxZPcYnquRf4fsWwOcFSNLmshGFpG5eTS1TfnQO2Zvo7Nzfbd1LsxruL15Qzi8Hg5QVyhuj3
MacB80zsV/G3rPPPZ/a3zFGahQ/jPf1NEdfPXU4+qqb/Ci+eDiV69oarUnbT7liKjMhRMRhS2k84
uWEH4jPF1hnwc2Cs/OapzZJJNGY4I7lrdJUjXncWHk0qnqcvlNr/1Tve5aW4u/K0dpJ0RYIQ6J8q
mM4XDB800m+IBgNB5KjUSMxOTT0L6Z/bTgrvEjP69cEVHtKfyPgKYYL4PokJ3LDsR9Nds9vFaTSH
Z/eWJpwuO+9Lmg9fAOWqQnHKRe+1wQteLGcJqvxnpIDDyDeWajO8JvOLJPsjOs0NrFcmW47a8cGz
lCZsOPMvH1k/6Wdw+sos1t48N/djD1uwWM3MHUCbSe0DV2Fi9nrorf8WSSdqBw+qbcpfFSMIxwoV
zfW4Kn2cEgQ5CqnPuKwCIOTpwXt0xOwPdz+PSS0n0a8FBUKuocsZ81emcZGOm2UdVH0AOBVGvkAN
fOiWreVLZiq4iox4m3Ved99kCG0nSkUaJsc8Vm8ITCzvF16QZGyAu/dvCMXl+E6jRA1vVT0Z6ySv
bSlB9+l2nhabRjyWteUqq9MKovyybxzggiiCY6TGmZYskx6LBMllToeW7P9HYKp5LdtwYsyQ3yFy
vX+aDpnohIHZuCfrgyRlmKbS1TBAR2DEt4+HwKE/Q20LkbX1vphQx+glDYkJjy37StZKP3G9bB/e
/l6f1jAnthKx4bgoDfuL/wW8EnNTa269gdvAHfQvzVnYqbRapnaD3QO0gqrTEPMVQsOC3k/Rg+qu
3bBtY4wvFSPVpz6dXrfR42XP5mIOgEmxPIhfF++0sI9eXeSlExlCMPvZDvbQYO/ymxa89TMT1KAE
rp1kWvILyf+u6bWOsESCXqA/eeSVq6939XLyqnJJnUZAZTip2i1r6tvun2nE5IWRQ6ZRtARji63Y
94m1U537jjabQkiRzMiVzPCQyQD6TmoiqwBUZd3ldKeTTV/4ljaZmVJZ2SaOtpx22XVOz+WPO88Z
xSzvaIaGMDjGrmPYqk73kGBGlC24Slcz0hnbv6/A3osN2m/E7UkRB2QDlKEs+bMHbGHW0OpOm+24
rwOkwbrYNlLGUIvXqi+GP3GhAZxrGqmcF4rCH1CyPuZJfEJhCGW5zlPDBKYoV0EVsXJ0qFsBer9E
una+PhTdebhLV39jkuJlqYaC/Cy4HWPWPHO9j30HJBbGxqR5cRQehDgNQElfzMqoSia1ZnmXu3oX
8WY3KpiVL7lW7A09nXRdt1JnTDSp1ijWmyH8dks6fA/vYQB5UyKhaZC/D+cbdm4S+K6OTS5vlRsX
OmDLXfiFTcdavIIRMt4O+wJWEyRQGt4zAdqjACKoBNPYLle290oBAJW5G3CfS1mJZPqMvVi+sVdI
hOBwYE45W0o16Mwd4/QBxYhsqNpElBxrJEvWO4V85/Db5BABiEL19bIwOhOXbZKFR5h59561XZoE
s+pbgxiPQh+gLqo3brsTUA6nqRiTFSFOIzSwM1z/eaBTwQgMGQCMLYJq8Azkdl4sOLoGiio/aOrg
8l8/uDDgjGzZbl/XMJxZxIC94hMfxkSDJPi98Oz3ZDrG2E3lweVDrSBNDCsjyJUmRUV76sCxFPYU
0ADHzaeythJKzic+X9KrbgaEWNFD2XgGX69NYm7Xup7xHRXIrNdTsCiisRq4I270kYK9kZX2aWpv
GvAkMui89Wyy0Vd+faBVrAtbXbEy1eHGLX/HM7ika76RX34Haaork61QPvw7e9PpZnfeM6vKAkDG
sXbt1a4Q9f7Y6+DMPNRyx/yXl66cwIv410cGwIG16cuWwaGq06O/T36O7gIj+XcbxKlp4hMrH4o+
hGaMY/33FWzv6wkNV8hYQUmfRpkBfrqCOs4vpl9GtOGGiMIZ2ddKCrsWTTWdUJyf1XuT57DJk0zs
Z0ZCWbwLYoPNVcBhA6Bn3fPzO4WAKRpmsr0G6/aEWD85/tkAdzkLzXwh2r4BvaHpEf+CC/xGYp2v
VkeS5tH8Wip16oBXdIj1HlVGN4A6YcCr5beJJsdgZRJazV5bK9OU+yJ7IaVacfv5Tu1kuurtpZwr
JAEUxcxl0BqdHYA6AOD7R0Q5XWmqzVWcncOFU/sYuAZdXZH1nCMNK2T1npVf7RZgy2NX2tPd/vEH
00eIWV7+oeISsg6mK1CHAUUm2QdyKXDCzOuRJbGuGTlgzzJImUVXTNS5fJxoQoZyuBu1htadRG0n
N7hy5tEsaXwXncyaM/aenHmBE5MExMo2q5OAbXwSuldPkMzTa1mlPbCGbt012suQY7ZhHxqCeeby
kwI7LJ7KqxXfbeOEyyOao/NFmo1eF7Pr25mMjdCCIEtvLwuCG/6+TtAXIkf0bRoSpwJhMU2qQ1rq
j3vubgcbol2WzRm0zxCqQrvZJrOaiPGnTVvxlht62weG4dgaxlTgypSnwPlfVXRadKdUbBUw+rQQ
yOthL3e4EdFX+ZsbABjdD6panGAuMo786/Tdpg+cVAqqQeSKoX+a9wsLqg8vc3PWSwXhtnITmzTv
BDBJjZBnjiHxFzjfHB006ChpJIFr+gS+LT9yE8TDRxmOsxBg1vpRhWCbFX+q56YuVYSv7LWEYFKD
Aqzldr4arPu6PNsThPW4OKqpG9xXe2U/T/IgaMoSfgVIDBVP1w1tz2lkS0akoAv/jft2xL44udDw
DeHIrgdm1Z7lrGYLX3Xn3YXVAX8uS4lpWMMW08r7XDo0Mp2b0tHW8kBCtAKkUT4C2MYeHptgkn1c
mVrhzpwA0Ct7jy6OOJH9VHqRgVSGgws80aNTy9Qz3rBcgalVYt1t7dgz46ijxSESP/Q/GixnRt8g
2kTe36WipAqTtJqP4Xg9gugLKhmy5Q09ntkwBzTRmlybPpwEDmJH0YbgqFUp4n47frh0FfIW3tPX
+jTjpcv1mTZJHXcmfmmcff8AVNVWg4Ga+9gYN8J5IvONzpAazyqO4PZgMzCmxp1dI+m9a+PydrUr
uKixTzADKVEfB4GNfja14s2vT2HWR97gfyV9Qhy/zaEzSosmglgsHINcUJQ5niHcdtQ4GrG317FV
M8G9TFPHFgMGWx/JTVaeuaB1EaCpxF3oQMTvjzMuwDoWoDvd+D9GMCukT78YjfuWZKmcntBn6il+
BhiVGlayHhdWTWlJJpdoD3PfhHfefCrkqCWuAzqvnXH+3SFn0gNaHjhZD4eynH5DN1me0LPr/ixm
w+35wEmUMqnM0Tq1ANmA7Q7PTr5kL8u9ikBxfBhZW1GUo4V58A9I8fQzckxEl2N9vimzRvr2eIvn
Tzx5QSqwbVuQ95rUstMK2jq4IIwd+p0ck0GIMa7Tpq/ldF49mhlClq1rfm9LiKebj/CgvpUgsdrZ
+8ckQ8Fb3z9vGqlLPARRII3ut4Ov/YsiG2BUpAkbKXFNLMmfQJlkLY02mYwF55WuXA/O7kYoLqpS
+v3QtTubsJ5krHR7rujCXXcl3YZpvH8SngvNzNnDe7XsbVddJpU2SnvI5opaTiZvli66T59lWFBj
Y5Ez+9qIfbrY37u2sJJ0aTbQVGCrKh4NbcgWC6mJQHthfe66vRmwPwYEqO8kw3/nsDehUM5S0l4u
G20w9d0gt1JRWS3867xSCDUROQRbDUTeSXfuo067wqnKSCT8jVkAspRMvy63Kc9Xn2H3honp2Z6L
LbwIDkyC1czmhc3FfCTnPgPnBPvI458NQCoisYr47JM1VhXSCmSOjnacjjKCeY5v+/MROJ2w6utw
e685M899lLuRiv3WbwuxI6MLIxP1V8R+vu3IW6YuoLYm/JJRqCqTK8210s9zYAxkRBBk3PVRQi1t
P2kBYwC56NmueTJcZE0ZA/7Qd1otQj5B+mKXFH3PspdGpFEDD+mo0XTYfhKINEmtzRC3iAgvo74j
D3VHx2lIJDGJ95ag8JcZg1WBctehoKTt2QvMLQ7DGlxiUSMoFYzDK691eYx6FQmpl666dH6v/lbg
HrTz0U5tI2NIFesKQ8cNMHrEZJzAX+d42A8o6HHi8YxDsR2ZML8w+C1nMYf0/uD6+PEPuUO11GrX
eIgzwAYPYYPlFyWO/mImPtyV0lACcYRZz2p0njO7SlHsgeN9oJlURfumUMmp/Sd+snPw58ZHLt6/
QwYP6ESTp8hekBrOJOHaI6R3HcDieohjTtegzlcOKyjFmxquFP5BJAQF4Fkh+0cZerxZAYTl3LTK
FYV6HhN8utR5tVKxEMysDw/ItBrrg9p2phFvRqH1Yt1xR/sI8hyjsluInKnuKfKKQDdJNGfOgDRt
2p/SrpBUwOvGD2G0szbBE65cbVzvUMWNN/45+a60aNGV9OhtYzuEKCV1BwvWjDDoMBkI0HITNHj3
PoVxWqtkpY4pu0u/aGHMWCuvRZi0wpBsHWxWKyeO9hx6oNU2lnplHONnRSBB5MfDZZXs7FFMoB1V
iRqeOn1DHL1VO4qANgE+cZmn238JfJojwGjVCWTeQtVH2z1Mxyreqs7ivcdEmTrFXsTmVzOr/vEC
33ybxJ8P9hyMYQwHZ2kW/9sjN4YNuJZFIsUTkDoE4oy9WK0vPEJ8qI98UTcI8ulx7Jn0SOQM4D7K
hebNfHI6zHs3Y0ga4Uf4F1Y8l3LeQxZRWF6hVutcl9iXQpHrQjXqVFMG/mjbz5g6aOj+7vttH/TW
CVh1YZ0XF1lLWxGij3OjUJcbnZGgULSlB+lz10FkG9haKlZONehqgbW6CyuzodZD9e8Q39cTJTNc
DpeTwX833GbTwsJ0uOz+EibHmGddLr4+ssvr/A3E/tjBIbxdXga/WpHsbfotjLK8YZK1HJduztQC
FU5CfPYXzldBCqEQpjekEASavDQHmcoN1iSMx82OVs1Ps35q1+stPS//duaq6pKCiUCOGtfHjup6
nd5+qR6f7W4giVN3c+q3WEJ2fclNSJMyUgzfe406IphNJyxiRwG8H9qkAOcz3Mk2RHrJWLA4+6J2
3aYhsTLUFRzJrRejrj281yOYmkjJgOXK5agP1Qz60DjAYQMx6yfWvAX022jJ6rzRMI+4c3rcKvGI
UKjzstzs3GCkxg3PB78+zOpPsbclbKEIo7OEscAqtWNnKx2sqT1C/QKKTFiWhmCmOMl8/NZMAWXC
rRuwJmYnVyqqbLA55u9vbtbwck0yTMuTP8KIeqmqov7mW1RKPJbrIZScitDGWd7liTWVf5sItmJl
HZUmX3ZDG3qH+bmKRebuIjyxEL+iUvkjnIeqwhYP4uMdPTCfRAQ5yTKf4OjWCmlOebYTTAPFW3g4
xQy+PO6A5h5WBboAuvsjdFSBTGaZVuHT8x1jmQ0upBGuBu9aQ7kMKfvwQaPbkPJw2FvKGJXPQb/+
g/hvTf6mQApYtCno7X4ohKAgpX+n9+xq0LqqhymSDj1sP3ZLBy995EroSGpQEJXiF12q5vD82Avb
rv65c47e9nQzmz+L8WivDhA6ApeCtv5I6rqkxulW/+/DExKEZaeObJrMry9s77sQN0df2ybbMWgY
7Y+s0zp5v3K8/UPlLG7imN2Stift4cNJAeLyuFBIaU4+DtUTm9WNSNsf1OtxlnRX6UvGhkST3lla
LqmrQ6eC6ouTgn7W+xgQ8EIejGfKMJS6uGbsdRLqfu/rYle75X6/qhqvTU5riFiQnscZj+fv98w9
gWVbNByN0b9dJ398+au2kOwxLcYMQQq1qglWwMCI3V4Qv8VGI2w1KHbXl30D8i0S9HGxLkGW8Mkr
Og1u8mK1HmkEvemL9nSUeuS3OvWpFxDelb2KCSEzua9wXO2xiZele2aCWtSkFi182ZH8QoB/UkAo
5b2y82kEMbLAa/udIWOYS16b4JQQn7o6xH5KWCw82IYE0J762lznEqnbDc0HDHELEul3aS5kWQon
Dna2mqfDrObi4FDI2MynimfWt8wr1t5fkmcOCatHXIkkOfsagO+reFG14+RDsESL/6qqnRMMVATO
qbZD2m6OJUKaa4RmAJDttp+N++GcqgdTx+46rjq/w8tjDTqcNwt8FjWQzQzzRo3kXeEfvClmDp+3
+WVFsiUSCJgzMmvTHJ7PrV4+e3haUuQ07MQjdqTePzQaYrTwgydpwdka4tvWsWh9VZbXgTeCLlDD
q0SYXxn5mAYHYDohhFhrnNbf9dZeKmDYJZuiuKIIdYFJ23N+XCj895Mr8dtAKAJgtJYR6/cOnRUc
Y6vY73I17AyNEnoZtRkFMr0F89o5D2208yNbC5f/GzHYR/I5xRpK5Mi415LFezuqjvGGBUli/Q/B
gZcljy2pWWA94B2NU8jLzLh91SUJ0NbKokC6tkIyq9JayBwGZ0TeRP/4ql25rmIwnuwJ+2cnXLU6
VpgK6PdNeCu+zqrY9HsKbBlhGIdiV9D+vRvwN7lbS3BezvJTqX0rdhE9w928OYvCrjR0m+9I4i6C
0jQXX81tSkzPYHK8DZOcag/u1jjNJMumtVHVxN0KOz8A32MOY5El11o7172wblRBmEfBTYK7rax6
TOB8yJ6uSwJ9q4GS78kiZ/IU8DyofGckZUBCfONAMR99lgIkMV1/5xXnQWHS3nOlEppsBCPJgR2T
pH2t8fudtUjqgR9sJUOOx6FC/azQddu5RPwVH0P2scDJlPO2IMcfpFxJ0nMHU0EuhpZz5MKp8qQ8
SPrW8eHEFtaS6yzhl7hJ0W5TjJcZ9QNYYPilAEh5Mojx2kji4FhLtv67ZZrFwSJK7AfCnrGNhZnj
GK3ACENK4NSWVEcUTJLfLSk2ndXAz/VBDdEdfMKScopUVvWvz8kGcktHO4vL5kr2VXjgUCVeUXzk
n6wW39gG7eDqUU1b1wq0agHPsMWeFkK1kQTvWN3nV5Ejbyuh65iyqKwQEBmY0oTJ/+L6S/BapWH4
ZJm1CwaDuapcxZ2E8dNxt0Rzx9WMm3jjDAU2H4V927y5J5GYmgVqzrkHcC34pGXHYc9cISPPEvws
K/cBbLwSK/LUMv0Y0o+noiHyTm0ljp72NZZNmXavHGt6P1nz1W06wkpy/9WjE9iEWA/DjDpynC71
AbowsjL8eMeWwI9lg/auJaea2oLjPC29TienxCkC+nKQGAs0M1wolH1MpsItjFy+fN//ALcc25z7
ujVtyT9BNsm8QOKkbVlPuYbTkPaxVD2UHaxY8CwL8fKOwX7g1fF96Lan8FKTBNNFbY00HxZ6m52X
NBucHBN3CIBu5pDYFf3W4gNZJJ6FgPUYQ/7D2dFABhk5MQp6lk9MUe9XWFxmd5pjRQxbvxFFmCJf
wj5Ubm17QXmks0TMWtV31E37XRF3inn4RLTWcvdvabBqltZTAQSh7HBeyXhbLE12DIBqniMn9oIB
QfIb3FmhV1vaufzmh0Erf38GHE7jK7eYwUY6XlDRa7YjJLW9RQWK57rUGrIf/CuZTnub/RTXE8HC
A++VUbY2S9NCtgkQQze/xPhRGxAqZkyN6TA2tMNO2IxgA7CkMe19/63eQQ4vgcT2yoUn1hPyq2pB
CJXCxHVFuDzROxFW5kI/cAHkRAkPFQFd7rKcH5le1IUdIbUPX8N+Kbt+EfuZro23dJcmNZETgIDw
GOxpz8JCBXYRAtTpuYylRCmOCkk76pnSkfyuKUivsGTzxJ3zczBJWiwpWKWwsXDlxIeb+zcmIw2a
Mu1RHVWSSZY++3csqJbS2bKNJ5l00gkeZtQ8hR7rMw0fB2HVBZt+SMj43ZeefzI82QLD84P8UOWo
qvYIPb7IVscAvLibaKvlSe7Jx5h35WWGXDv91e7riZQMlVKrAacrX5XwPQocDqSVBAuLNqosU3rg
l0+4050TNKTjkuA/E8qTGJXxlfbk6ICyRD7DVtozVCZPHI0Cy8wxrBhXCZHbPf5VX6xgzLd1F69+
hXzL5xtPyxEv+8nmxkBwvDHPBD91SPesbedEbR6Dx8Zi6/eRekVk414gfZjMCwMf4pQ/r77p+qKd
mqAKoMnRjOWdQad5EnO1+raSxminWRYDrF8y5BjmU+DP9Aa52+piKcYE8DVwYbT1kOWLL0hJ/PAh
yn2CAT6Jc04foJ+PvojlmXw1wX7fq67DV/FcekMGb8yOovDHxmLXmOsgObLUvtc8x47SSEnXPj7O
wRXcRcZS+w7Daua7IIaNy9OU6vH/TWnj9JaHCVveGUsNJFB+2F2THe34NG6aflZtUgyWYwyPko3J
YrjyU3ymJDtoNVViEUphzSDA+vs17zd/xhnns0VDx5B5t4pci0WLSsQlKOfPEv4/DrvlN+cdRIBQ
zuewQG7XZ7SwzVXNZPHHZcOQmfMQ+HOotFBEfhio2o8EOJaoP4zxDpE9WAzEzFAV+2Z0TIhb2cQX
/kcS1j+rHu0HYLXax10T7ovrhRPTcGXgDqnqFvBDSfA0QCcHLKW93vs5yqSP/TwNqebyZbweVA0U
digu8NOcncrgtePSr+iWCdLrnHv3ehIj/gzmVwYOD1RqIhF7UlH+Kz4BTFqXK0+/0D2du/BL9Cw/
Pfr9ua25CcHQ5wO58p7cryooriHaY+Ch1XHy4dXJBtceYMdAgLhKg8C0J+qsw4Ukz5cWm12e8kzF
fL65b1tiwlUmS/zJIhi7Z8q9PlrqX7MzCu+cXDJVevcUw+SPZWWeKYKP9IFtTG6o4GLp3JbWQwfK
m1WYjEjRIoq39XBO5wc7ZSYortvdoekaZva8zJmwFXPM9QsoRLUxRdcepJckyk+I1kOEzr66Q16Q
YFFZPFuIj+xq15ykPDE0KOO7aZa8cRs/0+EV5PTUZnyyKOjvhHUr4rvX11ADUyZG2nXLOPq9Jjtm
tQi7+TCLyXDdpCf2qmXNl78aTlek2cj8XsKl/RTEWyiG2iUwC3rUmFrKr0XDzbCH8o1IEVAhrEC6
nG/HasouuTKva/aV3fTjCGfmjp3nV4B2g0IhMdbctTNXJYJn1O7IojDWsT7+u2/xtfpxJ8snTY2e
14+dair9wZ9BOuLueXwSHM+4Ha+C5bw4pY5UVJNpbvCtBADjxVnvQPMWjVEN1Qw9ivdew8MX2FXc
+DmauGFYoOTh0pWxg/icxhqRBnExzuKyLLr54ksSYdZpF37iBG0cK3TxTnAUjpK2+uT4z88LKxPo
DFufoX0W3zxXFZTvzuRH8nqxuiiQcg5ShZilGkj0OXKglqki50UGSpxocSONVx6CIOBZI5RMq5k8
vPZRtSW5HzctLh0rpp8Fi0taoIPp9YfmEVXogp014iI4snuQ+T0LuCIZug6Gsx5YtCEfdPZVP2s6
SJF2SZAVkRLxjYQ2PFjA2n3Rs265h/v88weH2BImWyAu4Gvnjk4xrqSex9CiDNuJmxHNHSs+RX7t
DkwzsDdbpvTHUr1oam7hvIcPYi650S99RNLBKGJdhPTp855rAD3PRwdpAB8dBuaUfM10c7BiWLE9
rDFTdEtl1FRgIYeFr5Nf0LmAoqfr2YmynJ4N/8smWGjYwzSOyQn0RJStuFNaKpnp8sDJ0AO/E97X
jg3NB3b+ortK1l/6mEi7/bsY3QC6Z8fuiyXD6Juk7CRHxF1YqWwruUTjlEsl7SqvyANkICn9t4WX
XqfHAx0JSBKZUEeuIQBCrik1GEfaeP75S+UzSJVF3os1ggkC+c2t2lDfoeTI4Iz1ivmXsiaeLIwa
SAWebcwkOB0khhzE4LD4sedm1RNIBYfdr2I3iaf3cbZKSK+L0iqkidOstLPIcjjTS4oWds/Mq85Z
XeuFFybU3OuGYVeTHc5/oMioxdXM6+qK/xg202HqOcQX1+ZnHQH/vQR7WHE4Wu9zWBfYOtRzVQ3F
0h+qYlUiCg7aKV9z67mQzksn5Kf5FAQRWMuTEgSCiclt/vawC7mVqDH3OdFB20owVN9tC17dvtcm
Qc+InQXx3IobO7855loNEW+btUcLgxVQEmTKlko31urKxU3cATsPu5qp5KOMlcAUS8x1gH1d/3v9
pXEZ8TW12lfI4jwR5wutbnQ+8+DtJB22RKPy7guWCjsOlaAVBc/AIFfN5FAgGsUOZ4qGn+WQul78
A5Ql1hLscbb2aunt+TvtyCDRo2/F72wfDB2sX+wvvrzJEJM83vJaiFip7cF91NavPM5sGs5481hg
9F/EL8GHZUPLumwKOzDSJkOMof+P8EIeg2KmmR8sk0otPnFbFQpfDURuFtABGzDQr5Oe3imm6qiO
J2xxhve7X6+YTyycP82V623lcOHPNL+Zz24eThGFRqLQn+crQ7W9OJn+xvCMvB2EC+A2LcEOi3mq
EEAdPr5FDQYz4yEhZgWxU1XGmpO24RHuCDRFzI22WulIkbg/5Tl/XkimNaCJ5NHFpn+GZ8lmYkXw
Za+jQU7FjpkYHxm36bRypBKYwpyHqbp5/oIGmOtqx8ZLuaP/emKjUppw19f07YOUaQ6CRLHEagV8
9hGKZ7aYdqnxAaZUlp1UHlMO3B/uf+XZYtviTfPDEicpWbzbM9xLRroDpvqDKnTLX2xBLI7qp+RH
tE/7PjL90sIM8fxTZwe8qSdV3dLIDrOHHGyj/EUR3ko5KShccen+CrAJTOzI3QxiqynRCF4PuVMo
j8uXWkU+qVNSquwLEjkSKgx6sFL50Q7r+LA8J451BhCBOOyd8Rj8KpFcPdfozWqb8NSuDtSvBRlS
jk8wcEdPN1Aw4rjvxF/rK8lYu/Q8dUoBVbFb2uAKxvjM8rJ40u4s9GJ4IWFGZWIhqeRdaZ8kUnJg
k+6s+/m6Bk9O/hcoqakb/eQ2DBOycBG+HhrurDMmZyVMwMqgDV7NTqo4dYAFOxd+yDpLijpXNqqH
FdAxPPO793n2jrtmlQyjiWZXn/WCeET+NOT2NJxn8SG5JG8RuFfQp6ggcxa0KtZLggnNc6wpuwMt
MLbL2Z4FKLQlhBzUvRc+F0CVp07vlziT4DC3xG75Hb218zbLyZMzd8dV1E0cDJb4W0aIyqg7NVnS
KnENkSA+0rbpwpCaKMdI78rvy6ipsX0c2zCUxeT9KoDcM4mb6n/jOXU2liCpeF/y75Ua5S0Ov1r4
PYW5izplftsgT/DT77pnwB3KZ02v9CbzgBxn4m7DDCAaPmaRvy9BhwU+BtUJzjYiwEuqMjqPteJA
Yf/bD4/KeLcVkWEaNhe8H+6budERmX6yJV6c/Y8EtiWY9uPx9LeL2JVQ532ZcAOmsfj/aAhttkG5
1emgE0om5hly4RjafoMIIorvf8K6t8vwZBoJJ5XwnWKZBb0uIk47/p69DM3BnnXoBhpfEfqVXLni
o0lCmKDO2xu/auRO3j+IJVktvzYtWMNtS23RhUezZhsg1ZO/YJpIgYsR1657FOQATmVPSXOLy/7D
/hfoDGdJ+BDzkkfOQ7/LEOxbxiC4TZ/N4vz5CBXiELhNf9Aa6g9Z0DjzXkK0CTvmrLrRwQR0mIiy
aDvUODRfpRXZ9gSTTxRXUM4GH9IzNF2pyxJvpOPyteihsD2QR6oriQFgrvf3KE6IXrQv6EuzSAhh
fIgDc9PgtA8JdgR43Q+yJXGZVfXCveMplu4FS3TMuCn5aBqAT0O4pDQSock4F2Tqr3A6Kd2Cigzw
wsEY6pltc3jKWZ8HATNlV3/xX+WCHbRhVBLdGghxozL0At4y8+pGdDjJMM+KWdyiByGZ1kJHK+Id
CYl1f3GxjuyxMY+kciPKcIngK1+u11zee0pRDoP4GxVb4N2//fOMWaJyOO+J+fTk5gPqL8LEpEV7
hrTwmFmAcihRLZrmXSqYzWk1hRcYfxgVGS1cnGx9Mc9TjnvfPAvM9rySPqro15zYct82GUhkY5KC
hx1SO6eW9jxVg/yCOaNbd1vLImpdLgnV+Ti9DU9yyR7pPrtEKOOFEENryaPfxjAzTPHIegUfwTMC
TH5vWhNZSps7mDn+4XobMUjll+s+xB4TgfhujcEbgH3pM6nv9BVZtxZW4AuvweGPjJl8i8K+9902
keQnw7BbsNkJ8g2zhptDmJXkTSGmdV2yYTwYRji1ZbByvCENRxIwLFAUq6YZe4AUvq4m7fagSGow
be/3vfXQD3mfsmxKfPOFdm5KHXg83sF1DFp1LEceOWi9LC2EPSFPT2/jo2aBfl0k8E0/GegnmlYV
GAsy37hFxdjXxd6ppkvMZf17OYZQPCA7xZT/126Z+hktuR+q8GVrwOfwuoHH+fuCIoI0XkcColDU
M0j9Y7S2oAPHkb+vLTDtoi2gAxE/Izhw6hq89xUZDKaxh8ui092ENyPzcNhWg8vV2MDstG9A0/l9
ypfDsjeDye7b2peT/yzLrYywnwTIq3myXX6Zhcx0TFGEl/HEYpl8qZ9dilOETx36w/q0LJhXAgUc
XuLUZGltB7A/myhpemilFJ751pJ15LL1jEmszwOgmcfvlgUqWAc8xP8QU9o/3DSAcwn9a4hvOTy6
79i7fcYKOA8RbPLyYrNluiCJU496PPdCxdty81/H8C4nZS4kGJTYqZb0oqHUFOjnLnNPKpBaNkCx
yh8XmklQUTZvdPDEs8sZIFwhvEdyMQCJdJ/s+Ah5bX6UGROyF505yPRdlAJxsX6AW6/VK26RwtJ3
iqiHmBaYevQez18+ABbvp0KQzGoZ+R2ONiUQ/JX26dxRdOrTnjxMF3AzN4KwW+SldQ/Vc7LN8gF9
oJnkTj3kMSMhsnoNgOdJ+uBKeq9AKBT3IzY9c1iPYtkR1Y0t49SBD9/gwJlfS6qOP37l/+PkUOJ5
D+KznuQsfBMVRcCCveOSRqoGoCQCpVK2ckgjigccIrmLgEw8/vZ880iKlUG6AWtDPb29K2a3AnhJ
1SNWLTIP/Iff9uQpTjFSbxE9yCwHWztRl2YQAXan5HybBQCxLzZ9PWcqNf4miktbSMaBDT8fqUd7
K8FHP0kyy2Ce0XoFBp9yOhFJOqunQP92lmrAtJZ64WjwjsXWzK9Oi7PrxRPtzmqVd0hZ3+wouUYg
8YX/H7uw4teznq3xdoI/t3m6CmQZle5uhxdFhh2nWtvbVC7yePgIdkzucZM49QLLXjB2zP/EpOnS
8b+lm0h8MfsKyArFjXQoXOCqr0vYJCAxmsql4XCXq0uDbyUnvPgSt0Slq8cFsBAD8SVJm+RZPjgP
+jUkx9/sDBQfYl7BktHziQXN7P/AuKgIUZQgjYJRF0CtcIpZAHQdxvuJm14NqSC0ea0egAS2Y55h
2GuUc7vjaFfqoyL77Y4l1yzKETukaTsQiOp97nNgsxNo1dAq81qbog7m9vXfBM4AcB3LO6+wu/qY
PhOoigQEjrn0ZfJfVcqgAOhyHc8wnRN4cjl+Wj3ycYDHwySP6TXbmN+QzyOl9YFtHVQB/65qhGM3
kiSyJ2ICytp876g8m4hzVs3XfHJjAKacHTJgqMlP6SQjzmDbZmKP7yK8VFwuqG871Jyf9Ib4xdpT
mg1/2vSk/blqFeShCoZfm01DVxoglN7SKSk3YHJx1+rCfdb43CVjeoSOPu0ggmPowDwdsuo9p+E8
r+IakvAMfe20DWiZqsOpZxS4nTFfP/b0n0L5p539ldSmbKLRiEVt/SwFyd/RCZpuDjnIk1bB5CnP
aIqq2jHdmD60mIQTfk6bopvxVtVZlHS3aw15j4ehS23xrOFUX2Za32dXHKs03r1OXuAv3jU2RRQN
0So2sfCgSnnlEmq393UzovvAcBMfLPS17xMN7PB5WoCrey1xj4e8XVcuAJVgaSRuffDBg3TbQa43
OYWSqK03ba1jbW+gI8BSlK51TCE1gYHamwI3FDdmMdV/YdqH/GP8Y40SCUZFZnxvqnRj9aD31+Zy
URLYgKtFmJkkF3KOCi8LGNZHDUtF7KedmWZGJD9SwOG0kISKe0iTal+wT1z//jR2T48e+w9nDT3s
cssLAOTzcGE9tlqbHcijHgkj4lDho4xPyRIGZ7Gnk1c6mlHZzko6WjE5HOV8CgvL9TOD2QZdIwOO
lDb23cM2EXR+DBJ5FLZmP52YHu6AVL5y1A03KBUytK09c9d02NOPtAVoEox0eB0P6sSQk3qfAFVb
EBageiVUkRnSwwV7z4qK3PLVpnGUMjUP5MbQYYPxib+tKvO1mzy9FLA4BItPqhcllWOvkJ+PtnLV
8MtY7bDnsuHX2au30KARbZvjU2iUp0U/2jl8EiKmfgmEx3vnDQyBtC/fQyTiane0VJd/AydIpspG
m9/khkGeUsPIBzbE3auabhNQ34XDK2dEoA6rBsPYnRMFSZjt0hIRWm1bR3ER6Z8NoT2hQANWGuOd
u1tD9y8nLPAn8B+fnWzduiSAkHVHkbNrC1i4C8GtCww5nJ6PpI3ewa4wn3W0V7kruh24ZjRiabYu
0LXE5mxfl3Quh6RtEPE/3co3fJdv2cIbKXtsQSeWGUCgQ4YzS47DDj4owR1DsVpFXLXR+kEdX/7o
vhnhhKZ6hXXZ8X+Z8u7j6AKqrKznv6/dvgjNJ4zP4z8bsb26x5Odjd0obzBer62AQ1v2enyosjIQ
l7YUZWLIyO62X3z8pLTwR3edqw0diY9hXUEKD+iq3Xsn6O80UglOd/SvJ93DaZ1H/czvS4kCkhYr
bs7Z2mfnhoJroiFgSnuC7lAka8bLUaWwkkTDDnjaTJeyZQQGC4vrn/OBMZeyJcGLULEWqUdvPjSz
LaU0FMgw91NSdl2Tg2ZNtuJXP34MstwQnZQudF04XdIAoHKBWHobg7Scs3YKnKWDh1WnspK3R+Jr
2L//qxdOBheAFvyKhyfdd9Labf9YoxIVB7dM/mBmrCShUE9WEoWg9xZleCTdmjhN/BQS9iNYQx/z
/dps7kycZea2ojDCyynlPcpecX1HCngLRGREmi0167DB/I0uDxkdiDInTKstWaYRLGweV+KwUOQK
mPd4BdE2CTP/QGvaDiO+3nvpe+8D/awL8+7znBqyUhlv0OjDQMyr8dnwdGJrCH4htiWsb0j1L3N7
dTrfkp/KzQuKzijF54x58MVENObDw3l6FDl63f72BcOdTHUeR3/PICL+Ng+ZY2X1nbnz+tVBqyjM
weMBKMGl4agvg/Kf3CKBf4NViPZwQEbP3Yt+R4tsP1Rmk1eJuU4ewfyVJLBJ1ZCzal3IWX/xKoXR
CCW/WhOHYfjxJYn0cFzhkjHiCeQUAgoqoXTVrdHpC3duEDwWx9sw4aIG1CfxHx+FjuwcEQmUJFfb
5e3qLXunJUKugEEy+KN7erj7uXIjWJtTWc2aWXGlNaz0NDqKke7HQFJm38Y2Z2XDccWqeoHD65eO
+sqhYGcTU9+av5mqW0EEeg7GR66BetqH+phT5uw1BJintiuxt4pjdQ4efi7N5rXJahmu/dVqeh7B
hZPFo4M/ewWuBM3GQOaFvMRitLkTzeWHscNDd3HtgKPwssrQJdkE/vmkonJ/khDbSuHsfjAdtiGH
5T0mac/oSh+aVuEAWD4YUdDtVtEw8IMMz8i6yEtABx1NiKcvmL2vjtVh8zmmJ9v11yPt2AtCfsDj
gLwNR+22bjP84BSj0B102AhEoVF2UkEYXFRMnoJc6HB6BpYqn8AdpT3hHUfaYOLCMZhpeuOumgjP
bBf79mNefhNVcV8C7aIIuFXLJBooCkPsaKeLkf0MMjl6WRFq02wae77J0DWc38NWjS/o3X1YI/Q6
HJWxdvKNoAXOGqg2vXbImvHVCXtAsQeZe1uxyFa6JRQZqi4+YFjfICkARJrvpfw0hQ0XDx5ej19q
s/9tRVZ3ox8ugbTnzgqWJlbaNRkvA/6dPnxmn+xmlXTrYe0/7Mz67pYWMLVEV3WZLkc2FKJBy71g
32F6WBY7hh4kO6wCn2cRI9JpOAhvMhzliyUPmr2tD1r+4UWje1Tz42KRUeor7f04Rxy7Fw+JnuAp
KusK01CX06eDN1mcEOXFVlWIpMxc9IsOIq+lptzS9kLL+jSm9xqkizwJINUcJcH6cSXpihsUizwt
SMao/wd1XYOz52bZa1nMxaEMI6YqY/Yncdv6bfocnhVXRy2Vnq5eseY489Ix2FIGteeBYcTW/ywX
yRJUl+8mXIZTA1ClNqepFpG1/igTXQSYJGJqzsZIBEvxskWAsU8SBRlHV6/y5jX5HX+AVB1Eu4wg
TjMxOiNjGA9JvecudppEBI6iSBjAb1sYzFps2ew0riy6i0aYOlL6IquZYoS1NurN215YjTisSOaM
hsXImGA6SpuH9W/ocpU5n8k54+P9nYBZuX7+/VHIiohzbts1XHzZHgvPdoSn8qWh23wcdGb6phfP
GLa19ckeifoTECT4lbLFYDg3FqLC3B6rxcpSI2pNX6jxpWw8upTKB/ZVfSsy/Y3tBLmTgW93HpKb
W3mLJ4HYKML2kImrJXL3RhfUtTY8JUnyB4WGI1r0XkF/KdsKrG/St6kJN02G7fbpAzh92iLDCj4q
R9k88XXw8x5MA8K6045ydls8f1/B5p/SdQNOnLmu3wT4bkGyX2fEV7YIpG5nFHMiCpBAmEOGt8au
1FDGuPz9t5Q+IKZ/okCEvigPeRK8ydtXBNi4SUL9eZPrpiprCdaQvOBrkYKxq3PXdnvSOLVLEe3V
Jif6xvOBL7XybxS2x6J9tkQQ18BDYnQiLxwfqxhS/lDH5kTPtLGFzUESh8K21dqcswYq2dLxayvo
yOthEh6buVdqLlnkvY+Fv6qqhBxdRHZipOujvS+/XIdtEwdBSA9RLdAttyubVU4fRlpmz3/LMwA1
I8D+v4fkb8ilRh2ROfwU0NnJRb9IOSC8Crz4+TOIkXzpGg0JVzqgoTjnfS0D10uAuOXhZoweQzk0
LLwBJA1WJVv/0jl3qhJ3+judocRNoz9k65pfIPrFYl6T6WT24dW0RI16zMjxKfWhDSlJBQI0Vvcv
rt2ealIzqoLvFdfcJ39p8OXzBAunRbXB90EtrncMS1QJPwnT6M2w0IpHsljyMlWrZjbK9cZKTPAU
nTLcow6jv+FVvxTxA7xffjVmG5vHHpazejJZ/m/0HMTwSGHNlz8XhODXi/QTNj4yr1JndUByQ2T3
LKFAt/O+OdLMaAC4kSMbGAQ2MjiBr5bmvO02Bsfu5nbQa1ldMIevw4P8r0upN8JzyajSsTaLPBPD
IvSENVQh5BAwzeA3UF2iTq75Q5D7EWww/pBM5PViahyXnybQacAd3tHadAPr3uosTAriLzOuD1aF
8OzMVo5rCNj9w2NWLL21YWM6bI333NG+faCA8K7wllAl5KRzk7rKcjbzufUnQUuDMpEU9PEjomJe
wKK9iSt+Mmot6IQdVpVBtVvOTqbtFwZO18bkeU5zjRwk67IYd4+8zep8Oda3le0ONbSznCAKKuxs
SiNKx9ai0W2YKf8oeBYLOitdDf/RqldZxgzvd1kEnkTgNf2iAAtF5sSBP/rmKyora+SoYeKrnrUv
+KshYJ3bmXHF+66HA8UdQDMfpkg0/4SQ6dCHCOZbnzZxNPL+yBDq9fY8SOjF6yLrULBvOfUCQpaI
tK/WMH4gTDxqLuU8DPXVrA1zfI3SpAf62VL+3hndr2oJekWT8o3cZfgrQtfWt5nT4DSgFGLdTwrf
k+uAU1oNDx/+rTVTnwhNF7kxJt/nvnzz+f8898y0+OWSyuuJjQiX1UgS0XX4AMCdGJ7pduT1zFPC
S7/YCYYsc9+rMqZYdznRR1GCawOP2GcwMzh4PhMe2IL0IuW91tnuD1P3YfEkyAN9FhZATyEQzIOK
76EvKtrhOKM+GMnVDzDCMuI7mZgTxZdnVMHM29+1e2Suj1Ys3HGSlSnd/8kKmJdOZhqes2PRmkTz
9oo18LyRImvcsVht9avX2t509eYucEZROM0t4f+pivR8tn5QWklwFgz+542rrFgsOEDoJJoptE+L
ajpBtTbMDo7KrlGoIkS19WJRbZ7tWLnyJPKwHMVxp6ZKQjpVwpYe6XsOnJ2/Mbq8Nce0wFq6hk0B
VTmQ7vQVK1P77G3Eaad4UOGOAtjtFT4EcNL3Xki34+cctwz3mZ+B6AA4bSZNcDeSeCRF8gt7PZU2
mAavMrbMWUdLToSs0zwqGlnWcigIfZ2C6aMEieAWXcsiu7vnY/PKH2n89HvQ/+ZWfVl/DYW2fIGW
7tork7NqaIFGZRfB/4Q6MUSsAdKlFhFv1Tz/ohbbZdvKtdvxNb/HoVmBHrY1Gqpon7RZ1il2EkAd
pnXPJPzYMcMTsloNAJ/MMvMJ4G9fZCel1ONg5S1EGWMbkpkGSTKTytmyGtMlx/cbL8Kz8WGkbm4Y
mQD0dSjyUgLu6UBXxwOD+yAoTUU53OGhe3f40RiuL3yOGnO3ci9MizGo4rXgIYTS/nnCq+NNU/pM
upxWHnbQ75mMLzGFFMm1ZCthN6unZGwl8TxoKgYnc1kPd+U8eS3yzr2euGlz0Gu1PS5ss0tOiUcm
8fIEEwCV2vVIi43rZgk8xhOSx83U9d2ZLjqh69QFwKKWte6YkPA6RcD93TEJA92UtPu70BWox82V
jOMq4I5RS6Vc70AgMI8XyjPoacLBSjqWN76iP0jxmhjKmFhLU625G2SndJqoDq8LhyYsZwx/p559
VzkS+WncFSRBXV+BoQz5lrQFSV0G9I/LsDA0RhiaJVmsu0lx2bmiEf/wz4hXa7FSqvhJe/8hAwDQ
dZAFAd9EDZtJkbq0zXNQ++vP+GWam9yzqO+XzpQC5kyp3L6mSnB653nYDEuYnFiIHA7qaQrxyUHz
8OlSNCPXFbGzMYm42G12wHILDQ1njkkNZzpWc095WUSPqx6Kg97iUTknviRUoiq5rDTfewX8w9xt
j+fWWq5+/bnGXDFELsRLG81t74l3OCs9AkxcvOJot9GtYJBCEmmMJUrQ50+MLrvyuyn27okMlYmn
W/1oYA+jl8TYYJ6dIqkGocIbGub3ovG8Z5ZuhtEpUCvE4b0AHMM/ZQcAKTVHjmZTNXBbib3p9nAk
tjfgmJ2jhPKt4twVsAwM2sUoMDju47p5KWDxpU5OU325taY1DZP2MfZ+rETnfH19KN5ivEQ1Ya6e
UCUgLo2GSMAwlBHHphKWXPJ4f/Jp7yDB8D/+o+GDoHzMsslRjQDbZJLSZC+H54/oIfFTxu52sM84
ARI4InV9QAzhUdryQzlbqyOpWBMlQpIkv6rGcp2NxGJyMNfertbBFod0cVxZuwy4MaYci3v2Zz0y
w4i7y4GDJt+kxCIQxnouGiV0/KNHqEvQ0SET5xxzNYH7q0OxZSR0/sZ2KU5fDQWgHSsi+/kLOQnz
B4lfZYMnTcuXxcuzyTTbNvyQq24yFm/c7VxWQVr6a46hwhzlgkkUqOLi6DOH430nXPfiQWuA3L2X
8zGBJ/E6ghgq+ZHjCP9HCtbnXKxbqISPgdTU9JvyI6PJgmE+gHyTFfLLt55UhRQhzZG1a2BoJ/eb
TKwkH8YhI4MI1IQr+4H3XGEmyX0dq4qvttYZ3RoINTdLmoszJIEHYLVIgz8t0dltSqQScPJY6a7D
8jmtUecG5HHYt0PYKZr5H6bUcYMLZXuE9EY/o7OOq9Yp4uLG+wB3N7u6rHFktnff7alr42XkvVGx
kXRfxplfeeIXXt7uvAyRbbpI93uNqcwui8sjVTqRK0G01B+nHeK6Z27j2koedwz5YYeAoTORVMsr
NCNtqncmysRBdVOA0E441ACpxKu8SHZFp3lCxhPQIq+2/KUC1q8tg5rhHOoa+gmfX4rPih5nb0HY
Yp8SSI9mVH7sI2s9LhgoGnCCEDz6OOBZ3g2C8vDYctDDl4YalbETRXKsYBkwdmb+AjnznJ7fHRGl
MgDHtiJN4eh3ZpnbeC4SmhWfu8M+W5dOhRx1u6RchmA6iYaFdbRBjUS1lJyyFsYnBTM7+l4zv577
67cqDayWtsEo3ejKlNw2Cs2q0tdy5ogknHXbTbUjDvQ1r3C4QrzD/Rnv+k4vE3wrtzagH2kybMNc
7kej2jD8zK49jvB0S2tVQtNUbRUO+sbEEB6z+Hcsq5brzxrK/ydImzmT6kfff54eO7TQ5IIlPQZY
9yNE3XkySOTfMmjBwwr+t7BlndJvQUgYW+Be//pjjY8400ykBc5v+/93toTFCfsLYfB1GiV6L0Md
OKwoxJUePV5aM7oDTpqHPX8X9CLJU0ZSTkFn+WekF15VrWTlWGTBwHTH1NapkwP70HaXXxoBDYfA
POh9k1SeNU93n51lQWkI1ZACg7c77IKEa8vJk1CJChcezp3P4mFrlbUQvHMS0Kqq7g5oDkGGfiWN
3myN+537EbU0Kc0AsKFEUgdWLS3VKwQl8hcqY9PmgAJZjEe2LBFIjkYdvNJqrbTByw6bKfutOrXX
tjobPLDyCLlS+xH2gywCYZ2etEbPTJOzhcOXX83qYN637oWEer+nkf1YmyM6oDQ81AsU/DSJRBtn
St1f99JGXjuC4EV7HS0eje0skAkoIsHbHBSJT9VchVCEh2fM9X40AylrIR1k7lx507lkno/CaVgK
imt0D2IcUnLIDSmjBeZ7TSRtGIxulmIyp1PfI4rgKFa9pbPZ3DYZltj30S8UFIHCK4yuOn6e5/mx
J67XC0yipLS0MeEKCMg9mwxii4vaEMX43aXJ2kfxdq9V9bSbYEDyO4jXgUb5QH8evWbMw8+erCmO
/p7ZQrDR/fuSwpiHuqoN1kxSm5UyMYby18Rb/Pe5w/Y83MR8MRvZL4VWKzZQYV32Tl4MPoDHHNYs
gq8/NtGPhUrofKhr4HkFzBU8NEF7Z1xKYLUa5p+00Odz6G84IxhuRmuvKQ2lVaqkvssxbuh7SHAg
umVuMHi6+LL9JXfzGnxasYDhQDFyGe20T+2FstH5yrpksAtOMKpj3/98qDg9dqYrjaW1iLKsaIsI
Sk8YMPfKGrEkJqWanQehsL4ma0gKljAR2OMFH4YATA5fC2K7KQL5FluOTW8QOhjchVWfbMirKJsP
Ps0LIrtZi6AQN8pnHKiQd4Uqtkfhxl224Lf5Ey24mtNku/0CWmP3kkfKImrfiI1nzSTtnBtIonzo
OIyEc5dv1DG/+9yKT7if9yeV20mumknF4iNlmnlWnyvjySb5ezAENrG6IbJLWuAflBRkd9Ou3yWb
1pGtnGZe7UAVA2LghDRGvP68aCmH3GfE2CqVqG1NcDVpb8CTQaTI8i2fo6/kVmm32JLfCjyWiKD4
WMZmZVeh0+7VKB3BMpJRWzeHLqfj0hXyN5tLMnmw79ksRxD6jbTm95l/PIs3weAUAi3em5hph/SA
rgHxWEaAskGA/yl8TjHkI4hUYuWgD5h/iH2FFchFz6/5re9Bg1drvWN2r7Mwat5QoL/Jm2MYIjte
658IxyHJ9amM9JF6qlOSjp4E/WUEEAMaZhhly7vJlDbbF3d7Xoxdo7N4UInMiRLbbKTIl9oEiwHR
WDIK0l+DP3H7Q2TDXft0L1ph7J2MqO9UNF9lh+mnoICJMATpxF2Le44SsGtu2MZQ14GJIsbboQPv
JExkjTDscePJIQKyasAmd2cwjCx5CPlHBHQVGgxmgkiy33iXiToHG9e7UZ1cGupS+ErKBWxnS6Bf
YPdVXCz3HVu7OlB5Hc7xMNhj0DMuucyKsS+uvLvKVp2hFEV33ddErQ17v1xey0MUTCW36fq9kw7M
iieD2gEXF6TZC93YmcUn4Nd55eMzYgCXkp/mKFeJ+YWZM1XWLjuhZmoMaVpiWDqBgKTKQPUWteRD
oLtn1h2PHwoIeJU4/tZubHwaUNsO8jYB83iLjO3xY0icAt/aoQKmAOVe9aXyfr6HgSB4ar03V7Br
ImdYcrGvXYa9fjFxuJnUUag0RAkf9n5Lp3DiYmNk06Fy1nExYPqOzakkOartasiNbGMg8h+M3nJB
TQnFQqCS+N3VuAJqvc020Z5wPaj6RF9Uq8aM9A8op3i1Fi4EXewwJw6ENrvWz9t1Ae03RfUcQkAd
6Imave3IU9Jz088AaQ4B21jFDz3bMD4ml8D75oYSrja2cXG0cWetMDX00ZghCIlesuMVQNCXZ2xl
LI3Qez/IMFX/e89K1q2+D2VhrSWwHKkNE9OBJzVP4cfx/Q17GHHsZ1EMgV584axCig6HlJhkQLgR
hS9YCk3rIxeYzogUxZ4QYsViiYUj415yEui++5IEgJ+07/bj8kwIJzTn4vDxO8m8vLIvcx1IV3ju
NjfzpLcIxs4mY1nmhWgTmTbA5TRCJVXRXi0yCwcXSHdbOh7V5jJPN6VUc0J9kHgaAVCWW6KfTxPb
cQavXLgu1BxPlOAULepgLE7NDaU8x50oXM6tU80nPSGIOd/7MKtnqdVkdupbo5xgILDIhAu+Sd+c
iHrU21gR8UjR7V5lGG8xfpXZksH2wjbgM514ltYWQpplF8LDlsF/M9VgUeHJeAASxsD1yFEDB9k1
FJia0GUjJVdu18j4X5MD9KCYsA96tkEACUWW+mMHAGv/PMa361nWfbSd7+/J3k8BXE8yarEkgLhx
grrkDOrSlh/iFHjkPD6ROxJoKql/qQiHp8AGsV7Ht/VwK9f4zp6kwMlKePvOCSQDDsPSlyG6yFm3
h4t1vyFQycCUcCYmquPDRZj+dfGWGAbs5AVy6RFUJxLrwmwBuThCrKyJe/5syFsEJgQ7EQTwV+Ve
SdTjMLL8SsDBLmMAv93/wdnR9HbODQi99lEHvc8nY59CrfSebAKOmFXutm3PAJqVpIy0Xzdx9Atc
+T9g9nTnhY+7D4I/+xKLnlqYKktsT2iYzINObu4zpZCvzQQvDptLJXR9N2u54kU+LQI5DohqbqQC
NcUp+q+pbiQjBH97rOO9jxB8NNUACiMr8T/MxOZYw2M+A90fPTodMg38kRGRc/6f8f5ZUJLwgWwo
SzAbZBELA91EE5V0mt2SIhobGWcVxXWQFuTYwuTIn+/efJ9gD4PcoYOUe9T8xWKuq2Dm915j6Sq2
2RvYWShT0AorYBF8pBLQeOaoQ092+G094FgtzHMKu1DvkqgLuRINIOEIwFfVyItEZwNY+ES1dVUm
oyphBBx0cDaOz0U+dk6VCP28dqtkfgDZ6KsgCEuIzAwLcKSIrRUetWlL+y6+PPafr+pN/YLmIsjp
2VCvZmKEDDcWGxf8T2afWBFaTxWVvwLVZFn6bh4gjuyXayUr3+UtjS9Y8y0NgdRg3qmDJXhGGE+l
S33TXXZwWsQa+MVdx3pwYg12yGDxHY2aAc8u/PJKkkd/wtzxq4uonY1cgg4NaAJiXKkPpBt9rAIr
35Uwaj/ylHYWe3vfOByJxg0t8YcVKhWqrbN/ob5IO14+5/uWuG8Kq7CYmlk5HePuUBq+uFEK9hQ0
mVDXcIMnRM9OGR18tOCF76OjdJb3hivlUk+0lLxd3k13AZ9GfvKAShnCFR6ZW42fcvKQJidYSGs0
esFVcIhrtHAtJbKc9iHU+ANwTSWgzKI8PsUtcFMSz9iKP3Q9QCiG7NLRaGZ59L655qMX2R3bVLur
kYsS+v2ueIdp5fzL6S0fmIdAah/v7z/PzI+3KKvomTI0E+gqnUZJf6rvUz6ubuKXwUZz8zPFygLL
9bRsiuYc0Rh7lcFdsZEwXiSkfLAiuHUUY8GF5xCWsSkPVU0k2JWUAcEb/g2EGtFWZbLLokxB0S8X
Ox/n1x0P9RG+RvF/9faeOeK4XCcRxcJ2nCjx+yK3le4zlF6ARUkzYBheFHIwlg58eJH0J2AVKjVg
aMeneT/4fLzHSwQjUCm/UCASnpLuMNhh94rW5g6WSqxJPp9SbJIUwfu9woVRZMAd1TTNeCI9w2jl
Xlb2PBaLbxcEW0evWN6gwW8q5O+39Oa9XNj6WAVS/JERHkjf/rgQQV+TqCKzAoTZjOMKksHBb4bg
sTazZxpjzga40QxF7yqHSPEctW+aIPAb0mLmmoxH2I3sJNux7ZJI/s/mKiNB3xpkht6i56QGFR2T
5EwzVl0xox/Dl5HCb+v3ggmVgDJozvgGJMtAd4p3CCRVlKyiwyCpgDEG4j1mXwhXnmgCKcqDHbzV
hLZz+TeNoCxabxWI/RzclB/3QUg05hJUkanIugxaw7OOw4YvNC4Opo6pIZmMIOHBWG4u8nJ89/fj
NEQiQ9RgbV3+UCvTAyKq4QkhVEDODZrnwCbUeZSMq/a91ycmwe40D3Aiw+X7Ch1bBGdKH8olEyFQ
0S4umwpwHwMKiRpgEZODhm/aVRQbOrSu6daysLSyZBK9wh2a0OdBjUsDmAVzz0EAGtpkjK6zw+Lc
pq6Ykw7NIInLhau/Nj0xSslb3JvxqbXws+OXXICU84Etucn+tr0VKs4LUJp+2a/y+OAzh7ABVaLK
z5JcaKOLl2syASUtsoIR8u6k9GH0Hik8WhA3mI3rqL4T38lvdd/kj0O44GTocrhzzJzSAfCpTfxX
99pn8Yi1KspYDcWCZQlEvI67pVLINtnrc79bqM74VdjrgwayTFTCTQ+qyktAa+r4tUaxxROR8lCY
lHW5W9mHPW+BfFM1tMqK2ZZ0Yt8EtzbratTVhZYHSmG9kgidGLCo1lzgaMxobZ6x1IpLj3KaMjJ0
rlrsHEWPB2lTYxJScszF7O7vKXvI4uWO11+z9PjdcYcOfZ60ZBlWqoEgoHLaqNvdn1d6sl69rQ0f
6ldez7X8e3RlhGwVKcgk75SbaQ8sEVNIFtBGvIh17IGFsIJ379KQ+vD4K4mtq2nRuBmA6tVBB6m7
VDzP4jwVvYVzb2e8tLhzB6Fle7pawjs7RzXZWeCmzCxOs0ldmxSWQbSJ/lziqnU9tgrKVNugX1nk
ejYpYP+T55u3AndK/xnFMQZiETUk+1UtTceRl5PNrAIAFPmLLtfAsFN/8C9+gLLu2ydWb63EG0L1
WkXEbbg33qIoY49d8azsoDx1uMG1Duqu3kOoHo6v64wkWk8h3kIQQDDXcLk11v31Y5VxGDgSU6uZ
/hAyiaUm8QX8qxe97cGJnmcgDlXjqEe3vJ3ZxPdU1J3GpYeMbgCJhYr56M+7gU5tSKInVD2kxskn
1C2CcnqMIc6ggE/KnFZpvPY2F8D0kj18G0UlkWE4zo1sGhtJ3lG1oUNvlKgGdS3yQfe3KxnZyOjG
Q6Wohk5vfL3uYO9YxrLTcEPglcHHZfvOd1+Jhwvroav23itX9OFyrepbUvoYap4rpoX+dwzMmIuU
RFfV5GAkwpXyhbHjb0X+ucv09P1uFjAl93TyahQvLVpqhRkYwr7RQ9DZFiDX/04S7o03NOww25nT
IyhbxN9LkmZIuGZbDkbjNxJDQ1m0L0PKA80512Cu1IKkGL6km3iLaRgS+sAqo0SM/jhnq90puo8A
wPtN0b2EldNyHQSZNiwl+hqfZ31VMMzXRp+1rePDHdyoHQsWnPI1db/nZnt5j+2Pv0x8rgMFs73h
qSC07tOMkFVUuhZUkHKzs4hfU8/lEMhgUA0Q4h4zde6JL2cWgUuOWC4uEDK6olNO7H6hWWYMZfje
7/FLUf2fACoYq28COB5NJ2CcppxxnF0tlS7EqiA6mh2nKjZxvF9rMY1kB56npTjtJK7ANv2M+HwH
55SZM8UD9KopqNkPtF7+rglgeBC7c1zC48twQcKSmnz0Q/0411T/AEiBndD7uA9P1/6AxPYdSpsk
ZPqX6XCJso5w9D9H9YRf7dLEcPwKV1/c9dzdQDYhkjQ+duSOkPvKcXDH3X4iFmxkWzNkAQAQeJIE
XrxGSy4rTT0fVDaw97i/MyPjxvZ+4RuRd4Og0xAkL9GJ6EhT/g7DhDjOjZ5KRs5pP+VzPOR/4scJ
KfgkQBRhCszJpRoaEQ+YZKbnk72/L3R2AU4/ngkhPswW/jHOeB3Z3JKf8cTOhbpfhv482odmQnLq
ayiKlaYtRD/x+6LXlyQzRssCAjzdGWatdUATf8dYlvvMvGot0KBR+R8SpvwGpQIMf7NQT6FN1Vgo
xfOWl7lKxcoEh12S3QkN9/PDraHjWLWue9auTNAXCHytQ/Dkj/vNoQQmVv6Tf9hDJmCLq5lANIN+
HrG3Zpaexux9Rb+OgqjC2zri7H/AcFng9vOvMSWQxtDo7xdw7ks2UfbmiKvBV7ahjpLuwl4KGfCQ
DB0KVKqd+2Tn3sJT1D7VmaQIx1QXdTZ7BR8XIvSYB0tldDRAYUuc+ZYT73J7iakEg393EusTXjdx
zXUXKAcsRjtblSy2FoPUDo/Pb7oJRQUdY+Xvhflh+0wQ16uPdEaqAldKrwB2AcGYBqH0vo9kK9PS
i0WliRviS2pxcAR/6CTjgXQtgquGTYbNn/2IQPUC76vLU0v4UJMGnoXBhUPuxorm2g2cfjdNeqZj
aqlSV21ff/zmiSNuMq8qYDSxq8KyZ0OGWveDSi8zp6GyZ+gY5A+2qtqCKX3FMhZxS6TfFmyowzAm
efMKNyuWOoxae2ZTO9b36yYQcrq7IyyAafArEZfUz/TmlvJagwPgC3Q7b90RAzKC0/NbQP+yFhw8
LZGnZVqq+ObPoJ7Q/2uRhdnpYxabKN0KQUkP/ba1W+KcY8qjnC/LE3OHdDEzelwTpnipxsIl4RAB
pgqJY0wZ7DgOI1PAu+/Hagjt6Lt6oSFw8k4XYSJorncf0Q3egfu/DLDI6jelT9HTNgyILiV7bJ6P
5OmirVRSWU9Jh4is8vx2foewukm79+UlETi50xJLaHWqOaJjTntEt/1HB9xmi0CQlSAMTCKmW9HG
OsxMWYv77TsqpPn7yQFZLD4enz8fv05zgZiRmRYpaE9H5pzvrGcTylD6k9YfXCbXTCm9EsSSsS8V
0F/qc0BblC151pIT9k7Mxu5FF1fs+YynCHt6CF0alr/wQqI0mjlRSGrG95vwF3o0IcH0txYEakTE
dBts9Dtn/FG5UMR3pfBX/S9YnNTMcNPV0CwuRkVB2tH+xvg6W4pJppMiwYvsbJyCYI6PZA325gvn
K8IgxVv5uastnaVM8tvvVCsomuIidscSlj2LC815pkR896uxpill5jb98h4AoqY7Pn2bIuDsqJhO
L3i7SzRipAsKaXruCOaroUD4qBUBkoM+lKMoWyVVZgOrd5AA4QIFjXg/p2fEGCwFB+1vJs92gtjZ
7f2azK5KQOdzwLBt11J4kAi3seSc4OtZGHw/uJKPvZ+eHVMGWqbkzUNYaq0Mjdx4GMw2SsDZmWiT
ZrfgMm+2uiA6Rb/PVWYpelIpWXMBsnerQn4uf0zZTjiHRn84Y+GfbJQk3Q/wfx6leUiWnnfA2oli
DKJ34p8GZxi9XaR34NQd7fzV2chc00XgTaYvGTzPcIxlyCiSlmTxZXvpXET4RGLjNnymu7BHoHdx
GthaZYs6l30T13Gqew+M/PRUIJu07Lc3uwiuVW5sgte0TSsGWwk93dNQN8rr0ZRoICruTTGFMtJi
A9asBKsxBXgglKAHTChJVYU8TlCJAHZ7sik2lGL4apvUhLCDZ4THzrxzKyM6OGXsoZ3mzGW6I+O9
mRzB2Y/Q1mrcT/WTef+Pel+1CenrvWRT6iX9mAe/9NbhAUFPU5GQQxKAWi/yDRD7MqXqXYO10FnN
+ulpaaFyXAEQvPjb1Asu4NoU2pYs643K/WTad1fxCuqsj0N4reOGFrC+OAjQ3pKHVpn4QQNQ52mT
59PzFjqwyve7BDRNalSIBW5e6T41mzleL2PPpCnfCuvbtmkUVMtawAtne4VZxr/bG7sdCmP0sLd0
fPiTxSjQvUdfm/hJq6xMQrCFVKTHEzbmRtk01Y2E75eJnTZL2mCTZi/Jk0FkmtGmpkWMBdXSnm3E
mi2NVgYqb573XUOOPURjzJ9gRA88xyIojwlyULjXQg5rt8+ZapW4wSM3YXaGmYNkRAZxlNocrZYa
cbgd9N+1bpfoCOZbYC/FNLeZiXcqCaqRrXLPWhfTW19qFeev48DUUWZXLv8byyiOQlT3EelI/Ok5
VwIjXvf2Nt/+QoReoIAuvlPmIqZHZwJmGdgno0yJURJuCTumB24Ic1/FOAcxpoUCHsnp1HGlzKbk
N2JQ3Kpur8/h7VD3tY5qKABvStkGiBR4GVeRD9tIYs/JzOxUYtuI9fFKEjnqh/JdkxrxrjLRLt2a
o9xLiKaz3xdwtZOdffxGsAdrTZiT65fa12fWYG55d0U55PkmEm3y/Yl/leNelBKDEsbn8vnBVyq6
f8js9i+Pq0bD4g2RZS8pgleZqYtlb65IyLdWsnAbfq477Ht5gy/NzCUAnGewLokVNXzDGMzEIIeM
93ILJzN6Ezel39qYrfggX28AdBqY1OF74BgHUl7tmvmlUx211IcMBtrXgljYx9M6JarPiMCr8EPi
XlWsJuTLLKA4fPPHcRUsjj44PHqCZKgEAVjnSMfUFSpe0TtGCIc6DNrOl4IfqZWoze8sv1Sgry52
FgpOEYv8/pobvmPc2sCfwbruSTiyVIzdUu46lwlwSFwYKqgHknfDBUKd7sN0iJug8+46ikrNZjpR
vCFiSeCJavXvfaOPzWWkJ2+aqTk2Rz0SiVS9nnDBRQ4mtCMcKMakNkpOSyoqsbhkEAgyLBeBuvRM
v0dlFxzDX0Jj82xVdgEpELQ94TW+YaiqVW+aLi3JoN9ao0knmGqW3sySkacq9y//AlpWIE+yYE08
aPOVjSNZT8zM+HOrkqKxRbTeytxTZwvkkWXr80tJ6UnOwv6eAhP9QFsW65G8o8mlO0pa/HJ6L89e
uUX6WA9oeKAdKHoOZtS3rX39wbFHogsOb1cse5uMul0yobEzuni9CFM9IWLw48tQsHUju+1mWsNm
a/v0J7qIPQel0KDpVcrzL62jsReUevYE7Q1F6v+1c+pVt62LG3LZTdFBNPdW6XKkE/RQp+DDo4As
RwL7y1p4N4ytHYKEJfh56eAquBO2xpKvKEa04Y8Fsz9/fI9WHxsgfnt9bFsfZnWmgJ1l6gdpeL+w
x4qEdWNdCSqZaU5Vfyf26UgpE8z+xTjn0Wfzl1ayaRZRMcYr9VvxbjckVPK469GNoCfRo+UdgWY0
aM/+opK31wRdNIQ1gQ/Buc8MrjS93crMo7Oz6G9brlUsUvuF+CwXJ67EbEFZbD+hKWtR79QbKe/f
Stu6BH3ALJX04Dt3+SF9n2Ba+x4ykP3zBNDlp8amsCDEIqtUs99Ute+iYs1wSgnuVmkUr2MFdhnH
NkKBNbRZonCDG9EGr1fBbEksiRbn54V1o+VOdTdO7ia1e5cG+3VdxxFi8lqqtrsX1X6DON37eo4L
Jyyne7H/INeItYGE1llqbPC8azYHSdwEx/fGkbCNdZf8Vuzvm50MTGMuwUtEBOtFo+TYH3XmDrC2
JKjit72//PNoRxzrnpc0y2WOUgM/ZRMROR+zWMkLqYxbyCJ6+IEiEZHgOs/MetlkaQpg0hSs3rGw
dfZvBeYoBJJHgoM5UpQF5hAWbp62pH9U8R1sFeEHSfSuUoF+URI3N5VYbjYzxbU+ZLHc0RXAOSDl
kS1bzxJXxEPRiNSil3gtGpRdcIz+6MrWnS+Nq2tvJsB7Okj57pJ1AkLqLlQcA/lL8JxVDS+cIUJa
xF8G6Tl0lGMsYJ6bJlL3UYWzDrU+Azkpk/Ugpd4ALPmVE6H2ORe3yOCK9Nt5oEcM3z7oL1hy5E/D
vflGjj1tLg8hxADqZhVHpAvIU+kC/Vgiq8fDPk53eS0u8Nrbp4EWykCTuXKXCjn2hOrjeNps5a2y
S47XeTHL8aYqQRUxK43Tzdr7GBQu7nWkkQ6QG5deiCEf/RiIyyZGyFXIgLbc2By8bLXVkNYQei2w
CcBOCOcA3ekomAphp3wypWjPei0Ou/pQP7UJeHEhHPmY2huP/QM0WLENwBc0VDv+zMYtGw0FfH7W
elvDrj7Ih8GlFZvfb1BGeq9FoAR4udJnFURaulHWCreiNFSHYep2tK01zjRZsQUNX/bnVGgtfHLK
YHE73ZHGL/TZfLEZTa+0ZDDY1kCQ3WMhcvcoTynJ4eGiMx16OpVQ0sCyGPH+4s2Fe/29M/vZcw3I
sUk1oZCmBjXhblehDWl7wAn+IQ6xgxXbMbT2PMUZFBTqqLua1ToJ3zIWwiL2FEXbhqQyonS5bxPS
fcETUI1eGLe97npObm2Kl3httZ8cn+mllTKulce+zLnLON/aEI9At0jiQq7RZmeszLX+R28TgHAn
0GbLwCfFPuDbbP/OZlXNO4/iQh7kvSCzQtjVrtZIY0XpW8u8PlRrH9wY14/qCi3yvw2UYmXIfi99
Y9M6FJPzfLE9OCtZRjVlxAvSlGT+dICY4lAH26+s0p3DG2L2E0SB+VQYuZdyfxXB+jO5ADzWcTyR
CW5NgAMRlnfb5PeHhhGSrb6VwqqpOPGIZTMdpiNe113/Sv5h6r3dFPrJt9pdM9EYucufnMRXBHXP
pS1wR1UNckL5g5SHIbRD9ZW8v53BtyYMjhL/yNz9+4CtmhtU91bZHQpR9P0qmRQjoNKFg/JNwc2V
AEeYr9imcNEiKJXYwxv+1NHXmQlzwA/fyqiFVmmE55r6p6JLl+Y9smOuRezr0axl+TooleDfAAQd
XAiMInpHxy0gzWM07K+NXsHYrC4z7iRX64VUc9OYfLcu4b0VONi/8U7HN70fnF8XP77eBbVA58oI
NCZJME24ntwiUH16gELdO5TEqidKVCpNIYqTTNoKNogFP6vj6TwbrBZPqt0pbmpXm9mxTBYpfGI2
ziuIiQJeD2Ky2mzVXzhtz5gk5qJMSruF1pw8AnuWZ/Gzgk1/8Oag6NAkUsY6SYhFyt+BHeAVzv1C
mxyWzOHV1vtDdwEIJxeFJto2u/Td6pDFXOSj/TKk5K+XsCB/tW+fPwN8lO4dW3yfYYmN+PlScXAs
MPxDlZ6CYC0S4UkyXrOheqkmqCx90niWkXIvXxOk0bls25BQ9mO8R2l4GOhD/fqcZqv9La6gNhS1
8Q+DhxuvMLw9nL24QIczxU6D1Ut7Iyp0VA1wWKbWifDiJXtBBl42Fbib6/5bz2fbcjj83DmSJPTG
d8UKwGg5APPyNROWFWPUhchOxyOR3lBhiKBpct1CNm/8r0/6Lq1RAzN5w0CDMsr8IcUB1TboiE5a
vtk4u3vUf+hnOf5/Z9jFMLvCh4jmE7nIMPI5OTjgWESp47I4uti4nryUeGEuqXpOnXS4FQvXZC59
22BA8QgFO3tEMlCeim/g1eiMsfHcVc4JoSRUOSxlQHDbjcOZ0ss4ALVzJ2RYzrTuKcocKppUqvC8
vP+0phGXhyXZSPjMRfrt76hoauy4BWRnR3tSqKRdOE8afJeOMChz8zV3CUaj7ZCGYFv5Lt/Q00uJ
fgfzd89G9C1AxONPMtISksij3jl/KLJHFB358KGLpuULBc2Q9R38PJrhrfEy6qfIB8g8HzxGKhNt
2scWSPPbB2F+Zd58G+3KWY3sIonsxF8mrInO+R2jMc4TJ68UKlmepskH8J1mEWjpsX3CsOnDowt6
NB+REIfugAWRBZwySbxj/XjyJbGYa+fj00kaNf6r0+ZyPRCkgTnGlNKEmSf2oQYapKr6olgwxg8R
7hdECAEzHECymOHSZ8FBo6yZon/M04esb0ehZcSpzOzZQQ3JtuN9g8uNaohhoEk1pePrn0wFP+/4
/W2NsUn63qjMIy+K4rsRWHvfvc7PC2ewEk8vpxlD3ouE8Gw9+gGfsN8AGuceV0iJDmSya45f1kzJ
CZtYuV+GqhH4Fv7I5HpM+fu8sNIiY2bLgoAQO10sA8tOF4e1aKREDcZAyqmU655/S+cmkdYqNMVV
A/ZcM+wgPEA9oYGsGD3VXZIuU7d+Nb57rI3ocVjgAaB+5mBJdrF79x8jrVxcBoTLE1R2KthISA6g
xCIpid12FHZYXP22xUDUnpEPskshUFyEjJPnS24m/BtJRaYa7vMTR8Fu8lJWalNYKv06mV6bmxxg
cziyKywKKQu1wHOfQ7ujg+ETtjAD/wGU+9b9+KbNJy29CrtgFQ0SqcUynagIt30blKdDax43ntvL
+AHELk+NRtOruYDQ7NxjMpGyq3vndfKvdnJpJsMq/p1aVqL2QaAcSZ4wXrn7pdbXr4lCRwn92HH7
J7bktncCNW3WXEIHr6GILHZu4G68AZ6tjL5hKTikewe36aWeUfbRxEtKzH+VWMKQk3/wdqu1e1lr
YdFeWnaTfZ7eYlzA/ILcwbAdRGVUL2W1wWl53psjC09vTIy3A5eBL40YDwxuuVA4IkIoZUeYl/wE
0RntVduCCBJg02SvdLhzxgPbwD39duGlOs675AsGu46pmfOP8vhRTpfAc3rAkztwA3C3SUVnSvmG
22igunAWHBKHS7fBBuJzDVTf04ye33qPiC8L2VUV7ppWK0y//qWIEb1Ew8sTsoDBtFT3RQwijiyV
frPCG6RVMbJJLy87jAVtCdnw//MdGroticmvBNw01QF0Mk5aUQ6nATaF1o/Y+7ot2CQte2iqnNuF
uiOesCJ0+3SV890lDa4Q/tjky9ssZ/1YqK9zkWL+WRSAFmbw1Zs1zGxZJFhLrbdmqbShqh6MYh+f
E/OqU235aFKXb9uOUllFqmK3I+sv8NCM54I4W/rVD5ddHYQn9WVeqhs7lz4H+s0Vpb2XZJooNEWM
OpRjQtiR1NYpIUxisGT3CB1KCijngWXhfgXrr3s9xFrQVElDEGah2y13xrJvRXRoyHf4jhI4ztnT
VNkvYIy7OwqtCtZdIggdT1EP6Ytkx1dw9S9I3siMX88Ty6WTffyi3nzmXscajtTvVzeTl2WJicgY
edPYlKV8DcrHpVgQuDrb+Xb+Gxp4f9fSRjrhqTjV8E+dEX7Pp9cu/1YeGKn34PZwg1EorZfLFm7Z
MjljU73wr9V666n+WJAdpa+Tyxb+srJzvOdS2iRQVXpyTEMosU1/gU/F4eETELODh6cMRq5mBFlB
hloQE+uppGOLrBkdb2QB2ZJXr2O5VMi01s1987UyMSFvIey5GraHvXFon+hd8ismkEnNKvd0DcpY
Dw7N28AbAAJaZUVEfqwGW+/WqBW4GhUK/Vc1NJeiBOPMiG3vhrM5NDkNtkMovvY1LQr+U2HJc10h
QYitqtjmhD9DnK9JgPmwKGvO2HwD38q6yefCRsTaGIsOt614A+AMb5b+A8BHeCatJlmX3+4pXD9u
pg2YnBP/Qt2v/B6sRWKmVAmkAiqXGnUX+dyJG/fqPbE6vib/jw+5vHBdUtc29pPUbykJ7keWVjwV
mvnWVHXfAoNrPN0VuJ7yssIMVzkVXdfv58bnmdcnRrAwHJixxfTQgpQ9U+1u76hhKbFDXrE8IYAr
0r1/0rvVEyhk3VDdr89kwnGTF9FIIIZIgSgZHuC1hr8KtAC/ft1QZhWdub/bDfiqDd/NFnZPGR7g
2M1bcZyGxmWL2Dp7ZJBok6wpEGyvg7kP3GMF88eM1AoyTIfh8lTIaMMKS0iivIJGe+vhsaN7mzNa
FpRcKM2xa4KFdB0w4g1DfAFtQ69UKhAEGA2pCwCanRWBGFG0mLfAkgKQg9spt2T/EyAVgSZIxGRY
J5P6VZZT2Hoa0yDqFOKgPXl3GOVjj8Z/9t5laQVElZLu235tMfOPoxsKbLqmNxZWWzRnY6b6r5he
OYrgft82Kd6ohcIQrpsFJ1D2kmSg87kvBCzcxBi+NH1QBzR3U/em8l5uWDiDNO389JYNxAkZnOCK
mInTf08RjEmwaLVeskjWYhGqQGJaxTBf548aXYhiEyx06XlQfaBeRQoOjl59Yx8g6gdZNNgxpiag
9tRv/XlTlVEaZxlCE5p3GoL7gHC3O1kAssnniK6OizfaOlvAXx8w4jvSu4ptqSnKKhHsJlNZcH/P
mcbpd3o3aTjNx+LoRrY0gsPTXjEq8J1Rt3BWYOhwq3wedFbM32jptR2DpR0X+1bjfyhhctQkyoo9
L6NWoPCWSpcHim08BoTMEYIb0gAOgqnnWJOImKprlxJIyuANkkn3RfAw+UKpMYjXZHrGcSM3P7OW
vjgrN+GwxyCBBYvCxKeJVzur8FmiymKuJYvaFKjh/OR90GqV5JrcAwub2IN4OrYhxDeSA9aay5bB
xMZ4QrUwKxNPh0kwTyy8X/N1CLffTvtI6pZ2WXVrTN+NRh5KkkKzIe2NLOZ+XWQgX/t6D0Xdb0kB
72twOyCdvqKM9Ctz21qH1YLANDkz8Elbx1hz0OR2B4KEP3dc5/c3Re4yHuQ754R83Qo2WqkOBwRj
phgZAH7rjzJhHvsd0HoDXYz8XPDRMyq349kqkWfdCWcpGSBwZ5WOkyMA86ZxbfFVb36KSrdKWXQd
XydOwCDB22wkzHMzRp8+QAMpzWL04rB+Cp9iRUX/V+F4ZF25UXeVTrqrAhyfXxecBjqIfCRjFfyK
9pFhc8TR68gZp9L4F9Lrk9RGnSpsPgAWfCzFinyIIM94RrNG9gGkAx4wqSg6+zHSI1l9pvqEQVgd
uZrR9ia1ddYPflbQIZHRJ2D4zEqNT43/pqTlOgS/hnNhWTeM54BV3JUD2UzhVWc2v4xreMxUr7Mp
gO8whno1VegMgJDAli55uZOil8b1f8sqMKDiM7oT+d34QBYRdcSzS5oZHNS6N4KAQo2zL+UPNojF
lnhvVI3LHfgXkVg3EBhOGOZ3kELIAP9w/r3HDxn9lP6ZNrM2W63ZDxV/FcM61V8r3sFz61Lf01xB
yrGuer9vf3qnqQOUhxt4L7aEjoutKi5qBAyAw7H+MOwgeNnKWsmHRlfvVQNJbsNvrJ13imgeQ5U1
dL067i0DrQPDA8vLyWoLt8oe5q3dnLrI6QViJyI3q8M1gM+rIDSw2C6r4+XxqpNkCLXu7UZZWk6A
TU8NYtrCqwNZqL3t0rFmp/XDgwQYbqvusXJOZGG8+BbRXf/nikDvoIbUYgVRzpd5ZUPvGyeHB5Zf
Kux3TTRP/SrOHdjOeQPFFU5KgpjXsp5rC6ysYIFzGg5dHL3M9vR+6zZf18iksj2pa5w4ClW6Pjkc
zfrQIoJROOVo4+2fGF+5Vd239FBtCvnHfoTy2ulWC74E0O44e9AQRBYErIsSnncfEsmF4UYvi+sH
Nmq+tUhBrSNUKZlo3/mklK6840LSMd7fCEiE8SskTuxRE/AGTQ+9y1Emh9tKGdFj+Qi0/9A29CCR
UorxHBOsb8aICnyy+DpFOf+uJP9LZfN2WpHnjj45DEWDWD6cVhEaG9v8rCt3SVeWQ9OdLfcEC/pa
QhWTmIiEso3+PGRyS9ec6HDlwMA4eLVJDmsnzhAIUxcThMbC9q8cW8cX+D38cxnNoi7eTnXVn79d
d6/zD2+I/FLean3qKJq1j9oGC9IPRSchkL7XH8/V1fk+ph7FYrQ7WtCiySOrbK/lvw1rL/R2asLF
WrWIz9J9y+aeGWsyJ2i3Lux1ejBOe07pPfqL2Yr9/VgvxhdDVtPuj/Vmp+PBQ9QluT6FagKL9ZQB
MxiGNAUuq/nU/cUy2TKr0NBzs/jH1K3QXW25QXT5ZyY1P6234GeUq1z9DOMhsQ+lJfeaqOgYmeqi
BCX/3AMHsAokTmcOpPlpzEWFRsq1NY4yoP7yGrY1v0euoSoF6ufEj/inyaBeNlx78Hk3z8xV1KjB
MoMc+aEw7LYd4Hoy+IAZ6BsyIPLquQWDVpbELc13VV1LdqcOeG0Qr2Eu+7Q4y2I4e1uG3BJ1Z1TB
kwikqOEMvtsQtjpEmS00fF7XauMqd8V7dQi5m1azchGbKa9HWTR2mXKyzxuG0l9kjTP0CDVxILCE
uKdvN6gQm3JvXiXjD+lQ6aTZlA6qSuICU11uT/0C18droxt0Sk4hX9aqZjgxrMbm85YEGvd2lB4K
dKzQlnipgIQBG0olDossM7DNFLoWNrnwnZffBeihGDvEoW7ecSXtQc+MLeV6+yrpSLuDUYXgZf5D
vK+d5Cl1ujj2xrPYXfP3/0TNSxPOLjaNH3FTh+dLP+UtUDOa274UFR/9EZSQ2N+BQFIJD6hQAPGi
edQvK7Kgc/99OnkPAvLVOCe3qlig7gpsxoC9wOEbeqXRbl2b4eNNvborzgl5wBcm1R2Bu7xd2cwc
QZjWn2hrLZEpzglZsJjpjC9UqID8XzPspumBnHoA7mgi9HVWEVu277n7CaWb3FAlsXTcmepUJ2Rn
YXcHbHpiahBo8O+YOsVNuVhUNAV3g6CQTAu4dkWKk567sDDd4Uc7bwXJPnEia0rJ5XQaep1XSQhO
ZqKOlBVMVKNzRi/1HoAm4H+mKcagNVuw7H33qgwvE2IetJeVknFyEaRnPNCEsEg7lGg42fB6d9ji
OC8fjzY4nV+F1OQ8pLrgg3bNWs+R/92FF5kXShxOOR/chuzWiqoJQgqWOTruNrnyrc2FOh6u205A
qWX71PzTm6JXJ1y9vcq8HXUvD1aTVpzevIdbc6Zdc1JiVCq8bweJ/6ui/s9xS45aS7ZFsaTbAEPo
aDxm0ovxJNGPYeWvPYyaU+8bknmi6iAUzzzn3BjAFzYNpWqv/4zBI0Fo6cu/zyTtCqoahcFQpU6N
4x8X2Vz9b9PQF7X3m1Z99fsWGgtWt3K28GW5Nh9aRYcKjLcLJ5n2r4DsBKmqa4sadDW2N76uDb1R
iNDpLAwLMDaafBS2dHHf/Pal/Q9cizKoXUP5XXXdMQsFMMhArl68fqy4rMrP9rSzc21qS5x2mCob
Ftd8+wgjECn/1C66FZxtALk5bYh0rQVzD4uZne6zQJhDWtSvZhUa8rtuBXfpxM/pJYBkmFIDzFpb
S632QaQKn4DacFpEugY4PREHHy+O7ahPJkdivjfSQcgEiTMrdCT1E+Hc8EEgbBjjydnFRpLZBHkE
IS+VrcM2MUrH5DLwEh7m827lwt+5hkuoxhvWvwA9rIppMm2tq9Re90QvsYhCgpPLiRQzwTGX8JES
18ykidIcMqweWQD2VgTEEp7Un57zcnCvS1Ochng9tjRHXqese5UvQzjb6fmCj8piXVEoeobhwP+X
unC274cy+yA5pgP4bxlA2G7lT/KcR99BplPYl0Aumfk2v+gZzbXRwvyQlwUZf5oHGtbbvKvPkZtJ
XEdpjsz5wAyaf4L5a8Oteat21tjYByY+5O9hrD+l1sgXLvaHkg9vv+Th6A/OhOOJ4VqU53VXCTze
/pGWV6zuazaDKYwI+xAGiMMkRSgiA5nk5fH8leUzUTrNR3Zj7xfpXhDWPEnUlw80paZdS55cmvEA
HmcogjnG0E5wd4xXcGaIFG1HfxlJgut1ciTtQLi/YaYvS83YfF6c96yGhcEGwLXbRhEUJEB1ANCJ
/U2AoPawJ2aDiyWLdD9ZxB0CXX8bZ+66eL/mdcVotDyaE19nzhcmLRxI8RI8WclkjFxbrhvdceXF
/FwCOric3FybFFz3rquT435S4wmoqM+ilfxEwXfNFKycQP6Cc9RlqsYEdSXEku99FV+JxhKKXIXM
yDr+Tt/gmjlSThlFs76UgOjwukpPMb+xDJwJnqXwoxVQCXG95SXCcfG6zmlkXOmE5zZRvT+DWXxw
0nml5SM//20TJLJz22uxfEJbQ74IZ6K/f1zz7Odq1qKFQ2fdVkge6m5x6NiU52dgZG2e7NKNc13r
4ai3NzybtdM2CbUd86L24CozSjIzVmegYOwENT50Ug1MT02RbfgWMDVRS+fSMMx/qDlPUPP8sYqj
hnuBXfBNVMwIgThJtmi8zELKG5XmuQNtpJAVF41OSlVwl6eyL6VJOAcj+eyTJMRUfXElBH6k1BXl
7E7mPQQYFjFha3DgXNLViG7GAsJzEXQ+OSMJFkwd/ilPK78/dWw38MVhSMbFw1jNzG5cIZ2PZvNB
i9kl5KLgor6gfUrt2SZUkLCMF+vcJN++Abj85g9kgbn+DKCQr8bC+oJnmPdVrAOdhUD0ARHYdXG9
B1Zg7nwrjCj2pj18fgXozJGV9p4ftsnmA1rAsUb3h9hGyxzhTR2IC+Res2fPvNb4OQEMnGjh+Ujw
p+w8qDxMblbP1DecqFG+H/DmyCJqW34DJEKkyZwREfvMCjMz/ikiKpUYQIec745N+4IvS77jqHPt
Uypt+Tpk0KC3XtPqtXrSi4oACrw2cxLmU3Ua3gn24LYUHi20AosGZckgkc/aXJFXTZ40TsICS1QM
d/JrmaQJ71PeYTxkpzPSNggLgb8Yu1Xb30+dXsdqtNTJJ5MmnJj3oPTn8ManPbA6qLfroaVkfTjv
lL7KA80ml4mnKnDFJrt1NoAYG2mOiehJIhO3sZ82gT75Of7J0fhp/MD9BNh1CuxuO+Vg3oClSUZB
wD1e4ElwCVy0BNVB2K/yChTRCw7PlIvlMI7ZejCxVf9eCQGAf6pRiAUwS2u5AkzTqCVquZodRnU1
OVbBXFnXhlzk7rbVwk5KxiNQTZY3C22uS8Weg3R2YMSin3YIU1g5hF1Daf8FOEk8Cl0NxhL8XyR1
AxkUWcBmTzjIJHIBIqmSQZEY1bpDFSlFZZax0T8IjhJb6WlRyVcy8EmHcRkmCjalWYCw9rfzER8U
H9SceJuiX6ywA9BekbxXjjd++9psZ1GLA49GzlcD7v2qcvghlAFAPjNhopRtGdYj2P6A78I83mJi
6l9e7W4vc0rpDge/+JYCWMcqD5EwhgBMecxkvA2T8jK5kqrBo+95VS2v138F548/0+76JjlSIhAo
k/s8IyXGCvzmBY6mY3IvecCTV5A+bdiM6Jq8dN7jbCTl9qiIGPl7o7DhoVFRPe1B4AYt5Cu2W5uQ
IBKLh+yyS26dOBodW6pOwhvzo8ZrRK1MdF7VdsCvy5yDUfVPHoJzxvwo7lGJgSDwWPJzFlP30g+h
02mekPanGdjXA4I/wbIj/YiKNNcK4JAuUBXD1VTllwPeKG35HPTNjVbRi0qWdJltuYWPFDt2REIz
8h0WVieWcTebjNwXYdhBQshDpemI4jvx+7DB9VC0ZXgugSCcqvMH9gjv8MsU4N6N+e3tSwSwTsKY
qWflnr6cMvFp4VIAu8RFKLzYJM6mi+3EU6r/0QSQgO3np9FsOb9Km7go+YSy8QMmul8RyZWgr/r4
Hd5NH/CCU4MXVsgnazlipOGF2j5c3GmCXf0lNjIlO8NVCFmE2W8VDKSF7xr5N1ZhXov6qZPajW65
fq+Q3B8IO/yLwojbu2VIBQmdOncf5NkZoKHBqLkjA20WmyZvZ4r4DGpBWRPRvkOk/cyPR+s2JlE+
pV6vxAf1AXfXa5AhaeUS5P+VOzSeJfHqJG3M/AkGAM9UGRxfLCcb5eFSqcBlH2eJhg/bkxh7AG1w
HMNCt2lWGr9pKSCMj3YqCLYoJoCPYrR9cV1HnWVRmPo3Uy2mXIedRsHjbgUvr1oi2dmHj2C4636L
6joVlIfY9VI+DHtQPkoUn6Oi4geClm061Znvb53zRmm/mNXpfwGr4e7PG/tT8RCWGQvIpwx1Mp5z
HnhnDeUCjUieY4gW3TBuRLhm4AX/MKrZzL9KAJQU+4EV3MKoYNDOkjRAcD0mzvgbSOAZm0csJLP/
7Ip27CAeC445F+h7wyqbuw4wXz5U5tv1IaOShOmZWjBEE3hmHGcVuq4eb+ZQ4lHwD9vOjfeZZjAJ
ww+iq31yf0AR2NI9rJCQFXpr13p0Pp3cHqGSz3l89yFYONedutV65t6wwDDs4/iO4oiuI1EG91fA
LBOTSe1oB49NUb8BdaSAsElXe5VGdnOfs08z7uqXUYShKOwrkBypbU+vWbNED8yLbe48jEtJfFRL
avvyVDpTxQNefCW2KGNFcSCGaIQzbh27H1H2hiN6Txyy6GxsY5niiv5Xvq2tdRXs2jWe9N8bYSbG
ov+iVt9u/zF1qLKhIEUXkjoR4Do45oHQfQ2i5f1mYLQ4K90LwhkdxLXdWCO8UnHEuzSaOv0+WNmO
vciQ2ish6Wtd22WEwvZpbpVf2HJMdSUgZB9bg9sal/03MmbZJajT4Sl+bMXHO7eeRj/3a1I1OeKX
zVZoF8jeCa075fBqTwXHc/TE4DYIQiRxikezd5o+0riU9RoT/Yl60d6T/UU7TLkLCUyG91JZfZEW
vGLGW7+A+wPMInXKMiX8xsBI5JTwFJIsjjF7uq0Q5n5Z6aplvbEs4YAcddtDz6Wh1v+CPgFZ6pqT
vCF8txjFr7T6OExQRHf/1qK3w/NXUjBb8oOBXH+cxocHZA+JgwxweRi+Jcf5EpDm+HDMdfMT4VAE
ePKdvWChsNJPHUSjTKSF/kd8QrRrDB8nuOhs4Sb28yAZGOtcSJCNonU7spKfjrTw7mqNCGkAFUKM
IjqFuTOhSo5aU/+Ey/4KPqYoigZyzyUco6Ewn295GD1EAOKYyzve+N7UQ/f1mkEDuE+QipQdCVPV
MzT+R11BMsNaV/81/sc/FgEm8z77DA6y94C1eurqrTWZaD3KIGkRQ1A0HsYngtTVCbINvInheR/B
qpF1P08jzXnjtMx7v5eMJR/iW5TzbIHb+h/LdegvyEJ+4sCuGUFkOOAKcI4wnpK3WsJdWpjp/Q2x
yizdaEeQ4bZ4k9cdXcv12wlgEirCJ/ipEoOK9HZD2hhKcRh4w+idZelfwfWJzHzy8ppDefIk0dmP
iAOjq197FqcSKeuU8Y2x4eKio4PS9cdAmDLk1KpAE2s7o9hFenMRSfXp4hOx8b9xK4TbK17iMHqU
+ESr7GiLt2eXog1h2u8iYNFPxgcHHfLwoGnXnWPCyWCrwJe27vXuf0btT7amFhAj6O2ry+C1xJXQ
iAzOueYe7u0TjKyliFk4nfkvgufUO8R9syKO7hgIeVYmf1mGzaMe0+hLLCykF/cHnWF5MRSSECJ3
iiHf5K2e7+jyVKIjDYudW6tsEJ42HsX/sIDbo2MhTLxqEy/C9L1qz8Wv9VbXcZr9ZTAhwdBR3IqI
X3I53HtPyHx0OOOaWK2llrR6Mfpr5CLwhGuVqx41XsHlCDPEui8pVTr3i3eKEJ1FF/PLvDPj2ch5
U+amb3yuI3M3T9EFXX8QzjERw3qqrxCLzSte9wsthdwfmoy/+nMDug7xxinKa9yWWToW5GT4fjs4
TSGdNK6jGp/bxzSF7J3vbQof4eRvivWwkxUWW+gSsnwFOHQhGRX+KqwCsg4Un9iHN47j/LaWusIV
4ijExaQ4+rXPO882ttTIPqVW5MP7fGdEozYLtiNn4/gcGhRd2ZeeLQYe+CyZfh4WjLR7+fylCZr0
OQeYTeMJK2NMBPpwE6IggPEUiL/SMQZmQqKbGHNf6C1wAO8xfHO4KvaDm6Pe0FmO0T8Ia2mGIkPj
wR6lxksOsBOR1+Kd07eV2+zV13/VU4ooJp+nGs4iDYP2pLlDvDzbBVeD9F8YVJSCznwwUwSlgVkd
35V4AxvPPUdkOypIXFlT8khd8KQ8Be04HQVrzj2L0LmSKhrpCcS5TcFGZkbpw/QLCVkDH+86Wd2A
y2xwYzaVRdIvogciLkFGi/EuiM/ljRyytzhyelOtxF13DHiXFOSdkq3mo4Fv2WA2jYWBl6Fl3rPe
BvRpn9lfLXzIgo48vcio78PFjhx5kEpm87G3aBdwtL3Y5y6fHevZ0sAzTeuWrNFC553MuMzSoqJm
dgR2mBWRQEP3689fwgFUaodSLv3ih+BGTd4SxO1YweOtKqmNGdfo5+QXUMdwZZDBR5zy81M3+oFf
7C3VzfOGILGhtrGmOH1+wo6rBjLiMgmUoDLfbh6Ll8eYbxBY/kY3pagA2DldklADNaoN12OFh08Q
Bx5P/hLvyy2tTX90Q5NibtVb794ZlxIAHZPqeonF+5AtfzmfEvFnBpnaKlMmaWBQUFnH3o6B1bxv
Q8OawAlCsSKG24EZsJ5sil1S0Xb0yAmbHRwGeU5KIRISWWVxsLFt5Iw5xA3RfnFWhcQ6QhpehmeE
fGDuP+NBTMXMMrxjmRvxWxmVcMtMl08jm86hWKcbWwrPGKJiWnj+fgSTQz0IBVFsU7K5PQDBTRso
efaK1VIMSs0QLLKE9wvxu8hszQSnhgzKi4iBLmianB0QsCY19CjpNwPwjDOIc45JYpUsSi+tm0DR
nq0FxWwXWEHnNSpgLO2P27O3+5ugraXvZkOyOSPqG+ngPSYDllQOJ0mwrOHBSbYern0QlyYB1XOw
f4VZXHGWZZCJezrbWUzDH/RkTSQJgcM7/mIf4Uukj0aIYMHhtp1/vdWHi7kqH5CZiCU86NN+OSHC
W/Qxkh90D+jMItHjLeH5mdmX8J2sy6ufSOIBfiAuIEveNJPzEbX5eRKlkumlnKI7oYuPthPwzzvZ
Nub2kUWs4oWdr12gesC3igF3ai/KEPG0yXluMTcWe6nXIZV6PGBa8BCkRtQI85eixlCLbCgWh4Se
R3Ef4zm9J0CT4q082u+IuOi7w7t20Rznr0p65FLWHstAKNKGoQ5IALMAzYHj83w7eS38FTdNjN9X
X1PSgCRwXZSHbquiwRboAeQJJilhhauWZ2rVZ71BiuFFB8VSImfkNL86AfJaO3VtTHGh6aXYsdx5
bTU9EJqV9eOmfn/2dNQHBAzNm0aUR3En6RzFBGoOC4qvWq2RT5FyVyJJKFP9lHl68rKXEUdcLVC5
kQhoKI9CT4xSoW72rD/DBk2lJPRHxDZ5Reuyes8Y33Y21FpP2EGdeT7G0a8YEDcnKlKnvPD4RKAm
p7iMx0EuoFEjDjCygzQVQ9phLxCA286s8BpFlxlwzAVuiYQLsVb6xdUpzbRHziUTp5sl+hvFRa6x
WPrUTQYCIUzGhADIgT49biJWsfJ1bi1ZQcW6U0PGOKy1ruhNazpCw3LK3O3kCiB6XPylluTbv+v8
B9HSXlgFWVpz/kJgcFEq2jEzEfdC+goo50SaI927Hpz/kd77ZCZQmmn2AXSQDYCiJQtogy5eIFSp
4jshTewsKyMuuBAnSQwk3jCXj0N/lzsyI4+VLM1ZNVBWgF9bF/5z/aD/l7AFJlB7PqGSFarV3dj3
ThsSHx37cO4VjKpwDYANYeLiZoLJsZhK8f6T7KORRqPeXmQD0h03rLHbieZwsyla8EPm79iUkMJu
x3weKN22nINd41fnRa1ay59Nk/gHcKUAVaMxUeyX/PEkNvY3CcapbluMfhMv3XnAm4ynnEdW5zVb
toKJyajjEZPc0p6PamgI8ph9aePNjf+gkCKkkn+hfHNJ4VK/9f5DyWdvF47A2l1n29+9ANMs+vax
clFDxtbfO+3L5bySSg6s3KXcROwr2DZagYlyC7qfigZFAExy/m/zCJmGgq71dT18CdhProcqojBx
BDwBmTQLuQHXjfGU5Ety1u3kxBeYi1XYNJGUCYt+TJqi9is3HUDUQEB3eWrbQS6Jbcqt7Rwy1bvi
ZFaC2M7UQfQ+toRB3V4ck56T4HjmP2MVLZ1KlQdWV2LbcBoq2oeQsF7xfHNFeJL3P23RB9KLeFK8
aZS3WRZDtsJQOubwsjqWEMV2nAHGtCLSWhXgfAyDg07vP88ZsfxIkw281bhYuTQnrxcyy6az+ITv
z+lPuwxEa+aHTC7imHaPURdbG2BKlWiakXCqM4RqXDN2WmQFiiWJj51zS540qVCy0O+2eNuTrB6R
nP7RihBFEptx3sHAi5x734ZJNXDL5Z1/oTZCBiZ3ZgOfKiGd6BtpnOzsgR0Q428pRnLO+935Xlvj
ZNF4ze0h6yOP6Axqncd/O7I2zWW27ywtYNkBO5VhZ9NNiR7cvagmisWh3G+jaGWVFTaF+m/rHsZ1
8t++ClWYo08D+Addxzr4HSWQyonzLX/skbA/1QrkZUYMG/ZhusGKnQvo5onx/1kH6Dqlmrt0A/dK
vrLLpAULxaKIUneersiBP8lppeFiiR89m4iiBS7deK5AldtkNJf5OdOV747dvP/iWh5oTm0dPh2e
CyIXQu351tB+RipNJhTK6JMLrAh8iF4t1glv+f3s2NJr9oO8m/HWZ666Dnb2NH/xzFMYb/TgB9V5
bZg4f42Va0XIKTg4V1e8tR7qyirfV/HlHWQoqYtR7oKOUK0yEaCYfXTxcvcFJnd3nJNXiXy2XqLK
y7F638J5lY5POK710YLTck7h+FmvrpA5c5CacH7JYrpIi7qWSmS3yaWOBaomBYXiaXGLW+ESBko9
nIxTqs7Nr6UCdj+ZvQVdmXzwwIhJXFvf8VSWavjmq2Sb6lU97TN2ntZiEOuj97oIbnqg9eewsCfy
Ju6l/Ae3mzWjzcW3Pq9T7Sj8CstuLGYrcv1KulveZSlMGne6cZtQuDFniwLs0F4eUI5m3TSyC1AL
eYQ1JZPtmm+D/aAhqzQtxC4kykJiZ2SfaGaGLB2O2+2mOP9TGEHYtbLbESziS/kBpmEZjXW24kbo
2q+BDHbGXP33iLycWyYrLrFJ710KUS+2huKYt3RC5YgWAAttQZawTIJzwQ0LtOYH9a2Lqg0jynH6
8AOe6HtaHUj125kpo7ChOXeCwvksO8CBU0cohbbU9hKmZQFWYqn4MgDoIs/9208bPkq9o75yt6PD
gFlkaW5hbGns583QYTYSGMwjZuV5XVIfvbHFWW8y9KoqAjoH+kIxq3CBdMFx0sxVp76qfygVIgwA
MtTXe4pZO6nO8TpftJPBX1VL9ZVzPtrGezK1ptHjnTSlTg3WhIt0Lx9YMZM3lvpAwthQCP0Xz1Q8
em2lN+p0GGuJBIZ1PGNtzF4s2/ewfxuzYxNyn7gXOsxmQKfrwalK8iHkjXKUCtF3KLE0wRYFFgSw
bk28vqIco7Jw57IxamENZf7ZLKNG605+/fqT7o8oQv33ntnYVuazs+wl5y2dTcV4vYJD7qStHVvs
XHw89j2eGTbSoQ+uzYfORprS1bHAHtTDSAzWmwRgEPPpcjdHW/0XMLFcnc6Y4J7gPsJyl9ML5uYw
+bv5I6/2rPfJF4a/DLdouvZJJ1DhDZ7UfKNQCX6LtdbshI3D0zT0jucOxvz0hxnGieQz66nfuhBy
kZGZ5hb28zWI0aKxBmBgs/0vMIS6n27d2rTHxAQgsh3nbyFbzMFz46OshBex6JLKE0Yploj4oBSt
Jh6dwouXkF6P97AirEnKqcQUOUrGZaph5jOMAZ+GpminO6ci+az2cG+v/z3SCA0ib8+cR03Z6c20
gCsYZp0lbnAnU+oC7Zo5aMZjmm0n9I2r9QnV4fBkJruwrLhIW63aYjGHfgm2nRsltbEa42ojWSOY
uiMQsAQF/tpCyH8JWsJCQVHJ/C3PWKARcFC0gLk4wiN7AHaTWrbd8fb8bKkOcDVLFxzYnuS67t+9
3PrLvEgz+7cHXWgonr7jUymRBsAROUr4ITd3i5LkDSkob7may1DSvkWBf8Q8TB29KZIo2oOeqEl3
L3PbsByPxr94XwVjav2CU8ndLm2PBVS4Exu/+ttjcuJicgPd1Gsx8qJzi8lkmOS9nqAbMnXxLAh0
pPe0oh+1M7X1CJn7+TeNl0tkKq3ijHi4+JFhvKqtMINKe52ZtT9/o8jsmXWfoeCVJ8USo/qtxYFU
owLIELH89+O1mOIAqxYaWuXmYwwNq6xyhCyDfFtG3QwcVsx7WP0cDWkrQYEWFybthHjiykAAU3ul
FWj5o//fwR1YojfFYIVCl1i7gu0bWCLAhhGkS4X2WmKeJzbbHguMMV/5F9ESiPuHYJ5BHOXOEMKb
Sgj3KuVCJbQqyIWzc2K8pqHo9/fakgAtgkmEsCKYfvpr39THD6ThfOm+tUxx4Nb2qd7e+oFrh1c6
grzJ9ZhG6x2fyl4KG4hfzQTHsVFDK7K2oP5/67YhTA6NZWr7yoSThb7CBo8P8KeTxRG5DyA1oDEM
DoaBG87s1hxlBAXqSPW9MsHoIH+dgHZbBSVO+PNUkUIL1+yjhmMvgeTqTfZzmMVXYrYLdDNxJf4E
EnNoy3SS2LSicpZertHXZl4E8mUvhsVZnZulH9DivFSW1oLSpQWA6cWuFbhJyOaWgbxDiSwIBuNa
vqtymgvwOilBGEcKjgu2+ZSz1F185/Md+13qKz3FPQLfaKXe8YWDYbZOZwoLor5amuVGuLrcXZdf
SnEfI2BcWnjmlWFrwEpiiJ+Yn9orMOjhOvSroiYoBEhf75hywwkbSdpLJoIniuM1xQ50vA4T9c6E
E9ompm+qZsZyrZwtjfct4vtFH94rzalhbgZ+nVNfg/b5XS7YuWAFGfTmDm+8dkm4LWLrd4TKb0Mn
tD5NQdxuS9tCuO0wmJEKOyUFOOGQ62wEaKyLSSupkBusqtknlMxC3tZdvRlnF7690HQD1s9+msHm
0wAq54fnNjEZY4tEuhmv+0rObQFDgdnnniRCutltIrDsFoHJ2OLSVujLZa92I0I+IKrR5bots5m4
x28w3FW2k1GcWidrzeGYZ6Q5bhzm4x69UbsYWU7uV8L6StPEIpQbX5Z0fNOq85ELlrd8fnhoizWr
U0SSZipPSr4S2t6rAnBFa/JlZQcsrPJgnC74H2m+NPk8CXCK6utGJwidCQzBvY+ju0XJKgjrqijz
hlUdNpAZdQyj3+7fgH+1eCu/bajgcPCZBZyiqogYZksWVkt2/bqDaC9vDiZkXkcTU8dnLqCigrsP
B033sVhCgXWX21ormFoVLQiWys9+j58GIxREzYqAtIBrn8Cy6125B4po/xWwoBsJxg+AsMe+CpWg
/Od6wwkAQEDu5SgcKqzY5uAp8KB7prGpq3ylEe7UiiB8GQsb2OwVtIJ3JYh8f6UB4C0etVV59Qql
Wzr7kgkpf7+PHbCW6r030H9YagsbiNGGQC4Gozf3DPnU9ZyzgoW0Y5CxVXw8KPK1Vkpp/kZrK85F
FB7m/atEY4hZ5kF2N3GjJ785L+VCXClnbTb9jtEOrAvYskkEaySkttoPxDi1ldyF2wWmb++nHDaO
mmwsEJBa6E7SfI3RtFyPJNBwWGcn74tGJ/MqegnL8l8CeGcmpc4kw00ExlJez6H75J1shUSPWAEm
ROZk16NG5dYBlAGUbUsdKpgx7kC74ZTQHhZyyBCbrXg5uyf4O7oFRWvFub6j8jJf/dAIIhRGdB73
6/CyY+qJXOYrFKr560rXa+r2869cufqeUKtJSWPV5ahI0WXK2fxjKlNzCDDiVG0L/wqbIhLJtux/
tq7UIqkTrcAp9Ldj8+7YA7NrABFGoAWA5az7kQtQXDENMK96jRdFZK3RsADa5vE759fJVKWQJqr+
2N/MV09fOZE47pkXq0/3Fp+FjgnIwgIuC1ZB7e5BbUhBL105mrCJw84+JXlF3uem6qx8TM3PYIWl
F6zu6QfKKY8BL+ejh4WCmcv1ypEXdJ8Ze2EnVQ42C6duxNN6zQBT59XI0FtuKw6tdR+rjvfigANq
nSAe25K1sxE5J5/moHmH32AG5YLHYCSonzEoWHORUS4i3tp3SqSde5FS0lFMisRxnITntCMrGh2J
3ds9IQkQoltKj3oJx7LvbVozPsY6g9/E5w+5n0agjnAf/SgWTIVIHNoTPSbLXuhUmB9KmLwZu7WU
TonqGk443zRP3T1mq+Q7bWdxRTQQ/IPaGiAPAM2JaFLP4wImp48OKIINjcUWR7HwgzeUtNLtvo+g
zem0wYFuNzuXQfvzgH8rMP32ltrHCZMmpOAmgOQqvQc0eTcDe+yW6z8zXWyyBIRWU25PbPFkbsxu
gylDBJPf0YJ8WUQpMTzQ3wlHS/Rb8Oa4dlpn2edSzB1wRn5DeLBhRxRZJm0gcx4ksrjmoQCXNFeQ
ifykRrKPFetYk/EeYJo+/rl7SGZFc/6QgulVg4toquqKuDGoqYEz/CCNGolr7DlkBPkoKebRBs+T
t7b4jWJeojK8oYU4LCsDFGzv3uhYX929tso07BNIBt8MvV7H18QdDQckKuPE2i4SjnMlZ1wWbliB
VajXhWXw66+GGXcblXBQGMJVrlFGKWJWsFzWeVN+JljpleR/YGWjU8MP1nyfDGwP8Cm3QakmSSt0
5akcJY/ZzgzCu5x37CbScN6Dcz6AV2jgsgk/CTFbmie03hEaT6CVuYHCA5zUjrZbU1dmiFH+bqIe
kKD6dOh2K51rXgu4ix+mB6WpdR+FRT6mvr1y6f3pv3pCCJEPRVCrt/rbAyflbQUaDUr4U1EZ/QYi
6fcdoiQWQCUDySaNZ4Vdvo/gFFd4mMMqmx4BlJKkiyz0uQ4hzqXRHzw309m7ul+ipVHf9GPd0m0Z
NW4QvqEwWeBG0FLMVC8vnL2pZo/pITtvSMKUVWNRgAt3M6eOvnua08AO9/89wQhuwG6k36h9Dt6g
6h1dzerejpJ5WGxL/iWNgfPzbOFJ5/qipt+huJV1+sg5EFiGv2aVRPrrSC9PZLc4o2zdhlFNjwFQ
vWSOWIzXqRuNlSYviQHZrMugFc0wSwZHU4In3qSa9OyWgMCPF5PxAvJor3jQ3V+YJIDo02dQWMYL
05HwkYFeWYet308M9KTDiDA8jasKE8p4mctbkxoujovdsE8npnFBxwQEdh+7GtN4XEdHDwo8qqMW
KZIllGjnxNyTz9qhu91M2xSNKv8gHrd/e9uePkP3fXUVMIpiQpcH9W1FchOHpaPdWgSQCrTmi6qI
0SH1Ma9w0/8P/kQzFOH26+Yi9IgWn7LUN6SqnGeeNhmIh2FKZm5zjkfMz6VvAYaQ0MS91ZJC4KGo
mKWIF5+2D1FO0CtNDSMtGcBrcD6vGriOwXhACoOhvfFQ9jvCmwOHn+mAcAurzgEfoxQYVmv5jSs9
c2S1PWsszWN/ub1qu16+XbemquMneN3WIWNGM1+1rYOYK0Q2x2OcpVQYntlEkxHy937HRlJLsqt/
qrVUCBZf38k5Ws9WKVIhJNJKdut/1mPJPwtL77axH6eK+iPHufJJJS5zh40jsHb0JG8iRV/EIRTC
FssSoJRjLDdIotY2EYbu3SZCkOrR2rikIGORaiyF8CtlJcirovxk3+HDJTE9qzHAwgPQplgX6xHx
nViqCqHvUg87zS1jRK2DyCXbuHemS5dKUVZunoSQKX9tq67SlrXiuDqc1LLYjjWkGZnk9qzipPjH
NrTwzRFYQyfF7z0/25rI1fS+PhQ/04IQAicUdggzzpr7MjMbh+y8FFxaCuZlOyw7vtsf4Xe9tYk3
eMopcAp/d4rR8+sTtDaljUsQWfhEOb6nG4UghvmUsxdJr9iOQQDZSnwopkB7/YOvNjHg+qtiumVS
MuikOC+GlsygdRtN57Zb0UCn1StsiVA3r9R4xgyi+5O0QsnklvSQgz/3OtRlQypFfTEOsgTQNpgt
KDdptPEAulNyBeQDdJ++CFWmm4oUEmbT4IqquUJKeqNEbANHJhXpUiKIsqpu+whEYRzVYifOQHOx
7ri7cGs3oo7AhwjjWxwiYSMZinoIAk0yY4xlCW+9cGrNI60DV3rUbT/qjg/j+Z64PY4XGDv+Ypxu
3vjZmm1BCR4L9xnoQPiTwn/BP8SatJP/zq2kkg90vOTZ14CEOpUTiPe8Q2woIxDiHOlMeo8MX52C
gc0k/yO++jNlVLELdtQi2sDXmqwUI9PJDniQSrRuwWNyFTgujOUMNGvKC4FOu3GXU7AVauWPSpRM
uPKRNfi4K3srCXvsyOlvifEW5dsNT0mBD26FQQgD9bKUBB4ev0Y6YjLyGfbxf2ePU8TAELdeVUgr
ZK0k66dma4wDwa7EHQI8TgAfi7LjvHT5w2q2Xd0MG2+7XR4bmw4R8lOjwjEI+bdJYZgHdNG5C4sV
wM2LC1CAp9pwOaxhfveOC3CE82ukYxV4VsmI+ajApp/+4T1CQV0o/R+VUS5nUpKsfkSFe2NJ1R7Q
M9/5+cLn3wt1+K+Q0kP9c4ntiYpPvm3wJdU5lGwDgx1959rpKVqB2JbUxPo+0Z6CdN22pes2aXtI
VoJVD+brpN22qeZFBxiNwNg9oze+9lbgY6Li5CAf816o683D2FySm0zVVP+xW4uBFJs4WwTxus+m
SEIfhdosd0dtZhZ+JqFxemBkoLL4ZRbXoXW7EmyFD4SaQBYcSYyiIrk9P+FZqSvYqkxJak9tKH2f
R5H6XPqvHEQRtDQZK7BQSTswvFgdrvDloX+w2zaFPsO/hPmN069ePZvcjzVAqeKXq7wgf8an6GHI
Akdp+9MUa35M2Hh0bfnBIPZ+yYVli0mZWCqb280o75RINY6IuwBPerI5FQEqYsgdFqbDgqU9Q+ID
htZBmRHQkeZjcqguj4TcHk57xCu8u6RxzoyDF2S0BjHJSKY+5q4ezh3pKALFE62F8fPUyjAigKTx
aedodESEQ1NYJwL4JGHCdwQ/RHe8bbYuQtdfd5IDpL8rIp791ldKUQQZVTkIgoPppT1DqwdGUsmj
KsBOPPKeah7d0Jl0+BnWHbJrklQRXVJtrS2kn0umwrNWE4s66GClP8/lITDeYKaOEJ7TDprl8gOD
rA8A7HeuN/O1ULsLtS+lwIjXanVbOAQwSRuRMj4ljPlbFNWmL28vDSyT0fQzltCftbOeq3aIhh/F
hAY+BN5JIEIWNyD4aQcPZBRIt/OzwHi+vRLUX3oP211x7qnXFaX2njEfATlR5CNUY/h1i+TLD45q
ciH0K1gTW5O7lI5mWEji4VMXjuFUZutVGVWTZNR6MgkjZJfMY/mTTy5DPWxAtcbOheqmwX7LJIAt
ttTSsNYt9pi7wyhDxxB3qJz29PcMarGU4HmiEZULoNFF90ZrUJdyRzyBYQBxPSXz+aK75zJ44AwB
Eo9segqIYOPXQ6rvoVpBMqmQDUXRxcn5zjgw3hUXs6SifkmVR4zxaekgmEas1OzjXuywJc/T/a2h
4D1b4r3bpPNLnUlSbfXPeDpNXpP5Wz5jZFi7OBgy4wCABwrJDMui8cHtZL4RoLeqDvUMu7yhPcBQ
r/S7FEZputTMOYAGBljcMNIgqoS8OwnEelwe+bUHH1MuUiHEmPMIHOYb77A5c+GVA1Erf4F7bMlI
91WC1S3ee3mbuFCz0+gO/gbAS809pGNNTvqEUHPbjcuqg6uPIa8W5rFvgjX3vexl+LEywfUcy1Z5
nqS/Qm2+jcjY7WARbhncTA5Mopu+UQE+K4flHfG/M8g7keS3WH5nsWaFnQ7Vs8u+XfU3U+57RvoP
M6ZVEf0Rhc3smf6xidloRASAcm/aNpjg8v+zqCgDVRIyVu+uFMYFbMxmJTTjOGl1XQbOCfR0hTcu
0yLqDH+9HRO9eGZFe1DlweO1cEWczSKhRhebMWybK+YWhNd5i5K5ei1DcpH0QjPfazmCV+YyeH8r
bZ4t8fDfSbIzqAjcP0TAcoQUZuyt9JrNZlGKcjqHFw+6+WKFp/qRs3kZ8gJAR32xTDS/NbIgNdO8
6wOeyeL7zhXOGi2YmKWk+7JzWM4is89K6HeANIIzEJ9YKWCVglbiZIYy0QVAOa82e+/aHJWGhZDP
lG8F+rgOg25kFJxOHDqfBppea5dRBLhjmwMas4ODEeuNL/BAwrGEk1mhayuZa/B8oq3PV14SVmqM
oRCQmPRfXcODwGe4uhkRmYMhZFqIvHJnqqeBMtu7jbYz07ZsZA8b/KwhBFvz6JPpr29ln+p5s3q1
/xUwE7eiX6Z02UnjQmOfU3zlUK6a44Ued0jIy55VKcUK1+dqglgJ3292GFZKIik6FN0S7xkTN1bx
0rswxbPqnwKProhO6FOHjupdAyCZRLtzgrKlLGpa/2KBRA2qtKORbvQ6JG+cM1kNWPjSzY1X6JNR
ZamznK6HCQMzdY3ayNWDVt6kwyOZ/TTjrSwFJosMtPHzbkIf0m3G7kF7ln406IGn6QW6lqGQEqdM
T2sMFOStgxrgr3/K9MObsRCasPaWRJynwkAj1a2qesXMYtxEJAmZVkx+aA6Uoveib/Oed4L5EVAZ
olN/UIXBU0VLKIA2ac9iOtQntZyljMIE+j/JmTBNQaAucWRQ0c93QT2jUo/iRv7M7HZwR7PiMJPa
tOsqcvEyWesAzjH9OlUUBsMgO0vyqB8buRlfwrF4A53gNhSaTUJfAg4eNl1PY/Uzfb2/fqXt0my6
4OPwwuVI6ZHzfudvihMJGfwfAzD411xe8/JHcuHp3ai18f6q/bml52YFJgc4J6FNBoz1a3dXXc3V
O2k6xopOjdKN0VvP3KqnkLNhVWddNX+5vjznOSnUOfCuXO6x+EoOblgmt4Uqa6VNahlC4fZ4kYPd
HtgJG1g3kguau3BT/CmlAaKGiO8GZ6oCfZeD+QYM2MhAdGCVEvNJ9DBGMO56m/RjwatScfkvyhEd
FqKBKgY67IKZnJpRt5o/t7frr9MI5vxCk7MdoeRtl5OsPFjKW1iDf1W7IMqqZ6B/BIHBdxh8QUXa
kx4HlmM6s/xKsbte6tch9Ggp7zhNcsf/yaA7TDNp0ydkuHjZa+S2JSlJaxzcBzEBTOwUr8WA6YHY
dZ3HCTO73oqk/eDuq0/WCJtdSLPi6GqnAAQrKs6IO5z1gmN311K0pGPBel7a9nMDYSAS0EgZ+zoE
+OPvkM2PZM5CIX2PvPkIiZ0SukB8d/VcnUAR3FVF9wJITeqPQw0e8K+lzYGOTeSPlwQE5/OCxppg
yy8VEnLSLTGpqKnKzM6UBZvXN0+k2ENG6g5KxyOZIXQDegBsdk2fz+DmeAdTp5V9gziiOdcg9zKI
DLuH6d2cJAjOQE2j3x/3f5uXMD37ls7ksf7rJFEv2AqE7cubCaXwKcgWtjT98tbxpudPlapPNdzi
p72P3iM40nvVddE0TpwfKCqQ+twI1IBEGttuZGJ/ULwQ/dcFWF2U/+F5tFGs6SPYDJCntRfxARll
EazKSKKCinKnib+4N3Sml5G1QijU2S92FQQcDbtY/XZtcSVHoI8X4ZhS0jc5TdvTnR7YSlIv+S8f
oj+xamW5VwjuZyZo7LLwpbBeo4mc9fQ94I4cICRIIekU5Tf4go7MymAbThH83+e8LZ5kw4qYYksG
g9P+s/IJ8wRUn4KDwt5XF1vk9q0MRMehQgkP7oeWFrwLvDGhroHWrCxrhMIzFDr5rqe0odB812lq
LEA1yH12GomSCGgpN09WXNnBlEKgf1f3WVCS061fBk33Nf9dWkcVg2JVU02JpYlCXMi5puT2uKhx
FWw79EW5ieQfcTAd/kOPBth44Hn5f0i+E1lyBehUYmLWzDRkrVBaX7LECZY6eE/K6WQ+fW1W2b2n
fZMiBxrHJdOXFiz0gN7NT23jzfRr33vQACO9CktpNKnLtx2xLjKNfPY4d/cOHE/sGpjuav7iAZoT
NfYGgtKLC2ODO3ZlJBmYUu29Y++jyhir2evmj+GGUyO091e4oTrLIpEls8Hdmas9E2GPaDT2gJfQ
dLqzZnhbB0D+HZGBJeTQteapMmsT5NzOY+P4w3jX+bSKZMzJ5AaCat4d+jzJWfEWNpTU3vgHH/IB
biXj5NuPqPg/i+tEgzT+DGKSHFAipVyehhEWv+hQfWIsE+5XA2HbhunOvJSQmziHcE/yGpxdNxbo
AKUw9h+4E+Cro7GzEaWS9v3BFWY9k9t8txTwKouPIXJfgsl9bA3j0nN+S1gVmqbCbQOb+8Y35oJv
nfvK8As0R32dwAeqJYwkgPSGx0UXF8g0Y3m77BgFbCCtDylCbhdDqw0D7nJ506dTEOlE/Od1kO8b
lllGvA+BPHKtMu6ucqvgjz1LaDJdHz5nFdCzkLdeNsGn2i4Z3yA5N+6ou8x0HKmVAnguqUpRqKTg
OXkN7sSWBnbJHQ/2UYlTCKh6OOM7WZ1vaiXIT31lR9gr8TTZedEWZWB42ff1n/9p7KHhD6pl6McD
o1BOBpcmajvO0APSHqfCarqeDThlGMtRa+WF1+KoTTjOwodhAFvM3v57ze6TZpf0feCrJQCl6XP+
LpTOBM6NlhOGJPtCeG3TC0o1jZZCizZjeEAWhhhWAGQpo+tW5eaOC8azug1FkCGXhZqLQdVEgptg
hjlRPdoIwn81E5+WSpR/TkAbgu0t1uxbjEI7car8gyPc08+lTenIgso07TbZgS5R5bwDQSYvr+BY
GP6HtL/74x3d3N8h0W2gvKgJRCWWVAtyozVhnJInOmtxv/FBFMZE1ljh5HMWLJVUqMQ5swc1jDsm
pkkkXukclA7pFzkNh5Fhd4hY5zIFocgOLmlivZFsfQ9GEC8Iqwf2caPCzlS33L7zUu5evPsbWDeZ
EIZm96UXaRJbSScpMOQWa8glh6nSRu0nYjrRa+am+qaZVuQxmGDmVg2ajHYTjJIATOYE0buEFuqx
ELx+mz0MlQhh5w9uiAjazJQlpLTgM/QLI6wzN0EjjR2PONriUs/AhtfHD/ano2vy35gS61oc6n/P
TGo3vGgFYr6uNjQmHLgC8+yLOgqLY8QSPNIuWpOJfACNhIFTQ+OCKeRXUE3JPcAQ4npQHHOYCSaz
uiad5q/yO9gp9kI+JFGof2bFRzT+J8X6T3bf3v7z5tVkW/8+3O5jZvDZi/AcjhhAmLvzZ3l4S8W6
7Ty6Na+YIqb2o7gz/iu0sJu4jcPO4HPV657RxKHAFO+mPTeNKtbey2d5gPe9B4pIGs5YvKI/ASAZ
iFS6SsVqZ0Uuu0Y1dp3WZHITfAAlF6UvTSL/d3gzQ+FSbNYKFJEeU01tEpwmT4tDECeLMdkoNJeo
DWzmKQ7kqSZ7mQNX76RhVtn9tY7kgXpqZKsceFRxcXBjN74GXoO1p/j6WmuQ8pzcVAKVvcgcZquR
CeEgrDzGZ3+HmKV1Urfb9q/J+Lmd4wgWbeZ9mOqEo3MmUMZtxzhjGaJ3xAcXFegtl823UuS9SDwD
EG7Z7U9BkpdyParFm+FgtjAMxlcNXYPMQhw/HMZKGCEmln2UOLZzoIFHh6pBGibK/NmLVlQjazWB
2cX1R1rnILasu0u3rQ7nSAl4y7suid+F+CicPJ0DCDkLutv9yveCaH2Bn67oBqQY4yfDlu6NX/qR
tFVKaRAtjNGz5aWIfVDkz73uGgHpK1FS4yGGDdQ1VapMn3lQtp2RxICDkiN8b/xq6X8x7mNkPdgc
qujSzT6pmXGmtT/ZLlWGKL40ASV6APoag2WXesEUeSPC8P+yfIGJnSaRYOsg2j2jJMu68xoWQb0v
5VUC+NBLE7R4h9JDWxQZ/l9rVe2HffqWY4lC28eXp9GtGWcL2lZMeDUF62TW2QTZQUz8sza84IHV
yR8HphyAeIA2rUKHDhn2WPC9+ctoR8s5eA1dbcyINS0Thw2Uuni1T4YbvPHy4MnYma0QI1LQakp/
Cpoo/jWIiXOY1HUd2blDDjPU+uYu1s2mM4ZV/q/0uFVMP+7EhaGwjSsgfyGZGdGPBryB1viT0Idk
0U/Td64bs7+C3HX1wU7kqCkMMnpXVYY7gnPaAjk8rMYzMu6J153uL2z3cwc/wxhyZxLr7plw623z
7JoVtcEMIOp0BsAloY+0Exvb6pGDB6gBJZpLXM2A1aN47uJl4LEyYNQyt4VHlgDyuyUh+O7wVVfu
OrVVI5ZDBms0s6pGRrdr9aCZHgHUQJIKF1sd9To4SRxyr7MhobKKPKYtfd9LR/DuPFVhwgZNwEl/
F9EwYxKHuYi5KKht0spbYVucYUK+gixiL0a3gCT2wKT7eUomOTe4GVqzrPmsMeSrDjawVmI1fnYx
bmGb1Lg7u2V9gdnliuxON9jVHISt/iBE89/cWzGoWhx5Dyk2mDlwHghVpQFC0Z7Ikxpg3K+L1kTq
9A0wdn8589rsXz46r9tiT7DRJvB3MhlPzOvlOGh/UQL5Z5hdnX5u2AH3NvAdORB78zEqWlcZLWcp
11zPsLdcnB+NpC4QrnIJrFO6O+m+WB+KII65Ep4Df/b66OTmaIB9UEEe+LbvJLz6OgpJGNBoBMxC
UyYrTEdfv/IrIcFXjVgwxM6YYFmJnNGhJZOnQ+4Hy2ymJiBDXJTqU71a2F6uC/s5W6SAkXTtN8OQ
ApJpnpfBsTz6QR+gNm3OevIFevnT7JdGuMuDpX8q27W0uJLQ9P4BMWhy1qxm1Tke67HoYEhpN+og
8ok9/8xv+wvKZGER6eKFZrjatoWt7CUDieJru3se1sF4OcQy0JT4sroTVHciFJV9uZgq3xROMh/l
Vc3UVeAPhoY0K4yfFf+79M4BRlbEj8l0T7D0oGGesecPI1JlDv0oZpN5TBMr/BgIGYmyswtxypAG
5aIdrC837hUdnqF+WwgE7ruONjTmqC2zXOaxGI0mcLfv65kIGbuJwZhTsg3jVHRQrrenhhIGa0ay
9ciJP5gaRvuXtrtoof4NgQTC3bpMyAdvUp3ZEM8wK06zVlMNz+DFhkG4c24/efoC0zfEegh4tp+0
MU6QRII9hbIMCa6wE0YQSgMzDyblm/OGFnL5iBiryY1fXLaebThz2v4wNTco1+a9/yuIi+FgLKmm
AuspNXg/cCVuCnl6NpU3lAJBGPeqRDoGsnRXhxAZzwlY3ZSESEVvLPsD85ofmS7axQCMfPntaaWY
2hv2pkuh4AoO2FnOK7hHI6LYHyBqGMNloJ46ZL8IyclZBakyjeaNW4ULO4NBxKxAnkNoPNqnnCUu
Lyqv9ocyPPJj96sxI4iSiEW6YqO00kUWQ2vxtyFyB8ylBjRSn0ikXaJsJVDFUQ7wLzn4JNsSQDuI
dtIJ4oCI9K+f9Cefje1ySly4TF0NfD2ANQFRpWgGgkeyWbY9VArCxDkFoyxhSWCNXwCb2CXGg+tu
M5mj+EihrcNSu+0JYaIif/BYK1ceRtRbgmZiv+KbLYrJGRNWOWlRAZ5iPKm6GkHVJOPJfPKgQ7PI
3H/UXARoprSuOtAAxBi6v1zaaFq5B8OUX4c1qZi+yG5tGLyWpmOmC8ED1X775539t0rOyHwDe4yv
DG1nMd2QRRhlRsmn8uBiNHodqkhZ7MiITr2Iw4yG4ZN9/73lgr1Pomby7iIccGVzrq42HI6uPyMD
pbDJJkJK6l+B9YzJuIYc7u/3GcIr1Fpf5sdsyXeop8ftOuNVWs7oUG21Tatp/M1vgSXH0/x1klAU
VmuSd20WozivKh5v8hYpv0rBhdXTR5jdyl9OBi+P81IRZhTmomsl4ZOICrQLY8+ry/xOPBIWMTY9
sY+rBAz+Z+pWQoQzLDKPtePMuOAuibmMWo/YEc0JsSkhYMTfsMMqe2cXnBXb/+Wn42ZiInlHehyD
Cv4SC09hY8Cq5v1rQYzb8wc9FIPFj3RtUTwF/kE+Gvo9vzQrmg0UixQTppPV5ro83U/vLYvByO75
odeR4xRmenj7wRC3lDa0zhgWWwfRCZQ9xpGAPXNAu7gkIwp25VtcaHXTIsmOGihn85pAEC5xrG7f
SLjVMGTrPpeMtHPgdXeZbMzuNyTATZLylAcq7xPmvvHYVXmzhsY5w4Coglk4s5z5iltlN52BrdjD
m1fghtoSiq4dCFWwjzl6qqaoHHQII26CDzLGVx6mxPb1cp/h3bthjx6hHVdIBrC9y7I6rz5EiGbS
TPrrk9IhceP77derhINBca5ukcy1zYdCE7SmQsMhtk2x8BJpZjL5ildgWynhboLQFfFMfCAaOr7h
2K7461qEUVQxp4KQQAFyiWjlXWlIJ+ISu9q4OFnDWw296wvL1azs6Opy4wDDl56BFTuylPQN2aGZ
7aUQszXbXX0qDHK7nhCuytJJ+CrLF1leHbOgT0rMx7JxDsJZ9ERdZhKNOmhWub64UFwSBQqtR1M7
AiPUO6FQL0HPY9+zoszV280+E4rUi8lumngOcFj3c3/1dDNXL3DLPx8QQF5ttiuEn2ZgSwwtlXs4
qmTncooVq/qw4swyj353vitqDdIoT2xrE9vIBwL1F7DswGDJNKat1aRBqOaHaQHn9eI4aDMD0u75
3aXvZ/F1jK6BAI2FyIw0DrbwNo9kKSEqzGcblU/NYRyomINd0OFVBjI9304kh+YSN+fhZ3X3uxd/
QHEdbxMdOluSnbcc48KRdXwlX3pd800ozzCIf57qRPOUkwzU63qeSKG+iCYBWX/6Gew3ObqZVsjn
13ecwvSLekfJmg67ipNG9LnxujsyqH0aU18udGeRD0BLcxW2tsWOLOnYyFCotqqgTXYt39O3emVR
idxAB/xW9NixpOCdIwrqWMc37r05npXRr+m1OI8ko3oDDcETCwlwa8SwsuQv0/F9w+t8hmNQj7TQ
CwoGPQTNE2Tj1DIH/OdlGOYxUqvy27Vw/C0gW340Lds0lhGPSMckOV8IVhu8tbT75vbuHbm8LTOM
pidYxNJI9cWmBwJ1SIQBqbw60vVZ0bD00j2CDe6m/TcA8u68uLzX/cLWFKzyKW1trBBrluLUMeDE
kl2q7yzYQlhfyZ+6A5jvxXjjcGQObaRAmKySqmEDQrIfg99XPwp9bv21u36O6b6xXsDRDXVkbB7d
nEoYTDxYHP6Xc4VGVT3gY7gYpe4QCENvwryeJ2qWat1cAt/XK1pNAsXFgQdzQQIFlaZAsz0II55b
Dabn6qU5wki/ci3iFgG2n1/W/D1uBoqC6LOyLdR1nWT3d96UwvV7DX7uhYvP87GEFkbLez4oWjqU
BsJ0GPjctlSOUPSYFJ/nq7WxhzDt2RqFhMutNjmWTOZ9Pn4I1qGy97VtB0QZGtyun4tIg0PFEWds
pgEdzvAk32M3YeZZKOXAlQP2PNk76kCbhV+QRxkZnm8w7kxpzZx+WapE+FGGZekXGQoT21OJTNrb
uu+TE3tMdQVxWCb9HltHLcHfFeWSucghVqUdjh887En244YsUYWEle7mwQK7E3Nb/PqSXPvxaCJX
pk80UOhVVwc7PA0JHmn7QvzBSZmSw4OTFkt7WU1HHg6kDMa54slu0EaoSBsFxu8+Lftj0boEKSAb
64MVfDNebJSeXoqrUKX/FbW4KMrGRra3R0VPOJlbEY3nwtRzGjOed96Pxa4Wx6OeK0vln/N8yYZ9
5/1OAtYIem50TyXVKufLGW6dzWLEnzrFImHUGzluhqG3Ib9Qm63ijq1iVuJaj13SX7joSpMC+V5v
E/Ed6b0SUeAXHoQUuuNQbD9TTmlGTJ/o7Q2YHuCpIhcZOHou5AgOeL6c4hinSaiB8rStgIXhnC53
cwUtX3Erj6ZJfIxGAN0pLmXeOBmyqjFXacgAd34JKxo+eaj8tw8W/Oq2X23TQtdDn2jfm2Ai/YB2
hL+SgdhNLeRZ6GckDSDkT4l4PSUYKlVSGMpClA3XmPqw2hhdXx9sMCM80RETMi8RHPasBWNvo6Lb
NNIEVH4gR+2YNqSHDt2gACQhG6pTdawPbKF9MHUzjClTz9EjbJf7eptF3Q/Rfm5wvon0/BFy2LEf
x/1fARW/Ezpo2uAwO2LsGaeYb/RJpjfXry0JcxQ216J1jB1F8QiRBnUmVH9uSaa0Q94OjcdQm6dU
KCphiMb+J96W0q2oaYJwYsLBoyTFvF8+11i9prJrDeJNtlZLS2oju6JHVaHzIpX6+QnX+MPhX+zF
oqAtlcURLt/06UeEVSmFYVGw4fX7g69leql2/TMb3U6XYnUvcfu80igARl6Bh1l4Sk2RZ/r2QYhK
P4gV1p0C7+66Ps+hsOYnbU0MhsbLTJHyRbdGx1lwPZB3CpBc6AxZgfs3h/xQQYIHIHFBQ+5j5/Yn
KCo9Vf4e5Z9SKwdirHsR7Sr2jEIwDstjkhkvOy3HIVy3vqqY4r878DAZEIGo9aZNyXbOrGUQvgjl
5E3P7eUG5M7Nm7eL9BO99S60Lf8rG/U+l+72qxsu7py1bTPC5dzfGTrBoc3w+Hf/umMIU26TQ5n4
rPCA48W1MTbGzqj+oCBS+xqHDd+BS2ZyLu88NUijPuvS6flqxIwzS3vNljYZRGq2/AbT0lbkxkxU
hv4wtmHaRJ49PjPxZA+dl3qYgMsKgVVk7oUweJsz007Dwh+APlrnBzQNG/Zt24MZQzioo0Oyfkcr
Vi3VOxf1sUoD2TNriRjKQmgOP60je2rvtR9mg38fiL6dsVhYAapAg/Yf2sezF39z8UQ9PRMup102
NCu6fag4xDrJb1dRbRPu4oq5UqGqWRW8gu21DmLwtkhiICbXDniiYyWZKepWMsE1cI2tGSzHHnM0
djAtVKYmp0o3jxcRNjjeRVvLt+EKOx1WqplZsblTzCdLYp6VKwcHVo4S8LHD1zfLVkZtwnn0KNRb
5T7u36Apzejo70+IBk4LHIaWyuZ4SlI4J4SXmvYSmIsaDgoJKUeUsuCjjbftBr/SwtRc6zA/xtlX
iIg0E+oxhDFWiNpEJXWXRjT3LWiA29Woqsfqmo1tD0xlhGi3GJHkJ4aqmYcqqjvpLn9NdqmT6lx8
S8eO/eE57lYtdqKa8w3bS8KKUhZm0T/dgCEaghsVQoKZqY7s9X5TU1SNweFzrLyoBBcNWu+RKJEu
LGAIH7/Vx9JJGEZc4hPMlZl1I2Hcr867tXZdKkj1dwyGVSdH85o4W0hOpWzQv+PdAbHpsplU0MBF
ZViSU16am9qFGSVd4y4q11rEiR5ArYxTF45sKG3ulX72Ax5yX7iYwFEPmmipqjcgYWRuhlYz0ekO
RJh1rO2TjLyhUGFnrwqGaYFlLzu8nPrwa7YLfbGz/5zB4fLTsh08/eSOfC9BVy0yHyMiL275n5rA
uicJG9YdbDT5Cuy0CvONiZwo3+3hf4yZyxm94IBLMXKn5fmXj8fYNj1fXMfyGi6eH13v8Je3rRlv
FxtDdrnl55a2p84vPGT4UHLNxl/VPMZcd/siGl3DxRSRM9tPg45eeV0DHpC0zoSweGiVaXrXRxeS
Z3/EdosttTND+ovS2WlRsWubIrJ49WLcTz8TPym/elOjON1LogI29LmJbwJ2Zsi0FpDn6SPmXq8d
UTuiyY7uu6/48vR76ZGwma6aM/EtTQ2o4QmVZ3FJArWDK6GZXqbEKc3Es08U/aFM2VZk+P8BCLbX
3rtDnNnDOH6Vmzpsrf3XQum7ezxDB7+DIyPrLQ8tTu0/UjZXoiz1kKGxPAkhHI+S5pXOLSoRbnkh
HEgV86Sg5Ysd+uVq12khDA16Zu6uERx8ckYlenHXrvghcg3T/WENlcwt+XjUtsGytMkFpbzv2wFg
Y0UzE9Q6hk8Yl1UDbbS3CzcH9xpog+lgF4Anpupa+sShKCeWrCFpMQ21BZm6fTC3I9HjSu53D5Ez
mdS2ovov6gMBgSyQhqNmZnFZvOjK7KIhkmqK4gSZDTAbEiTEy22uwhfBaAb8zvCEZlgGXHFPXrco
w81D85rmfvEjRwtlRxcL1BKVEIBQeJ+QAcoSswByucsVvsgTG8gTQXfls0lNwAGnfH12sIrbk/s8
1OmxZXbedU5vW0WSYmTu6lh7ObvgviDa7kdKWBtjwx9mkh5EnQKoycuajjkvFQTyUnF0nAAqtN2W
2rVauAJcZYM874In78BOgwJ8RGxRxg4p3JU00EszxZijWxnitnL3zxJc7loNEHd44AbiiqM9JfFP
/UbuDRBC+nJ2MMOoWD84A2OkLmZgeBpnjPPqkOLmEiMaviEuhkn5w9VT5htlNeqOUWrp5bTpwQ9p
nUli1ZlkKh78giKrAG4KvTh/SbFlIIvKpA00g1j3FGEk7W4ODMWaKCKNZNEYsKgbV9b3lvr9rdx1
zqtULuyIRoOru++kOimuvpuNlWz7oCVKNWS0WSFC9XNv0lQy9GRBw62z5emSrxI1zsUYp4N3kgJG
f4lP/SJr68sjtT8364Wa5AZaRx/O26p2SxH8/RCG96YRDthdyvus9RqNcrpouFxSoOlmvar6OmQ8
xehNzNYWc+DMSPx5X3twmmebQxn6g9SRR1M34HjDxSUuI/cvgDFJsRUGo+0d6NI9iJmYBJ/Ja5Ok
9H8Bq8BY5KIMnoJoPzUHzmEOaMEPeVhzNKbsNNh9SgB/1heCFbsnwBxv4u3WXBEtIZbhlHdX9ehJ
bZIF+BdEFAknltpHhA6HigNWLP4d2idHXfq2L8T36gx0t2tk07spUk9aAHuD/4Aie2rse6KPDJov
Ix/LRLbetrNO4IrE2lgSptuCo1hnKS5mceYYI6vFJAKH1sircAQRCAkaacnO5EvOeTFBQSQ1w3f3
5hAN364obK+f7c7/PAzz5+I8vCtcVjNel7jb/be9apn+KVyUwg7xVT776pk8JkIYxgPyKP2Yaq+P
xTxsJvOltT/Inu7XSfoTRtElCiQbM8fOfuy9pBnEcfJY+WLHIeLIBiY6rWT3FPvxBzy0/l/tjcki
kviXrtKojf0S1VFSMw4aaFf1GbVMtwPOw9wJdX9L7CyPzxtseP5tvcLIN5QxtDFySA0+i6YYqMhd
kRPIPssmmAWe7BE75MGw8WgcpD7qOYxW9f4l5DwB5sjBrUgWM/Ou/HUN2aKlCTJ2oi94cg52PKsS
C2/xeavykgzLK2qik9hHx1YgXdOvZDoS/XWUHcbTStpHlLSg3ahFxelnsddSvJGcNE8CR0efzfkA
GkA9RgzF73YtlZ4Urw/nPHRByIqJdG0IsYAxkSoiRzAvDHULSoPXCDWOLx+GBsRj11h+f+5DAdh2
kWDsLYFTgTuJL/rVnOhZFJHuRuLgK/d3/ERhUMNi2Im/kfNqNCtXeS7o3QiDvEoBManF0qyz+Kp9
Fu1VA4gI76iF1JmpL+S4CXYmlu62BYzeuO/RE3a/9NtzWxhSFU3fwShzJdvQ5vl8xjnwywkJPVQG
+kCjuHglhezdq0pAb8dJXzWdPG6D58evJ1/V0UJrDQ62XKh6tjzGUhBWUjP90zyfPo0pB1cy9Ulv
Wulyk1Xl2QO5+iRDdqpCkElDhZDNWKFcsftXKE7MmPE3qUb99CS9EhZ6bfk/GKFXYpz62Mu62NjE
Q7AR6jgFuNSuAROwydW+iXzkf3EGMo5E8XD8URkbP5zsQ9f0jR1+3l1ov8ZX0phigJxdKDpV+bAi
wwLkEzfsDvBirSvBRrvUwKxGU5/7p9AwYNJI1QqrMpQt763cClrgvb4WI2NXVtHoC5a9MANZc5iW
cruCpcwKZCJ3fivhiEyPhiy4PEs9gEoNLyjqcKBXWR1Ua8dlDrgEfyVuc3KuOpz6mKZI/BGt+keH
umM/ZAPaQFzthw+Syt1gADtFe0XPzr4Jx7JEqwFAo/nwXIYOet8HR9LmEx0ilD2FXucOfI4ZbEyr
AxXfoG0VEfiPoT+VUvmw6ojb0vpqN621AWDTNKs1ayOW8JmNNScv3jRX/tCOzbbaQKPf8AIv0d1s
0TsasPeNZypVeV8BhJrId0O+8sSUM3lXTnsz/f3DbrgPmX3PfFY8gP6Sduh3+eaWZp2xr5VOyrwW
2saDFnzlikpZC/4s0yUYXXVzjatA/guOMPCtmf++iNX5Tp6V5lExFfU2FrfoEAbsARmNvLMQCc6C
8htytS0la3YPwsH7hxy6A0Tls2an0CRhbMemr5IDWGm1QcG2PF/5cwPo0H/VkLOc6fgsZ85flz4e
hmmyYmFS/CA05JioY3kUH8MIE+wGck5Vr+450XUYpWFSxOV6yElclX7mo03/7SBsuhX26JDoe231
meoYgZUL6c2sCLxinj18ol4JoDPtubPVuj+XvGOvgBJn0Gl8awelFSRG4MQv2PiJI37IHe3STKFH
3rgXS5ojh/A4E68q+l31Ald3UI+QE/fvo0+fmHBgQnZlQsQNS4xCR47mOTVt/Uqg6eBIRopaOn5b
J8jVWuArT1fZDYok/uDWwXU84FnOeeiH/XWUKW1cBYbWI2PUNKr7jA41PGpKjl2f9oYhoCkhGUej
yfBS4pH8ujIB+elDZ6ZaRp61Z9FFCPDuWeq85cdz0mZORzpKDRia4jdmvy+tGR/HsRx35+lb78r4
yj0xFXFVNjlTWKx4c4iY9a7cWlPUyxzmHpqV2RaspXtViXR29Ae2adVEdOVOpT4bDkc3zGKDNpTy
3zzVOdKngVgCMQb9mRD7K7v/n+ctzC9oCV/yT7b35RaCdGlR/q7CR6+j+LcIMEDuRYdGtxn4U6GI
TZK5Ey3VKoMkX/xk5c0TboqARXnT8ihfKcwLGPtBuMGVodTkBVTcuvwiXviLxglBG2ybT9Wx75WA
GBmuEZoDD4CXI4GMCDu4qd5/Sx9fnxTlLxcGd0radfDpvL8896XCSULeOo1BrNoeiwEbVFkkhxHk
VAIpGEHj/E6w/DD67MSW/w3ygbmUv0nnHgM0bg5a82O2wzNF45pWs665QO8PtmY1WetzWn7nDrZj
oD4e8d060OEV7seEywdJeOZg0NDQkH5uslJmexUixEQ+0oTTJh2ueeqfxiHHbCZokLMSDzNOfHLf
aexiSzK5M5XzZoBjzlsvRajqAhL9ZR9aG0RL3mqLAgP9wWq3zIZfYm67AWcXE9V09tTGgkuWyL68
Cv/5KsLf8fqX3ErqJ1zMrgYi0A57+fio6M6hwsJFINFDcfjXgpBwniM9okcs6Ue2w5CUl3moA6d8
V+VueK1CvDWKrLX1JJarm8nKA0awfZH8IXC5USvMqjKCudZcRSMhSkj5i8anq3fB2o02uM9gqjOw
xOCC3yXGj+eIc0qP5vIX9fVZUzIUW2F5tH1UZ/FDY1GbZoRrtUHcZos+wBzxxNUr9gMD6aKBQHa4
z70lwEzeHAl7fDHk+vLXe7gfAHZnfXg6mPshasHR++ImsaTWD1/QiCXxS26zcF5B/8eUR/scaKPP
2P9aU8c87qGgRoLYSZ+QCcfIViEB7GvUoH7DPTGq4LnsHaBd4UT66Vsvy2sM+fPEgJQhjAP9RpM7
cEFmJ9+fiI3a7m3puUd42O6Gjjw0mcI/i2EW4Kbxb1zvNC0PplytYvQVEwJwCPTi+M2OD2OrRZb2
fYRuNy16N6SBJF4lQl/ND9rerj90g0monk1QtynlhkgZT2vfgJx6KTdQq2JbXKBMKXSJinMSqVow
gAqMEDamwiN+fXFerB6EDH6IiePzorrtn9wd8n6Bwsn4ag8D4NdCa10MhU2JCHjrLWRHUW8KepbM
pdyfjjH/FE5p+3yWAla+sejmVioI14Vz8MidtS6JVfgmfuYu3+c6gKXq5BxdmOMbqQkj/nr7Wo36
aAUVPBNaXx/VULG69SSLXu24NlQYodiqsWbE/c3lBpWTHjW9958b8X6lYX+/XSgZSnLzf0Ri6XtR
os8NH192M+u5NumwHek5g+X++ZLN21a5DH4rGJoA/xJiyvEU0v3JqUXhQLyny99upxCoSVxgK9vK
PslV2R4m1k4Jvs8EWuv7Awnv6IZkUhSGevhvea2mqEYlBfgkoIrqUp4yr08PXRhT+MX+2Dx+9Pzg
4gG9nR6Uw8q3eUTgpAHRGsPYOIWMuW3/AMH2tSbuRUp8wK3YaN1FZogJfNcWQxlnJn/In9WduVj1
kfcGu75xUOy/V1f7hiymUvHJwxMCAhiOMUaptG8Bxq8qaStVuXSC07Uewps4FOzzMXkywAeWdeIF
JbztJ4YJVd5J6VdGNx7+07aE/A7k2kvquBjK0R2Tv4MCpkgZhEkD6X5DglPZ86V+3vU6krwRDzL3
YuplNeROfvW4XMD4SQ+g+3WD8aqG6EbkbhcmXbLfQcpO5JBG3dSLRJLc8S54O1yL2wK8BuFcXLS6
VpoPLb1lJnMKNRWieI5Bb/7f0UTrvJFQGX0tbzsrG2HUnMfCDwu5cbT+218Rgt8m+fzjrhb1Vtcr
EeK/TEC7CK7+FoguzYkTzNlQU1v3W0638x/w/o0Lp8ma8qQ+UWL6IWylZrwk7ovkO6I67r7WGkmi
imGrRDuhtBvs2inLlgfLvI8wrO18g8w/SkpfO1N4XpIHJpZc9kJjiSyFn6JXRwJoYUwoHYmjMpo6
g450Yl90Ugh+PFVFKUbxMmjANw8pV2rv6FLxxnsCAe275wctcckUxt1hwEWaKgz7sN40XFi7FcO8
LaQT5JC/mxNquccuedG7pVaKOnStc1GK0gF4gvL4FocO4uWXpUMqMwEM3k9EiJxKbCe17UCc2wY5
Fv6mD5alsQKqd7znta2ikG4D8O6ol8FAB9L3KSxxmnJGZnPYwA0EnH4YbHUwp6icr+ZyVqtANgQ1
cAxLclXjdWjvv4avE6JVT8Ni76HIxUEAPoX/QXU5Y0OOTNAHVuAdJ36rD94qFOhxCR8euJrsGGaT
pya49xK57mzckGbMcz3OW1uBRGIC2bfZ4D8DsHZjWSFIaoKd/33TDnnWFpMHPiIsbgCt79if0dbU
cTZY3pF+64XRjIbeJIFPeuPsQopsW2OwdshBSCUP2vMr/fbvB2XNtIeiMcC6bdDUE6EwWbDO+ucb
bMu7tGwnrWHPJY2z0wlSGCXlx9kS9XNkJCHLYCe3F+5FdjCLK6qOV+wkjR//ywlJi+Bcf34EO3hg
p48LhHe47EFqQilNzWylU8HnKJKaQADTZEoLOaoZGqMRAdBX7A9BSbXCpwjJgsSFGmG+145zCOaM
tvamw8/dfotS4x48f/Prd7qw9MCO0sI8J63MAO7ympHQRkVzVANh8ShMtErWer2gmKknIM0D5Y5p
cwqlBqNHX7opIbwXoT1yg9MQNSHwL4oKGWqAn6pBya3Kkn2mLQMS1Yxx0k+V+rBdpTSNWX7rNs0g
9JKpcOcCsMqvZrCtAgDJ8eMrqgrAf0XCEigMBpLyKENaCtmbIHrQc2W5sxlZveIH6WCpsOSFc4Y8
gpNdP9s2lafijHFqhIi17wLayx3hTN3MM5pqtWZdy8nnhF2t73qZ9ReIjHzG6AT7SHOzqviGUXwg
cM7uBIiH+JBaEMxcHTeCkwBbl7vLlxKbTYWEq2aMcUwxypGVNRxFnewjIAFL1mvugAuxvciFG1OJ
sB1LDHx7Mx2QgFAD4nkxVDdSILmmu4gFBuYFtT8p6zyQWRdHnqiIdllU0z3V4bIY0ZYzg/pnhvgZ
vn/h7qWPfAq5yN2xkkeN9gTus2fy6wRfHcGJTdDPpnSN/+mCP7f9WWmip8oeuesB+PMN7fCdfLPX
HwwkWDoEygTUF5FEHcnn8AZ7Vnz8E1xqwVxS6qpq66NE01FBfVyvcqu25VL0UpUdIqBstGaQ0+st
Jr7uCU9SL/t7D6ZMRaksqYou6ZTi4puWL53xI1ubmm17UImuBzILWeg6Nwv6b/gTomRRoObGcc3F
G8wNanokv5rAcNbnEoWKU1wusKui2vje8+mHBRHgQOCA0DcHNjET7Tkt4BufWsQg+UcSLubtj13q
Ky5lX72ndrnr33DlNlzuDbTKQs5MKqIZ6YoSb6i0FO/oR7D6U4dngyXMJDNAF1NObaXQ7V3rMRbe
eqZwLtEKBygBlVAdqc78SNQCA2xH1rQABDpivN+BlFL9ojHJhcBXJc6CHJMKX7ebh6JkwAPyaJ8Z
WfFhEKKMA2dMVcxQFJJF1TH0lo7pTJDcw79opSH7FavyWRzba9Rg9p5VpGmU5AeW5zypyD/Yv9H4
3HA4BmQNSI6uzLmT8S0YuKoHUnrCFnvw+TP1l9AqvnNJDLR+m3CxJoH9us0g6fWt8wVajzJs9kKV
vQX7f76wjGlREbkOa2dZM9DAS5ciac+TjL0zlMvm6fO/o09j4MzlKsAaGtydHbMNoMfBHX0qR02F
lt+J09wiZ9tOPKGSkmQMhk6+mjSimBz6mDS92/vEeIiqvZ3OyYUdS4NWzNFSwA+YMYIaRCm2vosT
nmg5PE5t9Yg6Rxhp1Z2uD8d519zN5+w5QFJ85cGvuiO8yN5iy5ej07eZY8qkfErxUDgTTkAFPlRa
F7iSDRoN9u0wIWoCb3MG9nsjEvNPmevpUBIW6II4BvOnWcygBqVQb2p/BHk2g9KODVkbFtr2WVUm
8G5G2NJUirfdZeG/Gih9dsuwg89kSyjXKSiGWpthc2+sBV1qkRt/VxQ7speI+vhXXfxVFBZs+Aey
k0yOuPPza8RT0jymBImFcc8/zjjO6YMdDkn+zAQOr8nenq9IXaYJP6jjlhZ4KCR2LTcG+p9Up0Ko
zEp5lcM/1giPBl4JCa76UqGPjO3/kOkP3ibnSStdLCTccJKDgbrwAoyC3+75VqPO4x04jQXzuX+C
npxELJFUU5kMuJDvujW3QID45x06HiPevYEIWZQP22Otj1lI1b8U8KALpVYEscJVlBisaY4J209B
kbQ8jjQuvCtbGMlctyeOM4IAerBEQC8HDKypJ9DDyrEaNAzyy/X2/oyyV2lNjpE/AwhvFKSvb8ZQ
CzHmL+PnaUwtiO5unJwxd5LdyiW5CuQM9hdGecON3lnkAdTdxYifD6ZiZTDbqL9D+f8Ddni3H9+N
44InxH84YhhdvXCW4OTE3GRJvRGBds5PPgl3qvQQ82SJApSGn5GoBAGcVq4eiWyDm5OaZzLbGQII
XEUsOfPxjiJwGwerDp9/mzYILWfa9v0kdoB3b8KYXcovFl6gVAeWmHZ0pYq5d7MVfhIQlvyU1si6
eXbJxt0EsuoA/tY6/WBTzsqzKBs9efcj59/dn1uOTAUMo8Q2r9pXwm2p/h2DUGJ69Iw+yT0NlvDi
PopQu+N9CuCkDWCogmqYxEXeAsp1InaHWRZSotn7QVOTBV51GjkNXh8yDtNKr2BXL5LrA0T6U33y
Cq4JsQecyXuFhOI0rCYEZbBBByNnAugM03pfaeE3Cqh3bNE2LsMXMF/ztxtXsDZA3nxT/MMpbtJD
bQNKyU7KqmVPJ1gYpeVHXCKfZB9nFSaSgKynMvVwUUrtSkJ+1mID2JPLn6YJ4kIHN76zAygdKIwo
npcCqF2ybEfIeMJSDsBeXAUYvUKOyZZb9MUQ+yi/xQSFOleLoEgIJXi1jseOPc5/WLlYSqbtfEhL
MYL5t7IkcpVQ96QrvxJz+AgdAQerpQNwJ+NgpNgioUk6ICeJEIJitUckAGeOUqO6Ss/BoAKDq3od
eJxK+PUSC561dfyEMuBImNThc2AbtYQQMOaK2lBySrTqfCqk/Zj9CcGlwm8cxGfMdkN2BA+kcjK4
i8/cMhLnxhlhuQN5wI5CD/rqC3mmAKgdOdfpk76bU22c2CliqMHbv2eMVJ/MNwaxs9W1poQgpf4r
IkLl6RalrbU15NDwfsjytYHD5ZrR+G/oUhS3G0nGcFA07ESLyyJuCV2iglp7c4yYHA+M+CuZza3k
VcrlxBxJj6Gk2j3kyppUGz6Fp+2v4ToTq1LEjSz/TvdH19bnNUvuEkA0UcQKwovhLlF6irS9BlVE
RGzgX8nfcDOjzqw4i0XVhQ0g4gllmCsYNaYWLbJYTZ8UX/LAun7mRZsDphPl+ZJ0jZTJzeG6vOcu
fsn65370NepJyEoXgYWTt9S883BrgNr91GvcTS9F15Kg4WdZKk/EhSCnlIentN50tcutxtBUEzYX
/60VNZZlVxVA5QiHDcLa/imtm4M+Zuq3datySZITh6PKIBjKAl/wDGD9Ua0mBQra7IoXQd6nokr8
2rud1TOHwsGUcp1+XwkKABExYOQHQvFzt1hP0UkvQcFygzavtzCehqmSUBIC6XJo14RoaY4WBfQH
rrFxVGY966Ht39aNl8XUxO7gQ7ZhGXD43mldQg0I5+BufR0Aymm8ofKvVecULGVMlK5VqY4gjbxP
3E/5WfmQs0vIkCJicfwfW1yYWQXQ9vuynMeds6P/d2SMRQRGgHHnda0SNXE1qZb3re+RcBHV91Uy
+Pg3viace5t02/7vyO+9XadK/x9Mp78F1afMVw7MV83A20nDB69M0OVT3c7Aj1RjKIc1h3Bg+VV9
yMY0/SwfIj19r7Ak58T71IO+fIETaG3uFRLiEG4HSyMKSZo6S3MWQnQ9KcYTnXGdQum62iA+gCZx
dXk0Q8IuxUBm1RwVFRW/xspz9iUjJZ0TdWjlQJ1vWdMwnDo108WxbZDLefhoWaxQU8onr8z+3ucf
9siYQ6R1HBFTbtfIXaSbnCuSqNaIdvfPrnaP0UVE6+4/v6GI7MsXTLXCgrfh1x2f2X0dmtVH1E8V
+9vgofnKrTNELgMzM9TkjuAATL/hS7wtNWbME03w5Oh9+Tlu1MLuHSgAaPFhthDXJ7yVlcsMVKiD
yIObLPfKSH1t0CjU6x7dtjh/XB0TsPNTQMXsKnRN9SG7HloJ1MgJjDk0/HAge4M2nxnlwXW37BIn
+UFWX3ou5nvGKVUrfcxnqbP0AFNypI59c9Tf9RjG4WziQnCrDK+f27axfLgM1317fyakv3ttpNI/
a3gXO56ZHd+/yZNwydPQAGLYW04VeN3lVkhtTdBDpuuY74HsqNYwAS7VPR3EC36UbobjCovoAISC
wB9gCNqgp3d2wXZo+A0tSHyFIJhDmUEByRPHexVlM4EIXUuIr5NaruX99VwRFjiSO6vMexrNQ4IM
s4faGf1TqQ5irqgmyPGv1KnsbE1ii9qCniKOmt+5M2MoYwIxCs0LK57P5PxvgVteWp7CsBh3blRi
y/L5awccJsY2yFHcoMF52oizpnLebh+wP0Yc/IhLMw2QW3GVhuxOB+UCphkiSmDCaNuEovIVDDwN
gAN4xcys2pKC4aeC9FHkcrImuCv6GfIwBo/UrGnV/PYHdYtc/JC6ZvqLbPjR9FkbMChF0kVXIqir
OFFMCrugZbzRnS1dRsZHJNjbJnb20k9Q3ytumep9M2jIu1ax9PBlZlUd9KueyVCV3WH52zK0SVHF
Z1Y28DmYYvM1rJLixB4Z3l8GW4W+tqKFqGg7xgvpoMmvqXTwU7EVrvpELfA/LTujfMWVtogYD/FN
Xm47R/iMZKt06/e4Q+VHRhOcJkqTWnVYfwQM5fPPiSxQqTSErPWQiz5GSrOYE7AHfFoyUPsQJkZW
YYLRQFkDvtTn0kDm+9ibPxcwxtL4+o9oHZpIw3dd6GreGXbNAEd5O+wwxfjr9Z8GxgmHCdONSzfz
Hye2xLn3ZHYkmrDOjFnxZdNOF3QVxN0D0NJmr7U3FemW8Lpg4ci0+C7J89YXrPd2Wapm726/QWD4
9IPEhKduODTvmg3QJXvMj43+CFP6FiVB3HnyFsL3HVTfZXboqNXaHQtQbz55xMs8LSGrx2mSuqlQ
jIzHyCHmqDq1laTmyUdb41SgFmkZ404NuNxlyvZQkbOS0jRtEtCgwD2juMdbCg7dRFzY8qlggd0N
zyy9K8lvYBIPgzqu/uFAs/P7PwqJmApQbxTL9egPXUgOEgFhjOBf8U98F/Z4YanucoLXhqJz9xmY
3uQWASsWdgPqOvsX7gM1bdLfH/1SS8iDyF+c4xZnpUBlrPRC0mFDPOb3XPvcVuPr5OjMXFF0PC0j
GAEuHFOBsowHvHewersaI9GAboSSxG8F/YskF3Q0ezYxE0VbCR11VmRMekH++DYGGGPzLmQ991C0
wcVCFbWW+T0TgEJy3jGgxa2MFg5ivTrKSI9EK3ANDfQCozjSifZbUQ8X1PJZzKlnmy18nROiBVfJ
RCPthQwYp5hIRBFfYYDCxe9HMZbeBRBdSahwdrO0WQL0wPIwQlihzQJ8Owvf0Glm3lls0i8f4Rx0
JuX5zY8SrFSW8/Z3iXDSvC2nsL6Bhwq+sbbmOQzEOH9dn+ZwGCgwZf/mn8izMKtw7vG0xGvwrVrO
Y25Jswd2uJ/ovfDVJXUmiFuOhYCnbEtxbq2tUqF76Yu7RfGWKj1cifFBbx7w7gv4QEW9CgCr15HM
ivm6+Ie8XkGAdvN7CoU2nedWF9ceybFLcQ1IY3gtuPDHtabz2UVDq0mmqzTx0TYT9ZsYcovtBcAf
shobmwzA3m+4/WFDu2VyMmeOa1w4FfpRTEyUuwl+imaXhmAK7upkJk8Sne9BS1M/bOEV7NwZ1Ew+
SQM3f/xMYbgzJ5lMjlusuSob7Gso9nmFpiwTovuAYPjztlfzklSv3KLv8HcDJ9GCL4w7CyiSQ1yu
9epbqTaWQbp2qKEgS+e7dUJ5U2xd1qznZV36KICDWquoAuXB2bSZMAcjmj9NC7F8docRczA+MudH
xummuGs9YtEEV/nPPArYJeQOg00SlQObnQitWs4zGVisd3IabYFRQkiOQe4ghYYQCD3mbWzPn50Z
hVTmFQTndmyVW8sXmWUUMHz2HBggW8JHNGQsUpA4Er/m7ruS6ngg5EMOMLXQQRidjpgfm02rrlVl
UPiTCdsHjiDKn3gQkvfKdF4EshVINQMPPC6Y/yfSoISZgOjjZGmMa6yKl0Q40wnrt5het1jNGXNs
nwFzU0tINfnZJkN4c0fXJBPwNwmypT9swiZg5TkOu1TXjv44cRBNbAJsL7T4V5lYZW2hLgQmZ7XU
d4MYSBVYne0ukZMI4eet9Ru1lxo18fUQgx46uOPvxXNu+AlWm68LDGCp3ZrhDkseHZWz+Rc4SUcZ
yleMRhZ03Im8drpBB0PY8DebOmwVNLeqDX70VlDHOLRog5BeXX70z7Coq1Fpgg96d8caiAnBhJkf
S8Qag2MNOhLn0SHsptY97Xabr12Slmqrc2F603caaWFI2L3b/G1+79z2I0fKnBnkN+nNHjwqYrT0
daTm1q8RQJvx1UH0LvMZxzoft78jlNYzwruV4ClnxIJb6pfX1RIepdl66JjqST5583z4yfO1hhd7
9Z4bsnRP5oxjzfByiR6WvFVHAuaj87sM4HSuruVyX3WmV0rjYnqapmLWlMh9yUzTJmsAQJ5vy/nH
6VLTcEPaQAc6zQSQczbRKJpgv2Cac0faN48wimwevpFFZPChDdEGOjQxgIVRIwcmpYrAJwU1a74/
3vOQS8ac00sQWmiIdvs0aAmQ6wEKkB1hzKeRu02mqcqx4oq8/rB6Ee4LlqtxlB57aCzKJu5NUvCU
tzbieHwUqwGlPMiRUC3LLBZ9SokQe0XiPQKkyuhOmlS2QU27TA2S4/AjE1+uPq9b6amZAvQmnVuq
K2JLT5L4G5P0T8Yl4pUD8fEloyhPq7x6rf1uKS5OFrXt35mlf7wGivcbnO2yYBD1F0FNwS+br4LL
6gIcMqO4UjmI5K+qd1ZM+58jg8vo0xj/QtZECtvxGxZ6o5w5tiDkTyC05Bjwt0O/qSBo0XMjpALv
eMSfopy9T8hvSeBhKA+5uhoiAUBCr7UGkB9b6G4xIY70U/hnIl/lHzLCecG5eccQ1wS18emaftML
+5Dzg+bzYA79HCqMiP5TkxIdDltIgqeh4UxRi2x9v8fKY+4TsXTuAUw30/f/YaBMghH55saBJ+hz
wUTXrNbNltU5Ig/sNIvi7b5yXVy1swXcxKXWU0BHlN9N3M1SKwmyMJHb6P9HNWDrifwDA3gcLcQy
E0iL49bPVtU+MMfMljBIuqEICK5ygP7ZTxb8YCZ/Qb2P8fYDEUgvr/5mkx9ulhk94a2ad4UCNulh
+MAJNCa0dZG98Osdznq3VRkoUwqXJGV5o+5RG2DUqjG+QR6HW9G51rBtrR5qs0/hhPP33onqSEkZ
Fa4qouz/0mqjJxWhSydyJ/u7gf6Lchzt1UsrKiJUmTvpnWMOy+HIkoq64W7+AtSW9BAdj0HWgGzL
HAaGN7dwzBMZ8d6254amJ92giLyPb0E5Jy4eo6oatJj3fzPqIlhHCW3MuvBRaoWwUgrTRbp8tYIx
wGnZRrvzRXmRFgswLNckOHvE0a4OddNQdhBgi+D7/l8pitv4vPPU3KkMRWuGNAWmGYZWHFM0wZHz
eYGXZKArcXsIDmsP03UVNoV5IDcYZr/Rax6yrExrjy3vVSQojdIUfo8RbjJTW4ngsmxO+jtTgw4e
voSPAAImCE73FXpzWnaPxFrd7RGJ3u7VDotffVNoV9m0jyiQ71CsqSZ4z1/8d5gMBw3ZgCjasFlv
aqtByh01IRvrQTgfhKrpC/TZ6xOzOfBwE4daBVXIGI0r6uqSvkhstDH5zACvK94sOUxLxR2xSvXa
EaO+l7WFjGR0sC/Ph9HvHh8EpicLNhYPNBDAfYYbPv0oqFiqF38eBQNkiweblT8lgVrr++prZBwO
sLZZHrZfr7H4wRZp4BIX204hzEzPJauXsCY/aDgk97Ck1IrYSxCr9z5u96kpHPjhbrZn3yANaQe0
Y1+dz9lf9l+Zy2k5zHs5y7nVlULFGWarj0hw3M8LIx/sxiIrn5F9ger8ijXWKgUSsFYfbVnRgtlQ
Uhys+8GuFiHzp2BhDP1VsOMVyMu+VZFCqkC238vcHnipy+PPgNyjhefHbSaQHWrtcnUs7Q/ld5Du
HHF1Th9fUegXzmlGIB1s/lmGUJ49bqN3wJFO4w9027G7a4oxAbUPHRsgh3Hln4SuWlKl44Di9VgV
tvNkbTqfVlfvKvY6vTyeqMvx9PCHH0TkmJWnsKNFaXMZpXxrFEqrKykvyF0n8YpNbtDsxBjxZ3AD
eO/lqvLtNHFFMxymsS4iPnhzFWBNTXYM2YuxF9YNmPEC8LPukKvsCr1M9D5tsjZxyxulfjM5Gp5f
f7o0zT+Noo/RfIuOok1CvjoCisSiomRHzleM0qsEqprMcOMhem1TwoWsNGZdu8Fzd7Xvy/h14CY6
uLp/EYfijI9K8PA5B5pwgBxPpWMNb553uUbeDd2YF48ZtLvfG3SS4HBhh6ZIKJPdG1TR+Qi1KIUv
2atNucZiFw4/sXVT5dlijbNShPCialO35OAn8y/hgpAPJ/Yb0Sz2NVMPzSHSJNpz6WIcKkOseemM
uAghJRr8WT0/Dub8ZyshlqOn9YSFCRlONnl6x+9ovXs7Cr9tIJ1x/vUOnJU3PfdMlCJ25FCfvepK
avHJk3Fm0ZEX8xbOPmgXOF1qu314S5R50Sb0lIVfpv4NjIgbKVOuN2BMdqqOa4XP30SH6NWbUEcG
DVEfwQeuHSB6jcbR7awu3RYmdZ+HdkuGlTqhrJ6FQL4kkI0Yqr2SMQRYhjanKneCO5MmLXsn2qkK
MsHl+oXWMPFcOXRyP50qQ51KbfSh1Tuoh1L+R0VPgbXtV8J0OhpzzXydBSSqm7i4k62WT0zwUaX7
3gWZ0QjZmWOHtTaAHcdKJQfpcuso4pEHY3WVkheKC27qjpj9r7JKShF2hh8fBYwO2qDDwTXQc3rb
HjtllerT3HisTlFLUKgcG+jCWDr/v7orQ0ON0CW7jMQ0jkI8GY6t/+Ip9PwK7ilCfEzLQqFBQKIg
/E22fq/YuYG+BUbac0olVgZjmEV5lzyq7ebTAlJRCzhspQyvgTJwTSPGIbbifVyc/dHrX2uzD7zI
bAZaQNnDZqKVf2Mo/E667Mr5xEw64gio/3iVcaD48YEe4OVs8zMBHUn2IXsWaPd6SY4XAkD1GQ4X
/04BVuZkaqlfBmtse90j7rh49EaOQkbnGJZnT51ASXpIzGKWW5Xol1Ym07uQmdeV/5FOb8aqqm+L
gbz1NK/V5xEVJYb3VFLPYWGo9+ac8jALsnnJuByud0WP/Mayfb7h36X02ZJ8dYVwZgPAUstt9tUh
9c4fqIZ66JMUfB36gBSmSAXs7WfnjZ8bbElta439C1oiCOq4pTmhQF4aeF8ytgcqQiYnt+NXZArU
mA6ygcn6U5O98U9UHgOxLypAcsfhWnat+uvWRbPZ8Fj4qF//Tglgc84U8/xhJr0dAQh0mAtnFOTD
ORmxPV1Ke6VhrtKSQ8c1roieIHHT1QL0PjA+LbzK4D1IjFQMdC5uYjfwd05HOiVZI0XTggVCizCZ
AlZ0ci/9GzJEau3xC1KQHVaJOusAyjcA1IdJk+LLRfrVXz43bxog3wQd2Kbw8GRohNzaRkiLBE5g
YXQi4e9K4/tvsDQ3xEt7aewQZUGhW3gQr8F9t0xeqieoPk0IKTAjMk3HOtT4YCP5RwAt13BOQdq7
yYm/f1h6+DLyA2Oy3CzHVjazJ+zP8K/rbpafEYxwdAJ+iFP0m0EQJ5DY5/7ncnOoNYCHLBlBvYZ5
Wcc5i6GQcxawZPYXR1QnH/l/0y8nxCPCtqAaenJrxPyb1biwST5wniVWnyBoQWwFckIpt/H/yUUS
d8LNPLXj7dsSlMezlCgwgIH8Dx4AOKBtcIVQvDF4QU4gz94eIvtI/fPFC0jhljWYz+Nl+zYBHjcB
Ou+GIhR5C7ceECEPAhTlkrRtv0At+aNJhU5TRLIERumCle4ypBgg/AhQcUFxk9BrIOJn1zeDDMQD
RiHOmtw0/KCu49xPNolC/9h2gd43sRclPXNLGc7TSu0AtullkPj6m9OPPsteqys3KB+EpEao5+vN
acFWXTdpfNmZCnPcAAtnOG+h+iWmaikjwAGd6GxIQSxsFBM+V3SuciiquVI0gYN1CygdOQAs1Wut
b2nIXlajlZBgktLmJ1Q/vSwg+iH7sPGWKGHIPv+yOFV/0VN/JgtPXD9V8jzjCAS82t4U3ZD5TOYJ
fKGOlwHmATJwQMaSzSWcOX10LjHd2pa6Og2Wjk3i+cVr5YrLdUe/U13tgf72K3qeL1VhKftGW+yr
hZlYsEzKMPz/qX2LL1r0soPhvEynwHWRxFbTkZ822RJtVRYWllhs7RH4zLMvc4NFNN0A4IL7uoRo
ajtSNJzgaSkGty2AqKIbcAwX0pokgVUp6gG9prRXRRI3z2h4KZ4E3bNCI6RARVExVmAQ5YFlGrZz
QC0OQSZ3lTNH3qwtlXwUElsz6JFwU9EQZW5F/iFAE9zkcVzLeoBUDjEDBkNm2ce7sqneUeyB31w8
8miMtL9Z4VORn3KRTcUCp49BTAXCPOXaCpdT0+8Cpf2JwIl7Gs6rjSgrmfOHydYUlWJFOr/luG+S
V0YFjNe9Ce3KOzCsEIlrDWMaTTWADMnIiqnMGZaXHEDnPD6DE2QPKBXuBcaurNx2/RNWAPFA/b74
lnwmoxBzV8M+OTiXbYd1BJopPQFMFIjKNxTVmKRkfvFxVoRxeiXadRdqezxx6sjDd4hiF4W6+NJN
3PzhKpYGJt4KrLrNJDyRllipYni4h54rkdZ1pgh08wvRch2iFjIM15OZOdTFhJmjfS2Kq/FnSs81
dPQEyqRsw6+a4nlIW4pJLW9pheb54GjYKDGh+Xhds6MlEqDiWSWlxIuAxodCMEipAW4jLnzokYgT
Dh1OVUZ3Avk3cKe43xeH3xsj3Hho2NMHrGIayNc2/674seXGDCFJlidOoG0gMWUCgXIIwQYYBfFN
RLreMw50AwW3m/u2aN9uYcPH+Com/5tPadDp9rodHAeSJwIMezununO0oVexwoZrw20sfyRN8EvM
ytdZ9beXuBkzT5JLDHjZS7xigZP+DOOh29wHc7ewXwOU6WnMX4Cp2oe18UTv2ZWOjleFAzsvrg9M
sIFzfTR31vYBJwNJavghAmVVdR3MyD5hpdIlYXXQ7y7E5a5He7ZV8fnznJXhpbnSNol8PGkNg0+1
swICR7HklXQpZ8yt/OsNy8/wdqF8mJlStGxaEKgupX2cRZc6YbqnPYrF1DkqSXkX9QG6hU5CfF/i
PF3fuYpfIyCbvc0NvuXYqxZtUjbrLMKbi8o8fNW63XCGoEH72mfBgBtL2CyG2gy3D1g6YtdCZgG7
lW+AU34+AlhV46iXPvzR9G4EJsojdckiDf1WbBzM7seibC/nmJOMPGy2haDLHQzCr2I5fL4YZ2Te
0NRJA2F7aySZgfQ+4bRRuItvRbuoGa+YZRwcieXziSn3GLErokMZHSfYEJwMsGTLkRHgGfY5asUt
IZkKDUUCB5GVA2awJ3kfxy0NOBdt5IXJOu+YzKkx3UTT1iIr68YUMv+WCEAIzh59+sqQDfZmhDCt
K2DQGoBzmIhExSyKlU5UI6I6yV4i/BgWLRPwSy3YIsmC4ZT0fj8CG9X+QefQnZXbtotxMkTiuov4
GOtvmzo7NAWAdhP5ZpGyRroJoujOUN5Dm3qAR39tvNOyIKyOlRyoN1TK6okvsqMInX2pLxF163wq
yzW+dfFm21yG7alLVz2BhKJgkSR2NTtcxMdVA0vo1/D8FVboasQsSe1EFgXi3FKdzqNGOC3Gvziu
YwqrHmm6VB2YakMRL49RKg82oZFSXdjgTb9N1PXwfsbTADBejhpC2VvSEiWiDQI+UB09bczZLCyg
BLNZONs8xAepeHqmhjTaTfH+OU9MxTcCqy/Kg0Dz83IB4CY519yWx5YVoaWTIBzaBf6KyvHWHrbr
sjevMij26yCIxbggSBwskT3XGlt/fAhDihSx2B3GMDD6U7L0MbTOQV6UQsnycFv485zqVzex8PSU
a4YGoc0dEiEb8FsGDT+P5mAbfAneKyRlps7qexpBLIQbTF73cQM4Lp3wEsSJRrTktJ++iveX+3G7
gcqn/lg2iSWmI5U6HvEuOGWw8+H+gG6xNGK2NqNp8ewJBgmSDDRsmelVULPw5g9ASF3KabIHkpne
dsz0HUg6a+iBnX1/scIJZtnwUInvA1ZmKb4Xn7VW3dvjEG4PRpqnVrqeG+IOKCQykEQJIP5pN094
iI4hjYPLAQawrBWQrLj5bu7I0x+yy321LvAV58c6mpTI9JsjZjfJurmyR9FCkzdRCOF3oPcWqHiz
hoq9L9YdORJsZqiK9hMwEAtrTAXjmr4JQJaz4MO40Osoj55Ps3/2joZpWa8rjn6mPEjJfI2ezSL7
9fanKSXe/+ODGsxz/cQdvs8sLnO6qCE7usAMAr0JF/RidNou9dgPmdu5b2URpW/8tV9UxOvAx7v8
cl3ItFzbEXuFfTzBtKGNmGyY2gcUnG1PJUuzK4CFzzecs302FPQCH6vOb3T9Dc5A7241XJzVRQ+z
cMPecuYgb3/Oo4mtG0daAUD8UQw4oKo47XIf60HanWVwFmixPZHesWLxqjLbFUwg3AwbJuOp62cx
CEtfW9Vt3wNujVgyt7G85eZ2Xpv/h8t3hRefbKdKcOdR3qdq1IM9+GF3f52D//E931we1hAePJ6G
6DOpnGUxb80h5YhESdOxPU0R7O6i86EZTmg+K705LOy3Upie+5HC5ISXMQg3EBoqELsXW9DmPsYW
9BBThUT4D2/3tjI0BvnSjlPqqnHavrmYxdX3il76CcWamaeaX0kA/KpUnRI09OOXz4v/AktDN+te
0UVZQB2d6/OMrSUkfhK+Z+7ASRoT1PBslZca12pynwVLuOvG50duaAtnOGlfSjG4lE4/XQqLZISy
XGsv+vHX8Oo0WoW2FCeA+S+g8PFpdjfnvN988A9c0jqPs2eVb7NhsKcp63fGswCHKlqKiVS3mQKL
WoAp6SYmllgmPt9D40OH2jTIstYG2/z12CJE+2BVCnAllbh+YRhRnGq58hX8TSq8tpQ1M1ICMYwd
sICjg+c4ipWe1z/YwueXzkd5lCPlQQog2VjmZKL+i7Z5qd/liAHxhapTurz564Vxueiy9QuaIpM/
qjiiXUNx+C35qCTSk+tJfVHz0DtYzO+fNjLx5+tGuxUrq5H5RvCFfNLiLGCW3gQM4ZFGfWVdI6gp
pxsHq2LY2u37busTBWaSHt4NzANLc7/ILBuj6b2W0EqADKcfFQVqag5HhI+Xe4oiMtCsIRjZ518n
bX6ZiplrjrS0aTiBwCX9ba2LXaIlEKUKuTS3QV9IXZ0/QU9S1duVVqNZ8Y9porp6qnEsj/ddHpm3
4ayHcPuKmFWW/matiDwsi8FdWk24x+QwXxWkmf+cnE/+WgCPmMiG0+rNhVpM0OfX6KDnxKbh0gvs
iWEv9AZsRw3cWwsua8WxAKcznXhJcqY8IYTB1b6wizl5DUQ8K4s9dYhsagScp85qR5CNt0w71ia0
AbORbF1nb1g1cDDlEJQ52+j1dDxx3ZyLEzHZBwq6ZiEIaiYEi48MSpQOEe85M3OZyuz10YTIUAKI
zWKyAK3Fo22UbZYP25k29b80QFYiK8rnoZb0REUHyR0EFsaZmsUjDpUDAIpgZACdf9Ml1eo4X69Z
/lQc/7XMuVPgxO9Y6Afu0beZmY4+l3Sk26RyJ0Yi3164HLoaD178Imt7XwVWfFYOjnElIhUPNFTn
e50EBg1WmJ0BUFmdRUJnhVOXr7gY/IqLNExlI2+foz7gTRBiJPc69MzFCj7orARZh63SlXv+j5Sc
j4DcAZdkLrFoBFbb3TK/dQyfr3syjwLROw5OqXsXCRbiuo2sowArqZe5VeuJeD/S+b475+74tdqp
6AA0ge+o8FKBqfdjf/ZCkldcBEFWJKG23WlGg4sfKNx/mLH5yQlz5P88qEyt10KinI1LI84Lu1Bo
SOQAyt3q/2CkhcVb8x0sOqbKI33qiM+GK6wFAh63EG8L1QMR/1sH6AcP5xArmTR12smUTg4qA2F4
/8q56fXUMmJJ6xcmFWmfUAm9s+K/MPdtK/Q2CkY2FlCRbkusmDZfVi8RQFtV3I1eO6n7xgJtDYeU
IR9BGPTdeQAzX23B2ADXki0dIefNYjQT5F/nomEIYP4Iw/4WfawleUBw15i3KT8dn7K/TRupHTJM
l2DKGhPa0SKamxfBNPD4BRV/iU63pMfQvTxldwR4AjxZ22Otvui6sPlefVPyKVxWPJLqlRwZRm8s
116snZ1QSVNv3AlLYmBJ98ZqIfbiuAwVk5ULZxLvxRYNR6OfsV8TqmEebWQNHhtNc08e3vOhFjNW
lcDbpvpWmiu3sZqLGeK7mdWPcQrwHpoTao3v0o86ZZHW7HHFZiDiMWcEdhRX+11YnW8XPsdbrkdC
sadU6y1mvw2kKP0X/4R3/nssi3TCxQcf8HRe8gpejt3KYN4p4w4m6PJjRQGQvptWLqrmR6uAwDyH
f/Do0v5VB3qFR0c0VVQ56+MXzdyG3YsN3hBtnU5lQioVfeRs7+mjpx5B9pwi0ACdU4LHLOhvT+SU
yCHypVR25vICPz1CWEDB+k8GnZSVLEgP6XVfc1ew16CTTtyoHXZ9SAlxQGmls2Oe0JhyUQ60Z8TK
8yrFOmkBY/E7WNJjFjH5aB0H1Rp04NDEdB5x3ST4ye+aAcIU8EJHSNJ3WDQ5nhPi9vszCxky/7jg
/qcJGCYZeznGwYgsTFD8SWJcvYVk51cxwpoH4ZXjz+sax8BLpq/6aA+WSha0JeSfhZtSP6WHyBCN
KYmJ7RphNY359Dzdp+uRqtCGeMJOKBoai+2JJw/QCQZ27qJhNjxSvg1EVk0bYPpirT0kTUoIIr0Q
othyBL5c9YN5B68vaqEOhX/rWa2bV1oxJIPHlFuJazYzDx8zm/VcFZqU30UbPzYYB9mX9Spdnhrl
bLD2oURjIlKmm/R59Eo3lQKSpQyynX9czARa4hF6sFNe/7xW4aOoDdePj05Ot40wljbP9p406Fv6
Dc9QzbXik11Tn/dN4yDooQwuAiTqYtpvOI9EMcQf9qCUXL5mhZTbuziaNeOrVwxRrqNVQudK+n+7
mGX3lUETUGzAAxAgoF8qwXJE4yBzPi81/HRKhjedXcXrM1umQJ3N+q+2FetGq4qOYMXOQKqQLOrx
1Q3ECr1n5KBrjHogH1mswZeEEFEHxIM09d+PoqWaFiV9dg5Yad0yn2cZ0EUJIV49l8LKEdlax3gQ
bKXCYYAhX6vp7kfGi5xPJAXLSDEOUfdgU2xFZDil8kuJ+UocFi4QOCN9rf1WrDxTrvdWe6BeRlAo
9GETfW+oUljoduRKfyKZID8mCmeKTgns4lBEOBXLYCCL/Jx13fXy5nUyHgvjeRxM7z8tgs5hI1QW
XifzT/No1EN5daD2LxXoEvTHEb8lmuBtqCsdvQITQJb1XiDxQRr2T7RI35FlfhSciKUcY+BrZDfR
Pp7rjcQ2dpikTZ6EFjgtNRAPxqQt6A6bgxzkIddja5prx9PPWfG3x+Us2PI02XziTjgrGiNiDRGS
9XGv9f5xhlRAQnAACI/F1nPoe2fnDhtp1mEKBCZCtRw4Be7k7DaEmvD1l0uVPW2y/yJWojOvxLtJ
AUfz12B3m/Tu8sPFbkR564R6DSW8U93lO7VyZVJid3nSRf59y2j6q30X8DL5F0gchEy0aPjNfgHq
qjGuckhJXf+y2x5z7QyCdIIqj7Q3zwBj1fqZ61TFyM96S1RErJapFNb5fKTF9s/jIKLQDrDUZSOV
BD9cWYeY2Xe71j8tOhnOszGCcS+e4raSKDzimno2dbm2cdPRA6j76Ni87p3S6vJFHtDUHBR1uFjM
HqYGmgrGq9HgH25PJNdUT/xSRsZs7oL60LG18or7HU30wFTvUujsKy+TJCAI0e2YK4SSUWHUEAe9
Rnz6cCcWits+SWL8JSSCcBvW1nW1E4GGXwVWgzUiMRvuGbnf4HBUixojD2ENbWZvxM1VJjv5GF8A
b40rCijddmGzvl/jtHSwV05cnbJ53oyxs3h3cZ1cmk0MR3HiuvDI+CdOu1K/rDswhze6p4iOtR4G
cNrDRn2McilyF1Cc1EkEEaKPaErXQnkjxit+8Foug9t5IL+2CrJqz/eaRvK1h9shcMN3fhQJSqG6
THbqXdVDNGP6m9Sze/NgBZ2I6kyOLvfnv1FBjvCxDsNIX9ZQ6sglrLsjUI9eogIsYrPmPp+oO5YY
xbUeSJVNovyUpDH/uGKgAL3SbMnXfOMBvMa2s2XQmgNXz0XjZiJB2bSr9ny0DY1xx1PlQ16C+m6L
8eJV+OFfeic13F+Aye6cW/Ee2wVsqExC/nYRujNALSli5w1Ka1TW0C4qp/A9X112N3ekQ1MpiSkG
dqB5b1AjVAev3os+rbKxiXltlhapkAxfnNlyU1uaSlKXypPVXvScCvXaP3Z1bCNXtwl9tTTtOErg
aWKZg/LYGL6oD8sym3hVJb+lOo2FZiyFrz92wClwaRu9HMGpiESx41ngNZJDaKixjx6c1Uccr0i3
O0hzT6dbsR/OInFMYvitXjCNUf8yAD7QMK9/ydxi4sT2jb2NotQUanNiG1Pr6gEbj3WMvqn8EmHV
hl6ZG1zyYBrA8aO5xxzeu5PwhLnBcD+XedIljc1oxYFxuTZ+nKip3BrDn0YcNh3hiHIhpHrTYhqM
VWKbC6Ow4z6dk5zA9SCgePc76Z6VPDwlTKOtmNI+75IX2FEyYww66tefBNpjJGUBguSjqo/+mh9c
/hUr8gYyxH0L4Ey/3R3QtxQatLM7QKEkz2fLLV20t/c5h9GYfkPEJplW5B/VUULg1CcMfBaa2/6D
XeU2/KvEplqIKXB31TYmEo9JCzHLojQlpTpyvi9MNaOpPwnI/K4/nY4OL8PLN4o8U1Hr40nWNlvF
Zy9ozleJgN6I1T9eDGXCNmZRRJFJwtcpryhuhHIisIs+orYYaQsGeZhokNGbXXtChiLxH8Htj4m0
YH8d5RQKP+z0Ec4pK1m5IQBbLV8WR177dzdIvgCbat46YUq6oI/itV03K46RmirHr+m/HxOweds4
mt65BfkaqMrRsQTwTrCnVhFGZkVa1FRbDns4CC/q2MvI0y/DAPl/pet1t3SHc3CvWijp14SLyrUj
8Ksd8szxad5njVTaW/kF/cRL7dtrJfEgNjvFtEcw7ItqXkFQnyXU+BH9Ww4I+k2YdMZE+qCxwQ5D
baD9eCii3qFrzdrPcbXfgDTCxO0yi9X8TO3DNxV0Qiu+0gDvu5zuVKT79VForOkq1m1CTqWUvaHP
z0U7u1KqXsSaeHWd3/Ad/QISdbCztgmgYf17mo1EUVGqjuxDzSVHQH7VLFUrZCcoLjFg42GR0rs6
MI0RDvOH6qsxNzLdCR6c1yfxBxx5wB6EHaX1y8//al+ey6CDMaRXmlaLwj9LGOz2Q/J4FNqYMzti
+Oa0uegxtKwhCAQnJDicuV1uKEtIkqX5Ei7Dsk64URsRxmwA92+NERWJWUSF94S5OvG9aD1ZzLKy
4UjoV6Irp/1aG8Edmb/xZquu3FOZINgUREEDMDgwyug40cPs9aIhmTkTcfE0E1iXqApfVwjitVIR
eEZrRNiXQaPZsY/tAcROHOiJ84fFWEBxalVCXkirPp0pCQC4I/03ssqKTKsFloxRs+ZM6IRSmWSr
F/sSAqBLyrDwCpnJa8j1xuL6HaiwFTuJCsqLNZxgN8Ew0BrEyV6Y8CpD0P32cz0NNfZZH2EjeXww
31ju64SXYzhzUJhgEPMEZgdmUgdWoN40MBd4QIFLQnMIGDnGkPzf+4gWFvW0ovgnx23dGqghN3+1
eviENduJgLh64kGy6TjtgCw9fQ4aUTqzRZ7ILu1Xe5g2b2+eFIgdxVhz0uPIfAXkCn1BzA0tcYZI
LPPpBQcbPEJtce4NKk7IA44bSYQsKHZxKyopwjfiRiB7lfP+w27mLgCScZG5wsMmc3L2o2jBm51P
UHhOHqDPRGYnoTj2fFqOgws2kviQyLlaA4hkSNq0hHPDrvj0lx6fRr8HXUcXliXoMMx5LXKW7yQ/
IXSW8neX7yrssc4CDPw4FdjZif4LQsXTwrEbyuygCP0HsQ5YMsVro9ckfWtLfLqOvAf2m+hNb2Tz
Tr1YaHW8eEc5VUqQIXX8RGWtAKXJNkA6u37V7zgKVv8OG5KEyO0BbStW7lIaDmu8VErKBGSEwG/c
t+1qcuAe9AZmXg/r8XMdiAr4dirSDPSlHjaZilxGkrD/Z72YOoNFBEreFEuS/54yu466GO4GQci6
dc+RgBvxc3YShhYmoG2REwcszTBf3xjBpzG5mhu+D5MQXrF++Ah/XmlsFITxcQS/2TDUL2r0eW3x
rysvevz221w+se83GrtReGHf5BYVdYHRj01EUbg8x+/ZJMTtUfdGE8vtUfRbVubL1f4dTgX1TLsD
7ZhjUf2Kv8582AP8G193eW3GluuM8byr4liaa+VRvDMic3frP5w5hVRuBtvmyglZ3aVF00GNlXqR
w1cXIe0GFCbAo2cL7JK/nASmhxjERiSlU6ZGgoZfPwalbzaUob6ZYUDeL9KIUlmsOMZSm6s+ARSp
2TTbU8yZsy81q+SFrxBLTy7LFJJ/FktkoDz/lk2TsO+P1iqH/pQ8m/ka4cZgm5PvPnGxN48A35PO
lRQeg/GnICQHWxLGtwAI42j4aL3SneB5HgalagxC9zAZrDqbO/XjqUe/sMO45TWhVO7YjMj4TRE/
3OoLUK/n7oDGEq6CLh57/qq8EaabYYl1LqMYBTak/N+uHkLb4FHATe7ccWmG62Qdpuaxxme12aXy
lowQZG7eZhjk5WW+0Rb6Qd+adOzsBGFp55eH3NdDH/NiZjaA8lH1jfA55C3JddsaR0JyUmPwUgy0
kjDndrKvK5qsVnRFSBK8VCrwP9V2FUR1gY49TDtgDJIS6MKfnC1ku7Jvim9EamwnaEI+WdrLTP10
FN1Rbx+sNR4jmKGAttTqzbABs8vVRLXSYo4BUflSxp8ibfmsd3NCjJFQLIO910DHVjt0BZlGTx/k
oPxxURZwL3tXQCCbXhddyYY1e47y7Jl2nF+3GCSefCesSmKUJ86ZnaaI4WKCKcLdrZ1sjn/DNCc/
AzUbAWNCvl2zgP1GtbZobNNZr1xna9U/faQ4gwQC0NiltJOF12Uo7RRCzSqltSA0ua5fh13hCg7N
Ag9i8JlRpOsYYytMlkCtsMjuDL/CAR0bkLMGijIRQmbHw4Lf8MBMX82VlkrkGrk1wOna5Vg1H4mA
Pbaf23k3N4oTQVfTB7OMbXIhPdzutZ3uq1bq5kzxyIoRTcMkPIVICUrNH2Z21rwfUzuD0skQwZg4
BDD9L+vUbkC+rN0zqNiGqFdIr8RkPGZVPyZhHnKaafwNA1yynJPCYkiF9pNT9IagnptyQI3t4kp8
JWx+SiI9sRv5WtzlHLgWWTvxMvkN8a2V7xoRoFP9YwCLcSz9kLiXez42lP/Imz0t3O6wrmA/kvjU
r6ieNJGSfbw+OWv0mBllbCEO0SgeZ7q1fzL98lEc6xADQVW1IMDz9ujmoQ49dO3NzJWGxeiU7SkT
mck/+vqmeEaoF+aO9dX9UMmNCoUeETHVCCTtzrbJfyFpaV8V+95uyiEsBudqErxaUQyGSnVbZINu
rVOKWRv7eCh0CEiozNZGEpYnyw4vrhAWheCLtQANLMTnn2jRYzoyc0oLIY86SICftTrCMShwi0c0
uEHFN1ONZ9O8E+56aoICym3MtOxuxj6SujMRjw35kM6fQiJj7NhA8V0OJQkSPmyGqoYyOXaJQlsN
CHb9AJD/UUBrQAabfizHF29DVQjvEbtvkLxNv4iFMlhLRzEhysXnAyUkNP+T9TACmB/Vs3h6Kh6X
XjFYz3SkEOt6nLL1DS9GODsQUqvs3LMRy5WaDc6zxsl9pb8LLDoJ92ciRTalyb7gnIZs9ELDirMd
vMnSgtKD8x/QsmfxPJk1VSJ2c7ZRyMt95GmajaTVIT0ePFYrEBfaXjOE90tzkMAf3AgHZ0EZexNH
SACsR/xUZESOZv6d6CBa4MQOnD5bXzMzERtpWg5BIdYMrA/D4KIHE6Hxh+G94zHOXMyrghU5HRrj
eXF6hf9Bmw++1jWbf9QOpvVNEa3sTcViRBLX5JXmF/Jut+fRnV2iXwFaz3XbqagqEE9Mb1nU7AOX
qBiePEYt7bwKlcBSTAxCDe/WXzzCLB0QBT/N5XVUlueHFiM9MV5eS4d+ImHhsBdaUKOcjRquT6C7
pcVfQ5Er+MOmtPGbi4Tu7ns+aeJ0ZFevS517jbGR+x2FLwtKNtPdSty0PYSXUa0h+xoeEK3u/LJk
97LBlKC4MDXe7oHjsRFyzFKsLmPEvo/JTh1RCspZH96N3qOvQ3/b210OiSUlYRRU5s77Mn1Rwg9+
aDHhQ9NwdtdRKSJq+pEoh0eTpoFoMuhG/qxfPV3yHr0pZeVZFZJDlmqgENmqihYXqqdljdFw36Mx
sZdFbgRRoEgFZgUMll8YaRupObfEXsyqU32jsWuLO+fN0QL19fKFimCMl7FxbWm4KkvYMqWTECnt
/DHQEJa320DM1VtD1ihbpbaNU2ecPX8suZ5+Zk7V1dIhiuBL6vwmsK8Hww0af4nuqSql3f6NbJaK
+MG9/f1jPiRtCcuPPfDVUO5Ewz0YuAhLvrczfqvVe/Ulj6ZDho+JGPSNqF1PhH/+2V305GF9/kzi
4t7qEBMSXvlnOhXZOLFNq8j063RThiAiOk/ITA81TNze6bqwn3lvTa04zHfwM7O/CrvU8ZI9moAg
9jrC/zGnErVTB61W5onKRBjnsP3booiigTql4rtoNQubh/eH9tS87P2FyAvVsRA1iaXF5pBwdaER
zLX83e0U9bL9Ffd/U1bF0qbywvgPXwaL7rImW/0s/CKrgT26DngiNyCzAz9Vk4qg/XdprJLO19ff
v3sTewMQ6sba3/LqPm9URIZG3Wx8vu9bmWuL7mhFbbFmV0lMhIh7dMZxxlw8dA/XIyElYkYTJYMg
06hTsRzwG1+4/mMG8H7K7+rfr2m5hFKcnZLKg+4TtsuEYsSLj8RZzbGLJgX7wJsN/jd4yjSkm7YH
OXZweNl+Jv43506iuaZ7AN51sBNyGDvAWLcrfihPHMpQwxYtnmtLYk3NmkwKMJiZPT11Hwb3gPQU
161sSMMqPubdmIrYhC6EeRyp2KiMAfMtUaDAmWqjhe4BCuEsx3uSrTkvQnMWPc8L9Kfji1yNCJyE
H6voef0CVq1b7ZLEL34sqRA23cKRjdc2C/u3CiK92nxpQpqFn4fZ3ZgKaWfNWBV4x2D2bRUwx4E5
h7dtONfXLDv1n1A7DJ8FYfvjZ93rHXrkyUrc8VYfOyMJGGcRvcUXJZ5lCmRiwoP/Efa6lkqpzU+s
Mb/qf/kHi4erufSoUGD5y72bnLOMbenyG5FXRpwQQs/J1t4hbob51rPiCh3V/O9VTJDzjBP6kyIn
f7VzvGuPr2AW5YnLuhutlEDJgVT+yJI9hRttWsQB+qUjRRN+MJr9pl4Fj2FJKl9nJlwZnNli9vL0
OjFag0LphObodV/i7NxtcwLqVaA6l5DebgCK/dA+Lts8Of7gn0B3jTLwkPomdXXKbKRy9NEzieOf
CH2O0HjNeJ8p/CQwt0HioOHIKEkhiboMoJ+cGgOp6fec2VYvtVkica9BM5j1ywTZhH5M7vipgKig
25fjiqRzZ4xBnuV1ECDvUNmkK3um42t7tntUcwzcSoCcU7a2ZGBSbjkLBpOZHChpwHVq1dm0ell7
BKFK7RPshGopHi6n8j73aJAS50ADaSk8yvb4CTtRadVQp2sYvT+SghYsigikEs7E1tbXc6fRWwBM
gZCpIkfvhsy7IVa/0FRt9oqeAFmi1ggs24G8mQFpqi2F2it+DpH2mTVVjU9CzqXfZpx3gmU015tr
2NnHW3+lvfuWK+cASwuMOdXQVWcUp97B3fOV96nYDEqpXUPIeF0oGqZ1flm7Es0gNPKi14UuXZmt
J87j8ZxOXKYGFweXkogZlcTO5sXl8k9IdOYAOU8Sh5A6PL9VLFoSScxLO046ByKcrnxQNBGv+5WG
ui/NWaOLsoBWbs/tFZf5JJIsM80Swm74VmIFJD0FOB9EMWT+xz9e2ACYPpzg1iv5IrIEZNH3zAOV
izIu/SVJ+Xzj9cGx8joowFfKsRafA0eUcFu6fc+3SHsv2rUeLV3vV/6o10gOeW+zNoqNkLDMzbT2
r32oRDR8Um2T20JL/+axq08MYlCtAW+hiRicvrAQiKPMmx+sdLHMOxjOZIr4dtMLOPjIDa4Q3FkS
cIbPT9Azi6xAb65pdQ8ds+0IVO42XV4hszU4miRSzBJCcA5nENA2txkzUno5I2xyIFR7DJePTDt+
NNIXGbIXy4PdGKQkt4D7rhTSejQA1t5UHcc2D3wM1SaGqb79ER1oTi67zv48Oa+FhT/czAo0TDrt
XBeh80zhdzMdbNo0LwuVvOrkEOSfAX5abVjY48Cy8I2I2bJzO+bsalIDizrPsFniZBwlgPoCE0ho
E5TOddsODM2vG9ZCSDLGMXE73GkrnQKTnKtFY1zJhOKvltQeKh/EMvbuNVwNHjhQHTi7ui5F4i16
b0IVHNc9p5qLyzJC47kwnDheQ8U/JQg8r91ja2Lve7sYYlF/AbgiNlOGbMT/ncELHGTG/jstnK2p
zSe52rcJrDhzOKvLYAgV8duVuiLutIC6FP6Xtl9QTP30sF10ZAugt+vQyXixOBu3krQRO9MKYL3+
vppUWFl6hvmqCC8EHoOt30THCZNESo0RHTjT4GylNBA7iOpPxph/W4mLfbjVRs1pCvvlJenPPq9V
RCPAlM+IFaD0qQVwCLPujHylcpQL9eigcc3kny5h147gNpmCzaatetUHeRRcurJHjGswEA9qHLbM
y4rv7zKxGboKMuX5vRdThh2Vmoz+9jhGO/i5abNkq8A/ZY07uxmqi37OhA9UNDwZK9F6n9I4DmPc
uOCA/85ROwcYFi1Cm6yolXFqmySjGtG4ufaotewSrOVliG+3Ea6V2lRqTynbak/OmfzS5K/ykwnO
D/cNy8FYLCFH7nNEqVHKnBr7qSNa5S3G2EyIWZovhB9Mb5zgfmoC3wG78l/D45FYriJjnB/xiVKh
k7W6/+dmZpS8JyoGpqf6Yy2+CtCKBESDMUph5CSVNRBQADFV6Qxp8aFjc8rGJ8DN2vZ6g8+NFsKo
Qqt0oXZnk6uSEzl6zfWvOEKPJBTkmZfJ2izXNKx4E3tKQOVxBOzumUm9D3tSPBrZAe9vdbjmwvTx
QnPrJK/EZ/DG6gxOsqsZeViYVlZ55z+RpFQEqPWg9nHso6DD2hUGwBYCwO3IPAZHiC5bNRtU4x4C
umM7uFtmCfe5t75/rnmwAJYRL9ln55GeADTOgWJ3D/fZ8Qi7WYldteRP1s/jD5bB6ZNCV5fvEhEO
gq35lnaA7GXB4JwnYO9+1USesUpQWzPKQIEdUdBuGmVyctO2Z8Mh/51sFb28YS5Ll0XYO2eommws
f5EEUJDKwNo0atrXCzEV5LLD8FBprmlzajx5OEi5tJt3YWqFhCgKP/Hh3hAwedgVvQWiC9UrX5LN
Hp3vldZ/0uvWYggwITqQOBFnUfWmNRs8EguLaDU1OmHqCuCu51GfxZYwifZ9DiBq+NK1Gi+R7rEy
fZ93f1CT5TQAiBl9GAdv1GHK3LXq64PTxMpQ60W+C9XApRHLrk9gpDx9BYY29keQlKNcupM6/ORx
P4lOxf+PRXKny0xOTr5H34MzPoz2ZZIxjXyoagTl0JIakugsfX47HPRNxU1w+BmsThIw028WZmX+
AOB6YouEyig+l0FURio9v80C9MZPapBmWC3K+UwoQwGlkEzxRV6yX0hva3ZlRAZkskmQqbKp3iTD
i5WoDhAynFHt6GjHWtg4dUANHeEayQ5OlAPhhJJT+DYk/L4yWO6JBSUYqF0mL0Fi3fQRlVZmL8++
P90P9QqBEAnGLmV4Q0XOsAyD8HuYWO+mfUYXxVIfxfEOwTkdmBcqEUAQF3f9/tBgfyTau9my1RZ/
lJKS0njAbKBLgR5tYyydYwcfdjyrW87EfTAvW7ehBhY/6MF4QEeI/bv0D/O0Ylv6e+3R/mo3t7uO
HvXplRDItHIfUbnYR71ZJ+o1HibxyY2HRJqQamYJTez0O919Nm4P3qE88FN+XFhhsZW0pZFnyq5b
x6gFIymYIzJjY1EYfV5LAEuDbgb6YhaARVTMX3iqJNjJ110Hv/+/6/Xx+0MmGGcB9bJ88q5xut0Y
jrxVBFoHP5r6waJ1zRU1NbDDTjKd+6rcMFIZEsRfW5zf/wccJJnZhPXmzMigd9NFkwW5M7MtXi55
kkoDeqo9rIdsnBpJeB72zbibS5fXbvTAb9l0DTA68JcP3DZLsCbsc3+cZZFR/ZHS2EWqA9GmChCy
AYbRoIziuOFhIS6BsMf88JIsBrcuJVP1/aP4iOTLoVqnAfJEQtYbCqpgpq5bY+dwIx0trH+6NBv+
PcUhSJ1X2uRLi+8BJqtXMn1Gc4T+ICZUk5QCjXf00sSFAjE+7ztZwmuHxCRm6zJoNENVujGTfWzN
Zsta4M8INCvLk40ATahf2vKr2Z1dYV67xFPwp692lwlpszkIQneSHkqX3609rEqPabLOlNfCwSaT
0jrQCFpCIJ/JxPOSaKdWBstgwfASdmhbmqeerNjJ4mkm6p22FLvFC/07z/qv2ztIOXB54ITzF0Gi
Tnj/+YM+ftwd1IfBX+jbQ7RclU3GgSd56dBziJtIt7sqFldzlh9yQySizKeS9+aWWNjrBCL+FLlS
W0oU1b6RYYcKDpRqV00WBA+bav0/Vra/2O8QFVnqX+CH//LLwvvEKN3blUQb4wlnQ5nxprj0soGS
o6RsdRijApgxeu6p7dU9ybz8QQPvqEH2+DCVsD8MH2ceL4Ki4oxT3NVfNYR7hZFmVJgQ1Srny8pC
p2L2IAoFg9YwV+rPD8DtNAvbNekv1Z7VRXKoJilwk+th6oLyvk2XnUz7CW3iidW23BeIMnBPU7Fb
lB1m+2F4JDEcKHYwGlfL84bo/wlBYgNbQnFo7O6sB55ja9OVE2i6Vr4RcDBMo2QfE5MifRPVxrTJ
vl4bBaQy7Nuk0s/rTOUwfy1RsHxj4WE8Ng2r+ef/wDENBHmHnct0kGh/Hpqy/Fwt6PvqioC+xNO/
1MReF2Gp31t1iHieIzXu3vljLM7eWznvkBthmufvcOdC/EjFTL7L97hdqNQGqFdSUjG3mxwQvDvc
KpJAXWVvcIIgxt5LLK01DKgL8D62lZnGZIbVBdRyd8HSgkFX+SdcVEaN7YYL3jgeNOvQTGfFOvpL
xCJ3s9wtEhDlL0i+GoSvUo03IPDqJ3oLsc9eGteTE4ObIBFxJ+ZOoxNGxn8cGmLoA1xnbX5mFZco
lMGbM/c1I1KxU5G8vOHejEIMmGEaevgBwm9TDAp+gftqG8/OE446dvNsyI64G6B+nlrAT0HSWFR0
lG4A9vRE25ZgYoJA1GMy19H3s7vzTCG5c+fcAsJxKa/LwfmAVGODh1fsNutJCGL+KumpMIjIYc0A
e7xKNbAeL3pc4p/tU8JsUmFSzE1nk2Idcz+ZXCO/nv2cWSDo2s6hLceBgqthoXhjOIRW506QShb4
O9r8TTHCX72AnNscfRRJipxUq9kaQR/ZkPGKaMFeZxZM8HGJjQSf5yvZOaiS4U0sDH5yitDXK5S7
V/91ZGqLwCaVzy3lYRxHJfTAtvovZFeCx0ryRvAXqi0+dxw9gZDn3D/ZGeEMRRCVLhyTKvAGA9H5
+HSQSmnmkvqTNWUhUTZYBMTwpA6E5/GarkZAt+VrkEbX2yxhhpbPDpPP+pSExdPbEenfK8fu3SWT
Fda/N5vOkXd+dnjIS8muq7dO1R9O7O9vqjsxL7MBnP+eKmOmK09JlwvnvAXV1lCBeHPARWOfATxh
jsAVRISWv/gktCmat63+nBXgu84+XG+D1csD0H2PZ9HLiMrbQ8m+k7BD6R/YCZ+i0kX8+oUqz9Sa
31jhiSOs72grqzTzG9fchuCD1yFetXxQF2hzqmODzonbNZwIRtMtk5XD80PDY2LgDKtNLv+d1Tkk
0mWGqFar7a/xOTvQVLUOnQSmMgWNUktDy6RyhUJnqzpZNux2bmDRIOmupZW2QHbBM3JnNU/uUxSp
IYuDv784b2+YjqW6SAJr7zLaGgt3TdhSZbZnoQCCarPhHXGaGD5gupVkoWvRJo/Mi5tbz4/zLtBx
8Vw1iDR8M78+tOu88cmf0/p+khDIGsjpOw6Yd46JmB0izGcer93GeQ7P1zx6MVSxXDvGjUponHVI
P6IDgGrn+rPTPdQWDpoHb/phQRQD7EsPYE9JDLeBVS3tbQyGKmRNeAub/xTPFlcBLFMPZ6rOXscB
4hwbUQdcb6Jr0vbL1g53qevuSKrCp8AoYCU+5g2XkJqWzNRiJ3hWJ09rs97gVd21kB/BV9jD6jPO
t6FPk/6vgOv5Nre6+isJ3lq8dW2RhSp6hhZr+jYxBnvTJAkHf+Ey672qPx3zPwkgtViuEF7mejxC
xA9JUtqkBU6pUOJRsLWRLBw2uLWhAJXbky6W0VDupDC0mDHKmh1b/Ihd6ICwrpblF2qXfZrKSHmf
qiu+ERN16MAzTHpWLKTushr2ih8S7ZFlVHDkY0X8H3aGMWs6GRALLy80dRcZ7qf9H17Bcyr3L3ic
NGNb85VIK9STQpj0heTfuXMcRMawtDQqVHOOzRAI+SnSiH9XOljb9a+1O5ZIE+Wp769yrqcf9Qss
vsKE1xnuSPTjNmbjwXRMoxbvu/kBwqxxThNPTo4e4mOf0seQDEaickmieQ5BXnrnHbx5ejUHFrr/
ns1YZPTebabwqPdDtORH0GbwjdVSoXQykL+90b6oPkMU9GiNYquOOhZhagXRkU9HzmYH1lKnR09Q
lI4AMDw+4YFN9DciVNGe+9hx9Z7cG5D071gpSOAiAUo9FloM9D39OJxsFT5fEmYLuf8slqzlE0b4
Rz1eZRq3r32bwldn5lLjFFpY0+6542s+XOV4ZorBQNdEhHgv95drhdAdcc82825vSvk1JJHlzfUK
+fEfP005qRsGsh+qn/KBRt702USNuzQezF9auTewnoV5iMVL43R4y8X/Eyv0xnvPCcLOq7YoYnm9
1cpKQ3po/0sSJbY12Des4TQLePxPuWaHiEzvVAHa6zB+37bl2tLyTmeDkrDabCecRUU0cE3hsgVt
1067SoXhby7kxhooh5BUDZ4YdCH5LTstR9ydyi5ak+y2i12pOGfyG0NTwGRb52OKiQ5wVnTxhQsH
mJdgmvEHU8v44ELn3Gf5cM12sfKDWWM+/QcA5/MznLrIiLDlr/clAAvF+rN8bGuoKtI1tCX+nWjQ
YZcxWGkwSHex1vluZtiH5mXf9CU1cBIRWmJnh4UfS73uwI5e0YMCrf5utrhIedMntONSAEq35P3g
OtOQ36ch1z8O/+jcCQbo1V9coDHYH0tquGFM3jh3PNjT6AJmw1LDHU8MIFmIBFsbpNAu9s1GM4Iy
UDcyLlmnRR8M69ekfd4HwUTlpEmPAjKMRTgHUix2884ebs59L5q1BLMEC+5GaBgCsH/pVUWPYPae
r3L64lPxTI5V8xgMOpWqVivlASzK3iJ5pJZ7JmmtB8SonXoGmTobfe06QO5qa2lH2gWGQSIteldu
d5mZu6JuNp7BsyhUxgFURVEcxZo15jgk5bRUOi0y8GnMVFaZjTg+7ddA3ny0ktMn20/9abQPLetV
lAvfyaHcuiY82X0Rj9RVlrvTke2hdi5ibhKJNxAnVbLo360lghroAnU7hFKOJHdzQiJ/BSLuK1eN
5kNsZo/xD7z2UyqbilkoYF5D+9hs4NujtSJA+xnLt8kMzDO10vBFcTeeV6dNG/oObO1AC5i71zOH
NQF7WKTcJHg8jwK6Rak/Q4H1T1pkKhlDNl/3E/nCfHRtqOOmEyQ7o0kmzEZAG0wUia4ffXAPVpD0
CvLd/f9OnNcHZSUAuw9EVBEqGlhyxX3VnUkjFkCFXK3WhdiybTUXOo+U2zOkd/W4usadR5FRQHyJ
N4d4lRQPZo1DEj/SOuf4oUDkxs5IccAVu+SVS52h2ZkXDpbyyrTXciv+rmODxCEyM7eV6EXx+hai
N4C36T7AL5raLNlrQMjPuIr4Pxfbov6pLAHvzmmNOvRNemnmU37quxxEPyYJo21bLAvo4cEKNDbe
8QbwpxMF0+QRtj/RpdtPfanrxEocdhO1HjzGCmKgCoPQak8QXYgHoV9HtL14oQtTVq3BGkfKLkgW
dfpU5mKhfHk30wwugV5BDTgBlvDeGgGluasghLVWTwIkOaIULsyZ0VvG9/+fQr6eO29X2kN54hCT
oCPdG3XvRGDp8yfh5rN54JdC5r8OjkV1iKoO7gKJq5gmM6ThQk+nC3F+e7DWaD9Gumhwx2MMrlfq
jdFNqZSHayQYQ0Yd+2fPK/O3KjHp5n+qmyLbxI50REAfQGRbla/QwOi4UoWMCjM0XUy0qMfApOdn
izwf/PlkvMEu6SpRaUnDoFUirmqoLaaFiNSzjqJ7DmjABhjiq7UhTJ+4vtciwzzWilbLkFYxLVcJ
D/OU0cdTFTQJJdOoU0CoX2AYHtaX41yzaqcEVe1YhMULzSq7e1tOsjQbBRMPraML1Ib+/6V9E/dW
578qkwIQeEdsA0+80xv26mzzoFM0pLQOUW43nyjOtYpTFwF5dCVbXbMRbqZr7mIx1GYa/geAs1jq
xcugkiiHw/cqRi+cBz7520um8hnsnrqSoa/68e7hJQujYFsFI1RDJLhZwjnjysMMvu2x1onhKE3s
nKBYDutdnhqU3IpMdJXUbEMk7SzIc7+lfwwgaETX9eXVSX9+lTNKP8OPDBhW44xGwHmRGGncuAb1
ArZKouqszhEHol7dQFXLwQl9IfyU79gqvX1sutxdPQPuzXXbmvlaSHV657Iz9rjaGrB7faSW/DG4
Nd3HrysmnfaNDuvjKD8rn5mx+SLyUYyqfXw8FADJviP++DlPBe7rFyEgl86axCA4qPWutsqpaqiR
iqq19oJgxTOA1PHxdxbE1Uqycua4GXH5Ey9xo6zsXHuQgagTQrxVm40GsbifUnreKLT320AFKBF8
QxwZQC7JQsjJLtiYSgQLvDUPOEtgmbBq+HP7hDPXbjgHERzuhFzzEzFJfA/6+ksRMfBaEzmdh2ku
WxQsg4KKt0wM2IfuY/1XP+YYRD0H+io+o0cIC8s0DRQIO7HVTmUuqL+0gGFEPfkNeQyaryhRx6ea
+TzVtkBBi7CHeILgN13tq3PYQz1h6HV+CfLiRGnvz2LjqyYxVCY9EzKIZ8xgqRJoJA6McD7jQfwR
0D3LR53sRadu+MQAq6gZ2+GbFiKC5TLLb7zSj3eddjnIHC1OLR79ZPrGZ7vd4/48NJ817Wo/v91T
rSxKBRS5Ab2Bcj5DyygzhAM2Xs0hyWZsFQN/rUkVoMcomf+KjcJUijZ3Fj2O/LVgT7+EnbBG7tGE
pcY60m5u8xYoWzaenaFA57wqL+6qXlGxHMWnxdyNhMBr63OPrliSp00RBqf0e6qqphELvLkFG149
p3674LXFj+kdDTHbzk9+gprN8nxxRvbmN9A1yC66/EHmzTfViX+Xw8Qn2w7lqaE7CrCl3dtE3eVq
bQnFxSv9VxE4I+lnKDTGh1UMtO3Gtby++nKTwE3EM+XIjM5GabNLEfIPlHm7HXNoF1DxjyNQsdml
afR5yhNbhG+3M2oHlG9L0N2mfJiPds250ctcqcJmzVpksIKQJ+p5ftJ6XrZSdgpZhlt2qX1PnMZ2
Jj8AGjIUSoLe7E1r3xtcYX5J32dvIRWpK7pnVFlauSttbjxcA4yEh15xMa74tHlhpAh9qpCPig+T
YTd46otOk9h8L+kLOxgpxDy+9blUSTtgWhb9QwewaWeibaWxPLnbK2IyU1Q+STAUQb0Cnw+GRW7O
LCCoJojaQR1dLRh+pzkq3ScQSPRLFt7zQCX9unXTm1tpAIqq8Sc/Ukh4lhzr8LRs0N+9CybF0GpE
ru6mJvFPyJeScUN9VIfEvFrlGWt21NVq9v6rmlL5DUvm11fPmlcPZP0qFukJeRRosvTonqdrXp91
I4dmpbae2Y5s6rd2SV4NuJBbhncE1UwmCbEWXR3HvQh21Voi/Da+hGegdSn/tqcAoUx/+X3l5Gzj
kpgL1LcgPqaUltIVUjEAtiNncnRDldZOX5Dyuvwk/apRKKtGRldOOLdNpQUhPvNFp2MQyoNXkwO9
ILfhv/KcaYZIH3J/N1IMWaWeBYVY324QDn3tcpOfrua8F2Zt9t+7aiBqFxk+q6naYMcjaIF7vfUw
44Mq/Q6McBkdQa8A6EAtjxn2zXo/bJPmkJmdNTwBr8o0eHBs3QxkeYWZxJDiuPbvhL/m2x4jy2PX
QFwvMflH3wOMyG7qh2GiHqRTIu8WfpM9Dlo0v8qxtKzTMXN97XFitvNsbdc1a3rHJ8OOckxuYdyC
xRVGV7AzfZd8L7YEtoWhY4/Ks+ltakzB039t8GV5LZ8md5Swae22EMsvgagvtvHqy2lqgvulv66G
AWo2TE7FcvFTu6NZnjcjKYVN0KnOyG+pxAiIvcflp+BCY94OyoqgzI0IG7fIE0ppx8lvRuh9VtfH
S2bsWVz0QgPjU+trVo/fKZ0ZwTICUaGTd7gJNSG3TQDKMErfX1k8q0C60JqzkmBnC7eLw0vienrc
CU1kZVtDlyts7nhhDkACSJZ0rTSFf1UPwqbblBT+qEGcqdtPF2sOLxajVGBXQP14uP7ayCUPT+DS
5XKmBN872dUGaZa0k5CEw6l0EpZgj8Np6U5+8rBl+T3HN8OCQDoQJRm14MXaHeRdvqbYy8VBwX0p
kRcDL8F7Xx2toodE5hzIs4P1JknQ2BIh8RxYK4nTVFqtPIYOjdwMgtkCoQkMa74+qw26d5NpC9tj
6FpsunB/U1mYmleSnJYn4VGOJJjplCi+jI7EXdk5HuuUphinxFna310H/x5fEBqynM4GgnZxzED8
+SfUOHRQmE8PpTOODxDQqXgcSJRRHKmydv1oh318tiKbt3GHzXRRxW/wtxna/r+zbS3zCcXO5GSy
O7y5DA4LUPWAomHKjHS/CnlIZNU1wAoGrSlIJVF/YupWEYr7gUGrl4wz9cWsQi/97SfEvPUGwvbG
O1n5lFCgcEzUD8h9KHako3s1vNjuPh95gxTPvh9fSF76d4bV9AdUD79jY4Qs++T+j7t1zQ9Edz7y
K18yue9d6BEaqpIx8OaxdJ9mH7RKEP78PWNVpGCJm21Jb5JG9dNppUpJfShYMwQfwBy2eMeORW9c
CPdscpbWnZwwNCAEjO37KZaPtUQThaAjJ1VuyJPCsKud6wE9cYoo6r+Egfej+VTypwztuXsgEgf1
qpmCjdCXnXmd3bthsD5PgFoC4etJ++gPhw4cOSRTYaMQatrkOpKC2Fqz5YTwIHZXA9PWt+/Y/AS3
2THvlSSilP8hLPFCSaqyAP0fkCOs5A2ibg3ZhhFbR/V4eHtFtdGZgOyAAzBkN/G9HthXnwY50sLu
M1DfNdMA6O1Dq1g4M33IADa8TS8vNHZXuAk4ZISr55xwRbQrKCUdBj5KMkPHkBXLvsVWVDJ9YcIy
sZ9+l4P6viGL6yAi1QfY+ayvwiaoLjDZ6aekP9sO4MYvqnkYcZPAM8SR3x6jZ8hTHhxKFeIjxVJS
/+h6Kq4717xNb6nUUjPNSrVK38AxNM69A7gg4kU2ZpbFmmBVAPYbEMut+Eqa0CTjvD4KBn2p3GGo
maSp429qrNoY/3euEzhe99pO+Uwf+NEtD80AukrbKC0iJVz+IWMdxgwRsqS3wRIOrIv6/lm/47w3
0cF/sZNH5CasTdv3m5nki66cchRSIq4snaKtA/6WZN925iMInWVjhsLmBdoG8bm3VuvO1lNDT3ZE
SIu8TnhqDQiranVjHUPdirp2EP09YQRVShzvfYyw0lPRav+W0ipBDOBmnYAdGG0cxULqqnMtRDFK
OGVN8yPb2Mq5QcdmlNA7tjaT8swRl8jSDU8bBTgsetj98zor+a5YWWv40MJqz3WnO8fAzYSi3P7f
iqOQdrGGwW0CP6PJ6V/SlJRdyC36nX9jIXav2o8lw8KNaebA21z6nHv8pt34E6L7EO1SMYB4qhPT
tzENH2wdwFEqALPAa1qEIpWUoJkZ1D/sXtTMylXSToHIDBq8EfMCGMN8Tuxs1nEF0L2rvLUx6uVs
cG+q9eS5UKRIFwUZ1u/LGWhDACkpPpLtQ4E7d7mucv5zxTN8w77TdkOUzd3bSvx9O5L1kKyPPk8k
bgK3d4mORILnzICAUh5ZZLeM4Be0xPYcEk36hIj9gSoXKgTuScDDX3mbVovI/NPXysNJCbnGa28d
4Nic79uREVcwxHU8eFvryJDWkoOpdxd5iHG1wJ7HuY+/+HDV6P4GU9agnzunWHLt6NDNJ4FPFdvy
CRM/bgpxaTsjB/+qcQQAWEVHMCt1ptijYqgmiaNO5Cby5fi9Z9dCbi3P1IPQjS2c4EtAcm6FqAP4
Ts9ATEUQvwk01pqTlMePbTsW/qaC/qlVoT70YO1dn0V4HeJccPj1TyJsRtQZG9ZJiUmTtM2tfFPt
Tn7Y0PLCgDvLYT0tfwQl61S1nTrJBl3rmlA6iM0/b6H3/Na6F7/zHjnwhRMJKCbJNyIIRew6gOFG
GG2SW3bc7qoVJhKfAUOEkq6KpwzvgVAeGIwHu0V6MgK9mq7qcuKAGIbnVXy6InF6k2XyoHUqOmVe
ysMJBsGLkuMcgdIg99S1xxXpHTRQBMWsl5Jb965AK4LV7h6CvmkgG9s/21tdJ2DicCxIUQcQmcBo
tEMTqwf4gUe7i0wwdmIe1pT7r5jiu1BN4A2g1rRGvu5lWteo1NRThLkomGxTUU0mr8/IGaesXlGb
g/+zvO489h0aYbVZSPNvVgytLgdBs1+C/9fB0pDl+rzATiHpH12Ien+mNjEAAmw4DuYK6/jjlNzK
koSxKr1cLCaGgAnAeGx3GjIepq6iDUVqHdaDJleVmm8E8hAR2YNiu5Yal2RTfYNvIzzxiAVQRXHh
c3t4EoXWAJgy7zK6l+WLCQRNz6a3P7NMYFZC57u4h9CVXeRfhqDGel5xBD0WsRYpvP9+unieqccJ
xwhRlYoJIfrgF3z2IDKScqv2t1O2SoNj5J/PtuBsTUBtaUE79xaiNm500f/tAnbvKgrT3Md5mJRd
1LsYbjQsL1TRcYy5aGt4s6FOnUZ1VmchUa2jW/63LEAwws4liIhNDuW0nK79krTz7wO7eSCjKmOY
wtksGAg4hP73y8bIA2if2V5IWyzHa2rm86LaxsG0sGbOWAANqj1/Umy5SHaBaRj3DGhXJZXlt0jd
0D8pg62fv8UumI/P9vz2s0r0V6OYKqAvvP1gycDPAsRkbFVIJQhLdcc13RYz0cLjh8vnPxQHz+qZ
NTsn6+P8hAhA93BJveVizQXEApV14yOHTm1+r4JggKuAXMpqKvnEaiTmvIQy3QnQSLoNpd8eGGOI
UZdBhZwxbCufZz9Iidv2RjEI6iWRCF1/a4Ee991Re/703GilYobcQsQJESjOuvjCJ6kPnfgTNS4U
CwBTfDvrxvdV554VCAIHMOUfuIAuA+UM2U1w8RZUULKx1boNbfGp0hAzKy8nsbdZXu02z4wdz1IB
toNlL9NWovNK4ABnLYBWB+HYuGOCwx3MyA8D3fExz7t29+Wa/AgR02mnSW8+kRtlL9RtN1+Unrg/
GttGSdMyV8T0RlFBjO/Q3a6P22+seTwjiSdPEHsiyKxdgWMgu4toyPGRbZ/j8vrXHbr6O9N6MuGN
9c3HSgyRc8EKex55ureZl/jDgaZlbTEmA0Km5a7p/vAYB1sB7Dqnf3U5tEjBhl5MZk8mjIoavP+N
h5QzMSBuu7dFeRJaD0tzDDlgUs9qQ8NvCy06UqNir9TDIghRHgLBuc8TWhnGoQsJEV5wcwnNoQke
RRpF3J7+xDM6e6YRcC81xg3Q4lxSqc8DytN+XVe/VVCNAUauGg0J0Mx0avzDtLt6mUeb1z02qJbu
BOUsSA3Vj8hlE0D7dM/NdGdDgf6XlUnE67L0scyaB7PxriuYjS+QBYB+ileP3E9gQ5gdL6s69BTh
hkzAdOhTlu9rHvwJQy1GkmoPqh0VCct/tUhVCJJiwLd3ndq6VEvIkxW5S0fdTI1iMcLTlPw0RsUG
Q572yCCubpbkvhqGMM3IeWfP7E8ufrQw1E/XO8WCIE8tGSwYJspCpjriG/xXML6hPOvlqw44V0Sr
XVaGvOdEJi5AotJnPA9ZzjovEAdK7j5IlB0JkQmUJFBsqnnunq/TbmHutZ1NQYSlxRPfR72JReUk
2mQGca/k+Sy4m5SB6tOh0AvZaN3jjVRu7m5wf0m834BmyjAcxotKV175YBxBmABt1gsVFvQBc44l
BZAnvqeO9POMdYXfz3tJMmztEEpbIJhR6eEiW+CayaO9oO13HK+cODRNjvtEcdAXl4Pg2XoM1u6C
JCR8XlHYj1UR07uR0qKrjHQ64i+ThyAD016BYoDJD1z54H2ehNaqwDPilJjW3rPkGUc0bgJdy1rp
ICCF8mOpkjXo9LzqgJno/D0fN+4SCFhmxxuTFag/F2WtN8cgBnluQ9u6yQQriTmpwhBQTPHiL9lD
O3MAjT2xTazViNGcQQe9Klum9QRpvSO0ZNBoIWsakZq+dlKidOvyhKVJHvgE+uNbemnZBJqA9tP1
cNG3/+7GrfSQH59hgPb1iqR1tjc0A+j4zfWwMT8KRXyTHkFxhRFdp0jUiFx+p4CYsWLtpl7rawoC
H7o3fhMXHWXMCFCvFRHAXh33ZZtDnF/5K+n4c2ta0+1rj4TnW4scw7wZUCGDIWH25wHVC5f8V1xX
MQxTvvY2y8N1fNEhyq3I+BBVKO4i4IRpkDe8xoVb33vyN3GyYZzTnniHIKIX7yWHGETlYl/YM9qc
Etki43LDcMc3AuBHEhh0jqwrGnrE+iOVH0sImG56IdWwUc6bdSuZ2HvartufASixermFx6z8Awkm
hl1aSvMHN5svmXFyQPsFA5jHv39rmABReFM9CwphNCJA6jRsXDia01Ja9rfNYLqfllU98Wj6DDWJ
ufRR/HsaW8TpLnsGBu4uK46jGimx2cD10bB1vd8Wi48oD7Jl7lY4DVQwppGcC+6hdMTA8VpU8FSK
uG6IMimqfdjjLWj6TaT8G9Oe/+HAD02m4a/oOuph/1RF2E7IiYTZkDSqkzywllsYQe0EzrpIscNP
s2QwS9fHcGCwmpdBoSMhOGANhQS9fUnQp8vFoR4l+ePH0qpNPMwNSZNY4ZX/5iOMt8nACc0P3+Oz
jvsWraRNoiRkzTlIAtsHdqaRX3yVnX335Xz5c4w3YRRq4450fGej+NHlrIeB4pwyMLDMSU8KjFRz
PQh0DexHhbPZZmMI9vDO1S0FOJfZzOl7k2+xgT4t2JUoONjpCNgFeAyKsmCwKHEkwsguzCCEDj1a
+F5pnXdw3wOnlK9kenfKqXWgwJrOhQm5Jg3nk54CCE8xqY1gmVTlAmIpMpOV5FIGu+k4Fr4xbUDN
sz7Pds3047iT0ixbjj2Z0B00zQ6sKZOZuyLMz9N0KsBvS428l/AC5pan1dypOaKr2GrCUwzosMRq
fFf8Ephix0LmL1v42aMMW+TYE+Zz9Dqo4VPMfUzZpwv2rm+La6dnjY3tpcJvjjfWRjzkmWKFqmeU
qJ3Sw8CWUotCYhuGVeOe7EWqtX9BPGEiAHBx2JMXpbj77Gq+eV+vljyX1ziyCazbY6xqj40xcNNr
WtxnbIz/+LsP8EIEIm0zhTtwcUB42yu1l0Zg0i3dGWDeDPvYV9sh0NfJq5wYarJZaB5ZNzGM64yA
fsgxBW62WROd76JgM+v9NarH/vkymH944e8onSo2Wi2zKsHxbMUQwFcHCMntf1oDlUFcWOcQNDOc
HtfOBloWEdRB09N0IjOqVIn6WfwlN7I40RIYoKL2n9ar8Odz+tolsDeJ7e+i/IcRJEADFXGKcYV7
SvZo0h+1NPK9v0quMLURJd1tu3EM7OddD/nnEsmxW6AQFSuDaEHJX99ZFaRK/VmySQJP/S4S6V00
vFjTZcJus7JLQyuBp2jzrZecnjgN9ce60uMp6onM/e38szNFKsdsA6vImhci5e8U9/vlfsrEIFGW
s2szn0cAfcxBAGlsXYovBYaNOzvURzWs8WtIXhiGLkMQqpWiEwQPYKQrbn2RPv2tW7StE2SdTyeV
bo3n9EwQFI7U3w8mhnE/inFzBqRNTmm64Vf7mUJTqwhm5jjCZrChnSQXEnh9HBgnXRBpPo5J/EUY
uxIBO5CfNF7CEMJXCRImP7bbvIxL3yHkXcA9Ot0rMmv9wOzza38RKeP+m8FyLwiuL78lEiodOor7
o++yDI43Qe+nLjk7JxGv7WTMUkCEPuy5FuYt3hxEkzkTfZKG1rZCnWfgkW+DiFiMXW1ML8E1nsEJ
vT/h2PkAzQM8nToMbhyM/8qRxdY9pl9ccEgfBuK70r+ZVnhjvQkjC6nfukj73mQqN5R6EQxNd7gp
VnDBiwShcZTlPNfuouB8cCzwVbHSnvbHIbj2UMp6UCEhzEuiDc6ncFaXqAX7cd9DsOzWIg9h6PEe
+fzmRkIUd1RS4rlh7a5gz9ZoEXBYrIw7OZyC9vHiswfoOZbRv4vQysqpIRb3as0KNFTcgWcNXRr5
mr4zfNzW0zDc8H6lrdQSEDsLv3EzBYCQErd2Wu3ymrF76v+nEVkUZU5Y+Ad9mVMR+ExPYUurJLDP
UN6zPJ4vT7N7FpbCsC3tYQH6JnfXbSXSXgjcBQs6PrAMpevsXt5/cdKG0+EE0Z0ayAOe4eGFYtNj
61n7KPz+dpTyaIpX5KA6S2Qey7PlJBGft9/1FmXi+YtGixU6fGbyfFZl4nr2vPfM/Yll1n4ODYmu
xEsC4OBrpMn6f8JxhZgmD3JjdSr/IRHQo3GjY61HwIB7PwPGNDyVZsRYfd83Ad00Zjq2ZEYvlLoa
r97+lFbZcuCbrtAJ7kywiX7N0YmwZnGvYwKEfP6y4XEcxCGjFJuvzh7lUhZ3dTamN6QhhFascFms
U7neuRp8vt2BZa12K+ZtCuNt5kMHNc2DrymFLnXauBV03wvbKYQGsgMS9wZRaTGPf59n1lUd70Q2
o/CyqhsZ3bdD/6R4pME5dLe9pSstZYAebrrd44K/jmBJrEohY/kP9e08Nt0+gEEX1JOMlxhZ/msL
NTe1DeLTAAot55EK+KnyX1SZrellKeFmYu7iLQP5WBRMDluXb4et2/6Zk5rHtuLcAmTf9Vg9yzJK
Pd8dKMkzP7jh2JVn6IdXZPtlhc9BbH7rnT6bJSglzlH5E0J602e8GEfAzY4PVOjeygD5tHKJFeTe
97l+mWmS5JSYDcS5S9dI9PrberuoNP5E2y8VpGO9GvKvobLD85eZeP8ttUHZrdBbFoXL7XkK3u1M
4QkNpYQXaRaHRcbRwgkFn9wAh97sO8Hsxz1CZ2nNKwhlWAR2O2fTbPoulvUrazcmTrrkDJUeendI
W1Yko8X2VA/k8ow5otIGGnCQVT08EXuA+cjCapV+VBOeiiKQNPoumRjKeuBIWtady4pE60RTLlU1
N96cVTG5pqhahDrCKK3mn8AC35GsQZR0CD0h0p2zeyvdw9ohBRk53jN6lupdhnQzT2TxKpGYB9Zg
ECdxBttypXf9rSILd3gRYa3JeR2g7g9+bVFY72lM0iE9LCHRn2+1EYWr3JhBpltH4qounAT+uoyn
8/XNo7mKdCc+jMwAuTIVHW9Hr2mqUsSDC5vl9hhC3SavUm9O2wwsoD8Kwe0kbOlyxJ6zW38Zt4gm
hv53zGqu0ZSc4BpuHUB+ooPXGdc7v1rQnNAjPa8rboZU76NTSeyc+mBa9+iPhKH4R2Lbie8JRJtn
jUPlUF0HseVqrvRETSo24xwuizfljhm32IVCwIA4qADBaTKZPw2M48nO4GuGe/XdYbCHp6u7sQ2L
7zkYH1aQXZRcHGl7IelaXtk0Nu5XYuATniMzN7lValnUzMkP8SRKMls8CFMJ1IjBzm1yUo7lEhxN
85YnXaUKdmnZwIDi8xxc7mB7NQIQ8NgF7kIizcYD/cSLI8qRdeJ96QEjXGSU4mbSIQgKQzNDp1GH
VoCuyfrwuf0WarQKzpFtuUV4iotINcdXejYI1Ocb2s7OeKFzEc8uRm7ICQBy+gEZuakEuV62vrsm
h5K1D/QffqyZK21QgOIOgIz2Nj8yWwQhPvqdObz6TWg5SvfAgVniMCeG/LRaJJ2OpwNCJIrWy+o5
vC9mhiAmzAlxbwL3EH+0GgaGC3+GNZt4dUdez3YR6wtaupkctpfiHr7XtJFFeB/DvaqCQWnyaBUj
gpdnaNV7wlh2sC2avDz6l396OosMcCEVvNExESWF968STIOhTeMk1bNalhNuHkdGsmPOlDKsIF61
IqVINlS+kZ+I68htcOiz6/BKcYw3ecXkzIJctdO9a9deO6Bo11zVomZdIiUs/qAEYRdGZBjiF6qI
USqr9uf8UiDCue8TY3Va4ke5Eani3nI+/qBtCgZuWjpxs33qHj/tF6hZuCYzoTsq669gW5CE7lpk
Rwbi9rsw/LX5LE/7rSzwrH546o75Zch30fwEQRTL5ZbxaUKMMf6g/me7bcX6d6nw9i+hNkHD7e01
0Z/0jdXqme8tPgWlfQ5RAMqiCzLfu7XycfxDG9qP74sqHULyVduoDifpYFQICwcJBsi5Co72BqdO
58VcUO6JkvfQfKY/KIzDStWHYj2V7JqeB9WmxAxotIE2MxKAhRjeUpKd7wzqHlTiQDkhwdrnqdI4
cqMB7jGSCc/tR/qjn2iqKTrvXQm7FoeMvcbxYJTRdG9IsPhYuIoDj17gn6OlxHvXOTQ+Qr4VScra
cGMz1FanLsaDfx5Q9JgspKq2989XWcbWwuFkvPPNc+El++qa3zO4oCR2JFZbRVk+Huoz4XwO9/pu
jiTw5CJNI0Wuz553/cORTIReaUb54uNv9e1eMTJaI0FrrXmYFeZzmSTjs51CIh1QISBAP0uXkr06
kUhw0xyzVDn8dlMwGy7j3BQiTqC0N1GU5QZKDDB8YuU7McKjcXNAmc7ZObEjXXfU6PQcK0T/jgTu
vLH7bRfTmy3QVakYdzyj+t5kQGJEDWU0DoE7YDB4b0xAyW47lMDBSZrUutsDNOdiBFw+RtICnvel
gDxAi++72cwaMf19uiBpVQ67IjxE3k26FNDhz3JLw36SAXPos+74ehStpLj5No4lKT5HKo87J5wx
Tf/9YE9KhOCMiAmITRf/DxudcO9MAgDGb/hvuo3m+qOrziKbGfxmXQRPTP3K6aytK2Gs/y9xs3Mk
Mk8oBNJFO4fu0dHmAFVtigldtJiSnsjfX70N6zVopG7WAU9vkVC6NaMytkveoqxCM/bVbJkYPyZ0
XXzJUlLdjBE2ES14YCHTSY6e4nwOi4PZMPFoyOokEkmsAd+qSQ7uZDyrRX/IZrVOFEVCWVyvwYN8
XgRB1O54SWeYIVyogtKJfwM/ehHDGz4UVPyd9xVJ1omlZD5CQdCM1qBA5pH2sC/4cIxiIbkIyq92
HC7kKowss1fK91RbRtb7LpnOhKGunjlUSqbT51Hhh5ZoeAZ+6+lJPXjZiSM13uxGcYGDLvrI79mR
HmleO1Dg6vZrEum6P3UVND9i+4owpIKN0fh6nvN+a+0Enm6Vn81V3ZX8RPvBxocJZwfhox9MjKKB
lLEYd2f/70wcsCwhWPqMBaozahwcFi55DA4U+KhLggiLKudFN0sOmqvuix42TxWvO9MBCT2qv3Vh
jzY+6m/wwW1qB9D/vZ/cgyNymOUAsXv/oQHsb0FEr1GOKaYLkO0Zhf1AhB+zK10F/z/usk7XApC7
xIpE5bWjlHvc8xiQOegHQhT0lOZp9Nmw6vldkKJKGbcV7FySJ6+StIKKfES80CEX40KDvbX+IGMO
YMBi4npaCtaNIrdUr39oij6ZPPo5Ev6vcI6iQtNjvqzSr6XxD3n1VAz+uKobrivpq2RzQSB4s+Xt
JSK6LfxwrdJoQAnxGKFFYnuQP25WIa78u1aiY8cZpZoRvk2o3MkCenZGnM2a3t+q+dNlMeXdbS0x
wfX55DjbAxImHsS6ZPHmOboV1eNcuuGBzyyFgzi2s8SI3m8hO8KKvZnx/jCPrsUD+e0GB2fBw3hi
m2oe9P91K4Sqm6g4GOcLROCaH+2DTUFUVe7uurs83E9QPcO74xDEk5S88t+WFfvnQT/YvgYEAgLA
+W5hU7qV6+RK1vVhYPZiMWAY5hp03aoGhPZkWtVcSiUBK0HyPa2zBvIAj5+XZUnt+xbeurgv/4cx
5cB/zXD1y2ZqZJSUQ9vJ4lfijtHaS65GvVMWjYDMsflKaNYrdCyahWNyy1HWn6tfqMr+YpbvXK0I
N9fdvuPsz8m/ak8z6YMBMzYEKbSSDKVJ2HFB1Q9XpkJfb68+nhEvLSh/8JNFh64d2AHh34nzS5vy
WyzDxX8zZK40YvnRCstCfnPklQ3GdN0/WtIjGTTcg40ojCwsT76CBl/fw3ei2wzmvvyuQBif9wU3
/T7zCoxrweB048kNEdbYH5gpEy0qJoqCTXSlQmZTVO7xCgxUvSHayjOgEleJ5jowlP/qvm3q9oc2
M4Hp4RWsu+tDvHZMQDIQwxYUO9kazYRcfzuEX3yqPWg/HqXRbkR/YVZErzSZuxRf4wLS61QxyiWI
ouGP7/QrJfdHw6BGszeNAzNJBW7DO5tGjGWDoYJDpfuS9Oq/L2ateBHeklQkGnROKa33QaQfVd5U
tssVjU6Ij4P7J4e8m3BoKJ2tq75UogtrXsdJRKjahxiYn6GEkB+TSwxCWyo4mOIYh8zbxk0zQhP1
Cr2KOMIt94DROk/F1tq1Gi+G97Sej/4vkBYddCFwqoowvxVwc3c6kMlbgJQy+3mrOdLYXUCHrjri
Taotj3NUFaqY6n3hpiiFHBcysj7fmkS3b7tjCsRIjWb33UYCl1THizFeL1OMb0pp5OX5MHnpvfNR
pxOd4AmbjtkWT5sh5dt+DXJEzjjanjGHl4Uz+/FkjbKZYLoKvFKIUCLtWdsJxCVXhvnaaBF0ARCP
y6qiEL71wvBcIfccLM20oWFEvMDvac+C4k9d7Pybn+4/UUOru1KG+Dqa3Sxl0445xH6LA7HAX0Pa
kR7GgszkLuQzUYnP/5LmJsHOqWKIfQQel3qlKYzEHKOP+ixq9W0yE6BeELMz3dPSx2yIL2PWytZx
6x3RV+7LDLi5iVOQu3Venor9Y8M+CeSILkt/43Mb40GMFXiZeiY6hKT2DmemetLdqIP+6xapZCn6
ySISsaKeqOZ/9yEMYrXDwK8HlgI4h1npzaROLOSXl7uGCOo9PWTZLiDM8wlH+5Zz2nmswjs9Q/t6
zcAE6Ep0Rgw6AFus4BYStNlRAxDgjAnWnnI6aI6CEDGmeOcH5wm+6K6uKRfZ/OYeOF2BMr0xBE5O
4e8G0aQy3MaIf67UZLQ0JSLR1YhXp3Erb/rO3rkEnoaFU/Zr+kux068iN8vlN3n4R016KDh/tJ5p
Pho3KytfJ2JhwdIc940UwIIzbE+fmRe4+2xw6MxWeVNLkVwk3++7kWqRtNlN7HUA7HYixDNE1Ju3
IV62IrNc2shUcKJ9ahKEIS1Yi4pRwuWqf3DAPRkywqDUA7j8pmPZ5CYIuoaoXB945WOGo02P3oXx
MWgH40gcsoQade9/dmUn6YTy5FItZakyIErZ2EsKtsI0h1c1wijCR9oljGVAAl1jCGMelrSKGy3z
uWIQk3sO+DQ5G4kgob8m710OwrlX7MaXvNfNyRulAfpep5YpoDEqCXWxH+Fl0lJmD/EUdlof5wL4
YCxeWZ2qWoqyVjOVatPnGvDc9i/Kn586k6tmH0+XPjk2zSZr94oj95ryWKpmH/Dcj8IQ9Wwo1gof
jZRLNwh6f6evLMRm9tCNpPap+QmXTE02jSREs1h2LUccl6sUFZHSuPBhGpZRigOVnaUGppN7s6uQ
YQg1cEfSPpuFFJkSOvCy0D+wFwnfnvQlvXNYFw2MsMP6qLtd2r283ZHSkoT0IMivfb4re+fYOpB2
lZgBEcEsUcmdleJWv+2AEmS8o2S1Scyo138AosqWyr06/diVImR0UkpIZYSBYuVgc+QNbiE8Sqwz
tXQveVgI3dtUxZlpkGMB+KFhX8bpMQsNQZiEKd9bOlde0mtzlkSr8wcfdSqdLeTTiV2lH2fI/l79
o3QixBrSM0O9t9ZfN51I6qQGDGDumdhlC6Vycc4zAeReI13Xvs/hx8+oZ6lXy1l5AvPnYlKq3d83
iw1Dj8dob4ZBuU9wvC1d9lmE3AG3d39Qac3JOfA3Imxov7PbMJw06l7SISWFnDM69Rp9hHadKmR0
ElnbsTZ1eBA+Sx5jmS5Sp0SqIvP8RINlnsV9bwkOIGZXcISwKNHMnvZsbHBUIjbJgOi94C/r4hbL
X2Mv3FVtyl4jjbzcs2qqYMtsHxxI6IYkoSRuq+XTOKILPK5t4dU2KzE9khc96gmYcYJR/PRqvO7f
/+qzTaByRAU5tU6BP90hD/8IOKjGKBGdpFxVVTnYt70skRj/CBck11adCOIxeSJhcdpkbZXICH1n
sG+Bz31MXEqE81k0T3r4PJjIKc02yoH/Vln6smEXUeTr+/dakZcaFhu8BZbwtJjE92C1XlK3YCt6
huagt8yKCxujFIaBjlAfi1KbetYb/PGL6/j/NuGsvfm9OTD2ccU7UL3NVAfZn3AO0/7sds1C7635
N/AxhXmZWkNS/uNnkTTTXUfGwXHRk4tOlh5E5SIld1Oecj9xZoMt5DExRbcFfL9V2P12IBZIO6wT
fsX4gb4xbmwC0RMYEDpV/ChKYi8z02XeRnBoHdeaeSCUi/6LxtrRwY+B8NXy1Dg4UCNWo8JZc0Yi
hv5pRES7UG3/pYavEf1I4BdkzWlXFaIy/QAGIjzquZcLHDxrunpeqkxC/DQt+Lmzth+wQdtIZuqt
Yakz+9mbDatKYcW2uqjx8uyVCtwkUATbCTTsx8j3reAq8vv9PS0YdzxFyBGQPWczeUnezEz0GdGF
uOZ1XnVIQdcXIWrhyYVwXjk5iF8ytPrq1l3yFXXdE3Y8WVsjuygbZ1x92FvKYNH0pmGTe58gQVXj
MSMtHLq1bKr9a10mw4bvLkwuzxYBXjDBcGJl5n6MSvrjR7UnWQCraAo1YVtGZvMCcd884T70h9PD
8nxd8y7hGD9u3cpJjQq4R01iaJxfeK6hry5vkNZhfPKD+ZidlMA3o0JZYdLoY80ZcanDaqM03To0
YHzJrwV89m3KN0pGqnImmhEl9PKLjq9Ln0emRmuHDJtahoCnKK8YvHXEqNXrSpOqUaszQ8qJ+NdC
DpueuousiArnUhpcoV86/EEDhBXC10lRgzn+8w6BDqcgUymgFLYEHhynoMDPmW6BVjk2+hND+lkB
mJ8W8EAArJQ4Sfu71/QywysXqdaFUpfwtGeczePZK+L35u4Vvt7qeowhF/ImaBJV1yJP8IDfqH9A
WGY/mMPU/1LcGYKxW5dDuUpOb2kYCB+NSGGBW2Cv2P7l4kGRj88zKF4o5/FL7E4ctFmlZZg0wnlj
/t0h64ZoFPzu3ou8iHh7o9LEQPMzMcHgIY+fbiGAH4i8/BfFnxGYS0fY5ZdAdqftMpYB5jwXEOMZ
+jcvFE3Y8njvpjXsDZJj3HUKtiSguNvw44q1X2IoXDviD53Hz9C83p4SVoNbzHTThFqnIAUGrLEr
0LyyaORSEnudUmi2/L7N6R/zSyiLFrR+vV5SJsH31H3I0HfBcko03DpD2c36aZxpKD3i+SRfUmRf
gT46GqeLT+Yr5TU8SM0xYFdhlRdUTgrvWW2R29yqwwTRe39KulFF7Hgn2ANdT1iij2HCtDdzV+Nj
Lqgp7s1pfI6rsalKnhHO/Jb/1eJCCWTxuqX0u+AR1+U7lSE4R2tzY43pADOAqbE1jLQSTWRbyb/s
XFBV2T+NBqWGk+DQIptOhewN2gPjmWYdfHNU6nR0UHB4OzUouAZsGU7cxbRWL7ctSA2zR4oXULGZ
NSyEbAj8/8UFfypz1t4sj4hkGi69dF6Dbc2lIl+QFgM7LjxP105mX2wCJEjFNEsFKaP+Xxu5wG48
TkKDiQ2R4p0kvfcv4Wof4jn3KeiG+4U63KRU1S0Ki8VzIoikHeO8WT4Vt30+MdgGkHFRGAr+TFVe
phD0u42B6uXH1eFJzT9S/9SBZA33Ko+5pk81csCrRpIKbWHNJvi6p8Q3RhtMTHx0YRkbasGswgQE
LJaA7GvdjFrLmf6Tc+jq1aMU67oh8RzNdeIASGgKieZjnHvxNvioVrYq7fXrFHrMHult3UBoToGj
Cm4tp4Yb+GbfFFFYiZB+ebXJNBxNyFxEmJcfb8QLCr9oPU8bcnFHVdDw1kvDIaMGCIMPV+qkYfyx
xUIMHwVnzlqeZ1IWIsDdugwUIfMaamxsWz9WyspL0YqYFzAqL8+rQB3+OUBGDHjeaUZuxFF7eYyd
x+bTFzcAj/NmcJNaccZvydNOUiGTm0fDhpjlkmj69rplG4+MEg7+ZcPdQ0OGo4yAbyKPSNZiBbr8
X3qdX4Cn9LW+NlT4yIWIU5xik2GcAyuhfIFsxrtxmnJnZcpreL3KVwkMDJEuPxcZo07brCtHDk3G
heg61MjZejLq356w4/OkEBMCpvClRDjD0RnpUoIQoXO9JA+uNwhEeAPwdjGqO5Bk4//e40xPAzdB
rsB/4Idl6IN8HznC41abeYAAfN03cVI7Sh0t5i52cMv2VPdfs7QQqMADkr8HpB1Bol2H/MJ2/IoD
SSbCUTPOQNPey5V4GqF7zgJ0SQhHfyzLJUQhMXvVfKMCfJ0J+8BUI48M65thuipz8slI4ffjw7ia
BdckP3m7rIVmYk1PdtOY7mMbRwzm+IY5cQDmaR6FT2T6YwuJ/RgLAcFLZaLYDl0nthNb2kKd1bYp
qmvwp+HIK3Qfcia3DJadPuAA6K7Ci3hLXHDj9KXrAi68uY8Vd6+JrADXh1nU+Lb0p2tfHE8EJlRg
zM77R3Ooo0Ta6DNZk+tnoDDkmBOuyQ9Y7PEACoMNboioVRdSSrQmjJX61hj92GSscMjorVtcDCgl
euIhN2pT6fEhTBEkQupswAGnW3bh21I/xfLpyYA1gNhWWux35guyO6JYB9BkkgrUa/1nDAoIAKSK
f4DnO3I9WeGlmBhZp8bUHSBmfQIEHnFmvrOi9VfK1iuz7qUudNOvAoosWhNTRgYA2TGOJRLd4/oq
CWm6ktp0kFYTUZP0cUnTNOzqucwtrn3q9UzwCGmWGU8V97EcVqK1PHyCPPCLuzNomGXa2pnjow5I
kpwH3KmszfYDRmPesqThz/l0rjVoOjiy1Si77LTjJdCcBM4Jr5E1uh8u8mk/GIhRnv1gQCAoipBy
3a3NBU01ySpy1uxsPE6Dx5V+40ss7GbY2DDIS+553BZLQzmM/jsywAMRJjPkhBsHLfI4RD6DSz1f
PAKDl7fs3jGhtWiafPhVHQ+G0YTNXJEYwCt6qnj35T+trOZwwfwQANQE5sOWEg01++M0WtfbA753
t4IGotwuha9j/LQ9NHCxCrVpA4Skz33XW2T6rkwRf6vPoXP7IW5zMq2wR0YYqxCqrFR0shfkXv6B
Jdi2k9FCKsPi8m1kygezNVoEK3iEy72rV9RJxPajqRI73Okzib0nzYh43lDe1mYrJCKqyrV8mcsI
Wc98XBAwMtQF5yTYlGMncHDaG1xQRiPkLDKR52b1GEc5p6+WDJjBRaOunafnEFC4bZNS7NT3hDKk
8GE815bLp/+w6lRqJIEyus7KW7XURLZMvupWQIUqdCxgQ8+skOnLU7hp04X/P3DoN7XWcXLqpQ3A
YdNLea/TSNHexvVVLZ3XyltZd0r4y9utn7TirkWQNZJMp4BYaC0puLq1Lj9v34ygmfMo72TX78ed
vn43wKDjcU1knD5CpD49vyv+ESHMi/YepOTBKsCEwUX77fIAtfVWwfahnDOYq4Wr5tUJmz3twd4B
FX+YDksalisvZmg/8fwmwpcwfWYB8jU4WKtBVyqRckipTt4GDgC68Yo1kE2OGW4NC5irGfyDY5JF
UeDwSHyWg6scc7TxPn4TC3WxxgzF3aYRxN00dZG9VgsYuURf+BT29wcd5O3my2eR3z2afTAbp6dH
hEwQRTRhjdrjiMam702WH3wyJ7LAvQUi1t1f/oi2IFtapXrNbIRBPwUa3BvFKOQCjjvpU8A0J9Xh
Jd4J6GiuONJXUiICdSBecJ8fACyGMTjh31XgHx5jibvaaRGYfaAbJm+INX45JPwPc8jFJAkUpYQl
gYcDyBGRm3N7e5LPcIZAxa58FHlACZt+zH0xDkXxjscQy4JXagxE6Rp7g1Fsc0Vde5yy0vs77HJw
Wu0EvpUv3XvY9QyeJ2lRBiKLL6SRkKQC5Q1o9VS/vPqD9AmJ7fDGOX2u7tnsC/bo/Nx7tXvlwH27
hS5s9xORmnW5Ewb5NKG8jr5QGn59sFdUcIhUykSVSdl7LsgdF8c786B6yUYGb28Gt4WyhGnUsuUX
n9KqU0PlwWDHtXjUZr+8yK9SLBcWF+LxpizqAsl0AnMlEDMrwaf369omRdNP3Iba+JsIIoVA+O5L
9ROrMtsB+GEg0Z5izAexLt2kDFg80ylYYoC3bIfKL+nuH4niimHKlfvWA8IbJtBWy86d+AxLXsqc
J95vRdFUDwIBiSqxlF8neXzxrB7SjU/X6ENpyqfNqIG6iPfdzm5bC63vheS65E6pym4gwS7b061x
4qIVfuFyMUQATYHfqKnQCSD/R7kI0SB4dywTVIR36RnxmK2rGllOLikXuZabBkCfw9J6bzd4hAKu
Zpvb3HPY51Qy5kOwP3/wElfDcfRzJuE131b4aJL/CZn1dzC7fP3+xsBM1DTyRxbm8Q6cQFDyZzxg
HdkGFmPZ56Od1bPL2u+wxnH87FlqLrIiXuBqDh/3HITBEFCFfX7YrdvzfM+5uq5r0a5wwYTtvfTW
tcdmO4lYDez2TqXm3OeqaCz9OZrXZY7ZwKGYAp/goqdvGmU32d4+8ZhK2Z/GuD8DxyjY0VNvLGrN
7J5AKYzRcI/vc0Ak8t7YPo6id1keqCti1d54id8AQnNneVO2WdnxQ1KSfTXgKPzFyuVh42eFNEUd
suqSQUND4F4EzMypGRUR8lF02KVDjjXSghKL2lU68xQiE1o9DmqmHtoaaAllPfEVkjq9T9Fecft9
vj6Ka1yh7WII3sl9R7UmZ5aFzvcJWccmBA7UNjxTeXlrAiqcXg8RRsj04FESWushITjPduI6DrZw
7bUPqGzU5KvqfqNh7QG4HKTvA4a3UYbjyqSVnB5JLDNXzCCY+1X7h65C4wjZB+9smtq/NDZ4BOti
7iKx2RE1rK25uw9m5osk2RSunU8hkAMOZIZdg+azuH92RwJMOdMewzND3x/JXNUHDHSf3VNKKIvj
CssjzbGRmggzS4JBPW0iAGQ4avgWmZd1J4kP5Rffs1UM88lBJNEpeNm+mwZZnJrGmfhouJYqPV5a
GNzKkfi2ioxgulidDHN2AGVyNbXPVzo9ixaFjryhh6qcmNE/MPKoxQHFLBfFymczA6MaJRUa1L2q
HKIdX/xFKrNOtJXqMfixtUgOqFo13SVleSJYfUWqaZGHhIWQpy3hNrpbrn0k3plWSvjXTp6+ACK0
2V+qIjnXdoT31yyVDMG0lGleph6koaHNWVo42twwzzhLb6eTQP5C7SAgXGnBhJodHoJf7NmWaYnT
19E2IekpcAda5Px0GTF95ES/VVWIvQzW2UB2OJwtGvQfMXgvjghn0q45zrozZS/MnxJ+Hn4pz1mU
iwkTAX1gPC3qxLWK5JQChRT0cii4Ia9+jK17SmNRisig+lg0zszrj1D3qv23j9piFIQMxZ4+L/r4
x/Cy2HY4hJyTgAAEfyh6JKX8dfMhR8blEqJ8i+B6WJqtYVf5NMJM/dRS12A7FU845tO9UPZMb8PC
I+6Yf2sRt9YVwBlQRK94rcoFusOUO/UaiwVCzOOy/he4DEZPuBGilRWhkEDmepUxiNWJgLaaP8ln
yr/fvQY6tdaecQ1WumDInU+zN9q7dhYVSq+CWUyASb4b6iMicKxo1Zob3NBF49deGywjqmT43yBx
C6T9w83W/695Yl/hRoXERKQLpt/D8zKt4jB+zK57ttxRc5aL4yOAdbR+sE6BE8uchqvSU3tOvZ9M
l+4eSzt+xymj5hGGHI3KPiYrFR7F8RgmJNgpSB09uWPOp5R16HKn0962lEtLu/UaMpzbY5uwM4WO
BTO1w9fK2TEk5qAZtzVsiMOh3IrV3ozaZPibVKNba6eeEtWsvpPE4x7t/foUWtFnWC6xK3LUkOzh
fWWMR1CjGkphZFSPClu0EQR66s4A1vOV3Ksr5reM7AV+nl1PaiH+THAECW8cp0nwyItXWIN5u5gk
FoiA3oGVJYo3CoMNeM5cj1mfDgDxc0NoXTTg7LRH1i6pv1C7oBnTpkydLnOJbI3QEMiGQ5FsNvHt
sVz2roNzOuJ88Wi8JfejssMvp+PP1H6pYH74x55wU0PCWyVlhed8HS0cJi7jsfDyNO1prHldUCXa
Tyxn9OM/XUg8XR/ulgrhDaNDsVqyeOYW96dXpmKHS2UmdpYy6YLSxRBZ7TPuLOwykVCWLksEeLGL
/LXBwepVrdGDNAqt/rVbilEAlS9obqD+ogsdjS1DUA/NZIBg+sjfmt2YEPWeQ8g3XdIJcAillSIV
bJ+DlXbgcAPUiL6CASuZ/xpEaLIKPAQezj8jKZ2GJsoO+ayZa39A0ooLEmBjOTMdpSdIJ3N3xe7/
Wfr/4Nigk+xyLrekIHDtWGTRJabYWUfEzs5BxBozH/o/LqUwNysKs448L34ybUyeJn4h9mBp4BHC
JzDBhOkc8Z3e/Nwo47ehkIrQ5wfVd3Mv30FIOk9BLOrHq6xkrsyU6fhbkCK5BKsq6FMNYVCWcLfj
X8hcSZYkAWU8DV8ciN9huhjNnLsjG52881TdGBqH3spYfx6OstMLd7dQfH6DNMgT1XC1dMgXyiz8
TYUQDR2n9IsoIpgiGLSmiKEUXunyOOty2UAvmRKWiv7XrUbIL1LG6foGqojiLFWn1P+s941OSWd0
YDLMHz4eZdAFZeIGrBFhDhtcl7ONcl6/Ju6TSW7zRgiL8b9XhapJYsJHebOVmB1QXgDcxBUTUm/I
wMgwHrk0Wup9eEufrEZxS9cxACDAIIErGkGKgLepl1ESU8VhLy4vUkYwgoAtb1f64anr/06LIlJE
St6MdZ21u/vB8xAKYY24HsNPqjkejhpK7mxoX1c1+3GqJdlXAsvtZdwvghFWOy1IG8yByYWKDTDB
Y2mPlQ+fuFNvD8efvcGvlxwkknRbZL+xYX2cps9CtQkfRhtPGvUcVEGGsKDXMzUz8QgqdX3jPmRg
94wW2q12RquGU+coMzzS7/+57CRjlehl5uDhHvwjpWwSIA6sMhYpGGX72QT8ph0jPXgORqnslaDI
pobyfIqf1pq3f4udg80of+wERtLDULmLxJNuXP+BSxkKU48OLDcdjPLKgHnmcK9jO6qqyPDYhTkD
J4ZtIH7nW+Junzw2rSvrejfiwrO8zbAqfmCHfpEWaPlF+Te1zkIg8xuwL3v2FIT9MgjjeEiXAnnz
jN1J8y9bIHuZA/3WhbzisATMd54vGp4xg8+LLouXvqarFvlhXbaeUGxMFQ9UPXFVuqjPUKKXx78g
lKXoePgTGeA0GbTdvqbe0bqEAj1CLcb1whV6olm+DL2hAHCXZ2uREOR3eB5vE3bha72q91hJudB7
G2uiS3TSagS5/YpAYyu5t3hWZoAfCl9tDfTP7UPoXTpZabNHuG/FeXichg/F0yWhFztivSGe28a8
3wYFqwoLuTDMDbPYNSiKD9zo4pMrGvg1us6vxH+B3DjHF5QZcPXLyi1I2aXut5HNV3lJcpWj1x+s
IIMhUbSjg35la8zHhsUdkmW60TI/iyDgUMynaYzNdncS0uWOus6aq+TzlQtM5Okke5QQ6zVv5ja9
+IxRNhCRw3JZXzEcgBGmP1x670vXm7mmRGlpHOgi/c4x/o+Ej64LCWX7K8mxoclr+FmfFHMzgRL/
UgeQCKTLnpMiZ16xJQpmU6MckMKTmxeK7x6PKQs9sgPsoau3uMGF+/NuBx889NsMYpoOO/oK4TZg
FGo6z1K6qKLaZ5OgrgfQvNdiy3dp057iK65NH6eMk9R860YeRWJRL+I9APqceWOvE1TimL8wz5A0
Wv6Yt1004sCCi9OzbLnT1hcDEJ8/jiKaC0c2J8m4vbyfr/bXp+aEqdgNRCcSVohswI21mRfqU1kE
ApGjl5zrBcnE8bBFuaF4EZ8TmFqKu6EkkfN0QqsvOfPzJ2GObtagTZ/HDobLCsiu/upuPrLtjz3/
ayd7r2S5emxXWwNhtE+3Uwk56tGXOzCzLr3Jh2gYsJZ3No7ZG1gEqC0Mn3Ed4IFNyKTOx1xH/1sy
D01zpYiyN1GyjoURxcdwizn5bjavurbFpta8h4XX24ii7xnk1/zvtt6SMXrXIEcxknfM4rK2lVx4
skYxGygGs8yaRtXSrS4cO7Jnb6iDU8yi76CwPjOxQ4mj8095CgKp2s27luZPjPuc/YD5tgixRkOe
CB2JjL28pLnBO9JQ220YwhwLLGeWoN3MVNVACU0Y7hGfv5RXrQ7720FxGQfslKkp0fh859qm/63i
kNjwHX+FKjmicZ2Q5nfOlRq3ELMVs4mFeiHaHMSv3teV2RhASYoe9JqX4sgZ0kylZXJnwPF0iCfT
UX4ejCFR0l4uhIleFFs+K0yZ93ABbTktx9JLW0WDlQdzJ6NXdZ4uyvqLenIMZFWYMetKG+r9gAlG
Ib/2uKzohd4efzYFzz6J+pSf2MsMm6LUtGoHW297s2b4U1dUJ7MPvNb5QRnE7xx4vlx1GOKrshc6
bsrKNLNm3L2+a9AX6sYR0Kq8Wc6oVIihmcexAHPhTnxFUiQqk4jcFOhLurFnek5KWCuDknQYiZZE
4Kx5kfSPkhzrHqq01oMXmVY1eP7Muf/8EN5EjiYhTatZPl8Qp84nunZbQKTsmXpVVzT1NUHtd+4u
l6z1LPEWQ+J/WCGR+C3lkXtBvVzIp5SbUqKQYfWdgjpWfWucybFZ7HmM0rJ72N5ce1spa0oGhq3V
sW1Kpd5LPdxCZzngQHoVXm/Bc7ebRMzI69RxOxls5togR5TrB+PAUb4ucjecSlu+rKipq9d67rUW
mec+R6/pkCEbDXcJtvq+M/QmQ5La43XsF7yY5j/EnmWgei9weLB38/KYLgKt0q9bzk8W3Vqldt+V
/IOTceVSIERw2Te6T07nzGx9Tu1M587GZEKDJZjuzOUuHd9Ddj3kdpYIiDQ26p4EV+cgpeXtt9Co
QZ4c152leo/BS9a/H8TftcaRH46gtHdZifKZyvG0KOSWu/W5xFDG65Z0sVEWYM26pJSGlM3StRyu
mDNtVbriN9EMuqn+z+Z5B+3lPz7MkythfFwGWlcPaWb3eRPLPL5moWVfkF+UEKN0Zcs0rv+BExLn
Tk/Zg2uIoCiNNeLkTNi37KOO27sExJOvvkY4/AVDRt88bBGsY3JYT9Pb3Y1AxyKro53de34U6WTF
1hkmSGixQimyf4uzA2K/MbXTXY28OscJMFtGnu2WnolDklrDWDpd79pKLpDfDKDs8AETSu3RG5cY
vY6EJJdmemVW7SBBRhbLkwSTnMKXHQe7xwYJE0yt+piZdQu0B4RMouAOWXtrQTfp2i1o4BrPAXqp
6Weze+H87+mWdIoSt6drm4abfycnl6apYYMIF4Jjqk6hY4nfhaxQ7hy1qTykg3GCH8QaYw0JcszK
DjXJuBJjXXI9y9ocpbsJkkT9UtbZE37S0sVf2zmw4vOjN2X6AhGkFkXxAGCrGikgkns0141mVXql
Q72ApbIJMtP6Fif5dMyW0sAXc1xNjJ9YF0t9bAgLaGkbiFuC8ZOl2rconTwNllRqme2672eq4dZt
sM0ryTy39q/3gV7qFQwWiQl+WGOZbZMzkpkJPsY0LUH8PbquES6TG4mlSs1YX1ZqEHWGK0+Uhraa
iyjBB97yJnr9GSTSCgoTjrf3ZI1ceI+UTw0ns62oa5s/Anrr6E1P/S31tNXGAaamIjaOkq05rzXo
L7haZ5wHRUDDB5kLMO1zA6X6gO6Wxa6Pg5AuakmN9jdImpWo6nXj6nYpAe+AcVUQ9YJgZZAsh4En
mqOyq9xg5HPKjL+wn/5ITzygbRs3TI/6na3BUUqVXmK1HUUE9K23gsioYM9yH1vCJn2KHf8kcDyh
4EZlZBeVfr/FlvI9fKqm7G9XGPTN+T0iK4ovZfCr8mq8JFG6tcB9c/sazRsMyXu2bAmPhOcR0s/L
2WcQBi75POXj1cXBc8iBMxHH3PdHib6AZlAQwCSgfo+Y666/d1AOiNYVaODEmWuHG/3bCRUhDxOL
Vlry4lYXh9Lv2qjRgKXjL31+kb0tau8NTv9yNdxr2P0xWm0RZDzERalVkFWdVxEn35DuNZIQ6dvQ
Qr0G4UA+efn1dolRl8LaqJ3BVbEYQpltKMIvuvktfIyA/2QZT6LMKN9+RAhVILxFfWTOX7b3/+BI
m5v7XEKq6ZVYyahGbOjtTGhdroy9mfL0SGeLJTw7/slg4t37lsnbKZ3rebRKS4agvRlztVmeNB16
ozarGvvQUOnVvBiFoEqcw0rPMIHrNRX3B+m1Ff9xeTN2LfAhgForlJF2NrX0iRHb0Bk+aH1+ufNy
RuWwAwxvY3vtQXKc/uuOCY/LziqrxlRba6RfmOsTs9cyMkSe3wI1Y49GQ0fB/6mzOV9SzlX51dKB
ZN2mYI4wqRXk69IKIJ69zopD5L19J9DK592097wQvGvunRkPoUAtX+iNg7OBbAC2V3CRAK9YdBZN
Cwkpo3RwDDOqT3mzsR/JF0Rn4Jqgh1fZJa0wDiiROeHyyVad5Zm0+19nJeL2XK326dxkHzrp2RLi
OJpIzbWKiop9IX4m61eNSSNVsTPDlUWumA+jk8ysP+4VxlkhvU8Wv3JudkoSYfN0FZHcGUe1X9ny
KCSviKf8fs9OJSvZBBo5FQEYvjUWIWWZ9icWZU15NVyh/CFMgV1+uE6hKJOwC2tBsK2c0Ai/Er5a
VcyevUYCf4HYKGV793ZrgScfiH6bxjpi5VGHGshZwkh34rb810bvuT0mC+yL3Utht8eY3QlSIp81
/jtonsmCb7nt4NxDKQF5CeyWdDjCL/uoaGftZlvKwtTGFGmNW+vOCkepS5/VwcFPsu4DpWN2WTzc
a7NhMOQDlIjSjShKTwurGekYFIZ0j156sghvIM5O87xRW2S8X6fRjRmlCBxiJoMxoJ8G1DGXfbz+
HalT/RbxhtqXsIFt40FJCIUpEvAzNS2llyYhYNL6vVcK5bZIyhf0OWH0j6b88RgZrgiRwEykURC4
OaU+mMgSnHGpQ9/wvdFKVlfPaS3vrPxnOMZFxpeg/9qlxAF/fcSQLurlFjwtt5nPYvcQboUNfd1t
z6wQ0934sZx9vH9JpEQMDsYDtGNy3iPsYbpBstuP1xNvph+gVk6UFiRnmC+0jJQ5taf5wVGUYsM6
4t4OjWdFb/MJ/90Ir0ZjVRPOZpSJfDOwdODPM77x+t62QBx2nj5x9ljv87TZmuOjmk+fIx4ViVmK
ImxftGVryxq8U/BL1Mxmb/OJhXiLnQZ1FFX2ZxUZm4e1cmvwjDWLqFeXSa8Co7OU1opr2imi5w5r
E5+0xkKbKgB4t7JdwdTgq0ybRDO3xgNeq07r7RP6SNbe58iDqazNaCXgULsJCo9wJ20knrnX/egF
hg7mFfCKDw7T1SCroGG86PXEWCjywXrngtQxR2+5QT56MHcdBxFHYsq9WB0Ap+cIlKVEAHyMnXh9
uIbRs5lyccH+yWU69z64PJyjdIF2QcDxbxNo/0v66rwrph142TyOT0keYwSh4UzaOHUnBhq+h/AA
BzgwDg2Zi7sZj14UnHIgE5AT482QyouOcb7k3AC1EHh9ncFBwSAwTxc/BZR333Nv1MPITw5gG8PY
0+wiIFHSQylmzeeWvDLLEqVUM6gFJQFKqQtfHVGi9jA9G9tngt7fBKWFR/OWNe3dDXkpfEBRAUlt
87bX/34HZsg9a0f1mD63d6H6/rtpj1uP/1O76EUS4/rNYMLpwkdeZ+Kxm7JClNxLxF+vHklqLi/Y
r8ppJLsL/iCG3NpKx95u0HC2MvfCNgs6Rj81Z0Pl5e40oG36NO8HeWWB8DX9aky3nbt7EwUdQbqt
0UKReiZpYsqq2tqt3daf/dJk+QZVNlC5z1m247z6zworwVZxGcQEiBZflX2ZLcoGzsJdOflsqHsP
BkckaNC/Pc0CoegKQTldrr+wOsM3eXllkIwzUSuiq0Ruxbo0JO3/+a0VSljaiT9BRVaUOv+FdPAs
fC3s+0Z8nvpIGtck9iV4NgU4C3rafSpikOA43/wAON3pUJelQPNXDzqN+KM/myal58nSyfzlxzxQ
M8SdrVRjJcx3mw0eAFAMVsvzvAX6n4w5zZ0KGrBScKNPASDwrbAw3gcHg7kII93BaWExZV6eP7lY
6tfJLyPrmO6P8KlWwLZm4g07Q6zKVUj/HXrHeIjDtKaZAS51nTDYXkB7LfwZbtbVT2n35EiDtYUm
u1/VDt4fxdXJwaabHrO+cjXlt2PIPlqNpBbc/xaDn0XyXxkkHn7ln27WwsDO3vAYt/LgG6kBblkh
zwY08yBl3s6v4kXCFb+MCnWoltXz+4fkrAOfQ5bRxSp/kcoSLeyDrN3CxM/6/RnrYXZRjRIu1HO4
+y0atxmX9xsRhpjAzLHM45FKfWskHAH2+din93DdRPBTSBXpOcD9SfSqhtjyRz6LA2tM36N8y3Fg
W7xmy7EM7JIY6EQUK1EP0+8vhjep4okbm1LcpYkj/0VjB12GJ8dfjzFwnp3+xD7C8y8rXlNoiNG+
/syivny+Z9bSkoeHilx5PkLzXoG6LgQDTIAI+mebFgsmkl2M7fQ+b+pcw0W9w0gJGJ6SUo+4KA+E
UhGhTWmdfICu1Y/88VFq5+OtQISh+qOIQUkecxwG6XGXPmD00vJ3DJQheGpuDqNEC46E9ge/9CWF
005GeF0LA8zqktAg9iAGVp1fXjVzznjS8XRK8/ngNq3+QoLWuHIikZCk6z1z9jStro3NPE3tlJsB
cUTyxGVfMuc3A82FYC2MWtClQduLJ4d5Jqm34/XwTmlFEV0dpIdIvaanno7Uk8w56nyU4p/268oL
ypu72ByEEEBRrWKweVFjBULKe8urvvNf6yF5f6LBNi5FI6jpp/Xabk5XgieJtHWkqdvGx0fE/SbZ
V5hTHQKn5wrAWdHu4U0T/SyuhZKPjno3A/VWTft4W1pUvOYYsxwBTICegdfep9TL9V34e96sSjeQ
yPd9w/kd9DKErclyuNUIhv1WZkinp3UkmY81vMiTCQSHKNq8t2xGuHbcyBU71oSLLg+idKA5QbJh
rKzsbMQhsatpL2Ja/I/ZHy13hBBRUl0ggEepitytoLx00ONXQGqQ+5sx78QpzUSNzGZEZl5O23kD
+b3S92p+cz4wKuqpiw+owJdLc91JsVmzyn1rfusJHsrpbybOIgftr+PpX/UJN2niOQU0Ow6ykMPx
34YYSX/Va51YIkY2xhTtwbcoZORbkJ/u0v50WYxaRZ8Y7txuqGc/ThE3SAC0LV3KvXYhJ2cA0Att
8Ynn1o3WjzCG0Hpwd/a9g1X5k8U5ypwqTf0kZ83GaNTqES6keApwYB8EO2dZ68Oc3Wco5qUTrEDH
chg5ERsTKMIpUIVl+MbvezGnVU2zRAcFmc3iVuYIoFMhR6PoPl80qkCLYgOI1ysSroIAKd6pak7V
0rBd59o4IQQPoKfq+GsEbTEGzCiBbLIMqYxEzYHMAnoYq+LRvhKN5cXS42wDQX6LulcPvc3yOWHS
1qv+PZMFTTExZHz1kWxo6/RLc9gUWU00+X8HVB5HQIqnl8IltEouYDU4XrXhc18f1nv8qupRpfdf
hUSoTau8Xkmuk1KaeHh4JXAPiRNjTyODQ4p5YCRwJozip9V9u6s79Ta83OUPDLb5CUSB49HxXqMU
YjcBi8Lnki5WFQQ7mecm+PBcEscpvObHYK/NPaw9+7VhgPi9dtZNn9y4McftENL841vhcZxGvmxt
32Pp0ciaLa5HovkX4nKT6d41jdJgY7Mltb2GcPNoz46TJvSuCIZL490kQszttZVBC0ZNYb9tA6Z0
8tLWeVUlSKHmw5xKWYrTIQvjWJLOqOnrZbE5n05pWb+j9kYYhDBjqk5h4eJciQCQ9iD5Q7FNMI8J
906424LnBAQTC4WlKpIMgCwriCHnJXXhbVzVAkv7bLgBzULZZkiVfFNWcR76KUqvQ290TkcLyfkw
z0xY342Zr5UBsuG9U8bbGQ9vbynMIkCzdt0YoGgCqceAhp46O5Itcqm5liN1K8ks5gWo/5Bn01VA
OJ43G9r1ztBo3VyUDivcRM3V9ppgBb44eww/699fLZ+PNmOsm1ZsmnoJ9HtG3RBp/hNErcQDCdEd
btZTt7rpP7rcklFlxTH/pPcuwxRVfs5K25DHWRSI/vpr8ZZG8puceIh0wNWN+8j9Uqd5JRV8XgBV
XbR9KbRnQdXKccX/prAeHB9428U12NJgSZpwlnzUaGMEP9zSg9lRBwQOfFsIAvV4yg7PIoFmtghy
fyEpEBlTA85ITvektJohfEwPl27aXT8D+0Av6Mi25Np+vdlG6kuO1K0x4QoinxYUFcgdQoTYqlPx
ANeE1vWbwdPQzZTmSjrxWyONv/yn4Vm9Q4H1UskENgvLWs8IpN8PqmathOknROVlgO8dMho57YDw
ARRXeWUr4ayD62DMQhBmJtDgmLnFWvsTQGRi/tKS4ZZJOcOo+SP87tNLQu0UqUCxyEyqilDlCdHK
/Yqb6PotgBrBZjyQgbbzhJxtBO9BXgElbci2HAjT9bOouyxkwBIJIAVzinrc26w4oXoofvnLzOAI
sKBk+ohv3ka6dAPJAfDuXQDkAiXzcRwNV9ErdoIDmmWdAACe+eQ1EZ0sDisEVMCPnlWdU+/pxsPx
iieVQ5MzbAXKXfOQ+yiFJUM5IBmnghNDuIGSwKKuA9egeC2t4gQ2GXgigtMBscPwRHvc+ttBACZk
nxfkQ1zU0x5xNKquRKESFf0I4WCX5/RMSLsHiZ3Ob5MhyAQxsuaN/yf1HTXJrGZXJbVgrPBPcY46
sj7EMULvJ5nbXboX2+Lo1JjYzuRv1GE/PcWEUnFEnQ8pgO4XuyZhWeUEV/LSNbB1iWYrBGI7AO7/
3KHCTp78w5MZTjh++ESn8WpRKcPlYA3EaY71ocs1fSEV4m7TtUjOcmHxlTYFui08feGnVLT3B3+1
lT4knI6ZAo+u6nQa9xEGfodota9PJF/v5h0BE2reZhGJ9RosSD7X5m+/ybI99OW1saRI03MmuMqc
pfDvD0zQKFWurNs6jfFNcTd2q7mhyiZXrju2oQ1ITBxD6VBRPvfO95IrWBlPW9TYjUdJiDpqORBJ
4+PEtCI6kf7jNfZjewzMSGpV2rsQEjWk7cwEPVb4kqKwFNXGMDxjMW0sRwwfGBOo8iD8Oid15Jaw
9QN3kTCA8/TG7aAY9zv+NBiSEdZ/2/eLT9aRBKzkOt2tI8KahfUILlrkLJAPhvtVgO8zbEEoHfep
xkfnREDxDgWgcfAhT33rYQzzXNyHFVVtuar30P7UkYOSsSybsBfZhYkLK3Hi//y0I2qGGt+EzMN5
OgTshimvChRpUco4Rt95k9CciTDSdHr9F//gXSIZTkQ5uAB1gncgK+rfiDKPa7YNtTaQcBaz80JO
nHx69k94j4WQRxd+6ZKuu+k57rnnzrRPAumUlP/asw+UscRtEx1nNQ2aMb6lFwK7zkFllh94KsS6
6fniXibBLo3i+zWhH8aNuhuynAS3vafjIxICQgVuyXeEdOpdsD+D3jY4MDxMXxPSSj47z407sIWM
lz7flHulbu/lPC1ccYzeLzN59L0HHBgBuZ+uG7fNwrlDRD6NpwYTjpWcodZxIV9R06ohJvAVOnmB
dlQjo/PkcJJIr0JUc6iPuRWi/wfuG5/s4fctgqpPPSmljmCr51757HPdTijuVKu8gWRuuGav4ZGS
VuTOU35qXXFwon5RXmOlw0rfMQ5JjyzGocWcr6wQbWLLrXf+8vDyjeyLeD0n8aiCq+p2vb3aXJQj
ilivQu/CSp4OMj5oG+XCLn2X9R+wx5N/w0ISQzIcQC1HzGq7d3wt1UIdO/csizXi/1FMn/imYcXi
qkiMdOgFLINU5ww531ZZsqvCJU24BaTQje06F4s/cpSVLu3urlQdsDhc8PN1owHfxwGG9So4Laby
5wJcWSr1j12eIgSR25dwh1DjCzHS/Qf8zSK3vgRwArAuNNRzUzFwkJheC5twUMuqdrI2WqTrE1GS
A+q384wS5Q8XNph2kOu99cFFdpcCf76i0Zy7PNTeddyv66vyCMIbt8ru+crFXA1v4lwp0ljGAu91
02mTgoIqL2CW004sTJ0J9egydr+5PXoWvUtP+hRiW8TSorFOq/9A+YXRuz8cH0Uo2rZAaR5EDlOQ
l4E9RQHl0kfJqwOQoPpoPlBwuG0iWAA1v0bDRQjnOaWlczYXme1tSlOi8p/yBbXIabboI0ebMk37
ybMw4GUe0ccbuF2LV9VwqTl1o58MPtOsZ+qGeohvLQ4Ub6KvDrY0d04NjLXdjJgeCWCYRKD3IEZy
xIcq30h8GzAmWC7QXDa8UD8EA9RDXOkGOnvsLOaBcWi+xCZ9WnBUbi5SqlNUBBcB5AJi8PRbbOJW
sVmDZCGwUgLqd4xgZR4xyWIs8SUr17BrbI2uq0OkQyrYe4yCj3zVPqHMutneIV6Qq5N0w5Z31k8B
7TA4HMNbJjJSQ78cQ8Q45LnO7v6xhy0vUQkxIw/Co38i007MgSONXSxVIlCPN7nlWB542L9KHLw5
IGfCnSmGG8tq7ErgVYgfytlRRvq399u6cPKIPcrw9T+uj7OSPLEx6lduVbBhtLJO4CVSzwuPT4lT
A4zro5bn7/f6rFt4S2rjd4eIVsqxRqAGK99ty/RRFqpu6R8snqQNXNAXSaIxdnfXAAen95gmJ0gl
HRjB9+mLcRDNCMy/ZtnyTTQbE02++oMfT9HZn6fVujoNhSCZjHPESmE6utJjZc5jr7LnNGBnYRoz
NvgS0EBtIXATefQbmbKh4uyOG549/FZ9b7lWWeMbAX4t7LYkLk+X9S0NrNMdTGTmI8rWDBbKAz/7
+UgZXVlCaqlGuTj43s/+sWCA0htUUS3sLMJS34v78D/aL6jMtBz3JEKgfQIRovDXGEDp5nXkTwlH
cc5/EZ3eCiDCCk4nG8t/nKDTcr2mhtrnCfEsRkAR/k/ACQaNtPwajHme2nlIAJBr0pNrMXogKpJo
0+9o1yc3Xcd0Mk63Ifilrh1pmCydWUWiLEwuQ/LGw6rPlY/qr1bpPwhZ33rebm9ZohDGkSIc3re+
gFFuqmczH+Sbm+MHp8UcHnERUKbsRPmTbWlYA5hf5HYtswbmE5wXt0l93uU7NmAyYn8I+JdyQ55Z
1YwlTrdofiu75+qKXlh1f7w2nMfmoX4DnGX4q0DPXbgkCPinJ8f6nBNVLuIVmutYCuUxZ+JibmhS
Ajm5hhx6HvcDJZuJetCa8gOtfBZnxNSPAZw7NeFgohHbqe626LlqiLC6l/KKcW5hcz9htWFMIyA9
wWLC5MsLbb3mADO8zmVCnAFK92BeBMtg/ZTKoGe0l4KGZl81ojV0LqKGHsSOoAz65PpDskYtGTVv
RGcKZLe1Rcc+0abxgDKY8vSHHVVmUTeXYpLk8IyQqLbhMylg/AW0frlcZ/cHURCyYUTKyLS4WSlI
8Khx60RuOdWCIVdu0l02+r47FrB/kn+LDGbd9XKRdtyDJ7q4C8zXXVgLmydATnAnP5sE/dkN5oO3
FOYvoSdDWVcavx81WMy8shxFdrUdslAjn8oj6cGKNdMnjXtucGVHFnY2t4nUnyz88haPxq0w5T5r
lf/2AQm5ajzemxMiWIXq1C3R54c/uvfJx1lk7ECmhTQXP2oez7DTyR+MywPGq9qRxsCELEkWbr1S
W1Kqbk5lqxXwuZswJ46iQISm43HZOCnI2dCOia864HRPMMgc/S29js/Z963WRNwsP34Qspd/eCq8
Ac9dKE/49g7jdM9lsxPDKY4CHb04xeGzhr68UOq1rzBtwBXv5FsZLa2pxqeAqrWsDGenRIugG5O/
TZW+C9jEQPHU/4/KG3KLeA6wf4I++Eqie/uqpPVLz7vEtgNiPFGmnYMdjc5sVETSKD0rT1Y9NYhO
MVxN9HGqmX6Wdy5/RoQMlSvKkbL4UHxuC1+e3bwtiVq+ZA0clOsSgd2k7D+xE8EMjmYMT4UDa3yM
QPN8/xgbtLzWgEn+gNX52akVYje8ICHRSU9qp09gupytlYBlbefV3hDQpzg8ezZsrrVrD0wND1MO
Yvo/r/T4sZwJUX9pxyprICbWnO0eLMoyulYbEjETLLLvA3mTY084bnOqDGFYsk30xbbRqpstjFkD
ISOtepLne5ORnlxSOWu4Hckf+qyxsYgswXVgAa1rv9hw4dn2SZiXybxYuqIdfAG5ac/mhwBUGrdP
1kLp0FFSfTqc+uypiepTEIRRaKkwVlKLHHnoLKxVP+9VcrlGT4bqah94mdnWJ/szia+b9p19gEZJ
5vb7DesTfwoZ4K8BMyrYV18lm6c0KB9XUhNQcFgeCzwGZdsRTuq4MGPrw0Xs2jpbiwSBq3oSb3wm
IUyE3n4dpDL3OJ6m9hr2XaKmxa0NsLDVTQcvsS8LYPdqQt7WV664VdsBW2E8aqFq3dKZNGb5FjcY
HF9iZCgBv7YHHh029cU0KxhGR4KUEkC/JAi38Xvli6h1QBoOIfutu6NlmTY7YdJeec8NlJF966Ni
eYWYmVjKQpPp9HiO1ziw0DpoOJ1SNLRFzassubMi+Dubhfbe2KPlKOOqI+lIPSUY7B2RnaEx8XO2
Vf9uS/9dDUd9jPcgT6PIIk1NKXkhJjXnbm0RnN5BMj5xp2WyDg31a3TtTHvUrlgs2X9uP23k8nUv
Laeb2oM1b2Rv73XavTQZhfBOM3HQtBdvUkuaLg/qvj3mJJWFg/LEkXqs3EsXQApSaaeYsVHyeQ2l
RtfZ6+m+OMzoU9V5NTk+fww/fO/JLkLu+FIF7E33ovMw5T0ExEDpFj4a3MgcU6R0C0Usf82L5OKA
PTAMsJCSpHOwVoyrb2Zw0dnXQDuHn7JAcXUJ3bk4vNbclDnjXtLI4FJTmQZvj9MIRDOEuXdSOVGQ
hw63NgyxR9cI4HJ7NscroXFdZLOWNcaUrocvQx9ZkcXBhAjg9bhglQTLLV6sfmLbVZus6TwkxSOQ
Bi31NHC70gQuugPWcof9dge5t1o9cl6/aAZ47nFXRg4RNaVx4wHvjK8R57/a58QeY2ErYkWR1bzf
4N5eZ20LnwmJyU3CG87IchfsDM5Oq8ezKgs8qKN+lExEIk21T5CdpQSGxxj2qBrNOWYat62goUEG
iC1kf10okEBQetTjzi7jMnaNEE3xiPO21Q2FPBdNfrRH7pGRKJlj3TWclgulgR5g4ONbc9pZ/d//
LBTd86J9Rf4cY36sFGnhxTaRSopnD61oprbArqyhy8jgCBWyZlYi9E0GGir9nD0gaEyfNmqjTgfm
AsNESrsAhWgFagFNM3bz9+UiuJQvO1h9ZLvYyu6pG5UfqGxca0wy0dOs2XWYE62csrYuEvOxCd/J
cBl5UaqY44MdvihwYy7JZ/iz2LWs/NbpCNJM5ae2HTt0KMI4f63tLS6M3J2Z2JQqXz0UC8n82hDY
yww2QCmGR8NEnbZ9VFWGof9TA1Zl4tJR31BKT9YdiyZXIvuynkpi+Y2RP6zHI6+kWiKSCrqyc1LO
skVxObYXAG9FuuxRo83PM5D/7oe3hDGqPn07M6UZdpr/wgjWbuIeb2wgj+Mjk0uwUkQ2s9AQus/B
L1bSLFLuvE1R07bOKo0jyx3i0Jp42x67mw6iFTXtag1i/qScOBUX2PLTGD9cw6WgvaHxaMo1XdB/
9u3T+nNlnO3/iU2nKv01JWiLMsk0LB/iSquZkcLEBZLsTFV6BAsWe6zIMn8wtEBDVotqn0OKj+To
DYYxYhEIE31ubO9cKIT4H+RZ4UwvyV4+ul12/++UCuz0rioW6WnZmD4/8HKfZmLQclUbbuDDodQO
7/p1Qa9T+1XFEDZ3JzLehoSsOOAGk2xJrz460PbtBAkIbENDJ9+wQiov8f40EikE/ew+pLs0o/N8
Borprsb/YPyusSH88zSeGMeEqcO1fZxgNjL5N/hnAteaQizH75e260+S12Mfh/x/pGt2HvTL6gq/
LOTRXhQPXXqo4exvWzy9d4jEjegghVhPlhiNnPsTRod7Gz3aWsUnOYGrcNkD2YCbcqoOq3ZAiFKX
uGbXEHw74wIvhXbhSBxV1F4IWku9ybOAaHDwjnc1Y35i4yRJhdTTzGkyWeZ7n5EFs5o1RHBq9gJg
kfTl4urVlA2RXj4O3Vz5nesesrRnDcYtPFiFi04jTTV7BH+gukY6bi6C1oPD4YYZUYtLr5jJX+nd
AKb8T5prwMGTgSVGVaHd4tFs2pCDAHtWGIusT6I5JiiQh2cbUN+HDu/1xBWGfn2p/K4SxaLIJlxW
W9FMp33m8U23oSwR+jokWw5Poyi+AKEbv0tTbwjkJlt8hGXtpXewlyld0tkYMuYUr6rN+SMaF4UM
4HmakYxuesJz7Yr8K37MQy/1pHarlQGD77ox4IBGkPvAEfQ4Jl2eRPnyBDMKWPFNNV5fNp/bcKmW
F5aM8S9Jf1GR0hTOaCEO2lvuBgHUYeov7/M7OeD/6AJiByWxaSLOXdHYOi+eagfO2VTl3BRNKPJN
WbAfliEVrerdv14IsBW67RqxS6BLNWr+otG9Yu29apeQmm1lNJ/UwVEJMt+4fXdKsbT8daeTk3+j
LA4E5pSAiV/q3hk9dYoyrExvnvn+CUqhn4V2aq//+zD96EJozqVGe+jyjSEBoNuShGNcFKlz5ool
uhnXLR8Wemc/YRkpGcBkcZQlj25gJCp3w3x7uhIWhjWLo8VKxRt/zjcfPOaJvmpM6ZQqA/ltIQDK
f7Hmqbmk3P4m0jofat846NORG41r3ikVmo2aAaksl/xU2yrTAt6HjN4TrOBJ09twGtuxtSap3XtM
T7YIz9aK44yqrDt7iUZqPevuRWpYg/nLkE6uKnG5KqQjakHE8oJ+ELto6Ywjtpi8UOlMR1S5VLSn
S0Xd4t+1CJkN/VWUnHRJQjNhUl63O5WIuCob4HbNdCyb0+dHhCiHD+5i6tTgNYmg9hejq1l+dw37
ZD9gOIMQtszMCBZLoytegQacLv8C7lODGhxXJkJYtoqg1JZXmc1F53WUC6ofO87PuPFho7ssKVBU
Xy3TSZ9u3BmnRw/4YZzh9QKVT8uSuRcNNd9DdLLnmhI7XhulmtcRJZZ0cZyCOtGudDAokOb0ITik
kD48hfzkGqneG4cIwP9J+5clnl0CBss5FPfhvyRywm97MYEX04u5JuxwOKtnk9gVifB8KnF3XhaN
uZTkB3YJ928tEXS2zF8J0SY2jveHdl06LqyJ6r/gv+eS6XEjaKD2GnyC3PYk/3yj+ytPc+VTyNMO
es30W9rydQKwBX0kx8ycZ2WmBkyE7khimxdY1BlTC84J4NNz/7MwiIjG+sF89GT5DO3RMZ9Gk17V
CCrJo3NWtlHTOyaMGNQgwUef5lT2Y3aAB8c3R58sXPqV/VIzcsQ2FfJripy9xMTgBhwRLicZUGpN
fExuVfn8nc7od2W76ilg6oJ3biGZZ5Be9Us/6V7lqzmzk0JiKyzxlaYgu3/A2UVorVmbX6kh/juJ
7okb7HdPXxGyBdBKPTglH83PA3q0sQML/q5G6vCbROFjavHPURnVLNp1H4p1rSilAkL5lwSFrT2d
B25IKlxqsABp/1HZ/MAYCKwRn6Vxdck7kRZoOR/4Wr3jFe3U0aK9OoM7cU0Xjp2zoJE3vx5Fj3nf
9Uu9DVNLodrpZXejlHRgbY7O9RacOYYxZsulwVkLM2/NpKjRr3ImvmBBuKkR5CQPENkHO6AIq6T9
Mx9wNVYp2jhxNzxHkKHW+sh0mcMeQ8ln4q/lA1WmA9li84r5TE7HkDHbmBP0Ed12cIDhP3ti6VUg
u/1X27paaoFcJpQZjjU0fV46j4JV5RlhgSitoM3dyQNGMbofTWOAtB90XCTATFEOi2j6QWp74uLy
NAJC9KMqdHL1NVcFxerr4uEXF9C+GbOLXvNo5hL374mBTQmng/MsDy46FeC3xYmxOxFCT5SzRwzE
nCLS7UGBcAM2SdOWLijeOKIwV+PA/Jb2rA+SC9V2LzblgCf82Ag6rjfNMFez6qE4wv6tigGDO5NQ
1MrDZfmz4ra/9agKoxoxn/DawD15CvXXNYEF/K7oavnESB4xHR2TEOYGe7Xy3ir+qgWV7xzI45Cy
uLmRbka2c1aemedt7O3v3g9CDBAj1cGyoRck+Vk5669th6v8DfU0+wpjkvLx4D8RYr6vNcoGp8EQ
8lEGSJW4mjyRrZE4is1Dgg3ppfgi5kSgRV/krNBUFtDiSdltFtRgJf6I+4zrdXb8xviQn9oCpsA8
KaMrol/4ZQoXIzbetFofUnt54xywsNdtdmjsFoJLWMUsiGyHGNUcnAyLincDkDy1zJrLvXZ1a7CS
2ZGQ26LtMJVu5LaqjKgt4PJFeRMHv0Km5qi3p4RDsh5nBbGc9IHGlZKa94jzBe6HEADbjdpeEqjK
ieWummH0/aLeZwF4lfHvGhTNO5h3mwe5EU7i4ksM7a/zoBRGRzS2nQKeMF9hpnZsOxEwIxgneNVo
fFsNyKzPxN67gkXJ/2aR5qrkjR7AOkMirzvQ3UW9pksVx0vAmvbptzZuxj53godmYGhohU5jWLgD
1bBlYGQldwW717gietQsMRRK1JxPePaqy2Bdg4E/P+11ie0WINr2DzGic9DRCgm6nj7hWx/QLIs+
g3vsH9itoJNdfvjNqd4vRDC4qdvhzMN9x1dsrSnSjV988jx/0Mk4isRnRkSHJn+BoUYmQTVEjJuX
9MDQfoSBbEaQa3WLoA3d2acnTbQnQMCdZBsh2k1R5okSr+2y87WMRusL+Bm8ryaFDXgHEc8e6ZQK
v9ja4hUP5qdcyPVIG5lY6Hnw2hw8UmnBe8x9eXNdciJeUiKFgJH2Oc+UWzzztCSAc0MwNA0li87C
tzdF+TcacS2n1M5E6PkOVxLEtGmCS2Rj8otqX4XAvhaFVGEIBk4MRqSHVrXg+SPkuQtC6dEFT+2w
VKvXEdoND9SXpz4DcHcVftEsJo79iSN2Non66eL+OveMgi5bcLWhvTp87fDH63TQDuflx10zyOYS
srXxjzxSsB2b0kXbC/ViiEhcCCj2TyJu1fQt1/TRvMBKH12ZxQmODV/RcmQvpCtVido8MnFsVK2c
oQS1DW6ISrZpUAoDf3UStVi0P+GATwv7mGIb9vsmyfpIRU5r8OmKGRHwa+C5AhXHGc/Zl5tPvpyP
0mn6dYiDw3H3qZ3rzKr6ZVq6GoI6CFZXrcpg7OIr4rS85iWWTmx7F1c+vdC1rCe+tsj16TRyvfhc
O1uXfseBVYFjUbAQypV5/vd4nXqEWwjCYr+h9DYtImmvjMOX7ylmc4vXpImHMZnOtdtprw7bMmVB
Qp795TsVcNU/V9EYtr5Al3r26Ey14jNfwwp7lPNub8/wYOsrC9IaBmmtkPsribrvthY1b+z7ZsVc
GolbHnbWf/8WAefi1V1l7CZy0e/kYc2RGqsGMJlzuNGCv2Y4wWF1HARL3ybvQgEzmmkdBykH/S2C
isdSm+OHe2SzC3pM8Hx9Qi6966WWBI8MHhOsh52q4GEi9/nwFwp1SVzU7TbWvywstJviz1XdaLBc
yYKdf70BTKLmclXh3kn37VjU/WQZu3e6C80OBNuWXjqSLde2weVqmhTTcWlgb8iP7Ili1tfVnaCB
RMpl8EWBBdcjUaekfGCXIszksklNQgb8Lyvl+hi9Nb1HKtBr3xC3spom9q9r4N1deJqiPvMPEFQ9
kMCLmMRuM1BJPF5+tYmBNvAvwkDzSB7JoGYVMIkH3ytEd7+nFAaMaJpPHxrjl3qw9fqLmM0ACeef
Ua6wzd2Jl+VZ7ZKg3xi5dRZ+/YV+77pygOcKySJ084OqZsXDS+Djx8jkJTJqISwq/yaUx3gHJIpk
+QKoWVzafn5+7mWwOpb0eyecfFBnLr5xtEBa717cXSBM3nhBfLL0v5TBKKJzxn9AxP6l+T7B6vEm
eKKrkN+5upo6RPHRW1j29cFpJTCYJyYehXWd7vUGLgwxb9wsUZy6Ys1GopikIPBu27LWSEHs4QAG
0GwS53Fegc/dFFHpSh3d9YQvcBaqCvxeJEJ3YTulIQYdvaF+415s6i+iivB4kZyhjdAaxDQIHrtG
rgtvueYOEvHVrwVGjM2k6QIJol9aw2aMwMLMnINK2Ioh15fMN+Odd3v3GVnOO3RYUNq5QUTis+Mn
WB5dhhM7eNtkJFYt/wep/SFJvxkgtJL3rUJzVH8CLeCARJcZGwxnsOgkpkvdMnAYcRHfYYnjHDrF
4R0u1M7jX3KMnAtu3FfIdfB8f9//ay7RhEdA/5WXv/uFWvytSdhamZp5Ewl4EtGbvRH716TRbT7l
5rzAKmH9OA80AoWqkgQtzJ2fPRJsRLrLuJcplCr5ep/cgpJK0nUv6V8B8J3jiKIA88LlcQa2QdpU
SpkKe7byHZVG8TFdJc0cJPJmFl8ux308q+/7FGHUVgLcQJVh9LWxmCM6rHknxvBbyxFt82iyw1BL
8FxydA7AnHCC7AyBCIa9yuVasbBRYUhw97n7qimc/gD9nFXcJmkIxUyxsVj1TYXFO50c13zoXBA6
FbUXImhgBnHfBINcfihXjbzOoZ32+YtPc6ZE8s3gqka2XCweYmGAaACLAqPIuWK2U8yg1BnICBJ+
z3elHEgYnxyVAf0trvmekf3iX9zjuGWIIwnjeaQb5/LzdFlPFMRgc3qI3OoQ59VilGsjvhNqMPt9
8SWTsb8iXaldOfXZlHxkgTB1pZdRA8oHj88efpKGYns+t+deRdX4vCCqpgfjfCG0LfwHRw3shBP0
6wUfGIjOdApHXXvvhlnFDtjWWxu8gqe538G87Zl66RHqDdTdFJPea9WnoITYq4iAVUYiuna7lVbn
7VGhm+/9vciwfbusiP1RlA2+Ix02ujrapNSCkGjwnURL0etLIvshm5B+FOnA01Rt2Yh5mmpweL/s
QJhsR1ibO89YffWkZ5SSXL3iRGSEoog38ybsnj2cRt2CbYJdbLhTuKbMvQ/OhqQBxYZCrJklKkgb
VLlFCcxfw8ls6U1MyWAadBFOQHIqlQm5TefyUNgqUuzfMzPsZ1xEqU2mQmEeNLkbzxur5hJjH+m/
ihdIiNTY0Spl2m3PLheuKt/VpwHkrlJknyd/PNvAm86NXj9O73VJjNLsGWDR+SlxIXAkLEPgwhjd
+Ekaza2gUDBVBeu1Xu+AHcb1rnzBixMjHZ1JM7IA2Y1/3SHUq9e6RfknRNJw786L05HKFKvh9MZA
QRRTaRElxBJlNPh/QjQu1ao8hKw5rib61Xx1CJUeJRqBdPanTjWfML4Hy31RmbuFC6DKMc4Mbsab
QzWS6P5IEfcm6pYc7DgyakzhFptFTMkg6y4xwk4eQ5ksK6RF8yUTHzXUn6fTr9W7fJOTu/AMuOju
lhICIpykXHBNSmH8LSmYY80bz4AlPYyLSBIV85ADZ7leU6XB7ZR+Jax/xzKD+8i4eTmv58x/3quh
XU7XgLl4FTdYQPrCJqNNgiMqY1yyJXD6OatXOiMMmRtC80H7jAU5Xu1gh48iTeN0KzAXRWTb3byY
YbWGhe4dfSw25bQk9CiXJ2OrnKfhysURxEYO4/HwMM3ecMRA9GlJYFUrLNGEkkVx/ERMlba/7MF5
xBCgLSg/BS1zn0xHN5yKE4IE6Dcn3yTbIBX3CdJZ5XgGWUO3iZw29teSQzU/XZsemDaIowIOI9wo
x1iYAyRH/dmDa0N67zsbMJ1kskSnY/Z8soxL3BxnJWdRKj1ec94ghmMmKSF5c7h65WqlWZi7s4KH
+b6baArYKM1W57hn3fGHw7TjdVrm4w5OkkuXcYPjLDseJO7h+6Bv6R0LCAykbwB/HhXxJ7Kjx4C1
AxkU6ev0lly6ib4j3QLfb4Mgwp3prW+S+ZSWSLqwbEcsatM5aEHTqB6N9991XdbXHFIICgru1roW
P7KnSuIqWnmRlHYtn7/2KYlE2/jy1s3/k6PD5jjkqlnQfvxfufJqe6UbpFt/J0rDy0OuEzUKnqbH
OoUS+0MlQudvcwQ2YpwlwMabuC+IrivJsuWN2BE9bPe52VKy3g/9+3LRlrRP5WCDjeaY8uGsT275
D8RaNKOiBCPj5VvQ7GkDhjzMQUJA8kwRK+/9rGzGoyURv9LiUPj5j0MxCBttEcuy+t5ZZnGCeUSM
1H4/3vW/Eq9dbH0LTY0rJfJLqTco26Oo4nw3YcUt2Ho60e4nUAKjUR2Wl0lYwixUG8wmTEtrkxDU
Fzh0vwJkB4zxZjfQKOiE5/dR0sseSiNGhgav+/lXL1oU/swxGTKCPPWBtx2gup+9mmLk4vmwOe1R
VQMldBBtslqealcgd4cbD/qmbgpMurLQVyS5jz9/8fQaL8yYSIahTy1ix3tXHR+Sum56kU9IQV1y
kZAroRL5BwFwtwxnWGsNpinp16BdA/XX5bspGt6720faBWTD9p0mJJehaysRBKFjJZtcsaXPG3Jv
bVnC2fTxffKZ/wNjAwNqgsl9O5lNC+N50fKGpPbiDJ3tgdLLx0bbSFciwXeVadjLr0FwM+F8yv93
vq89BrLnWSWVVm/ME26yBHaSzMfNlAwj85IjLqRdTN832pOtYa2Wa2JpENRHCIakSOSoPEoa/RJq
ZYAs0F1VDmz9YrW+OxIYBvT5gu2f+0PkUCL4S0wz1196LlqQ+O7yTWqLicPZ0aI1ZgbGp4dsYsfZ
KbiHTvjNmqLGAJS0Fd13RALavDLiBT37xbnCSgMfS/lSmsjfzQ+1/JQ1OI8lHvx6DmRFTsdD87QA
x1PHR4WTP6eqzl220ORLu/45/IcyXyduJb9EJZ1fs8V56o02F2ZRd4zwoN8jB1S8RbLi18WC7s3c
+T9SCEYbtAcSHqAgp3DGFtP0CtdbhSBV97gFxacnzRT7prd+Q0yXe4y7Vk4v5HYCWSSzIRRfYDGV
gMS+idqsbauon6pzUVpMnJLPt7eLZmxaHfx96bTWooK/dugiD90EnJ/3vaVdywPuTZIsP7o7W/i6
fT4HkBrfDrIfHLqMozlizfYjXi4ztWu28GZDbVVdE66Bh5tG1Fxeo8h0bHRJVYx0vV+D8c4U0/uo
JC1+NNsmdPdBCB7kIl/K4mF8X3VZ5jHvCcD2aWS7fOKzYz8U6NApJHZUJ6XaapneMdYJakkaOi3u
hsK6E3Ch9vNa+aKR75EDaXcQ+CtCnB41x8suEVuhj6jTp1uvHPa1FlwculYqcgc6FHWU+MAKWBDB
D938FziCvPB9f9E69zCJf+S9VCbd0xAd7oxYP5hi1HTUBWsseDyUZRTMpnsqjrzI6tjeu7hk3R8u
p9ettK4TAjdjNYMc4kGKgNV/F5W96uSnLaX6S0aZlS1Lr3sHDYBYr5d8Nwp11YtxLMoIrqsqFBoQ
GpsPafcp5She0xmnIy7kNgnAWYQmpaml/ShwFl1SC8cijedZcBoazEcoXQff1MV7hKVbmPJDGyes
bDp0gvYQ9wyLvBfF9gHd+b0wJu47pQmgjUMQ6KWDkZ8SdeqByLQA4RnTllqsxgnyp/pTDmqhMwhc
Osofx242mQYrnU551DHaLajJ3pl94ujX2EGPTqYm3vVJ+T3UDDZ6pqBVSTR2U9XGQbIU3yEUNQ/b
BAEC749JWL+H8V6/ByZUjIlg4Um0L05Cr7wLxIHE5anPAwjicocyG1MvWd/O0qfCByWUmQHSwsiw
gbhiy+oGJU+Vn7dpfjpHF1yemNXX+uuR6sQUMJ9/rt1RsQZECvC+Sd9GaYIPXgPE6vwJoTskTbdC
04TKJec9UmzKP3h1qqdqQ2jCvmyOkChkxIEd8xM0F49utMMbt/IffnIflT6RBWq58adlty2wBXoQ
nGfHnuriFZ4WHnNkhl7ZpqrgGqXy1ixJEKN6FnassiidElGuHFh8DpmeyACM5hDeMVhwltMqBnEZ
nENktw+revNfoQt2y/3NlJiWfDYBmJOnifGIxSPWAHsmHepivVVXhErM5lJZ6idLq35itCDGxjVL
nB5DSCVZNXK9b0VXHLYNlaa3Aa/jWFPT2+CwEoqh8XnAxAtNPGW51lxVaRwWeegzQec1c8rK272/
YyNe5MsnIQQvgndt1/LbbIt/ZPYZFCczs+yWkJcr9X3Nqg4yA3GvW23Fo5lT9pwYaflofDDhgEkY
2x4D+eBgBtk/NtltkaQ5NRWev7crM2yba+AtwWoNVWSRDyq1CF1y3GiQXwpL0pTJFqsFd+jJSsku
KfsztqtBn5gxR4+O3MnZrtCCjcD0diLHC2ya+ibBjIH0hOQShWsPTUkkDjmKR4NKb0+dwgrUvXUx
Kw7066jSuU0ywlklJFOQrw2K/w2gMng1UHeQOTZq85xzZL22kvU8++IgFAajHYpb88rZ0/oy5Z8x
HRf4HVZr+RUG25fAYlPJf52EWhhuK3Iz0ZF5FzuCWZRGfdZRgleUqBpxUbDWEVS1MYyxk3fqR8Ob
96htN+q1i2gHoxNNlR1MvEPPq+5obkd0wwth/aYcaQ/CtuZEq8JHkVSdYAHjEkUCNo6oic01CZWT
wp8i+97oEXhPAZzOlUw90D6i4jNrY7ci5NAaDP4loQgE7Dd+r7URQRScBRuvBD050g6IpZpQWdi3
Ak12MvY1EykteFNvPgoaBW2ZH4umQ590amREvMgMsj6tSYRTvHxtn+dWg3MSNIpCq2vNBnMr3Ddz
OPmHxr4FmwRBkrXA8Mxitj+iD/3zZkMExMa6mZ0pvx4IDEd3qndWrUMiOLPm2Uh1wniji/rJftwK
+sMb7amXepcoTgQFU9qQCXucC12obGkNeP7bv5oHHnbOKJjC6LXi8td/o4mclXMMrP6XyOtJwhTV
OwglDilo2K7Tf38RA7mLeEGxOc2umSwKBlvsNfcfljywRCElF2zmbJ1Ovj9gPkG+zedcu+gXy8vK
QyCUw/IEl240FNtV+bTJKN0ziCH7KRNcU4T3CC3QDcRSBoFd7ht/HdUXPUC5h3lJ8wXuNbsG13US
0N3Dvvxewsz0NLOYOCso0IkY5j+rXD2Hi24j+7adTYlKoKxDbNvTKJxj4G3loz+SRqjNHFTGa8wy
6qel1BKtloP0SE40AkFmfcbv3zuIJ62WoxgLeY9ebi4+vBTTt9VyYnwTiYlzNbhMcARkIr7HXvA1
95hxZGn9ziM41NwGNsGzVpuZu041qFzIReF1PxInU6wzXO6mPAd5sLCsr6qzewIeg76g3R7I8iW1
eKc6xIedmrdj+ajKDxzFlZh0bseZhQ4m1ofZm3zp4mGPBGmMR1begu4Xd7rPP54K+Wgf4uFIoXFm
/pzyae7a+VWRdiNWuz/A5ySEMrnE3pU4LXoJprdXrdwKrvzRXa+dYH2HjXI6AqUT54As5QYQ8jeE
1Rkw7y4zcjzs5CrhwBS6TBQ1Fma6Tu/7+hfbUsfVRed2szVueOloKY1vmgNx470vn6krUICZrseG
dozlOy78/k914nBeKh6SvYiBMLabQZ8nLKB1LTgCZZMj5OABnSqKZK0WLBCyk0MK2GXzgEbdWtDD
2uHEZ+0hdKbRBGjohJnCW0flDU+3FfP5ABOvlLhl3l3LZqSCZ5fSkGuNXCmfeFRZqJMxoCnMGBYV
cbYfMYOn7e2Zua7ixiDp8YxYfIrjXOMnOjn4po4lyFKthtRIwU0rOVlJQFJrA9PQwXnM6muZdCtC
BHgIiXhP+D8ZRKRAnuRnhMdhxLTRXn6vm8m/p4jmYxCfEzHBDLvJWSKRWUWHzss7h4mRWnvVX9Gd
n1CqHjuUUMv64ApfRXazfAY3apPveqyi+8IwoI+iEAFvayXiScC46pHT5jywGZaorHSSp484BRkE
mu8LW8reYJaDUtpVWOQM7v9OMw5VHGbPFlvOxahRuu5DORQjiajiVdJ+iEVIstP7wpoaok86hn3o
zF4cASZAa1gJ/sVMFpKVGF59QQGvm5FDhh+QAUbyLVHZcuZos5VUlzgoXwa/zOWgk72tGeSNrxIF
xDv7wfTgya7E8AiFvDdmoXEFAvYhUq0lBNk9vf6bWHd5e3XUShUWuRECxEB2Mg2Zh4EWXXYC7FqJ
nB3RjLvnPTmnVVNqJKT8yXYEpCe6M6TyKmlx2qEhKl21l/FdaPlc1oh2+GlASMDfLT2hhtrpo1m3
93PP7cHiqGOh+vIb9UvClbVgOrZ3zRqe3c/FkYwbePwE0UlETG8iN9u6dygdMoHheYNjJ3yoN4JK
SfjmBFPWqdY5NpmpIONf8gPgONSdEfR8Ub3vU6DHhXLytZf1uqs3eXlhCqFO6CzAQ3Fnmkks9XU0
RXYD8SunXJOLHfIko/d3x4J7AGHBRDF6QKco4In9IkKZUNc4BjyVfjB8/vK+r+zugOHnG8/0uhfq
YIvbsk+zrIoITLN7F6uOsX6GJ6+uzcd7CRscjY+HExOgNtPwap3ZecOQoF6+iE5Rx+sC3mgWYdHu
4ZMEk2wp1fGfIY5il/bTDo7oklOcuufrqZySSIGSh3nMpqfK0QkdBm9c/pTm5YgHGG9FYe10esmh
SZ2a3y5gS6t/243HfoM/BcBpY3lxSCvO6c79iIQ5ivWRe0RFjypoSgXCnaz92Zza1RLSjTzAjkrp
PSK+ejoPd148G4aEEb5VLAOus6UPkMnpjtk4DJImhSUrx+vJkLWnVNh6G+/cPvD3TtYRsVAepynK
k4J1quy3TNomhJvKjIioCM8VQ/dw6lf2XO+fJxTIUkuawsSA+w50sTXkAW5HO3CbAzbw9NHUDxoL
sTDAhRrPrEYd4PlMlrFXnNm1vCXC2wlWzS32MpRonGimXa8860oTE2MxvamfVU5qdrdcWjkMqxS5
nPcyzh+TJ8SwIOPZKEP14imTWo5/ZkKWRamAmPkp6M0S/7sZmS5jP6Vz4I10Xmf4lWAGWjq1XyJA
JLLjMdofsEPJzWAm5Y01El/21XUmhG5A/Nt6fLgrIWQDzKKGXlLVeWL9hzv3z0KNbgxzEEjasTRe
DU38flq75iH9yy3YxYxZVn6dNudS3lJNeSYeoS7gZyl+lJWjkDIElj08D3Mp88bvO98C968a5bGB
7nqvc1HB++Fz1l0E9dOipg/0uwy+wpZ1O8St1m/1Z2mgOaLjjNC1bOIuT9jWcc/ADsZ+OI8oYSIc
X9ytjQiYEZmNPRMH/FN7ttoeSrdCps2XiznABpbkQ0smWaKPiTf8j74tbuGFkOs2+ng8drqu87Bw
E1uUCFYv7/4j141iU/xAQFtM/+3W+YpBW89Pa30Mh6SbGTVUHBVXUHGPZPcNzuWZX9oDNnJ4Yw4/
HcHzQPseC4iFVslGvyD7c7bplmCF4HAhPO1Yx6ljEOiSKXiGesath1mt985bWKGIZHDroWRrItx2
ExVXncouVsZ6ViuM57HKWpHfeTgbHXmahKVyiOzz1VTxnyBOeJteVzWkyLFQk8GpUlcNo2LLfKvu
NXDMyTXkzO8gqg0zioMqAacekVDqyVdDrwcsXNDGNGkoQ5hUAh7SlxY26NSpcSMvnW/S25ik6yW7
e//3loBwkHkilMzKcKs8ImJhbt7MYfk+G7t8iyGu81ftftx4Rwv10OSMhQW57XzlyITnx52rgrh7
fF+ePmBimPXZt4XuwKjXVKttqTIXdLm8gh34kdjbsjVMkzRcxDF7rASLquKRlEwCMbh95FI5kysI
XoRodPOHD5cZ3cO9hJi8FJ+44JJVb6mNMIu6kcwaGlWjSrKUZqG/vD28l/8GHf5+RHpuEq/RAVnu
p7o2mfY8J+07DZZP4Hd19KC1D11imahMiE+qaUNb7acHgFAXj+Qnp+GdDzn1ZryCT9vC8GtjeSk6
5IPLLOBdZ3yW3MssPCjX6FXpaGMVARRzN84kpH/pUvNGph2e5vfSCOTwf4GRcEZvMa3qwk0EzJ4O
bM+44Mb/okgYBfYB3ahUUD8K7HjPqbabwwUuMajUG+uTAgnc+rblhd0v4qOKSgnFU8x5+/e2F95Z
uYgPdsm6arSYyFFfEPCIAJsxcFW8BKFylw45PTsAsZTqYmBhmdob8s98Fxin8JJZeaNQs7LnjKjh
zAmB/i5e+G3g1QN1oScEDn5hjJf5DgNkhandbuqtTzQvVUGCMdBhAscmHFQyjX0F8Rwl/uk+9prc
+3Zihkc0KUHtRXpmPvfRU4jpfsWHxhLfi+X/Kdmv3NLHeGyNzFzzc/YQJIVX2XIS37Qf4Mg8PSNJ
8vcq52N6E+l31jibiPgNuKSf/T81AXg2cS1mdGBVjwJ/6la7CpXhKNqr4X2IKy7PyEApfS+IIJIl
UOLE5/Cr7Y7wBy+Sakkj021WqSzv87CNCEFPNGh4EdAm1V5YxLa+nkJ97D8vBca1+c+8HVg4q/J+
FALHFPzT0ZuyvymGx0l1Pk2ggpy6CCc+QWBuBnDnHc7GXsh/c8c98r0jWrmftxxk0+jArSlzOVYF
7iNC2epw0pn3TKsi0OC/hGtCN7S5vwGnZjYKgauUnTlkpblDGnCctXBvJD0DW6Hf1N+2xWKHq/LY
/2fCbjbbNaNYrpama0WNY0rvN5Txa2Pj/G+jiyTiClTpZNwhElcUIeE4hfav+4+xcj/3HXBLwRhL
/VhY/hoVE9/Aj189Kk8aHhaP9lX8CRqV8QlVf7oz7miHayPs2FGNHMtku9+tV4gZI7Lwvmg+oCcY
GdiGIL7Tu5bCRKu0YguvnMp2rg7NSMkVKttGkO6R2vVwjofAK5px/NTwZ6H+T6iGwwh+q3HAlVLl
4rcuTElDFcZ1OngskTgsL4gxyG1kM9aY0F8FEDzPrhDmVxb0fkfHfrzyns8GsJ15bK7WS8SAEzqV
pYuDjia62pGAohxwWMxF15UVGud46KHuQximZVAcPJ9ERvx0M0c2WJe7RwkbJQHUF7DSsYW1BAyg
kVK4NNiwh0pUIemsoDYzIkWf9vmeDqqkKIpB8KpZyzeXXEO1kJ3MVr49dSyr6GHnIzDBc0qoSrO3
gPV6ar28R5oYhKF/4EjBulIecuN3hSzPlq4ZUyMKaLzPkQtV1KQaGj5rEDqnG2McNEfB6lcItHPN
8r0KdfLH8veRSZpGQ1huW+OWcxGjGNnd97lMNzkdiMYkpzDmdtkhJUSsSb9opoyWVdWW1kl4EyEN
M74l7YyQKDbt/2SK/Sw6BpahY7nI8h94Eajka2YgXAJ7u4yWyMgwfAxgCXQK0IYOOpcorZgYIbwI
dZmjQojpgHklIkbrrvzDJcQ235EySdrOx7BkpfQzt5ekwNQo5ukvBoH5cdR5LK/3XoEDOqoWRJ9n
jjPJBl4fNLFcdkjxpxiqBaoJ/YFnjCIiOTk8Qo1Cxyk9jBRv3SLs/9HsiNFcvx+j8SoIbjISBWo2
RCeXme6/15sJKNdgVy5XqVZlkTX4zLYym9J8YZKIMwh80yq82OKyD5GTBBoa0OGJDUhLZRyO8cZ5
1vLGAZRoUiNsX40K5hh8S8qCE7uRqEiGD4Etd84AO7pYQENteXaqJX9v1o55+UHZkIMTXNJ/Mmuz
Amf7q+lNuuJX8eZQu3hFMVex0Hkcmrh1c0M2ejwTEPlIDw8iL2MkwlRxcWIH/4tMk9cHu9SjHtGw
0VCSVfF4BbVoSBI2wOSMswJF0Az8VsDTk4qU2ZI5d380EYEEAnwR+gWcHdgwIHTcHSfMrvve8l0X
fZZsoKP+kZlzvbKXY1hdahzvtVkRsMjZlBgdwRncutrqEqhiGBVdI1z4NM7zE/NGWOb7Pw0e8XpP
KwGl5fMfLsmsOXMP4dvIYg3i9a0sdb7h/iD9pPcI7fdgCvONWeCaF0es6AlH/e0zbZuZ4U7HtV+M
QEDIfUGHZrLgaFYf77rDI4jqGcy6ouKBoGOWrsUU3mAHiMtYPTQ6SSXVenEpM0lp0Ny444yDE7xR
kszatyE8e0P/BTarvrUFyOt7U3ORcMTvpqE4OLVU90fu8qOz6haQKOFrBsR6PMYqUFUf0780nd6D
OHssTcJyIN/Z71oRycYwwUVEfPIHMLtek7g95UsViHum8TNsNk3K577UQ8lhIC0G1+joj3OvFWW8
29Q9WI/QHWQKCPTtLeRCuUHxFgHYLSJmAHnpec7uD7au1QJW7Y1DB84cq0F01XkvjbwUGWdNXoEW
D0sacVSfw+TEoyZSrDrglwG2BT/dkyHVtCyypFueBqOXXCCuE9ont9n5uQ7i6vWgDdVTxiQdigr8
XjlAqS6tM1hVgOPA4hzf17oR6lioM2qn3nXgL3TNpNBS+93ISEAsnP2RnzHOx5jUA1t6WG32q8hJ
tmBKwE6cSQaQw9jry1jgVk3sDaZca6D0L4OkOPiR10NVAf+bmHi1ytCioywJ5v0G+F10n51ufalz
J7rjjVOsA7BI9clpFi8Mqev46UbqtefBHnxpIbzg6LtWOxVhzIbkfVwWkFNSMDmXH0MA8qXlMD15
iyZbXIxgH0RgZh5Z9lqRSTT4NVFK/Tm3IFLsvT0cHXd8BqH5HWSz1x/HjWbRKRBOltyZpuyCQXiA
vrrj8qs88lrjlNEmudAmaWdHzelT2/nXV8qhCDbBL4LJqt8+IFvjt3EvCm57wYI4dcS+nRmwsr2L
bnCpmuQra3gGykjyPjPKG+wlBd5ADw7o3f/PLm1CsHsQ7ZM4jzz2AJFs+Q9lvza6rRbJH6qzUGD4
CXHsZ31UCTLsI1COZzz5J8G9EBGyjOf+RLuxM04b2TOtgt6mLxpBi3+ul4TUyM17rxL3ci2YemGG
NFKNbK2TIRJsrd6+Qq9JnZthjT4SWhEUlScHZLd818WDUq/ZFD2hTE78j/EWunyUg+cDxfvwAIkn
kMkAVU6rkLP+g1wp/xv8/5RCceU6XxJDUMPvO6ebi+4U35WRmAHtozSfk5Buu5B9km/zEyWmQf5X
JHouVVrliShe5x6xgTkSYtfXipMngvu9Skn6wXSv8s5vInpIelxi9FSTdjUSm1r4kkEq2vMvNLGQ
nvd5MYrToLsYTlgHijs3+BavuFZTgSbF3f4ltzE4W++pFSfeB+iB5jJy+3BGO0VU+B6kxLSPf/VW
bHVRyLWN2fJG0hGNcV8vI8fJXUwRqN7xw+hC9vzi0/HrkxW63XzcC3Zx35UJNY7X16+njSR5SlE2
+aREhJKVo26BS/1WgZ74OLAYoamADVhsZkbufrSewT5+IbvhjDDDpHOng9AtYH3YkjqpbMi3/B1x
N6LAAHHU9c9/pVLUtAbiRc+dWJZpenim32J8vhulHyX/3fe0nX+uSlHxD+T9+LnNuipNp9msY+Kp
N/VmAKiDf08QVuluqze74NiqErInkcO/rrdTPoF7hX5d19eTsKZ9FC+CP3l4uDUgfGx6+qW4hV0q
kARcd08tl65W/8moKlHhtcPAC2LP2vBmzyqY3QcTJZNgAAn2252WndgvuObykTbV4mV5v9kW2qRy
XOAhYGKGbx+Vb2CUHvqhr9/WQgnWTTX1fwEMrNSxjYY0w0spGghqhcsM1b3lg6+Fh8DlDTpn68OU
+mdaf+NcXvlab7NY+fpCmEYqodtY43gIUrMqrMK55R7lfVjLh0I2K32eWMO9LhGzYcY9E5fDsOlo
Tczq5AxSyMDsT6a6BAsqBccnldD7hDPIwMJkK6/rxtdv+G3AdeICdvDEmY3TtY9GdEtCz8Gjj9ik
WcrYgJnuZU4noxwhrd2UEH6PD6JKBfLpFyDkIctCElcd5JeVeplKDve9HKA9LajSXK1rLL+P5wbd
n25y7f5Ih/S6NLwiLY3cLBrGxeD5Af05Q/WkS1QsnkjytCCOoSZrzZbAORHTxnhebQnIzBL11UBl
4/8BfY5XvQay0ju3QzNiMwrqE+Xqggoj/h8ffnszl/YQOlooYFNkS6uGRI/B0btSvISo6pKoZmFH
V5/BPSYEqYBQ5YjRNxnPZDbRI3EMBIPZh/rvD+WqcjyPHsiOq9FkYZEk6FBG2H33U1qKVXHqWhnO
xEChID0mGae2ZaqH+dVxZtI9rKwdCGMeb5AThQNDVREkNf/ZhUYIXdYKcjjHIj2a8j/W3wK+v86Y
Amfm0YjfcrItvJkEmW5eYSMRfhKAqq4OAgIAGbEG++mS+7iHYaplE4eVUJwK5B4/ej5RHukmAVl0
wt2YGxLO31lNazebMCZMJiQO1X6KH2anij5Y9GBkwFzSZsxqj8NxJKrLdy5hMe6ZQOPKH0kVLB9H
zfk6LNioRYdM/s27R9bFtAtpYQyMtdrNfHaAZzdCmx4sjjvbBZOTw5NAPFWHDF+/dJ4ouJCJgLUY
IQgxWSFiOeA3gYwC/dZg5I7MPFk7whiWKFXGd+hZCJ6dhxYVi9D3pWmW2MOjgn96TpsVr4lM0Ebr
DCi3CoE9BgKvxXe2VyBH5M8qDAfVs+7OLc/gKjvz3xljIg+xv8E7KCSxtiPVWE4wVBtqxk3LT+4m
j8syUJ0q3X9YSWaY7mvGmvE7w5Z8vBhSoJoqtkaPHr8qjvtWzznPuIS3pmaD6yVZ1KVNH7YHY1iX
b6xNJKRWctA7GdIWGRGbuGBeE8n+PKGu9JJ2QPoT17qypQ3jGjO8mqJPifRhRzh92nEqkQ2BArIf
EV4SxajcxWBKNoXky2Pg7P7RAoQCpKwHhs+8mtXhhLZsZGCaBVRHF3SzYIcBydAlV6x/L5OXu/V8
bTQGKZrk6oV43Yu70gUooduRYA3yyah09VKt4rkaHcBkk+4LkptIzc11jPtFW31lTE4BxCzXwZYK
qp/gJ3VEZhsEbGbZp0x5fZ30sVM1Px5NDxPIwfmqxNfC6QvJ37n84f4IqASGhKb3rl+R6jRqAOpA
j8yH6ewCX2dh2JxfgDzQC7WrmxWXIwzjnHjjTnEwJTduKzvFj8gvPRt6JPaHaClHGqfDshG9tODd
+38150Vt2tMPp64eVDIhsSHVvFSCds6FmsRG94TvHfudlQaYkV5wMJ9vK3LK2k87OoTDBPZVJDr7
6YO5kEBrVnp6e7/wFdWJm8mSCX5u7mep5PN7VgSHAIKhM4VsOz7PNP2q5Iv25npRX81UFcEIF58B
FVP8Z+zsV9rZo0xiAFQjt0GBZ+HvpGo185gyLGK/aF0+ysSZdsNGzXLFuda3pcup5AOgnbUwOKmW
Qv2msF2K9LrSr/HnyDjX8yEYeq1HKnMlcLccXOcD9P0lPV8XjzOsFASZOeVntpnYXQs0dgHbngSw
8ypLkcVeamlCvhE+YreP3uvzBQWqudPKGvWcVuI18RzKxuR488k6S7kpMNx0lSti3iulBWAY5TRy
UgWlAP6BvE3ufGh8Uw7z0KbqFcDjZifGr+tEqxMyWznr/H+FuwDlR38l/exHajU+ISdcvLcXmxfW
vZg/Mdxr4waP0TvlKrjqA/DSOja3NdOYZUCwGAzcS3ie1GRWdm/0QHbbhIq9rSyzHDWD/HB0/ofK
SyBKrD70iFve6dqPA9XzUOhpwQdArr7G2GjpyGxrRojlkIgmfXKzv9lUjlOAs94m2xFbsWOl9zEd
3J9U1etaVvuVpWfA5VoGlssV4Ebm54lodSVnL3R5cQxTeelREC/w4mLhGat/6ZEqLqxFJpIgHGxA
Ci2pTr1Mbh/69cnM59bfb/MZtU09DUuKnUnb4YTRav4g4n1rV3UFaQArJlYRSY9y+nacYev9284w
1Xv1oDQCJe9NIt19urCKfALU7rL4zjr04qLZTGb92BET1d/dL5h7Sg25TyWN0Q71VFe/7gJaC3HO
lB9Evq7SI3v1Bo14z0z+x9TWp3bvaKW5fct+Y9YCB1afbIU21ADX8n+ipTVLtXFdcMkIChhokmIW
feOWiI3p8DlzShfyl+TXjJ7OH9LzRm2z2yMMGzDN82WcouAQz/5gV+Z40Nth6qke+9W2U/6UG+Jd
a9+uYxDb9WWBI5gW5sMJWrUOo6cTo05PzgDEk6P3T4gfOnzu7zEmglpKL18HgVyI6jX6bZ0riYB3
rHmdl/sfsuK1+V0XBASHkVD6W8Ewnjrg33gJ1kiDxcn0AH+YsO9zHGk7Ycybu0z2Dw0KKaeNHTYY
Pnpb9xoBrvKSkIGyqCUGbfgKu18aRqcJxv3Cx8prCx44RJrm5UOr9cuecqnnLiILehq7EZ+4NrCG
J46L8WL10/AyDdFnmAuI6vqDbECyKMu8v+7LKt5jsNHw6/saA8l7G+2yxL7deP4HWuXKQsK9jqdu
lw5IIRFAE380vBPBotTq7I6fPDJUuJBVCsnJ9ekC59V5NfAGQuY24tvFHt1biA1wP5fTgulbh22P
cvqdnj2rWK52RCex6WKOYiHeJriJsj5+ymFP50VCDFJq15c0HSLZeaxZut5AxbQLlLP0QWH8Rl+E
Vwe2H5Ng8Ox61HzoXH81mmJw2B5VZaUzB/SEJGmA+E4LftJQKmnk2DHbMyd0duBVm2JO30k2GRAN
Xca6aMsohJbeQj8X687ZaleYj5Ubh01PRhvq/xZGr1s5nOwgUdGWtlRdcSaRpby5RTAtrbBToaly
1i+qqBdpP4lSo0cy87JpS4cVeF0C/gsVcoIZ2etyQEXbykTdSG2XqrnX00c+UjoHkKU7eGb7LsmN
GWM+V3mVQBlYcTwHaTMW8xFowsgZWGTKK5uNeFeH0lqOB5WpYAzdRMtgOllHkEZ46IAZlqAXbaaQ
ZFTuqJJ49wSTZnkeGISLd8PYQaKGt55NT3nA9NSEFrs1R//z5Oo/FNp10USaDIVU95/XM0P8Bipj
tY+qjtwwamO/SmwL97xTaSr0Z52ToKgFRXeBfSBxRDzJPrv+Ah77QZdi2L25vvmWaRVTmmysMNr/
bP6YpXVS2yKOarhhEWQHE1k38WnveVvxIjEI5qodnFpuw/JUjjzUz4mU/nX56gOAfGTn3X1ex3Ah
cn3sUbYhL40i5ivfe1Po4NMzDFVifmyD5iy4r28a43f5eB3pd4azs79P5Tc7+SLkXihNgFrwfDbc
uETLfJauD/6fgI0lUQy03701mriTRYuZ13+MqZJJxXklwDODkRKZX+G6i6gWLweTbrqI/hJAh2eh
H0q1d10PXgZ2GldaHa8gHmbisW17+6EdxCCZOMWqsu/1E+Oo1nHMiNrJKnax4zV85pnMx3KcyV1V
dYoK9U5pkPnQjeJqqGf1JM7WY8f+loVZH3jBAj8EbWA5NwtOy/87rwx4JP3JBfnMy4qBCEkzZpLn
WDzcdPDJvoqljw3hli28dvNQfsJVq5JXze81nxjsC304jdezMNr+0M3ddWTw6veygBJAinDOykl/
+Mlc6Bk0vFhwfKJd4HDuvdDAaUwAPwiJZG2LcMaE8AL3TaYixjLsHhBHJCHgub9di1u8veTdOQIp
m2rSJLq/uxrNJP+n2DUttjlzIyRRn8BbaSGSf0Bmr9Suep3/McWlVZm1kA6KkXEXd1gZ1DejK5zB
qm/ulVPIPkxkwVDLu0Q5wtwPGECnZJhoklQD4MuWcDkuw8QNQ8xOn53sio/zZoDRhe7WQgUJJwPp
ZNc649LJEXwFy53qm3V68qDD3eFQplGQ5wSyI9tLaJ5hehc/N4y1vN1Dh3g7tqaXLoUMwRLnDdev
g0dfwvZbBLtfnd38MLZhlmEgVb5lelgorepmFy8+3Q+H6J6DthT866szl+GMajf6/2tvXfNK0r3V
cmPLPssWjTwK9BJVXEUdYp70xiWssKAB/EnX+bt30JN2ZLc4MU544gXlNdGGT4smZKJRLlCWLPpN
PR0RslSuyj7fvkIG5QVwkw59s+GFgmr7+Cz1dOH8HQAVdnYcHh/V6iWybFQMSuwdxbxn3bFN0A2P
B4iGw1iEcRn1IRHPJzP57T70ImJC8txdVwJB8FUjogu6p+Rb4wgiADIpCU0dFBegsqGrmGSKgSro
M1R3ZGcQeeJdw7Pa8N5NEKmnUQ1sihMdFFCFXSlhtrkq3hOkREvkJdUkpGcsWX3ikcQrFzbiNttT
enTOuzwm/SvdJVDsOSJqGlawAQ7DusY13TwFufQIbfhaVgy2c14RJr+cegGVQwUe03+9PHibi1Br
M493zx7nmlkRIXWf9Ua06+xvNvP3aC4piYV5/MCnY8C2bIfjpIvDUVThltPOweXrdZwtjxKDLSix
CmZYhRTFsHPvMCcw2VmI3DA+Das8B78uzwG7O1mTjsG1u67diI3sUTJf4eMRkzAjh3BrI/O9REqS
htrZ9nyuaFAUs3DpnZX27cxX+4SXY9YcjysJyoqVRwJLjFHQJlSmuAOM9fCMuW6VqLsWd5rFfuma
TLEdKNYCnWt0XJAONFx9BODXL3iz95aeDec9g25y2xjJtGmhMe19g0FQ935d0/iZqi5zeqahwsBa
qfoGOrwATHcPxVk5XvzG/1YOK9Yx5e6JuZyVz9tB+3UyQ/oKtq8Zy51f30vFeHVK9TpOXrNbYOU9
tD3YSRafJI8TFBNnVEIhNEgExQJoRPxHFZPmUCNPehoScrftyED/6gwverGivUcfvLo0Un9AWNxh
M9s22zmVBt0os/QEcp0TuvPN9NGj9g/kUGXAkpOIpw3uRb6u+cbXQ6dLOPUruRTTZJceb9oBmoxc
dZjuPDgCRS+jHpCwbwpFJIJ6a9H6jjdpWUC9UD1W7gcFsM2BrF+FZse4hNJONiNxYN54Uqo0TbEr
hNQmGULmn1PjXzJovmWG4hiRP7zst+CgdR6h4GA/njCdj+WRDdhyYCMkgPtPqch6h53HofxkWDOx
JXgfjV0WMtQ+Q4EfLdk6XO40jCDKJ7rvbVeIAvW/NUUzYOGXtN9HCV/rf9AtVR3p93nDyiCkyeYS
3OOkvxrLYDKUC7jA9YZxXikAANYvy3g8CUJdNW8CxMVpaEsA2E6fbXQJFWN25Dd9SkiyInK9sea7
NVVjOPIYgVGrJVJVapDjVuhGtyToWiuUA64B++FtzMrYdpzOlqAFeonesUj2hOtKRmcQ8pz2qc5A
JZe3S0Eu3CG8qfhDvz01iQ7YvEbqpCiuuMzEuKqcuK9bBUWikADKOKX6cjTK/zt0AoiXkqoL4tBn
ZlxcNVA2nA/JspZvk+autyrPFztHDQ8KQ1kdWrdLRoO6wEvhwFvqoabhKcrovi7N24GK6ZAyWigB
sWxkBTX+wgFGccY7tW8cOe7zC6LriWJPew7kc4albvuvRUz1oCZeGQDe6EZCy5KRYQ9iHNbYVxLx
LPUnGzEuGqEiSXje2+HecgiYAasJJ4DK9tVNZU1J/CynFV++0LFg1UEikgjxdT1rgy3wuGyEeLPh
1tWprA46vP9yWPNHHCFlKxE1koot8O93qQPR08mj+7uicV0+Jt7rZwea4s+JYofbUrUjc+fh3CyP
+GY43Ahe1LzOmCJHGkjMo3+ZOdjC6ZWqyX+Hh2axrAxuhlCu7daEnk6aWDUcdxlFucnbmKZv46Yx
wt4XQMlbyO+txPn+PDFcoXp+L51A+OzgUcToSJ+uuh6P+l8YXv9zXdeDTqbJelSEvN/bUSeDuexE
NWJ8xv36BbfcUtQih4e3z3n1s9s3I586NMHu2REQd3JHgafNegI2n0N5jVjv77ZPF+Lr3SwPSrBG
4vG7DP7pxiFTm7NVhwEL8xe71hKs2dFW5EHx6doxv+/HB4SuAZevyEYaJf6kzcOhxxkqBxz7cknl
NOkNg+/6LI7Iz37T1LbZoVF13QUOcF7FEazpQKRp7sr5FHe+CEmPKUGt+6YjxgX3t9SPqJEBC69H
Q9WY9cJc5dFmCSnET5sMSj/qifRPvyOR0iE1yyDtNTxs+BlptyTdTbmFy+6A/OPKSZVN/DY5sAbV
wggHEr7h8G5nqYR5MW8rZpsXvhB0s2BQTrz8dlCSQ3xmoJGOfH9Efez1lHZkSUQtxvbk1BmJ1RL8
DhNs+4sX7Kq4TFrRTwvuzHtHRakWNWW7dXJ44K+mqAOJbUpk88Sul2azkK/k7tNwccfq+OkRaaEE
RctXBsEcICMNKVp4GuEOL8DUcs0ocMLA7juh9lA4t0vkEvq6eEcfws6FnyLJsMbLuraDpc8S6rx2
eKPnz5v/dAFLy7WmjELfXghE1qldOyhpi37fS/v7EB8QznxuZ8e6H/5lEayrINBgLKTWWgxojUk5
pMNrPnHznJI6IMMdtJqIkCYvAwU0Gvi1eSZHrRgVtOSv/LM0QFd0wauP7j8kLYmn5xwe1Y19mbhW
yQ/CA9UR/3Ud7CE7GLH7jA9qTIsSlQq9SVRB2NDgdmbARxJABvfzJFLrLE1UBs7PRp1kLePCbKqg
O6EGX/QmXApJcR8YhWR1QMEhHEFLCiNkrOT1eFzO/NfSuMMFz3ulql/oBAdK4AGUxAQ9ALPvXys7
Z14Wd7KaQxL2lfvbtdzHpG2WN8jzy6oFXiEs2o3pK6zLjLT9E+nY6cHVuw/XBfis0TM4YYeW09qA
+KxpPOvkekT+hJcR5Xs2Lo7tuZTW176IWl0vrQbFcdCx93/7Jx/wKHITp257xkuUoE9Kb+hcbbsS
z6ZMhH+pI60rlgG+5wrst1k8lfxEHkAWZaIvvxr8IbsJPRxMN7s9ccSwWtfDJCe/k5j72EpckodN
fUIzt4VOT+CoaKmgvOCnujBOYSUQEWdMJQ/29ZZeK7Z8avKTnX9T2mERo22kr8zn1md4dhIOkWt3
8LYNMkEezdrAMRbIdp+r0WuW3doO73r5PqSy9M4bPMW+r/jIWj0fyj3Gj1SAk8Dyyr4yn3ByEcCZ
qZqaq3p+ECMYYscqTfwn7TIBZLMN2qHhRrWyHcJSa3EvJa0Zc1fnGmcGj08ggsCvFNMjHWe32gNu
MdbJmCBeVmDkqLKh10xWIew+7n3Az3QDgB4nPLC+pgARMYH2KrRpBr8gMJhiCiqgFrjkkN3Ly1Hr
JutK9lcnqcSMKe3UASlu//fBvqJkJ9BAZC+QTi4G3euuADVOs79kOJf99MwqgUA8cKsbKODm4WqK
bWhLv/4hesmGYDHmDwJtPwXsQkMpCmIRvQW+kCX9hXtG+jnIn/owIWOxOJX/f2X8a9sR2dFbGaZW
azyCOsJRCthDmZwfzQpPRIRMj3Z0lVcNMpVVkdvH06iM9AsrVQfA3r++7gYtuoPdJ8zwFEGTTZZA
LiSKzqDp/nB7nn3vk2sqlRUiQ9JzYd5dnUMySUViu3l7frHHvWssbVkeZkX1EPr3fD9CboP5KtMC
H1qp03DvL2XO81sc6BLy6bEq36KqojHar3mFTtQ+TPOUdYyjI/tbn2hWV34vvPWZxECWa7ObjHJo
SzsXQHBFKGXW27gLMm3HXkJL9qzJstbCsl6FNK6+tX5f4ad+Kqka2ychYlNg9/9AXCJ9YFz10BOL
9+OdZiOlslD43c+iN6s5XDDV2uNLy9tl4um4M6RAMMaAg9E/P2qs0JWNmBkGQ71gmIWRoJNB6Hko
nIXLY1g7rJu7/AZN7KBcPWR40nA9aOxsl5Vn8VzpvVbgNb131PEDx+92FnIuqZEmE8ym1hNcshAc
KjS2qHSi9xPgga1TLdH6P/Q0qLOFOP1mqUOcuG84PaAAkxYjcmEEO+DdIv4TRT5yBjIIfxdWtVvj
5kzkC3JwbQgSRZpvnfXFUa0+KZYgc+7o7KN6Gl7sw0aE0Y7UNdNYx/SzX455cb2owERQS47UESrU
U+Mk+YKKifrzO/si7V7uZwlemKu/U8tnBeHt8JNkOzbtvcrL3j12TDGKYDn64eHPPy3qLTCjMkBn
cabWbfLm2n2/Ym0ILjk23fbEZxLvTw/z1eKWgvokHgQYjRAjnestIqhy9wursEZ+i81AkbXalvkH
erhIyCH+uhGFkikruksApWQKoVzaJ5mCz4Q5dIJ0bWPBE7cnMIn1EwNsnfJG4nHkKjRa7BK7GUqM
V3MLXN72pxmIc4BFfh95ivg1ECurjtTc4fB3PB58MLxTgxm6+uiYYcy5UQmK4rNEXOTpvz2CXPcm
ZXMOFLfNTwcbdxMM7M2X5y7uyEOVdr2gHQs1z04O8PW8mcSyj73LF9GmkK0ICLHH8mxY5Vvw1x6s
78ZiVP1WEBY+wIA+nZQKA2LTKvbZgP5iddF00y2vHEOKe68VtQghKRkNkj3zxmCnbPV1AaGAb23Z
ex0dy5DOLwYW9gPCJ8/IkqZo2Yo/KkIPEeORPj6KnJJcskdSXGpy+zTIPJVTnlACsKM6YDVOuU1h
hWyvsUJO7sPnsfVYfSBH2Ns1XLlN9gYZQJqB8C9rC8en9rKGesGcjy87340fbPNVLlPtJ5CIStPH
e1iFA5g7+HDk6TEjyboFiCk5UKD7Zz8mkYwhIvDAeMQ5/I3rJ6KDUDQVj/rK4sF9j9gy6g/TPpzZ
kV1HDlslgsByOVCXMmsQ9HOxRpUDPogGkGQeH62ix/2z4zkW8VO7zOa/7EzimvdnGUOi93H+RI4Y
JcF72Sq+dbOknyOQzkAyLrB/coJN4fDqos4E5e6foW6IwICS22VqBTlKrC/tNtgBSyyy2vsmWSxS
Sai8x33fwFMvDR8AJirdlYG9O92Z/FQQ2b86Yhs3Ri0A1uKdndpDKOhVnupka+JaS4SAY3Ika2Et
wQAaoWkz78EJGzIk8hle15jXKCSFUqpD0v3Wlaq/5f12YQt9Fj1ydpnoWAflHt63bDrvcgiUAV/V
VMLx6deh62YLXSaIwDODunF4jPRCzYmdU6uVvGy9VHgMDLRsS0t3P+JzFtNUcaq1DnI0wLFKL1L1
RLkr6bk7zegVpjAAW6PXoILrsueTT7NhDgJON+r8lS0KxT+kYFWj30f0WsdHcQT1v9X7SN+GVNCZ
4AX2pK+NICO1PFH6+LgulRWGerMjiL7nIDp8O7FZ2Yy2hMHhigIItmiDSOnjEVSkhVZISOL2nkYh
xQYZfFNqU4vSS7AjJ8h9N5jJH8red3x9x4/cpPJ1quPYq8/TeKMMeqTs4EVTQ+8PmHSsqvxHSNAu
6O3KjL0T63eDNF3vQUMGcBq9V06VByNemlk87z4XB1+IhPz5O0/2wEPsrYV7qDIFEwyEslL07fpV
IvmsOO5SaI3Y6IktuB239DvbmJd/DokQIloOfLG2H2dQDePVI66i/VfxoPKBH78KHkPUggOI2VmK
4LIp1kciPQZClHzqcuGjZOvzyAb4rXCUe+oGce9ZaiyXdOlzlF5NGgHdCEPnRAoINKYn8axKwioU
u3YMdRuGrAF8e/a2vvYKXNcje2uU+Yzc9rHB1oCt/sWHruif4gUOIp8BmCQY/HLMTvqw4z6kqmDs
PK8IzestRvR4EnZOf0POvBx5krpj6Z9G964251O5mYq3XEJ7W6hu2intd0CWRnJBHzHg+5MGC6Tb
bqMHq/GsZVJRDHDCxoPDCTY25yBljNv+W9UhBK42iWECYlbwZyUgR8F9L0m3WdlOxaPgqmvOTqUO
t04OF7AtRpwCO006nuCwN2hUI4yWul2+2iCupTRlOxTzlEU+g8Mn5A6zlIuLHrNTXOaIAlbKL9p7
0xpWHLJ8fBPL0aDvrc2whhtVqln23jSqWT9PH7bpmy9lKsoVvKlwwEXtarYM9yZQP+kSRUsQHsnE
j+R+qFvo3DGOAwKaLy1njB3d7kW7a/FMKbcJteln9IRiz4KV/NTHbIrk3Gicrs7ym1Ij8OuvUQiZ
XDyKcxxr+vClcKr3e2kLgyJ/BEznOFCsdMxzX6GJJXCRv6b3iaqdUuPlcvEDzH/66lhpzHp6p6QT
lEVp2Peh55SUo0r3Z9zGBjz0a8DSC2IPbhPAjFlWrmuIYL1Q82CZMyqAYN0nN7IZPbf7ofOoxcu2
VhMfX71o2LSQ6vI6jXVIavkHUHDyFM/Lvhr+pzYKycADQtn9b8bWjkDxzF2TyNzDXofkj4zttJuj
um9cOYgRw24sUqIxlOu6cCUWLVS47OKxv9O6BO01OwaVpUb/NuO1mmidOt9EhW4YN5UBew88C+eK
JSypf2FFyjoAZ1YT9XPiL3h2tClhCHZwvsYpqATuFpblZiihLgyuDyOGm4hN4F0X0w6pM7odjLOZ
gxL2hs7ljp5BmMIHTwYrDCiV08Fp8Wlc/lWDvnA4xrO28LDbeg5PYZ5a31iVYmTAPblQM95NkS2L
JX1BAVIyfVoANDO5rY3TvmIfCChIxkItSePkqeLveJc4tyLXgl/E/Dhd+LioRqafix1F7TCVG7p7
L6dao0uErE9i0PVNvquk/vaVaGWq/J/H+QcLapenCylwkk3X5mXj1O9GUm1l+QR3HTgIzVbcf4qO
3xM2woLu65DUqluV2q3glLyo1VG8DziuIgpvRI7GRcmiLXVuyFf+o9lqGRerR9/68HdLGnL4fl62
2F74DKedpXMnLjr36VmK5JqyFUUFMzmt3ENP+c4daqMFIBagGbeAzQjDkeM22Ecac22pScctpi29
gE0HAA1ZFwHKuoL7xnx2HaUvhwPuE92Y8V0CB7tbGSrMw/C5Vmsbc7A7R9qys4Bf/BomoS/R1unK
LRVHbw+ZfbcOdi57P9w3VAYe0KrzUH1tdyzoCOwseo+6hywev81dk9iEH5MnbJLafe5Mfm50tUqM
9I6+GXlHbdz2vPMKBgwVGiGcl8EB6x04DOpHFXcfi21d086LqymFJTHWnepoBaB0F1mDChd5wf8g
+cabZ3TOoNhPgEbMnSS9+jqcS2jgdM7otsP0Gzh41dgYkAoO4oh4t+YYbwYxBLz3Q6t3NqftycAs
Lxf+qXUz9A3isVCZfCxiG+PdsJoJXO52QPQ303p3i6e1z0F4hAq+AjLNHk+EIwztsZkSq1zbv8Jw
l3raItmxL/8GIi6la0Rddd69IZERLybvB+m+VayGnUIzCD4pkKsRAeJ8HlDYmoT/TCG+9UbSgaCk
Crhk/HY2l7uwjtUPoF58z1ZzMKmbXC7GpjEBcaBGJ4hCR1H1x6H2Lzglq5UU+aSEmmp+FUczALz7
8v4kvp247YZDaTQsNId8F77WaUzggggVqSkRNo91xnFa2e2qVyxcmHKc6RO1f3kFeZ6HpnVld6/o
Qz4rfM96Ta0HXMwxv7rtTHtiFh4Rvn4zl2URxZIVxvTowQSKn5IH6oqqim6AhyvBsp7Hv0uW81Ti
8Bw6tax4QxkcIV0XYLC+uE+q8ANZnkHcS400nIoGe6oh50IPFzBMQveZl5wUl2+8M3RyQDSIkZVg
xqv0J9tnLVvBpxpAtSO27nfv+rvcdRW6AOmHl2QhVlNQATFK/D2jh6a8WdFyn/ltaEExpmLCXIgI
EQPXU/YoDAaMSKpIeS1kAcBM6kKZCWGtoeQeiNw0R4xqIxXOPsAo38ZZOLN3FBOR5o0vuXpzGMTw
aDcqpiZrUP5JboHz7th68AYLcFauAqD9DkQYTPPo/Yv+ekVb/OueOUcbuH9AW1mqFtSAOiTSV3ai
MczhpBPrZ/XaW9phpNjy/nwlSTlDaR8DLUOTJ1bAV1jS7U9gPjS77TsrbkLKxzDkUxFesJYanaFS
HtlCjMZggotyYwa0FTvSqR/mEe7r2ajrPgW/CDezqe6S8GrxvymYRVgp8jjOvOR0aPp7AZUqRN0d
6Uyzn3QAz2wYWONe52X9UY57BoEdJWnebFTrHr8ZGJCrddvifT8CMbAwBTaPrVzo+kAfA85I8oKf
WCtFqIU+urVvsdas6dMhgoVFHucf/jr1zLdwa4lg2Bb4w/xqa0t/LHiQIp24Ys7CzCOM8uYzihdd
UzyLATh7XVLpaFovum4YfHDLjbOYR5jvWuO4yeQuwsjs7XL1enbxq2wxzvlVkTOsLSLI2RmhnOan
2IglRWGupdOdTJTu6T6lJ1AQJUjHNg15VhusDFT7x1mnbzm0iw8bUezPNkBSPyA88igipX3fIBRW
xeXPXeJPuY7AwDPr96UaAGbXRGya9AWlPDzUpgqVVlHTBBmiS6zfIxtSZUh6EHYIwSl/V/IT+Dq8
X81TCMc8MzlWMZvcmlUvtIBZXZ/9iSjbgyqdmSCg1BOd95zZozexBd4k4WNp5wEKDw5xo5rkmvRk
RzVyPMcKyyo0mCtkOsNgobWCQX8kYfgXz1/sGKaM8SLCE4GJDWpJ21A62f4pP4HlneJ91SeYmFQR
PtpEZ/w0ra4Byu9tzY0TVQqov9RqNQ4OaSpKzVAUyA5/kWyKbrVO0iMyZsLKDyVr8piQsMXavrf3
RU5XlNwCChw0bs9oplBa6sUSICr2BngvcWY5zP2m7g/KG2tExtM/pqj+S9i68vnjvaII1+vii2py
vkMsHl+2K4tfK7cTj4tJ6i1c+hAQwieRnn6XxoEDLCXP0a2BLTijusRhPbUQ0nLifoAUUAGXkOuA
E1+XFWx2sFT5UQ8kmkgYXi2C5bwgChILRKH9t/EaovtNiyooR9J6YYvnIsvpQDEvRb8VEkK2b/e8
nmPuq91W8j0IW5YMYqAmqYKYCoSK+5uj1dH1Grq7qkJMqxakru7yaQdHD18bnGk8mwEj38QYCqX0
j8YZLRCO05Duf/c738mE36MT/C/q7PFHOuf3a6Y3RktDDM8HFmNpa0lKeMx5XkwgRaS7bsqjInOM
njr/KcsJtXlVxsVQuA232nMlJDfdr+BrWRpZMSLNb3KhBZT2i0Jou+IBAGdUaju3fe7ltJ8dNJVd
r0aLQ3S792ziqpsZ7r/zRPLKV7zKWug4SRxXtmU2FtFIkiSFleVe7GpO2v52RPLSMejdyVpoxBBD
k559ebqkjMMBlMaZ0saPXB8ZADME6NKfwA/DN+aqtMhjatqkiRyvcB3YEj+SuyOlkfsuJByh1XwD
DXvfyOehagK0N9Kdx9pQlJd/L2K7LIbhpp/1j4oyY0vSSylTBhPaygANCI46PV7sdDhVHc4uNFCw
UhvKJFzvDQaMzUGHrYBKwPfqjH6ZhHWyetAOtL9Na9eHj7ws7RFibSMmY7jzzVey67tjkrXATgRg
j+VmonpOq0YUQOU8wiAEnHrD5gWrMZYvZEDcKn0vSjP+CLdPmV4zIfwQL8TiGp4+uX0v/gPtpthu
peI7CCCowyxstFBNn2rbzinHPq5Yu4tHsl05cutmWXC/Q+ip+CbQIBIMXqSR0llkqq9pQl2ZJA4t
HPkUolswLJOQ13vpKIx8bZMoVjrzHR1eXMX2Vm/YOOBeLlEsG2I4L9/VZkjWzYURUlyCMS17/xt2
P+EkW6+79sDeX9IUBxaX1A6FfCDwkJM72F5LBxoeNUC8L3ybC8dAV8P56ANPufxM8kD6HTxZXY0q
LLObME1PT2hKlVF24IjsxcRp+Kau4E/sb2Q8E9B1paEgEzbnom7xdNZGLUSfCF08vcnMnlmEWAv5
+F+4rJ8EmHNpbGBHjcxPfTXC33ReSLkbJMKOz2xs3SNlpNY242N0l1SPs6/k1Ih3fyofEvanr3DK
CAZmzQhX5GDrc3dOb5O/8qspbXLjHq1CMYUZgLo6CW5xrFMwYH08hShvwLWiJezHa1T72GuBXcCg
X8rSjGeuZco0oKDFWTOW5u24xb24LxHX6cfit5LZFsopIiq1nfZz3nrudlIfRCTNpJrJQjZ4UBym
WmBgAKYaaGT/bkIETtFQOSBFd2JSW1kCvXZ4A29sn4D/fUV1eWDwynuh2eLY2yQChSfW00ZF7Jgd
yA/JBjDkHQzjxcMnabf3zlOJcJTS0R32L0j8LJNkBcvM76vwRzuOSiL6eJw7WNBDTZsNlnIGpNt5
8GlgcbM1Ed87iL7G8fmAqYPal8TTpS0hNnnP0cUx8PXd0rWSkCFMmxk/XU4jHhrv1nNJPrKo63vI
QzG86eJL5VPODkx+dXEDLscvW2apCpktez18wzifov8fnRqw0fAr7QMmcQ5Bb6ove3Vo2ipfptqD
bRTMQ4D5a2L7ZTUM6KTw04vtI/TRL2tk7Cqtcxxt4unpdK7HNaxL2eBQ1sdbHLFCYrMeEL+No2Ym
iDWsV5drSkdMSaOUhOLUGS1TSPeLdOC1wWylx5n0+xVuB8ZF2mr9cguLpCzIi1h5rm4X1VEAk8Nd
KZrZJNwPhyQLYO2Z0mfawY5W/Ju/0wM9qoMDRtPed16EEfF8rwCbqFp+pk8JKo46KkzJ/pw06pUj
zNjvCcjmQFs9/vuIlbtz8g+UHnDzgnk+UJ6PyGh9QkS+b6txwrZCN7gfWa9gkcVHFv0Ib5Zn8SbE
O+zXdK1+rr4TkhDSrQUNSWSP0qJNFAEkKCHuql/QfIUlesA7gwB9n05VeSUnf6OI198tJ4G3aVfB
kOc37qKhQtdhk8tTneiyKan3d4CKtMpZdNo4z6xgrZYgsGQ2S6RpDgprLZkShnN2NZXgTZnoUdS5
baRCb+FhgbY4eWMwwR7oMmVxitOW6QqYyw4m7uxrvMCqF3h6ni3+gX++zOFEI7ECE3OsRTnkqJq2
yvrkVd0mNbP5x4+RNNfX9TymK3n3Plh+FFIUumiY3OcgyXe+BNTSKEgGiRUSe1l4LOLr4Cypq0xq
nNvHbaVYDFsBt0eakFs6CAjbIGR8VEE/LokSHGAB7n6g4WnFLsnBYUr6QS10BrKeviuPtZzTHDXL
B5Z5BpJMwcc3cIdLrRYTKsEKkvEBKP6dtyk2lmtW2eeNzIPYDFPM/v7UTtMShd2BySin4FH5rhi0
bflO+YLLbzOiEqcIaPpYr9wYv8Wf/dptOY1EbRjnG2HsRo3myWGIVqhKXtON3phiP9EPdCXVqJyp
wB4MM865YpVWYX/m1sQFjM/z8vUhXsvhGXlCQ7jUVxitFH6hOy8XzhsLtwRfoCx4mZFqIbPRa27W
usgcj9BCchSq9nff3slPANpvlfItV9u5nUqe39SPgT5JRBo7ewYy/KZG0jjfjTbeY6KzyKGR0ZfW
OEDXxLX8eXMXdo4qeg5ZOKHiYfHhipr9CiRViUnTK8NcQ0tAqn+BuuKwsirNON1yxDVX3CEDD6nG
8iEhSXX7+C0HMdL+jccLg/XoRaIhsJ7qrhl8saOoyIyQUl/X8D+tDXUT0GPb7WaNn7boXMeNdo4e
w6PmugqVYE/WGZOT2ASGYhJdp3dDwpZZdVzUj966UnlmlsUroG6vYAA6Mntm00gukV5YGXuWwlSK
6+nezCEtYShYonIaTVOfRlae0vyIoFnOHhKJpxZ17bft7Fa+xi4MVkGgEq/g6ZwE4W/+B1+MJ8jX
G67Qew+Xgo3N58HrSotjhCYWexMVku08l67Zb+qdk5mOvimDobX60hi0w+KGLZpMSIUZBuYd6hIX
BMSDSaai/EyhtbrlWlQnAKt0rTb5JySrTxwlrHMAgDwNsjajs+3RMa4N25GD47zN5AboGcqjTPl9
wH6Q8WVT7EeYGXAWuJwST+BACLmvb4fRZUhpiHJSNqMVMKFVdlNvbGSL0BoU2C2k35BWGu7mbRu8
GuFuPEslBBbyNdfbcGjDCKaQ76iUJRpDIh3wEXoBgrdUvbEj2+YNQmz9Geo2bHE/rnj7xC+kZ49Z
A1Shuwjw75fEjhc2wVsd3Kd0mRM6iww9bgSonepNQ24dHMpup9Qz5yVvPeBM9ZOIqD6FqMpkadmv
d7pHH4FPv0YHUui+cwi+GHpPODMs1Li9cIzuDgPtFWjekaRogcu7UxMT/NKC6cs7f6RfleIUNEly
G7IJ1rGQkgdzQ1HmjpisE6ZMU6k18rFn57nIMRGVGuiOEaOMyhbjbNhFxYaj0lRBYd6DfPltqTU5
LYs8tzEalghM/+i1j/mKPF/7vVrgyUn0PwQA3QqDqwX8SH9wSALQsg3W9xTq2UaD3XCALeoPFlKH
HWx23byrj4qFYWTcu1Kj5Uv1D2rv9lItxvFSP31GpG+tx0r5mwAjhafEs+S+ukd4fTVbcRiijZfw
qLrzefq6zJ6YNrK2BUYgb8muG2pNl3WGDHtUcJ4H8b5AK0MiVBX/ac1Rzlr/evp9O3sEchOcyTw5
vsV2KdA2gWFsM7Oa4ta2FPWSeW5FJaldYEFGyYlu6oxxU4kjpNHfhDmyXFnOGNYNJUZtIr1yj9fo
jIKm4FYmV3VTpm+3F+QTK05wJ6hr3QF0US295gFAnaRU7KXclhxwhoohuBMfvuSm3PSuFPzZ5iMQ
cf6KsHeG7t7yUKHwzFZ5wrkh27kkkGWcGhKITXNS293EGOaVfqwt76hCohUTl49yg9tiCVMEwr7y
JdMPniwOCNCwQ3SaEQ87AWYCsrXxV7Rozo49KvHxCZnc9j9WkfL/BjnsmkK7I0vNdBnUu2ixBcFl
wCGGhXnwei7UobRPNZrNZB0sDpTrCmQNNDH1QmmJS4qPbNDBjYFtduSrf7QD0BibDth+qjV9Zbug
3Mc2qQsn3Eijp3KxjFuQI3wJ3f7CPRb/WjOuwLw2CfRdksh6/8u77BR6B1GmEmVhpMz/HddMnXsF
zh2zUKe+bcrtLAze7EU+Wj+uieaQcTzuRvOBKC3BFdCzV8k7Jhnzc0oqscGBcNOGLcCCzLy9VhbX
lRD8RwwRkNMwJGTaSaOrxrYarhMoMon8biO2G9zzv5uk5lhGBhns516AQoCW+EGtt7UV9MVsyibg
8ruwvZA2LXTglasnAP9s6TqnwBThHFts797afyTjKH6xJsz4cdbrZGsmkzg9Jrb3w0bPEdNSNugN
X3h5O0sjuRKpF4h8lHWm7DeCevaoTjn/5NcYVbg2Ns1P1ujIkoDjomCKJ2KcaYH/v8OdMKf8v+CG
py5Jk7Zrb2aNfO70hzSMGScf33CikBAFe29Gyrjyi5BBI50y9x9F5O/OLfOUtoSFr0AWFsTqIFS7
+IvBKHxyKUV/8whjhWtrNrd1VRfN8UIFnvXhToVjPhRO1TP5oZrGLAZ7+MCDrPSuI/vprWaUlAOx
gkMrx/62JhmqPg8KBbjH3TRdbMgSSvJTJIiYWXooVzoGNCc3EToUfhch9VR5hYc7pLmn8Z4VW68v
2Yab/yRntapaRuykZHjHgz5iLdOFTE/UOtlZBOQbSK6zxBOJK6+tWa/MPobN4YhORT07qWy2fSCJ
ZAotf88b+68Ib5keeZbdXNZoFLSJqOjTiCTZ3KEEQa15jgR9lykEvEgUui7ykSnWQ4IW/veXZSDi
Nn5aIYJqpKobbpHx16z1iNzkyeOpXdiLsAoBKQYNYyEVHL0qe/xO5Mo790E6QMWHqliVVDt04TSa
ySM3z97o+THPLrSiU4bcJBsqeXY9UBJGdy5CA1kmSXFerR/Xs5sdH3Zofk0Bwn6roxBSadFbx/rG
wVhtZiLRwYhnpoPiIGc+TgrFUp5r0fBQajGoexj65S+B3SczqsSFwXVRlO5JW8a0FFRu+DtvQUmc
ETRAF40Hy4YIoBzbugWVczVdj9CyLRhAqeYT6fHG4U754oE0JtS2tLG3OtIz40llABfalUs/qfOh
hGzmTnnyODvVt937XCtvkMLgs+2/n0zljOESmdpzjLgQNuWNmngdWk0uDqBpUKGOUkFmHDwMOHCu
eHWSfPLXX9k0CqMiYKPS3Yzl8dWqS9MdUBrUnklanAx0avcUs+Jxw74Jh1UZHGxdf4R6h7qcK0vT
KnGOb0GrMEIPorbiFtCgVK6wWGguy68E3iXs91UiJ2WKgujuWpKHdZkwhZDeFAxPBAOrxfTcAWwY
Hv8og4cJJxVPo4EFRmcRybsDU6wb9ou7H3KDAW8P7k+EJHA52AWeiVRvXLXpd8v4lD8GGjWlmOIt
XjIkdPPciLNlJnGk48AQ0mPYXkWj4smMlb9Uz5Ux/VL5Fl4ZpmFKV2XfXOfNvPWjfZn92c1e5zZi
WfELCWo6o30MO0HjF88OhZiAgTmGvtKgx9JjQWrsDFILkR4sIIwsHBZeLM8Mq5mWHK6mrSL7WHFa
7JlVaxBjzNN/BZiI7tir5cqQS1Rt1h9ZkYdlHInLxQz85w0s+tcD//fjmU3Yn5wQT/MRLdbrp6/V
KqXws9bzwA6KAcF+yseEyA+pk3TIvStrqdaMyHJ65C6wxhrmhN/gi+7z2nacvwJYyDDnCPaJtf9t
mnfEWGNzHRq2TaEx0OoVfmum2e+No7aXqyFjVIK4APPVWMj71Xihm6QiLAmv0FZuQwmEYReFaQaV
PW4pz16TaX73pki7JurgXFzrinpuBT7GG1QfRwMcMhPwOiPNAA4BUvfeMxNGT3A4/ouS4rjmfo+d
dCvxjg9EcOVeZxUQsgd1Pzyd0GySN1tMw1008212hKai/gSJkv0quqLHgAhErP/NP6yvvD0DA4rd
NIOTVA7zmdyx7O52IFEUOiy2tIUB0MFfygo2Fqw8rVuAl/txtoSQN8hVhd9OO4FjJH65FClOcQby
V3EXTg+mciZ4N1cuK7adSPIZshiH7zZ2osUbpQTWXOHkdcUDes7ETwEtqTTDgibeQ8O7SPOyWUoP
W932g932TTKpCJhuDecEGIXQn/sl3g0dhIZlFEJnNQyMoXm1f1ZtFwFeG6jog6D/J3hc+nrervCm
A8SRXeXe0jVKVu6ab7MMbHS0HPFSjallnwHhr/xIRJWbNC5ZswMJ2VwowNq4zhdemu/1mfEdwUx0
7fWmdFoA0LNRMmmm/2c5e4g+v7KYPKKuRXRJWaFT0ztKeeIORt2V+/R3E+8q+j4Zlw6D6MnvVxeT
eugT01JmKKE0EElgZV1N1+eOyrx/7Eek2pT6PNgyPfKGrAIsTg71OigSrPI0nxHMx6pEqrDtf2ux
+iCWU6ob3AE8j49TjUchzX9JbIP2sj8Van0v8ElDYZYjcHIX+jN7y8l+3TjLjPS1jh1fEyEJRNj3
vIxeE7v68XaEyS8i65gkK31b0uPK4eStBV3cZypT5S3+otAH1+DEunVTvxUpqdXYr3agPc179ERW
529/Opo+JPt65Xj4X/PcBSKnznSiacf5xUDc9MNmcdvjKt79y550kz2Hm235Z/WDlBkjuzXgK6ng
wtO395aTqPKJCG0GHVECS6Wy4SksmYPa+0jTpncU6yqhikuYMeyzIFOC+iZ6CmtRj6OGMxKduAfr
S5fjSotx3m58YSUfdWQMn3NLM7+4HJ8bA7JRY2h1TMYkIYb5fsuxiPlSymPyTq/prYu/BPX1+x7j
wSRemR6lsfMUDh9gOgPON29HKrkoXvos3mih1KSVCxmkmcvxC6B9iLGzU2y6r7hFZ8lnJQFs0eRx
RjfIXuD6yBwVcSRv61uXmVCs2f8h0GugEjMt/xVLe+Ago3J93U4gNMsPgglu0F7M0c0RSnvdECPU
/0m6Qt3M276llBhJB7ep4aW+rzWw0GtrMm1VDczSI318GkSswSlVyo6n1pXwnNA6goezzpLLIljt
cx94jcmTxsfwHpMNgvWx4JulkJGcaznanRfTPa+QCyHb7Sk7YJ05ALfcLE5U9STmpMlo4ar44rxW
KrZFk9GorZgHCXBb9+7s2Xy2Zr+mnTjIOFi6Vo7coPKgHyfvbDrd6mn1iQpCT6RmvEo1OsXRma+Z
V0o21qogvcCPPpuz7tfhTbNcL5MmqS8jJAMinuxmT6O9yjvogIEMCUKD8riuRiF/g/i7MoLgJjOg
jDajxBYd0nkwwIUqU2PKUW+/cKuNnIi4dtUte9adaT2jq2TqPYPO8hzlxnXSTiWexPewFz3hHWZt
AzCpJfSSplpHxTPW3MvmuizU+YHoOdG5L+1GHCqHyydV+pjlmamfFHp0cFYsEIdsUAgzCzZpYOTf
1GMpT9vcf9qynyfYULn2zlfvFT5xDoykdIM9d8tG1xi1HOFFudX9D9DBL+H+79XbAXKlQyExuEh4
QXp1Vhkx0/OdvxBFBKvZw6IUrs1xv0L9xUeuBouo/dv2xAxWzVaAWWUksKcmDcWVwgEENBSf/sNV
1Ke1cGS9SFboOKvMN+1JN1e01zpYVCFO9sT2TM6Y8dG+BntQ/G93mTR81gkfpM05NkISW/lbquKz
pI3wG6ZdpXKQNjmsYGzQMFYUm0sDZb9CzhqMdZZ86Ucp5kn2fq1mBIZ44ytoqHAJTsc+o/zdJVaX
88kP4AL81H/CDaPHijJgYS4mKTvw4iJ0jBAccNHyF5LY0eZR6wlIirljSnlp+u6z55Ql47qWjbX2
VjOkM+KqhByaxVf6emQcH10gAxbQGgGMMZH17Ft0Q8ynEhPSeZeZSBnFE0BC7SwYBc5MVqbJhftV
n5vfbzFtBBqMpDYzRXJmlQnyQzDWTqh3TGClcBROZ7UMHK9+1/7m3bg3wngVxCb9HI/PM4MqQRAJ
MlrN5qSzUVY2qclBq2++SrTn2NbVC3fEjI0KyVHMPPNLHcB0QPcMgBwMFTmTFiU14zfeMUfB219V
LRut7vLiBwtLjS3zRaJ0mHMl62TTipK8zb2GOEkjslda1xNYB+p/3kiVihNMsFGLsHedTo0spbDM
aVk5S5yjArcjHurEhTAOoo2It4hu5FT3A+f6zdzapTZpD3CF0sz8Iap6ZCUE2T+0wjreyO47mBC4
6NHy9BDBp2LAgaROY8Rw6ViIO8zwtPCYoDcZbmaYKnpdAcTUqnxc9q4rRV11+iox6AvN61hqpCLf
IrmHEK9CLnFcKnQCEy0Y9IRQdYkJmpVsZFs8412uDpqd8sLQcqq8ZGn5IEiTCTG0eJySH5KZXEhA
uXXJ8FcoTH51cgIt16gHFZAdVnP/uyh4X15SfAqbxNl/oIYWkhqXJ0yltkEsfGRHOviqvfBffW27
Y7Qd5t+7docGjaoYxRCLAEW6tZmWtyAGkBX2QwaiL95KEOtEuxOtTc5o9mMuzXiQ15RP9bJYZ88A
1Dwl+ptn8+CFCT1s8ODqvczLjqNmSvHEiFHEwlLN51EhyZ1GEnBCmTNdlCJNBqs9aWrgCOd7cRuN
seOKoSq3NZcOlBDDPIHKkaimSpObiKqGtthlt6ixn6C4lBY7uNPdt/GxuZtZPH2l1KH0zzfKMnMZ
VU7ATOPeYDo/oR10ImFyTXzmVtkY875I0VxTJz8tD9UCY4JPNaLTNJGColY2Qi5BQLfowpoY/vjf
1I07/By4R+7LwzMhBPXMzWBJG5FNhm6uc7kgYm6/gHgFtE4GHtTQUKOeomzPO4nZ0R2JEMwGncAJ
xDqYMaR0aqp0ntmH3CmXv1hGr412hpK/FUB5a/SqzQAtKjFQl2bPoqe53dBU1cB92J/hJJ4QRK2L
dWrK7mkK29vMwr02lqsxiyyKc54yPJ8ACK2zMR1I7NLnsJw0fXC30FD0K/vOWHozPkMdoTwJjTyF
vW0sOg/ZhTpeoRZ5/kKa/uamMAPaVkfa36BYnRvcSal8reNw6Aj9l6ZwvK/0js8URdHrmW76WUM4
lCZGva9dGw8TjYoZmtI5ShmPD/fji8u7zXNcwNrz/chCyqaQosHfX5uJNb2zNO2vGGmGdcrJShNA
dAFor2f0meJIwuQ3WNZ6wHiTyxp7qV+0/6zWkS+LTDnqKMLl/eiUZbbfehwNOVauQqdc+oSBbDqZ
SPerPC73XJ2YAy6xhbL7glMPquDqnXakADChMHg/jO0+SvfIsVLZ1eaxv1ZvEgV6EjnbB94KD/tu
+CKACxILRHiu4mgbTrV1l0l7jm7plLjxZHXcPKsabZaYalwxdBP8F5La+EjnMdoUex8QX8Y3Bax/
9IjfT1t5eM5Fg1xU880lLD2XWXnQB9OmaZxIh3XoartgJC6zecYQGJYr2qYBP+1MHJ5ALlX3KhCE
Yvf7GsKUsIW7qXOWaWs7CGkvtWiRXhhT7G8018ik4oaI0qIh/Cn7jPWS8w3eKT+i0ux3kyDl/aJb
x/CGBcj+BuQONHeHg35+pPRg/8SD51YQmtdF06xYe3k8RW68mMOLOFWBaJCS416anD7bDVwZxJ+L
qASKbfvudlf9TCWzfVv1D8cVXC99cPNiYMTy7naaMdIlh+CPQWKP1hq7Pu1A04G2DLQlEGOoabmB
d1cfvuhENaMGaAoljbLcSp1VSBXK+ZP9QeDkQtzPZcCike0hN4Uslhd+nxg7ekbTDVhBM18k5Qks
voAE0U2exKkEWzkiLn0toHWElK/BAlMciyHDj9FDZsiKgDOqzmuCWiF9InoBv05fp4cYuRKDR3Mj
ukNfeO9EHyH095YVyPmHcpG4stJg6vQkq4JXoVYNeyppHXFpYATOjkRbTJqjJeJ2EMhN8yK2se7l
/wnWsawTpBlQPwAEWpRDrcTqR9rTmWWqe07d8ddTd5uVpZkVGmQtB9Af9hKf32lO7d4TlwZgXKvS
S1C4zuNkyYFjXsV3P/dXH+TfxZ9JlK74n00cFZ+hfld/xQbEGhKi/bnS23NJqtpY3NZjSrOUdQTC
QtH3J9JgW5+qBxM1h9j0iCQZUpiTPJHPsefxgXEm67ph9G3bX8zXKMi5Y30dMLZJJRmDstjFtWzv
j+Q/Ly/ZgUQTYhXo+ioZwMuyc8WxbqV8xmpol+4FY/fVxtWxHgXnE6y08/+ltJ+u6e7qX5WU8dQZ
Zs4468LDe+TSSaJRsyMJe7nudJp40oBSNsl+DcbFVhzW622yYt0ixObW+bd8GR9GGx/lqwBHyKMS
cmxq/YJk2+pdO1URb/z24kNp/jIeMc9rnRxYC/ytAtfvJvyB4jbzH1PPkH2BQDu+zjSk3hA4QEwo
3CRU+RaXueTTTRlWKm6xSd0yoZDKLl4JgsZG7ZCUZebrmpMrmPIh0pxScYX5+G4ESiJNzOpzyOE1
jvIjgbFVJfVifsT1VUS5iMUXaEAKc/ZAxWbxrac8pyHPpElFGtHVDHqe/8rN5zXJupmtET4S6ndw
cfnTGZrwU1PM786yxX+Dx6bqtSL6x+0TRsVxal/Q7fRwOQa48A7qyZxWSIIpRVlEQlhr9B0TMfiL
WLbnAeM5GtMt7K/ZCGH1nGKCFs2zEvX6Id/eMpXcFyIGtDzAVz97SAWP1uj1eziQtlhwNHw9p6Xj
Rh1i+zrPhdi9l0kchAIcgDvYJYjej8t7xvB2Gl5RgQpu5vM0ivxj2DP0eSBMcnxJ9m7h8QS3Ry26
pSTCRQ+eKx8X5tqXJ3D+J3Bm9rPTKTK+oMdej6AsuEROPrP1V4RrXpiHmk9lKueYqMdsa8lvr8qU
BDx0u4RiLixskqI4Ngpob8PfiSPvSU/KOjFypayQNfA/nhGmDjfk02Dr42r92lASBg2+uetfxWLZ
fnukqZEBYDF6zsxE3yVxcy4WhgmurmH89fCbJMW2R1N8jJ0+5dqlI/ffWlt3UL7GKjhcedkN45Nt
i7ttWGT30V1YXAa1+D2RIev+5YIuWHplXqM/yC2Cp3BKKAvDPwBZutKZbnWZ/678kbbE+tSzxfZ4
039tUzdnCkKYhBN5T5iZI+dmmv+ha6NUvK6hWdnlTjuEaShK5jaBqAwD/ZPXuU73u9FFO/dM8l03
MBmSDUevyf31BA2MMDkflS6K4O99YBgL8sx9Da/SRvE2lBUUU8BMayELfsE9aTj6c6psdGxi82gE
nAHOsL3yNQlo6gBtX9Q6HH4DY1zPufo6tbynxZH7ScQGLQQaeKY1gS8mSe9+SqK3JVlrGjvZVDmn
kFiEGzzzLoa8fTTLsr+rZvZNpQJvGlWuRUGzRBuhiHG2+5A0lzx4VEhvbQ7vVLieKM9COPVkEsNm
9F1g6oLf+j0w97sRjtuu1de3nOicR5FDmo7f+SY3gjsQ6HL86999NdKtcv5Q/GgjXqL0x4XxBN18
W7A8kLWI5IdtO8YVnVcjJABznQArTxhYODqyOFMz4S0owdTd3tztbwnjkk078osDU3Sca4CYVMKn
xKtkk6/ED6k+ImTPiI3VoY/pRDgO3uycsPVNeZUbcgauZRfxmuZiTGrZf5Vwcv71YQ3nyRDmJ3I+
vxD9MHVm4qG4p2FM0KxijC+mwTktkF6S9n6o/Yp+IAbn5rgA5Cw/Ls6zu63eafHQzna9W151N4Jf
cqrBMmVrslCW8Ebahr44WFZiDuUUn6eiK+Shbl2Gpjnx7L/rgjIJkiclQNYoSiZhVrhNpA9m0QAp
Ho4JIYJ5UgoPQ0nAXQZTm8OZmsVcL/BNJXxVWk9NmcmSKX90PgQ/DRWehRzszu/ucPDQ5WDjSOW1
R3OYaHsL6IlPB10HUk5t9qXLWtSOA/ZlednPlfg89/2f/8a4T1OEo4JmN83B2uIFiz63KrX5cHa1
enkjkfN/i0frM0gps/2FW5gnUOdfOnKBXget/srZAdM02XZDK4oZSGCKVhm0g2Vh2fD7PUvWTr1k
0XRMC5Iz1Rntp+TsEKQjUblp8M17dMNrPt6uLXs6nvOeqQ/COhJMKXKtljkgKGPQ1ubqNsRWhd36
ZjTwKPk69NViklM4CQmgZBcPN7IQI7FW/2kczg5DyaeQWLx7RDRHhnvEGJdfYKh+jRVJn653RXaH
22kAXUFqMZd+5w/L/hyMEwEA8ahJYZWobth0QCBksg/QKz0cqE4ks2D04yAHo9fb+IEHsszri2Ar
yABfvQK0jKLdOtrp9Xc+283VBnk6twFr05OqWQEFLF4bWKYGrLRg2ARFSkXiWVEY3R+WhO1qBceB
8heidnAvti4164nyMUvEE1Cfkr/hQmmpmrxsHbAgt567BMYvLOR1lYt2bjba8r+17S1tgOI2t6YO
Ff6jF8EkV3rXVtjGpIA9nvLEk/EOVWy8t84wKnV4bGfXAF0IdkFqmA/sBi6raQBe2BjDMCFhL92W
Qpe9WNC18QdzQO5iQnXj9IEjWqrLPIJFbbaweouDr1Mzaqms3uBPYu/5n6LpLjZ9T2FMOpZOfss+
8HcDKUPYBnr+AGlNjigHYA2UbjKmVY4Su1pD1avEEOUBrE/V7pFwLjDcA/6BhNGEdm5i1Rxnw0BT
wMdclploZDYX6N14v3LFVcDDcuDD/V2kSjiprViZ0Bz0Q2CdxIs/NaA2YGtFoXJ+rmXxgwzSyymc
BjlcjkRAtuO9YwmrtNluRx8gaZQlwewygh5ZX52s2x10HDApt/7He+soKYf+mgG7WYqGBz5yUIOC
Oe+hN9MJ7eSzEk0E5rk2E/vq7ATkSlQvxa7ztPLJ6SHN0pW/QFqSDTg0MpUe31vw2u3LakxfvZsX
kStwJygS7HPjWSIpbGul8UnSZXvoGbkZQSaAaUQQfgL5bdfeXxSoiJUVZWkh5D+v91RqtlwH+tta
Y2WSGlC/a8KuLq0r1adIUxzlPp3+nX7cwnEsZ2tQa4yUPlV9AqQID+CkDXJxbtR+jchV6grtjQHI
eKoM+lMe4MNrHvDKlMRnxoU0bml/aSI7JI+Xkb/dVuwnPbbU69eNCjN8cGo1CgEe8Q64XYdyT1z3
0QgWJnxnt9B0U4iAN8q7N8f5TxE14iEHWHjvwko7DFilZxdeZESed/DFhIOw5pXMG5Sf6m8fsqub
1eyrRPI1canyg/SL+3aJ0JcbdRMpNctrcU/VT7dX4Wy0wFAe8zPZKmlPQX/ZLpKFKIfCOLjktYX2
eEYepaKD7VTJ+0MguXBVUcuc6AOkNo3Ryq+8BIVbQpE7Na4kmEI5u3+pZtROfAu8Mv9k6DMNyb6Z
ONwKTp3wY8sysrKOLqiaeOxbDXU2MiSkRk/Vwczyd73nhY5cMqTOLVoc83MgaO9U2QIoE28SZwd6
GGLONP0r4xfImscEDHti9wZM9mMbFNferlPsEuVIP7oPLeYABFaoTua42C6wuwAwAZdKUubYoLH9
0SbAWCX9nVX/Fp+SITnYhvH3PiVJnPcbt7ZpEl5gArmb491p3RWSI10yH7uOR4dpnxSHIohh/uUb
dCf2s3tz1DEcR2AB18ridhsugQk9pOnAptqiE17CY+dbSNy07VE1oCcNb0E0JQbryt1QM90DMG1A
RXrJrBRaTqazG3mRlKuqJYitBYOL+0hB/vIgGpfjzWCySJxUVBxlf5iXZYvYGSuMdaA65nBNP3Ea
dftia5+eYLHHE1Uexr5ye/W5fPhMAbzgFLm9j45XCeTqAZ+citJE9Qwn8nDi77Z7wyUqihixoiCU
mFT1LCwlvCKsgp2riN2StRx1GJhNrOlniz8Rszq3u58P11NI1LHVwn7cK8cGc1lP3fHJV7Xlguwl
IjkvbjQg5yjxArwKZwJGc3YSt7FBLsMh960K6Dx1a0yQCnGxegsTgIPJVFhfF/byuZJNPNoibyVE
o/8F2jPFDZ5sa4uauYZIFCrrixUJtH2oABJHCs7VGb5iIMf82aMppw2MKTKK87RPPzon0+su9MjU
SQbr2g4DfL5DIN3fASSbVQv+LgUU+E3wajBA6pyPLZNZeCzF23PTdj2iFBsOaxr6XHkzt8v5v2N6
OXe7W4+p0LJ4vqrzBQ7a1NmKL6pdWP/XrKHOfYKJFc/q85K4RhXQGwjOTvjiSTSuYopoMbW8KisT
+qHHQY8FlkZBrdiWA0K73mDn2tcplcAK2an30AQYAEz/8OG6JWX/K9mR0Zm/dlqu0zv7Dx0PtwzV
RA5J48JA377nADImQtxF+8/M9kl3tHZzKePzVx/2IKneGfDVYF4sNNM4bTWuQK/zltVTcErTh1hz
FCQfNf+iR8AhQgFvPk5pWMSBp/3p+1xjyyUq8LgFgtb4pQ/zeX+0ClPek36CX2pF5/Dz1vmVG/n4
g/23cLCnQTiD7LAQGuSQVhP7j72rXx7TARaZYEJwPVcmjVmZnkHQm1nxNs38RgM2AyWm9YyOaOgi
DYGgBjI1rnpoD3LxfLye9zW6ycjRPl0ixDC7n84eUKC8+qqAsTwADZV0SY6Wh0tSBf1QekampSwR
4mSssC8xIaSsGJiF2z3PAeigQH8A9i3OFyi9E20rMDuVthw6YiFkRKj+usHuFOvkSLH1vSL/hBt2
cvQsxIx4CGBz/Xhk1AhQWfA4i2euJNdaFHgO0KWNE43Up4NrGNCaELRCjJ1nfCGXKUAE/n35FsT3
S/nf9mu7mRH/RHNFZ1ZJC+0C2cjz1HMRpWMHL1tMO5HmmffKh1PUiY7HHzR44+++FLT7OMccV2Gu
O+mc0YLdq+oFd9twgWPRP7o/emlqQ0jkOKSwHjzN8yTSPuRDXB4ix5CYIbaqpfDV26fAoBwO7zeM
9MwTZjUL/m8X/DY0NHlFqaoOvWQ+YzWIRNdwX2L65X7/AYpdW3VbMiCW7lzABQHRd/GNDPsPQ9Dg
h4nwqFA2PnzmXcggBmNdU/dlsb8tno96bHY7g7UYTaOiNqtKUUlFyV+1++teVJhqB3zKdUfJJNWS
lzSPGiv5PaBYa6DMZc8QIUjSxXpGPtmcspZsjBVk1ta1Iz8vz0e0yvRYhleUKGtIYJOUEHxNRSew
R4wMCiJYP9Zp9hvz13udzQiLfMiZeKBL4Zfb3zEzGxxZ1FsV5wGLcjW7DynBJNv8XDEMf1x4ms04
2GAdQUMbMkbQfK2eIFoXJBQ2aV6zE1CP4I+96dfsdpxxiyx1gZ5a7hCNqCqgImdiwA/MRZ9V9JX7
fo+swBBIumdDxybE0c/aGC2PZK/QDzt1Er0XplAAvv0MnDVjyvX/XOUbn5qS/f3QbA+umRJlMnsI
chWnxYgjkilv8zxhl42g+W62CP+cMGCmwjRtfftHsGHWS3WW3gUk+g6uc0b9GQxS8z1uOy7Xxd16
cynrxsMqguF3X5wn1XVquElkfLhUab5c00RrH6U/+uiNh2Ww3Aupz94w9wLABmAbYwltk+gdXvdG
vTkBIkApTgyB6+17u5sOum55wVWJ1znhudzPWehOxGmwqLENrB13qWZf9b0CYlxLw3S1OPUJshuK
GlXqkuX8t8i+qEQkpI2TtYAdHR+lkxYTtBCl4+YlsfaB664EQajfeCfWf45/MHt4KcBsj+o6ahYC
SN6S2c5UVTndBicXzuMuTk6zhfQHwGJVfxSYGy6764089BDEKOV0Noik/F1UIeHj4WRMVm1A2UuW
5YtgrgCzBXlwqHTDCGtUFmI5voD1mgVkAN60n9suqT1SO1oEnqyqTS/LUGvK6Vzf3Zhcoamq5vdY
lgagmhIOANqxppPD3za/PZ2d9RyulT1WPhEvJzZKarhHmWjo/wS9iJ56BlF75znE91IE9Z9HJqsh
ctKgdcieGjOOIY2ddF1kFzQDf5TOYHFvbHkzDfWRZ0ldCsZekiwF9Q9d3yJ8alHIoLBIKD5qTiqR
GnRdIsoQkPLq1VbRC/3XgHTfmdSF1eq/AbdVWEvBX46mmizMzyB31QQYkCTTxWT/KsywYe04MqMs
ToOZpUebizU4hICkjupU/XEuQZWDA3rCw68imepjZp4kKwQ3kr3nteV/TD9gGQ7ePyCOP/PNCiyk
8uYiQdkHIcqGiSHAMRWzCoroODtuUV09QpxzIuVx+VEElG6qdmBXPVAy+lQ9AjDtioUG+YfJVvqH
6XJTs7UAHlMb37gIajPsQb33+vZLSKXpMvVYqUctkDrFRleZgFKYlmBH07yz+xJ/po9AlWD2oDaT
nKSVvwsmOEu1XeEGqQEo4JdDlBsFTUHBtn99woaAeQGy4v5Pbxl3s0j0hnqxeDHD2oFMWA4M7WAt
9BXkh9xApKS1H397msNlcKQYSY49Si2YwNRDV7UtXnfN0ZDrKYxeARFZ84aMywG26IybJBtZ6v5i
kY+sn/OJ8gf98CFhhwTVNL7jp+5DmaDJ74JqoDcLHsMOGKPl8LfIRpi2dYiItAWXqVPrgC5i5XyS
jJk/QIJQtYdfQ7zOJVa4a2uOeHGU1OhLg+Sn/Qt/s1//mUZJL1jh79/DWM/KGMCI9MKBMgSszDYN
j5IF9eDYbwLfG0THuCnMtO4BVWsbmpsqyJffzu1fzMzN8wVzqSythklL5Jft8InKbuhJGgg38qOp
PGl0nq8GGdVZRZ41UI6x+MQuIzcw4OVcVUSnCejcf7q0HL65/hU54wgd+3/X0tC28nls8YKyXcqz
SA3QFiWWzdSz1s7GhKG540tWlF51Prfp8+nU2xTQ5dEac4olC+KPtgO66mXYDPnczgX/X0QKMeCY
nsllqWVtumZ8zsRSYDdW0hT/uBPCEDWM/sC72sSHTIfHNBh1xNbZmhXek6sscFo4teJgJo6Tf0iE
NFZM+wQWAh8/7nbWLgrf1OrKofNbdbN5Tbj5upoqkJB0Hfc01ot4Bcww++jKH1eOWBqMzFwDVNFp
awSmtus7aKeMEB3gvKxmtQo+YqOPnL97k2xnqiY/Fl+rJRsbLJlLdnJ0ix8wywC58uZ2s3Inidan
+zUm0TfIlUKGmlPHRNp13gZ7iI8QDj9z3XxXe1K41oD+witZrwfofxxcQgsGOK5mvLkN0/JUN6n6
1UdgtQDCgYY76hCqHgWqyAewLUEWb1R/o+wo0/iSMAvO2UO6b+LZjZkdxDZJOFxqJ524sZJXzG+b
3AcSZmvUXxmtVJIRnAAe6w4VMZqGm1xnsuHjUTNjotSQUVB/11uLYbk6jupMtiampY9aI1BhhwbC
x8q5IX0A1tAw7w4lBp42MP2HTkl/+cGN1qDKmys7QV78qkBNrTR33kZOyKuyX0QaD7+JC87Drt0C
rpoxKP5j47Zkp1BWM1ttk5wAJ5dJwJZEZRVqu3UFyIIkZQB/OlserH0ldoj6kr6C0byc678zeYVo
JONi/PNG55Xk79hJNvW3q+dgIzXekqmR+prZvB9R1PdFThR56CqLCgja93JPvLHQNaO8dW4e1DT+
j7QQLVYuoNoKIkUEB+HYptsquUCzwF1dxieE9P+g3ea96ftRBKOWMcgF6STTBVL0IvomsMQ48sud
qX5N7UDOGV8efF3F+EMO/vwljKhNY0RfbyHURitwXFJJ7Gm8gGTnuePxHwSzjftblDO1xQb8a0jK
kSuJIOfO/bV+oUpv5CGYVovZsDRjU6y71xMgzTIOINoGMvKS7+aoieZXyN6e3rRR04Uhz6MJvlzm
6klvVanPPEZyXDKC2/PQxGqz3QwV2TqeZwRHkW+DbHGHOJXEbJnjf2yMZFxwwSzMLNfNzziYAxGw
8u4byfp42BLUVK83kHJOugKS5T0T5MRaLiyD4XnEcWzR0lG9zDyZEiNW8JxWjA06FVSk/6dr7Ps2
yhj8GowARkwwe7zmJj5YXeo8fbOX1C+dz0MG6JssCQD7SDBr6ABvAu9RDb2+1ASueQVAYh3wP0zB
xfVtGYs+yzFUliupUg/5MtIX2M57OnbzuY1AIiCet7lYb6UaZaMZPLbDhuJFfiM6gOS8v9VdRIMB
O1jQnb/xAFd+bBvABHsupt7Tax8/lDa4P1wi+i4ilEr3q8xBjStqPDteiETWK9QIZtRTfU25agsW
IE9plTAHq+4vuaxLa/IKVj62vcGZHD19haZsT5c1Jw6lkmq/CgZualoJOdnTt7c1hc+L5/5dF2kC
rvyufsoymxmY0fNizhbU1CU4gocV792CDlp95liH5EX6bHHQR3aF93+bqZ7DGAKUmbxpz6JWCUM2
QmFOyHUG4Zk0LiAhk4aMem+y70PZ2CiRxj10xao6Y7o/zbXNk1zoY48f73Am8yJqcDeDQ1cwx8MR
vWIoWsyq3eSv1Ir1JBagm7yxgyK3tMuDqRDFGMCBi5SAU3R6XfdZU2O0/whPnOKJt0HEhLQyDp84
nvG+Y9t9N5uFSLvEjVnRJ7O2UrJs9DS+vhaSfZdD9W6smb8RsgkC69laOelqlMTFQPfIFhzVuX8M
Wih66E6Z4iwqn7L6dGhEDDfEpIfAHDrQqp/t9VUFgQHE2UHa9j3jVEUy7hCWTKWX3uPhBhAgS6eV
t07g9dGJOVqF4agpz28s3Ozh9Ry20BPGhoy6kaeLYgmLMIy2sJUaCuaoJ6EUCvM0IHxVEfUXPpMQ
akkF8Ht8/ngFsEZMEtA1I6f8R7iu8GC8SR3LzvxGtyRDVxY7/nOjb+nGEYYMRxL8apzKqYc/jg0B
LaKEc++FtF6OqwXF/ZwC5SIkZuh2AjRkGSGBVb/437vbGfMBvHYkx9XvUoGYtheZLB2lt3uXoD30
RutpNnH7pmQKZB90IHCfk7Hr0xQh0zY7QbeLAYV0ZvQES/wJuMEehKEXPDd7CLbHZ+CErDE8oojh
dp8+rYMzBdZa30DRmSFv3xxu65U5YI6sqpxUKplZ0c0K5+ntmotMIy2ekVowD0ZyLKfjbSM2tN9Z
urVhLYSvFoPk84kKisxTqIzlN05zxZe7AUabTJOLtqR6vDLJKKozrvY7DWOhktqpV5I6K4vaDyti
Ry/SH7Gfxci42Iz4OPkYeQHoQtjppW3wiND1ZGE08i4DSFFUlr9RsENczv6Nu8HYnmuh6DW18ard
/jhhTv2qw1xuyY2zOkDVsp80TPl0mHW6sC81TXEjo2IevUN7WE3XNEjTjUtoIBcm7laTqmzd4bMP
bKlisTTm1DAoJno/XVhgQ+6AwWigiYH2UTicyjoGV8GpeLCCfwKw5sW13iUoYgOapBBiVJTI1Shj
udefvBLx928EVxXx0SP0Pi/GKJNzia8SuveOo3O7cqi/SwwTnZuxqQzbsFKasbJkZ1NKZQBw2wwo
2fk0UXro133f2cBsM+lrQC2Ss+sSMoTss4exNcezJHylVANUuVStrlnhDRBy6VZ/rRSsDLF/f1aQ
W3lNo+vnMKvFfIGh32KggA0GNjhy3f5gjTk2BEQzaExDdxj9u/VKeyi6lNAc2OhJdPZbWXJW4ONH
UOefTAyz+cwd6ayGxRLznXpidNXwEbUdRO/1Jx6ZHna8OzhMaZpdhQu22HLMULfjdwocIoXOS5B9
mEdUEaY6MNErsBd/jMHOfO9YG+UlpAOOHnzJ8M0izslBMjrkBOznLX66wh1fAOcMlRl7zuj5m4JB
I/dRFB88KniR/I1eLl4FWBuUrSmV76vTc/nKGuiiIOK8QU7LQjrhQsKkMc5DcRI/4ZldnD2ZQStC
XD87nmOc/juzlYh7jy6aD3E21jVD+52eeaOFUcE2r9T2uBYF2nE6GuLIPLWAYjmsi4jsHE7sgG2t
gr3Jpi2an4jsEEkZ/4guwL/xPZRHFiObBvok+UzFhSSk+t0jd1sU3AVOZiZh9vZK8+70GbbKgWPS
wq/nes/JtCubXvqrgyRf9C7Fra1AycMIwPNmlJw3YaNbrPmuLuta05RO5wd0NbkOmjw5Yaz8UyU9
1F2u1cFtOA0QlsJTrqSC5zi4U8vxxbUgyoSpJllYqOnpESXOF8dffQ03vZUMmtYkXQAara+hx7YC
MACcOquXET7p5huJ1HAcVBPG1g/nPbx8V+DBSCHH+vB4VgeUXr18fhUmM1ULabUiQW51mRE7cdVw
32tuALaCISUSBZmrsm9v2Go3YRV9n53sV9nHcdjjjRUBruxZLptOaAaT6//k31QYMyBdCaxAjEN+
slqiQTqgaydDaN7RZm5XXL4L9kRBC3JLThm8BipN6XZZQ9nPnSkxhXjgRe5Ed3unRR1PQYN1ISUe
JG/mI9xiDVWk0d9kTde6radl0unNK8DYUccg58Ql/GVSvgRXiiYPDN/tZ8LuBXqv/VcMG90zi87U
cUTvKATu/3clOMBwwi+s0n+IO9sog90Kd6l3LGq63ObOjSTPL7AEmeZayQ+M7y2W4e9VLlP1wVim
hzuOO68MeyqrDxZx74Kg0QDeD8x+Cjq8RMmrFKTaToVC9pYJemqznh02Ka1A1uGnV+I/LychBHz7
KFafCrMd4nX2yri+EjLpC9VucPAD2HrroxgH8nen5Wke4XsXPwMT6v1eR8nHEgxaFK081V7KHhEa
ZHR9+1bpAhfGNwDr3UguMabCYqF6wyyxkcPblI8B8jZbkQlJgnu/oMH7/6ZkbyfC3W13F2hfonI7
8PdAiqQEyrNKFUSS3psBC3BafoVXWBXQ5sU7n+lHiFhKK2JhCY6om7U/OmC1nUouWJAKgnCEtSGG
IVGsHJV9p55bIwL6phnxk6lALBwBpV8/T53xNp7sK5jFYP9Plc3eBf53O+zc7w9gFNoppdS6OsvV
psq0DvIVcfz6qAJV+28umzCRrbQpErgB11yxCU9IuroCznXYZ1ttLL1SuK1xKPNSRR+rLwdE7axW
AsF1p0jOnovQ1IGpy7hzH4DlhU6/XKTymbt38ubn+M4u2IcvTwemjikjg8KFzu3RLyxJK5SLL74U
nkKrNhyaJcXu/MqmNCAboZsduxt/8pJeQYI3jJ4xHXogfoKG08XuD7ErF7hCImxat6rmaOBH1dzq
34LMw3o2wRM2kH9Lhp8+Crg2q4jlFZ37iiiL1WpBr19teqjBMKi2SUsyFO9LwCl3fwaZRa+K7dOe
3gmgIqUFWHjj79wnOQ94x4dNgFOMzziUeZ3AzhK+jKgMsNs48zRxleAGl0GPMr9arx5agcvyH7N7
d3gApan4ttvrOiCDvKT0GqYsEYL7R7+ysxnvxKsshKsN83ie/P55CZ5On1G7M6LQfJ7Mfq5DOOVR
fvdf94r/qVLpwvLNbK8xsWPJcG+ySCSJikySn+pimZSeRU1tvbYF5oNjbnKgpp1Eq6hTy0aJMaxz
5x/CniWLEJTewUb2Dy3uOdOWzMS53HiBgnzrqm3TFd2mVfgVRyZLdiXks3W5m4PvTf7mAFBpGztG
YY1GIyRfG4awy1damqEtX7BLFy6BHpDDDLSqJGyws6xBkhnF2new2+KvHM3SOTrxz+/R6GPzlK/3
CNQVGTteoGMELFfhEGIww8Qp5fE370OlqZV3Ly5Q39V6jveGfijjy6AOmrUcK5jTjvtK5N6sIwM/
ZpNQaWpTYoMvR88tWhTMoKfwOScDQMq+LPIvKtJjMqCPbZugJ2f5IWoqtNc9FQpG+JxR3+cDxd3m
KzNGspmQ+bQdf3dDgw5eRXOL/GaWD8uh5DRUBuFUnIh4WZCdmyRgHTlD/szQ/kKd88Kpf7R1bEKn
adn74u4KPKawhC2W3rXvWlSN6no85njC+Vab/RuMIV04HVJOTNXbhADqig/AnKIouPa7PJ+BwRZ3
dzrV9CPTCZDxnHRbJE8xiPTeuguntiZ2Gtu9Qln+oSqzSKgwKxSZRYAD9g0sXY/j4KKkfkyYByS2
rXv+QSAw8L8HxRF18SMu7CVSr93jA+7CGIsjU5uO7t915RWMVNMMLELr+V067mvq7Hglp4loBNt8
21cEmcXdGtNwcou8gpnA77lE9zaafmrsW4P6hgENn8Ard/aIfmB+wgTauk5YPhbfwNW0MbSviwoQ
v3FoxWml/lfJmLPPfG3lFCrdilabVT7V7YEqki7k7Oz/aFNquoxeIJZxo/U6yCRfR6wGpP8lkGro
vL3s/ojzgMgSWw1pAR+/ej/flsWkPrzbX4V2fV5eKw8YVVu24RhLLXOxUbvouvkCOWEEJfaQGlC0
P1xXXBZ5cnjKFbOxP0AG5eafU/rtsTsBFozS0nI57T62ZavlyNJEJqZhuar707JmoPcFFp8CH1SY
7d584JtlZkQzUu9YjWT8e84uTz0PoFsQCoZP17k+33VM1ELokPKkMBUA7dUKAqVR1fnZRaNKPCJH
0EMoY4lcr3WTPTJq2gRE9ZoqHedSX0BNm3mYAlddjinBENQVLPBu3lp5eDdHc+tzG3xBbp5BJ279
DSp2d06WIbKbwmTQWF6keiGPUliGuDiFnYxFBdMrfJmZexUkk4iPnB+TZmxhlTs7A1JU5A/quI6J
rsYj+BBdxUSESDncuwf6S6PmXGcjhYxW/sLFXueK7exlzBoqOFq3n266IpXos4Qalx7AaTaJB5MC
5Pz8PAhvvGTeBKKORHdU73sYsfx2Hzzv8nYbHiwe9hOli3D5GI9uLko8aPfxX8olwh2LwmBH7xP2
q9ZhjX5WtSPgTvYayjL+FsbsvNqd8S6H9CWGYB8pFBC1BAZeAuw93l+Ee/PS4YDYsjXxTq+iLB7A
UONViIPSpbuFLiioG1PAwvzPjcy5jFwj9dyFcTd1ky86GLq23Q5jkc7ezd+FSy37RaNqTQrN9Y8p
aXP+cjMXpSNx2ECr9AQYD/k5Cs26weZKXUqJNM/nQLWOksMxYZ80ByrPHHIy05L2acIonTyaXIMm
V9Thgy6OCofDQDCNjlZX12nGFxiWA45RNzQz15hCDNbgP8ViLPPyX8eFEE4/+fE89sbqfO/czY57
EIAjJm2VnO4tRfLdNWYNL6x/+LvWSaUHX6Nmejsg3ULy+vmnvS43otFm/TNXCQ7X6nYHyKB2Yky2
yY5eLCuNO5EDdYfuNejRNrA6CS6jZNMI8Yz6D8I0WlKYenzCpocgAv9vAVjWl6RSOZiA163heX+q
TYGzuJvWR6QgIDYH/EKcgaTokmzjvmT5ZI465GhmFEYdVsIun8cs28ovJAJsgAb2xZCON2OnhmeQ
rY9CMMaPOKjsy+dqGJ0Asj4B6+TyW+/FSkkTsoBNwVNuR0htv+tI6nI42uemlhg6dQxmu8Yt0TQZ
lmrJCR9Z99QiiMmnWi9Z89s4yGkzi9pr3dBnpXbYVrJhmOgyNwojnS7tzEhgtZ/XgLH7yhykl0dV
3XN62UGlszuUruOH5Iwi9UD1n8wubC6+zXTQ3NBS7Q2f/il9rKjzU79vYcHoe+mAJ7TGB5TaPHx1
cHQut5vwN4oSyYDH0jb+sMqtzRuD73Sgaqp2qGPMSq9+kOrsYsKpyCOEP3rptMKFcn36LlebO8tb
/t5JTAVnOXUzd60X/q08jWRvLBfTrAjINV2uuVoHBeIS6BHBQbC+a3aXnquidKbu1rTxQWQDdYJR
LlMj5aX2c7iWRHlPMPC+nLvzDnNNU1GusflzDqpDQC1QzE+cdFtqGSFoqRbtHldoEKE/29uwcFrE
9LxKkFrHua126JV7rvQa6Eogc0/oUO9tTAcp4HqFEcup+rT8477qQZoeHR2hrFodcHyHLeI7eegD
xW/ZU7AOr1djlg4GM08RQ1fNWBdNMfIPr2A4OThufAIJ0UstAUIdOembNUdLCcb8qr0SJK5SZLhy
g8y5eSqO32Lp0EZ2wbpMhaJHeFpRJZl0SIOpQBLw6WIChbD938pPhe0o45YkU7P6Ti7NJ5lmak7i
GK9Os2WgKVZcoa6Q4RguNNohSeuyHxQH5ZSAL2Wyd3wRUGe2bcnQL+/XWPZ3AI774qecp2+Fdaf1
B2uGCqS/oF63OdWyPbBo0mpVISMauqasWK8lPFLhn+HVLiOr/fFXn5bBT+TQaPVaD/J7BKTHRecY
lMiWs9rkqLMJZ7kZQz0lceMgXSKCadWJ6qstK6MAcyzr/zoe/t+HXXrhhDuNovaViusY0aUY0c0X
UsgfWqZVxhSxZwytIyQsi0MGuodQwP3jz5U2gS3Am+PWl2FWcVn0ooHEbCfluQiSJuHaYDVPqm/I
BfNBW5bZAx9WmSpju5kKNQ+7vjqSY1YRy/FypUMj47F+xCJ5TnMaYsDFfeaeeCal5YVVLLUEEKoU
u7xmuUWdL1a2XjnIlAjG1p/CnNMf/8zCBC113oczgIf+hmPKGKMoekVAOPTecV/mZCZneEzIWzaD
Yv/8YKZUPXCZZo1X5RYjAD2f9CzdL2/B08XQls6fvoO3ij7VzEDkQfBdOpzPlMGA0QZzlkJQLnzJ
zdzajLGUpKoclqXnUT+M39YTFb/VvBV1+xQqseMsD4iqdnyqoPn//KECtr8ZNtJNBtFoUF3M/iun
2sSZexqA3M6AGTpbNk53ty2wAjUREDnIig+GAEjUlyeWyPd0u4rsSVZtJz5zQWt4zkLw+jrsydd8
nlCECuhGSp8MmkWYXAR05ydUw+0HOkPLyrl0uGU40tsXgWWd5k2HfGTrcrnqeM37Pgq5l3/9ureZ
jJv9T0AckKJoN3EZaMuwKkMyu6Wd43YiUY9bJbC//UmVt0HV1BIzOyt4tNzCngWWcjc7q46SkXxR
IbYH5sGJw0sjOBAgyigxwjDMUa0ZysSOn1sXU6Oz4PYWWLlX51Vdr62lIvsvFvt3OOtJA1DGxySN
v5Y4WbH3yCqbkjkZ3CRCZtt6OLGy/EgxI6MvJ0+uB4W9/nRw6Ui7B3bJtc4HVfkSCmiWska+Diyo
pQe0B3qiTe1Z5aOz4eah/UWW3ZHm/dQJUZMuQDu2KtQZVFrdYst+lS/YBDV8LimZA8XGuAKDkcXn
+dOU0bjQFc9+T7Aw4baFHIZjFyrzRRI9pWAyp29a8WWrN6aPLubL3pORy43t+iKgcIjlyUjn2zin
JRdSjWePACBqcpISyrbpuchDCGl/k+cxrDK0ku6nQcAMMn2yC4oLCqu5oOrW39mGDcx4vtYZAp3m
v0etkNpaq6Ow6rV9tBiN3qFsDRO+MNqlnCTJHWtMQI475m27r5gehLNpaXAcqTNL2Fqu6ImzBjxl
1i8HIwC3uH/j4o+Bi7O0WgztC0i3jjhwpOVj0as+EzX5WNubpG+/uNcaJ21xNDN4oTcBtMtUHFma
3TGlpKvHARualvOVDhhDuioCLZZJMzZYuIdZwGGs3i96FsR6bvIPqN1H3pXqZs0e0J8M48ZuR9kh
4FEqzEzKeczthVkP+gAEesMop8/duFPGZcJtsX/7EyiJv2LmB7bgv3SdFidZRsaFyMPVIiflikHj
SNV79zOhba8kIAg2psu/Du/AOwgLp5nwYSP/+zhBJIF0eN2OKZuyGxAbOoLIu3uhoOrs++LUDZWO
kxmQRzU+jiweLzlZEjKgVIsM2Zlln4QQgthuD8Jw31XfSXfYH4EU+XaNHWEBvyWWsl64CiykA25I
CBUNkwFF0r+rR8os/WaEz02rDPH2egApuiV7E7PC7Pefs7efItygVmxgWZmo+OJHi1TWOKVbik2k
WYAQpizoqN3Ru6rK8ktNsUHEb8kvPNX9e8pgSLRgk+CVuJeUdQ+68q8PzkkWc8JbPkP2LoVVcjgl
ixbRcjE6urvrXO4EM2YV3wZ8/1ZOaS+oWUTGDAfA9UCLpvScfdB1ay356rgNyArsfg6uUSf13ZHa
0mufqVFPteaAlDnD00SiI14PwspY3AUf0AkZ4g9m0ct5kDVNo9A27EeX298+IEQj9IvEtH4AdZ3j
dIJUWnaMfuiRGYuVXK416kIpyGQMgeg0bdL69ztUsiXUqcMYvILCyAg3806SnirYthWivgu8VSw0
5dcRxkoTWlhNErfWmJ6AGX7Q3hofvkXj7cKD9UBDLH67FCgsfLRkTFqdB4uxYaG5bVYRcxktCNrx
HKMAWr53XQvnpQvP0EArWvD1AmKRixQrvMUArogeiSP/XyhSbh6QgoB9cRhLY5aoCPMHq2STNG0P
qRoOh1jwEKB7K/zccraZk1Qa0Zt94utRzpN4VZt9DKns38C4u5LDxq9RBisuj0olohJtRTdLmGLg
kvqqihxBN25UzX51yXRPNnvVpzBb+pkTSEYgvrThume6HyTOzE1Vbey/X4uGKnqF46fAk4gqQV4J
I3uSjmH2nejD+hBCihOOLS3x8NoDMo/s/gja0+Ldwthlb/5rjc+IXUBaXg0uUG8EUWE2v7Q60GVm
4d1RD5VgesHHMpVsf8N2OKdteEwKyssH5OOU3wS0csGu5e2PCpCWbdAyspY+4PZCIzMQWVdkd7CV
yq0iFcmijSRrTIKq6bnsO1dASOPzbH4p200NwQorYkUrCcAceDC0AE7YT481EE2IHZr2KYXJrA9I
QJUL+xBk6CgUFVFM86FlTle3IZ5+JoZmNpBUob9mwwte/IhgAhVckpRZilt3LrbueoPs2HBVOQ8b
e/eYrKKnxQCEfUs8DmbAE5vqGxil/YKJrlMoOpc7dAi1no38xZcUkAuaZPmrvT3P8VFojq0PGuXJ
jdoif27WHHo35OE14rGggzXvyyEfFolXUKdgYoxrY4nbyOGlAmfpV9xYEiVvrtScG+qiZlyrYOQM
nmlhdhr4dtVQRdA+Nj3NtoCnZPKOtTXc63SciBh93zThNCa5JPSFAncQIDuuIzdQfAs2nCGXVZEq
FjddYO82sTGVzT+wnJ+pKiDo08Qw1aXGgnl/h2b4bV721aqZkN2FfaBXSQO6ji5ay4VGQGb4n3r3
wg7GXIdNAlqEC63bd+fA29t+7idFjyZ9uyY02aysVhzxysl+PMH3kxSI6uYHHufYON1f+YBRtO7y
CfxfEdKyeRFLOhIfi6J6nf2xtjEHJLs0FiDjN0AiVI8lsylvzW9vJNn/IgkhUMlK5NlpVhjNx1iw
VivGvwUL8WB+SmLfHldGRYXlxbrdzUxYjwMd42uH1PRKo2QZQ43HIDLdtf9reWOVDXS2g7V0sM8S
3Lf7E6DrBRCoNPdqZ7khx5aOIGWcNh8v7iiczcDYgMzl5t8b5bD3rQ842vx9QaIIUNCMHP5ZMDGq
EqNqLog2ukLoPuePc/HOoJRzVnwEmRzZH3njrgedHxmI6nQV8tqdjma79sOtqTynkzfCeOkR5M+B
Yn1a8YdjB/Y6TUJoKyB+h7aSkajGENNTpqLI0RojjtiFz0USqvm1MhpPPRHls56wLN/AH8cxzqJ6
m3/lu0DYJQbEOP5/3M4nl7/NlNHSq6A7PaPz6NJcNxF3jB+25d0XsRvDwIZKLav5W3ywtwhHKTxF
sjQ107gO5vkGZxPnDY43TOqPGPOPTKFGW72tIXArVCrjVzRdIcrYMD0NUxqFH3nZtHJ4YFEkFeyS
VDB3TjxgBIzFyzdxt4RY6xugSHd5vo7QsFzuM2xIMgQFoqheeqF4cSYnhN6XFXVlOj+4fLZa5z0T
cmo65MFL/BH2z4zUEZYJgGHQYrTIqlrfK5DS2OK8Ql45yhfTsPDvjUA93nLxR38O8syYp05uuz0F
L4qLRTazD8tNb+lR+ZdHzhE7j0JjXVOHqB5DrK9Ohq3HlXyW3fpfXhEXHoVRkoTkqLMpAUsbnNah
6tkgtWmP3DWZeHzkwzkhjxrUKBuzd0+fDUN9JbJYLTRMvxXJn2BrS8Iq4l9H/12t6Tevu9JsgDZU
J9U79A0ecA08f3hWrI9AiuKSwigQcrDMIO8jmFsmxcsjmHsLlKehaTaXgNwnIICgnnPA/aq3D/LS
A77AvTiNrSB81sY/1SeB1KbT0dWWbIAb8jFvBK68qjPxwbDlAKYOjmAiSMyiuTr1LP8mkS0tsVxB
VkLlNIOKO+LgcxxaH6qAHlq0Is93buLp3ziaHWbRLQF3L+Gi5Idb536BevF80ioRp6c+npfbDBTP
o4HPey6b2F9TYl8F70MPy2fcj4hhH1Nra5VC1Rw73MrdssqqmBMA9tujbfIS5eAjtgJZCkfiadFd
Xv90a7zJHibonBsFBsA1FivmDG77zeCtHKjaTVmdWDfAmrwue9wFNkYrrwkJv/1fkKPU7+rcPx0o
AEOFou4u6HaqI4a1jA+cZDgy3Uo5fsT6+dpgk5QttXd4IOvRj6cgnu2dRTN6DGihCYnwybEen1Qs
10vtYss9yVO/imbA0FEbooEq07swZZ1z719dk1N2EKs+NIbBiN6s5rM0+Rqw5tXWiYuWy4Q1jb2H
6NjRdwO/RocaCpkFRCnQ/uQu10kWwP6fZ+dZdcUsRVzUPW1+BuGb5tQ2nlPDHuVOAko3SmOXG4Ge
vF8l+b5FKI61tJIfiC35DCQKdUOSceQTlgZWBhsxCKTZ268TrkakwBjutLaEIjOE3pRd6Z4JlIq7
zBlgM3RW9X1HqsYzWQpAc4ieNciuSe8ia6AsWJEkAZBMDV91qKFFMlHe69DgrbGWuAal4F2+/rzh
cxlvli5IPOvnS2kXts226ZKJfC/Rh3cVM2P4I1UKoSJAjGn5owQ+wL4CGIEP89FFMH8qqGT12clN
Qsa50CB5yYq+rn9oAuhpgKdZJQ8QKji0lObt9pcF1TvyO3uzS8Z6IYwYsR8dCYfeqONU5HTRHAfX
AAeVbyyRZdUx0phSsxvx525wjXRxw0vZAywy1n469SmJyoCYd+ndOepUP2VO6yptdLcHnKhg06wR
UhF0EIMSYCquFZGuPIN2M4pr0yLCjmucXRLFeLIwYGFtbNe32/FKjwCn/7I7bUwNQ5UztpcIwW9Y
WGwRk9wR+N9VhDEZyTknTdACI+QbXZvo+hD+wx20J6tdsQaHWqAtU29Vgev5bSArQAq3hnykd8z/
f+3jAl10lEv9vmWvLsoMJpzhhk1ZTPYy8vzJ+rzE5oEFpvgPZ27MiUcYGmkAKMejZxQBAyst12R+
b2VbnpfrAP/7qluzDLj7NIKlkVPGZvLm/cZRSyqSevhqCZq3L/uQYLMdN3Vv5WH5w/sddLDTn09v
28tDVDiMcfoPFyuVj+sCwVh4/OovxAFzA1RSIG8/sxevqJhr+KSWq4ejHm46onw8g1yYJOzIpp+W
VfVJRVnLe1/PbpCbNZLTspM2OibcGiSg0fDhMiUqFlByC0n39+XfX1v14AxnBGY7MY3nGVAKljMt
DLNC30K95wuOWELbTOOAeK3hHyE0O8e/XXhMSdgflIHlAiCBrxl+zvB+KbFwJiVyvYl7/Mx9r0o5
AuRR0yOHiHi0PsTCs+L3yYAcIRPr1gIN0qv+DSy0GlDSw3YvkzLSeA17jPq5vHiHTjNyyaACkymz
o8Hxuzob0mRd14YGYZarRuiI9av094QOWIYT+0TSxHxuO24/c4d4fw3dKAbV+/dD/FT7mqpBTVNh
G2P2zHYuBrDYVv9yJKKznlsC5p2GqZY0B37rVh0EHw0+JN21kQ4uzg0MmRlLdysNAV2V8+sWwnrE
DsOL5Il48JD3K4g9y6WxXX5v39qkvYUIBXDz9QUiKCD+Nf0oEHewiMmsxIddbxwJ+SWRlKuSHE09
IvLXNy2dVKzxpowKOpubyvgiwjWxp5DeVCXmP1aUCtTjkIGKiwzOoZ0HnyfyxHJViB7neikWZ7kS
Z9/YkfKadZmFZSmUVfXjBiLppLrvRdsLcqbZtXtMM4X3/0dwFZYjtzDPr8a3L0hWkyTdMQok7RZS
vh8/vOffxP0iLhtT0yYKpe7fygwFEeOPPmgq+nJ1fc+S1GOR5hc3qU1781cV94v7jd2AVFbsctA5
h3tKIjmj1mJjUIbg/GXeyTpedIXwa9Hd3ofbcw11C41KuIzcI7ZjstFVkeT8jGY97hFdyNEiw1hB
pH07UczgiCiBLWcpUBqICTO80oGHtgE9BxFZa6rqF3uPaAMiL2+hOkaK1TqO4MQx1VMhU7KwISbu
ooJ80NdRoXlBruNVGNyPAgxv+fyKJwZl0bSUh6orX8mFzdxq5RRcQDhGCH6KsbUuRcsN5NMBC5Y3
X87GKbU+w+KiAO9O8K8PZwA5HLoZ3WtRT6PHwOw2OZR4J61wv01TcR7oOKnP8J7iCAsawC/e0s2U
l7D/tAtmqAsW4LU7cmxFKKl4RoGl5DeQbXD5P9x96K0pbZXvI1lQ9pfrAPnhJBj+Hmn9qbVeAQ70
dmbt20hFIFjS0oCbsUzHZPojR4eL//XkXQKlIzv3O3NoqxBssOgQTgFM1v4A1G/mq5bGq5bgLG6p
x4bXXTcwAAyQatFg50IxxMU1jAzAwbVcFCUaTQttzwSYTIUp4DBbC1WyI5aFHuJ3J6Nt65aJ6jbk
P4IDxcAGWyROYyDutBhsPQ4+rR61Q+O8zSicT88kr4D9Z2P56+iWT37rc7DzGCjXzvBmPhZRLd8V
GdRWRtjhPjpMdFJkLvryTihMl6CpfBUuttQJjZT6hhIksugJItjCPo4m5vv9+chUczmbzJ5npoVd
TdXgSbvyUm4b/wEcRjf0Aal7afz7wLIngZAbegaJElwSjmGUhSYSp7TigemzfKwxPCLolMtj7iBp
LashKDERb/yXAUNFAYKjok0QmC1Q/OAiOVub8pM3A/Uob6z24eeJbAnDLa6RLd3pG9lvFPczc0Wj
OyG9mLd9T991TEc4kH9Y9A0+VhN9hS+y2NbvkSyBijjkR0tpg82EhGHhDclKlit/uxa8/sTVic19
/GznsvsfjfQQoHjdggGUIbIPCnVjed6ygNrmKILZM6S+e4PQjrC23LtqvbKTJhkWh23PMgidGYE5
6ZgGcJSilgBrVKCqUkVm5AYX/176OGU91wubBCuTEgh3kXQeD0xnn/87wLt3NI69vKsG10iNSuZp
Il4RAyQcsEIVvXPwFT44fCikP6kQFyrkzuovpehvw2cGzz4jMqnNo/5C+uEKNiFc3a3XT53Xtwe5
6JgZOXwnYMI/MSXiBVAH8Dm8ddjAk6psm9Ui+lPYOPkgenPr01sxrKmqECw+tLC9XpAWqeY80E7B
zyd3ZX+cXpHungt/K8epW/XZ+EN1e9cXAmlJ1VDU97YSdqC4p27JPljY6Dr5hmUce2BPsMk7ni7a
SEONz7+tr1sfHdkpxiQnd3ACZzN+xlX/ldDRwEk4w9ABSVvlakb4OTpDY+7O5/Wtn5nfmHdG4K18
dpQe/8X7RY+dBTqhbhWfMh1VeZjG6jBko7uhTi5AQ1aphItC4/dt8v6kiB4ppepEKCwtwsLn8WPd
UNp/xuWck2NqSTtsfiJfQylk3tni5oJDeUUAGGVBwcMgplTA8IN/Tb0Yvyzx443aGk3Ob3p7+rPT
SuRgVrClAehgyn9U0coc9/RpVGhcS+MiY3a9exSzaD4vpkBTZRxEXiPSaiDoe3PsVbjnDa8WWPY0
S/zMVYuFhQFDY8YBwIMggNAInMvcUzkNfu76FNiyyG+ijk0STZ1JxgI8tXvh64LVDXU0IMekD+y3
dmRJ72KSD30YkTYarWLNaZz0ico1dacsZUvZ37X0JUGDKpD6uuYjHVuHSJvsalBwR8QCJzg1B+XJ
EF9EnEz9a9IhOKxrRFXdQmEy5p6bD610EYR4YGJxe8yPfLvUQFdB4Wmka1Pj6JXX5ieGztikpB3m
azN7HQ7Dqn2j66WcJqzez0MZAvh9op6rqxYRTDuW9E01PJZy68ObAPKr7YOUWdNX5I5K5PRxnrYu
QHZKsl4D+C2ceEiOm0/7U3W2CkXxpjMqJa5yL1YPACdFMfM9Upl6ph8hH8RquP2+FJlrmhfxqW+4
Su9Idggtt1xixPBzyAhOPwoF3bLjAKRGwEh3ydXOSpHL6idjmb9nCTTviMVsJT6bT3p2yPC1OSMw
Ld1n83ydIGQrGW3O4R2JeTnegLBHkk+2R2waGXodhDtQKotu8YLaXmoOzgZpCP2+64uu0KkK0/J8
k5UG+ygW+LDIEDWnKVxbx3q0IxK82mwWAtl60zdCF3+ZWusvZnaCFTOKlFcx+gNmD1W6k2NqyX1V
RAJVfCHW8WE1jHsfA6KMnC/vFQZLSUGitu42pKTZCJjmejEBQVJPeSdMa4npDDY8YUnjOWvT48H4
22H17Kf+obM06/CsZFJBblVLj+uTrfyFj11AADkU2HZ8ShV8QG5s4nPHVbUBH8fqRXf0mU+XS+il
L+n73JqPsQfuEJ31vdSOqZaVF3XkAuTdoq9SAG+rpFka6dDrq5kcV74nXPqoLfSxi4grSHXd04/m
AWzmQ312R7JWowGe7iW1btsZPAgwR040IRdcrDP+A8bk9s45zQ/L1Xwr4EVADAswWcfe4vUSHD+h
Tq2BLtAvCkm3IiiLXRu1RlSml9Wd/Gsf9WaN8HmimVS7nrYsU4XGLRaSLUn6wFLWx3qxCTXrDuyN
9xYUE6aHRvLK0U0FCNpedMU9+u9gRa7DYTebEVyaZPwksXP+6O53k9nHs41t+zUhwBpExCcvI4l8
J8MH8Hlv1t/PAgI1Rq1pljPIQb25iGBh0c2GPeaXwhsHFMKYLaYJSjHfRHPaTChG5gRu8KOAPEzB
XGw+33yrAiQ+IVtie/51nOl0FFrBCzRV/sHjQ6ZbJkRGoL8u2RRdaTYV3kvvYrPxxskAkVRkjcTb
bwe7fNm2oOPMW26dU1XyaRWH7KsykYQ6+AK82qBr7ibcVZrycQPY8qS0AW3PZWAXN/+D4usiq3N8
/F77au9oVl7fo0rS95vJOz6dS7AJKGzFKKf9p19K08EqbSO6BZ4Ic/6KjAuc12nfbb46yDsrRUt8
8S95whRhFkxaddfI+iDya043sGNVpL0zAbhPda0w0ZYEliqt4b+3OWiBMLOlrmxjDuRLYOy14xIW
GwTiVlVqGmAp2Gx3pHqISmpabD1+uSXQUZunXIzH0ESlnWt6P+7VH+RtGFggF8reAz5W+NClOtHR
sfEsEDKDJRlCaX0MW78Vc+SMm94y7jgWg+Ziol7aIqFQZAY7mpQWQGBPXxoTNAnhNm+yYxp1uDHc
rorHaK3HFQpShKd7cJnmrY4o9eIjELGTeQ3wyZ/nPSrrk9IzzP//UJnLaOFDCxoMxNWizT5D0oCt
XI9Qj4Xy4Abt2hn9p2ItY9gfpjwnzQjEDUGtsUIcmkzCGZ+8zXJQoZo3breHz+7/BRUvMWmgLUeL
+MOD5241Hbx4XEzbjzGAdXdTBva7b1raSng/Q7UQDblL3riAm4x45G5XOCyudv1CU6wCnqJWce1u
vvlO/AX/h8Tjc9KuR9kJHaOYd76wlbv2OaEaJTpeobQ1HOo80WQohAU97/VRdMCfXwJRRpOuO5CH
fv61jA2Mns6oF1og+/GKhWO6r79I2PUyEAsNw2JEUPBvEutza5H69BlE62VX6H+omzSPpSJ4f5vO
LaHB3U/PXsOi/efUHsXV6TPRSLLQwQsZu3QA5TM5/Dr5wSjSsr0l2Ah+ZAZpLirLboWDq+53JNmn
UgrKkwR3Dos+DeVWtUnSpkfSi6gZz0MNfpaknL//4ZKYYDizkXRZi8Oy7TCrc8OWekJnlTXZLn4e
RZ6SX9DQfgV2prpolpyck29hc2EaZAISGIzuREaS9Q7D00qOymOVsBSRX22aq3VvvvgvMeXc/3ST
UyBt1PxOItp+Y2d/cMvVfUX4MGDpFw0IIKtCmRVIFHi3sOHMf2M1Wm2AnPf3d/yeHuIsczjsNP+p
id9ag1NgB3fxUpcntxLOG8Lm3r+gMMIML6xXZ5sNo+BDKEPddSCVTfojPPnMtgslYg3bUDkAjt8M
nGxcZ2IXqoPTwuue8oi4yjwFYya4c/lLcdb0w57fNPWwExjK8Ern+4h6jm9/LyH8GAHGp2PvOoN5
w0RoKUaLsKoRGzEscSD+WyU/G6UHqhq4o10yB4mNaaMf+k/0G+Pt/pTRBANEPn5xN8+zHeSVsR97
PbSRU4FgesxcOvEfigrpVpuPnHXmk7e6A/lBInLVCMtIu1VMtlb7+ac6HblGzS7WxKMFIq8Xx7ZW
IDOmECxL38nEq2Ut0EMqlk5vQT21N5oJ9wbVfNz9bjmkj7DREG+hFmdI84g5ecUBbaVedgiTxc1k
gqjHc7ucosnVfbIe44E/4RlG0ZKVPg2XzNeBOfJ5J3ofu+H4wM1waFJFnIUJjSL+ALZnN57bBazT
lXw0PS9BAlzB8wX3XYdqfBnjB8rGd1D5f+dHww3H9/NWyO1mWev1SWi+MFnoExMgzviNJ6Ycqw+e
6B5kzgIgnC/wywsTUgUr0w5skJ7sK4YwbZ1oBZZbXhZaB7NwNj1liQklGAYJZCdW0PwMdeK2i8gL
V58zILlHTybJEdUHDmRkY6UCLqCdptXCGJHSmaMYk8ZdAMKlyEMmBzFNOf654d/s5uUSJB8FD0lO
ErXvnNx7eOfro7I6o94Nc01NPGcfkUrt+KmVHZmwHxN8KzOoc19AY8DTdqAynEpTztyaYv992L+8
GvJp5hwiN6Qql02uG1At6u0p8c7d88BKLDttIjyDAM+cNy3s2eeAnMTYCPFT6F63+HvBz+ibjI94
YTZmhUMule4nQFOMv1GImotK+JYO92olYogYBFhIMPeSB3uORTmM7eXnfvrh51awgqb9arlXrr9h
OHbgIFC5PsryjRifZfwW53/b3kgdAHY+qh3+Mseupy+dP/j548NisKj9F5ZYOsGCOhvBUAydVTV1
hSAwVHS2z7sNo86ZkY4DclajaBd4aarqaXm+lAlDmTWALRo6LKkbKWRiIdl/BW/qEzxNxsvfqEO2
rqUJJpGPK0MGvqXs+Kjw4tHv1a2rGw3CsqHIEjFUWa1Qm6CAUC7nWO//ldaJ5anePeqO+plI7vgv
vn3eXgSmomITKapWzkNGXucFCv3ffRZ+GjfPW4OMMwu+xJAY9Y49HkaC9HjM9OX48niy64731l0Y
rEgaW+xS4cFzaHpbyaVOMqKUq7xIIQn6/p7s8fJJ7LuE+6NuqyLL7AgTO4tsDQEC16nQfLtBPx6s
GI6ExmMft90sS2ai8d093a8gzZNb0CPSN96Vo6qAAgCMpuxJP3dv0odlqlWPSM/NpIwkk9hdF6Jy
Eiz+WG4G2LDZ2xG1RTAtQZDcwAxXl5cUQTwv35ztkZoGZpoFdac72qRBQ1DAhdpl7pkl35Iioj5S
IA/ekT2bGaeIy252GJ7IV2ElJ8T0+M3YQSGVEuAOgd/kkHewkf1YuPXblPToja4MBa9fEnRQdNAi
iPabnf4T1d4UAhkzkU5r4/1n/Dccslzn2uoBhMZI+0y6gUeOfMXBY3GGaU4oUX6KygCiB4NhzaYx
SGPLgvR5QuU9sJz8Shsu4cTLU0iM1A3dEkMAsebGBfVSF3yppsBFFVVLcp3aN4zSCOfr6lP/Wx6d
ZSIuJHhm+pDe6c2SYRKxpmFSJIjghVjRQiI05ETlEXLHFwYz0urJ7xMgVVisIZyofqgO8VjhHiUw
ZeZ+20gZlaUtvT03AcXkRJN7nXU+rePpll2tWpEB3uilvrrDWHZEP5Y3+lNe9KKdp5SkG4b1hvnd
DNoGqMcgv2RuJT/y5h94P5ku5TNv6KWToLtxhtGBP0gbQ9CJs3BZcIb8uIoeS5AGkxzim0JGldQs
Zp9sJJpU6PtWmT/yzE1XUeUOKyvfQVaHssw+DAlrnpQGzsv80PF9Y58rzgts9str27/mzdbN0T+R
vrMUQEplFlWHvwY47fAkIVKkqjYRDs/wRtDzjmdqq7cpD1jlk91yTyVzLlMisYD1thRMRTFJoWoP
8Pd4xMPscafZB+i8QBMJWFtr8qh8GJuUc7g9pSE/GPwCroVnboXxJvb9YX4rH/28N+4R3OBc4OiD
FPr7LIBeXdPW7FM/QsaQ4GWHoC3pEuD24s63tHSuIWcPbTe6IPAegt7R4TnvDfIuta9InQ+ONfEW
GRirbQ7Lgaj7R3xacEKfLbAvu2KhflYVzn1JjHOm/+Js3AgfGU37T0dfOViONBOLMsIlN2QL4+IP
zoYhWg2iFTTjLkGMqaj04/z3Jj0v0E9Vg3s7CDlDw5aIjnE84kpakg5bY+VI4JKEX6HJifiLG0MV
T3oi4wQPrIwFMBMNRCCpnXXxo9B0Zk+hd56kpSu74YclihbGRLjFjf3MPHnmU5FlIzD88RVgeUHP
qD+pN8vHbSMrvQLc98zrWF5ahMfs5rmJ0Z43OBEZSRHdXxlQ0N3LiRvJQjgTBJLtQqbDLsvhMwlK
SfUYdj2bmAk0gQu0Jm2GvW8wLFT7nMAmWse9Zz1cL2au9leGUPNyM2bfUNNzN/vq7omF1iNOKyWa
XMjIb6jhwLRmdY4NbjQ5o5MWcasrDjFWSeGpe3mdJyHJit+Dc1dVCwk1bd5lx6zYCjtbo9qJRB0f
OSwuH6M27iAnASWuk2lKa74rOQO69gx3LCq30QY5KsOR2OBlmCE1R8yWqhTYONLGsIuLswrDGvdY
GJZOAemEzmojvMBYTz3ghhc2Y+jC0prAXGkC7iwc4jdYDTAvaFTSuK6JtpE8tPWZLR4Y13aIpi7N
k2hvujRx6eHGt0lu00C49N61b9FnrKJJlObq1+tq1zO7H2LBV4H5mnjIFWEyZaVt0fk9ar7T477K
l3UhUFvZB3N9FbgKV3nlDMcL/Oa4dMQrDroKofkKce8uUR5E0KbYA8J6qR+p0Cqhwwzd5rdQNW80
YF3VszLDycBtGfFWNCpTnALmpKIRrGvZ2gqYvhSvjhbuAVz9QWXRvNcaMuEjVrqBVsWMh2sQQQYJ
Dgw/4BtMSmT31VrwjCYE5TkVfIGtGkqmanmVbKzrZzrd7MXdHbQOIgLpJGwf6eMw108RsaW2U5e4
9ZtTsBP/6X07+zHLwNNQsRdBAw+sBj1Gnf3qOD9JGGsgQhZO0eFLCc3fmW31KTLbbYMNRG6Ex+9X
oVZg22uJRzjedWqVykhwg897IlHWb45s41AP9aRaY+lt0UZObZelwFrPSH/76drnsl8cuk1SvScr
hvPbop0oviy3Q4shiVp32y3Erv/AVlFvTg7P5cBgaOcMvADO3Q0Wasl/HlOyF4JZrG1CVoNdUhFN
FCPBgDx4ahxTyIUhJ9eKHRUJa5DqLulcm8sHlJyPNUMWWQgoVpnTbL+xgigwz6kY4VAAlmQZAekP
6r4HwZ5nLxyy9rXXqbc3fZUQyakWQkMWLiBR6CGKQ0vo15u1nYZs08MDB5jiY4lfx5kl8dA4b3kD
X5Xp3Fr4K+tVF98FmML5SudPHM3Dc3SrBrLUEQF/0pm22i6amR9ngRPyQ7gl2F9GIl8GdmX0jp93
jSFym9XL4AgnaN7d6M7jQeC5iuy+jZwDy7CRXGGIqTZ3he60jR43ChFRV9eViIWDtODoUNq1TPVt
VlJBSTrDm9mvuoeDLoOggBQAeHh9sfcoxiE2qryhUxhF5XzGX0kbdrbCb3fk00TQgPBSGemYFe/k
HKrSZpV40d8tCCixQj9lRm3/AqXyzcljkhUgdt8Dsjtrn8nIrTbETfSTWPvCEPYdNrqkFhvi6X+E
7ykm2CMLaXizuYciMzpNT5FZLEbzoD/6Vev4or7hrS9IgO3SUT4WaOAXVKuAEjDBAYp89Qfm2JGJ
68Kcl740SslBqiOuMG+m8AFenZiYvsxrH1dQFdkK9ZRaghtTOG8G5JbNvQMez09Bj24GM9DMUCLl
WdP3YuuL6hnwwyHpgzJL7PkAew6C7u3jcjmuyQ+YgXYIVjBE6drjvvDwl2zjLku6Ws2Lsb+ACrDP
zYedq/f640UylbvCc7noX22EySut9VOWnTzhiUDhpCmrfLiuhZ8tKnxBCJaDlBiuv0Sp3wJ1FZeZ
nUkKK82nmj2eBwsu6r8Mj1uzIjSQvfetdhBuWQrzb2PBjr6ioiLzgLbXog9Kv+turuUubrEX5qeC
NY9GY67pnYIdJM2FaE4jvV3WGUPzmXYTPphUCcTkEEkqR4JEx+5nL/2/j+si3zmJfx1nnmjeU9Aw
czJrBKIfBAc2BwHykLUTNMEDGvKrvl/ZXpX0p7K73YCzmCkNqOn0H9oAlz4H6PCB7boYw0jLZhw1
sqRoC3DCFyiu5gxz22BTy/uxh+sqAfB7E/EYK1WCmFOM/iB0kAKRn+RcVsknDKHh0RdpucyupM0D
uttgrZpvUEa2i+T6FfmMfYJP3esg05WBGLnjELfIxYO2xKJbNuvfFdTCiUW9EMNrO2tALhvdu97d
h5Q6X48RplaybaNzE32ZJus2nOhVvYsMtMqVAl7ubTBVdqot2IOrA+TAFdn94E8XudBIuMDYqZql
s9+8afIeO08YhCsfcRV4DDLtkXoJWL1Vn6cI0lnFSvmyGMwXBIlabSZH9XX4qwhrJ2vgAXzl67fN
AsHZr3cxU4ob4FscEfFSdiCxiTkJ1/f4iRH0bupZl2q406Ih15Mb7csYkI+zoJf1tNs7ywDxGdte
7WArfUSJ9jsfALA3qrHHO2NAb6WMeykXd7M0frLZzk/6yPqUw5JkJnVXUcnOPB79vq1RvjteCczd
QN6Qgpi7exLQsU3PvdQQk4NsMBzxbKmYzANOG6b84W6UBUGosI9r+5B8HC8nrkLFRProG/hcLjyB
KjrLq9FnrGSDI1rL+pGUUVouYTdGqaTnuBR3lMl3+xjvU9ZWOMcTCFs8pFvuHQ9oCgKqKoCyYdo0
xYTT/3HEYX634mGBhVF90MJLsyuAVjLGzRQFXZyRXpaYo9cFlbkxu36AfBLcWnjadwaP3VB/rAXH
SauwsyOKtra83eplFuN0ntDZFYlIXxZW8OfeEsQxz5fFFIEVehK4T03zPrYdZpU+tZDDcTelIhF2
Kelojwj9n451qcefOEuLl5MmifzkYgmvnZkbq/stlPF33sx8pgLgmbzJGMyxjA8iZuId1+0wgGGI
uOHV+ucOoNGuP0PVSADoR02TlIltrOLmWM8jcZQrjftaGcmvR+7rEa8TPHReJM5mfCkfQ9qNfc4S
O2m5xgf53P6C4WMJR/sv7KhflbedK9fUCSU3oGvJ7xvsHp/a06r0EVi4MR3yR+Hfkm66OBoso4nO
C5Zgz59AfHurdr/NTTd5I941cvelQA2vmhvWaNaAmPFWuJhls3yEpS+hGLhgLYMvRRNoFb5NSCWg
xOS8dekTbcwdNE4MO3ZCJx2JpKct6jMEvoXTDkmt892a1lUDleMNRUklq6ECylVlNX56AsIJI0nJ
4/iMFU9iP9PCw68hLsPex1GUUjAKmw3e+y+CBl/3mwU3Z2aOpi1lc3Stt4CkjCI7Zp1nGGGmctbJ
2owl9oUaAkGSMGQ+roP9sqL98MDBFNDYQeb1ZO2YUsf2Wy95JdH9tL6SNxa3zoGFz0jN9z1RyqhT
XVSBucD+vJgA3KOeJy80Sq4m6+1SxaqDMnwRPrb6BXZU5uPKV1QlqWMQwDHkX91kCKfCmsBf5/z6
BsdWljEzKKL2s1UCOGga0t+wXu4u7eQtj7VU1bbR69gfSl77xo6qPhrEJlzDAq0GRXSO2BcEKAYL
QAbgJjQS3lLovuDx+rjqR/MUZ4bNPHAe/DwsOJkgAtHLlnYYDiRy9sNrJTRN5FE4uPoddIzQkSPP
LoBtpiRiMAYQ/P6CMi7TJVTlED+iC+NQngaZcBsX0zaIDoRqQqORufBVdKX2caf6iAgm6Gv6/BvU
KpOPDYfJ2EKF4wIBtu0t1y6U3nLIscLaOOOLqXr5zg2E9tSjLCiH5YgSIZWrAfsyjpCriKTscXMk
1Z0zO47yQiw8JXfv+znKwM2xmSNMv6UR50u+wUpVQNxTfMah2m3oXfNjZ8JtOXl5+lhZFKysk2Qs
1q/7xvI7ORju8GhRucIYvXhIShHi9/tzBmAAPxwwP0sR2jrMyvQ8A6UpeO8V2uuIWWOQ1dgzvsTM
v60TYmy43cIOfp54elEjLP89UQaeT9XmzDhniTjVIi3mmoLLBlV9vopyKZ7qQij27uWX0UbuIS42
vkfActLiuHyWrsorKwkfDPBq9bTRl1iKJYxUV49L6+jwDUy6W7v8/C//OhOCysnyAiAgaHlMZSXM
D5wKbpY0cd8lGdVzFIHjBjhlwcHw6hh6drGnPtOlJzK5HfAUZeK23hfp9sb2T88T9N+L2VLxlomF
Nq+Hlj6jmknIn4DVv55Rhyi/DT6McpixvAjZJrJ0sJ8R8KO1KYAwBOKTnoIUr/NjPqTvrVWUVmUC
lVaaXmoYuebtxFSlLmredlnGcqluPd0f0GHLd++Rx484KSNam48ccPj9+bqFameyQxC4MlvXKt18
15nlzqxDrJH7ryzzR+0nDlFBLKjlj3+MhpZ4vNFzzRu98hFmi+DVgtKc2AUAJzdvUWoPWxnewenF
30KWEs3mFxpDwy9lyO892KSHz7XreLap79jK8Q/scKfhIbKkF+mhPB2SDK14m4v4Nq2txiOF/27B
Dh1+jm1hKI7vG3xPp0jmdfhM6oFRygz3fRE+WbLph14Iiqy6KOURC1aA/rcLMdLm+9q0V3VzEUpp
Qp2EL05N5paHJ32DmDPdOJFv0juAQ177LjvoESGJUlSQKh/3ozgzURu6LJBZofTKr/6n4PtgPWbs
WhIaGRUlgA8/8K5qG6WtAgoWsCt2iEQdqyPHirMFPU87K8vRzLBr6TAAiFkSQHFfz7E3HBIiBtnR
kHYCNFTJGwiAVWmf9EsXAoa9rt0yr4OuKn3fM9YuXHWipiB0N6kk7IqTALhkq26KhRdTADPYJBAD
GPJZY9AduUY3EqQ8bSG5tn6eYR7tldwIdY810gUfSInf2wCkauQt0M+tp5q27LEdVJIotXkvJcWP
VA0l9RSlYHxiqZ/mnOr5rYAAlsX2xPXE+DTVIEYTmv+CSar+KEZbZoFwimxOIzmwekadlo11+VfM
IgomNw3lILw4ZEFrR8uP1rTFEcMCOTYHdjFffeVxEjmvYyUQZ+DUqFGEGJS0kk/MnnMlueby6102
Qytu+45v0L5ne0u8UctbmHtQTAsTqbzjqRYyh9WqtMMj8uPaVofeC5a5x2/qJsgavl2i2bn9d1uo
GK9yf/vnJM6C8tIsq8FpHTQpen6Ro68efnTWjeWoGS4fj/EAbRQM6e+y+VXCWCqSprcpDXI7J3h3
LUZrnLj/tWR4QLQyS26p8pyMndzEbTrJqtky0laZAohEwEUWNBhh895odR90EdGnObBYy/+ym+PH
komXbNtC4nw1xjvzuBDIXN4fDSzh53Iaxp7JgUnGZDQmcXdA5QfXUp0/lLlhWIkOZ0oa2EP5GQpX
BoTEAYwp6i3YId8vhP8fUExRrSfEDsYRQ53w0YUzBhgJ1FALjfpS8iulqCm7wQqJO+Dx+AKBjoqx
1grYqF8/zG0XGqJPIFdyAWswK1rRMKE8Rf2GRfy+2q7P+BQUN1BKgr49FeOlnKd5KEQm3a6SDx2j
FiS0q6VTWPgmhRNTPVTpUO8KEMgM4gcQU5DSKEZVaywpNzDaiZMFQpNXFyLMc5wkbzD8KE3NEPbI
HwKNbGS2bOpWJ1GCg7f462yEWBoQ8TC5Bn2Zw9QzKLE4SiCVxYD+9mnHGOmqg+goVH23zZXfzxlf
nnhUK/3WCah/foPflaTQ+7lUYPUmB6P13hP5h5Rqe+jShZyF3kbPBGnLhm++BR8zLwxAJr+7HIu+
NgRSxgFIg+dx3UqPHUGaMqZmia65YQJrhAeJB32mV7S66JkHOpB0XgZx4lpAwhDA8GBwYDb/XGbn
chC9nbh3x+8+90IePpX3HGCm4C2CKCf7XWYFZZSHW6QVKfnr8/QOQJxEKkW8PhuxrWoOHUEG5Etj
tOnlz3RBHMuMZ5dtTTF04TXIZNS9qifIcJR4UE6wGu9bVnMl92JM9+DKONt6SJ4GlMm1SY6XUzXt
iKrV4bV70vNzBhNOW1wjDxxYQgG468dYjP3BS6PFPJ03mKnRPM9eqkLByCE7K9fWXqFN8abLj3I6
4/pHCLS4rzWMrl2zuBMuZADbpRTlP/PKkeJX6fLYGsgh1ZHbAHGSIvDuMQpODu1DhIegfKAmnM3o
qHwL+4Qp0ShW53cIcM0Kh7XqFi+13nBkibaosR1F7eeTRy3WWs9+4/j34ATCa6GQKp2qUeJvjYYG
6/1h9LswxT4+IBcY9WZh7k36ex4UbWZ2hLCts0vPkysUX/E1bTGHueFT5FLzhY2iJKUw6M2HdR5T
U2PxxgOfIXg8IDF+IHuVOQtNSDr61nT6YfEWva75AybzKsyX3Pf3sb7NgtJVAR/Tr3Iq+9D7IFJ4
01yaO02ed3ldHvUpV1GSJiyWOssno+KhHzwUcO7gaFvaa8X0JUUm7eFqvG9V//ZRSGw7j4S7EEwf
HsCDIrXF8/qK0ngOm5j7ippkMiUzPEMu0EPyKLxANRcYWb/TZHklt+k0tUImNpNYuGINL3AREH2x
+lvO/CYPP45AeItd+/4skCaED0b8ccPc0jy8zShL2l79tr1ChyPbtrZpVagRf6O3EB4XFmAixLGm
jTQ3Wi0jZHw5/rFeeynursvglQEyvPLt5WDIBOi1l2uT8zTISRlNNJcL/gid7XSR5I12WTHuNUFm
4ho26zs34mr2JC5dFQZel9fiRboFxiErcstJQwpcTYp91UGAFB6GKmTCFBQnyT4PUtZI74rYWTRf
YIv2kxfRl5Oa543A+zolTC73v3/3K62Xyf+Y67KHILK+6iQZBc0Mh86zBqp/x7LTXmJKihYZnMWY
L1ED972boKbR8UMrggXq8mrFKDTGsw6/v6vM2yELXzUQ7j457btUhiHdhAFQLPlqIyXbpaNAmMhY
BNk6oASvIVmZ3p0QYxwtKMCywP0/ZOtUIVvyLUJHPgOm5bjXE2C6U2A+oiAYtB+Jbf7KNgAsnsJv
Oczhuh7RXKAHq7s75KaLBJBWVBix6LiTqfci6adCAhlDxpXz7AgszXmyplSnVR/U+Wj7i5rCuJ3d
3Sim7EA2IsHLGsrUARbGhmNXiPKNq0HMaXO8kyC3IZMwjveC42RfZoTw6PNMz8BVmV0WL4s1SIYp
uG6iw1MGt4Ss9UB6atmADZNdzIJJhEeTK4tbH26MAQg3blylj7NQxb58rk7xradaoDrA8vd1J2TF
6Weqca5MyH5RmCvu6POL8ev5YbL9fA2nPKdubqYw4fxZ/+KwbMQ1+JrYfgC+urh/RPNy6iY49FFH
g/kTLtanQszvnLBlhad3EVh+aKr/WXivOIETdw+LqILtugX/gbe3SX3FG2/keOtFngJXYneiJ2zM
ukTEqzXO6nDXskVKEYHef1m9s00gWAmsBpTAACSOgmS9NgMsl8PyGLJIoxxBSG5YT1uWKL3VVTvm
aMEVJwcrrt48zMzuLTntCoMJTcKfsJi75NdFoWswDZX1auVtxEMVh+/IXIwL+IfB3OIOA13dVkCs
NELOUiF4QozEUOndqOlAx/9TYAb+54/LYaxAHp6iU7KJwiMhUrIF49lOjzf9rCuA7mgkXq0GtVgn
p864jd0nieS/+vdYixDCCDQhr6r2nAsW4Slr64k02miLt7EV8kLEc2Y2ohG5RyInGyFZoPVEgib0
e/pp90t8blw8RHhTK5je7umWmRbtfEGrWAYH9QwEm7IUsySRi6ZEAOaZ+k0d2b1/6M1PGlJAA4v5
kKh1Mo/yUv8fxpofnm1Z8tpikhHBUC3uytx2BqS11BGcj//6gETO8BYBaMMw4acIG6m7Xm1wajKR
TuoQWe5U92GPIyClRJj1Yw1n6S+C7pjN5qE7VxIjwXADEqbpJuhkxisT1esLktEQavLK3uTENcpx
3S8/iUWTlRrPzUdp8cOtcFm1bBj0idwoXVBBbuk6AVi/QsKwSuSUJbQP3jpdpak5bQxRzCOgRYDF
hSPkuteGszoCnQLqCAgWBfzyM+7nuPCTDXrd1xLy90GNwje+kIWMAEAVZhIgJDeDJ1tjVav82XUz
24QidaLnYOfW+/3Rq9bawgHi9APYMp5A5Reeqhhr4OF1w58nIMS7APrwG67mwji7BKSBaEVPqI0r
o8929A2NIfEARjDkUBoAJiIocEe5YaoSv+Uk1//a+Pvtk7hLmOjPrMFYyuzaP+e3GfnpFBH/svUC
MjTEk2/ozaUkpKaLi7tTpjg42gvDx+qR5xxkDej69Jq834Clsywdxgc83S6ADjIcyUeLEfcTxT1l
Ss+lV27ou3WGn4aE8lhSsapXnmc6iND8dSm04bqpqCfoTd8LlrrswWHTDXU3P1WI4Tr3pUSZtbzx
SXC20FBeZUJnxszX3ZgsdvldEFAQla3A/Ow04thpFR+HG51A5PoUt2UXXfVj30XHy/+z7mbmv43l
NUz/gE80C0IMZZMIjhXFdcwMX3I6vnrDZ4nfGWGG7FHIiHEHl+cR3JDQYjkGaZeKqpJQIwUHtMGX
hpDLXaQaJWnTF0PNo1k8E+9ek+uF/Cy8xJi68aDQkzCqdMsdo+GB7udvzvOdGPsYeChJ8WJzPjKb
USbVeIzwbM5C0LzsI/OrSzSbRrcBgbwHIEVb1XVcPu1WbLV7o63dmMBSynK/xM6YpeL58U3JLO/G
llsWV5ISxy6HWsVGFU9U9RZP8eHZjw9C0SRlGAXGcvo4b54sSoibGrLgiVRgGlOAHuF+ZLGUzfCm
3udMxGPQ981/rydFySTsWgztQvjBZvrXZgWvmjWfTZyHOlJ0kjAOvLcw6N03OENLoKJopgJCpNT8
lctHact7VUkLr6XqhizNjYltKwuQHVEsS9AsFjPt+jchCuH7V4RZwqRcXXMkQsmzG6lHBWR/vvKK
u2KQEv+RAEelG9xPiVQYcIfjWq8BCOtHK86+J2pvF81vvcYDqR63ozHkuZ1YVHUGvsKlKTEvQz4u
dZavWn7IZ54Q44Jv5jwXVmwAHg9K3qfePbuF2OTBDlJVWwwmRddzbccQnFN2E9+l/1vJwwVZYAD1
xlNPYEZ4chUCsQos6+bQ8dY26jVRVgE4RoIndo5HnzhaVZJYWB1VCu1gKMqMCrni29f7th0hpjUm
xaG/2Qm2DDFo6MrD7hMIezbJ5czaLPwpe6Kuvn7lL1fjlc4Wu1+pawcu54B7yIvb1/jIpe2B7+PM
EZBlmhUkOgvoJvz4KOZJAaAwwP7FVV58ntiUCNdI+fNLnXhdI+EPwyTpNqzVJuNQJzzHrRIZRkVz
8ldOSEm7w0fum55ToJGBJFWG/8Hld8c29TZSOUnvP7Cb75kd/v3kNsL2FCKxmT6RVMU4o09aiRTf
i2LM7DUTA/Ohrr1s5EAPqEWv+pSeqQuF/9zzVzhJN75VwMJLWpIfyhrjcmUOCZfhUDvmCN77YjFp
PFBKzXQxVy7PnWnYO2eM3QjBi6rIWajxVkiL5Z/4X0S5Az2dKn7XbQ2J782wuwpGjDHIQ4jLLyf5
pTRWLehXHMs1YY950VdieULXnmvonpL30IQAVhrVpqOO/sPuOofmFUr40Idja5MkNg/D6+Ml+OrU
/Qbf1quYFmjQBLur2iRe6CjWbmD5pJjrIJDEPDJVW7VCnXd3Y3C3Cni0IS4J08Yyxk8WP2o0sYBQ
IhzYN/Yo6qb95iO2jbl+uuYqpg6Sdy7+QHcaRw2X8qU8s4KIBkLyBZASRlY0KTNdPJkQKhNo4fxY
vvUAnUDOOUgKjezVkPXwpSY1sIEQvTzTo6JanEMmsIcecxXzyzKbqvPPqcLoVfzBh5bk43CtbtKZ
Cmg1beExkNW5H2Cs21Bw+D9Deg4YwNnBkPHJxUY1YeIjLsWNYgfuoae4N4+mPt7SU6b2oWuKNLvv
e//cs+SiAURLK4r6weEBBBqzi4qS6x+ToX3Oxsj3+geIKvG3QfwmuwGcTMhY3sTGZtTId+kXYR3J
rGHUuKhsc2ElMhzdX0nr8tD/vL5vjWxXBYKvcPmuIh7hnKq7jxrAxZc7JZzTw/AAMxMD6k4Ghu0Y
/dH1eoJl9CFLeL/qxyxHtGt7iJ+H7DYRga1M2aTzPieR97qm0grR1aFpTBPAh0bhYyJeGQNXB0cG
uVGTXZlnssFfYN/eXnfSTonAqLQF/WDEUi41fc77yrEzhddBjnkMRsQRVi2hAm23sOra0Fx2Vmcd
yI/9CIGp+hfIMoXOv+HopcUpzf9XJppxAVvFfbY3Vdt+GyE22/soRjltSzUszh2uQfqMf9OYoTCo
unXz+UfgVz3RPTQcI1gdjtN237DA+aTFZQ9yIsLcyXQrjA7VP6KPkdsnKETG8ADXw/GMcn50LKd/
EzvTYs4Joq3PjBQv6mKOHAO6llN+Ok1DeB4CE6XPN2pllVfzMg4wPmUVR/AajW4DJNzcHB+qt9rC
ACGU9TTYH60wGXgLFqdLMr/JWziD961JtHZiZGvRAunc578HwxMHVoFMDRmcIYJ7OGuAMmIksr/c
cZC4YAXpIlEBfs7Id8HBui2jAkgIXSFwWkjDeUUVojF0Acn3SOCUjolbLDbPTJOF1QNxjammeSSa
PSsoZ9AfkGAmHBmxXJP0OiawEHKDJk/hA3P4zL30P1ae90o8oE3sj68zj99zyfJXegE7FBoJWheu
mPRRX7cDF75XD/dofD9bea1qz4d63AI4DBcgoEIVo1GCpFXXOaLunpO2mbQm+iRuLJBarNfIzMjp
m3sFthozCM/F8rToCPNq/+MnMYFGOB/di0TN7STn59vyzRHAkUPNQumvcsj+ataWu2ayfmqS/PuF
IV4P0+oqYeecgopuj5njsmYKTgXh0q19t/L3KdN19FpuqMGIQn5KyaQFALDHRRLNfesRSoF4NlTg
7TIHAq47RZZcvLbz0gw6nYQCXZAdskiKkF3PRuu00Z6OC9j82d6UYILKivIkfQplaTQR1Zj5kWl4
Y2L3hJRJJsN61Rrpi+QfT91r4UPCG7n8GKXfkqIt9bYMq/jNC5mtxV1IyqHNLIfs7pqs+QwcrJLR
5v+PXzKpwG97+2PVnNytOQWXPis3xXnycJYKWLSTPABlEaf4Yk+MtR4g/EkLWfVrcnDfqrKQctaW
HMj0KTj92blQLtuIwtUn981Ef65j3tPevGuGE0zFDOfPQ91qItz6jQ8IjG8DTfoZ+po49sq7CPIW
C7arYn90xNiI9AOgZ/kq/hnkSn8DhZNuL27EBVBbfUh/LpGTOBXr1muJmydg+nXC7P31DH5VIaZJ
a9NvrziW6YuI+Cts/JxqZYSqb53zjdir67JodJJxHiTn4nUl8YcmnOg1sXt/9HzYYimXyhJ5UmPL
XT04aA+pKi04c75sA+F2B1ROA8nrgLzUX3by/22ZU1vAyNH+dWq6R6/On/aKPtjLfUuW64K99igf
rC9GsuFpcVsGZK9HZODnBouUxxylcdRSbmLZQZu9Wc0o1Sfa0BBp8cRsOkMqu73zX5tFJq5P8w5Q
hPIk05WS76YZ8OEMveUr5vj3Wh5EuGY62tPxdKcmqlP9u3HYL9J65r8bICeqdW2a6BiijAsG86/f
K7oIwx5EhASgzGc/2PQGkeQWpit3SvTCohy5NFKGXaUWgrsAkmIWTXapw1OLqhZuSE9YIaiooBRj
QOOUenC6dJKK1Vt4suWJSoR1imh+Q6mrU5pv4mQCrH9xcyNOzJo6wpZCMVLHyj55QHvMpbiJ0wN4
RiTeZlt2ZwGPCuiMHEZEuw7iPrRpKwl4gJu9rxo+1peY3L6XYyhSD/Pd9hvUKZw6NlcI2s8j+WPB
VZMuGuiLFsGYmIOzWEBYIoXxAPZo9NvzvXhUXFyd2pZzvUeHm3MzWgamtzxTPJCuI2jhP01p9P59
WFlU54WhU3mZOdbWBqLmbb9/RrrD/r1jUciZsO+nbijlcqreH+m2AK3XB4mUXcy/HbnCMq8DKQdV
cSrwhCWsuouZFevG4AYWT9libiIG022ksnL2qUPK0ut0SJ1R4KLRwk5o1OTNx0JCH2zEKm1ximcy
13yT20Lt0pQ7EXKNDnhc0UDnkSw7N/dNMijEMcRvb/KKNNUozgvOcmyFrHulhvAQTIxKtoY4O+Mm
+E/ESzqut87h9dnxxvCMQaB8dpGli5oh9Ah5oTW0sU9UHMgN7z5y6fEk/YMN9wU0mKTHjg5VSPCP
HD71vtkYrXoADyo5QoZMrLmSdOUzihHd1jtfK3LC6YxdVJO7vGb4//VfmGUqC7rfHV8I8zZvu7XW
2qNJhDw8a+J+aozaHMn6MePZOOj5ny/PX+NWJhdETOF+TR+ij/s0TaKFnP+KRxZCDaYTv2JrhLCB
W+aNmIBDtS0U68BI7Arwv7O7Sphyf/CGzmgZHhCpb8oIB2XgPcMRPrdPOItGTNAGh3v7UPrY9Akb
CWTxOuWBNSov3lpBNe1QvP5AZQxqHFjgMCmehcc0YGGWHUZt2eQQlPpwINgMkM+ddSEK77dVIqBj
a/V9An7rZ2NGniPge6I7wHOGpp49IAv5R5KainisZ/xazYyVwKOPyaofAguYk2Yu6DaOkRWCTtvf
/WWFInBdqvk9C2ZhDWUTWz74KJLhlpne3f1LwK9luyxO+28rxOXp0mMWRZp7NeQ04MxzS6xVXz5L
uQXoGO3Q4W8fcMivuMFS6M3kJF5V0idhIixAp/QFg+E5YxPhljGsRzsDDoikiSDgnpkVQvVxgIf2
RynD4449AKC0k/UnwwULbloVDF+M9Q4WivVMm7vINHLqcjbg/4FpRHLLW0w9YfHIqVeQ+kJEPUkh
9hLUzreYnD85YNh5vCy5dSQrn6TZ/xawQ8Se62EFWnrXSgiDY9PuB2HP2qHzavc0Ahn9vQbL4H49
UAcFJaF47bP3tJ9WS094KaYWPVleNIj+pnWzOTBDZ3x/BtqKBmG4nUuhdWXqK7yRb3vY2J5bY3qf
j9KuALyYCLRSVykgP3XvIllPk2SD1ZEvZJBPbJ6lCoc6JFfj1k3wg6Rc1GcouLBt7WOsFFyuQNyI
GXmzu4sSfB8HCAp9K9WVXQseupNqiqka79IBCUqSdiUSkwJka3pYTrI7Kr4v+vNwAAgCVRShHRqq
Jxbo5yYnINzO2itUq4r7hUmTN9xvwraWpV1lDp6+rCY20H364I+OkrqhsiMU/lfJnAMZnjEwB+Dr
6l6RpKrlL7bdqhp7mDQmfdsrtLGDxRmUdJN7hH5jAb1kDK9/dfchfQesfUHU0Klc1h+5m0mX6L65
jkmwLyaTm4T01YLkBKMYKu+S0cZBlPvpJ3Nqvz7KVCrPQtW6PHrYG1xpBU+Uj0Te2VenPDkjskpA
ovrDjGzTK/iw4JcJmBuVjKp/WMTpEPtEoKpS9BL4Esg+i1GwK3rXjNPGpDDm85vVj+0aIo3OODl3
eXZJIAp/izaJvIy11MuPXUzszULgzYGgsoGtYF5ORwTZR587LXuADWmNVvP2ZGGnJKvqhK5bcPpi
+C5JYlunWYZhGiXnSlFtF3x9zmqgJs68sxH/3tNVzyB74J7L+ZnINsoQI8X6ECAjfU/4T3crbzjI
qCZjnN8kTCMIGirsIK+QY3lnoiFqsWMZ7a+4JRdY1VyOVpan0OY/+aA451YY6et0Yyo/kbAvW85s
sqF1g6ZcGE/Ux9I5wOpR3j3Whh/NFDg330pCssfA+TQmTPcrE/wH4YC0AK9hKie6mR9mejq99D0b
8Di8CZXqQwhVYy9HNrUFMcPHi6R7WpW7+sHqZALlsayyhj3PjlLR6A+ykXI2NaPq219M2kas5t+M
C53GOyQigpnW5FPCjkoWE+JcCgOt4m7pUdRmnimGE68JZ2y+g1RRPM+szh7zJZF/L8rGNYT90tsw
jJgJS1bt5YrmoYpvUVkVk66gvBsoJ2wG46lBLrAtisKc0NsLNz9Wrn6f3CFfzkhkNgQLyrvMc50K
17i/bPdLtyXjLnI/s+v5uWzNDSnXYvPDyP2j5A3qjGtTR2bpxk9nDZX+qbpQz3wgStC2FQwyPkbv
Ke8RyfRCw74Fh5bDUjxFWK7fAIz0s5WlODsZorFlhmHpBcrPH6U5fotZPBf0Y07NTOWz53ZLMOjA
vIiYuacjwWwYdgnTX5NCEZO98sYjEM6pUHojkPc4DPWCV6MT7ep3CY8mnbMCcOPMSssOwGCtOgSA
qxZMxhYEXA1qsk21siCgcY248XbQJ77u7ZPxO0YPVskMuEcvCSN0lM2UBEmKLM5Clzvu5UvQL6qJ
FxI3gz7pUvDL3YCmuABBPQk7TJh56WQ99hI5x9ECMe+440TCkGlz8Fr3ShhVhljizDuzvFKopseZ
mHRcg8SKWcPe1Jh54hOkOjzaEQkRWHjYsZjwZ4nTUIUFs+AjEYXV8ScS0kAdSl2cXntwvTTU3ean
6bJ9xKBJIsRaeI5U0MXB4TEplVR6DrPbAL7kCjrG+RKuVWlMcERiPmFrzyRA0D/c3qEfKFL8TpUj
mbSaZMsmpMxmxdk1QI6PKlzvrDamCSC3SDT/toUAlqQWSoPFmtWGAskMaunQsshgvrWQvjdUsIAp
zN2/nsS3hQ+JeUNyutlesfp6LGrU9l2Hrq0NuvcuvLquwGDgiklEeg+lmKT7WDJrLzDsVIj8Ltd7
cUhVWq+Qpe8MtT/kz2i0tuYBpqNTLFqnY7egxFYYKGbTF/2VxxqnjICrl3rltkxq2A15rPAauKgF
zesviab6ATdLaamcOp+un6gGrTE/ysB94/rj75ISeM8gL7iz/k+MPHCwYjP+0NxGUvumMrDrVfkD
7ra5tszekqHYaPKz7EwbDUPXOBRr9e/huVO7Cvdbo/lH8ICAP2DdLx5ZPqh/jaK4uIEJWsKPiHJ4
ueGBzCCRLI/R1+zKJI64KsewvJOcNx7QUofikChKWVD6yKxd4HPmevjM+SCsdPeAYupnwsnGM1Ei
+BoiFKp0hTyvw3RpJGv92KARI1zeupuiDW0aDwfHrFaiPmSKjKoB8PvYzM91VZX9+zRzNye1Ra4G
ptnI7Cf4eXH7eE487wFZ1DvePStHx9sxrg7R4g9jgc57TCpB3yCd5hU0RtWA5Brhakj7DCHl4G94
OEqlmi57lsV8txeMYpPoFb7YOFcxYCujkKB7l4Z/n03/JrRfY3I5mVvKcMGqgJNv0D6OQO9MiXWJ
a76xfpLwTqJJ5vqfrQSkNhGHHRUXcuLrvkx9AqVo9ewU/OL+XEY9eftfHildXemPVSJ+PSY4JRzp
cDP3sBcv8Dkxfw8fgrn2aFIjprII0mdp69E94CxezFSHlgOb+jcfJVykOYZjlnjYBi74Y9l+p+xV
wnRKilseHjfFf31iz1CSalHP22rqptIQN16WDTlUMUgfjwMrFfteRjHwMDxofn2vxVQA5kUZtD+u
BT/f1A1L+H99QIi/+XGH5ZkR+yMfuqlCgqeOtjJOWTRilqVLlYfWUdpxkKRNMPU/TYOZwBfc1xIn
WYasAPgoImR/yU68aRzEibiOdTSmrQdbzyXe64CxW6JAQYqd7SJEJ6F0c3BuBgaWL9zxF92VfKhA
KJiWihh0GOI+j9SkahoA8LCPbFbY/S51XAO+H+/TjVjKTngwa2OcstKP1W7BPHsa9Y2D9ubXDGYc
NNvKpgMS9R44QpDgUN2peq8QsNzhpqVDIoCAHj4j5fZrnIrgfFdBcPkX7lFzr86idd66E2Lsk4HK
F8OybpM+Zs2KkxI296iHJfQtsx5psXRGlAEum/jhh6B1MroQ7esDT4FKRJDpYYqVe/8mHa5of4PE
7t3j4Jj780t4g7Q3Jk4WELKbZ95VGCTM1NvUIlgHeQPh7tQxpL7iqbJXgSVjfGomzel9DWlTPWSZ
X67hZaHc9/Ar1wFTH/j8eCEW3biXF0U1pNPWh4qY7UwVZyo98tmBDVwF1NjNIBEsYdIdeM9eZXne
pZCh3+f7+7fmoIIvI66D1Yem/QlnHiua7W/33QaK7DN5+OVXH6TJQV3LLvQJUvk4mLMYAAkydLBu
f+6//hUEhJjuhcadAwFtp3ulLsbbIhclXqgo92yZ3osipZui/0L8ZGaXB3fw5tzdF5sCCitvOzJg
qfhZHnLsnG0vF0cKym3eUM6fHVGqSVhzDbgyRLXpB4ArhyVf19XeXfxv8SSldeG8Woh8XzvTCl9d
SlWeXGHWHBxh4mhiS5OsvcKn0f17XLRZQJO84aNt6j6Z8J0UX+4GmSObxZnohEYaY6DKXlbkTFfR
y5ZnJ1NJV4pEuU0wmElALdsfKj/Iyg268y1iMioPYXCn2bODe9NFKKI3fhX3EKZ4MpK1/v1qIv3s
6Rup6iSpL1WKToXcjnpvb9LN+6ZmRCY5KYh0YMYAjCGr1vs2gr67XTKPs0ENB2FEB/knS4Z52GP7
QrdOSiujwFHHwsXtguXADR8/1jCp/x1Pp8mkzXj0TUcqnR7YXkBlqkiAHDtns0g6DTX9iHY5tMeM
ko54qcNhBnSiYpvcf3IVxPyfkr3Vcdr1l060lu7Mc5BDbgPccc8xTYhaJ1CeG/W5s6BU9jKH6CRn
0YUls3/kci5IT0IktjCZ4NfsTZHF7xYzJLzp76Td6qt4B/JFI/WFQXS80CjMyZSyWcmLQqdQUuQB
mVcCjDjR+ppgIkVhrgfPtXHmiqvsDJeSNpc7AFntLrupXkj/u51GxHFA4BRUGXDzGTnKtnPcK1RS
ofYkBG5UV4ZoVRTpPRy1sb7ZFrgfDzySiwyZNTrVGM90kA0HfxaXZ6V7Bv/cCzLig9SPoYIIM6mG
x9r0NHRRpP6FMFugR+Gd4HOp5chowYZQSlUE833/nuDTY5CmNKIx7TM498h5ZPKB+FN53HRi4FAI
owi/vvXz/ZZY6X++ZV+WMnQllGzrO171a33X5FfusqWAXUzcJwkmHrSsB2VGSYJ+lk8lnGA0g9eF
n9UdlmpJwQpS6wJEXRMNWwm0XS8nkx3QxgFnscRiRo/AOIsiY4hp8bVK2T6VyCjx/Ozb5zseBtNS
4AWFpa6iBcfV7xcdG35zaEH2pYGb+MBERemzGm93VkpR5JVO7cr3XFguVxtKUXJySIKYGHVtZUaO
Whc/FmPXeFihqkFraKqGjVS6Orkj1H2D2CwTZSr6jOiIq+UfQEImNEyrUEmzEyDVxQd9krp05F8X
G1XKeJZyWTtU6qxgB1avYvImREG1pVpF+qdYqg2KafL0A4GH540GmApkrbugG/aq//VaDWonHPKK
wpKjzaJMelthKxw8SSQJ2F6KCHciIAGQhWeZt8Usbu5Sg24rMXKlUjDUoUzlB0LPjo93XQLe8b43
lh4Qn72PsLjSWAnirHTlr1T06NhOb3ECgjPOvSzu6LwTU8ecIo+YkEFy5CmsvkPGdkTI2cAHKGo8
ZmOEWlODpA575w7XqlYZWhgtCKDh5lI/jXjswca6WGuaIKefE4dAuJpj5ZYG8/VxczlDU3MxjG4M
Y+/3QT6gbDrZm/t9R5Uczx+M7OsHL+gcPEvYPoeY48shKf2EHRpWb/8ZyINh5eOm8iKY28xuI1bo
S0K/ojhnuzB65HB3m9KFz23tEcYOwConnfqzyaw7djeiWpmmBSJEn/+lbdgKTI9AQnV41qnYww0U
Gtep4phMfMZnusXjrOADL/1P5pYKqdrKMYIsH80S27TQwZZ2+m++5ZBAhAm77gqMAC4V10IaE7bf
pfAQN4o0V2MpLRFUKv9sd6B2gdjyHWlfEAKGj/3xLa8pr7n/5zSAbpVy2rQB4veMTkncSGbGV9xA
Xx2l90lF5k83tuOg6721adO+qL1CdPl3JUf/3eofSHxe+p9cAQ/RgRoq4h6d8Vbc2Y650LUA8+yR
+MZNcfql8+Yp8YFbbGrK7kX10CCs3weNnQ6+Jr2ohN5fzp1MEJ0JNqlJEIZlyHj2JhmtVsU1bDDm
+GOdV174bmkh83SgXljMKmRkd04BVDAoyADT1dL7Ksc7JUvvkL/A6z3AySpGZNAwrOmcqEovdNCJ
Qoa6RnwkwuiiOkTXB0n1z9fbII3yEwH4XR6Hoe39aX7h6fxsD0G79+qRMRkz0tVYtmAMBM+Coxh/
zBh5LLwMni0ASLxV6262pgp/di3pOJoEnFXkb+38TIfRr/zD+bZj9Gra7XvcpFX2rz7hBMqsa/wM
p91QCh8yI7kgv+2Pap0JmJI0wSYL0hQMYke9y8qZS45STp9bEhdrQexBgJMAnxXQGboqv0Xp5M1C
vvivNERCggA9hbdURB2/5uYzVpMhbpWlAo8J3o76NiHnJaFu3Cn6ceOS5BrTjE5jlw4mDJWij5qx
8+6GpMWH5IWBuf4G/c6bKgRP95LitB2tIMedTvDhB5M/3xzuVNW5nFVXjH2q/OOYqK83GVRLF4KN
8aL25pLEOgKMze/K3YFv+PGJMKwcpJ//U/UBpFnfQc5Fs485U6TyAdD09EOPBQRGQVYduQ1V4v4Q
douwdKHxcPnWLk8DzBD+W1zP8j6vFg2Hqqzc4LboOTqdGi+EX3BIir5EAsZLuQu6G0a0dWGa6/SH
rcxXDbBG6IGd3/dyBnc0xbNQZ8hxFwuGKRk7UFS4qt6XSxYOR10zgqRrPpjorbYVppPm1rbffUsy
bjkJlu4BDWMR1XJohTHSTrgMfqp3YA0yrqMVH+syBj04WDMRKFYIa4YMyTZYkffD1QxqcXMyjssr
/FEWfb7bwvnSSF6vTnIjN5Y/5B1wpfJ/PoLAYiUrMUM3kIk5Xq0/L58y9+Woa0LZ3g0LnTjL513e
D0XdvKIrrrrwZ7Anx5qK6UqSE91vdMESjvUtued04VZJ2QSQAOYIw43YfpjOztnInlUZStioVTBk
wBY2zstibubJ21LRyT8peG4wM9gGjTTDy8UF8sLMDXRhKCHPo8M7qqe+R8zzyipTh3Tmq/0sZVSd
PnRAplDOn2RMylYDPWZ6iRJGrOv9aSxPvxxxSCSmM1T9ibMfyxXvhRrGVWJzWLpjV8y6BLIrqcXs
8iD5fLK3y4B4rzSuszRTeHCJuRg6uWOAJdXLWLg7X7zuGfYD0+pqK5Ekxfb/RsjNsFXAYocHFsUJ
V3JTVZm65yvz0gdob8g7EYR6tZkgDMBbpvSP8vnQp7MvSnBw663ZZrl+Cfe/fxeLUeFSgveCA42v
SCv9eXHOmr2dX96l4oIa2R6Ek179jfHTeY8YHuI9gb1NyyfLtlsv6AShGwGGZSOxZyqJjG/reAMh
O4buS7XnqmbjijX4o249LbapdoWBYDIwKBv3+nzcXobKV1aBy/y7MtRaQ2DZKRHG+4lUOd8yTrjl
jODzEX+K2I2kW3DD3JqD2CGKS0Oeyxw2u6+kr94/1yvqJhrBj6CMoJWJSfxm843ka/GKYz6dpaRL
mksiXHsVm4FJ4K1uj2N2rIPrK3hVYrBjWOKNaqJ3zMkb2zXgjq9YHFPK3V2lLjWieGfQiwE6Xws+
W2wWSXgx2jhzzgj6a7L5VB1ZCNcmnXlbbOHTuzeDutxPTqK6gZhsCzQbIu2WKKJCxKhFUB6SR7aG
B3O7TZfQMFLIzTSkyIEc4ij0lWNIvSb0IoHePhT1nKE3Ft3Pd7owXLwBSrYWXZBMag9XXAPfs3Bj
IOdmznBq1yY3sMzz8TsGyu5ZLm5Xr6aVvYc5mOWqmzO75eHC5No/5kRmPkb1H1/STpSrAdntbiEW
uN/2j4I35Mknq44HO/iUh6XA33b+Ai897M4NqApBu1QX6y7fR9nGWz0Vhe/+rdRR6/ZFvTw0IZ+B
jK5Fmvbt0tVdFjjlYtva2BXdVvgkzjan8SX3NnaLi1k2D42xCoFaaaPGIKZqp8IQs44tVp3DKIwA
cNAij4usuylPKYsBSMVmqdQuHqfH7SU3VoUYAt+hPZtUuF98qsP1/4wXwnFT/pZCycQJn9YWOc4H
pIeVrg0NC+AQMjt8n4jbPatUX/ywnyJ3qlPIcSKNRm9e7qhw2q2HVc+PJMsiIOxmez1yX3KxHcIo
UxjEkPCNmtv/7LANmgBKPJUiNzBcbViOybHeDHLIHqYsKly0Wn5NRldV4Gq804EW8ktDb8cqyojf
aQ7JIHtw/pkUSbcu3PIfq6XFWgxpd67f7PPo+a0P0+P+rIVTZtBzXbK//xogz9pfXjbN9plng6uJ
sgkcUa0r8xOx1yijww4IvXcsnzQzZ8hJGR/YjfzmdRgYq0jSixegAaBeB0FVrfidoNipMTfpwd2R
MHO2YHTD+M6mV+THGUeaMOfXrHG9eDj4iF4Ryrd+IJcuuUYrcvy5IArDzXbEFr09ux8YB2qdMSFa
0zqfeSas6FoHLlWMwpz1TXT/ERAl7t5HaMiIXNvZ9ebLqw10pNVmjb2GIQhaJZBYYFiD24jjhmX5
iwQF5fYd8JRGBFXWkQkNmmMVsZ20v/ipzikI/OEhZjvD8/sH2POm6HCs+4D352IyqyTjt18P5UoM
Ak/kmSqApVuDSp2HvvznO/vYXdASEwm4PHCRZoXhhlvrLTaV1j3Si9xwtkY9N/HZcvV+hJJPfAIk
QJZDUsENRWfeiV4WPaytc0xjLVe6loXcVqfQiaj3Sy7Q1AuC8yGx0+WNltZX31E+v7Fn5KWZXPHZ
op68aFCsJaAQ7K8ASDP5dC3yfkEI41lXi5U/TrnwFy0vefs93+iExX1tw/6hXdnWM5V2F+RfF9zz
mBdnDEl8qsy9JpD5svdSmAkvOxTmnjaKDE6422TAC1rCuirfXa3aY7+E6qvWew6fNwQXx5cWcHND
qYG1GSl/KDOnCQv79tAESQEYVYZuZN+bWS6rDFZDeIIpCNqIvuTGqEwetO7EvPs18A4O7Vt6a0TJ
gvbPAwx+SbAnkr8qMxDx3s/c7pwhTZjCd/Y1zykRrUu9KB0YEMGyhvx1na5WOEDO5vWRyD35c1tE
1T8K2UZm9W0JkIecv3etnYd93upAEU//LQea3abh+4Sn7M/y4hJ8SbxIFVJCDcc67Q9o17dsd4D+
e9Z/3pfTYWmd9k727Nx3wYQXb7bvC3QrQj4iUm02HuHxSqEjWD3C3gOTPTrm2WkVg0GsNcHwkmLM
at1mIUh9CTjU3Ndt24j1tnv14UTPYPDdvdNQiemKC5EuxsC9lcHC2KrTomHH1/aKBXnx59O3nFZQ
QW/GVKJxxObSPGmjkTe4/Y3Efbppb+xXIxU7XnsyZs6dwkS26aDnOKDzZxBcoeoVWH4wdrVrv2XY
Xyd6/Xgt/NqE/JazyzBC3D+n2ePSMH6XkNTvanmssS7/GUS+x2FBMpARCiaQBPmoVQxTXph7XwLS
yyNMkA1XbqSQUGagDt56duo3TTojQ8CC0fO3Mtc3Fwpi4ieYgRhrSvOnExMoWp/h+tI2mwU39PYT
8zbAm20qqWDhwb24hUtDqZ94/zzC/1AUK/fCL5+TOz+JFO00kVxE3PYWwJYbTx9aCOmqS5/EeB2B
RcO2amFBUqmnqqSTC9vgCul8FvKWrW1vI26q/lEF7e7PhLC+nSjNKApF9xDERsgBOb2DZb4QUvGH
eheHn0GKv5bfW9WFFJxiVCEXxwu3j3CxdCSQ3ophQCuBez2FyRkxXsjPNSIUs7nf4ZuPYk9INZgM
UFrbW+H8ugWnkwvL4UFocyYGLTrbbMUXn6kpL+YDlIDOnBV4PhEACxVzOtAOY7oIlrqstGuowEE/
0QTrkvsdFW6GuyHzwFUe9azzj+iDfHxMQCsikQmkuldDu+o2qybSuBqHgP6rq/B0rXCUeHJXejw4
uvCo5EtkAYMdJGR/SCV+UWgsjYy+Z1eav/NyP1u2+pyhj3qMfzuqUzfMkYpvciDngLzStpkzpJo3
1FhWuKGjd9sWHuv0TnkG5S4FrXUtz2H9slByoXGUVejIXMCH8BIm9p46TgkccgDErL9H1+46E+No
Nota/PyT+jEpJHedOdoXR8T4E6QqUL3RaJ83lETkD7gA8r8mYulLuoCUPYMEBY2wcRa6dKoiEPKB
vC79QDVriAIvvKGJKLMqhECRsM0O9DFWNmZ1NwPh5Sug5z4vRtgClMb9FSSUtQFi2vTVroaESTfO
5OiWY2ZOPleixCVXEUpr2GabsHiNB3HVkgWmYrlMVxv7X3OROFD3N4u+cuDkfmDJCIDXfQ0cVf/1
yFxpY3z5IBOcnoeKMVTXNHwlpPrO/M5Lo2py7wXpuBhuxwX5ZNEE0JGILBcNWDzG+0fx+RnVODye
uA9nhu3DVHwb9w9nRTTXsWSBJ7pgEHwjv52lpzZZsfqFHwA1XjOhSiqFQbmTjX3fCAmXFFyGEH7e
kji+WAQUC9jnFlZNSLQUR/XE9LzUO+ZeWoF1pMGJkg3FgarLKKcP48YKzj+XXrt8UNkFZ5hFKWxh
3li/EzFF3aG5TQbvSa2TiL8DD9x5xUdMO/r2+VyBuN+za3LUokPfSJrBBCF1uCUou9xzxTMOXb0/
ApJBGYQK//FamqiNkZMKaikNZ8Px6ib4OWCgx57/p0cK3eVf6wA4H2yND7DMdx+dYy4onGRBMYJN
zZmD1fpNZEXmnNC/9I9STQw++NLEtFWL1sf0z7SGtlOSt9s/X90nXf/pznEbq/BondQwIuakIdH3
wQKRejcSPnTTl7YeWdtci3k1IOv97Hm8zDzme676E6uM6RCvoDDp2Gg1mC2uMUOF3gwWf17nvDkm
Zwkj6jPdU069azBm9sAh8OrFIMRLNeAM5o/ykfpTgmKTa5I70ptOKGR+5bsrIhp5/zjRtCz2G1gj
X33NKHZTg60QXv6V5YIHRMFDX6kzM2XV+oF150mE2KWkv3UFb4xVqA9DonG4+B0wxn1LuDzV2/fq
C+dyD4+2f+Tl+rmhiSbavHcWHNcWHyzQxUmBTlD5hXpbM4R10rZX9AqT0mu9J2H8b1vjZwhEKDhE
VTWxcThvtTgBq2fDnxAVjqB6wFBwQpTTzxDEXwfgRMG47Rzlvo1xMN9Z+n8eLh0KBNseUiqlxl+V
ERC/m8ZYB5YXVIIctagDloY71nH0J6F6vQDi7XNbZp8gqIxAAOsnD4OuLUAZVKKK/fobWtkriNTd
uVzpK0F2eUBRsbTkkC506RblEZCQofOTEikTkhUOX8it0Ow6YUqpgGEWRu0yGvcUH68qg3DKd68h
mBndn9+7kehlbkbDeMmXanEFhIx1xPgU0bSJ3o/aCJw7sSR4pdkn+MzfbFjKs5u6AT45ycJc8slo
drosIU+65q65qln+vrY1thUf5ZmvncISGopgB1hiHPfSG8GlEUNTNTHu3mRVvbEKFRm7BQ1zAgbp
IKxf1k1QW1QzCkGau10MbJ9tUB2IBuIqlU/Gu2gU8bnioZQUQrmM5jValMK2wvqDaEbn+ZE/AKiD
KeBx40jiWklNx2nxUntvOItQqn/eI3aFmaLgflXVpx5CjLP5MNAqroJMw+rL5ZeDb6w7zHYJ93Qk
2JR+0oFjNbnKL9ixp811F9bK90CE91EmvDnd3xVTlZ7McnI+V1RNgnIERfeeV94Cpyp3ayT7OACH
azOgU9ppOX4BW6ymi8hsAbf6vLM/fMbzmnfBVffDwC0jonR3TJezrpVM/0bD6QE/xDkuHLNQ/ho3
krS9x9wHvcBzeYRC0AZMFtB2YHrXyAI5VWPJgXlVp0/+DgUmbfKK+XnSu9pwVIOH8mlT1gnXUFDR
f8dT1PM3pXWOJeB1uqVms1F5uDazZTNHvAL1lXLhRMVbbmNERIbSmG3ykRh4J/cjZSVsE1YVrLV8
Gd+GBTPPgOqjG2CwaK/cqVPAGCoNlizYOvLUTTtQwh7OCTSor7tMxOFiLfjbaHNZms+FIanVpPnS
Ox4hxdNLaBMRw/D+UegU/hMQdVZtSJOrpJm5c/PeAXiQg6hGZAR0nF/nmEcO+FQlI9dRKGclIkDy
G7WOZLJm7PjewU6rFIgDao9utxhGFzQKCsHNWKu6G2ptOGzxH5ICiNO5bN5KA1UDT7VM+oDrIIWp
0oD30e34tcz6OEVQHp9TNCWQpeOJSgFQJ4d5jLAQAScBQsj+ssCzFJ8i/tDMU3WQPVROT/SmijuD
esOJWifWHSVdscQM9Dv0/vVym0FYOMbMEFug1HumuMWpSDJqq+WJigcn6iyOeE/Xe3joJ6jS/Ys/
7O2ao23tk3A61PJhoeApCEE0I4jQO2JLqwUQ7rUbUloquxa5NKOLLjLqvnaGGOrt9s9jGvuRW6Eb
Xpff3R7g0g/7gV1GlrYqoFTq/4SUi9U/672TvGu7mu+ihXrayeiJAuxHCJcKdSCNCX2iu0V+Qe3m
8iqY3TFVBmny1QieIt4myc3bz4tqT1pXH1Egu4dn2fq/PJZzHq5UKpFg6/O2KzRMIv6LTUl8jY6D
YI1BkEX6HT8khNXRnld3jMXIrU+OpfwIOGsPZIWz2nFS10VCWmm0kt+drXPALQqX3V+1BsQPR3vr
vZTSY/kIk90n7r4AIQ1L7NCidjzOIQl6hJnMTKZB1zZ/XuqbeADz2AaqpzVmxmk5yHajAvP9jiH8
9bAnoSWF332kwLpUhKJOM5UHWp5v6qXpMY2M/mFmmLdcITwIIEt9EzcHgH99qv7vy//nYUwXTAgN
ER++Fygmm2ZL5EqMDjXv+jPY62V+zxM9YZpA3GkgvukCuiH/bxs75VTAh6j8HpNwd6P0rP/H51Nw
Cl+oN46OtDESlIHItS0yH/ovzkd23LFjAUJZ1wVthorEiQipQ4TP61v/t516c2AX+DZTaup6iMw3
1+ZNgLFRdEzhCNw8eokB6YLkI9lD7meV2ivOh7hi6OeoznbsO/T0EF+MZWNzNI6pxalixPoIyGFR
2aqzlfk7cuuGIazEII8hhXIZHUmLA8W6KEhu9Eo2azwTGG370MQRcK1TkXHXLbUtsDgu3iKcRXEH
+tbSFJ1DuLRkS5wfiIIGdOllM8e3rcjx8oOJuLltOxZvpco9lKQ64+7mNLa27PW3g+a5mtn37MSd
g98hjrvfCxbXluXGn7862jLzZcSqP8tpYKZuL8+xhxzGEY1L/PBQuztjHY0508w4mc+wdbcDhtPi
DvGhD3iqPDKwQsFac5Nk9phTcWBHIB1IWCqtiYGAw5VzJ0OiagAqn1Tt5Rnp9aqe2LG6brF7rTj3
jvMurov+i7YEqaVcbbuFBDqO5hBYOEbH8bs6L9NYJ1LziGEY8rk+EbhEVPfOzd7kH4I5m329EcNJ
sYHy3bez684ahuPkaey3mPjlABcbT32G3PL1KWwllzft6CqrITyWncX8Zodw5gxzheiFEU/0tI/H
g5VEjcL3Cg8lQ6zl//cef5x9PBx8TffyCMK2kwlAj5IhIEUB+IanQ9hh52bFNcfUfCLUMaJnnbG4
XcxsHOiKqFxctw8wjPUSN1e3ESKCtFySrIcDk1clZTtrZvd+A9SA+ukA7XwR3ZRUiQzHebiR3kJ0
N9wZsVgoJD9JnWwvxZvqE02DLUlbl4w/YxJ9LOOJM7e4J7HDhr8HsFXxBdeJxMxywev4veY7AIMo
J5rHuVoLw4hreM4YAbGZYUG3N2BTAzpVUOM2u8dOzjunoXs7TEm0nuQUqdVxQ8mgGOhMHZmxSZua
iKjxSzHvZ7Mw4le+UZRB6nTOuoi002Ae6NpJimvsLA74BaslvV4IfGdVea0lcxBvwuh3vwMucFCR
+thqK+vcD+RFZLrp10j+5Z4yMET9Htcp/O2DFnqsWYdI5ytnrpJ2MruJye+JMRJSU/Zn9JbpWjDN
c6v0nvZgm3rvHWlY3EZeWilp9npJblu4/tBJWPFk+gR7AhkIE2eaqIzzwsFxeoRP2Q0Z5fmEB5CS
N8cvTXfZUmPlL40rB1SsrBgD7Qw2MpD1uyiwuTYI/SofFoqkvstvv5HifTw97+n9Llixa1731g3T
2FUrYPcvufW+x4D4XyR700p1sbpHGGF4sN9/4EEROgNUtb7VpTdqkZjEnByoFrW/xBBupNEi+H4p
7ltYn0xRK9FqrBVPnQjsNTYHSNTSPKPwPcjWd9VgZlF6tGZc3fzmtEIO9JbhQyCblt7Ldb1y788y
K4KFu8fJvBDW1Q+ndujQi241sz/1E5NoYlfjZyabFHSxR5ib+8fI89T/AIJTFQfSnCHgdSbxsMEW
Op0O4o1p0BfdY0HKifLUgRpA37hjLrJijO3TlKfiMuW1ARwhlRvZtEnTZa64E0dMGkjfL8dCaPwS
V+KS0ZRaSxtqMzNHX02tOVcbUPIUedYER+xaiZ+S3Bu8z7AUaRNzK+KX6L4zAyKte+26VnWmIoTu
I3c1twAgKyg0Kj1kboqcUiOzukfrUR85+ngrQOXV/ctpog8QrdyrMc1KsED7qlPcRt+dLxzDxzIG
cvy7hNZ1r8g0TLbFV7Ycmf2xvomvNkepXh/Yt3d4XHwFPI67DlL1M1qmzTsEChnZ3pJX9hv0jfhi
2FZ0IxuARETlyi3l62H7FEmOOYJU24BByve/W1YORCCD8Lb0pOYyWQW/ccegfti+ZDoKUf/8Fg/L
roNkoHtr5ln5IZ7/420moVJbhFgOtjve7qtK+DovJu+NHULd7WLZHBKJovlxAQ9IBB0O326ln/Zu
42B101jux2qHerr4VFNbq2mfEdpXyQ7GGi+VkcUVPWlYhpjmEAiUtgzzf08S4jMUCd6CxBLuAG8M
6HIN308Cl9MFXToZRGSQ1FYr1kRYXzOsYeqpn21LH+eP/ZeLHZ5bFMBW+befIIL8sD3apKa2PXpv
f4kStYS1T+CF0wCYz9mSRRY5zvtVoHFPg9ItPzHPwQLSuC0FG1kxBryQw65ghdhmxxKrUuFJsXL8
q85lt4nuAPSlxEtXLz6uKBn/U8hm1UnIEJDtvzyeW7Pl/EPkDBZslZ7SNs501dnBSBZ/GDiZ/eUs
7ZnfJyNgJfCFa02qHtXRWvt2VteDJay41xoow6Y6rLA4IqmyoHuMAW4U7D80AU98r5toODTD5kQ8
m62KkRcOqftUvxQv79UWxrqQHYm1xfExP/ODE2B8oZtu7XQcucn6TO+FWS3ytiH5lJs8n6emva6J
kqBnENrn12nWrVjkJ68AM3WOlZBPxvg8acjPndl66M8o9pe8rbiIUn44BJ8Ps1//PwfJDlxR9/iT
3R6YkLMpjZVlmnIJpGEC+0Y0ybu6USnvKuQnGdSy8m6HL3UtEJFFxFeIZzJC8zrGdOwmzzJc7A12
UGIWws2bVp3QO4TrHyPE2AFWLbtN4tnSyf4Z8P61LKnI25pYgzkTTHYZ4cjOPoddY4D+0kcfPVne
aRy3JqnWipRqWbMatcQhETa2RJmxBKJQ68xVPhsk2jlPI5KA2JYeYNFgQXBqTB1xWz4K14fNclDd
MeC/Cfh0IpRGhvvfkzEVZeM+8A+gzrloFmjHwMZ6jMHOhgvoSEx9O+fJhMGZ+KfHU0YUz+vHyXOx
4KezJXOV2KSVk4idaDulr3ed7km5RqMSP3rVMeiuqDD0rE3sOlFr+SSM1k+EQ4gyjMlG7EY3b/X3
dVYftFyrDA6/lwHbwL/6g2fLdBbAW/Q6wsiEAv9QTk0EHfNsNqlwdOpoBVby24C5Ykg7D1kIOHm3
vCbr7i0Py8YAKBmtm50ZYGTzLxlH181FHeyfS/ugPkpRsk6Ek0uimouRduEdeEvJxQgni9WkMFXY
rLek/8+QAJdJh3Rxcj3CPZ3svLR20uSLlgo6+GpzGcrt6wWhDJhwWMinit9ozaBx08Z3+JfgVGAt
Ra2jbUG19rOkC1S/9kv9t3AZY3cT56O5kamoVmf0WTlpscolVVZyqvs+AnucZJS8z3R4cG63ox7a
aGi4ginl+dXwTRqi7U+GEv+zIQSED+4E4enWv+n0qdzS/IKlyKABorhR9XRsJj9eC977X1fE8i5D
lpJ32CS3rENGLi+GtPsR7X8VyWWWecAWbiSRtzfrYV7z/65v1US9ggT0VNE9nYyWJVfWHc4ZcPyL
tkF2Z93//Hz3dU+mto7QpG9lJROS5b9FkPM5LsjSdBQsKxI7DZ/GyI90WTVerNE+IS8/2KX3ZEeG
mAFko2PmCGGX99AeHFb5PrKe9RwNzu/wLzHHTvpSuO5vn328b7h083chF+9p+cWdc5QsN+4fFmsp
Sb0QdlaUM4mJcTORwyWvMqgs5NNLnCKLW9dk/3SSyVVWuYGqwTQsc9TMVavHqRw6Dpwkow0eKAhl
XEoRUkIh4Q4JMkkyNZrVWKM1hCRgb2sP7MHt2xKZ3ydNAc8gnu87HbQrHepmSJrhdLpfd9TUQEyK
e+zNqj4W+rZGHQJABKEy9JIjyS/5wxjB61hL3Tvf11SmNGgcJC8zVBpJbBXCXdNqEMDKrQxKf7p8
hnUrYgXtsfqVBOzIDCKOnqT7F2bIDqP6mR392RfenKxWq/WRE18K8pYXMny7hE4A/SUaegL4OiiR
tsiMtURlqCQSOnPsdIzdMIXmAZLKIho67Ydt7ZGUWmXmO7LR0fdk8X0wbZFcP9onMv6bgkau0RA0
jm3z6o3xoyoud4dqFDyxxs+dAxVyOt+pQaGQLJIwzi7vNpWJQi+D/Y/2BFw9s/zvd83H+M1M1ZCr
qFTM81FfWk24wGUWmbEEWGnH6eR4f+R8J4TSCE5l+kLeLvTSs5R0eYqym1v0cQnXEhS1MKoRQKgn
a8napqYhPab5+ERt2BDqR6PzTB9/OssO1LOa0W/IugzqNgV1JgdxVnc6SHfCjmb/6RqS21SjKMj3
GS+bYGvQTKbu7AVn/ey0/i1XN7gCw5XMQ+8AmFUxgKeD3FER7fjJ59gfvSQ/oO1jf88gYzmJ/IOB
az4gGdbL3jKVLuWJHZAcaTcfdqg53m5fPZKuzNq/Mpx4MNMVG3Hwee6r4kosS/vV+szEypT49/K+
qKPl2Ldt/NMDBQ/flnO+owZSQWd70p2eJVRPd4h5c5ICYgOcuyDlratceq494DSyfeD/g5PmpeUp
9wadB3XkyQ3e0n7yfqXuLv92stPIfQZMq6RLOyWWfuS0oWVpM40Ik9fPkhBAJhkL6fzAu5GygSNj
A36V9w2os+IU66FAtBcnwqSwrvx9F1ibeVgsADWxADoOoTurIVSsnLNAPt94j08x385dpr3wRzed
528Gk37NiFfN3XE4J8kAVqLetKIZocsgfTt3Se5vE6gQtqgona2Z0kWtdnVl7BIozwBgjM6R5QU8
00xkTImxImGOJ47iN8O3CSBXnDnzhFPE38xm0vmtTIwNygr6DjRyM/9SjVlLK2BWlJ50t9vWni/t
wNDHnhXveaMkF0YCY5Yy2fbiNLDzZYbRExwnMw8Awz9P1EpWQlLLEov3A3xp80NaDgj67QlEV7zB
ozxD/SrAum+/nq21cPoEQZgmtV6N0xq68bPGvkJ62bx/QLxoVMGloXOHGh0NzvjuYTjllut0tujD
ndsZZpkYUw6vXpjwB1gCE7XNSTK5HNBCKmMZF82/eXkV6+a2Bxe/VVoGgqzgcIvbiRpl5Cr6oAU4
tG9VFprnJK/BVX+0vetKrvnOi4ujc4LQoN1vDV4RCb76ht3usy+PF3D+YWic5l8SsYE6I4mjW3XK
2z536I+SCd19adc0jugy50uBlXZGA61hp+1SarLQYUTVNzSrEG8pqHAAO4FjQ9IyJR6j+QhFjkgV
QEF0Q00j1sKQa15/FG8COQ4xQAn5iCEitAoXKaB7IxaiFH1IZ2vt9eC+7+vOhZ7PKgPXLjh3j5ts
W44StlSGaHQJOZ07YZuVbknu9VLAJBDNCASeXxHYBCL6S1yFD/jHrzSwlsRKHvpTAC1cfyAEyNJJ
BaLIEz+BgfComHDWOX/mOtZM/E+hO6+IZAnTT59GyUtvUyd/AvgCxv9Ehcg7JVbOEJwOYP0ZfJCU
1vpV4DRamPBB6GYYnFE8CCJqZVsEgEUvHJrcKcIhjDi4TR8jgREPZ5Ss1K5plQdqGt3h9SpjWkYL
EoM7frXjHtV6wU95pYbIq5kdudfDgtVMJNL4BdZm5BdQOtc9MT18fxu7d/dqbTfvYScDJB6YvSmu
bF5y7Fj9m+pTJzStaMpOZGfX2BqQk4fLlPtsFNk8s1pwmDMoLU5Kk77ESRQg2wav/cBFXvf3Cd4y
BaGZ2+07b0whLPGfK8IHiwnrdgSBuVlk6gZ38hv57YdLNLRJz1jx+SimB7zlOLTcAgy4lz5/9zw/
kV+5WCkHoHV+/SusKZFyyua135SATW/qWh+/0H7V5b9mrpCDa+rvfs28zOJcjm/pD1mxI6DE375X
eHUy3vtvMr8Z6htbVqCkhwDXQ99pmbrgqW+CxRz6XeDkfzV+eE84zRHmvhhhVAEWeCsropLCJEAT
BgMLYdrxOSAEo1qi15X+x29B64Q3eMyGTd4iVDqPD+T4CsqTnoGh+uGCrnHqHMQ9coFKZV7Ze2rL
MGlfQDnPBPBMpKWwx5EQhJrAMGwEmzfklVQDyKxzolGbawKYM1fSjYJs2VnyJSqHZxoazkQrIQma
+5M3qbtQig5lzza2oCiDcFp25sD+Kfj2j8o8qJMJVOcr6AXgMRSZtMPLaxuup5BYRsEk4UGbXOtr
S0TzevLdhCx3uoBgtVVeQTmkoWSURlUre9aQmk1zL6XTYOiRBuLQTCscrOxR7u4jK8//XvJPgwe6
8lyBy/zw265/0E4wEZdgo1Jw7wQIe+a7Voz5RmQKsr/zQ4Zwu88c9hm5rwzfIzq94G6J6sTHYnoB
ou39WJm0YRi/z/UmcpE0GKELnoMwrBRpwk/RgCWPxMFPTNorr5Iu8iRF55SkMQIRA7VxlCKHchpr
gt603KxoknRMKaCkcHiwv5QMrtOSsv4iq0edYHudzLL+98sAojPckPLGTGajHG92Yyk9sOXLi37F
5IwpPmaVtQFGRsO6JJXmzE5tdR/WUy5g3tLq0+QrcnDWpwq4mHwa8xS/hChepXgqrAg+ycdw6mww
9Wt00SFE9sfdIQHlF+4FzlDfz3Tc0gzgRzmSTISuiHBb8BIG2YS7WBnFCC2Y68NyFM2fLrbDTKeG
eugPjfHP+K2jrUlp7p11DvBt83VMASaU6Y1sQO4oN+o0UjNrSArdoEQLr0yHC3qm2m/D88vHGMio
EJgdHyxrqrZ1USmEHBM0aJahLNhAT7RdLQ+PE2Hyq/cAAnuaBnXFzDDQ8SNtPvJWWOQYNaxMPvEX
+q5ethq/u2NJK1pvSjHusbokhndU1gEXk8E/cMhn/el1CwwuqgGE4bj3WNvtw88IRiAV5JFsKcjJ
hwIHSc+rWXL7UXZJLCtLOWUwsqlSDJtfMa6HLKD/drLCRqUI2qk+6TMTfB6lkEDG8OurECe3FD5f
aOf4wyQukts+XfApEYCBD7nSBoT4Ez1lN4yEQQxbejKV7s/tyCCPM4oS3IXYSCUWzgVghJ7rfRTI
a2KlrqYaRqTsXZEUZqW6VqRoOpROVPI/UzVc95Bg0QXQa639Xe1TuvL2KvhzYNdkjE65VooTmzCX
97ZC3fv4L6MrcAuALuCQc5DcOz9hc74gRhcuF9jaagYAQbyQX9/TFW1aIpRUtfXbZQJwG7UacM8S
7ocShbRVk6ikF13DF4ZQJbv0B9yVaWOHO1x1txD4BJPeMWoPE3afjHopkbLJTHe0TMxItEgNDt2Z
dLfp5IOjyOXZupP4c3RyBAO37Zm2Jb9Ck/17Qao59NNXHUnOunBoHJKjA6yTkvRvRRqj1CVjGdoF
ozHD67tcqGtIHuAb3UkDAO1y6KXalbp9p9l0v8Mwno5uR+sXzu8x9AWziCmk0o74pNd4nL1Wb4/r
wIasl/jkPqAkXBrpuIWkj9uxiwoL1cZulbZuak+DPry2oM78axJ49ME5Nl9z5Rzd05wM94PslZjS
LvmY4zbJ1TatKNlU463HqIymGbKgt7e1j1k2U6qbChkgiMejFzV3zLmgmhrR7nGNjcxuYcpOo0KM
aXiaEvmnnMsRgsc4Auo3qiYsX3dQKM/1GBwdo3uBhLkpGkPm8toE6vpZAh5/DrTTjLqH181TnCwj
pIHquoZCihfqmOiKTdDfO/9sJ741XE6bwyfgZpxS25aTDWVcbEgA6nrUGfg5/RMBqaFeMVuM9mWW
7NSnmTJMkj3pCEMfO7IDpcTtzqE3xGA+3C1BgGTZMJwTBC99auTxHBIjOylqGhBqrwpUkIeXLZDX
kheVCdn8fgnuk3esvFEA0FeW394a17DDIN/XylMn3mZY+yy1WLE+ScGHl7a/ETcVIilrZIxOEL1q
YY+NCF7k8M3QIs6keyTMA/2hYuExmFlKLnhMwehpBdVBWxh94xEU7Xe97p9TpeafRcpobpBQ2GdA
Q7zochAB9s5MfgMrSRbXdvChOf7zDFPPr6cpfkL/SV6b3baxX2qI+FPI+A5OnKyCn5rfyryDNE7A
Z9g5U2yNLOx2qOv4kubM31JNotzFHCsFKMpPNc7wUSKNoCrhy6A0KVh72vyO2+7hQHKBkNoytG98
kql1nA3rDTnE2UFtir2zZXuiwfw7SpXgbrxpMuKUvCKaCJpNurYLiIA6QbwSCZJg6kfdGpIorG+c
+NII/MZW2k7A/nNoUFvf1lYGj3QYav6hfpZUOFVHnCdATXnAKYqVur72+Kid0VdwLSvXz+Ullrp6
iGg7wr576IwYlPNG4jSx8PKmZ/QxvPYP6wnXYERjHO+ITjQoltIy4xeAdbcXZA80H6mQDu7Fhaxl
ou4xiBonPMWuVnLMT1eiBvdYxHYURT1cIcdMG0c7CNA+3bKqC/TylDJV30rMOmiJqnbKVTCTSL1U
ll8dBx4UiaxtxjqLFAU1C6Z3MJAPxWABU/Bkml9GxByHERvEV2ZM1xMPiDJjCPYW5uXymZ23zL7r
wjvFmOraVI2wxZ4Qkcn48W4a0oJ2vSFDqNcV0EzZ2DDZbujii4BrNMTwBo1ByJwkdScP3q+RD8GA
Wev0boux7YUoUkQr/a2ouEI3rGgI8XRh1fDhSNED3p8jBXKKO7JqICMoJKOS1ubYTgYaqTJum2vY
UyVUDLqGeSSfGuNsICJeeEx5I9gRyjeakbn89jZYX0jG0AJMOMH81QOki4BRkpJBhOHDBzVWlQuR
IPRsccs4KrnEDfINt54RH1ipc/6M/hGYhheKjiOTqb1jh+S+TPZPlWusAZcMc+hzWCkVMTIkqubG
LV6Np9maE1tDIIbvlwHSr7ds5eBC3eRYfUNZCC6GzQsoA0aD+6F1SE0vr8XiPv+a4KGAWMrs23xC
MiqDDJxqv/mkHI5TVSv9zeImt2vfkn2gn4bJ1pcjtIKTExTf9WEAj8YnZ9nUoLARRQRs8Txjrga1
v0q8q92fEoM1OeQ/pmbql+FqrfnmYtmRueiqdW3OOqfTkhd/Gr5yKRNpBzguDM57QEb2Pk0P7lKs
p0NQIM7qeK12ERoJUrwvW1EFItubc9iHMM1dM2UydVabgnzEXtmWOgK1psrJQ5XsBTCWOHDzOTSU
hjpV6c79XOpFynMWDIa08D1cvQsQnPO7Nf1Y1wxFgUv+9aw2xY3uCxKjWKnFODoEelWGY/Ag8gmT
HTMSKYQ2XUzJ6toRBBZCJ5Hgt+VqWd4q9hA75gcgw25A5szvg5Z5dxKnNkLuhgaZRohCODVqUnSi
vr/f+IUWrlpT0B02I95o3Q+ei/Qd+gXcHfXsbxEUZOFQZBZbm3buF1EhJuRf8kiMWm2emoCiHVbk
AB6zOMgGD/zmyn25WiJMIj6eCNT29inyK43JVeSplgJV8UvqyNgshunbZFcPJqRz2WbK13COS4W+
5RE8jxanl+JoDpr/y3sdsFGb+WVyzMDL4pb+R8NL0fbYlst2Sbmx/kCl5Nr1TX9KWQb2jlIdoq8i
iOq/jir+IXuWDcMwCDHnFvl4eJ/y9O+cQeeFFDz1HV5/jtPQQfjQnhzQ+AjszhlVthQkkKfeoAnM
XibeuYeKwUZW1qrclV9uZ3X7o5tHrTUv0HXM70pXbcOSLfNlOVAsnqXQTt1/3/rwTBzaR2N87svV
7PfEkiFyFs9dPDwLc+G9XKFd99NQ/Z4UKRnnXViT9rVg+xABWjEooudYBYeQ7aUm8kZrXntxW1fC
zKpaLgfYL3H3AMXxaNHvX0epGf2fTDH525p/d6SDCxkfKR+lWZJv3ubmwXR/WTIxkr7cy1FTEuG7
s2+sLKEnpj1LMjdXF5zK0hqJMP3WP/CvkBCPa2+tWZgedSywi4lCk5v6pnixR+1g1UlIrkJ+ABGD
e9k4zfK/7SZmY/i3JxyuJc1Szb4GZ2KMC0CLUpljKNfJBJjU6GuB7oQDVA03GuIx/CB2WqrNZd2J
Mfiu+Vp3PW1xC53l/3ro7AWW9+6yGDIJZ8K0cauIDFbUr6Yo9sibu6yjbK1WMw9S2Z81CuU4VLs4
SpNH1p11U/web+i19+0Ikra2NwfkdKNKREUlpZtRv5BkbRc50W2bTwdJRuv0ANd29euA0MLZf9zU
1L56DL93CHuVi2kB3bKFb1Sl0ZaMX1w8fxRKruQNHWFRAgQYTTKmzcqnxJMlXsyCWnlia9Q+SZwp
YBCAxdbJM1I7sEUkcfUEkS4WYm4k/Ebs50FH8CVF3QyVWXjaDsjQKf7IBcNqxVoTAuAyEJAIU1MU
zJxs7o8PNkT5CMPwZiRu6HxE/2v2dHCh7g4QUNAy7dhqHLgQvtBaTn4Nwj1x/H715SKIRCdmrSs9
rkC/UhGbZ/r1xawvQ/DehZDkkVgmZeiSdzb1wMd9tkEUeVE3y8U9KaOlPrHzUWh3/YwWH61LASaj
5w7EkQTOhGT/A1Ch+qdUrFw18R+E/rF7uafHVO4RSMIh59opkJKycsIHAyxRazG7sT4oqmWiUmSU
8U+tY4r2fqq2SogBiFcFN7+USw4opzBaGDyQHeDXj0XFGdVzXXWa2qWSrBM43lNQQrDR9FT9ja9o
rpL5YU4bfKmy+i/bZ4QBY716qeXTIRu9kwfMKEhQbnZxiAFeV7xHzzO/zhlYbcSO+t1y12gFukJ1
qkAvuzI7mWx/gRyeN4zChjVXAaHYyqK9g6lq6t+j3jDSlF4klr/us4uB+sl19Fk3Qbkq+p13Z1Un
DZtVHgr80voHl0PnHnkaJcI0FkULygGbdkmz9NuLGgRVuv+hSSgL6hd6fTX1/1F+v9FvziItXdSi
wO1LhZzDGdMNwjSkB30gCdEJmG6F0xZBKy7hG89Bo5SkSxN3jSubEGf9Kr8GI2/P4SRH3WKqPNve
nM1KX4dQAPBcOROm5hSViAolf2ubsp07oK/9daRSJ6+8XCJIYg2r34ECr/+D1vxQQ1/4BgtKcOP6
9Dr2V/QzKYaO37dFeMQgbN2r6K7hIwe/tJkLQ/EMzjFmPYafKYvLwvkvAwXUKCNKYIf9ZO/3MRGu
fhg5GvxHORBwp/ipeCzftPNv2douDpUjgzEM8BqHwCBXzrZ4DM4F4UZPy2aijGLjx2pBY5Qj3QUu
Z9l8BMyGcegpUO2Id4aH0mdZBcqC+sOGLWp7z5DuDMiqeBzN8Z/uJLk+or9wzKQn7hPGWVwMi8vF
VUj5goNTr5tBeUM29x/vggT7ch45QnQQl/6ESmlFBpJ81rJColIdxSeRAZ7iuN0Q8SrIiMaOV/ls
gmzPXTvqWkIWtrpruDGO3rmQoEY5XFqNQGctnSRZ/6miEgGGPkBob3wyIhNzv49adZJV9PGm3L4j
3W4NSumKxIrHaI6kIib3VjmDYMisNdskSLvCma0lwpJAgz2B1h4jrKh1XtdDbPgqIZY923HrwClf
GCY52GyEumOnK7TBfNTxu7UrrtBabIN0uI5VQWoVJBzO0nbka13AZ4uck6QaV3bBXi903FaEZxC4
sy9Q49pryTSyhrGL7OK9gRmH6CZcrB/itkpG724ewiSqCANRIO9h8IKlRJVLxl5piSKbMx72zB9V
yESxoUnfJlXNRv3lD7JCJ0nkhpb5TQXa40HLq+1WSuxnuXSa3x7cRHuqcencYt7k1zLgY2F/eNml
CRbJTjjDv6EMjPdRUO6SHkbDhhA16tmeSBVtTt7YyTyBlcDbb+8D8nukhGJETtx6xcYIOea1bWnX
N+53C7v6+nXAMFDxBTPRuDQJOsnR6kA5VgU+9Wyd+MMIPaXh9v9PTKbakrXw/MJc65WkYdWWgUwk
Aga9FO3iMw26FTYeLbp+pkDfMyppmTw9gZkEiFKBEjGOATHoyEdh0P6l/gKEktVeyYUX6giZsllF
z6Ohnhd3kCQUPF2pm227O08jiiuH6qjCgEZsOqWq7FytRX11qW95B9vi7gea3FTajp6IH3cRX0MK
goCG2kM/rudozCvC/9krJIpT+Grm+SlxkeIHs/onLaDcIxQGETC/2I8JERw9PJkRu+aIykxUfNO2
VbDO5lolrs1wYuc/BcGsHD59bM5rI5WmuKfawOTT5auT7nq4KJw5NIAMgIH9IGfeDcS0Pn/Y2G1E
DZ6/18yuvSsiQmg56CJyFrPMyhE5kMCSc+nuatrzq9eHIJqCm43p3IimieHLZfFdgO+cRpS9VE3E
Gm/fUuukfEM9HOlPaa124jkyJs3sWeZ+1USre2CGzUeinHOWp3XJpEtX+RAQXQe4l60EzItbG4Qa
zrJYbjHCmkkkvm+u/szKE/03ttPit4iYibh2Eyv/Tj3EbyD+fuz2TIG3yCEHa//6Plbm9ov7Qr2v
Jq2gu5lgnsI9vOwR/C34etZchP54Ckx/eomGfKGxE0eabm/lNuQF6R9OZIdGRFWk7uBE3JyrJbWC
ZzhysLlmGOoAlIz3GiHWXw0ysOOKNN7dvfwY0xe1tqkQc6tu3QZ3C0etMglVx8aRc0M4ZJOlWXG7
c6TJyoZ/1LndQvqYMMh2fvaa0WGZoCt2eb4ml4YPusMpKdDWX20iMvz8JOCaSF+d1KupQFV6cRo2
UJfcVo8auPqvgD91Hkzh2zOQgQc+M6cIMG4vZ4YhzE11EfVwv+JzW+uS8SNc6hrNUcmwCpk4HIGs
bTorHp2QCP5RK0RJ+SChFZePmXX4onkO8gY7s3IQKk+YEPV+/fojn35uqVD/XNOPjvyaZbKRJbTf
ZMgbzLi0/lHeSRV91ErqdC3UgzDISteuSVmy90obRIL5JTWozBkKLaO2RiFJ8peZpMPc/yYyRr+h
mWdLDoZ/AAGg6mullPH9r0U+x7vrClvNKNB+1GXN1DUSGjCkEV40rVIoBDbxSqFxlC9upEyZcSlt
7CkCp8oWSyJlGbcxLvJ10GoqRhGBiEjOy174sp38hBX0Rbc5+alKp/L2tP6nZCDcin32okK9FCfA
60eVtSeQe60iN7U8oRZEkoeLgEJcashNekyvcP9BijSyk38Q6giIhDxLpXfkUn7DnSmQszUWmcNK
LR+EqRxa8nv1bs9GV1GxZRiaeBK78NaKjn/H4hk0TTlDvqfuH7790iAR8sxYcKH7uK+RvnJ+l5jO
Fdqs2alP8eOjncZUx2SaqTR4A0OOFeOkd9XTr9xAmQCMqtdUfSo7zmJjJB59nMrOASmax4pnPiit
Ie5ne17Jm3wrhTp/uXM+ThUOW4PWgUNofSpCC/l6RCkdzopNY6/GRMapFePR6LfkHetFz5E+TCzU
IcSnLHmJxKXt41AR+Gj91FM0n15K13/lBLz5e+LcasknqKr0JwFmYrrXTkmsz+ShlzTb3tdhbO1P
7Dpge3Vwz9CeiulYoiU3vr2ZW1F3soXqfjXhhYGnDL4vwzgu2ynxJTOXdloGU5Gq6ezTuy85bQVt
bD6bZsmQb4W1rl5oTq6qGDCDUT34N3mvixQoXi8LBHjXWJc7pLjkLvJf9sYkKdQZ2PvcNUXe9Tz5
rZZ8o37Jql2RoVYzSdQeS66N8pMQ8ilUTicPeOXj7zwa39fv9mdCYxCjpMFXauk2qURr0g+miprk
uZXlweLBzTesSsPrtDe7aV3hrmWE+P+UzBgR9ywQGARhHMiv3MBaxkTbirsXYJ+IUNug16Tb20qI
ZQnc2v1sGmu4+coUNKqEZEIChGR7SzbBLpzR7kwlwGw4MdNvyVNzkAYTmKw4itOcj/kRxQLV/8CQ
IpenTxdLh98bC6/5xQ7x6duKktR9NC34D48Mxb13/vkYwCbf7hKC4BJ7dsaCeg6uD6Y0OmQnNlfK
87XZn3S3ixl6LMOqSVf8x4uv/BzE1Wh7NHXrr72euTXVNgwjN1bjO21WyQSp5Hw7Ymwhz7vqHJns
VV0oIZ85yy5XuY+xWIbiBn8P6OhfE+XkLgQolg7XyniXf/Orby8ZYeq2Uyh4hcVrElHbqU5OkYFv
HwtU9ykXH4h7gnTlAdcb7gpaQfwmN6i8FyDFwSE4E2CTBnBnDvUqsoEjQt5oblLmkBMAdVICe/8/
x/5LuwL2CRRoGwdScHhVXKYhA5v9aB9DuiUrtSH5YR+Kl4rQESv2dnABWj+L9Kk5F5FQDPoMsvDg
u9xc+cM51NfZV/+siX3dn+tqxhMTaZROKbSJY2qu626Ix6IQBWYRe8eaFxzWT8IUKTiimu6IPOxd
0FGHpWYH47yM7i0vNnJCLm2zaCrWSJ6AYRAPMIwcg+s9wB3weWNZ9r+Ew7h4o+Q8iZppMbQvSYsJ
NsOiKl+uaYYImW6yHItW6NPqJ5XQgfCra2biM39kZQVzwhp9D1ifzuFGLldYSh2pKiBKWQGZ8LLW
G3pGWDyk9BtvEyS4FB8huy01Pc91i2s1oKG4x5wXn/6hBhjgdDoNS1KyBLzBivzgMTIskq4fs0MD
LpTrlFSYxleuTKlllS4VLdqP9dpl4DD1Jj1eGJsqKbmVXPsmsdDMM+WnVNjpp+5aHJojpJdd2a1D
9LyirdNCLj403iuhWBUIVZL2mmpsj3hFhSunXKEMHHpdgkwtWj82JgEI5pEN5/8nmd3ONJrr9xVQ
qvb+5iXOfQYbTmju5TGeZ8/WrA/cPTZS1XkVpY/m304Llw90CTd8hJHGrmpIkTHWtP+c1mdsD0VV
jHZJjpm8wnFjNY67rOSo9o3g7oiqBdNTBltBV6k102/ASyDqHyVoaSGtY6TjxSrmD66p5j4IG/eL
xqwfS/vSHWLMcGhRSZCPSMGMprvvTNacSUC73Lyw+aXmGfdN1VYRlMvAocHI8oPvLOS6gqLIsQFz
QylTMVuyEFblcVpqRhBG3IOSRPi40ppVmCNCdnyZjuomRd8CBYDzvFQwcGSa6JXn0Oi2zZ24QTGw
XnE0WX0aexYxwkOLboZeCRTh5ob8wMw5FJorzNexGzH51Qr9+9+NM3UUJGsJtdd0FkVk7+2DRrSX
hMKRyJeG0Mi6kdnkJARVtqvvgDvcCpnyWyMov/12/IQWSkwafnEgeHZs/hzvSeTVhdsl7KCRTYeZ
KI36kTl3jlQoXrltjjd9CJoOQxVJa6VnC/j532lgCvunh3a0iWCbw1iHlK2ss850jsvpJIGz74GZ
n0E3128lZbFrsZZufJu9VWWhRt1RL9+jqihNp0Hem6EILYAAjTCWqEJ2BEZrNXjKn/N5lESjBunX
sL/h7kK5Nxu0kdYVgVRIxJxBUfZdt7L3MLyoqrqj7Y9RW84ztGhTeK997wJV5CnqFTJf/4gOt5T5
oCJ0iypYDu6kEJmIATn0AoLduej/5KQvnxrZZT1fAbXag+EeAW46/iHWIM3dzOXBVXdC8ILIxg30
FHRVcHQ26n6wOgn9upsL1e92MSsRcMQaqvi6VKoolGpjTyvQ1o8K1is9ZS3ii+JfHSDj3BHa1OjK
nHHk89w0icWXIInluulmMNz7WMhe2Z2n9UMy5Zoi4Ohx8c3sp7mBpE14MJn+vudmR7QJcT4DDUW8
kCxSha6tbvczD1/LpVFcACsvMPbItaeDZOuCis8/j+SU3zOXXI/u1Hit53w6YEBrZzQrkiHUCb3h
LvEmNHaKMxDhsepOIuLTWwRyexAS5IAyeJF0Y1WyFOtIE2M88sRXriL2s4iLSUEwg3unRptNJpNG
jJuYzGCaMdkXRr/WxODslUGtoyXpdgztPP2nDPbJLH/Wd2OWXu5APCx6vzIvWoHVrN1lCKLWwQNx
Ld6temM/twOFQoYch0KOCM8N5ExKxbW4LzzMYNdJkQdgC2+w54QdjbbhB4Ko1TP/AUpDBVMPPQQX
21boGsfQrunjqX3Ue9ywLloWvm0mAsqduYjpZsQ+r0YKVlym+I7KCpCh63PLUlNB8/pBbVhtvVcL
Veqb6f7gZnh7saflR7RjxI6U8z+4r5+9GXO9T/INGF4nsY3FIpbvOijiJnR1RX3tDnLaYBw8INh3
KA/7aPCIrAv1OzBjOTnwBaGrxA5sZHW73vOCyUrOyYyKlIYEZNTjltVH/DJPrnPn7e/db9R6oMBS
gpb+wawVh+gcKzxWp7UMyPhwqR/pLGkOkrqrJpTBIq3nbDw3h8jVDhcYmYyki04m9mDIt2/9wP04
Y6VY44bVk+3Sz76DcBEuLkUjpyQRrushrjpk5oDgRISv3CGmDsIOwI1d1F6Wcc0p0ZXqIlm434sC
X775adgaM0SyUyxTNrOgDbYL+fPBY2Pr9oAsYO0ok+qIgPUDnoIsNrCX/g+GG+Ss4RMzhRzrMfiP
KUs7QKIXbAJP6FLpqf08GDfxaTOdnsNN7+jq2nDWorKD/lWtfHetp5Qo/TDmImbhS9OkPu4bKekR
QFt1j35bSrT9Svrd72jWROoOIO0kAcwM7iLf/9bJcsXLyX2dyWEEkm7Hk3mTy1AHIf2xgnXZVlfv
T/pEpCcHSuHlKOsf6d9P9uCzPasPidHUzyNt/+FxP7uZ2BkZjCQoQ4dtyuDL1W17g4zW1c4NeJ1w
BnV50N25u1lZUTpBbcr4yfora9FIxk1aMCSRLz5RCVJk0Y9wEgBRTzvsjvUDj1z/PnoTwPCcqdOi
IOgFgOOQpkNChzMrSgXLJMWHlFQM4S7dyML9iQedgmLsexg9ZBdiv8nh8Ng1na9ySJfgcyhPtv3n
vLSBIhi9vuc3061Cm8L1nMtA6uewNmCRnwH44N4VMiAwKUTMHT9nRqG/c9Ch4GTQ+Q22f0SpW6jw
/X9LYJNx7RR5u+9DRoVobDrEM9I2WlnXiYoPJ9khEON+XB3yT0H9nwVNnSizCM1lwjvlI8OEygAp
JPPgk9Sq/Oey+sIAbHTnPA0tUwDqAYvqP99aq4hr4z9hccI0/WDVkCeHuJt4TS0UIilnm4MH+qk+
Yb/+Lg/zzB7wpLFAD+h2/LHIPit8Gfps/3LV+pWaU4+qxzB4dh4jekINxHrWnY2S9oysL9Qgs2R8
jBfGTT8C/VivEEGoNALf+aVQ0VwCvK8aHc8VXC6dRcXd0PB7xrPtPEq3fqu8Gnp6K/DWayY3NIPK
91psX0eFW9vz+59IrC0x2xLWI4sXTHsLptv01y73RbItgKJ4sQmxQRAMjgl+sY2oi67gXGjKIKTR
2rnANUusP4R7GTlawtEo5crq/daI7UL+q+ob65BK9lEoiGehnDLF4157gNXxGn8QxXw8CQ5iOdSa
g8rDCvyx4KwmhhykcMt4JXpk9NaBTytoP6SpjSC0NTBoaILKJtxyQtgLtrJ21bGWX5i3UryOpmgU
6j2qa59w3C6+pkRMn+cpus4oBK9HKXTGsfOEGLdXF4FTC8Mw83UhsNvXVp20IltvUWN86QzHKr46
34IW2aInm8Of5HOelRPIXCTuhWgYOwdLl63Nz/bR8nHnemNkd/VPv8ow7rmJdwCkCKHcE3T7TIjh
xMxh/METgh5aBSwFKaIjCcMDXoyP6l+lc8jLzSHAr8RaeojXhiOObpXmP9M7TlyF+jAyGXgdqwaK
P2lT/QO1akc9y0yGq98keF6fQv19xeuVdilkXsjM+FL6HdmyBNQWfb7Ynu7LY67LQw6yAGYQyElk
TeAGUh+nbhwcv2Sar2wbo9vfMSQItHf6BjgVETV7nf/1/ovwNfEhMzX+y9wIJ/o95J980fgwSzSf
Gw8oN1vdRMNlkQXqIbC/OmuHn8ioj49uNHxL4Wq83Zlf+iPsRZOx1BAkjxwRc37xMWJKyDuR3/R/
jkLZrx7mqOroX1MYR1fvZkYN0c6dTGqmkfm9b3QcUxfLCnQmDkYB/N3Iq+Jc345pDZQ4tT3fespd
+7LRtg6da01NQa1m8MAnFAdItlG7SxfmVmiGBv2Pdp6dpmryDnM0sWBnxlr3vIoIQHYRgDGsMF6g
tWC1HYQQW/vNdK5mabnEkae4MQQl0ifZ/MwtTX4xtuiUql/+Mt2kQv7mQvEzF+ej2b8KxvA4whzt
KZ48SgHms3CyksmESwd8rV42eQFkRDTlW5RGS0kW57rSPq1xmHZed4cLgnFldqRVWpI8V8YC13Ay
5juQyNfglsmZysY+O4hfJV51nKA/YwG1HH8AQ9Eyoc4TxV3OobCqPo/oedVMH4wZa2pgMxZbxABY
3b2GfHDzqiS1jmdx0xuJC6NBVI31M+mSix+ja4Yt5dCiiNqPh46OJggW4IqXfnA8B5oGKSDfYLiK
3u5MH7bu/CQXbo4Xz5QWlskQbaJy6FPVyDf9xALz2AoWcqdiMgdWkSclpJEBkjS0P3sWCkK9Kpe5
d9a5IcRrKrpA3KpMIiyJivqGZQHP/FynItAKR8FvqWYXHZ5bU+tpsjaSUyZOmpXJ8SW6wzwxmjER
WxgSRsfLP0MMKfBUKiMAAnkoN/desUKnYDcZEntIaeDl9qD0qJ6KWv+zmZDorZbHY4TPEWKS8gzq
onq3SDaS585Oe30afgNjRTQB+1CNziHrh3eFIuENXGGOxUllCz+ItELBm0CYbsEIXQgRqwOyZ4hR
tffqi9BTEf0SMYfQ83w88LqfJOmYeP732fkjf1NVB4LrmcmXJMctmJahfTg0gTsMRgVNR7ZEiIkF
XrDoWl54cLwqmbJTRjUNrybI7bYcwk8l8gD74lZzzTHJ09rvGNzRdy0RMtKGW40lb0r7t4NTSure
lU7i+k3/Qp5ljksRTude/KiObmpJDXY/kxXGzVHH2TnXlD0v7ZeGJckzLf5wr27FFi0vtDg0rGsT
6fKt/DN7Jih4TbVAkghpWTZAgIFA2fbYMPgTnm2ykKQkxeGRscYpjO/gUgLWAt9Uk3DOdf3nWj0M
FMpyjgQC/Sd36l4CXbRi/m04aq3O+PtUNJqcfcdK8yp5/2NvtUbEHWFQ1r2eJyTNACGsOwUMOGVR
DTzHmSfIzokCtop3l+q2uXWZBc1LAp9m/rKEUjQenItgcsIS25oRATAaxPuwPrQzmxJGYwB29zgg
lMtdrXhUMUoAh2wxxOX+U05Reo45iqe8d2ZBNIJhbAErzhh43nSYtj/4NfgaCFSyjd4TPJVZY3ed
G4z0PoE1CSeLA72Rf0rwG+ccNnr95o/YFHqWq1n5/poz2MVEAoKcnzA9EpnLVJAn4NFdCDGH/Fmm
wdsINnzSo55+w8paJMODRYO5z6DBI3kOMTUQif5DkuIBiANrA8NzBXTOEC6Fw+xRjtQbNP2DL0WX
SMnOG2LZaddxEdy8XuqmIsoN0NP+p72QeoG9pf27+W7c+wPHjCnbi4KgkpaidoqQrd9nRWOXDev1
cU+0imokpjbYDm9cd0neqNepesYJUxiQ4LjA1wWTj1ODs3WvTA6lQXSpib3UY4pQcIsjHxjTOIzr
5VTDQhe3VCU2GNgtZXgXa7LFA/6ItJ2C+BvATMPZyrzUyPhmIexRoHDRxomHV28ozPRSFHy6vNTO
CXiwmrFW62sQMeP4R8GK0hUJzBm3GqYu6jWnKcjNzA8K575tHD6cJGC5LHEmKEwbVm/TUSBsI7FA
VTSFqXHfHypMhRLLVSz/msJFPIvrxuAVi1BlgbTd8PUcLwYghhkZYFToQ5XNvqPpnK5nj9gAHgTi
r4gv7+gBb7Zd+3JjzlSeDW2KGihOB7BcvL/y1Kx2I6GBIm0svpUrKWj/r7qtHKtjDKK69in83qP2
no0K+NUiQdujdce+5W066di12AWb+NcBlMf64N/vE36f6yIn9VJWT7R8vkUCmscAvugSN5ox/VJN
gCUol42A/mGSo6lCzn7tDAKsAmCtVWpwxLLbYqdGB+lr40tHppDulNeTM4CyMK91DO/VkIOq3TB0
HmR/Kc0awq0u5FoZHvLZRc/yfj9nLZkmN2aiC/Kxtca6RmNgiFi6ruMS/dejd5mACISFrPsxJhgc
U2sfSZppNgL7qNoX1xLO6qqSHoww5/QfteXg3iO28lOCLu515REFJU14L2U2ewpwHGdcJ4cc/Pp7
g4rpkraDRquqcOADUHNT7+x8W7CmpvbzWChQjqJEdG4pMUyu66RE9hNQz35aGFpgGQAhhf56VePg
qEzddLhE9eorfsl7Infx76JE4ldpacBuDFyb5k+tHW0b8p29HUYmjGD6PHew9bk5mW7jZIrqgbOh
abpEPKkR2Qjig7f0HN67yBAa85pyX/kpK2jSzhdPlL/gVV7kWDcP2jrJSQUnkEWBfZW+Jp54Irss
eZoYPv8VTEpxqx0MkkdJQ/rls66jpfLAyT5+AmIkcwjdN7+aJgxY8yTiJz65B2QO6Euo2A1lPe/e
IUErV/GtxEmp0BhmNSSOEl6erRV1MDmRTLhaivg9kEufarLotSUPPFF+HiIdfn1IhQrYf5mqNlDc
JCx5UlHU49DxUEfrmb6xLHRTpVNeCHI1jaRC9Hpa3Q6/BKG2LPQTjCvBOf9QQPZMhfvMJ+0BC/Lq
Quw4N7Ov4Xm57Iyk26fvyqbU1c2sEVWeQXmof30Opynmt9IDuzxHuIpzj3SwMMP4Rx/tX1uLWHrP
JTzG9Usp2hFyfmWNXfH3EMZgxhEut6heQFcWQIBh/D+S4XHNUniAAb2yEHwH5C8wTYlPQf96VSmC
GCKnKPEiqyHJPMzul1jSSJvshuRp3uIQifvfpsyHIgDFtJ0dkOAgyu8lhtJqkwa72iTU23b0BZpQ
M7BG8ONLhcgFUP13l9KB/+wXCFVHH8aH+NyuWRbqVjSHiQf++3EQQfN84006s/VnNyvyPI11Wr12
xsnQLQQ6Ll3waFAbaFapYKfjS81suFlQGRJUrBdghnVgVcsgt+NP1Ot8gbqwvWRvd8EcY38qprSq
zTWzcc1E++BscqotVK839dAy2lhBzEI+jZLbuJux+hxAvj0n/JZMtdWY2Tc8/QeG0GtBUckkB0tI
yPn9Yk41a9J6tni3UvzWDxUjkSw2H5f/6GZTJSwOXPJ1/riGLWOpxhrByYMnZcTK022kf8xtF4Pl
7KadtqaEUrNM9fc9lc/lDVl8CS+n4OYBYWS5IU3cIUqwltp72YoMIAn5YBGv23CZTFDDFIukFsi2
JsXPnr9qQTKSaPRnNAoJK/hEb9Y0ZvgsJcf54TzhUgvC6yJSjkkzrBBBSp3b5Iih+anf+6yQRTU2
+khcSme1V5RwBR3nqLpUPEpDbhfsNAoJqf/WDzhkvMjX+KthDd1ifPqLOzPZEv4AHW4mwQJ1SJ9B
h9dTgxOvzhP1GO+oNwxKw7MHy/KzXLkNAfb9Uep8sxGyWohh1MmJ6uhLjJg7YCIEg3Lf/EhJLJiC
roWutA2GG+UMhBrThNLAZiKLRt5suXYTNmCDKcfMmEQd1MPxzbG1XYRQmXyDnq8ZSSEsjNNW87vp
aHQVLzt4Oeyg6Iw2dhfPoGH/OiKk9AJ7TCPOnTtxZBCxVhwcJhxwv8kPyuOOzFlU84FIB3LeIonf
+ySp9qPe3sQ5GQu1jNLP5x68H6LuXl0a1CREnX8HNDMQdkhN9cea8e+G/fYRPQQNC2Ur8N5gY3qS
Po+TWZ+NxT15AB6n4gtLQYgDt/NqiXrVHkA1VEVIg2p7VjszQ/ZRmXOcEB215qnhjp/Z/y3LTn91
y5EBTkCMzIgwOP5YfSoW1r4hDvw9hbienQ6UudjZKjwg8GiQeMm+Pe+Ndwa7w/rEcocrbVaxYPhz
WEglrrK6VMsRVHqVnnEJN8awWvFd7SDAS9NeY6mcn0TLuCpa+kPSp0Jh3SOaQrhMvohcjFmL3Siz
VjgI0pq+GlCxEKZTkxvOfj7fWXmIlNQ6XWlvgjP+q0jaBHL/gaDNWxl3NKtyUdnmOPfTSsdJWT++
LpW/WAKagxpDY0mgD++vR763kTg7KKhJk/zrCEcqWL3Ia2haj6n04UZhmyhyEmQ6rvhIedzWbedh
HdzP4X5GlpDk3NSV1qSFwSvKmAUBZGhPQNVXT5yimUGGI5FRTzSPGVSvVFJ0Yzz1rRQYCsIKRnlk
hQ/dYk8Xornd1DqwqXG4ERs0anrve84r4yuzpcVm+m6CVNg6nyz1JEEhyFc1kJrE3nrzIsFueUcp
pdzFo/5rKy9qSxLUL6PXoQCOtgEaE3/km6J4vbtLNEVNGF+fCvk1I6+uJ40kfapSNoNBI4YLdbdx
1rkClxDbZ8L3umAIYhyg5j42LbnfODUmlBmi0SDXFP5/jZRCHKm9p7l6SAHESlLPmoYTKgbqgSCU
8vH+5NNvaXqbZ9v+0Zi8Hsi8VbHRHKKRJEKqngTccrCAtMtphFIEVIbzLTc4fbPeokljJUVIecvL
jZzlSGnYmbH5WlK13dk/tlp2Ou+g7Be2wcr7VeY4rCechJtHtuUIfCQGsEfJT9GNo2JNXef8ebX0
3i2ey74NlGfsRFcZVSGO7UERqRkbGSQV4v0oWyD3XNiDlcuudWH1cXkLmqnFpwARE/qitElnUa4c
slo8YzBaXm2m02c/y4SBVNrhp8jyCcpGwFOZBhHeYGiQOulW+2E6/zqGnCOvYk1k+eJwhAPs1JCQ
8mtWhQ7Hgi3nVPWyJ6RBdnHLigS98nWi8rIjkM103SIMPdzUBQ3t7/oFAsvlO/myKEZ9aIRBEeLi
NEwInngnI0KIdPwtwu7GqUe3GwmpJQSBTYOkb+KGo953z7UbO2M00Vzu6j0Zon/D+UbpEvgRwPWI
oQnHrw7BGi3Po4D5ZFJ3mMtTg8RdsnpsIdsD/FTN3tdd3nLO6X7EzkPqpkJVoZPApycSnqMRh5j1
7EpcGYgd/fgj9E7o2D6GIbxpu5dcSX4C3vxQ4E3JBft8FF91bzeCFhLoWNB0d7B/EeglE7hKIFke
WwrlSCvpQexoMKrhnyERlIlMzUXMOpFeRPRq8J6F0kVKbYLZ+jxpXBIHcbLYa1VYovM0V8C/lpWv
o/qxYwEz2wFOWNtySGlW/IpMXjPNwNxZMHSe7J2xo/BHMfo127wuvBQ4yeOVhw69S9LAfCQwS82l
p99PKzAcLwhzcmhzUTTvMZr+L2j3AAPV5/NPCP3K6oIdrmP6fuqkf7R3cmJpEYtxK3kEaofhtNyJ
xPMYvMKr3NOJk7olWT0vLC1SxTp24ZeI5fb03hLUG8JQO8rtKWCx54JXSXRsp6EMawnri0nTe792
Qv4Cxqr8Qrf8JJ7XEhlFQqH8NSDIcMu6AnNMxdx2z2oe/H/IY2Blg5Q7A4RvUlq0H/9R+3FvLkCA
pwPrqtiBQEyRStfmhCXbiJBnVC9tugKWmP/gYD/TiEPv1GY1mBE5FZTjIiTJrK6ply1by019MDmF
84u3Ot5fGzFV4mtob0Xg10FGgXlGYwlJqU2ZkdZJCL5/l3sJgQJ6Su0GQg6ZcediehByTfFWeps5
Cg0IvWQjQTgbhohCOzuUqvjcLR5YONgJAX1ncYWxka1MsXIQHByLo6GyzHWHVwFX5IQlMTc0SKef
KeNYLa7vlu2bAoKu99CLJweM4iwITx9XedrjxMMU+S+kJKP1rGZQOiz0BoIgLja9IYTr5YXeKIuH
+w4uuBgvQ0VuffK+2GYuN4PO5ajARN3tHDb3ZXYxq2JzDW9pXDMMTLNoKoqVrbzWwS/nHd1i1nqV
gh3TQTfVjDLjlvM1OFMl3AETSqxzBHUX1EVMjPmR8pFRxPCoqpg3V0a85hPu4fDCM9es+maXOknl
i4wg2Kp022GR7KsfIiY1penvwG4vwuvKKTiZqY8o0amSixFxZSa47FH2lAzMgH8xdJmZ26LLtWF0
PpxxypJs4B0DPWGSI/+zUSYtP7AaxKYW66WfMxQUn5Us3num8PTACad2QrnNB1radsKggHYOMY7J
JAkuOJxyKBiVEzE4q78bswuWmxW/dQ4tgrir92stbfMNChrtDBycrVkePhFIYrlQqjqUF+Y31MnO
6k+EJYuOgyhfkLuLfOOz11xmNbpGbCgwc2fobbnThsi8DIcwzrBixvymGz6QWb7Azdler51xCPeb
Z3CrbIh9S0CmgTfKm6YwBIlvXHck00bOGCU5DX3Zo/RrLUfwY5giL43UbqLABPrI9mKRY5Rmtgtp
nXFhxlHDic/t9oz9igrPGZkBwbU7OPEfwFaB6d/tMl+xzTbUy0XL6b0h1owi0QNa6rGJx4flfF/Z
IRvmQeRPNXWcNzkezGgD/G81C+hj9ipueCFa6olV37oelJ/v93laZgBr+ZFGxKSYzXKZvXKE3bN7
o1VP7XqEbNpBhdbelbhKYGc1dviVXTt3585fkqDFjtLazfuMrLEOfAh1dXeZOFnl56WFBnPi6g7G
dU1wWy/QM7uZhDOP8plk6vdNzQOlOZ3sZhhX+zL1E5fPESizD4MKvP7KcvdzR0Y+jS1sSecpM39q
UZbMwwiUKcvnY1ShzvOJGktq9xweEaiZ/G4XgidopfcOHcVe8TiJMMuApfT4Z2wYtWVd5quclSA9
crohAfOf17Xs+ktvKbUVYCwAVybdjDpnj0+2NwO36iMjfx6VUgJyVn2HWf6NQoEGKkTOKGi8rTAL
ZHqBNBMZSo7kZtHTikiD/ni5cYkj+s1QopdMc+d11sA/ctHRSTDNJSN+bOMkgyj7Z0HT2J9wwStG
ZQQJlGBKBSw02owWzno38YqGkDVxUWA50W5IVR/QG75reQu5lbps/dUH3fXe+vIv4L2bC/RxnZJz
ukC0ohWrtZzC3wBDCQG9Xza3OvVkKZN6Z9Z26z7B10uwwsxpa+Ey1KOB/5JplB9Eks0w9fry9L2w
UgmyTZiTqXd05o5BuQXpsWJqR0BcYvS11kQXPJjdKYKrateXROJ20zzx4gX8Fgz6zWrlqXyEZ9I/
XKfEKGsiKaP6SozoHfXRF3h3MQmUmAcSCCWQgatacXznLfirUkzdOEHT6dfM+mOYq0CIXJDuhbjF
LS4sx3tjHBBUn/7oqMD9h9Gf4og/lbahuDl4tHAIpI62EDTopG1o83ONfhLr7wnnqYlsFepsCO1A
J9NoaC2NIGhAbAXbeo4bwWUm2RAtFDfUCkuArXb+lJFOH3GNMKFhn11ay+kF8hRX4OPOqTss0E3X
IIRwMSxVdvE3Mj1KFe+dKIq8DApLTnLXzrfRZNKwyfN5hbl4unGrdsCxg98jZcnOuZEcVfbxd23y
gQVlAthIXeXAI+Q3xQ7Ph58RX7qs4C3jxGm8RrBzcROk75bVEz9DNk2mHaUqutltWWpVM7RkYE2h
tnnl+cBcEClWu1QRM6QCAPiGBT745ZRYMX7f+ryyP9julVmmI8Cy8S+64LuSEJL6lUbevXPw9nBC
aqHkts6oKyh6pPpqfL++u/X7vTEu7cvQqOIvsDUXkwB4hfvhBmEzAt/WAIk16VBBrj5v0gA2ntme
bP2JfQx7Zjk2Ej2pXVYlvra5KydGHV8GHSywnWoQgD+b7f8uGbQdzCHCzfpzjcpvvv+Qku3QjjOt
i5vuC6nKIvh+RihdkoWUE6Og06+4d+YmseWKbfMjihhX50+vrRIuWDYzmxcjTAptfnKPTGhe9JH3
yv8LxHh8Hjvci4M8U5ckvpIahUM2bC+Ip/UVZK32nqgorYeJO7u+gOd6pL/kNrn/C1OZ07YoUQQO
ehudpeKO3oRSVxZiaCHdI6QdCutK+bgcE5diepkOMWGxUzeyvHsTYwt/+FpkinjzN1mJ9kMzb+b7
cAxUbRKgv/mEXLrIqZIKJSKqCNJuGNZVRcvOhc7xFXyBausJe1Vuz3zfsSsa79QdD3i8pLAynjZB
Q8nHH3l6Y9zjtOUVbWQjSw4e6IXYJh34jFeyu5IWsELwgYB13xPHUl6U1FFWZCXzUaFMQ0wVEfMD
v8aYITBCOU4uZcrkL8PZmQp28SUUOd3ypc1+8GDTMtsJvEh3lCryOGvJovCM50LMBDFUiB6ErzVx
xrhw28T5qThnrM5D80eOQ4hqcIjs44AmzmpXDAv50sR6KiBxhY4em0SUhgaKrgbhSQWUtBMVntJ/
d/MtGpNWSODDL2z4INy8MFgGR80NPKZ6dklRg/c+JiI7EKyiGCTT3G8mjZ2QHzkBrz3291W2q9Kb
dMHOHYm8a3quCJ0PxyM95mX8nLL7wrcXcf0TJfRSHfjEidTf1G1F/1S9VR9H9Il46q/johQ5VzRn
N1OhMO4esOjk+qx3LHgx9ihv/1WoW0/c/cfxXLtdfihoLNfCq7nBUcQz7swrtuNe7FtppZp1+rpD
fTSq71fMMhrp4RyrFcc4GjexPwN/3G+v6jm8RbraS68P7TJLaf9FJXlrMLiPrbCMFCFoyYPqHodR
HhtkwBp08coNa1TvaBRtscti33Cc0ahI7VXyi/02Y2I2UM15M7latnvXxGyouQheI+lq+DeZSNDw
WY5zSq5Q+sr7rTaSEaXdOhSL9sj3fY5Eng7NM3nrqztlEUL7WoycEYVbjhpxoBsJePQ9XbCJh7Dy
QLifVuz9D327nFHlBsVC/SCLK7wZBrcjZ7+W4G063fwrZbsPDCTordk9W6Cbezfy9763lbhlMWnL
5utwL6mDrFNCQEuThjzfSxPHFDqr1BWVOGaU1dfZBwMtJJvqvSg3psRyxnIxxwrDuDZMqtWf+Rfs
kIr6YJpENXOG5Rx5h8MHPw2n0ANPj9JWH17sis1/yuZwCUfTEaHmXJ4UszFxYYrldmkEyDFQHu//
aj5wLVmDP9FlnXKEYgLZeWU5PArRUQoS5RseKOa3CJM7cCX8RHTglr7p0xt3dnQebLD1nHUWD3jJ
Q8uemfGWbKxb2vkSnAnethDvy2jTxC1MTvjioX2XRPcH5qg9m8WdlibLvDJWlFDuMeuvRGTlccJ5
u7cyPqA0rIm1qVB4HHnWYVOSBSLlYIhwbfM5Q2Or8hIcEOdzUKuD/8A/RnKEcDrivNdhRFoV2BSR
T3t3nO0b+PhuroL4AHEbQ9Dx5e7LuDDua07JtdcKwiV4YTMqEoo/ibN5UqjwM4t7TI9LDvEAaEmD
jgZ7qcHWAxnWaY7dWfBFkdOZSmcdF5oeMeOf1tadf4NYCH+fgyqNqpLbzlRQXo9hBrptDAXHmGpG
3JznyAGsdBjjpiTZspDDr2ElJIk9zATYApxRAsy0xgjDLw36vzOjM/jtk+qjmcKopuwMJa+EGu5n
MozHCkcedbhK5UYkdO1EP69EZ+6xzuRXDhwP4NSvpGBFRzmKEhoBmeDptDswpRuINK9f8iT4WDdR
UHxCOnAEPgFX4AIlp3/y5dHOTrAuMK0rnoAbfWERkHvzREnCoZ9hNBJq84ew2LR2kzCML7qHNqVi
yo1fFzoCsD9AstAx+rH5q9IHzB6++NjxodtI/BnJtqCil29+NYmYeM56O57/sWCkk0a4w2jI+gMY
TSpN+5ijhUJiueGyL6eY1Bdy22ifTmuVDSbBFLIQzC4NZ4wjCXaej4sukZ3C6l6CLVqXplJZbAho
8AMH8vy96r/cUq2OBgu/c8J6ZdMGTl/E0WRT0BjWI/f1OK5FlkChZlSCI5jfFGpKtQEgFaHGGozu
A+Sfsjl+puwG3uWd2qlIKUEnZuK23mI3RsMvMXyH3vJttLXn1g4fuVAJrGoNh0tpF1SKMK8+z+Eg
NOSmB7f4CrtLs7Nlo1sGBX0utKRGU+CXZRB5v+RpezRgosjoVqeLNbIPxFSaJAz7jde0IieMTwlb
C4KdMbDrXd5sFsRtE+KMm6SdLc2iCyAMKPNb3vmnJrj+Qmt0AaPk6UGnbYROZVSk+itodAWehAKC
eDeUqFzbU50P+g+9lp4cMTAbjzY8ISIDVAy0Ks2ElCPj4hSfYZ5WVD2TiUyPhp6pq5xZY7/ktaTv
V4CIwiyOwXALqPVrj92NaxpvtpQX+H1QHyfAYtw8uTqmH7i7C9YP1GlrMiOchR6efbIvRtKLddEh
pc+fH2IPTxmN5Hm1oVZFU7ARQ9OBlcwO5ztB5deEWfW9YgjGlgbGtCYDrk6Gg8Oi3JxG09+Ju8Fr
GyhB39cjUlHI2w+MdBGlhn79r6KpacXC2jMYCZNr+2EuH/p+jXLQ2QgOmtzCw6AQjHecZ3WImMLU
L9qxTRfPqpkkmxBZneAr/RirVCqzLOTR5xwmSONLabkCGOXfBnhMJM4N9HmTSdHv2Z827AeEXM2l
cjuKW4Fjm0PILvGMBe6REFhPkudtUN/CNjvesaSdsDMlQVmxvNKNc7CHnL3siv97pdPgcDuBYM/h
mSKx49D9WRFPeJ/VBOKppXGAbP7f4VTLj5LEPc/wTrgVFpoMnenMIrMjio8ZgDoTchDvoa1my6HE
gprHYGVIzEnIj1wgoNLojRNHL0NSd+VABLYSHUcrnbt3SMCyGW2KJWB2q1d+4+CN3QlcZse0CMae
ou8j/+pMNba6nJ0yzj19S768pUFFqVSaVQ7iH4yPDgGqI9X+WDYF75sG327g9VaAos/apsMxeJkN
fbW1KdTNpsQ2EykQssf9pjbZ41QiMmVrbbqa8ysv5z7ugYoVx/KAMRJ/KI9Bkzxpz9+uWtz5OR08
+BUKY+z2Gk3UuZ0AiLkt1n6OErK/+qiWRD6iOLPJDngZEShCVojr4bgCaR+dQslqXHPhM7au/tR/
G040NPiWJapv/f7bxGEFtiqMNcRWkhkW22AKf8fjPEw8559lbb6s+4Fk8VPbS1gVpAuXAJ0bkUBa
KV2JNaPimVr0pUYjK3FxecjAH/n0hS/HRtlmyLBtQVeozcx8nv4/LVKutwiCLbfYr8m/vdOFJK9Z
mPyGPpf0+0QlFHMskIReGtCqY64/vbGerpuhPNx8YjdyG092cN2Olk8iBA/Uv8wK/N4t0QzA3IM3
FGvLReofmRamOFOlrU38UfxbpZfsVCCBxPzwHcGr5sMIm4BWJgK5ZinIBKTjTdvNH0xR8m/XWg+v
VUl2xiIiq31uqF85wd7p5IuJhDipe7c19WkCY9GlDeI9mhjquJXIPQKuHyuAqk+LkVpN79f/neHv
DjZboGB91YJ/Rcx8ME+LB9hI7SnGZnW7x8elaXb4t5vUwK76gfmuD1EBjE/jxSjSKhRPD5PvRhLZ
dXFEIG8OSf6fZ8w7e0E+Oi7XHSwXT+G9WtmsyS30i253L02cAKSWrm8D3fFEz/zTZz54x9PsJlNj
ozYObzFDY3H9lbuMgX/G+lbkYIt5O2O8yMAWlNvSvDGykLKAXRYcHqHxT9z95+IoE6WsGcSN1gJ1
g9VLp7S35ouGIg/4NM0XrhNkgiZZ27TcEKATscuLHxXcdvUolGVY95k5FT2qx3BFB+hdm2hnYExc
dUYcf/AMAjZNrMcGq06b4c9NRZq+0ShrCqr1h1McbTXlXZrPI01WXvao72wwbfUl6p/JjgeBTewB
Ki3DpT5OuadIT3XHTt4LT7Ly1THDfowAxMqhUmco4v466wV5dO6ZXJ6KlOH0w+bhvnf0MvjseJ5k
9Hl3RHHIW8VbOrJoCQCjM4OQUkzjPug0H5kEGrcapz+J7dPX5q3VT9zXisv6jyiR/e8RzTTa46ng
iC4LdOWmE1Bmy23+rHBIiQ+cIfQZnvjs5yfIjW6eEmqYZ6ZRDC9hJKK4U9NP3f/yMtCzmlwGk8UA
4qwPoLRf09GDEECpieIgvTqmbRK4XuT/AIR9GAqtC0TuNtX58WCXkuPtW082sC+NFZ2YcAWSVyZV
izP0djMJxwn48kpUcW22K2Ep3+sdG3t+cVlivDkG6Cc5YZvJhMNHRppUp1ZfRJf32poqCyq+8e2e
3TOcobN5wZGct78byRUcvvxKpdAgt5U+dE8kpmJ2qD4OIVeKFkF8fpsKX1OSwNBua1w9nou1HKmm
/Kk5QgErHmR64oJf7q/hO0nANaeeFiCzCOoOJCYZ6j7IqEc1ZOwAZ6o3DdjGKlHpuqUmRYWyV1Fk
F+tT8CFXV2qvnaWuPs+e0Hg8hhAo5JrIooE+liMJI1dSjIX96kSq/ytYxSMOdQPdH4+it882BG9e
jwUaXkGSf1cM9D3fHf2C2DKC3JayGw00K/3/wl/geL1Yc67bm2cY+WdGYvNUsE5KiDzoAU5LdhJG
YsJwMCV6tTpuRA/ybWQkEUq+xCEDoRErgZAdP/QGGv3TzdYsLXuflHj8kVqa86grEZYHE50p4XRK
+nzgdIuxIbMqgmBiAAs0gzyMrg6gZXnS6Qky4IFUS6LjsTiKWlK6x5fkxwvKhMQ13TqDeNyweNox
+tG0eqkNH7ZqHdxuSbOEXVcVklx4owS1Zw7DUzzfdhZLjdZijHwgcCeEbhtq05F5xJI2ubAUG9g8
hp0zmhII4HNR6J92KL8JPPnn/85M5Tjq7b69sFLnk1b/bwCOJ9iSLZyCy/+MHkvelCD0kbz9Jtjl
ZDtwyM67JpS1f/gxmYzojpbGSfB+vL2UNQtNSnIaBi8jtjXt2OutzucTgSMlDwmb9JUxdYCKaz1j
AAwkgP/QP1/0Y4xGLZP0svfiT/PDtgwuKl/uK8BG0ZEcwQzwlP3vg+iurpux4pvt8K6DlSrBTZZ/
b8flwOn8FO1SYTK2etmwpt7ZkASU3+k51mZepslznAsNtWrkcwS3RG6mGFZULT/5IHuPrbxIAsX5
DueYnhF9dK7paSC0TL+juVMDWr2GI0OF6Wo0n9w23jmdwXeHLaiqaiDZptjoJgVkFSqA+Ym3jFQD
bVN6bB8M2a291oR0i90YPaMCf38qxKJ+kUjl/LKpJACzRTz/sCmdBuHFvXcgpIGrYl9bnodCAUF5
Hu4cUzHAT2ixRUTlkj96hINaGSDQFv4f6AweJDGg+f4T/uCVGHRRrodvBT1FzR7jG8ra5Vn057ET
Bn0AajSVcuIsGDTBn2je7K8vRsVygcr+dfwQZbYumF/wjG+sMENbdUyFJiUNzW9sXaH0FuHhOJNb
Y3CObdmKN/+HHqS8WZG2qtZogkvb7rKi/piUOWCtRb/iT6m91+co/I5lvuHpItF0kNAaYDJRN0/2
Xu/r1il9A/j03HFHHWtHqcq4rFgX5zR1CATwXC52le0H9YZ53v6JoJDVGC6HS0tFLIrN7Btmm69u
hJk2p+lLrcy3+d5iBVqhDolVyR1QqL3Exm71pegB5mkFM0f6RZdzIk3cF9YfiFrjjaupDpJ6vhIK
77FmXHzMR7w9mjlwqlmx5huHp02dL1r2G4x6C09qEx0ys1I/Jt5yD9iIUjamhIt/Z3x9vHRAtQzN
+jS3EpMRqFjRGDIOVxOur3TmiBpkSiMR1qyZrknHCaMeOXu4Xx7hV7UdsMHjq+veE2amnFVSwQDZ
gdzX+maTWEtPOrBpoY44Dq2qoVN5H+2xClGCZz1AqDM1eW5fB3op/JEeAm3E72CNtOK14r3XW999
9WuFn4I3kXbLf1GME2NHefLJuDUSIiL2xlM0GeQfPUAHRk2FL/2MlCGhXV49F/kMwTENreLf5PII
0boWbcQT+sR5A06m8cZD8SUp4qAAELzKRkxgdRwUBH4UHEVTTAPGYkzssfiB5FF+vj9laL0lAmWH
UaIibfRuoqQVHYQQ+IIwXEuPJpCMWjcUVAYPRr+3J5deHN+4ZEJuNOL134U+sD8nlWQ3wOEOnNp2
jfYXVCkHCrreO51LJ4hyCKyiX+pFy+GnvIRpWzhzRpAFIx9x+z29P0TVLyLhvhJTvVQC5GVQwtJr
eKxK96QU65VeAhxXJNcW1/paw4J2vmf43jCDwKqnNzs5wHA/my12JNlOfJCjfuf8XhuqOB7mghDU
nMA8qXEjJwG3rRl/9lPX6u1Tnh2tqUs9p67+7Lyuw4JE6IQcDKKEjYlR/2xXWOka/e20tp8nj+hf
UXLoKd1h38MqNAFIya1HNfG7yIq8sZG6YWu1ZSh02vaPPn/1hacuJBsoBL1DW4ZICggx9fTADNxs
+A1UpDMSqQP1fERORtdLO+mLIm1OceOyncfJpjr+26kCpFgFNulicdOQ6raZRrvZO1E/BH0yWscp
hJ+MTvLULEipJvHNEPicBP+Auhc5Fb0mHmhrN+MtQXCzxWImBPNMe3nJqKoGOdW/APjVQZ5LzAwB
BBKWE4ILtyJdVRrEiXhSs/BXA0arR9STckK9lyEsZ/pFSKbqW0GCVJj7EiJ04u/641eDLNkaOe/5
UKcpdas8JM//H3I/d/yDCXjhK8lqlhtVrtZ0ZvZJsvMxllRiKCmDjdm7MYDRxJKglUwj/5ko+RrF
G2vMsQWlrAiwml9Qmx4YUK48rjQhr08nfkOKL/orRsQUP3ARzgHQ6l+XOxFmAfZSuDDsKAApg0s6
VrBZQ9858zLzbQVdJo3zL1FtzMAc5VMWkq3IKONgDPoaaIVAzG9EWDR1cJP+L9nWXvk/Wn/UCJfO
oQ5iPeBlvZOR6MfHsYziItkQulxRRIWSIcIhVJm6glCMA7wBbTTl5FVoBUyW/bFPdv1w1Kto6AAD
FeW+36d44FvBV8sG5JVmHH9OkF0x5jveGTZHgmQvHgiESz1+nBtgNKKady/znn1f1yYeJ3Vz8EMf
tJ+jUEs4LOI1OiZ4q6DxOpEGRmaQdfi7TyTc+SEvE/SrEnF9mBgNVigGkvu+gCviSCQ18/Dl4mEW
mxRWhmQJ4mk/WsrjE8mY2CgIt/rWZWNhewXjkLdwjfSNLOsQ0tiKK7CS2DKFp4ct3D6dY3QgfdkX
7uhR/Q5btQwtKONL97waRNwj9uYFKHn7gy844EE66fd2VnmgWCVBoOXgymUi1ScZgWbPQ3qGvGKx
CpTAxJCE7YzlAM+3His7i6hVNjQyIBKUllnAPmNw27+IT92XjV69cElO3M2CKtYiajw6Os17HqQ1
35NXBSoowGl6SE9H/YOyN5hvNv8bRb10mZjJMCQE1eZwPTfv3g73m3W2K4EGVD5osG3r6cwO4fQ7
v8eTh6aLNh4Fr0dsKzKu0wp2EyMkSEYeafuI+SOHb6YgMXOP8ZBwiizVutrqayi6lT91SxRgS8o/
r96YegKmlnGvDasJNVm5TIdtkhXTTJrLIB4lMQE+9ZlJK0e333UJHWjZuBE789xWuvCG8RaCrZe+
UNj/w1bnJ81VPjIAq8jKoIcDPY/umCHpl5cnHooM37f85Tlx57zPwzk+WBz16eA0TZXV0mmRfLTP
6aBJioerjOGet62E9Uf+eoSolSptmTUNF/6CHZkSUiFrYQBMQnSbWhwWGEFFROpjQx4s+utp7h7N
X0m1C6YsMm3uQFTYxqTH4v8oHoREQoneAHefMYfKEXoNX+UBBCORRMWQwJHVSax2tt1+5FWf0EYa
FmhXEQM86gyt0QjtG8eBATSG1OxgDm7XvBhODbIBX/ceFPVTRtvP1Vi8UWBvrs40TD1rbYzw4g6/
GgNrCyZ53evz7ww2C71/AmxzBu88BcD0anO1Lgvjgi0iL5lopV60HqDCkgtBJ5gPG5bhAiQLxjZ3
zi1WtvMDxDboBPuJ2yiLXY+hIVuCQlkoKvMorEyRlM7UhMsPsG1WCnEAaqM6hcRkVJgM3FTDSbY3
JMHJ9t66dWshwlB9hyDnrBwL9hXwAkxxnG3uN7ey7Zkjf7zSUkuFOQXHpTlcHkgjYsqy5LQxBAXq
OlgOSuSC7G8LNMCet/f7J+x1cSbvQpHSFpAuYp3QesY8CehvQHJU2axNv/KGmsVCmd5q1RUpGEpZ
SLtZRo+CPVbaV49ak7ij9nhv/CV/0DXF1mMckV3H779Babh8A96OygKTR47qM8brm5raNBPW3pnI
3B6OJpHqBjR9buXCqoxaCXqiVRzbO8Jzx9tx2YTp4q3tzPCcSk81a68xLKKXIVsV4KKBd01L+IUe
p5Q4n5aFNRVFjg3hXfncLANYJrH1OFaSlUJUCZbcDW8gR0MbEO61suovm+ZL/HX1IcxDhaoXXzSo
4pDwycSB5WLSs9CDDAUsp/xvWG/h9uwSwyRW+OY9/LI0RKP8J5n9gaUDIq5ik10QtkCfqPCyMdDO
ptYztgnNaKxJCfe85rffDwYkdjD4tXpE0hkpaNRXxpS7DFRguUSFfU2IMbCsKlPUeQwKHfJoBjrQ
5ddAJHmfLy5TYWtU9htJf5wJiLACjjC/h4L3G2vOHjHpsNNThk7wlmDILjxN0yBeMoZJoPmFyect
+WeBz51LHx6/Xifxi9bl2Z4C8XPCYj1ofLFvalkyQkGPrFlwxeyiPVgcdvbohmFEWGpi1Hp6h5eF
fg4E58WVOktyyqq+93o8WM44C2DWWkybrm0dyTBBSj9RtrSs4oO7eGOV85nhV0I7PCazfHa/ub66
dyBaO6/RaxAeUyKoS2TTjGT3fCUAfAmUDodG7XVMKPOjFyWG02f7AoZkpDw7FNI0c0bY/pwJId0v
0tL7Tk5goqKbwZDy8Y488N2M/CWCYGz8qpIJQuczsteFZw98GShuilkiRZAHz0OPCe+ZvVC1pjI1
InuTALem6bStN+vRoMmuWAkZzu1UwWKZ1pyXNnApDscIBcexKPYzXDFs+flDBROc300RB0GS08pe
GJrsBQF1Fd/HvYb+bR0XsNTBoXp4AOsFRC310OIExT7YUlmjss/8jdsPdkoAvx5OklK66m91P4xY
Iy28dIvF3bmIeSll5ymdfPAPjHoL15GQTcl9w7JyH/D+iuouB0S60aB4n2utPPFrmmjYoiklWTae
8DibTpeMLJlAUm41lyHsw6ZtozvwhW7NgGcN2C8yIXC7oU6bngTAEzmZ0Gb11Youk/ziJ+pzheN8
f+1GSvX7tRwZcrZZoSM2EkB5GfB2LEdf6Cq4hPRRLZdvOdXJ8s7iYMtmrFiX/kLDWFNGREMgBH7L
81W6Kcm73aYaZqHOcXFJDL2mkvH8mKZ37awF1JGQ+dHTgyaN0rhnSRSokEqRzkZs3WN/dOMAW/0e
FyIbByponxywioVGGJU6Ekg8KLy03uV7fsaERN/m2zdK/ORdX8uH3UfM7ra7pRhr6V5qLG4yZ3PZ
U0aqMhJgZnSrGUhSK7vYQhuCEkQfrLQuhCfkk6vbn27UqtnmktfYZpkSjGNGZFvr+1XU6iTZeLAH
jYMNrICkVefW4kT7T5YtkNL11JWLuDLWWrpGqpZvI1Lpk32xB6+LckyvWO+Q6IjZjePxXJxa9p2o
p0jRSwxYDjEkJcvq1W+G4JXPKvw+LiDW7Nnny6nG2hNiahqe6Qbq0bnb0tB76HksBhh5L6Cv2K+c
VOqorAglE6/Oj2GpEg2nyQA06zgJGXJOkSmLoZIbj7RryYb6fMbKVzdQMeOG4FlDF/F+q+GQuyEF
DH4rUtWI1SNLyiU21LSFICKawK2KHAtAi26FNrJ7mj0CduCQtOOuS9G7/7vE+XqzQm7HaWmlBpvs
pAYRAb1iwdp2I4fm03IDO3GvN3vqoRBnPQ0qyADl1rmOusdgF260QFNIzgNHac4qirohPhBAhTHD
FITr2qRQP8hdEZPNzOEIVNkxDHNqsaWzSrzSjiKZv/ll2UUOCVJvYpstmb4WRgT5h9hR3k1Jfbxl
+PB3YRkO5s9rf4VtP1CqaL0OFPwWCWqfFwicE5u3dGS1Tm+lENhRguZ/lo1v1HWhCtLkhu9YyR9N
jjTKqeZXVRvNrtfdzVTHbpR+CK+0B/wwaHGQI7YpjsD54Uod+AG+boitqxzjXWK/1efDqlA2fg8j
0FMn47fFlRukBtRIiW8p8NuKBXV4sO7/3jjBmzhHWQQL5uqQjlieCE6JaT2sP3Ymft6V+sBI36qu
hThYyENzo7s/KvoRqCiIUu+mnHWgygsTH4VcXjJWGFG/N3hw/DLM7acTLDudIyYaEyWjgk8BzhhB
wJ5ajd5ccVnXL/vGQTToEeHws+mPBKX4G+4ySaS2d80Bph6nK24hQvulL9YS6c33uJohOUCMrWqW
fOSW6qmsVTVRd5fkLJj75jWGcOZdp+M+bnBaJ8fK9n+b9ZJlXggPxA6OBi3LKGq0lHtQYXuKkq/h
RGPhkwuQ1WB6ohSup0OfX4jsidHob6dzNHUiZhDjX+cnkLbvr7uFidji9fvm7Ec2gy6avIlO68Ef
TBp2tqBx/45Ftxx+xiExcaPgYRJ8r9Fm610LFZIu2Pwd/CLWNAzChfw9mJTdpMMqCumIw72E7ggO
ix5G9FBqrSrTnB6zENpB83f0mqgT8zQBlfOTSQDC+f0L99QZ9jvThASn4O32nSVmARG9o+/5yYW5
QDzXawEoVWwroavUCZL/BpLkGhHIb3yX4QDFbanIvb0gQ5UvIKAegoDz5jZG3bTZSYdBRaqqX9UT
BqmqrXGH6Qh6oiHrdZ3gz4fE0YSlwWMHjqFH6EQrvKq1b5HHAMKaxphrVOzfQ2HiZQqVtG946oLg
oMpACXxCY+C3mvgG2jSq+inrcAE7PataEFhhwBUf/erIUAitKA3eGM4y693SAloNbQpuybc0lUxH
JxxWcklONyn6T3YgDEe3tT8ypuL+lpzpM9/fpqAiO4wlsfUNcgHBIrK9t1NXKAW9RqGtbHmRz/z+
dEDztEx+Z3hczFJv3++GMV5Q6ucuBfuajtKk1uWpXrvKR7FX7khV+C10QCb+S02W945wNnpGt9vt
KCO1pAOGC8Xru/mn6kZDNp4VtlP0xc1KekzDEgovlqVN1zn+LCbpJVOyNvAQAmZ6iuCGFv2MoDmh
Bch9efK3dy2frw0ICYLghYghd0C0wxA4erthoZV7f8Xmmct+jUUgVArTvPxB/E8/93/JG4n9EAi5
+jpYN7+z9FPtPT6+ZnOZraaZKDf/MAZ7TXx+CE0TbydNG3GVJ9ZgS2OEX4GpVoWPecndL2lq4crG
Fj2T8vyThK6RZeG4TDwmOndKsbAIV1W8+m8FFF4xg2MGM7zlqN4H2fiQaPMgwUUM9yAT/z8iebWK
jOfEotje81oSW4eLgr8XI0ZKz1WatsnK4MbYJw2iQqIbuO4SD2Wo/S1bXu3k5tnAeBlD0VdNCFk4
onLbh3T+1ltyVkMYYjlLmtOtssqmlBcyfOqnbHX+B8/cHCa6+eA5trV0X3atE0dFCcEMOHacI9Hi
AYtomw4wMOhmb1rvE7GwCNrsSoYI9jBLlcFFKpNXEmkr68ne6ZkLCGKyemiJqR9sdOYilDLcfFAX
jTd5ess67IFx3nlUssIiyVL0VLI1vyVkiz1jQ6gjptexnt2bnIpLb9+byyfZSCvzRT0D0+hOWSOE
lbwEM82f7BE9pe+jYb1G1r6v6EXSYRgyp4qxvuxbArEaqx4R8aBw87hJDiVKA6vqgjR2ZXzjBkXQ
pSYn7j/vX3z/rBpIuwSg+q2p3Wf7gKNAmjpgJxw2OC83F/8xjmGETUQUXnMviup4/Q/penrMVZ81
LMxOhh0VqFz2PT/TijfZfZmb43A6BbbLrszxYebp+ZPC2EDzofFNhtyuXbRbUnOpNqPV4X/CK6mo
vyCxMn0V3k31HI39ZefT1yKuGpXcL11+y1HjsJelfa5z3e/1nOo1LQzqpwkRg1hrwmUAU6v86DuH
VfbCqXgdrxjAtfP+vOarBv8CZ5ayAgglehvtVEwgLzd/B0Pbi+zOLWpOMQY3hK0CRBgvtkKDBrBT
DDj1wlMBVjvjvUMxOMSCOBE1O/nhQeIGrv1WgtNjiT+GETnd/YplOa7ADOH11cxz4UjeDzINKwK9
/adOaraxUbw23GnlunKu9S8TLfadvlbuA8GR9wl/B+GSFflYdW5pebVLoQzrnn/infHxF2uNpWJO
Bs6IVtRI14ayqr9f4c4ZTpC5AQUg5i9YI2XfWf9sZu3+DuvBlyDo9bhqa+bbZtLhOh5zOTbP0CcT
7ixW+Kc2FdG2rsISjfE1zokx+EmwfslSC7t4zk2y5+wOaM4R/BgbF5vlM4kf5zhUQLGqG5bqsneg
35+Qt86ezcepaj80l8hIaARyiLL/mSRj6sJRUOTo/0+W8Hhk9vwAA0F4aUB1kRDWSTkeiwAkbQS/
EsU5wqj1XxKpyCqSojhoodCh/pFpoenyh1yMo2rctatTJ6YZVXs8iTtsh9DkXh5PSvSSpbpTFwuV
sVlXSG4zp9wIlHcz5XhGZTQSKTr+fMIInUnH9vRYxtff2RKRRReFO2P14ZdOcBaK3VtFPpQ3E5Vl
qoFvBln2cUDoFEOl94H5UD6CVn/QCDuu6b6RBReklyCC7AbzjvvJy55F7XGS0VkqmFYPt6gioLdj
i1eknQ5YNCVAI4GU+S8Ddf1JSFBYI2A6AD5eBeY89IFlvqPAJ7R9yDpuRA6AuWAogHVjAKXJSRph
em8yx2o8M9i6Zwh/pOFTWf7Uh1pcFrYnEdJX9yptnakadLJIiYZWy+BOsY7VsQQiZYlxQzPjiXCc
iA/YYCf4qQFDtf9eguhfBUaia7TIBUHTc5qqwnDa3/vQ8LGovnu3OfDmb3KzvmnQQ7vonKNJr1Qn
zawSbDWJjwCjFuTx/gmENhsbg5SNhFxVltR5t09nRhxOJjPjgwIiPlxWS9gbtRu2OVF/NGn7sqxB
0sahqxy0Lw2u19zMeekSJ1xCb++YldN3vHeZGs6A5zIUMhbOs/NNtPHy2s0T1NztvtTaO1+vJ3FX
mvJ3dCek3rIJh42l5I+Bsa3qVjeD0zbdLqNC9VthpdVXwXaWQeWRT5S/tFT5BhsIBq8WSjJPVl6/
aN23GscdMV5VrWUrUrt3r1uV3doeXV1L4940i4Hfev62r5iQHk4Mcv+jVvXSC4VmQumuQJRC4G41
2d2YC5Cvh91EUwNJ92TFYbqqAncX2xDEg+1bGwqlrw3q1aMel2CbpbNm9Fsdz8864QXt9CGEa0ft
N2w1xY4DBB6FVhuydqAvzZsl4KiXkucClnfRO6MIZsaqAmeJjkU3iBwD15R6qtVfkQMVGNusmnzN
qlNBrTUeV5nS73+PoegUJZRTLeImrWQWKlpZdt2IZ0JfpQFco88XpLoUTPM0fZA+TUozPxbrYa7/
S8BIRguUquwPXWWCELu6noCE55wQ0N63107/jRzw7qR8FRqH3F4+H/eq/Eolf6zJ7ZoahqjFcz7l
OkYgNJZNIX/DwgR7mBXXpmhKdlaXfXOpxWmvBtGr660KCPoOC2w14Z5y3ldY8NKtG9+e6lECAiVF
uWYgdswgpUx7iEobycjwu/UEH2gLZcajesrvqc/zzB/qCHgAHzYtHwLfU+SKHdaFoHx6UCzqSPX+
opgGdGckn07ugLsi0BlHhcHQa5E/a3eq0oRfSfb8nmPDTfJIEzNcb5BEJWq2x1FoSdHc3Dkx3DMh
X3meYh+pdB/W7KLLv9dA2tPDtkcC7i1F8yZ8JIQ2Heyw1A60MmJjVnlRrkqLOhNbY3AdzOEmu/eg
ARKgPWOKD6RsO0LiWQppd4MrQGjpdRkCA76fvPpoYLlosbqlggA7ryaHrMF0e/ywHpg9vK9TTD42
lK2lRlf4U8X3ud8leKzt0FzZMgyr+mZWuYYQxUV9x/Esf6xv7MK73JakUF7aKoZP4lXYN7ko04Ec
wdqfSOWmbQew3n7QxdSDEsTG1qbMlClTtvqznc/BqTiVBNj2l83aBi8TcJt3qViBQ0kyP7wpNNvm
FJ46n6xQDa223wCGU0fx6d4yLxmxp0mZnIglu59rVVVAqgG1FtYRudtxTplznHO6pLjM0vPtQftl
7RoDaHxPFUDKD00NzVw/SayoEeuDinFF3xWyxtExIsAzy7bVtg/5pMTBrxS6UqqJS/OmMhNnwTKQ
hmcMtFlMXA5rPvKwGhiavmsv0ZtxRnRXhEN3qrRiIRJEpbRKlQQwzaQcU8sZWr36U+hsrirB3eOx
aifph2QW6QJFm5cnawZqfyEH+Lk4fb32IAj6CXMlS9MHHHW+5C/7CzjsI66qloDthQunYANQ7YDT
Y9vHrTL6EtJkzoGgG9RpphyPOQxXUQc2mO9yJABmSANcUV3Ylifk9eGAS+jzxYOu0lkK65xRs/B1
9U8czR6Ib3QvHzBe6yeb76kopvoInMS6n+s171APDmYtsxK1Krp9OHF/7tCKPoS4+6Q5V/aZykaW
KOT8v02RMyXyQmmC0FdcH4PXhgjUc6ExK8t1euR9e4dL1Sz/yMxpLLNZQR6ggsT+StYvCPIWW8Bv
U/OcqI1jC/tdF2iuRWDUFKbYFa2TdwKgi7KTGr3koQw8BijRqD4PY/ByY4kKfhd5v/h8DVaSzROS
JsBpwENtGIyIirag3kqo3M7qKRwtrDIV5IeA3af9nUAoWNy9RPs9B/EjL86ezMYiZrEdHWW/3jtZ
KiK4KdfUhxn5IwhzpFSxPCJnlCArMgj+gBK5FHPHhS1Nx6h6FepuJlh/hTU1EkH/V8bVYvtXitMw
Bk2eJ9hYWAFL9nUE0P9DQEr6G8bUCK9VSmsuwYELa+kJYInvShnztuc7j8EWyCTTIvM8ZX68cm/R
9jMqKmzSf0bXULPghhT9NhZIGOT2Otj9K2Wn3+n9dUueA35BSJ2r+6ihCAB+BckTq05UUxu/IU/v
63JKPro4ojuklqLjHYBw9dUfdEFa/1R40wFb8UPy+s3QUPxOZYQ1CsZYhi0qzsJGnm0lhSz6Ltnd
eKzbDGQfL9gGdUnuLoVEuD8d3LjxocpeXRz0jXaAefCYL0Iw6FmPDbsBbyKb/ztTUER/uYuE5XEi
nAeXeZjenVJe8uLbuf3vBaklzdcH3NwoDPBWEij/0zXz+6gmV1IUEIgCP0cFrUN0dIsjP/i9nhFB
4tPlzcUN3JlEwiua+H06tcDiBq4Pi8HqlzGMpxXYNCH8BaXRGQ4fQ4E+1UssPvf0Sq5cZhpnRDsb
LKZzKlDnLuwG/KAltzpVH5v3zrxmg6cMy3Bqe6XurOfqhjwSZEWmWWMOY0XSXLVAmlicgsRYKiW1
G47xJGobg6YPkJCa7SSZTqWuN6U/wBOHIjMk7r8j+tFmrRn3kAV0Uf0+R7isr/iEMjNL/9cV8dVC
/LXv4r/KKjm47ZV2LX22oDU1lSRsMh1Pqkufb960YdpuVu+F3FWEsNUeZ/qGP1avvoEH/OJ6/ODT
E9c6mwlelyPbkENHISk18pUYRZzqUWaW5EwgqFq2vonlBxtIUiqE2pwJz7UhHh4Qbu1q7xRZN/bc
3RCAegK87jBqHHEIhG3KjdvD0s+K443T3ZJ9F8n8geoCzOA6Qo6U51SkNGOS2H+YFH4+40ZtOt3U
oIlwwyzDTyOovza8+8kbfcQLd3VAxMNeCfDwQkUEDraN/hjoIgmajrohK/TTOlVBUJ3vdNKp7J03
5ohoZNzypNV6g4VpUyQLLJPLJaQs/YOZlovxtVcpoBOFqJhUNquZj4KQg+Go7hUEvLvYpweiRhJ+
nrMdEaOAxioVdCwylWlmZpL41EJEwboYwD7P0VG0fM+a/iSPmnudq4H74KYl/MgIS+YggP1AFFvT
hNDPqsC2lkUFnCf3Arh8blk/BvdxBOSl23CFTA2L67V/gjF+1MuncA9gtsso2RKY/jK1e65BfHsX
WhesbyfwoJ1Wxpxvd5u7F7aM5CPD3y79eI+lFiCJmN/FeIr/B5nzNT2xz5s7RlHwy8IF/X44WynW
U4uVkl1li4FbHyGK4JvRS1sSgkxVXr8nGg51HGQ3Dv3ifdZmqda5coSSua61HMRfQ3ioyF+kuKEz
C3eYXUvISR9tRryBrjp82+BLaaPF4sIinhnVYPiAO8DMMyRkPtz14kVGRTP7SHS9oEpy9o8bhk7z
MIsmqVuL/ozjrPhGtRAyNBsKJy0jtSn3BDHDvK9DSDOywHxHbJ1FiV3jCfvUVRq726JNHrh9xGKR
XV4xI4hv85sBR9erhUCC8an/00szs8TNIqQTQ4rKe1YePUoOcj0/xG9uLSNj2iT7WzRjkc+tDtxp
uRW13llsp8lG9iOhgl2Wu53Q/Kye8sZd4cKv8WXpRmj7LvWuV7pg1Jr8wbyarkPjaOyqK2OB26NM
5NJDifXFuGDhajdxGZAM9B0xVc/MPm6GfTML6YKiv6JAM9co42eoYvpCQR+thS9ZqDkNHBiKiyWf
94pCPkjl0UZCyisOiSjBVJ/1R6GLIp1R4k8fWTQHJiUI3bb/I17/+K8yya3XIJ14DSLAKxFQJuXp
10pfL9uUkkrvnnCmDMNjMAgYErfyhUemYLtlbUve7J38U7T+Jse/fKObvLl0b+SP7X3SuyaCvMqE
2Ewx085egnwlAbW7COQPvQSfww0G+AOpM9Hop6RxJxvEJ46VHw6jA0BuAyyqmSSo1hoTQpp4NZ+F
GBtdM8ZFMF4spzJOygeU25ZejNsw7pCVPIaJVlFOF/Ft92tJd7RvDxZoHbpL2YkDfbQAixbVpvJr
6dIEWAcg6ON9unbBerOdegWmeVw6nOJlgfuBN2+0N8nXr/3CKMIiOf1u/UozZHgXAFpNPmhLdBWk
YQu4fKQCdzgIvKnlL+SSvqnYZi4eReWjwZ0eFXNLVhLRbqvy4hl0D3jtAH2iuoAa6XM1fcCjfNBg
DO+2Roj3WDY+2/CTNF+G9gScwuUBIhOHpRAvJYWnSbsyrF78/SFCSE0JWeriWuC92/Tv1FEpEfRU
LncrPzF2gYAY/uwW1Ny92UPdDBvK/91J0b8qYnSF6x7qmOZ+7cCIT5Vm35/t9W9kyPGdFSND1ZPc
h1+j2Lg8m6L7sLUmaUkjYyo2qhXZ7GcYFEOjKd4OjScuh55d+VbHr1r4w7i1rCdbc8mG5wIPo+zC
gL622/+2GZHx9vp+kFpquXdtb8Svv9vLkBRFsOlsbSyzhD5Lf1hpAzPoSBXgVxK5KMFQCWRKwDqj
1Y67fMgCWZXro18Hu1z5+2anVInrwR+bAwl6gm1PK/PZ5g0zjSP+GgfbKCPAA+WkyDVUCT1LzDWY
LMWkAEcAnxjCNtmF/AcyJKujIzh+hE8nPJpKB+SOfoN/9S5KytBkG9yQB1+pRzKK7kQLZtqDoaYY
LGwpaNWYZVD1eDV3wwZwp9P3pJ7mgGfJjGplP+GrPh0B73sLy8Pc/bNF9VOXlZlbcPGz63QRcQ7i
T9+d2tv9kLdwb3eP2c92LPQaAfvHnUBAOdDQJ2rnBXl0cFY1KoscUTnnJBy7PBCc5ZEe7YGF4SuH
exc3gzNPsp4+XLisUpj+RIulTqvARbTd6iUr+k5LAyAOgY1/nMXPQ8LIqROBT3yjBXHR6ihYtMKo
YMIAJBPdOxEqMMmdXNfX4E/8QQfkMkspAIzfuAo+M24x5ljmJ10AwDaWmZx6VQQm/dr9snbp8V1p
VoSz9ZRVr1w0k5p/fpFKMXmHweG0QzVG/YgvO1S4tlkAAvRyk9ujQsynTDMxmXNe092qg163BalV
Lw0LnOZTHlO+TecbkuYrJyGC1ysLeX8tTyGMypz6f5I3nRvfqBtHmaUqR/4zOOx0uCG6LFTz/7Hf
BVRKj1kFsZ95bukFT1N7lBlxJU2eTrGUUD22eFJHqGicZlDjALOefpwNQq9UpyoOzlhUupt6EdWe
9lV7BnHk3o+Fbpm9fUSKUakosiqAhtHcYxpJzDsR2ZO4Frp09yYZu7j34XAnYqHp4F+kbtmGrzLS
GMZn51weC7Ag0cTe19DzQRMzkpqHA3Qio6pH/NlkQuY7TkU2hdSj11MJZ7EM/2IGZq55o791nnFD
PqA15Nia9aqZKHmqgTOIj2J9xv4KjSGPGEPNiZOiMaOGPV2BunThMQQVqwslFKaG5ftPkxZqvh82
KFOvfxXXfzdkHWKSoedEjRfnW9K8FqZTu1TdDDcw9zTjNMBMkfKBjtNU3ppJO3i02CC7Rn8sQ0Mt
a64k0rjnxg7k3nfg7vq/gkYQRodOvsRr/zZhNhMzIddyZvjdcVyeli1ilcX/OFGh2++OjM3RfNub
o38Af+dzjcaU86jRJMOKTehDuzAduwMVbgNMyisFHbVZGJQQkJk+h5s340OuDGq/71Syn2a9tjF9
ddw/3HUimKfA8/WfifvBA7Bjmtp7xcjLKMD6HI6HEBR/G6L7UhHDpG7v4sILbbsXX5uUuU4Pokn2
LDCEYxY0N/Nlrdi9kf6+d1ClJ3Br8Ua/ZD3miRKj6RjSopAFPv78l2qVsOwmT4gqk5SAlGZC+o6q
/6D9w5UbGPtIRkq+f/2xEt0/loswYuF64L5WJq7gDQPphddX9aua8nPTAHp5xiKCp2kDFPh128xW
FapzCwlPID8sqBefrGMSaVMtX8kdrbboTijmDLWy1FNXZl+sFTvVvWTZ9yk+n/fVy65Fc/ge9d25
riBCA3YLZlKZGHScLpZfhsz1FyE9gExhAG/qLlKl/1kCUFop39ncJnnz9ItJFEZDE4JorjgSlDIO
ayfzbVOgvBV/TYazGQOIm1DchCD9yqaBx/dJT1H17FQ9gwiAGo9cweJk+2hPK98+Azyhp20mRmJT
6b98xDmZYem1F4osJe1vKpFAZwtTcuHmjAcEbgwthiaUWivfvjr/kefJ68M7yosvto+R+8aJV/dp
CbESUDv1rHAzEjbMDTI/6bdUkketxajD6Di50R276Q83B26DVmjU3vRAXI6X70f7FjUAAiMhzrnp
q6o7VhFgrPiHyF6YfRgpa+dTWporVvrbBzqcQEzdBY/aX1lpuNP9qbqfmZ0qGdhlneraXu5BusJc
IXA1fdjwLq9wWYfDd9b17kvDII2B9LJirtRP2xF+1LZGIeHlxdyy/1atOcMW8JmrVPc4mW4n9ZSE
nrk7r9lqz2OU30PyHDA7fZNdlmkye7oq3+f7xSLK1LvOqlfCLXOnqdESFDd73mtkBPfj5YLtgwsd
jSz3RL60ZakesrjAQbsm6g2VSItKZDRxwa44Q7eA/3C06qH58qrciYjAh5fF4Uu9uIYoMe5uT1dX
H6/KSIJQOEwnIIH7ntCwdNFJxefrqIbovQ/0h4zLdR0jDa4hOLf1TRPTGBhZ/9OMvLA44w44LJXN
GHlchgjHuwOW5TOI4zctRkA8Th9hZGEqtlpAfcgsgq1gzcUwkB3iQva64FWWjGdVoFg8r3BRbMPi
h/KhSa64yol4ZUJej32cjGvvb6K7LGCHf1fMOxnmIV6Jjtw2AZHCJbIYf8OYTAuLcHfBxGN+DExt
hGksfwL5CDd2fO428AzK0bFR/bJw0w5IAUf31gAOi+D3PXJpCNL0Q8XZGMwAfb0I+fEXobp9fpXs
DkjTSwdggVkue8HcW/79J8Q+JdwujKLjyBlnd5i0F6pNmXaXNb21I1anQB3FOE8m2nGHj1O72qzJ
PKeYhX1Y0IS6yxYXpoJE8VJe/iWtAvu9Nxf/512XRJb3mtAHJfe8qQyZyDewJ05KD7xOBGXkiBlR
hrckM0GsmMXU5M391TmYoIsWhHqCA66eSW/XNoKS2RsL29TjGCr65lYFNEb/4rakximWy3sXxd39
0IuseY615uhFCzCWaqmA8pvu8kqGrxXdjp6n379o6W6ruw4MwAg5hEfwJ1FiVtXLP+NmiLfHS6SA
FObgeUaZpOPSHcdNOHaA7+qQrs1merqEUriLqvZgtEnrVJmWA7hpvjlgLKKX4tks4u3ZVDk4+qUB
wQlusN7qfve8Xj4fei+8HuObIXPi/WChQKM5GQibNyxHmlJTUwsHt4sMv/s8mGmMEUMuLRHQSYkC
5yqIZ2iFH5kN6x0AXOp8T/lWvhMrnmR/ovXFm1QgTwqAwWSS0tLB2N8UGKSDLXQwn6L7QDa/ABAt
33G9+6x2G3/s3QSKSwG1Vk6tFpOX8dPl7nYt9/Cxb5vlUrVTvzxJd5qcFB1pNfLI39jzGRmEdW8P
lr7vPiAIU/tR56fa532gKdHNaRo8SxjOYW7lzq6f0GL3ZseCHRM13OHS4NVEmXB7LoMatDuPiHEd
2+MTpa7tLBo9IlqBQOeJB+sLtwnUagSXS+B0SPnnVynUAAm2h7YPzWlIDj0ft/paKf3wUkjMTye8
9wZTeZ45t/flVGQhSKcDwaTpUO80yxW3RbC+EWO0bqwpVRtlg3aRusf9eJHjd20ierFHycQJYwg+
UnPBZByvClJIO80e8NdIIedCAVtn3pFCt6WISfpo0oKgbbrZGxgaByPPStR1LOjeeGdoTmznah4R
wfptjFR4LEL4D5bmtvR1k4CctVNQR4No4oRxusQbJlkDJyfmg7jHyHpdu+V4FctWiVbfcGwSE8Qf
oopOZK68tjKKbToiBlxbFYDu0TacEK9qTFz+KRypqIwLElEHij9G23cqSbrliuc4qeLGSrqTMqtg
tynXJ2raQX39NQ3K4RNDFvKAHE/7MXSuM0rLhi13PAI5Wn/FtBMg5tbLRGDt88yZrbK2vRWCB40i
6EYIbeNz9JNrSkTEg8UdKSrkdQdISOGJzr+qRJObH33NFRqmzLquneY+Zg+ZV0/Uhs6fYSo93AVU
z61K6TkE862ZG+kX1g0V9FH5qVZs8s2YH4ps2HCVIWUiCG/9opW5cGBTffZBtJ3k3EES2Bnv2yOK
lXQnWoy2ZhSZFXEkeF3YpwfYWbteRGd7MUsdFJAEtqncaj0cY3mzxtVoBqYOPIkO92OiUfW7AEPJ
b4RNYhXfYOn5JE1IlAWllvIfBGjKCnJEb4vPQFau5BViaV9AgssbnmS8POkkFRqWHZGJ482QeJHU
aLXXP+kmoDn0IjQle0C6EkxAttGZTYR8SyWA48FVEb1gghMAoLkCfRgl1GI34OKG4F6OBVyo5/S0
Y4PpuBZRiVZzvAxIc9NXqoFLp0JlB55bxPmDOU21v58jMjLrYP6SDxGq4YuqpGMbtx0u5mi7mnNW
rMXj6EymRXoxjetsz4ImigqeRS3vjN31F/qOeo/UmLIlEGz4qPeWon6wKmB0kcYMmVF7155vM0ov
EzwgC9xqbyZEMTBMyqi1Gk2DAzkmTRlnjuHS0qg8hA7q73G99m5C5D4tz6IQ4yGsBYcdT5hIXzbz
xRfpGeVT0Hr3gWgVkCcYbf5/0AcK03pw484VwE8CloP1g7KkrPhEkhovWE1rYxKpVOylvT8D0cvq
nGIZhFhVJjgEBmM1XZuloz2OND72kCl5tk3I9gasfsodwdGd6Pxo2G1vXXYc96kslTOfmgoUHG8O
7Hb2qpbDtoGSqyWStstsqkUWrnI+fPpFsi6oVTYppvI3/9iXsrJeV/lyi2y8bBnnTP9Gc4WnCw5b
dOQPVn8fiGzaAHPAdJv5xdTTOPQUHvb6DueaAJ1Irt34EGmzoKKIVwDU9jalfYlYKn0+wZAEryAo
ZopDvPMbcQC5ovZQIv4tPgcjLXggLlB919Axq7Jyi31XGwzjDUO8gblCO/eILdB8UY81Om9Fje+U
Bh0QH1cLnSZZG5JO3bvC2Vau7IKwHUFgp4f8ZByO7mzGdP4WVOfJHYuXARfvfT/kCq7AgdG+Ry1y
dsqxGhdi8w5tezeM+ty7/t15vn+Q9PWY0c4Vsxp01+K9COkC3gBdVrSL/oVZQ7iP9RAB8WFvEA5q
ZPrE1JO3NZk1zCwaNYRWvO+L6t4zYIBGLixP3J+qRKwhFpvVGlFxHHz3mBFHBMTrrYVEzG+MIFFY
P7iqxlBhfoD49XdMC6Ow3ah26SKLTPu3t26VV01yB2pBfwLR+P7Xk94KyIAqlgbUrxOduWxITXsF
TP36Dwvmi5PF4HiWjbiBJ074Jwc3YfDw/WMinB1VXts23YMiud6nZtf45NbiJsj7nNbzQh7L9s8j
j/y+KUVIrewdhan/C2Y/9yQIAO7iANzb+Y1s9GSTcOJGcIm9rj82RF6Pi/4B5r3l+9pkXlFvSIDK
ZbiUddN211zLXGr/OHlAiJAnSuhgADK08DK4aLAcQHyy2iQQyY1Ksg3da3jjysb0layCAfR+k8ON
0kw46xz5yz6rcUbpJiY4uSauUfOEgAAh7TDCLkErl7dRoAzHA2+ceY/3E8ExPY1rfcLUriLl2sGz
S7tkc3+rgsv48D8S1tVkK/W4BNRZogWazUUNERcd+HXDUmBvHFLaYFNY8sA+k5Z5Mu1iDGH9r3jV
rBwmCwl/pBXPWZ2HZTRhRPHFrMOqVdKjZWx8e7L8kU3mrtRb2NWgN21rLzbgkgKDHxqQALSpICbL
HFuc4hT7W6vqplFGf7qYHSFls2djyB/p6gogStVHtyC6ZPboseAu3LuLrl254DQZWExK6EUUK3Lq
8yP/RATEr+37WgP/WGK3JKahSdVGjKcFBudixbKgle5Mlg7O9roSC9whZbcdSz/TqW/tCB6wL/v3
+7e4etdlbSwDmOEVmGY/I+Uaiih6Dv5ZjCdJR/PFqQt7vvBU0SHljXQgbjgTj35mbu63OFxW3J6g
OQv43dbJikEwDdyFRoB8QTul043vFyB509D6PkiQwYpj97CujLyz7TnpWtwhj/gLto01A4ILb6uw
iBGnPtm0tkRsjyTbaG8TYRyIO6vCgGGhr91sM2p9SqcP/NXgUsJRQLaqK7o7lZYE0/58cpA1iNJM
DUCjLM4/qlAA+iN620uIJsQR9CmmrWABeRgzvisviDgOV23dURGskWiTh7IZ9/Re/7ZxGtQw/CEo
APaTV/GryMMeX5+6FlSIf3xfmvZ34BWl3a2Kbn89m4LGBBQABusKadYkPCi74F/YGo4QSSLdffgx
3SP8HdinvxYUyBFAWH4OU4LW6nIhtyUSTYlRf3gfwBbjW7JQnevSGHgRmg/LLTvQTF7XwTRBaVXU
aktnYKIJ4tNwFJCYUCw9JLGW45MZ5dQZEP5yeJXrdKR4AadKS6Ki/zTc9EtoJTNZE/jKgJvDN5sI
82qktiQBQpuTNgTKVgXylza58+H9Q7qijtjBli2vQoTZP1FAcmtMCH3Mzws/hdU5mFu8XsT4WQDv
90AR/+mLu3H4AVP635UAcNQsE45yvKz1vPQa7ytXa4fjzD/zmiGPK0sxT3eVhkMXzUG9YjoL6pnS
8LwuCy2YtL8u4K/gFq5EL8vKHfZlj0b8eZVX1gC78UfMk3eqdpoirOr5B5WeADDydlfRVXhYCgds
BQIVAnhA0c8UzmQEs8U/I/6hwoHo1bfbzpcmsUwXv5G0sq71mr7O7yh2ugDpQ26Dp1ojknZbA0rc
k+GPoo4S/WbKEGrcIYBqisEccHRcvztTOYzYFgjs15dIIRoAhlIJxg1I96fhb9oXNx7WpG5A4TOK
n0xcqJDSy8T2VF8zQm7VXg1c6tffK0EZ0Av9kKiI0AzErei5HC69CxhXnt8HYimF/EDafHahfnqS
tsVLnAVoPU//AmuP5OYChw9StWRu4KYeLJeCTE3GkPtrYWm3Nv3yFKibzdsJXjjr+Dznec9z+uMr
Mr2kIkbgYhT9X9IBSeOR1jjj7vqM0pH4ZqyBAvPHMjsF2N76u/M0jo9RhvLHhUrjcggmfC4+Ok5N
TU0NJXuXCXueNwrS6cQsG1tZCUO7qmu9i65wsrkfnxbChXjS3kEdqClRc5g5ujouIq05RzQkzn4I
NvDMfujKX9Gldeh6lhoLyle1JhHO1eLOaOLXfRur1FqaF9XMjNvGX3NDUXzskUj+Brh6J9iRF3EZ
Mat+lh54SE3kRHEU5A31zqsmv4plvYDl3wl1LVlnLHKBNROmm6B0/WGjEpXKddmODGug6STpNFXQ
hNPPcvZtwZ8m+Q9THTXRMoQPIfd1Ca7MI5rMMAujFu0q4ZrBnmDiSjh9+K+DAmwcMtguScbn/dPJ
8Xcg1g6DNPL1Q2TXROES55LBeTdOBpPOfK6v8x9QkrJAgRVqw1saUm0C72eP+V7N+oxehUBGyftf
jJyJPoMPjqoPZK/f5HcOJWRXQDesAQNO7i0syl9CyvEzlg3719ociu8FyWcW9k652cZFyymyFUZZ
rzydobg9JSQzDZpPoLiWh4Xz/BSxROxZHAmh2AkDCDfyWr3FTFPQAE2skO9iaa3b/04ylq+qIMHt
+cM919wlLVICaOFta9kZkJvqrKA2e93ftQXF/IcNsFwqXtrKlzzbQ7xNQV5/8sXyqCyVPS5BI0ZF
1M0ia2pkKMj0hC39buuQQ7oXdUQW7/s+oP2E1/xb25F5xnYFGJrgnO2ZVJ+4Ks8vnpqpw2Kx2OcG
4+08i0JJezhEGAj+To63e7ABfwgrTIO96GaMlz2KrxSDW08yo9W6F39ResgUOOSFYsA9Wqc3j1oN
EA+kMO890ETClWMBqyHPMtMs3rWU8n+Vz/wpZJsVhPRdXNe1X9YoqnldBObwZihNZ/dnviG1drUX
8oqezVOprR9Lu7KhEiTnY8QFzPxmDxM2eRlmGqLPjLjrPlFu04c1vkEvZIR9WFLhpnPeLD6gdIo2
aBRSXP1moQlcbg/QJZGivZKf95jGzQRIGxeauEXL16RuCMvWQGGx9g76Nh8foTY+YYxz4JOilCqW
7WbvWi27BeZ4j9GatAbWyZDb4CVNFLpAHy0y0ggKILY56d45KfykyOJqWGTI1Q8p84ij0TslxQjX
jNZ/tqTD2uiQTGxW+3HfsWTsJ3AZ4FRHztJPzf5ngQNGtYZ1FqjK9ltqdKBkcQ176VHemTs/Lc5F
yI7cZQW93fPF5PEdmTaV4LlvWhfXxUWi9ga/JpHAlzFSOvlRfhOc3cwCqHhR/F0TKs7/8IA7eSnS
nGNTmvNnqF+hAH0mS060QeXROW233l43w6YWra9pbSsI7aXqOS7esw2C8cIsvRvQRf0sobITTKVf
siYeAw1LzKDc/0QHqzzcEO/ZJKqNX0W7cCbfi9a1lEeIMiWFsIhCM+XhcXXHche4oQcyWR55ZebE
WiIQaEDMDtc2qXKCMKXoobGiBNwNmjmPo14CHeqfiGFxN4zUPohRaZ2NTCDTia8Ce38xEMl2DOvb
dIPt0Dpzt2rt8bML/DA3rA42qyu4NQHftWcCdfbei463XqUlWH9g8+mVRJejMz6I9TZ8cSimbEVN
jzOCu1Bvldrg6lhtwYxA+I8pBhpQpmaUqtoGXRNeejMu8YF2ELtBfpypOcwCF+hFfjru/VfQ5rLO
dtFnkXrQqPWXbUnTH+YXcZqkEYhrYNppL47+TZVmOEN2Phq479AYgOEI8HZweGcxgtpyJMqL74Mb
MXQm4jyrVjJQFu4AWPtgfJE/zvh/TxkheqZyQRe53Z41ZIsMer7XUXUlcaCTi5gMGaeTXJO1B89d
CyXvvbysn91Das1KBsWvs62Oz+mLjs9ZwifuSt+t124uKIwPNn/BjFG0ZPRAJgRF+PiodxzFkPXU
lXJNqrK332ZOQlMMxJMmJKsoly5HKjDJSQY/SweuAyu0Bh2ivDLDsgB5SUUU1iJNzqEptWhngGKP
1YAHACxF0HN0fnTsyYxQ/fk4RooO1d2Y8LpNIeRrTHiYJLWUQprirKZ5IecfNz8+4uzvNl3YRyvj
iCnlYQHmHKRnbUtHOqWCCwZo8CK/jRwhxhkbXSuJWk8PBrQ6326C94xt+KWVoRAeGjn9qu2muA+2
/EGYVz+YmZZbTBBgIyb+PiHg8e4YLMtoHIF/+iahN+rMbppqb06Va7yIRLSyihyWcFWV/1yTtgpM
RNyXS6bANFEEXiuhchalnceqcFUUhrW+G9ga/nlcU879zoSeCeUd8TQYrK8OxeDPFAOvYzaASzsI
GiYpJo8fHncnj+QBKhYl6T5pijink+cwO1v/Uen2pjySu+4JZY8G9BWG588GvtEh3TlC5/nfP/kw
uwscWNPwkV7sreS6ijeHPfbFyN9Hj5R4YpAUvL+qHdj/YQRpJMul6jaakqCSxAnI/3xHDGscaLiG
9u3ZLthOIY9taUux3tfWG1NeSs657MdH6M0eX8M088ZA1n9u5gyXuz011YujelzqAdn9cwJL215y
L793NLPBadRC9DgHqWQnoa0+2eeye1n1spHiXtBzaPilYeebadjNl4b9RP9e7B3Z0ecx9IVsdT7n
JgeiNDKVcriYxvuhx/2xhJhzloyB4mHFGeDZTT0dECw0ZuLOJP4jW1A3zP4rI//oYp7hBqwm/gum
nKpbFK4nqx7+sUjk+YnEXVRdrfzEJyzM114ehNt5CuiwwmyiUu/f6wDZGh1XhDSBhcApN7UjeHTr
ydr3RCOPGfdcjQ0Z+SzKyGr1LNKU7302LQVQWiNdQO6UP+7KbuNMa4aZbL2TQsGi58JNDL+24sXD
iXDY+9gc5hm3MprIjNYisJwRXH5LW/XeLd98dA4/kCnltGfp3X3qYluZO4SBCHLie7Kg5HT6+Fk7
qP3I6uYhhvvYG5L/QyBoTzJefMteEmE6NVQw2dkD6YIO5YE7IDzMSYv3PmEAA0PN9BXYout6/WJ1
dswSsAA9w2j+KzPWZfAskZekJuH71D8Lnx6rLkaCw7QW26qEPrzPclj61BzSyvr8ahZM/4jgXq7l
3Ao5i2BKGE2TIuWzgMK4aMlTd0S9kA9+LT+KALIfl6iUvap05oUD6yEelKCGfFVUwYRziMZKNhyp
knvIxwETN3wtSsfIipvG1XzaCy57rfMi7/cP3q0/xa7ARXex7CliO2I8Vu8J3/g430MKRiPgWgwC
gRqaebOajV7FuCxQO831c5TEPeQId5cFKzEd8s9UoBNrrTQE/F9k2pNVu3cVstpOb2ADLx3cuhlf
IkgZQCGlSdKZgtZgdyVt0Z6ryVDPrDIFZgj6rb8QheZdIjD16hH8nhHf16Ay07Lvw1YfwugBc8UT
LXxQLBmH3y8z13ACKHkCGllAhYTxBzwS0vDPhEKF87fdxwL/6xZ4w6ZOUHYHkn1/VLN9C7NZ83hn
HM0LaV/uvT4BLRb7zTm0bxFfbPpecMA8wiTuddE6uspOrKjS5q6dArgaPKJd7ySBmuLztzUVVy+Q
269KBZKWZhuOioZOv3+BMpf5S8DCpYc23FqZwSnrCSYpzV31YriqtK2pl9BbNRfc3OSj6r7i0bSh
eXmRjGchmGR69XxFB8drKd9JD+H2bIE+acEG1/ZBWoI5xqAdDdsrA9tqb6zm5A/laWW2GKzGSnJY
N1D6fzhErmpO+4/sf5+aoO4LstCORHNdd0Z/agsRbTYFjtqNxTN9xmDSNTwEl6hNa1zyn3McVPgl
6CRlfnGp/lEhw5AghwFKV63WpcClmzGKhBFLjv+eEYjyY4ydWcWzv4iQMMhln4YjrO/sCpyDCvki
tg/XhznaFh4ZMTJymtNUDL5s2dyxATIKN3qbb8Zf0JWH434fmYHxF1G8Hfs8ZCGjvY/hZHzLSH52
S2RDNA3AYwW0qInpv3cXWdY27t52mhzPZ/OWx7Iu0lhOzzWIMAbaf5BYYEUR4uLy9jU/+aq/lQ5D
tJ7vw7Ly3hcg2Saoz+3c2SccQFIOHC0aMotxhieoVQ7uBSNxqHZWeCItidpbYZ6kJG3ibsiqWzOm
ViVbXzzVfrrCZOQflnpRx+HHmZqzeymoIdI2CVymEDV32RXTkwFMC0Xw3t54auwg0Y+enGgfRlgM
azZB3dgVuBoYmGNkeFgK0fJFwFmsuTQfD/5Z43kDpW5HtEipfnWQggjBjciq40R1i0KhyH4yYD+E
5KCpUkGNtnLrG/5UZSjKXkfKPOWSFRtGS2BCRPb99IlcGjJlli5kovCA6EqOG+BlJ9MyVJ22tEta
diYZmKkRjycgGdSD/W07bLRpwZYQwKqD0JtsmDZdeDhJW5AnqxgyYjA2F88CLNlwyZ9/WCjc727h
2Egb2DRBbqCCB2OxiGhAa60MxxlmbF+aN1VMRLh7OtE66WkSgSJ1vGJGytTpXpZDHYR0pIs39XAL
oB61hBFC+R7KSzLkers/JG8lglZjljtoMm4UquBTMAnFVcDcNHkO3LNAyjvgPUqpKUVHtYKFHPFz
ezGuVERAqEn6iWDD5RrrnudKJg6EkP4iJ9HeduoxvCJvr6BgqSSUDw1c+bmfPvxRc/Skj+aWyUc2
+KL1Jad2PLvD6cyeg7qDRda/m9DWO3V1qaAsX0kXFeQ2JZIqWdapfEkdmFlhx/0GzmgWIxWZYNN1
RkEYMcLtPsfhwfwv1q4tm4s2m/CgRYekwROZYjjHBUekBwM+3W6QtIL1F4NcayE/Kr0bYf6k7GkI
7iGxxj7mCjIfo2BACh5HopmL6c9eQ5wI5xTQHLIdOOE7pdJB8O/ygM7NFC8hJymqyIgPxHOh7cLW
MTwjHCXlbtR78FP0rlI8f9dgI3DjtRymb6kOPfJjfzYxTyR2DsqZGnicl5uyKDzOZhgLTNlPnXLg
3XGtDWtO6VYokbAof90c7E/GefzOdcMewfQKIlOUuQDj/mH/M7Yp+cteG1UKfOwMu3m/cGp2f6FF
LDztqGc/F5DqIaa4zx+442NtVx1wfNV31nGMYKNcna/7DwPLJ6HWgEtAnoD85bHJCdtD4AeH18uv
nrIaf5tFt9+hTHEdMHt/iVszic+vWJ3U281Knzx5aRwe92YXS16Cgn4olS4bQ7yI51hNVQrcothO
Hm8Q795r24o59loOevx3trlVkK255uqhwRExtyidv5FTT9+gz34HlaqOfrvfv/9kZI6Ze5y3pvVQ
jgHlB8Eux7uyBHnPbafL6vY77l26VSZ9CyptRHR2SVP2BrY12y2troiMprC1N/dKRGeZD2FMVx64
dlPOAuevEYfpmojNTYZW+5JKwhvazMfSoYbV+GtN7GIy+sD5xWFYEGUiV47+vqmDoHMKYklMf0mq
05ZyrllgwqF2tb2Pd7wHirKf8LEhA7lN9ptRldQKmG1Y/oQ2gkwk4Z6MrRKA8TdvvwZfMET75Zeq
niCbWC2Cv64/3EVIZ0qOE9+HcQAbKxc60I+alWtBZukRXUYVXRZMQsjCFDd/fSockX5BYwPHkb4Z
N3okgozdVC5mqYosrRatqEosjqEwlyufHTDHtlELPd42fSN7pdEzVXuzJ0+XJbJnHR3BmYT2jh7U
09G4uvi4MyGGWwJqg353l8B/6mJguq8+Ov3m9RvKZfUAAL2CO4g4oaxvmb2y5gftq80aiuy8MwM/
0H10L77E3Qq8kHrAkoLQvH4h1SIhQ2iIQrMQGAeWw6/YpKj6tsFlZTks3VBdix4Rz+Y2efEAT5T8
MdevVJf037fEDcm4oyJjP07xjvPM6+uJR1IXT3M4QkHIVMadz/8hj5Uq/ioAxCwEmt95FShH95Vu
Hm0NDst3UJjRcv/scMhPFJVYXiKVtA1z5cv19DEilq6EDw29EumK0G4RnzL6iJzJyq7SuQ9f8cNT
p9F8kUprpe4FiVXArLJwdAGM+UxyvCaq61UFq++A8AfatWucIbAPAvjuARpFZ1wlmSm7s69bRTiw
ax+82MQyUzH6Ul2+6/SF0lwp1IFbnkxwdkmx53qMlrwOhjW79mHi2PWiVZQZT8aqZHizj0SD0m/Z
TihYPWJPJggNbFmC9N/P+l77b4i37W7mhD44xe9sLB+7PmTEjNMtKrJD0ZvmogDx/Qu4zqUss8eP
gEZDoDAOPjsocXKWCIKaM6NRzK2Yf2b28JZP6iY/BP1kV/qzpJNGvIa1W4FkCnTeA1Gyysf3NcQs
BmWl1llIyUsPNDl3WcomFeh6ArLimEB8NsuikP0VZ3unZfuW+j/gDOi/dr6vEXbB76xc9gbDdgV+
5mmcgLR/QZysxL7SulsECxqA8feCWpfucZAB9vgJ42NAGHLsRWxInu+aa4QQWEg5WHBt8st+UYQN
rifhORl3Jj3ILaP5kzuRnHppX2AmzkEyPp2Yn2LWWbyLt/bW1jNn2idGQQfuB9RzhSLTI+6rPzmz
6GFkosQlw8ZRNCSHQncXqCN0mrEPZWH61WIRYUUmO8veyymBZW+vuh3sZ3qePiKxvrLCxVrzkgPZ
iDLYwv6hCZaDF/mQOrv9DWUpihXzNTZ6HNiCNv1ZrF2id0aEleHZ/ifu9203SRyLQNmisydR6BoG
NS94VcxRV868AIZkIdCVULqcLBEydr4l2uk4C4+gAmuF5d4ux65nIS56s6c7kTctv0pL5nR9iYdy
doFjnf9FzUw3PZYlFTS4LgsR55MC3TEfO1XfKe/OMvUYgT/KmHmMqn8JAr6NRuCn2uxyX027vNvb
nmt8iyBWehZJYkPsKMIDNYt2uLt6hnpNDIH7Cpf2V9rcv71M47NTzuh109y2cIpFuWwXs8thJf4Z
8JEDbsITj6IYpxovkfwfPBw9oip3bNyHlaJ8IsWfD/fyT3E/9Yyuh0Ga9M78oQxJuKMW/FZMa2kw
mMD3B0DXEVJZ+PCyklEuaDHPu9jjh0x/WUZGOnbTgQ312H5dbDN7Sf1tKH2dRrMzsi1+66ga4bZW
Yi5Z4W+nNo2oNodHJE/PBNZLzr3fh4J4RCMd6mnXtOl2snZ/63HsGe9+jF57cTbhjP5+VMtICFV0
cthhxgnKqxg3tOBYdmq1esqGSYyVGbsbViLL3Th6EshvNzjizDQimh6awckCZSOChQXs9ljGRBkg
JUkyNRJv/+jqfrIg2vIhGUu17Yp6oTOx4TA66IU5Mkg4bHZ2HpMvcMfyWQdFkO9ZlHD3T80QeU9K
iRnQDTFBuj+gxv6ha/ErqbYC2/WGxTalpuk2U5PHLo9kJbIOiRoGKu80PFeKRVjtG/i9N2mofmhD
kJolRlsS50FHqP6xC6caYtvrypIbfD/ToxH1XoaOSIwCxfMnwcoQb6MU2s8IvEo/ONgsgyF2UwXW
cU7dmzGpaf1C7xwvUZLbh0lLTdtPsrpMDJ9Cf8he6IzSjGDzlXSZb6cyM9Zq9sNnzToeQY6fE/M7
MoAF//PElS0uu1opBRTfyvDgfvZaBoPFv/cGIQxtRwpPMxGy/MeF+tOF8CSqE33tDxXCdbKhMMrb
7KowESGAx3NkxYmXeNv1dYC6P45ETtKevSZi3Gb+jk+rqievOs47x5KZU6ulY+9PXa03Sd6Z9t1O
Jjz0iodOr6TGGpA8wqRLrgOVXqU/mNJHf6rM6HN3Flff08jlNWMdOu9S4Rk8M82j4e5oN8nSnilB
YqvLCL7QRmm/Cwml/zH70LN7IEl3SUPFKnLJ/Qw3hVvgc0Udh1LSIS7oZXK6PM0t0P1rYjHKX8Nf
SQWn6pGsXO2oBBIGdzfDow9OEMtO1p60AM2uWE81o83C4bs8ol8rerHWIxIIjvUmK0nd34Hsz97s
M8RpBWSp9iAOq1ew1Cjocg9e11Q40y5fhTvYKqydq6Pb/L/M2Aj7Ncq5Q1CpgD8lAeYc1KpbVfzw
0jur1Qhdbj2tyvy5dbLnKM4OIG4hHvx4CR2IRu2KUVmDCNju9Y7tpL1cbiC4sa1bmEQ993I8DmtJ
HZhh9RJGz5NXH1OzBuHedlO65jFeCdgY/r5Gtd+6CouUqdq9dMD60jMWIrxl0YwmldQovRvH/PwO
Wmoxc0ihLpIBZvQt9osqgqYUlrKPdv76EsVwFFA0SiONYLDubp/aNI/qTuAYLdT3n2bD9CO5Forp
/tWyrZxwGTGiqUfkyPPt+VHpKtSgLX4qyIpevwg4T/2RRM746V7rzNhQ050OwpAAapf4Bjl4hTUz
s622C/Pl3CV64Jhe9v6seduYolrXGif3gqZribI0I9sMQNSnddzBAxywUFCb1/BiwECpnTbQNtoN
mdlmKy8cJ9iA1TiPhRekfEOUCj9zYZUuGCrq+1ei9zVVKQ+v6gSxTWcbmW1RmnoUWp12rGEXfWH1
VaijBxfe/KKZOn22exH5/WVQMpk6xpAtHmTqzY9PKux9upO5YP5mnkB+zMfzXIsXligD+VfTDAJt
CpvSW0f8ZyMzSS5jiAMM7R9EncZ0Zt/kDwLcdiV6aepNDi64b6d/jxcvCKojtV4GS9c51UIM6hp0
e2XqE+1PduYlWVvehZr1/c6Uw9+7HzY5/3eUZLeNNyPOZh1mVN3wmfe9+E6yAZ/sYNoTCDbvIo/7
v48YDOty8J8TfpXQ3eONSH4+E82QjR8Bjt5JMQhUegpAh9hGfxz9clnqorufVLk0DX2zpNNgeQus
JVdM/n1ntD248TV50JDS8az3IlTf8B5n1fjj1H83dNWVHuxnjIRpjHL/IIVKmMKofvYCmkr5mL/S
BHBkWhpDbzdUleAYKi1RGoXoCBkZo8XUKMR1SQkqzYoI83A1Fxt+FndKjNJrcSuO0OyHp+KtzqH0
y2hmvlXryc6//p/KMoAXqnGokLB5lRlSEB4SQ8hXfdXH2q8cHlEa/HlYP2+lpI0bOM7ecZF1Bb61
k+KjIz0OzT5FUPE2p58GpKtD+6MtEUk7U7vR2GzwuuSWhlGlD7Ej3pmhnDcPP2LPOMVtKCT1Dpvk
ZK5AYjDpvGK9ckbsCVh6MLT+Cb5Tv/GXp2VaVSV+UndZupyBh7FQL6vWPRUAa8LSC3muMlmUCk/C
OoGQzpDDiozG5erSWVWQ57NG1S4aZHmVKb/uTcy6j2CCGzRDlxcC8mwbd4u+OL/UJw987WqY5I8B
TJMsOnYAokM45L3kN0qP/MvAnJE9M+2d56xq9ODhFO+3ZDKTywpV3zq4AChRc/WhR53Xktz8IAX3
Lq9OYnJKZyRzjoJmKrA/7siEEAQEJY/35p81GPooygWFU+23mv07rjivfqeHTUuZ/F7gy1AlnX5n
6BYJIGb9e1EHP0oZAKzGsfLpOKNvRMybHJZMPYcmHNab1tcSFE58uMEj3PqwOjIOQV6q17/l6lpl
U30C5UOoe//90iEEiFTGow3s0buZsYFGWdfQeDl5zY8nMSpNJJNXnknDr4lVYH0xKLFoqlbdHL4+
ZRF0p/tv0B7ha02sNYDaFCLBfxfVrMHF0vD1y0NQK/tjiEYyE1c8oNmRvyPvXQBp5knOJUSw5wE6
7CdpDG/zr0TXQ+XdWraq76jWkB5CjS13SeUS8BdkEnBlN+Fdg5bQu7aFtA99zynXfoqxWuYzvXvd
D6pjha/B+0zMlpgNJBGHTHiWGdl2A3b3YPp8boioZ94cjG8GwJfYwAZz+M0oe0ZBZQcYEXPH7Qyx
Fz5GOdusG2SfoSACI3k4+q9NBRwEqkoTT0RofpT8uPBMF3djHnpCtDvZ7g/dvQUI1mzQYKpj8Jcf
+AKglqE3GkEuwMT32BFsbXQyLS+/By+JQamYMpxqL37Tpl+UQPX6kwbQBRf0IswuUpCd8j2XDr2C
GGboO/0eOnAJ8qgbhlMku+w2/XR2rduTvq76ofRY2LGlH3cs7HF5aCI7glPQD2EQrb/lBCa1DJha
KlTO02MinqAf72w+H2AKrlTxbVzlxB3Sf7G4sjNwNGcQPynlj711TKFg2JiI2jyo9i0hcHqKC3ny
bt3R/Xmdof2lHmJqXd0N8eukk+gTZWm+zM7eS33CuhXRKAB474xAprZfoWcu3yQXqcuNfIHindPS
lQi7hvpz1CH8E94a1JZCbOsjTfR8H4Yr/Ffz65YxTZhtgmGAte4D2Pr3aqzcw0r+nraBsdDgqZ0W
UIEYSYsovYsXi+/DSAm9IO7Y0vfkt6XBTmyUqcGn1CayMstjm2Ge/pAx2usIqiK0VCQ4KoluwVjo
5975AgxattdXgeQ5rW97ynIdODGBKntMwgH9Do2+9JYKUqym5mXT4HGg8mydN1Xrzft5kINQzDhu
sT7M3ivGCtNtLXPzXWoFRC8fm7mUP4S530rdFpUKtQdLYgE48OPFPRokk0RBazRxWDZ2rr3utozd
YN8uE0XEkjajlmHv7P+s/1mP5rUP9SqRbgspKdSFDqJQEBPZh7ldda6nAxpaEU1ApZ1JLzqHwo9m
ZA8VG/z4CDKv23BLphQLjDyDaT4heLiQmJrtKPgOxm3RjK0QRz3AQfSaXTSwgscUq/4p4Mi0guAO
nQXl7f3BtTfWxwO+h9t2FKZn+DcvZeT+hLsHKPhTTYYGgApm6RIl1eAFj1Ls9vDkQ5m5Wpkymqdf
/VBYxt2p5U4XBcO7/R5P9PesQ2RBmQdzJAIXFS2wM5TQRgmIReg+TVVerKx3xm9glfmHbp2T58qO
7jkCg3kvOegjkHhJm2mZc5BX6SzqMx6fQYiucDFbl8DXt1bPo3HPcWtuqjgiAE9YW04o9YkTV7Jc
Tn4CqA0MOg7K+5VsHbIi5sCpKTjzR37nsY3a/gqmaiH7WREf4DMk9fJeJWY1qVYQ9wwQfLXLgcCG
EvtSPQq6l6DlZN83IEI3Akm9NPX1cGWynQlhcWTTxB9NkjdMexwbKFXKItnI9LWPsRgdaR7ueNBG
FpcyaHZ1BeH/CS9uulLxEXjztsruyz5+0bzOhll8SaUcCohpYN9l32Eq+Vy39dmTExWyirTwl8Jv
wCte5IUNVkEru303Jx05G9KcR4TLyEseF3ILuLEMnyVX2AY4SXUTJLE2ZYFMQJW1UzcsXYEl+RIE
nwMcM2w577SVxnx+yd6Kmvu5rjs2M4jY8vaXeROkF1+N5DacB+30pNRCAhEAvXK1idOymI1rEn0X
oggO+y2HE9VtGCZp8olaD74YyBm3+kJXYPKllA5LsPnR1l23Wswkpl1Vmndeg4QsiAR66650w1Fd
zDbCutc6M+OFFck5iHfI3JtzODSKgi0xN/+9TOMjFtvyZGtPCiZkwKAZgAclzH624FT8vJ6uWuCe
9TrmhQ0c9xoBU4sMDatLXG00ofppRAa28Kxsaffmtv4lFChxEt9RA7/QVZtmfASu1ao+T84WwF3D
s+fp4dqNi/h/dzLh5kQ3NBbwqzG1An4n3fFB3aEPXTLB69H2rzVkfL2mtCZSGg2KdLtrdiUhf+K5
8wbL6KcAn/rgN0wZM3ONTOMgjiMVgoqnjhAZf1lp915BBYLzdkAf5V2n7xflkrUPUSq2AfFUpRT6
iUCRCIIV2FDWK65H9hsGysEuZ4Fx2G3i8J7AZjss9V8RzsmBfkfMLiUAQ7Jb2Ue+b9QYGbfCO7aQ
1lS0EsN8hfRSvr0E4UrtnVFhSmSDtxIc8QHBpabKhopF4RQADaClC+cZ/1GxPqaw9EjX4cm47Ree
bR23EYMavw9ArQ2+SdHtOXUAtdw9gq6NcuCI7FFiBofi7QlQGZkBLgLp4TYUnWUlpRfX4dMmuUhE
HnH1jGLAQVtSzTgcwTy6Xqp2AMndF16rS0WutNq/3Oxih2IVdhrltU74ubqPSCadArqwj3YGzElW
URbS2rRaX30tazRVaZZ/shc3BZhLqHa8SHptAyB/G5fe3AK0JbvrDSSirQc1VSNntcyINBHXatBe
6LIKjqD0BSO/L/0NJCSx//Lg53fumJdcN/K0qQARi4m1XfIk2g+/COOk7T/ARs2Q3aGUYEBUF0kB
+MwJNf02ADECXGtZsgi1kwW7D0dsWOv5fISy3uuWTlexJ1HVtaTUoOjjcQh6N8TD5gS2NZODnFiX
vKwYpl60Y2hm5Hc3uidRMUvonucO6Ug5tI2QJJLEftEdrNOJ9DfVHcMn3n2vE42a6r85EWH1idyb
9OnEKcpQvz+KEhUSrj13Z/ghyp4KNBi5LQJXnWpbMeUAObLYP9rr9C3FDBoOxoxZlwxlwPyt0gp8
eLuBRKZAfC2H07ppd0zeYYr6whL4UZWZa839KikWiOEcfwENsBRGe1FGUQ3k4EGU61UvFtDbh/Wk
pRLRWv2H9Aim7AefUzUXD52ZlWEImEO65HGhqnYW0xx+XQo/Cp722GxtcrAxHDsnexnLuYi6sTSM
DCn0ZsXLj2VEf9xOYvUg4X68He4vOSnrcahY+eWkTCvfvJYHvFxSMG6QbMq2atX2BTv+ykbCIKuX
Dg93P+JhFfWmZt1ndqcA9pZWU9B/VBZH/9fzPTRwQ0bveqwHBSjgnXdEgQJOvZJJyA4o569h+WxL
HfU0TJnzx/rRAOA6mKEMh/6Dr8d/L+92V443pgCF53ZpBBuPk6VjkLvh51qs7RrdOT2lsiyvEzAo
qIA6P5OdEoz8t2pg9r75zgbKxy+r3XQCiPOIZJBgl1pFA2xCumdi7eYtPauAu0I8RjAwYTkL/jz6
FxlLb9pGpeTop7z4ndiDjJafDvUOnLrcqD6/HqGoBq2vYwKP/TcYu6uFlAXhds841nC0WsrjRwX1
cjSaV+HxS6jS1YSsGjgGnnoUJzi131ZtMrRO0QKynvNU7qoJIHsplI27P7HhCRnDwrt68jJXendz
mRP8tNeNtkqfJ8wwIPSxXtRKVzA7WXv7x3k/HbYpyO9ec8Ofn987X2XA58yGWDDalXgDtROwnZPd
XczMw4KofRb/ugq3/duAMLd19uETDlynUyVQns87co8yQi+nxDFPPjdKmjvZG61UPqUCryoZs5hx
ZiefwKJhSts9n7i0ZaXLhqjzJiTBtwHt2KjidFYXKIA81X0gz4LMbwhZLgjKm+7ZhvZDlZAPV6sd
Jhvcw8QzpsgxqQ0d5vGVlI2JSrFQ/ILCgxl+rMDocx+xkt4vh56eqFduMYt+CsgAl4bV0KtB4YHX
HvlELLmzQbWXRkXMr5u2BwRy80eizRLbiGQV3VGj5xru7oOGLWIyakI+scLdCiKxwwzPbEzklhFD
ni8EKxE4Pvfte1Bf0KXG/+ay1CVLnfckc7mV67yeoyvrAUhnLbvg3NM6Y9qGJgGq/+6Y5hPrZrXw
HcXKM/w7mIXXAGp9+mf87SmhIr5Rx32ziGsJd+bAo3IfxwXrAgz4u26BBAhzjU9/W4i7kjyoo11i
NgvJqVvsNkQaxrFvI5VeiFZOfcGEUsjmiD5X10+c5gZ+/GetIf9zOXI2NzzllIGqtvL9X2eAceEl
ZuD/ALbO8jOfy/I7byw/ud42MD4SZJL5EtaaKTtgdgw0rwtuiBgU+S9FTKo/OBJwQCg5rHEJklwl
/X4k/L6m50ZgfzqZL+CzaW84CCO/GMA4KpgUY/A9fyas6Nrn2Da8GUeJdHT7ThIY836MeTXpL2UB
ssCFNt8qmtQPJRtNUr2DTGM8XyOu4aUn7QvRHd2wZxVJ0WTdnoKV5N7BpveYQKHX+1bA4aig2fzp
DYYvztHTEw/k3KxvaKM4ZVb9dvYZkWTAv2gb44LBOIffIHJ5EGPyc4DNgSB2uzjakl0gIBAIPtg+
AXeYu84Q+KfxG4LB7BCY31cGiAbVj5KRWa4hZ4FnJjcwP+Brqu7NIarMZyEzUI1m4lGUxzwn7lfL
DZ/Gv61Ys/eOJbJ+jncqYUVOnkB2M3Ubx64sMwbpR9fXEKO+VHSu7pTMFlm7AQo6YtHiv1EE2N1r
uUSCyJW1s7dPvozratMw7fhfm/fCLx6+UmIxw0t/nPcTJ2a/2Wtg00Dr1LO2rha9QuOI24F0F4V/
yCYwKmNKizN2/qRAQuMkGHVotPWL90z1IGC8xxXf1DMczxV12AXSxbyyRCQ7/IuV/aEnjsMlKKWB
X6uzM9/4xzFeo5sJgFNyMwCzrmQc6aKq/OaWC4J2O9MZ75Z1MhXsSb25qZa3RaTg+judUwt2ij4V
z4jUlhu1FRB2WufGQdfOzjyXKrcHP+m9iKff658+5EXKRo7vhJisd1V4zAJyMcMtcpw+lbzRhv7E
FIOBpPgqZdsMGqmrj4i4/pppYjQCar9dHULU/YyTlB6/poOpEd5sjfAj5mRjRPRUMTFNl8+dj0dS
DDEWghO7Acgdnp65t3djC56fm9yFp68H7XXFh4Bf2/rbGzZljvWaw0IgGHuaYLJO1C8AGuqu/Sqd
GWojaNznz6Z3yQ/yCw2rZjjUWS/vTsMEBwNGpTjpnSdrqtb0cv1HS7szVUZqJYqe/aybMPWSaZE8
RsX3of+gWSWXz4A2Ho6E0wE8xfcjcgA1Kc9aYRJKVAMQDL6m+NekHu55qJLmcYK1nYJu3mzbUGeH
ZGHNpFAXRbunvv+oTp5UHd3rrfxwANUm7zWyg5pmcP4ICKJDdnLYMlot3z2/fhCMxgVSxkXuAuFu
Y5ua36qaCuwFVQkb3KlxqE5AwOdwocotPNiHxbzHC/rKyaENmnz0cJmciz8SxjLqtE+f9Qli5FgI
VFjU080tBIX1BXfFVbMDiF3r3RUFErLGi8Sl0mq2CXReu14MyBl+NtYTAjnmt/T4VJSQysQj8wHl
1edJpl4XuwD1cupF5sZ11e6JQMjBUnTUiRXnhUFUB1dpVSgmnE5cIcFYUo6ZmWtpl47PsOSotC+J
NPaBdlMuyd0l/ijkICT5sWLG7A2sOXW2JSqDePSeoH2qf5JfeUCY5BlVbrUX9olJ4cDZr/kAwNFS
5/wZGYZd8aLYDqp8/XrqhUSziGCtNMJqqzgXqKsrRuCI1A87Gl+zt6BbK2gJOuxnJAV0prmOAv9j
FSJDGKGPADXggnJTvFT56R+UBBkquN+6RAccVl4/UULqBcz1mg8Vh7TBTO9t53peSULYmO8cPnJw
QxA7AiOXH2NLr+HBLUU4b4RoUFpFm7MMwYVifGWqgHQ3+v8Cl8ObS4LycYJ5OYiz+FCXOpy4w4PJ
YYp8Jop15m2vEUSo3MbcW8txWI2HhqNioWxbwL3kMaCxXfZyxho1rzwjg0UaDFqZCPv4UOo94UBy
N4ptClkC8RjFEDI9NaumknC4UR6pw4PqMoyQjD8wKB3DqYWrwvr81B1bJYKfQov4c96uyWI9Rcim
OlLbgQWiWgh3fm9U3bNfpkH9fVec1VnTYZ8x+9lbX1EH3BRTIFdxID+gsNdX3jJFXbx1+qb7ay9h
OWX/2amY7iN6Ne7gAL7djYUMIql8OdhpmycKPR/u+Bg1pJZIZrV7YL8zAuZZDo+8dybKFW5Zokbx
0P1dyIAVMZi02WHWjayeWrAsjBAFVDzPGJ3uyH+sy3pRbj/aom/p95pYtGVG6HAn4nj15ix87JIu
uUkUlXH4zCZ9UhjB7T9mw7/KhSxqcYsAVH8pt8SN+90LelCBQPBIhmJkjE0Q128R6omZJS7dKfk0
wZWNteuN6zIhxpGGq0L0u5NUKIGL3snmOL7qeQmIP2OLdC5T91rNWKAtwCvYrGHdFURthZB8hvN9
kkUPgu5ZkZd3oTcU6WY65iQvkg5TjuTusaGOxynq0/SZZjizuQaEWirp6/9QW2Y6Ui+CssBdybAc
XD7a7FyL/T2wYUhLgKXfjMl0LG6RO8kjZXByo8AlbE/fZxMr5WrYLnkSLfxGVcDE/Uq6bKCxYjak
pyXqwHB//WKAutavYygAFpWcDTyXDSsYvkTVSxcpftrnYfdi2gKefN6FWvE9B2RWfIkepbFGzuJD
ZBXL7rhm+ssoL+bMwdylAHMZ+mwd+LNHuU7zcoXnHrUJLCbyueLr1DqxlMOBZdYnBQXA4OxLO/Yh
308fKbVNDfbcjm9P+pP1wn8hP3jEJ3iLFmuH+MD97F8wq7LgYaHPsWxHLIcwyrT+ARn04Q2qEr7L
CjQofpz8b51wT4kQQlS0+7EjTTmLAtLIrq0dqtx609fH0zVeltGJB32S5SIhUHIUd+FDr0cKsTiX
32tDsVDVbsdXMxbyo4maqaChPPzoZiAV6Z0Slekw/a3VPTsfmDh+fBvnfIyRhNbEdgkC2biNyScr
vr+AOpIaQ9ogyTRF2CtmgMvsCZ34noOtXb2pzk38TKFQDNkhGP067nUB5ZDLntJG3/dP+neEMsQf
BtfX/ZSby9+setnMzrclCuVn2maI/I35shw7RCBSsgMInkhT982ztzk7JwzZtHdHGv8C1JT2sr3j
dKBBNONC/C3y+TvIw3Z+j5CcO5AA6xsP9iwX4TcGG7jL2GHBzqCT7QvkWpNSRY018X8KLdxwCIHq
YaNQVRvtqKCeD72bvocVh/Bmh4GnKLqxHbG0R7poNxi/Q/urh4hkjrHVDR1bq4JwFBNO9TW62PXW
E3MFANQk3oIH6/48xgefkGnQx1CfRXLPj5hAGJLJ8CzTbmCM4LAcPP56h33hxEuL+Ac7NBAbfUNi
OYVFKtdrl/WZ8RXVaF4pQlhRWULqFIUGl1wSiVJeG3rd5DZ5jkjU1LZgKi3KqGoJDrynvCCU3XT8
LCaXDwyTZ8BWDhbt5nD9ZowLainGh+UhQ5sGGhniZlfzpP4FqAeLXEduDKQAmbrWQ9slCD1N+y03
3jnCqDcGV76Ywob6BexJQvdzBK/U9ZlTZ9VQxkMoF3sBX7Um3wzmHfcVyfoqmDCblAEwTMVEcgh8
7WD61hCrFyD8PB8RiIuoPlKtesC+J3qwu/g0geYrGDAxrtASh9GVrxaA4SlFbgkZJzb84+5FlBkK
7zGwfns+BoE2Z41shcUvd89aX4YcgsXXPIW8nohAAAY7kxSjsgMSKww+wnjWjbKP+F43sFCr960I
5xgly2wbAFwMkoLiSnk3mGpR3JyuJ7gsFJOwNdT9au+61J2qoarmCl1CZY2X6OF3AJ9tAqZaIIzO
iAHDvjr/qNTZs18VCOo0nlWyfdXo2LXyQmD2Lq5kgRuEbns6BGgo+qqCC0nvnCXU0j8+k4fL4YTk
i0vsKpfU4xb2uufqCfRHaJeupKJkWcYWEkUDjHKXujU8j4WDnLIj5CEbam0fdRNAz4dOKMstqH6z
XbKGl6K4HyfkHj+6K+c51dslXC0FSm11p4d3905LZDeG/Z92aWIUNrFFMthZLCB6JrxsOmj106oZ
GNTgEy8Tx4b8eOW2EL6L9nhXujlAvkH4NNeXS/mTOXhApQneY2ZZl3m+8GLyh2cy3ybauLJTLqU0
DQywdHZQ+qnN6QF1GQfTi5LcoK9mio8phcVvj081nqsAUph/5kwCganXMBdtoBKixsNugrOvguap
9lidroimXQvHPVg80hqZf1tw20uoUuopsCVp6irO04l2cHPdwTUjf5W7jkeyCOx8WbZfwYq8+d0e
r8YJdRzFb7r77Rrn5aDME6+Xh5dLEpJ4S12RroHSY5pJ3HtoCHQ12i0seiQGrB2L6JxH+J1avjff
ydaAy4oHWfxH/M0XSdcSm2wZzsUJf/vlYAltj/Dv5MUBFXEBOdZpuX5WTHFd7mQzGFdQoxXpsXn1
qnLlr4mKBSDx7QjSCaH+XFzBIaZzReMAu2oQr3eke/gHOFzMYKnYDLx+nQVHAc5DgPi/V3QsT5Jt
WVS0KSbrKu6EqwlIo33k9pRRfX9doH7d8iYIsnGdu1fF5erTb+eUiyQXMpsmYuhm7u7Zex/zSDwe
iRiuWgkRtfyhoS+KhJP+Y5VQdW2hwKfvbGVNwuAecoypK29sJQtI5vLhrVANMU26vpTYrwTuRAFB
4+Ef8X2Zdl091hCWG+pd/EfXIXcfeLITKGmK70RkG6YLtTdGkwmYB4xrQd+gC/oQfDr9QuFoneqj
txkTFVA5N1ZyUl6ZsLYO5T3mf3G9jGKD7Acvo7nopUOdGVd78eL/gqE60oWVIK+GApOTtdvWjrly
MN3p4iX0bBq5nXj/QLJK5f3zwFALhumxxzfoW7JJCCu1euWolYNP2nl2aqMRbexNYoKHmhSBDASu
hZ50eZAZH6KF0wAUxJYqr3xUObjU1eQaWGtiBBwb1XOm0lPmLtpcyNqmK+CDoyFQpIluFQlUwr/U
eRPG6hoZXCyGrCtmL6s6MqVCMSMfQM1rzfWtin1oIv51JRcd4tBwOKXdaSjADVaCmgr4TEV+I/jJ
wLcYViSQD0g51ZGev3h58+1B7/S197g1CPti4qydQ38AaaoiP7OFcIM2DjmahFXLySLwhZjXV9Os
Jhedk2GLv7k6rid3p1m/Dv1rsGm2dTvQ2D3sNJy6MV5tj1I6eARm218APKEP90LtEDthtyB3oI9Z
VwKlYdqMbI6v5Ts6fEouhIYkCVdWdLhN0KxeAiT18WAu2S8O7l9D2QIkTPccKhzYGIU/gaw2e25o
YFbAt9FSRPwxKUU+J9jjvSorcIP23NOOSP0DcgHI7EhseicApWdCVXSuQqst1dl9Zrl2DUIA8s/x
Fq+s+6s6GlLuIvYw6sxy4RGax1Q7hNKQ9p32ogXaA6515bXXaWVb8gzgtu1xK5d08hYNE2fCWAAy
kzJAboWfFaemOzfu1DVO7nyO3zXShbXS9IUI0/3TtP6FT206g3Rcds2ZBcgnBqAAYzgfF4ZuWGiJ
6MdMi0CwX3EOiXSleZhcY0FbmBE2go8o+n+5E+Gw8LEtL26RrQM+nLhMJnAHy2ZC6YASALtNrZoN
UVt7DlI/5ntKAFcVANWyTDFMIz/03n4G/7lufx6jPXM+1bsn+f4wrWqhWFpihYe7Q/lwz8WLy4tt
NSHG6Y9wrX2hrZWGKCjRpdhyX0kl/kfUH3Ial7O39+h4uRdLA/0QAUQdo7xMrTUzbMwht6HKgczh
j16/IX6Fc0bgw464+qo+C5Fy7AjsDW4QGzkagodB11toZ8b6USbnvVrphV+6JXEHTf/iP/M0lLG4
XYW5lxylAZpxBQEnQIhKLPyj93+vklimxCA5GXGcQvtbf3naFWOf1Kej1Y1HPL+lZM6sBgjAyOqu
H+VC3SKeOyKoSOSzS0+2N9TTh07ko/C4zqiO2SHqGz8prglkLkQpt7oiD2lD9U4vPNerSG+WHEHg
ePdpSGVg7FqcRwEgzHJ3QNixs+2NEKKeMcDHzcMYbSMcgjzDi0/Of5ckSdquxsklNPo0WTRz1K8w
fJUUho5gwfnHTCsLD9/jqCaCcOSUIYee9EFLXL4mwtgCM4v9yXFBH3aLJ8q+k4NNJDlCBoWgpwGx
YsWIK5Ylmy+BCGgHtJlXJVgS2Fbua1aqApP/uuikPT+OIHSNv87A6OgizQPcalkeCls3+rpIxsLq
cI2QdVAyQV6CMnxckky2s2SPxcIknnrdaJohZ97edcM+BTOJUz2StZAd9EDBdGSsDFCUn/gtM/s9
z+JgTeQ28hbU/TCnordtNQGd9a6KdPvF3kZyE/YWoU0o9zhZK+GrqWG0k9YCEvxmpbH2QjnXlBx9
dHIs56NyfHRU7VybtF6xmdiKB1p9ivR1ovDxND/zEDlR6k73FNYuPqsWKeCj9c13irdfZxl3JR8G
YfA+CASXtBUGxo4/ciVrcFbMfxjvf5Kmmb9AAnFOpiMJHHUDIbPHUyf5AdT/adnw9WORRj1aHWGU
L0+77M6K4YarXHw8KigGGpOnBhDA63Y60XxISjZgb+SAU4TllkncMzdmaMfXFhX/9FsN/6Lbnle3
PqpEAMAnvRdPdPK0fGkqJM5cWp3ng2FTJtoOHrQpKiBirfM0GEOfrOmweri6XfsxczuWvfgkPrUZ
/4jmY3mO+06c33mRYkqxtqTuzbzHx/SX866RIQ9CA6O3ro3NLlaBsKVvwuAWChG8IApziNUc8PM9
yWmbctBG9zQg0mhHiBN8pmQpCHwEYd5SzPQDPXmfOYoh4TlHxp8HHd2LolX7UCyGbJXUj4rsOBbo
ItEY0fgT+Ce4iV3IOu6j3N+PvgCDDLbuTcgoEMTg4SmqynsGNJ3kh6b1woP1w6XSZNwg9y+gGIgE
m//PwiY79N9eRqOMBW/eiHITkngv4pkDXxpxd5+++YgBjgVYoCA+5bTXwU9SYLVemIllyfJoGbdA
14K742ZMg8yngTRptH7rSSEwkezYhacEsH2HgQFbnqmvIx7Vq65MVQXThiSU+b78R2NUlKhPHDBl
QRnRYVZ++lHdkXrxLjm2txqs8G2hx8XOvLLKzviMLzgBNOY+yCAh50ZaOdHf+rMgvSraLzv2X/5I
ep9vHBTIHc+PN+mA6413cFu+CkFzroWNe3c/t1/KofutU+Z4TpAgGJ1hgI3qZEKPMj6v5WeR9WaP
NMBhizWnZFFdwF+mNBFgdgZ9qf1LUtqUkU4wGN9YreXIgCcTdjHtW7Y24u/GrM9W8yOAh3nR5V4g
UKR78l2iqKkADnI+oPxMWAjs7uPfxlzHXMzGCfZ45lR96fsjrhNQjm6CAiF7LKkgKV1QWp2AvviG
Vj4Qk5x/EjRfzc4NuJniI+wkrqEuhBekmTf50q38GjXHwSQo88TldW+1glDBLm8XDpP2m+tV/XtD
1PXgAwcoRIUJ+CSOgxMtBWrvl6GchNgjxoXcFFrGKhjeFsx3Shnmecs/lkOzO2+hMZ1so7XdYAIk
l8fMNXX7SIqIuVyR1KgR9GMOrGLBWkv500u5I8VWqQfYNcDK4O28e/0Xg0gSBlGOPxQcq1VKy2eW
NI9s8G6pamYMOgU5hXPNdunXmRFA6GERkeaXxMPCjWmIUbICBS8KhICddG64OXYsKcRgIUNXpr0k
fpTAwQpGN0rBZV1qgUiwMYq3wgVHKBrh6InctVpS+kXNxpmlQlrlW4NLCugt1Z/37BAPizZL7nA4
bm5Ylzd88pyF9E7RXgIMlVC6izWNvaqs+H0H2GKODkjP4py2wASxnq0gMnYw0s6o6iEAlm15m7Mk
RvaKT2Wn2rpOWEFZxvN8oRWPkXAkTb615pgH1ZPRW3wyHZ8UDaWkyuLQj09jEOGtUbKiL86Epw7u
BbOiK8qod/Y+dgdiReyq6GS0nVNZW4X4+1gr/ol2olWMdOCTH1NwBve21mNj0RZScbccBCb1ClJv
cHUnzRwnJKCc+3aAn76sc0EYa7iDV/gX8pJRIcaSF/81csLBqhxN7Vepwm6mVrFAnZ7L/380SWqZ
cE4JKBKJtZr97ToQUZGInSI3ppHl1hcFdW4c32H32YSCslXBoJtPewr4GdGBTpGSvGbxYos5khj3
n+1f3gqqoH5Q7jkC6N/3kynatVbPZE8+aAbFkxQEkDqKQSrM6+5g00ypnaSEH/44e8qnhNdQkSOE
jfwfojHw0Z4EJdbz4i7aBt7VtTC9OK4J4StN6Sgiq0zBk52r3S1ormf3/7ILj8Tx0icFh/pu5Wl9
0Zfa/Lym9QXuaafN/oFcXCbU5rbfRJiBbc1hv5AU9YK1TcZWlXxWDuQgdHKnF8h33dIoKmYg6PsC
dqfg48aIC6fgx/oV/HwcbeZ/e24rHJccYi3aElHH5TZM8nIIW3V7fGvAHjqXrCwMQizDKQOAlB1q
/Nw+UR5LMsgcIxzI0m3cNlgP17EpX61oVI38KD+gLyT2EuPlSnAOhgIijWDqUuV36EzmHJBxSXFf
aTqlaPwsByafdM58U0UWWfE8FhKk8WrfcF1uuHBFMZ6FK4XWsR3JkBHXGblVutfMZirImxTkbESw
WsQEVLLyPwuDpkTLx73/gNoBUFYUi7WDb8/qmAIxsDDHr5PlIdhN86AZ+hWmaFToCsI5ycUEIeaJ
w9sH+y3vepjVmcClpQxcozvSVixP6HIlAQYKt9APEOxJh4JrmkrTSfQUkm0dcJmF0d22hDPo8gwf
KU3/P55x1DdEDOkDQiMT0YHWD38XqxeXNqUCTydWeVIIPGFOr3pfG75EsEajymXuC72Kgp1TYR9s
/UR+l+GEdmxJacnJ2LiM0PgqWXtBqOyhDeVixeMbCIbNKpYOZiJ9wWumLT09tqrlxWIlsrxJYIO5
HgU2i3t0fY+gAvtPXvYHD0z0V2pJEEiAyAlgprBnsdOQwezcqsE2JA2yWEUDGIn5wmA5Kjm7pKIE
mQD6j4ajvRWWwSn+idAh7AvDcqdd10n5cI7qvG6Rild9MOzXf4PVq9+tJOI7NeDEDHu16Jr1sqBE
R/oJlAzHdnvHLtMQEPiu7viZh8ivm+AC2rqmY2apQp8lza4m03j7a6uNDe922xYguxqdiiSif3rE
SM9EnrI1wjG3L/scw2N6LkBvEpi8Uqg/P4tMvTP56e+vxgL5hRik9N67KlSo4b4pDh7kR18I7ozl
gIXbffo5SwbD9pFf0YOKn26iRcmel7J3huyKH+zHn9OVRABqy6NfmZW5+dW1V55oBdME03WbwZ8j
P+4XgRCKkRqlTWLB2o/EttUGTzo4TLQzfqC/GVjHgJTdRfCcsrfoWEaYi6IRHsjqCfw2slFJsdSw
iuvB+C1kBDHAxQ3VWi0VOIdjvPGncVumrtglbVyaZALZCML7e0ynbzdTAznTcoj0i+pxRk9WCM0K
aCiHr3tV8VxTUJcFfT9QqvvGlVRwu6iMtiqKik7RGRIGuRlPLJtz2IFFfUj4oQYR6m38X4XVWijJ
2uoh9zW95bW8XOOWpf2003bgSc/7351l0vu8949W+otLrciCdaEbGo4/ynbtctAP2aauFlhT3ccs
t2m45rpFy+z6i4JvSgfJxgC6Fg4vHYAzgBr2QLDc7h0eKY2EiPu0X0TLP4+KiQhUH4oOr0z17Ux2
tHMtQs/iqKrhVrdVGjko4PGsOprikYvkngbjuuwsXWgHr3f96ZTvesvlfj9wToUkaLIkpjafzwsv
XQ2zTfegqqHwhFIfd817YOeeCr+JvYoCga8Dz2EuInOGS2oxDBA0QE4/bcLPIZj7A6X2xp+ZGAFD
cmdeUp7r1Exnerw9cpOAzweokJlaE3MixQCLA+JleytzVoGaxCYrfqxQHT5oPqCcKu3+k8ECiayx
EXtoF9FfQJu8tCR1b3kBIUd0aadQGZE/Aci1u3IxQmc0SOAv3DCzK3zes/xUgdcbAM+NnOR5qtSA
weAJwHSN66xO6QJy/X+kYbF+wByUgRgjnKineab9wkqPuCmGmjTniK9JSdfz9DnIgKJGvZdeupXq
/89afaQ5nYYhnkURk2fV1/AGH16Iq3FCKaZ8RLPQ6OfevApZUO71/quzOOgvV0ZS8o3XayUmh8XZ
WfqmDoS2aNe+gz5xLW11HYAQTtG+iPQRwhJsJD56GjtbK5h+2zFSFyO29cNEd+PIv1BBdKJ5zhUk
PMDcBRE5WAujeT3Vt2Fxi8m+PV43xA3HiQjOnBZyR+K1r1qM09raLkHixr6wHGWRo5ronbu1j3lI
6qsP6UXb+VJH3i5iCncMOwZxpknkUbMTmeImz8SeW1MTbpz4FaLMLIg7Pmk0gxhx0hjt8Y1ykx76
0ZtwkiRBQ2U2f20DGe4rFzXwPOXufiL9JmLxyEmp8s2vqlH0kixRiL1NeSZnqm+tI44rpBdCisyp
qZwQR5S49ilZPpJhPnlTdP36iu9qEW349HWD1JGBV994FkMFVbqg+7FwIxMNfcwklwnIXtrVfO8m
w6FDw8FkqSonFxJ1GjuE2hZeuoHy66h77dp4ZC65T55CvLyCCdtrb228ZIqIBKeTUM7jkCj2HdzH
CuYv7gczjgTksD4TeYp+eZCKT0vQbiB7YVtkEA2dbcHOedc3DQ1JNbwKlIvU9j9zUolnE4FtB2xz
KEd+9SZv49KU7+SxCk6t37eULAYnEzyNsguCLxolcHuOxMN1x/be+Uy0xxnsYO7xlxf6udUCqHcq
aYO9UPcDPrwcUIyGGhUo3Jkp8rrVyE4+MIXmfQBzERNXmhUxVTS4pfD1/ym9hj1uADCtgeRtplZx
sG6jEpGsoQHyU8y4KiEjFMqwxqLQRaiBRYy+Etyh5DMPTL2HjjoJcB0aFIzEedL7uRv5FvN6w/Nc
yprsi1DkHO4RriwWMfsBHbZskPwV+Vs9iXUjt60uHSIzoEz2tGJ2YYbtemQLlJmzRHXbaHcxDtF2
sT9kEBHhnOxAnuDB70IdzQJn8rIiJsXLASDMlnP/4Qm198E5yaXnXC2w1gXxXenpZXAOHdH8TFgC
QJZg9egdX0E1t7UwDKhY4S9kqha4+A3Vf1LECfD5tdOhPSyB7Zbrgk1NL0URlSy773D4fEro/cgH
A/59ZljFw9AEBWvJ24o9lqQTpA4ljlCj0/HV9HCrog5MzVzoT/h7PahJvR8wMeEX5qN0A9noYKOR
ViBM7lL473V5m7m8lQgRJ262MPsEs0snaAxxo++T6MXVlwJx4WM5DwdQ46MllT0Qt5/m4T2LjuIr
zC63f826NXgOvFUg+MtYPMsJulGhkAlVzCwWheEkOBuTYSMNwWX/2rW93AaEbg7zzK2F4Cc4k+aS
KrM/Vd/OlF9znNZeEpXNxsgPTWjrl2Z5G1KvaFoyvMssI+sqCdDHynpJ4uz8J8qhRQfyvSkd3wS2
pEmFhoOramkXLQ92eiAbxw2rfAJ7eaHoAXmEgxo+uOyNgUVNbuion9tut2+5+K09quErOa1dzqur
8l95CBrwUyoO1ftZQkekexhDV05oT2IhjCaS9pxmq58cGl8HMlfvMkU9eYDeKPvTgD5mlnYQTBst
MZZeMI09D7Xyad6nATwAalp4w+MiuzLtlRZ+k2Izu51sv7mj63D5mdQXy5dIqwo5c6xB/lNextfl
OuOqSjNRKYdV9eRjCM+fly1eSdqcbqABBJWGg2kHNlEuAT69EdMsJWq0shGk6GTeCcU2a6xqi7HC
BiLTJ01GwJ52PT5/BhqpJ6pWhGP7VZMgmSQHQpB8JiIzc/7WVXPvnsbrKyK1wOZMp2FkRP6faCe5
EHG2X6Vg0qu9Y8kdIBq+lXcGQZEqf54ObeiYZw6ZBgPKE8knNur5J50XU4qHiN67QZFJqrLj41K7
pAx8f/bNMfiZ6EXK7JfGEYd9u05VMWiMV6ekb3PJ/r4u+XpcSEh8qavW3nmE0uf3oZUfX1IFIeAU
8HjZVJELTWuKfaiUUZdtQjd4f9QfJr1bDP7gQ5kFi+dmjcHZuRiLXndRnHRO1Msobh6saw+tTkXj
cHw8p6LvfQsoD4m/jB6azppLmi+sDu90l2ISbYTupvTkRCOWtZJl3HNo6FJ0KkBTiCZy17aZvC0E
SHYkLugz196+qayVOBJD3e5N5pZJgj3EhrdxrLjoIGOn3tPaYurbjSE3aAN2lZwhWGcNHtMeTyuy
dzGIJn3jmSq1nd88SOl0VSuZZkve5HZj1L+xtNm5q2IJLagNHmILAFxKzgphAhZbBHqylGuJG4ZO
GIICKnOgjknsTrch5ySWV+KSrNAE1zHJcq68he4i7M6F4cnlUm05Z7UjRlNnYWOQI4VIxtL2VPmW
11011b2DGUMYhQOqYsJaCFoxJ1vVC614euXd5c618671R6kOtmlO9yV17/VWTQzVYPs5K/Al8mlt
iDjXYff7MvooebFBeaM3g5BmCzUFzNMLwYDRCW3FLystWmZOaSRBYc2kr6mor8Pm6UtyvP2xZIwX
rh8JZhznHHLc92mpCAwGpyITXpBOPkJgGvZAGyj/9HqGT5t1MuqSc3JhfEgnjpBYyR3EmDbDPrR2
AikWZCVWwmCYEscxsSQpAeUrtslHOUIrv/M/2uech0UB73pLvKONOdN1+ZuLX/eI2ItjEyrP5YSt
toDzcFPDj7MDQamaXEyKT6EchgxwF+uGcWsVvzuLCR6sBHuOIh9ffTNtIbDzNhtH5NKZxgsS2vTo
pZ7M7qdJi5/iLHXz1a2mYyMw6uSOUy031Hfbon2KjSomUk1T63gKf1JdmNn5kS8aLK+OF3GM7JWz
+fNQzAc0yGBaB0m/iWSSGrHnNodYp1f56J5p0/K0xswr6t635NiVyUzIBFoDcw4IQk+tkTpg8f5+
/1ff+d4oXJBgNvgorrRS2yRYD/Ifpxl2bMHrC9tGPwTMXEf1xTPF5zDqMiHcKBMdNbCoMwwSeLFn
6F9PVkm/ly7wdtMUnajlnouF1ii8eBJBTqbzVj5daY+771rlllS70zrnEluxNsoXmrXsLZLgGTQX
CIdncAY9NYucLmuXUbVDPEMpGCnaRwH743TviUIyyfRwu2dNmETvT3fu7WtFcLnceF9DYmz3owOr
GQUWog8QwJq1S9zzQ06kz2u7kssaArXSEqn0oIka33kBDvp4zfVwmp6hlRXWfiztVTh56MNkyioz
RmSjrtbrQZ2ZtNKVe2WrDhCgTaju7s387KgR6HYfKlkt+uWV1xU0Bge/rV2i9U/B8epEfpr0Kg9t
FJQWsH1TNxpnOAHXud5IE/ushepqGDI49jYTyHd+ohYRnK2/s/TBIMCLHnvzfi3y/p3GPS8BLHQl
fiRTdsOh9bWw/tK3wNN7rIPZ8vr1Nqc0eLuRfjdmbSqbeoA1/hhKttbAmJt7lTv/0lTJAUh4Y+js
JwkveYutuZG5FqCe0JTS3RRHUFOxQv1sR5TxnHP1HKGdq9Lc73yV2TDfxd58vegODxq/yTkkNO+i
MP/oUAkyH/SKuanOZdlTfcalAYMvk4mISuNW3DkQABiX4bt+Ym4cSrBOj0Zx/PwYEzUyeaj5ZwoX
2nvgqS6BagKOdIbPw44snORO5L+57pIGg5+QEg1BXm0u+NqX83Bo6eham0GdaYuPIY/2rsFYlWnL
j7mVetyeiNXbIVC+0fwr+mJxni84AVPbRzXngY2KIyXncsNZ0wRlI9pDN4SjNYLHRTb55g1kQLii
hsQDAzrj0KokMaYi1ZAEcsmBK3K07Dmra0ZXVsElS6YJcHGn/T19cGRNT9mRdKPrNCGbccthllZu
jtHUiKcRJinPTQge1jJYBTv2RL+5BeFQLQz+79D3VI8zePr11FUsnJp9Wf2pJ3hi4WFVhsw1GfBn
09HxCG5VhaZNbsXL5xF+povN9HeGc7M4uxOPKceaoRN/8dSsy9FCVzXMN25E0qqWWe1LrVsBsXv3
lst0zdYJQ7f9nWVc/Cf4TfB1iS/+Clp/ElsrTtXCP+/TxpPHo9HyREgLtw4YSxX8chHE8Q5bVY6O
SzgFXEFBSdi+5Bqyoc6FOkLFEyInfL7ET9xDYUHnc3Td+1tKmb33Tfy2+21DxVMxQOKA9fvOayhl
iaqu6ut1B232Eb3IUtVcN1H6KmyuJ872H/jCz+5pNj5G9A53RfquAnaM4qNvAXGvuIr+AQ1ShJnr
AmiZSDpi64ivnYwhvmEMVSey1NaJGo0dkJ54PUN6EjVQLojibqw+dqzKlB/yA/oBHdqTqkjg0V4C
twvfvtPB9ittfZBJ0CHbpKFHJHL3QruG+jSG6FP8XOuxCvX21WFW0DhCfkWYNiZyrgt94lBmUbBe
niykC5chXMqCnWLy602GYNb34w/DPSIDDZQAt0O8Om9FOUY3ZGWZ+PajZOH878pc51/JkkIUq8IL
IdUF5PcTx0duSdAExUb1yzea4AJQ6tIduQqNrTNa4ZZlp5pDeQpG4YGBeGYy6zV0qc5Zb8WKc4QP
27DERVJycUogBqeXkkWeF0tgnM4Z1Pe0mRESZpkulhZIV/tvT/U5lZChEwhsnH7//RmkmQLeDpJv
ZQbhw5YglABJOd7f6euYpR/+7eoKVRVqeSy0Vc3I67BCqt4tUtWO+cp2fxGRq28jysR4Qx8QxqSy
wYM1Gi7ZVhwvjcp49OxXrC9cvQsJVQQFDb5A/fOg/P3Kcf2vP3WBbrMoHrv1qwV6UQAnaxgeOPwn
BK0J94pjz/3rYj6D2MiOA+hd2t+yFJS5/ly72BLXYCHxgQ/hz7PsEEiOY7OGYUJyUiQoSVQE5LyC
Hh4XMZyfJzfkyOz2k6xZrWRCIkSOPjwM3wykYhWWx2WlcvrBvCs9p754Qk/teKesgR8JdlaLmHcc
9QHKFAeVJ1xkG+jFeT3Gs9prA/PsI0i8GodpfrT4EXhqYgERtQEByFNUH+nrBrNUYr93sjSqJvE8
aSortEDlcz9G0dNw1OQY0HG+GsReAq4kpFiFcGM1cmH8bML/rHeet48B7kQZnYCLSfluCGd6Egt2
p95fhi5RUhbg+UjaS2+qAqB7OYFH4ioGkWbU+OAxa/YAj2/Nnk2XStDrpd9VmOPTNkN9A+U+wThu
TREw5wO6G4Ql/T7TJK3u16T3/fcrWkmANTWMftST8vcSY488Ka8yI3W+LMuG4I1Z5OOqAt6cWzd7
MbrfjkbLN77ff9++Yg9EdxspwR9Hswvpsx1iBAuiC4zvur1O/xd5MYGYkBuQUZNAvcXOAcLxFHiN
hP7HUwqcMVbp8R0eucRW80+eXiA4kIQ1eVS/nrXB103iibvckPbU1TaewcD03NcVVsJfRGhuvomm
DqNMboflzmeO3+5kParWG2qUNmfzIY5ZMVEIBmJsoKe2jD66Wzu/oXMSyass+EnfTJchRJN6tOxD
HDUrheKrD74iiwDz3P75iP4uJM6R6MGprogEToDESwqzkieVgUN/Xy4l2rUnI//Y6ZZqrIptXh1h
tEgkDQ+4X7B98axQW3KMCOhJqlV1we9pfPagXmSoi5Oe1Ynd8MHW/Gw31ZjTwoJO80NW6ZW0w9MV
B7tulMlSYEFHv3qfW5J4hJcRGgGR6Pn/jFsnJuX99Nrlq2v5/gKbvoNjh5V573Rs/Apo2dySV8xE
nk8h1nnBIYdnKl9hXNRf/6mS83b7XnMc5TAzPr1tCokbs4wlMIzcvcmyLjf2o0wZfSih0hlL1MES
NJOaZidfuv6xw1wevwzUbHtI+58eb+50gH9FHxDuzOeBYRYo52DwpipPl33b5y9iWEeDTy7XrShe
RG48xANt7hgI8ZeKeMDqskNvsJQDZ9+OPxM8iZE8IFgtumDBLr9O5r4AwHi9WP9TMsq24My418Jy
Ufw9lsu+8M3oicbPc96WLxYzg2q4Vw8Ow9bB5whiwEb5afNbebEvCGBcz+bIGlxi+sSMXgv8tNfO
TdpFfuo4fXQEb8R966TfckhOS2N6yF5hXirDOi3xSXYCKvlMqo6BeTneY3Z/PVl9V2EfEYF976lH
s2KisjSMsvObkbhlMjV1d9RgiX4rgYFGqMjsFpAfIxraknBpLJhdDKVh1tYl/CqTV/l8+OytkjQT
2+dWkqAv0OjwSzYTD2YewowqJhHEB8BWsAtTQi9X+RIhLAhYeuwz059xCDbrh3LFvEPGajkaood0
rUf7Nm1E9I+MYMOCb1CgQxpBc0FwRnm97TPrMVMrtG1khZ5EivMqSXETN9SMu6GG4Drm0Z11Aer2
PVCVmXvFXSPVi+lWqSfYp0CsOAQG1bhkgb1ANsDlXc3dmqXClyNcm14d79DpUcHA4KINK/47ZuoG
LvAXrI3POUNTjzJP7KQc1zl5NIubgxWNg4aaNxewz46pOAK/sUMYLiedjpB5oWIFRHGOS7vqaMyP
LkQKPRm009mLSH5OvSQuBFwrXjjDZ6FcNvBdTPvX26O5kIyA3zkf8Nj9VdfwL0d+Km11Mtx7ZKa5
j9PeX4UR9OhVpFJDQTPPwklQOTEwmiKsCNlliYhghGUtv+trj+hT3aYQLf7omCIWGpvK6EbPLpHI
IWd8ySZyzpJn+yF1CT0+Oc349lIvKT3jIMxzlsT30ZmuQZ/a6SrfjBMvNj3hYWM8jHOBUmGFRHNO
eshtd9wyURWSSDww0KlPe5rb1caIA39Wi+sxd/1Rv6AGwHYhbW3nbi8w93aHMHCTI6tQBdOo1WEj
jOwpnX5b8RD61Fj+Zq3+f1UknEg1QHIQ+lOVqfhSE2npNdjR0dJuu7h8yllyBciqZL9TeKrZMoHM
bcwl6ID04GzK7akGS0/CgFBmUl1md5Y2msqchXQdO+0yGEHTYbyd1bCySy39NbPMZgZVQ0DCI79j
aQDylZoALXHyhecx87O5QglWBC6ZywacsRVtXMFXi6DMNBxK/YNKFipbgfXDgBAMNtkjzb9+08NW
4ufNWa7hFGt59KlqeMGvqkqHzmbA7c+8QNkv+Aj584T7aPDgf+44V523LclLsnZm3U16swM4+Kcf
Gr6bzBKssdXPcW789JWrogckAqT4gn87zRmkrPN2qUzf13TqgQq9BSwO7k9Y8ZiOBOHDKn4vPmaj
7uUeHVN1GwwQnrQohN8SfqQviqtf+VUPG5nbR/gliL7ZbtY8ynsYEA5EuMvvpX8g/7ViHssjUi4S
ljvCWYOsJdjbQyDIEdyZk6D+643jN9K/Y7xSycjhOKkMU8sr9Xk4geR5LSNYqe0uzEBd3lMuIuMT
w8UnAyHO/7MySZhXQJbOUofaVFtjmWEGIm87OlG1MtH3lfXMrmlsRqCyDgjhDkS4fILVEgWSWJJD
Hry2r6nLL3BqB2Gvg0SlqZlGn88uEPJSmdHanI2VkRsMf+Hn7OqR3l/5BUjKc0Y/x5RFTZr1hURo
PmGzanx98KbxrK9BO/ke+Xb1kk6tmupIncOHCEUaVw0k+6pBBpNqrPsNL+nWJ9cTusxd8gyiko6L
4J8QxEc0j4T6ZKZGc5yegkM0+gkNwbywC0nnygZxeMP45c+6btNFvj/5sjB7ArGgUy96rH7sq6da
wN9oYzK1jyHPS16f/ap8QaQ7i4m1CoqRbXItPoRFa2aqszufo8HXnfVg2qb4YJZaf/OrGNQEauCN
qKEpiejTk7546t766GwGoc9g45M5jA21gYgXlHGU/zrH+nRx2ApJlr5MwQ06RYkNgWMi52bYqFw0
9jjjJVeFuN2hb6XBGZHOhGO+f5usTGuOY8+z2AvApbaUbkly0Qidu9daBgmx42ddYaMaHLll4wgy
1Q5HpwHYOCsPDj+a0DLPrEFGusNgYdiOwYDpnnIx5DuN/l2pyObDfOuGDaZYYNQ5SxhIeVlWXLuw
4muzGIBY2dFB+BsRzkwPxRTIoLa/KnHru7gFoRFYYaDlHOmshke56kyFkgRnZcx5TwKLLbtQk5gI
83R8+s4QHCcMnR6j+6TTFC2T5aSosXsYCsLm/08fdKuL4nR4b3IPEOiS/H8Mn019qDQ3CRk61/GZ
AWL3S7XqCOXyoDjjJl6pfvuzgmRBghIx7G3wSu8eVm65bMDV8+cjK8WZkWKovjeQ4vypHmQ99PLT
nq5XtdENaHoClDXWE3zBUhsT6kC3L1+pfed3UGoAvcV8PksprX+S30L5LbG+zLvuykQIQzCeaJuA
2ajqfgkkLELeXLgrg5BfpSo3AplwDbNrkQaWqDG3O4zy4aJiptHBeuNtBDlUfUa+t5TL81UYYUys
OXZuOv8To3QMWUMIuO5+EogLI+JQF4vxOvqzGeNfrzFvdHGPw7d9qcguPZtI9+NuZ4IC+A9sCENb
j8mVtSpPIJWn6R0vsG+Q+5QYX3cYrJOJMNN9g4VbA4+8crsuW58s9CyLQWg/yZPNkm8rjwibwAVW
kTm9gyWwnBluNzGNA+oK2lE91MX3aX/vuYQ+xfgDKX7gxc7S124EcBdDLNWHQLJDhM22ELG8PQka
3lsVSszwVAzgoPJEH5rMTvDmn4sJJOAFKV3Y8pIGktKhhnS+LheOHPV9V4Hi6Zub4vIQHkDHtyho
qmGIZ6rZrIk84S6zfHL5C6fnH6m/uut/LdgU3V9/UR3tqUNJhsHrydX80NOBEIhTbBXu7t9GqJlj
4Ke21KnLa3lcc4eH2m4YaDCs2XQQlB4M29LpCdDoM0w1Hvd2RIgdUmK5mmKh0FiEUESWWocO40F0
bGMffe5y4LCW7b57SMNJKjTVAHEp3ai7YiblokDzjmyZejyjk6wAm7NONfiC0UmVUk7OaE5hSE7x
3vADP6jrwW6Luv1QOqSDwo9SUFouayBdJgNVn8qLqOqF7vj64PRlw/fYHX5oT/P0od1K2Nm+Ku3s
c7IveRrufg6s8pp62xc8c0XIlf4b8W/0ObH5n9jQgYG/9C+3IJebK12V5uhBoIIhIBwpRrpOhJgT
zx7C+nLBOJzuEKgCfebDXfXtzRdeqOZZ6pyUT2Art/Bg1Lxehf6up6x3UGD+U303U44HvRKBZ55Z
dSFaApMG5tKoKkYcgONrqRpWgbLb5kAqgzL/v+fBNjmSacVbjfsfhw6+8j2kTC0hx9EzimtsFKk6
hMpSym9L2m6zHarVQhlJT2cH0pDK5ta0dheTjDmNoOg8lCzINydeXA0O01fGOEQy0jz1g85Iiulg
Q678ztCUqZwgO4BqbeQtFVPUIKP1yjXTXLU/ADowbY92fxns7woR5ywIqm9qp2XznXFGLMJys5xY
6j5e8JG2fg/wugGUaya1gVJb+fMn8mgBgeAnrZTkK3cPwbVAG43JBTEIKoaFZ6htjd8EqQo/+bA7
QgCNwUH2esPu4doe8CVrSJGD9OUh9fUKLmheQQlGz2gCYvThS+mC3mHr4xV77Nj7pt+2HjpUBdn6
FyL/1aorEfMDmNeksciOLdzV+HpL5eChjZiY4fBuEk8MLQ4+5oU2sMcVk5b3QVbCAVVgmo+Vf46R
oC4AlK3Ho1onPIYWQSr/luUp1DfSnyvs+kEQO1Jc4siML3uplFNfP+YPa0cYnD4AMwy3OERBKUEl
nJ9ZvzAtQSgWxZYTt5tQfDyQG3SCe/rAq3yKoq0nz70qJN/+PN4HPbDSXvjwqIUUkP6/dIkKuOPV
WHJ99YmIqtwX03l90bHj3k+yP8ahgpZAr4FBZnp0XdEh3EZaouOffyy4iOwj0ABQpF17GN6PBn0f
UoP3qhoEgHU+vdWihEQecRa7TbVg5OXIe8+pLmsDILrMAbvPzB0/zzFoE529oKhIKqE8XXT8/gPw
MZAPsRNiGTmBFtCZz84AjIbpI6EWC5QsNlLZU7qD8/vx3JqhwI7Ht4iv3MjfGRoXIZJnQBvDndKy
T18rUMXYtyX3nVvWH+4Q/ZffRa1QOSQS9a5j9G2+x37XP3DSj3mmpgzXTtZYXwmvXI8cXBmhbEsp
VbPwAPPA5JyE8slBo2okxmNcDu4ffcBm4fSGgh5/Ohb5XIHgnc83y6z9vEbGHojsOE8W8kGswvk9
pO3JYYJmgTUOcvfcSksBsitmXUTZYeA282uWJMrsmj9LUNOBzQp4LH4hUVWCjYlmlWIIEtaGv+tL
scT5YQeOw5MrWlrLJ36iRMhdxu//QsIVyGhoxypYv3hFIEF+DHxVXkmbWCenwigbWxqKNYGomBwW
yHoFtkRwhjQ/i879j3cmeL4blDom9xsduWN1V9W5tGX2jTPvfqTRsj1mHpWLWvzPkwjmlB8rQime
HdV/tszWxabQzX48yz3OpX/b4SBJF2WoWcH8CF8x77eql6HRS4D4Jh5Zhql0JG5WdzIy1kOw3xdX
bNbSfMbWzLS4N70sX6Vwe4jVwNW5yCXtrK0jooYAi8EeBH5uDsUZNiQ3hlOqHuoYKhw7fxufztxj
kOiGtGrtZsl85ZFVw9/J5qpLJ6fOqnahTMNazU2ypXaZlGb3/FSWUdlsgqCOB/RXBH/xYo8PwjCB
gbjDNaHg5udf9XGN2JqklT8zG1zU+sp5XeXd/m4gngQZDHC+B1EfgKx1mPXCRk8qODq+h7lmaAq6
eSk3lJ6AshAuTjbwZpZjld2cvMS57pn7Zd/SSBw2Trr9CgYI1uwJ7Ver192xRSxWs7MUbfckGAAV
CQLt9uTcw2rjGw/BIoXJ99jugAFHnn04KrHtADWvbMtabR9sGgA4wxCCBTaJI81/9OGIIO0EIZXo
dEizZS1/DzPP1lwFXnjYtUezUdp7E2J8M6aHg2XKWV1M8msEe7zwN4Ne3y32sWqCubn8b2FNZB49
BekbjWq/7QEM7thThNE1Ycn5MKzdS1sCUVjTWO/lLZUFwaSgSKIu+SC/PlnAki8CeHl5v+9VP4a3
gcojzCmiPE8rPa1H5XZu1YS1BZptDHBDUUmrqNR6QjLHw801Er8TyiJ4cb4TfZWOK/gBrV7H3SdO
8yduEzrr6TL4aU9lq1gPqTF3qJDRiMf5NR5J+HjwxF/XtDOsr6JF29QNkO9QqYoIaJPBu+Q91Exv
2qiG64B+fB3a15E/9kdzt5/M9yi1Dcy/HOYcrEWct1T1MAPgYWayMz6gnrXIBL5oBkSzNpKyVLdR
J4gE8zWH4ED4o3IPHddajL6NW8lZBfSI4kezIcnFVsRZsMCH5Ct7+5O2L95YuggiC471Wr6uHyDh
+UGaqSfjtZWn6jw0Mlo7BSarlIlSfdDC+NzVX8gxPegL1oNONm5XhbGlG5VFTseTMreKc8j87UHs
nW2RDxhYxMAJr6H2Ld0J1XxqqYwX3ejXgTozOdCrqSGkz6zYMV1eHxlPLHTmFiMlcegOZjlLI4gr
koMMHcD4T3+z3vRC0TwOM6WG6pmFxm7jI3Sp1X5ddK+S9CD7KDJ1Ck3iGzDi7zDX7RQ47Qd05BPP
9Q+pFmVoFTIzpEaqq3mUehaWuaZWHI5RH1URG3vKUAHz2tpauFYInnFldC2w0dZ68xQfgVOn85JB
NWphfdF97bY3Sw5VIchj5igsdn7bfxfLfos+gJRTAh4pNWym5WLcXTmA6B8KUo79vgSwS2ibpNPS
/v6/GzXC1S1AiEf4nq68O4cmiUj8a/MvhugRfsf58dlDiN8XdtxztoPUFKd7b/2CkXPt3A3GfNvE
buQLUgq/MwdbYUtd/wTUJ+YY0WkebZ7H1cfMXgwXQw5pWqVvxoiVYg9CyGO6YTi9iwahgI5sKMfe
wYzbfXhxVGibj/n1xoYobboLR/cu6zwZCz5k8rh5U7E+ICLb9QOSx8Qf6mdMfkvv+QBpOQE8Uxtx
NFiR2g71ISTcFSgd/2t7yqgXuSAyIYv/mUOcZFGBe8GaFOcGeJ35qnt5GcJZn8J6wpa+Gp+FO6Pe
B9+/GlfiKXKP2tWKtIykTOejR7/JKSyLchwxx6T1XS2P2QoZLOoNOmzp0aw2/AJFAAohYcAsUeoT
9Wy69R6PqhXWG8plHkpeFuXX72Cl4p7PD+So7pFR0glFXWx+crJhxH3h30a32uCzZsTKU9wAmgbl
iYlqA6wF2LSFPi3NovXvHQd3OWIW3biK654sOZlcu35aMbuR0aiQ2TBOm1G3/eO7vGfzPh2U+vIQ
HjRw8afBS9AReNLAI5OU55fvfjjn6XIuNqeU7YFsWjuMYRiyVFxgA+H8VwgzvdD9se+Rqk4c6SG6
WIyVyvUROIwCCUkmcvqAibMNI8szduQux7jMIGLtshDRNx2QDR2Qc5Mos/ZqXHvqE6wZC1TS9RY2
wZ9JIeCcJlwpF8R7tCQzLA5eERCUteZr1B5kDV5cvDsXhWn9W027thX97kSrG08w/Qp8WXwl9c6j
neUXWozSJp3Pp+em2ba7I/XLypX3+Uzzi9qpCRHUH57ms7RGvnn4tofxGN7EdUnT6duEnLNPHczk
BwrREQlek0S/xiSWXDcgo05Ch056NYESdY06M/tP4NGg+rsV05m/P8Bf6bvOyx5dKROw5oiRsVuV
xJ6MGk8qquTNqmwYVz3Zow/PtrOUg5yfY8q2GFMqYf2I95Gn5zZ84sDRd5+CqSCcgEUMlEmr6CGC
DtBVr+avCKiMkDrqS+2TNctJaidv0XcfQNzsztoSTJDzqP++YcnOW4HQ5lY6UNxQPoPtkLnFJp0K
88dpd+S3Vd2AUV1cGHhWXDkdbSH7R7zpqrwrvyYIiWuWWtRXBLyMZkDLn4cvFwVUR1a+tKxtVJsE
vTG40HkcH90cODpi4Yoo41YThtXDGWomNX/w5otp8eHo53HyoazHPf2MxeiQZfQQtDOoBEYNd3O2
4jSix0tWCPie/7x+ZOXTBj2MNXifw9xI6WV/ALnSxI2lIkzKGFSc4hgPpbjaycNGSNV6sFLwbBo5
pE79mTb5PtchDzua9Oa7Eb00LzYlUK4n95WADIlaF+wBiRQt4lHIyvT8acrGeAICjHcRaIxtahcV
OSXbSVZW3J0YvIPtm4/8ygaGPdVG+q4IzVb/izNukd9deNKrh9yfYszLfqBxSV7cn20W4ZTCOkDA
Q5RQRbwdjkf16EsHfWHQbEf1JgQ1Xj9IUUx01NtjB6YkPN+RgA3EWG3WrcSvd9WtgMq8qgMhlMtZ
nd50JTxuTvXcgKoQzg7SMOzOaV25s6Ht1+jV0GhV0SUxSD9Jue3zDOhjv1CsTF3A5NERjHbSNMvV
G1hsrTkO042DdSXUvfVq6tTGAhdTlP2Keg2gCntMRs1lhAyrc8WbjTKSnPFr6CCMdjcQUofVdgxD
2clO907yLUsC+CeC6MZjYkoHCUgsP1wJyMTAEqXaDrTd1q2nfpW1SERfPBVDyNR/DOSLO8I/u9Pr
421RsLANZBZpgZJeca9a+ym0+vW6I79KCbMiWcRPoG9L3cX9v/rXQYeR+F/zPLUB9lp9AA5z6z7H
LgC3sziNRAc7daQJ5GHCOSMnN3dlMoMsapmxwhw2szUox6L+fbrOLI7MPzDbAYx3eS4iBGDSkzdS
sT6usfswWdWweYVEANM9eRJAV9VtqrlOuqn0XhmbB7AU2HTM53syI7+gPa2HHqKiiy0zlLTbTj0b
jvX8iCqrdUlv8giXkfeSsxKZaz54YCUqh3sV9W+XgwnjCFFUdUAWBUqhQg0Enj+8TBgb0AYVrD2F
BYPAjUNSi/5KwCPkC0h58UnyuGTOVOKat/STtYlrN2gBqArPSe9OActVyQIGFB47915tonITg4qu
1RTRgARMbglbWoeB90OV6ARVUV/TSWzDevmp8SeRmspuUM+WxZAwEBguC3Ez4yWubKS55+kpRB4H
vLB5s2LRmyRqPeZPsnItYDVzUfMx7uM7ITrq8QxzTq/oTFcqFqRpBu3vj9bnrx/f7lMkCo5h4LaW
G8D7BdsrcsqxcG2/Bf4S9ft6rNhVq+akGiHlmJR5FnQ0eH5cW3Gpvc4cnFE4abnuFW487LR5xx22
ayVzpTjkuu3UQZT++P9RxwJpGFqKbh2FD4JKX/HJBppo3ZUwqGtSkhs1sroYmpPexntTDWn0xB8R
ZlVcVacW0WUvGJQHTFCkf1L1cxV5CuiaunzpvNjQeJ89C9g0H1u6phyjIaa6qxSKeSSFMNEffwfi
kUxcuXht9D7MJ0ZDPBTIHmXsHqdgR499c4igsIoKcQL28qB5uqMntVHmUh6kzDfsvd8MQDkYAWK0
Ni751wmKkR2aIvkKxEj4kLgNSZ9PVh0Tonad988+Z0SIp04FOO+Q5vmRxoTyaTENKH7wVsclTUwQ
CUumrPoh11TQgXx31zW/k7ALjYKMCjBamqxvpyIRsnolvlGNJnvg2au2oVZFJijSvzXh31jg8RVJ
TdmoaXg2PghvVfcTj2TUxejENu+7kAIayIcta7cQZ9ro8bVbACNYx93IZu+/pDA1WWPSTspVptyq
4M1lKBsqmpZDA14lpXoeVuJ5l4DdlkxwNIpYz3Kgyq4GAaoIxt3tO9r7iVPNsG+/eB1bUMKtS8KJ
VW4b1Vt0+0u4ZMrIeS0onmsGpT+/EE1SEMmM2Kach8pqDs7RPNKTeJgDxnIE0/3RJBJggBfBk8TJ
swA+u9sq7FjmB65xlv3dE03GkQ9cZc17EIUPhR1nfBbuxasWXASvJ/k/eF+L6AGbcSAsWJsNaI3P
SmWzunQUkdH4EcDNXFJNIxul5D+7obfpAW9iM3dhUrnq369wYJqJv5ZiJNcaUbuUv2rdUjMLNdLE
2xgQ4XroqBLmguOQOr0Bi4ySOx0Esn3+CTDCifQXw82w1iW2yAWSZhZKeY/IekVi1glUakyoZSJN
UM/i02J+kMITcIWpmYO0gpn1Q6/Otpfpa7M7jjrY4KACq0n7jLmm76NwYmlaR4I9GpnmPBhXMAxc
YHm3VuVnsNqRMJATwN1+iVaVgAyy+EmJX+Higr4P6THIPOiCcbKqW7ggLfLjCGpuvei3kbSSZBTd
Cfl/yDLjiTB2d7Rh88CEgQv5LHe6a9/xlKwkyNsnaNX/0dBOdUdlRghs687w2dcBuMXfOy1pYpAN
CbkJ5KubxohEL6FzIn/4nZE5TQnzqA0jQdsiXBcLeX++EgHeqiFvaneT6P3KHeY2A3B2S6WTzHSs
vImFwh2DHMF0Dopt4t1Zmmau6SqEuGqfQQjq9PLizdnkk5PtuU8ctk4L96uv4EC7gzMfme5hjLOW
or9Rt5BemRPJcDR3uXmpf/ulZQiuyLhUax/b1yR7r6FbKZsGczi41Ow1wNSV6ZWccOkwM7ASQfwc
qXQVERgEbDxF7Q2lyJGgvdHl8GQiO13ezMvg92jMrcODpojHmj6rdorKCaFPAanAi4LPQcifzbEs
XHuReSBKCTi4QK4TJ86OkLD2ZMBUNWI5x+eBooZTCgn72wFtbkLGKoLDXS3wa+fNN6jK8/A7A7fp
tvMy54QCJr8wqi9qxhbfFRirfgBbHN5yiba/2ejhnrMZ38X9szuX2YdOHCfJuxFsfQqJtNplnIqN
U3ZHwysgdGtQaKPxBnvHK0j0Wr0Vf++ozHF00IG+CNtXYLFUbLUolZpnJFT2PfoXo1AM7v8+gc43
EFhSwKx+E+Z0ZNXdZBkSWW7DHjQh0hpO0pllkGyegP2zY3qExVnHnsaXd7uGRSutXRuLsyTLXnrU
qlgp7blMdYHPi44xoo4wir8ai1UKp6XJ4PF82+e3Eygki7qP/rd5ylzEomKgjzNsLkYZLGFb75Y3
97Q00CIRk8SI0JNgm5ISZJK0xT9MLXmH0SdbZXTgHKquTCH1Nfry1N/f0xq0VJGCLpUBOjS109P8
8WWKt3PxVTwdv4RVIcUcoYtc3zrGzjwqhOiZzAHK6IElJEKsNK2PBLf95XLyv7HwlbEz2Zdpfu0H
dXjN6Yy4/wJiFAEovE08pzXmgnudayeuu/+Yhet9Gf8ycDMUlDIYTObaOVm7PIdghB7YHitGAjgo
Hmy21/EGSf2pqeIPz6yaFKwVMz8xS/sKs2W/GGaESIi2iU00u0pxGoRUx1ND3vAu9IQX/GTvDxrk
c7JBx2WUzkfwlEz6uzlaIr6MzXV6nbhK/wYn5eawiq9RqIHL04BW31waXoUDtlh31ejHkGphx35k
qM8ErlqHi3ZocduFMBcBiAiXdwq36Blu9SFoYxNM9cSQaDQDqCcr/Sph5sER89JbsYaTE55Z81bW
xII0OvnCdMwpVNHZSSG1A47hHDK7vCdURTFPoLKqtbgwjCXYFeh61vIntsncFrALPTO77HJuv+t4
3sFb2GlB2xFeu/IGTS36SNTLVabhIulnDGmWWP+tvhp8QpQ6JgtdrfnIuyCOjoJkQcTAWPlJeANn
zmjSAyEhG9cCsWtmDWPhiUJiyboH1Pje8JhEE6dUzeSLZMmH+slC6gq4Iz4s55fqPbYPMDxsHKdE
yMGjVnV3RlEJ8gH+5GrjmbCyqzj6JGqGgQ17uKBDA3e2uLldMhYVnX3TUoRXLAGXgXzy/wg+rPLr
w6lZzxm7jCm7EfsEGTYjlgl4RatOSNSqb5AC6ea4Mn6fHLxs7SJWfG4vHkmLj39fU0yY0JK9Kl7c
0YcMrzZIuoqWgmD9UGTl3Qt7/FVHj83D5fbUvrU0YGwDou3S3jvru/T8saqg9T23xvAWD6plzNdg
8/miq1NVcQPtd1Veo4OuMxW0moqLgtCfMtrG4APWn9o9RKI8W5YVxls2S/RCEv8zVsP5VgNNJ8OL
N+T6LlDGS29JLo2d6pEzvGzSKraehlH8DYxFUYMfbwjichb5nXiJBlsGBvV+CYvMkbUPtac46Fau
AA9fJ8FF2wwFvb/Puh8S5/uyMJ5jlwxYIU4yzHE+vYD9R24qpRMXdqLBWvg9LwTDaOW3PN4ZJ3v5
19hXqyFLfLUl6w6um7qrQxiEKXfc4NToATX+iM7ij6Che1YfXFaauEh0XjFxI4J0phJfTPrMsKfw
Pyx8epaQKgteGe3IhDnQOvK1JfhoYCNQmLKZDizXsNQXIhtnkua9yybjdH9viG1xy6nuK0AmzpTe
Kiky/GpXn06f5DyHheYzRVbAXjIkbs1lAaLbQyoionMCausW98urz4t2oY2Bar/RZZ8oBW3aYsLy
IOKGqKfchAAw0JeAc9HfsBMButvBVHZ8gXwkRbrkHy6XLRiSoebRELXnldI2f53Hfb+bNCclpnnv
Byt8EagLMoFEhnpeq3i2NZzyS6q9eMTvt8lKZ3fRcZjPw82qV6EZwjF8UyQIDCdlfsTAJZkGRAFY
hHyi7AngcIjK8pQVD7S+OpoG+C74ahwZB7oywWTDACYx/NN70vwEkNcjPwp8anMqGhbRyYcxPNOM
UMGqei7VTzrq1UThvW2LgsPjAWUf68xGSteoTKGO8jKEyc8INBId7X5LfrbEs6aJ3LMwJzQRoHYW
qW6KicvjYLS+XuKuQ54j+bx/7WtNIwGG+gcl3YDpUwSUKYD5hvcwVg+H80BQmQIMpepD4s+q9Vqf
O0xmfK7+oy2Vl0k0ETtVP18Qx9KKmCBeKL9zteMhXn8FVXvvwfOxrNvMXaEb1htjpzSU2AOaZtZe
rw6rS2bPcGArnKaZidS+1rCD7HncYttNMKvymJiHJlmOIY2bYUXWAjVst0hI7llF/3sQf8PFqfD3
HUIR+zMA2aIZ3SEjdxHiDiJF+f2Mvw4484onLku0Mha55gWsQQz4P12Jh3+pzH23xXR8qDwU2jr6
6+4k0gnY8j1zsgrn0JwoIbEprCvf+wD6mNW4BSaEY1OhQx6bEk8YnTPAWYbHGLkQxylHvUFTBKdh
w3OeFkpj2nXBJ+erQGrtaODFxE6WjoUtFGF+lAQ4a69qP+QEeT3orqBliW0/zk4yMcZPvadg9siY
6f4XOKfaCkLQ5B+wfhkDkRW8RbjuhxF/G+AswUvet7CVO/vJEAsI49uGsEquRliYaRiy0xnUJIum
UeR0fLlskcMlrKqwVae8hj+aNsOSc3lIgwiDqrbfLZ2VU2UCPgKGKl4hj+rYPpBaG6t0JcYHa/fi
dNMAtEY7R5Yx21M0aOehuakW8cITN1MMQtR5EP8Qfb7TTO5w/Kk7BEqwHDjN3n2ADrp9Y/38gmpM
H0PT2fsZHtCmq72QA7JbXXERC5bIn+rTAjE+1EYn5T7AA6b/EMTLZblc79ESQx9ukqUNljBpieef
AgX0VlHp3fN/W3spyEfVuKx/KVvQaxda1CzCMCT9SkwiP06QqBOPCnN+qqCdm4PIHF69aErLkiVW
NyRLLaYAnG5ocyaJb5+PtgsoSjovoqoOlyOxIfXdknCqoZfZCfnB5fyajy8nZE3hme+jyxMTgIxn
64qlL1YP7w2tU6xoWgtEOKHnjDyZuBV293q8xrm0mrbZqMRN0QvEn0rNx8kGaQJW0eZzj4Fsz5Lu
v4sSTb/DljQGOXiOPpoCB5m+76IFyGuNsrzOyJ08U0FegRELUVNsFG2ZqaIn17MeZcUx0yqn+IWU
Jh6egso4p7kQsXsSuZFeBvPb55GVh0gSFc/x/OzjmlrQocq2aGj9gDagQ0X+p8iJ2UmcjVIyvN+5
Lp6FCQR72xUZY0aBm9RzzfQw3zzesx4h6MEWq0+29Wk193XS12NswJakU8MjcIIdOZy/FhOd/jhH
JAFVtKe9ewoQGe1YslR+LpKQYWLwS3pTBrUYpzwf55F9+PQX15xcdOSWfY7h8ucPKJe2fNdLRcoy
xMEuY1+Ur5VK1Kf2Aky61ci9YoGqBWIoUpFf5VcpyF8VEiVkOIXfNbGJUXlscY9X7fIA1ttXhm3s
934JOH570NCn2slmh79ZSs4sGH6L9VnR0Vql7ZvDoNiRRxoRyfNPhTlN40kwSM5rx+WXNe7WuUu+
RfgUmGUe+Rtat6mYtIw+7LSZc99/haR3eyYgiPKs+275DtqrKZopbR5Gb0h50fFmonGvLuXsYLUO
T8CDZh4e850zILrcRqugRRFotgvUpz8syuRR/taUzNP+Hul1ubE6QnJ6jRylWexcgjeXcdc3yM4m
HBKETF498x14RPgBrYbJ5QzVcL6olfGFcJiF3HHhTWeYnpwt/DI8BXAgNbWhyty3VtFXupSfUTtg
yhu96HKJp+DhJTSTtN/y+Cpy3tgY4ENqXOGbOht040RoniOvm6euMBK3+bshYRTotLJvLezWlTUW
agSSn/TM46fKbxzNIEkokIm31VS0PtmCWUTYq0+lk+HY2HPBaMtc5TY+twuxk/6va7QaGo1ZzweQ
YNXElW0/eyQJlso+KEWXtb+Iec58gHeU9mhEOsz1ZEE/iS+UCybD/Jm7KTNRzOZZ4nOyXtFMOIZY
aoFopdYpDvymgO+fIx9BYX3o0cmglUsIB5bGaqpcgZsXsnqPInK3hs0H/G5DMvaVYqLqzc6Y86Z/
IUCEbBtfcJO6nMhbo5gziknceqNLK3oF6IRYybyKy/wwb+CsWS2fyH7EBUee30Ne7DpKUjkHbmFZ
of+MG8117WZ+YFYhFnKG1wyscjScO96pG0RRZHZTL7rpwLpwU+ekLRjFyKKJkXeYtuEABZVBvDtz
gd5VvzstX73F6p9pByhGtAr19C4833ACQnONNvpZkUvhqQWNZL1GNJLB0RCjgiRPf/FxE9xVK5fi
qx6G5FpVFPEtz2+ijC5VNuXO4PFUwsPnFc+Xt+fK+T7dqNyzAB5Jywme/VApVsJHxBx+1YDbrKEE
G0IaX5yx43lEblMkTDVXWRt4ckmNIVPHGyFXSz8+5Zcuam9e5t6oMTMUpqMoJX9kSHHj0V15PMXp
NtetUayNUFZmVk3WTaB5XWDq4iGjeCvzZZK+5ybt2UMVuO4fsO78hQyZzJypP2ptJ+RRsP7A3P7C
9+pBl3Ba3i+3L6rei7Noj5tKM2OnhDkF62K/P9Ur1AlbK8Pr4DwN4s9r2qZzZkQgQVCZrJgLHlcS
/sONoRA9jCUWw3DZFWqn2DmQO7xrDtw4MmMlmPnRXzMjzhyua+I0j/pj4Wo8tBfGJkkqCv7V7LJY
V9AulG/vb8QOL75/Vk7Icec3eJsmZpUBnNKKDE/h114veLqdJ7zunhRl7ohPk3w3Zfvu3Jc73+Zc
MLz/wkTc2+iSkCo4X0h+m2fZPhzhb4uMI3gnHPiQN9jK3MytAb5hlWw6fjMvCmneBisa1g0+spQO
/0TE86+09eX822SKr6PPnBcieOdwOlcP0ihhHz5J/jlXmzzsdR8OI/bUhVwQMYzUkViV9zHX8wk2
DP3Gf+5kATFLQPlt7mOMx9NFEpe9Mk8JBuU78cMnoWbasB7RfUxa4M6xEMlvnWtEACETTBQ7MHR4
IcOeEIa6Yk+hEf1kX/Ojn7jyd7wk/MDuN/tMZ356T/I293UfkZFHsCXxIHId+W85K0yVy1ljmgac
Ix+IyzABOw6gGS1mUO8WOHt5cS+yeNHZYac8BhAP9qKDrkHlsDXvZ0zV5czDDutJLC5sVFuv5+iG
HRm9lwwhoU1en+PwqWsJpIdxb/9vfwjOMRmKVy2304XXz5OQvPczGASuqkrpPuKRGnkhqNK7TBfN
XC0A/J6+CXVh6uEbXB7yC/XUhQlpqQpHMIZh+coQsro2Od8tzmS+Kf79KCdG+33p1B2OzZzV09hl
4B5pmWSsZaSPh6j9AZIdQsNkDLvjsjFFvL7igF7zVnnfkwwV+QKIlMdZdRakBHmikGxrg6u7LWzX
Ttde28cm7hp5JVJNv99ngBKABvWXotLnWHOCodDQ/9dGFRne+GLj3mLvgBXcpkfVsZeNJmJrvt3+
QhbwdjoG8vrTf6nxG+3S2/554EIP5v4HW2ta+cOQt74MHiwA61FX9zlQi43BIJu+VPr8O8efKhjO
2Et5edepWAzYlOSNmhFmmiWrd95+J6bFxLYgPlinaonnlHPH8+XgMTK9LRHJwH3TZ/4LIXtksqCR
9uWL9+AUPoU9C292AE7FSM5ES+MLRbyN2SqOscObjSt6h0eTM6nVc4essRFdlz9D+YaooEPIcofm
saSLYBwmxMYDyDfqHIdmXsObC6FHrgoTefPk/y63aBe4xfIXPSvRtFPAWrva3guQJ7CkEmzOf2H8
InmSgaJLciMGB3q3RPXwTnxPaylemvUw1jns4Iuhy41xro/WUQ10b3oN+JTQEywpWRzo/cnh3OMO
eer6IoS05JcPY3ezQK5wKzwzonshGQl2QTqKNQJmulL9u4fTlQ9hlId01+BIMzfOuc4CHPzsFDQc
4PXiQE4pH6s8MXJ06Qb4PRehBPQlu4h0cfVzkGTiuFXVQlOyTh+OX2AFzBQYWdBs8yPRi7LPkuPJ
q3KnAsR77cCzKbdG7E2n+3zqNPXRJg24q8aH7gAuxWudXnMYq9v1WP2GcgcjwJtVF9b70LoGSqfF
ePc9Ca6mIrodasSZpQFQA7XBxG/2aVoxLSshlOYTPqc6EZawzJiU+sJP8FeGdVcDA5/e/FTUH7Vx
1oYusyAzUj0EpYlrWPZTdne9bOcDc+K/de6YzZEUV8vMn7vbWJtgu0NIYWkLlMIrvnRHtIkVKH2X
jViamOkalv1SMzV5PRaf47uHng8bmkSUeG3dEBNfnFhhfP1QCdKzOf4ItqEtcgsFtb7WgatrPDTa
CGjKoigcHne7oc4/n3tRC5ssOU0QDeLTk3qQxRreMMUJ5QHeQphsmhqdu47F3/69RdjSUYcVry36
0qGg5wHeTtuf6SMKR2HnDVghpy+bTMOZi0BSCpvHxS5bM2QfstPT/5leFpqHKlZOLdLEmf/YL4es
PRNnyLZ5olPcDKNt8PX8nOb10a3w+BaMzWbzSfMalvSoGobiySEH7JEYobJYN7PmTgYODyc9Q+PZ
5DkiT254UINfKDLVRuu5rjcdEH8JEkHlUio+KVWhXL43/DSospcyQnDXkxhZCdQ5Jqb1l2qV4dVx
1An/tBqcUdOfqzgPKLM32+I5gbivjWXnzIQCnzk3U6Kw/zFBAcO9pI2IAGOvw9haXCbDmw+viDWU
pBBsRS8VmACWzC87eWzFl7TiA4HjIaU4kF4xpK8gg3dC4p5ZZOIDTqT6sRXv++Z/M0UnQcoiYeCu
iMWhD7OWhYU0f4cLjj7UL7c91aeDDcEy6u1iAorwB+7WZN+g11+aVdkH+mVmnoyE7SZF0lc8JU2D
u+MeCh+0JZ1+NVB+5V673mTm3Z2wCiNeS1Ij52GrBhrhq7qN6OSQfLwRlUsp2yypULff7ZeMw/pp
u14aZ8js7Lutcv0Fgyyc6JSwLbdZeRfJKvCC/3KyLDIwcudCGY0F4j8vJmW6/Ek0bd852qu2sZ00
jJVWWwgL89Eb9Vj5GS3feI1V24WjnzeJfsPbf6//GSh3x6Jb/CCW2rv+8EhKtLof9LTmeq8wqkTO
xq0ABYZjQgbWf5ZdG1ZFlTXR4B+8xu4cthC6FRJ/Tye9kwBzzvzglHizUAbdg4ViqkH0jirskMLU
63eAnrD2XxoGI6b8u2tIugsSnDdq2ovfefU34DpI46I011j2mDce8A+toiT7oWfoNpkmR2lbu6H8
xyLBPNbSS/WhDRlVEYoh8J3O3sYjdsp7UyxdzNTkyy1IeoTh32LVL7dhT4/HjAAw8EF4sTzsEZeK
Kx1itREa216jP0hxUNQILURh4WWCyaepB2ar/ddLAH7ibU6bnWt5znghtNlDXiI8sFMpnv0ZcOKL
vzQ0ZqSARTQLCXSTOU/yJcNSDxTF8cQIBTuOxP5nuPCtR9IHZPLpDuWfoDgX+ZrkNY3tY3W0jAaw
uoS4Wr/6epC4zWJzBswgs0is0KJ3kaHW6MkRCQB2qYU30Unwbb3wQpsMvItD3Tv16w4DsTpXy8s8
Nl+ulwP0YEZ1pkrbrnKbO1LFXU4IywNgw9Jijz8BMrzr2bGx/ddkM9HPzM4XDHft+EJ668WzRXKF
2tKMLQm5wo6Zg0T4W/RAP9HswOpdnPrM6U/v4f1okacBjebAmTv9u+N+4v5kZSwGmOZPPvahqLQ2
fkLuqzQoHYHRM/wxWZJlwYrgLlk9TYUYnI0ugW4Puu8nMm3nC1G+DExbgFm/pp5qUTkD9w1l3+jX
ML1mTQd0QAY6W1ft94uEJXUzl08PQuixIqAF6bqnN2jRMnv9wgTfG0KRZY3fkalQCF4kAnx6cFYq
eqyww5O1TVeOGznnrgYlHrBJm+Ah6j3UTlY39lre4twpMSwP8VkoO8jmKqOLvMkWwtkc0l6YlvdZ
Qpzr6iSgF5dgkl0dTGutTM+Dw0JG5YdI4Lf50PfszX16P9V6ELpzpZG4vJ44flHDpYJTcvjI+0iY
Fmczp12tdYQsX1LLyrP+bivukMvYVc0R/Dw1rSZ1vuzgnQwf4gKSuoAxkij1/cXTSMYXIXBPhufD
IeqgkrVbZmrpuIpmX/eQUdJ1It08jOylADDdK1mCMIF6YKXGtVyBM3tdRyLC9ojAUC59pZrrmy2O
2ZlA9P4mXKLzVEKh/RpYkI/hjOcaYrAKi/PIPudruUYbwB9o+uADtdsVeBxQVIDCjb7H24wFn94k
/xyWBsSzDXL64Td8D+no7WrgDtD4gfgqGSyMTq372+G6OC4Z5T6urobv3KqJTbMKX3laYZGO4ZP0
KgoPx1L19MJQKRBqYoyEsyWdzJtgQ4S2y/AGsFuIWoFmgYRFweYxCtv1O2IevILS6DGo9WccyY3f
s02KeOLQhpOcS3w+l2uXTrlPDAjmqOnD/Ik0Wf6gwXyoU/vzaBQIKAeK8FbBlKEcNzXjEgPnVKAn
LJxTjqPsRB+4ZdFAVmKCZgEWG3oM0noAf4uTnl3kGDlH9MgFSkJtblw/1U0XKyomJdaYKObIEej7
M87oUdi1t0SR/nGUooGtTPe8solqwCXF9FmjIK7IkvBANiPckTV+c595DNNGoD5jIw5Iz7GDOt+2
Ggvu9Z9RZIHpbJm2T6L7DuNZ5H++S4ippc3tyoBqdmCZSJbQy4c8FXoSEU8316mYo7A7DRCc9TGl
nDMEdZRlbdmVJ6oh8RcPDMXXoLCnss6EI3cWYI/493ltPC3IuNpREO2l073ZwFWGunch9fO9b2Gv
epONuWaoVc6vPLuqrwFHm0Usf/ncaGrrmSrnY4ZLzyxbfURHUSvDSGroU5hactws0p9Iw2tDdRUW
aPddkafhGwqPjB9ICMU8XgYTk8bo+O6TptUg6EQqYjxSTa4BSoSjWJghGExEmk1e8MiRNdPSMhJj
tBQDjOL5Qvoy1KsVxymXk7KiGsSFcANxedqjNZPiWc22EGAbhWp2v7fc4715n94RTMYD3iNobkHI
vYBPCsLincim52bqdiHNqQ23azV4CxZNdAiwosDTEzRuxGajZvvrbBgXAy58VAoEju6evUp+esKj
ZEK9roX0T9ZNyWX+YQVs7MFKAqHwUaOmyB4+K0j/wphMGA92zL4DIfCzr5Y4WfxEnbB40Pgkfk3X
Gbm+goY9vYkkEJAW/up+zG3/h9JMt1LF53p9gWhplQiRJ15ogdGrZOGDAaYJwDcRCNijwi7B34L7
xBOCdizLqhS6mFSgMqow5YfX9TwLse+Sc+Qp7+DY1w1V3YiJvraotWpE0r7YQZNLdNK6fSdQREDx
ubeUKo3UoNyIIivbPhzhnd8SoVmxilZbGKlWzAYxziQAsgUDhJ9U0zQ8+x91rNDx4Zq/VP4Qi7FZ
cl5Jqb2RIG0CsH2TNpBuyoItfeKboLwUrisEt21GN3yzBOtmthAOjFCLj0EG4VJZXExut4WHQ6Gs
fao9+8zWNtl+qHSuSUuVGUgbH1lg3tk1O437BDF4W0E7xD9+qK8L508IG1b8YZ3/WljgPdhVvdpi
Ni32O6yyloFBBelJ9nuqqkqLsSfAUvoujDiS4Y3g27WQsFr98t+LOJx8q2zjWRyupIbCenuI8yX9
lLNNgOxwFlEbhDmHz+yrBPLZoTEv0zWv5CSZO+wGd5i+U342rjPu5wibf+kZohpcK/Vzv3paPk35
draC19TA7wYAulivzTHJRvynH7ec1UJJklXtcI2EIkeIL9aCASJr2Xj9Ai2mJbVzDCv4kdDjfvbd
7+F0tb++Hb6aiIjmFzgG4iYudQ/xz4iHVznJ1kXIiH1JoEBpesvocd3JNtfsooZkt7EeCsYq/5L1
gMpX7wlunFoRc7+IqM2x7S2H6V557DjwHaqP4ZVEc/uuHHVKYgFKX+2AUAhMcx/uh8X7sy3X9IsF
f7/Uj9Nineyy1zjlNW6p7M6lHQ0aSCxRTNOE7o3auySOy8uixRosPWfmgrX8DqcH08gIzdH2yGyo
2qK1AwZuW8Ni1jYmqXcx3rxDMLjwbIPNrwY5Bpay/i3c1QD4H/PKtiL17/tVY3qkPj3VOCK0t0p4
xgkkZraCHq3h05BAL1hvrqGqiGROe7wZ2Cw9ZuJ8y+2gFgOgfOuS/xjkevOY+1n1dxhbkW+emSgm
35iT+0UmV54x6h87ZuPzBxEUqeeuQzLaegZctjLAQxNNj2Szb/DbUE8hk5KkR9HAQ4pchLVfliOh
NRD+Znqi+saEfSy7k+ZuQ7gnTYFEUQcD6lCf06xefCn3qkoJrbh1Q0QGZ9nYopFqS631gbnM1ukP
DjF2IGB7hrR+yPJj26gPj3HaDgzUQGl3J8Oa2dM49XHmLnGTmHTzy1XTlU/I/e2I0pgO0W2x0qT9
JwRBzIz/rYMnsX8QVu0BqyfGQalTQDpHN6fQXgRuQ65s/q/jlfJuzR3XtrNhpH5GKe/Z4Q6GpDcI
p8Mpy/YwjR7lwnhlloKX6Lx0bt6AQxOr+nIDfdCTe1LM9m1yG94AnazcXIscZ0BLi4vlGOI4JnoF
npQIyaJv9Vg+AREU5DhC/Bzt0WYDXTwjYWZdR8PEqRU9aovEa/hcHfAKVcYKzLNjmsY0FdLFCVHT
ZV3suZLU7+zZa6w4BGG9DX2Z3cgsY/p9Y5vbHOQFheoSvwdPjGE568TakuCW7fRTV+o5JpoV7zri
c77yFayADKAu3H+Yd1eBc21gfYcWsvoq61jNQXbMjA2O+0Kq4IKa+t848xt2mElC54yH8mXUQbyF
F/2oSHmf8MlYvZ5wWoytC3s1/eF2WH8idpphrd0U0KblMza5ngl81TiLTBWyKF4bAFqrI/GrAk7q
zdlZkn5WYeXd8Pnzn+z6tyc/umUsxIJ5Rhh48YHrjvp4uJNdPa540Uw2wK3KM9SIOu1vGGpV1iW4
e61jBHTgHdOqVRyuWF2kw1mOX2CiUjcawQ5uYoREGdet02C6MRMnezPzpT+fdVnU44dxCfSd+2k+
V42chNn/wsBx3MT71rk6GQ+t7b24ogDuljYkL3EWsIdIAFY0nmXjFXjNrull0M3IOv9Lnjbbazlw
0Ns9VDZNmNSPnZ0c89Teu3RtB9DjOgt/gphhYbufULCNcMsk4ht4VAUyY0mcThAjhMj/1/AlBBhH
hr8zkhez0eEYJIQJhoFdvgf504gn8BJ87aJ4rjmFZMnYTPZeGVoi44b3tAPcpxOnjGz+NB4w/MWg
A3nzV9cQG83kFbrJrNnSJCuIvS4iMaE+fe6uKm2a62zLCydL00WcnrMMTDQi3ndx7SvCOhEgmVEV
f6kJg+T5ZM9gnhSGA97M7iRBfRGNdZX1SFondhakhF7/XUtL9Rupej9ETylU0e5owIx/vq5kYiuc
YTYSPgiW/s3PGyZ8p/ILSAPJO43t7FnhNEyPL1PRTzHshCS3QIqFwpFOm4mZLKK5SSnmrQYJ81u8
3/qTt1qdjhshTe7hWGDWzScwfSPY2ZHPnFQqXfiXgHn87uQYmI+VR0wujo79321Oht67BxjBYkJz
6AIqC8yD95iVQRT1F6yVlJF2SyPoXVw/ecFmrHvHQE1Jqn+1Futbf3TgV4kr3XJdhv9DCkmt1BMs
FnFu6ldaiahw5hCw0UTr3HLLLuyBSuqF1Z1qelKanWn5mA67TNtzUbzKxCmqpvVwKfoBw5gzg1Nf
KdBEAtNSYjMFHQMZdwhO11ppIlHFW7lXT3h29hV8RqL0cAKms/MlwU8/FdZQ28K0BSbaXcrTDMVw
RhjhXTYkfK+Ot1r2qFQyiGDUA23DrMqsaqu2cDdHY2UeV9G0Lwug/Ck6EQ7I5l2N11SKhUQwSvb0
5wcA1Ku/XWs5acULtnUobL8hQQWxOMneROaXL3FjT2I5rWF6QjhUJCV5ECudl1jmVxhaGlZ6H9Fm
G4bchg6CT3ss3TifSfFXnG50hVE0b51zV8+hVzRz8wuEkuRp+uKX3cRG/GI9Rcz5U6jpOdG3Ef81
jA67A3wCt7G+UuwQwiFwbLvoHwGMNtTe6DJXOZqzSw7LXsx7My/XwAVbbfdEwPn/tRQpajJdxub4
xnhsLAkD5ngT0AIKczpCLOI3GD3J76S1tFc4c7qTAGeJcvnSFvh7JTy8e1VBUTZxuwyePmCzFXeg
1VS54T5+K9g+I7Vuj9/OiIL2zvfLGj6CRQH8MlWlS3YUt/U3H6fa6tltvJAE5CAI5s796AgzNpQ1
5ILKUMYbCeCN/f6mlseDGj62toTwMbWEPXJpdwkd0r6jWmxMCwl6iyGBP8LWyvb9m92Faz6LUeof
0NQm+XhdiNpZWXstUK8hXceZaOwvvxgeswU03a1NLFkWEQblhDNzmxMDrI9P8kvEvh9b9SZykyMX
ADBVM3VN8lWypU6ISq78/op05u58gFkKMvV56gF7tRVxsJML2zWlXesle+kaxzcAGo+v4IBvODBD
9VUFDC+IJ1Lx6hIf/CfgM8dB+WW4fkn36L5Fsa8KRLIi/bDQQSgfzfViK5geHeNdQF65unF54ZHo
DZVfFT9bSlwbNcUc0tLF2ZUtkyPgPHaKYZZtcwYzGoTF61jy0WIs/IcpJnZ8xHBovBaysSstub8p
ZE9TIT1xky9Z3Lu0WG3fMvlVGDD2uZShw4Yfc98f43WTEc8ofujBKt2ZA6eCM/8XhZH/byievH84
oEJZfbnWMx4126QaOZu8vGY8sumMpXXwHhMeSacnuFenvJbmZVEjbsqB7ck73ySF8Lvr7ru5JuWS
Wcdj4g6acjhqHb5OJgK+fJ9iAjDndwY2mTd0gm5kYrinQpEiMExzrOoRkIQchDD8kP9zCQ60qq8u
PegWNMvpKNwufQnMzEWjF/dGG+CgkLO7TBqE9XzSeCaRiFCIW70QTitTx4iN5xVcTpooD5Tk5HZu
awZmxCzixJXHMBM+Ivy7XSA9YJk6di8zEyulKiAIbwvK4pc2vwaJ+20Xyj1BFt4AyNxidI4C9Dnk
I0GxEBt261cKfFricGtrz03Ra2y7vo6M85AAPP5JaJ9RQ2N7nlb83QWg4tuZZFUHk7SqT4qsxn5+
8e1NGS8B7u/jtZgPF/pSyoEE5MypwJ4FISrKZv8j+PqVgzWz1YY+2GII6TbKQlpQCVTiE0WSCKqa
60PfOc6hU9z/mmLMCyBab/tQQADu6Y2Ic6QcHoJo4ovaL9aRSK9IvaAEexUMayXYnulbWgn9TOCb
rpWqqGdtSjvLJqfdCuKI5m1NZz4LwVFURVoLhryy+iJ4Z9ggb6jYl8CAkTgEVKJ5afdUuK5+d9C1
ylW+qRILGfMbj7uy8VpQkePghdQfODoltFRCbr3IK9+awoW6oGkYZd136Ylma6pHvx0TjBuFetXv
QK4hmwPBakvRzeEwmrXA4gERZXAfgNfqtQpHk/8IPb3yPBfOhETz06VG7xr09C4U43+xQ5Y8j7Zm
aFKJsCILh4qmUnc6TQHj3agR57Y5gBECd1o2A5ffDgJPxEiyZQ9c575QKzQfa3Th6MdkscsDQ6y1
rmsrMWtW+DEJHIGXL2wAA5iZZwvP30Cy3ywNgcjgFqQyCEwawVhOG9JP+ns3yen2jsQUO6SYR0oT
iP9Rr39zyYuE/R4GITZIHk7ZALxX3MZezpbr18dOHuiME89woumg9XtZFLvt6DMbXaiyA3UQFSQB
qMcphoWENM3xHsJb0p+UDS6/myD5GkEnHWPQR86aKr3UZ86N4t5wsygXT132INmzuP5ZPUZFCs8f
QJH9d83WKzUrH6gNV3gxfSeSkMMgRW+oRKqPOlUwu27NKAo5SgafjIy54+KVfrb8KSQEOYKYyJFn
N6Pb4IMgJ/5B6k5cqI+sWT9phAulkHXv+zFvHfrl4WcqhBoZuik/k6zyA1PmGe4lJTWvGAhl8kI+
wt4Gj9fvyxdpUpwG/o5yBQBNwveQtfKSUGfgSM9QaublaU7Cj13MQqmlLSxHZGg4h0i296uRpALN
gKhd72/QZx32K0HZKbYyofANqw20C/ZZUHl9gl1wgMz09+9RyDNfa4RxTQqPbfNL3UZBFPXAVFnz
SWk/2sOH5R8jv55+2SLy1rilk9GnG+FtFBsQqV9zTj3iUDxWwlqqKZVp0efhGrYsY+iv6sH4Di7G
rAjKLfS+pGF9PU3NMYDAUfyCIaO9NYbRImCB+k0KLRP37HCOT1Hvi5/Y0zPOXMUQCe3otandcDdw
BndEjst2jB5xrqT25ivHE3rewPcNoL6GlmTk+7cZpRgkcdwFK3UJi5k+yQ7+peQGO9KA5wUh8xQr
oE/Tkegoujeg/9jDikQB3GNCBvmtFMQJvSjWjSGXVCbQJcxS2SfOXsRKyparNW7UVrMv05ZhwZaa
xfPYPgQzH9y3IpI84IsBUARajdsjCtlPdJkxgn5Auudx01uXiy8TAEn8xH+RSTy/BQ6U1tTxQc/h
KFt7s79FSAqXUNNpED7iAMXFJl91eflA6NOWnMXA97cLoXYZF05VCXQat9QxtK+Wwom5lgXV1ls7
WEeh5e0PM+deVrMSA59x0xGswc3tinBgYRikuMXG0LwtvOMJ2Mm1XmUDemSDiwkpbwoQVWxRZYQa
lMk4czjDgUR7SHb8icKp/ubJxmfhHt1ckrcDW+0r3dhFfu99qNKf8p18PeLF3X0ICvrpw05Sv2lS
URDQf97fu5ZPcDyJ43KISA39SnJJUeUN7yA5gfTPKS6QO/yXLZF/ZgTpo5Bwn+P7Wir3Qg6gLEmJ
TtVl4SeZNz5PpdLIqtfwKdcGV0vqUEu5JD13gXux/Jtw/OlaM1gf0WCssgbZGw9d+hmCl9qkKo0h
CtlB7P9W8h/mASs29nnTHXqRkp3wr5kH6BnnlVczEs5ZywkDlFsDjWC2p1mO9lnWV6ZVLG4qRW+C
TI+Anb93+77x14rWV5lK28PEun0TC0D6s9LSMQThouT/jkKD6mEsb1GqZWNSUfN8kVbuYzjrM0NW
gNK7KasG0BE2KCvwvOLv5LmRFfYT/OaQthRzLcgjGtA68LReU5bqTVa/UACr15oWy6KQL2Cgjx0m
IajmZryoqmT3VlMgubXAazCa55uixy5PNBVj2Fm/Hpdo5QTZD3rZcJBqwGX7ZfA6AltdGU7Qhncm
0tLlZhtPtzggUipmP7v1jcC2OD4XzeVI394Yehh9eIyHXatuuUnhBSmDJnk9jsjCH1A8Ff/JYUuI
xswz3ySPICrnuaaBYiguvWzJ+VVmcTEB1T8BWFSAfyJJsDQAjjrskHPg2D6CfQe7K+Y32ZV3jzEA
08GqFaaKrkW/8Lrb3oRWK4/zkCuzRN9RohjK4A2tfTAaXyMk00hAiIgi1WWyOfDwYIW19UvAZ8aO
xyF7JLOEvdqXRxlmhqC4e/5RgJz/ry+aHki1eprLga+ixifWgvPP90Sz4oYQXPdpzfEL24H6kfIo
aMTqayimcZJaOckRLIXdXoEWkcN1bRFndX9h3JHpeJTe1cpUoLlLP83Ncmz8hzYL4oHOkVCVVyEI
ZWZ2KFlpML6h7R30+dpt35AfY4SLmDjd7vl02kx41XpZtp6aW6p822T/pWsY4VJ0UZYdJ3WGrzjq
2Kw1L2/pQ/Ax8mLaQXPxyGb+y04aPiMY+5Ou1y9Gv/HORuhuRW6MQSt3S3dl1m3EAgEefHWxkiKl
kkUh01GOz7Et4nuseX76/qHzuxNzwF/3++97dBd1/+hWJ/o22iPCFyBmdF32A6SR1rNtbCkUA8If
k3FoMKhhkj3cZL+lIKGmx2niag51YQsNMBI8ANk3Ux/A0JJGjfeQwdA4grzYRRT1z1f4uT0kZcCW
rByPweK3cF1lrEpovFnzGG+qLz1+jXVkxS7cD8UFVzMlw7E+VrSV/EFwGOYZoHyMKK2pEJxReIQi
MfjiljrECOT3KF7WQOwdSy5jvgMKsdig9LT1ojBn5z6Pq+y3iqfm1jsyidurCWCVvEhmeWoMsbHR
95eRujCDfaDyrvLkdU+mplnOOF8bDZ9Ui3WbavH6U0vFQE3bxm8tMKUtpfcPiwnIPDaXAwEQrm3z
l9dFT4tWf8gJKLvSFC1BwZkWCjg1jEABGHdDPLBIENkb7KTYFNYL/nUnRQeKoYWBSzW9LWFb6n0W
WXQkqICQsay8Lhl3exlHrw5MSNoW72yio/ilOL8EnY3tO5RpiKSsFtSbB5F+kK6DIH69McMBHw4a
ycW5fv3nhIIjuCDA046JUMWyHVF3eJ8iQ4KhJvEJiXC6jDvC7+Cm42QTqcwzYV0NYxggaxUafjA4
LU9QghzlmkgM3W+XytcT/Bofq0vUauxmiUTXW9417jZu0r3nfcyJjXrggfBo2K1zk2p4Hsev5EDy
TFtWQT0mv2ILtxVuepVzfnArNlX+Xqln+40iP8ISeKec2VpQQV7j2l4oE8vI8aR9vpKFM+iLaxUA
XiCOdP2Ak+t9wkHcR1m9ZnwPR/Bcla9aV0elBwmjRa8UCwqHXJ7P/NK06AAjYBl3p64+8C2le9Zj
G5WUhlHBcCS1XLdihMPafn94X+UCExJM6lVWjkB0w++O3hKFp5dT8MPe3ulWWGgAYsoPJMAbERHf
AQk24LSz9bE/mpkATyPvXd4xWh+hCDw2XUKApnh+PU7BjSEpt4NwuciTdsylrM8e67/wbGVAQRKw
5qgLnNhRCz8eNr4WNFjKfPz2391j6jcAaVrt8oOBaIckZqloiq5CFJech+sh0XykPHOYd/exVwIN
6EvVpmYaptPrr9MB4FxwiOT/WwMd9xGxSLd4YrP64PpeZHoytHA6anBxo3YulhZCwfefA6tQqcRs
fEM5Hf5V4i3RuqndV5lpwkfPcXUUi6FX5UuAroNLRiRnD29tKC1NgGtaZPb4O6luCT0oiU90vJmd
zeGwfTzoeNAX5fGe3EyBnA9YtF3obW/t9xw9nTATkuW5BiLz2Lrk9lLNezZZp88mI+ZcWKqv4AA6
LdgyMMLqU/E0rnWhHlZ9lOvUAQTQm3KiIi4fQT5ElGt9t91cfAtgVoxfKCZzfhQF9Z895qAMUZEk
mTfk0LrxRvzyOkjRT8ZPdtnENj+GYuy+iTnekGgmX1i4LlBt9Q0xTfVsKEpaIymUdj9Qy6ru7WDn
5PsnBb9vGGq5eMYGz9Sx+COj3eI2Ok21vy+AZCgLQZULqS41aZTrLDbjYLzt4ki9H+3c3hlruY1Y
QfEhJVIqTe1e30/IMFUVQmyHd9ZhBTgk8i5geHwRySPFshP7We6UXK3HDSCqL+l2N/kHnTkCYLNP
HxIADtn05Zj0BtYpIannehPUBTftPU3O18SJZo6QRLZMabrWUFu3XliYtRkEmsR8zsyL4ozNQYLl
t+nVO42rDsYh0390VkARr9knF1Du4CkuH0VqlP5CLPfonzFquAGAzCuBhWIpXAqTX0Fr4bFVkx8z
6bbcEbp9p//RevhkS4+I7XWkc1gnBl+tbKTSMtpphZQK98AlT3guQi2E5t5llwthuBlsFS1+5OWB
lYpBgww/920+9pELeOB7bCg5oMAvFt5Xndpy0JsP17bvSVSsu7svneQW24eK9sNwejiFSkog0m7z
eveLvmy92PAY0vwQ8rWYgNhSPhqc1K9j+ZtYV/9dbToOHV5omUgSPdUxG/Lx6Woy1Gfla+6mD5yG
/yS4pGz1lzAoHzmGC2Adx4olJNWD4i80eS0uDIJ1lUgmUYzVgfFujljrtUailpbTEVnJsTVmdXk6
5mgI2kHvDBt9KieQI8WriLlJfvuz9tw2cNuiz1TZOiUIvOmn4YMBQsTSa61XngTf+bCpBqRizhuv
wtb2gHMDQzvTC5uc1vvFkAw0Ef595EO8TIFc14E8xWaJqxTenyc6pK0KzZmMXGD8qBlO82HcTsN8
1W+MIPCu7i5c2UyNhkQVXnVe40FZr+FtAgByyqFf288KBpTzKbC1IFXjfelaFlG2ZcD4WKtWJ50B
RCnx2KIgwIlv8SaCZLKG4e5mlLUbLEyNSF426goKz1Fur7QZo9lhvoGVePhiCtV6q0ZMiiVRLJ0t
rtN+PKrUjixbWb1iY51SgcDCOyQ4hkhZQk0493tB/oRDlkLGlg42TWjx6/Emcq7Oxu6YDmM8JYgL
lH+1k6fpQz17SNmRFvPA9+4hgxkaKbj3QkVp2moiY/3QXw8tl6Z+aOZKfMR3qBkAhfcTVUBIgbHR
4nd6KsOXPevmpCCJ3yHr+YiuVxmx4QIh144CmiXdaI0OmRMdbz/Km/RDskaFPZrluSPRkmsP8XEy
g77C16h+a1H+xGNmqlWenYcSedzLfxXPhNwSalgo/pShu5+a902f1k/oeuP4nW2yHDFJkUjWOaVm
PzRS6uplN+gRidiTXZ82rInDjLDfalsC7lypvCj1uxipFM1RtyfPo+fI6w1Oqyla3v5f/XonE/6P
VjRUzV1tfeO/5O+b3Y6az/Z5jeCYuTNyQK/Us5efnau9CN0wlsk9ivi1u8z5r7eWCa7WMykrG4ey
Ehm87ylG4MB3ry21088/r9roLq5hVFnS955CN5SzV2kLsc2J/z2Tl0Bzl1U/YoN1USbYr5xrCQBD
inF0tr8UUjWNL+CZ9ouTD8BwCmb1jm/JMCncJfVKwROBvKzOJrhz0T9w4qW9145RQJZni9vTRMqA
Sy/JbdWqj1NZB38tSTCGVKXJmoJa+STHcUyVP/0Q8XfiH2h7XBm6I57EQAAeLuNIdbrqyCxPhU9n
FF3AA+7XGPL837uQXR+3vjdj5VcKSeIJez+hYIlcqaPMDkdigvqBhyHMPA6Lgm1JEU8CtHR6rSBH
RISHJ6wF6gVVhWPI4ra9J/2GRMh/e6DErkL1t5zG65LQXNZUPu1Jf9yuSYPbmmssCKdnEbbPuRsX
cv1zLpmtylmjcBxIXT/Xeks3sQTQ6rGoJrB2slnaA29+0dMR7QAAt4JcOAe6qK9E2yS7UUGz8QGD
D4OMAJBwCMpepbwkZBCrQ3USAYUqyWsvtF45HAGxP96y7WHVRBghKE1ZR42TZ9W/qaPHVae7GSix
kK+U2Da3RtcMDpSmVFIDf6ndIc6my6U0cO3ltTEdoXvGMs77BgadB8fYgQ9taKiZ2CpZJAA7zz0U
T4zRX2tbiJyvz+GqcV1MG/WIqTHmkifSJK/iABQ0Rurx374d+WL8EZFph1EG+yf/k47hbYHsYmWQ
1mkQePrat7lc2RIg4Ce001vORSJUHelokq3B6St9n0BtEFXuq7vxhYTTVFJU8NtkytaC1qh4FNZ8
n2fKb1MUNHvI7IQjhh2b1Ztnvgd31fVJ6LGjg1tZ2nB00Vpgc0uPLbqPphfhwui5BtWgCm3cRuQG
353fvda8ww8XoWmR2x3WSVBog2CpfINEM8ZigbsJkbPtNY7Uv/jMFtQ+9+vzoflJVnnDMjPWo5c3
k1qOgg2r3+/wOM3bjHwBN8HqN5mCmZEmX0Ij6oAoN8VeL6SCrqbPVqXdaXDkdL3B1Fpj286+gu2J
qx6F+l24zNeLbFxuEu3xfEuyoOYjkkaZHgoYloLeA6HuJSYF+mOYqlWelss3XiAqJdY+oL3Rm6Qg
c87ICkckmlmCjfXbVP9iMugqxp/7IxdcjjYuHUj9nNfZ3Cyx2t8Aviw/UzAHGCKotlJ8MdVe7f6E
0Y0qpRC0hCHsITYNGRRLaCgAJw/iSbyGTSoQ2M36cP21++qYWqFMF7l/zDhsIKCzQGl9pA1nNFD2
2XXmQt/8AU22ZqZsGIkT3opiskpf8U6/3sLewqYwjCY5so8PUeM9FrO2ZKBP1x2sXHcM6LKfkOOx
ETbNcK2OAthsde03gMfDwSm71GyHCAU8xc29muutxU1ayFDKGrL6Tgz+KTP4EnnmsTDv5l0zPBKI
Dln/MA0Jkw4YnJ1CcnFbYraddJClnNR1tqK7EdrxeToiQDsbH50onpuxSoHjFtLxp3HiZyAAHCZY
y8lG14JFex9yXraSP+YZVVf7SQGEvLMfdNp92dHS+2ugqUGSojv/vCGbaPEZV5T1aaqwLJZ/jW2V
EVdXqXEMPyglSwAPYn2uiBnEil31ZZtW450owz3peGe/KDzTLuio02jHUofEDpFYAB3R2WUppq9v
2xYDdT/Fea/JU0ATviZSFoa8/e4+GxWiDFJbPyx7DqITb8LHmKuwCgFwEZRAQ3pvReNKcGgzBKKa
G0ILVZlzJT1zYrZtw4MkWg/mhtMZdFf5tHfsadnntY5VFnTHli71fXNdT+Iu/9f8sG/4cdzcC/e6
L8+mUExgbcW38dqLb1mkFlFSRq+pH5ngmp6Pkws+koUb6iTUPjY0tA/aXEHaB5/DDZKIDQanF3/3
E6yCU6fsVvozbzbzVquTVy9024ulCXibwmmvZC3rYZo78Fb6fKDyKH6tLYQOxMGcMR0O9BwnPkUQ
wBE74wUjxHayKMKzwnSO61CkNc+0UtmU1fqLS0Ml/yQfoDKeHOiREchrbi0iAV39WClMbVUTnZXs
rDxGbNiD5itnSeGnYHVSiZ7PUkvmLoO/F8ay3mp2gzK20kF3gebOF4kiRKRPHuRil4yQYROELsty
tG1FU6qKj4G3uK0CFtiBdndE5LVOxGjMClqXaFojcT1Hd+Z0k9lzLikewE4Rztq7tb7mratdLa6W
O+9ZqzZSnCEip5T4sKtnMdesqG7/UKhUpWTtQQ3x56/bjx8n/RBwNStBfFDgsJdcnun0FH/6EyrO
48AoFpqEBgQqgEEOdgFmn6vlJGTDp0GhxxNHFRs8BC851jIYt21i79EkD1fdizigTd6aTK/t71r6
hNK8s4B8Ver8UMQubWLQUOP22NbibBQLoVokk7sUEo0IL2F9I3FYlRqhAGbcWzts7pqtLZeTvXM2
hlRdWopdSo9ikCBEItqdyZXg3O1lWlq1WEcfgSZeg0VS/OP3Y/7EpAs7Pw0qBpaeO1tstHb+HJLY
p8roIwmlNkYjZE4RhxtvUYxCUk4Grl3DKKrGrHuKgwYvsuHBh1Y749O8xtGAcajYD3jiWiBDJG14
YN/ttuC1iNeYdYHTSsYr/6SpcHWRCDayc24Aakbv3PEwYzHaASPtmQF6AAcMcAc2HBCGLe84k9wl
z2kvkfJMZcSjQai/WwWr7HQGcxB6fMzNvJyjnEVcIZO8BTRK30HTiXYlsgH7LL+R9rjFyZPCD/kn
nl882S+XS7A4+BfghwWoK3eiZkQJj/w/CJI4Ym0GqaVHk1waTxoK9hzXHmkhXDYMhceuKr5fG9en
vDOS24OZxwYKhk52aq77lmW4j9F3pcwNY2Z3iRc2VwrwEfo1iKwtC98Jf9xM98JmueOxKjrnGiUZ
Fqh5iPzFJsv4oVJJhSglJiFs3BaQlO0eXOORWpHTKrts2iUX9X8FNlQFcziTKei8bRmK/TepZ582
weMZreTUROvgCCac8bvCvTc4efvN47KWwWUz8LkP30eRD0S3w5PustHEyOi5YrGSjiOC5HCvfL0v
S3OuJtfZAyiNyu+ZXpBOnITF89dx3/tos+dd2ASVh5TvJeE5X81hqL5BR5wqlc6UjWxV5ZhuNviD
IWdBewEEtqJ1GRnYJtGXtTgoBDnsDAvm/w8nnfWPnvbtNMl/+/jX7iE4s2KLXq6yvqYtq7fSOhGF
Vcc+wIuKlOJ9NimD38gBulL1tYBc0bfiBZQVzcAYy6R/EMnZW3pAp5VY5++P81kuPCqtRKDfokCc
Xu8bTG2zCgfaf7wmpSFWzrl3dvs1jKNsEoYElht2SEs//q1zkZRAkcglVbSyyjno0MizvdgTYM5i
+eevM60RC/Ko/7ASx8Bhv74JgtMBnseyxy9bX+MvjmGbEeQIhb1PqmUg5at71K09RX4g3ua5jDQ1
gjUIRmhVYBr0gnxnz8Vkhza9WScce4ZHRMmbG1x9WSGlmqYiyKJxuyIv5mWuVQf6k02TbGSGrRzh
4X8inzI8BmFUVKSg+XjKbRyHwh8IIUqNmj8Jmo9TimOstwdIgSNh3Ht8JgvlStzneSsm3TMr0IlR
zR1UgFX24uy5JTyvXt4t+4PizKoPKmhj70DuanKrDtGm0US1i8GRkniEzXHnwrreSbZYPmCSl/i/
RfQYeRUyj9dMOyFCl6Q34AE+ah9BR7VvETEUToQcZtKmWEPPFuBuO+J9KRAwICtGV2hpEtxCKtLB
TafCnojAwuT3bJCHscdf1PKct2y7/kOmOvNcbjPgnRoQ+ECSfvjnDCH8FKt/hnYN8JG21BiJd36o
42VMOEzbnWDIdlVHB1gWSPn11JInfUHa/Iz2Oj3gO/lP7T4929SsS4kVYY+6Fng68FWW4KrG+r/G
9P48fwa2pxcrsbV2LsTe1rouQKjKVscdM2it3Bb/yLju9Ed2z0GdRkKUcfdmToskgEbwSBbJGuXn
isub1BU5q8x9c2jaA1VTXVN9XXuq/FeprBadoDn+ThW+iH+BzK42JcT7hJTeLbfzZQ+veSMJ+xPh
3zQb1sCjZEQlwRzllfNChlRUXugVUFfAGBfGJ9MK1r2CexfnCKZF0C1DZkIXpCKDrdp/ZF7SeRyz
sGp6kEWEfN9nQDIk49gz4tBznlQ97ZJiA0K+9W/ADkAL4VdQ8iOpZa9DAt2ZzbdnTVG1/0A6YSYJ
nMgh2HLrkOmwOEvfNGi70nwLqR92Gxi+lHfJAVrQalKB/E5WEruOA8MSSAhvMF3MCwTPvi013X3o
ZaI1UAZwvNAELupG0abPM9dbxJ6wdOkeMBWgzEIk5C1EmtsQ82SJ+KQgPQNFgzPNJoGtOHRyZ20M
rUO+WXBd+LAFzuuvB9tggdne0T3hk0inL3ILwXvgm7JZJMM4NFrVnVSMjmSxbZc04zHX86LXW+zB
VyNiRmpbuwSlMtwFqwuS7IRnUHGOIQlP50fXQYqukwZ8+G9RWSjMxJD+FVPOcK4+2JRviQODmCnd
f91Y2dJUMMESb5a8czCWEEyWYEjpnfXUXqoiZ9147iLh0SGHoumqYwGKaIMPhDO8Ieg0eeAHGV7K
kAeER5De3eBowJFmewHTEb5CYioeDvh5jhOpkwEDH9ixQOBlQKR3F+/VL+wjvQ5LA84boY0dGZUF
bMI9vms9XQYRDLHbbhBMzlRN+3/Rc0l2ZwsRQvu3P67ZQMGjB7tFyMmQZBesTAB49s3p19Dg4p69
4axTcTvOkPz2kY+uM+xD+x+Zt8ko8RQqYIaHZ8iHeuAwliPkBgKzayspIGURw6yIhl4yKxJEwwDE
PKCKRW2H0IbusDIQGg3FJEoL29RclnqeVek4/fH9YLWeWloDSq873CrA4RsSNM270YIxkipUKVVv
9UWJNhvC/x9MJ3+Yoaog63VpgWWD4xOtJCUCwyAq83b9Vu43cfYbtK97tl+vc/14iUhjDNHoWRAW
nbeBpiTu2862dHsy+KmVFqraxbiorq3/DyOmqQvw3VAWdXyHTqA0DkGUlJqnkw3utCSEYAxJWUG0
eSkzI863Ejwpbzhzc/w3DiCXUdFDi2MR+l0yiaeg5B0C+cdWHAYtmQxEs1cY+9dY3nx3j4M5OJdL
HwYmQVHdPBWyh5BXD18ZoFuoebDrWqu2kEWiIPG4OhCBGJNMLx1cECY/6s2HXxJvU2OiQ7Mc3qwJ
gNLhnXex7JMOoUVV+KAPihp0MdC5GO3DREk9pQ/dPqppcsN8wWLI0py0+X4Wb9Nu3kF1XEcv/wdp
V34HS/Q+eQWu1IUjtRmmM5yTai2HAvPBa7RaiDwFI29JJ7FCujuqOTpV/zZCp9gRLGzJ2o3jQrg6
ozHZPZ7AFYHhs4IJBz5UTnKv1gbdMY+FzkDS0d+8lmR/ytb4be5i+ctwcKo7oA3iJYnA9i9ev31h
v1wMgkj2wMujVzydo8OEiZUVrYfsaFEacroG8gEGZ7nh0MunD9p1SOAsCK9XhXE6z9Yrq1LVQeZK
PbSQSMSyFRevcuy9gaOMtW+2eMHX/cQ9KM6KixntWv+++YqzCZU36OTkUzHwPGCTcMVdVabcD5O4
6jJmGRHofclY8sF2a9r74Bn7T3irJpOMoHtuUyQvSSgo1AKqf/0TUvWUytsqS9Z/slB+9kJZex9y
nrxNXHBYlo1lKKn8C5S3MfjLbTbp/y4la4+gLbhmC0v6wrQpTzUU0lk0auc1frjA5sU5C1m8e+VC
/5z44cWYz11VDmSdmJKzblV2wYnFaF5/MpVzwxD3OQKBIk6BrkR7E7h3695iTwJv1p6JX15vaUXW
pyVydwqiKY8dMzlJEgghfrupBTKC8/1A/3YXC6XAdGPzC//bWOz/1Jf51g08QQ/5y6QhWzzp6Qcw
uiG8JGwb4MlSvNoo/oD1qLD78kbxMps4KQHBb+PMmMq8tirF02KD13l2C7rLcyYGjMW4b9fKhS8n
nPesWFLjnjNwaSFyqkPBvrEhhlOq3oNRs61bAEYeVbRqetlCR8sX2PY4OpgDutzKbiKVS50jS7rr
ctu9dZmNsRopZITt5GEzrhftn3w5kg3sDBZCegL/ioKxDbFKpf5vFvSE4O6H9E8D3yJwRaGXHFBy
TdhrrG4Gcjc2lnFixND24J2ZpcdtO6V8LnLRfqhAG74u+7z4OV2dUSxDY4CTOhA2OnYdjsR6U7RT
pJuWn0g9uJR57v2YIyVk9VRD7lDa1nq3ZpW4GDBB+1kur7qP0ENhzP+kBTb+Xm2Su/7YQxCXpI1s
RRSt39MAoDHBPkW9khY+q3+zheLqoNYu9zxNjBmo/BiwG/bo6Dk4V4bMN4CkN0TdsghxxIS0IJRP
TdjTz2XdsXliQqffeqzA2YqonwV5ZEwgkibwkLMJYfagBW2scEuCfOQ4ajIhQvYsaI+2e3RO1l5j
83vH5k50D3DQSfG8Eq7D7YaR4yidZAM1ZCE7cJ4DeC3TxuYWw7ixY84iy8KDzLaMnc6PyFSbKSw8
1ot9fgcftIoocZtrLoEyoexfzacy+axwOuGOU4chVFdX1loadCvJwR4irZ0OTZonpQxxGNTERTuu
/X3m5qraotF/h8gniyYNjPHoooQOiNALPW6K2RfWAw7uS3VPV2/m8TSoDehcg7N1eHWZ+bbjfCVz
rtaJNS3ts0Il2/g0wAWEjX5sZFUELbqfCRDyqOAgy5MpPztHTAgfWatSEg4CRib1ALR6Ou7PnW2G
ghciDKjvBMrIJ4Fqc2pHhtOpsa9ViFjEep9/n/li/nLAqFWbafg1yhyjypm96JUN6FePB6MVM9rl
Tm1MNZa/0jE7u67wEwwfO2pGw+bcKGi+JR9ocPyMgNpBSirv5I57IMMQxep8pMygJaQPEHtERSRI
UDp73XQUttJ0dAVUIgcQhoq1CNrTuZPEKh8r1R2caDZgc2vSvaLdeU+Dqd65b5eM95R3xfXMEHms
yJwik+nzuFaGEpxbTFRe5N7hN9rPwMvnYCRSPRlNCOHZRxDPyFCcn+JJNGHi+vmPB0wcWhT3cHnK
Oo8d/CZ+qE8TlAK91WgfLcJ2m63zbX4ENTTZjyqnDyvslgwOtK2bktrKyHw4KgPiunFcjssTLRk1
ubIUrv6Ko4j5jNAJsJqELWfMR71KgDkpoh0qH9yX+yhp70YXkN7ZrtKDyKBD9OVqDWc6Lu275+ti
aHjX0loLtY1WL4pCOc7wmDw7gVIBK+sQmErPiB8xVH5i+QizYiffcRqaAZhl8oVjvMSqr289GTIk
fUIpG51EHBLzksqgOWDPfL1LrQ+S07M8AQA15SeEBzMz5ragkVApZGdtEoXCgmLFugZ65+9jt8tO
7iqC4r3sY13DesHqHafhhhmKdB8cRa5Fmsh/MXE+X/I6tCwKOdrFlD67+y5TqQwU/Bag6XtzVw3/
bMHAcQEIkMor6BYb2S4p3cVGrBsVRUgoLhxj9roJasVeaSR77XQ6o+nOb57rFmFZvP8R369019Cy
iWtUmBkXd0s5Ac1Yu2yzyYmAcrMhpNZgxPR8X3QNGkUv9X9blCq7fb/6O02ySxqh+yu5OwRJQB5e
uFX1qyj01zsG6zZuECfFSXfMK6v/0c8gnqWtOIDTvS83LMo+yZjP+4M74gZ2OHI9pNgPFZvAI+wk
o6PfT4QpF+R/TLVlbphdizipNW41wp5bxo1clYWmigdt6vSeWBIhN1rOqp2ajrZ0GOQvq8WX5v8W
Zz4Dv6BniUUi5JJiv84//Xof1zhbtZy0+jLhnb88Q7QcbhCfsEf8Y5ufZO4WFj2DFxS8o2L3ACKt
KGPezHS9eTgnHDcO+07AqU0MrUdeD1eSt26FW+jV3ilCqE5cWnh1/4ig+OFImuRl1bekOLPItNPW
FD0GO6JfWG5JoXOFMZbj99okEtf5cvoU+E+QGTDqKGpqtKnosJ+Kk13iB3vbENOIpndJ6FpZnC6R
Zf9EAXY4dnoQH91IBeJexUQwq/t91aM3SI9ImrtRdWC+zwa5zhxTsZMDDnlSixtH2Mqa6QaTl9wJ
jo2jC83td2XyopWhr4/h370l1uRJYdphYkBnb7KJP8NY8dPJIr/lZy63K3Xoq9V3Cj3z40DSxNbc
AbO8fvFLb+xfr89PztN3kvEmDdQFisJ5ZDsUhdXAagYveae+ko7wEbyZXl2XU4bAKSKptIlPQhLp
V6SlUYLIO8On1gPcaneQCF3wW9gUqIPGeDAX4raGlrPXZfoIbEZQFv2ap90n0N8qWkR7WPMcxKau
awILKlsaWaj+icMKINmooa6EE30GNgaiLtwuZnSj/Ar1cLo2JtKA4LWAWaI0wIz3DIJ/m9I4HqpJ
hK4gQuRqZIOMhaH76mV8yus+pT/XyCoVktqRvtj/rEv4kdupoAOa7/0gszhxyPhryu9iubwyVf5d
hWgn0KWf6EEyc5obglDvutWHHOxKYczxU/94pEfs/r/fl/nV0xCoE2YNaWLOIO5TWXMeJmBUBDKV
7mCjmoYO/yZoecv5WcS4KEPUtMX4/IeHJ1XkDOEJG6DESfqbJoDx+E7QTthdUH22Na/Zsj5eUIQ2
kFGoG47yyqAmaHD8evIUOmw+y5IybChl6I9tfDAX4fre4pFm5n1F9VsDEGNXSjvCCPCzrwYGXcBb
ru+NwRue1Al/uISJedFTR9dcnRelfIrOk43muWnJCG6bEfWoBFh1Gc6U27BsKI5WkdWNS2ZD7nZG
XYUdUYd/7qJU6PqeOC9k/nkm/JxFMOSCzWEFGnDqcwRDuWEhd1yeXSVtEVnbqKMpTtmWp+6jDSVe
kTgue0l+z0ItZAkRjRFvqLLWXmBvcl36VroiIjdvDdl2PPSuXMjPLmxvQ6aZ90z8XGa+iGROQSkk
EK6oczOrkpp6r/ppoUNtNHqyaQlWdL/XtHeRXOTi1tqCOrXoBI1KorU+InP74/w9r77nSTT4JXcD
pmPjJBc4YhQK0msjJxgBP7ObdzoBMkoVd8YpO4cIHE4O3pBt3NY0m76kuycqMYOnXKjwbJZ2yU4O
V0jthBPO93WiugDL5RQkX5a23saXRvz+UJdjLb+2vlSLsp0bcvxGuueuzZptr8neRdz6jUS2fMUL
iKkJefbNW7y4k/3eCtsngxGDI2k46RARN70qdLcXVV7cdATRs94pw1IzW2xNhxIaN3gh5NWD4a4O
ubORWZeZrffL8VF4BNRCvCr0o9+2U3NnKktAaXGRp8523ppAnKQhEeB4E+5JZleOgSR8phjZRRnT
DvcHtPg+YMBEFphz1SW817IA3k9K9+YZgdp82m4rtG7HarfLyfxrmkBt5cu//VQi3JJax1klRAFt
8b3RoUr7XvU3XGxhdz17Dp394i8UwQ8poMjg4tW7f9WzKPEGz61//PsXabF4mGOMwoHo9b0O2Z/C
B1nApNdNF/Go5zwnZ6GzK38ywE4okYwEg6E+ZemOBVBRhQChWnlHg8i5bZHTFBE+GCF6cW42fvbr
6wspLrQI5n09UI9mVreGsXo7iZU/yVW3gkiMm+OzaU6VI8pfoxB2BmU3LNLD0aypR7woApWW2SAl
gbRRA9UTH51aHfcLfWMGprUf+miGfctZD9ShxH/gPZ1uOJc42VvdvOvFRC9mod9SA0IMImivPzP7
BdsTy5Elxi958WjH+WcggHyTu2DhwjVtCrhqW9FgNL045vQWQeqM54kjgVSGe9PdMEAnVJW98PUo
UwA3phF+vbGyqF7itSh5YeOcuX07kgzSugsMmKJl8O0EQeg84ql5rjgGkQLiU7GzHJt0R0+HqD2d
XT5vaePPlce0ZQjSwt09ItLVsDr/lT3YrHBcurTnoeMWjlt8SKp5SgvvJShIUg3p2KlRhfqCGuBc
c14Y+2Wjsr0dmTG5h6Bd+dsI9pIT8AkZ8cpaOC1gq8b8xutWOyQvULJExi6LLpItpELOzvlTmm3c
aO93VWDbl0IYNRANkPQWLM4A5OPCmYrZw6uo3TaviyZR0ELH67zSrpXr/sstH6q8K4z7qZHRDYU5
mWz5ea6LdYxUmYcBMKBDtxJCQeE8aXXJNLECPrWeBr8qHDpDEQ6zx4shH1i9vD5Inswe+5RHrSXX
luREy57spsTBcS7sWqaK06fysa2YXBKs3lasqeJbS1rCKUbeHKAujLNB3bS8El8gDX8fUEy+o3j1
Th9Jy3XiO5DlexzGICBKytso4Jf9C+w7N7OSC+BdxAgFfGl/Gy8kSaiAqDdX+n2FVFYy4RUO2vBJ
YubfdJC02LOfG/ldsWxghblQ0k8yt5ADNzruddH9Mt0aw5W3qG7WeoZ783kOIoJdLkOQKez1OxTX
uGlY1zaIcdv2xdFEgMTtYnSEKZ482iPaOcmBizE22CYFAT8PNBz29jAvxz73Cab1AFl9aMdLUxnh
LS59qvPnMhwW9rW67CTONVfm/qgPjHbqqDGdi9UfUeUWTxL5VxNZp9phsBY9ay/dEKCqC/OzKrlL
wA6oAImwI4cwhLb+XSJx682RaTT3PNTp3t8Me7Eh+weaLuDlopkAbMXj2RaRfy14GJWhC0vsi29M
1gA06/0bD72kEA3h8pSiZUxJeGaMHZeOWswcIQMkmD4ZjDxLj2bFtH+rcfUSgZ580CFPOdr6ZFmJ
Ns/TpjPHzzkwTQ3T0Hhce3CDxEhrRhRz7C/WzA1qknWPGSPIz31pB/me8ZQTBfmkZ58zsTy7Nf/c
/Iq5P6HdrfxEdJojmp9cHTPkKM5macR73dJhB8EuFNaBd0LhQ25wQUKM7sH+rZne17baptAWM/og
+0i3GmH+WrUoQxuz9IN32+izSewXYU0lvGWqo1oOZYzf7xZnjgWg03i/mDuMMlsRayI8QDPUKqLn
0pPcjZ8GGMMVLONaH9aC1WpwVqgnT82kT7As0rZIN5FJWayN/KU79h0susNBQZH5sk2YFvqYZ3qx
jZmfvcnliPISfSAcfjAva1VUXX5bpqwOcr2E08OdkQD27+OdTkY6wAHVp85mQiyPSFxPVYPI/c68
JB1P2hE4FQ0+rGZGC/AIoJei0YzS+EcBNngxyqqQFKzFdyMVC+vj/eOmWVKAsFKspPGN2ikhX92A
miUHeYFmYT79zs1UrpKPzMnjQmprxJs99S3UAaR7AA5XCa7wWe8rMD7NVUXmch6Eea9YtcrtShwU
sC89A9c/IybIc9EVeSIj7HmYjzOeHVSHiAYiTBAnF8i6ssK75LS9+nIxIp1IjU4vBOTsLcMhyCoJ
palM1KzRkdxFB8DAVQlqsVogq6B60rb8OFaKAf1oJMa5oo6kM8p+raTyoFxfV1RQWKOhmAnMdGxT
vrunNf2og6+kQY1ibebt5JmWx1Dl0jp/rS4wqUGC0hVIJNVzr+ZN6x/HVfEgZkBuPwvKUNYp4Xb6
FpzGHKKBfxS1EmdqAK6CaMArz9vEQSlHOZrLIx+JrCBxyjxQkRVaDg4q06HkYMjM6E/i7pMUCe5c
I1kNWJob9xUOfS2KC15zXhR3fCxKmp31kxFsYuUTh0KkCqfx1nfPxSelYk34znAICuOfFsTtk+5Z
4H50hqsu535a4F4Fv7GWmhTX6ZnTSKzAPGyK5nMhETvuWs6PUrC0HofgQeg7ykcxkKQk3Wc06icu
xP1ftn2hb26fENI4TUE51oT38bn24t/BD6Ypum9ppFmN77Wtd2UIT0o79mMFkbOuJcOH7iTV0Vfj
rBSxsZqBpoP2r7w2tgoiAxJOoxeTp/UQcDrV112Pobz6WMkU1VQGyGh9uQpFZTlSQH5t1VwpWPQ2
FCTcVvoh3B3CDsdkn++S5LZFgVnK4CA598XSL+oSIRHPJZOS/2/6jIJnLqHDtxpfEWS1AsNTdCyO
V8iRAuTXLp5U6vFOF8Zn/xCHYCVp8olJlKQBXLoyhfB70RjVHq7yg0x4NLG7G+evT5rwABw5PfwH
OX25oulqQs481V6jEacSmOibosDIax1SusnG0Yb3KUvcXLEZ0XYERELCMmAAEsWdd38iAEvIzzrZ
JTNfSTMGNdWZGdH3L3SBLasiXL+qPCCNP5xnze7phD+eJGiI84LQaWtokRJ/lMf2TjtLkku7kMDZ
ZRigwPrFqcPCBCPu/khga+oVOMJupYPnG6qoKOXAvOHTuYVYs364HQajx1gsguLxVt1C5WRoAC9E
o+QeVbzTlwwsYY+dqCX/bmyAc5M1b841AUHvYRMM8wLYLuaGp1v+TXJHkuxfwmbUW2gF4S/FU9CK
0JiP7bEoYebueY9sZlZoQlKCphqglo0+/O4zZlW+d/WPAdTI0FkdFFfSBEun/oujCAArX/CIj82v
A9BLZs6PKI/R+acSDMCdjfCLoTAZv7YpOE31xUwt1A6DnYpIYdl+t1nIW12IgqmsVXz0+wuXQruR
SKok3vtFBLpMAWZnFUWwNKjPMFD8D60RQP+mZWQP1bOFAU3ftxJ3tiQdkWQ0maR/a5B2JRfph8t/
gfIZoOBsBIMoe/h8yVCZpXFmCQDMExIELJi2Dru/pbMGg5mI2PVxNAkeKBbwLO3j0yibvHvzgKsz
rtVRo5ZJrmVlgfkMaNPC1DYg9IjIlhn9BE1AlmQNLsNQGhg9nU7ScrTnYaSIm/Cc59hFqB+oj+bI
dfLm6oNeuwFw4jw3MbB9cCFgi1wzpJXMnIP0yYsa+rnJYzvbD5PUsxQrOG1dAbrZ2TJABdXpuyao
ufzKKjyxbte6FyQgfWqJBNj1oF04loSABaVU0NJ9usKaixfwsPeCtLBWbzUTVYQDD5mjfsrT/fd7
0ZRiE8edw1Da6og5O5grdkt7+fFzMFpmcJnSPWrcM3J4T/KY5oslgIC2t5PWcE3C+qbEFxDivBQq
+tQGJfX+64PpEjrOuMku8eNo5so/IqL1LWMTt5l3XpfizFheOXYnJeSO1GXBMAIWtFBY0jhxnGOx
khlK00WB3bZlOH4DXdPR/7wKBcX9U7mNknpu8AEDiIKrVv3eht7jV1+zaWdlqvUZbhOWzZ0jksUZ
5K+zVLV7pHfj9+DKySIReWWM9L5smJ/KNogZJaOB45yIkPmykeaELCgLXc+qkm3Lj2kww3Rut7Iv
q+vdQnoeboKFbUnp3IbQodhgEWq0s4PO3D8GIDqcuVbDfomjbCYIF+MAApaqYipbXlvyNo0eROwy
TtISXPm+GjS+Bwhmxqw31tjdPivkx4Sjd1YhYIptCKLCBdPAIBHmC/oBwA+mv/r0NicPEJ8o8oBO
emDIWgmO5B4s1DZzUF9FJP9Z/8Dpf4B1LK0zSwY4c0/BfQc1Yvth1zM2//ABFwCX2yhz9naV2+SU
WnfMZjjERORgdNexpsT0el56Eeuc3oaW8FO1tVoNMtWGSl7aL0n3PnIj6RZ6cmdqaw3+0+VnT99D
VXFSjsPA2ELwVbYDL9oMTs/FmUC3h+LMhps172J0/5rB1Qcy7zBEenvxkU70h3J9YLf6VABI8yqD
cCwwIYvVtss+f1B5SA4/aW4SEfd+lOVWW+y9hq3eLQeYhW7nFGZLhyktWfY5W0l5epOI9n94xa7w
Vg3EASRl6g6Fw1GGQgRO8Bwn7ywyQAjK+p0c+Q11SNMd0CE/7JePorlcwZjTgUZPTFrIUzzulGUm
KuTAONCzRxYpCYybwH9cmXWTKwUZr5e9If3Rf+R8YV009f5v2fsm59cZLLWKq+M64otQp5P1mdam
EFs4GR43u6zIn1gDikGMmwiJKB7MaL5Ns12EK5pkCAkNyii2p7O0dEETYb3rH2S+7X+yvD8eOti+
mFaC+vCz2r8xPyzj8Mkx3cfnppgqqwfRM+G3bh54HztnJCewzmDaMffYMiUKyCxsjDunxvh/mUai
odbw/nTMEbVXWJW2VNekSo74sdZUumLx34SP+YiUvqs3UC9Tihgu9qKXNlFb+OuMhPmTwDyLYLza
AGxjCyqlrpeuf0taZQirDzXIRorGcm7gArZq+fr75Hpu6Vl6AfqQL+NCrDMuZn3hiMgP7Db8TqSK
DJ3Gzz6RyBLt1hZBHsW+1Co4PJnK5PscJlcydYMxgAd2l80/J+7Y2Le1mVaG6PsMja9Uf6EZlQiP
FSz5gJxmL8GUIJsRboU608z/TIEgPEvi+eaujaVIDdIPsyqkRvB1WNxPEIUV+hJj/trViW0wYVRc
Ce71okrPtKax2wnII1Gvz+HLVzieCYwKErIVDWVKrst/8LwWHL0Z1zmtS1OZPhaboW/KReuQFZnc
LvRJIdMiRZ4urUEXx+qNnI4TRbu/DJ1nv7ZEtjn50cF6mtZ1VpbjbKhftLVFLDfLWW0abRBtCyFZ
Fr6wPo20XerClOYnTy2xnY4clserMnEBMtrX/tb5ETZi+tk4s/cA0qwS73BmToHnzyRxN0sfsZlA
140zpvkwncUecA5ge8O/TEsLsZ9R3L5qYvKiMXnZ7KxKUzjDDwjFhzvlucmwkztPzjlAhHXYFQVM
fDPG4nMZn9xC51I5Uj+Inb05wg/brwq3fQiDP8OowqJxH0CnnI9qVaUvFo+vP78s/dr3iG/A7id8
+B3q4PMFsjo5jt13loNq3mIVBIsVH7lGLXW5lQdDifQAWRqGdlQA6ph7vcOgJ+Re5yFLaR4UW02U
IdQmMdazdaKFttNPLzmTnfIpzOnYedMJIkbbdk3D0Bh+umEmKflPl3AWzEjxDV4cezGmNIF3949/
W22k9NCewWtIFu4o+e9H5MTfBthaKxShDq1I5z4bcSWwGU4qg+1jSc4xZq/YuS4B48Hq4Hso1ynp
ZLfaM3XyT6DpDlSH54VOHAs7a25bSbKhMCYja/SzF0HbmWe+TwKjIu0L/amQOzmg+ti43ns45q4P
JiG0wIePFL9mSYimwNegiT2o4xNtZw4Nre8NJwrqgAbH3d2a8BpN+1NGMq7orI4sCiqpDBrTV1AZ
RGRqaqGZnOWK/5JopmV6vLRKGcfKGVYj1EF65XdltYBOwiWfTpohE5NlWZo83v5rtAj/FPLtisY0
brN1cpePJk7QaScThiZ4NHLh9Yt3XFLtPQw5omCdyI5wmjkRpHEqhCqC7p0aqZxRxRjwUWQrZDFE
w5RhgcoFd4zyar/JVPb8wu7dJXGgzuqY+A3JnV/bjpoMu7B5OqOuUqWH0WmVz3L3xQwRej2KN91m
s5hnePGXFJKPSyahPTVX7OBtjC6cbjb4JZrisbxELRN/E++g5kmnAXFEnFLe3TGg5FFU2PULozH6
6kTY6MB76MekUhtkszmGIQJ6a3MqaFAvl534NGiMeKTbL7qByweUb7fp+R7BsTTyCRqJsM7rJA+t
IG0AqaRavxB/AKST2RUi/YEtL81mkrUaeJ0+ChjYAjloeNM17HvbMf8iqsATQrj6r1CRu16+We4Z
+WE0DYabC0qk5t7L5e8tJn5jkmLaGG6wMCZI7ETYcbLpUkYCZXGoi2+3wewvMlbMTRFjZmR8z9tw
EezfOXm1qtcDu6q4Ina5pvjMU6NcywfzwRFYj1PvBAp/Qar3Db3SzXcQjR8JhvD2IIPkPMHc68U6
JYTk7qXMN1Df9+zUfVTZv7vVvhuXtyeGzkG1moJmp8wihGJLLrk2WgNqCekNsmcBJq/92tVcyba1
cm2H+o/aHPOghCiD6S8DNf2jRKFyDghRb99y1+eNkHcrSvLy4VM4C6Q8s5ayxPW9y9ZvvKbhDsDv
sTdaAiTiZRheQQyGW7y9INGGVSXWxEwEEXxtQRI7WBrmDhZA1NesRwA5iIY0EXiRmHMqwWt8sLaS
7GA6I6SO64COlpGeeV+BeAe4NYTlaFB/b53s3+HQKEXU9hZrKiHpsW15dfWD2Qbs3t9mww32/uKV
Ga1Rl+2tDlfH5h2AFu5rH16OVmkaShbEoyws6Ek2ZbcR6Jo3dWq8zTpuk+7FtLsD5LVmB0rJA7e2
KLxXT7pjFN0pOztDncRhfenCSPZfr0XQVyjxecjogr+n0FonDgyVilaivCtyI5PTahzC48hKeum3
FvbMYUEbUXqoC83Fqr9n+5s7UcmAyzpZhpSQQM8lRWEq/NhdhMISY6/sKF0IIvzn0jJUB5/fqX07
rk6O87RMoKjDYY3W3YubEPCa/KbF++3q3vavPCoCD9IOgntVwrJKwbqNThh4rXlJ/8NJTNw4LFOh
sk3LHMNuZOOKSyx+dlNU1NeE7oyGaVwIvUYspzPz/WoQqDk8i6YRwwtHbqLvfVxvNVnZFJRK0VuP
s2TkNT9ZYI5D8z8wRXZ69YPGSfz5B/Esd+HKQTYlgflCphu2elLqDSJVSk4PAnKJCbDBzcltr23q
QODtQ04cSvsU7VvpjTfTjaxuDxArS088Be7Kk6jdIlf3mQtpEeG/gm1MS/JIef7Ya0mywixePv09
1NR2N6LQabrMZSJ9+AmfeZQkw/tOSqbBPo03nPf0kdSA2BFhXIRzBek8ht0VHyRi0JrIPlr+ibQA
kPeIzl68JdaGfONwwhPuoeaXcEsgS1B93TzMJFiFIUEMcpCK01i5uETheEvQjDUWDQ1E8lXNSH6N
HwTRm3X9w9u6uEI0eSP1FNTRtrwBiCO8B3TjZxCMDZSsTB5lFlHgdpLf0U975Qcvll6vExcWQ9Tz
26Mb8zHoYL/TYB9foDH12NjmNyRgtCoXv79wORBGhlU5mjY619H2AE/zp1KrCQcogz63dRI9NCfu
8a5rJJ/pU/m5x7UkL5Nof3toqMElC8tcwkT2R1DiOSAlREVVhm8oCqpveY6mUGeZtjtV+yCQNW/e
ukEyMLspPG/sud273fZ8KqK/qiiufaIhRhGNwQuRdF81P7YEI5and9KWR8C7EGdWSJ8X1/ye+cUI
xFNW9FDTjyDTXXjfD8+TiSUcQbP4eD5fZ18Y2ukHK3VbKx0AYEmZAPysZ27jYtPKj7PbQwc4p+gn
khLX2bcww7zAug7TXmsvd8yAgbm2idYsLRGwexrp7QlQwcMLiHuEpVADowFVo25RiT+1m0MmDbzu
dUy7QajHzZQD1S37+YwRwMeO/9hEVq62vXG6wdjHXLcrsONlSaoQnDFxnIEBoWbYaQR8BsVw1ajm
8pSEXOHgaR53L1vn9hgucJlpHPYDvCMqmSe4Zn4eRMoUcfwfvEWzibUCyp7uP8kCh9XFgu5NJ434
PntvThk6UuQDutHMDY7knlqt5HDxXIrAhmTVIJ//u7q7xr8m/itG6NO3UAh0D9gZELTdIg4Vu1fd
fuSY1j5hG4naHICTLvEMadicQa2JLtr1OdF/z3ZNeCAwECEgNkU71ryeGYCuDRlWutwgDOEgCYA1
b1aBjl3+7l/jKBuNkTJJFIvjAtP1tgl/sZWGv92qWF5Pl6C3gbD9r2qFmHLrdwtIpagP4R7piwLW
1plooYgQF/Bfoddcy4KDuBzfFDC/QaoA7xIOSQGA311mV+Hq7JLF9bq4FcHQ4VIxCeFmxyLZoD0k
DGUWViFCHM/egB3eYUFFybE8YJUke2HhzonTEjHEJxcQnRokShbUMLlO3S2kjtZZotJsxrpPOgVp
0Uvsphbk2t//NeAw5rToqRCaRetbGI92DWkJALj8Cgjfkf5hNJEd82IsroPViKXTQdJqqUUppGTq
UvA1Ow/DnvV/wStYnf7yVVEcBPMc7VNL4N+7IvZPjtq/D+q5VmpiQHA4XtLKyo8VBiRc1YQATDg6
rOX1CF+QjohXNRza23g5Q5B/TqYilXdeO4NClNduPsyxKgd4KR3puu4Vfod/kobACA6U7kklBTkd
JyBb+2/yJY6WaIJZhFvdIC2qYEG70aW4p8Jxh1yEHp66yzYZpSp8e6oE6zbH9h3HbIpedB3IZwhO
iYa6GhiJ/KPDU1kRqQeDTWf6/JIJHlmJesq2r6fAlenPTUKhXvrR0y7X2Qwl/aoLYqsEh7s/FeOX
9K8Uh0dsdkNnBzsP1bu54kUgxxarO6CBo+17mzacCX8gASGthdPu1NgYq9gYOJpSR40PJyThmR5w
jb9M37xX+vwCnHA4ZfJFCAQ2eK1ZsjZUIaOhPaHkTLZAnTW/O93waowBLQgVxtQ5nyr6JDMWbSNo
58YgeD4rdot7QjVGMJ50TWxhNCl5XOM8v3PFasDBozO/QbSFgzn3xL2MWtZUBj2JehFsykQu8Cx9
mQvxiLSDrN9bw/y7ciO1G/pHeeJ7ps7eadTV5WhlxyUem0HirR6n0abmSSjGcGAmtRqxkJSmhZK2
Gq6XJFnJDedt2Jm24lh9hKwPW1IgZd9EbOot9WMenJFp0eduAfEs8YGS0r0tQ7CYfqnLWKb4AZ1o
BCvRpisusA6TkCzq6sXu3j/GtzQNQ1PYaf9LcHvTbHiOuOAYQcXjzTFoQ7rN2obxRI0fNx9JMhXg
w9tOt5PIFjm3qrXsWk1gUhm0ls8rjnbDSNKdxXbBkwE8xX16T2oMpzIfa9+9l7vGm8I626RhkNdr
gQLO1l/2C2ulFa6VotFexzYY/LdSGi50N0jYZf+S03ERIV7cldoZEFL28e4G2XEI7/FRMEKRdYkW
SLDcJZH9B0OR9y8PUDiCCdA4RQSEOOjmaQ1zAIUDoiw30pDRVHCtCpJ1yWeNkhSiTESR/EDJQ5IN
cuUUSOvehaTsNxWFQfWUgiN9OWB7KGtx5nvW0s6/DERpK8r3RYVOnqCnwtKgNzv9NZDzZ6CyktC/
NzLDBeIfiU5BHOvZ69uO/1xU5/kE7DGEp5gnrVB11DgiJdisKp+lMtcZo9GSXPKO/TLki9huk52Q
p2xua9DHfgOLHrX4CIJeQnStyUT16jcJJCw6FdjX95FSiZuQjkvOldbRJ+9JYLXcQnpA61IxflG/
yWY+7XAW1l0AEcRVCK3TU/H8+33Wx7C/2E8mtfKSpna7GB5KzmWUmC1z3fqU4rv27srxJp1p5A5F
exRX6LbAU0DqVXztrCQvNys/z0KKi0i56bVxzBVDvwfqRXtd/ct1xwShA7LAR53T71+Tl4vPFDvS
nTXY1yUaxgRaNHGXBAd1DNmMHRN1RGPlBVNKhBCZNvO5u8ApROcWaWlsSwMgXGthB/YCdCVdEPvN
EmLnUuig27ChNLsTfU6rrZdwqgrxJit4rRGPMc78jB+llb+5+/4XjWT0x6krukED4vRJt52+/bgy
i9gqfTOxQnChkNdCAhVNjrI4y5naGUwezm5ztD3XU9C4JUDOk7d88+OQwrQFenT8OpGa+BeiJLmn
KKaSXl8Bt6vMGxs7GF26oNQTlUx64YbJJqfm5qyfH9zZ+nbXJK0RVVFCzSWH1zcXqJzBzn1LhlC2
NRQg3vTIYcueU7W4uPFc8kAgmu88S9P2zlzRADSm/Q/nJQNN8v/9ZIlMK9LzWzPfJuKVwHvzjlsK
I4Qyq4onTXpXtmmPsvpWxZTpGgoFBz+FK6WVqBl5RIUOKgRQgZUrcN2Rl3m1UgztBjgasPgvUiIg
YbZVu0lSZZ7JG7HOqucoa8+6J6I20nHCG5MK3mWrO2J9iSamBuzmM+i4EKL6hh/mpV7DajlgFUCO
gZ3BK8U8rhq/fN7yXDzVMHjBNn0RUegJXPKqHB1nwehfX3uxIl2O+Gr5GC32cpbVerXGcXCwIZXO
dsNma69udL7rTQg3zLNJZLS6yAoL+7hy4/Wcxn56gj/UthiXbfNCX6eAhzVR3P4fjHFfX5CC6qnO
IU7sMRQPp+h7GbTanrI5ne8iSKqRUacuLcpuyHj9abMG/c8qSj/7bUV0lOoA8VyOUXbXIWxwvIXy
kxn427T3QM/TLM4FQUQXoji8crapD1WLpoRBPE+xriZQjYnv3UgCfFzI1hDDLPa5CE24CNGKGaMm
wqZy/w90GeJxsEwaUA9AYZ9lajFncgNxyQwajxRTGHPdGeWioUPbyOMnZUal+PS7Rl4HLzPQMcIE
+yK8820dJZ9vw8T38fu1VgbU+6a6uzO6WBtJxcMFqsCvB8wI9BmHNp6bYQHysqjm7rESYj2nSTeM
d0kkq1OMP3H5SuP9tYoD3GFw/xLGpM2wbVhdKE2YgBDwp+ii4xqEstkdXgvD7l44IT7T+1JqQX8Q
0lzoZxhm0z9Lyn+9ggJZTXVNkflNL233bFdttAgduDNcp5bvXL0icnd1ICInuSxIv6ANEODoXdU3
7YSUwfwy9RQZK8I6Q0HV97io6FpRlTcQxCXmb3QaIMJGX92UBLusG2TPwQ7q1SdEVylLcCCS3K+p
wvqySgdOaJjPzTVybSAzMKNXJ4xJ1E+g/2uzH/KzJCWuZtEn6qF10bgC5yQnlP5uCgfcD5gXoYLv
qsQ7PqMxvo1wYch7QWMbbVZxplcfN3q4kvP/n4RdG5WLHhziiGWJpRmiDj+k6WQIKJivnZ9/Ps+u
QcMt7+KqmXlVL2vwkhnJlJhq9Qp2lceEkbEhboxoRRU41e4/tlPHRELfr0VCkiXhVkltKb4Wl4Zz
rH5hNYNGS+UXXo3bkPgcr4ljKOJstEEOwDoupMJIYZshEPDWR2fX2Tho3T41BeYL8cSpbS563IN6
ofNMWjK/hWRwaJ3olklKHDAsqhZTM/Q0+PPcU4uO+lwdjjN/Nx4CZ+JSC5y76GXdol5L4Eul3ET0
v5p09muAzhQC3bk5S6MCDUWEatYm2RyKWWoBf8APKiJL8vJP9aOOSGFywMagsn8oRO6S4SXXKw6S
nQjhqcNO3pQ9j1FXPS3GwbaH+tqHfxJpgLu0DCCfeeddyh8C6mrFBvJ3sqfS8HtEusaWrcGQ5D8S
X/21kRQeuDMbdfSsasAr4GkhVPCiXn9nIrylZYOBLze1kG1oLxWRTSDlCsZoxW7WJFHEuabsVdpy
m4vL/RDTgUJsOrTv8k1gneYUTT3+f9lGiD5I0Mn7IIPRg2jlg6lXVU2HbrX3B5AAMEvSQxM6qBwR
id6M36nVe8RRRUs0LxlZv4r1S2BvDMQe9JQ4Z3GcqhWWrgX9cZPSxUoLZyHAN7EpZPJoM2IQ2d4/
oRFLWm/r46261yJudRTUWKM45WCSzqfVZudCpeI/qSK5b7oWfuuNKENWYnxYWP/bOytVrKvNI968
vvteDwXOXC1NUL7DPCGXzNUblJnG8PvpIxngVsQS5ZlibXjh8LwlIvXO5uV34hileZVQI3qJkJWu
VItKRfEwM62edEfkz2dh5d3euDSMJWNV+otofzBwNwatP1Fe6PgOxgmlyHu4nkLz/hz/VuMCHZKe
d1MoxIXgWJSLzTWcKZuXisuMEyFIQXSQbZQgRhGuxNaNi2qrISqwfklylAr0aMYzznGQovXNQWd9
Wy67jv8uCpRtVgGrSeQQ2ojsCtPepcus3/hieA7b8SiwxbXBk/j+1I5j/iw2aHgGZq5kArorOxNq
Pi7d8ZV87krs6UozFUHqF0n3wZfbbPTdfIUMTIgQd2No/m40NNCF3tTl2X6bUDkd00ie8FybjVMO
4HtkQj3RS4kw9OlPceOf6n70J4K5scrP19uo0MqWl5XM+YoZ8rOPO5gnvtr29ux10mB078YXbGmr
3daSb0DsjxaNwVQ+UA7PddHJ/IkDqT5OhIVUO51pk6HvBigE8KAXScCCMaRoS6yjDPym/drEatIw
bTtKid0wwhSMYOxRlyDrxjBzfX48OPZ2SrsvGtYrDlfdBhOIHp/tP5RT+O4cTSyZCKGHGV+ALw3A
bCuECZhqGn8TXvBDGdE8N8y2p1D+ZbLv0c2z9TgYQXTPStt2KJkanedhbWeIPgbEHUDW8LmYw7nh
EO6f7vfjb1RGtJ1jw2BS49jrmEqT3XOntJvmWZ6by9Tqj6eaPv74rbutJEt42nRrKGb7zUpuu02d
+pvsZ4YB0wKTQhQPwbcGoqEDUwMkPd3t6ziUTU+1POUTEaQKD6wkBmYKEky8CeIaosrS07X1keyX
Rlk2K07FZqzWwI9+1ffY/Zrlrv2l+6KU8q9YxmrRlRwm8aXvUnomLtPsiB1RNzf87eQ+7FwFVyPu
XlQtmE8jGUISfVA9cu2ZbqzgDfN/H7BFaNrwQYxAtif7WKMGOpBsQGo6k7mGgmCcelxvvNGKVn3w
18FMsVxac+7hrVGj0wcgcWr5hwiknK2RSCbEA+zHJQ0r3MefASyZH6db8qDehGhxvMHRrvw1E7Y1
TSA0pm2zegQCArMUGIUBRIKE/vkm10bEFTquzxm2R1vC97gALRB7YygGr7vU8QZT92QsgudzHfK+
aJuhKHBYYKf/BeJmJ+TrxpWlAMX5w02xWehi5A4Mng5A1er6+fXeQuRoa4kFn0Ybg7swrQxkvgSP
DshKYor66Ki024Kf5zbBIF4vgAvpJ1dhFhXxpR0Yaz9moyZPrF+KDWthJurN4I/UxLa7/FVze+17
+MQm+3wCPy7cqDGsmyoSD+fw+HhR/aaP0NjDj75hMZXqqjvAOSkFOGUbZhRRuRPGqlYZ+ZTsxQMh
N7vlzv1wPibVnAagSerfLau0ox6WO2hI6nJg8CbbDpIXPjs/t8w3kBT5cnIaMFdCDt0T52ooYLq5
DSP6aoEtVJFPVnvwAyryf6lx9y1e3LQTbo9SLV0tclQC5e05/VeOOqgjQxE3ru1+2wn8LgpgyddB
OXjEjx3/tv8Nqs41otSh1shu7Q4omkyNJPjsVcB4yl4fjbVizDJ8tkG5/hQmWBAV9aesMkm4zaGt
BotlYu9tFTnjg2T36eAM7ILHz+38lSv6SEiV2Q3yqXxC6ikdLAthbRxRc73H/DcSVLMfaZOikuss
BzLgk95Z60zY+gV2XowpOewtqNiRxbviC4AJMLFaVz0tOLZvM6P+2RDuF7h8U9Nqv2TnTexmWenM
Sj3wwzCxCT/wA6rLg0lu5vDZSI+vt9quVzRpTuQj/Z5jXu+xJkw9BqOOkTtdunkdm2/YjpCteC6R
UE+LKY4WqnlCAviARhQXuhwBdMEA5wumYCq+YWIOVvNQ0nsOqCzfDHgZsGalkXsltI0k/L15QT1i
8k7SV7rIrRGG0t7NUAzTft08HipvTPtQoI0Q4GRCzkEO/VNfIZjLTjuVCIPlq4b3Pxr5It5iDBKr
S4OP6OeSIEN1GSt0hTwJZ09d2cW7h6o2ENPJZbq2LGHUX2mnNcMA0oNqB2vshECJbFavG4Cy4dZq
K9Tyxfs5DTWX9jAZ0YRPlSCzJDFN5vzoOPZVdqwuojCdsjANPQ2mQtx1E4V2a5DD7nGyDItULNQb
ldT52Me6MLS+fR0qqYmIBI4gkDpMQRJog7tBylQTyO4/GuzGtOoS4ZcIOCEV8pR+rfLq+NDth0JZ
Ns0j914xXIo3ALe/7T9GobhLYMNRcm89L+ttaIRuDFXJRGq/LYTXvzlMdFJ+qJ18SYNTLVY07UJc
RqsbjJIy4ulUZPwZHzBacidNCtHJl7zpzZIYvmFVz8hHhEC5KUSYni81jErK4Ex7kNEdA3F4HIum
SqUxb4tRJfCvJXMb9fli0VGc8DfSsjlulUU0/jiwAW0mj1d8JzE93iYbWem08lhIvK7zufclb+Mn
EwwiUoX+I+dtroUTKgCvi/+/iqhnDlYT/AIexBCJohOal3WluygMJKtX+KjU8isX096xTOfGfp3d
TTHoerq+wIe5mdzrhj6ZafKqqGLVJmEgChCcv8TEYmguA89wX19oxRmGhUUWDFY3AQcNzDIrwN0s
lSQzIzHi17mZ4MCvD4Uu79PSSbKTl+8zp5LtpdYqw2Ym2jYBJvYgTFA3M3nY1UhRwy5uw2GQHwCH
hxhwD4zpmrmgZPSR7TFJigg3y6ypzCaFoyY/0JQVzenkcdP1c25zXdtEBDvJ2GAnVmWq3gPP9ULd
sjan2eU07Ssf8CcU5f20Lw2wVIr39Hvo5fJ2gtIeKHcjUsO412f221qCqc2cpBDktJiK2EmtkQEV
D95jcdNx6c7wnrIocds/JkSatOzwBq9fRekZDCZnT1BbVMCVfclNL4dX3Nle5pMX7Z1eHydTWMuc
YN9QWw5xICYpKDav8x2L5A21+0hPnvejkAwHAwyN4QFjWRJ1XLZOyUikmJWe38aFkBBqJHkrnt1N
FwMhQFibSjXSUsPeOvE6cdz25NAEQT63nMQG3kVI37YmNWRRSaQYoYvIFGrdC+gH9lZ4O/RtBb34
00ZLMjagKYlacVG3c60VzqHIXN0sxIOeAwPIlZhA1AmiYW95Bf/lVqjh9EJekCjEFoU98Cr189t/
mgmjshDJfcSAhXrY3EFNy3VO8VP0AC/bbyVDD8GQe6zquad3BfoAWOiE8ezN+LbAi3O1855P38oq
8Lh+HT6rcde2x9WeouvTUYBDvjWuBeHqWGdbhGFUtjw5WX3FVZiCyywDhIr+nXt6lBBTuh3mZqGG
xrlUzDXvM7LLckQ2z6MdkOp3vp9tszfeRaVY8yuS2wPphQ9P615AhZYEW1c4HwWKGpGsh2UGx7dZ
VlyRC9JrLnfyyUqAy5mp90ASdPl3sxRRL2oByU67S9TY+CuBo2WfxYMXs2Mb7MUh+EEVuOzPwToj
tjhlxWwILPmUeIbuFEh77HPA3Ud7h2a7GGrPHt/MpTvPZnQ4kCSSDLAis/dT8wvX7ut8Uo131HbQ
n7sYC6VOsHGzEkqVIpOOXV3v/rctb1sUfiKD243XIHRENDy09uHJz5h70EopG3mjV90t1zhptdzU
mWblJJdt5BZSZB/zhp/8TSYmUrHBmZKJVwvEl6Z76+FdIm+/MyIoR/DzmpZIe6M1CmPrZnOJhcky
XSjMJZCAqRmyuRWkc9EZFt/cPH3YOxnGFjUtRt5Iue0S1/+whr4p+5Exd+UY3E/yDsbGhdWjVGmG
sg/0Ez00OLZknzXpknkyToVGSnEFLaNvwTdr+FWH7lsqnlqjUsFumcLixcuCVKBLdBUYkx22/+5m
bz4AuPGmpZ9soFaixdwMNawO/2+/+FXKnCgcXQqAj2boxAp6a6+wAiXsgsYDgP9d5QRT8DFmhJOk
v6S7SlM+KRyKa0x7Ca/2nOQM3SFMUA9hTuXyUdmKppnYDyISmdcjChSKybevu1S1+eoz8c+E3+yN
MGI1fdLnPatiFS1nZYDNq9+vLcUu7To3GSkmLLWoBBfuj4Px2RH9aGR9DUqHB9D411BQQ0ig4pRV
kVTErETraifKDIQto99Gbyh+Uj46kICC+Da7aT9q58hUTFg/Vz8AdZXF7V3oyFd6zAjUmVs1DIQM
v6sY+BM61JStGsMZxF0g+HNYYW7EnoLlGnCjPICutodfSp7LfzRZzg2X7LTH5fgYnwfDjsgvbTII
/8GEJs921KTliHvvqJGGl2H9RHwz0mbd+2qBTOoCgHN81EKwKuWhMU256eklkNopP5WkZdCzBq51
K8OFEM+6TkkEO3VbJ1Ehd/LeIaufKES7QSNPT+kNb35WiCuqhDT/V7oPBn2BIND6cZjHdjpuwCrA
WemtHfbJScaGaekci+uaFIeiSZ4H/UInWX5yxSlRRENHufkJQh5MRmXz6KrqLrwT4c7RIglWIBvk
Q+iUr9rf4XtsxFw6a2RKsPABu4/xYaAidPwWjhuft2TOWQkANW779QU0vC/y86BhjCpP5QNkXMLG
6wNfeS46dl4V/KzOpoMakWAGJxDqkca6jZF7icLrDO91c+rP0Bxj0Mgjcfoe/RNSDzxZsOdehdaB
QTMALQal099I8p3qmCwoIBgplbxiVaqlY1+CdAfQIvsosvziceNXxHkZHUwN5HrdbmLdpKxsciCi
balpwNNSfpQeL+zXGq52O7+pWz3ST4X8wAQJN6pPwA68BW8ouC1ducQkqda5+AvSYTVbVq/tim5Z
xncIML9H4iVOQlHVeBO0wo5UBg0+vZeZPFK/CBzsEWMw2l1OGVrFCNJr20kHh7T661Xygi7EHSpr
JhK8om8pKB3oapHkrduv+daRPhEXuIJT8glaWN2pdKN1C0pBvfyk+oKJHtzkzjqmrAwSCj2DcInT
792zfNYuFT1/fwsGtdO9dmGVvuhgj5ljdnvO9Owv0dt17Tot4TFwRUrSIS5wZpL3MXMxjoQFjI4/
+KBBkW5p7WTBFP2T/pnGgdMjewt5kiTWRXBJEpIyCCej+rb44OOWgkfYokWyuS/wfjmKtfBCTqGl
h8vTEvWGNPtbiHHVxe/oz4E2M3bxgVs4sB45e2kqAmNlgaREMj7vvumuKEG7TZB4FS087muobcde
LnTLCbgvUylsxrjX2RUx6pyqmlFLDrTPVAKjDJDpERzo6W8hOIj/U2GTivYOzTXgN9tQS5rUX1yu
hzkps78Ac1fAEV1r75bdtHm0BTfT5O06XtpLNO4qBSj6H93uJaXRsW+IcJ86Omt+ZKw9NpUJZE5Z
DGMDG0bz2Ejs7YDsNmfL7p2aIjoaYgeA/FYwZ7XmXqaUHiqOV9AIcLkGRancSFAkYkoUVrj7b49U
OEqjCtaYVM4uQcIovLmqFFaPD7hS9Y98hk7ALqi9NC+O/yeH0FdZsrlGiyBqYksrFqKIfhQiUf5O
kfPRIzkQVzwPnfHsbAO+mYY98lNnK7mss3g1TNM3M6NnP/jKz2lOcXyBKX/bXfFQ/dTpyqSGlulu
ifmESkZeHsJalVCOe30fPJzOYpBKh2hxXcXGe742pXFeQssT+uUmJ7DONlNdm92oQhtqSSS/URc8
j2T7617QHEAjFabFK38auOZ6UYJxsBCeGhE1qGEbDBpAqE3bgof3/0ou7hBFi9T8xnXTGe2xg1ja
Zu7dON4QdZ6RA7xoFF0jEi9E+J076thfuh4KJntIPgG1vw6CM//8aPmdDejJGhZ+rqURvjSYb272
MkKHLOOAlvnPiNNwqaFJM7RISvCnM8VQ4qzpiXvQ/gt85Vzz0irURQ4d4rU29mwbNJN+/q6S15XY
tTiMKpBg2JVIbeOiYOHMnmVJrL6pkHHLMqpk2TwrNc4jhY1xdTlBz5vlWAVsbFPcJ9kQtnbGBItB
ijLkNKTrboJk0RFVixRujb1vOLoswePIQBKJ/1ZiOLLa5ft6K37ZXvS8Sw1KlS6JpjlYqOg2PmWq
oOGX3IUwH7YGnN3xxSh7VWIKPQdaJk78Wv+G0mRo2XLtxk5nolAOnOZw+zWHyZ+e9dcSFRU//M8E
wrF23sqdHBX+4gl6vW2fXoTR2+owWkZrSUcs4xfCGdyS2Ph55ndyDRQsnUcizmbWZVkRquFPCwI/
wfVMbQFUWEXOvbNn6RI741gz67Z8UairDxHSrdLlUONSThPEPeo+SdelEiD4PEN7ie7BMkm+fyRK
qEPxS/JcYBo83jFm46Supl8nAf17ZCMPMhK0oImyITo3L1sdSVHpYiFbcRdBu2+pWdOKd1KXjbGV
iUd678h8kswCaoki2xOMMNJ50CbxkV6hJDxJq/sSDweZGotP/VXb/qfFgr+f/S58ZbRv+yDWye2/
6cdBhDMuhjhEHd6e5jvRc3iVsFoRhQYCzTNcax/R4tGL+GhdSzjeAzTr66D3PcD2co9fhKxPKxwp
KFPTTTdIurhHt/IIzBybDNsWhIqjp/+E0rSJuU5XmW7utRJAkuAtGRr1NeXfU0WYAVLGYBd+zxLN
PoH0rj2FOIZVFL3MVxeJASunj2EKqMsZt/a826eNwvjES9GMq0W/Sf17NOcBeCMbpap5KEj7zEcB
zVKtk95Y8BbbuJGb2caJEJZzLgcEg6qE+QrHww1XCujn7FhGX6ujbVZwhe4y9WxSra8C54d6Jj5d
1qTewf1UGOBmmEJvABp4MT/YCXiO8lSPzZXs+wrdaz+j7l6sr/RIbKz/okSwhIq51Zi4YROghct/
CjzkeNpZjKH2/wR9NiZ3U/nReURnyWj7p1OWinqcJ2pDYcQUYTT8SDuz6oeCAckI4Sw0EMku3VYd
opTI90e+lm0cTVmC+Tmg7hq1JzzUqzU60YoWh6Zgq2ok02F1hcDnZLnGyjRt+rx4gK5JLq60hz4O
CiOHrWLQgxfqSb96aSiqvsP/It0Rpbi1VPRk7JpFzbTxGgS5uQSQx1gMEzpEFyqS2kK2B66oFx0I
aRApuXRoEz5NnAgOywv6n73dN8UdZ311t6QPjOWueRwX9scQDuli6bKVZBwPOuTCyd8JJnYLUAQz
9jJmX237hp2+oGrSvnFWL7AsSRCl7J6KwJJ8qxGoNX2kaqvKmXQBDEgDOom4+B/QOnRwp7ZqK3rz
Bmk1hBHQDUzKh8JC6RxWvHPYyjMd95W5y8tghzT2ZHtXvj7wXdoJPzKKadq3/2Uz0wC7UTG+jybc
W/1hgT4m8C15tIYWQ2LathpW4/EZ8J9v1xUdnlH4kqoNK977/t86i1jvlAgoWR18vi0FSx72LcYM
9fALwe5Jqv9mLNiwKKLrO/QB62NMEfjThaZsFDLXSePgbzFVr0QngecTT+EUv1M0RISlbFAap98m
iExzgGgFJMIwcbHcQ4KnOFLdanqie34XLIJK1KsJlCVoWIUXLj1CUg2xAf0wSkJtvAmq++T1ggWl
ppfqtFHz5Qi035/5Ap9gUObZCdyOtWec6qyAlOSM6whhLBJ1sVDZniOz+1FD2Q4WJL8dDDyLNJF0
P7VV0vZd0ZZBG8wc5pGSinP/UHmsoHl8hpmRmMqk4+MPanxTELd+E5UQ9wzPhDCCRmAEx0QbpI5F
37tIvR8jHR0mPplQ0hi+r8COlh6WMckEJeizbOzcrBFtT/NSTj9CKTFXbcHpRhJuncUJAlcqb8no
g0E9kUkLKMIPC2UTCTU3q11HlQ+66D78q+1bRLmGDDsPCgCKgDu9bLBVHQ0aSwd9eosdHVaPAAzu
+4V3y/wVrMNWW49rr5tDMcsPEk3aKHEd6vjEbtAqf1aCc68ZLx/BKXnK8J1NZbYkIPA+ji0V7yQ9
mWAtxFJC7ay7zpw2ZZzD/jGF5yIj3EYnrbMjIoa6lkosi3dt/3eagpA6AN3/PMfF8ifzbuDky2ar
L14aCSqDLkW0bktjf0c8slxGWd6P30pnFxBZd1vyQwQcbTLg5ChkgdAcH9YH4N+hfYH66hBbOT1h
1XYemgLtWVpHpSyyxyBNVkKbTGYpbCEvvEyq8cYhRsRbTdzIahZFUHf0qoWsGjrcw8GNCXL0y8N6
TrQk9ein/tAqCpdz6VZiWruoYmnbXiXtDRWa5JQh91VAAzP3E2Hf5GSmTno4opNDqScxUTNSScTY
bW9ehQS9SKKO2SW9fCssaf32Qd2Harc+4s0iG14+efncWMHPH2hAzpTZFZmOnbObJsBqDLwTr0fD
1Br/qRNLvBbxCHVlC4c3v+jT7j3WR4ZhHdoEaWDWgrTAYnS4OPjIDqOCuhmY1gCTrjU0HnCtyyTt
o53oRI7D02feXbJ3iaTnoIW/JhuBY/3/IVZIVlIUE6KgJz+dwAGFgZhbI33qjNCVH5MscG/BgSoJ
g2DenDsDf6JGUTwaSdGnYz2QvtOvJBO+VgkTwEURYFH7HKy43adRAs1sglzRqajRaGagL96FfhY0
RTNTOuEopnwCwruYIApMD3svSt6KlBFgtxvD12jtgRJgE9oGHs0bI5/w/XJSeaJWCBcopeVePEgi
2osAslLHXizbZmUadhCXXNzkCK5CpUY8GT1TFU6uvttL81HpvHn+6GIgfsiurX7uC8UHpwcMpu+U
1dfQSRa+GjRlRzNhkpiOnHbRjJNhmjUuShjpZdoFTjH/LsqkCBtDmoGBB5768/mNhnWErqXfNt8u
tsXKrFyyE7ll5ep9xATNll+Sn1zd5CXNvP8o5UCr08Ks00dVcK1rLcLTfI4+9yhU3c+azF4tLSar
ClqifDEIu4Cccy3Hh/nhBWSO8nFTkbw0T7SbV4TOTY+5U4BzRr83xlFwDqbMYT9WX7xmgeggOu7I
BC27QVO2Fwci2MyQ5nB0vaYQtUrIj/CfBsTDfL39alzi0fCHEwkwqISJcWsmN8KfYvXF0wO1qWYU
kgnq9N4CoNhdcuOp42abRCW7AZH+Qq+YZKdm6msa3Tm3YipqHhztovoiIUsUk3/kdxt3VLTrNHmX
7KNbLhICghqby5ZHPMJYacUb279cdzutN1WmdsF5FisC0Wj1kagsU1ciYsQp3jFbE5ghrILG6gyh
Xvolg1iIuGFtlwrLCDzFQqMQqnq9RZ7CmRUe48Ef3JcbvScXdbaVZ0XWNHZcefkYQawkfo/u+Gaz
9sYwEwu0peXj0nERRWYA9LOSsgXaKALihIWyK8sQ4gevymWOLn0/sAhRX0dOkeRpR9GfdWuN4xQF
6mKFTF4Qbu5XhPavEo4MVn+v1hivYjuq+WwEly4kxC7lysrZFeSHSuXpTfnZSM4pSOBfGesvfAmm
2lu0RONI/WtDHwOq1W3qBFFS/AVaubx3InDhv6pfnedfmmVJ+0I9yvR9w6KEjF14bmOR7z4jsguP
2luMob163k0J42g43/AsRMTtFJdJXVhoFkJB1cKZ12w478C1ECIMSxQSLjqKcYzSmOUl9K/dz74z
HleCT0AKNOp4TDfdbEqylh/7JI6oku42ecktmYDvOg6cDC8tba35794pRcqWCItXZmB28tLET0V+
dVXbh3M4mbKCLbMH8O+s+1YG4136cb8DNuQWocjtu7Ak42zTSUHP2AS4DIOcWTMWPrvSFxbuLE+9
zWC4oqEDF+qmRFEK8nklB0/ih2E/q1AZphfnvY3GDy7M5m5R1aWzH63U5KvY6lha2JZNdUzNBF9l
k2HjTQhfo05iMvztu+RKRQSMZPlKSUVbVaGWgk5HsB0URN6oXjGzRzzq1pKonnav/L1q9nj9u4BH
G34OQCJBrOsB5Rgp39G7PNmSDnC59ZTMzAw6YKzt0uk6spQHbSq/up9H2+ZzsB2NJOTyVu50RuXG
8+WoEnuujEA5vleajGkluK6oGe2l3qzU14I9tSTBZuPfqE9qkD7gISvJDB8vdqhh5t3MlF+Nkhp3
uz4YphDYemQ2NDG18QWq0RW53CqVLkL4EBPEZ30KgSzzPdrNN0VORsutWtB0DNkfXRSYAPV2oCZj
X4pjaaMiFPy/fY7j0CurAssIYZQGlg42TMbDH+IIVr8G9iMZVpPAaDE1L+n6Ii0UgM0CyLiCQN/e
weYW8k93IehpwWq9/sTaf7vv8ljpEz63i+kR9Xo7kr/rM7UVRLTm7cr7GccoZ7nmIu9ZMj8eE1Ux
baamJdOW6LbIF52e+DIAdxz6QH9Qgh1voIaGp2J60yv5jKDuukIA3hHXkIO5j7/QnXPfukNXXBmE
rROeIvIWWbljtZyD2EQIgkOFg4XQ4DYYrJjJJvHIx0x3GdEgBflFI2MPk5rmtzJZz3nBAbvbWLEj
lSRky9eeyCJtb76taW9ZyDQaxGoOKcLgVe/npGFB3yaTzAuTACF4t2GV8hQQsptgT6zh943/Cd3X
P8L7bcrwDWLy3v/HLAbPslguwRFMP3hR7qR+oAQ/XEGDTrl9Xtjzkn8bTN3LBeU8yLldkZu8ZlMS
DQ0L+rk29hs6nuMACIBgIZZx8OdyeT29M979siYmzxp5YCTim3l59ks5QZokQn8TnGnhJVQ5GnG2
CQn6q9bpBhBRRxwqhPnlRSDGZK4kFNmiprTK4n2b9z2dxOPgGj+NsJJIBw/tl/UeUACgPTOPa5ui
X7Jqv6vTBXJCcnUvJt0Z12X5oLph3tljf/EK3SaxmALqXo/5f6+or2wWsPCBllMZ3VcMcmUF9i1c
t6SB15sgreyxvWJ4wGBmpaOcSLYXCORpnarQdPLSmlavU3UgAq4Y39nN46zYU/S7xQNQ4lAqIsMs
qiN9lnqZmSzR6EugAHx8AFGopDdywXN/YsxVGm1iPhwRrCLXDxDc7TNPS88AKwlP3OMFy8ULkWFD
Zb7EUDlyMymnUIRoSn7OUSMmrGBkktv2VtJSoMsqPwaIBTTF6Hwx2xpUfMoPWj+gajefXkZigIfg
IxvhTXYoqV1A5QZmWvl8Xvh4ac5nX5cx6hiefvWD97xOqdJ2quDoIFROBvKtBJuLPR3LjL5qJvUc
NMa2XhSpDjWCm/Eqo2w9BDiKOzOupjThF9Fg0FyvzZV09yvKhiWCq1CCLdfo+TE2/JPXB1P3aFKD
JBuYnYN0OZ9eue3BF+llFe8PO2JwLnhBxqc7hZYt5EQdiGBxpyE8V5Rlh3QhA8C9yRkpKWgqyrXR
J1yzblGw0xg4utoRjOdkM0dy/G2SDnKlSzM+Ih3b0XeJLma6OZhHnleHATShTDKDc5zoZmeVcG7p
xIt1XxIKn+BCjPLeeniSk7cKe9NkvwCVCjeTumEU/LuwpK81mgDCPVy7Ywp6zTGaMrVAHaA+5joL
DvWqb9q02QEyrbPK5mq8t1hax6LOb3ie4rev/vtY5WMEB7OVK0C1YLgDBdo1/OUdSp/vJE9UmXGM
4paHslHvn5ODszKAjKPMz0jSZ/QsbJdKMbLI6dZtZIP+Z9sHkPrScxkdqlhHBVEDDZoWDQn97jG8
7f6p6JBk2xr2/49HOlvQbCxUZVcN8zxIxkjsW91u4RqS+KW5wVlftQngd2r6tVE5DqjcJ0lbfFpJ
c6Luas9kuHiOPDt70gsosGNyQdvVpx53whepuIu3SZCC5hVp7/RUETbeYkHx/F0OL/uZUC3Q2voN
dsDSq+1Vcy05CVVoOvXQqYvUYy5yMeHyHCHme/FST67cGoY9Ag2ALTbkBjEmLA3IbMQ+6f3kmTe+
+smCwoImGl6SRXe9kIcYAg0WPtzW9GJo4Bs58WrKJuDzgL8RggJ/my+l1Rn6x00/93kVPMsBtikZ
HL2YbEYK/i3gV5wpffgzZ0fX9vsHElhfk+o20yUkVDzWyztiXc50giPTU3B/n6S/3lTMDTyer9+g
yEt5J4UgP+fOrPvh5Y2vIcjdFfNUIgNf/p2tbmd5oWZcqBs193BbVGFB5mwG/GFRDJh+/U15mAhv
VNs2pMOUibkgYwAil8cdVTwUGiBgt+2Sjt0+4583dWd18hB9xWFK50Fp5R4HjN/LPBcMBlRgvUbq
+gcvlVRaZPRgGiAUI0ioh8UzmOLIqL6gxTpe/0iiNgAg8wW/jGE3IuMYysF5CpOahFopMfBA7VjW
pKNyyG2y5PfJY5ql4n4T2+LnKILPPg+bwlSx90GiRuXUwxZb1nVbS5Ml56UnP+d/up+I/fucUy1w
Fo69aNC3m5TsWpLR9kxXM/aAL/1l8K72BnMA4WAvHZLoTVJAoD6I0csMabudK0PccFWsD9N5bknq
pNuJzNbuVSrP33I+g5iDa+awKIv7KF+qkN9EHE0uewl1kJMcwCSV5SgjP9mJAZS2JYe6j0tdxHY4
gE5l+iZKs3a+em4Xu4wmpkNRKq8ynI2kaVuEVSRIbELn0TT7RRtQayb4bAAH7405qBaNgMJzj8LE
CQYa6Jh7LxoKy51JgdaNKezCBAkvyWiXuI8MxSGjgddObFzzq4gSdLdNnYkGUPKbll/Q8/mKmhsy
col5boo0/1LSD6O3kkX+vh+DwSaVaXQcGSD4ntKkf1WRg7aZlqEBgqVUnMWcypkrNLrnykrrcHWL
7tq7oq9VO4FB9leFeH14BkzyPHI8+SkScrMarSMhyIC5vYCCTzmkj8Wz36kvedIBhHSXrjPCBshS
94YWRAWvpHlRrKUIC2qlrOq7TLDu4UmpdfCPL9BN6THqlreVRLLyWec1Yvcv4uieIqOCsQl0SlGV
5vt8km5A3Yhl0dEr8wCwXIH3WTVAStKJfYqCblhBczOmso4Ox8nI1eqVYWz3QgXvQ1SeOoUxU/BE
w5fMhurILsMZfIveuzK91BLOFWnrmbsl3V+fezmvCrOkisw2EJk453/9u+4PSA1yP2OYbFtO0JGT
LEqr+a2P4a5fSh/H8DqhUnk9A+DtTBGHtcT/CNnnj979BiOJNuulqD4bJBSGJR+PujQVEiAOz9ee
KAGwM3b7YXz12wmpAEqMuYhJBx6L+rLOvTq+sd2RILBxYSPxZfej1lirXQEu6eNdCvOJLyymFfhT
eWIiQpIlEWnFsRTxzx9IUMsZlj6WlXCPLH++64rqom5jCwfXsmZ0gkZOjKea7Cadk6CdcpsWrK8t
WXZqNJ9xw8P0agzFxVv2dE0lnJjodbfXdkVSpEHeAtlq6w/OWp7eV/p7hqtmrAEt9JdcOt2twnNy
oMmY1Kd6TCTOiZL07wBf9QxqojTTu0xboeDyZIqRMD5dEm8wJ0gfMtMre+hAYRMJqxNbYMVdblY4
lqFPinHemxT72gO168vS9odD8jPM0cpbdHHGxmBzjrGYEE7wSMl9vhGY74Ux6alhAnNRqpIB5yv2
E1DQc2gAE7Pfr107bptwaAJMmPpQD8m/M7vzW8p3qIeX4Hkqc/2L00pXaL/Vm91UJc9G67P8wecU
tGZrY9/i9xaCUseNeErO4f343nDbyXAB+FUVfG9gkKQ0ATykEExB3/89Uy5SqAXcXuhQ8jm28sEg
/O94zSAtiBtsD+kDGwRnpmeWFzSoJ3xuohzAaX9UQjY1Rw/ZeKbYYKcuqOraYcUS2VQy4jgDKbqq
bf9aSo32rlPCzfE8VioE0d4/bTnf4uwKrcf8ct0S2jWn1LTWYdMWhSkiiIBqIxjx2yxJHjf8haBP
RhuIh9ZViatkDNiBRU7oZ1jpf03PmOB9jz2D5iy1wtxH8eACEKHaHeJS9UsU6SvGjnJRb9JBVuyJ
dD01N9Ha5rwCoS9vwB6+XzUTi44P610VBTiS5lis+7XZAebSRhENOvBrVnNzGIBcon9pdHU428yk
qwdNVkSSogUkpeURMcmzDWfQSLweua1Eq+SRCtyLePHkYZH/5qYwXZA+DnhNHvylQkbWYx8JfB97
YLoio4MfaC9lJ5cjNhmLuyTywxBMb0OnF9z0oJNhO98mBE8V7culfO3R53BmE8uQmTaT1UG6WlfQ
kLvsYK0+mniE7HBCSZQTA+mNXIi10py4f6xVQ+0BvRdxpqIyc/D0n8/Cb6rQTq/k3ugF8zJjaGJV
ffzNxkm+lG43TJ1Ng+7Yx/fW3ARFtFFq452eKi3begOlvfeLh3bCxwZTfoGvq9IytXQyiXBcfw7T
png7muzU6Nr8qs90LCW5kRKlYWAmM1dkDZfkKlE4w74MSTH2Fi2OhzBWGX3dBDdilSIb2jeFA0OA
GenQ5LsJlN+3Sit5MujJOHfdQgzHh7v9IjY9cdF1er13RgMekZ5Ff1n8C1fXwSN2iwqFcDUsRy9w
qlvwHHuBXWzJiW70b2GwABNqsSGyX6cySfZDtSrKcremPoo4lHcMMBfOX4OfsRi7tXEDHmlP9XJK
Vf0wH7QBLzdKg4SwpwLGKnFS20mEBUysE67evwvEpxo0VanEE+IbVILhS4IaV6+yri/CwJD994gF
Iuhj0Z4sq5W39cMtgAZogLxKRRmYUbLp1zOXWMjMKTarYMmfgCCLd2+8A1pWlV6fE5LNBmMh33ni
E4QhYMT1s/zdtz7/eaIJRDN2hl5FxIY6WAf3RRyT7hjBb8uSAE7EHrOxVETtSIX6w30cZYHXmsjh
6GgvJPEfFAkCB9/vEYUIC93mrc1iUS1r6xcR+K+dscgsEYKGJkNe0jHfLyngY53w+JYQ2eD1A1Ej
zLE0c0lTiKxThM7KRL5/RD0pSi8m1EJQjT97diVnGMEP/0tIrzQ7jpg6VgxbEe5YyMPCEMbpnl0C
UwEsyae15TLUUNqsTkigNBq5+uZxu6SFmeZf6FaOAgMhb0wSPqJ7zSXm0RL925kHFhOQ/9PCEb49
ygq8LOXlOlpZGANM/to+avGz8ee/7/4VEmHaYdrfiYF1YzOcbuZOlPDbLTXIVffGMyVbuwNl5jHX
H+7sY/ak/XxzrHsw0/VtS0hAT+1wZ2qsqTPeK+OyjybJQIahwWvo1T/4yea5NrZ2i7enO+4dY067
BQOTX0fubE4e6O9LyuBxVdn8QugKGtcbA0qZeZylbIci/SayQ5X7ATyCcdXGs67sxb2WuvmVCVGG
ugGBe3AEXBpidBnFjgcmSxbR3h4OU/Nnsl2grTxvy1O4jSIMRTFoD2gl8DoQW75r2WWnf+lyF6bM
ePaxODFTmJfPVEqkvZmXH8jEXIvubDxxI+XkXwLiR7eaHFjhzHdqJeowGfxLBhwtGFKW0ltEMVBp
VUGw7hzMNOaNlshbMSHqkG6sQA9NShhu2gpcJPr3L7GFo81f5iUFHaALsOHtWApEOnsT/DaGyRca
6tdLBtyO8QCeOFOeuMN5UcrytjKHagi3xcHQiEc5rY91W+nKSb9j+w49x2q/zGgdaGkXMr7JA0ci
806SIQwzBvwudxGFewGS+GGGUBY2Y+kKxfT7s7eqqFQoyp4Opmz0SNBHPGD+SjnbL6mGk0WPUqfu
RpzDOwqmxZliDublH6fBEAsf9qD5wq7RGlNK5ZaYdrITTT85T+UXxOvW5GLk5XIx9/Jrz9T+un5Q
MXUI0SUjx0aBCJ3x9HOdJbUQYQ1/KcfZ8oJPv708r0XoUg6MAYnGNmJEFs5mxxUWvP2kq7Y1UGcl
F7hd8djPn3iIFFpq/yryztEeA2Ik9XXelq1ZxHIBUc0djZdNk42TeX5f/NNkM4AkyXd9VH2vrQbn
UsbFOCN6afG7js6VgDYhAH935LO173YE4pkn82GC+PsmxhZyvwXKsq/prEUMG4axH6/TbN6OHH6j
v3ngdKgxOMeDaeTjmq2L5Rp8gcFn3D87cD6uX0U7amyg5WABf7CIe2ah87xd4h59XJyMeiHe9OeE
zxZZNAzJ7jHH8KOuCCC0cI9k4RIIg5egb4gzvBM0FqwcK/ZwXYDSicmHJdO5h6Sm6OIANjYkSQZG
+WVBXvzDG2C90QN/sU/ZNNpC4IKXp562MgN+rwV4FBNzL8XvDSYN1d6kcci/iDIyPUHxeVPeFQrk
YFSyhwkrSFyXfT8KRzYRhxq8OUw0CyxX3Q0KT1d8OKoD2ifEW6pTOQDUYs8qHObzbcGBNrGZ25A3
cZEiA+E09Qg5jYdwtJjfj2MtfpY8CoJctmcuUObc/aHWhsxj3rijkjmrz34+4YCnNSvsi9xR01/I
xTrtfYB++3NlKnEL1ae3MfzVE8wIkVyhcFOXC+d/UJ2fNY6D8Jk9fIpF/Hbyq7DzzSGS1WOtgG17
ITiiZgAZiV3fmgeBoSkEtBpLNGZoFRB25pDu6EPfDeen47zg88wlvxl5vfPhWjtrIHV0zoDyIbNa
Vr0X/2IRIRJeF6vDv0SLT9izQNAP2UTq073MO6jwZ6oHlerSgXawSnVFOKrAXZb2MPyTqueDLLhY
VAhCXU27sjMstgLOOVOmPpnyOZaxj7N6JFh+hA6EF9IhRxC+b4BaECs6oc+VlM5QZlOQdLsthWhn
/z1ZYbsz9aFFBFP5gId+RqFKd9V4nhtZiY+UcRVojc6bkUzoFC4BENdMYzPGTgOUrNxtILlytTpp
UV/ISDwjxJ++bI2kpdgbdIctoByYG7q61qTsF3Q2gdhswTtAK24mF3OyrRJNJapFeeAXyGH2tzvF
cUJUvZYcA3oULDJVjnhNHAB8/g/GL4+KV61eN6fj6p4tDhxff8/eVO9/ClQufbyX8zQ/2r9K0qVm
uRsaAWV7xnZ6Su2O+hObWFKc8NaZOSWQwPib3ctA1M2sLbh/0xANHwjkSTRjltN+dalUI+yCbKIf
joTcPiGr6BJIGbzCZ9/aS4nhpBt87Qz5gd+rfW1YFj723QvYPp6PMFxzetkpzABn6kOZN4dfqJqx
duNFriD5vW70zDEYSxpnLhh0CqGV7znJHq3fLVLDhHj5ekPFUIg1ZACdwkRBUG0ibOKu2D+so1Zz
uMCAApX/SxUiO6lDy9As12pSJnKNOEF/nTyva0/nygma6C1dne4r/oNimea26Sh22c3yt93zTeyV
HcwXeDBAyi/K7lIhbtB3b7MBXO5JCkiwZD722FNTA78NPlhSg7PKVQA3FuFjZ8/f3vzWra4AnOM9
aLX0oXve6HU1jcEfhbwMEGb8DFgrmqGWd9+U2brj/LQp+9bISdjCjvh1RkqfZ6bbrabKb+o0lUjB
c9cjzwRJibGZvo7v9bq0GtP+ex4iC9coC6KCS6QIfEgAIU230Z8HD2a/va7MwUf8CQPFc1UK5IA5
s7Y24x8lzVzQTveo9539EB92zbL6k0Cc2GdjST5jXfHzWoPT9CsdPF576ZERCedmH7CkPXEWDM+s
Thwf5/ErVBUlAAKIlLHm8zk7YFMyqJcdS53hGMXNFxuarltbduCVHV5JxXXFRK2P/NIk7mb3delM
CqwU8/s+VZ09/1LTqHELVmdRNEnzWlkVLTTwueVcm942/twCEB+TxPY8fwHu3gYiupJoQ8uXp3HD
KPxB2iuMl36q3UzxvrID6bNvAZMYzDziXO31BFi5MYm3hAfhXF6UIuXeiSOdw0ehj3cO9cP/z8J2
fpUWU1DI9wl2v0HZf63Ne5Q4p3WL9QZi5Lk01/vsQpcolUJKarKr3F/AG3cx0XDcVffytqIQBJmm
BUq/BBSX31NKGTuw/EFNJ5+FxG/fmbal+4cinCoVC00tDWULVY0AIVGiI0NVMj3+MMX/rzIKuLrf
MsN2u4sef72Sxls0VzdfJTmaEM54MHJF+u/5L/pwLACFXAzqtc481Sf8AxKtKVwFXq0cUZtgk3GM
iTLuhcMCmcJd3hiW8No9DFZ2K9+T+z68hl8MASzA+fjxVrgSejRD7Ol760NGL0fCDeXAnWGLY6aG
Ab054vqwOEELUHnCSJinrrxSIwFldq+fr1fxEkTfH/Iio/zalLiwPqHlGb3CBi2qTFhsmNL5GW+0
YMx6DfcQiaMdjf1WCV1JNejkr59pnLB90x2PigV7kE3EcCTsaI2tTUVG2PVIwC7yKmGl50TO8NVn
sPKRG70slnntCjzMjteczww87XHzu/BhjR9E4irFhe4pnO2e3DfEq0gjo1hLF2EESBlLUH9s+Xmx
+vpN7r9AfBIqWnD/czL3960QoUGnuEg0Ool7SVJUinyu0Pl30XVMNGH7VYEJMw6FbIzeQNTNPoRA
eI3KfXGFPk1KFMeSFrlTQ5tKWwhbNwIGoX/wqu1SYi8L2Dus3VCa8GEN0DdOBQ0lB0SmazX3PBVt
/TKQtu0ez1tlzu4GTvUp7HWGNsanTfCSVbu+11qVbsdZBBO57XWyG+OHLKy9/DKX1wg45O2sVPkF
U47KfCDs8Fi+y9BQ+U8c/I1MO69sHco5f8mNh3HQwIxl1GBxqHTrDE/EBnJjxBc4LKTMDoMDw4YE
txp+fhaVtN0aAW8cm7kXD4i/GwX/E078uwx2YUrJhAbqm42QKk2gwiL2ha8pFpznlXgRJthqt+S7
tnRel7pUholjpNMivN9S7GT5RVN5b8T2E2it62EujDmrHlvY3PTc+pcOscBUm17Wa33Tkz+jCRiD
eE1egkL8gegCEzXAW80ANRZKkyWzrx2JgxRYRolAXN5n6HugjC0MaaEhMnYuylZtdKfXnAz9nBO9
6ujO3BYNXydzc5v2IrDJp14KB2yny2gBiBDIaM7go0FY8liZnzj5JIEn5qcRDx2rDYJ1965rcv1a
MAV8Daqn2jeuFvDRnmNeyKZdSfIIEBy3EcxESzBMGqChFcnvscqPnfeNYdYf8wKX678MQ3VB0MD+
fAQvwqRoqFWKGhx3Vv4LB52+uqeM/mj5TDfrrCnt5a2TnpX5emxY6/yDQMKsu+RArFAb0IljTkQQ
tzMuqqzxOR8nmOy8sLf0OhhNjJ/yUIA1jZaEhR8Hk97YTiMjrsQznDuF+jTNaSv0zd60EoXQv2iV
wciY1cZacc9t4NJyNgnOLgPqdQwtdmhz8h7r+lMjakEgSXmEIRqwUuAgC1A1uLIQmKyOZiiYETJR
ClC9O3LEBa8TTs1uQfjX4vJE5l4XIW3xLDfrNGphu5AGAM7ZX66KNCSIWmgm/TiszZKB/tq20GWy
ZBYeTC+piPGJdRS+bhS95c75C5CDm0Gr5G8BG1OOvckNGbhpTJThFq+NYzk82/7zU/DVlsCcb4fK
ixrSS0M2IP1m4BMOKV+sqmuLVBXj6XSQCe4Oiasu/s+N7bRxrQg2kpqY6LxnNw90JlLxNslqcEw6
IB4R81q0O7lLuwKnldQ3BU7W2Fpfelb41Kpc7L8Z9VCO/hUxJafEDt7M6abyYdBF1XHEgmtqSjVx
9pPZ+Dwxsxr1OLQdMXlz6KqhBCZZ5kovhnYxruyYsbDIrIhJdZ2s9R8IB2NHSuPubDZKK5dBHwzq
7a3NauPVvRua5Sbw9WQptFeBq1EVLQcjOzEHDCfuG1EDafODNuYo7mA1i4YCb34L/diS57EsNAEp
tCc1njkOvdW4riRxBg4YzWep4ofGk5LV7SxT3YS1aPWII3O+yzEv2VhsvBqZnqcx8LfG8uyQYUl0
dxuKu8Z1baVtLfUkFjDVWl3jaNjII2nSoFt4bmRWTQA2VOYZgbqnjrzxrs48qeTvRpmD44ApN0T4
xG/ugl4nQRMptRLL3uqAwCuBZgaYx8XLd3Sp4DBIO+LJgM7jjUBB8VqmIswKMrPd4pssNVrsJU7y
2wuzeoZBcB0zvRAfv3+QpFgWGo8oeE4y4rR6dkFcg72tX+lWyx3uI/cFv+D2eyAcP5IMZzxTtDB2
zvWnXYGgFsCgteNJVn5aKeOGtF+VhepoWZyoQm21pq5tSpPbNqEOYC1ZiFk5x0wGEqTxOzfRD3lL
cRcoEFrujeA1spbXu8MHfWk2obHO1fQEDKw+Grvm27EaoVhiCChYeo6BWAiqnTR2WJGD4lcBv/71
j9FOiNJxrginll1H2TxyIuLxDxpWpZZgyzIlJIMNAryxVeCFWeUgc1rT9ZR7BHt3HP1iBznZ+95i
KWyWahxa2A4jrUO/ZVUX0CDB5eBTHcrB0ryevJIz904mpDW3Wd2YHObxum0qoeMbNpWFTsEcciVk
U6Se2JGYTf2e2CSjOHPOq6hKo7nQ4NmEq8m2LIKLyFPIkEgLhbSjMCPKGEamtmc8KxDvUpplt3rJ
ASIXbxayNz769NirzgZdNJouA38UnYGHOtO5OYsOKyY/3/U+l/WlkfKo4sjt4JpQJbQcP6U5B/fO
S6qnoWaVjGVXteSYCdF8QfzWstu6BwMI2sPCl5eL48DJYvIkYtX89tWD3+Sgqq8O4PBc7CyyABGy
bzBwN2VhCVkjRdEvKtvMhR+6rjJ1BtWgaX00XvKCvD2KUArn1FzQ0FVWaZ9tFcJv9JiKvqz+pdCW
n0F/QiYaXJeBLESyHSBM19Etx/rK2JEyvQMaYe8cJfGBMcz1liPKFkpezhgbeQOsGkQ9pWCcPeZ6
kNbwFM0omxLZ/iuOdV94z8m+idTb5E0doM+XJ1yHshdQCNnXbGl4o8JigjO6POWy1yiEo2y3zd3q
2T18JoIU5k+NJ8QbkSrjjUv34Qj334lEw8PEkxhtbdQ8fviC5aKL5i0gs7ce1OijL6VVeawyYD3p
6CfRQXEtY+jpknf83zsUj2nlp+OqxzR7WE8r7I6dULRtzFRKrzPP7T6xB0AdXGVqatR/rFriKub+
5GFI0KVUrv2Gmte7NrzIHopsMnZ5yOvdSueUU3Msy6SfDBc3P2u7jO3shb8HeX4xg7COnT5Etfaq
15Yw8FvT1Zz14ATwNfN6K7j1ywugZYnFPp8J0bUkcNLj6MJoHGY86UOHhPqweBOJDj0cfvnm7vFV
VPJpkTIdPn+IiYr/xXlA11BSGbmVe8DcIPMU5bY/ktbkg5Wo0dveuEqSwxnICYaGS1/1DR64Wmlj
8yelTTCSXZPpONaH+R0byLLVX5YtHNSW9TuXOqYGaieXNmM5iidB3jkGtuf6EMnjVuRVYaOL1cXE
cyH/okXisXIxWbRhSdDB7CzTxGJYzHGc36peeJOYyYdaiIH39eytFO6tm0CJ3+eKqQuhq6XribPZ
W98un9hAjWSLpJ/XlLcqzCvRaPc3OPczYMdv+zRkhoAwBKQXXH8bwZXd9hLjmoBwAlkAldu/t5vR
Kip+WkU7qPS/TUGj/N0vR8fxtGy5gY1g06luVtFGDuhA9s/a4q1vIeFJtNkiTo9vG3f3BqI3poLq
cbtnNjfLAbl0OPPoO8ugqb1qs7xByg92Xqow3SnA2oW0KNZsv2CBawa2MEk31vJm6JPRCSFiIMdf
Esq+pbC+5SdMMSVkgPI6/Ch+73uX8CQvYoSLuY6iKg7xhHCu+3TWx3UqNYDTJXzHS4s3/752MMjV
C8cqhxIxWcmHKBS3nu+sS95dKMxU7Z8q026S2xlKw1YC2KpwtEKo6zPwe2My07FnUcJ2QUtwnVzT
tw2YQh7YCBWXWOOs8/kVG/yThjwvYR+1TOOFuMWqG+oatA4BvU8xFRmXPwkLQgUq98H/3qK4y/Pt
rGdvjsAtyEr698TOye0OL3///Z9Z1y/iWSSW1F96PNZUeaYj2Qg/bDn+ID0PcBU80Pjz3GpABx5b
SQh0eGeK69HwZXXk0+KJlJJkKpRQu1JHoXwm1sZfPoUgr5xcET1exs+OvAEVEYq5ZEpC2kpexwQT
aJ3Obaj09XZxhtMKZgHM+xbTZHXg/MlUbvlxtZ6/3bG9kIXVRCEuIQB9UXkkX1vrzh5ke1EqH4JI
u4o6TCF8WWd+y7GPKcUtwXV67pt68mkf87WT2zmSmDC3UyIKlYY8dPaqNJhthamIDmuMeUfNGxi8
+rJ95Zc54S0GNn0fOUfT53PkaHZ2K40OE+dc+sWgbj5nc3kCaG/Q4g1x4+nr9582V4DJYhvFQIa4
sCV1tu/Pg+pYc8S7tjVFwcymQplIiga1D7lYILA98Mmrpkep0nGuXVDti23dSyuJ0OXrJrz1SfhY
VEXgvzWVq+998MZd4L+ccPHqkSStCjVP0VLKxhtQdJF7JvUVqJOvdWWyS82+TPO4iLZnft/uOyth
lqht4gn1TIn/LWB8sR3JWrfIKVxN8EScxTCudyZ7t+wJRsX/oalzXFd3XvyY/TyuzF77Nsqk198C
qtgNt0huOipTj8KR1M7uyn1gvWOYnGZJ7ZcOGG0zFWQKKyCbFWkumDksB0ijgmNFVtk0ZAUyUjw+
tl1PrHjakU+Mncj3jwmKV0Pqa3EI9hCcNnNU2JZCX/2GTrXUzVAggAR0aZ2KFhS2totwIwp0b7Wm
1exYznR6t9wGtggP7IRpQVKSyIYAhnzp6wyut3+HSYICAsLk8VoN4g/ec56hOh91dCJxcG3d/5L8
cU+81vgi+yZ/yNf7fsWuZf0hI7Dx3b9ELoBMsZcbX7tTtGpNS2csfKtCVha2rmfW78lvR578BqkS
oYQ9f3FaKEKm1jYXKUW+5tJsO7NlTsNi2v4AkxiX+NWm283Ux1Zwz2ymcBm8W3os8rNqS1IZrGnV
PcK+qbslB+FGh/NOpvXlS/sSV5I47sU6VazGWxi+De68mfOQwkKyclQcvnGB6g8mdIYK/PTvqueB
7J5FtbDY0N12Dc1nDbWe2KONQcpi9P+TGxL69A9BrhYOvHgcuVQQl2ocfIv/Z2RLhDxM5XBD1jrA
DMSqftiFikWuamygaHm4X+Z+abHj+l3uVz8soHCT2XyDL1/8Ify53qbo3UxunACmvAeAzQmysSqq
o/mkne1CPMsLjN4wxhYEI0IH1+eRV+xqIBYDRmZdngoCgPx+k7XZV0kk0HTYTJ0Qe6iX/v65fWPn
Mm5FP/zvK3i+gYBnOXJ0JMazqmm9hubthq8QFhTII1qGAUlwenAlO4uclLbqZweCI3zFFHT8hLak
fmmAXxjnHUd5Oc5ONTnx6UDFdbXwgdZobEBauLh68YdRd4jfsxAYsaFQk0wNO2ktFXCQBRmW+KoR
sybQAEWJQYhICzpiKuk5SEThm11ggjp0qSvCYxhFj95EyrMz8TkeUnf760UCVs1IJSBPGTHT0bYm
TIlFLPOaWtDAwZvlKE/BAGCGD3e6IMaP+kgx8f5SQ9RPIHyDqs7F3v986aiC9pD8kZSxHCEzq4x+
VH6Zp+/JOlcPSaX+O9FRyD6mCmrDg3lZhNZNtOhCm18WHL4Vtv1oqdZqy9z8V5JV/dDsbeKcqdDt
dxiUXUl3cVkW3QII9Fhp5gPBfwrLLaRXqWNUDiwperiBDvm2fGB1z47C6eL7aujrPAoZxoMWmxHu
+XCsnJcKHQPsp4jEsrEblr3FtlC+ZT2AeWEnk+nnIi3LzlHQVZVcPf30BZKvcqMIt7UQ8edvPC67
3FY7ZJgPueF5op11DXIISR/KzIKf1cjc9FcQcrv3PpJ2yc6u+HjnGkfRc+isNodN66KxoLez8DjW
r7cAJuegAI6XI92J2d2+tThsxFeoY/03Cx9P/BBdOXsRc/zIVJFBoEiiMEkKuaFmG+DXEdXRwDS3
PWL/4HPe3SNneN5dAjGeO0CK1i44haPDljf4R5OSC3GJadh1mhkC8/4LK3hY929iaV3pnF+BRXJE
wSCXkv8wur9x41ArDlWJK8nCtGIkP1z4H3a3MdgWBUxNC3t+V9jaRGJrfp/2Iw9iUbLY9hpv8xVD
j7ov/A4vTo24x+2C1hcBU+AzaSkbu+NV6RkV9He5crnJN4DxBWFft4E41WwKhttQMFIpu1KIik76
DAEGiewJ6AXaVEJPGpPx4+PW9h8l8HH0oHcTOPeIW9JKA+KBNWkh2zpf3LNTB8caoFWFw+U2cSPq
rkRaCAeks+QKWJaAYIuwfxxWzG/T2ssed2y51+PgLmCCryJ4tLPbmUaDftd+O3SzuEZLPQQE2Mpq
i/eVbUOHAdCpxKktXTHhifphsb8KljVjRCLnZvHDB6UENFkXcJetP1RDpvSLvaOUPLWZ4wVLlHoA
2/Ie0Yi6jkCAZV1MsLLKd99WptDyGKG12GwCfwOIZi+DZmKGUX2deWfXLKptsADPeKVQ3er9hhYT
rteTkGvl1T4nlVxdKfBsRKzfx5VH6XcYheVaPfAmVZMyacnDNj46nScUkirPqk1PJ3s8sKE9lUOr
jLgInrSpyhcB8MrsPkTiUZrXnXoR/RYLSvSgttdmgEoQR+JvVnyi6KwzC3+T6uwAmz/OUQMNRbjp
eYS7QjY6bbVQXDmtVYENZ0RuU94cHCYuQvptszDg8aEqQIuZk4cfUy89WMvUmH3nKIdaVNbZdIKQ
R7hTRTxC/JPNoVYfZs0vnNdDega1ZY2LN4vXPQ/NzjVZJ0ifHL2UUzIY2Inhn0mSmb8Z1t3noN2z
zPYZsczieI/eee2d4avGX47RPfZuhWyuTKX1vhgZAANo2tUxklNj9NCYHJ8sZxNHQ8xmHQS9TaPH
XMDwzuEjxJ7WM3dqVIvvzN4dGeWHbbdDvLudXjj1ok26NBIwuYNtektgDuR4qTu8ghluJfur5C2K
iD/+P4ZKRTzkTObJEo0fK2gnzugh59wTknz+0utOZet9DwjVQ6Xhz5jCR0rJ7vDcC2N6ZxlcRiNg
MLVfxDoEBqKr/BJvet+bEL8OrxLgLc2UDSL1r579VWCoDlkhZ6cwW2i47eOK7HEtN0bqfWp+JVVY
ozsnSwNtTzOSZQBr8D9024x0xFMUbi+enhzG0kmbxLPiA0KrkOwaKEd2o3DHKoAdNJCKUQEIbo6g
Zi8x/xcdGkxIGpJ/8uls/XkAgdLDDGuSi3dPr//hmYkROqhUgDIFzofALYd1Q0v+nsCWzKeLvKFu
btNJWUO+IxIUJsqsiDNoQYQBj2l2JzdsJwgKqJM35VQV2dQ7uD9LKLjjUs7hBjmk8uoT4HMP0fw0
AqlXexlsp9rfX/zGaXhwlW8ctPUIZJaf2IfMT4IRU5C9zJjF6iM8wZkGpblP+U1Kvw5Gdn4EugkE
0xIzXOsFK7w6dFImAVbGOQW7q50VDILNIG8CaRMksPwlRISGhzqe03Ab4gefsCJ5DxvuueAJjZsC
DjvXruLOCb8ZHNZ4n60sPAUjwuZ46s3quzZGlyEQoU6VMM8++ErNgAwrkja8EHa0xVtR18dByfFq
YN2QUX5L9hQ/VA7clI68/KW3G10RN59Fpueno/6v18ETaoa+7OtYGeYxYmL/3O7/ND8az17iP+pk
labzXtuJEZEqqYJCc/w37JFbT/qhr/QrA8R25Qv8VT/0i9OH7i/HQksDH/ckUaMyhuFusutpmarR
6AaUGxmyvAquF096K7q5sOtmxOi5g0giUGCIPh8FmYwPeI1gxYLDOygyK3VMFzYijbn1KJ86qrYA
c/w+eCNL8uS+ztQNZrH4IiYAZHuo0n0+6vH5NLpQk8U1SghJ0Lj6YLL+eJQa7UXTxZMJ4jXmBMIj
bFkhuKvqeeSQE1/a8hFXp9BoKpIFCu+Gv7tb9B1/dGcY9NvcI3ZNVm182zIzlo3mJgf6crTc10pr
YPefKlL3oDfvGmYu7JEW37sp9dEeCv4ogiXxYnHqKzw1OQiln7cq7I9oTiz7Y0GxJ3D7xBBq48O/
JX6RAM0pIID3fvTM2eXQPrK0OJA0I20/IbG6u+o+hGELkjXjNamTm5+xNNdJFt1IF0VHi4co6Zi8
5GADgfctBBeV0WpwWLY/1Dt/Cvkm15zQsWpexB2x1jIHAzfUdgs/YVFvUU00HL/rJ97SBjDRBZz2
c6eJdPyClmKbytmlzsfudTCjnIIRHvAT5kHKulH4124PsQySYTGWF+vv7UE8+otVhAWBVwm+ZeR3
t0jFk5hndMFYPliWk6n/Jy1VC6qvTHPXVu6rRAtDi4rN1Y+eV70vGQFNb74oNl5MIjvYmXiV+z31
Dv/5KRJzM1MTI2H86P2+MvF0gldXNRanhYYnABzeRT4gWfy+Yy1caPJMAn1TddMm5CPwKaOJOXW5
bF6N06kxAt21qzKdp/ha8i04/57/uXkdo/48IhRvq+kt1go5sfDa2GOAKP2WJOkbAdxhdxTyvuqv
qc0ISZlC0/rKCSlEz0E8nr8oXb3GjYsRf/ocsGc//GwZO56Jmlac0By2ddJgOx6eYaxODK8NAte1
dbP7S5fzp1GU1rYQPL84FwPbwZ6tnjTUj8rxwqSvga3folMr7Q/s8k0ThZ7v6aiHVU36/p7oSR4b
jxoaVdvuakId7I5DXo4k5r29w260iqUc3/w/x/Ss5ojNv0rYkHqxu8G3R+6THVDoQTiadFSFRUdp
35BDyZ6/J/7g6ex6YGO8PKmGx6NbnLXxFohdHQ5tz4/o/paZRQJ6RephMyoZA60QB7lodnyXn73d
cQRXRaEJEIlBOzQrJUWFFo7xb/r9y7Xr36+vWMCz7AR6iwFxzJEqHMBwEYsFPEZdP0g5OmbkzeEf
+yG9plLHthbJAZNKutfz9+r9XiYiWZo9c7H6U+zW/hLaEl6+g7+GyfT+F3QTAxUium/HG+WDwdfX
gsC/LqHDYMEsCbkXJVxN8Xne61rIMGz5Vem4plzz3zb418rzcpxNnNJoLYOq6M968n781u0QrY+G
hMaF0RwWllHCitrkqqFDX2k0TwB2ko82Tsp8yDctHV+Y9ffv4EaMhkaVyR4nP0Us+pVZYpGavEB/
YQlbINbyzUfQAhhs7c7B6I3znVtllRATr9aGiyXNNnGwGzyEaARF7B5eokb9uqIpeWqbK4c+Qemu
6UJmA4kYA5QT+DZeEXdOd6Hb+WjBVgPM1kYtbTG3/iZMZF1lyDn/q2Ode8lAv0sdJqDm65MOSI/a
8itvlxvF7ejMe/NlfHCMO3cnP38rJ5bVlhcxXheoMGx7VNrgoJzS2uzULH9n75K+0ojNCei9TIZt
PgzodYBOGqnRHDzoVOtX+jLcqtRQlhjnnUaGYTr7sTv+sNxWLtO/AIIu+5/oFGfD8+rtDFKEjgdi
SwP5LkZJR2Ps56dezcrwq2vO3jiJGSWbT9XFwxab0ia1fSL7NLljKfYCzLoOCExL4Q0LazAjLQ6L
UJS8e4KS2rmLcLipCCy62DTl2FW1RpgJte4QJOiv22we4/sLDGPGl1NSvvhznJnEmBnmROPhGJXW
6dArE2hk5K3DqCfYaN4X5G3bL/mXZYSH7LJebJyrwiAZjvMKh1gMesGSW9d3JzKSPEa4WhT5+DS4
U7MI7apuqYJb5rQbOhjfvUR3CGGWcxR1s8f+WMp0CqHLWaElaTnWobyJATM8P9kemphPKaKFDGD0
ze1oEu99YX9908vK6Oabn1J34O3CtSLIaJFloMYD8Tp7zWZiuF5PPFwgtfVFCWwxPCUi4/4UGsOX
z92u4T1DfxV59XmnwuvQ56zmwXFsuJW21hQQEbcChepHBZMKQNRWJigbFAKYFK9grjN0Mub1CeGa
1vHLTYhV5Vj0v/Gwm4lmWfb59Vjnwci9jm82MfxEd2kHyKfU/JpgwaPmUg9d35Lco6/bV9ykAm6I
gIv63ce/z8r29pVfERRlUhKK6ngV0l4ZkMjeifdBK4gG5GBWOi3oDlZ47CyMm4slJ/p6RlDRdcBa
RdDOCBMANRI1cTAFO+dHQyAjP8umYbUG3oDtpdtEy7kqx+5kXCiIbXEifro2pIdmkXTlJZ4rcvnP
Ae3yUV2Lt8mD7h1E6+qsO4WhPGoHI7AyISDWDW9IavHq5JW9IbDNUsZHEcTfALhCduzKDNfMQ8qQ
Aakq0QJpBPMYElPkL2ZxNrRvt7POuUjnhdiFHq9K2bjKEy+HGmq5sFnIU3lCtbUs1f7H2rNGtWQd
7KBgXnmZvgWZNQDMMyNOwnrtNRgCQXwfAi+jumalu231vm1ejqpEtw6c1o5YaP5ALmVIHgVw5vpf
fppBpQq0XBuWTyt/ahMfFotRJkzsEUGk1In82E8ORjXsqwq9KG1TPJiU6jL7pNidmUn7fjIk6XVt
2zQAXjLieQyhkWRrJGev57bNfDbbeII8/2JGmUBAkM4IqbgW5iWpiUCQvXvEwGhdbpn9rvZckmbO
/SVtk/Euz1uCGHJEXGUDEWsS5z3i1D878hVl/O48gg028EDR9G0EWkOqKduTMqA4cGj9lOKK+hvz
f5fEkVWkUVFkdXQdfvaCVA3nvtwpkLG7KxXuRSARN1e0DtCBAvgr56HmWtD1Ca2mbBDgXu9CVgB4
Bd/qguSHadL+7z7lWZK2SNaBjagRx1vjpCCWxmF7DoNvyujvJgajZPT8/+TT29rjP6gg5uZEVT0t
eGMIZgmAvYJbaX9W/VfdlfdNyJnnxm3AmChc0Q2S7IhWrK84zdqc51gMTk8srklZyGcYnLaBVC4B
1HguTj8Yzk2d0MRHXY706KR8v1texXKrDeulqdqX90o06YogxU/LVzy0gEGN1uiIO3YmuKz7npF4
nDG2XHHnsexC/t6+v9HepJPEkWwxXq/peeu8YzUYPNIpzk1NOAqTaysBxCy0YcYNqOcSop+aWxAL
y963Uh8v5sj9yqclHJml1JPE1kJOxzlMcxKm2F6PMPomnh9seSzuvFjKEH9PYI9jLB5w9bhaKbTx
yHLkhSGksX1sQn/NwndlioTTOL+wXFcO4bjIWRuicj+l1vV4Sg3tpyZmcfcTIHyqx6KLncABZXIu
/wj74lNs7/YZuYcHUR6zTXfz/dPyi/OPPnN0vEF7aMH4wY2csS6UTrLU9z7p2n3krcjAmO5CWhpY
hWj0N8QgkdSfe1OUwbROGlvHMJgKMQrzAiHzjEyRIbhQ+FwfTsQFoLss/T19+nd3f+2xtN/KpyZ4
qrfXV8XkNrpgZ5ZaGiqmg0Pl12E/DTDrTPgW+Y5C/7XQvI32326cESrVYo3Cp+6mzPNa5HT6X7eE
ARv8Mmk1N5PXL4CS15JScwq2O2xSqa9vG1G7bOIlbj5wQo9CCAvGpsYtpwOK/qgjB95eRlo0bcOi
Hmd2ISuZfy0c3+9Mf+3MLxjBTnteWWPkm1rYwvWdZa+9yfO3p44zUSwebjw3vmU/0lA6ry8kEFSc
xF98s2akslIBjXMWwfbFGopEesi3HIBBcAxgKVuQnmYH7s9a1dCF8HonT2t8DwNXa3RDRiGre1xA
GS2TQUJizwWqCav3jnJDA625thifK6Ey4psdiQxblLJA3g7Ghkc2h9/yzHocPRNFmJdsPr1kNhgC
hWEBshVTUH9w9JWSF1wfRC1u0/2sk53jQ1S5kj/h/lNlA6RtOe9MCSSPN8zbkUmTHar3vMeief5h
wJ2Y13U7dL0nKQE5MQ0FSXOMpy++bZSsdNp3uzWzhxmoJZ8iSiUpyjIH4eeMvu5c4N0sfxCzoy5N
9MH6k2s7kEfXPO/PpaEmovw2prgtuV/B8gGyg8PBgCUkLKbnm5s0FfXGYE0+3+a3YqvXWLZVE6ku
QXDbCXGjEkA/Ze7DIZWRPgNJpho7hxYlCnrwiMO3OcV7KKT3WwneKiZvDO48EH+Se1bRvKi9cSLB
8tQp2abbHoKIRwbqiY9SlO5IcuWR8ExpJgZsaYdBlWz6vkK+ARVLb2KcTKGcEeewT3hNC5Lagh7Y
vBz4I9aJ/wRolLz+1vjR0nTz9ClCUDV4u8ad/CuwEz3epSlSw1WEyxmC9MZQ8ESRZBOjuB66EcUr
4cBJe4PO8EYU1QsxbkdAakCAxA8vFWIVkEXxvFe2Y3MIRkpY/pPtIbRsHTXb3nIcYcFUk26IwU2q
6n2nplY0ZEB64uzOjioGG2lYXlqLw6anseHssNeM/3IANiblW9WQAj0UBp+MiZc/6LTLcBbn+gNf
7C6V/WnO4FBdc9J3QwytiljjvvfYWJWMtpr2/9poCbcKBGeQ05VGG/P/BgaMpi2Cc6UtF+AnpA7y
ro6vTZNijY2+b5k5eqd+N+1/pOK/OXndTlz/0E4sSGYvQMXL+FADcyI4kBDSwzNVYsokCdF/78/T
KYdik2TNyYbKBFUyS3yPOD0PPg5cpu9T4tmnLitz5tfGbNPjxea3zwIEd6ShF1zUHif+YocUVcEI
n4TlP5DGP7cYZkfdhDrTl9M9+IbN+e8XoZl0+o/TyAcQMwEqsuwH91O7mJGb3nYNvdC1jsJbUXU+
1BffgdyraaYYdNkxQL2lhlaxrvqMrZnD3cGz7CMnNNYegd6aUNOwUHbsCZVw9GnkN2esudy34atB
R6TH+wUrM2r90kfPvCy/hDYdi6qmcZkz4tQWW7R6cch5eEDWFYxjyzrYgO5G2k/QeYQA63eBvRYV
IyGjJhAmLux6MeC0A+vJE0HwdyWldsvmyqooJ5jNHfIUIKHDelu+nr5OFR8TiJFvXzMfFGmARveg
ChrGrmDxyzck8kHK28LePrbT17x17dcoe9T6HJ2U7NoZ6iFbXoyx33GVjMDsOHvQutYAPjHR/6lL
bxIxd+H1s3AitnjWUjpv+HAPgiMwEQ4/f0GWgCv3xCkCuiMUbuukE8xNmllrWj1/Z2KZsrjj84nL
oaxKWid98MIvi9A6NqZzOlLbvod7bX65H5GeU4BcMWZ6+gQ2KSm84qR1ilVtKt/N+YxGXb9k1vfH
RSt7cvUAgNhsiKh3Lo3XEm1GByb+L9c52UhsHp3C7PbAVf1AOUWCD26rM1UJRSvRfznWuRyMnlgs
fuCMgrEHZO0dafltB7OQXYO7teKY2m0d63kT0vJ4Eo/9xEJzcBiT/nf26KUjSb9TJuKjs5Uwb2hl
kHe2iJuStq/KbboPVBv0SExaYZ+KucrjTVKH3i8lauV0LvtXyXeZQn20pNTfVMxPbl6T3NEDCKtH
J85yuopNVVztJNVYsmhTkiWACmpJGFxjGrdT1jnr70E9cIqs56p0Y23y4/qXfIRWGHeT9aheQ3mE
bmt1RA0BEPTD6SmLpPzR+NRuMs5cn4x0wt8rV8ujhZ+YjLrfhi4xzYyE1qIIME+kvsklbFPIkYLE
klqu0PJO/MN/D3eBFlrmIof+PR8B4be9CuceUEgJF+HBraMhr7XXHjfTAE3Jtm8WIBNfcvxQbRjH
5YWR6nvnrWGSjyWU9UCmvV9M2Juge4MzFDZJaC06YAX/Sf23ugO4N7JN3xR1NtGqDrFE89IeA7pr
gaWU5sknYXtY5gluzKPTqD0SqSKv9EOW/X/ViK0q02AmiCu0i4n2bp2RVAG6BNwxcH1H4YUay5PC
panmMiYzK8lZqaPykOa6bPwO+6Qp5lsFb2OYCwIg2ncfiI7RC1uj24wlSTotCmcWzvAvXmX1E/U+
pDRMv5iPXuOKEVCHFWR1Rr9LHswnFBJuEVuYVNh6iN8OynR9tZSCIJjge5ZPiHFOsHkUiDbIXZJo
CyYerHsr5VDwzup8WG5kDylnx4SqYCP64CIYS2q1MPVQp/NrWfLIkYQ/MOLpHGng51sa/Rg6I39L
c+IXqQg3ixuqDUaP8eBNZ7rT4y1U04FolA2Ox4crf2GhAe/XY0GvCLZmTjLl606GM8UnuLk6BYWu
wh/qo/jDDOWFfWuVpKVREQayFOVdx6bIc51OeykXwCjSQWEUS84HnfOYCufNekabdQtMa0WdZYEJ
YldPMBGiE40RpMqrzpI8EIQkvkOzOs+prdxJyCzvoWj2GLzAkxlie/QZfFmA7aAefZulMezkNsR3
eNwdoxXJ/wT8fu0Iyj2HR9ieMGmZ8/8XoylMpgym9pKsLcLouDYEpANVZMYrd150NdqDiWSIKSyA
lmDGKIGYsraFa6anJfKgwfZ/xpbdVcQRnwZ9hqghiGE8V8jHc0tldGXdk087EfdO4rKXSVkf3n6c
Sough3334Ti4uG6LAcnDpAZvd35s4yPCVBpiylHY1S8S5l4BqMSPs47n+U1UdvhRNkGExgLtsQw6
eZC4ZLVgCfgt+vdpTAPaU034LK9FD+j9kl3JqrJ4mBwvS/8cRj0NPGVV3fC9C8bSf22/5Kh4ESzA
BILHIJf5N5+yUeOmHvn3BxTVvnQws9ZIYpJNatR0SgCXFzER2uCbC5Q29Bv4rlD2wU9afjMRyFBm
wW+7EC652fUNpsza768/Z/7x8HkygihMuRSn/oHV53W7PiaJXeyyqvpquJ66kv/IfTK4Be/OF1Yp
9nPkvlr5eoaE1R4cNn8n1buUtMPHqcK4FTBwX3EI8AiXTlPYxLPo+tZHDjdakjx4q0b93lBoxrjp
xvH4JwsYWDnPtOb/oYkFbNkKz6OpEGSakoSJ5MHiaccIivWVcbzO94Fhrc4ad4tfmD8MMk9XBSrz
0w6sqlP4dTLw0Si5AYpm1eSnet6blLuZPbk9fyxl/58pYHnaSTCrYOf1EORa5iPK2CGnI8HgPcYO
nzhHHAzUB74HpnhpBlkXAPuK0GdE1Y85/T8EiKyqquqiYgeLOccog5lIRDmwJ1hGeFis0IO2eO1S
6WddB1BjaPh9eR65aAVkIoXGv6xxyXv0zyb5/k5QiKKaeAEkfN029iulek7LBFpZoX/DwPhi/pJa
Kth/QYK3SLy5wlBYQCf0eSOFJEnRdlTvKd7AppNxfIotsA1ZMq3jzaL5GSeJV7iIXENKcmc7w3bc
uKnNEfmRZPI2lzc5pWOS+1LEtg5Gm4axzvKy2j1GQx/4uZ38hvtwdpHO6ZrFwDD5lB9nOKLNdeNK
YFMtLk0bKYfx3VycTejiUh2uSoNcTo6rxtY2dsc1016trEOJ5V3hM6433y4gGQDfR6ucmvHe0UZK
2PF5TI7OZhOGig8KLeaLlTbpItglLb6b2jiq0vMaQd4sJhSIuFBqKpHdnp2vj4WuEZEIbaGVpi23
G0aA/BrMNCOOfMTNi3a35w9zEGfk33wqZHwzSeu/0M7SbgX3ABdCPZ4nbTNtQTU/DcGnceyORlQl
tQohOIc8hDHvf7k0y4GHPBC7z5W1zio+CM6EFedmP/JIpwaj5aiJ/A0AMjDOC5nKfKHSuk5X9zIW
+h+H03FL82+0s7iPRYyvhFkJlo1+suXSsrpAHLWqGbGY13wcayVfF3iuPwLYfxcCAH2hc6wdKnl3
QA2lW8BPfcHgQ4LGh4O8twaITK7Ap6zBaYj+NWMzQ9rwDU0U0QgmPVR9rcNZ5qXU/7VGQ/pb5dkJ
ziPdfHldXt/sry8/X63LDibLSnvrEUw6VYh0IGICxN7WnCBRB6t4XtdfuKcdcFBA989y3xBKO1fX
BgPndgc9pZXwPp5DflwgHM6CjnL3vep+XOYNeie6cLHoFh9YW7iEbeNFDCmXoYRsGfEUY3VPuSkB
Ke7n1q+OFdeDWRLz2CCnkRjlezvgw+DxKC5SkMys66QXJI2NENKcf+lSWbJ0lC6Ff0lF+aB9SVWM
G4KXOX/dwJRLk3WP0kNXjgrFww/55uXRhCuJUw8Z9MHhAIcszIbpyzx40SHQ9g1BzbmzhGj78hdT
Bi5vAauTCdQfdq2FvpxP7AxbXXVw1/9B0rPf/PZiGo2Hu23ixkZoAnJW9wFVmSF1AJfJAGcyBAC8
ZcQRw9iPAErIJvwjqLDdN84aEMjGlMxwqbUhP1Oce+Azje2mtd9gKFUAlHuXDOlxoB5FqCZyBV4f
scCoVMCYa8Rz0+Q4e22SthaMHnjSVX6PJtsE/yv/vzdA0YZynUv0XHlMV9y0ZtY0DDvjSpfDMP5r
6MRw8iVJSm7krqno9yWFUzKDg/VJ2XE7gtuSecIgNKQPCa+cB/M0+M9kB9di1mgouF1PLTqrwY7N
6ccwPVX6Gtk2V4TXrbA7QeVcTkVtmaLCKpgh5w5FY5vlEQHQKLXxg2UlToWlumI2fB7bh5QTHDTD
kuUBp6Po4JhmOhBdIm/wES/0JC972gK7e1tO8+VprpiUZdnsDk2nUDi8CURD/opDYalV4TBaiLom
9f84kESLKpw2L0XrVmMulsZmZLAlpbayQJXPaV++5NTyyHZxXRBSMY40TqrCQ/AqFHxFVLlJtwSI
2xkHEW4zjJFYF+4Y0xjWiKCYF1UdMcZeBHaF19YRgOTCtXq6vxmkeq4tlYgIowC5MlCoaeTyewdT
70RVR0XZd39YNU7DI5794VzN5GM477g3JaGiBgCGfuBxCk0MaqYIsRFFrcpAWJyDlq0xAcYnz5Fe
N2YKTYuM7IQzJdNRD/hTu0OAm+QHjaFSu+rGU7+cv7jQf55W9E6MKhAAgQIC2WM9gLpwP8MzTJom
BQnA1RceiY8FBFfpTDmeZF9op8ql/Ko9iDO4BB/e8XB6TzdYtmh77QlV2QGNJOydTbSTxXnzKu/v
auNLEKAozV7DI0LljM5CTY1PaRjvAuDd9GlTBuFq/FS+WFAnAX74PYrTpBwuftmDlN9qhe3rJgda
rc7ieOSXCtvj1psgOizo2DRDwdDSTnufU5yq2Y0EoknSD4c+BHHwiBCbmBwrsE1rILvPIRp0ie+S
ry/mWF70WLGgiwHGOP7zvO58cpj7oSNMa2Px+Esz4iLU2wbYg6qPN3WYX3BBVG2q4njlm/GP5GzB
QTGQcSB83mOngqT8kCmGqT5BHm3INZhe7k1YJzU/wNp4BFYKOOdL5iUpPO6wLBkHPWSOcNNrFm+A
6QPI8GovXr24iYVVodIKc7teKRlJs1Jhx9tt+CVwfJlHTQuSdjqmGabAYsqJh4apnFhrg28GZ+Yt
YDO+GhZX1fj2JpbUjl5xRL1ViuTOzOBqAu8oglSFscUtAOE9rgGwuaRTG6ltYMfH46cqIK+cPj89
PcmoKgK1BcsY8hd4GmUsLEivL9jOjup5izwoKjQ9NUX55GARMAdcsdsa4T/WFbtG+sp653E1MOuG
tfc6pvMYz9C77Zc1xflduX3CUdZFkkdHAbSu8mcY3zKIVdAX1G/aZcnhrOU6q1luR5DezG/7ax6w
cY85JurG2TLZj9PBpASKgf2s/cZMVFupPuXKUudTEMIePncatMBc8G42+SMqHnHqJ/w/ITS7zlqA
/KGkV5gRT6FPNTrWV6NMWqB/xLzTvVlS5bbh/4165oSvVj3TUpYAyQWgidVccvldjhWEnkJljaxe
nK7WzSDA7NZYn5NuoPnkCgVu37kQwdUXumaeNbIwJLo7BnrMEKAMfhQFv9Ce1f5+PadnBtHc2Mhc
jofM92f7B10oPhcELaljgE8mF3YaTJX4DEXqMfEmdeGZd/41TyH3cOw98cmBXAJflHdqdHPTaQi9
uVvf+BNUM5hnCxwJWn4hMW8xltQ3F6fXLjtFHCg6I7y5v0fyF21HE5sHL9VaMTwruvtuuFx9GU7J
vo3zgmf7paHHqxqSolWaxeb8lcd8Ll1aV0aH/sh1WDuqhHgclLMPJ2rezM5JiU1HZgdo5Ke26PwA
2gNIfsGiJf7W9Zbq/JE7ef8VHXrUvh52px+EEfK9XSctxKWWhgdRB+NOq/aQkZyKo/4967oH+FRT
UbmpUnGTKczjWculFDqJ/ghZahljfPzxPlrHV8I0e/gD6imRu/fJIaZs6lxqB/u37LT1ktTcB7Oy
bmZ8SbtADFf/x3zjGQNErj2Ap0dxVTQkEOh1Z8cbCzbiHpMGgOTlPeQR/qyDl8kBQnAfJf/5JYgh
R9N++a29mOSVpUxaXa5M7ED3vinMTrfh2aA9VNbZtc0MH2jleL5jvnJzWEXWSN6d2mkIJ0V0XQ7M
SEE9f1zRcrPDa34nwYMe2D/NNBGdwWT8wc0myqt9f3+WwXyd+y96rCGcB2tOMvyYtL96bHAblcUx
amYZmuVokOHAQ9y/cbALl6Fdd42s8sE/sKUZyHl8t9VIahyqnNzOmzK4AMktIs31HSdb8sL68Aaq
dWzI94kPI3tqMu/nQEil4/2qlDgDeJ66Y53E4IsQVwbH6CJsMMV1Md3WDpy4VdoHh49B4fs9n3Bu
tlkxECwVeHXzIKuWx+rt9u2wXrCLFXaquaMDXXzjXCktRp1EjVxr5XQlrIDfUUGV0fnr3jT3y4IM
wQ2gr6nNT0pRbMLEWmTLlt0hXJnvMYE09Ze6/farkLb5WqwIjy3MrOMBoKwwM5NDqoK2IsFXRKKQ
JA3d3vt2envY7HQ4MZUl+cmucJ0CUDmQHt9MHxiTIjRaY4yTSMHvaXBwwHvV09tpg2frlBxVYjFm
R0B4RieWyqk6RWHvSFIGGhRQJU9e+IMMueYx0/uF6ZI8kBFg84wcJWYq9LU6vPuNAWs1lRVYULTt
lKOFw7Br84dnpZqGwPbqU/T3xhmTPnsPmwdByzy7SHCHukiK1xDWDVX3Lx1Y5DccYpNbzTs88cc/
HNF6Fdy7Z2OMj9Q0xaPbZ7W17fqvPAxYaWB6eI3ukjhwZbAOGixf9ORl+POJifCbT3ZZkwkj4VC2
xZmYeipS/JTclpfuBiVwEPVT1sDNRg+CTXF4VmoB5gqecJS3CiuE0rzrUzMASOlPvG0zt9L4X85Y
bdsCLWoj858Y2JcWCkUcEZWlyhVQqA2f9C/i0Ok3JIpxhSZTXYThBRdYuhNnjaFqTDAq2+cB+Zhl
7DVbia2M1VaXkmf6ZdxXHH6dAX/WMKDqdSKgm4n3dEB5y3Ck0ui4yNrZu2BhjL8GkltNj4nW0/p+
97rD+QQczjJofk03BrDwzxOBVkiSLw5hjVtu5jlrTHn2vrcoORiFuAlAFxqcwI3iqhRg/cQ/bNZN
PchHLKDGKA5KINdOiKCO0mzuURpmxVhEjqi+XBlExPC8QNTQ85p8IdhbUZ2f71ugZRc9VXxsFi1/
lmI/Px9QfYEE3Lh8/FShNI41p0VzMqVVX9Wr9NWE3AFhk7N4RctdbUraMGbKfxlnhmQSbHmCzTP/
fIv6/bHp2Onnhc9WmwUhHWOybFi7wShi0o0V5KHAYdzOCDUXDCwGmCtGOOfv278fqfCbfXgjiT+n
lrgyr4MQDIILyHNbgN5tbVZn/G2vL5Ka8Fk1ext0NL99bzHRd1RHEXr4OTaB/bcQYM2okw1BUbGB
A5ZgEP7qlFOZ2xmmk+jRT+6NaeYCRvwUNVZcOn3InkG9mAngGpfMjGSUSjjkJmOO/ba6olKNsG4z
SAQYF8pxOIVd+gjQXtaZF2Rs2jjE6gTuzus+zSvZkM0uqpF4fNueKxqqZbsYAUky5UDnBorcWOAt
hie120k5y/DgGThnu2HJ9ZJ0AmoTndADJ19aWpDf1Qn4gj8H0cou8j1gnl6qrrsMLSJFw1yZ8Eg7
JcBHtiLHwRJttnMzFE81KpR8YWMjLF98K0YI5k5Pb0wnydWQE4XUDatHtGhx7VBdVfol2kSd3mE9
KZrIld32hmDvJHwWC56bFEP9uzxZ/WFZ15BVSicWxEfdP7J3WzqheabwWT4+qvfQigTSTUnHgKz1
vVSUG1LRgurSH5jh85QcCCgqwlg6xyMTBbeSWJtVxgFFvpYg0aKFloI681tAjm+QKBz1jHvWBjh4
ZJZO2xpcLBRcpQrKsSBTiJiiYUeMlsJQyCeAVLdMBUv6qcQ1XcqMhHQaX+o6m6rCTLYc4+Ad5cqg
JetUWMSFK784gDsOXJMDEGFWOvkOjve8UYzV1V2CcfWXexACV64ULPOvw1OppPMJNy5TKW+VPrBn
vhP3zDsJprWFtIPcte6x9YvlKlJaYMgwQkMtjh9BQPGSx6iw+eiWWE/5Nzhqxom87TEbjmsMpIMP
EujyEn3T9Vo0giFNCa5FlsMJUl16tqgzJ2LgTK/sTnzvr2hnjjMScl8WRWawAdPSWLqQrJ5IqL5A
W1Z/kikX8Y2UkLAf8Hyzu4mGW7e2a0Z1Hfa1Za8KRn1IJXveCCZ6zsO+Cx+bXbHoFJ4BvJZH7+IN
kxWxkL98vDffvZnpSyGnL9gt0GcoBAyrOfgQkan0CDw6RAEnUIIY92E/RLFJvQMXXupyxCAalanq
BkbaTnfHHp4XtGcBlI7glkqHUtrON7dNAT4OrqcOEsyDOcws97kp5TOqGdR1ecWcYI3wPI1d/j3l
um9QyangRMErFUZ+xXIxdAcXOD7JnuCmRAkMRRUIKJE6icann8lK1j55hUDr84FTRvArHLqWPCGH
DSjqTn2ZKOmvaf7kGiP+SuV6cEY93r3DoLEQdew42zJxQeyJ4TFKlF5Xn+pz5rnAfH2b5y6vasKp
Hix2C8bO/ZoCi8IFk8hvnTn8+tEC81kgPiqIO2WPPyYdqAGvU0Yseguz5Od9ShMlMWf1JNspMG2e
r1hUyNapNjf4J+G1044It92Lef02P4VTlaGC5+FPe49ZjNgOrOP9Ilv57JX/lQ95611v0DgMnRcD
hQpdzJnB/gZU4XI4bCMzSCfGq55sPkFM33k5uTqj0cNsPnmguJuta9eEKtmqJAnmo2Lt5xlpk+7Y
VC9qOpRmTPf3LS+RFBpksNQ11GSqzliratnMAX+QVIkdZP62ufCA0fYCAYFeFfkOBSYbXD2c/iNj
JAicolVETKLzcZ1kihbQXLkP/jRaBZ+YCbgEYNOGhA79aJtwQbxMWpJyKZ20C8ImEebpP4rKhYPB
eECX9HmzrfiLFtlmn45t/4MFEr12I+8pnCEG7hYtQ83UnI/IXStGWjCaTtuP355B69H3WTRAU+4T
hwLjOwE35AHcAYZXASfHe2xFrGvgMkRtrpDijXNKEENDUoKiwQmpCVeJSFjZmbef0MkznApwLt/w
CdERMHBL66raD4vR26gvC7uK9a2O4PULLkh6QJrSA9JZ23w+oGZQoB0fWlLu8UfpTf549URDcZLu
OO4SgXuSm+23yaYLD2ehfARygrOJKOVx2hpA3L4D+BjzdsYhwqtXnPy9QhWCFRRt07jSlC33YLXe
9EcvxynvTg+iPYpvT3mgk+rNcQRcffaN0bPhzzbDm9W7gU4HoYz4ObIiwIuzr461kR5hVImMIWIu
zf8Wkhh7MqP0CceOd1G8st3OwcN84uV/Nf7yChkVX//m2UTHYskdFqmLy/3XbUo0lU1RRupPCcCP
IkJ1cpTZUQ8xyKFPrGjsH8Bbytd4VQr7GK8KW0OEO07oAXo32VYidSNg9F3HO6ZqTthRSMRukeZf
+uKmv6VaXrGsNEMTAMLp3sgzGdRf3or7iSDybkZV+r8Qr4fvSc5/5adX/t8iAl973S+sI91JRGjc
oytypeUCHZ0z2fV9vUKptrfYpz7NS78sspxIwN1S+ZUnnLLvNAZ53BAYSCD11ROqWS6WYALu2kE4
d+QSgO4z2HKpzOeM8DjEQVEPoIgTkA9+MuqtfoujHUcjCotmIXFxjp+914j2BtcSTkGubdg4Kva6
ybUeVIfIb96eBOm8PNFG0NLOne2hYiUN1l151vw9bEszXDLak8AEMFuhEURireapIRjQBz/COgMB
14UB5FW9njOeLbrfNtmb6t0O2XgdGZgtg2lAI8sErxprC5deCq2valCITa6uElAeBcoSGtRxYjvI
cRMvUM2duI4YqdxuTqXUgPHXXacVSR6KLr7vxC2+tDNF9ZyqqLCzFmR5T+VDVMZaLwSoCpRHdzVk
AQYftxlOePun41FHzypGkRhHPiBllJdYUdHdQTBkCIMsnX05w+XFM+8V4Lz43IIvnDVbB2fD1Rsf
qL/OyUFJdZoYJvcz2wGqJpmF7YS23g8tn4Vly5HkXhHweUubS7Q0zGBhaF/PFKp/ZBeZSWghW9Ne
5EBOyQnaKUBbQvoEQfAqPteaK2vjvJkJ4njrPFvUkNxCXgF6knzSzz4VzrPbzc7nmtQLH4h4pdyc
7oMX2vXf6z15KxiAQEeRCtLehNTgIQeRaNPDdWDUjlx8RBfl7+gHA+Rvw1LSpaVXjg+ivquM02tV
yKL/XeSq67b1YjPllUw1nhKSAwmxZdW5gFvBIVohNAj9KplRN4ye1SSBbE9TWz/ZA47u8A8O4PSE
xJCQYQlBvpnjixLDVDP19qTtWR1K9MjojCSr4fga9ZTkl8mJ6QkKwb1w8CNraiSNrgQRL6NOuImO
aVbGVkm2mciENEDwKxrG9Az4IxLnWU6KtoxIf91qkCPfyrO/OSl9J9wTru5o0Kl+kBygVEnTSeik
JZ5LiLs2oWYnlBoCpEjiXpVQIVf4n5/Iv0ixB6OuRP4bIdMCqnKjs5DnaUO+MgB7AW6n5mYkdCir
JfkhQSfTbJ+VvL3oDiXkbg0YaCXNzWgjGcvztS7LXMrc2hTXVYEADcq0TIgXvtOHTliCKJhV1zIO
YD23j0EZ6jDhR7hC5jHK+CictY7SErlUx+tYWmZcYCZdTTwqcDxCfBEJUqLPbas3CNKiJs4RJlKy
NvMcZPvVhAMMI+F3H2nN4SMjWExFtGvW1SC1sM6WujZp6QQSieuwo4XNbRJjxb3hw4bymw95Tq0a
sRIACpBuGDoFrP1ztiMDean+7zfKqp/Gr1u8I6ZP20sws5XmkwUCId7X53UAPTdbIw8lxTlz+B6w
ou9ZrNdMd6xesds9er7Xq3iZ2pl5g2reSwh4Nl0BqFlu7JeBIENrYS+443H0aqiZo4JN0N30nLS/
toRLD+jGaMal4DDEdgzz5FqnHxO5pIoAZLuUdwAqbk3cLfaojWn+okSmCy1QxudFfnwCnbSXr289
mYaB8BBJA9iCZjgD/1vgf0E69Emj6AJMW4pBlvW4AUAi3hWcMHmAZojVtgtN820nGDGlsYKvpire
DxDrw++OxgzCM2aZ8yLSO4l26eP7kRS6wEPHj+lzDdZGg2oCIPN6iM1A8BZTHltT/dZPlFTIQvCq
bSHlk8WaiGg58Eiux0PdsSLoFzbomlRNUlKyMslqzCyqv4Ks3R9RWZwa25yKS59Rdg43vghhBCRI
mzb3Is+aM7MVPiznLz5lHF6ApnIDqPrzjLuNyCbtrJkYAN8GEjQ4vF3pXK0DmMk9qohYYmdyeRfo
ZnEvK8SxnYgf6KIqzhiOmPoVm4pU3XBEZhNEsfkDFO9UAzmqbzluF04VYEhjc8fWJNH5/xnQqY+v
NgNLIQEHSvZfwDQTj+xuhkasxU1RcsgFUPDP3SSozSLTukC4jYqwE1DTtvveJK5x929p2kESbIUA
I0HXp+yrWHIyx7tCdaqnuAm+pjJrEazJE0RUfiKmzXjsTlYNIZMco582SiTqTa/4i8EFrkYK/cEL
6mQJX/DFsxYp1a5xsMlSq1NqYPKixLITEZAvBxh8NDoEFgMZJs+IZj9JyAyF1vAWh4rt0rx0UlpM
Zs7MLWTWS2eDzuuraNOlqVH9ADq8VZxUVvOx34QqB0pDPOj1yp2e/THqJ+nTk1G5Bf63/pv0G6bs
N0GlRa4ML1+BYMn4xevWZ45uQJT7OslsfrbcqopNHFD2FUgXJSoyQWQjFM3FzjSiirgQfojr+atT
PSYzPUfTaIiWv+kK09scxjwN+9KudP2lvgVkQopcxhlUAYo5T/jmDsGekbZ7qeDtj4GipZ5pZ7oy
7qAJj7d6CsVBimzgZI96IkP7xnJ7+LbPswIoyYE0kpbc/XwvkiA+fdOmFv5xy0aNb2rR2BK3pqXI
ppVHiZUJXYc9vS1h143XSm1l6MgkKco9F7FZaSaN9Zo/3Wf7OxbSwQlX/O24Mhw3Jrt3r69Zos9x
2gJRxnM3Gigw+Cggrf2NN87pwgB96JWkdHHR15EdhexUblsMJuyvOO1aHl+ikG8V9oo3rjPOJRih
tx4fGgZ25QTm3bYAEGHoZ9cQ7ouhH9pGsFPdgDu5x9PCq29sgIxCCeD15BaQjtik6Mdk0Ydlul4D
x4F6U24PAIpCLgVHgX6/IncrCmVSzkJf/crOP/qRmJ18Oa/mDHN2Ze6gxMfG34JtSpTRzbHL7q2P
zj8HfRJMdCNo7rzmIJ8DHtBpklZ3CSEToqv/CB6RnMEqBW/4Z0MltHNQ6E2+XK+2PJZCek1HRjY9
LtbqmmvAo9Qld5gKIHDrDIqDzCqG0XXaLx9Ok/UnjB7IALAoDB5PrL3nT3rv1pmSSMAZ5GDgQP0W
d4yVI6MRbJYCF0JeOJxi/94rg3ic3IapWXh4L/Kp0pTNKwuQI0Kfm9rDmutzLGP36zUesRvlXCOu
BWlZEXKKbBJY0/Ts6DVWXQeMZGS2aCuxOS533ooLvAztLtGN8b3IX1/y+sghL6osjpNFppWWo/i5
hZyHMHT9r5JXmbThO05QR028DFhUSiahXAWAKBs+CMFPqZN5A8I6BZnN4k9Bpaiy17TR3FVVuMBC
XisSw2xV2CWr61zjUHu02tbjoBb/A/EmpQiyDAwhU9U36tYoOcEfuqQTUr8IMNJ1f9DZI4+C9wiU
Noltd0OUfUaM8ZzKOmWbte6Wk/X6011uGfVCQDRPBs9JQvEvaHbvU5BpjxQ36WatIWDen5rT5heG
I+IxutCsk2Q2lMtejr0f7R2pTf6l7Tn3h9N0jkPRQy/bE1aVF4W4xx6Iy4VEV3vNsGVa5Wa6o4uK
Pv5cp//hPnDkh/oIpzL7hdtblAbSNEAtiG/y7/iAdSf1Ycw1shisO403qbJnKQ/JNQjbg655anlb
eLId9j0ZaQvc+OFgeza1IPmYBrF0/qlKk/5HUcY4fh1o1ldTHImvKkJCf1hXoGJXfHMoFOyNOhhO
WaZPSXuhEAHMupsBYAuUCluPegw75h+D/NXUYjfr041LzAPEizuis5jLOurLAohku27z5gjA6zqs
Rrf48xQqtsnMAlwCjxndwI8G0sbYvFy3Rj6FmaZuX6s+ySGD1S/XSISUN8NIO2T4dn1DJ3dbxCgX
Z5lCgh/J2mj3+3ze0ADmsuCcDt8JwJBZwgl9xCttduwUvkKJmWgxwVFTxHHFpruc/9QIoGma4Upz
bz1hr1L/sH6u68gxJ3QmG+FnqJEBPs0c9fnZX7eedoqbF5OO0zd4drCy8xPjaDIpptYE2tpo1dbe
AmEpcKQZKS4wnnwrCu0x8wIIOrt8L6TK9iSd8QnPt3elIECfPGC6Cnb5OHxB21bwp7+1WNLDsqfk
6t3YO3TWYeqnhluFE+N8c3f3ORf4ib3HQ6MgwIKO3mo/RzslnKvLFbMTV6boFWzJkc3xAUO+I7v3
hAExMDLmZUNgFpKrY0T5KBhtTJYzufYL7suONICnjovul8jqAuUscuEPaYbbeKipm4C+y/Owm+sz
Z1qU3gAKSx+pT93dQ4v4Rd2h4jq+GEb2vKOurrPlvJHAa/HUQQnryYUFsoWceDhWQIkrFhdVnVqa
8/Nv0RrgTN9VzlA1cUc/nSkxCpx1nEpXpf1Z7cB6Iaho0hKsjdjrCCAvA2naPlTwlorHroY8hzkA
y2D3BhtA/qvHsfiMHUf1m+j2PIGhbBQt+q3/5FJ/5wL3RlIW0Y95PaaT9fwab4Qk4PDhuyLu/W+A
72WuY3arijhSFx/CAF2HNSVcC4rrKsaSU0ky+Hhb8Gy7QRy/BF5zIpD8RrAoSkhIdKCEIp+mDcwT
q21XvbaDJR133DEN0U1wd414FvY5835CJ7Aoni4IQ3mGe+yBQoBnAO+pn0MYkyNFkSWwTG7rZLC+
jC1YFSYag3lQn6ZEQN5ruKUeH/kMBIYKj1gzR2LMNf2Kbc4mNWcFhGCzr41RXKUWYr0wsLqr6f2U
KhS6Wg63nQFOTP3V7r4N+5EbNgMHBGxMXZXjE+XcAmuBw+IOyHNNOIRPRasXviCOc8PysMM1uf7m
G0661dyuf/VSqTIAlV7a+HxMU6q9JOWYurP2X7BOYK1bmolVqvA5yTTfeF8iNxZlsvpgquV4MN+i
Zl2kvagXRcloCYb5si+2nOpO5VyK6PKS2QMyLG3t3O6KInei6Ll++WwNPhwO/Z4bgUo9lqRyMPTf
EpO8WDloROixUP5HGibDyH1tJ6IZIkk6xE/qJtdmXPmzXZ904IYbpXHa7KC5CcSGCuySYukeY+C+
DBIetztnYC4Y6HlcqaBwN5S/O0fwpYpyfic1H/+TMB17aUaMXa/cIbE9kSBkgY0jXdvQeXFNATKM
55ASEUY/Zargmtf/lqiFPrbN+LK4LitSUp2PFVlVZZt3yMwslQnp7F5+001567yad9FUJ3faQabe
FCd03n+5F9bg0o65upI1bnEZ7N3SVl7Uu5pohCFWSdc0xBPftwuoOjWL/YzIfigWUBQkwAp8A51Q
A8pKe5FngLufGJmoh/V3hTvePWGxllrucEn3gjUIllDXd/a/fSPbNcjVYxD2Amhx7z/O83phOPTs
8KkL5HQp1XPx5Wn+1o56aOF+Vkq0z2F7Su79aTsljYNYgMn2T5XxtF8TjSa/2PHRadD9t0egD+dJ
Zh8sJ/WJScmSA4OAAMd0GASUcaKqhbL92qAck3/SLjnfuBfd4ylPKQb96Al483uyPV6bYn+shTTm
aNdjtOhGn5oY8PO0DNMYFnub1SXI1Cl7cKGIoURfVwge2FnrBdU4xKqkg4P9K/1u/h3oQlWeYZ/z
SWS+yRFgSlUALoZUg4Tmf+ramCCFGqHiw0yAt9cohCLKLv28rY03EDvQsSrHDZTwsx4O+cb5JHkz
UrQ+jE6WgMeZmO3SDP3IAIxiqsxTHYWuqZPuOTvpHfYVPj+hAcE97u843qUjhjn/kvbzeIdm8iwo
AMk92J8rn2FgnSTwQORlc1pGSHTbqVR8eT+YJagVx03U+j6fk2LGlYowTPPamjCXGIZNcRinBji6
QEO3SJqJiwa5Ap9frXJWHwJjr1eOhznULXjI4CVj+Nb+VyoCVguIAWMuHIQ5Fta4i+A8EXwsPHUZ
VzdCCyHKCDY3QDxhrsOUaKfTvMAx2nUbr26StiEw+z2IN62OKaCcamkuUbgdsxK6iUDWH6fWUOUL
3/RDo/8le790DVtL15Uu/UC+bIzOT4swI7YWlZLOSEGmQT7TUwLGRr5xTH95lTzjWMRuTevacRbD
qg3BgGg38sO3+eIFFODrG59YRjnzN4Tss807eRndiB/902hxinRgP/fmFU7FpVvMa7j7/XsDBKN1
P5ao4wjxpUkL1KllURdIU2Cug4p7wSoMEjY9Sc1uj7NNyqgRO34Zmo3/VBPU39ADCz64MevAS8g/
dse7FMbhYBKqYkXBsyE+GCkJyl39nrLGlfgjqIktpZTqxFpIzoRXbY8D97KEtnwdPzBhJG4nGA1z
SSoV6DhtkCXumQTOXqCev/qRRY5ixlqJ6ymC73xEyxeU9iRf+PsOIkBsQROdzG9ILExqBO/GkV6q
IRLpFyGFvNeV9oj5b6fXsK5lvS2d59A5IhGEnrHzpO8usvy8VcWRujZNQAMtazcB70jSAv22pnBR
iTwykYGyzxRY2FQ0OqRD2EzAt5+AefBAi4DpctFOVhH4CCjLSMmJ22uiucK5nW19INdzfb8ieWys
5/7K4C9ivTNLY32Tar9y3491gpS0ar3V70iwR/+Tn8cfPSllsRr1BvbxeG2T693eT2SokL7tV1jO
nSO7AtytMk0Rl7xhbp7Fc/cXiOxnT1lCsrfCqb+xPFoYq+VQ4zRztZISiF0nN69UpOV/yylJyRAg
PONmPeAFJhuqALLwVzyxu6YvgGM7psud5vuVS6M5s1t2rVCrIwTe4G9YVFuL4XeIx8mzP4unMRYo
Vr80Tt1b8e8spVSX0YXQe4AbMQxXh3AbxXUvz2+LvpYWJRAiK4qbAijtTRwHmwtYjiMyrAYvyp+h
sj3WHfPHJfe8rvsGy1Azr5FdFXa3KyK5sr49Y6AHF1YZzBwUZ6RcTC30guz1G1fN0T3ZJSbnKC/K
0iPuOnfhzNUrKxJXsJQJjA+T/tsJY1CBspWkc21Kp/REI/NL/GnLdfbc6K47uC1MCbbTf0MJybT6
GXyxTV6MXQCTeW3YjdjGKWArY3CiIWaiRFg8bOwj3rSrFIH/G8t12Q6iHkuXBO5MIv7rgoyj10Nl
awyBikPYhf0O/qXNhMAntM9nv62snXpD7v1KOlulghZGsYDBNJqGlJTY2zntalXIwhfnMA1ZTxlm
tfoBTuJKuQFdAiY4clLcA8ESPT17u+ysPPw8tEmWLkNMNWA/VxK66H4gzkojGggpJTS7oKwr4Q3p
8YuZaaMYYWkIVJ//QBI5iW7+axRuVresIyAORlvSWThNsFDIFwuKP7IWAzWiOl0nuh286OXnXrZH
nDzy220bmZ5jjdHn02xqxgCt9L5iZKGTmFrvQe3NTWhMhGTShiAZ0v6k10Qe5gj0AvQ5u1a6Gio/
/IuNfGEfMmEWvkj0bztSsL6vphPJF6lVfunV0cB4MiXPF6EdO5eh4VNt68GzNeLaLEMlF0g/K8e9
30jWPG71X9rno09wcODQK04LaqV2HgTmRafR4h2QU/eAP0xd9glm88wyv315bGJdZdba7H1X1vAJ
PpSrckPItDFPo0gAVVTH2C9Q8LLe4SmDtCELzDv46vEVP1nbgykTRacC9qgSnMH9Ux7/JsO/8YAl
SrhWUlDJHuyrjc78WOpqkvdZDNkAsBAlQ4GcLbfIXnVWJMW0VqF5ihW55A0VOb8geY1ADf/xMhGL
V4dhSPJXNoLeDEM9zPhCsBOVpLyD3bdAN/qmthOye56O9/cHb3FTOIk1rF8B4LqQCjQD5D6sjHMJ
DteJOq9Tt8iiWgoiwVwmB3sQ1BLSSzP4uprL/9iK2WWfwuB7RpdeU46j5MVTZ+Bx/TZ4Kddkz91L
1xl75KJKJkP0lLhhCuo1ElgA7NDwhUIGoanIKFkH0d2/6F8FS+Wptj0obOgUg44IyaFbpd0+AnnM
AabaGGRwHBunIShmzfhc8xQ6Bw0s5xbtXVG6a5Uai2+VdXuhC+wAJ11aw7vyaGKlEVNLCuojKtB0
tQWD4tg8gIATrxXMT19Rr9JeY+HmS87Rd/BUXt2EMk1zG0bEiaJ5akrNsmjx3NnwYmO5l8s9PXed
MIgQM5jipimwMkGBQklXFWN6VLtznBfWLt6F8cdkm9V7dA8efIjQOOG93aSyQ6MUl1aQDocWIgRy
2gG0Ck6Nv+foRo9tAiLOMDS0kvnw1z3YOn65eW6T/qVOl1N982+c20LoSnryD5zkVHJpZKrj9HIC
GPWp7IZQ30ZDwMQcUZr9gKvMLwC2HnpWToYTdIwLqdMV4TZ1BdYcxCt83emvMdb4yfNew3Srzilb
VNOYhu1K89bK7WFEYJwzTaY0Ywf+OjQ5Dpq7gX40b2XxeAzpY8jGnT4cFDA/T6h8UURsCOTU9kNI
rLfqqugkYBy7P2IffIBZx92HEYobqAArvZQmE9FPoZx0GokCTU7HockQXJJDCgAlv7G7d7Ln1bk3
NH23XnGQVzjbmcX7SZOZIh0tzP6vSRQx1izazJetSE5XwONxGnF+9Wfl1Yr0GKRQi+8IN/xBoDCb
gCF2jzrudsVjC44macqvV1qvk5q9uDF3Xj++BRVAoOSxdfmn+Dhl0QpXcT3qMy597KV8iRyReJjg
5e16eb8zS/MQvJdhmvShvEBEHQ0TEEruWF7ZHcwPC3v7TWsEmBNyyM8WnJ7RkXg5liJUwTZtKLv0
R3zEePbnyxJq0lPTE5VbcWbY8mQgTOdTd0wWN1pvxNUTAU/DK8kJqM2eGuXs2N94M8/NAnLSHBrL
d0l2DRP0/awpzIe5z53C2CWEXrXKXqZ8LOQzf1dPpyVDndUNa7jDiIJnnR56qESZjOlCB0Vnpdm6
YLDZ7NsJx1meiQXY2wLnI8ms2CaHTxjayzLTFoDIajXgenA7oKZMSPzS+3Bc+drThmqr2+Oonohu
2fh/vigbyONkix4jehANbGjVB2tKE1JuSPApfjciSWUMUcYd4sEiCVRaVcFfTvRQfIPOPqyTnCi+
ekO88aWvr6JuZ4thumjpThuQjtZrsrLiG3yMh8zqIIlGOJ8dYJT+xYSsG8FW2QOwhM12R86bz+dQ
cfhpXKrV5JmiggBGkr1r55lXiVFKd5tHHm7vmbxeylToJsuTAIud04idsV7G9QqsVQBafkqckMmO
HHLV16e+jTAXfXb6gwTfI4xUoY5oV6O/3LWVnT33CJYchAYYMYFLZvTzqQzXXAKJ4T221cYjcXPh
NxrT6PzPEbiTG6zkFvuXziE/OL0990KRCbMIDZQ/31FbkF0o+LdQbz/Sc1rxZPPzTcP+3d28zW3E
rw33/+qzsKfnFFtu+hN/+HtB8V+LfSRgMM/N0KjA8MLsFfx+752rtbewWjtz670yMYbr8wxPb5+v
u5PQz915MBezetjvWnk7R/mn+q4FpZgZXFHNvvGt5Uq4yrE6Sv+xscTDK3z+zNVjN3Uv85E74pWy
0xJrKSoyyhGx0TU7GMLU/lvKPb/Ss68oxFBxRFJTCBNF2ozHci23Dg2g+uZHSHXlEgEAmV0Vt+ca
XC4mS+bKC1QYmmaaoaP/kv3DvS4a3PyTuQGJll933pztt1apQIYCZD4bbD6A/r/ZQ6y5LIUWKD6U
uGMBN4HbsO+x0BW9tbXvsBCDV/ljV+qUf0uUt4QC3KUDGkmw/Og+H6bHii5XqzRSCDBNmdpmyenx
mKPjCBgknxymhGIltX+w+dWImbP7pGKY5ho2r5u1oEIyHg+RVJAmKnnWJ+gMQmJ4oTQhi787H4cf
ROejY8VBYG3cMnPYQU9vdq+BmYLdyMhZitBmXS1bR8ufzCbWQY3Fn/gOTIm8hTJN1+xPJd+ERGHw
kSab2ILGWA47sS/ip1qiBT62GTgCpgNDZI6MbynU+KY6ED4e168g+gLolTShvW39hr0Txm3AbDYL
zwAryatcRklSB+6hyxTmcfrnH1i6cVoKFpIZk3StoTvtGqwr1NFio1DfhFkMvl04QEzA6jiOTAI5
GL2VVldB6TG9B+BUJHsBo1L0o6ATuSpto19XBq63nbWg3JUyNRC9p65aUUgd+Ym+mv42TLTajqqc
XOouQOGqtaHNgOC12UIjzXsQUCGV7OAE5P2MXAYE3VHsS75+JGmwc9+aaA7WmkKLSdDJR71kng4b
PpVLyMK8/mG/xDpnN3TwwWMjnVYsGnc6jCh3liWSd7xk/vGCeNMvk92fOBOL5BJV2uvndnM7G8dL
hbDayWLWNmtyWa+wqbNkuHk86lNmZKPzR4K7Ks/EdAluIJ6TNtCP9YBRrjZH7nO5UbeXCdU8bCxU
L6YYFqZ0q9mNMC/qGWZEli0jOFLDNuAIip+y2SRUWe8TClo8Oz8r5dv5oZ40NVVxNHB+qQ0WrMTD
YX72tDpixZLR039CXgtUFk3Pt1uQYlwQyDdaDQM2PdDO0AlLpXzRF3DXLvdvso8/2gMbSnjcCd32
5FICv3Ojg0Vi1y0aAUmwZvuJntHM1WdFPdcCLYTZ8GEFDtC8NXPSNt5/naqLCudCq5fvcVnd3NSE
Xc/CUuq3eCa8ZopfhN8xU9lXkSGWyHtCk18WynRwRdZHYd8ymhBrYlObWm4nFHlNpWCkOdNkQx8H
lJIuvOjgH3vCFBCfvD/FyPbkJWn3WjSaYMfP1tWhcIh8FinHKZ95szS9FJkoDX8YBk5x66Dkx6Mz
5QPtC5d8fcM8ggJ+ROU/C03CF0QWmx1T4EO0G1wlq9UFVSWoSn+D3uAAfRSfAN/NsDKUaLYjQviH
lgro+U9Oj1pGqX4/0KlJmec5ZXuMoa1I8ygdmi3lEAwftbYt4QOfssHhTcZsYm6xqnSF+23yZJv+
XSA9yjDQW3ZhJCgB+mQk5o1Z2l4u5E7JPA4jwagWqEUWdVVqaeMt+taB6Ivg5NMpf+Tn7Quazc2n
IIms2+DVxGT4xfqjKFtfEN5zDzDWn1JYnb1S1TUhVyE2Bh71ba3YzYUUA9yIr+pXkE3nJq9KkKnh
3oka2/SaQHu9HEmN76KkvH4t6XqSTMrKAXW7V725rWdVeF1dS9Yo1UNAmE5P7n9j8a92cq9ErVab
tg0852ALT+OFJKrt/G57MxGWdUVgkr1z+hdsEEcDA7xyu4wBP4xAFtx3vi3OATTue5y3p/JIgT1O
WhaGFAnjBs9iSiB/s0eJT/BmMzxqOXE4M0qwu9dlhXW38/ANgLmVftXJO/btXhX8zkGwRaunJQXy
Os8iicyegk+TEMz/Oyi2rMEMMiVmh26USrrZ2CYbeUXlTLa3FeCIuyr6ikJwDufYWfsmw0PyfsCp
nC2BeOk4JYEAbt1q8mf0O0XgpOhpBBP/Yh725TLCRbqUUUyflAZ2UfJY8SI1sgWFH+SfI4jUY/BY
Dz5R6SgkXf7lDQ1vSpZBt69tI8k0/b5U1GtMVlmKqxqSgt4Bu66myWfvbEzQXNYE4MkNwaE1ovEg
0DcUIB82LQSCieo6r30yn7gZnaNnSCcxTucBYwwIWyyuSiTrYjJ7dvXzR2RQjP98Me4iMeLENH1v
R/C2RTMuB5hjG7gJY4zw//mYA5ZwU0k+BgFGjrKs4Oxot9ybi92PPF8VF5BkQ+K8gwrdpJPR3O58
Z2fQ+ROtDhV6Xg8FSE19NEdvtKa/zGwWq8YSIilfaCcxS5x1mQMJqnEHcyo9KvI2wrXtow3GaddY
Jfuqqwri2bgWmvxI7fxY3X7VCM9kf7Gppzz3e8x19eFkh3bb63vhf/CMeWjuWkCEEnL87u9Taxpr
bFehE2ThF0h7Zpz+x4jmGJ5dcyiuoeIUTwvKiwdm/3HyCAhYkxlRSf71jo0xr+ak8NnhMTnktf6x
IEzZKw3WAIH1Ww4g77qyOi+IO4QkFF7bOyo+VCuuHcNyohNbtUmHe9Lf1D4sAEeiZwPtT/XofXfM
2CPx9EtnjspkkfbyADhbLe9yln2QJoXbYwginoq7AMWNMRmGmoSECxmF1kV8BfOPyIcURq5CVh0k
FvAu49B1JilAwUTphwfjAH79uUsNw9t9/foME98hQj8L3dPov/T2YEn7re9KZWakqdsT6g6Y14je
JiLKlvRSYjvfZcOqNp+77ZuiLN6/pk040LD3bYBa8YYdN2iy9JzQgT0ZeAtfFOLNH5t7krKFq3WP
JVPAJo+U8E+htdbXvmjPZ8Nt6bPd2ZMSSXgyPNBs+1X651ORGw/UnIPhigRmtvWTyCq2cJFHkuC1
V11kgPBrU4+bylDshmRnpkwhS168cF8jYXgzeQ2idkXUDs/R1afTy4tl2JfDmkJ5w88tt/tJDz5Q
xW2JeujqO1LKdC3+Y+NMXhZF4MrfTJYba+SKlQSlj/mvELJkH5H6Fo/+OGeVzTYJfU5Z4nfoJq3P
fz+rFxT+ZPQ8o4w7LwVNq2pf53Z2KaDMzkl6esVml8v4SNh9IoqO7/4IrN099K+pn3Jt/iFn3gtT
GLMeiYFecWlPGW7J0BUf7qZpcKnlBhtYU1YvUSTs44JYN9eWyeEqxEa3Rs5/UOjjXsGkP99GTdxh
avPhh0mPl0pY19zbfiwo7frc1JUTUhHc8HZYYQvKYnG6Uh13TBsp+NW/zCFwBp2gQfRiIuEvUoWO
EXgvPKDsI4JdV6GLxNipW7wwAJyzDKBG54oZ1yytAn4o9tUi0pKvfYtMYexWxiaavk5CWAoHEvsX
VHLqXX/85ccdxGqDKrGHdOmEp5sIWO2Xj0raPWRdtkPdK4yc+edhHT9BDw/DCVwZWQntKLabXNG5
rIXYA1T8WqFYseZA1FUBIDseG50BvwRzR+CdXM7AD7h1linbY1ksUkfHIZZTVukj7kLe3udXbTDp
kr7NqLOrTMlk2R/K0oPBGhlXOTQjBmD/CWARI5aAmRdOU6Cyog6UIs1RryS13A+lCCxaqHl+HQBC
gbYQBpO89YsHSL8q9X9zDrnFNC/9gDCvBVWiMDLhOjjH1BFKjr2Wza3t9rojqQBm0kDoBe60CZPb
buKtMzOSbqws1nOQi4+Rb9hRm7rSVO8BOqzSRIuHJ29mUsLCDntyTdswRzrOivySiC84KIic9zGl
fQGAi58XIs7ymiQXU9i1mPp5xDa31YkE9+SuDaAjIkXrmSzC1Y6+MKFVQFGa4BG5WmHNt6kWbuIk
Jdpi+LL1p5r0fW8x2gyUxDwfLLBxc566rM5Ld76YHXuLrWTE/cK/QKsseWAqxOFFdIPhu1RG1/nX
RfLJhkUJV2WHi/+iVBSNHAwND3KGTyPOgzSyjKXqZsaDQjqr5uFHfot5jUTeI8y1whskt0Q7P2QB
zxYVBOQGVDO4VT2dDO6Cyijsqy8wzpmJ3Rla8qXTj3ZchYU/jHRzCwmPeCK9RfGJbb+VBck5WPtv
cTSI7ceVCLMIOYw8hj0IF7W9mYX3QQg5Tm6VM3rq9a78G4yC5Rijl65/yPLE3REmEVt9bb4+Ndoc
7zp3fx91OHoS3kR4Kv2b6zXxTjjoM4ali59OqC5S/zM+CVuhmou7q8YsTgYxjYRJdKl1fZBOXIk/
WYSZGxee16Te7pCwBtNcuzL5RjiNdPmLnU7DeVW2YpH8rtEAO3nMPaJHW5PKRFneFRWWOcRsOh9G
6eubnksCW6uGAmPY8rj3Yt2CwqoSAcQy2pDGdSZ6s/83lBd5pAu0kuyC+3Qp8XjLGkflQOWG3Odp
g2Ismcf9xOpH4gsmxdspwFK0RXq0GoMDg+zNevg7xTLmENd07C1yyQBf8orKWC+gc7tdBndbVj0c
NclJfIpYWY6n0mOm7fhZvtiZnFwsPEAyfNH7r2GxgGA3fy2OeZzS1qMpcVdohOybiQonGJDexip1
strzAl/Wo8uxwv7wiqyZS9seDqOzMMhkAmjGmAnxc+Zc9boaqizhGLdW6p40TaYlYcxZwrOPuqlK
f7pixMH9QnpNoTzmgGlhucwtVyK4p+WIaKLNhMYRwi31c3ofs/JhphnBNsmq8jypqctPiEQYodgJ
2RJ05HX+ehUjM+RuTo9Q+gkNURoFaN3yXJMSDvDBRvDmM8QcNM5The4lPWgTBORQGInldaHofCMn
xJV0rxfmkSh6XOHQt0Ll/w5Q+P9aCdJXiOKEEm16jOGCKQ9l2tt+BLyKWJ+YXFYoZVGlBpaicBTN
r5xpdSfDyRl+79S+Ayy0izs/jdZULVX7rMJN0rSjcOb/T2B5WY1SxPrApvk+IZlAbnB5BjQppd4+
7/o9RVGVVdlYxuxX72M7Yu7DoVI8JmnKghQvs9BmT261cOpMD+dK/1G+IFHz/tSBSyIPrA9OePkQ
ZV7MDSeKgquVp3prABeGrcXHp0BtuLWyFxKNbvBagG+5urK1S2aLwbxcHsIu91ZCCYKmcahJcR2h
uUj2rvIxcM60a4dhOxSIU+6gEbzYjosvUtpqkOE3VADEH42uxlz0zTyvipdGOt4B57MwkTTvh12U
bp0/HLfXGLrfqnq2MIkH9Akw7vsvaFKeQSLH1Zkj/uqo/60vduZh9va8RUYW2FRXD3EWpY6z7gSf
8S4R40T1jdP3d2b50i3k1prPQsOY0ATYkltWj/Hg3ZzRqCl9LsYFsaWzIYn/9ieHn7azGXtv999R
uMWiesTiYN0jAQkyaUcHuDm74+0mW3tCsnwDUewQ6PGFpk3m6UwQjES68uECHzJGr9M9CvIv+J9i
oHNMFmJl72xtMS/ac48SLEpmYt4VzkKf6u5UWlPwPVXqTkh91wJTaub9WhHSw1/qjsm7DerpyV1l
OEsns5lM06y84Datkao1F0x5RffV67NW4RwioM6PAkcRAPkB15Bg8bZQZHdF6YJ5YwuKhMaPO0WB
MqTQVOUISRRT9TGXuMWejJHK+kSMuGHLRIy/DLahnFq02Gi1gLVicEqXgMAn49A1xIBmjW69WHVx
cIKuvE7HfrSwRv/1xdZH6Q6+TpxvYpvBAbvBlABLkORekVR43IJCbrmGWLXlpSmdSZ43w/e2g/R6
kd91NJUM5NpcINFdWeZdi8LtLQp3p34CBOB0fL7u1OdWnwoEXlyu/uckL/rmf70cKDYRcsH7urBN
4jnpskRP1myCX6kQN0dNNGPihgzAbX+Do4p7XucSc6Ss+ZA+AeQF7xQfEu/tku+tK4TOizbGQAtI
muo1MmxxTdtR8MRsqFq7zOWCQyBa6dAEnR+oTo0tir4MDXOB72Eeykv8la42cUHrCKgsab7le4MM
6Ypeqsy4iBmkSi8YnNx+n7TUWUdD+BEBDINY8S0yhjN8oZxWSv8752Sx0TgqKA2e2kntj2LkftTg
pR11vtg0d+DcntCkWuTb3Q+5nJt0KHpiBmD1ZHBXvZ8MMwKqOR1BNJZPc9/mcv6gPwSaAh//QjBX
VvESWZUm77pRj2MwS/Cza8j5VPnlP3/WF5tP3rdFuAABkYrFd6oOb7N27fuuTDb8CYRbiVbEIsS1
qjZJd0h1EKoZWjUez1bDwU0q0DxVnchT4aMuEd5BlHDy2ChVqnZwzayroekbQ8bUsUavK92oXYDY
LWkYL1u4jRNcsVGbmvEswXc/9ScM83XLhljeclhOnDdzBVj8pYzLEnIFtBIByuM0Y5+tr4mDWain
aWuK5OGz9kYWZNBrSZrCmw4RNZqCvchp839NmVwFpBxFiH2OMFXKuuYwDhZSloQ/tVQGoZy8h2Ce
YZx3ku1VP3bOM9gHax+AvtnFneHcrcNx0lSY/SeIESa12ziv9EiIXiHFolDO2SsH7/OBuqL/dbq1
hQB6uPlTD8uxE9AYMqeG0c1yCPdlQcw1tQVruTpd8mzJwSOQSTN1DzUIMmcENQUNdc1+y7HrMe/7
G5Th3SuF3WQJzstTO+JnW43W2twfSOim9R4C+i786opUPc/niNuzifH8WLRH3N+Ql2HncBB64C1d
zsVrT9r94UyN/+BbsE3FvtDoNNaCMyGL5BpZWIescBOGcVBiqJdNNmsiZYXTeAgUcjZ3ZQ4EOHUv
iTYFlBZX2a5C1rV4AlizX2bpGzWrxPAxm/LNqDqF1ZWA0czHhO/jMAaab+CajufQ2DCD35a5bmLx
yngvl6nVSQ5UT8VNT8x2Erj/j3iYN8UbqF28jBezwy9ZUClEL0aMjmfsUi7wwD55NbbMCGxRIZqr
x3HikThxiJOCPdjQdrVCgSIwAzJZpONZ093SUIq2dfh6ZUgL5cKclyrz2srcr1Af9oRiMNHudgIN
KNT0Ir3DUuoIfDgcQyXa7OZ4h1MX7f5kQ2dbtShvIQofVkW23hZe/tIqVJXZ8gg8TgOQCPY5dVz5
hXb5Unyp+6PKlzO1lJGRroVoCP8q0HAPWnGTWOKCzi68NxbLJTlepRiOsj+Kj7wdWdrzmbuP5f/Z
mBhzH10kjoHpMjJUXy0c3H1U9aR/lS1rI7osj3AzPPlpNDl2YzQaFHu2ab6ceh8qUiWKCl8w8J7M
9jYObG4e+oxGnR16oXTRKKze2C7yAZ2yyTx9rsPa0gNuZt4zNHBdHQIR/uIguF0fMNn6dU82bW7h
3vOayqbjHCpKrQg5RHudCIjP1x4OmhcX43GRlodj6zHb24zEdnDblJHqRdLwgUMKhpdqriGXYVH8
yelMw5yfZEymwDaS2hcI2XbA7oPIx7dtlLKtO9oIMjFMACUMBM4iyCuCmpGyKKIEAlg8UgcheShv
NXGhYbe2uART+VW8C4JPDKhRTtWYnpNgnkIxd4gz8989KmVCU4v3gOIhyIsjXmVX9AdI8+0mzbFY
+i91ZIwQhWxYBZsQvBqRuHpgyaflzieyZ5pJzMEySuE78v61nc5M8FNrseNYwIgNTw2bsN6GIOJr
istivoQUf6yq/46rqkOOIlZgv9/Ob2W+/lc04y6C2+uUvFNuyw8PfZ+xYzK/mg5Ip6mJ1L1mqPCq
fWrqn8wzIc832my6ekNi1FTYQPABYfFBOnCsdkQ5M3sgTpTUrOB2vg2LcmRI6qN+gBPXKaLLlHHG
Z/+Xf7HqRiga4Q7mPxf+RNY123wq5PuUqL3rYgrgeHY5ZHU+nx3P7Boq5qUq/UYzgRR10KoqF7WU
QJbzbzWJZtKm3QNX4mps5skpG03hIFjWZaLPoGwyR2EjN3rIVmmjlr15la9N0+HZ19+bE/sqXaqY
Wswukwe/N2sQG599H5DArzyy+b0uz2b/mcWnLSB2Apd+1XN+GKoNY7Qdeae1AXQAOtUx5Ux6Zi6w
xkbtNQ0Eka2bvS5w7BgL7D0PGZNdIfd1XzSXmwYR2kXsZ4nIpPVZ36aFR1i10DOnJM7xSVihTkr2
RnTnGNihXyMtzG0j5r84rsxmbh77JIJ9PeWoGcoBgGsRBesTswjOVuFXxkpOnkalZU5HfIaU0No7
RrQCl0mbY+UND5+t1ZoAS5D6VSupiebp4sPF/NfnD6vqjeRivA/7VHTvakPMbRI2cmwQ3gezVeWX
OwUNEKcP0UXt1+ZYLIbY82yrC7fQfrdlQEoIgTG5Wt/le62XWUL8H6brgB09lclOGVW+DM5kTv2P
433JjPuIHz98hyyVEPIyfVI4oldR+1Ic1esjpk6awz6Q56lxQ2x0k4kA7V9C9C+AxXRSI7SffdY3
O/BZBr4Q+cLvbjkQFsI7ZokwwwT9DOuL8Hkl477HOGY7QacYC0tvbwduJP9YG0xpyH3Q4fKYV8LM
szatrULf5sfzOk9FpfVxb0qeqcxtmPiB477PVFaBeBg8GD8unqTQe5qp370/1jrlumC42FoKdyja
pl+FegXlmo3nj20eGGb60jubzbZok42VKWihLFq6uSUxtrZzmtAYPg42R1FlQYWvXOgQ1FT9mrqh
CHOsy06/+NfW/fBr91NknL2UFL6AdgEr2oze8kbNXYfrgp7EC2JYeY4Mla3k2WSyn9fXpB7A1sgI
1sZFoHqg00rB2lqIC78LvXD5XXZ9O/bNDR0Izf2VxBclIkZHjElutR+kO0g/ig/EdT8sAwCgChNk
Pp4CecGCpmqG439KH16epVkE7M9DPS53ujVwitBXF4FAfzFxbPVVWk/fbqLkV5mv7xxzksY221Pj
NgKEfdNRBLAqKmiymHI1XxKnoYZCneo88FocGKJ6ZtcMcUkpHsLB6bR+UJpi5Bkg1O5e7BOtNGm3
pheZCKSaeEBiIA8Z1RLWCGQTfd2/xGWbu77Q5895vOhMotjJpCi1t59Lx+SnSKC9jj5spXhjAlXJ
PT3/MAG/PUxBHLsIyzAo+RoJ2MCjip5F5FKnkvAaXCNlhv+6tS2fwXzYoEJRH4Q0CC0lpD2t7lB7
8z0+gdeNdpy09FzKBtUI0uYn1n444tM48bOz+STpx5xe6n74r+jA2Gq3WzZ651pYIxz+ra5q86Jo
xv2nnYp2CuziNrF8YBN6JjseaV4g4itUsMqCqHM4nB3Re1P/xwzfYUgC5Wke+mQXNKsoSWXPlgnw
2TM2ZAu4AFDo2eZ4VVilHWKMbiBdXSuGxM8eymeYH6YQpCCLkKkO2MwIO9/Otidj8bybvhUQmajf
7KsBK7U/zY/g54cV0sszis8sEzZ4rQfYJ55Fz6rJnUfpekVXGcganNSK2d1q9TOuxC2dELj5YKVo
P2SrPUZccZeYwdtJnEo1YxGVzqlDrkVnxDkUUEezLvqSrTJ3IoXRtd+2O4a0lOX9+AYSD6w/NlW3
ShRaJ6ZzRqXVzRAsSnJK3P6dXqs5ASD7EGB/gvVReJesVwBdhinDtaRVqaXaPM+J3BATFYYh9jzp
mMKFBHPVvveui3RAOA2RVIJGCZGyJRpbrOjWJftSq4oUw7QsF0pqprRBdf4m6jPPqQz4NIj4oZhj
BuAU5gfZVpbAzNiHUP5SyEUnQBTsEiC+RuF6UISR8jsK6FTuVyYpUTyrOtL1kJkETcjIGAzgXIga
OHvha5hMDA7k541ovpi7U+18AtgySdFmvjjThXTCbVEi179+dLZHatXxxUb3YobjFGebySibFso+
HYzwSCUydJ7P2kgRNlkNl68x08RPgP03Qa6ejKr+NPYHkmcaLyXAf5gqmBF2r+qda4ppiqfpkYPd
hHxdY7G6ARDV8H7MUlhP3NX0UzuEAJrP7sGd4YJK+N2htfCPmWnq5nEZz3AQY3qkCVTLgJNmx4AD
qxNBpy3fEl/pMq7sYji2KE5CamaVaKwBCa2jqQnGXgCnOVcMec93EMP2XKzmbW1YH0q9hyvMTGSj
E+yItLPDp3WLwBL2G4HjHgz8btH8WJYCr+FTqdhrrdeSRFcTtooFkzQoYslcqC1f9q13V/J3BTcH
KHLEfqD+gswHWtw9oxP614tWjbqDHBmeX70SC2RhuOpxvnZTXn0ouk0g1qRpMBNEsYJ4BxNOt3uo
/hXqdV7cMhJJNFxCLp4FC+So8yg5PI1FltkUCbrVb5yKjkVoCoQQk6TzXGJFrgFI0wQCKkHV5Ijs
+nscYbSHaT+mopOzk1Cn+G02bWpm6iychNyequUkXQIg4x7ivgZETCWu6VCM25B3kMh8HCmMAwa7
u15Pl4G8yVYEK3Y6j4akMqhf5fB3p5D5h8JF6MifoYqqAOABbQupuUMEoccFSIPEhbgYmoHbBsuJ
fP8ihkvFt5cFBr0EOI1uffIGpusPNWjThMu6omXlzaJK7nHROvFYs0lCNocefVe4rtweuXd51WHg
uZcutqXxLUWL+fKK590nkEm73wcO4+I6wNYHs4vzbZjSS6aPS1N3SOdSRmwFdHd3qS4nPQRMp33G
WVpyWF4fUdRbq056jNBvaVhv5Tf/a3+8EK2bn6Hr08GFaM1p8bZ2/HzC0j0NHgkeC2a38GeefVdN
zwca8ckxDr7+ur0v7JRL+kbEFE8Wd9dLAsvfOi6FMC6sldmz3HQybH52Bi6bmQP3FJKNwpqEF4o/
9Rd70sIAO/HqvUNfE65v0d65z7/+wyXpXUIbNeS32tV6EyZVdD1vL6POjyH0PJ6y/rFg7gFn/dai
6i/Tn/IPtkDXL1u6WCkbat92Lmu5lxdwWoHOohNSHft0nmWzi3ZTbhW0sihS4+ns9uuaRZ0R+sm9
dIIldTA9hPzj1KuDw5MFOoiVMChaQBDsSpLXkIwom0LgqwfJvbajf3fefJRgTKXENLYo5QksUjH8
mBfZeN3hlYdIWK3B7MJtyFeRYYI35k6R07HXxVWXAuo7+M96B7BC0hkR9OkkC01uPjkdK76Iga21
E9hJoShuAY6LfvnZY1t4zuFMvVWecPUPo3pdrkQQFrjKDfg5lFNUZ7BiBSxS+P4FtoiP++iSiIOd
wMbyzpN2if1BfNEmcALjbD+Q7jxYxHqOeHu7eV29wxIgUpl7dIHAToqQsyD+1pZ5vsbIWPajEdCc
DhgnmiWTjwfmN6hQgrDvlT1qX9MLbbQbpScPp4i6aJe6Et7/L4NFQjKD29DBH+qArJ5Cf/4Ir0Gt
LgY2SoM8cHQ652geSwSNWvIA8P4bbZNvlSO7WfeJ7DhTHCjmD7Gm0It3eYdkN9tfcbdsPbqiFeAj
j/Icp3jc0xZqcI4cDMnWWajeW3dOu/ka7dvQ93Wgqac4O3gc0YiMOfj8dfBaWI+xHYaos++1slRh
IvS24pDUVdCmWsISzCix+j5lKHUkwg2UI2E3r+h5Z4qjsmNIDyudVmCDpKYipFtiLBYiMZ4+ScHX
Rr6qKc61+1CajPAvuDwrgTHvhA74sSpQq6f5kqlWYEeOAPrZ3GIXrOHFyUQostVkGzXsroIZkyKm
tgmxUOcxOTw7M4/JhNPem/SmR21qv7XkOjSPI/O/bNIfJqPg/y2A7HzxU+2xWTQZT0+u8tJrqmqu
XoV+UuckQRzYJwMfkoirJNuTfzXJDF9FtfQNYEn5TQGYfzQqUvIsAp9MRbDSncn7HMWZ41zwCOpc
W/bGwKrSInQx+aw2tanYifH+Cw0alIb2gg74g5oD15h77JpOI+VI5qxJJgMu1cd297xYj5/ziRYD
BdffhmApiJuDVErKy2V8Egy6b5OROik89dX/Fyw1iVuP0F2AFW9Xu/TbNBH6t6mZozKj2cgPhV/t
J6WMB4sO+R4IPGxcpCtK+UNuAySphoIe45q3AL+fEhLQj+ZIRRMuFGsSTCEWXCdcURPGoegH1oN3
dLC791x7aOEmef0GBfC9GBVEh3GtB+nH6QfL1Kj6sPXWqiRduO9dXJD+6euxo26rocKre9nI45zv
KZR97GdL3OofoG2trvDAu8vcZRQBu2QvQ05z2GVutgGby5+wYXKf3xHPpORhKBtDTlK41LCBYsTf
ecy+XdZQAZGF7CnuB5Jwr2z3rEd2Yq0rLL5/k6Ea83X8GwxSs32sEtpyMnOlf5o8Rs+X6FITovyn
M6aoisoNfGaB8sqoB2WO8fgM6tzs/atRVzxFKhPflddzjKrjgDTYlgavEeQBoyokb0H3S0RWnkN3
wIhszKrwZwy8ZEo4rL2xNQzwhOT/Y01hDDEDEG6wYsmrVtdNddvZad7Lbi+Z5H/EKyfDv39qs7ri
tO4xMoyrRfCIbOdEC5SqTim2uLl3FaR7dY1ZAXf1B9umxCVS63oTQOgJtplAhYi8UuPMBBQJuQw6
xGVtUDLaga5hG6nrIdCSJzxzytWjABURieBRO2DE2EqK666MKuL2pbL3z/4mRPI8I4OnAW40gsyx
dg3c+ILenMfby7wcxq/k4rlgi7Jt1klfOm0tV0VaDNcHAmi6BBH9osQ2IniHNFuXKJqDImMqLVHD
BkxfduGibA8DLNbqk0OOYfJH0yG19Hw2Dx/boi6q2N3EvLgLXRQQXJXQKIk6S/aOLrPklGry1kFH
cF6WyZFvlzMopiprjM3figllgsz/ErvBocv45Ajvhsvf7HViOfOIX35LHQsxTTWtgMgXsUiQYbK3
ovyL2iRkAFRNid5pBckqyjLlk7QKAVPSTZdFeTB3/OBEjB+0tt1BT1mX9xBNrdunZk3DN8WXsA3g
c/H3mwnJmm+X3F5wxmPILyo4ykVPJGUgTp2Uj9+FLpVarOYLH1DFPZaAaz8DEhyzg55zDALO9jqZ
Lh8AljbK5R1SUUBJetyYhkjjAhUKtRajjb315v2y/PSECBBCoKbxlGuBjj0IMCOqQk46M/B+yyve
G9/I5hcx6KpmogsSsjKRqyp6J2sdfPEBoKx6SMIbfsjCYzLV2WCCN0xmZNU/vT++/2Bnya/zn6+Z
nzo2mMU94/ejHCXMhecXjKOcx0KsAR2VqvHC1axb2ylXrjKmEDY2/ku9njgq5zGgDSClFp83+F3P
rsbm+Ki+ir0sU08MOo8N06DIvDG9LKyja1pyFsKItviT19ErFbh91pvLPcZ6X0XNxDnmoidMtEWx
4yYiKv0CsjUahJP3eM51Us1J5Khve9zE6a60TqHQbAvrvhoaVCbrvYjiqv/TxhWI7ZNWAkmc/uuc
b3oX3xdD18AFUW3R/7wTxZ6NNpMXIJS6oKiVf9fGG6yZnjkKumYNCwUqBuSUllZBT2vkPsr8qypU
GyEMtCeHHLZBqCiXz9qQhGl5AA/CHrQupqZ0tkBre/BRspVQqu1h2tfI8hLeA/JV6kSxAIxss2r8
BusyQgTF82dtKrheBhJjNTq3D94Eixrj2loIYC3ri0GD6GmD/rnbYEyM8tnuup5WH8HzTKTi3PRo
MU7WjxoSUaMTIaYgeBgM3FZr7/XMWexQtNxuO1s41Zkj2aX+FPESa1obRAusxUIdpmb6ojPAdDIA
+DCd2j+WhU0nBApP+tIUqUJDBsEWyANZCMMTWnTwZwXevgKl6bs+/0JgLKjQh8B1v6yR761X+cmB
WXKJsVRgpp5aTgeA7jG5VRYS8Glaj0qSmDcuS+RbTb/5di3xPxHj35CMiWFGtVffFW5nzhOWXGIc
PhwPLpS1DhW+HwVS8FwIwWq0W2oR5neM22OwYY1wV6DiOdUqOX+vu1B5xy5H+3vAz+ns7UoqMs5+
wnHxdUtaTAEaPzwm0i49kjAcbWzLrswB6s+5Qe6ym+pUmQQSeF3HymSTRacwdJ1x/+h5Vs3s9CTp
YS2L8wQRoCo/ZvzGj3Z3DVDw5TUQdcgUEKzaRtzfX14TaHc+CWO3jWrckx7H1+ylpbJL6WncOGxX
HV3ks8S0ndjaPvDEAjc9JE7WGvEUM/HdEfzmrbiHEj4X1nFUL+w3u8WAhilZGuKBy7mGsbOLDS1n
gvILs9K+6CR0E9VFVhFCmlI4SgxgYvD9mkHvby7hfrm1c6w0NTHPV2VcjVJzqVAqlK1F+dSwbQTn
THYTOpft6j8LGOcJqD3ELiNU0tVFQIphdLjJTJm/LVtApgmStVTtH3ilwmR+Z21foUg1mR/JRdWH
fnqMZFH8uQ6oJt5PZiTIhIIN4/u9V7CfcAxzoQ+nBdn6C0cXLkjh3Ja5bbo9mFqUQKWS1/XDL4pu
OW3+6HPPKE4xat8Xn7pNG2Jo054+QWey/Uvgav+0ddmvB+GwGHidyiSq8TGLSbGuUf0WJxLokiBV
UnPuJ9Auzui65/NFJjR02n97dN/PxxmnSUaNnd2u90V4TGHRnpGhcjdjAwdxdCZae1LLsk2diib8
z1HlGUnoZpnLrSa7UPvA82uiuPj5wz5/sj1nFt93cqBeJ+3NJGaL5JRms3TnOwyKU6t0ummu4NyQ
ep5ZnvzB8y+MhfevUSSq2goir/jF3su37hVsWkmw40EbiakLmMuZeSOiHjTFSH+BaDbLeVdaTXWA
MdQ8ow/pk1+zYh8p3s6YAjwB3yNByzWc/Jh+e58QCC2E93cbZiIrOA5lzu/guQ7gGp/Kfp/SCVeK
AGnun0TTcj+ea1gM15eTaQNmdf0dwCMDVOKQyIz21qP/9CAAi4RTqtyjU/M0t5afhC1yIS/ULMJ2
xmipsfH5lL2OjZPpL5OMrGKAmC2T/kNbUfn5RqCuR5AyzoiOSblZ9iaHB2J0SIrXmq7ltjzv/prh
iXc+GuCw1PLLNUAThiACUtFxEE7LJiruyeNPG2ZVxly8X2pNK+L3yqMW/EcUDzMBqJuzHacIYqEy
D4K3dM9q/XOxv077g/NpubheHbMT4nd27swEzM5GwTdlk2ydIM0HhP63KW7yivL+7QGc5eeVzlB6
SCf7PG5gX7k1vkHIVKwvyfIuHlrJs5jBx2/e2F/znpkm8qV5cKps/OF5DNFNwFyLl/2sB2bd21Vv
SEcecLqIUydIBGYiG/ENY7fuMN/FS9kBfS32ZE9wBtCm8f5Bl0iLn+dpKyCEppruPgCUXKlwR5wg
r4l+gKDXQODgj0eqXbcBwgt27703tLMU+YyUAz7QR/bVK01Mw1V5TjFGDapwtaRbzJUPGtSqMJH1
xjvvXl8bWiM6+frxFqaE5RhnFKiKocHz9HKXe8RxzF+asVTF2PdcaD0AyuTIGqHyYEQ3FYN1es8b
b0ttr4c7nM1rcgh6lyqhacssRfq4rh5FefRTRup4XoxA0DIBnghq2iwqf6LQSLnj7vB6PRdTVkmi
hSNR1hpIigoygV+8obEOTVLyqx7jvwXcA8HRk/5N3cxweBhjSQwp27zxeTiODB+603RSwYuD9FXI
XDD9h0a9EjWrxwFOjtOVGMCYQw8aJlHzXTKO2LsTNwhQI0vijtALmw4IxxokkhMjMVe7oI7qwwWL
9fZsIsHwLjOSeu8moeQLtH0qtjmlUsXF5woAaEX3MZ8+0mjaNs/ZzPnM+J//IsNkzCSCX+wbpTg6
DnuwXEgDnOyZXmM4HQKBUC65RnTt5QjBU7v9kG/0Y+iL3d0Bx8V4WP9HGUG4EUM2WeMDVod0Sa0q
UtXT+nfBftzujREyRxeKinUmRElUYwJNI/Qt0CEXtd/JZVCjyRQ8wPrIUdMSuqMReUsBCAFJGqOi
NumbYn0spN4tBBPZVhHrDTvjmv2RSpJMwPM1C1ndLxMAC9PBNSYC+tOicmai2MAcX+9upQ0l4ZD5
2O5zbypheVNwc/dx2U4Ah4ZT10AD/1gpA2xNrRgBrnDqq2Ggt2IwJw9/PbfsevMbQoyio+Q4vmDP
ZfTswO9XcUrjyWKkxEbialW4a6PNB0+vylj6IRZipS7ZoaaaHeCXyrLwM0S6UeNoTF2w/1j528mv
ufoA0fpHBBHZYznlXMuiroSUPc4iVgiHni1AqH6L/DhnhZMEqEeeLgvUgT+RghW9viEMbncpTy/X
oxlVyNAwsSVlDrN6n25V1Et27onkuL4Es7oRHKB5Oi9QjoV507GjsDLNQOMxK4jBFS2Hgr4/fSRS
YQhfBibHgUCDUXm0Gn4QLUPlsW3INRAqxfH3Qm/tQ81/D3kJA7LPMkNWbJ7jmXKWBe1ikf4pXIhA
TSnHupkc4g88G8yBvQ+fQ5sKECU/sSXKqUnvebZryBYAfdITG6eDGgsuSQG8044YiIREpHAGqZou
a6+/wWFrhHDcX/qC/aNYApCcpICLmKYNnsV0nQjCbdxYefHIlm2j65+x+gWOaUYjOZdHLnifmqyF
yDvWVT1xEHIa4aySrgGu+tYr1cvwKthZRLBXN3ZjvRx1TazVSIHcWbaht7lhWcsWHjX6yb42hK2u
u43kC8viV77yQ3kOze5zijAb65nFh+G8acrGvRbxcU7Y8cq0GN02XNQFzIWXK3BFz7/G61kR5mKT
0bE1TjlRlQL8ETACKNqTf/Umh3QIJNCET5k5en0FK/j591zRMAD3uXMUFkVftkzJYGaFPTLiFifZ
+w6Ilzi399ypBbdtGq/pz4n33LLImD/BDy0fG9Eo2cQZCxyGPCttCUr3uZs3LiVMsfigFPBFVV7y
Dn1h42bHRu1wJ17qByVVuvKU3UmrUplu+m1mRyjgyctVBRpC2e1jI4z0vcKDtrXscK7YkYN4+HR7
LptZ/yeo7Jh8tuj4rPlbybg+dDMZpyydJ1OZypoFefEyvlG1/gxdlMXxQNbXOFyAE9uIKxW2O/Fb
9FZyKPbW7IWFk3brpE0SGVdkCTFUmbNRgdMo+trO0MaYCpQ1HBE7040R7x2K+HCVBJN4Ruy2Cm39
otUiTa/qN6OKqrwZCdZj8euPhqkpsTa8z0DRtzwNF/Ou2walYwUwMbJ1pBM+QvcfpDskU2+bhsCd
DakVdmYs9f8UrMev30kuTN5F513eQ3LGsgsreWHWWYj2hMpdVClyzHGIls45A0GhUP0YKEQfzqhp
B0oVgU8PDV/fM+qaQimLOx75gOke0AAhqNC6qmfz5PYYXBhQHb1Ou5GMWf51jNP1GPLRpaS1MGeY
Vcp91SquaAP/pDcTHQQ5ZngjHqkTPXJSjiwWBaMf6GUczld150TMXiq5gxQepqbQs5UXRf2p3PhB
RQwRVWfCKHHoxdtslu2FSDsF2dOZrk8a7wiIzblUQbyPR7T6vfERKrXykLqAHwJb+yiPXF8ljz8e
POjkFLCvS4OSxxtNH8052LjkQyeLNyYAHHKHGvq/6Wi50WLscFA9BA3MS1PLBXHRpxeu5+a2BGRS
Lu3g5SVER28RqJIgGKNEkl0ttcu8uZk+4CDbfTTwAFNloD3XoTYZXjETWIr7ZtwBl7dhDTkYqc1B
MT5XZaVivPLs05mqNzGXgL4RX/3P/+eLi3bRSHU+SD2USJ5feXa5Fg+wasrn/N3hR6Ci0ojvaLJ6
DB7enmi1/y7EPxom7lbycch7Hh0HwshU7KS5uv3IH6limDMm0azMLhPEPiTs0Y9JDjExcL+fSwt/
9oZKR5w8UHsRPMv/6sj072BXd+RdiiHbDhdmIFzouU6hMNKD2yg5a7KOK0I8Zfn/yfmCABUIY18M
Z6MybfGUIcGNN5I1Tz8CTo1nUdfSVeO5qqs8mQ23Xs9pOkdte1Hqx/adATiAtXk+qAdrwAd1WSmu
vjjirwvFq9D8wQzUO2g348UTgKuyzqVLgUFgJR9SX+6RRx2HTnXF5h9tY/TdSrI6GyWnFpuSd1HV
q+iNaa8xobHGz2me+iHQS2AgGEwfUeKiwDUzonpd3pq3FUcEcqWSPciK9fzWR3DvL97Ea8ITwrnu
utt6eqKKPDa53850HjEQLr5VBMHKRmHv87bje1/s7lLsVFspeVL7RpNkLZA1oKCE0wj9LQODtajt
VxfYJaw2NymAwf+gsIU58S/LZMztIuLp9LB4kWvtQRY44qUsCHC1ZBe/WfhGjT8u4GW7+nt1gjB+
a461ISr8BgQXsibsgLwE8pSniFOfTg5MTh5qvpCGaSyFBKGiKqYD30enQl90rKA9+bgFMEXXnNQh
T/BpKPIndnKvOUyesxilcB5aDNz09Nk8iEcfReZPXb4i7RcQ7L7PyRyapMEEDM1riePP+Rl4uq/v
iNO0jJfg6cWHnjPnUB9HucD8o24iVQ59gIVmqI1Xo1JPodEOqD/KTzFit1CH+ZSJBWBEL1nfSPIY
Qzi6dS8/BxCloYzmlgWmbYn/uN2jYfQYqXWNu47FK0WjWRKbjraMqhK2TX60r/XrO/8nxo36+L34
OvGkiKaBQMeFtbqp1bkVvfKF11coUTbFykqVYTHA05HBVAO4m7koGLCAzXYKHsUeHvOevYsLbo/N
eYQk8bAD/oHSamOiKCOvYUOVr+jDnDDNgD+DSbOeCEKX9VtlgC6IOU6cEbNhdaYBGB0qRy3FEcTw
GJS6izh/caD/hvT/jlwBcP8ga6PStOZpGigUIwLJBchYeaqJQHKDoQj1OAQwjsDuDOo7kNYXfKeu
vPL+UH2+9FTZe6rPsvMc1KwkzNGe7mxVdpR+vPZLtZgkKr7tBec/HEMEwh7WfFyCEKnKPqmHZBQz
OEt0ew65kNs/BFPpKuSSuW3CeVNKRpnahz4nep8TzXcK5ec5a5g8vzUoSnziXjaMZ6ShsxEaPK55
yaXTriRITxBjYdp2N6wZSblsnO7Ly90Bo2g7Vf33WYt87YUKk8On5CApRPNIlGKT0gvdxN4zv5za
UdZIp9YFWXOu9GPKvBgNcx3pZ5lfHkU076jkNlxL9l+IHKMqlhaWKCKQ5agjnCgS1l4EngcvFgP0
odgZ+WTznlvYH87PbPd3IxyuoA0hX90tvWvI37lOYw87W3aXzytO8H1H/sg4B5EvMyhEAjCRPffi
+r0ZfJ7gn1oFy6gmKeLEXkyHJ2F5DyUGNVxAlxoxskSIeWUEHy8UHNIRaaJHaarQx7Nx7SueXWAd
AtbJywWDrVGxaqPOxSAwdEdJsNej4NtvgA2xRzM94dyfGg6Av1vzMh+mzmJ8NTQfB2QfOSREbNKw
aRntz6r1RkvxcKKu2espCRnGkcmujLfuc3R2tcIDZckZ5m0vnES5pbCO0jDAv9ds0nL+EOssZ3hB
DOxjpnt5qc6Z5XN77l7bVbak/6N8rUaTq6I3wFotPt4Xo7EexCwF0m5PXuIoPahOZhjojFu/s9vb
adMcOQpZVZFCFxu080fNlTnDNRLGoWntGfxTUe9I0IaO4kmrPCgQVohGzM7YymIOeuYZDuBl8uV+
nOlPo0XTMp999zW8seIIiND/euVJsmfumM0IhbfZuPHf2X79cyT9ACn/zSlKSPzeZDR96Q3JFFlM
UamfhBvLtgKPAj7iIR1gmP7JGzJod9p/7WUs6IcJZXaJLp+BVcRpOghppmHafgRe1R4uczUVeJes
rZNILGnGH8j+tHUU1GsWspTrDRplbDb4YjdNoJqZUh6XnxlMRIRMm5/ij8H60H68wC5pspmwqcq3
3Fj86FEwhXGFY+BUmmFVvTBnZmPSQ+S8yoggKoIIce7SuDoc6kYRiQf0dD9X5Rsm7qGKHPzkS9Fc
GGGqLDapfzYNPZPmpdIqlzrdxqDqTATSFjbNV2Nagay3QKlejlPa06oyG8UXFjhS2DLe0L1B51rZ
Cxi77f+5R6I4qyJE+77QEvm8J//d00LWQii7fesrl9v9HuxOp2IhEQTwINFcwKAwfOxdtc0E9vaJ
ZtwXhSC3e5X+UpgiGqOSej8glwwjTsvNwkWe8aTZTZ+EkE1vwRlEZKWNhu1alqK2JtQC0kidRxhE
UTlwfztyWe1jTiDR7ZCY/vgk0YQQSUezImj6z5P+tqIuCFGAMuacOnYKSq4JexVtDrR8NX6QZMV5
JlPoxnavIa2ZA8X1X6Mw5lMZi/An6KsfcFFFM26xRRi0UA3fR5YPDK7ozmfyKieKpmAOTuDVhjMo
MvGz9XtWOZMDY9t1A49lGwjKwN1ZRWoMrVTaraUjFXgAeB0tZoBmTdSCvVf3kOIoIbDchet/XIZg
802o8FCxsisaSyK1OP+bbE6qPX6wLDjOVtsTDL+8dKjeKsNIfkTI30PQpFSelTA2acOQEs0HSpBQ
Eps1KwOKEq0FIwPpBTuqhLJ0H3VgWpUNkG/Qdk2I/kPQ2PbxGjxFjuPdvQ98CAI9HNB88VpF/z9t
1z9vdfGvoIcN2UC0ThRi3C+P5aQH5i2hEx/RInzyzFxcHfY5MNofWKQ0Iqer5BeKFDFLf7Cjw+zE
8uZTrt29GKZ7t4kcbnKUUvUZipNUNz5gm7ZXkohmco5r5c4ubTlsWwZkq/ftkvxnSfuAkGp7wOet
RsSVnpBI53qmIQaMKptynNUYXNrEaLvwnHGGXLVJMD+28AbHL6TLRP04YRc8avZpdIgURF5Nz5nH
PwnL2HJNR4A4RiitvLtJUcd7gLbBgSYOdOUp8KYdjbBn6U58ClrXzjUmo2Rr9xH+9eSxunkZLSQW
9bi7qIp/Wlh9GkWmrHLCEzAhR9NaQyUiH3rBPfiezrjoJA1Fn2S+e6XytEK4ErL1mrwIKXWQwKPU
2ZSqFfmz0iYSN3gXFP/vy61V6ojaCFbIR3hnwDGfy5nnTexjZWP4sJMxIRk6ojTc14oDcLY1u3IA
qnR2zps807XT5PjQ1AgFHPcmBDk5GVF7DPqUBSM2qIXQumLOQB6ZcqJ0aBAzQRGPCLOtGesFoOLQ
o0d2fdWFSmZgHPZ8g5a0KU0BIY3hjDPX8LpVaGX7sgkYTPTRj3zK9WjPbm0U3T0KFYk6HG4QpB9b
/vbtw3cX14ViXsGNtlwkETW1n+NEOol/v2qmbgtRC7+BKsRWmHhbQ1SwAHIioOgS9As9pTgLa1b6
nTcrjX1rVlXqeh5vzknAAgKRSApaqlj2+IwDuwdQtOo+v9wfOQQkg24nXfyW1Y3chItGS2foxAhC
rq/eDZU6wAK+t8aJfBTJpWUJQYf/FP2Xepstqot4B6Ro2UON4fDynLy9K6pQoltuDbV8MoK1jcY3
Pl0Ah2h08/5smhyVd/k/0iFo4QSBCRj8UefVwXjWbYUlki4C3ZBCQ/hJJEzFGCud7rss/V1wOo/m
qLbl6HXX3VDruOyG14xWTZ/ashRc5yafBuq0dxSDVWZOSBX2QBhzlvQdJlA1caW169OyPmv4Hol1
da2DJ8ma2tSEbphbdgerHb07Tk/t4UGQLINvNOteYhkrakrp/vlI9r0pMF6prUhiIkw9S32glXAx
vRC9/1ksyRUMujaL7rCuIplIkOmI+bnuBjcfcRX2ZkhmKs9D5kgso5424CmwxfhmVO7Od3Ja3Gbk
dWOQkPE71QoSpkFtmEONOA/uPWeYczLWHxGcbh5icdxHryOpiLUAClILhWn01zWFBToiq7PBrv2p
sTxarklxL51fhiKzB8RWHMMgNmhKTp0NjNt8DUdmk6gsrYf9820PmSRlSBlHoXDI4mxLeIyIe31w
9wIcm2QbIyjLFhpPWiIauy6gmMpqwvCmYjHDtH+lze7xxtAfuD6C4wBPqliLM0KGQSKhjDMBHy99
KW1pB4sZQT1XKq76Wa1S9xx6XDHfUru3QjRXjEDDmcS+qWOsuWGLS1xZvHOpTpii+plB9VqhxQa6
MgmCm06wuJXnyermfribAmzm6thOmm77SjM0EVzSgkW3uOoRTMSlTiC5Kp2kvlFKudbILhYDxuRN
4eKXsansuT00ltITrDJkzMRn8UmOvP6uXLb0lrS2nq4C4xNC5czNNr7RCuwj8wd1QFdxj2xx9rJC
c9agVWLBAWxayKbq3jrFQ5YCn1/7P1pjPpcEZ1itzkJKYCKTj6uFdIQW8pLw1QDztMBKTRWU5oSh
vKr4LJXSRL6vM38I8op6Z0FX20aPh+V7cQpY1RffeNKp8jguERT1wZVkSATXtIaH++4XMu7ao0Uy
KrfJWs/FrZueZ+xta1w4AdFCtR2Z6f/Jf5I5yf64xjVhcFDrnKgmH1CXu1JlLhmFOhmjYcqcKVHA
W3D7l3z4poSHRYXarHDxkl0IYQQpoeWu/wVSoC8VD/ROStC/dflikKHUUHTjmr5pkJBx3N0mVmkp
z1z2CCFHAxmRggjqanzX2ikS6+kCmGLYzUf1KI1SRIN8MqMFXM0TOh0S3FGg7Hht4TM/64oqoTWx
5v6qxcwa0uQdFqTFNoz41TYFsVA/appppuW2KmdtsXlcpialNOxc7y5GDWfj+pDM3SxtNy3zDJC8
9mqifDalXfVllLzpDZF7A8fA9p+jbO7iicLySwBeN03ItaDxU3sVSFWdJ0g0o+K/CH9ZZcDafdm3
s217Gd4N5bMS0EZc16dEbz7ncFsdxCNP7zOh4GQVnx5Mef/5TUcVr2hDXZgfXW+hE6glqdR4SUC3
PbTv7x5wc0IVs+sFDo7mSajmFiegXOI2Ix4WeBh2oDUbLMBV4LB/6f7ppe8VRSHIX4K9EgiZr8NY
6eogOnR7ptxzvoYOBi8L2Z3Uh2SABco48nXJ11mdIYw/o0lNkw9H0Vr+r/HWTWzaq+d/lzyeWsJQ
BOPTrQUsLM/76+bO0RS4XDBiFQymnfxRV01/WaTHtLonN8rJllY8uqrpubKcJdUfdKOf6cBiXHFH
KijIa7ZTqgimLK1eohWHjDSpFb6hZDz8YJH9yfRip/DVc3OaGjMOJA71sFI3frPs4jUXyCdMWt7M
2a0q4Qbcoh6+AH/+6AJO7RJj9vKbvby4mwMZzB64AbeZy5pUozE7NBqAvZ6jxVX+aBO2OTWclNfe
DFkHUqDiiR0blUO2CbzJfqtaTWPdgRtWAbAMyANHtl+qSeAJZHDB5MHR6XqYqcqRFwr0wBtj+eAF
+1RtKPv2rWTXFi+HKBxytJp3Gt5s/HPgEG1PGrK+Glkb+G96ou1vnfNvCQoY1J41s2EKZB1QHFTz
cOsrZAv1/3xIXtBuxXs99sfPYAUq+xX49Ki+l1VavsPIkXMrGSqfDtP0/YxiM5zn9RJX0NXna1db
vqhh2jQE0qUwlQN30VSzbF8b9B7SHNZtfl6fzXlCfk8R26/i5Tj1bd+vXy1qAWFDlNxxEGnnbFhV
HaSLAI9+Um+GnMgtlr8ih39lmVwu13VtZ4bZKlEKEd+nxZZ2Zp73NSTUhuWBRLVu77Qg6SB+gi+j
9fRTKRDx9RcOA6lutHqiRKfS0i+7uMlH2C3w3Zi3muIeDShnvs1OfXFbhxtPnVpgNEgFwFUWf95V
BhsuhJolNvVrKknHhz8VTsoM62CNjOd1hY+QPpJIR2+lblmHTZjqGBex/DLhQGQV5lH2C5TcZ7i1
Exr/TWB+Vxa0dmlyhs6BTbwq+12KAwfvXDrcUi4v1DWx+KJEWp/Ypk3OLSKTSGSrRLOgKxY8I7FE
ychERFvUwYMlKj0h4xGtZ0S6nJ0tutXOvFzJWeyJrmz02iil4xjkhGrQVbr7zdwMmz//5C7dhr6V
wsX+lsrA+PF98MPu1ge4F9crmPFFHEbwdTNMxZGZ6Yl2r60Gxp7O1sRx4Y7/doEeW2cqElWv41CN
1gQARco4EgonZqfRK6tmnf1uXF9v6jk5xxyXI+snElPUyTZbED0xEPZN1shDaNzqcdFr9A6RD1aH
N5CJJeGeYehE9Z48rSiyQdEJbiWre8LruztpnDLHMBwjWI/1znz3yz8t9P1ShD2wsx/ZQUuMLZJ+
mO8WYBKLW+gcdIH9wv2ESIQhm+Dq0AjUxc0olasdV+CdRbXivyeWV0IJtxfu3dpc1JayBxflzvjV
VMHKenZlMOvL7gyCxnmsFaf63Zlr0SdkG8SsuhW5E+yr/vf0WEaeGzAuU1i75MMj/CzWmjUJ2CvD
Rc65MrpxclC3cWU/5qCaSsqnAqN9AnoanB84V4vv+PoGb8oihK2XKogUfrzKtqM1XZZcu4MayVIo
XAKGvbhv3rpfTbPKYtgH0CysIVYLbAs1egl57jd7oq5Ccs43fyvLcic3f6+ilWe/wEyoAD+Vvn8z
9bGoEBA4vqwZVBmpant0OgCA/wRjYaod7HLLNqWaOdq/RS4Q3z0FJLSHYtgSGeQfbP0Uj4n7LcdL
5yOA6JOAXMItvhdGceu5Ayqp1UzAukL8Bp+rRU/8kGonxqrY7G8wzoITX+cj2aBmc86jHUpf4nZi
M3eXqlnzA2Tgx05pcrwSjDOjAPEtQvzQQ/gumjy5q7hMxglK/IMUNUQmklWjloFwD3DYIeWgVPyK
NKRYhKDOMjtGStOIdj4GVHuLIEofiNIIpNDKGTpI/X7FgF1yC5pB8eFHkJF6+3oyhc0KHMa3W1oF
IBQsdW4B4xirsUsdLDPkvfsAJWsLHV+lzeAQ8gIunZV651yX3hwkFiK/k7NJm9BH/zK5O2Bmt7Jt
DHqTWkBiXt4n9UK9PjkQu346ABkGMwW719M9sBOtZn93NBDbREJkvdOb/GdzOl0Tb0eYmEtXVjxN
p1r19BWusYpow67ZXmSgC+KjBjOrTTVVEu2QhpxCtiAU90Klj4B73LJZWYzZkz2QtvZi+2fCQKcv
X6IU68DyGaQlpn+qPRgyhmqcMIkrE97//DlwV8TU/8Xlz3qjH2Wj+RWFFvTHGb7BZfh4Ld6uElX5
XFWZ+AKDzNxufXiOlRzeqLzsnQOog7jeFfJu80GL+wC6yswZsVB92q4qd1Ifb5H7VkZmoX7qPvLJ
Bb0nyu/cgmelNnLJUgSB9eiL5OS+flTFJw4nRt9zfiyw3prAanLK7TpXJErHkaWWwbCDMmregmR2
7vg/SyileFlBNAQJIWiUp2NZpbFtzzzoUSt7hIhetikSYDnq7FErJ2nMImWMJYOicZnQkmjd8FmW
A4YE+TFw2w1ycW6GGN/H/RRX0GvI7VmfxEH+vPky+fOUzC32bQAXgY23Xk0Q0HyJfm7OXEYeLAm4
2wRVI6nm7ZKxyexlkWrplIojMmSmHe8wf7UaP3TZG7nft/ZXMHFUQcogjMidmRt/sM+Y6qATXOmq
kXXu7hIb/Vxyih6b8vhCNRheWjmUjgM8ED722hf1zpUUqoQ72aYBtJGW4lAfEOZJ6JrVl2RFqaOm
evkLVQUenVnBtvAylUrvahXNb0O1w/P67PVCmZmFsSi9UbBKFaed7tniO/4OGe9nZBFlbmy75Xes
2dl3hwiB8EG8s38S69griuDUvIq+iNVq3iao0QI3X1dc/GcuabGv4FQfMMkeAcSq3k6VAD5/Kx7J
yX0BIb7t/sM129G/xwTGgIfT1UlubV6fwbrjICEyzZh5ieXuvLfcGYvi4ArjjAum1cx0ohnkbN4N
kFPi0tYZtX7L5785beYrCy6A46hwZwvhgzALT9Xibo+mryDk1hK4TtLSlhdi1R4YQWUcgpjklNUH
Br9GHcjdE4CyPfOckqoF7MA9TSnS+nTiXatsuXg6kMqAAhWqVReD7lE+rIhYbWeQ6Qg7lXzM7KN1
fty/zPEWvpYw6GsDSENdcZiVe+AxudX+Ze+z7sFformQPMtCLfUqyHrAym/NpT9wGpM8AFzhpPbs
fwJqj3829D1CUIZ87BePJpapFfBbnJ8FZ1GZbS2O61+xF6btAtD6Pj2iwspKxbeYjSqz/+f2APAq
l6CgPRqV1UccBixVEjizw3u0BPWic+VrFndT73B4qnAK7WKGwMZ8vKrgguo96ZJ8844lgT3Wprn1
rXoEflklE6N9qr3W8M+ul9qKwL/+e3dUrXPElOsRKYxYw3Ypz/iurpAEiCCiqnM3A8u7mTVpbivo
o1ojLjuekPUJ876S70fD23jzlWjC14stngmqxVgyrncmHkQ0ZB5dGuaW/jnGEcEo1yjjU3aupk3z
dai9snfYpPhsZFqnOK+JlCpb2PoA78ILLd5rD7Oz02SDkX2p+2rz1OvCltlCLF3IlXJ+W9aLtsxS
c6lPJ0KazPJKpWR21V7D539rZsaXY6STcU+XcVoUwiXh7cJOWq9aSKAzC8iAa638GGfFWyroFNGI
3rYRTMOXgzSsvpRWBszzTtURZngZ23z4gUGyUCO7djya6KQ3BqJqv5xEESzwyGf5pdnrdlkt7X+K
DkN4pPlrYUBd0Y/kmCMFrRc1755hvZzlg9k+r8pd4z9rvQIs8AiShtiamYDJ00Ln2DZxkVRe9uc2
AR1g4J3Rih7PCSwx07xoon/rUHi8gmvDmkClBB9DFbGyEZz8/SXkkOfpUIOvmG6L09DTi+usBp6u
XYWcsu+hyYsuZ3RiCohLKtMxie+W5OBd6CDNORdgLXA8GWcPPeBuWHukoL+AtLRXG0OEJKgxgKAV
DTNccwpBeoGa6b+6+wUo5mXwiw6vi0dQtgXqdie/WW9EbbShDvpTpstZeCte50WCBMqGPkb8RxQG
Q+ZfKJIFbKwuraTB8jnw74f4tEN+Oig1kSFOAonErygHpHfaRU6lqSDDshiunV3T9eVihfbK0a6C
sEpVK+Ju5KBWugJmibZQHCMluG5lebYl/WGBotZ/5UZVP21jg7Z93RiYIN+7Hb/Bja7wW9Cbrkjt
2KwuwQ52/OdeWhSKuhZnacg7n3TrXeEVt/rsvE2rTkyazvPUaBlkEuld0mVtUY2unDZjKFTJENWo
twwzW5CjFJCtDtGigBtsRJ57F72Sf4NjTCxGYzRqqesxyJNmZLNI0o89kmDneZwB6W1bQOdxKR79
pk25wtu9To8QyO3niYPSUcNwHDSEB4cUMhan3IQa8X5WUfPWl46zmBwDAD9O8t+uAqy5ygaEpHNf
1PVcdy2nxC36iFgJK3jsNEYxTpJi9NztfYNYktwJhwwPM2brRPRqrpQ5qGqLakvUVbMPHBE+4qbv
gWLyLhuUkc8VkFkLjIZchn4Pg2YvyR1bEg3kmD2JcVW4y5s0tUaE3bVEluAwz+zMKKgU+4SxurM8
27dWF0EFlpXQCsvm+k9HeUzRk4bGP0kbpodOdov1tIxE5R9EiH0GxbY91YzMW1n2yX/QVCyr6/2X
pqN9yOO6mGYl8K5wIKRUHmiPqzHF0rLqkedLESlDD4s997GPu944yHz846vED31zk7GQPWfiTN/t
EuBiyGeWDFJNam61nCTKC1fm5aVTK3G3ifyEThms6FAcNfcWG44c+Mn+BAV+C5NHRbpo+sTOKbiy
qiG9p1UrwxN7NvNwd5+VmZ4/TNP2QskWNxrSztGjXy9QUU0eVhESL2wXws5mOXEwiNRU/3qeAQWj
pp9wUrBtuiiBsVn6oS+9UwanXB/2gowiRTmSut8p702q/2wM4jR5CIa+/pm9zoFYxsr06WahQbFk
p4i8Qztv6EZNMzC+Up9qhLdiBnRrJ3Engs6JKLJGk1kjcQggmUhmBNJ4Zzhhyocuzsq9wI80wFeJ
kYNhTGKAi++k/9FvCJA/jkZqljAvH9/K8yAF9zGH7AWCiPV+u4oqSCuNbtrPW3R6I0HALB0pTHvv
R/ojNqRArCLK/CaLVZib0EbFgdT3Hf+Me5SVd7OnbW2PSIKGzTN7DwYRdKh9CgJbaZdj5tHjwUIW
LhhHxd9iUyd3TO9TgVkNNnAL+XUbDgT6lBfiGgM1NrRFFHcbLshxQL3Sajl2VhIz/6aMmKjm+lx7
3meMBKWqpZjzyYU+Ep64gbvGz5Y/xTmk28hZsfr9BTV+gPEIww6tTxE3RtHiq45qKLZhWeYP6Hgg
O3aHRJ1xTxQQoRewIV6NkuRJdptAQeihGVpf1KGpYrmRGwmY+wHRKNKA5SB11aXTFoLFeJjXy8kx
jOH/1W7Ets9Z4tG2IrUyy7UmW67R5XeR3HU3fYlWNmOIw/shULPmrwLqp4gbQiEFyKybcOcx37t6
RpW4XBakhL5hSqhWh7PWfmXHCQkfosIc67lsWtrEDRRTTfqyZ/C6f6CWOQGCenSfRDsnZmREEJ3/
LiEysMWnpAe4ZUmtzuowl+vkARjQJ6NKVvRehHwUq4yVn80/fWvvaOKTSkBCnFhmPPfxE4uM6nec
enC3fail9u/Oqb4oZ5RqSzhwcqaMnDsu33662nxjHWwlvo01cZ5eCdVhkLqXU66MBHPeRxa9TDYJ
EyBUqss24/XNOe5JfUQll83WvUYxr0gaMlfHJK6KUalTHT1VHm1B6Jukaoapq9qtj9wnJK9gqG9S
sVprkCnIZZXQffXJstOAZ3D0nYJV1lpL88fGbgSyF6QuSzks0eVfvbNZ2bC394R2Ugw1STpP1vAs
DPAHscd9Tt/pPn5ASVV/6r46//eBZzv1fdOnBPpp7wJizU4Khy/J27iTJ04N4h6Ct2q78yovNyks
AE1URqp0kc4tmma8JbX59jGMtgQOvn57PifMPe8XbaLzKfWGq+tU14E9r92X066a77FV5IP+FgOi
ssg/ZG9fnvxle9BQXpM4JuF/UBrtDabLMys6FsUkPZEPmr8LCrH3whBbSniee9ijnGgLBkbqjMyH
daEXllUq4ndHPWa1xwXsYpqlv8mVv2mM/tA7vIG7pcbz/270Blukx2/Os7b6bNpWOuqi9fCuDz2z
gjAeWdElYyNJCfuSPVbS10xneBokWHZ0M0lF6tHgHXaojAUASryudC+TKwWmy8T1+OTCW6285Eqb
X/j+T5z6DMBKNcG0mrh3pUszZCOqAJff4kVKYm8lcCd71lIDHCBzZvwKI9yQk75v4Rjm0//frBgH
4LiVVogNqpd6dTnC9qaAFvPunlvSC0Ww7TJkF4pu61YPwguM7871LVydzWhW3EJgoAOnDIahCZO3
wmAtHE949mFtZWx8FK+j5adA7FUdmw4o3CKFQi/WixHzROVzcPjZt1dRDkSubgvUm9Jbm0AB+wWf
+nINcrv7FgAWaz07QfeFJDe4Aw4sRKVkZtpfV5N4Bm3nQ+8WK7kgsoIAJP5DXK6TI0OjYki5CMkL
Z1fJjZqP443BSE25dXY0iiE7CrNurlPnVmtwBw1dDRKOOXUpYUSgbnW7sp4Nc0cPykpETd36A4V7
fAbgYx7FAWSw4XS6qzrvPKXle9F3p7ndKdp61UJRrWmzkNoIBQyH+bW418zUBnIDFSY1fhn5pPM7
KNKNd028MununW+8mx7/qy42Lj/AffifReOvtE1lhjn6Asj4Zmjy+se8hY+DgCyeZ/nTjMcweRFs
GP1J4DN+RlgcEigPNnOhYZj8uW1WzjjJpLQo81bPTPyKDCqyiDbSs409mUbluABjuYsOKe0DBlel
3Ng+iyXUNopdCbr+/lQLWqDr/Lt4Rle3MDRMVW9mu7EjCuryxMu3cU3Q5EwENgoxr8HKdyy0opJ9
9Uuhe91kWi6ojpd2wkxZ6fCvQs4QGwXAqc8IYrfAKdLJ8Yc3eKaCQOjPPPSONInBIkZyF++Ayr7H
4qsfDfmGeK2c2aEOvmHb1kwXqWrpkR2RHT8IxCAhK6rx6pvpkOvGfrQJxrECLC9sHDG0GmDMHlZ7
Oe2eMo2CxNT8X4dQgaHOzG9ogwoo8aqyvFy8/FMhBYOp/PjOOtGrmpaLWx7fdSIi6F6Sr9vdIMxY
Vpcwa8AAwil20bMX0wGXo4gjDE68t9Spvu9PHbIakGTw2c9J/4sxrDKw78/KPw4lQaYv+sITCbtW
SIg5thFTgsQrtUJLHtEItCQMrLkTxQtRykGNThWrKltfyBeQ3RMknUzE/+TP3bLwmLQmxXPHvLoZ
WUt+UAGsFRJsFedDhDyfINW3nD32+sxCYSxEHhDuQm0qlv2XN+nczIRu0HkXElsySjkQf2L8s8bQ
pRG4aaXGN0iC88/6rIiweHhVgLBdb7agyygz4qTE9qwUOH4I4bEMyhuamUaouTh4+RWhuxsQvp83
+fHTXGuozKbNzrJ+Wo03lH8sYF6bnobaTBrewCpdfi2PWP83imeGw1FVVZ7tCljXKEQMq+q/Kyh/
GsHwyQo8xKbijZoDG+XFFinhuprqqKYno40zuiQTWlo736m1JQM1w+QC9F3uWFT4ei1AzXyqc67w
NK3krBqvOAl4Mi0sB5LWpeFAys6bMuKep1I3FHoTl4Mlb5j4JevTkD64xrRyi5T0PBXIOsOcF4iy
abj8lkzhWyS9Xcidqei+lJXwiqHU9zrEaUjfe+QfSrw68n5Y7APnc1mAyy7Ff/BNDW7OgrvTKkiH
AHT1kPqfrKUtSrwqhhz5Paem4OXFI0tVTorX6F4stD+hk+yLbefMpDaqqC7F8BTtQ000qogaHSY3
8aJ++40F0DkXnPy+u+t1fkIvWMiHEMNOxZZPDRa8Ckcg4P9WCkU0/csIlK+thyaDc4N1qI9wRwmS
vnoo1bDH2qhsmKMN0Krc1Yhkldosvs0xBVm1XB6hO1T0T6ismZUS3A/wgspIL4E9BM32PY+I4PTG
nsUXs2qlzhaYyXr/XW+BhgHGKHu70Gwg13JEPf4087d3ntOcEiO829H1YkOU5FOQ4U3hD8pRgycz
wi8xxJT4Qx9VYtP0q8WLRRDzM3g3CXDYDPobuIK/5IiID9u445uO71o/zyVm6mNSsA5Pt++GAvA7
YHaxyFWO9A4ax6NKcg/bR2hYxl/Y3NavsD6Oi87pknhRwz+0Gd+eUUmWkzZbyesascS4E6wr0zgt
7/ByH5aYUQtpRd9tYuu/WCjnE1nGrnM9BluLtHU3oImXpGwSyrHRaWzSCnDnVCE294n+527+rJNB
lBI5MlUCXADPSwis+v/xXkG/9z+dsL6hW7728yO00FkgoXZC7oBDfT6O5AUAGqWV2iRyE8BJLntJ
GdaCyKD64QAcZH91mloU18H/wR36GO8lt8Jae57nY1arjT8mhsgk3BQ1hVrDd/Kpa4mW4QT1Ycxt
9xw1Yq56eoXir4E8I46ebjDw4urxly6GSw0QP3zBIeBJWDK/EKeDIGqKNV30Jx2YKFNUVGavbtav
ZCUV0TW/fx3a5xMZ/AEwngUTMaRzd+XG1FtIkMfdXS9WdRMTBsbqKDyj4GU1IoPGI6BJwuPvvndu
0Hm2AH+adApjCoBWn/zLpZECYykDlAI/oX8n9H6+ISs09PydLBCVWkMrGg9ZQ5x4EigJlcO9dFA1
VX0mk80q/G9zZVfaTYe94p1SljK86l1aAjqHIFwJWWWC/HkgnbU3wBXrkqzVsdycewNPyYkIKUKJ
tuUmcGWQxeuMsoWhfVOOzTFQfRT88mQKdReN6rD2Riv3uukXHQmJW3z3WOA0MyKs3VLzwVNt50Mu
A1pTjFGO0T+Yhym/22/nI1T4hVbAnI0ha1yvn2APZ997tt9LXO2obLiSpviwfAC/3na0Mmp9ku/Q
ld58q9+NAT/Vnx7yCNqsRg4Dccmxzf0QC+02QzGeNtH6KfSYe3/3LZCg49ZwMQE9n9z3a4MIHqd+
Mb0htjRCZZJHwyseNmD1YM2AUUs3/OhsJ6EyhfFdiZz7OnYobRrMsXLSIV6SzFDL+nEGc5gGnoRv
6dA+CBMmhjvkfQM1cAZ3bNDf92nN3ViBZjxbtZURs3WQkkNpYTW81OkCKzT8WHKQTHUsn5pLvwDO
Q7CYiCJvjNI6e9Nzo+Av1cZ5L1x7MrDYTJuMBh1OnCA2dP1mLEUIfboK4xGFO0Iq2QrM4oBBOKBe
MmUhrWz8Nhj2qRLvX3ho00xW6pPsTXnYb/RwLiGvbF1ZoD/dgGqiedTXjnIGpFq0wm5ImcF5yiai
18znqhtraJmeVGFbOW2FBIk2Esfmjr/y04qes/nbzPqkI9sU5cQGTCiotTRC71QUOvxFMarK793J
DP1Z0np2Ty0Dk+bfv6N+qPPHRS0oSkD5anfAELFc3OrSs+6mhEWaqCa9hsHVgTz4x/qEUtrQXG7N
Wxz9uG80CPUvvKrQjzuLZWfQVS1dllFheg8ZIUztVowEEAMU6GUOMm2zcRrbbi7N/K1w2JPUrBAu
xY4IA4ppcbgj2GhGVX6F6PTo16rF4eAr9OqSsXJWwwXAMuczQFo1/fSbKLV2TDmZhsT057s96Y4q
G6/xzYAyzej66kn4qNwbYOglZz1ACWsJ0hSt7TiORHNwb/iuFLS984dVHGAb9wsO2Crh25tuAdyQ
Uh6qrJN0WY2hBl9fqfOBeXmaqQjOeQeXYC+SVCoLXOaiw8faNdRVI3Biy1tx3u0hj7eNHD6DCCcF
3gZYcTQ9Wmhp80kClT/InYccqH8LIaCU/Fg+q7XR5K4lJ89speNTmZbx7ndzRZRxS2Cij5TstTS5
lzceZgf9G7jACOmRFLmbbZlf7QyOI9JuWQyPrC1UW0veiE2ypJR85QiXFYzPjqwvqXsxZm5Tch/M
SdQyw6/48XdqNH48w60uJaJ5urSxnYS4RpeMEZGSMSFVOXp6ogrUjcmrctMVSAwj2d+Zi9FaZksF
WZBQJ+XbaNDsYqK46m98UK3tFkJuaWjFjyuX7KP12k12cFBqjlQLrqoJBUs9wyAvY/y2l2aEqlML
GigflvGIsGbp3cwz4i/fs/GEHVJvYvHE4jhGHj47LYaSMn9A0AZ4up01chgncsxkDs/eZsQ8atip
h7sxFsNxt5ZhBg/2q72JtrcvEtIs7QujWI/PtQZJ3XwkXzGD/I45L+LnrOAfxQhmvSLKDFyNrZCu
Of4x88imMs7dEa2/ScZyEGKyWc9EI7zzCks1aje93/MvPVzPDKMD6Xem/gCwlD5pSgAtbgSruIOf
TyWh4LCgkpeXRNo3bF3i/xDFwDNhTZWhdNttZtBXmSwuSX+ESf9lJlEJSH+XAuBDjyIITIg/hz8T
3ppFWfdvaMZ/C/HePZVfX7oJ89hur95qccZQXOO+YESzTC/8oGKKogwhPuxujrijkLXMMKeiL5rf
3PCK0g5sxzAraiF4cw5iGzsZL/P61KFTC4CIUvAzjkPjMBZPJLaFp++Qe7jLvblyR9vzZXkEi8Xq
/TctXQDSYrGk9p3CuB6ux+UUdh3JwXqgPUcPh0/bn7pEKGzHQHgg16eiDg2QYuf4oImBRuB+9BCd
3bVfBOrAE5ot1TvxmCr2xpeHzNK5FW2Pep7cojz0HwdBTByFUrXZnsoxBcitb+27BA4J6YkLZeEG
0g8o79idulDQV5hBTGm6MkfBgE2tlV4RA/z14opzRSK/FB5hkJ6kf/Jew2jqJTO/HQ2boaJj4hx8
Zd0zPKQQQlcpXifBEed7VZ8Ju/SJNany+Z4bt8iRok2PSxXQR8z12HqYjGuEeoRBLr8k9ggHY6D/
TOAgZyEPENJot3axM+J2SBfpJD3othbBv8rjrWI/Mgur1clFd7ymbI4quABENj6JhTpvhBUGGbxP
lI3IlkZm9DnYsSN5O4jdiCWijSg2vNMan9mMxmRKy9ZM1pm6vOyQRqLYDGVZwWzrSEbROMPtJdtY
c+uuVV/TpwLU0Vyb3mK+I5fC4bIW8x8Ncrg9YiN5xmtvDqaBJSlXyphmONTMPk0Vnqhh8HTqbz93
DucpaoVH+rUgG+LUGHIxqI/LkFdD0SrrQg59/nOZjHwihn9Dh2V0I0savuavK4Cs9a+KsAaJf2Ta
USFVuPnFm60c3WMgcq3TTN7NvPMGIvszcdh8EqC/OVYsJd6up91WoQGKnXcAMNJACd+oTXhMPMyi
NA9qBbzsxbuW9q0pQQboGJejd8m2H7HL81/y2J2wI8n79AhXWTpdTjnh9+tcripwEVhM9/a++GbT
iaVqJ94FKC/7jE6mbkY3C6Ey99c50E/wQzBY7jVERR+xAY5M+jq/74G5yoe5ca6La9zsW22oGSXD
Mw2HnSxZIZiFVkB5zcMGgDs1eLMa508xgU4+URXgQRAN5NvZVgTO2Rl/940EvigFr3HiECYzSTsX
q/qScengY9a88ZszjQUyo6664Iojf3woV0O6jkcVoju6x8+eqV8bfDOHQh/cR2isKlZoJ+fyLUAb
VyZmkBWgOQqCeGqRUXwHTv38xj9porLFiA44NhOxsJTMRBrN6AFbeylpkCz7DW81TH0t2u4geG32
A+OpprEV5N7p3v5Gp7LKC8FT/hCsG/iVpYkKEUadS130Ej08SlnnD879bEwuiAwIJKX+eVXRVMKK
FE622ltjcOGnEJIwIjbvF+NOrcWbo5Cdr45ET1NgIHWtfU1conugKkgv+MzcHta0tgsLXqJ9iPbR
kJlIyS64l7joDgsiHJNaPmWpPc4JyaRGjVdw0HfdZoZUIQFuJSjrB1ZAXqLsAA6qy6T7V29JSGXv
4lbasnqT/vnQCtco/Hz9NkcaDuifQZCrUkTT67oG0O+scVwBiihtxHvFAEOWzwygMIhnTnPw7TiD
eW8wFnxwOEQOJmYcl/K+e74cvpd+kxypvEo/P+W97U2YHyLmYaji2sBcVP4nZvoBDrxvK1nFoLho
GLmMNQGFO9KqIZtPvZQOvQyhqnLgpjlUKpnGHqbuQkkq2vigqI3tYtD9VSIesLbwcsu09BIjnUbj
tELNR8Ktul+tdRkRnPQYskdRTU23Qld+MoLdSPBYuKE6wLPG8glTM7ilAScQpd8A2y1KZkSVAGVz
SN7iHa9d5WjmwkLlQo8r2lDXIr43j91PQF4/ex/tLIrQawaK4GC/VgJFTaJgkgv52pP3/yUc7tIy
6N6MJ6pGQU57w4FAgi41ozL5rTo2gob/LBBihCb7kqBc0XO+go9ufNHoBFR1ehrhQIpYmbc9O1la
V6pPHuaB+iTIaOQ+uXfm3iIlW80KPj6xpXRarj9hI9kQmyAAl3e6RyEoaXwz+0zKASUb8O8UBG/V
OoEgY2xq6PphfEm9fyDOj0eGugBKACl+tw6kcoCo/7iOadjkPfC6hTH8gRK4MwB8S6UM7hEl80xp
1MTDdmGR0Ct94M0JYVRLKz5SHcw0AzHIVy4EtSHh/fzM2Krjp+eMaBanvClc3xjoIxJigZgkwiad
FWJiTIv9C/vycHXf57Z22kp4GgTptNcpjOWO8uzkg+1j19hPO8ACbSAA13Vk5e7VxC9RFYhFhtJn
ytKHKXiEoZX9lDrVmN4wNDZo6+ZnjQ4z/2Q9SP2PZ/MC88fkhKGL6iX0Ul4giLHpuh14VzpdtvsH
vBhUJQL8AnfEqHO5m/JQzsfW9oP9SNRe+H+5BqBJRVu19NguzM654Wq1DrbbvEInn3PV9azIHWym
2SObYHrOo2lPixEX8VUIJEK92pJizPW68B/cKtYn0Iag/2m6SIg9kgkrZYfqxtNwwWQMGw5VlDIU
qvry92HcMWrKv44Rsbw4TefN1u36SL9Rl+btq6gmmQDnLs2I0ptPXEzUOxWSfqH0HrjU0ImHNEu9
ns+cdD1TBP4MEsR15Nj51jUAcux11MTDTDTqtIwPHWYgVSJo1KhGQzoOOLuzUG/ja8cgluaAHAho
RxUgs/opHT1xHuiY31wSSY7Qqcosv2etn2Ow1/JaTX4zZVFQBYFHmlXU9cktrkK0Xk7W6tNtNonp
neuI1M/hGpu5Dzgi6E1+Hx01C+Mn2rjIQT+0qyZKSr8YQ99tO+5ZMZoi6PRL7PACb0tmRta94jEG
XJ2IkOzhs0W45Ld1zt6+Q2mbY6meuDxnst8zKQsr3F9tVzBU8gBf7LFMI4plTxKw/7WrA+PvVsdt
M345mh6MbqLTZwkOBoM9tRp8/5Y0n1VAd73ebnZ4J44dF3q44Ql2eEzXYj5arXRvtxihFT4xAEY7
RDc8178dyyu7VH36Y70dyGBG9SNgP28aPjThc+0lBXzTEI062O5Z+9RKtMSgBMTXVhEV46J2jNWf
tRvVLs35x4oGMXTY702Lo0tupq9Dx65LXdGe03MVfnjr3V8Co3B8ahz/OaFgiTNQ4aedcgjgU57u
0lkeY+gYwtsE65ASrE2HiyR/31GCg5Yhgy+vql/QRJTJQ4isd98aUsDVL6XPXNlIug9aJtoyRZhE
J41QobGPgwaDsClylwGrqU3DCfz6fxxGe8QOycUERGsPwxK39LlHcBLax89mFGgLj49db7ZhWMcE
HA7Fy3GFHV3sXKKHAfaz5007aba/xHbHWW1LPdhEW2FgYNOpDcqnyMPNAQwpFFLkODCJpP2LPBwq
oVoeuuebHr/LbTgGa2rc49cjDS/YKiM0WT4taS+oi+KT49vSMAwF6EvABRp8Hyar7W1xMIdUtgdN
yuCGWv60QtisxaXIbn+s0U866xgkV27B4ZqqBQTnvwFTFogB/MXRCXSrh1GmvFhPE60aRIY8ULgM
JwAJnDNyfa3G5dX52RJLpB3Dr9zJbJn/Ox+6TBzmJzoAOyDf4b4/QtMtxzerfGvEmXuMyffI7zw6
2uE3r+zCvRDJ7RcbxzVOi21yHNMTO+lilI/I4Z1waU6Jci/LLCBWz3jHhg+hT5W4QvD+b9UKKo39
x5xJxAJHOK21pv9Ao+/w4opQ0NmdBYBRep65bieQkYwfLuBJP+oG1UupWOUAsMK5QlKvHmr4OJyf
bFKqLQ7yob8hyh+FgyjBq8B4V+m9FAC6O9NAimiHFY2JuVwBB48ctruek2CftP/9rSgJ/qYXFl7e
kfVRsd+Z3lLE2Rrc6T6uzyRtbepfMJgDYYYWfNt16DtWZELVG8zf9nofUiNL2b+lYi3/D+qgQnDX
1NtPfR50qQIHcxqndl1ENgPgbYfyQdnaTurXSPLzLcCZcdSJn4Zq+OSzeTrZuyhc5wO/7BfhpP3x
QDpNbS4JCk2JFd/FKH4sqMr0rn8Rgkw3Qp9UwF0TxxHpD05Bu5HNjVUWKRaJnhtvVVko5bZEkgBg
WKwyIz5t5/6PPvhG1mSGtEX0Mpm/UOeiV3BA5i6BcK1tZKRMJu98mvm9Qj7jr2eF+gw0WqwBaHLy
XrOt9OKy29md/nAGoWSV/hZwtRNO1HyYYG7CWQlb38L70vslCWEIF9XiuAJVJ3TafKQx+6fGXUUQ
wNX549EtnpUkT7fOsj5C6F5p7SmwKEGXyVj1/ls7heGOJZ4tQfDBudeiCJHdeQMTYJWF3Iei4YjI
8oHDH1/gh+EUBwpZ9V+PmCtJMdr7Q6UFltXgmHNiOu5yaDnsZxOXLNK7T4eC9M7Hg7Mh0iid7pfS
poehCF1P2aHSt82r6dzU+sSASi7CyjFOkH9w4uGq9TR5dq/C9JK86CJfBErrftuo9qbUG+/BXKd9
+sUofL5eqygb5E0hjYlzZZduttnGhGbsGxJbEo03BHy4IeP0ffevWreTkHkaQDqJ4QDsmRm9YFwp
R4hH6Dwl7zztI8ZNDmUj9EyOQor12tCulcy8MVXF9W7wDc/h7pbBS6RARccZioDNF+4EGLa2hSdW
K04LGw+WwvUAnS2j+OPNzlgsAkN5PbYkT0OCZydfICaebUNUQoYN4L14CtWjwtUlI1yFUhaQ4vYh
kPgr87nrkh5VS456e7GMg8O1wIKItitib5hxWotxXI6UQZdbzq6VP5FR7H1UyseSVIo3lOkg0rbd
bNreYzTexXONuScV2AlyfxlKJ8GXEm+rzV/xI7Cqek0MidRYW5WqTermwAA91CJjPe32P9oixl4y
pSlssljEX4VU+bLvSIuasK9wZ5cDmr9VVv2PAOAF5ow6DQ0vcbbMDEs4RbBk1NaCaot1pevfHQ8N
n9cUzs96UbVxKH6jPpYEKq5E1ShTi9KDBF2n9/lf0Ob8ayiw57Uajw/tliXunuNeX61eUfLWNcHr
3AS1jvLIDz0qjEOlZk2mKLI5788wKczgczcidwuX3aMVf+1ApnRIk/87a14PqQXllcZhl0DqYk7g
SOzqIE1PfzV3BUuw/RSotcNgVq9jlGjf544WlwMD6bAnrA89pvY2hDcE4E62SM2GBcMgU72yY7pA
fqaonP/dHjehNogHJfLtZG5Di6GXt8WwWAGIULBRiPzCG45q12YFyXfudXqFshMC0u+umXEKdoMa
tCDGKUB+3cmey6y1oDRKqgBCkqAgQF5izsO7euo9Q4Ax74P3/FgIIA4KscyUwAVD3nN+PT5GjDan
zT9j9oN67nyxgEE4k0DReMq5JGY/SY3tzbuMQM4In+Ev5Djkk+HAgx12xKUYtx6aNkzZJ+bWzDL4
v1BAUbinDCQNTRHS5RV5hxjktLt3Z1wT8kO03YIxDXfcbJlGR720QqmXNLbpeQzW0KHx2qcrDimp
bzzaXa+iuhcVk3prn13jhb49aqmvkv8GeR/EOJvWIi0wZitvhIq8F4lfy+O/7TDbk+1HZPNXWrB5
ziIydesFDa/SLGnSk2JO85EAr2wi3rMKTeMcgGLUsXD5jLfk0PdpcpMzUtnKMnt1txRw74fjGC09
2fRMn2bEHsF23yb1deby6ukfXB0125+e8G1aNAng10Bs+dFmR46wGBJy2wyxlgk5Eb5JvZQW95NM
Q4wLcC65Hf0j6WdvBM/ti4hXDiCo4WG3lEE4KZYGFqSGHNGb7H9jcBiXfpQQQCXgUG2ZFqIPD2ru
ci9OcgzJkKGN+xScXLqQnuBnjlvc9t/C/tOOMs8PifPAnD1Re9Z0LidzsHWUbzyJ+BjaFoWMJfGm
qQhflTrAqlzk6s/VQG4rHz5MBYXdIlwcQXr/5Bf35c/AFZ6xkHMVVdLqSZe2JaspepAuiGpqGMHZ
4GQSRDQP9sydld1K6IbUpe+4TryyFGCuGTj8XyAaEDwqNL+msNznBLwd2B8Tq9sH+Nnt3rYgsWy4
/B184irbTYq5rXpcwKLdQ19sCTp2RpGnQogt/IZDgXPQz95FiU6oDpKy2UD4szHBY3mi1lDWg/kQ
DkhV/3/PojVFchiQIh5CXT3FM/JtuwibofSoeZADjTOeGTvDj+s3k8KpRQIJNYCn5R6+YB/OaYof
nHNR951qbkvkf2QDVuJgHLOqabopSAIq1sMQfA7hyyTBgbqasV+stTOrYGwIWEi9228a2PTR3BCV
yqHyFPKFKhjTGQeOBMv1OkCV9gGXF17yjokAxJ1qVh/XHjxsnHS99lvci3C4TpBeVvCgqQSDcUIU
/IVSv1UoO754Wmva1PaR5yQ6Esw4cflCvcPGQT98PZnZdRqrAxojOs+I4zEAla63zrcFE374a0L7
wMeztu1dIEJEBPrHeLrrC+YGwHdu3AVnac+J3JDSjl041Z21+LEHKBY+wIC/BS1lhMCdBOGvoB8e
6tuiAEUabRlcR/4oc59aMOZOS7xdj0dNV9CpPT8lmNYRDrCL5xexNHDboitLOsgMFr0SU3Oe/IDH
ivQJEc0G8Or12RbjgLJ+VYV3WvyvPYbxpngfy4vf4qXusCAhWhGt8rW7Hk/ummUpi/IvL9AFNDBw
G3HqmKMDb+m8h89CW/XHqcn2CFArawjbuHoJ7tlzwZhJyictOBf2rIWr9ORpr4PBLsZT7Pycgg5y
a/uXxCHzWxz4CCzzTfqE6Ig0Sis5cBJsh19xOxJbUHrSju7Dw9HPHHWbe6t88fLICA9z81cPGEvI
UG4sZ1dGYatSKe624ZZion/zdTLXEF5bs9rjMR3e+doCcNq1bigZx4yhqATlng7XHGCl6YAI577z
sMVv9t/hxX70TS/sMVFsDQXrWjiiluT+b29hDbBFZ0PDGmGlz8a6BazhdYZ65Cf3dH08No2zoJY7
juo9NdyCK4WmVQDNRf4powe+gB0klNmtML68bTENW4WGQXc8W3UfR6gAQni+i5MmPqQGcmSCgQgi
eP+WReyHJPgpoxNl47DeGnkbsqMYjwdqMv+f+NMq77SBQO93KOQGRjjkDfkgozSaXUboW/jMHgG0
05RWC5auKOZIG/ma+9lFKvfsa58ko10ZDWq3aApQq/qvquViZiuB2nSIedeRIP33n58E8i2ewqUj
WDMluWyxIpFQhv8veS9+LYyhLrqh/B6eUQ5yDVeeYWQKD5o80FouDH2JRKTuvU2lWth0Nd6LvAI+
kZ4I4MwQx/VJFoMmibcheQtw7gTFx2Vivg3QqEUH+UNaF6uXPWNGRDka0Vj+H7i+aOA5KzTR3F2Y
O/o0+XwHTLbk2E3jyYcZOchsyUCOMXqCr+HkYPv5HvS3u4vVCHufuQMYtdsOohqRya/z7Zk79wAS
yI2GOn/pDNvQYt5oXbwrPpUOMlHTE6glQCzrE1SNCeg+yCo58Z1J8KUZB0Mp83DsKXUmtIdlpI1l
SnLuhqwX+5hrNYNxisjoRiYZXRAx+f2X7lMpqT0NWcESHYAnSA/vLZ474hG5tm+mTzzaFlfAV2Qq
VqCj9CsTkZtOa5R32bMeYMat0HjwhapauPcRW3zTy+iZway211taqopDtf98x0DO9fJMMZBrP8k1
NVpbRGvNIxL55RHVHs3BMPfdeNCO0281kxSSKsylEz0+gkmEHaDyNvOQvX6xo2Me6XegS1l64fg7
tREs3IBJh5FMpLhugfvP0D19FEiigBGJqwKkE7yaj3QDmO1ciTK6TRyEL5X3PiS567by7JYI9GtS
PHDd2Gu7ISVWgjHGfi0kna6N40b0kpy+56n9arAyc3DbUuf9vnBjqLESfRXhoOrhxfZnUHr4SNGk
o+20BxaUjqAiGWaAUDnQ7CS63ASMsFIgcVwNa5xxhbrmd45OTJMXpV+TI8If9uKcVKh5gNFx411u
fIvOU8o+IngFqFXVZIL4QrH0JMQTsnz8p4rr8krGEWCoY4GBG6UUUKTHDCKuUGNHYjDLJm0zMuU/
qrmMLLXE0b14fiqNpUYZBN0K18J3nRz5qsur8+n4NZmzZ1lsXmfmumU332hwFoRKrY5HuIQ1VYeo
ruAWlwoKN4376PPJbVxCdjOcGWDqca3qP+C9Nn41AIzF3Z1OuFhVjV4tpmV8ZD3OmRdqydwQWYzY
Ry9L+ie29Q6MSIVXMMDHK4oMjFwiJJrfBroFp5u3+nIzFCLFrZygdQee7C6aZHzEzBz1jGOALcbH
pEYeVj+boTZCqKaib79AmXlRC3OLLiPCgVd1dgmfNbLsFbjV2q2lASnWjLXS1FPHdis0UnmgLPmt
mB2UQCitiNRlr4mwugvpST0+/YpsCm9xoxaVRIwntJkXcW0CY7sTqp9tIZPUFXL4sfzobRwTV1ue
AX+cWoQ35QPUlpmdos6d+4c5sIvj51VLWTZYW5kVe57bvP5uQHaoeVgTzTtm2UlUnQkwI0S3DVi2
Blx0gYIEYcG4k/iOretKzue64UTiNJRfjms3XYx4S9B2nJF99H+vpogQzZRyYXJzkLv9oq9ch3h8
yCZxfp8NaUawRXwGAEa2iU5an5Ib2IsHigcE3mAj2xuty1N66Aqznkrqz57qdY7AwocF1l9y73VQ
YXSYSEwejVgDjkjrKd2aNo5XAzf3bBGJmIaU9JOsvJcxPaQcV2ajafw/lQzn5HdhVQg+8c/P1hGU
+OPDrq028oE1N/+a1LgtFyG0zfceRZ+KNuptg3cA1dCi5XrXTbpV1GWREzTGR3XeCLkGLJjU6SKr
RU4Qt2p1Tbut5/4xiijM97GPxtnmVaqtSXAiUYkrA+bUeJAiReWnINrbMlj72BS51V5PNy3lenT4
YpJn2IzkDtPYY6mleEnr6Z4dSvs6Fj3JZaYgZ4O2tMzb2rd+04Z54V9t4UbVmAbkIIA3DsCqEsOB
2EyVXWOmRi31rdOyZfd7QC3JpOXgoot9gN6SkjnR0AIsULs2cUuigg+tN9sXv8KGsxYRL3KSWAH/
aCG24GhQi24JFpd0KBHL+HoQgLKWPyRKyzvRqOeO1xSqVsAqraCt5SoRQkHHKbwCYHp9fXD2nQhu
DsPMkICMzK3j+7ig7zLr1R4/x2f1yheh2jpRbFD1txRMUNEeVtsvvnkCGnMtVMtNYpuPS6Zmd67G
RRlDT1DcwiM0QeQRRURgFWmz2wBCPf3vMlS5jC53lSKcyJduAy+lFGbQvwjC19HoYUMxyVpU2Vv8
m3QXaPp+oncNGFWHa16Sl7pdpEn2bT1ICjYwkiC664Vt9CNHa2XEvmXXZLobryQa1J/a6E91pGT7
RSgPN62iWk3oW+m2Bog7cVEdPD/h8/+zqal0QxGAfvjUwEe2Mvx0/zUdiJlITGG5YLYukmt9bbzr
Rnn3blkC7yrZQuV2VEfG6ghcvVOsZSKIEhcFgrzcSEfGH/DbfjmTUY/VON1cac1peBqbNJuU62O9
b0mgbokPDC5UcbuhupEMk9bSxeJLUcnfgab1KsRf/JSkfnGk9m4xKjgpJzJ6VwiptceqKTEOLFs9
1tDtlGlIPHNc7j6RjSS2oAwRrUDDsAAOxB7q0YVfxMTL4pkS1Jbjh7T7k5K9n3whExxrWRofW6Ej
Rvy+cwE3t9T2I3DfYnfOo3i3mMyKP/n/FBKAMB+RCUGIzF3IQynM4GwgjIhNns+kANLzKDN/Qwyq
G5J8npR281ZGwdhaA3uUxcqPkPvqgAqFb/vh8J4PyHhntyDj3c5D4QieF+KUvQK7x6D7khHmphv2
cm6HQlgndza0KXJaNN/ROymnBuRdpbf4l5bhOeshGjQFcySM7TO4tNxnkFNAsq9vKJNuK5xNDWhr
U4b9nQDFZrrdplJAxDsZLsMwoIimy6ZCz9J+Yl0QCUQRJzBr3SUuuTMpAbV0aD5EfdMgE0W5ASrZ
hPhvLNuT+ZZIkJio+QwndrwfGJBh68kp4JIF70whwo1PclCdjY9XKBp4vQb0wx9luWIa9KxhtxsE
KsSoRShVGeszdyLUYgWSGbyCbNNAi0Ta5kq923TkltzNGXnxJb3YLrIBXY+eBzUXdjgKZr2SY9eX
iE7r+UDOOeUrq5GokHCsUX48YAd78d6/DdcqpHjLpFGwEFLaYh/a2ysf94IcKyWJCif5D4zwxR5d
Jtr4JvCX6J7LcJYPsnB+n/iGQgMa8q2OtCcqpVwas8vj4ty7G8qxqysI5NLF8uFhUuaX1Dz8AWuK
ugZkhwzbZp5fRnIMA6SuEpDQmFH9mII2nt1cziG7dskfG9FSz7DYxGsp3He/920QhNcW1QzZdMKy
fwAcgu+F1qn5Ac2uL91ejz9mP/Wt/LomehENDhXlZPkzaHtdtsH3y+Ac6uk/RQumCqRvEAE7NmQP
HZ0p+tzpVeAnHx3jiESKRffoN5vK68d3MRkF6KeylY1q1AaMElB9OUybDqIgfHzKlyEsXUohSbE0
M+PG/yAjhRGRUqQIkIeCmO2r6+OO8zWjknZOnVetEn6k2FzqYzW6WUJrshZKDpVYDe8GiMScGnVa
wOCqWHYpcWhEPsztHZ9Q6cAjyqbA11Ep83O+KrIgjJi+jBCncSeJuZ+bjZ41ot7Ua+MfgKlaNRsf
8XNrND7HiaN3PuQkeSsvhAlRNyAm0FeRROt1rmwkHtCNxV7TwxzZaEX1Bm185K7oaXHt4iJ7hFVw
MvNyDaO+1cWIfTA4aCIJmB4FbbWI1pV0oGACSCIueZwhATzHlas6XyBbfTSwDVxXFzXCivq0/FSv
jwf44XB3z/yAaFzKomwHTK0LfgX78N1H71YnlE9na+5rFjyC6O/47UQ7/DOOO/Wc1ZOOXlAb/us/
pKAWnfOIFGOfAHEPMTGWbU5+xrtx4uyhjIVOL3UX1ndRX1HZT/mrJflM+NtzzCAzEf/2yUf5UGAw
gKt+qF5xvBBLxx1WoijTao0gonD//NYtegJrQ5CSPp1+nJj1w1051XHUM39dafzKP4AukjNGtQ0+
RO5M/prO2axirtW+YGAFr2mkrJAvuIT63qBshifjyKwsh3Y/fQph70fOAekFWoEEaYR07E/hVR2s
V+VRh8RTuWbhnG3IFh7UsY3x3lw/nggJa+ka7cT+iWxl4N3NzkiMKHMoEcXmPNpvdkC5eQgSZvbQ
g/NfKD079IgnXHmCV1y8ilfWbnSHgrg0He3Gp/5Fw3UbQEJfU2qknGOWowV1S8eXqbQGdn1NHTME
Rq6u+O35r5Wc7k5TGkAykXCJDNWxCUxFqHCvym0qJHqedilVIO0sVrrgzHEYY/q6IdniRgnS99bz
a3GVFAQlvKarBJqvD/XYG0ZMklU+SL8FWqXdkDup+4QOUAVyPd8xHKg9MOy7QJI/KYxusM6azkgD
QmI9grW4L29D+ViRpGd9HHbr1LV8q+eAgpE4lgiXVU/6GokwH3+ZbobdvR93fS0MWPFd0JqcYDL7
+TjOIrt99DPdHjkexRBVewXavXDrxJSn5Rm0ekoR/WEWftVrqRV9SWRrEcq+PLjtyfxM6XE7majp
vVBZYtyczC3pOT8PEahicAn8xhzuEllGc7U6O31HZCdJD/e1hQa2rgn9tSSjGzPlWHnlISmnu9x0
GcWlIZHNk1t1xp2KMMAqPDpfGhY/N0wpVEJzCZ+PuEEObh6KeSuLjkqj//Fdl2zF4X00PsH3d5LP
DF5gfJilZD9QIgR0BKNvBw1oHufYyhKkZWPUaGxJDOBp7qa+jxbAPPDua/VHCalln3jQk4YcU8mp
uNHktD31V7izTWiWpbW7Nog7p8iL+CnjlpreTKClj86jmIHCPEjnvNf7vaTxpUpp3z3bMBVqB/aY
EOa3F6Imgk24917+KqTGERAVfhz9NNoV2eKzFVFd6Yjrvp4+WEStq+NLUei4oIPidIxRXlipcgib
8a2AZ7WyXApwG5nHfeo4CO4tbp3iijRGSXmIpma1hKafTig2j4GI3rxPGw6ZCKjxz0dSHA/6aWqB
30OCr4yWpjzmZ64xJqygrHTYYbtDV0cuzyv9vPuP33D4n632ifpw6noNSdUWfEBG3s8GemxOvM12
hkibvJ3s75hSohwJ7aUMNvq55cw1WMV1De1eCqofhM2FIPh4eoMzKMcG6RdJrCdZuPoGPS/lQMQd
MWveUqP4x473i/GZv1nB9AipiR6bJY8Q+nBP+RS1Vg6/z0JnPDWio9H76b2YYSa3Y2RMhsqaQFhX
ZJytcPhA+suu1bZi7fCWThxa3OtMuxXBArJsJV2QG9sDnPo+HJYEDFQNFatxrw6Ra8VecOX2Ol94
3Q39t+sJz5O6/FOrTYj3tI1xSftU9mZ+xMuXVs7wKy+YsembuY691zg9NS3d0r95tfLK3I3lLmPz
SnslrhSrtW6vp4+Y1Rn1aKzUwvHrIO82pYIUnrICO8Ep/prafiWgBiyvVjoO0A8xGKw0OMZQdLhq
H5/anp5xb7OmKJeonldB6zpkxAyEOvMAeyHA6mWPk2xpVK8HN8R31WWEtyrRdHNBIKJMZra28nh1
7ghvsbTNNpY106XGvlpDl9d51Z23uilE4XR84ucU0Mw5MIam0WIJbXPx4EkkNRyvC21b+xRtG9Ry
7D4yvk+XL0IrxvcyiT+CftVjP/aaJcfbzwOoYV51CK4D/cT6kJkEPrtyZG+vnQWvXPqYPT9SowTe
vBaAFNfyvaNEkXumJiXrMMess/z5nzIZsGEyh8zqBmaSmRTerv3aXEBOyGkOBkSIlYobaDg5sIor
lGmCsKwXF1rLPpsO/933nJS6JGcCGInKfObVGo64wORJJnBbQQiL0z+I535RppwvkEXezgjMuxPL
LRDxwN4n1iktsPEtrjTZb+amKW2JantdRvO0bNO+plQIPXIsnqnkeieznNVzMWmJgHyCMl95/ZBk
NK3gowxlMMswO8bcRVhu+N1ZHRqIrg+bV7n6adJMFqBn3PuLSgbh8iLV9xMl80MD9oJLy6jMX5QF
s7C80NOeFmiDJJnRHJByStpsCthX+W3CwC3EsqVave2ijdq/bE3VhtTIIJYOdm7Bc7HmipGEaOA5
5Rs1TuXpo0QKn/KEQuf9lDYQyMPVTX6uNUeVacWNgEnPjAsyQLuqSRP/KBRPF6XgVk3Sx3NriXrO
wzT3Z63b9sVLhyATIWd2DPqspcT/VTzOjO4u3DwdIYdoq0UxaksUfWVRFnAipsD+qAh42d4HEk9a
4q2hwTNKFR1iLHW4Ex49YWRaYbWpjFdQbTp8ekZxvmaNkv/GRqetBxKFeu7Bui8f2YRLDx0Hcrzf
viWO5PAF9kNiscDK3npR3YvcgDaP+ERifHqELmiJ0GoUfRHpocyN2ioiCwMuv499oU7R75oTgoec
60J3bDGDEvWsCRRUH1ZaojsU465CTIal/Y28eGVCL2Q6KdAGxDOG3wGyR2e9DDPsG9SqsBeVRk3p
oqqnt57sIN0trpAQQClUEhVhDuv8xm0HbhMH6W3gqZYWLjYT0Vis6jrlNZPBq/mSnYY2BkBkbBtq
OHZaCmfmNwJxYqK9jVnXkujzv72FVqUVsGoJpM+RXg9CcH3QDWWUYA4ZQOubM96klzFZlFBPrCau
JBOImo8iidkxrsSSuDSRNT353InL3dqp7B0CKW6dh7hohqiZiGc6zEKiYDe4LwOBMj/CHlb9/b7P
v1KZFC8Wl0bZnc14KYkA16a3j0ntQTHOU5S02+cmlOZxZb8MhNhAUZWs6APOWpeG5vJ9sTluMVKV
8lIuM1ZHnUBlzLm1WxHF0F9LF0RT4xEivt911MvhStji7RPAVACrfMxGwk6Tniy1DdnsRGe4VdkY
0rRe93wju/19zv7oS43qqONpCUAtUGMmJUsc9ja23/y8T84Efz4/VhIuxzem8B2U7hS5yIbd6a0n
meWSTnJN4N7ZK7yngwTDD9X0mhbxMdj3JLQJKKKSq1zKRRqzWHhMXxx8sQ6kjE9vkMLPNOM5RFLU
D0yl250aLRruGqPr7BxeqDXt8mC/QLsWCqkkjhDeVVC9WQH2Bv1GlFvQYPNIb5FF4sbHSujCu5Ik
VcxITYIH3CV2a02zGw7wQ7vZAD084vJfqsdoPV91ucUKspCzayLwmimiTyEAd4894MIRpjINg0Ja
Su2O6YSEuRxiY4jEZ1JBTQWG8m3RZGXz3z8wlcIvKIlNh6SRmYSbaWZR+lKwU0vlLxgcdOjYr4Ov
srgaOMan4cdghbKpiNj02nqWDn8kYm848zyOeZzmd2loNGf6oA==

`protect end_protected

